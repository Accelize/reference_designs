// the following constant contains the activation code value.
`define C_DRM_ACTIVATION_CODE 128'h079BF34102F9A846E56FA97F63D41568
