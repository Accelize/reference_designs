------------------------------------------------------------------------
----
---- This file has been generated the 2021/11/22 - 15:46:18.
---- This file can be used with xilinx tools.
---- This file is intended to target xilinx FPGAs.
---- DRM HDK VERSION 7.0.0.0.
---- DRM VERSION 7.0.0.
----
------------------------------------------------------------------------

`protect begin_protected
`protect version=1
`protect encrypt_agent="Synplify encryptP1735.pl"
`protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinx_2016_05", key_method="rsa"
`protect key_block
IHSBEaQtVt4FSbSgqeAWnbIPQqxVwsftKqOP1AXl6XR/2oH9NlrK84ylipQcJtf/VR9e7P1wUZmS
F+sZMhkbEfWVqkBp+30cfo7Q0Go1IHvebBNKelQj1S2wcNM7j9FhGYAU1ee48iZjOTbepdxw7r+5
3GKMD1IoCueFBbRp13WbHlm2O45bVJ37tEV00JgyyUFRzDocDGpvW7pH3C3u5e3RS4tM/owuHNqz
DMfUJRciZ3eto40QANYUjr1v1Xz8Azszq5h2xbaBaIMsDa6QciIKpovCm6WpGyaleHZmVkFPTwwH
LYr4KBD+i8fJwrZmKDpUdzgQ8Wec4kUhl4szFA==

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinxt_2017_05", key_method="rsa"
`protect key_block
ZojMyBwyjW9K1UbPRHunalcXYMlCwZOxR/uak3DfdnnTV+JyJyG+Q/nd+JRkRZSCb8vUakrY/zTa
q1F6TF5v3+1bjwMLvBtTKvK2gcnQtzc2Lop0JqD1EWACLC6hSs8qdAthPHzMX48LXN/JI+W40C7c
WqaQ3mAbhNHtsMerMkvfZ1wXYSLfgUX1a2kC3bTv37n5pTZKpSL2JK8qk2FeYQej3aOHhjt7jIyg
3AAeXZh8enDBbI0ivGhE5TPi0TIZqXgQ6yyJhJl2H6MO8lvGxS78Rt2t2R3XwKmfCTMlBKfQubNq
zgOpF5pyYNKOMIs+MTjqNTy2XEwtV4VqpKBO/A==

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinxt_2019_02", key_method="rsa"
`protect key_block
ZrvI1aGDqt8PzGGsPh5T1g5506bxb6qvAdFcCrTHSb32St1/RGVefqql08eQb4IHJ+2A6Xkf+1XU
GG+KiXLiRJ9Gyso0fvevM2bxysZqTV53SoBwjDuHy4corbgsnOfpgy0cJ1lf3oWeuwIEVc+J5a9Q
3hYhNXNsFYp2RojeUG6lmoITeLPAT2dB1Tgv+2skwjHHPhUDr3fCADOP/wZ+0asOjTwOXHT4wvxk
yazufWWlm1V0c74ZSfVHEmbaBdIqFQVgKn1esTz0VWmfQ9QbGEugCqApcvHdqcQqp6isvZ6VlsJZ
N0O6N+fM2ESXsRpdt6VwRcfUsSp7h2DeaM8GVQ==

`protect encoding=(enctype="base64", line_length=76, bytes=873280)
`protect data_method="aes128-cbc"
`protect data_block
hE34nKGWCnFfwu+fARoZSopG9FHx1YWtD68ye+7u3B76EhFMZXxFBU4YKqCuI5BdeupVbriATCiH
CrvLeGHWmPr9yJXevD1PCfpHCrNzTB7pT9iPz84gaO6+j31i1i+7r3r0aSqR2qdkoe8fHuEHbvB6
G+ncbpUsouasVJffgcgAULCpzAiXTen/WLT+D0gB7cpTiXhjrGzbfqg59bGyeqAdcLzMJD76r6HK
QLlirvp246/8fSs3LZ6OvuXwZzy7yu/upRXgoqZNmMY0vvVFi14+9RhnWwQkkCDsop9OeuiOcOIH
cmW3RV8n8e6TOvFco+Oi1gO3josV3hkqC1JfgCPXc+ls4Dsggfeq7qWHc8LJfHsKVKnZmEaOD2rJ
XtsipC260XFlfxTzcdYfk7dzDzWqEvMaMZn+iycMJi1G/LiAe1y/t77cfNY/S3R4jhiehSVlmIw+
4gPa3v4E2B1y5Rjs4YQGIz8yjWDes5lsIXPVpRne07k+FPTKu21eDeCwbzHo+RFx3d5pG8mde4hl
E6myRQ/5vPY8H79VtUrcIktVmu0CoOmm/cbd7ywLXdp0fewiuar0V9NQOw8L9S4TiwdNDfk/Czzq
2lRhlqPiqbL3p2DwoyVL3+pWYqDT2NfSlhSEDNXXsh0OnFm6xg+vvPLq0Ur8smdfyYDg+i1JoXVi
742o0xGbvpDqK9bL+MPdboscr01cEf9YfCiDupAej27wfuzNjeNfi/d3tLamX230vEkOlAMaCUjx
Kxgl37SYuGHXSM3gJgnHK9Y8J1B8V/S5aCZeDGRKcoer/Qe0fycAwlh5iHqKDX4W3bOgfS7F9Kk6
GpTJhq1zoBTTX0L8YFHyEbAN+fWThrmqLlyCeZHTYwSrcZj+0hns8QA0ARrlXNUIABEa5+B7CdI0
j2/ZuP2vJ2+U1YuVpY0LweYByLwg4/ohGjpmK4ma0cDs5cny/siFrrYlcDVLZ+QqVr+LwPFfTpjp
9kc17BBWPt7GZgGJd/BeHW9YeXMec9YcVEb8yvt5wZEcWBY0SLStuw3eRtEtsnGwtwikL7GlF8ua
uOljRcuCobwHcucbLtZNXxUbkFSwL1fGw8Psmc0nD5yg5MeSTwYG2mpH+WJKGuyGqrohZnPAOoeU
uEYO6qoAeR0n5GFqd/ElirRxNa8qT88kWtBHp7xJQ0bf/dQO4kEiBniSoKI6ugXuZBSELcQG21dx
YwdIbTJ74xORYiVMzQyu1w7kncBppDN02tHG3HilVL81fUSoTU0OLqsWNe474ALTwLHU5keG/Mvo
t7RT+TuxsLcfrGCRPblHgonRa1XJWtJauf5gzZyHz+LcYliDh1lQU61iOkCqw0+wouKfM0T4i9e8
FQBPGwgEzkZu+jAIVTJqUvNeBzwVi4oWIOEy7a5xI02ewWT5sxqf+AIRSrhaGfb8DFY+MVRlSxq/
vF+YsN1F7wki9ibTMLEORQSmz55weqW6hmOF1fp6or3Q8vc45C8GEIjIhV2eJdsyVB2vwAhbJaWb
coRoLue5oq6GGFCHt/aqutNw6ZkKQ4oZeBydcemtP2hW3gbOvdbMRdsohav/6dBEIbiytc4jdS+N
9sthR1zsC7RLscSDQt7wb4qrAHVqQfZ3pTKixUcVARwTrtZmCDhcTZ1k8Ixcph6tf8/TPRSyiT/J
QsgzYtOejDr7QkBKyl4ATLa3sIVfgJsAISGoUNc44K7Nf8xsiWF+KQX1TxF1H5WfkBmHQic4Kk8H
xmPmdsZhg7P+Dv0EH45QQDpACApnWAn5qoEkCUzui33vmpqvL9l5m++rKg8oc5jyJjt6KBsdinVE
H3Ir1o52q2dqz0wP/PDc72wD55Hkg0YKBTj5ns/0Km/9crsm9K4UKQYNiJRX2H6BvZJ32uCSZPFL
M3vRfUEqhE6Tal0QUkeHWzOdvTBDsQYW1Yi1QCE0gqzeUC+uEE5yirrIA3nr6Q8LVwwlbSyNwCW0
kFZ4XxQWHWQIc3nQO2Ge/2N2MfCYUMW+PoJHiKM1BqsTd3McHhK/qtqmLy5aMJBulrcrXpfSADP9
rydubxqxt/c5TtMj4vFb3AOW7azDylc9lH/h7ONFyB80aDitqDwugCYOppw16lW+jZbuJTJRCfBP
tBm8v6jDy7iZcOXAwZnwg6dzLe3FTZExEGIYd0/urpecJGwng1zT+h6Y91FMgS5y1XUrBKS/U+/d
eoZHN/N+kO5Mtgsko2aToG6TIagBK175DrRePFOQuusPBRMXgZ+KumLtrLg6saRFwXEexHvAkAaL
qK4messYr//zAW6C/3JFXewg+CXSJoCbI1SGMb30clw7fXCck+P3fub35wNPXt7n4ekgVaQd/iKx
UYIHCMf7H4jqiOxOzXSGNNKo+7Dx0yD5o1K0QF4ckVZegkvgODiVR6pk+a0fPC4c2wTLpaW9Fspy
UlQr+0qbw1OdJNoF36QwjJQp1mf5iXP3qn0UW1mDnM6+ijy1aW8O7oWJcDEYPDLF7GZ/9jVQqPm/
zZ4RcgANVMSi8bqfoNd3CSp/UGp6qgVncq8f2AzRBJ5SRCiRXXA5Uja82Ge9PrwZyM6ha3pn06wk
jeeB8zlN43EXDW1AKyVqPm5c+rEdQURKZLSCcQJ2kLUirCUJppM+nRBjZTJXOxJ/EVg7c84WHjLO
7C3VU9Dj39RNqbY1Hn2X68Z3tCkAXZXCtNcG96V6XGDldNSFsaf3oDv8WVGotuFh/4EFlj9IObcT
wxdAH7vPzMV3f+KIAB7z7ZqYMAs8DMrQP3fSgUh1d1INeCDC6RoJjj1Gaca6K/8ndhM/UFlr6mrD
aEsIC+0zB7O6b5eLIdTWSVZXOvSqlAYvjP9OYwEQ4eZiplrQYdCaYuuJpCF3G7L24K3vWnTX0ilO
d32+BdMr7q/9Ane/NqVAwuh8mlu+UjNXHkumlfy8m20L7eNwww2418pV47Cs7gd9yR/acdquzvn7
TQSLbBKyQJe6x5vJNoK79W4rvpI8pXhWrSbrCE8L2cZ30DcvM6obXdWVwl14pRIXSE1I0me7t1F/
uAnmg4S1tuVxdBJ/eymDC/HDqdfMul+VZ7nk7x/kCJ4SEFmbAZ9h7RUuJCysr9IRSTjJa/NQR0R2
HFGvIkcHK68DkDCitTKMykDxIa52evlF0huPTl/08j0PUvQ9aPpIet/C/mArFYurPl6E5zodR4C3
6hhKNh7o70OZ1euKa5WX3luY8IGV0uj0ZqJCznt47yfAnDjrDvCnnzAcZNMPiXko3oSHfLJtn0Pw
iPh4ui/T+QDhBNM/EcqwTem72zy/kS9WwZBRkh6XsTTp4hOtOvQKfmgAlEavexDFZZw3+MIS6yO6
bg7TwdnfNUWFvrwj/SVy7UwZfJcc6XtGFCPBjHbSH083n0CA2o5OniYXuWZ/dEKT9fOr43yuD/QT
uSObOayWtRPvIBxovAPR1xnc18ZE9IvoCUWfrA1meQ33GjNbBhQ6FPRd7wu2KWa+J4LNBvrCU4uX
EeHbxgd84/zDzbOuZtrqhq5eqt5oSH2vdD/uld1ZSY4QWDw3Dkj1dVb7ccfQI3ehw/iU4qQQB++7
WZgaWumJUPMMZ059lzyXry5JggwRXim4cSgOZ8Dz0xR+C9nhY+GWzus+EB5NMFQDf3OnDXue0r7o
pzGnL5FYvX6Od+8Z7tjgZheEHJdMdMo0X1mkJGTrlHZQp2BHjRd6o4ZzMXdN8RFY4TLsAm6Dq4uN
HgWt6683J4fWG+H2SSId3RA4ibX73oUC+blgC2+WUyq4ev7iVFfAQAB8ked6vkqk60OT/eHqxvuA
UFb89kg3r5K48Km0p8r6vxp1fEUjSPL+BugKWJcrKUle66MkNpNqtkWVhd7EB6Dmog8atIXNid2s
Nflc9e0CPexoDM343GzXhYtaIAmWq9uSfxOzAsjJUlGVtStcM2AvvGE7l+OD/lTV5L92ji+x5zCE
/V350SYNNNLnvUrOM/Mc70aAVpYbQo49Is17gjIOeYEg9TK3vB+Iek1HfxAnBkWQXhthmAP+UgSi
3nPXGbTQbhZtQ1HNv+3OHy6mnS4aCF1EesQRqTfLbgDeBlS9wQ0YMQFyC0dqes7Kq5jVAIjvCEji
ICljq1JGVpvo26RDjpK1/uhggoIcgs0rwc3FIEQDnEJkktZC/XobGWWutgmyAUaAPh5e4lzCcVuM
gh2Kax9kG9qe4jnM/Z80Kt+9i7gLih0eDvLyZt/JSf9P2HJ/xC35z0+Z2RdlCJxsow/csBTRTFqh
B3xQa/xCUGsjfj4krf9eBs+9jabJE1iHOH/TupDFtu0awvPmDgPq6v2wyB68AKDCGTJ1pfdO4Zih
ZtcR3ZPdCgKXvXkP6GTChvjHc2V0j+Cpk4C449D7q/9kbJbS3M4YbXGQ3e/co84aGZZ/HZhtm45c
buLh8BIdcA+7ZsMe0wqhd01VH1gK/+dQbH7yEJqaksfs8cgEd45IQRGLIzv+Yd0SjS1KplEt5SaQ
eMb+JNinU6Mhsw9CDCYnA3/V9NKvNUUJTtKH1J/+7GqB33Xk1/7Iczw0Pxbm+w2lPcrHxrc/qoZi
61GdQjRH4/ITlnDp+bcZ0v2HQCLZeRbkgrhfUb2ZSBFb3WYK1+FLfrLSdQs4DLC3DCi6V2s0bWHA
3ysk1uNfoQ4CRCSWtkLml51GdsZUqRR8Pn0k0q2+7xHjd2VkDbXsG543KZ1WYFTu5DnOcCVkVNnN
TkZ0pN/RID61+S58rnT4Q1M5rsZIHETIB+I7In8/Q+/l8Q6ohzk/BEaKRsXBVc1BNd0qTgubinnp
tg4II/kdREUr6SrJxU7PaUPumQGm8v7GiG0yJqKWRMb0edoaCLOCTpn4lCTqiG77xyBZeT0hYxxk
FXnaAoR1GY0ZgEIB/MzplYUsFPBt7CFsgl5ZzPtEwPqHjtyr191NVK8tWV3Vh0vI0tmRfImDxLBW
ev8dB+kaVSxgtwZIZWRWedHiIPWr0oteF+mQBuQpSNLx1IrT8HlEYwgCVg6Zc9INKM4RcXeZPWuI
jkT/DNxXjeYLDTYgSOsfrt7J562hn7ero48B4xBexU5xtE2/KdPj34mKmZ20wXl0zKsaPgkdsG/I
YVwd+We1TUOcs4ipiCp+LJUyEgYuODGMxmlbG3rhdeX19iKkHD+vUOGjp8mD64rjUEdqn0u9Hdbp
0KDH/PGK9PBFtHklvZ5OoWQHWNtXbTpAvsM2jHfOGm6JOdtRzHespXS3OC1GsZn5+CQBNsUsnVmj
v9IEBuyRCshVabQTmA9ONfux36HddYSRarKOON3/Rog9zJwM5RKB2RHBZJF00U1xtEbvqexJJImI
FOY8ocfZC+g0Y0wvGL8PKjoZJEl0wgWEwDTmV+RGQZ0pZKnVzkTcgQyVNLDg5Nu43Gzt/KHEks/s
v2QsiHO3iJecr+m7jUiXbzaW2xnEQkquK9umRfKlem14cJI2JwrS3AVl9wO+1L94x1EwcfY03Iv4
JHtB0mCP3z7R6C2eo+aKkCPMmoTK6an9r4tnke+7jSISYX5N84LLEslYsNIsAUVsnL6EPZckZSeD
VbaIQHGtVbnXAWJlbg5q2fUpqJlAgqdbBI4oUIUiwWSuQazdUlSLZSROLxR2fuCZjkYZBeDQjd54
AzB5ZM9YbrDlS5scq0wOMow8x11jiO8mBLc8yHkOfZJgvwKYt9WZYW8mrpp5t4TwpTtIF97hgP2A
7FnGBE8KR5y3qscN4cMAjA+iaxAKqoG6Q67CNyB4kLyMdf8NBqMSZgv2DxH3MMXbeeEtn7cgDzEh
ecOhOj0Hr0WG+RKCRfhOIvEA8VR+GeYmf75ETNCOaDJEczP2SrzZkdNagk45vTvMjaSPxvDIYsvv
u68WXiOuhKWcnlCd6SPsGOUmIKfREsNwTX3lB6PcP2nI/kWR/BbOjYhzOpLWnAfVKcZWo3c4CLGV
nr3g5cnQ+M/I5ans7s1fvarCNQCvXwjMmHXcL4XZo8uzWkhFvWVKCgSpi4y27e/1H0+UDccpnuND
ImUgrGq9/YZwptOtsFAB3SrsEsIxGWSEt4cqv+M178K/2PN4iYitROfVTSXvOBmDhVkA8pbjo6cx
+jrrddmFv8X9910O6J0Vj79JYPMi04fQ25GcA3lgipRCtQ/bmiDvg45/v+Yfi1aa7zfeOAtkaOst
Q/qC262/KwmpyRkeYaUbIHfemswU2W3vnypuOn7loixRoAHa8wles2uygboqPHcJSMBg4Ov31QdT
famCmj4YWV/BCVeX+u3EnuU4ogAXKkxWXQoVQ9PyGEkVHDCoJpdQs6a00pZIFiThzRvLWtnIzTGl
5SpcxGeWmbPuK9yWBvgzWqukaP7aPYCWzimW5GfDuo2Yy4S1AsmrAngNDMIIRykijzDwu/nXKPRI
0o+UtI+zvoEHhQtByL0yozkZ6fX6cp/iff5QS4AMTjKkHx4qHym5FxV6P7KqgegEHsyrT6RfD4e4
9odROhMuFiskCIk5HGiiMQ4ZfNP4qZ+DHEpvbeWiVHTTdtbcE4tLE9R7pyQOlg1bAy5c1ZMZoMSR
VEJrYufmptA6RYxToCG+uP1BmhooC8Sz4JsTpL6kXvXCVjzRL2Y1OTi9VbOlaFDp1lg59TDcc8K4
/YRUGywEQYurJmwzNNZd+MxE4XJks+flwA2SomVMDsj6xfJ8wc0zGYQo5vmb3xalmL4kcNmoBMun
D/lj3pLplrK0pKWqCCXTIKpNX0wvLCHUsug3ffAPs4JzPkcwACC07Yf/jw1u7UhBCZ+BcmzI9lKg
6mBBfnQ2dmbZStPoABL+lfeBLr/CPjbCXg8NeVMu5RpUEx8I79r0C9GPZhQ6lpXJXOj9XgmtDk8Y
g1D/7lFYX4zqxjUcpbJVViH3YJyJxaJ9zYISlqFQpfVZeFgbUujcF7L7WYX7FUHmkjqyvRApkjgX
K+PQZ3HACoY+AteftD541ysH64bZMB8EaRKr6V6QELo4fu0nh9+WbynUYchkSWYQhF+9yCift72z
XU+hGkwctGGVhzEtBKeAa2b6M3DO/8Pb2H4foaXHvdH/R8ElRTlCZAySuj2e306yZNQ7pSmlhfZq
Lk8G8bCiMtnun8IUG1b+ky0IWr2NgRcbPRKhcvmpvuB+vsFySQTSRCn5xyBx7q1X2ZZb85D6R+Bb
gqhqiNltOy6iqQ/Fg+65H0ePCDmdsBuj+pKMSNXZGLmG0y0+TvnZmQso6gYZejbScf1R+RBks7kB
YeC48ehdpQVoz0B9jqKupBVEny1OwOGSRSy8bQJoS1vnI0XFkZHtIxqGfsHiw+WQSZAiC4m9jtMb
JMCTQLNBJFgiR0SMREmMFZujz67SEEi67S1elm3iGqB6Ug9vbPcoiNAoZbeVtQmivUJvqsJ/CWH1
Z/GcF4fc9/K2TqGinWnKVgRxtCgufm5cCYjL6QgixSkbfD0bC9myXqetwGWTdNNUpjq0/pDkuywX
U6OXpW8T85sy19uhwjP5Z/aaLvlYRKAM/1DZvIh3dvaGJoDLiBDPWBIgSozvx9Y04eRq3pvOBeGy
lLNLM8D95JR/fWG3kZG1aZdJrjnnZS9dWhPCAKZY+mabUQ/NQsSUwXLS0Uzh2hkC1clXVDC3cHvp
nRK2rksQdbN+Kpo5NfYFH4h3aOnDkar8q78lq6pnw9PA8GXdpp/8m+3LdQLMzncICSaOd3ytrMa6
C4M9vsTTlnbiH5GQLB1S+dKFab6oejVaaFawHQ4vva9gL+Ojb/WElW8b6sbwTmBlVjUtG96co7pc
duVaHgvZfT1uZYwAHDHAUhStORaK73FIVBXQOQAk6pLUAYWOQcPlv9HgFWqAumzocaKK/bUFJQWi
YZDrOjLFK8ZYuImqbEMjcxBTpbkDvqzBDPmho9DH8sb8mzRRWnwi3KHsOyDN7X9OMKG7vl/t21DU
ggMcgx9Sxs0MpHVmN4PydDjZL2WIBDsYFwjisklVrzXtAL1aE0UjAfqE4iIdHqcFf6S/gCspGcFb
4MrW9RpruzghNXD2TGxPj8RuxyS/ROYFLxaAQpLtn2UUWkams5E4i0TWcVHqMmnm/G+o1/g28Vwd
3uxw2IsOkpP1iMzMBs63GL9pVLb+xtzZlOxD6fsaKEr0O6y3TgU2jejyYAc9hNnsomlwsYyvYbQU
7rKKCL0tJ3kS18hbcffrn/TQWibanY9sjrHKIwc2od47PHGOZvforBRjztC38py2RzS91NM66mK1
265h6fqA+njrBGOGtz52cVhQm94sj+x70Xj6vLtBw4O0HXQqXf4dbHLilqUGIYwU3A3GR3y6N3dV
LKMP6wzaT0YldwsUm3X+/r+NTLGsDxozajehk6slLy+QhAydhMh1cxvIPXcJwNkWWcgTgb17nPLY
8r8yZxJ3FokktXCRE39bYXtB2FxnGNoBrxivk+JdfHSXN9YPhWXlOYQLsQjg4bT0+wYlH/H7c1tz
I0SCbl9A+a0N8HXr1t7AePCPmYMGDDmumlHjswWAUkodJPH2GMp8W1dQI7/93QHoduYt4qfoOwUU
C2R26ilJ4sEhlt7xdk+HXc081DnpVwR2J9IVWk5Vry8wV3CqixKjIPXKAJUsIMsqQ7syc4BbnZwx
KdRJYK64Mq4UDhP3eiRX4MrWanD5dK8TU+F4lcKy+9JNy2+MREr1zLVJtapbttofucWRiHhlDcdW
QlN/kLSgTgO4t+HVvN0844E/pMOfvdzmRdLNxWw6TGSoG2N3dlQoAvkfp0M09p83dmdyrmAOYL7o
k9mt0Qp85+5FEa6JPUTl2biaJJXmtL/ruF6zItDOGwhtXZfT3hXwfWHyKWpHgcOIxv+d8I3xhWxt
XelfCjOgdshElqylglIJdA04/jth2iIoxgeCL9tSnqzCagKyAscckBWICDHEhIZrZgAp5pE1qe7S
Jt+Y6dSUv2TOYzUnrjT50YrzNiiK9XwvnHXEQeecDuuo396Kk6RUNj8ZDqDKfdF1qlJDmc+3oLMk
Qo9xF9mdCp8TlixH8piMaL97IPpmS8C08hbF+LmNPaOOddJ9I2Z882qt0vxAVuRSoKFqTid2nsiX
g5W0uay0txIlbVQOEB37PqyJNZJNc29Iy6L/iMnf1zvQ7wJqJupcxPgANbHIeADmxPq2+bGlG/Uo
FPjl4hXoQJCp4djkiiR1yXmi91coLvhxjX4DMz0xzRDBeGC/n0vLUZPDBJ/ZD6WwuWe7ctL223on
DY3IxGx6EXdwgLCgJlIcLo4OijI/XPLNhxcCIev+PGBCuyCNlONnZMndpip1QEcicrICrh7c2qr1
YSf698Zm99I5rxHPIWdCkKoM9FqlRxaGQZMR+A76aUSKXc+wEtggxg1NrcNbSRzLKP5LngYfPe2r
9CkUEBS4y1XklK2pwzUs1Y29uxa2eAo4D/QvAUAm0xy0c52ND94PRTfgES8ND/wWk5lZ14tEhn/Z
5xME259hb6n4FuL6Ccs+gWbEb4kbHXdAQ1CDYQsgLGtVrF2vi8B0sWaCQqGSC6Zfu4oMjxCN2Z90
o3TkOUTYFgmh4TRYinq4YySNEXIEH36c0JWQtWUwZmEd05V/VSq+7iSHcDHzD4ENm1naUZUBO3qM
Aj8KbCsL5AD+nBzTszMUQwnXaLKGSkuB0NN70He6ekymvTjNAU1TE+TCp6GCQpEnmy85gWLjB3kE
NTcH3w5VR5hQrANTGD+Y4nu5AvHQHFkV20ORS+myZz81U0S9AU/Z6sy5MHijpa7hby8XoBHPwb5I
ejLGYiWn4FrAz9jVe/YPY/uC5qz7FmIgeePEyqtcZ4qJ8jsqMBMlQLMoCEmyQ+MjDj3t135gOhiu
AqH6cVBS/45UYutTBmi+Mss5iSVn3mrc4hUxzOFBebxjV7TAIxA4zdjnViB0GLgO0UUpl4a1Y2/D
iP5i9yTamgdpZGwuLMETjlVtsQx6J4JYpecIrinwBQpfLTBcTo7kv52FRBh7oIPgeBFTYW/fAKYO
aQXzXAeIXsLAbfR/isN2Rsi8LZlfIJbUBqAgJXloXkfLrsi1Qqt/E1auhqHwgjYxycoeysNhkUpq
xCHpDNwnjtyaJkWtLf5ueNasR3NE3YYXt/Vl3FxZqtgTjyFSnx9BXMfP7iz8o7M9PB0lH0qfWEyR
29ncxMeSBeYUiRi7MypTPUs1+EfMdd3R3RZc2PjczPcx73EoMy+eLMTGCsJeoghginRReojNGwhW
8O3zd9JIQT/h/vU17Fr+hYtRpH3eRZ2/Ggi47yWFt2pSq+RmGTBB2t6KY9jiGirjaTM7k4r+lh/9
+W9UrF/O3cU3WAFw0GjFsyrJx26S74h2c7/N3KT4vAbLxdmplCYnB1xMGxNKZYziSKCNxPdc2Kuv
6aZwl49RXgEPRncemApwhSi6ICz/uoXdniOtIKUIHzx/y9rgKYk7CDNzlQttL8kvVLmy9sKCr+gm
TZoXTtfedempFnthuvOiLnKotk6BVwAmlYEXEhZMZe8OqeR+V2qALmVcGrIrO/cX+fRDM3PfImkQ
XIAnqJOg8+2nfT3FMIp3FOxovltcu4uxx0cRmVc1Gh8cnvS88qew9usoDahxfjTvFY1iQlxcqf2k
r+IG1+F6PtlYkAMPGrql/bmeVcogNgjo4/8tyBOZ0CHwLbLFUo490GHZhs5cuQEHR8w5aCYG+IXS
dD5ZA9clqBxMbHAhCh8FRR7E9mJ7dkr6uuxlI+O42U8Bezo+4cO6dt67zn8Pdrt8PaKCerU6mFqe
uCirZm3XGr5kTW7rUGumgVfxs08mS//77s9xiQwTO+fQKFXXOYKMXFIvl/D4PYnfKMRFbWPz5BfZ
u2iNqQOwAQ0CnM1wF0XjJPKBsRP+2Qu3i4aFweYQrmYNIAEd3HKyU6LBrVhVgyTNJp062QRuS5Yl
CSBC6r87Zr7i1AUL25Yko7E5BOgzfngEOVp16qYdbXf55dL/ZQ1FIRMxo6BHukdRNZ9zIyljH/FF
8b0F96l67I+np+OdWgoLAHj8uN/w7+pe0YOSKAn5j9kxvT0h4kKYHXw+N5g9VBO7lHdZPzGvVdH4
lMN1bWctbU668Gph/mbfY2ay6qX5qQCYQcvNA6DEON6gMPiii9ibz2CCvEtZhJNdFYXO9D5Jwo1A
SUFgruHEyQoP6+poqEzPgE8J289Cz9n8KdaVvxS92yytX7OagbnyifTG3JBkDHjSS8tunjR8xn4f
jS4GOPuowzFTtoDiryo7Ocw0MismVg76g5QmRti1p/pOih3ozjMrENw8t1nQD2Ee5sDX8Z+G/7B/
QsZXjWXK/6NioH3bquhluSYKUbpIdsUAG1ysA5ar4vR5WlcsJ2X9PV9kvn+EBBCPd4nPt7YcbHST
i35dpHKQnRbzxvFyvefvSmadA2MItroXQRpR05o9hnkqYQu8EJAKbksY78eZ0g/3ZV+Nqog5lmTu
8FG3QTB5KyuV8wgbf4kIxE0SRUqMtLHbvZ3dAtxFw/uO/6lzSOmCIAg0ciE0cYvsmQ5uF+W6YsZ7
TJaUypQYWNxJHMYf6aYa+FldFvjewGjuwIgrO51jrL1sLdmZFXxRxDgWBnaoH14eZ8ksAmZtECVS
9G6NIn0E5ZKkEXfyGVdLHiM95d/QqXxc/960D4Cav5QJ3ikk5LyMtF8T6mCFag6LBxVAy//HZxEo
PFezn4wh6oYeoMXwr6ASikQBHWVKsy5qXc5IpRIjnRgKyO0nZuE+1l3ppjcJsmAmlNzVteuVoi+V
v2lnfaNhEBdpQX6e3IuU73CLqgyWxH+HSWeV9tnyG1iWsb3RkuBaU1R5GKgrcVEDKfMW67AmQW+S
ceO/6wpepwOT57hcP6YoULELIz6VE5tfRP1MnBrZnsiUM4l+xgbQ9kUOqQmovisk2nuTQME5v0G9
GVWwnIqxA+Z914RGgsJ61ph1eLv3kGkLY5QUnHViJZyObczID2F8Kh2tJaFTrudBODD/6b47w1n8
xiGK1ISr5EAO0ac6zravLEOKeAZyIyuocXm/PLclayjL6eOvGp8MupC3mp9gOUQraCBMfmWGWjY3
vHJs1S5CCTJaBJcZ4vdTBaQbhVv+ZHVUkKG+ndFCgRhHAGc+bbn6WA1rC86Qapl/WzUQ342MU5/z
/mrsyvdQkEzg+pUlvlZcj3euJLGiZmVaBO/Rvd9n4wK7mehp7WtJfyrxp6NdEOgU5+NY5ZilzQL9
gJi391flCVn8F5bI6Fxmc8HkpOy9OEiXLSnaUv09WsNRL+gZdxKhSsl7SHop+AgqyTgZMKYH0HLf
mzfW+UgAbcTv0EO8OLbEJgDy6H3cqfhami3dPt/hqTL3PZusoLjevu/PCy02VSP8Rc6HIY09gRMz
OOwWrtqP6Uuf5yfL0jUgdwRaxxctpeHCALGLBYzkMrUTqWgMacH7DIgAhAlGBfh6LAiO8oYqJSjp
ZKnUBdadQRIztWlRjTu8prpWGWToF0196hzeNCdN/3/U4oDyImKZ3wqzeRsqTI9fsMkuCDChi0RY
jd749qced+Br6/cti7d5PGejTWPsdU2I85kS/IPEDG1Z9At8xDrL60T7vL52ej8tiIwSyXrGNbj+
SUsC291EfbHcSNavaqMEwTt76T4v4/8VgdTQBDQPBAE48/OowImQlJ56h1lzln6vEFOzXsqvzY+R
HEyWwmq+wl9juzlIRrOR9xmUv0HA7lxLMryDO0vL7L+ZLgtMORJ6ZfwmDYSXpIZjDqaEWw5RGJfJ
l8xhdQDa1GqmsFMV2ggLy1SYDQZjMTNwXOaMu3iHjJC+9FNs33XTFE5EVQOadWVU3wfzZSuOAk3T
eHKmHUOx5sqEQJ4zP507SzpoCoT3bBVsHdn+1J2l4QHecOQCfCN96TeS6IPzF8XBQOjdrinHuepE
utGKvgfOogqgbofxvxxU5zdutTf/2CMwLcnmAv1/GrsSRM1kdc+DkB00iVOIYTink7FgIKLIbC3K
O+8DPfHAaK9rXWW9HhwEis4Yc1czUq/SKUE6d5tvol8XIte8ILoR1f5y9xt5JSuAm3KsHOiXgEMV
FQXxyCN9rsSq5Zny++hAXdbrfKBqXNfq6eGFtw9DlKdz+jlt3MQ7FJR6U1NWrEAqtgZwNYeEFDDK
gSHhUma0KbIazeulKh3ATEVF1ChJQE1bjIXQjmeYUtsRXC3YQKqQkKVdmHn1peDBuY2R+ji/w6OO
SYK0satJe8cjwlxzS5+5mlpM4d9a7/o3OaDw+FzsQgdP3wx7YAQgTRFHbMoMUlurzXfcm06GO72Z
kK3gmctDZQq8ihhq3Kknz2umSSWs1tMoVbtBwn5tT7t00Wuwngsh/uTz5XwsmQ2v6JeJPNvppgaE
4AAaILgk0hk88iCu3VIH/G9Hjy6KRnpQ+gGiMlsExKIvzE+g3rgGfnouAzolhtbftYPbSNmzvgTG
Tw7SUT84w619SJu1WwKiNqqJmiV4iwajCJRxsvvRoNMZrHwNBmba9uXcEHnQsHq8AB3eQS7+G8u7
jxF+/wyaYnhp4pAHVXwqRIOYRKKt9VIeC5+yi5t5HCSWnObTp8iTQEHubBpphykWzMkyQNprEBYP
Yj+QcNg0MrNiW8nM6uiRgg15l6cPtnleXy3Tq3TrKkdzVwa11qagWk98J+aoPYX7BGVFNFVjCLpq
1BqIszJTr7dAdLXletwITvSVAN+81h9kkdQzLJUD9u3YSTAGoena3b8P5AeJL5AirqZR80OZjalC
i5cr8GhK5AeU4Ll8NpkwsSW9BDR6fTEr6jtjDsKSNHGjtruN3299msI/Jq80iYs96FVNjVb5fdT0
uQ9eFO7OrP75j1jvhT3PZA414wRqcqFomnU+44zdI5XuW1/B2lz8KU6akfoVJo25i78K/OfMedvi
GRhXFM/WT5b6aSwaMxmWoYTYgDD0XZ128T5NGj1li6buMZQoOUGZVEjS+bTDLfZBDUU9R8h7aOAU
iVG4mC3CEp+jgIXX48ugPgMKh9UdkuitP7tLTZUv7xnnfLScPkX76pns7AdXvlIpusVI++5fxtPo
CRf2Tkosmxj1r8IOMnFvsyLj6AuXGhgi+dlRS4yJDKWqxsvQ8k1qpM/87UG7idcrH8TsyveDVcae
20fhseHTcITecZouceWcYvTqcP69w71X4cDjZqLUxXwqb4D/6P1bD2k8ZrDSQ3bUyHxSakbbR7d0
uStZ1oD/rxc7108OoHXEKSu1uPNWy/7Lqn/iLxFu6uuoa3CBWHVYMVyaAsIxRMnK/hH77rPjgNif
wy/q+XtQUwx56DvNLUmJeuSOWp9oyVGXQAoblWYZOrJYUwlBRWov1NSbG8FnAL/Frp9epcF1Vdcn
/8Ee9LxWZHe70mLzdkJo31rTmDyqTQ7QVYd6joofuqJCD+Ve3gjRDrH+mES4Px03WKjVGt4HKJyq
9/uOl8FQj9QzMSDl+6ikNWy0/We5pwSmo2oh3P+YcGf1d3JFYH26dGCmbAyqSqjoH9faon5DC1Rk
x7QyCsm55HAPmuGFj7acc+SEL5k8u4JDSijn0vvElwskUuq5LAojr7UJXxrKj5hQxTox6Q5JRgsA
2rpp35IvHDA4eTyXOfZYf02xhHc6mdHRecdypceRa8ppzgLGORP0F7MDqvtgzZZQTr9nXQO7ePD8
KKvDiD2ljqqXdqXZfLstD/RgC7+po+/3dWpSvjGNX+Ovj1syK0keWaHziuD+m5aUnbVoMKrpHkzV
9kwj9hNDFoFGwU/+s3bf9yhHsnNk4cKD8h7IOOJy+4DRO/yofqO/x6b7Dm4xT1CCYNaHPWoiHGEQ
1YCqwv9A+2u8l/J3cgx8zfMj66Gp6bzovWEKBGguG50jancz35Qw7PfazOo1yFNR1ehbUqOfa86G
jSdv4aJiUpN8AnKGSeSJoJVlL83GoB/v++KTVSmkcThN/aqtAw6k3N8gTeFcPXu+1R6JgndeAw/M
Ez8ecAqFvriFcSimdOQbU5uFiYWYerhls21ZkbwnNsMB9lJCXe0W/rizvOGgS1HzDRLS4SzZ9Wh/
2Qfmq8S/p9AJJO60/Oiw2KnSkl296nsupuuzANVefKAHmUEHYYhdqHafcoVG45/aEEBDYExvVPAJ
LZdM7LKiPOCbKACpOB17Jm3WBehtfDTCJODDpkzfsT7U5cc54TRuOo5sSh8XpnWA3HhyZEbIQBeW
jG7wJ/SUxiCxGzNHBHlub7iQW2rDwyD/eK6rj1H+b7hUnzODEOqiVWOP2JVYjJvxEQBwPfbQl9Yq
AiBrLn0GFqOHdgGxNgZpAeX2Fkm1hoBdyHCZiJBKBN9kiNEecZyjhW6W2wQQBnLw5D3xRxuLyJvA
exaR4RZZqmQ1gmMt5Q7a/FOq+tIHkKjdMmLo3tDQ6SH0CNb4/rD+gbblIUSByjIX6V6qB0CxpJSL
RlH7+L4YpuuIhJFaCCBu8L8p0p3aBFZgfF11q1DdJ8pn75hI/psp5IQjjHg2a+9OWRnKY3Vwv7P5
pXP/4p8LrSLd4VGI09sIHPgKc53FwC3AWCm1QKXmfAGgqMcPbk0yzd5YO/ix8ETgatRP3wBwOtVi
BVahjqDKOR/ye82E6fvMnm6BKsaPGzwwj49AgL1varfkHczIQAI7wU6YngSOelWkfEj7uHLsTdJt
6ON0mpz/3TutckLKY/4ocaPJ5Nr+E9S/d+1/HjGtckL3r5xzy4WP5RdPwiSySB8X0UX6niBEWgU7
P/pavB5tn+rr+x+SveGzj2Avm3S/VWwy7edSYnlyAD2lsjezcVzuULv9/VAp2RSAH70a0tRm4jGB
jtpZxr+tRIoRsBg9ydbM6bx+3WPqmF7adACAU3qIaxeeFhZ1CuDWv43djtnhstqXEIZOwRB3LOXB
nPEEeAbD40jaLetiWwFKlBktkkLOVu8IavB0kStxnF5FK6fih9y7BcolXudtkQkCMaZA0enz0+qL
n2Pqea3oZP/1qsj5IRdSyBao7ny7dNl4fPNCNuBkFTNXjyfEgGGUy2BDXz4rC3/0Y8O7mMMGhaoM
SpI3zlNe3Lo3gde9vAIEqlRTK6cHv5P9cJqazueiZmFVAzmacac7avreeOOwcxg/4SqsvlJc+PXc
KT3WRzbBsIRSNbFcdEgtuluOwJlG7cf4uDr4FW2qvIqdImkwSyaUNk0tYn+OBsR1Rc8TmqkzaNNJ
j0fNG1wjJoDPvXcGnlYF9cru+uj6LDTAXrq0U9h2KIi6SYVpqdDu+aIYy2HkeUKtwKNnwkdXu/NW
K6wDQOgTncazrJeoUqA+7R3tybuZe8Lg2nAwVv+/Xr9bggeAZ7LVjqROOSaU9PjKIz+WhqRQVSdB
tkvO1VE3AYf33euxIw8Z253Q4XZ/XkaHUfFl4+8DJQ9t1DP8hJryehjf5c9xHt3+lfLtJz9u7p1D
GBx1NqsdNmPmW5LVubMti8f95NKn0e7lWuDpLfWmzFF6vOZmW5WevuPVM5kBSoF8oruKZ8c9uoov
VYZPtt0C8+O22TCZCdq/bfDp2txZHNFaQoPhqz6tv8PYIsHq9ckhF6TEwOL55PMXFbAE1tV+J5/u
DN6aN2/Dp6Cz8ZFTPkIyZEAFMf3ivt8hH7ZvGjxGiEFqwTI3F+ZHtg+bs/oDqyTGGzag0bSSnj+S
8FJC0zlfLqilwZXQHLwnJJqyAv4mCcKJnzHN36OaVj/DkhKcc9OvJ0shsB9cSvCidF8/1aXEu97i
LNqe54a5wP9swG8qUnDg9xmgRBtr7d7Fcg8wZNdgt6cHBC1vgHvKyMWRIzRETXVGMaSNxwjbovct
m1u9nWiXmiaxZxLXh4zhXFwTGcZ2Q8RhahG0qpS9861Px2GWkWwXecXsm80tkifQRnDPKQJ8Zzzk
pZx19S7LU5zFDTZITBkG8LMLrF3mKdHlrVcGv0RHjCgLk79XGlbW5WRn1yGGCFFlG5ZY855qydEk
5ostpYcw5lX7hyakmOAywKImRFZakfytBh85Na2jfrU2E/D8o6afq2MjEJJElA4XWDDQZRPdYvzu
sO/dtpP+rk+UrehqZz5i/ZZSNVJFuuhZyybPPO7DztPpdLd77j9A1iswG1UB269d5+GC4RXtA2X/
lSI5rpHhfV00HvoLmYCRsGr4xLlkf+v0+8ygwy5Yx9nL/1NQuYQ2ASQ1irzETw9bVC4XGS9hINZ7
6MIBn9ZlekvumHNPvC/eVpJ8O4cs53gJiABkDQzAmWKAyng/pwsNVKZa9nx6iwXNLAYSW8hR1M9S
KovKK6H2GaS8bA7hDaRC57vA0y2WhyRm4TdNBWx2k40Z8ptbxlcBbrpebHhr9JpuQXwlcIWbtduO
oVwbtBE+8an+ikND24Q0G+SJ60hjaSwxwAdNE+xWSvxWyceRzTv6fdRhlxlMbsS1ePl4pnwvYUdY
HDZgslC482ScjgZ0kIf1SbnifeyuXkkb5YxvWAjmgBeG8coogo+zwSiytk+iz2qoZHpeapLnOCp5
zs1WQAqCNH0RqIiGlqhCCcrOoRerO7LCykzt4Tvhe/0iNNfjy/o032or3exuU7eoPTp7pjgsaweE
IVfY6u51dEE0iIOb3vb5NhUbjJfN2TGlpoDnzAz9+A/qgXdNSDJsOhur90vohWtLGrNnhWaQNhEA
UOhHt2Az19sZTPX4HwVc+1xdNPrS52HkbGBPwjAqBr4xsOL0KaqhFAWm3ZIqCvTnZ6kkTNDOp+vt
tFtuDf2dsmVf7r5E1gfQyOvdYC6r41aoDp/9Q0mxxqExC5/GaCdJ9xMi9jNM4ivExOvhHWAEiWvZ
IkIS77wbrbOYCyVdgH9HvTs/XXDCzzwlX1gC1VgS9qrbmBWQa5+QVvsP1MCQq3FapXmLaasU1SK+
8p+drUjYAvNyWLYq602gESNFTz/12TcYcmfVfJC5tAKGX/ocT0ZVox4GyC/PH/0ywCAGou0XvKoP
8w68TzR2waLr23Herf4A+i32LCa+N69lAkPzxZB/LazDkX2iYgETiHzKl89HHlsktKndo97wNcV7
UNT95svaWdc7g3D7JDFkQpkPY8qYLw4lv6uSledeMH0rrBlLzSCVuET1qvK4StFuuzzSAzsGuxlC
d0+TEVoOBkVO2T+g9ynHwxzXunsJ9Kt9ciWG8cnh+DQXWUQjN3c1GL1uQCBUT366jDL9e6KFJBdR
o9La/6RbjVhJPYpNwn6eppoE9wJE8cjQZViaxP9jf9l2dVGIy7FPcMhnvmO5KjOw/LVqrACj3/2m
x4p3qmMQ6j1BPUeI9ijcdSeisDRGO7uc8ZV2Ji3NCAZ3Aq9pj88pK5BKn7LuhOdVJ9DQcw6WnBIG
UQ+0BbXMCOG1/oL6m5YlyaLqQUQFXUu0yFFoRXSPrvRKA2TXXrVD5KUnI2HBW/es/7mIjhvTVqDi
tJevPsAY+pFD5/RfH0UL1zWjPxo3TKY6uA5md8lOp824Nl6BjokpTES7f3wuQTcITgedXlQXwAmJ
wkVFBIynQmaLYY615RFjxAhEO3GtO0rv0DuqVo5pKSICXoCE7yMnI1AOt+ABVS4hSBtMbPkztSfa
m7n2RXBGUCMX60rAQGUKtM+irQ6/cUVzpJRwc+SjQAA6fVj/jkcapJcp3dms8w5LJCdwNoBkSkoe
7nOzAMp/46J8y1Hs2wFRMD/NxjtVfDODkBcYgUPdELz9i5eZTKWzop8l64IZIDD0cRHwcT7FUWWQ
iYPrF1JTywr4e5GiL1AMaczoMuNu4r3l2Q7CXGeWkPXrxqsRJq1wRp3jFE8iDoy96ZkhczydA2IC
/QxNtPd9d4aEnPAcVio2OissdFHpxrZQcIkTqQOj3e4XKtIYWGhT0+b9igUq7Vmftn0bJL+b196K
LkqRTgpUXsnnxxgB6f9L4CHC24TG3jKX0spd+TRDNTdJ6OkOB7oaDT2R4eui5vJWo67MgOJsyzOZ
9Gwknom5w7A90kKnSGg8yZASMdF7wUxIjTpxFEuVVYEFJqRV60HjEb201RbdEaR5rQ2YSNJrmIDs
BLBnHmA5A7FgAvr9rkmQ2Ke9gOVZ7LvR1S9ImCqEmALUWDqR8a0cGW+MQ3zTYRppWY/v0YW0lDK0
7GVWxFXAUTR9TmHy+AwTPcWuY/bb18/JfPtcQFeRyTHvzWtLNkuc49j/VOJm9yQlMUtYvQ83iZ6s
w46+bG6yfUYXB/BJb2TMrY+KDfh1ULXE6W/YjYkA/ZmnZ30vIrQ+wuMwAebI91gBtU+w05wfJcmi
M4uVz/c6iehiiWVzCmgYtg8PJxAgiOtVGo5CHZzZBzsGHWJsOlgLwh6Ds+ELslXHe4dEIz6M1R/T
szi1CYpAkXV/ZL8QniSnPFbJ0Beldk/WVcTl7dzW4qNT4oF/fW82DCJD/68/evz6DgMb/+9PF1kl
KJhYFWu0+1x0dlGh9C2RF0bO4WNmxgir4QryYrWZDstv3hAHb2V56hKZWVnje6R+YSEFoxrnh85O
IrQg/rpPnHjI0rwY0ip3pBh+DSWVzEd5M9BcO6yVl7nRuyj3ruObHxRb5+c+igX1Wf4JfTsfBmrN
/D/HQCaKRg91uHRfphXiPpjXsaPIvo45ww+ak/CaiVjbfrhQ5wesHMy6yR5dES0nZbg1Zs6EQyf0
+wK3RBRjgNYg6AP8S4o8I2oFj7zD9q7nSYQzs7huz5fv7zcmDFiNei5omjxvdvt1rt6cFuDMUnh7
d2ic7SCYye3+Xhqsz0NfgM6ADfhfj7/OO3y5w6BvA3eG0iMFYHs1GKiV6QGExgzkwpi6GB31whbW
xMr9HOHv2T0shskcdtGBgNu1Kq1zvOznSP4l3/Da8GYr5SxDr7LwweY+86FLNGKZShdmim3+vzl/
vGM/fmvwZwWQFpAtWNdhw16ouQxF2llZh0ySXlX7z9IDj26dmdhyCkde0l9nFu9FswMJtPuBxYuP
7Cckw0Oes1OSdr5wC9afLT9hiqqZcsL0hjwizTxuDxA+rhedzrnHIV+43C6bLk3cuzN9Ub3UZ6cz
XZmm68Lx9kOx07Ob+8DEfqyVNWt3u0gbTLdz+HLyFwXJTcI1sRay2H8pM7C7RoR7YeOaivK/eJ/F
wmVizpoIT8zBNrskxXSGHKzB5NjZpT8uV/qqJnPCO+64Wbacf7zJY5yLTZ24c70aWbGyVW8uRodl
0wEI1CRggXHguxlmfcEIBA4CYRsRj50ykEh1gBP18aZwoX573ULLZmjxQE0a6MK/ngv1NQ/O9Kt9
3bVWcj3+4OW5QyQq8J8JLk+OrW3RZcI/Ap2MCYR7i1AV2IkGSixe/8OkS0/wHxzx+MMxfT/ghBcQ
xNTELOgoJUX3GajhiNMfp1YY59+VufZg9TxlGLcvLaIWG+xkWNEiQ4UrJ3D/YJYgtWrH6i6u6CJ8
7qRfg1HAy90oDCwA8k3IEU+koqTxr18PIPZ3luxQLCgun+3ex2/VVZEOHXIa3iiz+lUi5QLTHWgt
54g+7XhyR01hyip7DFp8jUy7g/kZRb5jTZ05NamYnzprtM74NQPFBlTCjPC89v8oAgBMekFnlErf
/Qu1GP41ienoyc6HJWakYPFniBycGmIh3UaPtnU7ab+0oH/DB2t2cBVLbku9tI5W4MeAqCD8GZVL
JsIyxvXBUr+tOFoJuMPuVAx7xbp3Vq+scQNQW7YputqIOkcfpw16kHGFk91PW6isGOYLHHYPmXcD
h0zN+2SO84IUtFEFprR+/XP06tI91z97Za3Z0G5BUcmpQ/a4cex5qvoiTNW6M7vPdLjlLCpwuJ/G
Lw77SbfWHFe3XPo42GhqNuio/uEPH+eQCA1J16cqRPcYXV9PQOq0rDEYmgBGW7UdSq1QjahfEk9Q
d5Qym8HDGK6whNiPm/gd2boB9u2JuSXO2LDUQ0bNmjekY2hWRMuHeUixkjThhLyxqPLN4EXFbvos
7pSGU6aTZfzq8wbM+rcN33ipV/+8t9aLt1xZHArTY341zM01EzeF8S2ISBXPB3m3u4WnLCkRQXxh
vPs24sSFet1B+OB+X7QYet5WsSIu9vdrN2gCO9axvkL/2ooGJXfQWUZn44Yto5Iws9sWrRM1m+KJ
sLwPcauOjGVaQT7lOzfp3XVkb7Wz/jg+7pLswEwhiM/43Ekme9wOHStzUjIAOIO9XfI6G5THo+KX
PInZHdj+10079h4SyX84sIUeaenTkkpX/mqYlT48ETt06m5xAUB5jAgztwNuefGU6ndYE7/W0r/t
P1ynrsFpqx9GukGA1halgbBw7IAl0o9vPVEQPWlQtfYHKyPGCr3rucRq5dhx6siep32w43BJxhBt
Gmm8UQV4Qt94uCZ1TPznNl/CckXK7iDFv0mqz2jjSoJjxdLn30fzUtYOrCHHh0nlLKdvhqAwU6AF
CC5Q78rcYJoAUfnwXxjZIP6Sc1sf6PCQaOP0wrxDG7r6syY242a/hhOxRQM1iuIWjquE825KBbUk
m5nd81tsFI8C8sAg5+CzO20hLEeUdVXV+pTTGEIhdiKaPXXXXRSEDVtNdqGJ+AW3nmjAb7SxHTmw
9G5H2N5jt6Hh36QyG9zjxCOEaGUTGFJl+K3nVQIgqfocqiXq3CB0C0hgufgO6m4gD2L/DMGi2tWt
o5VQGMdEKhCtTVrvmXNDkLVJW0NnCaznrYPQ2LcxMINXtBHnC0iYgG0p0KA5ElIcLlypYWqbUx43
N6SvXodVV5zwlSrrbjBZBeLJqf1Tubqr9q8Fc2zjiUiLD7pOjxaCoDhOkX3WLRn8jlZX0XEXr1Th
vohC2qBREgkzlTrhm52GfXkY1fLzWpFirWaMVJfdk3dkNV0lyb8cqfOQKGbFc3qca36di0cQg0Ol
q5jKWSOxkUyMb1UMxjdUUq6tny2gXe/WGIVIYgZxw4hGXl19k0Vy+zCF/i9DeHBqx/hQSQc18ig1
4I2QSht1iIW9LSo6G/iQ7d0SCt/ysbnSKqwl6ZBxOheRozwurQjDKOwtWS9ev1vrGCRSJckx7cP6
ZQBsaoAQkifrnUELtJDKmjDGxXjnOc6k0RjL07Nc2tY9boPv09qqNsO0aFaDHEevKgVh+UaM1Ji5
M3MqVjifXRh3c66ShpINrXPIyCWKkX9KQQ1VlvhNFDv0jJG7kDJHshtNX5Nx4mOeUzkGV08RKhNi
3njig0GuFS7wpMTxjGuY1to/wrPN6LRWf5otlo4lOgbFM1EO1rWyX4ddwmyfVAwL1WNIVbZTRzYd
gQ8pd9RhJawMHsxDn/BItqFjqbdSX3T5cER8zoki/TMd66Dsr0Vp+/xWqgGOBv+cMz9wXDoO3J7m
6Ci1mjff+5WXCnyypbUSxtEWjRX9u6wLh5Q2JeZwk7R6AFdku+BiDMrY48CuVhmpEiSKInIK8q35
aIP/8qa1+peHWUVjSIgFJZFATzpcU81wrtU/SHXyLR5vRYh+yCfgE7eCHA4l/kE0liPVEaMKy6E6
oB9QzRmF1Vag/hQG/30wWLYdNw1tbtu/SzNm8/tOyC2viWs9//dnqEPXvPWz2vEw3jL+Be7luvf1
M40vnv2ou8kKia8Efmmgrtjp1iQc5aoMFvm1MQtv6DwapIIpG5Yr2PDMjT/Z56GRknuYPdJ1r8sG
uATGwj2o1iyW6G34tCTc3qUAfS3Kl5THirKMdUO0kzawltFHMxhEEZC2POS7W9AQia9wW0oN9H1C
cOJJWglTer1G/iCusXAsFOBXQAPDZmUyLukAo7+Bqifb1bYSJ/OAxxZBpyjtIbhVz4pyDZ2K3b3c
DglR+HoW367X4L/zM2kdSPpired/IL6KhrfpFBTL7fLoMJ/uFwMPRdXkPgHU3orD34BP2Xg001Dq
11H+t4SSEpCGL82GjHkYKVty2ctb+XnMxCy7xPyI/qVjAIeTqXSkYi6AJBGgMckKx0VIgsz7tkuo
d+7Sjk4oP7bbBWMCfSpct70aE26nHZc5rXhiR2rmpIfXG5V1w5qL1SmGS/pg0qyJ3jdlYTe2xJJW
dyQbTq22roIWcHmne9z205kbCbP/PAzyOsX4kNIhdtojGEqMmZm1v+KgPDTCFCUx6Iwc/Yjnp0bG
9jebk/ptkbTxKsJCZ93yHry9HD/PCWiQRAmcxvbWA7R1XF2mTL1gHN0B6NssApqLjPB+5oFU5Dr1
0stj6hoyY9uMhcUbUQ8VrXzQDslhmMqR+dI0LHvI9EijVuBmqSD38blKLF+erTFW29jlTF/zCurS
lCCGK9AM6QCwNXe+kQaaTQG3U04w6VHpHjuiXjRrZyQjKkoto56ieovLp047NxvTLnbb46Vd9f6H
8qSzDVjGXxSSozhUoX1m2anjsGt8cS8fvQWd46kRcafrmAGmE8QVWigp7mLTObkQdnpTZpAi8ks2
NObEOZROZuBtqiRFEypAsgZEHRErLpQXUoxDVPH3YU2ivUQP8exuNiNrzuwz3OYy0nkE7V2f6xyv
EX8JSo1axulwczFfb9VQRDCBVsEQRuppOyHP/9Xpci4pwVjMFEvJ0OWKz8YZ7nLxbmt4GMvZKJf+
+irePl48l3PqrVhXFMX/eCN1/FGTD7yoRv5ouZH9SeevqmmC4+jcl6aVeRpJ8TEdxdrgSCCiok/0
GLpiXZYZY6jENPv8bUZepIECnR71WOKv/evpIVG4CXWtHDA9psmyw6tbL7o2cJQrgZ0skVEVGqr1
J5nDTj/c0Y678MpOHVYKlhQRO0TlYH0XqvFbLkQu+3581zdu1LwsiXdKMlJMzTrMbYjBZ3+IgzAO
U/IX1cMA/dSc+i7rBSEg55b9UoJsOpYNxXTOjqnlfz0cQlIPQQ3ZDgok/BswxQjv1A7h7qd7dqHc
+KOI6Ijs/2hUnXTMjUL4mAmczsCpk1T7jZUlEF/tKhaHiK64AnZyx06Ilw2BRWOzFulo/FhgMaMR
SlOElCW15gX9kcNwtLZMtZ16b5DhdTpCNu4y+nsKa3qWWk7oP2NMMSqVthbnTPBXQO27/6rlsNPh
JHBSQ1pKNLsPxWNsiRlFagHia9BQ+lIKtmjwWgoIQUKpXkK15wxv2mm35BCScsVY3D9mkeMmuF2m
5qF5ktcq7/WIg/GD5oj9ZATjQyk4V6dY9pU5SyIj3p5fKEQ7+5huylWE1z5FTBfwqTSxE44tytN+
nhGCfmOLWKeD30jLgWCmYVmXpBW58GN2O1fUgiwU004/yo6Zoq5ToB0e0Pkt6NqXR2RJ7lYsN1wO
SNSD+zpECwf6j6YfZSX4OKfb0Cb1LTdCFBqKzIKpZr20WWROtRMrAdykL5DX13XmIcNAfzParLBK
eDMAdW8SpLH2fWDBN5BYVuulZD70FH3GRghmvMf6Pk+zoM2TVUG+Vkhd9MV8t0w4XwiXi8/nir87
rINhQKm9Zj5TeQNlO4GorFEmmT7upNPjndZJ/+h0MNfFEYA6i7UGL7r24B/CFI8blx/dOkEy4ACA
2lqvFboDq/WL8nqMUrqX9sOByzFf4uU6/NgSMGE+JaYc/Bk9GBJV7j7FgLvrtp/stkPvjYW4nTie
wQQS3Cw6ra3nGgqDffHxQUdNQzp+yy4t/IWs5tQ9k3hJagv57GEo2ryWx27A22quUx+A9HNOcO+B
XDWJNszBFyeu+iNahjY2NEiUlvOWSPXYZZ42Hv1Uh5Cf1UDw5IsVBQTYn/cIIOjpEbftW03xDH1z
jTc22jANDolEjuqjqutkQGaSHa7nQJwklGkj/0DVmsDi0glWp0diCGEsl9fVAudJ7kFkEp2CHhFc
WDlRayMxj6FgE4gCrWb8Ee00ZkBxHcNN4gSj9kf/9KymXsdJtkrSMKU898T30DkpVG6PPWeBGDsv
8icA6vxKmJgZVGscaOJzVt/Y6eJQBJUjrOZqg8PPLAFsKhGkbBaOBnM/Efs3h6/yfSPHm5N0NR1p
Ecd29AaTU/rynTTYvVuWQe50EDAwBh2Lx6HcaQ/K6RFXp5OPT+FdOyvuGV5qn+a1/xLCl3YDA4p3
WXV1w49eGQH3sTQFbF8eoOKtLh0qO9rWDLTzAC4hBB2irB1XOfFKWJdRqNlJrW2YNNPSP4HnM3zG
kCRr1N6qqAhpaT+GIeEYKJwzMtZPZIgLdqpu5zeL0cVsIzogra/1ZpaPxWrjn1Pqz0NtxFTYlWmA
9qJBw9aIojFJJWG5TUCxz5D+41EZx7A64e+MBIUKjLGF0HSVXPSWD25Fv4aveC2ZTzo1GP2ZBS2p
92OuenjKVcyXiBRYNz/olYqlfaKqAYSSbHvtNeEXcCltaOVlFcGWoE5Kr30BO5+HHIm5BJBM0FeS
eaRCGUPmMGjedaAILUd+sEiJRdqE8775XhnbpsofX5OuFJ6Ue8VEnahE8UtNCpWbifqO4DWc3phK
qJH56rRUDBdDHvunQMjJnsX77uZbmnOzWhdLG7JpmlwJhkVC5EsvsXEsLgzXTExUvC7M8fZ3DYu2
KdIUvA6mLCh4C3PC6xxYc0jd4Kvehdx95kPWxvy0FZDfZjVNwlm3RhtIu3DPfupuPXjtBOxk5Bdm
onZVIqvcIz/K+LSPIJwqxOMqMpBsaqNdx4tTyPDUx7zfeCT3GLdKiKt3jSv7RpuiPnGgEFSwV2FD
zz2YspaPxkBKJ35P29uvpROJa3jyrKEueR+ardZSaPa12kka7VP7KMGi7uMujgaYletY1KPtfWNz
zylUz2pQeQ7c6rCF9Ex8aUA36evZcff/eiNtYeKTWorpRb1/QYbljgD7PIJRe9a67cimKRVQsi2b
9bwMeHFOCdhx0lEBtva7WeZsDNkHN208uVobrXhxjnSzqsZYNrDGKKXbWmTyaeHb40Lwzsc+/CFk
LdKhudX+7G08eFzyjQ1HqgP3MXpZ9bnRAqrOiKn0IskRqjh6ltc7Jur8HBM+K2gHtFdlknNRLPqB
d/8HKi2KnW3P3Rk7PnKDkRepsiBMW4fJhYEljZfLVlthm5aARcI3LMP3qVmqXD8qjEW3ERuhOmre
Lb8bkRJ5PUuw5cM+tSF7ID4vlpkcbZCIQCOeqSoOMZ7vARvYiQl+vf0AUwp71gh7GR5NwSw4kX2q
1mT/SDU6qJeYZ4sP4c/4pYSsrpC0SJ+/knQ6NYPERa92XYlUqF1/jG5ixZrntV+rQi9Dnt74zI5f
fkCIEt3sjg8uMzrC3oB4L0wi/JU6/XMFNWh3RKcye2KLbbvJf8fCUFgwKDrTyQsnZL3Wplp3gaPC
yVvNcs7UaSCUJaMhqZhPS2GnLXAWqZz2QJEgc0uDuqAgBjTO8BHhEhnVK3qGpQ1Sm2BJTdOhWEu+
5dLyEHfW/p7NaaD4KyzYCQGdBTDEEOkeSjV0cxgEawxcv+nbcFpQ34Aac73r6KGpArdv94qTkQHk
3fraEpEZHYxdf4tu7NDo6Vr8a4kSHsEAFVUuOQO89IIj8Zl5mJDw68CR6AW4Hd5zgq7qztj6cyWQ
tEPmwClf3ce0/ZuhdYvNn1JHyYGvymJjG92EDKwmsx//GzVVIVSZOW/UyM40W6asgCCoNg9MRaiK
xTrd2UmAtWHagA7JyoIaYp+JL+U1M+SLon/VvQuNHty4nt98zZfv5XKtPFksU2FMYEjApTWJUoPk
U4R1nUdyU+CkTRHYR2HCZO4eqGI7oAuehS1UIqTz/ouQpmvzKGS+Vqc4DTA7Fdlcanx67Ip5jXt+
da1MDbfV8yXyEXg4k5uIv9PxspCg6R+WMpewzx2PTbTWWBAtyENcbmWHL+W9ISpPC447gb2JyELT
wFoKNzFw7ut1bQOm0MYQbbQC42ZsuPO5VmIUOTClUehZi68aCgEbkad9Smpx0aicRA1NFyDL5lFQ
OFQQQgwBeRbr/SO3DV+4/v4DHce8+JoT1OlQUD/axe1ORm7aTZ0rRguvk/rpkpHVp31bHd9FXUY7
3r52pdBFtv7cCPc+uMNUV8FROEAunwcjV1QLKGUCvkM+MboOTsEQh9U/zGZ2skiWvX6YU4lA2Jyl
Sa1B4DuyAXjE2adWgfZEUpubhKH+D/q9V/Uq82U+i4gl4X9doXzXehULvwguYSFVzkuveR7I4n1V
yeYFVTuTkp3aav+9ZC87NAgytubFPuAppmpGj3tNHpETWXBUveYj0CmMD/rLPpEUUFTOoEh7e6DR
A5gPMigTva8H3w0R7HekozlMAC/E0wa/SjKklYNa6b/hvTybHnURB3PmMhoFfQgrk1i127XF8ZhO
DDP4TO/uBOpF69eH4EHPZwP4t0YfE8GugKAYoVAHRkOC/vsB9cdyjzOBTUhxZ8bp4ChGuNnCCdz7
lu6W3skfk+u4dJYRwVRFLMnFoRLbv8+D8Lgh8/Kmns3kd3Q7orqc0TQF7NTr4K5Q+L/KlrHrMHOl
xkR4l1eas6TJX4XYZe1J1COuoyGdhYx6g4e6snZjSVq/bSmdyEv9l7qTUd5bWI5xPU2/Z+RJ4kSj
kleikhAM3NDbNFCNycGI/cggGPbJk+LSl8tzHIrVM1/GO4uhr5OAQ1aq7CtjufPrMNRWh5MzmZyf
VxufTlFnRw+/aZAwVaRASh+CQh7kfiZ6PvmKUtEL1LLChzH8D/CS3VBxN+bpDuG0WZH9oEjeCTXS
xxGU51DhOCZ4ja1NctlHXsnFuGDm6XwM6aljeYdhsooc2khz3JIUOIphuCBUXyLXupgcjblA6BbA
K+KMcIXi7ZA6g5JDorSFfqQCmt0L07PxEvTpSmtu10Isw5lVViETPv8yTzbfQsgE1+qbKDPQX+63
+ZXHNnyiLypjQtuMdMLgXT2TB3WjXRupq8Dc5QUenO8MdejjYYuYLIo3BA9z8Je+xGhqE41G5Qog
f24d5iqvMexMhMYbU1LZjvGGznZrJiGiODy8sc+2fAgtNv9tsbVbCgEONMU3nSCBjeUEA9zl3onq
JlldUzgvT4j6S7CxcpKTuxbbCks3VzwdkmT29juLunRJuG0ebJCiXoJ14Z4/sgok6m+1j2JsKVYY
c0/ggdNbeR7sBTI8KCVw2Du3g5ZK4idZjX+LwZjt1RCwZ3RDKsk1q8QFVlXRMCwRxKt75Gd1lquu
VeLEmD/hkJGSaloWn9RtdLrYeoIXA3pyQ9zzV++0BzgvPYir2eyHGmHdL16VnpVg3N1BPM3avYQP
UGKq+857bF/2DZ56IL6JjF/RvBAWj4epW/32UbkYP2m5GyK7a9a8XqmsW6iNVL41hM8hoy/ZNjwU
NRWkjuA7jS8GfvQRqxAzFhFUWXH3R1hNwe8Dwr4X2awYsXnnCbn1QO/XduGUAEkXDAH08QJ/nnaC
iX/cVNnm35EtGITQDqds6GX/qgkO5xX7ecKhPDm9pXyl45ZbP5vgkMQ63XDP6itVbsuSBVgzgG1B
CG5Bm3J0FCnfO+S+wMMiYMpTzLa0f/aIChOvNJXtnd2u9kR0cklU1m0z7euxKaJrV56hEAeuZBmG
iP0oYOK49/9amJ9QAy3qBETmTHLH7o3J+Nz04DgTnfAi9pY2G39nsnJuTUJaAzsK7eq0NhVDLAf1
ApM7jsAJGGAD1HdvJcyL5ZCPHiNDF7v1elugLS2OzGeW5fEa+rF3Sllp5bLUzMoBH3N6FlDnyv5h
cwxmInSEpAyfcJkzViT0po02IxhFjsqMvnNHFIP8rIotHF/XJKwB+qnyLcHwe3nMX2YxdhM5zjXj
VSsO+TsWOYUQiiv/C3kLDJtvevCEkB56EWe5Fs3Jtl4bYFyD1jJwoVeAuyGtwNDkH68n8M9mMxbT
/O7g6MtAAPEDyCafAziMOuOkNsqZpm8VNvgrg1WpCVBI1N0+DtSRyoSZntHq0+qdOl9Yy8OQ9JLO
264f2Hp/zNDp19WAA7TzSEwkDvDckX/TKSAFuUORkQRNXNRk+NGfsuAMYvzhIOMkMvbVWwi84Q7w
DMsXnPB9ZWzMvWGkolHFVbxwxEO244XtZKIyTbtE+TXdmJFstI8OwxWtQh8aSMj+dUi87U7wj7Yt
EljpQg/7xaCNtc0sxKfI5zCTjjs5HsWthf97ni8ujl1TfZKpzhyppzWw3Fq6SJcYaVeS3CFYw1wK
O3hcSc94lJsLraDntKozF1oPy6NOPqG4eb770eoCt+Xu9CUnBji02Ot0Axmwh5SpDRmAtB3jmcw+
cxXC4ARzPnchP+4tMxtzdb+stlh877wQ+aPYjfLeFWUjEpGNbapN3J/pNChVM0zelMTrp+58wzhL
tgoPNI+9SXR9svocJyMhpWF5fKLcKgleEMKDmCdZfGE7/Z0OTF6APxsOujCMf/0T1jOJnuWbdVm5
qLSiwYPNywNqnQ6X9MHwBXz5Ikoa/IzT6aurgY1tZgjMy2ziYje2R7qvS0gUcSXHccfpbpJ+D7pW
yXr8RiNyTqxD2ej5znW8dZuaW/qepKcgk4MBLplMpvwsJadsitbmBj8u+XUKoYpCR0vQ4CDDekfM
kv4klNcV0Xr0Sd4bK0ANJMPbTxAnu+D8l2P0waTEnC2Sxxtc7BrWcqjRpuqZ21Olqq4gPRvaJZt0
CO9sS4x4EdV0fAkeQzEmf/DMrPpxcrQXROj7N743d/XPYJLb9+S67oOBpGDaviEU3+ijsti6V/wl
BjxFpHJnGrPh/7dUvawQTzTuyYTtIuXuQrOQ6GLoBKmF9uP+Njlca7UNKZTrUZbvVJ7tkXrFXvfo
DyOBQxkdbhUIkKymkUzb+Uax93wsaoM+eFE82ujyu5RdEtgtojMy9cOgRho7Sm/8vXjuFwP81RMh
1ZQWAtNOmR8JmOGTouczcDztQp6C/j6JpluxXpbEGH2Jn+a/IwToAEkuHmnyL+P2eeBzQcIfs7do
CpFdwikw/g8kiZwKtydFHoo0LZf8zTZHSKm/48dTDYmgtho2O2pTyXOUFjRN24eeHQzS40dvKX+z
jDyEa1o+GAh3a9uC+IBBxXsNRajWbHIBiS+n7YK5j7lcvrhatnGwHrdThzOrRPjkEM8QE/i8gz76
utddV0samGuuctm7BT2qxp0lWQPSaT4g4FmGAFkmV0xdnj29ufFtXsfIxIKDrHukuADwtdOv6Ny8
xisUPTHkb7P94ub12mgHnvzrxRYaMcbmohkgbNx0JgcKod+ivdVpdiUwm43QAKZF9pmo7kQzO/el
CV92q0pAROeje0xHBqn969g3u8nXsTyc3ZFuiMJIi284olNTlZSciwdmz+uw6KSoEi8XvUTuxRDB
+PlY2I0hYS5SVrwBmuvrmWgbZhklru44yFWf/zExn8DKovCi4ZGGmAMOQmx2x5kGcUkUzk4mkQcy
TywyxfgfBbgiMgr4OI0Vpdr+1vRc7G7EjM1dUFn6KHaff9i/Ymye1OEfeao8FyGsOpdxmRgiLpt4
3mqtfJZ2KF4sXcTL0wL1uJ6zHamLM+tlsZZgUmBkiD0eaPkUtk4/pGg5MjJNtL1YehSApUErmC3a
QFtSnWR5AnNeiCKOobuha5bK3fIdCzfmziV2rKqLiaS6OAATUOCj4NsKNPkR/5M1kBtUhWANjW1J
mPb/6vTU/+njcP+Z8I7NDjFLiSaQDVXkTBPhDphIy1gXL5BeYJB2hx580OiGXMuY4InXlo+O9Vp2
5e94dCeGplXMYIJ3CEPDIHljhga7+1b2pHSnRozyUmKYn5Cl5xCrPfOqW3LMbO2oUGnXXXOZQQuG
RHQglLMR2Q+Zn/kcu0pUArfyAJ+xQev6NY6UKmWfJY0f1ehbWMhxaLhDX10T4IABPMing6JKhjvA
MbGlEY1Gv6pCb9hhrv/fiX1pr3+YCCeOJFvIkK+LzzeSX8JM5Mh+zALsb5dktrbgakSXeFhK4aDA
nlzDA+PYsTNPNiz8ro9CWUVsajIxqFRUiX2PAtx/GbkBsQjlc01DHN/br2sHTTzPh/QG57LxT/xm
9iVvCBQ9H94o9Iqeu07yxm4p7lWBY6ks27p0Z458Chxg5OZbptxCfOlbbqXiVtKubkjHqz5eF3Jd
BnDMvMk1S9ymm7YEi4Ddv9WJO8QVTzOOaAmnxreKq6B/GjoNKwBpaibGt2kmyBTNZ8/JUJYxEdw7
fWJXKBt8mBM+mA2UuJee/19n9Cpc/NlFtzENMoMFWBM6AE246GwXyAwOptYzeT38v3E8fYBkppBI
ODz45GFThR0mq+1A9s0HLQEySKyg+nt9CBSUnC1aEAZVxQ1sOGdefdShRVg051FZ/ExLtlB4uda6
JlwXtazVQdrMEqqsZG+jh9vFkORzzZBLhSz897R2vVIkFgEBq1ph+MpGQX8xfMHgRu32QdCqDrHm
gbvVRiDzSOaQY7bWRrjeeMQ3ldexKn316UHHGNcM7Qmb8K5JVuDWKbP+s0L+Tpk/o5nXXkyj/19H
Beqv6HYooIzoRxJSGhYhA2+KvOpM+m3M5ijstm5+Wlyo8naGjpTGxTLpqD2M/zEsquhrq1Xw/yqI
34DZmve2XcBQH8BdDRR12WCQaPZ/+g0sCBpYMsa/SMHl4QbqLkSbuqCg5eS/CZhRz6PBxEK/rkwU
aAtbl2igDK2aNCV+r9TUzbALIFRB7ej+b09kwGunA0NW770aFkJs/huRa6+qSzxkDykOyzXKctov
enPAabk4UT3vJuTtOSFaMETz49Je5Z13S1QHs2deHbOkV/ER8lx+4hsy/PR5LToFRxrvNtmAbpWl
l0KJhSGBG51UZSLGetZ+kpxbEGCf0J6D/BJ9p3zQO6WatysJrbzwg5Auasgpdv2mDpjyb+xvcspU
hGWlViozDFsHB7LEjWWSEpwrhy7aBZNNVR0Vi1Za8beHe/eEdEGXd1jzAV0uYoxckfOtJVkPrHR1
mgzEDNHw3934fvQQzbU/Jp/1+dVUHufHbfPUvJZjOAE7R0eHGi+2PlTxNilLmpAjSOJ2y4ksTrS2
b1FLaqlJ0q1hCYnc6OkbJ7+Sd5nRBfG/kSGX5skFkrJWFPKup+FVTpfGuytrkt81fccQL86KJIFx
OdhVtHHUIQFjINNstpUA4BDBfffh96Ki7eG0jFQ0/Lsx3toHTvwOyO0Dj6rWIPzcxtb/zr9qbW5E
dJuF5+MMpUXwQlWR5Uj3mcaQvqj1OIxxjNMf84pTDqTqfOaNesKxbeFqxRsQqxkDcUbl8l5yZLd5
UmewJmi/v1ClP7oRgERt0xnugm33Y/IdwnRioIIVHB+roEf2LeCIN8YwHVLM71bzsu0oXfuURDro
QPjwAqE3qY/9GyawfgqgSc3QOvDbEAJ36tIEsHOHAw8mTbCOr122yH4Y1VGx6M9FjQ6Q2rbZGFPW
cZ2X9JcXBS/cFX9LNZYqtW/Sm4nwtxl76T7zvUXP5siTpHBOwiMUzwjIhf88EX4Wi0SJyJc1m0tp
rqwsqMP9u3W8cTkmEQwVIACFUbN+gfE/V6V6NK8Xxni2JcVtNDLiR5d3LgJOwdirdq9X9L4OOXCc
0JSHnbvABLVLM+cFr6S26mmR79geAaqvVnXykSBDRYQApuqczNsRr/JWFh0ZDdTY0PxO8wNHQAk8
vRvvykRNGabGarXG2dMtTDSmLiZzEKoBNn9Cd07hNs1vtvMpYwnc+04qEnHuyy2UopQq1i46OaTg
7umNd1kf4vcJ9HMP69VDkCWuSsttTNn2KwY5CkquN37qnw97xN02L4qpA/0mumq6hcjf3MTwfEkd
Fvg91xyxzyweaVmFWn4pQDx+5etaRdZGxI1eFTvnsD5epeyWWhTG+ym5HNK0w32NKNc6h7w9RtRM
PPliv2zDOkRg1Q40YbLjlm7Y0OjICX/PomjfmjJ/CM/pNvEhx5LOHQAdFfoCwQFY8gE50etQ4mzx
RfrSIJRBRUQQOUhfWBKMqBPiT86VGjF+zEBP5Dw3C4QX+42QOa/tUGbF24bHfx/GZU4crhW2crpB
ignMlbBbO1XCqD0IrGSVS03TAmHdlbC+/wt+iQqR9l0OSn7wCe/NF5ez33cm/3gjZOIpgT/sOa/E
NAWbl3uMHQicRYSuzGr0oyVNcYWi/jfdma7Je2CI9yTyla7CQT7ylcSPyPQQk7VJJvOwWfm7kHyl
1G4x/3IujdQq8l0sQO736OnPqpJ+O3hI6D9gU5CdQhsCa7m5D+s4kQoVQXYroWylzDmbMQQCAlVG
9EDoisz6g3eg4uSLFeGyAPXEgWNgD5KC0c7HzHZaGOxYlDaKPJZiOtdLGzvF5kqzQpoKl2BEqNMo
HaWpw0kJ61dO1MxAVMp88Vty8YhMQJJMFPw0ImZr/PVDC4GzhZxhtVoffTR+xtWpma5Fy08NF9nO
V2bxincEeDOm2s3FwNBnPZev86LRZhMJyNK7gRbzA6vGXzoOi89yR6My1TVWqipRaZJHhrjSTNyA
LWuDcrwZn8QZ9Jko9/exh3xWUDob+nAKsfwlubMbraQvYvuWdvEHxe/MTm795mIWdbDMWBY7sA1+
XRxr+CUIoLxqgUTlqhqn0avUUAdZ5HvGyIX8V7Tw48+Y9oB/4Ql+OaT9Uu9lV0V+D5XXC84GUTVN
urYFEb9jSPbOFkRGKK5VcEketq+OU/xPWaxj0lGwxoO5QhdV5YZpxa4pLkmncPLSmvinQX4cQiBz
bPEgw/1yYYPmlzu86+/v8XC2vJKLQNmuCmg6+rmq8416Comz5mT+9pWFXs/yA5V7FPhSlJX0O5d5
QX0UGQ6PjPKkT49krhJtgQvLQsAPFdtPBNwlSN2Kfv0r5mqI5pnxHps4NOI33VDL4023Yhd8GurI
YEFeZxLKwtyn0jICeEkKlEVuhJdU7RrI5FUucVxJiKlS+kFjxae92HRiZTskdzz5PgvVKsgo0FLv
GL67KCUVoTihc4lbYVnoP2DqN+EBf74rvKWpF97WZaM0Yf/llmdEf3smFWJ8CXzjN+EPmgDv0Cei
A/0c9VHX0yv+dFrkEe1gZ68ZGcdmbykeoHM8gWqpVqkAnyjpzbqUjgUtoJBkBSFk9cjSTf1e83n5
RCIQgNhR+S0ZEGTlsdqLYPXgyBV7b5uN8LQAxSt7dvyzx1aeHB6tEdAJLEhqIxyF490VWCxSh4Bv
s+X9hNq1FysmZkir9j7eIu2qCZLt8oBikxg5xnAgoi0szgy20kjgZCCl791VGP+PiJ22FdQlJ748
lWJQ8f9D+AJrFjEELqInn9kFBIAtZfIyvqRub/w4cA7WSlnRPqTWrXnRUynoNYVWOsOWTywhNdqQ
llTX0iJmSfJYrwiSObp5tRZsjLLeRuZttivgzrZabrLSVadyqosXT6G85/hEA1kn9njgmQPpEz63
mRHFhA//ulGSjgiUSVy2A/9toYmZQUnyVEosZTySlqR0cAgYZAkg6djugXPV9X7AvbTo/iRQ1fFd
OeWHJm9m2ORaRT+E78m5J6gsV9Q4fS/kQJzVT6AQHB4LyCWgzS2xKE9lXfnPpyru7ePE8jA4Aapd
sJYb2IHLwv+RenyZLEz0xN8xHdRfX4ZaDSE1azft0BJbBwI/hNraLdlW7VxTiFkOBSQLA5m58mOA
1KZVsZtG9zXq39pzRAPjD2y90zVsH7uBb+5pQ7hvlsRFWmMJuWHLt2PbEejpPOq4pEb+tHAN549J
+1HMV8K4ey16LIsWbm0HhCb2V3mlpgcVBDtYh75CBsTWsXepywMWrLAQSK2RULqN6Fw4yrRcS4y4
n54mspINqZynOLvEICWgzxTkDhcrRr+CxS63EuOSWEfZTeG4G0L6QXqdleKXV/08LI3B0P7ldMIe
Cc3PQ9Qzxpb4uwYULk9SVerFDQlJaMp6STbXBL1og6Fg6HyGZEg4e9ynzcoCYumP+n/MgQVxctMC
R0Izal/wD2yolDKkqp0LKfE2KP+3yDbHl8OKAcFBuJxRPOGcMId6/iwsyz2PWl38sk1Fq9pobv7/
7pdJ3gtafwfL20DDrGtjgUr/9f/aHpUD/wPdzPuZU5Wc4gUVbbVlDDiIZC7ztvC52tN0ae/NetF0
Qivb58yreSpQsmaxmisszaWj3z9pGtnnmIBJhW446UML6UeawwxoYK8Xqi6O4dBVuAf6s2QAIA+c
zefs8UBKlmMQJ25I7mOrWUg7glZxWO2OV/otiF7A3QQPtkNOfdA2BhWz+phomnCPU6zuYC0jrwXi
GHUK1Bgg8S4tuvkPvBge5Q60vAzqMzVNkIu1vV/AChokIA8ZsyEsumQDd2MsNo8vy06JGzyWw99w
y/u1YDhzItIlt0BQrXPJgayIZ+Uf6JnlJtW4mCREeYX/eFQTZg1a/fjMcvXoe8Dopf+BXkzg2NpI
oHspUHVjLR9OCZgj6xxhW2CkkZHH7QAuPbp93Iy7xnLod+YV/+to1mCbbCkQNeg+TwsmCddawOan
bpBxdM/IwyI6bH+3JnJkIaMouCbmEzVLx/xS2ILeqSVPygP2TCVVxbiWxlDnxAzjqGCZAN4zMrUd
CM2WrVDMPJyMuDoVKl+3kK9MoFCiWM5G48go77rR784y1lHT1GBmbu56jmF4AO7AKs4nCBVTd/tr
E/WyAuX3gKQE1KvaP7oMHtNW7HtP/BY055LVEbyItkji/n/A+yE0KY2MyjG4wSIMj6vJQl8Ggqxu
Wdk5rvwBEujJc+AgjHvSGYopGw5wIlCXnzis+vj0aEsImYuNb1sKdMlDeiaRoO9CJM4eVnY1tiug
K7B0Udp81VXsz5gBr/LnGM4Gtq1ft6ujgQL/JVEaEtVki3GZUTCbiE7vDlFpVt3hmwXIqzdrnEbN
tlHVKLN/AlV6QZQVCwXGeCOFVeR+MUzYl9zyc7a8qRQD70Fl/Y02joLp0Y8ddwuGk/zqu/Rr3Nab
0grO2rf0wXfjkHbaNmqQ0YsjSwQU7jmqEg++Mtcm4bCei3Q4VBy/Nb5GJWs9Xjj3Js2Jqr+1L8Cg
0/RNO3iPTs1aKBTj7tS9bWOPfSS8OJDZrCx5oXw6CeH4M0YZaet5yrl1UmqNEe8t98FWSVaJNv6p
ldZu5XwoPYtjm2iI2+Z6eL5o3myQ0RHKfHhP34lmcotkZsBswDc0qCiA36WUcKED8WbMigfQpEj1
E4HtoC2pQNj0jIrz/yPh3qXO6ek8G21KHKbVVgCgIh58IW0LDHd1xZBWe/zsuX7sqpUHSB87rTkB
wCvZoWnd+RWt/knjpT2F/VgYN+QGB8KnRMG5SBsSBoGdzmzoYaTQIOCT+si/i8zW3Wf/95qIF4Yo
OMrNuGLgV8bd2oObxqpq+5rnrUQQP5niSyK72NZ+xBUDEDTTieVHlsBa2nAaZSMyJyUXPchD3dP2
T5s+CrsZHXmZPKuSFuMzXkzXVoILaqP8IEoHbBrgk0L8YpyPxKwkgrjcRvzB04HAoTuVtIyeFl1D
yOLld3VxGA7l2S+Z/jyAzMUBRZzUB4DGT07JpcRMwIyPROjlCaD4VoKQ9+KfOhM5WPyGrGL2KdLO
CVKkbZqbGPPSCr4vopR16IhcYeV7Z+POCFZUCkDFfK+07GqSFvX9U7VaBSqkVwAMq/d0z1gZuNbo
FY2SMqxrV8eHFYue6az1ig8kh1OjkzDrOmhEPSu9osono24YzQg1rJ2vDeu74vc4qNNUBkJ+0N5V
X4/Irw2ThVNV9ZRAZFvkK+gsb+mQm/0utJ2Cm5HUSldr0R/LZz4nTN2GPGcIPXstd65qncmn42D2
gPutaiVx42d0Hmkn9rxzcF5OYcslIQKl9L8315yPRtcrEP9aYgrnAYLcncgCaAgkb08nCIbeOhsv
p++9b6imlEim9iRffPuq3mwERqtrIlVuNf5eQmroRXeNC4oDZjH/E6vGCNhEgKWNewFdR4UoBmbJ
neHxh6YaLrscqneOrA/HoTKyZnOvCly0bSj30DBl7oV8jE7hXWt+HVcYSdbZKPO22ZoPbJWsg/j2
VUC8U2teKbqJLuG389vmQAHcB1jjtV8tTfPNREZlVA9E42vu18QInYcDylVdMDTiUFl68Do2TsWL
E8r0o9SvbYttWDeccPzEMXTG2R3zoLNmfVpKSbZVqQyuVwroOu65CRNGuU3uv6PCWEZBefwidwA4
hEhQxoA7bHrMbN+CNx8dUyLa+wfqMyXyyk8J7HNIZIHbhPYlnIQFEnoLnY3z3mZpig8uvy5p1p4R
VtNQWHRvNiHMwMti3fGOnQcX9qYDm0dPIXLb1J/qCy/zUIKgt/oPrCDP/6px7xkOZwDAgJxPvRp1
WXFZF2HvL160cG1uvdaU2l5qkUaqQPJrxVmR5jdTH6bu4/vK0a1xF1fAaa3o0zxxDb1y/nxhymYf
dHFCiOaJhMNvo0CzV6zBOENvv47JE9PYdrg21X9hYnPuXZiQ1zS/K5CpGcf6yefsgmZ9NREY+xEK
dhp9PdzoLktI5AJ48CRq/CbsXQEazT+TV77lYEfTFbYZuN6s/+OvtDJ/6i/XlsCRMQsbvB02KON6
9hl7hy3P4gWI+VCHnZ6TCJRP3Ul0uzPXOtbVstYwCiz38FSUIAuggIJIzTIebO/q42chv9hrQBC2
alGwFJd36sheTRQPdDwvwnhDt50Py9eXx/2T50grnOM/amSDFl89kjJ4zfnReUC1SO7w20Fr2xl3
2iBn+AKaU+98SAtf+IpDRaifdqIESiEwTSLRt6XcRcI+7YbYa0+JOo89JwN9Rd/Gaj97PwKWsYE9
cxA6Jg/UBInWoC+8qsQrrQ0T6kBmJSXNyFbI2R+Ts+C+6zz+iAxDBWn26kL454HiOj52vSshXGwv
4Kg1awFFpoUTzggmfDUkjLGooIWg3TGZBCawv6bhbPkHd2Amn6Cc57T3qol9MX1pWNSNnerv+Rfp
FcXbocsuJGUxIdrFVEHgERMoMMK/imFTxm0aKePXcz/PpaezbYiL0kC1/Sau2Xejem9bGrjmg5iE
jxbr5mX0v17nvp4/5kWlOwThLR78bJZkMIEJxiO6F1B1vXauFvw7UOIDmEdRV4oqc6nbIZ4KwIwh
CiUmTzeWYUuckpFkqua/Ad5bvrnC98qt25/rlyhTmvNogCPXypDiVGuTJOmT4w1SU5wgewwDcHRl
On2DDSZ64blAB4XLWOrijSQlnZG9nAT+X1T6oj+qKGLL79VEsB5PPWj9TVkr/vselsLsTitoPvBG
mUnG/vRY5LsfrN+8hRO91onzv+Q/6T7dtwMIVrsMDHit3lNIJnJbXVO7c1HA/AqLBJFpIlQTbbkJ
OJ4IuG3gq5Yh5esB49a1jtHMUGwAqWJY3hYgBuxihDmqqxiixYYbrgyHCEVwN9B7ISonhozivDUX
6bXriMOm55MUwwhbqN7bHBsqPfEupgGOSMSIxOWdnAj4SbSMIUnVCMEedmRc/gcTLY8iw0303SQ2
8fm8MJURAyfOPznN8L69NRtkOWHTVmmkUSeHSCYZS1buwON2J7CSZyyZU35ehIqZsJUe8AIqr/bL
avUWEMTbs9S4uhNJGNzwqtyWMuPXKXbICRRhRYRTgKPWgQNffqaoMR2OLOh64HFvNsmIYafbrFzV
EJjpp0zn6w+SvsAucs1Dbg366mEAHjo56cpLWtCxOhGqk11r6iEdsqnJRqsfeMUQn6a3S2bH+UVK
gEXFdlMD/dOHw9JUTYF9ytM7/9rcSHo6CUJxEvOgq+ki3dvgBKYnq7pn3sqOKPsWSRPtU68gjC1w
jsLgavr/pyVdfHGv97M/b+gyoUU8Fgxj+x9o4mO1K24UlhUSIXRWLlUkHP20mlGctD/pvbMtQ+3/
YlYs1mHXA+WerCFylxfmHcJDZdYy3Vm8LCkRqys6rK4VF/dAEbYTIzxZNrcbY6arWVE69YKXZvW0
WEu+CRKVrYeNS4rJp5KYwrejKS89kmwIGCpAvXHP6Sq12HuAN+kYmKxqsJjpG8azboBvX0f+AhJJ
qpeDsRmqsXg9wZe3VCT85MKR7TeVhl6FV4cP1JEAyC2X6xLKleuH4pDBuRo8pPkb0V5U20vmLUCF
E0sUupcQU04J6YmtOeFdEXbrncCYHjwBKKZ0FiNydZkGDnytJjjpmYZjCOqaKq6eGkZgej/6u3jC
e9ZH3DXxpzmuvopmuQRinteCPHVW/gYsBqgPqbahxq0mt2SC6+LUOjWDkhyC6BywCXj/EifUVshu
LXsGg9Y1lzf4sjrTWK7dDh2QDQ86F4Y2T/8/MaZCvZn/5F3fJW1nnlIjc3mzHUlXNUmNGvWsQhWy
gSNb1xoS5EZdhd6yn4B+Zm2EgbnOt/0PGumJBzIhlm7BAgep18vFpHNCS73UHzq78bnEh0fFDsMe
Xm7bltalX1V/Egxhz0q7d+Aq6jmsgZDRb9p97HRf5bjZuErmAMpNU9QGwF8ThBV32AGwDdN2Oong
DsKj1sYDV0vPnSlSklEccYY5pmb0R0qO3Mhy6vsmTFXXcxH5OT7RSYSwI8mILQb/tVSB5zbsHK2O
GzbY5LSTewUm4RdmRJvGUEPnwlhF6A67mnDdarEgTnLWyy8b646rZRBvp22X9yYvE1QC9vWzXCxp
Z0QuY77sDim8IL1xoZmq41L8OfMdccprHW3L6y4BzTmSsxu0SzCtfMLJ94KuZc5ihDL9zlDkO46u
wbTgrMS0Pq81/oMlFaRooYaqZRDHk4h4KQmTnOjH5JBXbZUXPsIlts9cFv81mZB2V0f+P8Z/zX9W
0XMqRKTA6M0br3WIR8mF0gVLZLZdJKhXziHu/5APe8AgVQMQczH6MB5y94nWFobDazEF3LYfvZ2W
iSawdg/QuO7ACARWRbERtFVkJ5FpLpOUL6I5NlXSw1CsrK5Q5yZpEs65tn9cwahlFagqJpporI5w
aHiMODMKD0T+IL8aHm12crHAYng0cMFTNPC7SEISaA5VIixZ9xTfJuddh789Cy57b7fTqi/N23ma
AeNGv67psfZeV1fyLGTI6643+USqNyV+fHr80UDZ9v/aXrwQhr7LuD62E0sHoroCdWwYZ5U1wKsv
x/8oUszanVhqtWhOTPjcSWGe0NfQRmj7FJpwZuSMyPFtG9hpSDnBh5di3CvzGJ+YhC6HixhkbfsU
IXBXinAnwvvknFiRGj4KSkcG8T6PbWi85SxRFu2YlMqvRc+AXA0Jc0eKh/4xCU5VWO1XcVF+mnvq
gOp5o2ClyU5o50pFwsfHHR2CSQOHGFAD/rkzMbUYjw1vL7Ix4GyI9NeetlSgDDSSGz9JkqwsQuKN
tXbio1/7ES5WySBLJRuNUjjfD2A0+WG8+GP1M4kXrO5xLp+H/Hfdvg/tXojOlnTurnOE981Alwaz
UlE4gX9wk92UYpWenoFqjXYmOIS1Tyluto5ps4MPR2MnpNC4wEmtgV84FGwgItHWMk/6yJm671oN
wNl5PcUpBTgO+WQDOEzLtSq5xwsVjm4AQr2NmRCIMG2Lf3ZrSXIesVlXEfC2Ri3yPIKaqNdTik9u
Lmh44yfSbGP1/XszUSG+5PuPhqGCzZ3aOLNMJ5Q17uEFGeQ6I0JYI0vuQQsDSQUvOGUbbLsd+zAg
/gidy2NQ6yaYOrnsPwIuERNgw8CQBpd9cAyaSCRqpUG6fi5XbnkAWDIOlQ6R2jCv+6OHQ5Uy8eGU
jrp3MYpn9cCuIGz0RsLbvv+5LVAUkWQ+4szy2Wj3ShLUs3/SnQ5yyZMtQs44KxU6LhTkyaNIXWxD
Vis+dz2frsohkvnzJXKbWrCBgbaE1XEhyk7Pry/B5JDKjHtjO6FHaSQ8yEsjycN4tIESj6y8p6qg
30EPKXxzU49NdhDufCBvFKIOHRDFeMk72QfAqoRtbhBKzWrNG+mSIzu5NaXa18zjmUvojGZXTd+3
qJBFXbtGbyzYKh1m44nH7r7RMJZHk9T+vJQNbq0nXpEyjF35zTzaxzLjq8ee9S0/dUz3WYFyiSC4
o8rySS8OWgOdhGp4exQUCe5yKLSpe4Td4AFvtEtnUXwFiLCtV+L0XXfRO/IksH8cKMmHcXbIIzkv
D8qtOFE7D/iE1d4QCDw6rEFJlPG5z5SoatFUWyTlSqqKVPt2AOb+49WoNPHP73OWp1yYpQan9k08
xE7jkPPU3uiVqzIfdjJMK0tlZl2lZdadEH4Svl/Dq0uXZm/A1q7no+7VXdABPYvXsu15rMiDNA8z
7lr8u05jSbgdEY2U9GzHqujotH6wv1oo/rZOozIMU3sT8vsloU6CpPK08lXV4bXEol4x8AFLlAQo
rrsaxAHpFeYQSI92mkChPYiakpIyET436Gxg0Ca71GumV/Fe4sM7lro8r5Q0yXap8LQ5ZBPVTXh/
0GL6OVfYqZbGEHtqctQlT6h3lpk6Nzf+g30rZl+8tGkcK6QtS74ccoowBnOrVrwWHDSOPahEAra3
V/3muvTtOD6Por3AsPGnKsSlsbpOW3NTKMyy1BIRIH0a2zAIh8P798rlawA8kKQmw2H7AKCBgwpR
RqwrL40QYBI9ynDuIO1+Lzd+4o/TZ/qE0LM1QOgBz8IWDDmX/Of6QCx286QZIYPR67fUWyLA7jqb
5xyl1lGBZ20cNnJZaHjZIrg2TEL9HIh/pFNAA5/PZMkmkO6QK+QuYgwcjesbaKW75Q9ugvwOWUC9
APHrUehdAN/7Wc0R8cdIKXD9YBZ42AwtRHYXNvwIsqIlVFW8HJSwkq5cM+frXMhVqoCabA4aNS5P
YW4H0PiPiopvB1Cht8qsMh9+rDL0iyDzUJwx5lswMltXv/O/FHofctKjTz0N71H8o9mwX81UY6dl
vDBDf4hT6uDRxy65/JvxjMUZmGWb1rK0+nR0X+PkSVnzZRugNqSXcSkOINmBJi887HHSqjI429VH
oemeJjtb+KP+QB1nZn27TQXSN5qKXnwclMRupalYhg9sIf5eXtwldXrZImvokTpGgq7UBwCKq75c
ZmLUZ5oi3bnFfZxDTzh3+RfCU5g/HwIzAG3dGWxg38k1LACSEgnWaX24RURBMAxziFuDgtkCRYqk
Kagf/4+KZRL+wQFOK6F/J6xhFm6eFi/Fq1HDQoCzRHKfDAvcEUD74F7nm9uDu+SMJWERgLaPJZGF
G1wRKf7tCgb6hPP9CUlBoQRtoopV++7mabYwK8nNuvnA5s65B9xL572NTTiVwN31cDDuKWd/aqoQ
2+Ruyl8NREKv7VK4r1v42XSJxFfPrKLzmx/tcrO97qLOwaDrUL5avZSBtHEyjh2Z6JaRoNvLvDfZ
6b4vXUwRrkaQo27R5NfkFbbTn5kNgqM0pdsD0OjHaGwIuxHtJsZ/alSnUzPAGLqHnwWaj8UKPo+F
EOWgHectxvlZcaXp0qZVy1uxP5jp/+qy2MRlSQ0BjFo2jTgMuQHgwMffjl4MibzWYXYj6ymhnu2h
dzZWjA6UkIEUzjukjNwxRPxgQxXzJxnpVeD4cZ/yaLF+G9imyGww/Dg4uHg6RBP7U+AEvs1w1T4h
X3vB8f0IFxfq2MQ05cyBkM8aHUSX+QZjVZgx7yz6E5ZBJc7wPixwLhO1auQ6X1NN/KCT3pVM0o0I
5Zd8ABv+qjHewFItRCvA0l6HHV+47V7tSoCmTNeadXd4sFwgq1/DFV0a1g7vQXGUT8pEADZABDNJ
HAUZl6lCIVFErCYL22cx3x1meh1nZsYwRcPOjEE8w7ZKfqx31MoxG7nptGkmLYckKinbZZWH2ClT
ftnZDGxUzyXPJO89sG72C6F0srQfT7GYdjCbd7AbmrbHzmK/J1r+GFO8VjoKHkCYmZlDeXMPZBcy
H94Uk9riC70YafwsBADUBuT5BXlHudAnMBbXGirm6W5yVwqv/y6zaoM8YriGCEyNotlmbq2B5zTp
lzaylkeav/v0H9deuEWjvWIv5vjINZqAmo3Xb/yfbAdU+Q7P1Ob2M2/+qr4MiYGRT/A/aZUmcNXB
3snFWIsLC/2Pvm4GPfJMHPlBzPk+JVKwdhmmn4R41rk4wsnEURJJfOzvaG/bfbm5r4vEwq5GNYdG
pUUXW3ly5mNkcqILeVjJE2J3CGk7vmNF6jufIKG9F4gOMr91RrVFuc6sHhRJ+lpGikb3pNZPC/hb
LTqqNEybOpmqaBacY58QuG/JmkNBcvzLL0+Haz/1dK4oNO/tqzZ6FWQYm98X5OmYl9nKVVoIJH96
utYFmPFbz7PeoHGGXD5h+GgtxHIKd7mNAVP2npQADTVxsIBUrgITA0ffH/LzyovqVs64H0o5lPHW
6dEynwtS2HgqKaxnLAF3mpK3Tlafp8is2khgBkJsQPRas3aSQzzOyX2aKRwNnGNWgdxWyTLH3uyI
douip9h3Ehwznl/NrSxfanZN2NMxneFDOMXLh/Kw0oyxRSRHRsN8zLWOCC2X0f8RNJ1N0ZSPk5fh
XtYH43E8neczmOGTzxFXnrlnxFaziS08k67Y2Jm5dB7bFe3BAUt01skQDfSaF/iko4FDsgYQS+uH
zY2YiH6uMq9DmpCRUotg4RASf+DeYj7Z0TIKCAABmJdjVSyJJOj7PHeNXviJddfgiAyj7cOLBYR4
2+vDhP8nS/Wu8vwUFuc5eYAPnNf36g9kQ3jSgekDLvYYLu8drkIuD3d+8Zf3Qi0SehlkGRXmVVNp
Zu5y73+q1DaMQp1C8NdEomkQrTCI2icZcpFUiJSazkgeJLiMCP+Cj1rMzoXNyrj9IR8lAy23Q9Pa
+ZQOp3RogGzfsG1ih2E8/h0NFVa7t3okilF2sPmkKtGTJBhCpjHrhwY+7mgU5haeWhsIcD6J/l/y
4yTupR+mm2jOcKN7382YuomxD9TBFT77V1Gg6BojFrIY5wMXzdyNTdPX4AG3qUAE5MvCU2L6oStA
IPFIK/A+2qPXcfYULZ+FVEk+ZuZEwtdzSjR3orgZO3rWHD2PEFyHoJmwWxwkzDTz3xZF/Q/+XV4z
2hn8wq50bZwQyPWNN2QRDvbvDoWrQvF9aET2Lq8YiFPNyKRxztk/zLsNsTG5PkeKXZVCCKklAUwj
50OGfOFU8SbQ3j15RclMFUVoMd9wWiWTXIEPm9JB3mfaJlDQkT/ZnNappHyttWlOMid8McA4SXMd
Awh+bZcMPrj7Lc7y8HyGuYi9q2Uh/b4vZgyfKk/TArJf3KpwdgqA3wiIzpnoHDG2YYiZB2GOWsnp
aZ62alAssbCjWR1pfCmtqs+ELxdh5PRzw56anbVpbRqlnZGkAPIxWE2lEqjI1JBw9mTifQUYENLZ
eu/0msLtbCAYf573KTnsrWNb/KGSNyoODPyYXF97YYDeylM5+ifrWWnEBqcM2qf+Ze337inNXdO/
Xj/U0f6LhmIc4Es4I3tFNLJ2gPSALlNRg3XQyYvQm2OduODDpwNKTzsusZewSF3Cj/x3mJgk/G7z
bs6H212HJmJnOD6c97j4Y2ZVpUo3twgOxUZEsBU3qjwxDHwKpuEEpe8c4p0i/F7UmWP+v4MkG5lB
hkJUNiDKR0fn7bUpC22ltNJF6KFQU3ToJDU2ikGjh8OgRElFIKy744cHxyVxUbh4dYrMpuLMUXFl
DJFlVLoizGg8t75yUhly+mzNaYt+UxBBjLXSrmXa1e41Fk/N4qQ+YWmBhyO5eWpH8bChtTLLaRBr
ZfjqsfLIBc+48PrIVj9zIbqb8cxlde/nDNiYhucXIiadDTbCYrHr3FNe1oNFbMHXVAJPqDpaOl8F
KopQ1wyppyAwzMz1D6d60QbxrrRonHRrlpF9Kj1rZWqPWwYqYSRIbb2ybrx77IijgeZEJmmH0qw/
QkejCLTLnsevaBL9ItOwyMGa/cDe22QwBAns103NxdYQ1ynhSB4E+x6/GZVKfvvxhpd+S+GW8/Ko
MGkmybqkq9do7pw08ZpExSceRuxnWMkChTREBgvzfKYN8Nzuiga6b/UOAOd6tF29S8ksyAP/x3lp
Xf0axKRqJ1t7rBefUhhbzlSkNlAPqdn0VvjNbRBCd8D9apqP8VIyU51S9Dw3spATQQ0gk4jqQmYV
3EsESroAcYlWKC4QUjhvQ1RXCWmpEO4chz4w+srzXtHxJFJgnFb54xS/jJnUohieed+lBWBlDPiL
GFB5jj3r6+l20h38khzwM29+f81o+72+scZ53s79JJWjx+uvmLR69+8nJ0WqSgiqKV56wBmWfYjp
/sXB6ptWQKsmSaTO2lNaaH3DRqV8PBbWcU6vtnaO9NZ3lKw8PCyAyP8ywTrO1Kn8MXC3JAPmBE6t
nVOnNF9A5u6h5yEnBF3gUOhcFhCZ9MRNK2ILUpXSoLIYzQ6ZAG6Lp+dM4u6qiPgVM5NhXGgXiLEZ
SArgOiBBp1u4PclTPDJd1Zn5fwIn/dQb1YjsoXDjdsqxI2dLsjZ0IJuzlIlRv8w7z5yX8weFmnGc
HlUi2EIvMSl54goneYxPFFgd2BhNeO2AZiWkl5NqAnfa1+3ddi4oC7GnCyQUC0MgAe9CxsbwG71H
aczL6fE1CwUWNN3rEOBhSuSEafn1q3w3kBbiD3bXES3KCLjDTCq6DFymkduqIbiQAWo8G1IswM9p
OjA9MdbepYrO98aWsc06JjkJp9xrcKy5HuwbqG+0WTNV8RHUK3MCGDfITKFyCbTwYJKUx4Sxi4Pb
t3elEbV2wD4DjFBKUBaP412tR7dseFZ6kRrcvKNLVscY1gTrV9QjDEav1n1ybmb+hFgc6vIEHC3T
HBpsoyQXJd1Xclzfjd7hsWAknb5JEnXvZn30jdnRieQ+F2gVecWMpsUtWyB8yAHJSW0Apxnfblc8
8IG7qAR0sJtwd0siAA+6OckMTuWZdwp0ezlQqROUgnuuTAmlkTnjqwSpLuDYrcgkb4zVTE+MDD6R
tpPoJ/r7zZImxlsSWqOTEjlNLH71pU1IchOEDvvpdkEinuQDBX47wk/UL8skv2VtbwNWp8xxoKMX
7mb5MZr+FBEpLvvm9BJJURf3BdfJPDSwUjjNJAvU04UeYcPq7MroRTfe8zdpN1A6Bn9MjGhQ5Yf9
qiyl0q9puBVxQRfCZNGPYuR8Cwex7aaBUbf5GSwuz1j2Qq9vHFeg2YZPlkWlVLHv3Iwhqj5oNPj/
IlJyKguj43idRdpwUvjE/fIeryLHemN2AQtH7ymtwkxWj7DkrIYrQxwcNtQYY7iKZ777zWH5FxpU
Ld2p5Al/OQ2773Y2jeye37C+2CXAk2t1saKYJCzQuYmQahSudWXEOgfnb1RcH6oZtys3Be2lQt/m
SsE26OyCM9JOGcVLpVPe2ZbwP7Hm0jsKPcw6tzXSdumXQ+SOTmfW5DES+7kpMIuGNt0vCVOKVqvE
6QTw0Gm+Cq51pAvt4BvavllQOeFwVeg9tsndM6/y7fbHRNelV516904zn3UT+yZHdfyIkSND99rq
xzvI6hsrynilvlrkcfBPom70377MUXbiG5SuD+3qNYyCW/YqdiOQ6373/DkpY7eERMR8scjqthRd
WdnuQ0rSCz5TxFrcq7tXu6DZdMr1NHjm1xf2SeRKzdbV1MoItbWC8cKnCPRu6YwMicsBul5AFBBR
4Sus67oaa4aGYbsB3rsjtqXGoEfsgItkECbgo4uW9DCOTrSFlHLb5U2k6hAmkBn7/CnAD4F4ak/+
V/C1kIWvtg0ID9fKqwO/0IdKgrFaJsFaDzpY/8pQiILMOwIZvxVf2Zd9yMvQjk/uT6okKEj58xPT
X8peIjiyL9Dc4LJdZMWbBDaZ8/cbtz/5aSKOV1Iej99h9k/lHkCQGdSkZN/UsQ8lKz8l3ofaT+yb
l7cs1IXh1h4X0NV3b/vSqg0qfBebRUuLujm47B3CI8NZBAohaQikgyTIvBbNuB/fI28a+A9rgwbv
KbGy+j5QAZrrVmwglUjMClUgadMsR4OcRZv9l2WKl+gZB+vqxkU+QDoFp+SXgiBhUHq9mGheBMEw
zHUJvlabCzTRsUVB4RvBEh4yj2GQYwR1hTQkk/UbbLlnDSQrhjChY7ahs3dq7jHw1jqWFzcqqTXU
3rGaWZ0qugRnyGs9ePyzfvNXT1FkjjN7wY9DaT0mAdywE3V+vlIM5e1Y97QaZQ1iwtcO23f08+sM
qTmR8aEcYRCoBDz7gGmwy5xrXFg3Se2ywWIch/i4SHB5m8eDENrm3mrfiNBK284y71ZiHKQeeyPE
38ytzhWa8ZGbKn9jKJJvmYkHee8+JgEY1YwHMfZFW8smS1cD1pqS0KMgykto+YOer347zVhrCvXX
OYer3NM59EEiQmR91FSjTIEmQvPSLH1+t7tNaDDSIU5YMyqC/tKekEZlIWI/5LHniCM1wQSme/8t
9skQFi4eCo4hZ4OtUZxA9T+pXfkeQcqP7vHb2V9ZAkiUPc5enTUtGeDKahpzVtLyz8NzTVxYni5H
BX+jaPOSvyB00hSOOJuUlwq5T40R+Kzfb15muofm0MoeQuuB9JDHTeZm1Bq26omw/h3DV84Y5jZB
1XyUOzWpd1urO66pE8ydb33E8Kt3dgJo1ce+4Eo6AlMncI8TRNid6E42/LKLI7RyzLFFaBYb1RaO
VhnoY/GuSDvnnXv4rhpWnIUh/DQn4QVErsfBiovhxxIkzt6klQSIJI37qF1Iqg4YfXd1RwJi8sjc
//5U5t1ysJE4TBIhAFZfuHFxnXEz2582F6od7+oVCdv1ph/zxIhe4LNX5IjGF7145q3TLZ1IqWus
IWjkIGN+ZTSGMsGq9tJrebf1oesnUv/Om8suB74mK1LQ+l0wgMwWQCTL6AxXPpgq9aifJ+Lk/Sun
8D9LvUV15F5GLz41A6Qlzqu5Vh+C70AaQDoqfxbk0BuaamDJ3M2/gSvwA4y3Gcj4TN/i5852JwTD
b9irDSQy4k+JOywbjOhF4t+wpKhF58G897qqvKk+PBgKOI5xAVH2YydUAW7UbDN8aDRp87u2FkpN
UwBJj7bzaSLjL1dz4cMuCO7iai3jnZjpNSVKHwXGu42c64Lmp6p9ie4NDDEvJy+NjifPJqciwH51
4I0DQbiOGzsbzIEsHL1GamjVXi2LacW+njqMAKNVU2Ggv46bnGPnUe2F9cH0yZKJDJ3Iez3A7ALO
tNEV7SnZzsvu8rD7FM07OAWg54qaLn7t0L7WFkI/wnmA2HN96sXCwD7rqUhYoxX4BYiK3fjeJbpo
LS39rw/i2GGvrqIe6zU72qtj7lj1IHB4QwPqRgjlfGiz05/7dlcOB9Msw+n6K7ERwHVXrZzzadux
YRKyN19o7h2N1LO32LD8W4gDAaZvnxxue3RMwXYvq6k4SRbu2RMh9WssOQ+IQLNy3vfHRf4fU+rT
tKOr5oHaDk/yfPLiSVd9npzQtRaZ/Yw2cXrKmJmwSq+UNYtY5XIg29/2rsJO4MzkbXbIbH1ue7yv
/hUKSD1uSgkf3htkAJrNRbHCBpf32shwfNbGQ1QQ1NV/dwODszagp1PcTPBcYURzuj9m+CwPT65R
dKnIYeWIzbA8gJvwEO4p6A6cmAHi0td6ZC+iBOfNtrByKOYEQH1coTF1XsbbJASFoY74ybFgS2zM
iBgs+0MWhccLI6Zl4ktOhOfJbTqqFfqowUwt7NV0PX3RrP8C3xp3i50JwLbgkEttWYR8UweZ9Rie
+KuHWlSqgNJAxJULXXF9tztkWzIBrNv0dtzY8/M1//dufdQlI17OboQQEzbpJumw8J23F6mqWkh/
PDL5zexPQ+gueJpksPaeoB52eMN3pb2v0kYbWj7UzQylKfMTBNSU3pOtCZfvJBS74nAzPi7zbNNW
a9cpM2Y3ukCCnVZ8YDTBdn5Lv+XupGOAw+NaJma8QgQq68dSedhj7DMv5ogq5xpFafSTJRFSJJ5L
+fkr7B6CxBzFe83Io7FLQTquWSlN/MOoMcmNzvKCkPq8mmdzsHMQ6CePQQgvTG0/rCLaM+55681Z
oev63EKtz1VV/zPK/Tqbse4nL6vhoNSBBWr6R8cb8jTZtWjB7Dcq0ACKqbk94c+KQ/LTozZcruk0
OyXGwEoKi6AeGVMZ5nxPbFlNqqyddGfeZt3SOdr1OYvXaFFIC0pL1EEzKYLzAuo9oHbxutbeDq4m
G+yF8VxUhiTq+DkUrufYAmfb9P42vwNYR2Cx7tb3shlo6/qWvA3nOyESBp6Yrpea67/CEK+2nFj9
jHK4uQCH2PoAgNpGTpEO7XBUOe4sAqYkpI5+2Ray5EsRarzHTCFqVPSOXxPQ6qWtDQTyCv8lWvad
beFrDZMHaDv8eGsUYhPcrN775cVO6nZ3nqWzXO6ZWus60npWqcyaIZzB+KCxl4EX32/M2ZQU625e
/lYhI0ptVZhLQ3AYmQF7qcw23f9OmhC5uVxuo03ev56FCmT5RjWuMarDfY8Vf6AMelnaSwqEqrz8
u2aaN6cd4iEFyxVRzNkfVJz2FNPbVcybAcZFfNBcxVodLPmTQVsXaQ9HdOHzE+zIReXtYsLJcqbQ
cn5yy+MoQX3rU5cmMEKQWs/ITmJoNZKWQVr0mLOYLuf/LaKPgdL2wWLqL00T4YARrz2eNG+DVCjU
V8lSBJbVCrKTF+Gel3+IXpPDZRvYa5pKBgG0AY1WkE651Vxjcfk5KQq2YE45PlUpw1dJ2t/Bq26X
6l6WshqvVSOLAh+JOyEg5TUffxytGrebDliY3DGjBxAi0qUjirhr3W2VIiy9OLZTRpv+8XhjmMet
YTAHPLFqrrGkOwA/LvWcgNI0O+I5GhSTbjxxVTulySBsThW0mPPO8agvbMYTxB7M3nBM5zyKj2D9
J0AoGQ56spH9nFs5h6g/nSeCTFAvWGAPIjUJowryEGlAuFHzzaUuk+01X9zRVbbE7jJATU2LzI3V
DsxUW/RHONq4rgjVbPrW8k4C5f6VLNFyoS2zR5cOZCuyyq6arHMY5YNsdpg/UIP/r480q3rS6VMr
C9FSKf9eAHlQGVuxH+FhrBntPugUsdTUaZmFNUIQ+E8KEwNyeHtt0LOS0M/ub6f22EuzoWErFMBH
l3pnhApo5OWocwOlGjkFsfHUHgEQxXf0xnSiISTRHtDQ6jFRtwAVbRabCXGWbyw2sk90+tOWYVY3
n5hI5/RU68sYTRsa0q3dxwcMoOtb0h0IeKc97gZcjVMOw7lx6V0VVWEU6G7LXRyG7wzJMiZ0VRBm
EXdgNwxepCOukumYBBrUzMT86qJ2LOmG2gCyTTM8hp6D4spdhrMpm0daMDy06WrG5VTqkVD/6oWk
HS4ZW8lFFIEUPSEjV9VI9/KWUlF1qgMau/G/DW/Yi7I7dtOj2N4c01asNahavmTQfE8OZl9d+0Zk
Jplg42FimwdvSaqYUM1w7vVjHEC/LeeEeX/zbVh571lPWjRqpr2ED/ZD/XahmXTp0TxfYz62dGEd
MBRuOho58c1dhsGMJUisbi0G0eyTRFb16C6jzLbmrlVQWf4vESQ7OGbveGNXgSKgj0HyeSySWmEe
kvySF1YhTrExNP+bpEfscqoV/tEDla9jartonMbSsPdIxYFiRjbZsSpWzMVrVvSnsyNyRMpLwZ3C
2WUHIrqKP8fnGX2aBRDb+cU8fyuK86J0P2PMFsb3M2tb9G918GWhlikJFvff7Q8wXQxvkWPQ5928
AyVdXyYeUzcX/W3KJQ7F4j6DrEKGP91J7g3eNhK5GeoUI8/z3jnY/rpatCLTabXBBuZInBo/TZAm
WFD5+B0XKpAXGpQnpD/ecimmKOpj+9Hgz9p1MbHaqLcn64ecDyRJSw74zJsX823nMjgTNOjOO2zY
AR3slkaOxpqVdOJjvfoeS0J4HSHdzf5h/oyBajKCvMO4iBe+BGRMgWIYRrUTm214WD/bBtOn+E4+
5Rx2TjuM4x4jzCIYSm60nRetZwTSf+slds/8MnJK8+1uwfkxBaFf9duedqjJLwmVxTqyVjgePxHH
gnPs5bfisIoHMwwtGX3OCNTHs0PE3nf2PLARF6+WXEd1axAAtCGhLHYww7NpuQkupf54uaB4PYqh
UXzJD2JLe9ih6TwYqO20hcNxQ/jQh9GVtm2bffRSvnb655g861xepBHsQq8j+Qw8R6TGYe6ffiEf
ZyAisLgO7u1rsFtoSvGJ/XW+zxp6bgmvmt1sIyVtR9mGG/+xQ5QJiDaw/oeHlSTIf0f5ksEk9qGu
BBjtb5UjTyxtyemzdxTpXy7SqxDOBvnWecQeGx9tepxifSKMzayPOn9cF0bK0otGohGHxOtLbPgg
A4xIbWITjou2ZWuLyq53D7XhQHv6TotO1RdFlU4Xj6eYmpxiZDiwt/MCzynx0oWhKgn3IO9VfhdV
7C1C2bxEwscC+yxoHCKXShY8xxQFN3zGxXanHGAPOJNOm9MkRnC3bYuz0C5IgNwP6XMzXj84fDny
uhTuXPwW4HdEY2rA1y+HcJqnDksZ59KEsY9P1ZY+nPIOgEx9MO3vp+WJjA6zTTo0FY8Qopad/t5k
/1tM8TdrZl/RkDWDXffAAzG7+LDdXfgT7YJrsPEkN77GPrx39or19Qd12BQG8hq46Q/6lKtuQGeD
AfBH8K/8fE+HKG2xADKZo3XGrvKuGzu2rliOrTkWpxr2y0puY0xCKZ1I8butEniOWPlz4FiQOGng
gkHhiXpFTGOnjMa9Cd/exhAe+4w544cfF7b5lXuJvfaTn1rWKy3lWrRp1EUZp8J5Vkm7uh7pMGFQ
pkyFNDcAd++H1c+QiBM4efbzHvUIrelAi3d8AXIHZElEVtknr+YsjZia/DCVECs4EGqLqhSpe41L
5PO/eF4hadafDTmcWmmMIthtGKMm05n8ApTKRQlmIzu3kH5QHo9W5+AUy3LeDu83XLiSPMMw9zYV
l8MiA0B+0INGx+F/3KVFaF5diWNIVFsT6l0auFnMuwkEGjzDiRe5YDSRTZKAILLEoCFU4ntVNYwz
qUF3hYkoYRPf8gfDaG59yU7yeE7zakc/LOYQxtAgNcO4fhHVS4IVI61CCVTjZSIAlJIo8zVY/Ayc
YHmfjHhlyQDii4jhcdXGPIanIHHTKtgl2vn74vN7PdoF39xuikJzvgpXVX/eofCfMftIPYQG6GsY
OzQ536rrveBavntuc6OqCFZ6PHksw5WDHbPsKTHb/q/swFgWPPJtbT+pvyC1hBQE5i7rSCH2I9PS
ooRoktFNGN2qoVPjGb69eYCNDxB3KSAnobY0LZObkWth6yGTAAc7Ql0m4VVYVyhGruohLM0dGvph
1wyP+qQrEBHwQX9BAOOfOcLDzfQrGQ4bTcMSE50pMhn9vzuExQmFhtRNvBmdcMkxUNZkkF8KK2wZ
YPRq8J1W7EX2t9d08EeTuRP7bp+Vds88oKaMy9lvDwQfjJNMYWD4rryWz7MVyJYC3LKptz+Vk67l
5YPQ+TYaAAR8bELgKHmyCHC4XzY0/opzh1Eja+ckBP+bAO3++ZK/FDbe0VThzw43j06NEsi8ZcqS
wPZdXJVUP7c5/bTlkWPvbdIR/y8RdUWGITgR1dKs/Dsw2iB0aM2NBcRN9VkjKHQYFtvj6Uebr2c1
yzhoz8zWzANkwe1A8ZHE2pCddVdWQsMxrNgXrjhNDvawiAQIFIHla7irLtz6MCuIsGnyGEfDw81E
zoSpX9vNKZvohLS27WcaixcapZ6rpr/KXVCjmkKBo8XxsDk/EB4XxQiEmE+uG8wIvVToSB0/HNC1
oMAk0gWfxM9rX1aDQ6qfvt4iLbLRNQk/KFkWf+5XkEG/XC82ysGPaORYHfp0FOKnNPcMhjc5I/Ux
bpId8pQ5t3grfBmUeCe0ErkVSG3ZogsxAZQRhbsBt/Wnjx3yM8fTp88APpX5DSDTB37PYJIVCESP
eio4ZR3IGBR3ayY+KotcaECoLuzbgww9kmPxMpw5gt1pu9k5aRycbWSHajZcnQrvNSXjfc+UXLOT
ka1TcvkmGmfD8O4RLNGM5GxMu2ib5WvVT56l6JD9YIBHkqWpBQbJAx43xPeGvPQrb7kN8Adflx1t
onIhLsQtQg/WPQk/bRHnKOD5Q9mwk3tNPSRXDDqMJSwlV+Jb8RvqtkECBWBJVAjRPiGemV7tVJpn
4Lr+hisF11VQbF//qxAh6Ed7VFB6vGi2mlyP/+CU8Qi5VlJXC3zDu/6hGb7Rrfg+vsm70lhOuobM
xHJg0MG7baBoIh95TQV6Sn0LUXKU3NqJNWfg6A6Jq01s3dbqNvsA1HzWqZWVqFOKgC4HFCvE2veT
AR4ilm33izp1q9QOIyOE6M8ECID5Bsgg7F+pZuuQrdtgFM/aUmrg1HOrhAmhdb6Nmb63PTSAYCQj
nqlg91S6MVN8gTTuPt6uxItoq45/Ch/5wWDJTgCOeBPhFpsoOUXWfllZm9p4YB1HNArxLmKudmbK
5L1ZiRXzurlzlB9PJUaIEclGSNaL6V+5jqwIfxuXAYACROmy7Y12gpa/MoXFvqh9hHkwVEUfNdfK
7bQDt54SJIkH+WXVev5pfhF7w2c2t52i0hRmOR9/NuRVF00TT6H1GQuenHrBrYK+oOUEzRo6Gsk+
usX8vTj4FwZX7A1WybNMKRD2aWwy/L1GFgFGeNd2mdVJl87FsMXMprfimRIFZz5WIM3h9kqndwri
gPLQ5imzonlyjPXK417K9uU3hXYPu8nmnZqTZoKsTtm9jlmNnlexrIKfojcWjUDzEsNLzZveToL3
zSBwB5BGbv3kPraXeeC6PThxMOKvV6Q2035klgvwYTwDWacGO8sCSMBmMCC30Ittw9WV64TRtCAg
YYr3FPpi16HnEAhYsp9Mx1BJ10KOz/CR/kqMpyYe/ILfIr3OSvrtbHAieMaMq+ZAliK7bYfieHpb
fF59CUNcfeQdbLGwqE8vvpQGNHdWHuw0vLcVukp1XOKpmAyDUy9gYSr2/NlfGmpNInHyzWJANsJ9
It2HZSwftZ7ubqxdMZgYjgFGakj5KeYcUq4RRLraFslbThx48z+mHz/qqjlMFZ4m4OkO50fNEhAG
lo+n7zVdsdo1T16SjZGgM7IoQxXohq+6JxqzX3mv0ikKWRxkbqplbkMfQMUEoEvAKDkyvh0WR3Gg
i809Wc3p6o24/FU1Cq1exN4fO3YHjZgOCn2cIe/KaN2Ty/mZy9E1/Cj0AEku5F3O233/sH4KeFqb
z1Ab118EfMF2VwaBwMPwkFKDoF5zo1bXYPz6hRW2xfDB42kAFhlxgVH02p8XTN35b8EgZlDQWWez
wtVyoOG/QGij5zQaqRf2KPO1qBDIViNJu/ye93VBiOpsPomuA8PH/MiVirI8CPvD0lXC6bIAvcFF
CAEz6Z3tj9h6ul8E/3yOaSfvy1pbPrYAreTf2wqgmVdUOPx9jG/QKz0SoZ1cYQNNPpMH9dMo1HUg
R2pFYssMkySuATWDOHVONzfW9pgk2TkAtnql3HWuJkgV1A85RuoqtZvCBHdwST7rEI647araGOhq
P7GDHAWjo6zuWqRzQKc2WZgQhCLEo1Lr2NbeZpuhXqpeGfjvVUwLAogr0439tECc5Wot/CNmF0M4
XG07puamXAcg3YxY/MoC2cvpcdovRzRjt5MdggFW/97A92C2gJXCvzOFXHal5vTrICMYnuMaU6aE
RCjARCY0uIu5mG4pl9qYzAynU7TezFDiYO89iMRoJvdSlFtj/JKUVoawlFQKMJGwnKro57UcszVm
V0B6md6oxDkix4k02YnoLILDs75LJts2rOwG8R/kjomNmus36oJp3KCWBzdsH4/tAS04meUJPaJL
E+IX0hylMcb45STDIloaiJAYR18GQMuBdR0YnUKDkZMeks/TYpxa0KqKa1STKdAtFCZwWSKL9eek
t0RGSiIOLff9wdwYCV1LQwdxvuma77FOTC2i0punstxj5eqOKlJcP+2nWqyGaMwWwzQaXhbOds7e
qW4tN1kRAZoP8uWbdm2ohMW0eex3Jfwy/Q+TlvJxzSqdlFLuDPxD8CJ0zucI6upedSAurxafoP0p
NBINW5PIeFm0JdxRf9WaiXoUhKi1+MnNvzdTzQ1NJRpR5A9rtbeTydy/79YvBDTmZGb98E2MWJL4
nT8qIZdQTGp/iUvpQa9y/Q/G7MVP8rQCBSouy/fweMsBEwaQZX1wPyeCuU75xBow4QEQMFD3qBr5
Yzxv39sE4AHDfNbImvdwlLhAUJLMLnOGfxFawKIixoIaD9qBZ2NFe9XRA+Z3Byha57Idv2CNrB3b
oyLarxsFXrCW6a/X4RHIFFcP4ZIeCsO1ZQzCtmOM9CUKv6Qs5wUROhO01PykV6jZHwLUa/067ijz
sOTDuzmmbvORBTydI0dA1TPE05KxtAG9gy6b0Tl2PGVHQlj9TWJ1/+nNxkTfBffzlg34vAsx074j
9R0MLT6TVq2FuNH3VtpRKY4h86WJRKEl2OBb6mD5a6rjkCsurKjLwixKwgWFZ09SuzXXygDiMmIb
E+7fKseNVXZPF9CN4XYFQ4lD/DNUG/5MC5q7kBM0bcn0DnaXcoZmA6L+z8BEpDvbW8K279zwUi+k
HBYS7WHGySCsdO8xa7bVNWDLH80Sdb29bfMc8LgyTB8dVmp33oZnTgY6pplel+nCPoPtlGg802zR
7YwjxMYXOhMsArLDUnx2Ronp13S0c9DIfGCLH5C3c097mwqKhawCtI19snPv9m/D8qXoxqjXeSHW
7kiNtQAGrvi4Z8KTTw7WtQ9P4P5lPfhY4Bh4id4RqiPpRALk3HxoxOd7wmcnRai0/xHoD1/IFkm0
FGclSotOOpRcFLbHjjhGE9XArVP5IZzjwmYrmmSUvrkrzUgfo97L+hAk6kjaxSuEIMJuDWTpYC79
BCyws1uHzwVsN5Y39iDJ2AKxqQdgF9dyR456QOCrznTDMi9An8LbVlx2gI6BkZXF2daRXUd6ySmk
/iNw07NmxZacLs4jtDIVVtUQZz/Dp0hB5sFLflDBOfW9zB++pXew5QAt8jWBV/d48RcWm2Cr0lkm
/o9LWIMoqx7Xh7V3gF5zx+h5gMcIM49empgFfQ8tZVPJ1wP4cuH3CKH1O9ilpXfZG0DNEhPgxjnC
LgdUeb8NFNTC/DN2OR5xamAo82DzuVUxmC5GqUsQFhxqUq5D6yuJEyZX3elyB4Dxp6weaKlyu8X3
dqQPKWzslwLJkl11no6sLV5NjFwCLb0sm12KqdHy3VcVm+ZuGUCUHWcs7lXyB/t6NntRgNn8qpuT
NfOMmp8bb9KV1Ug//PH5h1eH6NYfOzrFFxz3QOhUgzXHYtmF4YtQic+nYDS2kxGR3uwI9sr2x+cv
/6Lm1RZSQyy/WHLu8cG7O6NKhSmdoel2X59EjfwHaLA/+SkOMO4REfmsZ9lVPo3inUAIyvFDbMF/
I1S5aw5hp6L85fUHDK0334s9QjljeZixgqE6/tEAmQrJsfrJzMt6tTu4qXWewCm/J+d22Jts2FNM
1SJmazl7w4H+o0toE5lyEdSKsXRVlk9FvLcLvD95BeU1T9MeJlKfJ6QsSMglpK2SN8TzC4CeqeLb
Z4YO2niho9hrG2uR45jT3xXT0gu5fkzQn1kfi3S3x8gfRFNod43lTa0DT7YRvFBZPdYvCwtAvb9y
5P0WO6A/8Re53OKTSog3fb1OZHYqfwmkhbQQ50j5HYMwfVy88MbuiaoqDjk7dowfBZcIw7OZa1Oy
VYizq4AjIg2Uf0+ShJzzJkUv4cCOdlVjJ00Lh6+TkoWwg6HbEE4Mnkuo96ve47NHChbWJoNmGfcp
iBrohAarTckTmgWbX+OpgPQ03qA5qacf2Ph1JO2qJ/TNBnccxOL9xwI6rS6SS6KUVCQr6Tk0IVWT
NLXTgfq/Q70wSwLxlsQ3oTxMM1vveYFHPKZfQPUAnY0DxbJfo7wiW75mJuGXF47kGH9usfNtTrxp
XzNmXKBrfWSL37RExA8S/VohteSnww1xf2g5DPnyUYGlcjpyHMS7ow/9QRAK1Mzd3LRCT5bCLnuY
wd3In7B6HRIPKzC7SHj+msDSaiV8nEM4XpHK4y4jf4OPqAV94NZL7qkASA75u/gi6Peb4wVeHQk7
mDs7MlMZLkDYHywQJ2tPRs+wgii7VMUZFsdDMFGpI39mzRMaCBEhBMJTKvsXoLSYek9BpFRlxBOg
kbZds3J2cIobZgpYjPBKsX8qLjTLc5niVsUgR4W4bM8wQjJorzenQSXtGiYvCosNbvj3MJ2ZO9CI
lvkEZ5F8rfXjx2/gy3dTkrU2fE5Gw1jPEZrhTo0C+O7GqEP+/EyGnPyNAVN4XzyBS1BbclRADhc0
+pBRv/0CYSccio6gwdz4BbutFPwZjp1+ywvbDkusPLohHCQgEJfddAR6ydKOHrWov6/vhNcruj8T
2KjOAjEsiBo9UgUJhfR2Tz1y3rAUJH6TTyR72xTC4aOMncJ9znnNyIyvczqiONSwXgpeZLoIsojC
5COQFFIoXodMWi3XiWV/JfBVixKhRMIGq07bU+N6YCNytzMtskz52RUaAEm9chKkKZJX2eKIosST
Ia3feXooM3tiMldHSg1XHPm7kwwHXXLeMJRE6whxna0z+PLJ23pJpo21aU0Th/xl8Zb6gbjouxsX
xjoXGB9Gjl/7eW4MyYzbFiZa+TlmB4/QU3V1Ub6fYkkL4SAe3V3itOZ6I7SuyI1wjHzvhSKjGaxF
zIwTVT2Fe4MphycM8CdqlaIguN/SWhgqn3lsjL6Eo7vecoHp5JJzvSEaf7pYHpM8sJnjMP9IAWgh
rbMw1r/plECDbGEecJwJbL1f3IX/pY+laRPaDcZ1tLvfV81J2motUqZgbFFd1FcF/hT4SzlsyIIC
YFemP6yWYow/oA1LWUnG7xZ0pCQlvVq/Gx4OzJgI2fbDRja4zb0HRXFDUUwZ40k/cNfSyMG9Zwsn
oIT4da1ErPHVf/s0qSDb6V4MJofXmKjx7P2W3SzC/Z2cXh/gk6md4NlW3TaZ1OVrk4lLp4gjE9Dj
5sCe71HOZJ/QI274D4dlMTFPZbxUAo1I9SppeB1CO3CLa+q6AVP8o7WRXV1GYbJv/iEMQm6jTIUN
UHQAXegAxaUc49SDCEwBlojC2NUzhJ7ktve2rxs7WAfmpkQTVOPFB0/MKCPK5R7oeAgnG3HDC2a9
a7aqAZs9jkutwVB8gzhsgNklZ1KpETWDumkyJ2sGZoKBcJ/TV5OayR9E7pnLJRFW2AIe6p+WtKwr
XV9rVJMLR0DV9lDYndLqquoq10FS3hseJnozuEsJJqUQvBW5w8aeISJ9++qGBqNdujrux9qOVNJ2
g/YroWR3SsLtgG3d3OFDEfTbD/ARmcc33cM4i/EB/JxivwSh6EGrCfVIIznjRYUYkHGNze9wkvd+
piENuRfpw8cA4RviZDCiXg5Z8wut3b5mZ8pc2Y9LFd7PysRiocvzwNTU2rQlEFrs+91feZoHvR5B
fLdYkUJODFow6dt23nIOpBhYSgGU6ot0S/BsfJ1S4mPifLDzCPLefKHNDVn4wm9PeNpkRxFegeAe
W5RdskM5vPE2crKqPwst2VIiPn70W1zx6D3G+e6GI0KgEf9Oiu7QISdhMz2cdVwd7S0SjM5Az1tx
cZD/vUkzvC0cdtQXOffygxy7aaKcyJvgoWjffuAZWoj77JUO78RyhIaToVquM5JvPf5t+ozFTXvX
5xu1L3I3oO+cu6EGWngKsFKOLk19dBBR8V3oR49OfmlQu9OLgS+LZIUkqoMx5PLoD2cxM16MFkVC
U/1xUP345iW0HoOCtXMc3W6F/XK3k6pTSxT6eg2JB8X+fP9269m74GTYja6l12gINCH0D53J2X+a
2PW7Gg/j0wH59MrXpEhSc4bZENImwEfhMPjRS9nm2PnrndhxpCHiLny7APRqS8qJBMNXldkbpzno
/UXyTBAiNhWRmbfSc+xYDgtrqRhyQsJBoTtNRn49ugsqOn2tAsleAShwLPNukta7yG41KGPnsQfR
IsYoPVdRvbFgLxi5gr1pmIJ9XGIyxQpzBjiqVsBwVlPCKeAANv9VXXwD3V9Txfu7955fRVH4+3K9
zj0XBeU6/A8kAULqVsGRRHw1epGTSvztgODPfwG3ZsXmNNgWlKJrpj2gYMmBOHyaqQ0rQA+fxvc0
1xJuAdQgNDsoQz9jbiBocABqVmiGCwbz3OOdOuIIM11a2J1RmL+H/koyYfjuIdH+ePzLk1YZ0t6e
A9f/PygwtI/Ah6t4x2XW2RWTZjnRsVpq2AyXgKo05Dh0/7nh1Fzq9p2ERIRvsRiPDawp/XkmOvRt
pUqYnjXY1U8U5kWqFHUf75QqzAw0OU1voWJaTQ6ox5KNQvFusg7MvJ8OCpuMYLompsox6kOA9tmG
wg27MuFJjIWU/xOuO/LankoUEIhpevrlh1x/um31uV+NIWAgUeGo25J/BxPwvi4ETSLlUllRD2jf
27I5glw1BLB1sesNPJh6+AebxKtbuBd1vN1aLMReBq4OD2gHo+yMnMBwC5Bp4RCoSehjPJxgp04g
QyFqRRObA8dpD5Ifq9afFBtPLhFOMl4eOBlXpB4mRNHISza//41XQ9NcCAm7Qt78aklvb42ZkBv4
O0zmeeOzQuQL1+/Qjz5ToXqK1Ri17mn9G+FA2YvzMAQBzEkqWhkho9kQwTVHwU01UVj+d43bOfCp
enYRId8STiZhwGnRz7rKvLcTU4c+40OeRBpb72Y13AtqpuxXufw0baVcxx52lMh+N1tuFWXBj3Xs
kQ4ChHIdVjrQKhRJd+I3yVSY7DHTJ0EUaFefcfZ+vUzqxEudoaO6MrSieuBfn8a3Wj0Y3ejTcS2J
8EX77hGM7rnGsq/5ZPMVgDZMQe1tY5fTxq/+uQfVWrbAWC9FEO7W8MK3jTcAALw5kVwyqivA2ycG
95EL6TpYDj/zx3ODrdk1ASszhFMgnT7V65jmaCBCdJ3gzl51PAqfLY1mQxd4cUupr7DHbp3foaVN
tqwaUr4dVUjLCV/PDx3GzURR3PFDSRPBDLWetC50ubfifkuanoXDg/DJGydjmDOlCz53EUBI/7Lw
emMtBKKyjBcqm5yveUZBna+rOsHlZxHyXccKjmZdkJehlphlaA4yJyuasiA78TEyBCR7xtFGZV8T
S+iRsx1KvlgavqjFxx60YH7BZtD2dh6W8abE8Qwjuso3Jo0pNl7Pm4QbQDjZbulZU+IPiQxDgVRm
LVyyJIVVS2IuxGmyBpJITiFCdzlUjjcQTqgG+XECMU8AC5DH7+ew8mYV2MI8l/KHRgRMHDfCaIYN
kw9UstiQ2htUnc6QPWirpAeBweU2O0OrEHrlDeAV9bhG7UitPk4tqq7odYdavQSAPmklI+6t3vZc
tDbTwDf5gUfl1vi6ZTxRDTI12o0IGDC7IEj6ludmmMBQ2A9QuCrE9Ewd2ErrKGLuyot+v6kU8KBt
HM5JQG6R8Ep/2sUl9euWtjxHN7ZmxVMNHn9mN2cOVEkl15tzFu+N5k9mYojYsslLDb31zYUOx3nH
jxM7mUP08AwEBOaoMTSw0aBe5em2M+VpoYGnKbgXh7zI8g4yt6WENUdxfoC8K4o1t0EWN58rB9qI
Zcm10P3Mwh9mXfULHi7GzCStlWO9+oT+u6dUPpLMRzGup+d+e08cXYzZdcJVDZ1VeCjvdDjH7xDj
n5z5CUw4tJdGOfoRw/Y0YkqfLVkayJRpk7qkjyT7HxFnAGulz8IuemMgmxZ49Q+kbJRUGkDbviDd
zIbwLA7QX34SNF6PyC+DmCa3+TK9M+/oeJDC+XozDmFajpFAX0JKN5gbxTqUhdupK4QJmaGcdXHm
+jhfxxl9IDzKeWj4k29mbXFJ6OUdJhVYpvqNvp/rIiHJrj1LVRUPsFazsqGjSD1bNcZZcqXn7sM1
OV4+VZAaubQMnqL51lHz/voZoEWSpkQ1XcB9qh0fqW+1jIkYjIsPoYBCW5O0+JiAagOn4cKkbhhQ
xTJRB1Q6796KbMqzlEdgH8EWNfwqU+stdMV1bojoacNSh7ULqPo+nhaV02QQa7X/lf7fK324tDmA
eZ6dCTwJu3A0qRKaBKRWCapBZEPzCicCEAgQq6W+pqQYbFQlH2tQu39pXFH7ORW92LQq9zE5je9p
MMTFwoQS5tv7LeUMejp+/3n4twvBTpow8r3HD2AyQJTScwin9o2hXS6GWONuIWkJfO2S1LpZjyH0
srx55ymqW64zGWdeQh3cjNc8RKyBdpbGB2Zswf6weQzC9J/O5cashEFoutAA95nMOaMTla8eC+/2
NvXAF4KbxsUwAPwDYBrlIMaVanHyMoDxc9yfcPpGK/QDm4xwpo9DQk7633T+Kuf8JIiBoZAdlErp
M4zjYZF+tHq234n5FGF30PQZN2sU6L3Hd59N6qABO8zZ4RFvO8gSofsJRMccnZlqcKPw2z5bTtJA
Q7zllNmhx0zirzKB+QuyNgHfYmG3xWlGKtDGwkdCi68Cci90vjnZ7bdL2Rxv1jtbrrGc+SsK6bOt
8ErB3A6q/ekTPLxS3KTWkygomYJoNXnA1/FWwXq0NOo2WfKRLnEAurW6/UZ0Dt7ouFfla7Ng4N/Q
xG1+KBfTjCUAhr6RxEMWF4ADquglVEEHG7HcOOw1klJNpAyL/20O676ZksgdiwjQXBTrt6v8Q4Cn
p0OJ9Ksv38mT+TjgtyJ2vPCWL8oWEd32OyAGyInLXMsb1oVAqUJbgX1aS71WN7CaJmwexkk2FvMG
eBN/w1ZY0U6fI8m2AsNosDLbozeRQUuj7vRMhgq9tg/gg6MQmsNrwHR/Ow9hoBDG1QPy/xNTGVLM
Dhgul5wb1ydC+ThcGOrkczQ4LbfWKRH2L0A1bh/0xica3QUm9BCutvRfrh+u54TG88RSDjy91fJh
gmnIr3HjycfOLJN7Y3fjXuo5oDoXWqLj8kedWXB8zd+VzkWE2fWbCDnjz8oeXytMHNL/7YPR0zmV
4CyzQL2ucE7vt9szulksEOSxyakw5MrFWY4FRqRurme5bwF3ffG5TqT0FkWWiHHH8FnrZl8n+pIj
hcYE20CfiZ7PrbnutHCcLk64lEWozvHBiNE4FNIidbc5zwaiTLr9CsY9Ld3Jox5wI17zUXJ3DCBE
4ekFnbqoE0x/NxUk4/GGaRyeBKIsbnmc1rDGPw7au3nt1V/TAjGLlKwPkQurvVSYg8sr6BlkR8Nq
TcwnFYjizKrHyGU46NFD+BRhVnOXqXjrzZiKnQ5/BRTfJ3n4QKjqVaMtR52qq9EuKZaxr8FB3oLh
Zj9QsTVUIeYaZIiRzjXBsY6VN69OnU27ZnxT6CsepjFzYWwXUqRD83JDYTaPUsIIkIjpRofeeWjg
C6r0E4WIkIDE22YUGkjUuyV3wLmt5GX74TRFbEJYb25eZpuwxY5hOP/q4JR9FsXRDmahCTYMKKfD
+54pR9+UpG2UKHa39gyUJ2HwxFzf0AejQtVYe/M/WXSsfAj/HiJ7zC+ysFLh099JHOW9/9zoIgfX
oMdXl77NvKm21ZeVQBkvkdFxWnGFslqzOyzLxTP/VIOMdPO1b47Tev96YgRT/iBKnPh5/n175UQU
6YsgYNcs38I2kWnrBM1sO7dXgzmxsfB5KFfQ7xzcZMwxdZ4z2Blc64WZE/AiRxDYI20Q1nTDQb9y
6nj3HGt9bsdaqIoH+jvs6o/m3tZPF2cRDC3NyCF02AmT1kGBKA26LmZ0yyR9Pt3WI+uPzxgd9qD5
+vC8F1xUsyjTSamyYmGHwtVBrD71Yz89HpG3ZLH2tS1CR5fyWww0AxcRH27mH2XOX/7KRglXU5o2
fbQt8n2boLgdXGX6v31llU889xl018Da40r/MXHcQ9YK/CBq+KC1K9dsY6e9zuA35FG1JJy6jj+g
4wLhN73H4ng8bu+UoXSF1NVbpjUsU254YOlZOjB4p3rOgLhmdcpBBy4tEOzQyOpKuSemtJH4OAx8
mMWpJLCqFZL/TbhbQvvhxJ7p7Tb+Xhg84+K4riy6T3HeWJyUn7kX3O7dYw3gL+T7YxlSB+TKG4en
sA76MYGFZsPza4o8alX/dUKE5TryLXGfG9XwHyOGRYwY8PKggO62rs0DUtdYHvTUnMU2oTBYu82U
nX8LVIATM6u60+LZEDfb0tbxRVn+O6xr3GhsaBeuKeE5CDhpM8NOBK7vQfRyV+dEzRnnGkixs6Bx
lt5O5e3oAp5RCfAfiz00tYS6BQjbhtYvIB0O/hGJJVrd0ddNFffaQChHfVfTLu3t3OpqrIkS42RI
nfygF5pc4MMfG17A7XCYK+ulWYLNHnrOUKAEtgfSFI2+BC11L2xk4NfilWswfbTGYHmbN2UQIun0
PJ/uuy+EVcoElbm7HSPyhPSJeS3uy6/0GRys2vNhx0w3jKQ1eO3KhmyzaJb4DZhbWUc/EIutYz6B
w0yCP5wYsaE+PKpejcttQqlxdQsr2J1a0SqEkjjW9zS8imkdMEqoZERiy1JzDcM9puczwO2G4jsB
bjaF2JieIFMxhMG3sNNFxYOMoZPihI390V5mrEWtOLCyCJduTU9LP37Q+9p2DUgoh2VPl0rAWUQI
2eR7p8HYhaCyTqOrTSVECKS59gNdfsKgxVcxUBK/eaKf0D85sApTRKUIt9FbOOenGVrmWey6bQG1
000dKJkMrperTNki+C1mWifgfQLcZY/XgX0g4CtBVGHa5NJaAjv6QZmF89yFPx+zW96volFzr291
5g180TvPbZ9jFvPwEEICMCwldYecRjMNptj0FRmKuRklG8Bh6LzsyJtPsGr5Xvra/Saf5ftERi3p
yuQ3g2wrAr400tHjZEh/Wo1Ug5ndqGCwTzd5aRnbodaWAlsnUjcdgTLvS+NKpXzIoHeQ2krXvyqB
i2I7S9BLrsR5VLo/w8raGtoTjsZOdxZ6mB8F+nELY2ZIXgLw3YQmKlBz+EYWnXxdvOLg2sAeQjXg
IuDQErqy5mQzmNn7HdxwtVogkjeUSCee6XJjH0gug80OCpMmdvkBHhwIrltbgLIKSNhx+tRCsuLD
wtagOQc2RdiLXSpot+TcSnISA30TB7cSRh/MRRa5tno1RsVU3dEu6TNCFXI4xPUTU9xetmWnz3Zd
LCyNIzx7f0sjrRsBxsKvftiNFP+iPlTNBdFzeGxCYbCpO3vH1RMeNNkeoCwsPevyEAeDtwCDC+9s
BH5mIHa7cdtpnlg2ZxolZQdR5U1ZLgERkV4oq8GVfp5QiC+ufX1MqJiLvFYU6xZuqrGgddNRHxrT
TYISEcYJVbbwRXPnLGCHJ5EXzuojQdcobVCTAYcZdyGmfk4do48KU376VPLJgXYSZOXE9/bm2Grr
4bPDpbMUlU6hExFyIj/C0kSH4txrOli6ufOH5AprOPyFBJzpV2EgmFrgt5UGknFiWEJMZZiHnXGK
B3v6GIfwB1rgH6S7Y7uuxCjVtsvgI37DDFwR9P3Q/Q0eGwxZO/EZErIFdpFeW/EZ0EaIylCyvAk0
jc8vEc82Qc9hvxzwrOwJiEuDzSazypcuoxRkJ1DeyLqRPEwAonerziogBzRkdgLbi7x33E8cBJ1S
R10ZsyLkYBcRnTEMIppuycs4KCe6gPe6GLs3I4ldCHImH2pOcs4l9PW3EiaygRrB/iS9+ehJRCFE
uYhQEMmcEmgdzD3eLIlR6H/aYwwdxwwpU78vZIPbnTgupFiqyTp10sT+oMVFakmtiOQNu9agtNWl
SRXkomFum7mHU5syaW/h23e1uRxDhhLYTRqYVbq0LbMSdPkt6L4ci6zGIoEAv2ZCQIF0Zhf4TwdH
2mzpSMIz/SIDkXIM3ryPr9PReI8i2Ph8rA5EP1KEyAMLce8oh9kJY/Ve+FQip9ca3MPIsRJSr/Dq
BmC5u1L6RWRldr/a03Jm+W0G//vdvvpJdr2YqBYNjqisFQe28CpZUMqonaAAxaYjX7PgMozMe2Fc
g6yPhZtkfmoFiAnIgV3g4Vecs4UEtMpIttiznAFdtoZKrDBy61G9Zps1HfonZHHkR1wwekIvjcQo
I765X8027YCUtuyEy298Udy2WmGRGTuvuIxO69gMj1eS9VQ74WqpcpGt2V1o/CrESEUcDpeMSPIw
qrqBN7qv9FsIwyP9Ie/aqAJV8zYCLoS6wUIboNhuJ7MZS8u2oVwjmgXi8nyPPt23cHHEMeciXXK8
UJK6VuFGkJHTgoDfFtFJY7jdBQHOjxrpQ3TyiQpXXaxXdIkEcib6phRHXMswltgf/ZNawZZmf2Cq
/sVXVVcYBNRL7zAl0agZHKe4hCDR6VBspytk0q4pHpLt5qXVrBm16aeU0ke5i6zox2JbIoBla6tp
Gw3zpwGrJGbEJf2s3ozGjoThtILH0O1JeYZsJGp4pK5Bd66UhuMv1h4XR+OQP3CTeK25uzmrsFG2
gAgXC74Xv/G9yIFBONdj1ADFIsthwsv3qxkD7ILLpUA06DwIqmPHNfoqLdW+76gRIshglhdp5EjR
lV5jDIctEMiU/VA9daAkSXyY0P05cP2cIjGpo9LmMfUHBEr1x+c0b+4slD7ETsm2910Zdw6zpbPc
eyiyZ9xQC7jBnsZwDutcrtRUP76Wm+A2Cv4Jt3eaqvp6b9VdG0QEYmtSr3kWg4avTpt4Ok72pKeQ
G4yXx8XAjFnPApr7wUCxOkmcz/rPej2RX+ZDSu68H0/54D+x2G3Ajqby5N3D/N9xs3ElMhjyYJ33
eAUP3AmJLiSZ4CW528jxKzJVxVFdxO8hKAu/tLUu8yNVlPlV9CqYyCnyWOXFCtDmFVR7SDM/59rK
QtfgNVx2dIBkN8XTukf6a8HobG7T9/qppEYS7QNfgvUEDAgTdOfQhajEXcNZKcdQt5xrHZuTxdYf
CP89zJcuc7sBBd6rWQ47ARCS71xngSIGo/tFmjSGTQebz7BHha7P2oMV4aVSz3G7qucOSdNeWmaM
lpRuTkRVRxA63U22OTTdVX+/PM2e329vWvl07IY6EXML5vshde8FNzn8dDAP0NUh+WaO80+9bG3D
xJugHqpJg3qPsrAX4m7uxD2Ew7KXxhwTE5WLjLoYejPIXWu+5eAGhA2Y5ZoWRGW5IsyXW7+OhAke
8T8KSf+6Ht0L0/IYsfeZ09GtlyUxo1W0jh5UWxA20e0FXIFP5GDa22j4PqK5wamCArM7OFuTiCKc
eWumVq/kgxQKYh5+RbdfI2q1bWk+CP3z26Ob81EH1LG0Rm8seJXKqp0B3xr/5XU7XUOU96fxcPv8
m/gFgeaE0pTfP0LVi488BxJ7EWIRQ5hKZ85xoe/6npx4+DFSWLgh+/W1ZjoGrP4XqlgBf5Iwbf37
4MQpFGJBoPMm3gLo1VrEEsM6XF74REYHuf01Ohy+rF01/KcdRu5IZ10CFTAS2xobDOrnz0XL2LLX
gUVS+6bsx3lD+Jwz18du3H2hf6XwhCGgwCUVjkcL55pcwbK9y8IHy65b7KEByP+8F9OeBzgJQV+J
botV0NCIzcuPzYaUjglNr3gQnSGslGGu9wDgReUKRyEuVepcXmSeiOoh7g9A6aq0dbponvPAsjEl
ZN3g7TPwB+jSmyYsEyJIbqbb1omUPno0dLQevgrSTrcjW2Y+25o7YLUqCnw4W1QWMljgc2xQMemz
SPuyL2x8ail12XK33TanovgL6vZxxTPaf6ktkFmGNsYzmRDMpVqCIgkjXxHBaJPO584I6hiIYb1l
XsY7hwLbTOVQu13JccXh5avzFPN84o2ETFxYIMGIyAVTfTcIB/allShUIKKrFoPI3wGAJXgHCtGY
PV9S6WBGD8CwdmBw0gCRcYQAHkvR2FOppwXcwLh2DGjCvLs63zcCAL8/baEh7IOtjy6QijrJ1Ff8
3SVJTs8jLcfLBsfDPXVO+So6b7yEw9MMSmSNsBl9QI1EMCyZde/FYzvrWOQKHCAvtsFYLSrIMioU
IfJ0FysmthEB/U4ytNejH5xe/2/LQaFgrKK3axpqgBTf9x/uXqqnbQlU1zaceagVe4NYFItqGSV5
LhYCaHBzPqRMvwE2ghPPVb2RR2KJXClbBo59scY6P5xdTXqIcg4mJTR94neOhtaSaQ3uZ9J0vTTg
3KXxH29h8laI2jb98mJp/SPz9+aR5RJToWm0QKkJ1G/++al0iUdbLNGYSDW/dv7Fhd/N8FYmCYYm
EbMWLFUX4T20yz6GJr+Lq/yfb6R5hSMnOKmVF11cpJK9MMtxneS2JF0FXg5i0Hu0hSYvgf5cFg3M
jaMnfH6feoEIvGVku/1729JZ8YLmu8jeMvldnW1esEaGM0b9AxR1o+s7MkQeXnSGh4rtIvEto8ss
GVvVhRLwsAJYlKKPzj+UTdITky0bGiHMQ5zwqlVesgHagXgrm3NbYAbHiBI0qiKAu23jYx/UOabX
Zt+yoMcsVj8NiB+fDxfE/8beyJiqTlYnrTf9qIutH0sXOraXiYxUj32byGQ5hlOqzNV8tO+ifKaY
3UffnrCfFuqOaLeDVVGROA6GQHJBja4DArUBWDNRxukBwSAxtu+FWSEjDn4dzgjtbqnOjP/Ut6Sd
7hNs/4/sho9gS+Pyvio9r4Cj/59li26XS0DwISqmIhCR1ENFb8jzbdlwiqixZ9VxtIvGMhIhqIHk
w27BhfdV6jVj8gXIL2LvwOc15xnMso5MchVwK2lqNaecaK0Ai4dzmzW2mGq+nXsb8n2ObtKWHb+P
QU2AAPqkawjgMnQcXmDRfIuw2DxBd8j1THePpi0UImqinTFRZe0cRD0U8w7wJT66EQXIVpDomRAw
Vho7gsYYWiMRnlRFGNT1XMBEo7iI5UOesrpxMrCzA9H5oh9j5ssqF6ppymAZ/xzKbDBEyINBLwsQ
RVkl1K8VO3oN3NyX5RrBLo6rmIZojNpOyFJRYgbIaXuJj8Vr1/JlUjIOxBMqDk3wLXoYnqUMmY7p
OKSwgCJtOZ9E7l1122gWjU8kki0xbdZ9PNDzJsdvUc/uX09CX2ZgDZXqTR4UTN6ayKue7zXvA6BS
kEZFKQ1hhAuRr0HGUxsNcGOT7ktuQyiV6rrJTIKaSFbP5Ibg7h9mGzDjg7SUnRqoZ0dDVK5cyLq8
MTanM1ycz7Btek6Eepna5MgfpW8SUKmflY6J7V11IBeb5knIIixTrQy2hEITXPch8VAuUUkWXDnR
+omrnFluiX03+cVB49aT2c+Pb8QPKmtZfUV/uMxC3oXVEdUhx5aZFH/BscEN9q4AEz8RFO8tilCe
i5l1J6jNLayC/8K9Ug1gv0I0SgsVj7P2DoqGw5ullC1uJf3J0WpehVOsMzNPpqY3cACxLdPPOJzg
5I3sk6sm0GxTj/9olCYY7Sx0WJK2mdb9M+zY2hlfVM7qD0XrgOha9/i/yVZ/v3D/9dsiYuLn2C/P
9u5ZLkr79MZLxvwMKKy2uDkFTkv/ziUzIhH72RrGdr30zRK4JzpYw/MGlNTH0pwccid8Z2JEZiOH
yUhs0WMVR2eHSCjtBxVv3bSTIo8Qrrz7T11nllKp87LoMQWTxnsin2C1zi0871HHvr79bRE/IG0j
et0A/XIzAL6eZ3w1qE8ku6KA8hXxm4ENe3ImusPYCyXt6v/Nm1dy3ir6oXZtVQQh1jMv3kvM6aQb
6+/Bg1vCTpDBd66kgmHRZIMoUaTObd77c+YFHH1NJaEZAcRejQEHwRUeNPwgftQbkBJ+d6SuYLBL
NtU6FiqIhAC0D9g7HFO5nPyMz9xhyTZIPDwVcMKz5Uzr7Mm6oHi3NCwcxNKG3yyvirhlL63XmrXm
OOn286eH//4ajkZLW1gwGn0TLutErt+DSqfw1bK+8UT2s5bkJb+AHriJJqYKLTzg3JqUaY45eTm6
8BPHTrcUcLR8IodCxmH44gBFw2mLiY4OLrF4oroxzV4fseHqk63VB1qfeAYty0UliUGTkdM5u6zO
2ZKt6PMv7qLGa1VYuoXD3xbR/MeV3OEkya4UgwqGrjYze3SxuedFJtvaKgBkPaNBAcsKeHb8VmSK
rDUAfnSG+8niQrztAlvwguPL1O7eehuueWCKgaOylWBrQe2XqienVM0gfk/N3DTqj2de3mEiAByF
xhq41y5h1G0toImg+es/Y01LQ6BxhQl0HABxgQZbJkBpoOyrltTT9HuEXaWBtSyX2m9vtp36woDc
ASEsojBLcQtzy3P2R88xT/cCYkEcusFxLbBjjR7oNuim6lKFYY2NQawLD8pPEBWyxYp5Dzm9pJ1M
UUGA/y6J0qOo6aIRjC5PvnWAUrJKdPTmQSBE7JNjogcBfNNihMVxcm1fad+rHiQ2eqRlx17HActq
ETcxcUQUZwVZh5pp/tascvDiz/DqROLAdJDbhgn3HpZGKQXl3CSQ+sFnidn+xt1gH82X8+h1VH+D
TU5Vp9qJCtXxEqyjFLjhBh5jefm7QrLYXAUfc2xOUjY6dcq+gPe1DV+gftfqae9lRmBUg9/VCcb6
oYkHE+IZ2OoqkBZ0fckr6uc3xliIKObWXN2J8/wr+BO697osSbITyhG8wacnGExn3hsy0WyVC57Y
vmM3gwSQLRncsJ+N5eb+S1bLk4C8UXba3YhRyjU5oE245vYqHZg6rxlH16kxckl4bGHNOzCMpGPA
0UMBunAOAQxxVPDP4YChc3uEoege/UX+gPhi4KCn+acftqFN0GfDSBi6edtzuDdQrjcFUw+IyXJ5
+a8JgnNEmATpA4eOGGIQ9DvQHnD8Q7QkXG1WDN91I7Gro/fPYfcwqzdtozH1dKF9Bt9QBREWqB46
uN5x80WkSIAp3Dpbzo/sLf9rHk0YW5UtPLExiatqN6hUKFqS/nQY0mMBB4T2lsAWiQeIF8/WIdHR
bNzG5sVbFxVk4VwoXCo0l9kObShZNxLSj9bCWbKcJpAp68Q7bh4/iRW813tSshueSFdHVsj677wt
XRqFme3YZM9bp93OMGMCUGxuWxa0zbr0ix4sjMvSNMiZK1jaxbBMb7c/Avbt5Mvvd/7T9O3Bk8yy
LXGa48NQHkAMwLMK91CIHcXhC5hWJP9WkcfdBBGBi/t4L7gLUl7NxOkqV1/H42lwZTomDfgKKdhD
xEjO9TN5iZFjVFmhTC9VFk/fcX4/CG2BWBVb0CbyEm6IIv1r5R76GnE0UVEgPNsYmDyUlpOlUF/G
S91ZuefwPsAKEJQd/JjQS1PtLqXbnC9+Or7Kdb9RmlTYrcjuhoe6wpkoXhkKonXep1aiRiHBpuyd
OBRzI+Gt2raOAW6xQalfeDLODHZTTq8hXfpvkGLhe4OecwRmyb6iUy1BBaS10OCC1VdApp25Q577
YliQ6hRANZLttMJFsrk57AlLnUtuPhZSpSfO86RKpYEFGN5cGMSf9nMm7IUAoBj2CUVfmdGEhiX3
ZJJxqUkil0HEV1CScCv0udOuzyd+rB17XkbA3DHdbfIwaE8lRUT2o2tqYfSovcyel2MSimSuLi4j
wVG8qsSdDK02jKoCnwBuvTwLrGpNppLJFzqVzxM8WJ+YrYi/gB4dUYz0tQ7UnTChe8+5S0UOBusu
CeREmc2sM8uLgGWqW+Ta8BcTdxHa4KSkvEUNvSDPkN0MUewBHJXpI9SkaHjG07wO/HVHjzS+2Shn
d89YB3uE+1sM7QxFVeCkxFybVIMXsCeg/qdbKN9UCStgYGUlFLh+lTIdVGsyuIOUvromnYw9WTSq
y5uGjmZLb3ussEl8ntw/s5d9QD28ShnfbsUolVs7rR9aCL1CdaPmFgfK4mdV+Wt105De8j3H8dUi
zdcwRwqBUR7NrniBPF+zR9P2Fh5RqQ95WGubUboY4cdDCq/8nZPa4IBQzOzxOcXkbsBD0K6a/jf8
i2trBg+jpvRMEvEiQ89sD/B8y2NdNZ1dwvAX0xt/t3j0CuIWk2qxYPS7W6N7TI4xOXeg/+oJMeav
p+TW+RgWA/tMQwxpRLyJCZc/G8/BeFpdF8GpHKsKvfCYoIzu2LcdFB0fFKQLbqYuuIhJz459y0X+
Q2bOBxiCH9OFzhubRT8KMMeX5bJOvbRckA9KNHfsFHkQ5P8WrJQqo6G2tE8h0KDA03wXVucm2ILe
X9RWH31x4j3DkrsvKvGrz0z6GmEMmy7qu/mrx9B6ciKREA2U55MsfeJbLq+s+UES/R+ef6bHTyKi
rUvSy4bJDXnvB6J1iNRCpFGxDGXawWidRXpoJbz7i62PL6PQbsvUqUkAU8B2QHZ3xMDZ2BazxwjC
UGNs0RVxtvsQ5huL18y3jCq2kP5o9jMvY4e13LljShKsLg8mD0AagU/t1dGpz1/Gh2Thfymk1Oc1
r7x9sVHsUBgBtgwGn2aYEOlNZjxEPyUGzSMzS4rWEqPd/8y6Rhy5XhmrgTtjXiKfvgvjmcLUDN4B
iCfRXzAyxSesSsJtUqkR+9Ug4Zmn74CCK1lEq4jwEUieDvcf8tJ5hKHmZZzvJsEq2nrXsdheaYsv
amW5gw+XRu4pD8g9rW8XYFeefbD2Wu+am4VLUCyZR3loRJBNvyFe9VHev6yqCdmjMQEZHgX+Y/9h
A1TV8GmEdJmYPIYI0tigvEy7dAg2+jL7aWEyd6g6WtaOW7wwuiqnvibaowWJlJmkde9MH89k/iCj
tylpELPubmZhqHZgkUZTiiFcxz8VUp6/AhRLeuia5H3lT50NDRfbQJTjrhP8lV60XJm3IMGURv48
TZXVwLC5N1bP1eUEaqIrX71Ge7nxFVKmceVutLm/pp7JKy+JP2VzEsdMxS5A4Gk1N7ZRonirtJTt
algK/K9DFSZODv8ZCk1yqh92AHUpV77fx4YcxbazQnT0iw7RwqhdNb/0a1061u8nXHV3qwI3hsz9
/XUuo1FVfCgSGiXgKuk4N4uT2K6/vZxwvHvzzQCeo0VrFPJmvMQ+BoW0O78XtVJpQm/QHK2dhfX4
QIGrWWeVRPxNR/aS2ZFoEnHUobnTd1HzcyumKjYpKYRj7y8XS4VFLFFx602z/HM48JrkgPigLA8Z
R66MH9W7VoPHmoYZ4L4tT/NcmmHrmf/BB1+RuPxGhL3Q4QoV+RCLHtomRk5msXFyF/no5t08VqmN
wgeyEd3plrwGwhR3LKb083z7LXwFgMlPR0jyOGRlZ99Dj4Y/12ETYu+EKm6DNA61sNpSJKHPFp2G
09dEX3jBuN520fYESfWVp+a6LOzzxQiDgFxHSGRX4N70Kz52R0rK1N0hsAWn0bFpyb5phzcPKvCS
SCfmfJ3qlyZZOyUPPIVrtxSOcU2DViQLnQ0R47QUvYP6fRe/0TqxY32PPBxNL15Ps9Y6Ix09ETfG
Cz1fIsc2+SlFckBPB3+aH3wQgJw+rm3gIvNSFvtD1nL9vMwyHOp6s0TSMCbSe24NGYQOCV5EgwVy
izNv+xyPFCl22hHEtIrummivOsqQkB7RlJe3E2CRLh3lRiryGl6+YTBfalNefurzqZir6OAWNMgT
jDO9a7SP02QoI0pvBGta6zeisbkXEft7z5UvQdGqgX/Ie2o+qhDjgkiIO6Fh5sUIsQ2u4lFnv/x5
j6ngAIaQ7HBx61I/fs5o9XE63iu9uCo9cp7AAFaa2PQimH/+/eBhzrkQwCOQJraYNia8gMAdYaZO
2UDBLoVaTwicZ56+byu/s6VpJNDugScyBYaA5x4t86q6x4apNLL4AfByx4VvMGNlbp3/Gx9tgLsg
0K39vnSqPBZdadpQo1BHBL8C1xPFyrXOYg3f8VPjmtU6yZKMc010k7UtY2JOS4k/QqRsvjfT6ziM
4tm76M9u34FxgVntfrTXEHvsJ8NPctlSCwMzwpCv/nwiL3AgeKH5dZspLWhXi4DLpg5qMusV7LcH
VSwnGGEPW66MvvQFclxEEsvygv2oyvaWo4RIs7L1surqxhPn3gg9KeTjPV5ub6XjogD51OtPp58d
S8kyI4SgtkMRDW6udcpq1IT0EvaaDNv5z6VKUT6/5TOsIYC/BCGdQxWqIO5bL9s/Cj3Y8nYeSG7y
u8/hR+CB2QpsmxxB75jsSpc4cSPWApQSyCfqUE+xc2QidzODGXHHvxY5LmdmsmTnTgOThrXASwXy
PwErxlBqpY5awl4V41h/94ZAUeftjI+k+vtf+7BfsBRIzm/39KLQMtK17KDwUlQDPhQWlopd9cKS
nOGkJTgjM98L5GcS/WXMUlZqqNLNpwLNT+bvVYaqHdBwUs4UwSTXySuWcNohmlPOnLwvdkQCiBVM
yXWUuoWOYyE9oeFa0X+NiJBjtsvL5G5Br3wW2A80pKAbZFgyjYe7Biylfeo7lRbGCA9CaFlGtLA5
4pasKqTdwkHyFSHUNv4+TskwQonpT7+7TDvRNTD1DXw3LvGRhToqSHEf06EbeLxVdhjR8l/gOeNx
juy91RFnx/ihTK+bXqWGcm3WOx30oNP1tSvAIR+dSaLx6Q4khNLSGSdHI6cNzMtMFzJmL36Xeofk
s2iThimFiUAVvnrReeXaru5MrUMvLByFpEcqXuHw/3X8pdDM/kSY9Eoey6v7Kr9EYcaL5e1KLU1h
8bslsZTrYXSE5gfvhEaOC2fj8f25PCX6w/BDNlaJxMRyICYNAYy9MAKjI9xKwc5tiQDd9XK9kazQ
G1jgwxPZMu2u3mpo/AvZ0DeIXzTiizavJLXluExN+c5OIIJwVMA8z7DIbzoaUkXSZciDXhFF8Mwv
4TtCGTnJRqHnE2+vwjGlbrLvstx1TI3a0L+OLe2ThfAkkUbuRG/pfGbZz7DEpIXH9rOJ3K/8w6Hz
U7UaLUHI4/cVwZOvESmT9cLFJVdcijbi/be3FvgzKfo+ifdf9/j9MyoJH+ii8c/OMrnZHmVa8f+d
q4jAB4vzHHRKzT/+ZW3iSvuAX+qtCvbfWhKTLnYoImyJGsLM6GwFf52HJCJQSJ9HRLQq1a09JFe3
f4ftU4tpE/gIX+mpjxLq4LLcjiWTIpgjWEmiea9IJX+nZAyOKqhM5Qx2yLCauEXL0b6IoBNRRZcV
roO/O8t1bSsLfn416L13+XSndh+MDwhg37UF6ylVhboRrQPyKI8eK6PTo3DVC27VOgCL9obIbOHf
LvjFCbDRTllUPtLqjP6fOGr8Pc8fD/PAzK/Kw+6iZEXduZEzoOVf/wDj04rEOHOnN49IdLA/czJP
9hKs6+WeRztX6I7gzxb2vbsJDuLXHkmjukLb71KT4aJfAG/63m4qEEXbyirrPE/GYkH8VpYF4G9k
IOIe0e5dLJvy00LoqnGHz3I6x6PgvJwD/yfvA6X/Vr6Xk98coZAUqX9V+wzL0bt6GZjwMfnfCgMY
0OxpHyz1DfwwtKPnKAN81E3rSU0/Py3zozyNOWZt8tXUJkwqxvUQYLl3uSnskK/wxHJRV8h07ZH9
6OJHBZ5aWB3BZ6koQujK8rc/FdL4q3KRmOwyAUtFw3WiPpmOvFNGLa8lyCWFjybuchmQ0PC/OFPC
4bbonYRXwdWXUxfwAaTz8dTsLXipWlPbPNbQvudeMt8nrw1UIcBd8fkkP5NyOlUW6+olr2izgvjc
ViTgkbBPHhHL6Gi5rJrggJ/lSmxbSOEIHz3e6xSkkVSCB4cCLWlyedkdSLlgbtEm1xcFc1be6JRl
2cOQrcHOSZncraPPB7OJeh1lggtaMKiLe/DM6H/XcVSBS6UUFNKNYFozT1f57BETRsxTQl3IRdos
fKwPCHESSsKjDhXbFJQoX/2vy+PJ5UiWZjBGECC7MGT1fMHTW+BeBN8ryICYk+/Q02/6yF4EmD2j
vOFoK9Ur3Pvx0XVU5Pl9S8sf9uKt32REFC93rYumXTr9Eub4jeoROIP07f+tGjt53F0Cfm3kUGRe
xCsS6YWTNu2UqzG8m0bNkah6nwqWttNwG5gtkXlDtqxSK+5eOZdqvxgXQJOJ5ixoVj1tgktKnMGu
fv7vptBdZ2NKbav00Tcnh9WvvMWT0NIfioWIi0nAUa1fPTG2TGgZySLm1tTG1CKeu6EUZ7kWYGwd
vZKA+bVj1jtqr70NHZETplGNfTyYKmgL0JAVsGQcnffQmPBphOvBSt3qQmV55p0bH8hijvfTrRei
NFoymVJ3+gw9e1C0BDWkEJhs81IqTvLnnn4WUuEQebNiEDu4QvQVApQOzkoAaRKay1HKXjBzJJb0
D74nVCpgZ9JaiBnQBSKETrLqZQQlr4Hm9KcjnpoJ3baNNLkLO6gL1IldLn/AWZW0lFUJ60YqrG2s
aMuVQwK28NXKLrMzElgPnlzEp9tNw/Q+oqsuRegL+yUTp5zGxBYSB2uEg18O+mxu/1tmTyNQF0nw
cEUvE31t8ecWtIMI6HnBRVvrFZmPKnaPez1V0I0RaftZ9p9nNAvolRlKHED7QCT2D+P26rq4Bo4Y
/MXtfoL5c54JMWACZtkkdQBIOizZ963C4pDqGp6l1QJeIjzgRUWkWx01p3/WF8KAyuPwbj79lDES
oM2rbX7YGfqtBPbCSD8P6M0spU2g27PyarUF90nfz6A6K6+TF7UU6JYEKwDviiqmnTPqGWx7FGxG
7/v6PA84w7B2GMz6h4cyG8MDYjGNFfiRlCdVwd5eQcPFQwbyEsq0aoZ0JXD03RsecoDA9S8k6Z4p
ZqMAlsJoeJp0EH/vOY06CrbawRGTOlzzXchba7GOSuTKInevnk760o3UDadYQ7re81xAKJSPMPpt
P7vI29KZGQlTrleCsXT52KvUAC9Dh1lyKSOKL67ahuAPxr9Oyp+/eg/MUdkmoFxMMlJ9qWlHxi77
/rirYa5fzUyDjq0PWYBjF6iJ5icPpxpjkKDSrP45BZX7pziA9110O7RJCL9zAcseVrqZYduqT3Du
OBcfEoI3ewGfhwqiT2HC1vtpZffkRdRw2QLHB/dU8X/UkPs+bndxw45TEZ2PLMNbdpcJwvaffsuj
vlkP8gYV6MYXHcGrjYH7Z4hJYQSa6hyp2WaevoFy9RYdQ6xeIsjcxDfcyeKAQTpmb6w6lKonIKEm
O+xewUXRCdChkbYSH3s0YMb4Lob22xXoe0V773GnwhxNWdxiGGcW6AknW+gERnkeVFjxcwzazBcG
la7Dq2yQtzITZPrUw0+z3/7ehP7uDKoHOVp8HBec+VbRxhvCYr+Ru2LI2n8x6vby4cHNw5WkNKpc
AfxVHYtwgb/c31badXgenC7kHpKTB6i75LuA4tVDmtP2IyEJtdYHbzh8QKSMS9WMHWtWcspHSqj+
N6TPoRRlCC4lOz/2gdF9/GA3iTo0v6aFRboC14UN+ONx5gp4KB7ECGXxnuiS9hTb5gWsJqYZDg9p
Edj+VN6gH5/S1mPdfatSSOof7COJ0+ySzkrxR4AHWGJQWI1cX5dDWrE29i6nspb+eFhJBGJ38izO
vd8uyZBwCH/l982u0UETCZw6waoDXM3gv6HSmLk2pu/ppMCb2EwpHgC9IdFGfdzGp4TNcYBGTQrJ
EidzPGOPfVoryNp7cR101fwmRwL3MBvAM6eLsM41UzrgRizzbsDMubhqcxo7DL/NUPP0GlsvpVgq
Hz7/RHy6dSgTzSoBv2J/IV7a178gutiqNt1LwniMPXtJcBZdxbDxA+94h4RnQ1+6ZZnHpnaRU8xG
L/aP+sM+kQBEkL/C7TBnBAGsWsit4/WQdA6VQHhA0GEycPRK3h06Bd+3ueR51UoCWb/GcBGDgTFW
vgLaIyK+OXOMBweDB8kSkX53400xU38mr8NMYTGxGtdzQ092mDFZWgNMWMYb3ZUK6nNiLHylD1eJ
nUnGojKQghBDXPaXynbKXp5KrF3wmbDaOfdInjAC4KWRQ5jKRROnGhF4ibH2iLjSqL1w8oA9swWi
OM3Ctj+AZiJGi3CiG7KxPcc3yPjJ7QLtECqrbMf3fMl8QyHgLcGoKx7JRnKKLBF5p432/EzeMLUz
Rz3jWVInD+mYny7WJe6Rir7QhYV5egzlwW9l/kDxNKQxdNUbBvD10EtUGMft5E0tz4dnJUEmPkLA
pLmCYTYX9IfgQfvXRVQeJZNFOi/33X9b9vzxiL6vyj5YUVrjrIgzehBCMQWx1f0oXfpcmaGAdDoc
FSqmT0maF/0WTP8hbb5qvACrDUPwd6TWt2kDIfBcPgWDr2FIQxbb684XVJHwDU7/FZtA7t/jf0xV
zQa4bzIeVV+3M8bQFqEQRuC+dMBuxYwVYuPcUcYK5Fb5YSHKP6rC53aKdLC+N4pQR2NOY+4DUjny
cxsAdFrcGDg3Df3nvIRcZ+MkdZcA8sszAptmrwnevPjGBzCbLu6pG8aD0XiLmYwzRqYDBoPXpnCD
eRzrc7LNPa+Cnhme5SOVUp2WEptD7Sa12NYjYSdCLyC1UPe/STrumsPVWv00uZAuPgkeHz10y+0Z
yewa1aFZyt+btrbvpS2DZ6Vk58z5RmafyPVF74Nol95CgJkyJZpxsRjPsbN2hbh/FE+ZW7VMHmqM
bAiyCf8FwDlACZBtjmZaNOYda9jKSsXgTVpAiZs/WFhLPjSebrKv7/EiPfWNcOOxq8VmY6vinJxh
c0ldXThmQSe6s+4GrKP9nLs1QVpvDnW5BEwFlnMrOBOqS9/mdzuQ37tcYup7NHEIv6e3ViiHefUI
tSbp3H215L49879nCYIzVo14zK8yBdU68NisHBqdfTTFmJcn+wU4AmWLhFdkPaKKtmRWB75B6vht
8S28ePj5aVwzX9WgAaChYrQ982bnZlA5vO9pkE7m2Zrs5D+jUw76XV6camlHyieCirV9jnxEVqCd
VsB9MHNRXidXy04VSz4+vrez1Hiw//zYz90wQwEuiym0HmHRxyXr0vBrepwHLpdPZkcRbROAZRSv
wByFHqLQyfGless8u7LU/Cnk9gWCD+6JB1IgIuU3HhFCMOWIUjwiCtX0Q57muUcXGl7h1GHgyipc
uAJxn71gn4FAi3QYPTDoQ+aikDShWMLNSxSD8ArR7Mxt0eXDCuWX6MuTHOpGq5eDgqmbzulRiI75
yfFp6w+AJfuTh+67kz37KHDJcxyCxLj2nnLk2ob5e5LEcDvcg3+/yleAOFAjzAVx1FkEqqkU0I9n
mkJgmKcHQydM5j4yFv/IrvBbWSwWUdaUiHgYv3ehpGsBZa9UJidSBcRIXwZWwoMuapHxeffnP9EA
X99ebBVhDNB1tAxtjaqEomxgQlThRU3lZt74CuJxWerqMD740v5YLTPpuZdHvmxrf/T5xTdUICYv
NYL1hJ4mHYYVmM5BDQ5Jkmh1/76cuizvcwTJilXhywHZClMT0JCOiTco6S+JpJYgJ0zd/8dL22/F
LrSgLtZPwZytF3y+8wdVGkySe2qBBiAazrV2ItXWrcRZiYVvYPMeQuA/b+XC+oSdJG/gYDHP538h
7xh4E//0pFqxxs5TxSJFSyh0jNAaeVhI6yUH52l8TSkFYWe6a6yI59RtwSRpPALtY0nUi00St0y6
RjzJicreImJ88TngMLJB+f4WaazGXEtpWh66JRzmJVFSnTypSDZRpuLPBKmRN3hqSRTUkOSoHVuN
324t7PaObFD8poj8ikefEgtMCbz8vC168mZmvR8SllSkS3C1+BcOos+CpOp7/VEtFfnxnF3n5LSe
aWhZTIku4vxO/kdp6MADRj0HThQZojjTpqukL7TaWd7tlRIZqGg2quA5MysQj0X5Kh9IyHhhtxpZ
5JB44RrxbVNo19x/dqrqAWwKPfNAOt3ZpM7ElmWnN40Vg03NRkD/YMECs4dRLosPv5W2ogEoxImu
qtwPMzgV/DQj6JOrEbJu4ZtjmPcK1n8/iePebyw8wLguT4sz2Z4iVJ8cww2+V+AlHn7UTzADpg3m
zR90EoLX4At5VfWYqPK/tBzGgs77VHJ70JumKzbvHyIrvp+aV+znXnSU2uXrEPQ4J7wmPB3OEwdc
HRkNJmOsYdtr4f2TGYhRZvJwOxlR/72PPNKRnyd2xN+5rV5lc/dqoGsNABVhU/IO1wtvd64mdT39
LJUFYzUQPrb99EoZ2N4DYVe4yqhai1mGwHQ8ivy7xw9iOR2AMb22lnzFbZN6AUpDvKxeRoZHa8pL
toC0w5EiNp+KRkK0MTfmpB7QDZ9s5onmxK0HhxnbMpDdtkVPKMjlUjUHUX5xAcwZfJErJ46RIYVv
Vin0SHxb3y7Q1rA2e53K8xR1zWzJXFQoR9pIVI/YIgmlexEMk+bzSiWOY4JtgG6MKndMlrkMrpJe
tSAktYcK84+kVcwXHvCg1X9bhyhplhwR44K2vuc//JwqeCOcxrF77iMhfVAkxyl0na3oJINdzp6p
K6ia4fOBQMtXLGUmHhh+XffWhMYHXhvrU9+6+pssy42Yv5h8lsQnGTLFRJX6mvWp/Jc0zD2tc3MG
C+LnZk7K4ApFrlNQIDS49kThlZ8ju4eafQSeTgU5wlilC71XoYCDAmqANldE2F6B+jb6PHO6fYr9
81y3hClNCwEaSPmG1OQDfrMwf2u/Dha9QRQve4jkXgIp3LAsQ1cX3uocXI50yqU72iL04UkTEuzf
NzgwoHIN+F33oVW6k3aID/SfDvPWbhyoAhuhEpBajxFnNx5cdunzuEawKo0uON2YFJp3AQclmPVL
TB6Jq8DKwFCyhfKwjU/vSKAjMtj2oxerXEzPwt6GHQkc1mnhTuBbc7S3/xxsIFyhu7jwYYWFnH9Y
NO3pS21gVOjioGH/MizQ+dm9uvM7ODVSmXXgDxr6ljljCp5EphiPZ9kvCJoSZjmo12Al8oW7zRuz
MyeEnBEJs85NCSAWYU1Lm2YJ0yb2WX+7QzPr4kUwMxq6bfUMWZHTeCEHzbhytQu86LWfBfGse0fa
BVDHs/9+WbkoAEjhE4ElijRrUPUqDWE50xtGeXHYc5FOzfX7tlpKIkRzL8+2LV0Wcdau+C0ki/iX
gJ2oxN9IkSU9WSvueSnLH5TRPFowesSwkpyEJAZzzoY9sWjoVjZmd8K4SjNCautOPQ/Pxp+/fiVf
HINTdH6SOw2nq/2HNv3XthD9/T5gPplPenTczLa6tqJ3x+2MrdJdAKSfniYASiw6SaHx5lPsEYt+
yE2p82d6cWCLHSZ+tEarc7DPOSEQ32HlixqxqUdHkD4vv+7wKi/agSxkGQGp07L30iFoyaOSP9Jh
7lIqBjn26h9n9qxkfGV5yo9WbWmZdxOXLjFVs/Ldf1LWuSJ8VK/xgRPO4jqvKrmfVBApHcV2N6r8
FLr1pNtQO/zD5PY72QcRIDzhXU2L5bY1nYXEVCwSftGQGS6Hz4Q9z1+9YjVI4NXR8nx60ekwj6nw
+x2P00QMk4DWa586mnhlgCTrBr5+VBddOQlWLDWJ6srm4ajttjQJSLQAmmykThqVaTSJrfRiBt4+
3Y3qEEWpxi9IRqYYEAV4RSZCPrfY2Y4b6allIH++YwsxWl2CXbBNnOAiCLnu8Q9OTC3q5nKEe2+h
iyEoDh48iCw7BPLQSgXmvNegIz5EwZZk+D5WpcP6nY3EKix0Wa5WNq/6D9gkZtTYvQXsnnIKw825
qiPXC61HhubC+Wo33qx+pZ73FKujOFtjw2RGnODBMw+DQ8w+s3yzJQTmVIOTRs0OY7I/0n7v5nRB
YsO4f3XPibf1Cz2KLwX0sOoOr6jJ0ABJ5s7TaUa2K3XRqgxDSNEfyPZk5j1eDCK/Gwwuczv9qNI6
MK+aFu5rucCY+uy55soL5LjsKtsFGqrYlwtBT797VYB7B/7Tiwey6oWLtdU0VPF97V9jRLsvy6tX
2px1EJEsChgVOqSZPju/QWlBzWmYsK4CdHqgS++Tl6tMmD+raG1zUbi2iCqKs+64kqpZl90xACYM
guLmg9vTbsEbYTh/SpOFpTR1qUtbHKGg69uplyLDK69/V/2PHM/pu7ZZLhZAlqqoA/SyS01o2/9w
7sM+TVrGkg9teOq/PTs/hqqyf6q3uEoFv+FiG2CrZowpBPFhTYyArivV/MWC71O/6O1Nq7W7yrVr
Ubt3TJ7b7DUm+7upkalRdOSV68zpy5UAAsL8ctn4mNl/PLpbZqNIQfeshfDQ6Z/Y+MlLiWEpl+VG
x3xBZo+BLSurL6O5lHycVFuUDyn0ZFL4wx9qbv3hyi0BXaG1hb2vikx98pPenLoTHC9+xYBmH+JX
jX5Hk8gT3S92vlxt0iX2O3xhl8f4J8nUmIxsUdfN00ei2u4eFhNgEXjW4sRoBaI/gVPnMzRdqbFR
y8G0huCtm1kuAX6lD5U3vlMjhLG2WPotZ8rPm7Pjv5AHERT8tm2seswq/th6Z6M5eU4FVtXwihbQ
S/c0LRe+xjvLO/YXbhJ6oHb2BEv3a+kUzwJPO/be97gwrpNBcDkoCxYRMLmY+jlbsD+MfvkQhnJY
3vR3zPKTkq6WT8Dn5IbaqP/hiwLgFGaBWrtH6+BLUhYelDHXFYWJuiuAg6uWj18hh9n4gmfN0p/l
4ndjQAWTgvLZChwtSNvdBiHMHTSmj1KVvjHgBfxFtVuxlg+dsDrG+2ZEvUWtHd7M9XKHIAOnBw09
3IuWfCKUGipjCj1a1zzkqH8jIbh2e7D2xAI/NWXSwdBHLTVrRnwXKVdk3AlQlPhx65V0CmB+fE7X
lvjoTh+coluncyfV2AzKNoXP+FhY2Z0pA0WxUjWjioLejLmOCbG9ksUMErkvM/yvLzLSoDf59xA6
QVyhpajc0s2jiTH4aJu+DQVw5bZ6q8ImC+M1M1XfqzO5U8Fo7sVcdgT3SYdXx8fvpSPiQcWwQ+6V
t1iT9Mv/rbHjEQQjBLdAUlbf0NlWQKd/MpGkuQys3iX0sbRUqpPfqRvVCzQnkV2pt3NY9WWCW6cc
mfiWcyzhzxp9gJRVxZYl4Knwsk1lOLPxFsA2imJymeAQ0qkKopKCzMphb7O9FneSDRxRJV/egi70
zbDkK+WA+zRIxG+0II1wGSbuD5dTGpekPG0B5SwqdvC9lP2lXjpmSTV1w6dQgyXjASYgCqqMLafG
8LaCC+pLWpf5Wm4TUxRNtXblQ05zblj3ZIK8OnS+M0jZsA8577S30PEttl6YRwgIHWYWb3j0sD4i
28cGgC10KoHCDtSLrVyIfFSzoGTUihQhgkl2Hjvc04tqnlvEAsBqFOftPFcIUg4ZPt1b3Gb99+VK
mgE3HkhXmFfG6cg4XrOSfTBD/eJAZoN9Bk7wJZcZl31PbdIRKtoBAM0bbRf5PSYBfKYPTzru6+0I
5ndmkHhXzUPEFTw3iZOO4YBBQ8J6L3WBsXpZ6LikxoHDpr6AKEV5LX2yAADxkPYKGix24svjEPNK
+jmoh5Lvm5wpREBjTEHXU7aR8MyKRYziy58NfiDiVuIZ+QRHlP2opb2CR/S5N23pbRJMLqVhW0yA
P72Ie4k8Zxd9/Tca7P9UTToBYw9Ku1v5bO8t2sl14pmlTWR17AncvzCGvXUZcXvF0vGVcyZtO7Wk
oh/O0pmBnX4zY9hs7AwMO3fCRwkyNJoqLRVH4wZuJ+LamflabOZtmOSvrJa3l+0I8USC5Nyr9Vgm
tdMviLNL5fwahcflZO6I6ieVdNGP1wlcmP43W0I36I0QqTjDDMSdiVRSpIL816acknBQIU6YbCzF
tOQbc0XRQpC+DwMz1u0RjoYoTulu3Fus6hdNQH/Q6FWEWvYxLoVBtZrDcdst4YefWIuFtSq/m9N0
vYvQg5uFo0EZHlRuRvWIRxdhm4VFWB3KLbLViERFgnZNislK9B1Il50Wmjna+FmQ4wQTcvBIaqFa
ORTcQxlbF2xrB5J6WaRx77qw+/VvTcEhVOC8gk1lnWP25h1hmtFJAoxPpwn7zmI4utReCAW4rEZ9
vhppZakIc6S53YFH5B4yWhnCkd6akt/+w+SoFkKNYqtcxBRz0MJOsB0vyuSa9kugPIE8XcqbDtzn
dVCuAGUgn12AzDp4NvantQS1uT3Wh2wgIqSCBzZG+pLrluWtNIzZB28jW7T+VDQH1V2a2q/HyaFq
i2jDZXoP4lwFQjAwigPQAGxj31015BEicZBxJQyYMtylZkWnnoAYvhLmhh/PsaXRawqSqp2jGQTt
AQfhHo9YY2IbwS/8Anvr725z+G7LZVMRcUNpctqmlGuyvsTZIuuLNj3smqjTTCcdzH8gVq/TXC7j
lzNABUCt7KFV3KhyoLVPylLMzj9OJzNPy40tWHcqZXtxaWkUtBRE+9JJbiuNu7o6ojBhz7NOmDFd
4fMivagYi4vRCuzmPfxaPdPo4K0pRAW51crkxhu5KZSfNnPweicqimPsstDIz74YYa+3OWjGcmIy
/JYHcUMZmcyp22I9Vyv9diajArN5MmogeKa4qFdHVZCB8801zBZ6t+Y07xlf+U7mwuTJrzMWbdqS
w17JLHn0MBxRIfEmpi0BZBNO3be6vkHvdx93FDVKCtEX/eNTyVd4c6GrMnw+hNXZWxmzS8EMHtPp
QnZBwoN6jjFN0A7739/s1PO+yIQqRDCYRmLZ+A3tPlAanASJTUFWYCgG0PWyBGTKGv1xp6lIcBnT
ityDwXnf8r6FuB1uUZgFWj33BJxFpu1KWPs3pIvMy06BDMmySlfcTGjWehuPoo3yFmt98ZirDn3L
KmNkkFGPYDoEN9Vk/dZcWTYr6niDugC6Jbvt59AKMea3wo4RZCkqkjUaAegyV3nwJfnofWPSPz3i
qldDpSWo4Qv7/vMMLaamXYU3DWwgeLvBGLkpAapWLDED94IgsS7cTlHGWRLleJ/fbF8jzd/twpKI
BDlCwkAmXVLjzN4KjnR+iqclzp7y0DJmvDSTc0B17xPTA6zis6q0Vl3imSoaRGIo+cLUQBzbuu1N
f5T/mruaHcMfXfhMLB6Hb4Gv3g3HB8s16qrhS89IpEJNpe5bB00Ctf7Ge4wvQPwqz8lbk/ZaluGa
GFnh3xnYMw5ExyeujP9m2gpjVeUvBAnUyRzEC3EBB6gF693tcuCZ4v+3RU0aIqA6qSh05dikkHw/
5uvio7F73mM5zrw8zs3oND0XiM6ZB79vGxLeeXw4H+IiMY00s6NtLfHzuYtXg7X8iJ7fUe/mJSQ3
cCvb77pxbMM7JR8zruSP+HB4igzH7yM7oe88Nso5EN10u9xQKdL97sEfCrs+BIlehvxsPeABGFIU
Cmyk8xPCqQ9msw3hE55e453t4X5wpcnUQUVi3ac0RmnUF54mOkPwkc8zf/TUTeP3EMuYW7FROClK
/H0bYpQA9n1irr6BhiKlARy0AHSKXHbu8RsG80R4XfqHJ6En3TF3DG4+vfrH1tjfov/aJsl5WlMb
RjnlsEn1AlVU+m0ezxX0LMpajKgXmWnkAzG4rXv0Iony91ztEi2d+B7+p+CHVa2RaB+UthFH3ZrM
xlkRlwGpwJxlekkvn0KtswCBmcV+hxUylnO3lFvratnc0yuk1uzzQq7GAuFgkO1d6Lj/Iat5Fzsd
J6tRzUefoJhx5IgjADkcXvj6TFSoJ+5teBLA/rcddklKTPEdELSp6tyt9C1xHNQtOHUHF+1QrG7C
bfi06pm2W7FlPm0VJbpcI7Q3SgKH89K8PJ2AqkoIaxSb0N49JZGRdw5CJpNgf0ABFLC2vXWy5cOh
QnlEI0RnLNczBxFGkFWyAjKZX6/Li3akl4TtD12ptERz9I1l77ORVHYN5TfWQTyQHUs3kDKcqLgY
i3l3hzKAefOuSx5JrvvQmJ+RWoJRQGB0/diNqLtcoLj7HFNd/BrfJ1TarirNIij+iDJdmGSIX2QD
hucVxAIsordsbMSYAwhBTdK8n1OLf7sO1evYz9jjwIq9Vtb90bdh6QIXfbIDfKDO3QkmwATgO0QL
HKGshH4ttDvgR2hMf8QYC6akKnq+dhAjIoHHzXbnBZs6J1GVQHxX3NSijN6O/NcXfLaw7XKuS6MM
N2HoW4Yglt4yqo+Dbmjs8hdOVI7oGhcRXm5N7hspRaJkF4PTDikhSifJGGVRu6jQYqUMwcQ1kGXD
5gHJVAfuj/pVqnBh8DkeQh3qKdrg//QCIgftbivWGsVdnY0q0NR0gz4E0Kh2PH0HorhuK3z7jSYV
2qsH7J3ezKLwiXHgPq0t029T5nQdoFbdzRNLDLR9ugieXvoww4/3pM1bMMFWrZ4Q/GFw2uCpWoK+
1wS2z2jPbLucG0N3b9ksXCjU9uZ8VCS3EgYpi6VKJApRyg91/AQW3/D5TUrCermscgtG2XpIvGG4
qo1WYH+32yNbmedmxQD+0C3GOtY7Z0UYOJIrMtMxH6yUCcpQs35TXwo9gvD+N9jwrjVNQ8z2nmKq
EXGzVO9n4+NO/FhD7bOL93ywTeRhb574pq/6t2AediDeuii8LLCweaDhCRSLey+NqO+sEJ9rqklF
E00rJGcgIFidumV9eBUw7Q/UvA671+l+yS2VyfPr3/RrSPZ4PO1UepPY85lBBs2mN4QBob8RQi8H
k6rShpIJ9mFIGLBVx+wwxcP2ipplbeRJqTS4ycTMsgRpDXCI/T/3Pgd+Hj5Lw7vW++8sZCTpjUjB
Pj7hMJmS0CFwwiQS9JtsrgbQizk0vwQWb7z/Jy5JAC02DH666Jl05DBPGzwCEKjAJqpCatznFbte
bLOlIhx5ttpw97GNRfLN4ZqdTDoJBAa4lrGOWBZxuQry/RKqalc/mHn1GffWnUaDIghaqzbAjoo2
AvD/mjU3FG5ITu/nLjui0MgVuQxgBzX7rn6q1Wzqaz2CS9GhaBHjljrlwLNCtE2XRv3ZxS3idjGH
HfhK6SsSVw9iuQC5zP7EC5Eknlc6btnwkYmND/RCewrOC+9DqM80QSvjGYC20qeFNXddda/UFVsV
NanLQo7Spy1kvGFwH5HSHWHo2w+WRyh9FcTlt/+zysXm5l4h9qt0V5s9dbwWkPytthoELUFL7md0
J54dPz74cpolelYQXcndhLEBE1yZJvsQMIwYWZq+o2XHM4J2uWcicccv4zXCJqhmDVPn2oKN/R/V
olCm1UngSYwsWbIEkM8iZsuQfnR1OCCAndi+uidGMZIv9Wg2MRPjRfd1msVtri1iz8vNzq8D0SsX
Qo2y64L060AKWOU1XOCbsDbaA0qzeGHDeczjF/Kc0QiYgaE4chu5D9K/ZI2Xw9Axexow+ZQusX0y
CXUxawMhR3ajvRAt/JJFIxofTWGP8AKxoxUjm7y9kB5B6NEG1xDcjDvHk/Ovuu79gBZknv+0txQ/
W1ORFkuBs3QkgldN28N213+b1z3itpoLe4Vw56JLVHhVUbtBcfqmhMyZ/ecZhPS97eiTlgMhAPuk
uYkqSxO9QwtPKtiySFSGQSg1yp9HwXadvwt5x3AYDksVnWXhEaVa4VCHkrJY2rp/kQP2WJN+nOmD
yZc7B/iF4geOZBoRyZHGMXmQZVkLYYD34aS8I3PUVuUuGPKELR4tteSRP29l3BLzckPmqXbsBi2q
qI2yeCBhIY/rGVejxN73I3LmOubcGcvf5LhDfc39M6lSRdchWFZN3NGAPwrAZoZkmBDfkVR9Lw2t
D6/pfeSv2OFMLhrK/3gqZTjvey8AT3VeQaL1G+LQUG2vwYS6hHb9ZrBfwDlWEKR51bJdgJhIZZ0W
QFMRPlJIVLg+/U4gYHfK9NIl9fYNfZP2tPArs1tlBwb5ZY5dt4p8UXdafvMVkFgXd3YzztzymiFH
xC+rZr/PRoLXaJSUFY+SYlTHIGbYeUqjTUny78vBWqLt+W6BcJ7s6WzY3P/NxPpWnUyPXPbN9xN6
P2FdgN4tceIql50muWzWqigxD6WLwISZvB70FlSF0S6/tKP9Asp/jVSoWbQVghB+3tjBYarB5Tfn
wKaq/g6aPk7K27nm+Zs2xNybPOvHxqMZG6VzGsCcfKbW+Uqkm1kr0ip1C5WkKPGZMX/YoeWItPxe
83XE/iQKZPdf1OeoJ+bpovwibkcpaD/6+UNzKVMbywxk2UQrWN3C0Fjfh2Roo7CxuyMoxRpPrI1B
0ejORcLGp0HNmo4sTHcb/AzVaSxa1XXz00bVmVrc0jEIuHjhVITcd98gyYYBVQYPMJ7dCmfdMB5g
tvDUZbKQnKhD/SMi6xiWLXyfOTVZgCGLNlXkjZOpxj5A+Gmj0jX7QaL9EKrx3NWLyo2UyCwzW6fN
q3oOrCqO//wnHxxuhRvULSMrjkrGI/0vGNTTwW+mFE8mqAjwU2hkmoKZmi0jkhx+hClt+ToVkz+t
QoyQYk59w4RolXgbI8QWdDxALpJDez5TcOcXtvST/2Vc6EsTKvVUc/GwqQtur1yQRnLzvVzatIM8
NeWXZV/qmrGw43ibQXj2yQZuT6/Tb8DL8niM0iKzagjmraZHsuLGTH879W6rLY/ogTrUEmFRjsLo
be2pXE17e2X3+fe7C1VscVM2wMzt/bJHWMbzJk7DHD4DhN8uq0ACvjX+7XYS4dD+hq1DYVLlaOZQ
KUo5wOutm5ctODI5pObtPaeiFjmQVzrL0PFLwvzBDBWuvhonZ/u7vacXFpod0CrCDy87eMGnMcAr
WHwwB7/yRxjlCOxe70+8Cn9URrYyWVB/ZqYZEyXR6iPQq/sleCRF1tysUxV3ZO8GGBJow6tAuQqd
L1P2gorUBHvWkDs6ADPJBNnohK0SGL5FsKNMyZ2zOGMxuHyn6L/NvSlu/sqvbiHdlYIT2EgI2RBQ
AHnXSP4XFkhjGVu+xmhxV/zw9h2vWii1vwYaNVWmX7CS/woKqAdEW4c7pP1qd4odbgCCF3hpYNbU
fMM5aubgxC/9gI+VMIYN9zdXa3vUaJZyfiReSD22yyhDjjGZ1sQLkj1PHeRKlkYE7wHzP7phHD7r
Gf02R32vqI+DkPNJ2/wuaF/bdSbJaqS9/s8k+JCYb9e3M6hyggCIyVXIyOjulScKKDearn7zv9gy
RcdwK9Os4L9vkJ4KKMdawGZROCpTnWforuLSZ0ioILw94b0AzVqRmp4DFv+CDGvaKolBK5Z02Wj7
g4zt+ls7xAEVBrkQoKGWu4wGwXpdhlY5LkJFBXBOy/l+kH2Tck77LyD38EO3ACKTl1B6xPEeVgSw
ncheQrEYx2QqpiE2NBu81Q5zoUITwhq3T4XTjUwlpBmHPxVTbOLz4nmj3eAfK4z22Lk21Z+RIwaV
4VomW7k9YX65HDptjDhRHWcVeAWddZ2eaeJtzffTGwy+8wcxI/tFduOUcbXdBQtvJDO9GHX6qTgi
dE3lOwqvtAqZNWzi6pXvGlVpCF3gNFIYIuBo67KayV6sOj098xSs4aR8c2IEqmHDNorXjXydoGOq
S7FipdzlvSJ4GWdM/bs/H9tV7VJHnP5CfJnQ9BU+Y2xU4IQ8yNE1kIBPevo31qFSsD6JJeXWD9su
mrzqZB15sUZkYM12F2I0Tj7LSNE8kxYvtFa/xoun6orWFRvxy0OFFgNV/ph/47v7Ku22vC+67Zu/
Oq3LUrhSjAXVMAJucBxCFGqlpj75T1Llbi7NhSMBmqtYyfq1yQc8Jbi/5bo4j4gkIsSxjt1GZVjf
fGnSBQatQJ+fz/bPLk46/XNAtGhOI5f1st//UjT4EOyicuxjnFCgYHbrNqDb6VFVMMWeLKFDoHeI
gcufIsDknbU/9M1UAl+IhrludPgYptOcXrZ2ztMoNj3jNwfHG+LxIjdXGTix4ObCk9KMZynQQ98l
1vcw8BUCs3TDbv19hZABkTo5TicFjmLGW9F3CaEw7zk5yC6ZR5ExzH7JPgPfVyK1TAuutyhkCf1x
jesSMMHls8BAF/GEoxNF5xNiAtLYqwp/tF9sMLu+mRnZM2wpwHOWTq/49pkcaem8qmI96ZZwXXs8
afURP/d2ZPy18VtMe1+EbJXq97jhDmmgiQp/ydzMtHO97rww2PfrD2IAm5S6G6UCEYIkxISfIV6a
6CF2KDtIZP4QvetAMFT68foGqFY/VmX0QDxRGX9wKlUNgJQKvQM0eII5ocDRkyO4y4rSTpp5nRV3
xiF1DGy38hs2FwhfQM7i80A3OR64h1Pb2qiKsg2bAtB7sgXXBXqMyAsNtFISEO454kfBwlCZsROQ
/gaGjaJbODxZApBcgUV8xeu9I/XQmbooWzx86oAmfXxedpg8M4JT1r44Kj3Ze0nJqmToh/QXJ4Vz
JTJWKF2HuzMBPnXHJfHTyAnHehyY+QVy0iH+WBnGtGFDlo0riKmQboJfU6NiQXfkFHoe3hL5NoTm
FBEkMbUX6m+UwtAz8eVtNrCrcr5OaQPIR4W/uw02A3qSNNCJWF6nokL9lEQoRHowv5lwzsLJC/wv
Owk5kLBWiwurPAfg0RaY6gZHzEOhdQ35ZsKqZ7e/uuFUxUgwtKTv1Kg70grMvEkT+q9n4JuMXYHU
BbvmAVtFEkUlvfqpxCCUfrJRKyPNut5+THjM91ko/RTVtBBZrogNoD5HbMQHJulRF3j0p4sWeTuj
QajAviIGl4A9GJzDMWYh0hwUVdx/cJX7LC9HnGNOdO5zblyWhfd8Vm7LR4gIP/AjzMFzDCwBLiRi
sLHXzM/kuzH7VW9NGeHiXZTtlUzF2o2+AwrAsEG4VT+guAqHIrfU+B5dNUP9ZGrcrACVA9Uvhw/M
d0yBh6Cl4umqdO7+UVev0ybRKL+FBS8rXaRr11hhJCznhsTJ05043yhPptFWbUddHYP77R5StgK9
6O8F3ZlZBjiNeo07dfNyaR+10Eyyf+z2Z9FsqUuCTMx8G62A1Vs8MbEncpbipYPqhTx9DPVsJLr7
1wKQqIB3xgNzb+oCsQwYhKLrRidwFfzUHTVU4iEqiXyxHCd96+hDbMtTH5aOX/WHypw/tHqYCuyT
DJusLwCM/noDl+ZLbYnFEWLo9Dyxj8sigNWYhB8mlRS7FsjkX7lHBdSqrZCyl/UzOue7t5EVu/cX
/3zRsFee3kEYpsM0GgGOj1+eNrBt48sHJBJ5O2z1PR0FPkl9RMf89dcGnNTXQHjQrDhm2bqrr+Lt
fGQ9g7kFkUdFVGTCaYYCEmAcORh6GB3zxF78FcCVpQWHnhWCPauXO2Njfm96bozBSH1M7IB3Loui
kVcwS5TuMfu5TGSILoGG1fmhl9P8xEMVFAVKA/Dn7ulqbF1uQLKSuMqoQImi2jDS2XTSXcNdMKLe
IVmS20uKkBeTGcdE8ZxZ+3EEyiqKZnRtMV63GyWIWWlCUXgr0DWWTiInPTWbeHvEdVufAfjG9SsH
6QwKzHjNt/JjsQ956TamGPMRyC0eqR/sADnVPVeBiC1vU8UQrZMS6bt9TcZsYRf769KmptGIakUu
ziY9MV31xtQiozGr73gX328dmXISelVJnLfvqnb2jw5f2Nj0zLtXnxZGrLGXubiqNO0tZY98/WUc
rfuutguFIpX+wvEoBNdyPAf35YmBAMq9SnTN6o5cx2JUiWYJg7hmzzxp601eFrpRBnLhBjFFORwe
XzFsMxPrRw6NwM2+mguNaCb76c5nbKvRlnMTaHll6BylfiiBFnZJR+OxlpQacs9m2sSbwvFUROnH
68Xc4VM8Li5Q1d3/Vind2JsPN7WMeEcoGAAOoS5GFuNpt2c+lXs4OOf/w04Cpk7rwsRMW1dgoV0r
QHCZj5+bQUTJ+JVX0pw3Y4eBI/tLD2KqjJRQmuNp2dFsdbOx2YT3QLfXDlzRF7N/UsBIfCAeSb3X
RwkPzRCMF4QAxNTVXXiEwz3ddxSSKsudMkh6/A+fDoZTAVf0PeZJ1KCGN3Zhqsav3cGiLj2KFRkX
oPwUFidWOmP2stj6U2Y6o7rYTPe4detRgyYM5KVGUR9j313vP4ohSwG9bap/KqW4z/ddjKp32Qvp
jxeL2KeISFJTzMTsVyMWR0km5k/Xc8o9Lfe+OewjK5pO5iWSagAPVclTFKEin9C6yazOBGcQkeSF
vLNQwSMNmxIEZluNHsj4Jd5LEI80jX+KCvx4Y125MktO6Ez46WDNMb7h9lGWRJQOYdX1/KBTfmdI
etZcRHolofBpGR4HpyCHtr/YtWFPTn0F5+s4Q3o69B6b2tVhTO3Cd78gqvX9lt0N0BqjJ2ATLmHT
0ZtGr0siU7a5xjrikp7b5XnV9MM3wb9lNbeB5Y5aL4BsqCPNzeAgG/BbaMJOvMnkdyn7BuuPCqcf
2DSmMiuwSvJ/7R/61B7Ha2jjAq4tH1IcF3ijX0wMirlNXL7mfzmu8lscE1AKEHTQZXTlUrOTdJKJ
v0dCo4J7LZLRY8TE4VazvjIM+Gs8643KmNkWQV4mwfF+0kTwrWWN6632/cM8Ok5k/biYRt+HwqD1
ZgTbl5LBd2OeXogDS2OocUkiXy64fA6DjRTXOakdKLvClPgMwXDG0X1Ik5NfB9Iyalx9WnFuK0xb
aZSo0coR6t1gJi2Y1/Z4rWaAyvUnyBWJpk4sDNmAvhacWHrSvZ+4wF82bAu4A81+0XRc+ruCfDT0
KAVqrw9WJuzJ+DWKu9Gin7vv+IcLsarcp9QtutSMx1yZ/+qEGAYnfmM0yljD0zQVwlxQnttfFALQ
Bcuwvq1BXDx8MXfWM+HlFiKfoipj+5C/hbM2iJBP9MpmIwn+yk3UY2n9zzCHasvIVruY/l0MJwau
AfQFVWacPolb3VcK7HdsjaySNb+Fg97c8m8djQUtI7SA/fqlETz5/Dr2PyI/qKk33nn9s++5kK3R
CoDHHZ0wmFDiTZZBuBShD+GnHEJfLxba8K3OJy1WWmVh5Zo+GDwULugtAIP4bcRMKgq3TPex6QIJ
kZeo3hBMruLQaKFFlxG4W/asojA7L4fxrYqTWkWFisZH6JeRMVhx5gtUoEGqDRlaz+zXDbSIhPEl
B9w2T124pV1NIwOKPiMgk1f+eDqr9i6S4aLe/96RWiOJPSft9KETnjie/20BlOmlBKtkWnXybEZU
Wp2RIlN6+/jCDPBEJekzyB6G2sQyJX1c3uVX6vSCXtuX8+UxbZsgJZCv+4k/nqS7C6qn2/JG1O80
blW9ZDRhGXzPDQFFVyFC3aLHBYBg0i3OgIBcmS3y7fRnlbovhyqCGzZwO509zHNWWUYf6SoCT8lz
+0aWhN/UyYEvUxCZQNYK3qKfsLQ076I1KFqWa5zZMomDYX1EXhsNqyKRKVb1DTOu9gTrFdxrok0R
Eq6HBhGSvYOfVd3aaGnmqgrCicIdwZjmn5J6fUZqzKJN6QgnDmxqeiPpNvT/tOCRCPqPjEC4CNRN
hurIVuFz7j/8LIPctNF/OU06wrYLrJzRzAaZCkc9SkG9aTsyikBWTIUpjavSZuutuRUceM7PAsb3
L8xJSsiylV5j+MsY01h2bZVzdrI5EejyGsGLtE7SnTxx43buXRfYHZ3rtE1GVmaQUGR6SGgpZbCT
RL6VH2ucCwXXK7jlPRMoEb4P98+GuVBiqwUQSaoWRzJviXQqdlojt/dtbRHGoeLWZk5XbrRrH6/q
UpNWfXVjl2u+O/GwThrfYX6/q7fUnYWhKWn7igNgYfHF6yixRJtGJ5JcQIXTyBtmnNROhVsGFGXW
eJoIJldpJstot7EsdPW7tSmblMh2rMOTHyMQJbryaE09vGr//B8SGnY+k5AMayey5F7Mq/9Kq9qR
j/2ejD1jR4atEmeRfXYhwCsmF+7kVfRmdyAreg7vQbREydEqmYVPvpFz3HLeYW4JpwfTe0MDx8ND
/etK2m9hYoVCYNZ+XFDaqi9VJZ2L59TJtCDlTERl8hKM/XF31P5zYSuHOmm8QCnPxvnfYrw1anU/
uf0InGcyuR0350w3/Pat8EyHZTIV7g9pxzkgSzXl8cABWNuDWtqN8xdHHrjWuXrS+SHZyP+ZWDCd
4IYqLB6qKwv7XDm1aZ6YlTRj1akSKOFJMbzxW11acWAMeoczc/xC1RA5RFwgg3ZxnbATV7aoJSp6
/5sZriBElUAx2Or0MuTGp7ORSmkaxB/SksW/hqvfRfbHq5P6VL+530iwkZK4nrz9MTuRW9DPtRpn
xpZEb9iMwbGc/u1EKsP29vVh1TXw9wYaleFsxH/tX7BPDdgYEPvTOTmjH14wZ+7tEz5oywKUqO8h
3rUpBavJpN9bNldOYpKWMAxQD7EY0G3ovry8xdBL2OkraBqbPECpzRQGf0D76I4qvt9xjPoIH9q5
tDrZxcy5bTsew4o6vAN9CEdoMvyPfbKKS/WlgaC/QEx9TfX0/S+HoIxdlPl0LGAQjlpWFwUR9L0i
x6IoVGYIuLaWKQI4Ax+gtDiorHPW2ouPfBp7q21Qudy3TTRpUs8nVrXt0NV1Fqj6qJHtdVaOflzy
mHk6L11BS0uUhxppq3/1LhuvT3SPIK6NRVm1z3LfGPIz+hDoKztfvrLsMiTSizxr3xcQfE8J43V7
IKMTQ358JYfVnUTfVggn7h5ncLuWjT7Vlip2SmdVXQdKc0kIjHP5oKEogNtvvgELvRgsRpiHdIRf
ByVQ5z6oe3ogtZHi5d0oGMB9C50AqwPAWNRPE+QVhxSy+7xhcC2EgRc2KMm9KDK9WgmYVavzIEOS
BYZyUoPH04vvMJEj12ep0ktix7MsMSksstBuOPhh5/TR3KAKMZ5wblZSr7YaSSZP3LCkkycCZFsb
9+be72/BmbgETgBh7BFGIIks6Ywt8/U43f3OZ99NTlNJkV2K1JgOVVil6tDyJhlZyjo8x+ce7wJt
GPZ1UgfGyU7KK1RjZSSU2aJtCDiU4WKhQKhVu8ZmEyURzfE24b3unx/QsPjzl1cYqLkqf04h5pTU
HTd8A+i9Cl8ExYClaKNvs8g56fT6AlTt0lha3oMzZ9JDNA5Bd3JrQRyDqthwihVSna5VTaRYq7dk
aaDAY0fPDmTgt2Oc5g0cAMPrIbXpVKgCZIYUplxH65Th7FOt5cwd2K018w7VS/tY3D6gsqll8nAe
wRfSCwZ5QIRV+2pMjCBSFdhT/slTeDpd95CoXx+69gZ3savjDN9F79juoQnchqN9AXqcyaGOfkSq
AXmP30ouikHOCpCbpUsWr0Mp0EoFiBIX+0QWsiW+oW6LBxlo41DutkB1Ey+g2m1iCiIPwjBBAjYD
wMe9Ng+TX+fTuaVCPOgPsZPIET42ecM5USLj98xTXK4itj9cqHWGz4w08V2nMPPK+M9IorJ+vlXV
HYtT7tC3WkaT0CF0Jfc5rWQqYt9pipBoIelpyGjX1Q3RC7m5Wq7HullLAdiWaCYxYU/CxTVjYU5w
x3ofGLGZ+0+cx7pZzRSZUNynXaK9bmArHLlUtHdLWb93AuTW/iDag3/joVJdcZ7+QM/5AZjYhBSb
zEiljZdPC4RzjoxHEzFULMBW4TcdNmwSwsfQ2Lozo7HgWJA5IV3zOf2Gg9rq1Uf5EjF5Qzkk0U40
1kC2jG55zipvkKU7IJ/AJYpL5sfFGJEwK2QEEI3Qu0J0BdMZWS8ycMnnYVwtNHqp/ndYaAimp6tx
geQCUsCHX2MqbNFxmU0YK70uR5Vh0RmPDhBGqonTRekO6VmoORzdDzMLcyClPiiZl1ed04ysDm8n
2RF+KlA1xoQXosHj6DilB5BMRDgXtPUPeR6L45qn2AHrglwu2vqfqkhp0IhoFvzvfg1grw1ecMqU
JaqGaM8pZMpcgR3kyh6E73Dw1bMdJspBX/W47YGnkT8ZKsJKFUyDg4tz69Om0m+qYdlHfUT8V+83
wPEs6WghIX01WBahRIZZZqPC/hn9woOuwevIZmgJICiTt2XxUDH4N1LvjcMU9okiQTllOFnm/wym
GXTyzZmvAG4YphJE2BR3TvoLbpczuAcJUKHDkqd3yqh5W+BkrOmhthI3o1M/trR1v2lrGFC1+ACC
9kg/lqwF5fgXN9EXPtqbHGAEDHUqZBMy2YtKCuOGTir4tvZ4A0+FI9f6bEEc0+j2b821MF8SawVC
XPI/jqM6CDnTX8IEOyQZr5CQM/WRQqdsL/63yXao4S/5rDzQkaMhA4kJzlNaKzz+c3ZfQFsjPg2w
baES26s0PlLj+kB6E7eCc+QC6oLVVpqSc1u3ej/PviSt/PtLVjyYgXrp2EZzgyC3AlYwYQozB/AL
Eii5iCadvDXV5Wxo1RbBEcMiDmd8my6w9gFZk0hkG5rZiDNwUxjmD7BY06/axmH1nC32pXCEWFAF
DAP8R0GefL/AcTHvg2J2uJHhh2YYZ5EeJwt7KfjdqdfIRc5DLpMMU0Z7ITc3p+GYJPisD3WfijdJ
pkCwfNtOxSnfaKPlttaXpd6g4FtMU2dV1X1qinQOYN1u6dPcf5nE2ff06BQj54LS6eVZIOLVmf10
DjDTdBHS4bkY370qOHozn8qtMG4+hhNGiih+5Q8ZVdrVGlVDedgCNJuw2LxIrRgsUID/qyxDVik3
lb+N+2+JmiFOx8rnBCCxumoonHsFQKfn/QpUuX5gHbxzS6bmyxv+V9BH+qSSzsme0EMbok/aZ6ka
Fi4Dd7axDX8GgBFfivIYTesPaHQ3rLlGkTCLXX6bbJWjAT7Ld1sW4Db7BcxaUWuY4Nbf7HXxFu0q
2ofdsYB0rO7hwOqFHM8IGQbGi2KB/Hq+Xq+8X0px/lrM983UWzWarmr79dB36MeBpNWopqGNZ0zc
jzqwng3Lll+yBM01kX6zYXv1K9gq8xt7E9TDj4VcWSUOMEet1Bv5OqSngSt8ESMbeXyl+Q/Z5/aM
wk5ARH05706UO8UbSBOj0VPuNIq+eX+mXUN7ddAvbJ0G5NdK5A1WOD2bBsy6F1D7x+Guwj4DnZI9
VHSnUtsDR+pFug9zGCPfXsM+sB4f+FKjopbk17OZoAsJp+XiPuwP19HgOGJFDMnMHHbT0jEruWtN
s/nJmYJ6kAVrPCb2qXS+1N4CO8mbDhhXhc9Z8hqf6LAntXcsR5TCqHJedXntLEMi0Qgt1tkYXkwN
yNdLQUmHgosScRa8nscy2pLG5ObRC8BdbccJejyuEjqDYjve/nCTRS+LIT84gFz6Kky4p/DF+qmI
d4u6iv0qzzPIRHGYWpSUNQ/lFbMTAxQcCgpB6NCo4VAA0jKrDta2TSnXO7+MPOwW/HYEaGQ+dqH3
k9ufw7TUzhEyE3HF+IAzEgqJb8JLTjRSbUV4ia64hHKy/18b2/cWCdfZKOw0koUqt6dJRoGaGA2L
rAwnsjd7Am4P7oaH1mE/FmZY91V4nLXbHQcfz7rlvZm9/CLCSPHiLjkhjuKbR/rz3+Z7l7M8P+Na
dHHxg4lAbLXbBwxUOzdR7172AVIvSdKmWhjHswdvX7/davPjwQmD/Dnoh2U1ihz17iHmx0rnhqBS
viUpfjqpRW8BjaGOw2932pYSlCHTJy+WoUlSGoC783v5IuCfapHg39X/5arU2pEGIBL5cYZUkqN6
PtCBdbiZbSU1EXgoo04sTOK8x9Hh3A7GApx5VB9yFvsonGlviKFfucJh8WFULK+M7wOtCDhrqiJ4
Lf+MeOdLe2inVsPRQjU8qJLxVzMbuQKwFAfK/3Tw9+1AFhY+sjADMX/yDPHMnKH1WFmpkL0Gm7TP
OPbacbG9m817aynlOmtpdestbTGi1FngDlDkuACpI/MnIyX3jB5xup/hsUqk/00UAidUYOtjfp4S
9Ajr6hCi9k82N8Yj3pZeimepMBOrI7KfEvfzjHu8qqBRGI0EMuk4ncW9XJUAFsOvpow51zmnN9ad
cLX63D7xVCX7qGHDwcefXeesfrYshOW+4Ex9Bcmiv098MPDKgOXJEQycDYY4aIp+D6CIi9kf/vy2
DeE8A09jv6Sb2IKxBWYh8XheDPCiGZAphyPilJ8HuVPk+ZLOEMSQOyFHAfk/FekctsW8MSPhyhYJ
nq+T+BPfaiKkgIIxU9+VYOK4niSqiFkKN2WUl8vrXeyZkbQQ85++DglHaqPQNj+51lLkoZBo6O16
zqp5UBFfhdkrvDHt82D5Wum/oFyzZUoNwJeP81VILG058xVNz7VRNKaqUFeBmIt9xyxXlLGSdho0
F8XGPgN91oU3oQXNKKg/x1EAX6jGblXvrTAW7y0kOLdIdMKHgckBdO1imcFjZwhsM+A1sckwlzAG
acy9OSOmSnO3PelXpv+3jrW0J6ZlYl2jhcxGahaxhVSfYXIYxLCvaPc0mw0kKtaWPxCJorZajRJa
U3PZ1+aVG6ALHIUaT7WsxuLzJ/E0BZL3pboKMwWSLZaP/U/faFEMJaO441Bf/0i7J4kGl1U3Uu6Y
8GnHSGszYD9KMnZAuAwCDQrI6GS0wsF2wjf9OZwmE5uYL21Me9KuMJrU8vZZKI4TFCjsawPkyrDk
6W3axgcUttCYO2GJkkuZTiXa9IGxT0c/a9kib/5RwDBY2seWlpZbeLbC6t+OvW5BBBILL2yM76Yd
/8zARFgZP2q5RBZoa1bGdFDq1ORdqVfwXCI1bc9rXq50rF9JOg+Wyy4aj7sdwTXvXQNiy4lMru8O
1pmubW0le9Z3CX7ITthlB/kIVxlx6xnGZDvzPoI7uZP/KBbpdBTRIMR9Sniys0bHk1Y9KWUYITwR
aWTs/EXsBlhJg3JwIWFBjBtoPDw+iwLRyawsg0juxpLrxYoga6HYNIGF0pfkZIKXqzQ7CEAZFp80
v6oZGxHF3HdUhlxFTtcOk9GQg1E9+t8Z7J8nxPVc1/jupGfAr+0hB9yaIvZkHWV2S2Fvg6oPOTgz
/E4Il34N+bk/Cqa8SOAzLL0CUAxVBJR+MNEj6Htjyspj06tcg6zKqdmfWQFs3qWU2pg0W4RKiW4v
y5o4rx8iQ+ByOocMHCyqYfKYeQ/EQBprDJyyZWxdOJOLufwJprqTigj72x54vB1/g5B+NJnXcMia
Uz+xk503UhWZ/uZKUXBWtzkTcpsUD6PPTTWN+qNQjhiUQcyFhrEx6fbSYJRzxmDg5xQoixIEnhKa
dj/fUm6fRBYjSkEyfm/k0wv3EKc6itAJuu3yRibB1/jgwadq7OUQRIdqS8hSWJ7xfjoVc423Dy2m
LT26qftnivpa/c+CYqGKdjM5JY72KiR5EByHqdvQDI4tOuBr8fz60xxTPanxpIvQTIlBOqaD5Qe6
TU4W3S4S22wQQOwK13KgQvKocKnPNwOXX5i6looZ7dV8mULiUuIhrmrmCEZDWF2GFLVLj+K6R3nU
Z2pGrfhPCS5drsq59AuVjuDcMJejO9t9q11dLQ2bh3egLu7/1X4N+jjx9DZQjK0r2nOqGJcBjBzz
CvNu/h6YtOXhnSsrfUo1yCf84GK32SrUTRWg3112kPT+4maereRpEojMMP0RtM7Of4nKtwtD+IoZ
fBWHaD62/AKrVTXOfkwiO1hNNemOzjvKcrpBJc0tfW9UwusIYwrhXjFm7NU/a/IbxVSnnTNfo2/+
uT8E5TU2mN0yo7hRT59976azMjrCOsHgMo+UQRklm+wUbkNCifCuq5kVlZaHmiu+9sg70U82zjjP
zAL2OLu85MN32o2jHVUBtxBdzEehPBUoG7Fpcm1hl/NvK9kTSjxvgLX6L7kQ/U/v3m4kD+PH+PlU
YvvnRXWFP0mCp/h+TyS8/hC/Ky42la09xieZbKgcBDl+UkePiLx9LlLzuqlDbVduBNALH5spWwJg
6MkSz/OM71KNSzrurirHhM2LVh2jRcy4/BFualjGL3XhNGTyJomeh1U5SU3t5T7WxXViWdAr8mMB
WrciAgi/xPCA3kUMMU3MqM3hq6uq9URzPQEY59Lr3ZzKErYry6v8NIpap+AVCLZ0/zQiw4i6kle8
sM4B2hl2Hf/LH1yKOmgIifCoT4cBt6RufG1yVCxw+rYZcWM1BVQ+mIGeyBQ6NKexmV0PoNcrUBgX
22RKzNLmhfvejOQn3ydUw5EIU5LU2/7GVKpKHkQbAJ5O+6miFtSp2q98uGJR4ojihtuvjfgVHD4n
b+2r/XZzYywH9DnMb01BWLzZ4TWTIn28me2ApNB9/oC+H4lRCkjruVc2zU2MPD8ffny0knoK4uGj
DyInZdwjh+voVkMN46ON7gfs0CCu/0E4s8q4LYXVt8LJ1tup2xy1Z1Y11N+BNIKR9OQflEXmkoAU
BLzseYAb+kAONvPIheIjGHaGNlbsXYgmbLv2NPOi/1sQvZ3Gti6jizDqEq1lPJw3DmaqYeIhAQEa
3yYGTl9qVqL3EgnBWenurT77mPdcOmNw8lxLBhAWZ2Xj2s8hLlqzYuRhO/V9NTZTj/kYCcmJI0zh
sUbfzcBSd8A4o6sjzX+KJQhT7u5i9zk7JCMtmY6/jLj+f5MaqljEStecfulsiOQbB+AnAJvTjwgw
O2O7Cck27q89sBIxlNNpCAr6r9Pe2HWGSXFfoKJv7aTDAgAGqowuMovmGDb5Rtr4Tam1xE7c0eSV
ig7voKp7t7xc6QxjebvHPCYkpdJne8ttCYir4ABphyJFHjX0WlRepmtYM7GnHmmdhSN16X++Uhb5
nusPLfqgckHY+F6veGZP1TK72bN+ejnlnG80wRvp+Qam4W9wgWZp6t55w7rhnHKB1tfknZPE62MZ
k4g6xQchgoU0pnZ5eK4/E0TZuGl6jTqWV4xHN++cGVMMqmlpFXKL93bvoTrpWMk3FFvy3I+97z7Q
3m+bBrZXUYhwRcQhqDGYgiGxmRJMzldICZDFPfXrOqMsFUHI+U0rCRFlSELRPTVz0UggtRDAzi42
pDjZOg1WCIEbYI3N0wM7xBxcsF1PCzy8TSJLXc+kqaQEusLyXdbNrWOq8fIWuehl7pdchkxtCXTd
I0uioPpo2VebJ0FjdpvLG7AQ5cIOpuArKYjknDQGk59jPkx1KssjPkMM911icaFNIPajCiR3PC8L
ezdRbRKjJHzLHS65VJLGkYMTmjx/fuHwCUWwe82onz1ML3wjtO9o1N/HWURWCnIoyOoy2899ESB+
7VVC7ZPXAdGHQcexyVZgYbyi6NX3EH1V79QKheKYfx88fuU3wRUrWkpT3PtKlkAVN5yBeSfYVrbb
BsGtGaMaW5lOlaUtQBW48jUqT9jMzMzPXcswwfoOogX9mbO0mOxbDupx9ea9kYdGFB24ESE4GObW
dKJEuemx4avbgU7yR4OcKXX4H6/5Vv1Z1BZ8n/T8wZ9jTKYlWei/bhsh2bq4jfCV4mZLXwRkXrsD
NHaN6Fc4HWLK7hNTsksKZ2a4hignxjKRnUjErR4T8S9lrSTCD+8EsGyXvWO4EJBWDpzzwdgR+n2/
wya7txWEdcKyvhQ+3E2VzglIuV+R6XyKaxjCcBZNWNvrkbi32COd0EGZZsd7cQuNuMfVMUpa+47o
4AIcuTvhLV0zxw56CW2Z0tK161aiQ0srRyJD86y6az7UrSpYpZLXeX3Wpvjks7es5RjJhqcFeVI1
zMlSoER9Gxz68aLhl3VGVEuWMLgTcLISImyWfxyrFJbtgaAZtR0kWDUw4SjRKUEu3E8xTJ1e4tSq
y3+diwjzUyGWTbFT/UujLCoOyNtJe/DfbnTi8fUiUeOd5l8Ew71auhdOmvMS7wCSZMKEZG9A1zzm
KdK36RbaHC8GVOWKYtnYyJLPAS+no8FDKqRTowvI3yC2X9UibuK/RsuF0J6efjC7iYEMrdSWP9rl
ufy2EfcJQf/btBO2XNkZUobUcOTcf9T4qw1uA2Totdj7ALv5aVLZdh1gS5i5xrB/sVYWr6vnUCOK
f8rEsB+3tM0BcbGMOT/H86suOg6B7Sfrr38wnWDZF3WDzTD2qNkRtaX+rqzPyx6Dy2HxBCPxpSMl
KHJtjip0nQg3y0zjme9hNhVQW41dLRcwAFIy3YUn0+VendNboL8hgUXydSxbjoEB5ENcivrdauEv
r162iPK374gihbPSXCWpPQpAim1zMmuvwTyxJe1ZnSytzJKyj9y0tdULPf8nMTZJasFFIJr36ZTK
pmaqbRZ1KOUlkiysckFSwVTW0TOawy8kj3JfqUT3YKd2smPcmt2wrwsklJ2rXbfXADDybEEsgy9H
FojNsYeSbIFIFFyh+Lo73c3kV9NG1ZagImZMxYn7+qxP7MGNFs/a7KJt+ar3Li5ds3bUltpw2QRh
dqPGqyb8NeoRns1vqNjmu+8eYikLTyR5kOydQuFNDoIy5n0zvclxZYN/fgKJZt4gSnCZfiZo9wjM
+MaKpTdKqUVr3pRVW8Ws+sVJ97Ok5TU0NYrtjf8cgpR5tVid+w6/UZmekc9avVWazqH1OC4lNMSD
qhnJMkEy2wac7KOk6+XWbiP0uNYNqu+wr+T0XRLJiOals/kp6QxuQ6/Zg0E995HqpLh4zqzbexYr
pKXEj+QZbwSb1hl66hmjkV79RUFFrNbsCh71mcGEDW8mSC976pBE+KiHmVzWpGiX851N7i6giAfd
14oB0RnyuCHzqlF9PMdszm1B/qar0r5Mm7ftpvcGu/LFr7qjWmfSTCyg0Sdx3QdMU4QHARChywTW
dLk6iLbMFdUqkL2kzhLHnCCFlJTJsvOres91UcHAPfiOigmDioD4gpTdxJRO1yl+kPk/6Pae3Xb0
BdrRPeDh5ka+h/p2F6TG2/PC9k73qLzUq03ydHeJaimOyzr2rj0ht1HaqiaxjhTljIi/RfrpCFrx
98opvj+4ZSW3lwfTQFrZiPVw7Q/L7dKMzRZyDF11Hk8jmcxSD+MLtUarc1T+mZrU8RiOY0fIgTu1
4r58HEXQbBhguWG3WGmRLNchPg0WCTrL7oHgUcnOOb10bDFbV3yjIF+f9hMpwmSD4rQ5QAE2xpuE
vom+s7QdIFri13Cc8lR8uixxdKuP3ikmsGrjpo3g+6+GNdQiorcQDCO7xPWHpwwY7H5FVsZN+ecK
Sx2npA69JDY8dXxu3JnWq8gSCS7UZrJwuJEF4vEOjzluQcqv0kO560YWl2TbL7JRivhijGIba1tK
A/lfkRCKSfHXeiacog2w1M72xnp7VrdMFVs3hg4B+XhFOYd19L5zay+XFxdrvU5EgA0nW4bOlLlR
Qleusam+o94xTACWyNimBW5B+jNC6rmPO+QX0byLhNJG7D/CZQKowXKfBemeM3KgBs6FegJr+672
iBSaMMcZtrPz1MsdR/7x9goLaC/HXskPgkgpCs3YzeNF1X8qkOjw/64LSwfoDzCz5PBzqE59Fmmk
lTkFL5jtW0h0gjACO0oV85PGHd7TQKwKM0MCYeH03n7FTi5LzTAqGFdiUcz2I+Vc7L5LeSAeis/6
4OFnbt3d7ep55CPZmhmDoVckGwmGI7bOLkYD0VukyI5oxdpE8jAKbgsTVYaoHIqHKatTt7Z09FG7
VigzVg4QoDsIMO3W5jCfOA9JH0XzDTNmP7xl4R21QqJMQ8Y9f3cDiJx1zQ9OeppBGIJ8z4Jmkouq
GIqS/eFJvbYpnxKrka/bKdOrNQ7ZQZHKrcxXsXUEwdGtSSNviaaPp2WUOpXFme+j15Fg60jIH20Y
P0gt0U38BztpmQejhvRN7a7oyAKur6EdvUbII6e7iZY3NeCX6FkswIO1ihvNaIkICZa7yCpZCUFu
MjNr8r6k+udYKkCbGsDIGpaxkPy0IX9om1+Y/Q1HJfoDKBOIbL2Nm6lXbeBdYVJWLHv6PLS4QERY
32Ph4p8X1GJxlcqbjzKOKHp5AezX+zJZebyJIdRX3YOasHvPmVWRqdpxQHg+zm2NHLUNBUb4ojLD
e9EUVTn1uu7uhQ5BEMIJafubrPqDRbF6H+WI7A/jG7Euqfu+DFVgijHBk73RmYXIMkmXJI68bAUN
WLspwnSloiPRFwlm74KUluCVQEzOPeCnjfu/jszMNxfIRzlossf8OnD+CfGWgM5IOYkMjKAuWRmv
NCeOcQjZoQjzCe6Rp2cAzxsUlcJtRFWhj+fWRLrel5zaFduxEebWqS01w71FXOZ9lzfO5yh/fxLs
ZejCkillKKYxB+tKEAV6/vep1DzSS5+NXno+IERle5C+35S9C/kAenKAgK+019niYu1TLfeigKY3
SKsc38BrzO4OyW8Jubh0+hd6AaYZ/u62ltXtAuPICUbvny57x0h2f3U0vJFPWUl3T6k8clF7yMTl
1mvkkPiOc04+q6fgOwraomqUeQHHdxQ8wx4ajk4XwiyM+RHrQ/f7xZ4+R0OW3L/l1iVKkL6A6HnV
Xlk65BaQCnH7gp0Ry+JEX4kOpemOQVIZiALIoq70ogQAM/J0oNb99KUA4Ov0dWU0sggXWalGk1tF
CR8Dy/MIanw7xEAZDf538GJ+dElRGbE+15eltdObaOI4zNV9TYknOHxZLa4QliKHJLtdTaasmvrQ
CRb9jNpGbIDPDo63LLsYSo4QgCm2lINZA2Z8WN4eUJed/LkDzWbRvW1GCMwtusKL45LJ3y3wr3MN
wqXlHF+Ru5ngVSgD92nIcgoLUUI+MF0b7D063Lh2JAr2x4x67WeQTOPWg+XXANBJqaxxCmLALDAO
vEn2SmllbC1H3Rbn69pQxjcgacC3nHOyR2Z7SpM3JhxlcXSiCDd9anM3BNpVCknCNjHgoJBr0FgS
ceN9CZsKTi05QT7QMgTl3aHf9H2YDYnKJLDE6NLLCNbIAfz5JKqzlJMSFaZ75n17f6IC/12ovdVW
AXqo7AmTy+hfvVtBljn4OmUxRZzwNtximC1zkFYae7LaJOv/at85WmgFZ8Asp8K4qTY303xiSYP7
MNfZRf75twiqgGld2OX/vnIuk94v9xva9LNPAjzHmQOfznBJboX80F57GGF1I3vRW2u5Pi7wESod
Z9LC+pNfItZXAvJQNIHUAr9I6HnFnNJY8z4byZpaPRsum0GzZqQI6Cc6RMi+sXT1yVeSoAcwl4nw
4c5Wu49dtGsVVqKWFT/bBVc+1PiOlGuBHU1nn54v3MSaI3kjpR0RUBq9x3Ao1nA/4X/2JtrrhkCQ
kfy3OfMZUAyXAkyvFWWx1hBkugtK8amF3+807lP6g3LOeNnZj5EyRmOX2bYKeLfkgUiW5m5mpnnq
gkN3LbDV2Qp/wpSH/msEy7vB1UbnX7pP5/mpKsKJyl7U31SHbTjFB4HB727/dmkkoTV+dyfFoOBr
a7KdSJbkXZjCOIkMLWQGayB+5KAshgwjhO758xABgr87PZKrmuaIW7OK42DUhbGL9RO8FWTgaFUZ
SRkVumUPou3GlP6/lREJbL1zC2V89b6DOYPCW14B6AeLSU7KVNQWXTI3CULyRyQ0VLjXlMecyv2d
yRo9JYI1GvMKtewF7x61k+scMvb/cuHZwVdJrJPWcBJHWo2jQjAtHrCifEEorb8/hhF4SHoa3Swj
OF33Svvjgy+WTD3XpPZ7Mv/gdWeNyyxZJAGDBIx7B/dvajxF1DkX5cpRCKl9IGF6smGx+sVtBp/V
5BNJ7od/RqiuVPy2lhsNzYgs58erV0OjsU1Ik3mmXIXyUvSMX7lWPlquX4SF6pyvwYljPeLhqxnq
M5e803WXvxyJvIKphT7BZoM89ByYPQBDmnhPush1CssCnm72edyELZEDa61b8TmNogNvH9pvYn4v
hOWhtsfWWcYgle6e6ajJ4rGkTiB9ZEF7d4PYP1JCxtIxPhh6UC8dmKIUt9eLhsmR6SazdOjIGokn
4QMTRnTQ5YyuNGVYF8JXh7quBm3LOL36toXPS2J5JvSnEqXCVjB5F9tlByx4gI9fovtMN2yCDje7
L5pDfpwBjYAAVJROLulnUiaTjG1bNPe/crD3IiHAxzwPURnItQYrGj91NZyzkMylJYT/FOC57sC7
N7Xd5Mji/7GjPhsvLqd0/fVKfl64+PotUivhhMgjjTBT83ET+dHPLWvkucWePaor/7456zQ3h5/1
oj4a0Fz2bCmmAYytPpaD/tBd4rFd2G3GDA9pLUvJBTlMGXb8+o9Y5DVBfljAuSwi9o0uQ+Hy0KsD
S7DdFKkq/pybVO7PJRkpQ7WDA0KQCYDpK5L9/SzOYYNBvZf+/KtgKU2WWnFJawLcB0ElQm5uP9OH
5jj1Is22alCFAE/3EXaaiH0mR4XEeJ2Gkf6QZqy8/tocCaJXarfbD66YyazXYDz/ak82xu0ITqwf
9lQVYOMJQ+Z273I1VB60usI1lSXSh7TAvEmzvMf+8EjORybbTEIgMpX0sNVuxcg9z1n8kFjksIMc
bC1j3VxRTYXEfU8rBF+W5f7sItf9TxgqQ2Z3nPAsBVBzzKAsZcnixIBaa1k1tmEigPpg82jCvwUx
nwZkftfyK+82M1KAxBWu+OVkGQLTFgAjiyAMTKLJxBj45SDuD1mz3VE0PZlGD+IZeVFwIDqYBHt2
VFXE54TPEX/kmcqzOZJj8PJ6HwFLgzgrz2aYmjoslvI9WieGqsBOUf4wqTqOF1n0IM50y2q/E1Ln
q0zenU7aQ33QOiT8H15TzHfoqVky7YeHKz6kwXJHtMjhl6bc5hVPmMpkWKhgW5mi5OkYeL8bx7iD
cYFTSCedmsg/7LKSvHQWYHXPW8/WYNqack2nEF4cKYAnOLVXMCadAiBe/iPvOCikpKc072OAgkpc
Abd1v7F/N5z8epzGU/CuMpioEwl5ATQl23gQWfT9KmtH0u4ZIVjtgvyQLj/sRFkE3XdJQxBH5BnC
vxqMWt7Ie+VhV4bsTTQxsqDR0v5IJX3i5z3lzfUyyVhi+I8ZAGUdtaqNclxjxfuGXWGIr4DRQ8Tg
IoaBsQ8gbpkQ5zAYD6BQvHDQMX2G2qzH5rKr4ulNGwBZSnxt0Cwdy3qe+M3R/uZsc3TeDm6ujHv7
yPcLcorRz9txzhvHQwk4LaphmjqWjaOZDTmxofWltMtWzKXKz46mFyIP2mCvF1qZS7VaP3mDUEyI
wFtKkJ4sBWwU+2ojDgsGspvnwMcS5p8MAAq0+HCSxyzmvrF1FNAXo7gbP2NCp69Mb1IvBUAll11u
AVIVSBXWN8NRPkCIb2PESXqjhCrsKki9Soc5/5k7jC9DVaRXq/3px9JkL8YrnySh74DxEaF4JK5z
fw0PaP9RQ8GBAaSp/Lpe3WfIk9XV1J/yDBthw94cDueFSrwp+RuSAsfJFB4Wqju4mPLtJWWWItsr
wQnZrP+UXaL27t6klEkHz5oYgFPc+HLjjgxZ6hOaxvORPZyO5oNHfbYefXfxmeimswryz3Vjhtp3
qQLH3/0vry6EO2FeAfnLlfSxaaG6VEK/Ob9xCkYjJZSFBeob4u0ati4PGMrhLQuSk88IOFooSDZV
oE5u6oCv++5FQpMcG+1hUE6Pqd0l0rQP9FShoE96jyUusR+MmvYeLbBgddfH7UKsui2hah67QPAX
rMgvxKb8I7Z+0J87ZJh1IaAlrZRlEXKj2eZ6iblM3KFi9ol5DHkqb7pZp2HXD+wzqddEdV06XpJf
cmJu2xYda3e/IT7EDVpSwKjPHfUql1puvaKRNnbPi7vlYtsrqScBcNIJKatxxRKXEUdrZ8KgllU6
xgkmNa4gEez6CWAxtnzqgLfakajKUoNsvSq0zJMaOR5xY8AIK9+f7UCmT4JOo8pkbnswYoaI1v/n
21dXXU74N4KXtOgZ6Nl5miOduHxP+NRHXljRpKQWRiGr3Q3rIoND90nDmPKwlLy1DJwQHRRgZt8O
ZisHEOeZsEVNbpEIODIcMoKSlxZJ2mGKfk7GU9PTxVbkJX747rqqnay4bdRBEa6t6ENEFciQy3G2
7DWSmP6+/sbO0wRBi0suSb3E/lAUhLEdpzldBa9EIEtqc7ncJW+Q+NJeNHSVmJjfYR9IHyC43eBZ
sGlDTRDk5l5KvUvDSGbHnzfzRXNmszCTRcqUwWiryc/l5uBbSEkmNV8trLLJa5uYPmu4quFvD17F
M97kIXNOMwkbdW04IS+af65+WrGwZ4mShFVRTgmvN6kYo2SBaYdsKRQulZvzGXkttxU/iBJqOwtW
pZu9Dy4BzO611rfT8Moe9Ph5S6LpY832HswerJMy+T+fxDD3Ec5pC/zs2+Yh2aHgCLfrJ2trxIua
FjE0aqw8w3N0JDfXyPug44bJJe4yCgDw0ZyG6nweLnaD1KtSdeBlm+Y9RJ/3ELb1hSFsyEgpvapi
ePvrEKciwO4Eu0xOFk6+gvuVTZ+MvlAzP6gdlPRIsbZQ8d6Y5wIg+fUHD+l3+sQx1zh3wXi1ewMd
B3KoWaDwlsVoSvh78VWScgdlHqXBHqYLfTRS3pXXHarehT07alywehOHGqyh9OlgJfdgj2R1IhFe
7uTcOej5nefEruuIhm2ZXNouunfEId14AD/AmAH+X0vmAJOMH5D8cgj6CUlLOgX6cg9Kr4dAZp+T
kAPaXlIAuzfk5Yrf40+38C5nMPWMObumEPzHm0mkaiXGVtPK+ttlV3pOwqnbfn7kzljxHs92wHNh
GY+TeBnxzZSpfic4CK6bTvV2E0cStXvD/aiLvddYt2Z9iDx0AzFvfJaGuC1ZBUCpAMWs9JCLsI1D
f8cFobwBdvw0VQlXZ0tmqAOVxzp0Gq+7yhx1ycyLv3XatULiQW6vmaE5rjKiIVA0HxLMbWZYdb64
/kWHQgK24YfwrnQrsZVsf2fOXZwTDHQw9UG1pBLVa9vfLrWsfBOFuj47hg7+tgWClM99/lzfHYNQ
oHrTUKSr5VGbeaP4Wo42xt87dOB5cuVe6Uh3ybQ8RSVzwWnf0X5+nr6UW0Bzmay7b8/CxYksYgwu
rDlETJbH+m9di52H95tLFlENUDFQyX+Mea5MRfcePcjPhPnahiq5bnSjW5v+YlHoARPbZGS/OOh6
3RfR6QuJZfNgfjQ9R4FHJW0xBZbwqP9Tr8U0zQ9ZOxsSt5iMVqRh/kVvkyua4v2/c7Ps90Dj6Ssr
tUjtT0s9Jaby3RVwsmlAYbdhtrPdQ5YkeauBlSsZNJHp5b3LHlN3p8qSQ4GTBKEnmphdVyEcr563
6BDbX4yIweeBwjSWOlv49Bw6gUbmRzbXEMyTtnZBGDCBJutqoj38g5vAGZ3SM76cZF+c4KK+ZCC8
I8IX13IyGCy7oEweijZoSNq8WH3+R/4LTBwpPQ4g9Im01HAp1XGLNR4GCmkQHKq3rm94V/reNKml
6EhbltdzfP/ffQbWCQlaHGfZpC3vgy0dTHUknwK7miqSC3X4yDVflw0OcxvXWnqBVRKkT7cJtk+w
uMgiTsruRaJJdkdzfKFVoihccs7tYHPtJCzmVutflqSZLZbA/b+18ALM722Fr96j/HnQJCew+hD3
R/F9gP9KU4J9mBsJWgCc2PdXXCvKz13UAWOjwyDiMU4DOzS65QwaH0onk/hH5zy3KRCsJyIzrHJ3
PM4VfWmFt2EnFbBcc1+zjGty1BtbTDr5oxgHmX/AguPmIPCBLaxQ8KbesSOscpaUX0uqV+mmama/
DkPTkgE1YgGNY/ivKH4++BgTFjekznai2ewyKoKbuoItd5elg2jvjdmVMrYzeGokFL5sTTeiy7nr
JivILQDibZzUNMzefyoNQVilQ/t0uFNa2Ceuy2xIBpsZwfvlU1+w3h/eJYbO9yErlQvhDlcQrR9u
TJR4juyQ1ime1mc3+QGtWRBf9Mvu7/eZM70fPUjffOnmrkqjvUImZF49KnE96r/8/L9ibs8ModLs
sHSeR9LohInS3VJ025K/fWmbh/3rhHOj2/TceC1UbAuRfK3Xedm9vdDgd24+6BMaruzT1HU7DQix
lhMt+4a6Ocu5CbtUIHuUuGw2toztn6lS8t1iIJ5OrmHY/Bk1TKd98J7OjLxDRu/ehMKK/HhfZRxH
OH1udfTYexjbJ6IxvhANgIbXXrf3hmLpUvTA123p/QrHgmF71kkGtE0fY72sMcreypu7d9cmsgG/
RnVwdfL5aGK8VHUma3Eg5MOse02EDg00A7cVB6eHVd5y98APZSlAYe9xmVAHXnrk9G03rwQufRh3
KHM66LlkcNveouqtpWzTvcBKtsXwsyt8ifOTzJp2h79vWv4T83/9xHvoo/8L8LZSP8ACDD5WwcYA
pWlTxt6xzr7KA01dSZs3cypwkwmc2m7IK7CpBGhEhigKGr4yutdFQUuJv1SnAUr1EmXWszyYp71k
WFusMrwPIW5J5aaTdTwbLE5yJcNhLJN8gZsA0QQQvTW+Uvza0ewEy/CeVucPXNgyG2VrRMNeKmOT
5BdAbYtROEopwLoD1MSGlifwImm40IGhdWz8L2waFnUOPwDCM/N1UQWjv+B7l+sEJdChR2/rCIJl
DHCeIAsEXkOB1EF7y0wOlxZ4Zu0VjaaISAj4WEXCBGfMDHcEbPWZjsUj+uWhD6ajCymsbV3+fej1
e+REi7p5lDNfmIOBuZ8f6Pgj1pkEsMLL26WnhIT7AoqN62FiRk2TkLpfBnx4XO+zObyPeu/ePCgT
jhYarfEPOfKUxs9S8ubSGHIdKBWxqGJ4/j9w+st6DS+AGTI9zaAiXCcbKCw1NVcalTVAjTtLeAHt
wNQz6uDtGuDDTuMSf7UOD7eJUC8xN2NuE3TFy6wVfdoWInwi5pO1d0Av51LojubffSz0vHelhixJ
fFkYBas1mkkDo0Pzjp6s1p7UU86XpKeOnTvYD4eYlMo0MEqruazXhPsgvsQ5ODh6KOBKYJ5mGRf5
AJ0QYnOZdhtepxUcHSSKx7jmkfUQN8mwKJi+4f5KnNdOsVb1ZDVxvJwYjaxBAA0Qn7Q2M2pfHJBu
33uoIjEJKAXLMScGncwB9T2eXnLTrPlXN3QrXWX+/lGZd1+OxZzVeh8NbtQU8PGTe98NM/MXdglK
zGmlFpuaoNGdOSpkve5Yvq0nBrvs90+UFjL1tkVwdtWwsAwzPgzjQwnzoXfDO0tFXV1Li/yS+dHi
V2iBl8Suh51bsXIt7vWImkhRdJR69sOrPt40lh9iynhwQ7CK4cYziPhw1S6cN5rxECAEduPMfJ1m
DhfLWSkv7B6a5xz00S1rW5aND4dk1RB9EGn0/VNzjt0Fkf0I26oF7s0FQZ3zWeVXdkw/kLYsfOfy
rlqyWnJP6pGOHmdP8jFaiiVToaR6Cy0+tDMtoQxaZfMx+29COBhwQZ/tQ/CI8dV8bRyk39KUh4vl
yfE3uwxXOPfW8QlDZ1Q/Aa8bt7QvHDAf/MQRaU+1t7lTZkwuVnC6L03ief8fO1y/Xuv5OB4K5Z+E
IzR0/ZK7oB2wofxScAnuyj6Fn2TbBUTMqePbBr5h7oC4hTK71XwJPrjA80FIkAw+iYZtlt6GkgQz
ZQ55HJ2nWZUU+a0KQpYpFQbdJs6hX07lAgE35zvHsN+oRc0dA1zRjxPOxQG/kUt1++oo51EQADzX
J4xqev63kDCOXG5CFMG3Orq9gZkZsVF1l0yM9PWj3zy/Lg229hyh8KTivgGROqjMUmRuop/xLz6y
NYjytWQL267m7DHQw/NXFT6bGfVBY7GbCkH4AunH8ATUUslm0/mMLGcJcPa2r2wMmqRyo1nGZ9/z
fIL53EpM0cprGr6obgdahriistR/Z354o25O91cOSEEffw+uitC8RqH5UAziHDkfedmN9COuKmE/
zEqH/7Y/Pc5fC0p8smaaMciOzEgLas+CDKyl57fuIE9J2jlu5vABEJfJBY9/+1tyRYpIdJ6AtTEQ
6Bja/Qewww622f5rpaiZ1E3DEmfw/+ltgV/uEjPAw3DCCUs4fCJIUbRqWIsiJQj+uN+kK9yR1V4l
SixnSsXKgVfF4mzyTARaKvrvgYbrqneS8yZasyjdcLlo2v9bb8kOEVHE7dMJEkeLTd2nw4oA2RSk
FioQlFQFIMrW+5q9Gd0mxrwlWkrCNtDHa+qg4qlBUaB12b4oEqeraAKaZQbgy4NXXlaA9kfVHkJ4
JFsGX6xUtzsaB8sx0rn8JfIu0I2sxVZG+LQcMUWpgsH1ah7PU09hO+hy9rIrdtQZXvl1DKrAjE5q
0DVF9YpkI6B5DTCPXqluNn371KQXQLZ5kT428poPj7FuW4k9e2UThn3M0L78ioOiznd8BhZ6oKY9
+zmdL5eDL2KZTXtEyKF7AkqklkWkfTphywkF/0cURB9kyKe2lKS2WnrL8JU5yDk0qyqDDAvfdk51
yCOhSY5+oZ8gUS9wMWJISiEL85DHWNpqV7UCfO8UVHWew9RXblFBspu/OW3vLC5jvfp30ituFW6L
Ikt1d3L6/3aZkXjTCf2s8QNlchSsIMUhf+TYZyU11Kfq95M3VXzLc/HemFLBhfwMzpMHOE5Kufwg
4ouRPALMCny/s5BBY0g6+XzrjqRZ6nCF8KwPs00lI4q7WRWM///PyPkXILhcyyU1NZbvrdk2l5R0
IfLTuNY0F9ZaHAuWeXU023FCIsKP0uAPGVL8BlNY4inIz9lu4KLDOJTXUoiz36cHveJzmv5pirG+
64SnRTbnTEeAJqyrHCWwad8g1SF18qdjgyGsKQQHQLTP1d3aPEzbKdZmpGEnBNto3/QzPITR6kLr
767Uss4ef91iZCfsO9PrlqPKAv7mMCfLv/cpI1P4YmZpIFuzbsc3KHiAU3ggUtPBIUvM0AJDzVYT
xkC8McYpc0JSp8hsHfIbbb8Ua/bMD/sLSjSXLlTKh7KuGjZOdunKkwVZ6hxebVIIva5Q+MwYK/qZ
jK2MgtOwVSZX7uwwgwwOZ5X2gLHF3uwy1TdZwwIFw0iUqZiY9pvEGiOUBu6NTdyiCs7DUflvRkFH
eoGoR+zPbnTPu31Oso0m6brvg1gBDt6A8dXiZg38iEEo8NrgKL1sVFGwyLhTBq2vR2v+tkh0ooAC
5UBRVNpKwHmEcnoWSZ7oy8dMGkg/AQ9RN7oexCZnC8BiQPhXaIdnWo8PCGmLvy/0B02CsfQplIgL
2r6gQsk1/8csJdBDOsxXJyicei3P47Yp2+G+zbQKBwJ3xVI6yT0KTAPHXyo1n0/6nF9C4PhRLOjA
j26VJKLLltLUaE/jIOIrPqskpZzP0BQb2cdFOhRfep0pS75LFD23CDknxqGH6l6//VrKxkEElof7
o/adHQecxv8lk+/XN3eQH4sV1ql64oDkgica7Uj1koQPmoN4e36zAFlJQ+RGjdB07JBEcp5sX3Vl
5bX6Oq/YB5i2MFbVPf3fVQ1npH91B709z24c/vUWK4P2rD3Gxy3P9wtToWEL6UZp3gOwEzFujumg
91fUkmurU+yq7pg0EvVd0n3eoYYrIFsJaxiXfm4y8V9KuS0WjHFaWUEmOiqJTypBdxD6kQ+fmDtV
FSgfPIs26QJUU1lscoCjBX00LXbo5ow6oY2J+6qbPd4PEGAvCqGpgYN+29+xdev/IXHjhMCmP/mc
v4BRhu6oLiK5ht8KnEExmPJp1Ai//jn0Lugp+4wICVH66F55YIVSA+zYANqISgl2qtjVkq3UMtCc
epnrpMEEzH009k+Lma0wP5WC+J544N+77JQF5cmWaIUo8rfZN2SZXGxWUaUc9HI7LLZiO8rmxzuo
9IkQ7SBbp/ontd3UH8gW178yXfRKbagyQxjn4mOalrs7rHNZRKxPnVoh8dLw/IkyFLxyjNwvz6sL
WK8vx5/frmHkWmnEMwhmgo/p8kVUx39dbbkRB8s2EeIneRyFCeVIB2kWI8gcV6vdDmnwD+F9W0UI
UbJLRQxwxCCIfg0phs++XxKnEaP5S6wT2r33Qrxg2X7BsyFvDYVPpNbtESq9XaYvndapih/bkL6U
4EmXK5KCxCQcKvP2Cg5OXItysTwbpspiJ35myqc0HoICeSnks/5FU6mJIcbHDCzH3xF2L/GD6Dr9
S1q++bk806TtWZNyHTiErhaWyGKF1VkvhcB+m+7qtopn/HRx2VfAtTlXiA8ptzRnE0CsBk+qXdEL
jbY9znwznaTFN1UzXiT6Kg86gGfMecDLvNBvzC6CN/G5NuMkRsXu2oS+7BKqQE5mSig0HhrZRsur
p8ij8HHkxb/eHeQS/k8eI7hmEObgM6EZoCkWxYCb+BBz0swlK208r0XUZM+DZQwfk/QPRC8DTvis
Q1r8GtrznU9dmne1RuuSNBJPFo4F615oiE90v7InVbJWdDhAHf3mTRCw5Qm7kL8MPUR75cQLbW2k
SZvPg9OuoFFCYmmqKFNxJeEKy42XssYo+K+QNtP10gQYt2htmr2FTNM5hbn1KwTJuUPyYzBTqBAC
zJHlHJhLH3O/oxJUl0rN6GCAv2BCgDAetcVS6b5OQdHmRF7eobMxvIpiWDuy7qeOV9JaLIYIXcWJ
Yupb1t/tiOytViU1x/xMq17XczaCcHZNPxZEPRXZIyJdHb98qRR+IiNS/agfm9pSt7InORmVOFtZ
mbSsiM6+q1QketMiToZxTTNh1iMNCW5MVy+UZlOGb+6YagWkWQ6huv0JRehSvP1tfemC/DmBWudP
i0ZEvstOVqp9976nFWG7T3QUCi2OvjJjIiScfi8x0aTOOJYnyZ0W/o8QMHxW+luENzCei+Y5TJIt
V/J3Q+l9PVuxKEAzO76IC5vH49u615xCFZm/VQIfay6QeMw6psIrhVFePOCBsUd/BBWEh6Gc4Tlz
M4BpsNtCD7gkN2sriqWKqefsRyHlBmLtmROEujotwfRDkx8AfywgmM0F5bVmd+Tvs5fa3NRbdalJ
bNfSOvSx3JHXCBQ2ffsFPZ/0FmNCpG0au2VA6XagxWqaVZQG3Pcf2UUTQybVlQkXvO3RRSsk2qvo
ERVFbXTnDcx/GPskxsNXFb/XO/U4Xb8jo4nQKQN6ItvpOK1OHFxj0Qj4OgcQ9Nd51ORlUD4Qgwhw
/dEc8fC597uWwbru5RdmhRdUiQUYluYpYY2pEEjaVREy9XFMqK1CLbcI5FfJ2mGpesal5NFjbCjz
eWyFabpsKj7hNUjwM1fuQ29GsmJcSnnrt4iAOZhR8Lz6k5Rsq59IBQny63agwb0GeCVlENwc8ef1
TiF4dVNGyWhTwgaCy9d+hDkV1pkIkOR63AgI2F9LBJ5e9IiFVf59hU3CcJxbxxyVBTLCM/5hbhGQ
uPO14wr+EjxEVzGfoZLEd7NVYlxt7g1XG/JKRlClWW+Gx17m5Rx+SZsNFzUqwqlhQuhV1PbsJHlC
q4c3kcoIdzsXn6k33viBYV7JVjNGLyeXjyIc1R5jvLTUUadNDTyGAJJOXwuaIqhPN9/SJyM4Jg59
9Z2mPCfSqSp0/fpBSRZLKTzwpeSvxfveAYFpNxNISOkypxXErgf8BAlhYySTDARhA6h9yorC106s
N5yw3oTwqHc1HuVQ5o9MUUwZDmPucrG8ebyv6dEzkV+6Wa50RcZ+ng9MEiZqa7DoLTIRv1pPxihI
h7ABPuFVoxN91H5Ukdh6CYhRP9uGIUEzS6Lc/KL4KpMLl+kqEbyGLLsDfg9WTh7dXYZCUVmVwpNJ
VDRswqcGWls5kU90jP+tz34Tj16PjJPfQkGPxaSBp1UsfdDYYnMxjsPr0WnEsEGnW/fkUecY0lk/
hNy694SD0fy6YQBEDTjj15/cZY0DvIrggrf9e76450qmQErB/RsT4/C/gQ4KQ28VyFh4diqT0OiA
3JkdGEvBnfRXs5k1dZ6VSu1kqQaBV8j3jA3ms9dKAYpqiCYHhRShob7B4AfcU4Ke/dVf8ZN3XiC1
0Qm2vbw2W/Ibg2kFaJMDaSILGXMgXbkPLLdTDDTedL2P92WnUCWySPtciiFnt5yrUysGm0Ps6A2s
30XpWNhrmdDiO/LiMdVnqp4dAa7ONlyAhWRQK4DMCevDPPBJYeeArLzGLECtKK1Ifg33B+iEcCFJ
hgpGzaBAbRT6GxvGrV6KHJqrnvIqN7a3ZhaX2OFTLW/mQZyWEu1HWas6WT318ZNFD5j2FmQgUSjO
CMjTMEEjCdMxcuI4QFaXlZNfLUwruTHFo2h4gFTp7Mt0A/5N+46QyssbiUCMcZz0ohiwKVpQx9U3
HCJ1fMfoUXNCfDGpFjsuNgwu89fOYqnzVJYd0L0WYdQW8FeSqeU6RwPPFP2o6gJqtDaUdxvXi+X4
LOQfgVGt7JtGrp8ySg6sP+9XasvBzCdVYoLfTcmrJF9pWDSXo0OFo/UToBi03B+QHmP51OiBMisq
o0VB3baYHKpLLh9G0FME93sGxGQg9BOeNoNIdAQMEpGTGp8GQtTFo3pokHkrAE/2xbukhnOxuIcZ
xnFO526fvciW+PW2fBhoeD0vs185Pq9L73qaiHY3b80asZXz0CAr6vV1y95S7s8wBbXJPVL5Ucx6
Zd9WaYZS0LkS/LSBR6Rkm0Wo3j8wwkqVEJX+3m9a0Zwvi4Db2TMH5l97oSYyykWP9XUcv+jyLSN0
rNeVnl5bHOwqFeH2RHcPBtuSL8lKL+jea5kPk+774J2Ffij2I2KuREeKl1kvw432xpAJtRpeMHr2
swNTbx7oqjzr07bJfcUKM8lo4IUrtMGcRRJjENqga21htjeQgWijW0IjcN2SrIYAGv+DgyMmN5jq
hK3SvLdIuAX5YsjXmLLWKuXdniLpb9rDhW5jd/H2ypHiQaijRvIN2YS5Au5hNL0NA6XDXIG6PCV6
K9XRrZHZQkiphMPrQMvSlwJMZfbPeDjo1GQgIye5bWxzXPdXFNTiS/BVsoVZ4lIhUL0AMnMNi07H
LoIVYiL8meybOj6oAHRM8NuYAG4rzHtdb2jIgN05V6OLiKY0OpT2cU/5QV0i8XplR1o1s4rRt45t
LgEN705eAzUTe6x5KKPeELtixlm/015Q3oFM1WPBe6jF5bPTTZWx62maeSiPbLkxBvOXhQwAtfAH
/GcmdY3dnNKLXAoNkoYfsbWYzjiWBjnHUPTUSB79w4jf/RopqOVS7REHq3f9VLOXNLL2VCAmWyzf
CCayXEfoYQ6Gs/NGEBAXuKhdk5sX8txbU10rbp14H7yfjbiVDcNZJE8JzCWxB0/6cp0wM/AtTWct
W95wJhwdTk0g3wdl6LfszdDH0+yaBRmorKayWpQpO3wcKZNprT3S4tzuIoirYld1uZSK801m4aJS
5M2SAmvmXy+WIeqE0IeeNPmk95xz9PuA/tcs9Pp2p/t0eag5R45Ys7DdzF77VTbBm5U5gY/bx7r+
vwgOA9/sWzXuxlQL76Epx+6WtY8etarCZxQj2o8+3iC2aAwCkspRjwS5JSudWNkeak1Nj5Jj4rwH
85T86e7ILP1NDquR4907/pP/430oUKce/plDKXvLBdMZOg5IG4JB3/fxGlp2nEcfBd5wcEEfnV5A
5M1MvEogL9EVK4lokvI07Jrz7vcp+RLwH2CqlItMTW/XVZScVJWjSCMW5GbqLwcvXsU2EnhEFGoz
z4h9KwRX4Ig50OGJSnNLOV3FR2U3ZMOecml5/jxyiw5q08nwq7NIvL+NdDfmVTggKpE3rVLhNFK3
i8bN1IxlejVlFxEFQzoTLPvavCeHECUTk7rriWATxcTXwBygSOISRQSMLGLQImeLDabNkB77ymjv
8UnH5yANwD4+QenDAvB9g+qPV/x4dcybbwKCnaNHqOpYZssNlPPpiwnns3kIi7Bug6k+DFOqHpjG
sJ/3raHYiG0J20cMCbPY9qwSHLOGqo3M54m0+Ox8RA96PHNUCStPHXBXi8U9FNE6toz+lZrNvpK+
EoAQVd+jGChHcnH+OiafpEsVr1Zg07WSf0G3oPMLaDiaNTX6jiH3oaNJQZL4jzQrfrLVXib7ZAMK
NS1Md84eKXe3iCVchTSS9ZgawnfAoQQLI0aCstTLvIo7WW6LZ2W4zkCOC/uShNAcJXqUC6/x+yzC
t13N/3bilXDP3lz6MW1RI+OYecuW9CziGU7M8Ip6z4uwTZBE9xLICHv3Rx2VEAdgRmnY74j+5dkA
dsI/7Lxe6Bv4DJ+90pQ/3xbGAmKmvrdtPIeDBchQl823jjFnR0ywRrxvNT7HB2lZTntJF3u2W9E0
MDbHegiuUd0v0fGEUztl9++LAWjw1VCKguZpr2ZrEk93LZFcjUbtFMqkPNeHtQVLHSqstHmcKLNG
VV2ixZ7J8vF28bv1Py0GLolv4K9di5/UZXzsZo8+FHXsjVvRsH7gPowDRvdO7EeTt+8P8aVpeBRK
xGzsZ09yLdKtX6fx9BLunByU6S5OdJQS1NK/pyr6FrgPCCc/GD0pn4c09fhxszVg8t564k1HXs54
+kDukZ7OUPmmpvorqFtpKsIczwmcN9dHHQ/RXXxh6Hyggf8VLGD34DJIBwWADdxFbyC32+9C2fPI
WdjOj9nRH/We9T1me8rb/Q19MjY4s/oukAUB0/gLTnOfNs3xTZiM2YSXRBXainuGx/NW39hAnx77
K0e9194qOv8opVBJTbXA/lOTduI4lGRuf0KWcbSzKxKbN+qFERowLqxfJ0FhLx0n/vxdqZGI6lrF
jOx0FxoG74SexROsQ8NrfC1cmLMm/wE0GObbJ7GnFK8bRJ2io9LHgBKqbGX7HFWAfWK8D1jz5m56
grMYHrHeuqao3TEsf4ZpsmsLbpXAGijBnUEvhPuldr9dNHv6qOC5fYlJMzSPtEbfKzQnESDx7IfV
0oS8fJHR2LF/OFYLtGfKAUAOtmdr9ylKl7ijWd4xJktazh6CbN6P0NCuQQVf/gOuJCFQo7dsDp8C
DGT+ld0quiPNCpgMftQzNip9TLwR+W5BIEJleJD7w4frcfIEKjJH+uQF52UhpStIsGbWJlOnpsZ1
VN/wJIB36K+IyD74gzHIEc2X8Rjhn/oIZmg1AWyyoP66fTAWmM417euqCi644p3z+ingTi/+yPdd
RFPt1HaxMZh/y8t3gd7QK4HLiQijVdzHPkzhc11ygC8ahMZnWyp3sqc5eIRcqtjPWNsQduhotcnE
ZCPUq+JRd1caYDC0BCky3JJAZD/EJKW8ibdSdf2YROJDkO0qGOy09f/6JYzSUjbTBDCJg1UHogRx
/nKAovH5IWQH3RVX/Yt1I1M686RxOSbk1roq394N3c88U1HP1izufcxz7RtL/rDeZWm4Gy1sWlVl
zYBck5ucrPYE+hVreQP8KRQ3QGH1B9W/BDKeGtODC+q1tn1AcZjXlBKIPquSfEy87zrM3Zc3beYj
eipYNr3d/BIKbN9wOANRG8LfsRJAGwDUgJcYw+mhN9MREfN5mCRrucTgrmikpMqtVgBu0kWatHgX
whcDMimqycnmgP7/Vm2piUj3r1fTjealEeV8uDf/UGj4i+miWVRvIm7Q/Chl0yJdiTfmDezldF0r
RU2Mx9tOEaFfJTarqvJ4bGWU6OMZW6wZcYZ5bCjA5ncpNNw5DfKJ3OFB3GtTTgCTNW5EziKnYoUE
4ckp4Kc7lb+E/NJt8sc6ahzedg2rrEa/S7DUKQZ38eLNn0p3YNIljcfZcKMULVVSFTecUcDK2NiL
SBMrqWjHfLd/lr9ku78OpbVs224dhpbRPLOUT5Kjunlr0Ro1ITPQ4QBn8fDwfQ8+Cg7hdE23xgHK
1LekbeCFoSj5WXTjJNmcXG2d2Je47sJyjI1wDASo8ka0CaWNnr9YQGBSNEL2AM23JLi4yH5ZS31b
ktd7PL757S4b/t2SGQC7lerofitDvGVb6qeSTFSqXrfutxaXQ2kUue3aHHyoAicfhLw9ya6WqPAy
PRRLfs9kj88WiGOXZWCpRmOhHji/vhfQfkt8KGnXmJ6GJevP2KYbA+kHyj3uXFqgjUXYpmPk+ghF
gw5OlAzB36AY1ii2byCjRs+N0wBWDwKWvkXWxcfI+I5yO1Wa4SXcGl/IRsZJy7FedhqDRaGvpJRT
NETayNa2G4ZfwIUYmchBlXAW2V6+VBVaxWqyTCTUYzuiGqZmAC9nODzYot1vy8heuzITFZkHS429
KQ0MZJkvTI+061aEQVaHgbyiQKBH8rmqDpWqE3aSaiI6XKl+JdO+mfAKwH5bKXiw6SdL+02sF5Av
eDxwUB1aiDGyBbTIIkQ6p0XPoyjH5pyFo8bfmry5W41N91MwG3mAI+ot1QWhJnKc2Hqrzn/QnYKk
I3I62z65TA+bmh7KVDfQlwT705LiVD90Fk3SWdvhdSwMeNl2KYnhe3D5WqXEq2ILzmyXYuqtE5DD
+6Ag8lusDIZavU74gGFMU1TJOl5jbwsnEf6iWFHcJ+0LG1HRkXTfUjO46eLb85h982Y5TYPyhz26
zf2myVGFyWJVDiOkgNfrLKNk1K/TeNp623H1BwWBFd4qquVChaJzpwdcpHIvrHjjp08lCo38HVEh
Nwa+PPfKyWEWLXZl0TGI9fc1nMtNgEehLpsE4lW3LOHdw7/7QFHqa7Fg+3iSlh1G4j6pXKNvuREU
vLmqiqa+J7iDI04OTi8vvxi1u4rsTOjgbvSkofYN8j4Vl7ZI4JBwueAE/S3KI1YIPBu7paVwp2wY
nmCkfqqJd2LYO/+TpXFHmFNwYSV2Ismdjn46HKpQVfhkelT+4JDSyCwiSN4xBHSrc6l6jvjPkbjM
k7bpuh9tsBnLVjYun9fYlQmFUCFS9a2YILw/konYJ5T4RjiLNX6m4VAIX/9Cwjt6PnnLBvSG4Ybp
/o/Q8uHZ7XkFdt3rJeIHTCHOndmm1uYag8PhaDmueWR3U//h3nC/MLn6hvXnBGEF7P5/vmd0mywX
4OZcfIYCmYM61zm0q+PLQ//AQZ3id453P1+d6P9hIu/fVCd0Udp1nne8DxNPWl+DzidjOfObs3VL
ex8r2jVpWCpliwb5ZnX748sEm1MZhjYiA0vv/N0bOZpkgvfCIWv7B6sI2GGgy/JS3+U9ogcDcoDQ
ETn1fuxdVedVY2iu8lw3lSQ9ol//PvvVeaORoksMgE8Nw2yf2n6ByuThNMV6NU5kQN0B5IaXt3tx
KEyFf//2c+3rRaE72WEDIGiNkszpqz0FarBb+CqEmAJhgVgpvEHEFRXANkXdEbS1Fp4tlrgyiCLo
IWnZGR7L516g6yRwn1o8vfn/Ipbr4GFFi5Yot8n5+n8b3wdl/gNK7epJc8JV9t2KV1X7cU7eH9rI
kvXYijz8p75gZ0bk/5qKqRpY20w0aaQnOjyHTIU7pg96qPRqVc6PvUN2PQBNzGLKkw7t9+cFMIeZ
b1lTelIYn+nhGrE75vXS56ygrJjyG1UeLGLNJwwCsQpBZ7fuVLFfAJSM/cgrga13J7YyQLRylkGR
xgLlkQOnM86fomqEJpKbcLF/SnZDezlIgqlEOOen6FhEEU60vf4eHgwC35fBsZb4R9nfk7iwquwJ
S+le64ndnimEkvNlzJSGC0QYV+BtDDdEjH4Cl54Uq3f2haKer+vhj7TpDAhqeX7OLic/wmhpiYVC
8HMd0ajpENB4+xESbbiXsewhxipKiEWhtdmUwozbhy9OXXP3L9kiLKeary6Cbcwa3/RkBDXBI8Si
Bz+8onGMu1PfIdZm8TdeQyLMG1rfThQgECfxfAvSdPDQ6vE8tM7keRWxLbLBSjP0CaZ7QR7EKzXb
ugJCt7W+VWzZGy5n3Co6k3j4jy846YjhuyYn0SBjavHbha1UnZQfl15V39ZrOqoUGp6HJKB4GE21
8/sCm6HfAifchK29hi3LJky+rAToY/beh2pBiNNdL2VF4ujlB0BrFo2No7QWgTx70ywze/oe3Nuo
mYckCAJJMpDzyai66Hlmdl+esYzuYl3VXyntfQu45Pj9Sx3fr8H0SVmAoISRsIc8TdZ3m4llvOWY
htlqTchUptsGpNtLRZU5rmuYN7t4XTEd+XpcrjnYkagUjrg1/WmC/vkbZIRC6Fm9cAqd47g4qAbY
7swH8/JARrWCuWfZPFiRIWDMve1RmKfa0Mpoogl9ZC3hEPohkidhXExXDFWB4l3RNN0AajEs4axa
9fsHOxhaFkriAPcmTepHUIV+zmfZhsqAzYpq4synEmK0+xktERG7yXnP94SX61Uyz+XLReNCh58g
1RwxWoalXG1kIDbOpbqxp+BeR767EDm7FwM4kxO8jiyeQCOcO/U7xpND2SjOcboTVjp3FHhbJj0f
ESOBDdyI/U/jrLK5Z0vHpSUWdc39tqOUNNG0dzZbkM995GNdz/tsemWjbBVgr5U/ulAFVNFqZrFY
JmIKtN993O15RcfEX/QMEPzrWAjHbi6lRudOLSm7S7JN12hAfsZ2UTNAJWCPH+ritR9boAvGZgj6
2VBUukwCjq7Hn9MN7n/5hHDHjQ3quPg87WnleeGriXSl0hKcT1uBa9IaHwIb5oD71xjS0RCj0Ab0
cugsrrS9av7JNSDUeYiTdaJPWZ2e55Kjihh1UAJReb4cw7H5g+lXTDKLvAL4lODLs/RdbM8J072W
7rk4XXzU5LnJS/MdB1OId0o74iCKWJZ1lINZdK0d/6XfAdhRArUd6u85EZX3ZjtXkVmVd/1o2eng
Egh+Hbg68nuqcFk1HESsHGeZ2ZPbUT4aEc9zIRjtFEUA7egn4NcpG9II/i6W9WwzVLuTlzsz0nC8
Zne4xKbKo1VM8cV4FnOOPlf/dc3c9pl1u4zsB47PTtdoyUN0LJ+RKul5AxPPC7h0RdMjr1y/M4kP
iG/KcGKu8pZOudomcexQ63+VIJdmd+if25/i7hIcnq0J1epPphicp+UektaHHm4kiu2EcH0vLsir
q7/J1vdYO+uUuwD/3cZNCU1QIsZ3Acw4rS0URyrVI7QD9XAyvzLVsCAZH7jITL4S3wBzLrmRfZk7
kxf3ZJdzN+t5quKFtP/LccTG9hh2sEWhkQaf1D+uHih9swYONphOPrIzYdWXsAolh+B+x3MAS1UE
cvYOeZpxLbI0lkfsoYUy19m9Yxw5wOV1QgJq5x/3o/g/vq0R+vdphLmmCg+CrZmph7TksS0PV8iI
mmLp71EUy6qnZa2G6iQhqFmWR3nvrTS0b3jeyx3rel0pAomB656gXM4eij3a/xRQQD75QFc16BLN
vd8tVJxw/cy8v8dl5ohF7gZPWdMik2ENKibTSK9km/tqgVHR91Ub5tPbibnH0Dqd1xVbnQFeOAuD
abfZvND0lD9/EeyLeXG5W/kuy4iNBs5tHLI/XFjIhWkqNz3S9bmXk8xNryF5Pu03uz/zjcltjY4J
E5Y0YOevrt1GGp7bNZLaRARjGDNVlTE47DoVj3YNcU/cP7BEkVr7T70jBro+nzDOyZYPPA6JGAM8
tXIqFr4kCp+rNQGJzhJzYJ+lo4kE2j9rjcpYeEYW+JJik5gtAdlXOeuTR3KDVRo6jM/mlUyNGu4f
vsgYbk4U2eTpknUNh7Uu4BzxTpvHWn5PkgcmNszgLxhydnmLXi0pexCvxX4Ue33LKDu3pIaIQ2mt
6CDC02SXk8rFtLGrTTxjeQeoGHG1Er+bfyd3dDtOJIOAYqI9vFlAa9kihF2rZ104dypzOiFLUjRS
1hIqz8vAzu6ZmthRn9yWMIXpl/4GfruA39xSscBPtEeljX6Diu+yJ0zQkVQ5nUkGZZcyVfWcFEA3
0MFRgZekmiIfV5eVX01izZYFvWARo9MwTVxHC0rajIxTabnWWntjN5U9AhJa1yZvh/6jByJ3UyrV
kRuu2a/TjGAwfCS0Z1S+GflRf6Lgprl7bwXr9AYrwelh54TtMCmjBzzz6sDRjxh7M+CFRg/M50r8
SYoekcKmg+rrzw8SnyU1JuFWCW/OHPIwrM0vDBOQ3KSRXQaA9jV3Qmb1W/2ziDQTL/AxsaWpvMQy
qqin5yDBNbUzPWK2fn9shHVTGA9alK9XyJK9zg7fCilvU8M/c72Aq5MNTT8OtjRkVZeNeuzrfttc
bNoAlrn89/pd/IcPcs0PgNJA5ylMEcMLoA1WX0iL0UZZGNReDCCu1/x6pT4EN/+Lb/sQQk1DPe5J
7m0eVCq8L5D1Wc3zVm4i3ZvuNm2FIfURHJsrDuqR8STuSL1/uFF2DTA4oOEVjBjsvYweNq/M9oLc
SKX9q98IwKxLrElXY068FDto8VpbsnwaGSk6T9qufaHkyo2+r60eBvqrEz7rw2FNkdOdHtD+UZ9v
VdOt4w90SV+vpywkHdo8XLIuZj9E6yzmGHZ6MC6jGQMvdZ56CnBx0ooPOvFSWU0uTByetyR4mqfZ
PYodq5c8HJFoywc+2JcT3u/5lSYaZe1Dd1IL72wauvAK3TDxo2/KhYpR6jIeZpV2vuRcyA6Yprqv
ZtdSgYiqgxGgYZyapsh8//UWjUQaRWJ5PxbnUzCtjiGkp+aHebNstU52hYHsFpdwkC/0g+MwSXNF
yJfQ4xeYFy5J3AZgBniM8bqL2vQUmLzPtIle/Hm1fPtTMyxcHYrTINlA2MMH/AZFgH9VUFA8tyRd
9RYRnppji0WZ8J6EQHrlEq3aqOH8AZO5g7Vs+fYObWGNSzm8N14Hlpy8xoMxkgjgRzlEeOpN65Ry
wPxlLj+dmw3Oit1oh/uqxKHPD+xoKvT9etC5RU4ts4jqRtMP/JHigPR13MS4exQ1wsZk7RoTTjYi
fXtM1Hdd9SwxXRpQscpf+N24+ZDhBrfAReC1wKzwkAH36UJIeyU3soBSIw4PVG1erozK8cQy0hiC
3q6zMgANTu2RA/UiScYysGliDn2+eUgSipUvRl1FuBK6D8EzwPIZ64xCuBrrupM29rVaP5G9MbmF
vKsFoPu5beKF1a4ws06NevdaJCI0dZLirTqo7EGQ5nJ67mbKQGn+7HA9CTEqoZ1UXt9PnH3OFgiH
Wc3Qdj5+56u3EdYIYAwJgRAPaGE8ERqDTgHdef4c/U0o4uwd9GLb0JtixSRlAY+g8EEy7ndMS8C4
eS3qIUdTqlpTS5r0V6+XA6JWLcm1SKo99iaeo3XQf+pn1GN644FEKSjaG/d/obkbP5/llpfssyKD
rCM9CZ1v8ynCnl8VZOqPxvw8RL8groK9eePy7I2aVdgce/C+9RVCEpYL0fxXT+0C2TBSDdOVRbGJ
t6LL/xYzaokMgevZ6XDDra+ObIocM0U2wMJtyvPcpnqmnFoetzonyXzu2+GNhwCGVmHTwtvhsyJB
74hAP4/Vebf42lLxDeKdhHJDo+KeOHwK8xofsXCin7vD7PCGbP4PFd5ZZzPe1ZWakbccej0Kk57T
3yenpcl3PTDaW+ir6KcYY/JTY297NePHDyx4JphhOorrCCz5NtryQ5EiufqiHiZKhPINa851amx7
HgXZIdPzjDjpRjyOBhUoH5d/qPW1sps4tCre2NRLWDofuSf+Rrup8VY6jEyMKmQvK5nONiLertZs
6CGEEQ55BfZto6YqqM8HZER28yU+FAOPjPZnNRldkqHGmCXNI+1pbFck4G03kHoH9PdMae58pjZY
PqZI45q7fJ2WovJ2dGWA5lKMZpQkh7SWS7Z9PtDqGh9Kk4H+yDegCTQ8TgOmpKGcb1kIZ4cVBWJB
azupYjkQskxD7NtDPNB8J8bi5Xh+MT0vvE6TXTfVahfy5h2dC4cfSC+RD6TlEA8sA0JcQ5wL+pJl
WD1a99JunRPLA1AqjL5MSXZ85w+eANwLZU9hG6/yzb+9y5W10pPbWpAjpp4Bgd+atlv6GMBJ5zZM
AyAxpq1s/V6KShxe36tU1r5H5WZNFg4x/BRiXXhxVENklL5aL+MuTxxIzsvomD1faLDcQtmOB0T7
ht93cuKeTXL28v8EZf5iZCA8ncvZuvCUV4Fv2HAB8tgCCEM63okesB0w0qRa/PcOCUTbprOc3Ogv
HFz5MA8dd4UftwfqyUQIK6D8PGj6z3Cd4X9B+pAMoGg0aXUJzGFfHDlkEBgxdCg6xJ8QTOFXwh1M
rh1w+xECofVxbFLESCmIBrHuGfv/i6137N73Q4eeVTnUgPHCUQhxAf/kW04zJprOYp6HXwDRUnBu
H+uU3DiA8zqvGmmYjFhGW1NpK7/ls4fwhFxDV1jp0/TFi+Jo4f+r7+/3qKlbQAAp9lrKdpf+1ZMS
1EzEFTSm2Wrhxhye8jepM3jIP8lmFtftvevbxIAee3mps9ycGQorNNEy5qcaTPbMzkq4KXh1VjZD
1Cv5u+wxgundAiDmh3zd9VxuEi/mw2KwhUuTJxLEQ37nlkh/YTVN/IoKGHyHjgxG09qZPQH8Gduj
qCfhNe7iQe3GJ1OFhdOoKPRsToEfcNqioBoR7CUNHX1rwWZuNJQH//WI96imfBITpkNhfRE1Qs0S
KFVTw2JV1rWYvUBe9MxF4Y4JCoLwThUA8ZNUOISc2XVZDvKn2WNZEfpFVzskx4B/ieE8qvnRyRsj
i3/PFmK0R3e35pV3Fn5uTW71ojo5NNnq29Wid5R0Mk/Cb0pVF+5IgkO1hc6VvntEWxVrNYpiaw94
4sjsh8jpDQa9fmA9ZVMVyvdjbsPMiJwP+CoG0wzN5zEii2gxkdxgVji//roGKSCe07s5nBZOS4c7
DZNKfac7NjVT01gLVvqlXmXlnVKVXEFOSnCyq8KgfbIZYG4BMQGeL/NXoZSu+RkWZAzeo30FG8Ro
gvzae5tsO+m3F6IDFug+HMkfijfh8D40RCP5QNnEDiCsFIG/WZstt9DuFRvl0IM8k/g8kzS2f0iW
8+2TtTFFra4vTzIYzZXSO32CGUc9cd9hFT3abxCHjn1uOlHKCyvUn/fzg+gF+uwTrvwYEqkBE5ti
Le48sZ22pC+W0akFx/fx4Z1J0PM+bUoaARzjkQkOen1CzCNlu6nMRNnSgseetBJqBDebb9yBuxXl
XZw4eeSbmIYOiiijgyeR4FIWe4QGy3+lP5F1f21HEY62rBbZR/pTCGK/pN73N/V44wWGAFclILEG
n60reabXmE5URj801wSenU20zir03a3BQ/yZ5/KcNsJOOV2nnhK3NCaC9wapAGJSzmt0m9lfuWaE
cadAHB1kT4SWy2yAIqSeH3C1W0n/GbvqKFp14jIdFKkJupuAxKkHkN2cJuj/siiLf9g/7Eo2k2Ky
v1W2OVp8Hpf3UbIoCsA2uPbJvlnF7K0i+GS03m6YloIJOVFZpENngTCpTGR3fvfarijrxUlLYLcT
KjmdLiN6uN6NCci6a/Rw7+Bl/b7OX4bgNXpakumMGuq2c0MMYtzx4Iui9dxKL63aRRYckhwqzKrY
uRBjy6N+IIftG0EatlX6VTdzlQTwpzDGqyxyNoNNY1S2i46IcYV9iZtMbrYCCGPRo/dOxZcAB/Qi
0+BuH+TNx+b9ZzGfVaX1PhnIrEEHAU/kCLIatk/mBaLHeC8PHGAeoxvUtrqao/HP93teOpiFt9rz
PNDTQdMMKHYd80K+N3W/cf+WoxJLpGNrEljzy0gAvP0tyLendLAXEHKFLGAklBkh7v3Pwrqwmq/W
EQ4AC9zZfZuEQWpiJ6T9WT7/GdqWpIQibBSebzd5BKirXMEMgxjbNMiSqNuY8XFRYOnbjj+fqaHt
ZP/W0CFWD6K3bCHkOMkSxo52hDLRtFNOvJRHjhPxx764Iy8k1Pvp8hjHgjB4YNYe9YsWGz1K+TJS
Tqdwv5VceWsffRJ5ENNgrDYh7rwo8cE4xjgbdpl5FyM6uIKtmuSmq5e+sPtdzKbQjFa33aH/gymF
wYJSdJP5bFqQoMi9ZrknBIewfTIfXRabNgpw/0G38gj08hOqJJlEA+CYzv2KMMI8Giik5da3tK/0
0qdb5sJLK6uTPNwdBaB2pjXJxKkD9SRCB+unBB5NebA1JXF4qisyTC2tTIeTl1ha09LNNApk+xXX
+IqN2oL8bN5U1Tb5UTIRU76pOO3hJPIlxzp0vwQIv/q/3OZ841jvxW2u1L8CjrlvOq8fLpf7UuGA
4apIXjteD4cRs7wU5XvMd9aMftCH31Mw4r0tJNT9VeoPAz/A44sbThfKF1ZCKoXBOhS7h5hXyGpd
6LayuLZ99eFgz0VoWzQHWr0TNS532rRZf9K+7XxiZSLkEu75Wu3lobZ0UcGAoP6u+O52MXIJ+2g2
g9cHKsTxvSNbJ4xzv3T8LTwvCBo6hK5X0RqY9UqOcuWbs0mBnJfM0H9WddN6tc1fj9PD8dLJQV2y
EgUFi6AQU760dgLB+qEA1zF0KPIv2B2TiLg9dqLkkwRgxt6NLzKJ/disGyf/8zzczFUcEZ1p3zlW
rqCpeA8FjpydKBOL1Ef9011JsNTwH/W5RGzxgjlNXGtp63MOntOdlzJGgyNkejHWKNhtBTEEPVA3
N7ExoKvUVMKTEwlY+hZBAurYzb+mJlsyxMPFwdYrRzxuYqp+lGjL6AWLj4+1RF+kG5cXGRu+tcPz
MseHBd0cipkeqbq1Das2qBTUgo/ECud+zhX483yavFPL4TQIR/YAbiLAVvdav+aRtOA8RQrduBIH
YYDezeW2f0TjdYY10qNjsfiHoeoJhS+w7KbbpKG/iIQzg70s0qbk1+h97cLOeTE+XggxW21r8yBt
JEY7V8JAIoZbc1Hj2YWIhjGsdYAhs7m9UO+EV+d7Oj9k/U7zOLhL2/kxYeVCefjtfQWRBlnqyY/I
VK49qrQhkL8qLfUxpljctrk1bAawM7ANOVMSQpxv125HRpYw0r28CwkV3jIBSZmKjAWfzSAe22tk
MID93M4my7QlSzIgSeOyJik4jEJMiJvmvARJHqJLcXVYRhp+iaZ48yXXxqneTe6bAVXqJ3WaXYNC
3yh6S3AxO96S+JI5kEWUZXQzXjGQdxXgFonf5wwBPNPtXQNbqiZ63SgyCeTsC/nsBOr4pZUorbmg
dvZHmB2+BUYnBWgdEFqG3MTaCdKIf9+6QR7qZtRF3WO77fco0LkIL3veO5/xRGg+KYZFyhZO7J6v
NJmnX1QeTpPGjGt5vU/aeuU8OnkGaaZ0/v+Qzmt1T/eXPbzPREkqyhVASkdfYw3iHJ9GbAh3r0B8
PcOLBhzGY0Ql93dfZrU9IYL+jJmnv1aiUAwj242hWqvo4tTAE7lJkJIxtGPjb6UmkL78CJJtvPav
hAZnzFj/p0H7+T4beqnjmGTG64efUPInLaFl11+Ns1y9Eld+RH9OH6qo3OR9ZkPkPumgrETXCP7V
n2tpSN2MqQXyWzr0k9s2CBqxWzruB0NNDLjhapnkHsMuBiRw19/I6BpanTcFLj+jskDWXrs4uagR
NuRkqp8MOtR+SPYuvAwaSnaRZnePMxiZJCZE88PCuCaD9UOCHBeSulX3zx2IBmjfYRK97pCtowLc
zVZjLzb7fu3gTNiRO/hH1joylB7XVciyxzdbbDYS4LmnvfBkyt7mlcKslqcufkaYOgSjO2D8yo2y
R88KuVzo+zJIy8LLsIb96OUTTcK/Yaq1g9w+mqzTwv8yM0s5wbyxYQsPjgMCkRwPiQMeHqM06+no
27rGDaBBo5Vgdnm/VsLLhDb+/JoSs8r9cn94AwdtqajhV9x2qkPmWaD9PSDiT8GntAWbYzslKX39
FziUK7leGvyTl3AWzC8toL8yoay8qgTYEOK+kkLLD+EVMPama85MCWRhgqBNzJSrs24is+Mn2g2i
V/FLxZoqy3CubHpUwBLmJr4F58J9sXPhUAudrJr5Dcq+/Xft62Tlf683FdrbEihgW2XYuagpEGju
ojTU9M4QbvlUccC9MSd8bJm9xCH0m41cujil9pTOoR4aJgjYePRZd1e1DMyDEPn1lkkDnYMbBzyN
vNFuF/TgoaHw7InfsxG3c6Kj/n7Ik0geQVP57EI+71xcGY3uRE5zShOShppmtvEuQEyas16Z9Nv8
+YbbcxIdCfb0D7JDTNgZrjSRcABw3EXhCeQCaV09k0Wo1gV+iwRD4HyhN3e0EFnQVrxCx2wvtt49
fXE/it6mh2THJLN4wUcs+6greOs/qji24e7ppGLwcFjGcZ/9OCx7a3PkbqLzMnb6M3PQIXkEdyGp
cXy54bUyrGF+Et+fydxvZvFlPGEEcrQijG/2LNbJyCfFy/HdKbYYhR0AKfetwb02CwFLw2NDkIj4
lzRWk8ue4tOmKfq/BA6Q+r7/NGGKMhHspCIo3pCOSu/5fomltvhPdEZUw+0Qlf/jmpndxahDUJie
qCgJ/JDJ9CF4vlHKU89vuzbdGgGYRRK7AKkT5OnH8KkBZ5aGLXn3VXSl5matT7E1gtYNnjb3iKRO
oCp+CDxS0E8sBP1MPVsbmeQ6Gc8TidiTj1Vrq6GknX/kFLdexecA2BLS7c9OQGUOlzDtPqs2HIs5
7hYj4AEJm1vSbx4cd3b+hufytFrhst9F4VfQzCSehoGc1TY2ZacEVgyHCPJux3LAsfME74XLp+4e
/HPpzraDh8xNgg7S8bpFVaiuIoBT4gGxiVlBBE69y6HZUW5Xu2ESfbxhbudjW/JN3DzoFcJGsUzn
EXyrRrc3X+EcttpFBktN8ServCTOUPskAKkvF8St3IJ88NLbHSDaU347LgdVgqfUEI0L2uTZU3Cv
MhvjLB5UVdmt8h35LfbCStAecU1dwUITzrXedNt9d/SMLtmvOv+wESABYoj6OU+krb9LI+P6sVNi
OiNK2rfGLC/FHC409zuCga1FLSxHWZ1HGMu1WGnP0cpLQeNLmHbVAS2NNEE+M4UVpqW8eXsMMUZ/
9YY//N8lc328WoeznJCNyFApz2VfAwne5ZHcFYIIjW+IOlcYHd1BqiB1Vv4iLxMDwD/BcKyRY5GS
V2xUs98H5epuMSjHuFkpJSUDUx558YK9R+sI94IOtXxLPVT7xVim5h9aGo8t2zNM473iKwfYCpGx
BNQKOrot53642lQugKsSMco/zZsMNdMnycT1gHw4MJzd0GEBAb1QXqGBKMAR1XGs1bA8RNVKgJEQ
tRQSA1XK+Amvg/Qexb3a/YIr0x9eU3FyoHVkm7xJTLrEY+PTGlRzQ6hGFhgZaIzPFxLI/ZlO3e8O
FSzD7UjPLg4QPUbnw5RfKaFeiayfsyv1Sv8Fh+a1L8cV9Tua046b7spx8fzyRDm/iUlHdBb9V2c/
QAs+ZnG5rrHkr0Y4PRfalHxXlAL1UJHPnRTgakvlh7AjYxOF3+x9AgVZKATyU7lcZU0r48cjj9N4
A9HNBJE3E7H0yUtNv8gPr+mbgKtSyyjw6MbYIpDlr2hHeJ/xGSO3JOSApYD7tDzonDvp867nrub/
se+DMXEdU2yHMMzl4exbT8BJt+Omh7z88GbF/001FCf/kJsQIDml5MhTFYYWWVYUL273LIQs4215
YW6K4pIJabotDKuOs9CqLD8Xsp5rB/nDz1dJDf1NrSpdlW3ECCIKNCm+u+4s1zWCxmikWz+Lrm+/
AKL37PWp5ehxpWuA4J7UJlGC2tfzJkl/EBBJsNGbdaw/q1pzcBz1Z0QdHSWHZHGZlGzKjFUHCQBq
jP+0g4AhW33XjYTISW2angzaPJIuM0/PFEIw5Xts+PWvUNfKz/OxZoPa4lPd8Y89iR2rc+l5K3oT
G8/kfo445Ktcuh3bs0A/5IgekDoAbDs9204C8iXaZ1/4tsVthe/6wxUQX8hiho8QjSNoTOLUImpr
7slUxyaBM/ZfeOwIq2SWYhDwdHJrCla4e479svo9Juc8akAgD0ETG/MGn6BV1Zgibt+BiteYXDRB
qAIQ5Bn2n6LHX7G8H3DPz1CiLfLWhklSxn7zxQNNCUW0yyPgz5xvS7xuEbeDh9uUuNRxADpSimmM
k8acxT7pJ5XeFEChGlf+5e2CwA7vyMX8daMH8rGf0z/fJQY8SGCSQJkYVrDG9iVBXtf4rTYd+0uI
uikNE8DzXbgFye/fhaLlhjAUTgpLo/dOzz5ueKSoZ/RuWeTctJfjiXThPD6RkX2+5RX6fcwOQa4+
ZB9ZoMtK/hhc/WNzsvBIvMEsBaKEhZtnspQbOWJ+IDijbxHKiA91UHE+SDkhdDiCFmlaKHB6cRPu
d+ncB+Dr+F8VVNLjwH6h3WRvUp7Ei98U6ewfRg/Dxc8QmL5l9trLy5LBSYiNVb5cnzejtgrxvPV+
6izjuZOzDr5aQWbyXFUnALuov/T/pPm+IdcPQpNlSVJgNmYT+SKTs11HogR4JlxlvLlwURWfH/Ps
UjFSzN0mXu6jz+2P44Kqj4s9ZUALBd0MB29pEBgQNqEuhfmEsLEyCeg0Qibb9pZpnHsn6qauHNKl
whg4/2vxnO4ZQNQphuEH0OE09cn+7PgicVwvFyXi1lRkrSQVWXYQqeWg66tiPwBpg2cjD+zYG39h
fZ3K87t9+0Eme9gnXqczimWHeyKvjZexHeF5kMDAwoaU6IjtU3jj14ivd3XJWQpZr+DERyTwgBfn
J/EjqHzweJPLSV5fHo3ZvsR5IhBH//y8eh6V59i4XC9o6v0Zu3fmJmeJAZHafVHbTBdsuGCtrJsv
TYByo8cUGV1HH/GZKNcntgpVoGhNlRt49Qky9e2PtS07jx83iDiy7+HPnBbDK2uMIe1xAn2+wMbJ
h8obIILpTjmJoiG+wx1G1Qk/U0iLZ5BVf1OLG4Ae7TCeCVMIKNrS6rw3O4o5XjxHfXtjNBuT7Xfl
6GRpbZ/ca+1FNonU+O47/ADLUAWuR9EIzEzgEbeEeexaJo6NnaY137imintfBiiVokH17x3Jb+3r
EZq0rCGMnl7Fysypx8GiyfjWIDUVLN/sAThxF1S/X16eMLTd9c3j7yfFbxhXW37ekpBBqBkrTKKP
XJRka008US5x8PXVHNopLjlfz1xS92RFj8fK49JB/0kDRuXaZjKMyizsvQoO4sBcClRireoAY3To
591beaoKlPipu2w0XNafD/wJ/W5VapDc4HMMaBio1kcKaHIo8W3XY2XPNnTnELU/jnAYeFZ+boLP
gDwoEpghVzMI/+lu9H2F70Vxnd9pjEmbYf7ACCIs+NytUm7/ov0XBqbaBM0JAhhfiJIJlDeTX/HQ
1P2RZEbS2dw3f9SPLD9NqHBnwLFR0YwWl+3wJrpnbhVyXfE/wZXbrFiE8Va1lx8A+pGDU+yfM9n1
xrPPULWNCvtFQu4mCDMz384+K4umZv4kFpe12hWEHrVKxqWTB59XhRs9E+RLoiQi5+31I2x7cuQZ
2+Awx2/k7oJw7HfovMzOResycum9t+R1A3xcoWT0RO9DS1qDMQ/pTkPDNVFZkHOQKn5aEpKbNqa9
VgEvHOr+FbJNSzClerqLj2JYvzIB4w6Adhp7ew6X7J+eXwGuuBuNkrPa0JpYMVo69jkGsjDek1PT
kbKB+w3uiPUcke4Pf7VFdA1WPLxbOKWtH2HfAh3Ib+vMIm64G7/MuR70vGtE4WCintAFiLobGvjg
Z/JTFFMu6sZ8e0UHWnxREzGoA1nPpJNxrE7c0eI+6QluDLjeeeNSLkzzu0sHWTO02wELq9Cp+nRC
DI1n3kh2X9pntRDG7zJEkRGtWubBcNNjJuhDccXSdqOt0CDx2f72nURgybHLYfl06wNKoP6djMIb
NEpbzIe3R7+k6BEzyMiJrLm5eOSqg/hRAAz12uuYDD/QHbwHlufAuexVTihklH/X9GjFgsunDnYT
ckAjQInx7F5qfFmnPCYJGDS/PBWNYxqeAyTFWKSiZWcsz4WEQAm/fnavolaHd3tMvEEGQmVhcySI
R01eWuEbv0lkWs2O6VwuIC8WAa5y+9dEBv7UN1PxTqJ/sOim7SGtE7IwXPXKk6U9S7Jc3hz3YijP
vRF99Bh5C4AHI1vDSgFp4c2BxHjXZXY7vFUQ7EFUCGx2wausl/3pNWsEtOjqOMkyyB4ZPBI0bDx3
9nrT50tzeE3Cg6b8kcFLN7v2qKk5cRvDFcKu7UBA/VCQdmfJHKxcR8KVYaIZSB6dYaNXzYCAJb8H
CAfao9hZsGawdg9DD/iX9gCxKmqia5ud/y9sRc4q9BhtnpF8kCV++NDMjPBs4rIrqPhnwlmLrerN
NNwoVoSsQtFuUCT8EVSccKrEcr/cTTZd5c/rXTNz1ibe4BMSl9ifv8yHo/DsUUHyQi1z7RUsETGI
JyE9FLDscOlbOddRfogXcV4opQn/EALmiw+p2jeaM202J0ZKphvH4MaqSep2Omr1M/+F47Abw+JM
6mCV3nz8IkHpWaDMMSRaIgKJueqfGXeeRU60kuhaypGGPGLKaG38rWq9BCxPlH/CKJfWbdRFEXSe
EiISJO/8DsCybkym7g0T5HRXp0Nxis1MYgNDb2Ap3FT3PLsQ6p6oEPlW35/bV2qU+kMa00ZBeCS/
3Vv7qr2E83a+Nc7GPgJ54mG3QZJfAM3GkVCS5YI7l7MRSTW1yggSMwfF9M/9bx77FkL+8ng1r6sd
GJ6pWbfAgiTw3LGT24pNyFa+WAY9d6QlQLOnpVf028sFizud3pADVGdCEclz2xmxh7NNcjOA5Uex
8INMXn70LHJE6pjnC2ntsr8u66W81TURSarJ2TgcnpunbbGSJZ2eKBNeReFOtE4YNpUjcR4cq8mM
PF/eFQ4cnI6K8SvapsY/fGDduuQp8CCNcPHiagniFn4FXRE73UGt+ivLk2mSYcJXh1k8BjPUmN2Z
/zw5OuT6q97iJF7ofKEGApXg7wHjVCIdTiHnOsilwlgk751Vrxp4VfxNHcgnziS24o7+go1+8bXE
HMueI12cDQblw2EqgMlt4GzKJeqAs01/2198RUAxAghwDtqhXcvdZEabBg3wIZ3nZyeqScegqrFn
ILn0Ywerx3NqmEKSJ1/RtZEZHFNK1tit2DbXox9CZ+amBrx+KrWERfqNknpsL50uWUhuk1v28zmx
rL4XZIB2A3bEb+5CkZUqsjeTwYXdsPjteOpqmt7UbTPJIPklnc1r2eXer4I5e3GUOcr187uMpAfb
wcczN3QSyW4T9xW+z8ef092x72OEDcL3z1jFbwqWpMOpANpobYh2Z476hnuyCWTx7LlHYf1+24dX
eVoxORewX9tKkknZkahZcq/IdJiUpsNJP4MHyDuYpT1GjQViC6VWoYoJl2JqWTFikP+YSU2F6QjS
D55AEZD4hlonmC2RdB45fl8egxvkjIOp8BWHhFwRblx+KZ38Tc7gBPIYevgHJv9Xc6K8/pefR2hY
NeFCys1hIaJ7gIAzhBYiwhrqeKb7MAc5gwhaVeKkc0qEX/yWbyh893iKd1/j4XI7OT57AwX5zkas
5iFuUJmIkJ72Yd3cJxxnCVU2X9una00knSBWA3dVz/351u7TtRWqRu9PruVW2FohERdVJiduoze+
FPxqKHDVbwvl2UwqBkJ+qdaDFsMMoZeWGp/4gGZrAHJHzFdI62BseixDc/NKL0JEj99p8FLkEJRc
dP4+ppvOCqvWytMS6CqaH4z+DOlmQKJqBD+2kfRFkvYRYt6pBs+3GstFYGViBGm6+fecRBDWkSuV
N0CZHPDn1AC0QWwnUFv+SvRyfd6CF+7MiF1H+Q5VObQaw83sECkGCIyLYZ01ockdISekQwOxMID7
WSIqE1X+y34IJBK0hNFwXmfnBv0IU0QeD5FFdNrUVXPRe0m1ujm748Z8L2MRMO2CfeSx4lnYgRdf
MmXDkeptXWpdJeezBuh8sNsR2Qq2p4Dcs5uV4Ro1ak0B1JqhwuRaPsLrlyd1Q/SJgXbxdktlesDS
BA/QBWUdlLQL4hMbNhyefqvSVWT0uCryGZDZO/xmfu9F37lAR99dEdn/kKtdf/xdLaG9h8vxiyAs
GfoCUqX1JQFazFlQcLynTbwi1L9N+bWtPnDPsUAtJ6mP8xmNY85cbE5X7x8QBnL6CCsFlHo1/Y0J
zeT8TjZ8UqEpNyjmovLzcLFgIjS1n71KmEzqhwS0q4UkIKda6/Ggc6v+SZvhZfOVKHWR2D0v3hpN
dmMi12g1//u5OX78Qj6mzRyHo2rs4qsDTjlK6ioPnID3OQIY7FUg8PkPdh853Iyj/wt2Wsg0iBMu
MmjvFkp+RdgPVo+qmYWksRp9V7uPnNl6Q1qcxEWfCDht3pnTI9FGZjv9ePP70LOvt9NYry2SIqUx
tVZ3KkTfyFGzvLmZpAEvGC7RSeUOoJ1ss7txXXEttvLHOfiMoQpFtcEOrxDqg3HgQCNn1vC+UgS7
aYcuw5ELLgoHRgB+TEexJLkRCNSkOeqy+ILPZCiRl0yG2JvCluqTN5VxEiUuovyaFCMb311HwbyR
SO4WWVniwzck9ixGSMbtZZ4ChOTkUKXvQ77da+kkxBjAnzI3RVGJjonCmJ3xEgv7z3UeOwcBs/LX
Ag33xwkI3++VEW6fQf9ruQW5hvSklFPQhzOuaEcbHKwnQ8h9wj5NC2nyBBXm0vz4HWKwA33ySt3u
QCJlrI3DEk0BWNm5Ov0XR2QucbT95vw816bvsQ+5XzvN9SD0xuKjiNJplwJhp4oc6Eg9i4sgjETV
s4LQB9vz64Nw+7D7EQI6FJ9aoH0qOvYeffS8QQkigQQL5ArFV5m1Uu/+jc/6rGKoeBeszBs+OffQ
dSpBdxgdGL5FA/b7q0Ln1xKRC5qASMzCGS/jujPGyCLeBkbzEedHvw6D4r89W5QyM8aNxNX6jb4o
O52oVA0WyrwgC2f8rVKk1jv9kkG0sgVQOOUbScuEgxrt5TM4khLqKnlhyty6HIUxf0217LcV7iY+
XqZWS1hA1oDuC4TQId5FtQZw0+INMPNidKW0Vh49oJh+u36Z/MRet0WGHwjxpVcS17aHaspeA9B8
tcByRStpA8BlUoyp8wjj7qRGnlQI74hJjYAoYup24FGOvo6uFnylNkYSzkHaJqvM8GtJ3QNK1cVV
/gVS1H+F3UGC0gl27UvFmZ9ZK5sEQmD8HENDSJ2MrnWo3GKu1j+NRNkYxebC2ylLLPvuH2ICIOIX
EEHhKIvpjkmFQIHEfFRLDQQ7VX+O7l2AMoYNxm719MwKFDNa5aT66Xs1oT9PMLLds6jq08R68QKg
NIKZquLdm5sk9nuCe1CKusUg56QFPGK3i8tPK5SV3VE+RnBTcYG+6M8cLOxmUNnRJF5IspzCcM60
JUDxVVVImsMgypjM+CQA7w32qM234jXIleA5yqsgb6z8LMUBibiQ/PAk1dSvPb3GWm2U90ehcd5G
MB8ziLrVw2rr25LgTy42Gh1GUYXx1ZVtCeSav9sU6xB71s7HPz8rhoxRsvjKRDxVpTCQDWcXiDcl
diQAel+SuvFu3YmdPOY3AeVg+owtn0a4ARAMEwzQeqsC4TLLn3B20v0grKzC5nNxjnI60satqg+/
W9+ph/ZfqBd+DVO3fOjfw/lPBbifFg+Y9OfsMSRbdYLUV6nogY8RFZl/VMGBvTPQFbZzDA93ccCx
B213OQcDY0IKS+B25NMENxPQrYD2bIHHH32JGSHr4MTrLC1RZlGgbj03nm3V4zPZ1uAZFV7VcINa
8Pjr4VBRe7uycgyf8n+J6nSEq8FVyIxX1HWaenyyUAUbIWztxKPYWkExRLa6Gvx7na9bmL9Vfaoa
tbx13p4KEcYfSOQftEHRihttMbqXHTWblyiEBHXP0lJgVSbHzxT/1vgWrUj2LOKUvVuUpTpr9HzN
N+D/FxgfyM/o6EWUnUJWIkH0rkqu58+RwKX/w2xMMGnt+9NlZzbPRqDleZ1N3FSgPnsKJskglA8m
g73UrhJqcTVjTnSy3dcVCW3HRnp680rAWHaRrrWUJ0r79JO7kWfrMLla/OOD5ABlHjG2CuW3p0u9
STqN3wNYvjLPCNU64lMzUa8OtfU1nEX6/xlq5iCu9/pOYHpR2cPIfylwc1tnORdLokJLjLcanPUX
UJfu9tiXnNkdY6A9Vnlf2kBoAVdc893ZrwkHqZfRVpcMOHjho5ljRl88J+v53KRKgyUkt3461zGl
vhpKjsmyXtLW/OESX0GO6NCQD23G5Yrfr5BAKRv5+XknaPDzYzPLGFrUroRPPG1jlMrz2ylJGLRW
OIS13AdNF74R4goBseUAqPRj9Y5fyILqNS07yUq21wOreQCZ2BQooGt4fH9KxTHa4rPrZ20IyD10
QhI8Uh+JpVi/Ag6IRsJPg3sX6AqHk+xVLYPv5LbijEZlE237Rda1hWWqUOL5/FCfBoR4ympGAIGh
6iqnXltvSK/6U/4Z6BXkAe4LxFMJae1IPsEr0J8NZSVjheoQizuKFbAxNWdIpsJCzVBh5QJOEpk/
gPyKwSdQS4EPI1Yikr0W60KPRD20ILidbla5DpI0Fm9kEfxfbEQi3QFe4SjetkpNvQ7yztqkwNUy
jJjhU7lMV2vvx/QTy9NVbbfzEWzr7EeCCPwHIc1Rg4vXRaA4grEHq2LZzxV54j4+3NaGYpNZ+fqK
M2dlVrdTYkyQQieDmP48LZ4pOc6QP3D5MqiFQO6H5ayD9ilGDf9N3GQp+09AH4tRdGSEJPMXwwpk
/vhLc76UpkPmInBfPXPpBv7ynzoZ/K0UtX1Q1s0HL4E267JDDAQEUKJx8Y5Cp2hWOPtlo/sIBRTN
2dnFYEj3EHepygduP6FL76VhOdzXR1w2CndLVciUWXnngwozQqVekot7ra2qk4cluNCJn17CG4zi
kjGO4gIO/GdhD/fEhSJRvXJlUXP2B+DqgjnR9ZOwUDz7xcNxmPLoJhSZLQLiakaPxKqtuVq1atP2
EVDpOVEuH9ubxyk5vVVr4TIDf/eYG/DsvFnNAmsrXskKME7hWwXHHHfeX3HQhwKtDi70BTvTX39f
D2foZ5hFRknlhfMsQr4zYNlRrAa3IqGwWxVrOWo8neX2netaLegd755W4G2SOyjGNa4lRBkJPpiF
o/sgWJBw5WKmfUJ94YjPsJqm21k4UINL3lKONQSxtQTZvoDt6iQJqOj4Rv0iMcLUOlzQmpAJNVvr
hs8g0st+FhBNRDyUUccYC4mytIcr260BqC9mRsiJIHbTp1g8ERRCjw7oXk6WYeMfQj8LAgEgwGit
pRA57epRgi1lcuPWNcg9hVZQhX04y0qTU0rB468Ah7xs6Hn1MWBpCtBXzgut53NSqYog+Y9AvQ0F
DcuDqBsZ6e/nVbZ46xri7AvIvgaRed301860fvwMVZvU283xJXgOWkzvJu8hGoTvnqI6+IR0lzhh
tlL3bbTpp6CTehBBdhuX0paALIN0wuL9uWKjz1wGG5F+LVpiwq4/iqqsbm7nsInb6ydn8ZRrctwa
M24IOHimJ91hwIj0+8Fi1jwnxhn7HrdFhhe3K7XvsixTrMYv6v4Ww8pp8ukqGfgnqw3DuLDeFSTO
p8FdBvLGejoSkOGnRms12ebObeUyivrc4vkjn9xcqPFw2k95Xojn3nTmJwGbdkSJNKYxoEZZ+1oa
nCWsldkwPWWUqPTzs3w5Oa2hNKTd+RBW4CZ/JpprlMMnaAjxsjGsBOn12GFqMez2tL/NZhs5Qql6
rsNvzzmKD4MwPZigtc3Vt1ueikZPYyC1t1GqB6VMxtADZIMyjv98LCVEoETTboLCkDBExfCBN+B3
6BJzza1yJ4twDqqvdLsof9/85uF++PxWv6r29m2OQfLb691wirTuMNNC5yp590xyKNgY/+ZwopVr
feTyjkKCMGOuLqWAlJf0fOjXdlpC+PIZs+WEfaf0ndMNvsOZU2/g06TQ4u8mdH/cqM3bwsKN2JG8
HHRQoALtU8ljuOEUqNig3OnJATUlffkJz5EnCOvqqx5llBnifG4ZYg2+6BUpOevWfC1v6EVggcZu
dKV9BavRqqbD2y5nh1dhneb9TkgdjSnX7smod4CafX8posWaLYPMRNB+vRAG26B0j7RJrIUHrDZ/
B7qTitPcpTyb+dFmca4jtXsumDqn0gUFWID8ofZvVGbCwA52U04xHBBIS/nMXFvkwYfe+zISrE5U
MYWJR5lzWTwQyFyyMlOyhA1iKYrqNKsJcul0UEov4VQdyuS37EYM6w1wYMacOEdpy3CU44Uyx02z
B3zzNwfL9PN2P8q9gmaraRCENiHKU0bibGlmnHb8RSWR/4lt75pkkwAymCwB1jdkqZwag4tNLOce
lgnh9ikinbh8m3lI7MtVueTJYMgdiiPgj6xSNPWmLDuYEwcbU5YWLrP8lqn0Pm7oQM0yzGH7BePH
rjpDn4iuaDKlHd5gGKmbplZSQ9HaHEiT1obxKm7xH8ANtl+8G7beb+7CmyIHEAeONvwr2Nwpyal0
2IgfuL9BxqmdGSIi2pbraC6si+o4lxzDJkgrtypaoA7EEJwIIqr1n67bkBHfJSgK323J8YL43pw+
TlpZkYq1H1KuIECywHIvHfTC4vpjsFwT6evxMV/PH2GYAkkkNaYyVa7HoefCo4sVDD6WdoANFyaW
gCNUiFJCmwBmRV0yXBVpM3a8NmazmS8lpRRebCerwUQz6Yp47aDMaHdmtXYx5K9OK09eYgZT2ycl
zCAV+ymE6pZPBPgwfj4Jd8N55pcNOC+ZvvhEZKpFy2f6p+RwNnzSQawLLpl33cQR07lCiCbeyNv9
athR4JflD1Jq+qu6bbg/8gEcUw5syT9UgwdLN+JA6qJY4y0YNKd5XPdGWxR2pJby2yYREMFZ4KuF
RUU6UN7wnE9Po5V4H+YXWrd+J/hRUug5OiYFTqbQIyGX37mJ/suWr76vpaLIkT/fKLJl9daBUdDu
DR1qs8oYBK+IHTIa2CwTNqvA9SLwprfLt9E8DbCS/oB1PBAgukhDX837EprXSUCY8S/8c1/GutzW
UAIKkHoVP5AAUBzmXp+SvzBosy/YQLXSmbZkkqxnd782D5MBfR2kMB4KkUu7GAMwc46rhrAT0fgQ
8sQyZWJaRf3j85rFo4Wy6zMHE+IgcP5Th87Vpfw2/95/leAn1Y9tFBexAFN1fg6W1HaTETQPgvvP
pGFHVffxu6zK/spsZ5iRywiWYVLXAJ9WdfE0bsQZPXPQ8TpkIsCHB6fBpXyt2oaaxOT6XaE7Kmcj
6hQBNQpFNYbNpjWji1bAiMTVIAZ+pbBuJN6akcGOUp929HkW+0U9VfvDTIwjJw+1FXwVA5rZarQy
alky133q2pbFKjX3X0PqBWjRguv8svAaxfLgtd/CY4t5v3VtvxVxmVYYc39MYrCGUlmbgWo7bpVI
oHPxM5NeMl5x5rFxPX1B+JjboYGhOCsGYORZieWbp3q4q3aiIwg7QTuIAcgQjlBoy9R5EJ5QHWKw
ZHJDLZ0FL2kYOG1IjsyN2sEu/+dHsPm192SkZm4DKz0GC0E+Gy8IwHb4Jryd17l4yd/4F1HanJOy
N6Jv6pjP7v23D1LTPUEhlNfbtlpGrYCaPEpi6ai2pVVkgGbibxhI9CXzAYdcf5dVmgaedDJoNSVS
ktq7kdRk85h+lpMpyR9DpuwvkvzKm+BR1lYliEZUGQDiNnqA5vtkXMiFp7f1gg933IwaWV7ifn3a
pEA5VLdIjY9UC3oQS277lrvPzkvjsMmj/BXaYkNxZ+Relw0P3K9yP+qKvk7lwODbJTHIcC4XnFtc
M3fB5rnfX2qXOOyw2+RQ2oh2VBFUKKRk/3Ha+QOcxZgHG4+ZkxgPf2EDIvw0ICCrCE4eiRYNp1df
49xrkNPL0RouJbGPhYVX1j1ZAsCNgqnIS0AaG3Swbtmk+bjO2ImYNaVVXp5PlNhC3GfxpI6p8gi+
2RlTirTRTwImfsxL0qKl7SpdX0KcM6oNtcgmw58JrYMMfIehmSBgEaxg4H/AEFn/YzknGVMV3e/a
euvGobjornNPjmNVd3FCVOdqV6+hKySqaDUxUqn6zkcT7ehmAu7P8m5teqkgJDcWCOOgkZIx95Ok
Lsou21FKyNO5kFk6ybZgByZGsYYPQhXIHVfeah79BFj93wjaoanKqMSukacps9IBABBjPAqYTjOJ
sKD7dIv1qfsKdFfu/ypQru2mBHsrKxDBCX1zsboxrjIDA3TGt7xzwi0N33iQzQcoPqWMD3hT6K0Q
yrOXba+2w3ZFbXK4y65spBNS7QBo4NNzHUZtY83GXzN+byDKTYhyG722BRI5kGt0pmjAEUbqbXz2
8BO+CO190zuiInVKP/+vbLb5QV+xQWtJqlV5f20+wqOYKxXBzg4RLFOac1NB4UVzKUMtp1TyXOli
cQScKFSITVHJGnI+8UQAEJb3QkzPtzEHkB2Jinou/oXx+DzDq3dUTYjhFKX6O3HU+5z6cTyu1zwu
dEpSK9yq/5s5NoQt6XK+n2ssMOYYNtUoh6NrOeQhhAYwJ40MExT3Gku8hHMAOk4f4tuaabpXEz4m
srC9wVQf3lTKNWgP1/gJDildIlszlRlXT0bSKP+b/vIESD21BD2xZUduoOXQ7I7pAwaVDkn+ZEo4
4yvmq4II9Zv2y6khSyZFFA7JH69QoTMBo9ZjNyFfcLz35kvIkE1cX8CiBOJaGU0ACQ2msqVytQZo
5YSPYfXWXQl90pT1yic/4317KFkiKWwcgDZ2qeRMm3KiCckJT8aHf/gPrcjRm68BBg4AADb8lge1
SlI+jGGortikXAUYloUg7PvZ8ycen+vRJgEzro0HjboP0PVsWotOLgTFezOnVRTr6p6NwqUfvShe
S19oo5mAEKPaDHlVlBj0zH32BurrBNM+3KcbKm423Q//GotdJZCJf/RNjoOXoniniY1XkBr9+qe8
Sbptu5r2DRdk37/+qiR0E8GtkOOMFwvvzq5mQAC6+qSAXikZzRr/c+RKXlUSTIEBIrcPNcTuZL5b
ioyDuixdk6/HnuyUn74fEVQfCofrLL6FOe+6eYCSn/rbb0UfYAdLyLji5ZNSsoX9xPD9UcJn9w7K
Jk79W0Ec0+YKAS0ErgX4G5WBLckhFO0W7OflGdV/blnSH6UJMs/L0AlJmr3EE+OYphX1S+uzWQn5
eYO4zEhDqZmNp7Fg2xUHCh53i+xM3D3wdjTrmTyWJbzEiNp6JrNbI3mQmLvSIIcJ8Bxbgzx041XK
fpv6p32ML8JCZGyg5bTzb9YLyCHQGl2JZTy0ryOSEsi3sWS4vQyZ3JH8l0GFI1tzC1c7ddcbSh9i
qcmU/05ByINqDs3iUgAOarppEeayEk9VjYOQ4oE1O+Xled5B1YIBxaz4C23CBKCYQwC3j6yjt8DZ
dvyyAdq15cSOSTOoJUBwkS+pA4Ac5lznpy+wTCAFOALezsY8t+VXtroIciCXAAMr2SCunbU4bs31
xHiKGWcadvSw/P9vwv3tq73aHUG/ap9DC7mNYxCS49OXzqd5roWnfDYYNhdWmH5XS4wFXFSt5pr2
m9xdw7IScECrX30Pjrhe045Matznsy4tc6/788aSRKE9IDamAA5rfHvaok69Vmth+BUI3wtslGex
817ZIQa9P3JR1UZ+uOucJ6GQO4/gPkpW75kq+vPX/WVDwK6dk1mPPjWS8FNoBKu5KjfiNYZU9PSA
D7xDFeRMuyxnq7AaPGI7PDUvx5vdYEDFfRzJi76WsXOIdo+r2WjxB4W7s5GOHhrsnKTFti1iH/P0
0Y2WRNtHktMWc4ows06KvIWDOvFhnt1pbNoddVqckTkmkp5B1nMmBOrNfgjFse/7OOirctoyME2k
TFbUU5SyNC/Jj2nETDc0pHj6DYpYr3RmtqrGIuczLYnQtggDeJT1FTMe0lVp/cSTtTd5Fy954eGu
LJa4hrCCuTi57OQIMEKCe7QtUyyaaQ8cJWXlVGpAzl0GjyefdLEr8n8FC6YTfK1vFwqqXrJvZ9W+
h+yPTCi2VhiKEIU3Lb28EXj2jQ2zvy+XZGTxVL8GQ+rJhVM1Hln7JmHcIBkFMV4/Ab79drkZ97wY
h0h4HMGnipX7+VvM5L5oXI63oQWkue7TyEjBHepf+xomftoQOa+Qy/5wdCrupeZrjdc4AFKr8XeD
zGQt6LEgEI6U3qFMLXX8jxpPuGcH62YXngkRXLR15Q6HKIHg3sBSt99afI5qX7WLuqKR89EiCNEp
7L14JL9ijjk/d+ZRpg7/Ds6QKT394g2f8yWGBC2MjmcMSS/mgvSQWvCVQ0E3AxAwTPHbXONfju6i
Tzug48gdzn11bXEyWsQISnD5YG8uncjjDIPTdYn2hXk5mkOLmwwXLdGqa/sSVWb7mNSFw4r4j25e
PXzAYL+yVFBrltxbMlRcPK0XZFHGdAtsdLGkaIXOQYmrX2CEsRI1Oo7bG3K97RzznqpPkS5JY46X
tvWb3zjMa6dAlvqJsuhkIGwDnVocHZFjuJAuB8oJtkOyznV1NRS7ogKX5rcV4D7E56vdgSwdpk2f
WSVfus9Ial9Q1n0fLYDToXJMLf5RlyX6EuUo4hpy3UN06UcdHHEtVPzT4lai2zbpWUpg+G2/U6N/
xrFsnkoRs/pLWQ2T0LSERuO0p7njwzR/Y26uAzvdCIrWwmYJwK+YwGqJOP4dmrYl7sPA7W+4GUD4
k3h2QF/+tj/KSCRuFUCEmEPjOxiNUoJuAK6fYHKyDh7LSwWErRsA+uKmvLcO15+J33+08EDLVkFH
yJqYlNTzYgyN8UD2aeW/17A4Lem/26jeASsX2d90iyraZC7hrL1clSkliHl1w5Oc/3H7N65eWo3z
xloAryi7+3vDjZ/R5+HGFrxx419wmuWaoTxQkaQz8nLb2P+0oe4MlbBSuX8KX8wJjhD3Kbn9cVkD
TQztQKFqp8JswCKXrW6hRoh4I3LjqsPZZzgYmbvN2MnTxwQ7DShAwNGzFMy8R/iDkGT9jksdVYyq
L3/lWDLNS4aDugsrA2G3piECOYZTGTQln1LJ9/NVhp15fL2+4ucWUafKfuZqT4LFImuWultCpl2M
aYyg7sOHYCkzgdrp1OLX1/Yf7WWkDrvkIXDP5Nh3rplWaGuHFh/WukSqvTWqeenjped4O1Mi95S7
ii62UDOuiDLYp/8t/RxOdydbS3OZuij1F8fBoF6mAioTVtp3+BmwLxrmvVyZewiFT9LhPFRq1Nf0
PP2D22hzk8IPtZdKZh9qSpPBU8k/gxWhFs7cqEFRlwBlJS4I+l6JtQwfVlfHZoP8OX/1pmzfaw2o
0U2iKQsT5ejInS9Mjo70FMm5DvgA4CLnEbXRifDF+yAQGUOoieMPU8gAfRl/RouIrJIuJuFVsF1j
Zir1KPtNZANtn1g9FkPpgZdDpkpa6HWd7wUXx8FFbX10kEgcEcAdur8eqZSQmSleeUjAWTVp6Mus
kkIJMDcOPKl/Q9GJETo8eG5aOJ8/N81Zqat/r2xG/OUhMf6uuLvhQnr1503VLmHEDkOnZNuUprdV
6jNvDU1QsIbuxy4w6DdH8j4+Hk8PVPOjRgwNxiBAvvh4gb3rHkm02/F9PgTkIo4DKGl3yWfqirmC
1pnYV0RqHjJrhmNLZhRAT5izc7wswfjlfhaJMSnzAu8klbYQP5LY7slqgwTUAoBvNDvsLbVgOBcs
VVR48Fh4IKdvHCKlUd0bECQijynPFzgiFTglWw1SiWzcHldoAi/YIlXBOk7OB8rBM8Kx14RoM9yM
I66Ex5HfcLsw9ielEU/Muh4PzEe1c1nyuR+yTVu4u93gbAg5C7CirbNUXF6tPRnO0l18P4PAgI2g
wCnRoWhdFnfYzwH9FR6wkAURjmhhRZgbxV2DHrV7E9unnZzcK77CUOGmR2Jy+601++OCVZZMzYye
0ztJGK32nat0RJ4FDQlQVqFIJ5hf9CErgoFv5zoQkZcsfGKRcEijfOg4cH7LGSOH9j6BzVivx3fb
yStvqqLTI0jfurDasT/9XS8fTRnl3GKB9Ig1KxPfa9r+5wn6bK1rdD55SNaBqaasv+T/AA0XY2ld
8Wn4T3aVOf7aDIoYugof/hjG6oE/NyDxerzszB0PjIG2eJZ3kNmSNEB6G5Kc1m/XzeGq0uPKDimT
Z+HV8rAcTRfVZt/NAUn9UcwlnpkN7064m2P0BGns7YyCGLrCeACLqNvUcEMtGI+DMH4va0AlBrCf
EDkPtSfZXZyIPQwfg9+WDgoZEs3ZBFJhJnLutPE0kJDeBWb9CAkUUpyDLrT7WTyO8Lj7/P8MCfEK
kbHLf+c9uJ3UbF+to7MDOX1DDh6cyLxfZqr/PtBCHqb11c7fgonl+caNMVro7xB+SIaOmp+hsvMi
ZP6ItriD07tlr9QUlsCjNi3mS41wXfVTvPMIThtvlc3yA4WbQwGVIxGcked9T7bC8gvKpmzdieLJ
Jn/xuulrrBj0uyyMsHpM+ADRnv4dpL3WHOsDnpUbaOGpAcXWKNr69rbq5EzH31IJH3MxXRPSyHiL
YlojgIh5u8nMkwWGF9ApIZdCNhL1f0LHNdUAxICcK8qIEO49pPRqe83Vdng7aMLO+LevGzxDJ6J+
ilCRV4YXsOQTr7/hkqhp/lns6H1j3zG4/hpEz5wpWuJA7NXAhvGFb4GREWJBnNJ17TUhHjB7yqan
q5kJQYT+shPosw3jHol/nOWHYlegtrNes/eGqxF2uYVWIonQZcQCOx+pMm6++olrJlRSoGwGrOpY
XkRBvqjftX/MJaNoNy/xlD9GbPk3HQO5GILrbqoOOz1d4lQVmbFug/3424SuIT9eypbdMFbwJN5W
LmLPoYXguETCTknatrunbEYtdXhKIP/qdZ8/25mJWsfW76+w3e4Hawn9E5JdK71k9AkZN0AmN0UP
EnIFnHNHAnIsOxkEDOMU31CTpC7UBCpOBzkvvBr8Spa8/lz2hHlINHAG1fbyktaI1vh7k0g7XQkT
g64LTw/qfTV5HsCzfTCLtuadRlQcHJz9YOD/4UnY3rf8fUf07QyGiSf4QAgTNdiQ8bbUBmlYHTtl
CZj2wIgtfLySqkirKmp/CpSL1tF1tmQuGnQ62nvXFHuHJGyiaIIRJfrF7h4yuxP7LPHv4nATf7RX
XyI2hvY0Pf8dMnWDZ+RgzQCisLRMv1seDekRVoMUP7aMAVUKmrTLUV/C7rvB4b0hvpU/KKz5bvup
rXIYI3A33I+gwUWCnoHkvv1fWHIZ13pi4RIpF/r/S5ht9jLTBWgeuhMMsMfOoBNIzccAj5icKleb
+BOOGR+wP/0zCPUxGSAvSeP7Y7u/RRzZFztJX4geA21zIIMtfPTucOgmHMQKPTFuDE/I3edl3U4O
kW36/eppJsf1KLc+wWMAeYuC5zbXLY45kgdQK13mho4uCJ8zm8iIy15vYKRkH3u/V05c/XdWJ+ro
1+2XDWsSSmK9Mp0SVDQhgKSAB3ugsau7GL7boFX4ytRsvwm+EcMIgMkE+ZeWyVCbWT31iPTBmFIV
Re7StDm58J3zdxuUhGeuaJt4dEsjuXjrYjQZBdsLcBlAlc8MkVOxP55ftqBc58tNFIvpAX9OG6mh
0fEbDtyACyNa7RxYE7AZF4OT/71qvT2EgIrQk2fbcQ4045+vj+eg5vq/9Nbbyzv8CWKjHyQBTAJ5
PRGFXEwxuJOfzgchvI/dKk4M9Bkv+ASGaPWuRHUBigVODKkRTQwJWNreiqEVDjSyqv71v7GPds5a
aoMVh0E8kkaG4AaMvjZGjdxSvDyUXY1ReE2CxUd1tpwb7HIfKEYre7LaHrdC2fNz6QvDLphUq8qM
09qSOE8blDKwpTot7n56wu/WdYOwilGq27qffaabtDw4IOvC9fsbEAnltx3chUR+zvtZiXCMiXDl
gURNO042wv7CTicqixRattGBaLaCLVZDKWSY/45nXGZ4ycgv3FfP2cyzuEBoB0f6yRY/u+POImC9
+nofJOuEh+0vcbHBSY9yQ1fDmqguy7za2Snb96K8yfg3jiBLvvi5DiB4WL99MGYUXtJpe4h/O5Bx
SL58FCetUZd8IBd/a9kphIwMXf5/Dfo5FFa7psjLA0oAzUlqtkRbTalCeuyejijdQ5oC2QrvVZs9
0geKPfj+TQhJGc69Ym8JMZCGwkoQtm4oaxGHEGl7bY8bW5P7FGQlFBDXBG+B3y2JnPZa/LMZxHX8
9VeH/uVZTIg2vRmULxYDAJk5c3mmrPyM69Yto0HskgTij96zEup72eX35VhITaAyq39S68mEFt6i
V0Lb5BNMfYfscVtSvnrPm71QWmppw1C34ZETCuqF7DA3U5IHffGvpP5eZd84/62VAKd+USw+QbKw
4idyGsophw+/zvN7wjDCGfIK5PzjRWeCgtNL2Hnqg68EdcbVIDmsRH66K27IojY6KYjft/sIEnbv
uBBk7F7iTDu/NOgtq+rspEkqmRtl95HkrjQPgRt6UDwj/rXuZ2l1SqT0SWfR5F/tp0rrR5eKDfNs
M9Vh9oNJDOcPMs+UbZTI0j/chpMFG3nCa+6bIaeLiKSjZakDaFi7cVpznDtwcbT8X7GNUGW/THqb
OHDQ4k6szy7woiGhUVev/oVX8VhDTrBXfmOq9gQjqMDdJJ8PS8fZGNiImKDyND98G/sKGkMJnwEz
yy7prCSsR/qwOHeZINlT4qVCNKigIdL20t45ya3adYDNffM+7YWalTAPrgi4PkWfJq+O+Y9xFt1k
ff7fZNGrD2LdnVPkhvcg/Wwb0P+HxxjsNCMFGTR7tqPROplnWb0ueVd3kEuhVng+98yWtJF06yTR
z6cNEpxkQCQ04iLi9Pb1X4OYh54kZvIkp9zVlFQvYzZgW0b9w4bX1PDTLtef+f6fBkfB9nzl75vy
4hrARzbYU+g+4HmO9M1ZjUpPO1PJvbVdT3Je5v2I01rOB2qhIK2ape74yujn70Jf/7rLjBKfqNDU
ZgUN/KlDKOe8YFxHJ6gnuueWAjzNJW4giPdT35dwN2FiGAnGTV9JhxEm43wU9exbH0NMu1HmQEZN
ewAsnofwFdEzWbvh+K/ofv1BwbJ5mAHc3PwYCmdww9WhFtKK6bAOKg5LX7Qp3AjSibF5z7Y9I2g8
WxhpRKspDfat+Up3NxSu6XjDb2NFRTbL1R6oLkMU9AdZvWCQD5JddruFVCyv1pwQrDwbj8Slqhdo
IIHdBgEwlrc/C7joo+z6A3UFk+FAzT1Sdjx/jpMEtxrJJa5YajiZkW4+pUDVxHn2nwS++p9sy6nW
g0CmzLDg+pG/nphwL1GiWziC3muJEXsymajqAiDRwlqfMuaKXdWLk48POZPbX40yZ+xBDHkFduoM
RTyOtM2MA5giFtl24AcXHVBvvDf9xMtohz6Gd2nuZO5f290tqT5oOPo8sQ/0jKwYCVKAKkfT+dq2
Se7MXdWHr506SAZHg+KFSa1kYhDt6F7laLEP+xDZs+7keJ976Nophaqrj5KR3dTCKZNzkjpKQUCO
HH9kDJpNeTwEfGrFwkkHKSjN/dG8Kk8n+sz2MSLpyOuew5JSI1bKIuEWFQKXkba6IWLe6eo6diua
QPErmT++gICv6O5pjOOJnbuD3tM0wi95ld2KQnDyZfRFhHjjURT9QKPfVKtnR+SovvVv7HyvQaTK
TxuUYFppTbRgztQiDrQYbcaNCThMo+CQcykxnSDRgpVcPeHN9l7hVq+VSWgQSsyQf+yhxNev4WI3
CA8Ne/C8q5xfUSXpf1gS6++OlmxB4J7KYC2oMpMbqHit6ndzZeCY+M27sEJWCufayL+V7EXFI0W9
uEQEzgdfJia4VU9bQ2T+aLHKJGsANfZRVTzHA9rCsQ9On913kE8pBYRnaccVPzGGLkVO8N6ABXgS
zz+yZm97u/mAVqe9d6ZtcxfeVT0Wz8I6/m7bWEqVtpRnMXU0NEzO7PjrV49CbH8ZVt0AIc3jJ9je
SYZUi62tUi/j5RO2FNvqgeRToNB55NgLQT7NWZ79FAmv0pZMlGPMzNWwSgdsrjbRcLNtk0hAzBdK
qLOAot+zrDDjP1QJGvRIHaDIypDgKtdu2gKVnkEKaLiXspHSjOW3mKke5dmgTlsDVkbjtk0Y7+YO
ciHjyU8QdEVckOde/m51lah6xs4aNDKKY8WZJGdhRkjjNnRO7TyLwB8hpLq/qL1PSEgvgPvZBnsk
EijehtvqWd+Ej8iB7bLqUKzCRd9MZLl8VYW3T/ebNAhgDU3P4RYH9y5HacK0wE0DvHvDlLOZQRaA
mtVhgYbICmtyJNsvX4uUoE4IoAWVqZWmAviIhSg+AT48TS5tfDzVevBWK2DYySMkqeTLjvlUPPiF
sovQfNmNSFGkZSn6iyhBpPFybCi/ls77+OyurKerWVhU20FXoCWFW4vuUFbvJpgDKZphPXHhSDso
8cDZEIYtyF9DRbLpH9ikXqn2/NzpSoFzvxVwuXUVaoh4mnT2boL511I2QnnuTfgpUviQjRHmdXoi
KApFPjfBDE2sCJP4CQdpMA4sv+vfjYLSjLIHythVTO5BvsYRg2hhWMGwl3XIkZnw6eUpUbhseOHj
N57cyznun+mTBHFijYOZ7fEz1YuVhzS0yM2aAieG28pvPOa/HN1TyhtgOx6BpFS7YO6oDzqXpJ3P
CjRDNBV1PnNgcdX3VO4m+MusSI/fi3Keh9ApBtxTqjTzRERPChgzOPgVEPUFoxopzogUB4cDAR4q
FCnvpZKSVYsnjNOj72hj8Zhh1n0WlomRGqFx4JJdGG+s52QFDygABQUHg8Z+6eb38/Abr8k/ODMV
RExs4I4soAHkvJ/ez+hCSQ6Nv063nij37V09kaMcIhlGZAKz2SOgE8PU8hQWtArFq9mn0KxF/UlZ
XsXZvIZ8tUfn3G1U3RSBejN7gdyJa71XBMWSkKH0kKf/WUB/7wh1c+aNYw4cJRrnrDva+rxPNS9P
gdfJReVqawUGfur6zMQ3YuXxoi0alP9rA+elbJ8dGTFsazhKXRt5U2D4bjWw+LrXLdLj4Ef9JHe8
7EmZt+Lh6VySkKSEXWm2b3/QQqB7qqpx7Log2OX2zyumXNNsIc4NLt4t66Gjd/IcwjiyJI2KCpAv
aiXf2yK5puiAAByPoM5eQpb+j9ecaW0zzkSVpsMOErskj+fIq5PWhPj4SLI+4Kj+CYv5xrBve/QK
T7N3QFINE16P6LXbFvBpomm/K4ZSgoMW5LS0yL9HsSLI/6QYYP+5Gaz4J+6HUP01uk++28vVeuNK
LlzWH+LZX2QBI1uuDuH4dPIBYOEU7SVoWv8BFVqsojEGOZiuFgr52fArU4+0DuL3gzl6m4ubWdZl
BhYXB9DstcjOwxn0fbV6shtTvgQWrMlx7g5igAiM24HwUE6cUzg+Aj3hyCOVNHxAT3Yuh6bCEyM7
WKvlN0/CmP9FHLnYkC7lCJAukjj9uMN09m3xht2GhXHHepoWvAFXCxo1PrNzDKB2PA0wCN4vaSoU
r7dxKPH8yh6xAYfwNeXHSsfymhSY1R7RrBbHoE/ZJ2gpgrnEIuQe1Of1c67M592mn4uVjTCXVIbL
BEFMWdjWQ6wT6330V1PA+cXSyEKTcnaC2dTJUKBWP9qTr/Yy2Sg2AaruO47lTpoYw4K7P4107HNx
hrzJ4kDbaWZzTZ8+CG3aIKEVAW3KsZ7NSBavEIbYLpxwgUSjcwHTnkNUmPpoVTA8VRbmT3jy3Ttl
Zb86ItMe0a1HylgobhF/N2fgsT6S2iMFK6w5CrwV28cMKz7iwcbT/csX9RKlBx6/8xeibABsI+RF
CseA2wrwuruwk8yR18WRRYvGb8xuoTTgP5oxnMPG0mxiIhf2Pedwditav66GRl4AtgXyz27l/auN
PFU3KEwYak91hruTWiWCqJLxzH5Z44qEOE8aCvQnuualuxXZpqkT0Uuuh4S4p8lAjQNuwepnSvmT
nZc1IOsDbjGituxYKRA0LX13QdkQuU6g831myyng+nBqhnmYiJCjQvEgfuTt/DlbWr2/KNsF4Wcg
wTMywqzIjaD+RU0cBJN+we3CV7UER/5KfqIfy2Zo3bUFG3x3pbk2JdwGhH5MtimisTZh2w8m+2mO
ofb8hw53679BEQhHX2SnudkFaG5mz+qBm/8sZrjN/JFBXyqg6yr7LhjdnQT/vfdtNrIcO3V9dJ9z
JRE2zzZnZN4vs76q1y+d5KdPD7mzbt1Eb1uBGwW/kXrdtCnN/d2BgVdZr+lGqMqNwc+my3Pr6ph7
c194Ad4/HFrTPl+0eJvAhuigMTeaD9kf7bYV/vy0JSdsT6529bcWDv9w+Md0X3QcDyKP1G3hsNgG
vADDyDJKg/p7wQ0m8t1DIjwsuvKSS9zo1/BRlKhRrs4sNyqXXLmfK9grKXhi/qMJ9OuYm7I5DA8g
Qepuyiz+Omk2kb+BI89x9EDbW180mid4YjvfKbCLpY64aWBigsZyPA7l5akbckoqtt2vUuAP+10i
VlUE3CohNiCk/nZuipBG9bJrM473AVu0FucBJwr4LQNv002253ei0SZ9Tal5KngXV9QRGKU11+FQ
bS0QLQGSRLcnLOqiYdI/lnsP050xHKaRDLYFM0I+vCpfk4tpfTRPPKRPen1GP56iUdWMKGOCBTZa
MkEEyrnvaMZWccPq94ftcOzFfqBXTI7htJ5C76QIZQykfLugANX1NxxfrZBp5/0cmHxTHUcdvkOB
i9cPIV7YWuYbybTJURxtpYk4FjwfxXBBdmyTThsnx1+z3HFTsrLc1E3QhTBjtoMxMFJMPMQGIVk2
iuryUY61zM4QqOC5K27AA4aAYmSSgNkff1Dh/y6ZyOGJvQsWsdkVlRHPI2zA5P78UvfuL+i/+x5R
hgkvp3c9d4ugErpLLX7REvd/Vx1a1FTwtik7jfU65EMQhNpKFmqWCgnIRgTYpTSU1BR6SGEeRe6v
hKsUJgWmJAfwqGM8mEBchyfQRSddqwc8OhUgQKx7ruqud232yqDc3YHMBeRvUmRlixajwhMSKCC9
/ZNC+3IQcaAeGOLEFMC3JA6L4AeJTzo1Wc2e6mkcKFVBDdgSrQNcFZhKwB8v6nGnD15Zgc6sCUbU
uF8igrVUx6hsbUw9rdvu5eT0AZAwNKwlTSQUx8VCgcsM8/lZsgzB5Bin8klsdyqhzZa9Vv0bsnCf
y/Nr8XksWBDw9i0h3MDllDR8qNtSLOrc2IU0Wr71/Io/SJMYGPTVP45q+GwbMwfKfQ7ELEi9UvWq
zS1xCGj958uoqBVJhGCoh74Fs6vDbmd/YA/6+lBOMdlwUn/2wEVKbfmyK6aQ1uA+cljK3F/CX1/j
8hoJCZMZERb+zyXQaesrD6eSQgY+qtf/EsRBoxYqdqLtS14hj2KcgzOjy/WpanfmZl+HiKNcIEaS
gnbk/5en41iGmCw0ANOLW8GD6EalMBEwJUEvtIBrZquQo/Kf9JFNOU7kVc8vfi59bjBJiHLib/EA
DNALGd9y/u3kbo5X8T2YHF4pSuclTfosjbQDx3ke2KV/lpABYehqxEmEnJa6ZgzSkN0hvaHJv+Zg
cpcqwt21Decu0q/wnDH6FJ60TziY4QeWZmkVZaPkNfNx88jUEh/wYQwn4XMZPUurDUebyFfPhNuG
j/rWj8QJ3RQ+0oMrW53Nn8B3++/M0L5kNkRoza0FPSFC2jAqh6cReudbhI63b567U8rFOPNRhka5
8Pfuliw/BjZVNR93QJbNMnrm6GMarXFPenlv4X0S25lTcVGMJG/jsZrlyl9IQBYj5L0CjdykAG8k
dLhFd5EM3UxIGpPBZZtJIRg1b8nUIMoJ0gUO+Nxr5G59yq7PzF9r5jUBrRehU4UIvYg9qvCX1Bgc
9UOLKXJ23l5kkZtPvb7QUfQ+TusOIFvDsSoiCeAu1PH1fmHa5V2XCSaYDr1qqQOBFxqZugDDknF7
LF/fqEwjuZHpwy10qvwHYQDdArfV6Mek7G1xDDVSdzmrBRw1llg3p52zVPfbwR041wl4meTV+zZb
FHP71ZfnF2DvvX9EZyd3tgD7pABP8AWYlbjmXACSZwb8ZrG5ozrSfoFEjiPl9JfI1hyI9JEy41CZ
qjeIZnS3O8nRdvOTVMntLDiKqWSIoyaknzyWdCR3JfS1n+bHEF1O2Nppt7BuQJas8fwfXCZwbNlh
4vDuScLOxZJhlUyiELplzdVV2RZbUCh/1L5W6TQkEJYci0KaMpFnMRPSfNprl4jqJmUXuJSEn5uT
lBpuy14KqbwxPeQoJA8kTWAIjEyyIDdhBrfzXmpRXlaDg/cjjBVTTUbv7kWudXhITr22TOz42x4b
WUhS6Lk6Ch0s2rHuKc8/Q4ZRtR14Y3NPeUwYdvMK01Qrwir1pg289ZFlMs6NrfK07BgqYSL/kLcY
ngKpP9tDtnqy3ymnKr8Lf39T3xSk9wZW1Nv4R9CTLb5NwDu2kmKF4iH3eJOk+iNmg4jIx6ZFdAOD
ajROc4tjBQ4h1MQuIEJevTxGsmfiiVLUqZZQonZcIm6PnAIjR7Jhe2yZknykR3QZLHOEhn8yD6fL
y6fbLrSH1EzW00nk0sbzm+q5r1UzqfkicaAJPyUJZ2UhyhFoKsiXoXBwKvddF8HTy/RA6M6zxthG
GStoXG7YL2RJlXCFMtHTrvT75JZKRaKJsGeTpMsCIlVs/wv8NPsNDfhVj/EjGFAcmQOr4Pc24Hvo
EYrSaqsy8HAVNnaAIe+RxyzRZ9Ctt7ZbyPtwqwecsiz1imXM5A4B8VntfIw28pWUZFdc8cvW1H4u
jzzvATm7Lc6RjQLMlhY+irre1IwsI2KSdXB6bZQxfAHQCXW/aDRmnYrhrtmlPBEpadj5O+rdrg5S
rBhn9ZUiuMIsjx9iQ+QiYSOrzX3fbRJln+s8dI2xb3Yfo7c4pc+1spEA/bSjm2zfDTOsvmfrJKGy
4jljHBDbQoVJLb6zo691RuyCIv9oyKMVGqrKKiSCkkqsl23pbDpmuSfEbW05m+ja04n3TRZ7I+Aa
W5mLi4wNbMNtJwmWFFQSapymMnFUDIcmNcI0K5d3N28DcXMAMCNRF8FXHNk+8kOsWm95k97n4Z5R
8YLCe4nGhJ2j4J7pBHAw496gefv0qsT8ySLxmcT+a51XkPPifejOrwdyAoIHpE6cdeYmnnL/1rGw
8/QX056iFuBZXH2KEC63EO11eLXRmzeqG7m0YptD8+2yX/NhWiQk/nOoR2rN+FfYRKitiEjhIhOi
l3CT5xWw9aIk2E5jtKPTDWISX+UuGoi47wWGxsfkvVvsQa5iWUq8wFvyd+j8fBa9ZUToLabof2Vh
+5zkhftGNGdPZYTXJ6Ou+psh9jrz3V4yv9omgcDGeKgW1roLqQVQ8TanSV17aS3TyIxzZXZ8y7dm
tXEbAJYYtaf9uIlbOT9qoYH6PcZoCJ6HBv9erU6bfR+6skhAl6va8yjTvyof5wEzSbYyAFag06sG
f+e9OcgjleanL80wnDqZ3iB87HxZYETPnE82NzsLI/xu+vfclbEHy0lYGMGFSzK6JiG+COh+z3d7
OkintlvVUGc0RyoHrl3v31JKc3kWpPMxE7jEoJWxBYKhOloEgXehO0Mdmu+oTHvhUERdawgQ/j94
gK9D7WbAouF7LbZetqs/aa9cym1ZbN2fA68sJ5u48d/248y5dj23sH8aC4Rco1Ig5I0PosFcCrHw
WDKcDXo9xUV3w0yWetEFxxqvENg8hJJu4Xs8Rt/Qaev5SMra7AdsVcoUKozowKS4kdKUZxgebMWN
ieEDuyejJmOaRtUdEy81BGvpI4spafT6+4tnVe5TZ/45L+XDe1p98XR3EVYWScCal/kSCXAiyhRz
N9WB4Sxvf28gKQyuuLuW8AvbEyelHzu7t4lBwQEwD9Ydq4GmozHRYgA51qhlW6RqN53XCNZc8Pya
sFl0csQUS95zXPJCCO0ByRRVUyqQAESBFVyj7E/LN1IXbxMxgej59pEcFWwYYE/iXzwxPgJ5VRRo
zn3ojAYUlaQF4hVJmczxNCvCE8G9ePXWSluYKEqViKvZfYCkcG3J7VyX3UFNQgCLCvghB+agKP1D
6aWTpN86Wc9jXNtIi5AbERYP4EwDS4OVDPqSzwFnL/OTUG+s2ifhVFrrKd3hE7/KyZgG2boLNGQG
LXtmzaL1qcrREJtDXdptKENi/dEFZdNBTNgzQEBuebVY+DezEAQEuV1tvNNJ9WGo7olYQmviIEU6
gj7TLkncYsB68FEwKkc/ImnJHhFD/tURVUjvSpdIVv6wMyjyddKfANEYPLvNqbAeZ4tBzOjns9BK
hffxrMAPxFwiW9BqVPm8qLauZLhownz4ehDuU3A3H849DMn3S7AaJGPIOQd07qyoIR0YivOyv7hv
HqXG/gxfIuUbz0MeskPvWYc34uh9DdbBpqt7AvRi4ZrMujUqxyvpHoZdzn7EThevx/rJMlf2RPYE
1GjJGznQzcYyX+AuRVKzVDeMqqjGUAWWDrV6iNjCvuz7Dl2DeOpnkXP2wS0wCQdetihXAJodYjJ4
dj7+j/RQ6sfxY+5ibqd0ScqAc/T3f3YYnZ68TpXbWOc1il2MxwkwzsuDGgjIURJBVeQTmVPVI8Ha
k27HnnqNZtmtI8pW7uLZ4TY4jQ38zX0JfRnQsQNUxaSLadNqJ/1RV3aiN7ccwRorEHTefcQFiXGk
0qrQQl1sXcB1zLdv/S0hoSXfSFiISv7aimHWlySqtbbg6FfSavNkDHFJiJKB2yMVClKfQGgHZ0/J
j6N0FM65w1QVi6G9uMyK71HqzEQUXNwo6xbv2Mk7mr/nGHEPhU13pkRTEgnsndCAc/eiCcZdM80z
R2sQZ36cqaF1EnL5lOtCJB49KG7idUohGtnOqOjF0YhEA9FBMDzrwkuu8DAiK94kKkPhjDmz4Uym
e4crTC7OwaFRBkmreKlQxID7R3eVZPLpl8a1VWbBR8evkviDmw4HCkbCKPPk5kEsoN+Q4El+ix4y
ItDPKUio4jkodEPcd67YjSGW1Mdiyyu+5Q024dnBpE1iIkFokSz1O4W3OKX6AZ45PVWKUrIQLEh5
WShThtPqm5WW2NaOFj5ATap/HbgBP1mXJ4xO8dsCrNmH6RI2DRm/76htsrevWuMa0YZed8AaVTk8
a2nAn8mGmd6OVLd4g/ImrSNFzeHjQ2TWfARkdclgejc6lYaAFJRxR5T1aKNmAqEXEUGEAYnAQE6a
60oEZzqFa3GZ5kPXiukIoI2IupOf08M6g4MzggV2quU9A3aefmrvxlUZV1F7RuolwfupVz1XlSJ8
9bpJM6IRfTgAqHfRLOzbXlnIySkVgnTRo4Rt35PH6nJtPBCBjQc7xH/l6lErM8JXiuEoU/LkL5QB
2N41aziJ+MF9dRI+Kx5hx9b3l1AQ0Ukwu3TBj2asnvwmTvCL8EQ4MX1qPVPlib/JUYC73W61Lr4V
YYDfiBc+9ZUQKIz9fpHGZaV6RlDtyKbROHy6x0y3xHCGS3c9So9OUuGkv8gtaCFwdke7riCEg2Ee
ARAlkLS07jO+6dnTsndwsI6VBjp8DEstGjcOxFNBgLyyoTo/ycU0J3Q9H6Bg8pzOdx/zq+jPxRgd
g8NVGkf+BJTL8PnSQws36EtjE+nHF0svOo6mfCVB2Y0DrLCIW5jw78gxhz8WPbNJ9clQfcJEQc4u
O7QXf65JvRmwD+fqPdNeFpC1/EBgPzrbO3BHmnU61JnWv/gyoSmi5FO0Vi381S4L8AITZzBvfolW
7V8eNIH0yODYrgKMXH7QWzUfiCptQjUFqLm/6nmBfIFk9IzBOqOWKBWxzhf3K2suIgWk2BofeyI8
fJ9PwjCBltdSNoAg0w8n+sN/LRwSFIP8c8lreoewKVMA5w6Egojl/aHK5fEA9am/QdCEb2ymF98W
RBtdgDuwI3beOQvBorfn/VUZElpUEgFoLtqn98paZWaCrRoKKsPpiB8K/Ip9aG64jP3IN3oY4F+J
E8KnoQ3+mC5FMsHINa+FxPgrj5FglchBz9Ub/R9hJFP3HcUh83MQO45ZgtHkElpwgPpeUMh04n4k
fcQk5Y7quLLafDbBRr5WIO68zpTIXRCHRtcGfj334bvbBut6AIaQMC0enhxy2+6IW9tNBd7/jqGg
YszA6pqIAxEfXEBDo4Dc9onTwOHxIx3aTFOioKU4p0ovX3VcU9mGDW7rl7I+yojjxCVd0h7lKL+6
xC8g1Lsii3vMkBOzwZTTyi0S1Or1FPkdKRuzPyI60xeN5bM/aypOimMS4ALAFZHCio+14czGs+vY
1NCgpBZrUwKMj5Zy/BmzObbLych7Z86a19afefoqqsY9Oca0IfegP9vAwOZkeIafqyWgFcSS8SST
wBOd8WyKnynjNx3aNmD7kIgdyxYzdjukMpG+lBjZBaI2GPE9nmDedjPgvUyBcjHOYEf+qyY/M43l
kRa/XFlxi0h/emPECcslmKnIFDOZEfMTLzxdSL/+b/Cod7HhvqOjIc9af/lDbLahi0QJzPUSWsDO
K5UttGbeh/A5Icv3GOZJuhwremo8SVbzfNELhCmM1Qhc2cpEIOCFsxEMjxR2K4yud1xIVg2LCtWB
oht1Kct5nH+JeLGqvYSEhdn+11+OR6i1Gna7yAhpKKFPeWG/3xmeReCNJZP/axMree01vtcKzhvh
WfGzu3MZ0mTv+IgRt0z3By0mRPDdLZOlsw8tnZ2HpYcA+z9fH1Wk1pjKDAmlPbr/A0eStX0AYoxI
KkTInGQVf6e+K69kwfI/J7GBFKsiEMFWTLaSJg2jcqxIo60jo0kRPJI1MzWJL3NvLkBzdc6gFmht
fE4pIC2nrmmZ5Bc/N4pmOK0kLo9vvtrt7JQQRQ5EhW2a2HcMHjU3zKWGKZ/1Gq9Xri58PD7+F17A
ZhbqSHaEy2PABlgYdekCYffyegamg+TvCDhBDWxh5dFuFRDacHLXThLMt41Fz5bJ2mIYR3j2aPx0
tiwZecSc3CZd03PfHRYbuBuOd5zyDSt5O7XWE7I24q+dcAKGGXvkryXyY3jp3zpx/r9ircYcysaw
0ewVw80pEJxKLn03pHgHHKCX0HiJ/AWY9Ef3I0j7Gbumk9q/VgtphO0gQvbyJeco1RANOcP2aiiv
bLcpQXBGXaZofFy4n91fA2AnEMVsg7K7DHQF9lDOtGy84P4JTecvPsS/CfOLbv7c5p/xFc0/IQgx
NUZFcFh64/B2cCsWFLz8OqpgBm1EBowssgX3UT/AXca1swKeEwqh96mDhOD8IlCXf0uZRWGHXn9c
fAjVglJn5UkoHCUOHdUDWq9CNXEoW664Twa1rMg7+6yfSUtvpn3vMaNiXhgEEb8oYZDR5pnZmYFs
2uTwMchwOtfOIt90pS13btZ9yY7Nm08zncxTRk0jpN1ttre5TCWKUeDcFAPtD0FpoE1PN+IHtpr5
5jl/NMhcfajfjqKhs0qZSNrxgcXx6Pd5eTaB1RGwcnpIEKeSbpYl/LgI+ChgzV/u17n7ZHO/mQcE
6lgzotpiG+if8oCPfDANG629OYyuiEAGCieOTWpyIb4+wUnLvSHzOx9IptDfCIK+DAKeJ3E0PY8b
sMn0m20GJyMrBeUcDehUchQL80gXWUYebBA9SJDZUxx+e2/kOeBaot6Zt2uuwcccMInrbB8LXVTj
gZQ7Hv2ZSoM0VQzWb0NefeQ8FhIYZr14Ycrj5dY5I3rSHWBBPFGfTkzEg2adr5So0CsT5KoX440m
y0sIjP8XhRx9p0uIVmGJViRzpo6sVY5VTSbKhX9ZLm1DrK+ZwWf8tLhNkp1Rp4FiLBQCT119/OXA
Hoj80XM1y6zhSuApHlDnayyWQjYnx0/0GxXOcZsKsgViVlnUTD/oOwsbvvEXSK71g8/ioQ59YsBo
q0GEzk0vmikqnjenhmAhSlWT3R+QJRBSFrX5h+PnTGbYY1/3Q7ZyVPNdLOVo00EY2wrUH6hnNwHN
YeLYHRA8JO5m91KGqmThNcUJFWfegvlCC97y+6TZ9ON4b9IbDHCwgKRB3dD5vsmtX4CZYAtWfFBw
PJtmWiKqc1Mps4vT9lg8ICyFh6CAYeMZcsGkzECEbBJbmcqCv/kwqJ6D9jQP6+HxroQLQkqVjNG1
+cP1N6HrQbtF/CUgiCNMll0DdiRSPYS1vTK60L2FNwJDWuv6AoHC9JZ7pkuGphsKCShAvQhu8XoV
d44vH/hsfY2gsPMolqTamLpD9y2w+9HPQQUp6uJhSdAik3LPq6sihrzNfHLHEEyqDGipgqsV7Lqx
BlZ7I86922HfY83KqyveGj0lZq1Tcjowd7Y4WigdhrthYmpZpKOgTpozobOAsASkPFUNph7jfP6+
c2TlepqWQnh3L8UU+TNV6DRF+qiF9ExN3qyc3anYHJAAiY8opNxIIIDZe28l6AAPPPBxwmu358xU
R4HmrDiKE19hZgHyRtoIKAfzAfLM/qI5GV8xdoeUaIAo3ns1g6iMCrqBNyGTWdfIPT0C0kyDBkTY
fo5Bivfb0cgL4f9Uopd5KVy55/7svm+YX4Md+QPNrfp9iD7usDr0RxnDV4+/teLMek/S4ENZh1i7
UvLNbk34Gyjjfqk8i6m51ZmttNcMFZEQRokafCyANknTB7Sl782BjvBgU0Qk/4IDcsihlU1F7Rik
CjcpIdd/eGwsn5fmdRQ5AmkeQ8ZA/s/Lf4PwqqUE6e03XaXJbcmMT6TK/gtI3Q4C6Lrxp0NNira2
dRc1RJ1ZoLRf6+EIKsoAhd9aSIMVgiIxmKVilCG237lH2bJUEhiqFN5v5YNAwX/pcU7jESW29vjM
GdQPycT8elVMlOFIxPpNzvmNxf1irUpOPB5u+PPI8VWWaghkhlpB4woQVcJ6yfT1ZCuTAhM6eIA4
sUHZzXRxHSlqZz8tYFPAwiH+lE/gtl+sCNO328uwvkKdPOUMxw+PoF0Z6Xa4iXx1rsI5gpTlrz+5
LM9/VeV3zxpvlZDQMcaYigK/6kX8DanI+KYOkC4n8+GSHmtn3ZPh/X34MU009XeR416iGGvOc37S
EVTC9elcfNGKPTAum9/BcCB2qS1n18eoPcXEbP8xU3FEPk4boJ34f8WZqutljJeYmaBzCAlPYtig
774nnu5WYDZgSKeuLysl7MAfMDpnnFNjpJQHoB3FCAdiInyw88KHmFKKt5eIPlrFxrn97eqqAgpm
edziuLntfGX80YlaFuUQOx+1kjYJGy2UEnPf90jFpsscNhpCiZ0J7rHKH/ZvcuGvWAdIaO8CZ25y
e2ZHj1DYp/tcAokVFMgrFWrSWmKky0fVV6EExzPV9qmD5Fuk5eOU5t7TpGNwBg1V/+sICjbVl/ga
a3W8LgF6+UCVlb1YY8DaOqArdxUgmJ4LovCcZ/Z31IiiP019C1L3+w92NvV+agPZBXGszJTTWOz3
J8Z0XBHdkgAPsYEvlGr1RsF/WxI0/5Ut66Y9CTrqkrSIyY8qO5C29IhJ+fy1ejNNZJdjzgvwfv16
LrBo74rSJbuJbicanCAuqXOmtIFFkTOJlxFYuu68y5rszO+f5SK+u5jGt36vD7+0ciKCS38MCC9q
i4Uu0R3xCgJ6sQxTSk2Bh/XroWwv0yAUfHGEy49Cw33NNsyY4nr0guMGf+bKHV+dtwfJgSbeanOt
ASbIXqaS1W0KZ8bhcG9jgffugS79OiuWCyEi5ciMix48dc10xp/p6oT5n3/fRznr8ZlLmzBy5VaB
V10q9xTfBRaRyOV5upr40g4WhAYXFLdH5bMiZdpFavwX+wl/Xd699kMQTzYWa7J44o9Z1Q5sY01u
OX0hlVYUKMB5bGKIsX/3skI2qtAC0dSEKGlFbaaJ2ZQw8ogY205hlqs7o9TLPdYG5lJs5KggIMDs
25nntj9KlfWtce6709ifMJvAFEyeSbdZ0C2FyB1Fw2Vyy2cIntlJ6URUdiDbrN+9b1OSQpwxlnJv
TtyOiKjs9VO05cSqg9s31gzn5p4Kta7TnZY2by+LKk6y3UHMpHtStrMGl/KkSODKP+ciYAgK5Wv7
PPm7gDgxg4O0XtxsGsFZzMd/5ix61suwRa4CqVITTCHfvgBHcQNnkHkeFX7r3IqzClBaK1NnVif7
4Hzyx0RybFV7yuSbH9juFVEkc8NixyqjJMXbGQta8jxfwiltXq5ne5t7g8wWlGGU9zdX02j5YnIT
DMbXlkZ9w7m7QYuK9CVLntr3fMB8Qh93tVQUAX4nCPirE04LeeEToizwN7eEbFVWe6IDUBjsh+8S
oCrEvUjqdXEqHJqYvonTRU72W7UXRQrKdUBfM0r4Dg4OuSMf2XohSTRn1EW1jXiARS2Fa9zC43aw
9a3lzwM7vKDiRxFbe/Zh1Afq+lqr172qzl5F1ed/uuHuzIop+4+5qbFvdGIQFwKNojYnNQYXr9Zw
RyLJbR45SfIUZS1BGobHKRdiO2dsr6L49ozD8b6iqLF43yCc6RnDshL535CcJ+qP7FfBXK/3tNmB
9eRdS3j7R9RzRhR0OmyuV0G9ZlILxQ7gRXZUSaucrW4gxRbNS+wYWqBZuLV/Jj8wVyJn/BOG7v/5
ZY989Zb0YZz8zcM+JnHErF9SQ3JCBpkyxDHh5SQfJYDky3vvq1Xd95bFBwmeuEnPXFZJvkSyq7u2
bNqW0ZoPCJSWcJ5Zwn7UAv2yZJT53+rVpUTUNj2tBdKxqpK7B4LKIFIFp64lowMMxPnEY9v+cSRh
YrJfVXK/Qr5hCTJ/7e/u9+uSvMr1x+ZX+RWGwRQ23FgrPMxEsD1juD9L13PczuGNbT/fQYfNvZWu
fy28aY/SXOacIIF1frbynIRrhvsTvT8VOrNDT1rgOUlTMZRzthheHMZQDZiPTg/n0UZRmv0ZXzzz
YGmK+V056d1doeNKTDs2Zb4SLCfVuNoaW2UWkmuQ35fator0B4ITT9tFujSYJBK00N8NcTWIm9vJ
cgHG1VXxrFnYqv/J8m14ubaEkN9t1ZcVySVwslmLTSP85g3qDYcJTi71SgYKVRkEKCm1AdrpKQlf
YnEaE9e5w/K77Lch1iur25lPD6TliQHB16ksECebty1r3uVBs5bIRnEeGeRCFz0X/Cx85A8n57r8
9ClHm8OCPJJM1/WLL55wVZHArKmksHPxtiGrt7XMYXpfBJpIDUAI+LmG4mnLKY1mH1lHrBRAtl7P
KLP+1o9HIN3fkgUvZo88dw5ux1ekHxLpU0jQr7QWrFHvFbgo5WyWQo7OVZYgqI/JvKecbZmr5BKu
W24s3GGs0N5//4XX3k97+BMf6gBfbIumE3nxahiWlvh5emQ1dMHCtIt+GKJ9RybBHpDvqNss0Mat
D7IwUSdcJU2EAxDDay8KVpJXwHB42l4C3fV0Iw9ukeybICozwQRTWNYOi+1v+8vrP9LTaQRUchv/
dA/2Sgq4F/6o3cPJw/9eAFoPZMJI8D+9i3JgvGjX7HOSncLpY8jJiHY+uQY1GZmJYDblytO2ow0D
nNl4OTXJXSQBY+x7/n7GJK1EPLIZHw8CiHAQCf04c88a2S3BZQfDkI15ED8/TC//ttMhlWJp+xLI
u15FsCdkrR77/QjPA0oNVEQfKJFpR6NhxBytgbCfenTNbtjshRestd9LMvbkSZqSa/vnPS8DvJOC
AzZiu6gSZEh8UvoWey61TkAZAhk1DFBuwRDb6apeTtuWyrfzyig2nmq/Ay+2HGgcHU/qW4+l7nrq
AKv55Le8wPMKovfTs2Ors3rCsEPRP4e+WlzUUYi6bfWHzt+cjTF87TkTfiP4Livzza3L9kkC/imA
mtwzlbpYbat+5LfpUjVynYk2oY1PlNjVXbSYXY/uBTGbxubjM4uNJ+q/Cj+rh7C5AeoRv46UlQ8G
tKO5bSKFGTywGHfK7IqS4dpUqlpDFAcTOIkeBLycHR00COsgGghsLZKMZ+f2H7LTqeUQUEEGGpuY
bLHLA6v68jGqtR/uoti1ibhtEXdyDIs9wKBehH4y+IXPfmyOHD+RHAromyWEQXs+OU+tvzuvKyaS
ZHdzAkPTaOZMEh+IsQDKvQlbQf+0ZHyDXy5PM93fCAd45Q3VbIp8BYkV8rzy7nyF4Q85Tl79NesW
j6V03KXSBzYCvrmd2Inkq73TErqU+CcgOV4zz8ajs1UxFI+0zOWcyHbCmfUV5ztVy7LkjXHvPdyL
nJy0Nxr0KARMYjYguHKbatAmYJlxpokPJD5NOGoLDUQaB6QzqmhFqzjGzFBf0f9NbAJymdmE+ZJc
qnTwV6jma5je2gElMa9d2VmZHivL0ytf2tnj7xv3YOenENaCo0BeCdsvE7z9huKl964blncQObWY
ZKezC83V8Uc3KWuhvQP15H9EtS/vhV1EXEPLb2R8n3wSSKxoi/XRFIh1ZFDJ8NizOopwXhM855UG
E+oDXAav8ygaz25XEwJtw0Q2NL3vYt6i2HH/MuWdkwT79wQgoZzt7IAn4bs/rs0RfpumVWbg4+Px
yfNWlVawdcTc5CASuz5rZV24xXctuWGny8fo4e9naqn3lHJid/VycYE0cOuE0lKPmDtUbWt1jkB9
gHWDPca5gI/JyB0WYzDu7P1NLCLe1Y/SJGv5/yVWTq83SjS7tS+6kQT+1mZV36GWTHx+KiDEHdQN
jihv/yBBNhF4k6RaFh4P9i5qSQmFTeVJxDPHa5n8p2saWHYmFsfx26pyntZPW4j0kLoPNp/zPsJc
4HTZQvemrvIrF1g4rh4gNAvY/48zKnaT08tV8Gj1K7RlzDw+NkV9VSimQa35GnV+sp1vmqM4CpV1
eTnb2fcyVQMeHI/h9LOJEBG9AjcAwCFxXdd+mZGhU2cjyFfuMpWUbLLGBxzQfWiUXLQ7beIX31IM
m7cXHYy9NkZbfcNhUL06p13GI4wRKU5Qf0i6LhSJSKrEg9SJCpqv54LHHdiZ0ertqab2jaeK39jx
POJ8uv9arIQM9tfjxpTyoKrCtnqintqki4RVjk7Nh0il7elfn5GjPPxVLFlY7JZXtkoFd95QJ1LT
dUnG2CtuBaINbDWlKue82nzAMDfSABepeCcfQgg6Cg1XeRWcZLX8/S79f2i1rr+wrsZTvk/tXGo0
/EY5MPJ/vtxYR2xZD4cyg0ZEDoQWJRLe1VtwwitGbfRpG44aXW7VeLjqbqBMJg2ga/xlhJPTQ2W0
M2ugJQURES/8ZBlf+kPpufHSZkJLjn/4KRRS9e5k5T4ylumw6B64OzPtcH96JJ4RqfBGTKS8JRiE
Epi53XL8lWr3QaIjECSl5rAy8wg02aMtoYoeSDE6K76Yp5aiknM43hWuYMisx36X4L/f1wigdduB
eYq1i0oQcKRcnozlCxv34WVTGNJohyq1tnZpO/lFjm8ogiLAhYAn80HxbAu/9R+veoaQyEFbVweW
leP3ZB1adc5WVqMJ+9Pu2+vetgKtqH/9n6e5mTXY85RZklspFEtL/ILFNtipLo3CsAS2HQtySXxC
jWxEdreJJNJ1/kWRbbaCYAgSvW3Pr5RRsnPyNbGTvduWMZzlJrIOlYOjGcvV2pqstgVeaIVb3NEy
1W+Sgci/OraGAM8GXHy+JVkHbR+SiP5ow5QGZMoakfmHVgdEkrfP3RAUD4fjMC70XYwx7F91WFso
sO0XCQQD7f0dnyD5yfjD6efmChqDkSTNsOYoYI2AdW15jRVktAqbyp2WB47OfMRCpFd9blo06I3w
+R8W3SyuZjXlqCpqWmGjx5cgmkc95zNfl8Ty8D2rz1wQjO99/gRth3AR1OeCwetbwGzyr+s2QHqc
uSBaCfCsTdjx5f2UfD9VnRmACNr+ZMTD8dhlvL8IHMr5CickQI+FNnZ9Y0vV1OK9Rs7S07eqAgOu
fan0C96n8PpLEjySK7YpwLKsIlT4dGdQNr+WlJMeVZ9lOeQyvJEAPW3XBhgxGDdILNoSro1I/pLw
1nYCCBlDneNy8itL13f8eL9vmkgMoniPB6UgYSKdPJFwKCVTOr9E6TrxZij3BFHh2DlJec67cHHu
VSpiDDCBJkeGbQz1ma79Tp6yVrRHFcgvJs52uFXcrlf3tNs/HwTKNBObWE+8X7HWgaHwtbqrCyZy
yDqsKVix+HpDqUiaZ1IsaRssLQP/QTtR2iU8eiowv2AjxJ+LiBX9LPxEKq57J5JdwROPxXEw9c7w
q+o76OxBNdk0jyVXXaT4ZtCbKGUGo3ajPPvehsQ2F7iGl35jJzzPexOUI2/Csm5qHUWTzTIbTHT2
7I6D2QivRZxMkJuuyzqADRr4XhvsdQsvzR3HpshSBrxFinpqDZN+Kk6QkegbLsFCQW6ywmm5DDGv
jr72+n23krXVqcrCEBxQ4ydC8+qZkD0i0jw7+D5H2V5sTKpOapSMo4ZDVHs7EFGXjnUMF56Ljxl7
5D/9wxGJ3zKo+dNRSazZEmalVnpsOArlIkByJloEvEu9i/HunOW/uoVdDYGG9dSIpFAMpCMqkDh/
QUYCcygBxn6Rma7KtGDinlWR+LJ07Q/GJ1SnFLMh/o7IQXKzHPL29VY6wYy6+esODo3dnE5i9JH7
beSMaLEjK2dbhlOsQ3g94maI56M8DMz0ULgHyImnUsyzmR5hLXr5aJsshcaYcRmWJr0OBMBau9B5
IhgyFAHO0ETskQgkYNHxWWSU19TkwYqGfziquOA/xSbfOhcl0fkjFFgBZU29pfFFyaAc/Ic9ZmZR
yf4w2HIuoipLGl19mGQtA+1v7yXNsExt9UVXjVplQsFtjcX4Uk3DNNNz/E+7NaFkgUJMYZpVXkAx
K4hchyU1uRH8Xg2y0s3OHr4Lhyx95et9dk0BRVbA3Eg/GB1oEuBNpm87IRHL/34ChrbuL0OQNsSh
XZC7fFw5dFQTCEvajutiHga4PSvclnQJhtFTyCKVvmBnhZB8BQ6oS4PezPXNM7ErU9qNkytFpta/
k0Hwy1TJId3tyGeBqmVObdLmar52z0og1CUFoSeF08giuzleEOAxYdzJgqTKpiSlKZeThLik6vU1
KITdLCnK6UE5xk0ZBcvlmdMFafBJWed0fLiX5SS2P1i0HchTtm4sz7I5pdp9LJF/JwWzv7Y6Fhcw
AF/tD+0hNb6J242P3DZ1aTtfU44q7ihuiZpTUqP2orp+Hd/xz7upCJHvIaYDFv2RGFKwA39+jWfR
XKVgtTf1cEbSlEkaIBd+apPjIArBEDbWwmRoHWKWW7i9jNK2lG2o/kDTBD3KAPe5t5xWrFoy5//E
YJEUS/nl/FOBpadL6Lrmopt9LHw+4IOhtQkDHXaSZhhcuUJIYE4CLYSxG92dHOhtlx6WHFz/nVwm
2wZnMg1aemdbf8Dw0aZtyF2EfHYJTQATVf2dPvFn4h4/nIG/MLcfYtW6Hni9X+TJsSoA7T0TtHHt
eGp6ab45/hgU/QTWeY9AOL5pkzYcIJ/7a+SXpdorv0rgM5mi+LbKmZFfchKv9gjuALQcSnNqih2A
9TYm6bk4SVFQueFocfSVFxIkWCmmlMZ4BcsLBrPB0cIxNva3iLBEP2KZ4FvMGD1XfDzjDz7gnTs7
7JKaDJbo2a9tHvrsGp1pra8AyjH3uBYgeTyl3/+zt6xWPx/eB9zBW8UwvnFpn3ZU09/abWML/St2
bzy++mF5v+TJBhNiT/e0u2vzQTG7dnHbwaOzB8ZwzYH7lw2FAf19O8yCMZKF4NdOq8fAWEdVttwY
ng14iMfI0X/pG8GRjh83uM4BkimTLnGCgRaaT48nyfB0H+zP5WPvZ7OMI3POodAjydirmPlXdqvL
KaWdWlDi+5/BPFtBMu5EPqFgYSL2jprD7YCfOTNIMaUHjd4t9V9LhiBnsutitvCStVJ01LONy0r+
1s2WJJRllGa8h3b69zqer1eenXSb9RpEkn7+j/SyS1gzelSE6lrE8gocpz4coeffug/IX6GSHNTV
SNADWh8NnxqnnqQ0FT5HZiSz/rA28fBy/XgoXMcCful0Id2viJyMi4p1SgBWbb5nHBT1QT3zU2Nj
6B5lKWyI/Ddw4gMG+SCgnXakcK8Wz7eHH8YXJElVv2R8H/TpZ4k1gdZ7WeJvX7bnCoQ/UPjG7LFb
dEtZO3y6Raz3LMSGqzLwxWAQZKeGIFsleGa3gcnOdUjTUtgjZWo6NXTcwYk+FFCqTJgLW22chBso
OSQZ+gG2CB2PPaFyX/xp9++lTV6Hmdnrr5q6t5Pn1fZJipeTKemwPAVTP+Tw93Wkui3cO9ZGLJYc
cV5jCalcsypwipwPM9AV6smScYZkAkJW9yeFLzXDhbJPogWXmKZTiB6eeNXdsffioZ4ccCRQVc/q
IA4hIoqHUTwG+igPQKRrBU3l1AZNyF22IqQu5XJwl8LpB3TrwujDS3FOj83bDvmzJQ79g/lP0X+K
koOwdU4NgDvIe0H0SmiZNFcyk/EaS8WRJTtkJnTza08LsxjF3ltNSEitiOGkfYNn3vhqSsIPJAjC
n3eQ/8679qNpHudkPuLEesFLr4PGRUY8+WNh3ICKi8NcQTjajrxA7Jbe7qW9telKFqp/VHaZg0bW
fTahR/DW/OyCwmXoDmPMm96Ikbub5sWR9o4zi7cXSnpC/8F6BHzeH86JaOpEmgqwVnNmgx87PCC+
CKkSf27YxJsvDKmMlzt9j/yfWYCkRK/zbgYsQ4TrRHkgXMwincQt7zD0HalJhsCCkuQ0Pr0pSMxW
EUvAoKaeaKPHqF08Xho5JXHjoOPsKakb5pHYXTL5eewsQVckGtph5PRfkj+rvCTcDoTQXww9Ds96
vaGH/hL7OBQlypREidDA5a03L02luGx0INHZkKv5fOclwUPTcD+jKcyAPw8Cc/AP03i0kv1WCpHe
Z6l0xn6j8LP9pt3nIwtReDMgWbycJ9g1Izwsq3DPRlEsPNuuhfj+nvoVZShkmiHgO5euWRPU/65T
I3zzNLUQt+J0joSe4nXrCFsM0iXsijGEhgBkb4E4xk2mqyXslXcotPiM64iFEQisv0ZkJBPycAQI
zfn6NI95Y61M4MpQP9SQy/TamsfmOybwcKzq5eQpv99kLEV+hSJMkuFkm1CWBT3tQvidlOpvvrvn
Jggt9KnR41FwNOGSi284VnmYrqkBZKKp83LdnzFcBkjhRCQ9ZS0lYTyfUoARSOZQ32bR8hF5ZHP1
Z0cF5BtrZ1ZV9vPFHeksFdq1DCgbWrFsRf4jqXzsvnrS0sMuq3Nglyu0v6B9aTpqKDtZVMNzIgKe
kUEKspajFDtd04lKWClh8wj1kz52yVm7rDxmmZvk4HqdMsBJHSrqsyFJmuDMi4MfzfKUV2dpa8/x
OFl22j8GuziivYRJOHapmPe5FGy8T7U6VMNApNPrwILguj7hQKhqDv8ZF6QMxkcwguJEg1kcGs1H
+jwwggC9uuVnbb18PipWEVpr6rYtPe2b6F3+yy0ftvWgXOI5tQlIrA2ubGOrBTLSWVIrh8M6mB97
S8zgABXQppDLS6CaTl36uu91uzwTznPhkjEnZT6LVIvjvkPZ8WC6pShEJreO/ifNHC8xAQcK//PV
P1dYpXjjSUiLwd/nBRgouwWGGfqwbv7xsRCSfpYqLKz8to0JxPyE6eE6vAKaK/1lVBakGfvGks1t
mPmvJA4iu1fuJ22gaTj+slqLwLTRJiXvhOUyaZNWIm+FD04y851Lc04fTfXO4+AVk3fo4u7SwT7P
5IrHT+OcryZ3A5UpoTvidQCXkI6hWcG8Z2fOVLdbs09rx6RIRpIcX7XFuKnr13UU/e+2pVZDMNGZ
d1Z+CZQvsmWwErhPedeSgf7RUbbqkHuo9tzihoFjC4L8mqIDDbq8e6evddY0OBWGKoP36s1/btNA
3tWRLUXcIGT1pNd+ADqHK3WG8gJlZHvxkO4RO8t95oEiGJZB0sI2Wo0t8VFf/qKgkcPEBKQq1HiS
GJA2uOhZs+GTTw/KjOYm0UJIGWRawOMjCk3CTzCgXByAxlYKadhiaTJnQOxIw/c+otzdvRjitOfe
tr0AOQDBnWhh8eEksZCU+fILpffDNkq92O6empJOTbAHcn3jd4xn+on46TqTeiwEwkF6waViMu6G
CPQHSUS0H5j0zK3A8ZojnIKozeD+/wC2QDpRDHRUFkFR2sAGjkkt0CwFt3FEpqEBylEXfAKsZP5Z
GaLeanKQcW9sK8BeHTWXfiRBBH8zprs9rt61iU4/3bL+zQzRX4Cxm/npXfTdjdgVVx+ag7vFB1tx
XC2DvUTTkkORZqa0lkq7nWdQsz/uvSZCSNzxjyEEE/HQprMsIXUiD4x+etm2tsuhGQv+GAu6qx5b
Cvk4H40oECcMTh3GuqjZYmPHqdJaIRbDtuQw48zBH2Pugq0cP2sZxqEQ6Zu+WMgPI4oFkRosaryW
RTo5Pcvx0mrZMttWzm1VS1gYyuTMoAFsAGz+JvIC61Mila6noTWOg26F/J2/Rmvcd4uOIUtUKnuK
HUCzFXF6tDL2UW5L2lComBqbZ+xeqjmv7dVzCVp7Ap8fY7WpacwJf+0FMqdKbBRFHDroJvvPT8E+
DSBd+/llScLS1+eNAVQT3RnMr0tymHE5DXgRHwuMkPW6IyCLcZfmLP65gqQXrM73Byj44bTYTGIb
e1/uvoGHPkUeGR7Y3Q20klW38Zai7pB8GsUTToeqMc3qGPDwXtscg5jce7lF58OXUvTf7OmSgMzo
zEm1p1CTlNas8ydS0ie2uLNDPXfjGAK/JrXh/46IHTls5qsbkZM4/V/ql8qRGMzyMqfUjFVtRpcb
zrkTRAZjuDtXC7DE2pB2+3pmNsmUT4/6ZilcKzFvF+uI/i3bw9Oazfi5VhcZ3DEEA6+jTXGdeqyb
cXmkaWr91D01P9gMm9CJKaut7P7vPI/gHcVh8PWeg/8/YSGP8WlPDFKiiUTGYQLJfxreQZZ2d+5Y
RJAm+LpVtLdrSgRy3ZQzQYptdfUAOLGsvIdm8TfH32fJQGvT7nXbSBANKmnN6elcI4dk1AtbQaaR
me0qy6YMJe0sAeqfXqSxwLj2ILk+0bpufMnZyk8Ow4ao3azXA6O0erq4p91VX6AmaUYFlZO12CZy
7TN/KmRSloABlKqi37aqDW1DlXZpkOyElQwsBsKutc18HJAacK7d5oSAz2r6HNaV1QexP4wqU4Pz
ZsZ7r+7XYCtXjoTAyoB2IcIwZIkwaRHtopwIGNkjUcRC0bzzcvZdhzPJyyLw1/MFo29UCu5l7dUs
ItOeX3V/JdaEfKcqTaY4tVKc8GPAA0oic9LGeUXGYRI2WseRBvp6BSIogj+j6IGyT2RUsx/0w1xc
kKwuqv33R4erpjuuNRPGdGjNYYytO7HZEdYn9nAUbbG1AsBLvZhwR87BoVPRYMCYcPId02hc0Sh3
mxANIZ7tMYy3IB8mSn9DtUsAzl/XTitDkMJymezaONWuhPET2Dd+4eTHB5heQKrwfslf7mSKgchG
caLumJgP4XpX3kaY3OIpbk/IMPQ3rxTqwUWGXLF7JaIE+QwYSe7PU06VSJcpkbzm50G9o1VTX1/1
ZnlLXUK96BS3NRd4yjQeDgXtkGQoB1BfEuM7Sw4c8mFzeHPnQrraDo1jlzcHXBmZ5pka3VhxiSlg
waZNLb4JCkPMQd8Qqxkv4hEqQctvZIluRGrBdXNrq9m8N3KStIu+r+HtXiNLEyMwxeAkAaFdxF/4
KU85mxDx1kI5OZnbXD0AMk3yUWp+rSwtr18c7q94bLpo0fa+moguCdx6808IsW32m4v3JkKKpihC
94Vg72MsfMbY3GUVEEBqfemUIuSN7XESrfBtiqfxc2fbGJKOJtXrQE7jDflUWNKLbXnH9a4RovkG
HrBpYdVPCf3MQwvPDY6ksvtqyvB3xraXsqsxUnj8Nr74tceTrK3YmAf9dU04C04t29RXkRxmX2hE
AKRij2n+CJ5K6Knm8LlhrUsg64O+WIlEbHWu1a5Qp1Gu1osVaUNzuvky/GEGAOU6yVCOiWuJs4nu
qAZDIoc1DdUpaIJTw3swUng6qC5DquYMZDx6SSm6sor44atkai2mclQS9dTZDOxtQfX8HIi12sF6
HlVO1hOwTu+wY1g78Wa8Wgf+Iz+s7NZT9O7AgwxNR9pEA4vobZHEgQq4r+kw/o0s3Ay6TcujCsm5
1GCPzBVFU++byfMHBJrYr7uvI9FG8FbKeMzJtVOaTsNNFl/4znslANpbpr/l0jPYHtZutC5oTrTv
AavXiLPQ/86dkC7LgHE+n2c6BPEeQqMuL0uOljNUCBXGXgRqar7gW2bvOJz4j2D9K7Op69/QfWmV
6APtR27Tzusu20HeFrqqsLHjkj436fi1mrWvO1xCpd113ctW1QcVAFj/7ylYyG3wisoPzBa2EHqc
00jhVKxFwRzzOfyA9p516iTbUWjOqihfegaSi8jJRmSfykl//Prl7KGfeSbsWlBpeFEpcdgKWgRI
Idu0H/m/2l+MzRVB7s/On1O4pVAgEAUz+k8gNuINBT4HXc9Yes9/p9+Hh6y6KahTj2OWJHUedW45
UnMyF5KyGsYzoq1NIKnArC4aYnech+fWm1zPaRAcNEvAjkOfXRt24s3RVKg1+yAjzxJ36LqJdDuC
kn9NMJ+V1da9KySD5LNwlN2YjLMGNx8yKN17JxOkOdLtj1XoypI+uDIGnSiJJGfPneSNwTy5wf9N
MsfwYTS+5XnkQcpXLn4I8sGMXvXwbu6v4ZNYYEocSkwCseTy1bY+YebO1A6SuG3Hf5xxGidlVxTk
6I9P6HBN3/yQhCt8PVpFc8E/hIm8mBAwqpFPD5u1a1SvIF/0logVf5XTLph/mCY7J4NCGgAE8xrO
KSqcweWqmW06q/m9wKGtzfulIk/WTYGbgkFSUMKJnKWuqd9LDVXIFlN8RWRcGE6a5GLE+ucaL5aR
RVYujtQRj8MIOC7b5D3uWvXKW9q1Zz2Sgc1E/u8P8yKwP46C3EP48i2TP5PFK9dJds2ag4REGOd7
3Fp8nBMaoMDcwKN4g34qE3qJRKZX2fhLymdJC3nNaBhq3zFB9P0Oo1NASDQRqaMyQTctSEOI2Cmv
BK4AmuDDSL5/wwV5AZpHPtzD1enkRpaBd9l/N8vQeoCS9PgmMmUnKwEd1wOZnHPAy5GyEg1Gg5Fk
24+mClp9lLNtplHZA5XkHGfLHJWem9f3MFlVsO9j2lDcNDIhHL3ozQN7JCVLALq41J080sL72O+d
XDPZ5i6pYMGvZO2O8gJgIAY2m6aJr43St73/uTBtCYs04JwZCJfM9kaExd5Cu/b70dI81/ka4UXy
itIzo3NU4WhD1PaMKyp06XxjGz7m9ZblZncwtgWJkTxm1+f9IhlJa1hV43iQA3yy855T6Yk366yW
Z+Cbp6HoY2HBLOdmyfFd3b2/6+eP8Vw6sDZi2gajKvbNZanKCobY5Y+KKhQvNlrFQ7jV9wJE4YsZ
XJ8KXlZf/+LyUsBxSR2WNu//omlT9wgbbZPwkQIajqM+b1/jWNDJJrt8iowGasQ98lWg7yN1uU5P
H3C+9o/nfWOQRF3v3NRIMYsnQUBwXOXvnAWs8rvqcHvk+waWKBbW+TZNfXnvfnWbDx4NSQtBF/sF
h3U2YHppnZWtlPKCPZkoivT+jUW5u+DD4PBQsosibBoz8jyXB0mFUvWD9/nEFr3+D6OxcBmeW0Z0
qBvp6PJxRrltpOlk3Pf6vz+wh8FTVXzKUA3a0WmbRv8m8zMz94IbB3PXo8w1rm+DuoVF4Vp96Vf6
61+YF9VE0r9ZY6g90tWyFTw3ZMjf3QnJRUmE+mE/XcBGKlH6G3bkAz4NSRHIB73wZWy0vBzg+ZCM
N+rMlof/u5hA/9/u6Cdjlru46tuLgq/G5MF2u/v7l2LTNsLGVocdLn7n8AtuaeJUeKDTRAUskkk2
3SHqrWFwr9U0wpqgTQH72uXiuOqB0ZHVB1zsfvtTQhN2pVRyz1WCZ1LzxIiJaPec6o2fNfmht5ZE
xy0i9RVB/ZgBrTfMH1FkFI6hqS38xBWkRGzvR5odRlt+lmC56UGufY7FXTM522SoUHtuNWgXTQjT
kSRvpo63X7kupIhHPcOgYm6+vzhQ6IEFEyeI8/8J84IKyNQXfUUcCZ/F+gYGwFAH7L6T6Qno8Cam
OaceszcFXpbWE8c1v186Kd3+rRwEFM/zBSYQPqkWl82wYSxo2ekQmdzubLFglZiLAbwU0guf4pob
aYQO3/932jXIZuoGOtYT9AvJRj6Uy5zE0irNJr7rERawWTk/DIaKBGNFLb/7NrmoAD57lmoaMuvu
+XoEcgCHq/hu3DFMYjZoujZuK1FK4x1mdWrV48QxINtIX2rc9Z1xl/N+gwDbIv/l0tVrjsn4Q3eC
//iEhDrQsE1ULQ57ZcR1awD/yOalUrcW4JIP46jS7j+eftJdhu+TK5fWXzG9faYrZHVuq3GJxuRh
p3TjP/YWrk9UdPJg33aQy1nGAoQVU5cN03zY+Fvfumzt3NeWoUx4RbcTLYnJ6CRvWJE78voaa6V5
j0rVt+x7L0/auuaR9t0Mmak4IcMYxBn7n/gv9vG/6+7vp7V9nE0NxvI6TwqP8wZ/MKUAtAePQlO/
+y+9rR6YeBZYdxkqPUB9aSqRH4x972EQdqh9ZUBuBQv8IXOFWZyvYd075fvp32MffGo2LVVdDYlv
7wyOXUutVeKCqN3bb/caciiDssf6SFe25OGDEX6i5fHJpNHaRH0Ak11EPYA/lvgcrlbArg4xLuy/
8mlngova3i21eXxV4lWLpe4G6TN1/92zJ/s6a8ux+zv15qaKMAdBJDYQh5gJr0+Q7vXsdUqbMHxy
LH99PWIALV7FPkagiEBF74jdXHesJU73CX/F4OF6Q4DAcJONu/OENmsyO6g5yv4k4zGhv7LJtipg
zn4tAlIrWJVOXENAb9nQivQFS4QyLyXJZfiSDmgZ6D+O455+6rhDX6lY4BuTVBX+itoaFeoDs//A
Qed/ih91HC5T1dIEmQaqONOlH27Dezkk+NHcIUW/KU5NH5vr3bR94UJQKFL6s3ZJECohGUSgYC0d
B9znm0/fn/jyfSHo4g15oMledvtzDhM0NFYzK11hXfWcYR1Fzh/iQ4UTGSc9gh8VJjskYcZjG2Ga
R+b0pnFRY/9S7dlCvbkNEGhhJ2hXqbEw4kFYENxcySs5tkdh8fR9YDt8oTq2pdH93IckES+Rvvxb
Um4O8oYS5rhAQCJQtADl32hVyO7DNqT1imsmDS9ew5LCgmJ+YzbiSCWfsHfb9RAcII/wFTggVlgd
vVMOWvNUpeouISbZKkgekVUDywB9IzWJrVTpPr5kCHGunS4zrkFJmVSZyr2Ni2yjmwTO7yg1xUGb
wAc+VnysjvDb5rps+Zxn4O9P/KsSqjKUp9cyHG+H7kPhh6ZCb7ZKyO3y3/60y1UwNFlwSLWWxLCw
FI76pK8I3yRFqHh+D4zekhOUBk3gQCv0WZeW79FUv9yt4eQl/7msLJTKmAdETTF8bPjXksCnR0wL
jsPRSrEWL8RoT54fgtEWrbk6V9Zhz2bwQldNKKg2LHifmfduSPAN17O/r3iNWgq/Oldd4VsPGVwl
2lcf0eocRJKGVsUAWZg3m7ZZY0VX7nuH7Of2MqphAm/7pGpSpQLDBMzsx/gQE80mXHvpxgSpSaw/
t7LIdnSItHJBzwSP4NOnWktgsdNUcc3eppYsu/rRpRJhzmA6WxShQETGk67K6BscXsUqZy9pw1iC
wkSETQ8mjP7Yg+GUtymJpN0c+NCmHep/KWwrCUHdwVRfcyunZSp2PSl6WJ94FjBBXI3F+Y4Bnkw5
+tw+MIEqeWkQaenH15tHgWhBf9bSh3pAyqwebNi+vXOMIWJsW0ElRcbVFMRRSk8p/3edrblE7dlZ
owaMsRokSGAgFcCBAT4Vqnx2Js+nP2l9y70HT+RantW5wXYuW6pWdNeWjpgzlLojtSpRh8sFVnHa
N4SxW5Lar4EtqOMJHU/js9SkvARxQnrxQG3nnR3QUGH2x2Hlh8wLZu3Bxyr06tuWLLVCN0rwLdWJ
j//L2h1cgJqesk47IxlcDt/AT3sqGiM652Wo+FtCeyzLxzMI/treekmbJB3bch2UAvZPaev7O+4O
RSyxha7oesFM2AoUoITAUIt/OHY/vBIl+t8iLTj/OuMkkqEokHo95gXBrKZHmHjdJ503OxMxr5kj
BOoriJvMTsfv94gijo2jMn1xRFvZKJ1EyeqMRNQDWJrOX/yUEJq9XFD1LHUGaCCB0iOIKr73oA4c
LHUh63UPxCIxvZj4ZzmNk+0uoDbuyy+yD9sMlJkxNW28ZnHvXWYPBnZYnf8QPzmzt1g67Zys7pvS
eZuEzxeUM0yAuhVCdKGaQkHUxhA9Nd7jDXrykry5mApdibS92Ll8Xh3yAM3YB34MuU8WX6xAhe4h
4PjxMC0SAwqiFD67FGNQdCdmfuBMElQvMdlo3Xuft0GEg0j0liOiPQ9hEhkewWjUrD0e/P6b2HBA
K07o4zOUzmZO7mEgkE8vGN95MHEShyoi/j9r145RW7wojBoaeCTH8vK7sAJozgBIfybn1CV46pmj
gzEMz+T1x/fnYmluKJ6HlUA2tkpvip1+k5BI5gqr82i8fRgmQ8mjuwFJ9L7a1IEMW9aAsdKgX7dJ
5bEU9EgTxjKZol44FQoqXW36K2+GB3pRUEbKs+J/jp6tL6O9Tlcjs6KTpwre5EjwnT7L2HOi6xsR
GqavWEXGpV2ZXgu3WD88KJjKg/P+xruSGDoNYtWhkDMojDZuR1mVnwOn37RKy7Hxs4aIO2JI5sDJ
0oIue3cg2Gv/RYOiebRXD2sWSOm8R5Mm8/axvxZxV57wJq1zeZyTGtIboDwuxDGRlE9KRZoqHm0t
y81S8lMxXvIPjRxNRkMvcCLtEoiWJ2wSkmTo3Rvb3TCl/y5BbCmuahpsJ8nHLfIkeEqFSPw8qE0E
j534jUShjWhlH3Lcr2lTJ8/4dEWVuSzaUtiDwUn1Ge8dx2BE4duSBJ/fggBLyu2mYSLnnwHoHaSK
sDJVN13GG/IsMe653lE8/4TRb/B7K6bauF6NceXwdR6UKLWBizMMS0UV4idJeqrWYqEVOw80ZKlQ
FO53BzsCH7fXeeXAqGRqdA+yIUFve8pOIq899J9zrxWAvwNkmvs49WZ0UJ+bs9j5sw1cxblJ1gzl
6KQyH2iLwbz7tTbvfzY+I19MQc2LmBSOP1qzTd/9K/9KFBkyINieIebP23A7kRWKdP8BnKlZPDbW
iki9o/WCxJMjRl2GPIX1mWH+YD4Ph91xhfm9rqqNVAo3icDhMKE4jrG4NGcO1nGh/i0wkvRs7SEA
gaqYxyrzpf2h8bscuPbmqq5UNdBVHQA0yDvpvI/vQ/723JS0L1I51AMYHRFHCLrPZzvN3UjVwiza
pL3fPEI2HZJ50io5QaeJV6BkQb6VG4gJ022G4OMAxZ7V41zGWGjszxFP6bS8DiZMKzhmRbjSelVJ
ZoacKEgytGZbuFedMDb9w7FiGWbDaQS4/dKNScZZcCra7gQsBYXE6tpPHsugXoCF0eBx1DTDKNEH
oooYvieyvE+DWSpeOEIXotq5z4dNXBLIVeaxNCrdJj8ufBCfC+7CtWTKcQ2n+8gT3C6/fbZaRj7U
xg2fKlik+fB0V1l+cp/JdoShVK4kKYG2FXWVMFA1NwJAOuVCd3zqML8eEN/F9MyYHRSkyFv5F36i
4RbKieOrlAiYCTCiJfetl/3E7t6kVCGXgKbfluk+TTWygCZk3dtw1wKaRLz+nRtyZB91H1wYlK9+
pabsuEZVniXXNsrdgNSEsxlohuUnElm8bOqrbLpDX6KhrpB2u7qRD0yzkWM7FJwDyDKKLMdEYdla
e7tx3qfxfYfUq/Eelo44/7BXZ7MfL6laktgL4uJ0pyIxhcxObyyp1L261cMgoiWGhncQ0BvKeZTc
pDr4uo6x3TyoNtMFDP72veLZeHxp1oHSaROl2Mlrgx8NfMe4oozhryf3l3/DWK8HMgDU56cV7WUU
UpIHeibugAy0EZGwU5UhDRNlVbOTZfKa8VNPePBFgckNo4u3K4mgFjN+Ga8wv5lvIhVoPzY5j1Xn
dXSi0JDW0z/f4WnQQo+lKvmRATHSJwyotb+tCZE9i2ZKlrhsd7vMZkygV7bKncqHBdlTyON/ku3s
4cMRcCUogNqUPE/X/mNOmTbm4lyd6PMaRbP2nmYPfOG8y0BpzclBPk0anqu0lXS8k8H2Y4FX6k7C
5xklM9GMEqI7pNgMLmdIJo6Ujh+5Ln1lf0myaXep/0x4c5VTC/+BhwTYhM5uBQmh299oLkyMoKYN
gAF+npdH6u7pr+8iM3/Fdm2Axu51OrEXpw/dyKpt3A1NFyQULHczojKWvIl+2yBvwgmcGKtYSd24
AN3mqTwNkafIed+psEbTvaH7NlIJZia2gaPxSemUXvbjRdv+XWkqSM4TeD/FM8fZveGjWkieFsnk
XbpCnoCBMN4GH0nRPtgmHV2o3Lz1Plj5KMPmTqiGwhzzDgLwSFTpGRrBhz6emiWn149D3AYpQJAC
LB2j0AFCzqg/LA4FL37Bma6hgfMrOOi/n56x8SB/XeAMuuMELD+kmllAsGfSzb7FSZktxDKMWKPO
c4wUdFTYg0leNj4X0MeSeWPBwzER87zg2Lr/J3Pwl8X0WLAfVW1nFu8Hb1ifbO52u7M6uLvN73LY
7l9JhPz1gp4AeSN1L0Rzh/0dUFCDTUw+PLrC9sYDgYHKISYPZS/tk9NfegRC7d5yWpiKQQ1cYFho
W+zZjCWmisNfMs0rcB95uf4FbgcR85h00McjFS7zgjbHbA2JXuBbFXOzBahABIeBoQj7Dfbvfhzu
ryTmEUJxTNPCXzGN9drtyftFgH4/BVoz7ZpdHb7tGtWpPCs9BQsj29ofCD3ihXn1xfhJn+eQb02v
J3nK+ARehmeF1df0w8Ih44z3mO1k5ZAAY6mwBddNHDJ53RtDNy5J1lfCjl4Rh3m9J9QHX9Eimwo6
FRe0Qo01WddyENDpIck9zFvXK8s7r2IOfMtq9o/4G6pK60ee1csS6CgT80Gg77JtL5Oy8EwBWhCG
983CehyaAddG1Z1ivaAN8inI0xo1xbfDxj4LGtMYmx/Nso3eLzrbhj3HPt6Y/cwp65xF6RJZ/SJq
AjNPTqo6jmoYugk04+if+PzxngoAQmoJbD7GATQvJM1Fh2VUQDWkyd7OFVYraFbZx9gAR1ZsgM/v
XMOwkoVuHwRI3Fx6PEXZXerZmhgAnBAOTjeaxivl3Itadx++yh83el/r4lfjg2zagk2Buw599grn
Ov9rhwEdgNndfcRMEfsNwOZnJCvQwT1j1aCXNfdLQ0dV1z2q2RGHwfxKXVVCecM0vmhedIz9l8NS
HjkbyZYUcHdXeXUnFNnSELp7U3WE3L5qenPDnbbx+pAn2NAxxARuEA87WVJQ4DvBesfCA19rq64J
lN5pXX1QBuSjnXA6Crwm9paM3uqDWsnxbJlY4IVDNeDTflaFqDGCYtgruF9lhuQkCfV/YZJUZFC6
dK4qePPfVP4BYjat4Y8e0BugYk4VwQ/lQ4OM7T4I8YBXgLD39kwwcuvnG/kmrNLHKi+ukTq8juEj
TC1eXus6jN1iqOrOFiDPLo4QJW3AUMe3sd9Qf2H5bSuWmbS67Dgs075NWkg9fQ7YHtbvUdz/QpnA
HsgM5vMj+GxARlR/NCXIcsZtCoJmE+nL+722JmRWYeuVEpywrif5HGg9OdEiN9/TpF7uZRju+tnc
cJ+0hgYuG5S2E9mtDwzS//Q5b/VY+lYm+5Gb4bOaCfOdVsaRc762xd5kJ1fliDcN/2Fwsp04KYjM
JORdtTP3+dvBiSHwDentrp7fwVaSpZE3aIUQNCInafsvwAgI4WD3V1PaEVrJEg9ka55mFF+PcnzI
feGpNa7v+kCU0GcjKjGUJZ+kLL22TWmVJ0ugIeYWLiUGislio4oTeGq2c9ir8dphqqcwI3W5b1w7
OM9ZypDNQsIKc443KXrNJqMB5Mh149h2qqeFrnuuAhZwEj3LkUWs6pzA4i2m9UUct/Sc4YdVBFww
C6MAQe6uMAcm3R4dQ0CISpJnllcTTQJIPOR/NO1P+wV0k7ZYbE8c8e/ZpmtrZEu20pOhkz2WYHjc
dGw3uU5HC1pvx92WRSYXr+fz/AM4QYMzgeKm4tFFOVEkOm4mBChgYUiSvy8/OluZFK+cJBFKOdmZ
cF+yBaW1tL+JjFdxrwMpjVsOyBLETiI/TFZDNRSHEgIhgjGGd9aFkdwF8EwBazPN4DbpKJL3s9Br
VkeBO4e+7PPagDGIZzr+Xv2GPVQ3+mHbJa1G/ofQaXowMFExOWe9U92Ra4X629Qk17lEo0ULfnES
kfkloBe41aNLrKITg36tEkF/fqzSq8STQNodkAMD6KhH6aHU3pKajEDk4bV2XGJcVIgCfYCvEJ2t
0yqjrmPY4Uc9PgIXyrl/a+p8sEkkb00Xb9v+S7PMXqjA4wMjVvnfkRFRz9tOL6vl2zlQYWk2ZHL2
tK2CeyKgbrTWBmuQpr+rbncIxKucMnqNebrzlYAVQs7CV0arF0tzWJmO7C7Us3W7JJ2yI4lMnbT0
mR4ATC3Zn/xRcsd7ApHfRbu6dC98AXvaj8fkE5aLd++7lXxjVCGTIynL9ryhSVmGh9WVmd5Kg4gu
qzM9xrxIj+cJsizcm5NcFMN00Xj4RfjQhRaMd4IKvuqc7Bk+IfUsyVeY8tdw0MRbAvBnv/c+ojMD
K3NjzvYZEwTUbgOYNopVUAossf3uo6J/0uE0GCdEIThyaGR3xnPEr6kCUFQv6zWTf3ZiVq+bdxg1
Rv0uLx3r83wENFYaAYjyELP97rMhwbe0LsrBnVQwHWy6YRVLUKD5K3cRAooEf7r2D7BiOwFNdut4
/QPbDNU8nuxuNcjGtmlVHtiIijBCtRiXgWVqITE+pdl671qISjl5SBa6gnn5lyaUjtWU22zXeYPI
r6Tx603RP2oN3fwyWGW05URxZFKal22F9nU8NvGqjYxsGIVq/X0fvsEd4F9oMc5h11TKN4BjJFm4
1ZsyxgkoqG2hES42AOQkjfj4F0lQ6wMHs/73SRsQWjePMcdUNP7iwGfjfRCLiE4NxmVx3iiu5Qe1
tTRq266GZ4hQ+Lc9RGkMvnCV35voZmNA3lHVmy30k4nS1Hkl71Fez2ReWrFobzZdenTK+ecF+Ih9
3hfGriBTLt5YFv67MN16xGRX+0hQo9LT30nDqEeKP8LKGUDvKXZOq+18UWZ2x9Pamk/1HKMpuTeL
OjJV75n8nK7JWZ4cFR3JBx5/Djjvfn7vDpumrOfjsMZMKt/P738I3SvlVchigC9p82XiYKPnY4XH
7IuVakv49lVZVXXSH5d++y4V4JCaOlDb2qaEJL17SeDjnGQUmJDonKEceVqY4VAOoUSu+TcvfvtQ
SYFWFOudKk1SjxxhmAUV/Ebgl54akalPLoiiUiVMashkA5mq1Gp5csHprLkrS5mNGAr5ILY91pN2
G7+0FvpWM+OrSTIjpJW688LQE6sWYsh4PDsDWEEA7rNstdNrtP2etzF0Qfh/yL0ljcfi4dy9huFE
e5eHCn1egm72ZSHqBGvSBA4Fmafi8wOnuHeX8r8edKSr+8Mqha/XmALPmfH/aOgpzhiiTjtxJMnr
bRUpA+eN1g9VYw3bF+9UhLhiJB3wmjur4FL3/nGHN0/4O9c5CEvcOem3+niwrp2VoR9qa7DHv1jA
2NUvXCIQt+s/XB/F8H2HifVpfi5UGdoluXcpN0sej/mCuX8V/rY2iTQYOB46SuuHr6nrJS7Yq8y7
pPogKMBLUaiFLrjtX/lZNtudsS62kK7hpog/dgx9Xanep5p8Fc+keB2ubmP33Qj7tu/r2fcWyeSU
wg/dha9pfERRUCgZloS2BqjDOZ/tI9lABobSNjaPDx/o1xP/XH5XR5RCBkK9qTxtRzETbHmrlOuZ
FgTbpsJPMUXLOyaLqUgb5ENugaaU7wcRLPo34IA1hWmHvmdZ414rZ9qQfJFsF0elH1aGTJRA/c2g
RR2FA7Ei0Juy+PAAWZY+meo45BzIXSnWP4mcvsERr3Qe6FXd60H8pn/HP7noofMBNb+XueeS0Hqi
L4s3CcKE4i7F9PnmeyIkHeyZTcLikZHz529z+3wnJPPoJQj+mTKEXjhD4o05X+f2Q3Z/Xs96MYNt
U93rqMG+6tWcq3g5c1gOQgK5wUHrY3gKQ2z98Yt+nQ5cpX0zsJ2bTMpzpTKX54qnj3Rg+/GgqNLn
tO+SqPIiY6oVaz/oHAEIrxgyBYndezDMriwLmtRvI3j1FnS8wP+ttHB7Z2DRAmY0+PxsQ9svtkWc
C+NWXy1j2lOpGFT5k9YUPuvFkbIYYO58736XdhlMf11omncl9EZ57tEaAOB2ZKNgF2XDuf8ucDfN
SH41LO+D2d4D9KPd4TfTqfpNsZF+KnV2WnOOzjPsAH/pLajd4mhjaTogpBX76u6DHHfygdXrjp+B
wnfVmFJq2iBlJjTfJjGlosI/B9UEoIQO6V2a0upN25Jrxr/N/2ywAmXqZdrZN32w8ER7UNVRc7ze
sPhRaQny33ba7IT+xXjVB1Uc6d7W36v69GVhZDIbfdecKB47zEclWbUIVHIN1Rg6UlfzpRx5L96J
nTKx5xjt4Si7skzl9NPZ6/E3DcHTK65SX2hIPBeAr8txgaIQkPW4VJqBTx4JVLvPgRUM1bS18gWe
+57t8HEqll6nb5n7vzcEn2qX+a48t217QVifl6hUDwo0RhmEkyJfm4V5DaoXnilKxq9DIKWVLxt7
4nMs3iUqWpqp4XKi/lIiFCtZJnPFqhPcCTEs5vdi/igGfwmZhtgPLjkhp/rG96wmt0jZ5qauT6co
l2ksNAXMlttEGtfL+9GHOhSD1TvHpCwyAhau1yBNNf3yEy/zsTvGjhiqNmR0vdadm80GmaUvfNTG
LNgyWqKmg9D+eSCYZhO7ukC31EAN2AsTOGhUgmQJJU9y2KGfF2ZAoSoP6FR4RkXzb0vUkoNcM7RV
Wi07nhApNnKNjLiNiqo4bstQTGhBMTmZ/0fd9YCciZHaARTSwKGUIRMUtneq58uYUN8+fkGZtV1v
vEc1H3ORJ/zW/9rDtoOPtfAZvbVlUQEFuVCP51Tvk+rVu/lmeT0ow8QBJJ3Pdmjd9es9DQoKwO9W
yfNx+JCdqQ1F7nAHp6zsMUCDHDabKzWliyaC1yaEk7op0cy6hgBaIg6epNz6SX1326wC2HGT2DMK
brmKxntKmxcuJ1lhis4A3KmRIqrziFbLkyNLU8AoXbS85E+kFQBQp9frPA8l/KQ0obysMz0h2iEN
24ywnZ4jWhCGHx899RXIMghnjwhCmoU4zYo+0pzAWmqHi/kAWNZTtIL90bbJDB0X9YyZ6jjXnApB
0vNgAnNY2Put+KbOWFY3vRMvBpdFoD40m1yam4lszVSoSY9CJqZ4/+w1iwSJjfTCRFOkZtVD0khJ
hHdpMVskXxHVsoBA9r81ln3Gs5GEGwKKFeYJVMTNPppsxdNDAvnyiymgGDLj1zAsTwDrHORl6iqC
38snVeRADHn7ZSlPwKkkNBl1ae35G1PYXeeeze9QO/Nd59LhvIjA9VXz5XHuZcAtwB7untJ7j3cH
PV9K1wIxZ+U/Fxd39pxPr8uih0ZYkKmP0cKGKP0fTkjrNlkdRM5gqH1x5nZkWuu4tTzn2zlICgXm
qQAcPbfJdQOzoIGtOPm4ouUMv6oNsWEep5bCboQsB28BOoer9wyp8HREQLDnfNk/w8Dds97efuKe
aExpnmBniSARA7UPpWVKyxzaFoeVT5czK+7B4XPZx7wD615/DU9BVW3sNYDoOrkHyPf6vK84+hta
PRmvhA1x4QBbTVsPG70LMbL1WgVWdKuwTvtQQsdQoj7RMXt21gpLXMsCYNv2hjWN0UVHNoQNYtHR
xTqeDykH4+BIKGBiQRuRTAqIP/5Gpmwxpkmc5Xw80Eu14IjpEBTBJfpcGe5FmE4uqJV3QuLDpW0+
oYRdd840RILMWSEzOuEpd1g9vIuXVMw42IzaI6p0oE6QjW64930iaVHmAsn55RvxId/agLM5EZd0
Dfkp0PbBQQ/1ZhoOm8Utn5FHflc4rXmpcun1aQiLqietC/biCQTalpHaGmWlPfIWRSNdxj7jbs5h
PiWUpMReEZs9axgFPw1lfuA4lBpahrTKIVhWqN7+Ht89Qh/YABknqi2Ue4qZ+32dCy60eDaH5C0y
yyTBWBJWFtsChQ9juDweHIm96DLEbtAAoXTJwwpte0zDQX7Wd0ORdvgExFynB2adOhMhXWzihNmq
G4xb8+RaqudoYDkCKLt5Z0fVij3G3WFysaOGDOXvy339YpuhQcwAhYcB0JCeSSO8u0po6Yc9j4D2
xXfdXx4jI76CYT34htOuHpWRavdZmg8RwLTRkhXHzH/Pc5NRakuGvUcWn6Za+VXk2TNPYprVACwa
9D5mK335+riinqEZHlG/dPFRvty2SJp0+oBGYUx3V3baKaLHoqKUDPz5ALlcoEjHyqJpRRqkNifk
k8jTCaTbuvotXrGOU2qINOvEsbQ09gTnQkjeQH82JADYbYUiO8BoPoSiUJcOdw8taOYlyD9M+SbV
xYC8aF/6fRrxEPQpgdvAabsm3IXHJXfSjEmGkO0KLUOanq+Ca5hYSCxcfxPWk1XG+nfAfdwlbPrN
Ut0JjWHZH1X5y+msfDE+FwPVg/pkX5qF8WRomuVWCbjmMtIHg3Jer4QpIofQq+ro4Mal8lUKUWBG
bvqw4wtXX0qaF7Bkt4GqhUFPwoHrzn+Xs99hnv8iI0zykQVuMuR2lOw0pKNXggZi/EPHI1xzpEf9
8iJ/1Awt6AkBP3eVlbKh31/Lv98PgDa3un8+GjFnDevkGs3h+X20KC1MHqlZ6M+1EDTo1HtEIl78
9FCNs0AoLjqSmtlMPfXlkJz36JccRl+QUNXzGHtzWH9fEVcHmkc1raeYYg7DOOzqE9r47N9ssxqB
C3Td0LvI2LfU5d50wNDPsF34NxTuuNstg5nO+B0uz8VDy7Yls/HJUZwGiO6W2YfxCDhG1wsU3PBz
mPn/edh08NMVBR7PzAMml/A317Cf8jhi4mQ+4q/PL8AI/pfT5YKioOxW3nfsRhyccP+1xiSsaFVw
iRaSac7W0MB6MAifGNvqCBkw7Eg4tU0tk9+O1URfZM7KBlYS3BBbNZ/2c4auzRi+JJQXXVtz1wPh
TRtl3eOQgZaEKPUjUaPfv74MdofDDZv2MMRNun1Xpw6nZ7lXBIMa/N4iyavUPASq7TV+rYuzJAUW
uzqZZTz6wt8+0L7dzpeeSAYW0cQ1HUf8opxvsRL9M0GB8psWgmKzTWu4jZtzvU9JvAX0NMUKlamJ
ahPfpbtRKoQ5p3TL6Kah7gd4R4NTtVAAf1g40rRTY1UFQsfKoG26mkZ1JB/vPDyVDn49nGMxJW/3
v2R7uWO5PTlp21PeGekYEltrRq7uEVY4wEfp6LOhAaXTdwRgYcQDzF5m+JtviFLBMq3p7hLDQFQU
vPCinE/vsMVVyWocj6B34oVELdyqZDYzxdWObgMpXscLTU1lHNjY+y/BJV2XmX+Cre0ZiZ8rEsIt
SBCJ1afTaLUTlFE/c/pPuU9edIOrpv313Z7kxLKIat/eIme6TXwgeerKRL8NZ2qEj8ltva9vsPsU
l1bb423dodgntJftMaWXGzGFdLdbWTktSSXiSL/vcsIueruX3wrXasPfEwCgr71l0HOsgnWFdp2b
NxytUs7h3xUy9lDtLTJiXavW7VZvb89sunisJ+WqQw56lu/PJ+TK4CZy1p3w+U3jtBRjlnTfpMcJ
pXOzwR+W+36mUoZkMNNC4KHtLYhFz06pNgEmVV1BvfNEJAKEpmKCAGvBU0EDTw5hyprhNa+YeDnS
vN3iSOT9rQgkHkwiisCmOlJuhGcWRrBUry6aj96b6ZjjgVRI3tPhMlublARUg/KAPhXTDq1+IlXP
q1hvEeB1UeiRWmshMqnAW+3J6mGzr9h1vUXh1J/x6haf5KWJVo+CoEFxmtjGwoyCxee+g0pLp2/O
VwC/C03MX4e2HgZ0+Am6P1+mGVsxWXQ7LOiYknHpB56fkm0M33mBGW6+frwo/sWDvULFgLj2b5my
k3LWJ4VjOjLIePrU/H1VTui9Izdv+1ebyupPLZr45TFCB710EDXg9Ta0vnd7+6CL+VlOoaDp4kUp
Nzk44L5eZccdz1cktvsVrCBiFNh+9Sxq59ynbyXc9278L8X8yorp2KRuNcl9WUIS2oiKVSEQX1vx
KzOhnGooVerdt9nC7y7onXtXXJX6Eq4KIDfqIHE3yt87IHVfM0z4YNgRwUPo99iaRWOlR/BiIm03
qsT7RhiXvL4OZnBGMOu2wWNTWNYwChKnpAmg63OeB1yByQfHZ5vAn6goJUHZoCVB0nCfKRA0OLlK
Wc7bGEcC971PqC/do5g+MqH3nqeV9kHKfNCHe1SnJ2/6lc3Ket8DcuQXeWshs8QIYC3ZUeoL+xsF
y9U3PR2fVLAEYDdg4IpVvl/OGHRwWw8b9J3DuBuAX9pKbpI1+3SupzqFIdwuZV1abzkv3SBIQZNM
rvstpyq74j8+IYC208IX1ie3y7K+wJkFzLeSa4Y8tWQv45dlJp/oMJIvhc1n8n7AdURNMTHC8ouY
pt2LFByQYNRFsnfU9M4ohvnc0X9D9fzkpw8H6nc+gO45mKMKPhoeeQGqPYN6XhJ/eD93NPaFTkED
p/guMTmOuN522MTEJWUT4hH+peBTropTNk2zIuNUHOqwlBGR3LLVJRF4/eDy4co/33ynpYpD0TcQ
aWoLIopkPOweC+KHxIti8Vjc8Qd3otnKOrOOz0wfVqwlRyGXFqRD9+0zUQxVukMJTRrBcpoHncU/
2XqPoAYG4ydotKAZIfu6OOkvzBU3wf/Ehus35WvNuOpAqZElAFzJ1j1tCrrzybgwABczZ9mOq/dv
6sCmj7JgTh8cZyteUJ4o7UFFSAOz5kJCZGrk63GkftUgBzY10ZxNsdFxRm8ht0GKCnXrwqnEfBeY
SQy710EvmqSbXxP0aDTRtIz0worOehY5HK6hhNy9zr9ZEKVP9RpdPsWBRQV2guAkOBb9ur+VZ67W
OtDf2KcqVTNHeK1VeevcKOgYVbR4+7cT3ZXWAexVZn05Trn2Qsc1+j3AK324GqN3JmA+T/Z4pkTi
Ka7IS/I7yBqloaJLVwP1uUJCaQHoOvQ54yTsA9oseNcCOcoDxIua4wq7orzgHRzRB29Ifg/uK3JV
GRra+B4Ak4KOWIEbcicNvidzCPP/iNMb0/fynKiew64M1sk9SyBgsaAgxicH0Lnq98iSfm3mJLQf
FUDuL0Q5WZX5LYTrgW4rMTZjlp/z7uWut34nwhRfF7mzCubvutBthfCVVQoNchnpWJYmYobdRm42
3zbBNhrp1cDhbS0KBGeoQOmhFULvWiFso9jKSVVt17LXLIWRktdr17JJjzWhj4QSCjualMLIGw6s
MVagM97gyDRoRVo032Fr3/VqMs07JNQ9D7rtbK+aka5jVfeSIyS09BLvT7LHgbA6MKk/GvghOZvh
obxocBWZSuiVx3PEP5oJzc9wqTqT2tadpS+BClwwhj+Y15aN3+fCOanP62xgkw2DmifBL+v8i92V
+x+6TnNXW5gPjHpr2es+NmtHDw2+CCXeLOs4lNM5xNC1RtR7r+NASpNX60GrMrpn2Z0DPoM3SSpp
mP+LiAVLxj0MoaKPI3F1NXSSEIjGkzpJUOmDsHxai4OxSqOkQZsH4pFdoaezht/R20B7MYhMBYhz
HRF3tJa/9vjyXeAVm5Zq5vLnN2wf8MxS5mlRjuyP5F/TqBUznF5wVJtSf3VDMOyV3bfLvRVEAd98
cp/seWOx8D0RD4ikJoTO1ACr+wXv79lL1PyKYuHVuwe4byUBH/V8HXUp0nxxGi3Cyd0xDtLmsP/9
uTcSQPD+ds5r4Y6OWVk/aVHTVNXzIfXCTxhjmmr4EWGm2JDBDtcsRg9Lddsra4ouSIF7dztdpfXJ
gIInjd7b6qhM/b+bNDFJfQ2D/RKPayXluZ5WYC0SMCHt9QNyV5saABnaKfyu/TUGLFCvRmjRN6pR
nQSyHx5ROMh5FBdSzm/rMRkpNy+wr5wubCaQtu8LzRSHUtKPWrO/j3Jxob8zrPg7uzNjk4jsYwNi
Yd8qjkoLsuNDe3WTbKJjfM7ytIFecZkSvb4zDRMHLLl+14iAwki6LU19dyL+CnTFeAxAr+W+u6kU
XgB/h4sHwyndlNSmQ4bqk5pX0yP78jCYr0gSis4yCTfgqAHmMXi2SfixF+NZ2EicEDKoifJTGvR8
nacdHEZ3twn/+8AyglB0HakxYRlUPMoxrVOr7KruRJiCVQcZ9MWOiKD4qoyodGHrUm6QsGhBCp5c
1OexYRELPJaPJaT3WCkIRYse9eGXdQghGDafJPQkpxDy75WK0iYwWArUIAbTyKVFvg8yAc+cQbj5
2o9iiF/NRGkqGy/5SPL9QsJOaKnpCrw8gQxIXh4zKqoXHFX0XUb8XHmNnnQDYzOq3NoFKLK0XvnJ
xFPlJGjgBkD2Derev5apN1apltsLosq1aSz3QSBHqkGdgBtVGMW8Ft5iPLq4K5hvNDNchlUKxy3D
bhxzwdPstg3SV1HXeYawNNDpS1VJOZbwTQRCVJPIFzQMo1qu6OGK/XjjBOZTRO5VFGKeQGso7EQI
ICKzpHNclv4oqC+uyQwYB/52PdzHN0Zhd9u8H4t0PrJdPlkky5oh13ZwfU8jSabP4+79eqoUWKqd
+XZCPkS5tZhqLXQi4RQKqorLAJ3rXshAqGItcB0cY26K2FpxSVfsyd8Kxr8mVzthKB5XQnwskm5V
4XAaoRb1cYXH8xQ6KXsX6RHJvRrWMXOwzh3ptUDm8Ue1ganjRVDcH+wYdlpD3P+gbf774Rf8kiAJ
wiKROycNDV9tdNq2zHDZmiLCpjYHJC3DUwXKCErII5/9h6TfE4jSmytFDcQ93XXBopyvUWU6NTyK
PXCQdMmwR4MpjaaJ5g5v0GsA7Anr7t54PPD885lI0BqGwC7NwXOEbMQG8182F/+/Q6KrZQ7Kyjbf
nHT/QsrfMGjrZPFqU8JEqC2C2y0GMY3/3BYZg4vh9t0mLLtGHhXuG2/5icDrkSdwM44kps8Q9ufF
KVnjp7ajR78XNG1g1LF6d4u7Nexkl+xJpXfnwBRHMoiAkr/pYYredEYZZpQrpaF9UNiZdO5GOIKV
lnwFjCnwHPxLrfSQVWcWRiKjEdqIkf9J+gTMwheKhOaq6qc9+7nUlkMLwV3rQl7STshjaJWzuaGu
tMwEojfpOhmmp1M29is0lw4q4VVYrwJSLTZM/p91nJ0UlaJJ60BybXs8wKwLAISazqxTssr08fkZ
7/tk1WuIOv5y+8savoz3eaIi4+yiVaQJhJQhukqn3JaWmTps1R7+Sdz90Sh1dtS8irQQPM4hruME
i1VcuC5zO2WUyQqtezU7UpWH1qE3G4InjnlomkkXlXleI3g5cH0Yu4dOHFEuoPwd8vgwfiGiFO9P
sSWqvOazwp4HLWaA5mZdR9yz6t7VaLVDhypMDg48To0JWObBctw1/Gjx2uGGBqVhSK/8FFG9Dc4k
2q1/0BLZ9rObQukbsNKmufHf9aftR9xLDlFk+PCrb0CSf3JHXB1kk6lwhRBS4aataqUZP2PilzAS
sCsu7TdXU5+hU5Hqe8VAzdRyAPj7WWMrkgBz+n0jP9rqNYPSCfhkV6ee1ibYGniJ9uSTd3WqlJH5
LrcCHBMJSLFf5oqfrLrvXB7xL+OYZyntnNVaDielbft3yq88jKdzlAspAPFtmgZzL5kdRTH92zHS
5mDTq93xhQpjVSVzYyEYZgtLjn07pcf9bcQ+0NEoHqM4pw+mqzuK/HkCQ0Nf02em2yUFQzAgyuy0
KkmdOOrVD8V5SnVJjegVGxF1u3GDrZV7/79ofWEdD53uWu76oQUa7z6eCbhkaFop5PEDkXf67JzT
89DlBl1Yd1CFqw52bW5KGape6B3vj3Bic0kWUWd7lQ59xKzfK1dG4i+VT3NsFzgQnsxWpNpUHWEW
jcTn6dhGaF0riG8RKBaAgzuc/Q/mN7LsPtnXVNJ01U87bCT5MxRECWTRzpa2+ZRTbtAs48y67rcA
Xhk/Vg6nKVz6xwMPSqfT2NZv4sozKGGpWNR2j1n64/RuKQvrRqwacuMXn5l6/m4rPIgSQNMgAs31
IQhlQuksJy/m3iMlpBWQETLLcjz0A37MdzuJ7AnZdZZZ+5BkWrvSe9BIjSWhl8J0tFuo2nQdh5MN
+lQG4v+UzFheMyEb6kVdT6rUS4Ivc3t3p4Sr37jCwWSI2vLx9zsIj9XiEIlPsXetU872lcnAo9+/
PyvQ+vFw2mY5T3ALi38HmSYJ1V+Y6wPWJrApxfr7XyG7IXm1zAxW9C8o0lRAZS/6xxOvAR7z2pEW
GKdJGHVWoKgZfiuXlzR7AgTmg+6tCaSU450HYQWMwqruvzB5iuafSECqfx83jb3lrISeB9akA2j5
t2wGbzcdHzSWR+/5RcqmgIN9ZVHh6r1KrlrL6Ew3UITJakYG6RltihLQxD9o4BM9tn6eIBT7yNQk
K9v/K4d0ZCHacPjJXm9mMODkSfERTB9dg1HdS/TmDVxZiEnSxUwoOjun7cpDOzbeEu8jTkPBOG5p
Q/fPzPaCvxlWkeu0LE7zf1ic1/wUFwsOCUNKGFzahUUafUCEIeXpA9hVlsHgpUgUsIjoQVMgIDs0
hSWJl4Ejx6BorgoBAfOK0FteIub4BIqE49hiElJqjnLMR/f0+CWTQD8ZI73tfGZofSeg/hWBBT1Q
OHeY2iRdF9Fx4MLFZlmdXyPenASHhaAB1HZe5mmhd0svNjdlszc4gQDb6duvHtX3aRY5biSPkREs
PW1mH77bGtU4Uoou+k35lcnrIFcrYdgLE8JEYspPE0jfADEJs3bfNOezQ/eK4aGpdw2nLbkP4HzW
z0H9FzzziyC6j7vRZPWLrBoZJvjwYZR9Q3QiuOMasxuf/+x+eCqlfEWPjBcfbilQoJsprH8IgsvU
a6t6AJzTbjt7Iysoy1sbfPGMNHLyDeeFVlN2Xoij6N1t4htZv3qJFblyM77Uj9k3MhuCn2zeJR1R
09V4hMaEXnjAkZPRj2ftL5PfEiu8B8xOu4AVb7tyNiOxyctDRI2gyj7nxzKNprJCD1j8FoSf1E/s
lYxyRD6U0JfPdkjJqioLT50LwggWVQDIZIVbvX1tfEHAjLI+avf3ASMXE8+Oq3R+NTWyVkAHLJBx
wnSYxotJbHNSykhZs83xmIXYaA+ZuoEi9bOmZxI8vZMhuqzhswcPIOscXcyUKJO7RpdLEGM7npQQ
gYHIo5ydPkkrh/lSKPmiY5eVidvP6PhAfEBXdXKf/WMzIaIlAwWUyhM7c4GnSovUmrGQzZuBGc5m
AX3rWuYuAyD5fuGUworp//5p42AuV1wfSF+pOzlBl4ecf4iBG/He1UG4/Mm4YlhyypjyP38W5RsG
9jLcO8alN/OCYu/kpSX4YxtaDYUfiPfXpwouuEqF7moJqnBx2P9KQnSU5T6czsd1tFocCTiqxf/n
I5/a/1VLtt0jAd3rx25WDn4Sogy/rTex7l5PRKXa+2i4/xZR3xFr74p0dMaD0VzwMsN5Mf9eGGF+
VgK67WsHpyaKEv9R/FrUvp7e2ghiO9ENyHjBI5DYJaAxfmYWv+3q0Yn+m4M80nySBFW/vCsiri9W
Jr8S/5LIKiqW9oJPzTjSE2kMnqtYmeCYZ7V/vXbEfuxrv1+QAd+VsdzQ0ZmiRkul5XcGNt6SFR9R
GKFP63HmTVBfqv5I7gGLAhNj6+aAtRh4pJHFU+jNnMxZ9pbU4tO1Zu9LdoVOTW0mFuweoYMOIJJd
AYG75WP2ny0A6HXewGhQFx49XighfRiEzBJigGfjj5k0nDj/dPkurcy/vN82ZUnQAkxHmvlqIAHg
BllMq1Tc+KGF4mNlNLAkA5tbtJtewGDeBalYMf2mZUb4Z6KMBSWKfNHLloaSw9SpqMMtxxSXbQry
45UupidwQIgMTqCUiNKVK8U67Sd7VBpC4pRLi17yz/pTYraQ5WPVuc2IlOMqJnaQsXwsokFCz2RP
o1+7UAzIxDdBkx/W1rBAV4tQi0OsGHAQopiSQgHk0aGBjiGtuEQ2URSFptEqUS71vSWp+1UaDQMf
M0cQb61VT4FOt7heOcr4zH8vgLtziKVJjL9hDCu2ZFicB/PxOcrHz+aTdu9iWH662vpGtfMeprbk
KfGF0VW991ZWO/LZoEFYW3ekZmf0D2uzjf96yIiPHWAl1bulOjGhAMuND8i385s2O/Gp3CMkPlUR
0YUG16U0tnsTVmAfZ1KbQbFnJuRUCV6OcddPxQwAaWAQN0L9WlbLPobZAD+cpqZKo+I1L9nxQ6nZ
mITcpj/6CREJY/dB1XCY9/ZAb4J22lTURxBDw3m71VD9FJuzST9o01JnBJeK9xRL0wSQDoF3G0wL
5fUygCbgQDH3xX0Mn1o97ik31PSXo7eT3Oo5MGc3R2J872Nqq6UwKbEbm7hCmD0K9BsuMMdZApW9
Qc0r21S/Us8l9zH49k+xBQKI9m8GwfTJZ1P62h3z63D2ac9sCdBlKINAaUqZnXO9sP8rsD3/U5xP
jKX1krJaEEcvIPveu++uWvo06EekUossfMwwC3nqZrI41wJUwOpITjauSWDviaXi7/9Ag64FLdlM
GiXnwNB+zv54mZRDCq8c+tNKSXfhIRBKK5frH7U0MGygHuNs3jr7fHzPbwDBVOAH1Bw6yJW98cje
KsrtMDOKNAV8N3euVQeA+0u0d94Kt5HF4d4S2zCrVFpfmOC6kAFKNO4PeHUxHSgT0Q5/ZebhqGGd
45xhychKjUcb5aPFbkDDKgsopdDWzRhvDiStYlrzr1rJREHxiJpGCixY8kksWnX4pH4VE4n20npd
7us2++DCh8Z0iYe6In6MfJheINRyN04H3r7tf11t9EtjL/dmgf0Q8apA9LmYhondcska/w4MxiJD
7R6G6011CaLZ7Yo2YiDn1qArpKB0BKMHzEHIp+lQwxRF2rF6qQC1qkEhcM96aEH+tfqzlKNuOaVS
4ptVG73k1Ltt4M6bIDUs0xcfvQp/YT72UqA4uXgxz1KA8tL/R+4cRDg2/2CQQgRzkge/WZE56QL7
F4UG9fjeub0QrPM0fkr6U9I7iQtAoK8mS1wi+fsAKpYom1zQHlwVWpelPsVLN0+8C3r+dKa9Hb3L
dvsIwLC8j3oSaBmbN1vf5a9XnuiPcJsR17l7fOpTD9YJbf7WHmq5hk4EupSmiY7BY7wGnxTzI4BH
J9MkNtQPZCW2UavP9mtuz+n0s31rn2TqO2te3LErp7hxzRwjs3j0LNyzh5WX/i99omvE8mrahZig
kCphNLd+OKkPgP9QXUkZlCaLCwS2Sd6AG2z9QNo/DXTcdMvLfFCGAsZxyL6Hm4tUD2Qpcz4TImw/
w0GScvTN15yFU4fee+kWs9scHw2V549wwqIhwL+VFDQjd/5/VitJifmSvmVyT7HFyhPu79vKkD9u
mKJVCOI451W4B1UfaRDUY2/pm2g8yGsEEgOEfbrELgpqfcHltn0ANOY+hlHtVY37bkdi48SCY/Uc
qk4sWbvfhDnfsLUUOhFnReYroOMKZyQB1cY+S5iu4wG91clx+XTRRqvyXjnDP+F7wU5lBJYXRVj/
J9AMMVZAahWWBx89Ev7jODyHpZvpx8avQ3l9RMQT2FiH40c0G1B40rfixiH2ikUkF0cNKnrNTJXK
7M8EZEeP1thDixb5znMIPrjSfV5JlXaqZE4OvmqZ4CaWECm9brFIMLnpacw8XFoX+RyiN+jwwoJm
0pjicrBwvmu+LOsfWrWoa6VRmulloYLzIvDemsG3OGeVbMhxLf4DYJJm0v9U+eESAOiU2JmPSg7r
x2N71Z00OEqKYoSQGzyw/xNiXoQJFdJDe+ahsYTyqjrhawC/stbvV73cx/WL3eXkmW+0xLtpUjL1
mYTBfPxBDuqQD0cDSJUFdJsaE/+X00rU5Sg51efL+3uiiy1ncqETVJM9fBet8ZDd5C+L0YOf8OqD
e1cf1nmMTKvgdoHh5XP7bOArSQcmwN4vV7CaN+M03GfavI//NcPRz6w7FHub1k8eknfE9GnlI+Aw
nvqF/lNfKuYYf8NJeeX43tsD6PB8dviRHktpHBg2qWOEf0txFwA3hhhnWtox7PxVgjrXwVYkwnOv
ignkv+QlBSFmtvz4wBdVzAjpUYvignQo+2LIun1/lbsxdgun1+uZ2A/GhkeSGq4KeD+9h5gHsy+n
ITBkx/6rHqOu3AOMVI9cy3Fwer2FcJcoCPUaINgS4ncNEAw5IVwSCkox0EAqEatGdRTGJPsYrjs8
zed/wDBr71tzrpL4dOyl27CW4dpnNRp/YRNo6MuGw1QgE3lmX6CSbzERiPmHwSNThWjvvPFAep5t
IwtrcMUgBCcC1cpPLwSb/1v3hju4faw0OJzlrOG5UJAYoptQRN3sb2uW5XmKmbzCQiZ+ZolhwNiL
oBnyzz24PQoV/LmCxK6inPGdqa+248l6wLluqSnuMd8FIvx962lkDOY5X18gKXLm3LsMyAQoxo91
cloYjDrn3cvRBzyIb37Kdh6+rH95HejSLIiqAw2iCZQfllht2ObqVoenqeZHcHt8lTFBLVCe21oH
SZlIpE3d4/YMqrxTBdQdnUG4Cmc4VRTm6IL1/08SkgrSHbWVIIfODR+QmlhzJe+uLZZWGNlGKOyX
OBYoJN/1yrFJWdrbEMIAOvkeNODSUbMcmrvIjzIQ9gxPVWhZsHDwPmD8jEoc2x4vzFQO+3Nfzgwn
HwFZYs/1xOsuPW98zGAm1OwXr4BqNO/SP9lY1LiRtU09NgR72d8WR5P73puEg1gTW+HyIO9D6GNL
pKpX+ISoubbjwyo6cPp4EuUD63wc0pSb91Mob1J4xuLunYXk6vikkcEZYlZmIe6yHX6qTIln7Veq
st4onukvYCmvAUJdI5GDewo1zUGOWoomRAdd5v+LMEIXmOeogLQywUnRp5bM55T/n2KAZoYoIji/
ifm9tbYW6uAEY+MDcHDDdwy1eDLEjMRBVWEgk/uQc8krQ7goxZcjsK6vyedPt6BEMNPKtJl2CdiD
EH4gucwapHRPOK6tiim79Hz1qcpNYeXg6lEwUGGWNlAAaE+Ab4BD1fNiP7JbY/rCReE2RK7FCjH5
jWzDhhcvSkmXTyWcs7923nlg4oqITOHgDJTnUEHoOEGvJC5Nr+RFRDAjRe4VTTwYjtm5d1cSBzML
sNpNkOe9wh2zNbYBlbKQtznRFjoBNmsOuw5vwnCC2OA5JZFREbsXLc8hIhvEN+tMTULxU8prK97M
1IjEIPpaF3QDI5j2RPPD27WGf4iB9nbdCHU9vtgPmJ9f5crgoSQtmmW24N1hJU1nBAImHc0BsM0O
1ZAXJB0fLEXaPa9iQF0JfcLTZn2y29g9u4qGUBbcT4AJwaA4QnxLsTP0ECKFUDaDbfqtAPaqe5u4
2ZM3byKawoU5Xpz5Jch8st5L9xqLtdCVViVxyeCiuzkeejao51/ZrGBg3I7tHeUG+2/94lWWkVPF
8xanC45Fa7TNmhdCOaa3qTgc2xBNYKORXJwKKWTNuo3ZzKBUEBQh9KQagF7dsg8jZk1dgVnxtszM
emLJ33Jq84g9JLWhE5AXUfg8SPQOBH03b0RlClWo+k3hIDq4Bm6YNAxpcCIW7RE6QaB5aKHlWy88
1PY5G7oZgHPRHBqL7FfiVhauWJspoFxQ2LctSZmvPDVjiejTnGtc3RL53vKkp/WWPtjN0eiycojz
GrIGdzO+F+YA0nJJ3jpjbDlLHcj0UNbiV+82b5SF7AcFcPMBMB4vJMCsIVuKNfGNVbX3HM+M9CjO
+4en5f5Ddmj9LRFxWyi0VYQMBbUzl4ClGBX9HlyFpcmDORw5hiNo67CUjfg5y/7yyYUBRWmxgXuj
GI+gaCdF4kHCbIxyuGemSq3lq13twSc8wuSMPnjteD9e2ZeKBx1ptcg2nAhuLGADRTSmW0PVU1ON
/Yme8LsZeBX1U7oYRp5X5p97r7KMYqyVOGtEPHUrMf9fW3P41glo+zfeBTBl0S1xhufFfmj5ipgL
2KfNS14aaFjeEpbzvHW2YMHWnr5MmdleIYS1Hm6osvV82ENe1pRfvtpDjEwj7EZ52xTZV0A9xyKL
SsEqErhaINcc0jXneUjHw/9a4dcL7kZGL+D5XsvQLGv5mBpmqlroLeor/T0coLjicpRWRnK9z2vX
nzIh3Z/iBcr/OhYqP9ia2snIpPwcStY/c7ANMBehjthUflBaStvaCcYNvefO7F3IwyJo9uabuHS+
N5mZOBkA1331SFTWp774K8qP9vxK11AMRYlla3JCDeTo3hX+qtVIwPE7o6eJ9oNuyamDakYNWKSZ
hervFQg0pxqQTBt+VguuUP/fKmsVg+PSVFTDf4rjiNtiW+4pEHttlqB8qnOb1wv9t8lS8PDSLaK+
ZbzebYtbKxp57eaJhFcd//aJXprssGzsnTk3Pcsi1ysZkKXIxIi4eXrzDkpto7WwvBoTeomRo6Tz
a4H9yxDNsT2kEV2/+11HX/ayB21BChMf+eea0bjs41K1lfxFNZnqbi6DJI4Ux5GZOc+O45HIPsxe
nCKqdGB5AK2zOWcLKKX6PhJkCvAdqKPN0V8LDOO3JwAwTxfgp0dvn6k8L92VYXcGXiVMDovcQhqM
RVAZI1MfKiLH1WCiIP6QGlOJuDp+HgQbjc5tBaJYpGAZmuf7z/edReZ50tnNrIHocwQfS0LLRU5r
fVBA2xzNFymM3MvcuW7zb6bEX770QJWtpEWp0RTNd9Qu4ND934ltOY0UY2w5Kc9vth9+6fQk2lR8
s38lN7G/LbH9KW9jF+aExRANYWfYzuCYAbQ4/CoUKu09GkXgcr04yJw6alq0SjTCt7z2Y6rITd/Y
pp0BsaXt9HQBykGOeRGjyd+cknkSxN/JQdMB1WABLdEpouqRCWHCpEfRzlanqeH4bPdvjtXN/XW0
aezoOTEJI37PsJ10kUoVyJ+BhbSsUfqbuBqkWWkij3OqqG6bpkq45Ifo4sIHZe/cRYI2lTleun8h
PBEhEOVkk/q10DZMblxlNqbfmU9ECveOyrPLZ6PEZCvQ9xY7Ao7rGd6Xxygb5uG+FXp3USJDzu13
NFCUs49Un9v+O6ZuJ6SPRRo+DhbFDEKveTpe+0ajzRTp63Ts8kZuJCaNa6jJ3Fxaw9m0G3bI8jAS
GMdtSAJskson3smo/bVuD5GkTDjHGE8WZ+oogWWyMBi+bxosz52UhLr3C0RNGKBAcF5C93Ie/zeJ
r7b9IOg+S8xVF+9KJqd3VgHzLPkKH6xvNlwTZFh++GnX1/y1cuiCIByaznw4zHOOt0teVC3VS4iw
xcvDgjBcKAHSCNVv1uWVXZADXkApuAUeEfOqKl8a3KsGE9B9mup3LuTqEzBsd/HC/CK/HXVtdzRH
pDiQhk9StjGPVGvktJAm2qo7H/0/DMk1PPANKdEj2FWXQRQ0oLNTY7YMjygFdeXbcEm0C8aYPT32
DAdDiXVzwX3FcRqhPX3Z6ucVREXliW487307VdUfKQj3q//tha/nKxhvjOLgHZULcN1CtNntAyAz
sz+9GDc/njGo9fZch70Z/+uX6j9zwckRJ38NwLuGFBymYceoBzjxPQxiM/ub0c/tPmUP+xibpjye
649UUQ83QbPIELornViw6k1//7EqKxcd/kjAOE0nVtx11lno2M7GSkVP9/Xjdkyu9/+6hnmjHzLr
EZifK7AnfNUNoFTHNRmTvLSpmSyOHD6gg1MiO1+ijelnA1pRStB1UMgsoPoqJmL6bAkKOV3dSiU0
vHr+MsZze1xTia9gbCAadt0Q8q4+gqO7vADaoz4MJc083/KZMxGq3pisWvXtqGP9rINndsXdwXU6
H1V/373gZAHoGGrjhnsejWEXP+G9waxJ4PynduQ7xsKaDL7yCfACUnuqRU7yHApzEHSqh5IdG3R8
4kF14eEkPymTh0TqZA+l3C0OHA4ikgymaNVzu4/s6KagfukEYwvUkL1DDFtxMx/vumgFsEunlM13
R3prQflZ+Ww0xPm2o9TuFS0v7p5HsxJYWpPZ2sTaVWPYGdd9L2hFfrQIl1mN95ogR90dgWCjCIAc
5bj9kAORcjZjva37BoUBAtvEKkfm6OJfDJP81Tn3Huy8MFpsfko5+tozfiv6M+fb9YvshC7486Bq
E4DQA2yWTDPc/sbkB3dYRIRNrgSoYL2dWsbBry292E5joszMYdmVuGIhzc8M+I9dTL+cwV3O+SPz
joGpe+zUL8ZXE4hAfL1N0nojknhskR8405VH0dv5oXsXsHH3TKpOYk823dDQD9imcm/Xq4aZ8zf5
dqEYQpu4Ey9TtS6W6NcLGLVYQKM+vnjdvUjgTsvHY3CBAIjhxFM1i2yXUAYNVX/lpzmq9IkXjT8O
fmjN9bn/GiX7SqzfWpP4dfzS14iuZke/u1hkEGw3pjkSaOV1rHMit6Q2+JqNiw5JjGtUsTY+LIcL
c9U+J/KFgoJNd6XBg+1u7mwpFGq+97I6o4QQ6T+dpaEwyYfXuc5geFasPlhZpTSnByxXT8gVUFn/
8bGWke6aGB6dwRPLBxMdWVWYigWGFuQEmchmEfw1j3dlLfHFQBas3E/otNZs5aTSSKxncIL8JaUr
P0jSNranypcvt7/Byea8VXhu/vM0c10pQLLfNUrZNqRj+alegxwGQ0IBe59WETfhHuheMhNeNNjh
YDeRaIOkVAs0VR4aEWzA7Tfxo06mN7fyNeid3bad8QoQbKSD1y8HYaAES0/HC+cE7PzgkiT+BKpL
VeVOzxcfdGuMpZ7yPNAqA0P2WAna99Ej2kYyYsBpcqcWFL5FgU3MWtD8shdwQlm9seoyRhrx76Nh
JgH20/QS+wP7HB6akPR1pCmzHvZv5fuorvHYqexMU/ZwdPR5srdpk7Axh8tIn/CrA/bpc5epOwOD
xSNEnd0/dkYcs0INb4tX1VVqlg6ybpObKjqBGtnm2qxgud9DktNvsSjHPO/1ntfNhU6z6Ls+sFsp
fFs4/U8FFSQuh5l0qGjU+ng+cJ44atG7hMj5RgMDPQp7NBEnaNVfwSAjTUDJA0DjXiaky/CJ6RA6
/PJ3P4qz61XBtp/z1GIXuggXMJE4GCp6P560WrNez2In7rHTLJNnUbPOaXe/EXm72rQe9Jp2XeOs
xjMNi8MqppqhTR7CXY1TROvj12f/SIDbwe1achzAWVHT25FCLJSWMJVbEUDu9aU5u7vsvKPTaWHj
A2jmDebPMp1+foUzWWY/mDPxtM7iGVnSPYvcdrqm3BDbqAqJl/Mblp3cXYh7u95PTaGBMQGk94CL
mpOPTt8V3kNIbTt2SZF/c9EfHEcskaEjfxwSQpsFPwjmeQ96utelO/xm2XW8UqvPgzjAWf5emvbY
l43WO0blfDmxd51n7yJAx5Hel45cRbYR/+eMXd3Oo3TR/BlLkPDipP6Hn19U5DTc1pDCd3n+Zsjo
W8McCmNv6U29E+gzQg1NnVU02mAeoFw0Xmqgss2bcqhjaAgQDdRPES/bLDGk3ufd7sloTxBXqcef
15RSK0BxqNtBKWqBKxdYo8gfrXLrmx8iF7J0Z3L9DqovVUsGr2T9YlphoNk1LUd5LHI0m6kxdTww
ej6jV+xSfLZ552uG1Van39LAPki8cDI4EPjRwPlZ3KhjT0v2ymDfYxWMmvQrZ9ZL8NbuYBxA2Nsa
8UUoJrxlbuIfYYd/b7N/CR4pPIrYYniU2J4b9yQq6mwcqGvBRLfY/Zecui8RdarcBh5Vp/v9mxB+
9eQBxb3ePM31W70v/qxzA9WTJgf8CdsMu6jVdK3RQLCs62N1QirqxJ0xKkGT2iWIMEnc0d2KSHmi
7kwCvWeq4gbqhRfHlOglq7SoIyGTqqde5T6h0CLtLcuCsSX5w9erZKH1Zkkamss2du31sKRR2cpv
XgSVY+oudqnYD0BEMnRFUwXkzLc0yUg03Kszc5Jo/b5IpCdlJUrvQ8rnBnXx+Vh3jrUC+hzIt9mE
Nl2tj/Cw1yM646hjKf6O1B33i+5reHyKD0mf2hEPibcDtW3FDXV7Agowx077igeteLmK7BLA33dk
9OmqQrgI9077xtdvGUo1l8bFca4sELyy45qGKgrbc0SfTEde5dhftXklDXtMqEjHBKNmcZGqhKJp
XrZF5gQuUfZwPsimJk2CZPGgnDSjh8p+CVrKsWYO7jAohQ+/rcN2PXgfH32xHiSWhPzS8AlNIsA6
gGJWu6fjNKOoox5p+nInRGMHwFAiHUIImejkYD+lXXIy8VhYqGrRR7EYGcxCE/6qfLftgUggRa1o
37kX7TEVicW9ZGnQ09jnIqbP6WIfZueh9/pbziOxjW/uTkVAra778pTlT8ICnMDxtL9z+Qwaniv9
50N8MnL5PLkHzf6DfLyoO4FdHICG0rAFxzxpnWlCi9/b3GC/qutCMSQxRLsM8R2mjEttlK+A36KA
mx/Hdzfxac1bACmCzLnUOXsjDDX2vEnNrwTyw6pwJPp3ounoY+TyLP+eseylo7i8CR+5+M+2Ai3O
vwxrFsuStQnf3omckeM6ZeMrVgNUx8hBhsA4LQqhZ8uw4FsNqGfdPiVq8pR8BCxjWb5JxOhKqT8X
uN7NttagWP9NCcYldnDdh6ud3on7ylNjdXWEpeqoTkwexChVgjm/w8O5Kn9hdjjpyZE4Rhz62Ncd
BTrYQQEic7JItUvxX3png3RcpV9H0pu6ksNTFEkntdK7vr5e5nvsyKmlOreJSzECxyQNkbMWCri7
Nl9AGP1dDE71Z9n0cRZdu71ntNHnPyAjGs7sM/vdg0KXSmthMGd6zdidGxicpuWCe4Fq2DxnxzFa
Nr1bI3Gm9+vNVQDHg2mi+tHlava8cGNY0J/bKYNyc9N7VM0jTANJTyMu2sdxzEF5kBSjPpSTKU86
PANlfcWrL0DZmth/fDTYyerOawZTgyDzWhLsvLr5nWWo25PI1/ynBZgxwTNAVRdlRFRVhqfCcKmc
cs9eKg1gpkoom6044G2poovi+8FF7u8+YQOtUP77e1qZY8ozs/kP2BULVu14eNLymB4VogwhM1MN
U9/pX8as/Z4qelG25e6xEF/jz0jaul8VnPvd207bpRlOLmn6MNzGokLOdgEe4Wb3nAuDxbhVGUf8
xrDPSKvr825hU3RmDNfdADyTe2jLylUF2rqmVGz8qaawL/liSE5i/lkLQZQT9H1noaEVtstY7fMb
DCnNodlNWm9VRKdxtVXqcXnUZOx52kd5qDYB7mE7jBrJOnsQ9iXRhpY3CQ13m9OzPrCBQTCY/IkX
xZZwd309qexoJLvAM2uZg5E2XMTk/rBrBV/0oQwsMPdhGTKfFvMpEWgOfCYHsbzzByJq0CyfBvxn
QJl4SgDEo/hr1kKRGHxbRY0pfCEKhznTfV2N+wSAflmxb5lAIomVAp3zqxbB4wErwGRG7JsBONHL
YaThFrAnLmhWO5R3OxayxNYY4CIukaLAW60PETiSuoWc9o7TeboTGjU3JHK07LCfh2GsGfmLaHzG
cT399x0vcmnQWBMOy9EZURsaqVrnOJKon/1ZAnQb0rKRAJ1m7P6P0rkc3nduvgqnwPscVPkIBfF5
iDDy7y3tkr1hu+XMEBDHOR7IzrZ5pDkNknmHYOG/zfSX1OWjV7c070EdaqLl3d7xA0THGPzARpDM
UiibV3gKSlBlK6pmZObZklzuJxATC1Wp4DMdA3mqLbuSosFAJ4GYx1oFwJu6GqA1ISTMIMtMMK+A
MCyR3eBMZSspfVQ88qApvXvNfgT1G0L+85K3YJjm9CQira8ctsEPxYgPCZsXQCTvc44Dm1/F6W4L
uxkauu189ZGkBHYzajge8cEgN/dbLNq1ilxW4syaax5iC+iXF8/t+qXZIbj4rZkdpbjXpTVMyNXf
wKAC3CVKaMD/3Lav8OL7H8T/G+JczbJqbNkEe53Ge+3sAeF7qWZk9DnhYzcStjYb4nL+Wt18liAd
pZshHhPXrQIOd+sykceeXlBhcLw++liiHBsps2FE9bBFaqWxb54NyCYbiMqZWiJzywsuuoC5AL5H
UAt/4e3OSWPnrVD1nPaBpdEKetcYmogk9G3+KE+kFdZAzMZsqMw7SXFS/XmqdP88vxNOusnqVuX0
IU643ivzAqXzjrtUN+2N5tDE0o1mAVzhQb/hl+9joQgWGiee/K6T1LbJliJFbv3mKeFIQyi5j22q
nbx1Cc9kLN3LwGXQUjKfW2op3gUXYuPHnH2weukltnZi6PtU9BtnKllS9jgX4l8BHRohZpwwlCX3
VLOBZSi+vyUQ7Lwr7S9/p18PeKIWOl6jxOXHsajtUMoYPW26FgahiGAogZ5nHi7gQPbWoR5598iG
GH8AWzgwwluSXiIy2M2kp1Fe8Whvq1jOA4gUCZK+0FKl8hPlgHRaRdBUykwuApgPNHk1Sq898H/t
g0ZCS1LvhAHcQv9gTH99lVRbzgiFbXhb4Zwve08hjrD2p4N3OUCPggPRZh6hITgVP/F91Jmxwmr0
y1NpvI7yfFVUcYWqo4Ydr0k0DC4fgQbqQg9TDXncOMv+T6JkhZZp/x5mbVF6roO94CKpZ1ERwlXl
gzq6/BEqW5nPVob7GJTnPbvR4BllDNWs1xi8j5EgEMmqOfmhcWkUWmdZPUNbrETFUwaSDvtQ5Stp
gUzT56cFzdEERh4sPd1aUxnAytojvvkTYj2qqS3GTBx8Z+hy6I0Oh6AI/8wKs0m2r4g9xjRixy8c
mROdExXbK82vTHiCIwt9kv+iXZkM3oFYdZDI+MkVGz4NbUpsoAZ9c+mV5P3e30aElHHJwofrLMSS
aeYyFMT8caVUAb26E2VmhbqI245UI48uIZ/Nn7pWea7OnTxe28dBcrv8Ux9Tbyo0m+aKvCTQaRgC
NFZEISyA075A4bRPMSH1xtsMllnt50R5VZqEGlTyOPIe/iCZwJW9KYH7xhbuLqSJLQDi/YNjjI4D
ef8+oJyCdkMBTGYFYsfQrifKtCZhleXdM5QKHVg5QxHTBQcmbN1ayZijuRVYzuOWgvHGQhPNGizd
jXfC0p4/Ur1eBzKE9ghAPs0idbtpibTex3Bz5TYq5HJHv59x9zHMUeF7KCdkV6MZFwuH40DsB7SN
YvZ3cXCgXQLi2IHGTrgR+p5Ul2CGdx1hwgaN/FQcm8wrsWnms0nepO/opbUq5RzoPQNPbPzhBTyP
OtHeslEMwpcXd12sWrNuYaap/01axx0mvHOa90M5Waz4NP4Bfds8BsXJQY4Wr7lQ0My9UZ2UdBpA
OJ+Crr7AGVs/m921OcxaIwU3bmLQzos2cB+S86AUa+Iha4UqpdZzAufOxuUph8jHoMPaQkzqnzN4
Qf4U4Xi2oR6EG4TyeUyLQY0toSUVmljtontQHp6UK0IWYELEZoZFpOKodAD1ii4LPDMesMWWozSW
tdb6aqVDXPM7VYn5pGu5eWb5AXd5Xr3PQEJnDP4bFO/sxfsGTEFrcfW85jqjx3cppHeyUQEyFfH5
iptWtIvoGFtZNqyvALOeXQCBoqIzksTA25SjqyvWjbUtct/wpCr4XeWMRcE+nOsEt0kC2g4TZyOo
VSxbyvUSRVO8JsRYD+3oldCIHwB7tyI9C2NcbGdoCtBYhlbvVq0GeqnVtkeNEcRVJ3eu8CsXjCA6
7PDyqHqFNhCTr4xePhxV2fDNNo4JQ4iSEgxqseQ9uOkG2xrsCLPwP+r2iCYKQFbvZdkYT2aIulvH
HErtAZVLRmxh2HeLeP6tRV60EPnI48b6+UNQx+8czsKcnKJSTd/pUmYTmGMHW1evz+fNRrDIO4SL
1f+9Geq0B8vZfz8Fi67uhgWDUZ/ZB7CumRvxnfqpZIU/ba/Z7HAmCCiz4VcJZemAmy2FJuCo43L8
5qQ2YCPU+BvpnNM1+z04IrziZZ6yesCUl+m6JqMTiOzkMy68Yhl3K4htnsN4KgEJvc6hq2xOXi+h
n5d2YV5EAyrLgMa92WzIaIFChlTQ6x125di4MFjPO8yaUl/8JMf/TJTkMLD6VjanTQIODDIeSB9F
x1IcwXpLpe3FvtKGXfuCFAGBUVnODe00bwDp1JcvbWo8ek4eT62DGYlLxD7IQR0Fhf9BsEnZHWUh
wOsxWnpyqQpWypsHavENniviGXeDBnRKSTb/5FbODzcmr1sZElTCsir5nu8FOhmcxoJxx/XpjKDi
CDZQh9SgARfU3yJAnpgKkjq2tzj/f9GveK6ICtXy3qOuQZJpet5wKQGZklgKBrwUR7u3YziRGWt+
67S9SHbPji/T6nYCULWU139QaBmj5yuwo8q46LEyPeSgD8uZfXqCb6TtIVw320D0+i7yfcIwxpwk
MNC6QOWu1ZBDlr9BdNz366mhhpCsaZQEyi2onVEilvunssmAo2SZSElKfKq3kZQD//E9QHYzP50B
oc3x8YR6nluzAri/StYgoO34h51BmfX57wIeDzklhcRBZaWzkrNEyWBSWPV9zLOsafvHx0/zT9EZ
uQGROCorlWW49dJxZppXmWevzZ+YzsCgx6CHg5xKJWbWVrOjpdMrsRsvWX1D7mXcEWUpfjyrn827
OBZ3D81YZ1pyknxyt6epUMDyt7ufdyvRQ4jBEE++ErqkTTucEyOvLp0KrpA8Sur9BINVCehPWKh7
1vo+stb5gRQ7EJqW2idTGke7XzX5upYj1OUTbc3Kq0nQnQxl/uH7H+NVcaDR+ubX/sPVO205oy58
LAYr6M3LHoXlXjVEQx/eF+LVJ3oxtiN/giuil++RaJLoX2IlWrJGsfngIVrnko/juYrbtXz0BQ0+
ePrWr/Fn481U8j7pYQVrkOQi6471eIhKFcR0f5Ua/hvZHqfoI1Vj24wSiHCuK1AupiWgDUSOonyf
+SLyExIpGKXbh6XuPBGQlD5bJmP4EtPrXFojE3kQWyWz+67KkuOHLomAq4JnaLC3XNyUnHO9HVXB
w9RuwGwH7wNNbBP0H3IR3jBx+D7yKvbXYVCqKcrlYXAPFgofeHITfD/0N1aOleQ8sdKf8uA6EIj0
/H7M3SffHuWgObmgc4+SZwZbZwY0dJ3OHtM2annH3bfHnfaqyOu8cxyQ8E5ubXW2LpH4Ehy44yes
TpcEpEbAi9CGwhbo3SMpfTWug9a2HlscVjJOdy9IeP294RumXEBiKk4mfODdAYivM/d5HAd1eKXA
HOd23vl9ZNPV4xZE4YLAzDb7zvutxhG0jfYV0iFMG1tjWKLxbRhAriJA7JCF+V/UUG/zS2UwBp/n
MEVFsts4Nf9s6yDq2C/MQEo8dN9LlOdBfsaatjKK3G6ij6NLNMgmZ6OThIrMJf+XyV7fjlSRbmkp
kR37IICwRbPq4IHbrSfx912SmuKwyIE2MlKhVNB/KxMttjEEzqC41j4kMOj1u+yJKcFmdlXkn9+9
nRRiNQxA1xGjfwQ4yu86FQDI/dQcusduaiE++2FvMM2fFlgICFCq9k98UtqJ2/bnyDk6Uf7C/XTr
QVHcHKjbfgsk09WHiAGeBTGvE+GWnov2SYW2E0xPuNV8NeqLIAZtm6krfJOkfrmLOonNDGI4m4+C
9xRqk/FgKpur3RCvP37sLxCR9h5TX3cz3tQ6ZI55wLsdquuEaXx8sm9XheQngR0f1sMwSR+zMN9V
Y6Y/SLvCwsGUe4Sut1XMTlEMYqxfpkgvVrKyAwyNjX4zftkP6+P7foPdpegjJfrnhNYbQ2Ojg38Y
vuMqtcajYnNrD/yX3l2yihJMw0hE14aBz/kf7AZXSPMcS9rh+JkFcKlkq2/pJ4Z0IrDZpkjIG2Yq
VXiaiKSaHQHQbyuSm8xqVGud6IH34kwFh8RDEqf2dslaFGgbxu3ORrFJQkKrpxXKjd53C2LxJngK
rsJmdEB0JCw9XLUvyd0+kXjmwgFw5A93jC6Bp6+n+QGWU0rpIg4v4qqSoPcdYULhF7bHLo6KZohv
DQjPQvOSa7Yse2O39R2BNz0JzoU2AafIKMAYYC0QhUI3TeHdJOYS7O/lhu9aSBafwM3al2VUx/Z3
Tf2Gi9hxcWaA2vbCi52E2ahdTfXqiUmBYUm6WtHrSMCecwcKiDGfy8fQc6b9c8mXmvg3K21dcpAi
lyGBuvidCfuU3ox5jLi8Qg6NL7swE5MhQzoGiFCaCGsRoV0xBes85ufyyrP4/4tU+//3mX0BxZPR
5R6skb1i6WqtSF2oIbYHQxI/w+YaoasRGNr1BR+14pbhM8QLgFE1dvOLdZRZsTz4qt60WIwp13Im
B4i6chUuNXeywpfXZ9sEwib+7DM/oOkWzwt/0K2bKa5Q3Kwltq9uNP/BrIb63n4MkV4irPPcFrPv
/6i7xLGX4aBl4A6HYsmm8/rid0ZiWjBjo84eKRE9l2txwlH5f322H0Zv7s1LDNd6gQuNbMLVlxXo
uIQK3wlQ79sQAJ/6+CtvZvyxaCUrQ1pFJ4dL02HWHZinV3ZkiYeb1cUKS8nhnAjIr+SQsT9e1BYn
sXabPwiIicaS5hSTL759mDwf/4pVXj6NZ/xd8aEomd93ZOGQkuZVjby1aN0kleG90/BRRBzTtEX8
+Ya9AAC1lR2i63AV4iqr5HY2juYS3e79iRiqkiIv/nALRmZlmpT7Lczx24hFtbMgBgdffXq955qp
zD4l3+nY/GnBmC3g3mEFOrQIlrvJ1lagSCwwKvNlRk/jzd2fKOvptfUS7xnEdbix3PEuP1+axcqk
VB+pSw1um5B6ofAByQ0YXB097wySl3KjT67dDwI1X6VwfgZyzMDVKyWCU4QRiraOPr9BkrUWMMue
JAU7gJOvG678Gy4pOfcz63QjzzUpn+YLpN4E8w8mTcna4ZpUjzlC7pWcbDsiqJ+HhNxLw9uEMEc7
09RtZndvGP8C7IpERhd9beewQc3kCFkBUAi8dpKkTJ+YFI0ICaHyKrjxJkvcvw+UGr/L7J4fUC0B
YLcu5jgiI/wAECPZUYk7mFo5nzeAGa5bPH5nuA4pxmhJjEYL7qyrHc5YljJJ4NIJgBMK+SlQbP3Q
zR8FQaYKjq4xt+Eu5W0vVE9yd2XBj6GoLT68c+joVd8bwF4uNXSDHgoBR4BP/PAnYShHgCBGLxCm
cNBO43ePZHqo9Y2LZkEnnPRmIO1wEzhs27xf//yZlDtUIiSSH+n+zAOqVO/zz7d9AAlDL4Bmvc38
M5xrTxOltrAyQptWQ0+WD6NTQFtUvFtW1GNUimNJ9r14al9Xubpn8HK9ATOKu2al3Sp515EwLDjL
V9eATNrBHZu9b+jAZcd47oLvfXit6bUNDQj6n2A4TU5FeFgThsL8XTDHfJUXurqSMqmAjizDgUZ/
ieH4+bbBzFszWjWC8ihkNByM1C2vtEFYoETKlGNHUo1O2RbWp5+r+dXj2vwRAGXL1kGgCZrohqdv
KKncX5m0z6acCK/7QH+pz7WSIpWqoC0jV0kaWQhERZ/vL49f5LBJcjENGiN7fywotw3UkEE5sjJ3
U2HFI36XJUvyD3vzq5U80c4OVcYrgbP92Ac938eoqdSXHFPhSnWWA1KjjiXKo1VGmNA589tMA9Z2
kTSvLb4EohD3xATSxfKs1ihbCgkq7O8NokXUZEgj9vJlXuxFjYbohMqugvlKPEiAWC1XnS/UhhG0
HyfIfUof/hrhQ8DtAPWolZNgQzrNUnknZVRjVM5IKSMl4vVJSi250JxN2Cc+hEAMeuP1ZA6w1m0h
qE7k5wKJPDj7rQsm4BwCvCs8TIhvxl5LMIgyezYVyTEEFRAoi3pyICiK3KxX+DrYUP5MWvkUXu0S
AzBBoEmE/5j6f+SPkPhBT30+juCbzTWU9Z/gkmwSFSVcEWJuv2webfc/JhLGJe5oGhJr5N5/KPJF
pYkyBqKK7dZCL4XvN7VZpv4mMmaEpxxr8RUPqLWgzLMNGy3BqervIzta+QbQaJEY65VW0Le8sMwq
gWhpf0C1uBxg2lxaxn8SLv04wwXomIRytDQdKuhw1usA/DcDe/J3UcedqVFbXfAxRmcXQu20qV84
7FRdf5xHX1NsF1BTXZXfDHt1GKkVGGhUfA+3uK1MVX6rUazLVIdoyE7+LPOeUpnf2UDCq4o2k+jN
ooX50Oqt8+xd7tmUEYB2u8C21O6vcHAqXXItby//fKJCg/IeK4VTaqpaOoZ0VIiiPCGtVyDUCu+1
7XRvYYKCCKwJ001bksgcskQVzBgA15GXK53JtRB7aDpSbhntYrnGRA3lR+z6Yg2YzSnYmd5jIUPt
dScOMHhxAopFUsqZOspdX5oSzcmmrL45F++HmPhoYCcdwKyV5j/+qc43gX/LiFgYfJu3KoF4ML+L
Kr8Nv5mbvDQVUCxJTS5sUAuUOEgFMLN9/32VKYVh36DXE0ftsKXzY5IRQWmly07ZZq+fbtNWbyiF
2pYdjgmO8+U5+IY1+gk5UVxaT5a8hNs3Swa/7pUdODRw3hC5LBOAM2fcC6+k5AThVjIiatI2c0VY
cF7QPX2wnhJJN2oyx6RvZNJ6nrMcopz8DRhLlHc2u92e3Naka1imTh9xzR3naj0UKP7Jov3l6nfk
mAH4ygoAxzaG9ZhlHNyHZ9p+sWVrHr6wJ0tisBGWpTdCthzt7zVy4KPCnkazq5E6o612DF6ijmjN
bqbPTMGO3bzJOjyiD8JW3LhIdra1/8jvkgGT8L2LmIc6RSYk7jHqtrkULiv1Gbw4NoLlVeswGELO
KVj+TE2owO4S1IsOeyJEW5iZaGNpFpR9TZT4t9+fkoSfJphtkLfNX+OEWPq4o/2BwYSAsD24izOM
mlhK6BRrzeAUOGIQEvDtUm+FHdXxn3Vq2MZzgpQwwreoj2xkinVnuG+aeT41hCM3hNV6goCQg2u+
Ng2TJLSM6xdcOzF+9Pb0S0YxvyHsZsSilp7GMKi8H/0DkTWaHhAFWHzrpHOzk+LPmu9HNnuOGbME
i9TkYlAT2SyC8RbfLVnQJYCozBnaG5R/EnDkX6ySKDMEcf+LH04caXVPH8raRsEog3JDFCLFXsXV
2w9LS6aEIgQ9jxiZpG9e6/F0XXFZ/1g9cEtX0xNVewTTYhvbbrw0UrKQWjGgDPNl/RvHJYPyNG35
9pNPdkY2LLHR75k/l7vmPeMf6TCFrBRYA9QsXEMofQCYHoOKnBXfpQc2k03dIXuNT3xxD3Wm+UhS
Yt30fURmDpFy3XNGp0ISwKFqnh+LqhtHNiQBgKMWJg//TvSsP3Z3KIOQQcz+IPzsR0xC/jRi2xnh
qLXaabEkHHVfEycom3IOjX6/MF/Vof1azyc035qQmf2AhDZiBxXZGZYePSHw/YPNeTAYpTiuaPHH
GxMth1R8J+fz2oxfE7o5FOrCAlu8MlS/Mg7NWxH70hK20U+TY0YEQfhMiWvzOGojk6h69zFZmHBa
+nIZvgHPUaZUT5/5tVTjBXd3q3L5AxG6TKBpuELLXu8p8zIeeo6ZHP/HmRxO8NanIoA+FeA6qMo4
s4uJjtgW0UPgj/p7JaDZMSeWfwnGvBl1M48wk5HzY2wSJUgDU30W8W0YDe8FQvShp823npKCPqgJ
OkTfbyjQ4/xiGsRo9lf/AMjrocL4SZDu2N8B7+juKWmRwPyPdCvqlaqK3Ee6Rd5+vE4yU2sBEsy1
77Ld+DMXSIuBXYsYRIYS5TF44nmKZu3+tbam30NUjfAiFLJKwWeHHc+sCnrxWvCy1D9I/4c0KVPZ
12L6fw5OSVgJXzc9i4LDrCKy8LulBTppCivEPCYyqMz2BiDeLcAJRzf50x/GKr6XB0l1QCgmYdT1
K7eR59Hm874pDn3QSSXmDgcY+yioMQ3pPG0CMnVgcJIUG00+T+Corv/FTTFH1MUiCBR1Sl6LFzcO
FVgwUmd82ZN4aKn4p0yZ1gd7mLxBnIX6QNwzj0bfWRRiI1LSkvbquHmfX2udXTiXYtqC/SKQgjoq
2p1a6inQyytZbKRtxMtUPIRMe85oWRC7tvpCBWDMHFtlGnWbq1DKPzLI//h4oPvntV1cPN/FtOWo
oG7ABKuxPqUxUdy4GucSTMRvOcHRu4D0FFFosbbjFuqn92ryDeaTHuIEQSq/UclsSqFJQnZ3wcMR
TqEfs2IMZnEfw4i+hp6LhCpU6HtHQovGJ69HBTEUtGPm+h/Z+Q4amzRY8KAwsyN5hJ3CMrVfar6b
pFIfu8EI9vaCpuO1NTxJwTKXk7RSz5+ywtMgWqf2kkhCvyyVdVYo95PczmY9KV4Lz8UK+eYJqvDp
15yqFZ4QGrv4RQtwClAzixD24xlLvw1zJ6tvXR8nu4tv2A+6P26TfDyv7dJ/Cn1ou0MQ1nGpA1yv
Nc/Q6oZFo1TzoUTBiaeYRRg+LwP8sRHkeDvut8nWf4NH9xGGvPIYVve2RC4Wsm2GNt6UukgK5CJu
z5NdCJC91ZI/hO2dTAtI+p66FV5AhhmxB5gmMMYaWKh7Yw06wNv+T8PIaIo0JPWyxNZmQHWi3Gp3
Ue9izxApYEU8HU0ZQfoL62huLGk36YqaaE8LguAR5yS3TfpdUxBhnhlkQbAp3otgEk0oJfXbUrQv
9Ny84O8EubzXows54UuNqLN0C/O4q9FDGJWsZNy6oLN2XRzfpWEV/vGW3/D2Hj4dfN6EjBjb4Qwk
HLwTIg1ja7sSt0qCMXgjXNdsywDNceyjb6ZnW8GMis6HitrSqy0gI9RGHKjC5nsH5qNInK2lkuRo
wSXLHosv0UkS/w+KF5JrsV2JzdMK1iOBjAM2GHUeGyzQROP/uxy2cV/j0hQ3FaN60yyRLFOyqJML
KBgB0uFavdgYaj5gnj2tZP3+jd5rWLeKwsi70HjuCheFq4dwRRZZzGohQ/vOTxGG4c/K99AK2zk7
gG68b2StpiKba9Yybn6wSB8uGEHB/RryRJkNw2wntLaAbaAF1/gaRYoL9J5x/GUlH8kLbBSH85Xg
1j0nQX5BMRfO6UhVsbYTICR4UdPB185g1/cPhWPCjoptBZPTR0ljjnIeSG77RZdUhxh0yNgwNW9G
RdNYS7VVcfir6QWSqgPdQrFhzScr4gB+V2zpJ42P9qV2l4gmtxolqLv7vbXVehylNX+G/K1PlsT8
4nt0rDy3LSjBNhU7X/EYQyVhYW4FwygpTje24NtovCop0CsTubquD/0B+plZbEe2SVbXrcU2f+B9
ygV7yHHHp+OhLcke8T1iskYVHJnlPMOWWNqjvanOtOZ8uQmfQI1wU9wylnsaOMnDOj38JMpyNKB6
0lmF2Q/kIX/zWm5QhO0ub3MSJToiH82T5pd0ZgrAAiOMf5xx2LQeNRN56FdDtIzRLQAYjYm9271x
dDV032lnRjp1oBBdO/pnchw5IdBGspSs4hrHuWnylxpdtOLFmNbAZrn4/gO3sJpviUVgKUIjgghz
Qz7GA4LQv+oZ1qXN7XQvOwDkJZVwDGVywvIGKAHfDf/fDlv3U5RBC6aPVeXGsp2QKi2FdLSzyNmy
+rdFD39AYm0HwRiw5+M7FdTixZ8xSAi1vc4aKwEwjhp1v7DJSmN5dLgA9lP+bdnRTtQRh4fPzRQi
2ty46m+B7nuGfSJpFTwigBnVAqxK22l8yCICgUrYCqSR7Uooskxxel8syLu3891WTDY1TlEqZrKJ
4gJf+EhvN61YvOOueDp5Pt1byDx0oG6aTvemF3cEfQm0SoweR8P6ozYrvWzqL6q9R/uRNzNElQ+n
fatPIUlIEFIJMSUcmi9PTwLlH4s/emVkHQEasjQnwhXu3KTUm5wQegL4SH5UL7YnNjwXHHTaEYtU
Q/SQ+yfa3uK2sl0rc4n0+Kc4ytFXzu5vTfH4ItQ1pJru7l5BjYxVM0S1CWSKap/0wCJzvNoOrx4O
9ErBpj4CYfBiwnGPxP72aus504zNLaQyw/UvXtBnzIf2GWQFlXaGsimxHVfd2qhUST/ZgcQEqxE3
1Qvr3t6LSgJyrBCXrDOQDmez4ewrC1SRpqqfs6D+wrBvRaZw+d9s7dq8x+UVD6qZbLR8zjn1yRAv
0RHYQ5ss7WhWAuZaM77Zm2t59+bqC5HC7BsyWeJKo424bAQCEkVOhWYmgZREjhhVxwcRYp5WKRYI
JMTmonxvfX5K1rVsTuwVCBaV7oJKKEg7IQw4O/0PdoyIyLM7ovTDqVQpksswmYjBd6uCiXGtyRzG
scWo2oAFbHv74Yzlrc0kwjWje8pNBFLr2XzKjiKyAc+V7TkcDi7mxDizGMTSNPKCsDE9DVRM/U5y
qfLMXlAuzV3h17oyMZf27gegPG1dErr/nkX2pOj/B9f6GL328/ZO4KnrbIufGNcfTjSM8f77aR3F
SseA0nACYnTy1tXoqjVjEFIfkwiwgEWcXgMuGYWfu50sq2rNaB9A+XeFZDK9k7NmOX0Iuj/zd2N5
N9eUcoQQ2QWgTbUaZG8m2PSXvnHkGvwPit/pMd5GR3/hVKKeBRn0H9oQ6i69/uoQ7jIurMe69be7
BM5uUiO1o/IIHY3pyawpyR4DKMh9xLJC2dTb0GIyB0wHCXjC5WIoe4X6K4vpdkATXWhFL+0IUmzD
ehrtbScc9PlDdLQOVGx0GTKfY3gWLCCOkd7Mw/qRLxjc5yDlnjO08VgI0hr36srerQZmHtpG5ode
U0he8XwiY0uVf6qe0yb0yH34+UnCDc+xpCruBdiD8lcEZJs/dbngmXr758O7xavxoe7NC7zL+N/i
rgmOmfBcXSrdpu94lnMXgqS0lyCWdeOTywwCsmQdE4ZPmbUP394Iih3uqM+zQHC146VuTznab+mZ
epOpVTARidJVGZmSqvg1HplqtEM+XX6VZBqzKpCq62ER4oTp9wp4O2pBZf4wQqbvh2JO9EzBQsqU
qYY3rn4U4A9VaeFFqYKrRgSvYojocnVZfnG1K6tOG7rBNZgHK9GnujJ4TGMxsMwKNJw+PnBlBNQ1
jwxvfWgTpKuEPO6VSxwYiQEEzQPKqKL951AsYe37tq7qi2a9L+UZFzb2vWFQzkL5j77Oj86s6oos
XZMjC2gZ2aJPS2GBlw3GR3oEgKqTCphnbXJCgdtL4fphdV0hXLyzO/lfhRoP1NPEV86Zq/3e5iS6
VyU1xC+v4BKPvOV+toWqTzX/vsAmzCZq2z6KB1AzSWRUFjIlywpYeJXJkAozzGrxQZRjA4L7Zxte
4HKFi1zPDnXm/2eB+csFH4Ca1I4WjvqZ1Il7yNs+kb+GskdfpPT4qM2PCbssh5a6BkNuleDscbvX
7Us10Np+cFj8iYX+pzcJTkwRVBug5ymUsicUUbbaQ3jdGs1t04dqu3WhCnKd5usQMHCTPGhpyAmc
vNvMn8HlR4Crys4BRh49yZ1Bv4vwmCbecFs/ptDozbLGoEXabIeR3OmhXQ4tliOpRVoRDDPLToqI
CG29QuCan6LTXSjMcZQRZ7HMx2OsH9bjf/xHsrCm7NPNMeTcubHMJeYi9N2zTRjznFr93cvfgaP8
4FKq+zu4YqMWXbn0HbmhZacoBBeyrCbxgtN3PDLwIiajSM6RcUc4njKo7qdLyUP+4AAd3fYJNePq
pe2jOBDDBB/fG0GFZUrytTP2+q6Al2xjkUQ+kIo0kAiW0Q7YIP76uPncg1bdNsPyGQaAsdKIqloM
VHHsbDgGj39ls1kJXlYctm2lAA7809hRLIYerefL1g9d/qTDfjRwGLFTz92LJvokCSuCLZQcoqN5
wE3NklVC+Qn2l8egtIYO4pcP72+EHWyP9/LhoIJOOmbXlWYPSCZXX0GZAR4D2Ua9VE2dKBj9wjIS
SoucIkf3KvohRBMk5Zpg4a5xbse3i9CWapLXrvXBWbcPpbm+BH1dF79UFjkUs1kirXu+e0a0W29B
2iGB1P8g/qzwIQWzNDvaCPejMDyX3q3dZL2BQ9dlcB1GYBYrvu6uJST6QfW5pGLWzokIJbggfCjY
MG1I2OX9rOJQQ5QEG6pjnu0n/uhSHvc3WZ9bcOFd12Ik2c5EbtKH5MUROkR8sOnqsKL5nALWDxIM
I7nVKUj9Heab2r+pFsiWTmziYjEUu6PtB0DPIfpnHl3rQ9tWdZxJwSESl6qpZRmsvTtCCo1HZ++H
mYT5sBXKIj8QvSvrD2CJ1TSWJfcE4wghmJp9UWzsWbbZGrLuKzV6E1w5pjl7Jwd7+63W74vsLlWH
DYk2DjHm5SXZPJfYaAWlvK2qCtsi9230STdrllWFk1dNOIEQm0ZFo/y8ORStFk8DseWhx2UHxFQw
BWA8q65mFQoV/0GTL8S0tlWkTCa3yHMYBLIpKalhb9eTzP0PcxcvojTp5eKeWGUzoVe5Zdmt6dC0
xdQgeXfwDtnOLqx0al6cZ9h5U4qP+m/sTturc5gfJ8KutA6XM0yF/lYdVm+dfx1qihO6/N2e2A71
c9BqvIqYeRmo9VgE5DIJV9aW1pSm5oCBd2T6gJdVtIu0CBKFpA8DFpMbfAdJ2Gqn8UWtcuERXhlS
BiWr+ldYVjnmvD/ul8EjJYzunW+7T1DWpGG7JXwzgm8jtdqUMWGcRNfNxvOoDgdraZvkofebJe9n
lPtEkZYWvwNagshF27PA+GVvT4YDe5rhr3a8MKK+7Bu8ApAE3UI0T2glyIKc1o4u3Re5++OgtM8r
mbjfU7b9GJoSUcV5nGIEA5AC/z9ue7DvhcPtQ847BY5NNNnLf3w3qhwsHSa7bwINtsN3Vx5wFp6+
58P2rspACmiJsaKPvMA/sASIn+5sIR3KMEsCOTu+4KGa0Q0k56uDDVMZLOoZjIv8w8HYiXYpWC1D
Z+wrmIvmdugvuXEFAGStL4bzc7jZ4BOjsQnCf6VQQNUuX3G2ekMJ8upvr1DQfH/681lMmjHOZjIu
zYgfd8F7CyqIpI/YyiOMs8aDcKX/TuTrGOUxklSoG7UWQH6ZWUhvL9oVUTZV+P6QFlXYDL+V5zE9
uW+7NbP1Yl8BqG6/WkMol9ypd4g5knnFQfR6XNP/+WF/Xmu5LcnTe8ZYF8L69ZA/8lfMhtpsUAS5
H4UwSykzPSmpgH28ohTDMTXxe3be7dX0qRBrWBoY9OwLBoc/pAIfOxOqnbXwkQHGft0hXG/vZ9IS
yn+KiBg2ojeaAW8swYFunaannivvCV6cUd+XJLe2Jqgv2hUsT28QsRNwaCJSiePZbxfG9Q6gFeMe
19Jf4TFlDQzY1iKk3z8+hVDvztE9GM5euv1wpXU3MTQg6NWj/qFOeqdKsrT1KQ+Wefp6Is1Qix//
31MYUfRLsV/DGaUpDQTbAJJ3irmej40b8znfjuYAfjqwApsHBn+V3flEXjNN6+vSF+ehbMdROj9P
D27s3+tVoH54Xn3DeI5EAbdMy4jpdLP9HLDw1L549GzLrAjiDtSynI77YzU6EDDkfPNkV4KmFUv/
OK67ZQSNsmo4Z9JKZfJgijSPbOHMOH0xJb6o9+wXeetv3L/WWCpT5wG7mVJz33EYtC8pNZb9wR7n
BrnjZAGgSFAU2vZrd6N2BaOS8y50ffgwki8+wF7S1qukXwXfWPtdaK6DYuEgfUJSJDwdnn3JYVOk
dfKQDQbxcd3EptlESzhMZQkdPtd7yp2/IGvBUsnNaHrYLPX0QzzqIs4cOdsrACi9CDBv6jS0EzdV
6pV0aIi3dzhxf3I0l+um4j6VsxS0bCrdFoPb+Zoqc56HC19zwNxXB5tgnRvDi6K85q5VSv8SQYR3
1vknkSF7nkHOOBOiImgsAYre0QgtFdrRzvI+EbciuG9SAm7ZYouxA3G3Qo/tvbqqOePF3aNnyCGY
Ugdpv7VQNbDii7dCeg6HL0paGazoF/I9RqfzFceSO3XAvK9RlseOQW1uYQE150UEKqcn9AqwAIVE
/FI1g/auEtCfTiZvHmaP2yy2YLE2oF4c9on4g1Zt6fy2/6EK1scy3FQZp6aLB374BHMv8LS2FqWC
EWHnkHDtCkk5u9p72M7MOQ7TXF7jEdDmUVSjGbHoVUlDnV9MJpcbzCFqOYNbwJltAe2qfD1zwqO+
aprcqKpKhqSIjbcqogwsaRpbSLrrhQH7EUl7uy97jQhY+0ZDK/H6105ECBMB310A7qpbj0mhM6/c
Jkiu+bNuUJsCgR9WaHBZky3aVY0WDIOSimk6mpa7+RWoVzQF1CYFJJ2rfIkuJEQTyrOuK1vD0C+G
aCslm3mpvYgV8Qy5kYsmXPbn+UzfhyC0+5wGdpwUf6nUYNyptrb+VNQFKbD59+Z029oLejrBuoV8
Fbvku36B++ueq2+Sz6l6gC7P/uIxQ91Kx5wjC1U1x9GhD8FZHXki7GmS+hC9bkQQuGtlwKyeh6Hy
pRkuF5rSakUeZzsr+7viYoz7xDCgsL8hEBHw8TtA0kqMpB2fpRyJbrgzmXKwIcROuY38vUQjyff7
r41AP3A8QU+Ziq5n4OTDS7J03031QytlEGHBLc25HjnTzFLfkQLHnRLnTMmYrBvwKu2b0gsq6T8I
dMbg91ajqBCCUzgdY0DmbzNg4HEsSfL5Cg30HD/wBftXEGjDmTIai0+8Rz5qeub5U+8GQd1Sc0Kc
bme1IY3a5YePAikS+xr2wjUkaF6Kr1FzSGRzjQlGbRfgu0JpoDvwKrwrw8cdjHR+pUB3ZrGveoll
YdQGGwRTC91Ku1Ih5M4mknVBZavQzt6/fh5MOnTFkMVQN571L/nnX4a1ciJhB1ZCo2Whgk8W/1BX
qqFyon482sU28RyFiOPF9KgasYaaAKvfaB6A699NDzmEuIIyc1r/NXCefsy/Lw4ymQrYz3xv7mDN
hEScOFfhCPU/VmpRZj7BV2enjN8sQ3WwaT80Dwu3FKBmF4rXnZp9BCDpAi94Ip7jSQHrs4wko9Hj
9oBqtvuuq5CUt0Wm1/GbjKxwNYI0NhHDFSv/ncJgiW6GbDfzVTbigX0YTwD/UVOJk9nd6sTgoVPZ
FskraitNu/TAYp3wTIT5WaXUl3QcB1D4zp/LeNhViXGCPPYBhAzXKIWzqV6NgAD0yX+FEvT/yW13
fFJ0+CCMjsSo7AKta0HVroz17bz62BESKb0//f+w/PfK8XO4QUQXGrWxoVJzREZKLGvlt7psAtlL
l0LsmbhFF5tKY3iEURZEv/DPkMNaO6ofUNOkNFupVu9BVnA7blcMk6MFy/bmj/jKHRaBI+8aSjsk
1H81uDkd5uiGGSuvVJvBLdiuiWWAb7UFUD6ReJ9SrwYTBg6sq8etVDG+/Zyz3zc7b4M+RCxbiekn
7WnJps+kMvO69vfDHxs0ZtWZgWK/JWKFzQFsoWjRNURfguDQHLMmSihevVtP71kC/f2eBfO3sCLl
pQcORUj8SAgVXwLkdfYJtpLvoem9nmoW7UzQrj3zeC4Cl+cyMABB1v4ZioiTs/+JLsrlB9PuAxTC
3V8XmBFARdNBO6cXGDsY+6yuGkDPuyzgy4tGMpThSPfPPE/eX/1coS7DW6zRmp2Jdact1d6AOmkE
U/bmkC5hcXM8fLFF4O3KEhchR/+a10uGFK8ff/EQINLRA74c14ZuRJHgDMLY5yItr3BYeKZsyZyb
i0kHYU5r5wGY1q88CFIosEuDXCHxj3dpL0sAZLkIZXq4zabigK2QcEWw8yZQYC8RVnlLcacgvKvD
S2UcMxjjWO433fHmnSEur3Y1ynQirS+7o8HS5aVG/djQQfEB3fRoX7vz6ZRiHkrk8/mnbOhqJgw+
jaSCdtkqh2jCJC6fgKQBjw1ZqJQg3rT5m54pivZUNuowWv4IYiAvkHChOrN2vu8+D133D4+hf03S
pwTjS0ya6FhmwVG8h3cTxz0Wl1bT53jJx1bG8k8fmzvR/VAQGi2ke5UsY+xXwTTaUhcFQq1CABbP
AYgpFkUgdPtMmScjCM2TNSRqSLV1uJRqik87Xkf332TaUOGTZTJi30xvPID2EplGUOHFm6Y4YnDv
2UjXpHoAU5IZzihsGG7ftxugFlU+iXnwjCW7J+1sdkLhNY+ro6ViOuNDkjCpPa39onF7/zuBLotW
sRc3MvmuSICV/AQsXlu910jWTDGndA+27Z3Tg0nvlkNHvmShcx0dCno31MFZYGj7WeAoaEsS7C6v
krzGp12Pe1VbXuLSYYqD6VBKaNxNl3Lle1DDEl2ZEpZQRGEe3o1S6c0nhkmFNWxO3hpXzQbufJhr
z3Vkw/m3fOUc6YzrfHr7N2ZcP1yWoj/BUoRxs1UJdec0Ir8oXjRT9BGpWvJMRsO8zTLmEbnoijZ6
bXDYp6gbryXuaGTdmWRt1wIWxxxCtSu7jzLrfsUDSViyT4USrjKCYYgzyu4MwqFp6sihLcxDOCuX
Rm9nx69AO3U4obWk+x9JWYv/OAANxzWvmfi5t0YjeY2zWVS6bu7dil5z5f3I4+jktjAMrT6Bh/Oi
40GP4VQJNAb6nCRveKoNqQaouD7SOP2m/wovuOIyzbAWqERrjxtjAcrXgu2i+UnOqoTbH8wX/PmE
h8K6H8quPPXHjMrpH44UscCJdaz0xRcc/IVopT7AxpseuoAjRabBuDXI5dyxeiCHETeKUMsovNFJ
zZQJxZxnPyE+B+ipivd0QbbjK3VucB5uhGzffu8HlpsuwXIbnDaqYLn/WU0hzA7Tm3kQ3q9aSKY9
mMOX3TQPL22+AGhlLOpTIaB+43ci6KUdqKZxc2RSENF7oVOt1vjNybj4a9j4mEfvGEXl5P0aF48B
EYvP0UReNxd6hJ8Rceu9zJw2YKWEJRd0+0CuL9qdfY2I6eGi5zGN+88GL2KSlEZsbeS4rMT0dxXq
bDmwQd83yJRHAmvoD1CxHXQQtWbVvCeY9I3xryHfou9EB4N/Uu+X8i251F71CxzYX/ZM5aCs3yA8
t8QwkDnEwzWgt17Rr6/XR5VhSQ5D87rc+SLtinhjsk4dvE/6P3oT66rxinUMM39b6YgbUZ+tR307
p72OsY7QTVT9GBARMlZmwmJ/e0Zpoi29b4fCv9eL88Y1ra/zondhru6y+zA/q5cqhCgg/2SuGdII
NbNH35xmsn0JGo/EW614ENfC/EyzvjsnWM6KUtP2H/xhs9pETWVQ21KnqlOdHYq4BL+u7AgOs2IY
OYwxxqWwjjJbCWtwvTiyqbkPu9ffZuv3M7S7ayLlu84GulQmH8azOQdbIMIsPZ9+TDt5pk4Hpn88
dz5wxHIjJFjOgMG5FXdQ88b2iJjt8+CzAClPfSUfmp2o/n6MsMPyMNfAu2iHrU5jLycMyhy8G6nS
cl+TV0WqWPmUdS4d2U/DHGuk3T2rh6E6z0ROHplurmogsCHkkKz1y5CGidkR/QMH+GBHVBIms/7x
/zZdXtbdGSu21ZH9UvrPnYys9iVxMkVm6b0f4GMMgmVaJxVgKjv12DihFTn6P91JQlsjfXzcCDp6
/XzGhuafdc3OBTKIzYL5F6za9XHaG3oDFPvQquxcw54WbmPLMcrtWpu8T/iFoEUJAwPr/IfY4GJL
/Hjh4tnYE9AE/YaFjgFeOWqb0qvIPaLMeTgqUnSXJutP6gSzYQffU39wHYG5Skg/jC6ekh8PN/IH
KWqqm43khW46ljd1TLxNqUSnnk6psPIciKz/AulKCzupr5KtW7rp8XySj9VQgsXkUX5P4wxcciJG
ZDass6r/8nE6KHlT3HR2/9esQO8OGOOMZJaK5SYw1Iiy75F+EaUdBmCQgXxJ8t0anHM/62x3BSQT
Et5Zo4XUS1DRL8ZqOXiOf1yCLvWWjWMtvzSCpU0icXi6QjAXCedka9/f6VKtjewVbBP9sylhth3x
Rj0d0+O1XYKDvTO5aiWa7zvnsNPvjLlPGuXAoW/rhIy4Fsx0qLUAwfRMovna06hePETJgFYkfAK1
NFSEwbctfaiEopT5Rqf0G1Vvh7sDwMdjuR107ZimIoHBLBKVYf7oGGyMevQ4H1KsVu+cHpu5PXdg
LB3Qx5CJN9yOaAwcs8HzpqV1wp1nJqA0+M1K6pnmXsBqARDihZJDNl1Zqgm1zT7RHQMS8uurl+ue
+vuDYTuGd4gs3AyLkgRgoap+fgP0yTJtVE4q5UQ33fulWN3Nppazad6//26REzwfCOBygScLUgKb
amXK83SWzHPsrw+1KbN5BSx4mqLM7MEmJMtE4XRIjTXhGvoS/TdOz/unhJsbU1u5eDwENpxCb4Fk
w+nXdqFsKxKrixK0c/nKzR4fKfl74PQzJvVm/lL4vIJZZefEbuKnukR86aM2v5X6eaWUjw8JBDf2
9yMJz4t6q6ekYH2fGG4vhsJAzI0pWJEKoBWdn43EB7obCG/a3OYIroWJkPs/jzDHfMTycjhmzybq
T2AQHKXl+590NFInmeHNEDlISWSh4se62q7IHoEtd2A6MrmzLevlnEJO1HXr7ssdXmDaAq88al73
u+GcO9e8EsfCotVi7QI/pK94XHFnImh0VTtPdfYgi64ZzgpdzSE+k3WhbfEZFTVQBg3n5cTVl3dt
QSyBxxgGkjgqE8nwu3kJhvh0nPkGgr1e1/bKxx7pQXqianRytykIvw0E4+lGZCX7AlolJ82ZsoXx
VN6QOPe0SoHWrSR8V3pkdiTszpjG2sPccZEnc+mn+N5NXLVTr5orvIg1UdjHCMio+nU8PpXQfADE
8NTL2JJ+OVa0t7paENsFlSz7+OiB4rKI5+TA4cI2HXNpUSH89Jl/yfJLKZDzB0wt9AxuQc/wyRCj
kN0GczRcyZruENAhPA9GVSCcb9wQYVOCsEX5qShJNfpKzzHxhhvWkvsk71HSKsUfUnubm0F8g1hj
fVHPiY00xb4bH3DkbLSY8o1Ju71RLX+/gadklm5LGMIMl5LE1LaciLvBhGRXXjKIHx7H9J4ztU7I
EdVJS4+Pn2lZ12SnBV9UhsAvhj3O5DhEPtmwfg60CFU7Ax9rYHWLZo9/zwfOrXnFTx1BbHllsjTo
pQKwpouClsOkPLfAMEU5TQf7A34zZp2yINlQDIGLpIrXGOpR/nNNIka6kd/ts+GJbY/HY9yX2kuy
d2bG+v1nFKec3pXEhNYcslap9tiUUsh3BJlRxPJ5hDRa7pNq8QDmIK6FBLNymeePzcozg2hCoud8
FukbhnZ3M3BxhUU+5WFjsE6vgQuxxmhxw1WtDpi9+I+PEgnpkDAUWwh7fUrTvrnVpKfJncJDwgJX
X4V6Zu/bXTQ826Hg6DTZ3Zg1YOESGYg7x8izxsVMCY2RaMPukMASNe0610sv5Z4+6JshAKkekY+s
009W27YvWO9BjfXJYTaxDQz3D83nWwg342rL0yfv2iGMqY0uk+AL37dY6cZEuqYUm48S4WsMKh6Z
7lb/pcuwwbncr09gQmYlHuytNev7H4x3j0lpnYaXL+vEi/jH80D3eZb12pFBsfZvctDQEckazfGq
duooO8nQ8+zaV5uq292hbqyDByXdm5MX7zdky6XmuIXGfrjkS+rGraT8+JuIfZfbmbvX7+2Gf9NO
/NW2aCvetszPisMDStGkmo//KHgm6FvXktAhgWRauRbDPUZGbYxHer82jgow9gXnvqCuOc2Zx+gz
hynUuo7NA7Ukag7GwFULTD8ne1qrrvupMuUZoa4v3E5jLVC7vepUElWCuZ5iiZG4DxhHCCqHX+oW
yRrUeV3MiHPwDpxdOy1h5CIePeSW0p+LTSgmjTmYd2e++NtCCS/ViN25rFXe8M3ZBA6WxMTb0WWq
0Jf8z62MN12XyOxUyKBmwV1paUthZdI9oYuOOtUxzDw5eb4wT52k9VbWqk/hhiH56NtNHNc1v0GQ
uOqlX1MyXUA5HEqLE5rmnFnWxNfK1EYaelmskl+nfQ6lYraCYKEOO0kTUKXDrQQixO7e7xbNrTJt
1qxtVCqJ/Cim6GbIgIkVqhsC9MGywrwkbx/aQmC0ICsyq8smPZgPkxc+eWemjZltUuWUhjg7usfv
Ld9K4eWJ/CwLnO6/V3GCF2dmLikW4tttvH96E8J0gGgO3OxA6lNlx1ngKY+VyAHvHR5luv6e1c4J
275ncGP7dQONHQJ8mxnpOc/nUEPhBtPIHFRiFIWaVNhYhV4AvN4LgCO4iJuAE2kExcABVIAY+Zf1
GUS3sOPsifo2QGa93CMdR/qzlZ8f+Xt0/u64gtssPuN/ntsvqlhfl+3+zcDaSsisiO6aoe14OgRj
St7Xbnc9dNLcgZDKYWKDcJUXOUi2dJTTry5ZjWM7UpcR+dmrCA/1aHdJ6BuXi9PhlnkDFW72rzuL
KIulzD/eZ1+iVMJNjdSNeKq0/tjIkPx6AihTegCSx35AtzjZ0DTba6yDrNB2QFfgD5sV8YGjYppG
ZWFaWZLYstF4u/W3fbUdma/n53e05fOj8TrNa3+kVA6uOx7qgi63xD8rwyai4xPib8ii9rQf3eWp
nGSQNKEzo2kFZAG0Guw0dXaaq2KbOv/T2sQsFppCzFqRKo+RUpDhMWtL4j2Lyl7/vLnI/R0G3+3/
L8Z5X/LzDN4KK1dwghig90Nphrd5CR5GZeN1MorRFrmCWQT51WBQHpK8qp80f2x+5oOd5H0FY4B2
yOXoHv9DX3jEUtOMs8zzkkTBz/2ldi6eEjOQaKNIK7kTap1hx/QUWvvSNZQ4FhnODlUOkDwtQ+eB
pDC1ij8Aym0YCoXKTy+NstJ1aCjyDNF2dn2mWfwe5upIWSKxlV5g1ZNESQen6gw1nFJrBf2zdLb/
d69EXFI+ztcssOvJQZTbOFgdGkRat8CneXZwbI6h3rhELU9RkRG0Dq/3Z1750CNAx4Ol1Il7nO01
vcmw9V7nbTv2DLRhGAVKzWBu//vGjWXmouzasD9lGPeGfC1zPLNWKwOWM7wPyYsUtO8XLEINU/eg
mfBxDDgk88ln0AMw3u9XUEdAYNogBXbuOqGn69YOBwsGQoE+ShalAvfMXjS994376pU72/Ogkoxy
FNXjLc/2bYd6ACHF+G6BHJOdySdIwX2b9WYW8V5o0eNwNPpEf+8vZFAavJwgA6F5xcUN8wA9FbXe
mjFrw0oDF5ZshVFDSqFr+aJTiQi3w8f1Dmguzxvhg1CupCgr6ap4ZA5Jt8fjAEYeavxc5TX3TMJ7
lFsGsno+Yu7nrc22GJuagm4DyGsEsPvYRY6ZZT/qgTuBMejPiY02dNl6PlhaFIflANsQu31+U4vH
Ww7MrdfGLyipALoWncMsllwBrbuckyFJ7kxVytSFfNa0rgIjjJIAvUri2u189Jlj1nfLSmgZ/Hzf
GBcgoBww16Shww7s+RrMkVYH1VTyNZJGjIFneXAMaSLAcZDN1DMAvDC22QkJx05UBfiCMNJ8hvnh
NvObadY6ISu7SkSVzHX0qxP4hSkit7VWN8u4Nrf/OpxE4/QxZinms+mZkEsNT8RgSuI9K5IRD6YF
JdxKOACa/P4cd+uw9pHO9NB1EDtyl5cQ1w8y3YWkwGDG0KS2h8F48eiqsjoMLJJu1S84Po6Tw2uF
T5vlUaYWfl1C26reci/520bWny3QbEQsFrIcTucLiXsLsx1HfCSTE+hIqREXsnnSIo39QOT5FLzz
L1lXrkDToBedt+VhEdI77/N4x1j24XvlmaRqp9qSFVHJdSTHMxuMqmsjtWJNIuhYr76ZAzE8nQJ7
P1a/ePd4qrNoAd6OUumFizuoNuGl2eQo/HL1KfYuiW9jBDW9Q7bH3xcWWTf7o1k30PAlg7W3t56B
EpJ3AbY3PQsNQZmduWRW1Ext5rCDshMG8CIkHC+2hQRXSUyLAhxhwcIcXaUOVqWYmjKUJDvQ6rxp
335xv+6F38P+h+SeFdRY1UiKQVZ7URsgql4XoOPtlu5RgRPUmen6zSFyV+1g0Qoek4wIgxuQMCoN
URlwTSBZitTIjW+sVQ80NcvHNsYLEu9nfst1LxHZsbdqGuZCpXZX4b28jieFJGZMzXbGcxUFAzGJ
VjHci1zFczqTGhXgU9kgGsbjARMr+LCXREc01ZkWHdslPJCD8hbbH6+E1294BdPuwBMyaPordW4y
KGihW/QLuAPTPvFdPeOfU8KhzqeGLCO3cAi3OLPRdegcVMe5oler3cH7dJZ331+VZDUg1kVOOioL
WEBkwqY4s4Tq3WWiQJF7R2RFo+MUmtQHl66IxaPYfSQ/HA89DL/gjZxehbdDmuPv2LJ4xjZY+UcB
1HErhwZW/RD2nXPc+h9Iy0eRa9PGDwOz7qovgtTWnPp/cFl7JKjbjpQxDOi9/MadN0SsUS140nyB
5WI1V+GxXkoQ4WZKVYgYvCNHgmkyVmZBhCiHO8FFg0bEcKHHtOjc7WsLUEZTqiqfkK3kN1gMZp59
G0G7o/kw915qwzIJwNBfslBz2Jtu12Nd6CdWtMyNm0P0ss9DJig2r02hiPCMORgyhynPNEvZfwbb
rllBwyVdwIhwxbqn0cHRSfDw+stfRolA8FT9kdvN6nWD/EHGbbkppRgbA74j3iRcKniSz/27U5p5
nMrbuBnW+b+30bOlnIdhtC7sHKywKPS4In/m/Hdkjnc0yNeWmadxSW1qQiAteCAezlxQ3uLhTu81
EfcrQiR6mpybdtGZ5ww7LC1uFuXMrsoyjFg3AdcsrpFkHToaSkXf9ULdm/7ZpF3wVkJK+QU1DhjS
gaCqc7pZD+yU7GK9JwbMvJW+X8i0F0AbyDFEylDdAbfQzWz0WcjXwQemWFBz77bmzOpK0WPxP3ei
JjOXX33gCt64NhsrlCuLMTeog8Z82euLA/l+VmTDVfcaDDTClp8wGHkSVUA2gru2BhIygoL/iL5b
FfPY+aFCB1j8qh/wfte+1ilwJDmDGacwA2eznObEsLewhP+Q/4Y/QgEL34Vs+j45pJ08kMgHRgE2
w2Lggfx5ZnKRSutHcTUYxxijWdVMDkU14furtMkUnLvkW4i5Rq/whCuN01B3JX3XK2pIyq10a0QY
fgiSd6QH0O2BgWiy28UCBqOVYAJDCoFX10vNWkiVM35qVxOfcUqTo2QBS4A+SxFkAmDGXoUhFsG/
+O7m2JSNiR9i9T0HAQ6z8C88qcOykx51HGls+AHCmQRUOgX1ZSov9JHhXfryCsL9DK7SX3gs6JlW
rynI60C3kEz/Fp+4tPFpCN0Q0rLqFAQ1ZJhJa4w5x58nzyXOFCrGFjkqtYeeCG0tCVYNZO5F8FGC
If1q6Na0g1tiPkipn6Bm60x7Tc7y34VR5Mxpwuyn2nvIcQ2j4eR0dRsVWockZIXZKBI2CdPxcs8w
gPZC4XZWaufmrgYrcitJOX0LVeKgzK5CLN5lPDcJaw54/Gjr1T0j0DZhF04s21VDkEpq7CVWoEnQ
rOSvg2THSSx2OALiCjkhsdHulZLh6pdCEObsr9czN61CWkYd/PyOWyJz1pLAxcrTeqU6HT5QJmig
9Y/06+6qck34j0623kSQ/+NEIx8dhOIUsuUK1tckiB3NVQ5cmWteQBMN0J+u3DmKkgkvGZ7LfI6j
DZRHPl26gdGO9vYfS4jX8+wSK3jTs3T7FbDPYm/ujZ+KkGsEwFuBp+8LA34V4ds287CqlVRTwi8b
n8uUm54T/3GdZcaGdo5LVxYe1fVxnJowyOetJgOOPrM5nXjNi/ebzoKQTlcw4SiGm4NC+3SpLRKb
F4yw1IfI3kyLsCUZ/AhRYeqGxDJi4zgtapYlgElzGBGJ3xLbHrTBrkKhU7yEKJXaC2Rjl8DqPK6S
q+rdOd/7UJ+04FGzpjh9tkep4t3rZCkXWEhnjupJBoEIqnqTGs68ASjLCoqyydDiWZLLbSj51uKF
KecysmI4DFAaBGNSYM65a+SNuYQ7mNOypIVNM9+a6UPBjAUfcrLHW4o2gUJVZDONGPpM0qRowvGb
dEtc7zqKmEIhzUbnsMMokxQ8GJiY5U5yVdszq/Q86FshuKFWpf6yt8THezaDtm/eIseUBFt5GOYQ
vsrgfQWPNTHRmtxAKAOBe/4UzaYAaXMdblVfzzOgRj7ZFiPaZt0L1rqC5lrPcAoPQwTUjPIxN6j4
A4G6ymUrOpU2WSGK/PhgyE3bYjjv/DA3Z5PPkuhbH+P90SdIrlE4HdKZx5bk4PQXh5jR8k7Ep2vZ
dkC1U0KsFbC/jBLAb5RuYRGL7Gs0jYIms66K8MtpVOXsMaTT21D1JK4a5qPIxuiRJ+4DVjgCgPKH
Ld84YG0S0DlFinHF/0q7v0S1OCQyZVmRzOEbnPp/blmSDSR/Uj3kGrcNoaX5HhsVMP2hoBDn7Ym9
/sG+WH0wDMqq8p5HMXJYxjV7D4nEB8yBBG1iUUDoFFp+BocLinvmO9q0eTMpAahmty82FXJ+4DcG
WiQRqR8AdDYrMyrIufvdekwb3MDHs5+2DCianZuV6no7vTQ0DYuMR0KHVyUB6tU5Oqvay/4IeVyb
Z2Q/LvONwB/shYuWa3oh6CTe1msli3AE13xH6eY4zPVVtJoJ2WewNRBn9cQRiwJHQL5xsl8pcDuq
yJi4wLXi+vwtJ4LXR0ZGpl5jmC+idwZk6PlEzZUdbaQDU2U2ZZYnAuHjfWEXG5s0jZAll3/uwyZ9
VmN9nSY+JbStR/jkn+7qR0VwIdhkCkSEqgyYHXBvK1heutppmbC1NfORZu0k46dGvjPUHC4DkB5X
kUxrkuzg2Lm3BlNncVLZp2LxwzracCTNLFhov67v9DExPv40f1f0dJh24eZSeYPaZDwUOmjTPFk+
YlngicUt8m26bVRhwQ/99kNYvjc5A106l4/A8dLUDcOz7Bz1K7hbBJEuq7rXTFWGO6gRtRlldMPW
Igner6CctQ9JgOJTyRA5sm+DnvpovFPaLCl0oPPlo19qWMeHR4Ddy7TuPiF1m4TMckoiWmNKyqEH
QiNVvt3fJe8BSbZXVb/aTBqWUtHVYvj1UEz3VUaIy0B1A51bkZ9YCC+zVLVhhKiYfmOJhBstkZfk
c3yiA876cojhuROarOGC9+TW9cHLKKM5QCUDjvevXQ801WbUc+gdXzfCKgr+0psjxL0DkJTlHXSl
Ut0eV+cX94VEvWsbltjYVZVODNP5zaTdAWTIo9ShpOp9OCH6dpx8cd6lN7bC5V0ZsFGqR/SL/95T
MWgazLTwu5lhLcntji6GHvnhtVxNgOTOdF391tJtA5wTsBjYdobtz2s9f8RRw3c8VXvisiQ1Cbt4
V3yni+5AOLTjAFeBz6S2E7ds6xdscJip1o5fiig1jjAw0+XkymovQ3uVGlxPzhmGDhPStdHaIkAv
0N22sbpv29C4S/uATnweWe9NgWhOWxT/oo/tYW4Zff22XoilGZQhmfvo7NNzgOMqM9QVGNqry+G5
TvEMEa1kGSO+KeynWFu8G4UKk8sasPMkbEpTXO3RyeV9xpvFjuCTBuW4I5Xw7Yf9anpNUv28t6W4
D3jzw7Bs79BUYOwmEAcJRS43WgUX97ycjFgEqhWERk9tkv4EPYVyyFHZUthhlTmToJIYjmtr+Oek
5SprAKuVdbSjXnHPhW8RdhAd9HXdIgfc6vDnxaqnydAqs8fiuRo4KAXdiTSg95Tla+9u1xIoSUkf
eDOO8AhrKGYqJuKvxzNp4bXgYENrbjl65NKcRoneg1UXXMMaFaiCsqi+OZKb21smd8K1aMcNq6Kc
5nxrumhPsLdLkzyXWx/ChmOZRGPnk3g4N3+IXpdKSjywltXEDREoxYsBP4RGqtfQStpho1ole5rY
la/aCNPRtQ59BLFq/HCP71n7iaHZk6OqiF/P4Elq2yqgqGxo5psrpNwDNVM6h53JHxIBe6+O0CE4
IiRndtyAEf/D7CEQLrwPdM4AXU5as5ozRyRondNdAizFLfpcCZiFaoKXQVekexADOT4t+LE6QV5M
Wip6K/Kx/SbGpZD4obEOYyb3J6pqnTAdTJzqGPn929su33+vAThwEzLklKVkyzAExvuBz6v67LSe
KQcW2oA6tk5aajcSCDIFRjOEtTSNIirwUCzhbQqKHiLt3Cn40XSP81Hy4nM5zVO1c4GC0znvIYQr
UlCCqhg3L+EGS1B4coNYTpj39vacpboDN85wNoJPkqOINrjbHI1m8H80AEkzAKMdleTWKVPBubpd
BRwsHVMwEJwye05CBBfm+GK0AVHDWyK/JjURuhOMLUlLX0ijBK5aMgYeSnQ1VDfq1ZWeT+rAaJ7x
GjwH9Ayg35qtOr4SIVMGEiXCPWToU1LWd3j0iXHDUlqK5+qQ5+EfU7+bdenP07AFct1GB6mPd7o4
yjFHrWU6K+4lMRJJO2q6841EMGRjN2+DiHpOhc56HYokRP/6r9Jg8FqnqquS6qE8d0rs5Xh6fc0K
nmdfgzGn+Qvd5i9josrhOoY2twwTz0NCRLzld57hhwKtkaD102Gw+CyCCjj2wPGYl0rbdGLpcNON
0u6chdtn6CrcYV6wL1JUfvWj5TrhZ1+1jMxjyNXNnLyP6vFE3FmGt9EvRtI9QdeZysLwlE5VUtSy
5y2kFbGWLvXdUMiPUCMgKqH30euX5iX3L6QZum2Gtbku0gl/SMGsKi6/r2vN4jGkvTy8aN+Fmumf
JVBRv1G++pwsbxNrBdWZr82Rs7cSBnhZ2aJ5fQ8y/0j4YMkWTnnKXRTJSGS1Qt+3fOp58aiKcyFq
lzwp/kYYbgbF0DvnRFEdwXd+u2gI6n8nzv0l9e6yzMR4vudug9+RsRFxV4LIjyAzxn69V3c7/haz
BKsAmc+mBhzCmCt8B4VOUvs5/tggUbZRZIXMdtX9IUc4UgjydDvszKGoQTffQpGxSRNVusDWF07u
djAV2luxqDhh07dEJtGW1pTxMRfSDfURjFpWHSqE4WfvKVStJfLnGey5fSehQ0DXPgHCYc0FzSPC
QaP0yhkztPdS+kQFwadKd6OSTdIqAQ/GzZXskf1ClQWaxNdOfwyvHJ88t59OpYA5J6CRxl3Vz6Zb
ae1/y5E4W/HIxpxt/p6o2OzsdKA4ROYiBXoK83HHXzyS5sSvWr+97zxeVt1boJbvFN6DefDkPg/1
xtxdkRU3+EjedoLTRIXGOJB5TrIR1+ELCmct+/WvX98LyDwtCuFR6sDM17DZs5ImORi3U4xbh+Hi
FtshBVoGgG4eH66OcYm46j118jr8Sk5J1V/WYbKt9+M+0gR/p5XO55o3FCx4oaH7ta/K8MpqXGfI
Y1/rAbJSKdibR3Jpnt5WnN40QET5GAy01W8bS7KwGH/V0Vl8qNt1+hI4MvmJqUgXIq4ZeYlY5fR6
KpHA12P6HmXCukqYqHF9VUNZ5rOncuzoR+QGwt+DL+h2tR430rZxHRpqR/u59Jfbm1WHprHn1pct
BAY0o+G3g2xVJKiMQ97hMcp98ed/p/Mx31QlLmq+lJUT4oUd12es4nKXC4VN99S8v/pilJJGdd9C
knGTVtDYD5p70WCsz7RGaR7TwFzTA6mx61C4GBpRZ+M23Zia5dfEg2wES8gNBkPQRkTfPWS/T637
A67/DCviKJ7TIqyFtyQqmoW/1w0uq36mE1Qb1bpjm6g37ZcCwkxMBKpPd3/mgpddPZnKpMQrmcz7
CH1ce1hNjgxdJ96I22wOfHZd/VXWW/x6kUJx4kcEAevGavFDYNLmpnoscttkaEqM3bDrYGeldWoF
TMwb5zJTgjNErYiW6Mlv82jprXPKa5Ifqbrc/0jIsVc8goxWMZmFTTklZBZielzkCi7He4Gd9Ldi
CVKeGrnUWePeTyUkr/wn3bFpszjT9uqkpxlSkPMCpWf4xoqOUW7uhUFE17R9mGz6mDtQPe3PsOEv
h0Ir6YM/9WvuY8EypjH4KlSwWvU2AmJ4tY9Gism6xjF++MzEEYUjPOO3ptBgCQ7xJEUWXQ0H+QRn
nZylbRCvIph2BfpE6hgu/iNn6cC4l/8vkIB2fSerebrElSIZfzAZUys02SHM7A7UQ5lcgKoTLYDL
6YL1McCWgyQbuknodwCu40fKC/48pFsiUXsqx4WmqhL6My/1xXTtCElgVggVDRBcOXVrAmY/VKmu
Rggy47ORnn2m8dJZU1L02ZlVLXGXtj2QpJkZ/1B0L9okr1NYVQCefEKliXqlsu9X+Nn9as8nE316
x0hMxtIOrBfYAnYQY4tOURJ2CjFxefVp/i0st2Mp2O1vdOB93XPugRFazbj+cuLjdfkM8r9gzUot
wZWaRUBLrnzvNIdO83/C+ZPFi1Lgz+NCUX6Pvw4cu9mm7X84cucbfJnMCcDZJed0lHNrlhSClutm
TCitMUHgl0eHqLgk2wc98PvFyKbc4oaKlU8a1D3nHgf1K/JPXOeBFYXZ29FukLo9Jaco4JdYNRe5
0RlvQMKxxO5NAt2izXYx3IzxELO3zMVxocuAMfJ0wOrxuA1UZjo4vpKUewMSsESGgejVmPZsq/hg
GW2GJ2j/pMXiLfluljmcPZSc27JXaC1KtWdHuZYOoGTH57SdV5qjOKk0aM+0DtF88+mT34i+L9Ru
3P0ilz7PSdBefXdqIxdW2r7LDcS8cuBge4HiUbvoHSoujxL2wC+1w6xHnvclaGP8UcV6GWHwA60N
QbgQTiHqv/ERsHjcKVIQp/H/l6GBO4g6suOfkn+egrT5AqRFvVVfJIIq7NHPcWvmukDlzoIkA9e2
doYSRgU5gc45L1Nq3XM2grOA+p168T6lD2WK6lNIRSyLu6kR5PJGRFhoEnTQAY+hWGqlkYreYpFc
EHRRbHGYjBuilVFOqWhowh+sBKVnyz5yXYuQDIPg1OJoAtu98EAKeT4M8sTh6wZr3RV7gbO6OkUT
9M6UsBXa9ml/ylFRqRHnnINMKPiOxTCzUDI3KAwga/k0jg2D+5l0yVP6LpKxBIeB1uifUc1DW4Nt
UxV5Ha4ECN1cJ5TzdLT9HMbBlwKMfdcxW5xL04IrMuooP0kl7R7y9V7jdhhijWxx4SjbrWlygEBD
u25UHzMfW+26lzcZvbyB1GHWntHeDsllJs8XIWvGDRezs/2UqpABdfrDURX7TkRqQIA7/obqV8X2
Fl9XiC5nis7+a0FSAvMSlmzRLzXWfYRMwI2oFDpVQttJrjqNKYibX5+gjCqbtllSzbL7+gFu1NgI
GFwuylWuUno5DG6aFbWjsg8x8aAVU+7LBHmoTu4KUpcEP8GrWKNkLit9EGLHXYwWgkPwvXp03/6s
QlbuhgS1wl40pup3HlyvU3uv8kC6ydnDWNIgh6GzMEPYvRRTO40TqY151ybw9rVzjl6/aduRwkcr
ZIqeXa+nsp1lZAC3ki0ep6ZsT2EQULPD7K0bMzjZA07nXTG8kag2qoriUsJMlNdyi5i8OjOo1AUw
KZv+mNpvs+0QKYR2ib0hKiEvJYxdVk0VuNkmf2sIw6AQqIUXPlWUWq3E/FKCvWye6niXKk4qsqtr
YZFE5pHbpunaqq+wzEhYSOIk3FGlSimbWDP03RnYD+J3887K6sGfDEFvKEJXj4VNTuvQq1i7fB9i
w2L1gVDdh+bsu7B36ighHr8ipIa8OqHeb+JxC2b3d/xyB6Zmel/e1krBEMZo5gzHotC8YelpiPMe
uXCnr9JtVumugnrANPhcPf1lJKlqImfjtin19rnPzc5cFlN5XlPYQczJ2QHfO6ddNXkMYakiVVCg
Ia49WMmSQGKtW5ohbFRUFeS/YDxozUmHWkXGMGGk/4ANbYo9Bwt2DHFQQ3gpy9VcnrzGlHPSi8MF
a35fb2rNsNlZd7EtDnIl1IYGOU3lji8HP0Z5+74N2Bdf2Vhuo/xbGD3Oj6RNxVDDm+TkJdI+JyL2
9R8NZfMcZ0jd03lZaNF+uXbvOekISKkRgXfW/QplptGM/4BgwuWEJ3VIH8vAK4qVwAYlY0LWV6AP
+yVdrbD6aCfMBR2S4edKWohA4JtfJfAeY0xfZeRvjmpygoIKvzqwh1gsDSU8MvCxRW1BhRmx8K49
I7I8UJHosbqL0Yv5z7kOUwnYYMV9w2wEkcNeZNtSW1bypz2p7neiYGSnEUuBpgr8TKePaA9zy6Df
TvazE74JB8npTKVWxcuZMNJYYrDEmNTZ94VJGlxTZjWoe9O+LsQCmNvE38NscZJh9nwQlZbWHnyY
Azx6eCnnfpQAlSNz5/7cZLrnPFLnDHLnq7K81E23OB9q2j0AUs9aMWZrstVchAH62+t1Lu1qE85n
TxjBp9nqn9n5WieEguLfCJ6K1X6NoBuBVyAc0tvEW35idk6dR5i9Mru8vtobJgIET8Zy2+FNA5gS
uLc6wAXgejEuRpgAZwHaUvNRLzMhkcPQDOnFvgKVKKE0Yc6n2d2hMZ8nrVJcTQVDWJyz9ZwTWpIc
jFmr2aIgN40Uxxf+oXFVbsiTOCTIhSDQr7mixohhu43t9VhIgHYvuYzLC7hkqfO9uviaU+Wh8q95
7/fBf/IHLeaBoemncjluyvcC0uL0ro8yWQ6orrbQeoDKGUoqyvctH4M1TJRB42DyKkIUTTfjkRpZ
Lfqgp0jRKgTFFEcQnYyKRsIHYiaugLTzwfHI2zsWEsWY4DOXSIcULhWN3AT2vZjdpz82PMz5wo+e
IN0jEtdnuCKvmZWA5PJ03gZ2Ajk8IroD8XrwhR3mawJGkgRCNfD3Ww4LfQz0RH06/g2qtXDid/ai
UB2cKJNt7H3UKDLtXpfbCpWPquigyyF12LKJvPRGAtvhUkzHg1z01M0fxZIoxtwY4Ty+IT+OW9PK
RO/bnTBF+NnrJi6ST+5ZQss+deFgmveacysV+rGUwVxvldhbis5l9eTPvLZH1QbdNPJk9lyGDxXX
mSoATFrRlrpfR+3yBPKTqsXujcd7doaxXDEbIPqFdbv1zWnxlTV1DmP3wyGEqzpjRyEULN0cgQJ7
wG1ygfFClvjGcVETSBN6YBCaeiGlFqeC4iLupAQU/0lx/1kzun5XgRFYwUvs5dVG1BXZRDpbcWw8
6EgiRkXc6Z8WIWmWVcUredFx+WqaKjV4TFh12P98/dz++UcGXWYkROcZ68C+J/OnLz9j0w42stA4
drqWMLFmGIkpp+08cWYM8Jd4VWH+H/yErqKNP3M8FuyUC0gvOaDCXORoTv1Y4nZfpltGMDfxLeCb
JMjXrDoEuBe8m1GOZ3YHkWqSe3ZaHNsCBlc1zgilJm6JIEJlp+yaPeZN/S3xgkLSm/nyumm1IgZl
eL0fhvfpbsnu1CsRWEbVjqUwwvAH/8sPX7xPuGl4PpOVZo64uWrXUCmAqvQKajcu9FSOYqPkshg+
qgK66xSmriOdagKNiH3oyaFu0noEOiEAsXJ1HoILB96pmdsEQ2zpFmicMVWyMvjnvXF8BLc7C0Ko
RcXRXuC0AooVwiKcl6wOul9l+GWWqVOAoaLnFtXK7cwItr8jEFklPqRHqwXyBKLRjP8WThGnH1FV
VZOgngOb1dsNjUPUGgmBO23qyrze9az9RFQ6HuCxyMGdUmnAXXMu2R4IsIrkzpYJuXya90crluT9
0BQKb3G+NeX2c9mjbkuAviBiuVoK4ZVVJn5qKYzPsDCg56FmgCslVfv01G6Sd+rxwCH4vG5L8g3m
tTzpd8gl+is/BDgGaXwk0ciP0oVcynuHk9agaaSRCENYJo70Ezcid9HRiBM9nUg6eGv7tn+sICOV
And1IA2AismdfY45ohilJAoa0EXLqMEBGUvpKejosM4ufzJ5acZFI8e4zwuFg7pgkcFpx4fKFvo+
47sepHCckluCYcEPLoy9oJbCUiqa1VuyxQ53hN/oBattPFcNOaNaHlKi4lSjk3tMjfJBCAsnqE0s
HEbsw0+U56QG3+PelpADGqRKXMlRIPHmIy/1qVbEFdo1lzHL59TMOifaM1jWH8EuEcGRNgyZGF2U
p8UbV8ByJTFS0OWUQxWIQn9Vmr8hhNa0ZfOx9kL00SM9PsK3b8wUqh7LBe5X/TrKaRy/gpLEThqP
/36VfkDAkPIq+L/XkBz84NjbX8eJKqUtZzvtvNJCGoBHsiyqW5RfsnQSSKavNvOtxvF4B7aE30jE
XWuHSyqYXnOLypA+0z29HuTeRtRTJkI0oNPi8PxTnhB1RiFBLkcDGjnA/Zh168pcmmnQS7PqCEF8
EZYYRb5qKvp5qSEE7UlMRf+93/OQVSWgWrsoBuWlguszCIKXvhSsOKh5eKIK0kbTjb1VVaO5h8R3
PxibwlZ1X2wUBzJjpM0Uy0JG5IdnEAfKcdw8ot0QuPNl2onPe2Yononlbq+sgSYPgW5agHoh4MzK
YZ6fvFTwVnCcDHMrzstOslBW+yylqGxcZJ+HRK02ex5pIrpwEooHOTCYWmfO93E91gkzphDwt5oT
qDvQIdbjyp920tE/JPKL4ruaemG5/6/82aOAgu6hYUNT/7K7HUsSc3mMFJCQ7H6EsDhkYF4g5SnC
bJnQrY8uqdT6F0SSFCIxSmkR8V2n2AJYIZ5s4COV3we0p3qI9+t/HmYD9h+cUNueZsrw38s43Ihk
jGdvUS1I7Fba3lkDFpSScVs8j53AQomAqPax/4i2XtQri70gSAzf62hI0/bDcP6JorjHX3a4Wjnh
tqxAFaEVS5f49gF9mKq7v+9pOBnTLRxeXdiQKHswOGRcIDZcgbRhFcoXaihPxLhwM0MxXcPBfXzs
aTAhzVXr/KXQhsgOgrkrgOOLUcnKLfuc4/egrY1qwj+u/PNoBBn4qkcesOV2nGfbpxddCz7kp/tL
KcEANJIiAyLngeDCp4qLNYU0UxPd4fC0GoPLClCVHSjmKUyrrOns6+ASpGMvQuM0+90AvfwBubP2
ZdlRVAPUiZzdviHVbMtUa6QuXA+nVHBinjiS7Yf1pmW61BNbAQzaImyMq2h+v7mvXZZ/bRhCtkL9
h4hBjGLhuQqtvzKsFVQzMO9dSx6uNmYcKwcH3j5UWFMZfu9uhMz8FjuT3GBc2bDHlFgE84ZG3K33
D0T5tumIe827FPwNaQEebiKSLo7Ilcw2ozbvn0tKu6ZL1DvsTbshk7psKXupPpo4AzuQ6yCxgp1Y
WE7DjwC+q12GT1boPzw5UCVZ8cOUshQgSV4fz3qQvms5CnwG6ySfrxcu2CjJGyADvZ9aWVkUkRDU
jFCmNjmWtOlsir2Yqs1uuPb6Piek/VFnGXiKohnRlVcS/HkihXZL3/29STJUQ1wUe18J0uDLdiDr
B+aahpvEQFHtKmjq462yXkJJ6wkDntsY2+vvQntNA8L4xrd/0wcUu/zRWyADS8rvRgmp6y066eia
1zp1gDJ5l+BlYtwlcPw72w5JFFePLWmEkGH+WPpNvcVDkPRyuRHqKtpVNZk5wrvDJxf6990ilJ1+
mfwg0/TJqYdp+S22kLx+JBNxb3x7f1Ro0/onUhyuVi8J5ssRIjuroLttYSuG4IroTHQ+q2pjp1Dw
I4XdtAw99ZsX5XeBgXkpBztz3Coxun2Az/FtO1tyCEQztNYN+B1GCJ7yzyRMbJvM5IudJ00JlXew
+Qo9gNJ8XdSuUSuMVZWZ6q6LC+TMzV5W1F+HDMeqvK8k10BZzY1PQhfFCDUg3ayr2MU8AbhPUCQF
vObLhb1c9Y/4fYZLJdmJL/uEmFiKKBtbsiKhcf90ShRwwbvuFwlpDFO4LrtxDQ5fYGFDnDfcOlWc
IOWU1b1WXxRZ0MFL5yex8Zk4P28IYTjjCnu36jU94bPygJ5vhBxP/C2FwmocUO5HPaqKAT5ikp9x
3L5+3/Tph4IzjskGecimSqITQrZrVp7gYFI5jSO/IYtNm/ZDPAhqgLaV73va6gH+H8iVEKuSlSM8
TTx7EzUJyaSE04Bj2jmx7hzEy8r0bybrS+4K+Y6O05PfuSmvds0k7hQOuyQ1xu/fQ1COkAraptOj
YsTWO43xGjkXooX+fDKakBGo1ZCahf3dC36miTYd0Ufp2cWq4vqKlcALkn/ehru/a7yeV6Nfu2xz
kEk+sQUo1okTP7F7ccppGOESIwEmabGngkRK8KtM95U8xVqXNcmIHvNY2YAAGOU3Pn6rLYLkNher
vimol4F9xwSiVMnJJdrwkGxUxwk8MWdqFVIxEG+ZSSkZXVxWpXW4vcWSv3awELQTuol+uz6HX48B
w5NJgeNZkqBqyLCz3lL2G+kDV6wmQopXqX/9N6zUGI4iJhp6X+wxFyEt6CEMnj+nPyhUcPekWTJ7
RKSmY/QgDP/pmGz6934zp1TQEZHiVLHA+7nwOwKxLXAaRyDOdJItPk5pPrXQE4uwTL2QWEXRd6pn
ALu3uwwIeNx95v18q4X60po1+lvw94G0lxiqyUHPbuq/adEuR37lhC8toBx32U18JFwgOLjl7/xA
+QC76XFPu8tfHhTyJleE5WBRZAPLGQgFHUrUsp5F6yBKhz60SyZ4T5nBhaBHrP1SzsDht8Xur1d9
t0/wKdz9vFONjtXXprQn9VCZpB40yWUTNrMjzpoonYfImAMWUiHCgc+lTfjOlAK0or5du05ZesnQ
8rhVKR6BkHV0yg3GBbbd3L68ChJLWKfKdkU2fuJNi8UJ4hVgL8+XT8W0zPDWQMnPqtFNOLFsqIpk
k69HJZtnEPVZzcPbNaWTzjD6irBRlpULS+ZFKIxGdsOjlix6/PK8KpvJ7GCIl61UbalUglf7LCrx
Mvp93mNN86eN+jzHqbgkUkPqTHrygo4lu/UjWCpXxZS15vQj9Kvst02sDusnd5KwHwJWcShXEurY
2e35m/3dmYCyvc7+GhmVCBu2QkD8NoplVdWiy/hV/1u1AuW0MlmmqfvpfSAF/XJG8zsijVk6tZuV
HOXAAhHhSNROT5uR9V2Qc2CwcwoJryd3MpBwKhEwQgxF5LCpZPK459gAmQLEZM5ml/LLWY3IOfQq
KqA9BCx+U+cTmZMp//MTaL/vGKQE3kljfC//k7DgULG7Anqa3SXkv+MBYSvrZEX58K2q8KzegsGM
44RHs+/0SgB0PaQ87Ozmsw37c0j1lzmg4x097p/kg7UjP3kALLWO5DqhZr8nztsHghB/b4ZO4gIG
9F2BQIOjhmH+oC4Vy3w0uf3qow547uNQCl/qoBBspRCosUvTtcoW9FlkfmVGRvt1ldTJ/mVx1PjR
amK/WPO2MXAh/p5lcmdZJSwYNpDtYsFbQ/j1GyV0qOs/7pHOSCOpqI+SHQ2P/uapavnkD+xxuQXh
DrvxjTBZ0hTWvGHtxBTZ3ugwnCXXtZbUnXcm6i34zZ/NsMFckR3OvDMgX5Bky27rHfi1BNrnj+R8
u05jMR1xpwdllCEfiyvuSg49vtc2IR+SdKuZI0A+9FX8eqUXolCweW4o/i88snRzaJdIpTKeAydg
eGhv0P+T5qsDFYOp0Yf8EwJUdkRNJHx8hp8AKuisnHlpHKfMuchwqaKJHTYDvnLV4r5fxioIyYQ6
dqUjmZfORCBYJKz7eHNEdqZpe7FZO77sQ1evKfStPWyboa0D56jVLsnvlm1Ek6LozznxRASz2g5g
eVcaIrZ4vpFI2n16bGcKnMB48Bid0hCR/GRIBabCKZHXbDoHpeMz4qPDqxgk2dFJuopzyW9DA39c
8aGO0SARdvNjetxrOKU0oHgXL5yWdNnAbORjNzgMfBvba5Agq2WXzinW28EgN0Jk/sPuA1t654EK
t0n8oJ/IZCqmVCPcojc+BI1UqmGDEYzdx3QfJZc6C7tNCq481TmGKoVuUmja3iYhz0DwtdDtGfdu
M8G9UADgAny5E6A104TdHSvfwwMU0cdwxemaGtY/P7yvht3r+ehykh8xxB5MmdkOyjmWxXurWg0q
ty0JdGXHc3McmKbOsCS4N7MUfv5gCDincxnlDcDEpxKBmwC97YDFnh9eEvWTtD/39jN0X9IqS9N1
Wbmy5qR8nQFjE7HIJZ43xXFVf4Au17tw/hf/dxtfKrRD7N0ZGcSvbO91WMUtCEMqG9gba6NIFpKu
loVJiLXB5mQBaoJZKdbQamFs84+7472YLTNusTj/mXHhqMMMbfNaiatNKxJ+GVh8TV819mhWRSTZ
ven2MLpqjMYYxc3f69R5RwyLwN9aQpI+XxKmvYybohw3cebiGViPWikrtZRn16SjS7Eclk5Reqsl
kHTFRMk6X6XeUpkhHa/iqfPtUxNasIrQV80aHtYCyluqQyiAv21mw3thStAQt0ZkAsSkznFHm3DT
1xYZ0mNq82kAyide+Og/22GeFWok0jz4O1raGNQZ0T2KNk9XQwuhHmoXea15JVp5s5FtS8paMvy6
YbQkAtZSBfF2CJaBl+KIYZuFWDYXKH5DYZEYAyKivO7nzWLSZHUPIeUSOGzzyHSxziAFQmnzmxN6
AMGh7uOUzpHp6l5b5Taqs4Dp9QcX+TbM+VHvRzsBnudrBuPaxWoarPL9rrppS615UzwNlvi9miyw
XjTk/pb0y/iHLrwjKzILqZobuSn67CrGOmPI35/GthG8lotSUbzUjF7lysCkwON09B5fkxv0q4ap
MCKoMkjChEcsO54iM6dPuIzqkWgXFnCCWxktfXu2iDKlJbxRULYnpe12TnsyN2RvqZ50lgAurnFw
YK4tlP8SlkIHB8wcpap2kguMvSCqVO+ozHW7xDaAKSkc7mKy/TXog/Ke56XyAWBIzb2VsTlNwNSS
nAJ9qLsCm8j/NFDvjR+rjrtGSvKfbpAGE7STXTvzL7Orqj0AFvqlXhS1eiHieSF5ApbVTbE7ol2C
p6nO+unxXeyKgqYyZWyCltHRHN8LqMLhOAae9D6I0uzXR5ZWuhLDqi28VGcYnHJ8YDojXTAAMdXH
LMcrQGWBRpAR/9e5LDRb19jtX1aCHd3z8iXGOvXG3kmpMKjiyjmC4CiS2T0C6C7QXPrUfOeKF/LX
lzwPDjDdwIIju+9Cy7TTSN9/aizVlxj+Ht1jPAn82lkp+KG6uTdmNdvHCJrZZFfbhS8jutb06VHi
eC7koemLpodSkyrGeWRGfD6C8r0L+N1wst4H+EoqDaMfBuI88fdnj0AX3m4I6tSGNc4rv3PbFhU5
r/FNdVqXqfuxFyGInAb/fUqtFUcJDEwtLBV73PhMmcff7dhtHbWdCaNB+GNzn5UuZ7r9hUwU9d/j
j8WRfD051Rt87Hb8pPfb+Cg2helwkTyqwn/KEDq76EKjDrc5w0/cTwCoJt+DUjskdyIUarxipcYI
dNESQ4+QCJky68iOF7Qzf8sjvO8LKLt67eACFb0oEfoG4X7QVsfOl8r+fBVUVTOnMnYX7uvjJAzV
239uP9EYP87xNoSIOJRTfGgvsnnzzstzFdgt/fuwhBiBytpVKTTtycLvjFeX0+M3l+OxPmHTNLsB
nxDCgiuMmMXkKtAlLde3es+A/4xlUzQWJG+c67IAmdujz1dpa89CJSnyOrQfthMviIjlW+R2DEk8
aitogY1ysJo44WezExD1CUhX0kf5n0BcG8juno882UBk3eGktbFg3pm3tx4jD401tdRc7YuJ4fQq
sIurlcT4xANu4xVxh/MkxcY3giGOW3ryWl6Rf1xTAgI4KBsCN8RmYeenhxia84yY5yyKy8sUbIBk
+aAe+8Zjm11ch7AvZI1lArg+GnJG7dF3y7Rx/K1Tkehy0MMD+NPSXPqkv20k6Nmc/pot5vukM0tD
NfaHp7/fJFkC+qd1JwNvoFWNFMXqGBo6VTZOt4sQ33TZdmO+Hw811DkKtK35prLKPFZbvkpMVzVL
i2wWbuZV+Y5yzrazQ23497hZPrywyXfYI23w1C/oDsdT22nukYSjXK/TWrV60Oz5dtY7SYRZ2SXH
NFuH1VLrzKCByM+fHm2YejWRvRHX1rz62YuFdFBGKrg+sq/cABZXRWxMkgwipo3oe4DOrdoteRQ1
FkwHKeo0IrDbJ2KQcWraZqB/ufsyVjeOk3tJcievgb6g8myhTuQQksvEvNp8EBP50+zFujBBKF/+
MHWaR0NmhluXUVKpo8+jwUomT4BYwRj1pvlBjLNW2XKOWQ0EUlzKugBcKVzP983yMLBR6sCYlDit
bGxbHe16Fh5ozPHhIcbIv5kbD0BWZpRSKnvFHfdXdmjUUenuMYnvkJKwL7+PnqhOr9V2Wn9LL3ym
rWA/+2xU0sqDtwjAakCajvv9mnQXs3xylda+kFZ5KK8EscS9uWK3XsxKcjMvka5QWOcnW2VmZ2it
4oU/Di1IFTc+dNlWpWYJ/D2rnZgNwPZvz0kMNcgnsnSI7TQqgHgMXmD3FNqKm8cB5D61OANYw+bK
DeI+1/OV6i2FEuH1ZZl9l1ILqZSlALmjkVsd78wXEXv+8GGX9jZR63BwbhonZoV5+GpfgRlS18iV
GqYmIuxLG4aZ7NFQo4G/TGf78nz6nCbt4WiejGe+/8jzV3cjs7Vy7YOqilj7vL7blWFav9ZnIWgY
5RH6euqSUl5YDr0Cn95AD6ZXw8CInld8+fLRdl11WsSePctviw4059YHbjm8Mr3eJpXiqlIsAL/W
m2VvnVanj0oDaW0pKhiFNN0ap4GqyunihQ6yPpWJFfRrXat2o126Hk5Q9GrQZo6a4nAqQRMLrgAU
3t2e+vF9hfygPEpT/0yVMa6JAhn9IRf9G7N45ZJ1RjcaXZ92SFM30ihiriFvXoZHUKpym1U/QOzQ
ucv/7aLZ56kZ+9mmkvBn5sKZqjhWGj9hmCV7UEsOsOrDpbK/a1fu77LAntprXuR0Wg5dmyn0fL0+
jpNtHlLczPRfJfIvVlDA6OVoely7NhowNKtmjuiltSNIRGGENLnxbS1VXBp48QkuX9w6KZCL6QBN
AOuOWJT03AAXnNSGSrJV+ppWzoxdlMemkV1ZOiO/KaCP7YJUzrdmoLiDUboc/q4isfhssGBlCYSZ
IRsQb567aFmwDxPdT2m3m155NuhshH+yuSxKZ1hhIJHl3CfDlwJRtdbSrlsyko3LksHh2JoSKkPB
XK0QeOr0KbEIeygorZ0KlDt7Vet+ELa/4wHR8WcWJuZFs/u42XJnJBdBDY+Ma7gv9bCM7PUx0ybw
Iapkp4778i7x4k4BobyqV/8HHdA1+7iSALiTItPu4+pQ2Z0kcw7nl09fgVUcaYiYC07e33TVyUMu
pqCGnN3WDckx9wRDCnxaJhvVYXBIJil206l6ap1aMmPQW35EiQWTV9FM41EvO3jDx/A18U8jalmV
q4kbpENzaVuzd5v0f4xm+Ltrti8Oa00a4miEGF5gZCsgXQqSDcXSHCpcWazHl8dj/YW7ikoOc5fa
6umnH7M94t0uIZ+2yejDDfD8j5zh2IjP16w/1U3nlSWG+FhdWLPsIjkhmy1ajYaIPYRD58QArw2I
pUIcCya2l6z3GqZrT6aPuBAdJCERJHgcxjN61k+3wQZi/1wzRdxwwjJxdRtM9x8x3DPcXeG4sR2T
7x3E0GKzMsOTka4ub8iBKRqh++dCiwRNjlavlowXfRkrLEW/3dUuzknm3luLs2/ikMparLGJTxE4
kTQzqq86V2F2CyEbRCX6IhCnFYpPbMnZXgfwhemFG5/9zawaiW5rC6MtvgzH7j8M12WiaLicGqAr
/DdBeDRZsKqzXmee6tdJ1958qjud9a9kbRe8SF4i+z0rkOz4XaItwPOXuNoQOCyA8gLAmx+f82fc
5g6lBmwt765Q7enYn5fLJgyWSmu9hSyhEu3BElsdQEBx8vYBH9P7dWw+o2poOWAC1jVFDKMe86xn
5JXXaSoacEBn129kgbFewZlNBIx2PwADW6XqN558JZtmklgyF5fKua1oXNKh/kJQotvbpahzzhNa
eSGWzsIM60QCmFg0cOH1a30nG4YYlHp7X68vP6676Zp9Iqhxfubp69ITpwbe+WS0vNo7nAzrNQ67
oEo+MC0hOupf1dCI0ggcqZu/L8aSY5uP+1dAl8nKCHFts66pMBQsjhf97KxVIAN4m1OLTw2uOPfZ
+oPA7gjsAjcOQdmcBxgj+NbtbTTW/9sxSkgZiEA9SC1nepqvEapFv69WyBAVv/IQEfI4T3XAgh9W
+Vlrq3IuE39+/1kOCtVltXne7oVtDlCMiPESTuV3CKNSzQTkJ8xMqG+RegE6FsEaft4hDwGzwO01
CBRyQ0e1ID3OpETY4sYamulsc26u5N1CXKdIiWHxRnCXHlaYMLailwKyCknLvkG57ioPjVywlZsz
15QA0gT9M8F36XjDQwV1s/BmVE/jO02u6zGbuCc+ayCpmoODyb2gTrmm52ZBCqKN69309X8H3HBx
itvlVv8BKNrZHHhPb9AhGqmy6E6rLT73+ddVLQN8fa1aep2ZqbFqE4DLuzo/ExP9p7k3SDZt+s/q
Ppl/YkZ+0Q9dezOY7ec6ZS5iXGwCj41lQr55b61EURIf0IIj9qkjTHtuRFmtKLifOSUgemj0M7o9
Khwsf/JqBq/Xk5DwV9t8nWqJpYm4Q9NcBFfa6Lley7qsiWT5J9xQj300LuvIDk4mwq8IzOn8ORpV
ZvHWmZPc0VeL8ZwyxdIh2j6oFcju273/vdKs5RIZ9WXT8Zo1r4fFqjTrJoqkXE9T+3uuiip3M23v
yTjIUrT6ds+OZCs4Z7VHwiQDVMKkD2RwulP8LoOFu/jg5Sq1Pxp2tCPXRAjX6+1xKgPx6kmjrZIH
7v6eulTHzxkkJIEt9pbk3i8G0oE6TMGRv/sWKnTo/BXcsfKIhTTcUMUFGE217OSPkiVUTKi0u6mP
cZ/vQ+1bHUZIrtIOsgl057ayJdbWHd1bWIIHL2PjJa6As47If30++MTp6wqywFoJ4RhInRy4qtXE
cbJdnD3uEN8UyLSFM0lFHWOwqbKHBbA0qZ4QneXK+W1KJc1AcgmTGyXy9lDOnYx7sz3oFBnwtJlZ
Z3SCLsw8uL56KJnfbATnt3Vlfy+g5p9YQ60enpvcF2nrpaIShA4vZsxEjGXx/Qlq3EBddd5BEiPg
D/s7G+u6I3obGjdOieywU+8J3F0APikva1gcf+S7ypem0+U+2tTgDWJ1YNXhQ1E0wjpKgwPVq/Nr
t225nW1GLgszOC8EjRXTGVCVA1eczSawAi64f2zieQVD6xlVQoZNENqNY+KG5Wa9pn8z8CppCEFi
k5Ghgfu3fT1gy03O7FSosGRPla2Bns5Czx2V1shg81J6TkJeMFRhVtb75p73uuT0EMpVtnct7BrR
46qBG4oaPKsHSjWTOdFc2GWnRUR1w1mX5VMShz8KV5nCb6nUdv6vDi4AIQTiL6fQTlyohn48sDQC
MRJNfnJ/D3qYyhz6VQM4A2idWbeVCUC7LAJ45wXzd4jvBSEdIfqvLskZ+fNRebwABcvsKk/4hhIA
/hTV4A+wHOp5wHtzFwxBXNXN9d9HM4kzbkI2x0f7eFlwS04kLXMJindhgz8kUTSV4vmPvWbBz08E
2j0aPNAlQloqrso7LufcP9VFc+xFgKKjT8JNVssZRjwvKuaFxN8hurJkb9CoL0ClfTJabw9IbOaG
lmZ+EKY3B78+AXaKq5ayNv33TjufXlq7QAgmXJZWSyJ62ykcdy4NH5kbC3B+lVPRLZX9/MN/jlU7
8Ei6U9sCN3PCwVeHx1M9jd8cZ0U1G9NFlOf7ofbo2a6k1OwbE1q1PZroTHBGsNE8F5X3/IUhK/UM
/5wQe5eHn4hfqh63JfdCLbAO+gAHC7jmhDLqTCjvtwh/jnhEXsXQNBNxvGLet9yzzQ72WT3HHgCA
w07XOPI33rxx20rl9XxCi9A5g0p35/glml2xc3HuIxNwd0aKtAS4bEI7E/MPaipauGMViIqEO9Qi
sQhETKFVjmajeaRbr9F6Sl5b73rZIwyFW9SBGSqZCbueu7WKUMdvM0s7kOI25vaHioZTFk/GS+Yi
LkMgS1jGtFPLH/3TaVJStgvHrYP4c8hxyiyOzdBXu99ZcXkgx14fDV6wXxuKf6p/Z4q6Z0WGfFH+
vEb1oAj3MNmB1ZJl0y6tUNQb0Rhj8caW+Cuf+fN4pR3umA8Bkj9/BMlPV1XgAgh1BuxkGY6Bs/8l
9n54nm3drsaCNZqCTSSa7GYq/ad+/16qxr2JkrLYDFMsyhizV3RAuOFj1ctSCi2wcH/K2xIyun5e
AcnODUgBPv1bybZTK02R3I0JtfKvggxmSOgnOJGjKfoANKWeGrjKlJtChJTKWeX7xRBmMK3lkJiz
Mmt8/rB/KP50uossU+ZGpAAFqwL5JCj05gRcjQR7PJLWd7rZPRWi0gSMYHpqS1rw2dik4BUjeQ2m
A0grEtSwD/drvfRMl2ZeOM6k9catCL5IZSGrwD5GSWkFWLEsYR7SQfBWEH6zw8VpzqHIflyDiUbA
1USRLJIBjs/D2fU2ackCQ40igJBwq8dH8oPSBRpfNkTS9CjLqs0nEgz6nADNva9Pna37TEO+nW3H
Ox9eZsUhPPBnBJQ/GV1xjBZAoWE8PM8nYUHA3aOdI7rqJ42qL5U6sgMAOyENJy+ogibxJntLMjJD
lD97zn1rZrNFP8ftY+avWnW3IHdw7CsijFQdHvxZDAUyMdEPwauUKolry6wM+57K+J/aG7Z32fY5
AZdN2BBM+4NGlJU5m6hEe/q5fyeNvn/DtmUMMJB7oMb62lAGiS4CJBC75NBUzebvC5bUJD7gEqlH
jFSFJ6KC9BTT2MPczn6S1bjGLib/aCAEjkXB89dQnYkWjbwcfUUxG1696e2JqKTra3ur246C+1UM
bQtXYm+wzKBSjqszcdV17GPaLjD3IrH7QIZcH4YqY6NbHCBtwWnQzd8e738Tn5ixUqonlM2YUM+C
rgJvBxtRh7Rl8Cmy66LIJrg0HJ0+hvBKC2MVcUb2/N+Fyc+iPcw3AfAuQK5ob8IA0FfUseXOkWcl
fG9fdrXo+b/vof4ovyO9z9mlX5fIgdsd/zXb7lOx4W9ntW2f0ryeHGofGoPiLt+Bu/6HDqkFTk6i
z96s754P/nhv32vI1czPyqG5WHtQrff+KP8eRwleK6Qxmpl/4vB0AfQ5h4zf3ILvbC69VyfyJ5XH
Wize2Q52QlHczjpPykA8qZN80hnJg4HU69grplNaY8NA4ZdzzXr0/FVIXijRNVH//APdKiChWkgG
qzeRb47rNAs8vabUy3u4IKyXN8UeBhu46Lc1INg9XhkhAmcAs4ZtH54C/ziVWVwrvIvm8XMiGot1
T1dWUwMhy4jca6dZ7s6HO9pZGHavTGFPJEM9DvnhRQeFJrnZYi8gcQer+FQSRkpe6Mj+Lhi8nrXN
Xy26JYqMzab2JlL+HEnstt5MIFh+NwTYKe5nOQ1RuHKG8JJC1uWMbg4XdobT+qZtyLa6UNkPi2Ij
PE/iVy/T0nX1eNhVcyKMclR/JqFOPUbjBIa7YLGNL1jqT2Aq1Yo1ideGGJ4AigT/kbTTNATDF0D0
fqedC45dS3ziQ8x1STEeUXxt2RTFbxHLVx93ej1Ne+m3fGCgc/vptT6epycbIiK50W2Rq+MOI9Qv
X8wiVpur8TR/f9gn/bbmvJc6HCgvwu7hvQRds7+2wjMM7Mu5UCG/HU0kTdttis9QfbdyowWKzbRg
g5dWSjW2CQgLA9YWSgpHev70HcHlQtPJHuu1HSCCIqDCn+lzciPZn/l6wvzZolSjainxi/GcVRoi
0mykWHhnE2H6FmQz4o2WDUet39eQVOG7a/5It762fZMps3C1AMumWYkFZWRxvYzO4QuyQj4xUo8K
L62G2pxDLfEsMCr567L0SaM8gHLL4l7sPGf1SiEoWY+j+iO15IGYL5AzLoppKIsT4RFzGe/Lsips
Jn/OQsZ/TjW+0hqZ8ojWuonOptYQUJ9Eopuu26vw0FQcgNBrqNuvjFpSvG3bBhelrq1wyfAZiXbt
NLkC4SB8xJaDMrWsmQvfaCUvu/Awop5B7sOafbRkbej5fB9VGGa5INgcigeWUXGY/k+Mbf91pjtT
O1T2e7C7PFON00r8vYJlbXMG3rsc6uGMH+5z3No4Q66XYH1cV3+RVuMhWdySRoMI9zRbMZdn8ZV8
eVWjgcwH2UfYYv8ZJOXBVxh+eaDPfo1FsefUTywEA33HZ2c6r2P6IyiFb8QzBGR5jBO7J1flUk2U
iK54QxqkYXFKxBpOh40l4f4CRKl5C9N75CUXygpW9WzgUg6WWPo8EpssE/lbQWa3VluaX16LGxcE
HNCS+7D0k7Ts9xCy7V7mSif1gJNuuza1ptWQuPOQjL5LRTOzmCwvHYGB53A2+PfJ7+EsqUpx7fOW
xFuajQfAxD1BQxfigE4vW1yGmAHN0riRxkYkY+apFDF64hgiBPdflgc/5IfxVB5Y8/6DVzk2J0Ij
2dxEEb+1PtjQT4QaMbZmY3pENjKbQoe+2f1tJTOYXjjdRv+N7Ohb8ypDThy2f7Bm37GRniurSJbB
wid/B7nyBbIWlwFHhmz87eeYsSlhX4uPgW9b9HfeCSOP3X8n1efeDjJznP7nRY233xob1lKwjie2
xK6pGgyCJiChgaavAy5l5kt/dZIeHnhfgjnfbXrj0JiZW7sQKGt0wYGB6CI9LAwhkw2r8b4GtGpS
rp+2czTvJ67AIBVBYWfNk/8isqmu/bGEzJvQ4lbyxLOksF2eqa7amdy47ZOPr7Df1wKRFYTeSEvG
pdFjsmfNxkiseQlxO78AjUv9w6OpCXjtr2POym6m6Iw5eoYr4aF58ipi9WyhmxPwUO0guWm93x7a
6Bek5apHHMM35mWGWEGBWaN2aQDHB3z1ofnHN3UcjMuQf4pj/vHwhockK7ng4EN11zZtZxovh87P
u2kfUdQYOj+vqeCq38GC1fFyVFL0itrtX8j7EjfD8QYplqu+0BPUioyPO2Lrbh8uXznCHJJK3nNE
GT+/Klauxgpp66p1VZItVIk+tGX66bGCSNJd4eiGwxy1lpuovCsXhmwN4YEfU5RIdbgvL06yiemO
y1BDp2NaxwTmU7averStikHbK1llFpBzDohGUZQZxr3IRsdqVpR4fmznzWTqlvGI+DLEOHaeGMWD
FJ6VKDAT34wMFCAV2K/rgznXP2JcMLOhKnAtK9GkjS16cVA/i9u6BqLn+zUO+eqvj/bQEGn8UTEw
AV8pxWo/R6lrUz6iHjN/IlT6LQQH1fwWImujhKNYkHpQeDivLtjI8V+28Gp1J03rA2dxoWe+3UFt
zlXm1Ep48CckA2iRjyWhNHiwEAMaCT4Znwz6fUofltATLSL/HpkJG+GXsItDJY0wc3QATcAYydBZ
fdks5My/dkYASqixBFS4SS+ZIuv3QtlaHkP9T/K6OZCZuT45LMqT6EKy7G5/WmqTo7xS0v/LqsI7
V5+1evxVuvES6Z02tcMsH1OOscAQYJaNLAJaQp6ha0sboLO7Y+10X+6FVMPcutKFeabM9gX4+Gbz
iITWOgdMTPVJU5DVZbEOrmNHtiUzik/cAo+eAvpBAj3FXrNtQcAWMaP8QQ6FSsIY8+4m8kgmk/92
GhoCO3s23HHVdDtQgx4nf/vvh9OtcF9T6xNVaXUmq/PZEksHgnqGd0cSmTxdMKmGO3ti4FEXKi4e
vHc/HlvAT+97ILc+QjmjeZAxg33lvmwNTr9Jqh9bNhF3P2GtrRPpdu+HPu5a5W31WJyviDXf5Vy5
BEhtevLFB/3DOPKNmrG7fuxGeN2fa2wLtA5AcBcNRmR8dXDWNkW98nY9gNYoayNJsZfqO27xy4bP
7McSrm6xFrjfQyZ9xd2sv13m1UDgYDB1AE4fOkqBFxbu0cFL7kEFet3DaYoZyGaa6KqifLRIRclc
awVoWx27tNtRNuw9yMDNCZm0KHPUWw+xhFP8gWUN2n5fpMYxK8v2rkWDkBY5AvaVfqSClo1NDoRb
e4J81jYtagh0Hg7M4gDi9m4SrJdD2Qbed3D/ucFApdzA7hpBtnIfQC5IooilIyapGUbdZONAcFV2
28Hz9iGmFgpe+L6LZNglOR5hqtzemdWOQXD2HeZ6Bh1X8eHBETi3uVzJPrRfNTgiPEOPKRGgSjVs
8VIM55cYCgZnU2DDOV+Hq1ni5OJ9PQsT0bbw3fPlLU/nYrOAl7U2Gz0qCNRTjK4fLdaJ/1ntGKEE
00gKl57maGcffjm5FHeonbEmwDT/zyCgjaML738oRE4ymfc7Vhmquz4d2Hgs7g4iaX5Wh7GDQtnB
PuZUbwfWmWWL/k0v/GsF+3Qjd8Kby/Lfz8gbAK72jOX7KzRAjvrnrCg+YZ/18cSuyo/Sg2+7Tubo
PME5XbF8JehzfAnhm+paN5I7mkmbZ+ctD0fxqx48npap6iTC440kA8EmaYyPiz/hMczhb6+Bsus2
p7xm1XGWQ1pFkYs9IjQJIbXnZg0GVFLWvwKz2oLUmLRTLuPtPSWe/oqPb0a/AvdPcVQ3GmjODtCn
LIqfdT8q0EQzSKsjENF/SpoUk2uJ0G8YJIqqprjd87Bznllm95kk4Wp77Gp8oxaACJSGOks1BsKc
PGiCjNwhrVfpC7eu1cHJOPoSKsCCiyhCM5tMCBesFqwUvFn6I5/Lj86ZpgUfgXZ5WgKFAuQyS9lR
CvVn2jdUeFh2y3C7u2sGYsqC/mAjQrbEgYvlyLondhYH2v4VG6sxqrHB3Xh6zIVICDFwNTAptn0i
4isCSZ7ig+2KOm+S/qn5tK7iGO5lIAMhs/fYY7cRy09TgN5PhXW85QgcWfWsOiXTpHWaYFF5gCcq
DgBYRiotulAV/QGpzfikZlmNMbqXYCHby+0P7hjqej82uW4ww0g6tPAozr0+Dw8f/S7aKbwOixhZ
sgRHHsfj6V7h1sDHj3v22tA71nt0IoqzhHhIh6foY8VbKE6aWQNO6AZOIrkH3XMvrYHG9nueVltm
px/m9nBJxrCLncG8MuYpvkEpcLwnojvPrUXVD24vnN2TplDke8QN55/txgoYuC+5mUcz74TOuYtD
dahcLks9+13FJO85SwDRumslgAHY2mD41ScklU4ZA+c6oGINqn2Sf6lNB8xgUgDRgc4XPUf8xbhg
aMAcfoizCtVD0MWMiqPElBKetmuQEZzxQw74mMZ8DXfR4HYxhcu1VLx8PPP+qCwEvkYT7gzGJq5r
ZNLiQZW8TXz24HplJ0tg/N13f+8cYZz2AIJk/V+9ljtn9Via3TSI+BzSZ/joD4ZWv1u4AJ5Spita
bcB+QWycX/lE3EAwbjKsxJkVOEMdP0boqM09ze3Z8UzxgvWcP7337f3aNQebOkJND3y6Z+5Gagf6
oh2oKNiB2soisMK5x66Fjd/KnihdGjBg9RPseiT2Jtkk3pDn7TSdyfc4SBaBbE/5hvmkkhmpNK+S
O31F6hJCIWN+40/TJMpnZrqSaLV6egfKAjNwp1UHZnrC2RG6/BdvKtM3aVaR12nyYZ7+fOIKzPQD
2RDnKYZU5nXCf1hMiLGf+56kWasDnkxzyw1hsrQ+pJEf/Yowx1PZ9u/og1Z98sijQetQJbGKO33G
IjCZVWLBjn1DFMSI3lQTM7zzjQRtpBTvlM6EJHP3EEC9U6Ihl6kpItxmfJ+cbNfvC/mtDHxY/KfK
AwzwVdNJU2ISfPnZ5J1b9Q+sVJVDPPoL79B/YuLAw1QGg1HcijZXtCS7e2riNMygTe1zpeGY1mO6
7m/mVUy4fW0osczTVl8Ag0JCE2xpWwXXIgoe++ihng4Ff53NWscC3wVENZQRddjksMfkCBogPcqD
uUvLha7QY6CygCfOO4rF4IsJRG5pWsrkyYLL4u/Kf7TDE4xgVpKxEhoJ3X+/OCsu/QSU1T80uGJo
VT2NePFhUCvYTfnnEk+o3cPvJoFv7OBhxN8pBwxFxEA6PzWNEPFuFjFrxhwumkYszjNk5VSpwSI5
abeEG0TUe7gBL3uze1pMw7pm6MRB6sDD0nONFfRT9lq/xm7rYOSJ/Ke2ki9eHM76vJi1aq3MZjdc
l9h+6bEK6YCNc4uR94+Z/uba/hQTPqS7wfq8bp8lx3uhrVPkug0jmAk/XSseZ9cJJKUXePvW8ACX
8hhufWdYNztekOT4GnrBQEYopBrDLecZCUbRh5SQH3ddfyydx2FE4hfHf1KYMzklWYVcmn2yQqfL
gfE6AEoUeeKOAtcEYTCHe3xOup/Vjlv9EXS2J0BoBOzs83rtvQ2V87lwsCVXbLuBiOBk22m00Hqa
Y5j26Zrie9I0rze5dmtM7eJkX5g8PRgJP+ZtdBOcfYiUiBcjkI7lBUBcdL6jxla2kaX0Ec59Nzg0
OGCxK0MRou2MXMkq0Y6mo/8IUPRRDYahvPS7rLp9FPOb4/PWpzPGS24Nmmnd2W+iVoTswjvyKWlS
tSEQB7+U59PB81MDpkyojJMHGBNHglIoMgLGiu4Dfr6naclK3l5u33bZrhZFBk/hwbd+kq37RYgt
cgy7lo4AjhZ7RPXrWPqvP+QL2/Qe7OGlbJiZZRPPkK5gXF/IiGRtkOfekMA7W6YFub72mvo+ZX+7
vYULf9r7uJ+CA6GgKTlS+ZDvB0S+XhpyTGmCDcIN+ZRyLH+FNoAgr9eVo5TzXhKe5WzaMkLs3yoK
x2/5YbmYlbL/L/s9tkQKrRDm2P0d8kWFw1PZB4Xh7KmzbyxxxE7+5ID8OdpHsTloHgxI2O2wdaBD
Hbg+ItZVRpTiK/vZsdNRXeX4ZQf+6gLp6xNsKfXGvZ846X4XpqpB0taK+NcgWiDeHP0D/ghDy9Du
KeKCYGS4zwNer/hQDgZYBVt4yC9jc8zyVxJWasDUM+k2PwBQsN4MqDg0HbA9iUDH67Vji+l0Y63d
ZqcDGxenr7kYO1VQH7SdQos4gTU5SVOjJ44ptwvbYmVwZXVXcBvkyqQhXJxWblM13644BSeYvcaz
x258tWe7Yfsi17FjT5XlSUQD+ZdIN5GKuz/6ilRPieNUW/KF80heeX788ad9xfZCrdqohGr9T59+
h54zeO0r6GLwYOKPQHwXeG+qclAtpoPZlJ9y6JQJgn3K4GXXmFG3Bxs83mkS1q95knMJ3Bj9zZLR
/ZiIe0ci2BqKzxkYp6ahh4QNhV8qCHt6f3V55AaguEWpoXjmKLptq7LJ/ZRCwTlWpUQQG2Vuc4Gt
s+X/9+WgHDX6+2kIkjo9/vS9483uaJV8di4ewGz99ljIv8Fk6A0d/Dxv/5uYKdf1deH/8nunUCyJ
U3VvCZtZTM5+7sdBXvzcDFvzKLX5DcF2MQzef2+ujOgQg18b1o0RZMpdzRK1KVIgGEK/7OzAoNz0
xc4U3yE4QhxwtR9XoEtj/2pgUjZNHf/uL0eACZpAyyhI11Nkwk9lIoo/ypCCNDpV96mS0IEqcsAR
bkDOxO7QnHcwFxWd6ixJkNt/KkP+7rbOpNuSWZyPNOjjBWyjjygftbuVdwPsEQJhhuEYLNwFOvWT
lA/AowTn57yU8059y+RDc4El8UDedJx6D0i/ueUUjwQc7UL4/moONIKK218E55B2NIXba2K/9lbl
VbEZuhcK46Z8KgaYHDjVsI2QaIa3+yKikomuNbQhVYTxZPXuind5Z/gwQ/zKS4v3OfU/RJY8GWo1
m5pYC2LiiMEVJ+KGyI7zl6z2hdCuzw/sPczfzQJE/72gIClKvwiK1BDYm7GJt0ecbXwVFJz9XY3L
Ai00BdSpht7jxjpnf+zjRHGUVWHjTVDN/34WFdZWcLleOyX2LG5IHm2Ymf/aaxpcLWPfLAbFHAt9
6rGhDfqBex+Ondg2L4vCKh+1P6He8QrUUx7bnh9lbvpi4OtvckykM21V72OuonqzDdOCpL2dK+Ow
dMJPCYfrom5X7WPPSbxXeIoWNp4au//A5x492zKUTO9Ec4/kkUAiAkot3trH+koSl48iwy4PVTTL
WZjLnL7snBzUSDRlX9JhxElFVXBXhmY6v+P4+GcgqmMabVyanr5vj64gTmWJfxArsMdx2ET36cJv
RkW8h880LUTzWmV6WOHJHZ246fXC17a0hVBXWc9UpEx4LLGMEeNPp9Kr5Q4IzonSqDxV/CH3n39v
qabKfFK4CSenLvS/8naL3VdstcVseTpDFdY6XhyzXyYQ/SBhl0xWeYdixXcWAX3CiBPDg1xi/t0Q
KvJGLsv3Eb7FN2/guOYVm+9W+IViOCCnPUEU1OmacXyU1t6mOF65px45JSQ21JvaQW5zhqoa5M9z
oZZ9ybTDikgDxEkUuSu1OUMZei5TQdPoX4juWpYTu6QOOqoXtoqCLYaPxavAW1oddaQWYdmaqo2j
XyD1cZIkC8k8q37bS7yqu3880wt/JLnZgb2SdRfSfGFHwlfab5Bn9eD2fmozLIWwLvAEplQ5mb7C
YUfD+/+NitGMvcxK0m30pOzhD+K4TFW0cYbho5VWQHQibqX9r4zXUD3XY1xgcv7Uh1UkvapIsYjt
bNpnnY+8WkOffvsY8f3Mb66oUFVl3bQuszJxPiH2yd+9CUyaMunVpNtjM3VrT0RorcAOb05/pMct
5LEBYxV074ZTrFH5BV93XTn3zHfEKVZvw02WwkhsmXTcAxesiuNORhDv/0kzYD9CbukcbwYBn1iH
qdpVLIbgFBMeF3+4ri+U+W6CIUmM6mvcTux++YQjmKDiN5b3l/TKjPUvT6s9czQGcD88tG/zfUXM
PVy1iW0eNzHBmxP6O0ZoRAQwAux5X1PSg+zUy3Vq3/Gb8G8vXav3ggv9yrxqn6kjMnOmP7Hqy0Q5
J9L9RZEGHdQKZnXxlzSPf9w9eW3KzGiFgxMmVE3rJPwySOrh9qEMyHBBvh0bMxtwrX5xRVSVwYDA
hCDbnviXE3zY9MIlOQQbmz9WOavAzN8k+0i2VlyVb8wwZbJuG+U4igIJRjaRsYtpc7l7zi7dgbTr
YexrFvK/HD2qwnvvuAUDvu1wQWSZ3mRAFdLio61ZM/978KvqhvR78SfoxjGDqbrKOK9ccJl3ERU5
DVp2CF3dYrZusJE63hCxDDAET3W/HvBuFG0gnSrQ3Jt7XbL+0j7qKjj+9PnZsrq4hd1O/PK6+Jx3
USqC1gDIa4rV6nTsEo+R7JNkE5sWgUo+g8Fc0LhRa4oAT2m1b9sPIO+DZUiqnIMXgcAwKMHKuOFp
CfE+wbFivYlRpags9LmnoBfEAm5ukYWVCJbb4KBiZPF7z1iSV3P5ufTD3cnQ3s4XKDtgXvR1DRI6
gsUEOshsIp57S9eA7Fn0AsS+3NF1Eedb0tMGmn9Q0EuO1x5MjsC8x6p9lXz0+FsQX+l6Lx6y5K5t
iPhO8StVrP4h+IRaBXHVuGslgVaULxsa+wf12LqS0N8XwmUR7vWlJlb9/LI6QJ/8q4id5/WjXCM3
YX29CZixdr9FeeVbZ/0O5kPepn/Ysi4UkfELVkGrrbw8fXG8oNOl4jJx05sc7+/HKzGPkB/6oboh
o2vjDjWa+6kTcHFm5Zu/xJilnbPE2TlwboWl+9pcrERR8MlwBL1Ny32YPYjkfpE19df5bXWn3Gzs
JHBwaAjPMOLEscXkkxKCCl+qS3uwWiXTNf0BvRBA8HmJPLkwmtf31p9nS++mHRzugtAf8EDsg/Jr
OdFZMxf3fZcGMgLl6IQ/kJ2NKR7TGQPL80Zzk10TV99eroj1g5zl7SBKKTDvQYeQR38SeZfH31pV
OCGUcLgC5/L4Bdi7vemM3Me1DL9nIzAemv2x8f1X7/SfX4igIxUSG5cxn4axXpo0DQR7+oneL38U
cxSzbk7bBeNzQw+TMg9dRSXNhc1287muin8wCdpmNLTq84hAR7Qf+VEShXsOnguANSD/6UxJsBc1
Sxl5jGKeOy4BwBIhxPwaK35ebfI/JYRdLlZjAfV3pi447kG6i6Zmp1zhSXwExCRo85T1emHjERv1
Q9zBFZ69kO+6J6gILQMnIZt4pw0PYbQsd3qBNmiywBoTJ3sVg5opNn7SV3eJiy5Y93RT/AQu8Hua
MguvCY+ihmGSr4ypLIhqWC/FgLO0GK+aOkZOq72xRsauaPRVMEexo+juYjJYsmjyOYEvQ9e6LI5W
84N7PHqs6Ea7O/ENgi63PrtY2gBPARSAB/LjfxG0UoS7gI5WQQpnWKVdUzqh2gHOyZXBky2WqJZH
EVdVKRi/CEpjlDso2P+FSA5zzYLlelZZUsyTSmNFQHOh/3r/241avrgjeYpeRP5nkmZiDA3xzzFa
e64cE2BDu9PsYgHJ1FiuAbp74WoxfcXNGbRfbDpC8znPyPcJc1+9xAwStX8imzNsd2pAu3RKnVrN
blDWcaLikbF8Wf0hkbnlRN1PgIwLMbABaTah3BpAZHb6mpEokcXxomsEvQ3G4eKbAfFL1ZuEvysS
dB2ePoxELUibVSR5SZvAgts221QwAARS0Lks+YmBms8v3fpcrt6P7vLhtXNLujiuS8Ofi8a65oa2
0vjVE/z/P/w+eOJ76MKuyxSwHNLk4LwanSoKdbzqzsCElhMB2cBWkWmFQzAuabxDVNEDC3aVzOdN
/GirtLr1bw8EkG4ORfJ/14A1EHWuCH0Y/nhvGVeOWeRIQG0i+3AKugxQ5hHKz7MCOcdoJxBfL2Nk
EmRlxS53Opr2SpWPFuki4tAUo6zqy1u68qHB/x1eSNu1T7iOeT/ChAGF5GczH0q7NUl1HG/jseC1
ZjJ6AEciaLQd2EtW3F3KqybhelySESnI6+WwMuF4HV+DMduej492EwwxqN8Zvw/4HyLONHRpQPj0
oLum/Wbw9tjG1pDM2wmYJnon/AmWRONJ2kjQqASh68iPUNM54lhQV6LtQXWMfJD527qD4/fnRITy
F9/4BHW7IHXqBr1Hfhcokt4jgT8JRRMWz8yLyyWWkbFDB1KHI9Qpi5UYa1DLpJRDbfkm5s9yXAzA
wSeS0qS5xg+E0cV17Ufk/eob4BAI7/Fqpxblmq9R5VRuPOoy2JQLQK2RdhYLh2ym1lDGZlgOJJ+h
YfTFEiEiT6vuakNzT55/ZbZK89ONWQLiumRBXlneKtlK+JGBnpOAMI4keV92tCHCI8cXvXMXabB1
TgtJJdz6X9tlDiOxlFysF68DxwLWUlENHFZ0FnO2Gw7HPZ8Tmlp2s7kA6KmJ5Xwh9PEUe/AA2XRP
0+xu9Lqjn8DEWwVxRopp4nLaI5YtIl0ovDgjd0BYRKYo0t2lD/vid0TQ2npFCWo2NMugsb+CToCM
HsQiK0mhglKze47NOfZyi4h6P54/NMJywmA63M+w/fGUfj9mWClQnUpesFg8s2C7CH0vanQXT3z3
j8Yq5gbZqX9v5igL3tl4FAL7ffYasqjCfFeVX6GA7mUaPBM1tM43NI7Nh2ml0PfpOhEWp5mboHrA
jYYccZjQNRYIK/8yaHP2ebJXY/jQ8SONRPOp7Cd7YEu+rOGTF2LDE9dfyAhHKqXvNM5oXV/FkvhY
xIKepKtNw3uJ1sjOIOgB36KvDu0rQZaf4re0tTZdr7vrIgNE8/KyRi70H4mWGnP6nH+RbKblNUvx
bJJmMBmQF9c3xQ1dSz2DKkh07IHEc8ahH6WJ2PCm1fSgpTKtFX81dRQcbRhVOvqeHDT3wuz3WQy+
OJMOopzQaRzw/4g+0KTfSZqcH5Q3qwqH+O3dzvtiT2r5f0SjocJRpcLuM5hDjYNVjZf2wA3us61g
Euq3yFtgIZ//2h9hobYrjbF0BzSNdhDqtJb7pZafIYsrjg8JdrqcGntv0SkEj/+xIMX/SnTHL3fv
OwYJUxokbTtLdv5Uq6iVU4V8GJoQUKjBMoz8T6Idy5DedNTX8hUed1M7M7ychJ7jC9LtQdKCkLAr
/K6KURyhZ1oZsEcjvoaOi6D8wFwUnQ50MP92kASInIMlbME1N+81tgQ0AlGj7oqoxn8LJBF/X6oe
BGa6UP6ELgKngvUT8U09u+2SIFiIS9A2ZaGn7IyoJQMsbS/n0W+a+uAM+a+olsoyFLeVRcM1SIBQ
vjbUQ3P9A2IH9bUbb/HEdjrrMXYbU1swSJ6qiKY60B4+LLaLiJAkPQnsFQWZre/M8rcXx1uqQ4B2
zQCzXm7uz+ymUaX2NRIfkm4J831xyPKS6J0NO7Oh5Sb3lnLpVQP67gTSpPHvKCM9oH8KqJm9ZrxS
5JL0d51/buZXBaW8xq3aOD3nscqgBHany2WPbEax3qTre8aep7qHmd9J7k+U5yYtF7LJR8Ws9cMl
QRld/x9rcI032ZOOg6DxxUdQ0A66kR/iO3ZDZSVDfwpiagwJq1Y07N21+Ypzspce4A2b0alcfS+x
jimEwCBHGaqoxlXzMJGhrOmilJOnWbl5PNrWVYWfmWr6pqZl46qo/rg5h/IJvnJtRS0pJa1/p4il
+oaqYcAC9hGx+Ts17mKI6axUBc4IORGueZqV4RDcMu+5kDyH7mRuSWsRpW+C/8LPOhLD97Jszy6P
M+7xpfSfSBxLq5a0RGk7doJOVskAdV328pgErXI84BlGNQG/J8EJGaVHt4mVgiMqButw11CAHr7h
aXpkCa9Wv28eKP8pHjr7MkAELYIMala7/Tvn1NJ6whrz30H6R+nycRseoBtKPBCXr2ohDCifNcsU
2GSTW5Hj7PXG4hxRPFcUaCmubS6n+TNvDeUVqWKdd/PyY6/TdDnhaqafd/1PhX0eI7hyk1AMYtcQ
xzbhOKH4lewHNRTKV2XvlpKwqoc051C5sjJFHcji8dQYzP6oluETIrJ8JFcg9PhNFfE1gYiAHZ4i
3mlyttmS7kETtqkdhBQbbFIEJxAAR9GrNheI8u67ogVM68y+dtGWE93O/T8FSKe9VS9ocGi/Va7g
cXgqEeOgdIUE4p2v+f7Jm5MHkEf+UsvQOXvKQxuQI7QIS0aoV0HwXIc8DwUij1BBhX6Fn4GSL0A0
930mcnEdUxZxiotwDKaJ6eky6pEQ1tdOLTfpnSfw1hqWtu/FIQ+1RoUZbMaFYQp+cALmmXubtHJ8
BmDRylpAVm5mODgXFhSfxURVP8fDIpV/NBLUq8b5DiyL+PBodnfFWLCtdQvbvuQMqM8NEpMcmj+9
CNL5g3mtLFDguPRO5qWk02qfg6SFVgA1kJ8A8FgDWdiApLg+LXvG/K3pzC2NtlRTgJNrVspirelA
w9bZo4bPiePWZUYW5SydWYFhOex1d03yDCXCQqbCWLquqdEWI3lKoG6bBe3glRhZtD0fgLoZptH5
MakNRYs21gSvaPf75bjWEONLfDccxgJBktzODLkxljUhKEivNQzq8TUaG2rT1Vwr2L9Zisx+Kawo
/P3/Mj/u9cLGMuwjOutRUpDXZaHgiGYk3v5ie5GCfvvT0ajkk+aEfmUx8y/qnwAbJ7tMhsAXRdFs
xE32ratoQNeGwfwvitgfTr0IegQsKGi6flEFb/I2DiyJEYB5EULDs/MFcnpdp60kk6qruIcjRZbU
V5k0vyjhRt7uYERwPBW4/IIANQbPyyggUY+QEKOnuOj2wKAtxNIqnjlhuvkc/NvtPZIhTLhL78we
QCUZOcfA7Zx86QQjyTHIgS9+dtpDi6vntI4iaanIvEkqGfX7WEo3VVu612aNxOSSVLIL33p+dGV3
aY2lpdg+LO3/Eu3Ds61FSLCpMiceYZTTzVBdbXA1kgORxwcc3GmixAyopVeUHb0C9CuczNYq8L8I
Nw4UjBf9fZtzCCr9i5+0aH+mk1/6Nts1AElWxOZ3ZWTBkv+mLw08QgRCToz49yC4mizkzl48VVrc
dGig4kQ7v2yEWlId1GOPXIxg0+eSKPC3HHysGLqv8YZ29RK2q8EHr6u/sB1KPp4tMj3wOQjjkqkH
EZP9imblb7Ek0WI4t9mF254qYhOOecVdxgunsi8uA4uZic24BoqT0ot3nkIzeCrL0aZiQ5uDS1ST
E1pmgTButTleIyn/BXU1rObPNe3gFpE12zeFbGtezCypCbaPh5SgtEtXpTz+2Fkhvgy4uaNu5wsb
zMfrzoSivIUuVa8C/PA4tEFSy7pdxa/ZybybsoIIx424iUkzHKQPURg5hdwGu0GMEcDwzjGWe4+y
qEP3dMx3yiB+mAAA6Rub5kZVOHavuTo4S4SU+t7RcWxVsHtJ+nfZj59jHi5DLro3z/HJjYLhYavz
ztThBXW5IcyqrLNcs3u++CDJK1Hx+xvzPyDvG/itpSsQh+++iGs2ocR8rt5J8NWqhxEYTKhpz7xQ
eeTbPpx3YPek6VMU8y4KtTEhH9Y8puyCLxkCNiWn5w45U7ha+Ci63DLecUiA5IMVLVd/3e+d8w9b
6oh6ZHMnj0lKBLwSr3+b3Jwf2riRzOHTW5vxJ+WnXrSrraxOCHjcW4d9ry2jMxOisiE1Bl51fAVM
a6v6PdWo8apNKmUtT74XuIZPBMgTL7C4uTokYjVKx2g+/yWsC2Szz5KGIzRmpuSEExSBUQVvjXo1
ui5vJRPmOkN9gAwmAwTx00LZFzOsNV6KWxZWM9DKd0GIl0+xFWew4yAyG46foY23jyCUM5aVQvAz
+JD9IOt1kr1VTk77KPtUuwiSJ0zOcARGJl5yeiaPEZ7QkHCn2XUqRUcL9X23mGwQAzKsvyq8DoJr
s8XzeE9HpOCfy3dXiHzjXHWS4mkUcXJbyTwJb/O4RXxyA9kQu14cRctbIPUh7LqWDnOxRxLome/c
fTXBR7IFz4e3vqzGeI6+ecHA/omX1ljibLQI3fQ9h10ZPqipbN9NB4bOukdBZLcLW6VGLUpHhWzW
hkXSngSRU/UbCkkVuG9QH52EmOwiW3PA4vcPsJKDuxSjPHNrGHLIBcCL1EzDJdtI9NXsErYpPqkh
3/EjFI13LjtnQc7UjQ/JVT1t4cZuWTlxFalZSiKlm9SG4Fngw9AxJxZ7AMUX4ecM5Mwxe4Uuf8+T
rl+e3gkDrkKNCmRZHeLdte9lFsouOmjQISC+kNIhzZQLgNbxTNlm818wLat+lW6CJF3wMWuNdjv4
QeWX6V9QIiMceYEy6hf0+gfOBLK8U/k9/Yv1BktJ0Zv5Q84yrPGUZOmFaY8wAm27QVr2suLqqSQF
xAeWtSSEL5AszfLVzfibSun2ZAHUG50I0gJnlmpc5AUPu1ulmagEVIi7MSaRd/Tj4oTQmSdU9jRe
de5wNGs+7bTuupP2NBwRe1cgZG80qye8lzDcr70vYLZdS/81iwFcRIwwnOkzKEtRpv9EeiaoOngQ
VoO+v0E3LhOIYJQ2kBZpmLvqYYC4nkmYLgH8BqvEaoVbgE7bDEeyjWC4K0TRmFrciojxSJI67Ilp
nT2QegRjV/JWpbTiq3HCyNy9biqwDiPrY2eV3oooqkisPPsSg41hvpSFer1DLf+k/+anW4J4r9mJ
6YuDJO2sKaZ9jmnJFVBd6hweg4xdAROF2t89BoLif2hwkRcBI1OXpvzUK5IgZmNjAkpHNiO5mOcY
iDfMnm0KdkyW7ezkNV/c9kreurcMacFsHos34+0G+PvhmV0i9A6a9cVDVXwGAjcuJVJL2bHQ1frP
dW0GDct5H9MGX6NltnqBXDLmrhho4Sreby0Oy3ZHD8wo+R0Yt9ZU6aCiqcWP61QPmdHAXz4cgVcK
/BJHE7hXOS1NeOX/XAcx2VHPaCcYCa5hVCfhhrVG1aaJjO2rL+R3v4Iz3bFvViaw0KnZaAAxsKJb
VP3SgoeoLq65c6sZC7Xa8ZJqnXSCcDkM43FzgY7YvhB3jommZxZx1SEuLqnPLG7RbZ32dt/AnTv1
fRNueosgwt2OMgLRn3iM717LOmWhOEOJa4oQOtwUL6g0kUmWhmZnwGup8WEC++4/ti2TCpqn4t9b
ngl5xaqjbHIrzJl7hFd3PTHWa5ZkGTwssTWrsKT0asFNDUjhGHuLH34FSgXySOG5IC4CFWQyXKLQ
mE1HE8e9pF/j4JZpwkMbaPzmeOB5iSwzBjLRSCRFnLdvX2iN5DjYHGKA3Idh3F93di3gZ91OAGwz
3c6JSftT9iSLWd7wSZr75AYheyL44jSzfrSqSTnZU0kKwUlBO0sRcrkuuJJnP8l/p24gkjLD1+NK
Djb0S5ZvbWvUUJydL6nH4/xe2QAE3K0TQUrzOHAgd1FxjwSx9yfqWy7THeaJEKVAxkwAc4t569YL
LsgwsZegPE+tvW1uxjiW1Il511FcD/elbYRPNPUYTDenKFXmIoi0UwcCdEOtANzBkH5WW4/woG6O
GlfEywaf19JeF51MH52tM1n2XXhfJeuuwOkJetElG0PN3NeWIgOLXpXLklfayzmepJYqDa602wwa
8EE/rZ5pDFY99ZvTb+Jl/9vnraZ+jdwrLobeu4vlVJ1xuZi8jJgV4YcQxm2mDp8HDZUBjGkCjgLs
5XdsL1+LiV4D7+WguwSMJo3AVePSanAJrci8TWTa8i4a16RCtNl4f8tpfO7gkVhYxadqGGiCbXrh
ztBhmVCmeWEpHW07qxz8mzKmRocSoRS9MR7GgWlmDuL6SBJWNMa+O+yeIYCpD9gvidQMPSrJLOSj
rVChDV1aLMtrUYPcLHczWSImFXtxJe0ePZgbhzPd9KUAqdQ0ki5yNRIjUpHA0kM7+jrMQWsJ2i0u
f+IPIWEqiQUvaaT87Y95j4lEWjAnqpiua9GdC3/luOoQMo+nSlttYhrdYqEwVTixXx48dzARyBOF
u2PcwLGeAkZpO3sQ0U+2uZoZOo5+oR3M/23CUgPoG0/6KMYIm1ujPQ5gVIOopaDizlXEsUy764z0
FBddJzg0aXZH4/48lzMMfm8m3SPX62WRuaHoFu7m/byHwppjatw26/j5DUsoc11vHEIylmYD1kvN
jQs+w0Rxi6CTVUaxBo0rLlWCG6n5W0SPhc297WlVE2+xTJQT0LOu+D4xqZp7irOG57eZys7SePYo
qgw0IhO0TJYFJTzsMFcIvhAiMEPs2NznPZT36EhutEToaNEKPbYvFUEkJpzz86dw7YipRhr7tQhW
7p7KTmXJCkYjecfdbhYDwH9ZnROpT+Hbyf1EKjKfJ17PSfyuALyr6uRQzGCCClCGTNFRKyw37WR+
7reg+ZEBr/g+VkUQRcQwENoJW8X8qw73JwE0apdpIeJMhHebxULYt1pRoWK4ALJoc+nu99cqq1rD
47Z5N5s3aglRiJrh4jt1mzvDgxBlJpvyJyFu1jtpGSbILXjPUT7XTuSAWtpCckMlly2D4aZY9xIJ
p/ZW6zMnOOgelWVzoxkqNy/+oMR5w+pwlIhFrZ2rROe7KdqLY8SrGovp86S6C3T7gLuOrtP/Ohcm
O9UBMOixNCnEgUT/gQo8wN5Pbkax/Q21rwlMoF8KFi9rvz3FOMSTKpIeIBr81GhWapaw2R0rywdg
0iuPZjvw9MX+gB6Pu4aY+urW9mfWOnwYQxGg1HexvJvWcwK4wHtujZ0UpnTCoB5feyAevG3pYgrf
tdJo9gmR/6hHjzenDKq0e5IVrxgYI35YyE7dP4eyZ4sV3Evc9LzX4L6kf3MYKQX4cSIsFW5zdakH
AEUEu1Rn96CbcEXvHpvm32/PxO0HEK8xFC0dQP7wCC6LWpm4YuL87dOUXco65PckfpyWntdrmsfi
u3K4e8Grq6HZoPVI7Bso8GDvPHVBowUMD1GMtxUleSXDYGpdEobTbTG7y/EQdMUNlzRqLqS9UkSO
J7SkJ0BXPP0lu5sWT5/up4haNKeb5rxAUaPKky6E9lH18dY0Zn6FhTEmeOS1o79qnrsITdmcxj8N
eux3jggEwz/J8Sdp/hOwp2SLQJL5dWXcudl6XOGMbcsexHcOgT7Wiu6gWb+AmLghMqnrP8bdlTlV
lv0ZAaeIPGrzFgpcGsg5lIqlTUmZ0Bv5cvjrTZS7QVusucZLEGdyn+6W7WTDNl5Zl/cbQc+CpK5E
eXSkHUAixPMeO9AIr+jyyOj4YQWMObZsEXnY0+Uvbw4kGKpwh/e+qjsSsuVGqb0Q8OA6kK331Kpe
ojb00haUg3+GrYKHtfYCDO6ijSbaTQf94ujrHouPW6SjdtpHy/5aG1bJJV9+z0C2G46Nc5Bqfbv3
zHRq0QnoffFMSkzuXz4mVWKw2PVUDQfknKXzJw7JUBupA05LleP3v4cmS4URLFNfI66sSDPbVGF3
01aeZtMmcMQ6bBNIbpWZ3VTIc+o1RSIg51pLCWsBBCAlsuD+EPcW0e1pghPVwxZD3gtMfo6ysdJ7
pkXJp+GmEkwDiZGJ8pih/OTxoBuBwT17RVI0iBQ++ZpG1aAAl5waI6tr4LqjkWSxr5LNBxpG1TID
CsbcIlFOH0sBSW24a3TcmGUMkU7/XGYxCru97DyBlK7eA5s/CCQbRxkjlMc46wf1NKIcZPMgT/Lq
faHOyMKelGEtr0cXJ5PRSZheV7jwxuZQDrK7MtH/cKvyniQWXpO1/9ZTMNwsfIjXEWITL7gHIL1y
cTOsjoAJZtFjhkZYSPr+R4mTKw027vlSxMOFosU5zZ36/zMFJ6RFZXSg8/vDTsZ+WgwAQE2Zwxvn
vU4B7lYxXXJtonTgiorbFEKwv4hh0wL8avfxvtZ2l14pnTZRmlnH2gsK/hoPT4H4t2ttRb/LTEMy
kiGrTer5Uqt6+5Vs8D58EwZWVpUrRLj80RX1bSDbQ1YgwzK+MAqgk8nsiUbW+4uZG8dmm8M7XivG
EzjJRjdsA5pPSccFUf2mLYJ90ZQRp9xTOw5qePOdzMO5sz7MmXtjWkhBMCbKO0pE0rkv655wYKVd
0k6LfHZnnozrQ4b3MWiigCRRtig1reYqbxEbZlKbw1hcjEQUbR/HGeuaBc1I+nXypDzy5rJblqAo
nAdaMlMsMPf3BgZUS+XLq/ZPnvIzab/z1rVW5M26bDiC+GVElFbKp8yj4oRl5LqfgVmYBacjBcMa
MiG19uKlxVqtXNq5j0n9ZTVErZCUDE1MQ7lhJutmyIObngpkr7QV8EVDNHdFXZzbmr1aezFf1K//
LrSBS47rtlfDIqEOBDjI9+6ZS4Vcda0BQaumqwROB/7LhQDjQaTum6JCkKqTamyB+LvV7X7eTDQn
VX1tAC5/1ZmkxecE3QQX6wL4fMZWAhNQfoOBEfyOmv75/CbD5N4t9ztgdI5368CgOoN2kSWG2LrI
D22BB8eoOE6WoeLaIoaddZyfRmvYLB4SfOpDHi5Tw6OoXwUUkJPNtc5PT35TR6AHbMrTF3Cf791R
Pq3w1QKabMG3RiplNxYe5ZS3LDNZoD8F6VJIKDRK9sUR8vMvq64uAqT9Lli41H5ixmSZkCYb2iuV
GwWC66pV7Kr707i2J13T2IJbamMTaXbcWDcQFUZhAVX2PPUcys1iBGgmXVxn5xjtGUafhmyba2LN
K5qlMsI3mfCcBtbVpt9WhQ8K4SXooxh0DgiNLfjfGwZz3XDpXNYkqFNzskyHuGs21i8wdNcU3JHT
yNvTJKP4BcbcdtxJNJmiwxpG9hJefnqiSiIn6wJONLwNOD4er0bUv/75CnhZIHjQ+q5l0G8D5aKF
UG08wanvXRV/1u77vSs+e0R8W8bncySydpDwgvGRaTAo6rPk+F2CeYQ9/tJxB1vVVoQTEWARQlej
XQiJSe135YevCWxziwUhGswHqVd+80luez/49sgAuY7wDUIsPOIvg4OZjE51RV08H54RpTgjPvAm
seq48vG1FwuSGT4t63Ebvf+zf/ZTF+W/qHxkyG2qx0lIzXOKRoUi5EL23ulU24FrJpfgYA47K+0V
txdjZ0aypn96Kd5OMCAxef6lgTTDmvRBgdU1m+V9OtVWamOEmhxzzY+G6Du5brtW1+b6Hz9lgXCe
zKjIOB4BM3IRWFeSbdQRZ3BegfGq5q/mA9X+wckL0fZWHjbfxMyOmS0cCv0YCu5YFxLhDlKSK98M
igdGZmhkxCHU11WTLqTPzJ4YphUYqeJBoJgeqrj102p0zO1vfWCh4ggkwZhHMVZxPugmByH9tKUk
oWcKO4+F7fBuhwiBAichK9Bwnw3P/pY2JlKeIc8sV5/EpIrSO+P/GJ4aijgtkU/fW781wIDonG9g
0M8LmFzEA82YY13tlmADq4gix5oUY6ktn5Y85sV83/cvnkzikprs407PXQdKGvaWoVy7yXMjZX2f
kiuqwb/Pw6mY6xqxtLh5fmoW4ZfJoDy9zyFT3s2t0VtmDd62F8kr4bfzkb7IO2G5uM621Te/aX1I
HHRzRDVJLfULWZeerKd7WnSA/FkK2ffL4r9DdGKDCn7kyrDKxLaRjw2bih4+O8XHiDgC4yNtjeQJ
YmJRjK/GTWnJMGJGOMs9k3cAgWrgT1yiX3yPwet1tTYdSGw6HiCsTgN3DDobweGoo/AoI3t8zRwr
PpZDFHUIQLTFT6v5jeL+jphw5UNxPSijlCXWKFDWcrCwrpqAjETW6BRNIGXBT4kBVCPf/xwhxA2m
6eKONDW1FgS7cyRccoQq4JOG4Z5haAkPGrcbNhGb55h7PLb7avNWRv+jS/90EoYPrNVTU3rMfX7Q
ErTl0EJj55+/03HaYi+oHQ3J6hVpHp08wDgIhzCdYvDugI3vfDR+YU8qyaYlXQ3zO2hQ8HldkCzB
1RVm2gya9UHCQv6dnZkfKAtlBaH3szMuHm9/mXY5lgAtc2xPlqHZu3QuZyo24qzirPMJJ4uvwPpO
mTGRBGV2XMgxGsBEwur6nRFIvRaq38/fMb4od3nxvcixe9CRsAM3TGKqfKIKTO1XTJIvCgP1fffg
4Pte1VljazpmANvn1/FElCPcL1izMtnXUNsO1V02fIfHEIxt/VmvXzaSkLprLWuaOOTlZccUXEpf
uJ1C2b/4T65QGk4K6vrgL6zp9ROKgIP4XPfAvwS7mULr636ADIHDhQrDo7MFzO136zmbHIqt+c1I
vy12f//oVakBIvA+Ak+lncZ+SKp3V3UJx9mD64vbPVBwWram+KGh8g/T/8y54RyaWPL5Na4nkr11
qF4a1QxRIy70fbXfaHZ0WFpi7cc0B7TLkGN8J1gMsnuVWekb4tzgNA5eEiRv5ehQLZJqobOQA9JG
CaDTUF0LB/3SQSQeAtsOp4UDU6mPaXDJ415nwgDR9y0p5K9T5tswT2H2H2vmQqViKcHF3L5zW3Ps
p/xU76iC3Wmc0qfZo86L/Ahzaftkpnq5iXwWCMHZ0vB4NgZrvTa0x771GBRhYHhXq7ochxE3cwQO
1zhLqnW5/TtEOF0BTjhGhyTbTIXrl8l/r2wV6NerJqznPsL7GvfL6/xL5QrdMl97z83xQRsfGhuc
GhU4i9kquP/NJbY+22gERjjZta8+Uqvx86rHBs9XGuDgQ/XhY/LKHuPealREahm25NGVQxkjUL6f
V2ldQzK7P4/pXh/I0AAJmZQgaHuUoTMVcqdyo7XWaDFtBPqhp4iJJiTsY05ra2GJGaliJjMKepMh
9B6k+J10wAHGGLCZ1dKS8xbxQbB7qMz+/SDBEoBCtg6hnszevkyYWnvpqGt8YPYDiy6A5yRwdgDR
bsrYj5Xl/CLalVeqy3cYUNEsROXtIWutTLmUWOrUNsqjXIZt5meubqWHRMQUPfmViWmzNhM7uk9h
3OWn/2ulukH2hV1bpBhA1fODmByvOg3g249vhMOVXm4iqbxzlFpVMIxWuginKr/8RNYo907dkRrN
nQ01dO1vJWonP05mk0vE4E0UeId5ME1FHC1UPyOr/nvuBhyoyZDkbVVWdWrD7Bu5HYGyvRNxjyGU
bCLJ4gyZT8olCrLIg5txNQpmK74N2AAsf3Q9PCOf36MLz3Jq/pMHGbmAUJV5slFl4pzEFRo1vZx5
uVDfMnkKkSGp1tlYRhdHJMeOE5OV4EbNpRrsjArLELpvQ7c33Y2ajeSreYPAc0+PnMRcPk8DNzXV
tODilAZVguoquELD+hdobi77bnuO0o9Ah3MxolhDrHjMySUsMqGdWCQ5gOjE/pvOe75WBGP4rc0/
kqPczCRK9Gx5aGf3lQPlh3ya1WL60tLa24PG/R5itAvjw0NtcQ1Z6opNZBiFURd+PjTrfqbdVL0z
uvl0zPgkD9m5kOntliLE2ecsTP6urGkgJhCxINAg8fsqAlIii64PWlPj20mmdoCneRNntCM/gAEB
GDpqVNIysxkfvf7UREH9aSj2ZmlKLW6l+PtpBUV/dVsulTS64mL84pnrwvKCmxY+YfEsdrVvjXgN
N4ea0wyw4akWau3ReMiXHMbbGpJmOk8WZgi0whidodROxOCmy/7s8PnkWCEwhqJNBJcatyQXer2Q
zzZngFW4KmzQUXx4WiagO6NKUwkFV/zwg3GXGI8Vj9dw+obzTgEF5WZUPOnZyVQr/bh6+2wATsA/
jt2+inOUWWDxj2KW7Y1zW1aM4F+fX88R0IjqmNNNQF25t3AytZqjZb6dIzhiiN+PeHWdVp8vJcsf
USJziMQFUROYMtBMEpCB/kMv2rwoDNHobb/RSMZ7OnDL2g+p9VAKZj/YeIyFg5aDO4+C49HoEMAA
YHBHsmZH+PIRf3gOba2RGfeZNysLzVd+igD5bpKuviuY/y3AiUsYlLNRtNxNj7y2GLhJbO0Fg7Rd
2SFPm/DE9O5latZeg7T4J3RkVmskD/tBXI4zkdBoUH2yIAwi3qhJ/iKh0d26Njmg7YGccki110+Z
B/UZoqlH04f51Ve50YayBwsJYbt/w8uNZnv0hsXq3mF1Sxk28gFjZlOU6/fI/jwRnCN7VTkf4fl+
6dY+kVh+ge0yh4kUbFDzRkN39CY9p1bqoG5mlFqpn+p9w/utfJAwnwe7Qb2TtUicxBo/XxZnUu6r
JpJOirEAmGrXRr1NuSazMai5v0y4VBPiD6Eo1uXVMKSoGiHDcwu7xBFcA0lNPfyLOhK/IEgAR0p7
WbEQDwAjfi/Iv2DhP9KGhG9LTr/V93No0yQXZ+N37s+ogQZgFHpBYMDPPW5ik9uzttXLS13PgfiY
4NvnHD1zb248itdI3a4lgfIcLgpvjQpeviasfkH+eMhSvCiqGz+Uky3el1awU+Z7FOigyv5YppiJ
dUTBMixznAKtOUjpIgtQ51rYpuRZNVsULm5TFK9R0fG6nGIIXtQKaRxqJdPkAUBrEmbcjeeKuwZ6
cc5Ub5qcxag6rP+XB6ph/FbuG3UZ7JIlXMK3+JzU8tLd8RUzmSw6ZAdhXoheH1/zaK6eGO+HjCdb
uUQQA7i2kFXOLJfF2pXxFxbPNqglDCXJw3xpBPiHUV1Sb8stqFMf4iHQ4DR4tKW4gioj1/uVlnKy
sG6sDe2C13WEHAH/6v6nevmfTAxq/ziXUfIjfqeUsoS2tgtsFOXANzBR7lOQpJZRTbOMlEWkbqyq
vVctRP11Jayf3dnNz5Dn1AFYxNk2FeIdmVmPT93iIaBKOulD5AJBmvmVR8MCKUIxMXV2kmhbctue
B0qIaVfmrRfOzfPoIIp7vQm8F5ykLi/37KGR6Pc8JlF2wKgy6c6DTQBW4anrBDbIeiSQdwV8gqEi
PMo/0DLgVAqD2BhKkSd6vUlC3QR+QZDMfLs6YoHWIdi4CoFkNuGLWWMBLpbA73ykQQJs3qmWLnMp
lYmBd5TRwVeaYjcLh9/KjjQaTs1WMMA/aKNfSfufSwkI9UB42amyYAqy8YliVOwAlH8XrkxMCVrz
5UzjQBtryYmgKC542fqLSx66yI8yElaUFMmHxDzzhtLbNTEt4H2GgyYEljvo9e0J1bNb+WFtUM0j
dE1BPPme/hBtRhKHTnB1NOJHoznRjLZytPAeMWg/0TTAiipwRtwgJLUzCIKici6IN5Irpu3RMu4L
sddsP//u6CvmEudAR1LS3VrsTKzdwqZVbcF+5UM7YGoAf4fmFGJmuKZXYar/GLm+6Xw1tMruuDfV
98rsY+6ai0g9pVV53K1ykq2oHVvXBtr3oePjHPygp3NIhqcytbCY52m7YL7+pi0Tk5uXrPTI+Yw7
vn8qAGtzqj/AvcxV4cwLKKadpIZpzauPS6qa+PhLKPVZ1rdkrDlXFl3a6JmaDw397ahxtzBVdap5
4Pe+Ez0L46udFA+ZO4f3ttug69famfHtgkLbDQPuyDaTPc0N4FgTS3NPzubwKN3Y5PONE1WZPgjj
CddEltXuisPyF+u4yd7VFcTt+LDWbuxCCrFOjyceDCR88kJeErlsLMi+ddba94unjOjP1Msp7809
UNgJLzp7gLzi0k/BLvwO4IVFstqUFNGOrLMo8MoMwaMM+Wq2efvaJhB/4QYozWUj9lzKkS23d+yi
x/qnOIx16NmooxtCwCmyxD9IBdl87TydyM7DDQVbY41pwaGHpguj2X0mT87ASOTHVTHYkDI/14Ny
/RYsEzUAJRN1D9ClMPGbHoiA71g+rd3snak7BQuht2bmLkJql93iPZgRuAC/1h5ZGboG269RXZkO
fjF4k5fx7rBAq2EsnEK5NAWe8CGCUEEuy5ODTb3oAxCwQ+WZStFA3BP+mOvJ37ZKf5Je/4Uw4DUv
ivd8BJlQndXE6t2lmMQ4gAcaC6l5mlyaEe1rQ8cYRc5FCMYkN6xpRJn2gHKnmN1/uWzwzuezXAQR
SNsM5w/4HpwimnObqkIXeVMsNDRCVi5Ir8NA8sbP/a5rsRZIHJlezSKNS5Izry4ArMOnbHjAp7Fz
8LQSuJSTtcYk7gggN1MOH/LmFSmA+4lVqL36AT0HnddAKQ+GVxYEiRi9B7nqDjdpLy3pPhylqQYq
hEmppqu6rOsJjVs0asdbW4yqDX00gAqMCFyQ86y2KteWTPpNGb11ZmeDNUYkZFXENLGUHFv8w4N+
iodf8lhZ0fJrMWMg1GAYb1oUIaHszXCagzhnd+CpXEfrAggLDkIh5SFDHn2nwNKQtZtAaFib8YyU
PIYCUyXgWcPlBOPs1aUpVrVjZz6YzRXLDz1EdanogAxXUI+JRPVps9CI+yDnOZYe6q0+7H7afIRn
PbOic6LE05y5px8Nii31PicQcvaoaFzj99tuKB3zkAshwugUUeXJhLhmwIvCdoKTRmWfa6SigOmG
ninOkWoulwvKPx+r89IstL/YJ8PUXTMGxatRU5hnuav/njqPREC0WN6bRHlB43HQfDTUQYlmgOBg
9TNqhb9YwdYaS+0WpraLArBUlqHDiT25HLEHZ9u4tTshFtwHnS68JtZEqFTK7yECOdGe739Rn03r
uh/nYoFaWrq/anun0zzb+8Cl+Aa+HCsgGKMlimEyj71Fk3E+TLyaKNOdGY2/5VcW+J+dLSj5TBxC
6a3TEykTaHpJ/CsoLiZF5DQHy2CBYNDF780hKP4cMr2NJo9a6uGKTF7zKSavH4i0xx1Fn4YUTRq+
S6n5SQDXpm88RUiaA65WcKoF9xvqkdGpr8x32gHMZk+EV6EHBU/7c2zxK43nSiB5rOlt/9BrzQqZ
YRritk5yyVlcms5P1SU7iXJAT8d7KFa2gud3g45QQz25jc3unCuefY3vV5zTE47OC0OcXh6VvJ1z
kY/M+ANibvMMaas+bnaYsFTl1W1Wq6vu1eiQ2LiLFh+cFpuG7TNQ2gROxcksLfNbJMJ2MQodwJTe
WC16+f8KpmnLl/BL26Rknz4l7XtPvHtNkX+ZWWzHh79cruiH53LboDvWT7f3DNttTxxRF21alrr+
4VCpkd//M61Yjiq78OLFFL7ZeY7ET2OqaVaL6WwNvNt45OTNAKl8okhhEGWoANACOCOJ1z8SMIk3
Z7sP2PWsZiaM2KQPjWRqrkLXArD8WZ9TTRG4OVGnCiTqlCOlrrQdsoaePp0dzAuxIOHFLN3SXsEW
xBoWQRr9LEw7fZzJoGE2bTCxNT8wee7TinZqlROpAxHZNYHLju/nnHl9NAC6Ix59YdqpLx8fbEbu
vGZh0cTgmwkb9gSU3EB+WouesXQhMTLTRlt2FtNKlS4u/xZNvPrIvOwrF87vu9s+UPh+xSKm/H0O
0pFLKWTExHHUxyfD2z/U7QHqvOcL9B3mOaMoBSgF1rUEiNeA/OAxwYqAxCnRKcxbk6ea29L/tvkc
vwsMvzThdmBrSr5aXd+Sr/NeFfSMXTNfTv8h/YalieWcMfPdSk1MsnztZs5KpckoCaAMyXkDCQjM
sfvSA5EZ+iEt6YZNfqV2RN149fFnpXGKlv00wk53yHRYWMxKFeChMI1T9RTuo0bp5jS/8JOajZA3
9vM9WxTWgfSC15cDUcPCkaZYX0TPUS3fjEjyAerDzHOC1wx5pSWp3JxCMkzABtfIiaFroCoM1bAq
g3iJCfkm4g+yFYPAL8s1XmkTxjfbQnn/LsdGlvKMTs+BppHgoUhP4HT8AMJEs0q2c89i/kAZ4YsA
t5yNpqUETcxoUw2irY+LGSo3EQ641lK/MAJdMHAWm0hgun9R1sz1lZ8Gv66gk+GfxGMbQx832jyS
tX/hT868iq8tXK/Y6Y6F4+LqoMEZ9+0dt87oXF6bs/IjsDzwbJxvqhAFUCz6EfelQ0SKJxyxz1na
n8Z6i7ZC7jFqreDXuMXzHu6MRG3e88PxZfxq3F3gw9uTbhHev7TDc276tk3H1N5NdpXVOgYDMHkE
0aAx3hjVJ7nmticZzGLqgFKf3RAeZZ8fcUHXTiSDmF7EoKTC/fI3sThgu6/bF4M5aG2XcWUyTu3i
kuvy6a7yOkD3vP+2TcT11/bmhngqO8fLPs2mMRMhyiJPQWRPkPgvLWsgwdVNWog4Tt1o9vPRonqo
kosWVjTYW0JKkiuDP8PnC/LlyGoDpw090nCff9eNbdzwWd7Wt1ANdprwdTKpNczQciMA2VzJGygB
HzrFFOytxhDMduXqFpdgkpFXDzrsUP0djDGzbAOoUASmCD+6tltiLiJBiSCZZvwHbA2xBH8e8wIE
x7/n8dWWSOZdbnNEvEBgmNjeK1oRtuf4eTZdC2u5Oa98u9DVJcxarEF5TwE0WguyeJAtABZPlVK+
aFm2zj27HKVFKfwHxwQv52YLQFZPVUTxEntfBuCa9GTVaAFd01vwRFvjmkNtSEH1KB2y9gNgD7zE
VeXIVIs/djDFFYbZzYcUPXRUDbkJmzljDmRV4NEZy8AC0ngdXWjjnKRtEC5cicxLX9EBai3den4X
jftuI84yMJNW5wt8E7ZIt8N6ogXOlls4FNMW2qlCpgUU0lI6uwNOO6WbH99z8x+hC2NN7ePyg8rp
P62oW2p00vBOwzzfGITU7Amp6Tr9dxXz5rNZQp6rX2mBX58/viq+Gt28/rS0UHHsASsuFwBiFkmC
L4qcQ3TAvVbAAmFA7y+g84fAfS3pE/t9b42qcMlCNUxXVz7Cao5nND5tRzkSiwIo3NKKuNNpkyoH
eInE+iGYredDWo6iT7NJ6p9qlhsHtjmuRvM7GpHZIM2sxi/T4b9TbNrgIjI6jBBjAc0YljTvRRhe
0xSYNBVSWBRYRdbcLYyX50pFvB//Z2W34YUI6Z2EytfGgU3Y0VBWEqJgHVmOgnsAbb0x3ULgMcDc
DSEaFfAtBGM6E+tf7NWTxQf5hlb8secPMAqcEg3kLYtfyoKSHCyk+jAUZm6/52Dpc8xy5TsNey7b
oa59CXXs6WXFe6hStFYuM+Topl1M8vP8Tn405eWabDVgvILsy0ho3+pmTuxtgPemV9uXTIbCNnQ+
VfTyzipPiRlBjp9csqM19N6yriAIj07BQzGccPjz58vvAlbpZftKaQIxqV3RbxF9qWorojaM2ljh
CMOIR9HyVp65WC3ltgoRth77pJFPFMHWmM+7Iar8T7zUwndN53lPuFxO7xw0Kt99sZ6NlzYnBQJY
d3TyzaRWngN9FguoxCmH3VwCNFAISvo1e3YRNOgnLMmgrh0EOom/OcoUROgsPTwnYY5G8/hc67Bm
ZEWVDgXgCExXoxhdiL+LxmQsTjZxzx+mjwnXZxvrK9q75NjGMuzfcHUazad+d0goRP8nhTtffDPG
w1Yv1XfKkpsIMVxSDMMeyncgFOUN1yRF1RUQaRxOkI1cR7Y3bYTxiXJnIWT14oZg3R8CL6nWpakt
HqKiegZAmkgVjSYt18DjQUGv0/ma9YFxEqPpsOsz4Y6QvWJto6SXQgJCQw6MAZIcUO0fTo5AcliD
OnaTDWzAKu3+wSswW71eaGODj/IihxYXprV/HaJwT8oDqmSvG6LHXbjM5ptgLkNHQZQP0YGWNLFJ
o0NkZKX5yoeXsVZXqm+sivbBbqaahxLxAXd7fCJf3a4CKyvesWUSfTHHegcjxphhQdcNP4om76MA
g1WqN8dG8/bg9qVNiEhqa+7gGNFFj6blu05H2wNeN1gIHrrpfFMMZdt7y6+A8k6eJYS6lUOqigZP
M/N9Xrir2GAgFw5MRvM73TIEZAHWYArQYts3IAkfANBIccSlMfTN0o9v3bS5KJ0vij10uyVQy9sN
4tXH7/eYWxENErIyCizTyRG9DYnF97geQQnRIYD+8hWlob11AyATkvaOgPN1RniGEBGqAC6bFGrN
ai7Vbuce416DzR/19ZlmtYjF/YinN/0VVZ839Xs9W/Qsa1I080ox7ASTBhtM++VnGVaE0z3RgWMW
t13Mhx9G1l3SkcCfi+RX1C9N7qXjMkzASuT7pA5dMRNL5lzqG5w34B/r5S2ThXKEnlTRSdXUDfVr
whXelrgC55bshIwPyNZswJ/pL8oInYNBvNgugNOGkNdA2k6+1F0/DWPhF8ZT8h/kH01wZp5nsnZY
NXyURBwGHTQjQTlZHm5YQlspQyzfW5I8SvAD7uR5Yi7FrZ89xzyoffDTM8SqzBs4X4HTeBH7kneG
KBDNO3Yar4Z0U2lhWmlBpO3y7ECykixM9/yPYVEe9alZvMfQgX8WX+wQaYJI3pcFlysquaNJujeb
3C2LvYC+2hWje/R667s8Hk0fJsU/Qh6vTmcHRLy0n4qzenDQK9G0f0uGKBhg5AjMm9vANx3iVXNp
+0uYZlITSI5AsF2J8dtwwiyHl4mE9peH4M9HcbCjnVpfOg5Hl7amQcv0r8pc3O1KUBBpk7TrPI/n
QGJyynz9SFcsLmbKml7qRruaSLWe5X7XGFdGOY36EM8aRti0fV4118iEbuv+B74Hvj6mVv44MWJy
ilnrnoEtB+hn7wGbH3FWyDPiqJ5VdRoeuE7GUjZmlSwvaeWHZKE6t91J7YQVUOwMXDaXj648SWPG
uJWKsyMXYN+3EekygyFxyLIEkS71fkiMsFnnPDzPt0DGsP6iqCWeJ8sgj58cfJ/V0j9LRWWcWL8R
0cKCuW9cRxEWPbH2LB77F6jNprKoV9/jaq0z/rfwJGDKXzEFCVmZ6gpak02nz7NwGwvxrvSooEDD
P/Bqn5Ube2vZlzO1F+sjbGnDf2FDJPnbQHyYfwthk7p7Sn+emRqiMT35FJvGmQLzBVkV4FHi6xj6
A/rOIYUB6kLyoNdmpNWWsHCcBMH636ORAbJzy6u0e/1xmLI+ZTwbaTa+ck/J9EoTEasmDwMyoXra
hGQnOWwf8c6oMT0d5ahkmxjayGsMxhV7TgHbsKknqmIjmhOpe28BptQRBnoTwHidkJ3Kkipvi9/N
qkyddjVQc196NIAvgt3A81lvuD0rP9YgnJtBcvKRFEcdqFu2qXvuz1ROhciRfuZyxFntAtpHGNQn
36T5dXghPWJqjBRxZxK5e0lVqri43udYiioTLuNGxG+eogJyOqIHJtgdh8XRdqysanGCkI8qae2t
EGVg/o/XjUVmy5ZDzF+7K5ejccnIdLvke7JYIJyv4UxlYBWPTuDIM7hrudfL2upqJvLR4X5lu9ML
H75DL03LXvkpJ70uTyjctm8s1FCG1s8PKrnsTKQNia8/lkAUIMuzwexZSLV9AfkZUGLCJVkL3MH3
IpQaCW+umBlxwGFPKE6rfjIN7iA1e0Npc0tDlAkzPtEXPcevf7I2rzQS4ky+rjTSQnCBjv6aZKFn
CPJmgTU01p1qAEbcBFY1sxUYd9pM3SQABPGSrn7BkfD8SWSTMkkH+jVGOwpVND7hr6Y66Y1vioyt
W/puSgh17aMhKZ2asOFvtw8sNMKNctfre7oRxGTGLauT7Mao4Mbeqn+o0w+SrZGKGZk6M1iyuhNv
YARS3osa3HOGwVdfgZjU1EnRNwJdo11hmXFjU0OmkpIUUq111UILO49wLmqjDxqUimrPzBz37Stv
IdGjYx7ZV8JNVJPgqToKYur3K+QecsZU9PVt/3EUdzd5iRQymK+BXbzAgrfU5qcEwyuUQ2qerGvK
YKA40mV6uNIGpOuW8TDsGccGQndOYms0lXp124hTOWDbbm+h1uv8Po1a7H0fSJoRVCsyGoyZZPO2
8u3QhIasSBxTEghGOVq0q0VxSIGDsElVQH0bMZrDoSA1xGvWp/mlo+dPVvr3J9FIMx3qfntMyOWt
FlYaTmmDQYMAQgkd7gUfV5T/TJ3uZg9aDqVUcoWZvhpJE5vwDwEjZDp6YyPmtnWXU3RXvsx4ImwR
qX4hN/utIT1a5SwQC5lreb+G0nl0lU9VrkMltECvyr5Mo1oLdfvyOnMI1ZkoMpK52Mo5eo48LWim
2Ha1GlyaAvyV4iURQiwyxvkPif8iU8xmi6zF2lrTzKf3JtSpWR4F90eosI6lYutLNSs8+ejA0ItF
ndfBkqKx0FFGlLYLr5OXGlgUS5VB7zRVbgAG8kN8WTCNWXmB+tiW22ynldhG0KYhG6PsNeNjRXEa
EsCQze2A/RMosCQou7YpsDybrXcKYOOc9B/y0N9VESDhrdXDipwCiYz9fvKDNKoKjTQ5acA1GKOR
J08LY2kQzvf2RBge9N6CtVr9WcD6NYBKrurXxFAPjhovMCH8muwXcQpAXexbYQwuQmNOk+QvHbG/
5SUim4k1ycaKodAMzv10LrANGtxu2qzI9HgeKWfwXoeMY3ejom5XcdyoF7LFlAF8iLUl+3fiLZZl
RAmyXhZHWWnw6Ho7bNbmOJurcBOqeUjeOQoLWiwDL9hnqD8m/N1qFpoQ1TP7ge6IqMCSYSjJtYxk
E2s7OPDU3MfH5wocFsosktU0G+vVfvDUYKe+0ABjfCHPbZD1JCAP2QH+ti9jzEVu29FNh+LlSVsQ
Viw6jDrZ+aClIeHctGrL3yJ+bpbIKi+CiUBKsxPmsoLTaz6QlEUz12hiwJfS24Yu2vuBIdLZK5Ht
kikdlpUqBXn4NWWcAAC+KBlrfKxTrkFe/VC2CEGELIiQ8Zkcfz9TF5Y1MAkCV7MMQQyUpQF3S/QY
fAH5OMTsIe7tv8eSC8WkjLdu/emXnpLwcZRJJdYbaEMAzWZfoVu1LDDMvLerhcx3FW9TFk0yoj7x
RQ4iEdbQYeYTsROVud9pMSmuSYVnKVyiGFbA5B4b41cn1PxaYZHJ3su1olpFlu9QSF3+SPTXBDAh
TkWfaWapqa4+nVsu6+luz6IsFYkXxmIP4yYOcPjRIy2P+IZ8hlqbazFKXGVOOxZNULLPnkXYOxWB
j8Zub9F8sPZlz61w4JjBysoyKaY7JhoSzOap5tQ5TeYQx5zP+xD/l22ThwhWvwMHRBDspmJYiKoy
nQNgSWNtvlmDF2WzSG0FpeHS6aSabeJIaf0pFlvVbmbftuXeMQZpfW/8OEjB1lCX+QgIBLKVa8as
o9l+EwM2Kj8fAbkSspSs/w0IiJKSnZ8NYCpyszIyVLD2n8/XrcNW2sS9u4Dh0JtGf+jklwxPOA5p
vskgC0+L+QwQrLatRzo8uU74aOi107qiAiW25pp7F1JciQ6GEpNGeBDgBXrosEJnc8H2HxFTTyGr
s4tGKauvbjP5l6Zlb1yD9iupEd0MqWOi9EM7XOcgqOpEDRcs6TyzmGv1RLtGINeuFEplsBLprMIg
VZ8CzIoiNxpUiDpg8AVt2aMLylTV7Q9KbVwR0T+SAKHcLrF/MB4PlLtPlnY/T1KKtKJfWMy6jowU
/L79sdjTJ8lh2FvYZWoGED6JPnaGEFWKu3mv9zdEM3/JywSqWLeKcvD1Y3Ms8rxIMKD58IP8R7mh
GLD8r4eux+m4LnIrvBqXrIEZpxupfLHD8S6116MsecSnijievm0iiJpxsYZA2wNKaNQXFKKEc6+j
8hODXnT6hkn8c/Zpp9TE+oAh1oVNG8t+2Rfi4xAmrRZ1wklFumXXUyaT+xux4b+oS6xFG/14T2X4
aUrDecJTpmx33sthdY3IqjxraUlvhKu6aFDLE+1TqMunrVEEZKia9K1rGzfMHVhos3qHImk/Eth8
4CK1RGOgoXd0gvxv7v584ARZ6KZaf97+o4eEfSBvzPxqy5UlZ1RqRWzOzK/sjS+S3qHe3IPNO1t2
c3LqoHPBBNKQ8+XdBFNAPEB1X+GP+EiUIo0aJtRlLR3p67ogJqs4JoLJNfrDxSn3cQPTB5j1yVve
iEuXmPOwlFv88yq8KRogh+JW4RZCsP8l5AA9e59WoHutvt/uyBkhKNvugoJrnLyrekCaqzd3pqpK
I151WRzir47d85En61/MNXt7Yn+GuvtjIHwVRHPuI9KEWBUguUMz8duM9vhkBJo7aGfR+QywyNgL
RAn0WMzPh2cALXwI0+VkIY4HdLG6jh8wQH4aA6Qh04GMUeDY970XclzBHfihuLvCaRrsVOiazRW8
UJY+1zeGEvqLy6a3NvJaR/0GRjj+32H9v3qbRz2d48N5HY/4gwjzKq0fHcmJDj44N5zhvFf9kCV7
ilyGCzQVKjKXz3Sr0dp+8oS5BwOrs7JAHlsYTqlByawAmbvhLzb1sEa6bMQftKqH59CM1Pn/aMT/
hhDgW6rO86OBy5Eqrxq/rl+N8VdeXQ+syQ/mPDs4/YT7Lq1Wjz2i7mocutKfQxmb5j+Suee7gWcl
Lubq7rQz0pDnDGp3BB0fWPFo/UYbeBH9C6YDG9BRQ25Hcdm/de7p4LwEB30oissKon4YxHg2IsB1
e9y6wIRUOIv6IjRQ0EKqIEj2BRezbeXEPKU88heuUUYS4RdLfwH692pCfhHXZ0HVvWqj228EjrYx
pXZ4KYnQMQnXsw7N5mIAdGFDg/Kkx7Mbf2mnGpIOA/c6kwuN7AzLNze2zjdkWYXkju+besBcuHMr
rIySY7LrjIvbu1GT4XrkjoMGT00s56rV6sCEnv1IlCUilfn9HGvxbLuIykHr7JmMrJuqLStrTa8/
ubT+UrdPE6OK1nrG4XqhB7vJ2LS9llagjTIoO/viqbeKWE0o37mez4ji+LLxO0K0XsXFL8zdIf07
4Lfku0FuWmwR+O9jtKQVVDEf8EW7TOLf6bvUvRIxyXNnY90nxaHea3CvovjtD8IPw5ddD2+kBeOU
dGqYLGmB8UWg+np7NvmMabMZGSfuDGksQfgb+h/pBkpYBK1EG1JuDzKBET/JnVxf27WN8xOTinDA
ybGKvPb8WEpKX3VFzS0B66dNbMhH7CcLZ23vMRHatlSdpp/s4nRegILIVvJllIimxAeKafnh+N6c
TJZo2lpLUKzEXp3oQDH3HQGeY493oMHq2t720pBnTx5fRMz1MVThy9725Vmpb/hfse+bscYLK3w8
FAvNCwZN8BC0TaGD92BS0Y1fpekpQqEPyxn3Njt3WIbD+lPPS2oIt743MjniAA+4gLAr4hq6jLaX
er3fKGyuxCs+cTZ4rN/+Gm/wiwKNMma3GXv6RJ2txfEfUIb1gzr/KINsuno2jK86cHzmLBkPQB9S
6Jtp/rt0CjkveLzcjo5HTOpGDAEWtqvcNtxXAmCqGsaFoVlguDAhamLb7F7WuNuit4VbWbvG/2DN
/GiE9wA4sjQVsPT7SuhrvVrLu3qZ6ck98Nvu/RUVfw3VXhDxsFm1SyAgaRxxv64lUiALQt+O9nM8
3xMSdc3WSAJ9DM+qKBMVDCGRkakBJi20nIdpwZO60/hN6F/0+tkarmSME4YHSNU2b6pQVuF04JRk
eZQSgLNAc2o3SJfWrp8wQEnAJvvsvKqcD6H7VL0EPzFTtQ1tb6Hnv3s/G6FRC5sPD/W6zQCevWMV
duZxvMG6fM36VzoR1ZiVW9PFQoVGDhVAew7dLzRgHTVGS0qBYAgB1w/UAdSqbNvXh7xXlX6McbaC
att82Yjs4qbtiX33I9qp3/QEsikpzKWp5huVjPuU16qMGHmO3InaF8gC2PE9EdQUGvG+NvrZofSp
UtO2wewF6jlOatWGdkP2Yh3pQwtWod6dmulbawZ/5MPIINDAlqG9DGSXKND7x6h6NECwty1Fr2gP
29ETuIuG26fSKIjOVxRY+l2AUGLVTeG+f2ZsT+NoQ41MUtdfv9CO6PXL57G1ga8n7fVtgBwbCjuB
2htgLyjMSfOvPz8pTQwB7xLPvAh3VP1jgix6J4eWTdcxm5BsXcQkrL71K3+rLn4t6ygOTwQfUE/B
wzVhKWzIwSaFeEyPDR3RUwmeue88Pe7+giG6qnud2duMp3aLVlXmGMchg2a4QF+lH0ZAmD0F7AFg
zgS2lVj/4VtPdyeubZkJB6skwzCJuxWiWvh75ufoifZXQqPB3VeZOhgh3tqZirUoeeuR0ozbSsqW
d03OSLcI7H02SkaxIlib8tjJNK2vBnK4O9db1pq1bGe4qK5BPNBgclBESl+pQ5/e8h74ujcNWRdu
dqzGyfciuTy6JKJaLUgns0hrfzxKDaYr3nqEC5JAYhK+0bdqVeXkpaXZYq+JwERNbtnxhFpJI4hs
UkPGBatWmYt8K3kRSEpkrSp+vEv9ncZvQsgN+m7ctP6N4OmI16P0h7c5gfCzbnEb2mrltMHCwDIB
j9YGGAGl4C5nsD6slDLDVewKlAlVW/9J1rTRWJ8UqIBxwTmOIUJSHAeH0NYDj239gy9J/iJ9Fp9P
8LQ1pGfbLx6lKH2+Qphxz8wRsmGOLgAFBVh1pKncKaPdRTrZ4urhLoo/3OnGs7ZaJC15Hs8UsSUg
I3Fwg2S1IkhijSd/qrcM+YrGEVdndQhnQZ7unqPyAbp/gUFqD+Ah86U7nYkRMpPhaWErZKSCFn90
4oxSBo+yE1lXta4huzaaZcZ/uQUV79as8KYdwD+X2ewezSQl1e44SiQEmKAZLVWhtzAKONrlXeVk
J7si911Xjabv+TzOaQ8Ys8qK4Feea/4nnkw2HkmsuMXO0/8r2zQwzh1EKizHrI6y9PGZ7AJQDLWk
7MBfl5xmc3mAFP87p7/gkjuMbHvUcrDCSsmPjYNmgecNnHZmaGqahdDNCNj0R+SLES9jeflPLIXo
jY0Xai22jEW7QeUoLldbQCTaQ7jTWPTJ2mGFtTPAg+gNOU1KFxERXIvgwzFICKO3fdZIPee0i94Y
t9r6vZxxvoykmu3MTYP3aLFKshqx2fC1pIpVi+XC1I4CIi8/DwOg7ZKRnR2yX7cedtpfZ4IdhsiH
2biHr1l7pLK0OhOEtjD8ZNBPWBiO6pKDyfrvnI+ZjHNWq1PRXpxMUfLEPDJ3u6CMwR5xbSk4IqcE
szQahCRxID6xYMn7qYEPTjkENlvkmemxwXqWhIygUR4JNcFXTmdCWrnEeZdk0tE0f/m30Ga/yfb6
vSleEjuU0fVX21gllZ8QdPM6uor3SqRxRZZNRCHD3AlKUY8JrjsNpKuIz95q7IaZKcU+79OgPem2
+Yn/c+lF9pcMLb01epo+8+97J+cqei5zwoOlKgnMM1b3diYnPrs1FPw/92pOtVnPnWSZd8tiJzWd
pFj/Vx6YwpDVVuzqA1BaLvGGUmRswDGJlfE7vGn8Ti+5OIeARLJ/fOn/9vfK8S5sNYXKVa0DjcHb
JCemXzXnvSTLrws0RiPAdwZ27rnu4Q7wwwQvilDBu22hbDhC3ki/kpD+/V/FZKad90a+dhhajPEF
1pMdY4N12jbzeK9aNLrXi0yVcFj49P2hDlPiytsP32AXf3LHWS6efw96exnxDOyU0Ce0mxpNcnCc
/zkeUrbt0i+8qBRG6nBIFRM+s/mF9u2wtEc6scf6d7IM5ZHhVeAQOay02Njd5M+1i8kDFfTlgIEs
2s2rWt5NayDZyFffu0K5u/Vr34eO0t1qB2aD6pXqjoV/j2Fu3Of9MnzCIA/TYyNsnkl3HMB3/7/0
CaO+Y2USlRq26oDtUqZTG1RL9LB5SIgogbqkJGcKjEDiQSBSBPnga93sUGxt7idztwveprKkihVA
sAiB1RP63/t4prv/VbHv5ZSukWSc6wjGpp1BsoAUryBfo7p8VUXFvRQKIowk9j89m72KMLigIaR3
MZaDDBA3k1bMa4CaadK3o5slHZDzuxcb/Ac42dV+q587ScUurRayTGARorD8fJcO0QApDoT/AaDT
QYM6cmmS1FoQ1nytaXmPgSPYrTDlPARa5q2Y5CIEHKnuMZr1j0df6XLiF6FA6NQAdWyFPcKpJLPD
sKsgKq2OJoa29KbW6h2XGU3tUrILupTUv3c3FBvNepye69Sgnx8XjpvB2TR3XcRv+kLw1SaUyURP
tUZ44TA9cOUcYc0EAqw99XkdfPdXxMH5wZ0lwIJ79Nhh62qwK/wH8YxXpaw/at5xz3ehKACb2SXt
w7Y21le1THSWCRkhTaThU1F6Gur6Xt1w0b/3MW3ri7qtka+NuY2JblARvT3xqU4KbClHWymZJZx7
PhPQklqvKBkIosdHe4tislQZsGKNoSuzxLpriaiFQb3Lu4YYm3at/yIB0jOYKaMLuKrk1LSzAWRX
VmSN4Ag9WQL2LbL0Yd5K3tIg69GJ1iQwoDsnXwnLyxhH0pYaQ/iYKrZAMeXfxGapUKs0eC/pbS8r
cRpbfITGhm8Iz7oXCRx26I/cyEJbArEPVXyKE8cdiwrVUPQ9KErHQklIdBF5D9WOeSDxptFDk5OV
RPPpWqxDUI/4wROCYqLDiRLr5H32UWdcx3CONr6C3hc7Mfd00rd5Za2F2Uk0sLyP5ZeK3H9OujKH
Zkxd/cxw+pwC8v06h6ovdjSEAKlgFm6Dz9gvS0R7THIfqyOz+GKys0v4CLksfTCIdQYMGmOdiz8v
VSJBEjsvUnzYp7skJs/pEFTWLF2IKUi5E2FgSCB2L1DpCIPbE3i7vsKC1075F+lZjiTngsbDqIL4
3cpfbJK7hWvbuVv7KSF0RDKv31EzrvQgoh7Wtnj3XKvRTDmmELsEVkm6thK5RLSzG57kJXJWrjZg
PuhJHPwzU4CtB/XEebehmzJxkuPPpiAK/DYUmoN128IYCt71WP7WvK7UftXtw2GnOe6bgHC6VAqm
oOJWzdwiIBRssfQkVG6u0XAi9fNRKR5mY+hBot9tIq++qzxytc/mI2Fu1u6mzQXkwP+MYeTiboEZ
KgrYDU+cTjX+WQ++F8q9pv+yKsbfxBn97YWebCaBALU3pHh3DvZabmJjnBLHuJX4ebc5ShSFEoqT
A8CzsMJWbvBVJMpaTKFKIkLwmiXwwZ/RJcmlwdARhsHKwzRsdVZkH4pJBIL0oTODChA2y3UIco1L
Had+WexEEbYf+1kDeF+GhMk7ZyvAzs9p7BKzMivmYF82AInnGBHx+Ovr9MgAh80TJr/HJi2c61tB
GKqr+UHBXveiykA1cQ8nFyrILB8KY3DR7iiPMSMtUcMAzC2k9ZZtYspUSGrUQaDPikeJB/f6ofit
QCovmgsCxeN3VQL3oa3eBj2QInr5XnhhPOp3FqqEWy1on0CqdairE1arZx1Hv68gy8TEzSSXm7OU
J6vSNqu/s4OkjfM0AIgRt9wd8b7Ol4CLfb8PRzlIPFnwQugH2NUeVuOXvOEux3QfnmCmVkkVLAGl
SOC8MHj9neQ7njK7vOynRS4Mgwj+f4d1EBT2hSFvXR55XJKkICeWOPGuZbjgmhbDd8JS63ifIpQg
Q07EnisYD19Qenep7P3bWW9rFdlsMcqeakUtXyBdYqrxgzdU81LljQWZNp2uB5I+eIRGAQQWXeLd
/Yh6Cz70fpwGFs/tDX6dG+1dqIZ8+dc0eWryuMWYtZ5dGViYu4e/oR4ddib2fL4LkOmY0mLEc8Wu
b3RaveOmp6y1y704bsu9LqNwZJRctOYubWxjE+LGartEKwuiMLv1j3ScEUIMnZTZN7EjfiD/Ij3B
vO09dpnQ5nynppBDJtRK3189eBM9EW9gvZj1fRnwjqe34e7oFeB2xgctIGhr1LxStA6T2b4Hquz+
k//KdDprE5S+WeWUWx1t3pO32FHYu1prsGOrqrYSFnjnDlx5DnQHv+LK3045PUK2cMFHV6XgEpTW
8ArhR/cMksz1bcU/19dTyOjtYhFugaAWJecIfM3yxq5vDZRzmPbRe10mPjlBI72n4JX/RinO75it
Dli3dZuQYOMN4OwAp4D/v/JiaVzial/VUXXQFNQs8KkQqS4QM8vd4YE+2lC7q40Ir1wqj99KDkFd
VinSZB47Nkbg27+w+B4eFv8FLo4yAYDLbW2XezwYdGuZoRpazPKp19MYbsGnGc/RkfeDtVzQ4/MU
xgXyM939kvyk4SallJ4IIDvyOAni15aeGEtkki999w0ean+sQdHKn0C/VXAb961XgMBmOx4WTrAx
6c3fQI074ueu25gPKtqeVNQqfqe91y6kE1tiWBDOjxcLq51ex9tbtn0ALvTRtaW7FcYZeQC/Ou+K
1Uhd62lZB9MzZRhYuoCOf57wVt1iUqUl7vM17wycJ9D2Q4JQRID3+ZKGQjqVuH6SugqCia3URqrd
SRWHZW/yGdPYf2gEi3YcEiYGo3HAmdYdizmQs7iIrTnVVEvrdUSnkFLFUnAwpvIjfZDhTv6CkzLZ
4e3lrFQPg0KWM6n4bbyTfCIXtwYO7j8QcsN8+a9vQdHhjPA79sznYDhDyFlklJbzY+d9mLRAEtaJ
+io1FLDsjQsMWvKaJurcy1MrqUT3I04hlljclipkVDigGpi7wkdFfaN/aRj3OJQOVbuTk1Smb09C
JV/QptIkxAwlHjlZ6IJKnaXnUw1j8SKN8IoFWCokN2LcuhVD221QOYW/0Lw5Ai09dtJzazgnNsRS
rPAQvSrvWNMCcsSFY/kHrn1w7D9pE7C7W5ByEEN3J4qg7vgtOdGxuiFWXcC81ntzZ+OI4HRFnIqs
zt5oCHEDVgIMjCce+sM7tIhhwg9mTNfZ9iJr+KJtbOOa9rDBMbCXZz2MNRcjMPKIVTW+SdDf1iIz
Hx4kibKX5QZ4tli74zWAMklgzVXnhjzr3WhIC4wryujRDZexUGqpFgLyZGzDgEbZTW+Iiy1Q0iJY
bTcthbSl3prFmJnzhtKokNoYEKYURGb/0yrvgFMtKBqxQSsBqKQj4sEZCTqmWW5z7dv4SB+rtpov
6G0sKaxV8PDn4tDFwymPDYlyk6HH5eHlNaqGCG1U7UJeRBuEusvzNzXOW0NtY7KsSbWA4xNvysSP
7etf+CWhHGrGYHX3IB3QDzolLofb5QApj1rXUM06MFQuc/kdoBNEnLgTDaDrijNRO8+v4ke7Jvtm
4isK2taWwekfHwigtDgBs3/wQ6wtyiOe3V5L0GrhH9yMoRkjT274d31qwY6XSMei2jY5fuu5VUKa
AfyP+9Yds28crXIox0R7zAf0+FjZ0T5O5mb56+yoXJl+3MPYR3hfd/c9TXD72g9NiSAnZWQhcABT
Rp/N6DUXyca2ts74zwDMXhBkqqb/0xA5211EHB1WGvO+YlMXC+1ytb06aTvkLRWW/S35+Qha12gz
Upm5xDiyPPoXhLpFlJR8Chx3Ro+L8xj/E3ObJIrKrCkq+I5JAsIX+J51hObGliPr8uO53zAJiPeR
tdzjuGc5Ufw+kj9BmyhmIzZ2mdod1hfZUkLtvvH9Z+BLSmsWPMQ8tGpQmlf/thwpaHQZDTA31O1J
+v8/MwAy/RSGZJXcLEqSnf42zkITymLUx5THaQxLXM2DsNs5l1kscFihQLIUEEKIRT5bGxxCr0Cr
/LrB0BBrvnR0hiLQ0bIOwXG+RNlSA6ZydPbCMlOTl8sKAZpGhDNAvXaTczX70m+17fJbDEAuM9zE
wbuTXnMlB0Mu9eHh1Psf07eLDRys4ILfWYTTzKM3MN826XBajhKQZCMR3rX2mcEtDkp/cdbaquB8
MAl1dOiwRiV3+y6v7JVWL4tIUg2YkNVijR7W03i3ZYB2PNDRjKeKNaBnOIHxkWvSKklvdycNLxEc
67nz68yhdhZQ5MCMpony9378KMh9KT3V/kZTNpaC+5OmBJBQKdwCJGdpusI2Xr8abYBjz8gyi2gT
X7PWHO0dBw/WqvR82komkB9i/H7BPxMitCV248M2wHXmiJKKOPszgSgb3SQZnpLeRnJOhNxwRZPn
itpFPfMAF+41zRLCxZSksQ2Nud6fO/7J6MBT7l0H1NTfrI8Aty7euY1NHAIL6KBKDBb9K3pEgNj1
d0XAtsQKp9oEUtQYs21J5SX5Hi26VZjLrEvrpKjWTutWHmnvMdFVYi95tyn4hlCFFFehLXo1d/UL
bSXiDYxqwt7udynVUNTPzv17yapPHUrq1ERQE/XEPZMnWrluFbum8Y2MkspIEAYbmVdZLXW+a0fJ
RNLlQacfkN3qAlLStXkJQcbTXbClG5As7noUPOrShE/xdweAr1LgLJjg5F6A5ZxOpdBUdMsS0qdc
eLpz4b7UQXqBMbUotPfq7XxgQOBSPYl7zQEo2wW4reOkdzMZL3Cmb5Y7J7lSYgnKvevdcTkHXZd9
TCUHVCAvQfFFqT1g5+prfJLBbVjwcDf9Xjex668PncwF6/ElEq0fkrdxeK0IKoBSzoxaIx/pvuEF
6ptBg75CrWvU9ehaHVKz9GEJg32h9tKcPcBcIBaHUOkpJuQqTi15RMpYx3bhrSXlKy+r0n2uTmUH
EnaCdNrVxIA6O/J/e/SDkf/y6Pr9YqMIG80a+ilsHYQ6LnpTs6elEJujKOdfFU4IGjsWI1PEmzC/
lBvxTa/PChGidJxDlK7fY5DMwvfChthrJWoxYTDJ1YScazhxjxoW0NW5eM6zTVIrZZN549Q6kB5+
hplqoiIVRnYwy59ZPJrVDmaGDrYZXzkrGoHhgBT7xRQz7E82ZwQmin2IcaT7aWZGTSB9xUqUa4mX
vjg9iAUeVlupWnvSL0/5o1KvhyeST/5U4vSMVREkx6BQs1ukmzHgPeZQpRI4P4L+FpG2c6u8adW6
zumte+VkxmnJANyA5r+qA0/OyFR4DPLh/m/iD+opkfd+/8a++PoK/7KFSMhrMJBAfCKb7/kA7fQS
BsW6t4u//wAlhRM85BF9O7DsKa2nUUatnE2Fi2fHpNa2ZuM1QuIZXvMI3pYRwPG12cmtTKONio+6
oz6t3ZmfZqBv4pS/FHPJg5EXNd8Ivp98BEHFeo7X+DQi8tVAlRcz9s/weWoQFLsAnWQWctuCoyHS
hQoPko5gOTIab8P1OKxTrcgNoXSZebm6urmJoV1aY7Q+5K8gHZRnj50ERG44HdAZJqRNL3lZ8kHH
h371CtLYWjUE50ReA+DqvMwG/vvTXQK9/RHAyyvk2iYpu3spiqRKOpIzta3Aor++IAvYx8qucSK1
wlY2e68JzoqqPez3TC6YxCReH2MbUarQJYk/6kcm8g3vPCKlvLYO6HJ9Gk4v8qmwj8IRnABow4Ui
8O5wZp8NWqG2T0fSlD+iTuV2ZpUM7quKUp0OPgLw9E4/9a5XLNLVi/CltzzFo1l5xflx+M03I6H8
YOprA+C60/umbAuE4MO3uq7LFa6Owrn3alFCua7bn30qpR+yQHtitURxWvKkefvdSYm210A0zcG8
WCH9TCgk5HLuYYctHqIM4caSn0L7CjLPME/hCqxe3WkRYb6Oz/P1YA/fWKR3KYa/10JSu39KeKLv
mYAeLCB+/hvzoARCP7WXihKmErdBY4ByqSllYv4kuxWjbffutoupDIMGxTfrg0ts++UfTOkarBVA
JMY9ETRE/sJmntgXMHYDLQHJSfFheKUm5lE5d9cYoM2EUUDPKopo/bMvac5P7uKk6Bl1qlwA2XWr
lCvObQYvKu/PxYB1P7xczABa4ZZaEKMATHbVzyg3witX0tlhKtP1HcpKiWeHAXTfFz5Gd6bPsm+h
nwslxUPH8IHTWKPVUzFF8DNOao+5x42B/nZLSnGGKMCS24X6oEYYAeymAqvgFGbLsa8748eHAEHN
pK4ZYvXJsyw8VZpMn650IiY7dC5rPRL4hQlYB0Kswx1InFTtItxul2DrS/h4e5L+xtGUl/J5pCwD
LhN1iqr3ni8/wfemzfAJd73nmbHv47Cho2tc3TVgUcQg2RsIAvb+YwdTTS5ELZaHwGMndx+IGfu0
/2PTr8rkuHlIQ3+0zEK3NPiE0zezFmY/7sqaxtcZY+jUvXWfGkt2mXdM4VpGTqqraTO53Dwj0z0B
nPNgJcj4BQm6M2ff629eEZ5/UQ/E7jTwGnr6jiJrAANwFWOShZnG8utov7CDqT/GNKSTHbTRYhav
QXjnezqS8nYbGZClN3qagMlNZz6mOa9sSqeHmv2E/uEX4tjwfzeyL1BIU9BGVX1QyJ7PEO2YyJvY
n3sQDg3wKMKNb1Pw9GOo4XR3BXjSdneehKfk7x5YYjZL7ChDXrcCr0GCIRs4y9UCPgwqZETsmmsl
3CnIUqYN8XDyKiTcj/pLYYeIp+zHVbUnpK2XuRZUxJs6MTihOmeigNpQdlEsCJoOEThJb9H8OkQJ
W9eb6pCzhDlZoQ+xjdiYOPZLCEv8z3hOUjSv8NSQoD6pFSziQuwj2/Fw5RRS/uiFJWYH1CMWG5jj
e2NqeDqa7DIe+ymkCk6Xcs5DElBcR94Q2H1t7B/EaiQZK6BdaaQcGKtipegqa0mHH0MjuK6itnkv
dH3IndYZvo1fWR+bP/2aiPS2LNwhGblPS8BjpKPj+OH56rj75QB84yPZ02AaweGzoJ/8gWgJ4kB8
JSNp2OTMynNqlomiCymzJ8mOWL4k+EwQg+Fx2OtJb/WQ/hJgGJW4U0i3JFdmKu9uDPyZjkxIZH/b
fK6C8hmBzyg20CJiUqZQDm7Xc1PQF3RaJxJLjekM1Ff7pYy2Q8FPqp/56ZcEQB7gPZESuttDj4tu
K5/dPZRNYs8T6svCfuRBJdP5I0n6rPYZ6PA/3EK05D/N4rF4TEg0oOHrla0bLhX8pRZk3PFlSic7
YVVkJ4mjjx21chE9BtN8bg3maWeW1Am9AVhXxYIkJeS96D82MN/cUrzpAl0g+32d8WNa2xiCTdiy
qhqkgI1rg23NrhRSp9CTmxPpr0PubwcM0hGWCD2TfCeo1KXLYNqZWgFegcVPJTqm+7nnqn5Vr6bX
Phb48+30RfFWXskXISH8IsAIbPGqo/Ofx+4wUgAzsaYYj4/V3Sx6nC4zs+pfK1hoqroEcGPAbXsC
70y/yO1P6JDj7L4ERX1tlhINPBUfuBpFTdcfMkwEnoG60xzR5GUBQAGRd5A+fl217X8Ki0DwqMPS
yY43t7ZsXp36kafONQi2ijnSTtj1Qj4ngN152AbwanYvp+vvkZdwodExYOJQJIl/dVkBrkR/Fc4S
ra0gXl5+h3lvt16trVOYPSbjrTydie2j6UovJQ5oQ33A8DibkB3AiZrXrb6IC6MVXHtfELwDJpLf
DQaecyYFTCf1JXHzTylCvERInSmJMdQA3uOWZMNGqX4nangpxFKc/4aeThnD0+yH060Kk85iG9qv
GLP4jCLpleg11eVR1+PttHMywluWbnB3ZWDQVRanVaLjEHvPAS12LxR+w2ezG5DohTbfuUdpNvrS
A8AL2aVJNN1ZohR0N3gYzMwcnXKglEAJFtWbCUrVheDlyRfrJexmdbZCSAZ/kQhs1hVCT3D3ejqt
TXxJuM1Gv/0ByLSR2dC4iJf343ojq0xq+k6qt72jbS0zoHqo8BDdc1Za5cyLSjCESwBvI5zq5jwe
CUtd+G0ttgIGmWmQ1BJRHONR42NEgvT8ivBv/S9u3PtIrk64M8DbHxhI2jUShWGMxbq4O5t5RaD3
IfPz/dN90GXPpC2PbOhqchA5XCNB0VnAx1sqa1IrgdOizTAP24XctDeM/In+128ZPPTTcNzCoSty
Bqw2UdmnfBSNa3CmOXbsTsQbWckk6kvHAd2QYB2/DRac1YNhti317Bfh1iIdFrExaxif2L+TQWkA
ngwXMemBj16pnYmDmO/mCPLQcNR3qB3pYeOg2ajjjpu38RAYm40ju+w5WVw1clxtbFf4H7BzNrbg
3BKjtjxFLS6wgjCQ63UtQabSh0OAkLcxUL4sg+LqfdFBI8h3UDDHMT7SKZ7DpWUy3XG4zs20dp/y
4wqhjQFdJPKZwGPoz1byAgn2+dKzAX8p9MmUfHLiXBw1nIpvULFjhPCvi/GCMW9ERWQXQe4WAcIT
lWZR25Iizga0wNfYxAMIIsGBOgTAF+oGxpPISCO5IVMrPdKH8K8tMNLhjU8iEPgeq419f0A5Vfd3
pS9KDtvFTadKPA+1sUmudWuUwi6w8miYk1lqHQAqX2qUWz8zidqLs9sz5pR7e0jAEiAspiHeXaZj
GHFXef1j1QXtF9a4A569DpeN0gZuIlx+yWWiTpe4M0mXKZ0SUgwOKZ4nTwfJEZ1Ll7Ycd/G5EUOI
7b+/cRgogqFbE8dak1/wNRBN5tgA2+vW6bRNDVvtaM35gTKwHBC63hJIY29KDlEDbSILQvNDarqd
cjD1oTpCLq1Orl4yI3yA9+u2v9WdKMDqzMo2UzsPvhdKTR5WrFM8tOekxINgVxUYwVC2w3MCAllj
iGImAN2lrN9ZKRfvfNt4Kj8V4SCbrNdetDc12GyflS2LPODnFiX54d7qJgrLjo+QVYlNC7GvwWjf
l/IG4fek2nFmEJdmgU0r+LW6Y9Nby3wLNimC3+7b0NNzNEdeI1q/pfQnQ2EXvzN4fmAZTPKOdmms
BRjbr2g5TUHUG4i+puxFgHsHenNeGDe3NFS4QdWfz3PWKHqjllkhmLuqbJk6coV6978eA4Jrqd3t
b/bUIYvcQduzGb2IK8x0Vzgfx2g8K1uBaSCf7WdYUpJd/XX0xW8fk92S1vNRqwv3H+v8RuQnHCGt
3Rq17rIirrNDNoR5JKvAuJKXUmzkdBD+g9Zwvi/jOQYJ/biLN2YLaNOz0UWOy3mzYxotNC0r4t9i
8eqsRZobjCfAoNx6PEjOAXbhIgSXGPyYROoJR7iGQ/SitXFRqfhehPiX2sFm6WtLyU7OuJ787J58
N+mg7LEQ5HzkHI7G5kVCQRm+D77HLZ9YHbiY1XOCGG/txNkobTJh5SJshQ/d9MMffBj7awyjrBLO
FR1IlPcxHibqTEImtzBxnHDL5T2CK3jXjwah2l+qJqXUqf1NXwBUsSROh9GJxeCFjDlmkrEjU4cO
wTruKysDjRrpNlaSQyTHKqcnyTttOqIQh2gJ11aw7KGqr0hUSeT4lz8kpFCh0PLG80D20lhMzENf
97UQN/tN0oKSbYQZKUYpVc3DXwVKBjY9aB1GtrhsFHDiOdN673iRkGIJI3DrwXxdbs8va1NbwcBr
LbIQp9ZI6PY4TTrKYZ7TSK9Zh2k9HHJB+BFzHzeUbDFBa2YhCyHqShn2NH1d7c3Yd7fPZYnjj2oT
XbrPt1NIl7p+eHjh+tDRDfTV2M1zLeiyuLs+GRLDFGXVooo8peixdad9YYe2K/bU1iB50qImc4rw
VwRmN6ZdpMg/g/risI7JqV/YDYE9+P+aHN2xWMECHKA0PX5dU/M6rIiCoOC5CIPjRs9um9Az10Qg
ZNaCufuqbpXFzdKIhc7bfeNRhcpOWdjZIbbveiXFwz99vo3Xuama/u2I3O0X6OWk9cor+LO4UMvv
ADaLQTgbeodByK37LHGEzalA+NT9OpDWFwy9c4KReRVAwpjQjwl6UwTcvYX8TvIg6RondkkfxbEB
IwO0cmeIVXwB3oR6Uw+Czikto12Bpd78Hzazg5YPRwRLeVc0quWizU2yHtjHxed2n4UYr/zol9Ab
WLp62UthyIAmuEC2VSQ+LPBTnOyGC3OWPT+C0cuPUKHPUp+zg65kEX6YXzFVJb3WReGri29QaDrt
/cTOjKMPuJnba+L5JwcCxwQBbnM3eCl2TA76KlhQt7C9ico6iQBNu2kPxdDAcoS7gqLFwZg/EyDW
o+NQA7j5N2urz6aJKpkIBih9Vauw5nf/uKNz9RSaygiijQtIEd8ibZs7AJMXqpc10dO5REE76GCj
zfLil0u99UOHcSdla/9YRSBGL1ZsQWLbgeAPxiVh9MoIVA+zMJFVtVCFZlSOfZiEPniDLiAcFveH
aTBGjmMQYft2SmZ6F1KGfocklSyRrgz3X8mMFPcH9aVmoTX/Z372PRp2nBitJdHa4cPUW9jGoIXX
ceQ+10VqP73sT6dTdvt8XsDZk8yT5K1GOXoC44LEHAkRLVfhW6vV3KgwYAJjhgPO10m+tngPmqKZ
KPLbaozCPHoIEM7NIzKqrmiMtzkPvX7Lq3vXWG244yEHvSb1oIr2zPeIYdIPF+pH7XHztpXFXxfQ
/CoNuWTVSUpLGPtUjgb7Efg1iqzdkdF8YAy9Hyer3wFs4j/3d6AxLSHCjsWLCrsR77SIXTLfYwsT
Z8xlH3XLcD1Vr/PevGCYg/3AzjRQDABL06VYepWgxjW9v9DFkDwn7ggKDf+lXk++H89ZS6FYORuE
arnPSlV4YcS8le4Nl6/LHjeAuTKixPZJpkxM2yzbjopb817mZl5UoMFSz3kUF34f3y0AVLSaaHU3
b3V5o0HOBBM7J43a5rMBTdZG9wEPD65K/7cvbJvT59PbPSjNHjpTO8r6UPfqcJdLIAOqujIpIIiM
RSsLJZzQ2CVqX+qpW8cSLC2IETOD6zm0OzGyv46KhMXuRDWVBwDQhT5TcIAPNTyaRx5WDqxZMWyk
XlU3gLQCoID420su65Vwq50uVH5hg2dwswPZs8bR4Jrc8nozztmnQAxZKFSeledrT5DVfCln6evj
LlzVVF8QzCTyReBLTmjMXosF3W4U5g/O7GHHixrPi3kvlfYS32A5+W86HREIUILzSm+sqiWy3i/L
UtryDcic8l4aorxjXFkJLpT+I6CL8LNfxeTIK5LRD7mwFgQW1KE3XeNjUZW/mVpG4jAa9lq42W/b
YvYJNRyXL7E+YDGbOd2osAWt37dG4TSdc41EKMbIBpSGY2avfHFX+uioiVQqywgmaUETU/b6UeR7
csE7+GCjEYJyxt7ZonSK9mqhFUptjLp9AetvTQbnIYrotO3IvSeKwREO7zsvD10h8cAdKtXRmj3R
mNQ+Nasmk2YXVVIU/dda6A6h35ToaWroyxecp1eUboiRIFXfzO5+qfwMh59dZJFmQp2OYUyVMZHj
xe2tKNvNH8LPVL1MKo8jXoXurIpenmkq1lu2VBfV6bPe9kCUXysDDgPSVVFxOig7gbtaUJNLPgkE
bWWPxTHjLRzl3MKgNxD4Pmp2ZFZesqsbcSCiqz+ryl7MHDioFcqWxiPEKoxurfamEZMnf6J9Z+ZQ
S/wjAjzf2QZnWkVUUI0+Y/U4ff8AmTwHQTjkN6xPvEqfHpxD0uiIP42gKTvSrXe8aJNxdfpGNVXd
5b1OXJjbHbYF4coC7lXnkbGDf7GfKTE68pfU/CzoM1sMN8FZiykYrhPh1k9hdfdwLGPLlexFVxHj
UcCe0pGZ7WmcCl0ij3FgomJlOJFNqZkSbj4Q+VciX/TavvNFcLhadRRbitlx46lp8djF3hm3uJFx
9S7SpaLXGBvnw4eYTXdkr3nDD48PgC8WdMhk0r+HoboZF12M1QIEEWAQw7THg0XUK1r1FebFOX2q
jFohCWWX3b4N6q+yPRUw2M9exW1z1rBoyfnJo98fZ3y7Qu8geBc1rxxCdOH9ZDBmr5Ol6B7QFkQC
29N+JHJt26TvwADH5ltJ4BVzf6c8y+/3uKAEioCH5m/mu0u1ZqgAW2Y8faZUaP1lN6VeAWg/ozsO
noq66KuFJYER0HmXyrMbZJ1x0p8psiTSqZhaKnyNW26UE0vde2lI8V7kA7t0IGslMT2s7cTl+w0/
s5TpU0zU7iTUXuGtaKnEQayqtCw/cluG8xodAVew07+6JfrHcT8T1hoFIepa0Ez9NfcnzUvmqPxC
Ro/BwrcRf7yU9tRMZfHjYH7ug4sJFOWGXPAD1O4D6ZsaCGoIYzy5vDcdjxEU5TSVr99dPUF6Hq3p
X9JQFca40uJDQlWVsU20bxjCXjH3DronqrbthLZR2VvT3VImQq3+2ErayztJuW7ljHbV7n4FDq45
mugsi+W59KeUeTbBidxnXkGMU+Smg8AHKKe56VKElzCo8cQg9qVU1Y4tHatwUoI2RX8PRKx0SUM9
lYGjCRbdVKuQSt2OeY1UV0flz4coaDtojz72D3QZty4CPdVLbuMhdfrkRinxXUs+eT+YfJX3cGnF
g8ip8ht2gh9JbxeJcnqcrsMx8+w6StoUYFwRy4DNHazPrEz0mzicDnx3fG0qJzUuWizREKdvRjIL
PSXL2Juel5pi15YyZ1iQpiNlxXCLqALnNA+po3QCgl4VzfZKUkLysIpUEqANRfbT7taFw2IMi6sD
3OpcTGzUn0HJvD3W3WpGybAl3XsPWlygIKYq7lpfqrkvmbECfY4EtyapldB8YNXFTfUS44KpLo/h
lFqnNQRqYiwCMILljnn0HbBFJ4a/I5Ynsabw6RkNf2KMr5n24/vetObZEFpdmDaNIiB0gxa/j4d4
eodSccX4Qv4bdlgkMy130cP6DsrTgGpfBGx2EekhU1xMplPiDE/Yp8unCRb6GBj5FdfXimIeuZp+
4Z6cjZHf+jqpqO7XLRkp+Kqi7ckIRU0kcft1fpGmNhtbQnClREeRyH6x5EDCIT2ElolhmwAFRokH
4p7enYpl+OEVOk/Eh6uiR/xiO6L4W5hCNbiywmYB2g1fk/Kc8noTNSKdVPi6T1tkcyW3JDHaar0a
jljQwSS+83aI3zVPqVrQGtPaPANR4hPA6h0DnlQYnwxvr+uG96/T1KXcpaXpZ6CPR/ZTraGSQgpK
jLn0ylvG8Q0ba8ScsFp74imcjd9k4vNY+m4Qj3XWPjSmsawCBL55Y3CZggTj89hW3SPsnGis928W
9PwVqEovOSVWHGrQv3WTKYz1jFzL652mUpeAktUhb5iWuFvg2QVl1PwmxZWyboVmIHbXKPZTCaqp
pKfs3/+6AZ09Jwz/mHaYRXi3l+pTUY7BbEyUTXlloHKCE6n1jbWdCn5ElMMhE4UvxwrAgZ5yB5In
ZFqe7eCANaxaSIARN2/V7BXf8Yh48sR1lyF+EsRa3Aepy6Ne0aAbvrDrgkIP4wUmf2rjiWWbT6/F
l0Y9CVm6ttBfrzkWxN7kLtseQvedY74IPNqgnkB2MqYEA5I66V/L4Kk56viM2lXWVnXhJGgGuNrE
kFl4oL/PimWrRyKAPdoBng0dMp+k132r5Ysm9dYNtph2UJ+6I1SGohF4hLhQMAv+Wnh14ys3O1cj
a+ypZmOIBZHy+QKA4FJz8IC/F/uRe64P38LHCk5LP7rDvatfI1SaptpS/OX4iGBdFTSaKkH/mmo7
0KCSx5dXPgJMazO3ALLPyZoHRssAZJ/tze+zFXBooCIp6c0J/jKnR2njXH3ipNciwXMbnjC3j+b/
GgNBsWnVcl9zVKv52n8jIAWSuwu7AaaQaIhSFW0ZEoSRsk6yI5gai9UXz8gqVgBEFjglTZxDTwO0
vVMY9cehMrWjmhkcarQy6JyKurCMvOocwgA7pphKhSxqIrZpHBM1p3OejDNgc5rJcyiV/H8sMF8S
5vA37fxU24yVMF1kSD7bIPxc2kIBuoQgjjuChPwSgUWWXE1e/zyFxTYsD6XX8oHVAvQhAY2oJWgL
YxJKCYxtBzJcak9IcvzZJz0FpLNVlpH7BZZPyWoo2/dYze6LWmClxbNbEf+sqJhWkdlvgckK/8mR
2H69VSc3Mn0w9Zrvp687/jhvn3FztdROKx2AhjBEeKSVuJLdc87689ETrNqqEmK0bpMU+zmWrxJR
Lsv8PyL5apW4xzLiostFw0ET9ZJpZiYxCsek5qZJjswwdQn5rDFrkDMqH9DSbw9w3yHKMpkPN6tR
qJuPtU02tv0eN9eyQvVQRymOgpIr5C7tNdoEBdtj2xj5kqarj8ucqLr+yZrkezPbNY2B3HcCvZjl
lSMLz0rdgiHicoAQ6EcLxq6+IvwrPwAVnk3Zs6nLOpzL5GIGAW7HvBF5vxzbPiXJERMYzb4Bmfah
yQt5hIqcCveKCX3etLnLzwGH24TcqHIJK7E+WQcoBkIAiZ5XXjP35HuNTxiKI+y/W708exu/w2hn
0Ra/rBr0Q8BSM2/CwduGF02t+VVXHtZ80rnFwgunrX/uILy1Dcss54mCJUKQyRbSeKoKLRx2bLFG
mmveR7yNw1fMIC3Pj7lfcy362hKgnIdHWBNQ6ii3fP3yiZXGktXsk0bZUE5WommKYIdQi7XX4YUk
N+GAjeUCQCPF18uCaH05b46c59onP0t26ZyvWTo7h09Q47Qdmo1rM1/bXQm8XqYWhQtSZzQD9zzo
yyEAwG8q6LaLORZtZGYMuRhSqYMfdJsy5p7BCoXPi+rQhkmhbTle+DOFxhZc5teOZdO7BinG/Bxs
BYsFToUk1JcKC/VIe0X+vNZxBoS2LuYgnpBDtYSNijqVmVdGZMIiTDLF4iajrOydyGOeHDuzWcSz
73cn4TkxvkD2umcyecwaytQGyju6iZ3pDu4AerlQN4APxD4xeqd1SOsuEp7eFLCRbekCkfmVGsjC
Wf+aQcIMbszfvlOv+w9ahIl/Dz9W+zvVJ/UNznJZuaasBxwbASZMxoIYA7jLvqPcU5k1/AA5wK8N
XQRJEtCtGhm/HAZ3AcUSQNeZ3bw9WMlncASWOHe4BgVXUH6EIozdj066sT498WmT89V3S8j2pO1Z
APS0xyrxHAghiJNDwuDo7ms0zJ5suP7BmkAugfR+xgatabGRoA0G2ncQlYAIe4EyZms3J6ZE0z9r
QRhVhNvSEhzl4YUW3WFxorSPKtEL2CQC+ijOoJZ9pwxD3DQceb9lPthayyIJIcaEZcVaAv9ulnJm
b/Q/gxHBSYZFAM/esPKW8Xir9bZgEjQElM/2JqjVkZJRPqAvzdy/V4cLvtSuepc10r7ggjJmpyOw
sScrYltdhfmyfiB4PpeczJJEqtuKw6jM0a1mDCzgATqQUaSGKLtxa0mOVMxkZK4np6ep6N8OEHgd
ardlSEP+mZIxIUbwbwAdHO/+lSQHf86oZxShGLyd9VfUK7gm6DbqSZ+CEV7NJVcEv67bi3p3/12c
7qsicHyqtULemGdZtOtheRKtOnSH4CGM0/klcK7bd3KO8TFYDD+2KHkVfEZ9aeKC+QVF/Nbv1234
GrPYH50tRwUcX/8NK0z9AXX0XmQGOpXxgRGLWuiC1zl8v0aWVlHVJ2rmtSq+5wWnXueU1OSNc+fI
GFo0GHVUoGkdH66GT0lWg6z6zZ8YXPeUppkVHqXNOY1WN7LdDTmdG4TZdYd3bE6HPOZ/4O3cIOoT
A1m00tJVxiyB6JFuowyg9Q02Ao0zp1/8Czif6QSF1sTou3IQQPGZuDeDtRIdC9ZV3Nf06+gCtOdp
CFpq3V0L6lItMTSD4JI2q5UW/WO6wt9AP9tdYKfZ4+Gn90GKHOkjRJFHVx6JcmdrQFZz1t2nJrqq
fB/zdh1uSM1fFxe4pK1/YPjYPL4I6ekWEXNosTARN444UFsYHmCUxwKyIT+508HpUjC/hOONH8X0
sHydI9A4rjf8pVP33ZtYULMoQzuuqeePY5d0gH4drAgtEpa90653L+rn6SyCXve7UHHZclIANAvb
RLM00xXiDhoKKXmY6EQUR1mkYGF+7MPm/uS8Y0r6y4vfKX3dyo/QFK1pi9j1jMd+zrPBO5UIyfoM
5X5LgA4Dc/iynssWvyQjd52amCdM7Fnal5D8SZeFhayF7c/FkDqrAguQ7UFPhKz5A1HFisXErHm/
EuBAnXeUIAyYi9/odmab1etTR5WiPEnI9OHH12A3H/VlzFdLI7/5J2U3kriAOTDbvS5Zd9zBP6/y
wCZxCT0cyJqq7OJtVx4fdM8iZlWOmltHI8dRyg4lG+ljHhaET7843MgLQwfXwG+6t8pURna1ZZNf
ZySBtgLzkhouOWVeTAZpgkz4NLyGSdeDYQcVS5sYMddzO2xmvBqyBVQD7uXJYIdqitu6XoU30vGj
pjVCL9rFbJX0rpy2V7m9ADtRMIpkpviE1qZhxMi+fWB4uNEEJp14ibQj9MLLM/8XsV/Og4eFDdEc
cnR+lxOIabFwdTT90LN9pTrFH/C+dV9TsftCW3UtgJVCxezpnVBKNlkHWRlGzP1P2v22HrWtJib2
//seSMGi0tqSMLB6sX+9FDChHf9X4JOxzppALoTOQrEnHUrdhHYzdZAP+xLsx+4gQvB/GBtZWE8n
zja5XQjXjVTTpWF60ECYjzwr6GdgrKJyW2FjY6B3MEVihK+PVC1Ux6b0jb6tLsLSj7rROSKRmecH
rHwV5e2CMazuHaVUb9emACgC2x5hU+ElQT98+P6dkBQOYZmnVaQUqEu/wzrMbPBhEJ9Bg8V3+8EX
4UOYFq7UA4+gFN5DLDnuFlDyP/3jUmWJtpSS7dAnePe1mXPBuL2appPGOOZ4hv+vnfHSk14gtMA3
AwlcI21VYyzT87aKqegbTWpmhuWN6lnDoKpiV1qSf+B0Hn/5hifzc9wjZ+LWczjtHvrSZWVXKMmu
6/Tc8BzvnlVQLRUafF7fIi0dVOl7khDTpw6LmR5xI6iVnBYJ0Jd4Z8URNngsG09akB+sWCnFepQQ
SBidxp9CumSaquP2cxjU30IMerHy1GvocPw7lomEHOD1RZbsdA4mdN/Kk4GgtYrByKG2PxMLn99T
l2nH3bMzBz3rC3vM5xhV+H/LDS6mdMO2AgBPK3JBKPjdRlVPmGhWRllZ997XIdMPI+7CjrFDwb1S
GYHuV9hNDiZhzJA/cdTDxyW4L04RE7GlQ+zsWM26eJWoc+yrYSwRjaFi2wlGDc/Npzn8yoAfxE35
bh8ekSzKJ4RIlVeKx0tJMuANbB1wgGXCPvVqwo14npTDSfSzL7RWXI8AQkuSk8vkP+Obpi4EDYhm
oR5PDP8z+3X28jAhh3ouwYCqdMl/f8K+r6qVzTTFOPW4UYJ7Nhqyr35EcU38FxRVixBzYM9wCL5U
CF4kmB+WS0YI+9ysuBkYnYPkceCJ8LvJQf1SYG4b137TUR0VMoUxYiC5204ArqJFf0ODtqzQ9Y4o
JMvRJVwnS4pebfBwRZj1cNYbDMb3b9oelmrqFM0WTHyLnKg8oy8uAKtpOEU/476n1nVV9GgfI2GU
jCKtTqx5/5LWVaVfp8S3c+JxZUBIzNuWwuyRyr7yhdEqdW9rIlYAZcuAysXHilf8ruHVZv5v6BgN
Uvf+Ftdk19x4vWdm4A4PcF/0QmdV/9QRa7ENC83d6itL1W4z0WC1AOCK4C6/HC8PbrdPK71eDtrP
6khmTglMPjTjv95WKpFjnlnISJr8ddfyqyUk+pqITi/jG4+TxSmY1YCdulV3U9PIzD3W7JQ7tGDw
+qZQKalnT33mY2U2Ensp4Ib40AVxrkIRWweDzDYvw8zVUXorOCXLxqJ2yrXIRMHUid/Xq9PcsI3x
a2B8O97a/VWGx5Ngkl8kuoflp/ZEjG2VIKBu/D6PzrRDQI4bl98epmpH08Jan+5g1p9W4CWyODP9
FSTIMr/O5frQ6p2rabLwRDkthzWKa5Ipb0V64AraokuyWHlUPJZIv5NaygVhC2VUseHzc80j+fxF
j6oBSxPn6rqo2Y3L5iDMW1nbQSEEd0kyR+8uoVRQDfd5sREsNrwruZ7RG3MaUxOMjedxBno5tOnp
Y+7oNpDpkFOj5+8HT/hS1MP9+jOdU2wRNhS1T5Wk7lfY74OydklKbCymb+OGTIEbUJRdUhZ+OMb5
574i65q99dnTtAHyn2u0nBbW054ellvzzS5Ot8ne3QOUpr1rIaitI+EmdHppKAmu7eyXVmeHYOLK
Kt1Y/x4oT4vwcCmRAOI9okiPI4RRNDY5vWmE8s+eYn4FjNHuPFCfO4OqSTu4pIj/5fxurn39LWf+
ftEsCvnWuGBfKTOCvF736I2SEGLROfrX/sC4bqO3ocCdqT+jeVvLGSxDeB8WNYW792x4ceE9nvG5
XLzSN7OGFyXZLZtbkP/ucvV3ZwK9iaz5PJTcg+C3q2BtFIK4lY2Y0ZGb7BC4Qq3CkCnr+dQzoFy2
BIJpadUslMwuRkLHSJgcBuzrRmkxfHpY2ak8lrwbsx3VRadiqrjm5WHv+pF1bl+VegxNDMSGCbDN
ghE3wbM9L65Tcd3mCZuvzON+ObUpBaXIaQwJ0uAY93J2DveyZ1MgAO3EVknrres23x2Sk9UinJcG
f/B+Q05me+EyIhw5V9N9cjj+VQFf4VgxgvPLLe1Akq4MNbdSOu7ZPaYc+59itl7/W++GR3KfREVU
6ebw4n2fahqPZdtWxipvdo6IAmnp77m5cY8f5GadWsOjg2VtRXiv7ILICc8yIerwJkppncsbtj5n
tEAK0NEYO17S3rRv+APDfYbAilkOf5dtWmVxeqJOv8VAW1QCXu9Iqj5vrm92mNKVXP6S4Q/7sjmb
Zj6SJNetxaDR9u8mi8qeGFh396BKxbHWONksGM6pUcdmZMmX0tvskyOPOYFwlfMJkTOu+cFr/W/q
ZWePWNTMwdWsF7OxU3KRZmluCiJVuwpELTbP/QyykKaCswEflXfJ3dMgh4ISf2j2cSoq3XNJpDjK
TaOqfZ4EDN4GG2zSvz93fwkmUNlTGI10HYZpGcZCLeQTP+own5Tk2Twm59n6mlUK7WA91hYcOypi
Gz2hmnVH+lxHrvDVOXC+ba2HhcxZQ1PM/xCFxoowRrze0gvYYprdej1OM67DxHmpyfGDsgiJP31c
pseSnHwKVCSoBmE8my55WijTcbEPkcXyh9nogcQQMQuk/MdPbjrpZyC/PeZtmmn6zoZbQ9/6Fdmq
mZ3N5TgcdHYLt4rr263QUllb8XGi2cXXNW/cRNYZAO74Xp2bbkrcZMqIEMnjNsaPPlpCOU0r2FsT
yCAE+OnP98OnZgTYsZHmPfB/qqxdw6faAuunZBL4ZaYq62OLPodX/yvYjGsPfy6JBjt+XWFhB4Ne
/S+fzU80hMhTgowPJh81rv5ENgis2LxEicWG/fbP2Hgn254moOXMZrMpe2/Ot+Fmkf9YGOkBhObX
1crJuH8H7km3u+V0fwnbHtTz6W3DhmXCQFPAvA/tu/GxAZYXwwQtomOKZIC1nNRkg6nH1Ui5k2bg
pvuCnKdwrvf8orezBU60cZC/2xXMjkENsZBCqfX84aMKBtWC/tBloCrS8NjUxSWdRTBcAkGTaHEk
d/8fE6FW7btd9BSPkDuh8QQuBePIlpdNIRozryKwdbFt1AJvc+0fkyZizUSuNp7AYiui+MPTC2eV
PFfaOH2hxS9+/LlAISjOv6p2HtfkmnnbRM3fIi/ri2kp0uSCEhuhg4XdN2VWi56gC5/ZNPfD1o47
DVJBo9YH6pDcIYBzzp07u+rB51ccxGVHQ89RRun2p3Of+xSu5PXe/mlME2SEBkrAxpCVNaeSKiv4
j2hAw5iELdZGfpYwmQxxzNnvJ9U+Z9HFnDTsNSIFtBB8hj2+qwV54ZAIsvtrcHleokJYE44RCe9S
/5dwkbH7eKfdUl9BDEWDs6FQk13Sld8LhqeQJNMvgPuHb00vT6XGBJNhHuFcDk6ltoJrnkT3AeJU
uYEjOTFGvAvo+ktE+sEzUZFSm7l9jFzSuWBexhWg19y6s8JGPCWZebVQwbc0YzGaiy34MIQbJDtT
uSAxhQwRmo4tJA9pSCFxkD5DfmGAKQlnFv7ma3IAd74BKRYrBYg48DPCJwIzqytIJYjez7o72FJA
3uR8yMkBA2OzOgzHg98E3niqHByN/FHfGDUjmBkYzN6aOVEyEMokR+efoziHwDuI98npMlLRXOc9
fqJNyijtDH4by41RET8mQI8XNywlBTuDu2b+ocFvCLBGn32t5vKLbP+AKA/TYgIABuUr3fs7tr+l
EZwHdnKC5z0WW350mE4B2Ov5iPRuWex2R2Lz18WwsaqpUJAG8nzyL/IUDfKykEoRQuAFr0IojJUH
E1uIHQD1Xuce8/qiuFoHAQCu0DKAVY6OCyOPepzXEiQnh9oECC37O/8jIhPGf/o7uq+ZFAoXGzVy
TieGMPsYwISzO5x7pCEv49A67WldZr6u0UqAJrYqMYNm7WDRhIR6XojpB/9T8huDigtSk+JYYtF9
QyJkE9SYtzfwfnvS75ybGs+FOa7F8pw76iPsBrkB6fJ937CG02paxqrj5g4i+5FakzwSfFzwb9U6
xRKDhSOVSjhHtVxZReUxXrZIrsFvNCNZnt07uHJiESgPmNnhW/V6IFhiPxAOYSgoQJAcNsB0VjbR
4/6z89YDglv2PEHZR3T3maYuptGbi85G2uhehCFfP45c71VxsC/oK9tVQUbXxyVla5DDpTsBuwG6
Nb+uzQ1sIP3kY+ixOjGdn95B0u1tarv+XmoY7DylDrtZw7SxlUVkyRpLuJYFxnKuBHEvHq0ezkaz
9BwWDxxa/jul99CIqiEhhRCDKdkGMvJ5u9is+eouwGQ3G0GpmKguqllPxhX0FNCKIY94/lyHY0Yz
jlHLZpFVYHh4KegHZZEdQqBNF7fVTlHG/j63VZS5N4ftYx893BgoZ6BT0sHWbU71G4nXHEgw8sVm
m89Il+lIRPF7WDq9SaFZXXeFjaccChsYVjA1lIT6r9ajAvv3yUBXaSyr/iwQKXP0+JfVewM7FUDp
Kg1K9LLL0o+DqFoEfS0hGSBLbhakyJbBaKxnrXt2kzaoJxVIpiiMX93vtN9YlDej8bNjhXisqUOi
4CRttnExhR51DZs+bJrX3fd74n6gaqHAy1MfL5nNYzY2PeDaIs9cGpcJQXVZ2OLjCqlgZ/JUuxxV
n/pjTvrtp3tnBtWUj+Hzcwdua6jV4hr6uMu8na/aVcY+gCv31o/CuD6nsm2FVVoBkuuliPqitblQ
eP470Z3+Z5gpBdPEpoIRo2r4Lfpito/KbdS6GoHVXcZj95+NeCsjoAjoPWYVw5AfgsqEUCZY0dOR
nukBTHehgvDDgg2TsscXls2o1fAKhueBQloXMwgl8cerCgVk3mcByHlItiJ/vimrma0HHp2+mdOm
LkWeziN1a0n+bDmwMkiAciXMNo0JJY/VDjF/mzy0P9f0iTyPiGGi8S1c82i+rI1L8b3Es7Y5fekl
ftx2JhLx70Af0Ka8ScCuzPZu6fR6Jq1TAHpAKNa4rZTQGCCcnF1hWdha64IqHnB5fy15GMp7RjBj
grbQnSpK1ThBxiUMWOnALlm4g62sPvr7aASt5D+a+z5rnivcNTT27mezJADliIxvl7Nx6LxCYofJ
iL8MTP28V4LKGBZIqSdsx1PsOzDjsncps+mO2J4NJpNNtqX0pyW0qu+h8nn7KlbSWRKh42OpW1fm
ezIMBjcATxaMsjnKHmqxz6tkteiVcgDsCGYFd1MDqtpMsrP1+GrJJnxLwm+VkYDwGffiNUWRTP4/
sOamZhr0C097hoiTUj0IHNe+9gk7YmDyZhQ7dNfkZEaiQGQiYmOzieNpAkzzNBTer9eKv9ADVq/n
qptAnN15ucr9v+2GaFoDKiyZoyOpME/Q7BKU9UAvsypDs6OmwO1aA4l88Sjlw7sK0LWORysUV6Ui
D2iGQPgYNkxREoSxuafNTsa5jhztjt3GeuwkptLmHGA1yH74TXHs2KBDU/Kyc2xjtzOhCgEltDW+
Qmbu84JCD3GCH8aPNnkf/Qy+SBWWMOPcjKD+N6XqR1aB8RiXxGWxzJdLK64WYuVNODlPouijTxCI
efz2OA/cmkxarRqiTe6l/jATsS3MdeYNEi1UnEfnhaIf2/SL46ENQ62CdrT6qlK1luAuqtwi8iwv
KfuYK270o3hiYh977/GFaRZBUh/JVj1knrj7Nb/8xEyEHPC0Pe8lc/EQd7fbWiY1A4wIZOW2sVak
CE0370eqNKpuXQgcTBR6Lu717CbP7iugEif5R7M3F0qZqhniufiz4QeOZnJ8Vz/tMOpMDydV41/E
M9oDL40daRTk3ds6EYrW4amHD7ZNZjXuuXb4KRJ3dcjxaY0dX61+qMYX6gAtDKJ7wzLTXEdHCqIG
1l6Cy+0aNYYUexYKNN8ieGffucoGg+gOFWd9bHvDu1YUm797P1t+L2SoEGQTswL9zj23Z0inU8M/
nU2hlW2OhgQ3N7rQ+u6zEsDFvrTlnQH5TGtJlE0Ukv9TZiIgPqDjiWIwt7iEv6LiwpSIPE4+3m3P
oAUMClJobeCRIzC8ai30SgTuYXtiJkUi39cTcCuoF5Rco9m79XAGU6b6Ye3lE1k6cCJv+GgmdiB8
piIjeSNeMNyCtMBiep058oZOgsIu9EJjhBEOXZAh+NM7mtiveWL61ux+2TkxpDnd9uvVV/WXnxZS
CYLaaXjeG6T+tjKAXb6aPp1rLzhYKSxeJM/98PKmXQaf6z70ZJeH+8moalRflfCNy+Cg2pDsmY+1
a0iWu84M0NE3OWjisVmcignYJri+u97TUDSs6jFjO/fGeBqHB8URBxbg9OW0NQfp7cS19gUhqrHQ
3UpXVLEwwKUrDCXm4vEky80Lr2kEPr0tWh8KH4UABcFd1Rg240aVM7q8ezBeIpJWUWt+j2RDu5nx
O3Sl8zn0I0e0kibSHDStSbMy8TBg0hdUmdutmb2QQR+5X8COy9x4uoQXS23IxgizvFmdosPEVCh6
CNCT5/GzWkVxBrpEpFuYFqbnlvoOIaeKpW+FoLLjJulZV2RWgaauubt3d1fq2M8T/vrFheSLy9nB
k3rbkXi9NRDfru5JFFLoHjHzV1Ss1RQ1OiSZ1vjPeZiak2D9mFCui8iARkWcXwqo7Ln9mTtGyjdV
TbYkWlegiRJ+jkC19MgUX38s99uY4nlxjTWQ3iWWtqbiiMo+1QZ8KDuM+mjNNzGV9+yQ8VzRBfbQ
C5C9TsjJfB1MEAhTDfO3uGsNamvEMWFa+VscjLoByAS9SUuaSufJwIveeHdWLCB0Ge45h6iY9FCo
N6Jg/jr5G/Q2aMH4DoueT1EQEMcNoo3Cu+UhOF7rhZ76xGBvJwujifm4WclDoUIvAwtoeqNicoKD
xseNx+F6grWYmaC70cpGPQpVDqJR/FGe4n6Hipxf3wMbwe+CMntOf9L2uoDOdI2gcNUsozJvLLMx
bqXjjHbjqpElnxUeII7CTFzZQ59XDkc5FpUmkSRXNSuJpwyN+v7FIhqlxMCasyRbZQPgeVnnPCGf
K5SOcgnvilJUv8zQRC8cVh7aKOf0N/y3g5KLzBbo086izLjHzkRg4v77pXO41bHEEjYtiPeh+mlZ
IyXPOBMWIJUBJb8nCOMZkUDoEcL8E4j2AXHAVjljc2OzXs5lW2ROsb6a5n2VeJLRn2eofauvNBPt
VsEAuW9jrWeU7kcxarnjVvxL6VaJFQq9yUTzxrWDZXWI/B3poDEM2T4J96L5296GY7ueOe/8p+PP
q8I1NDAwOf68dk6JRZIhgmPp4tg56n1c3MkCQPqwPhU2qeMopwN+izqHbL9nGC+utzwKY0SQTfE6
ahoMhLJUsQFBTGxHQsce49/SW3CwUZVUl9TYBAGj7tddDrfCZ1yAzv42DoN8Iy2kPEsezokPfmYn
+UHiAYE72CfefZ3/2Bkc6nKQg/eiVVbw5hsGqVVumrr+0FLee18A7G1gkUl1+NuoOvhVFeKRXuTS
8foZUE/xNb6W+CMqdsdXh4v0dSsBv9pl05V0KV8TnGaNN+BA4J4Mp8cd/ekGSlr64jdAcKCcbmyy
zXEXPntzFBudRsUDsj3CUcUHB63I7xvxjwZkcuMBxcfFi/STbr8wUnXwjSsWlQM7sQiGR38XSYxa
FWImJT6vWIzEM5rx3LYUOx/DWj4gluI4Pf/JDg8ZLnLbYGJI0TefGv5YzRtSddEN0jGVIMvRaIkD
yIFn+PMe1HYLVDtrlG3fZYpbE6/zZ5rSiavVf09Z09g7mLoXeXURZLbxeO5GZR8EGC9l2NGJ/HTf
et1QNVxZJ6GVFhDdaKihTvUFmcIDNIKi0L9Zg6RYN91Dq+nLMrKZ71NGjJ9srekfLHVmnn6b9Egc
/d7i6gIf5hj+yMaqaicwzamCxIRIaXTk3v+qBU+lX5BDpV+iaaB73+d1WI09vfh1/xb1QYcE7fWX
+1nofgzU3wO2rZoaV9fDgAcvyRYl9AmQ57OSPiUm/mCgH35JaKav0rkRClyWdlSN0HUCeNc/O2GW
cOv2jP1soNvD2wxhJiG0l/bGxTXfV8muCbB0cpzIfJU91JpliWF736gSc5w/Hvq3IxU+bOcWJvWs
gVyQSV7uGm9mfJcxZFeTVZB9ZtLIqpow2s4ayX35pQHGhnIngN6+LObYTM0QoSHNjkrnGC1ZCGVA
gW8tIE+BKmlOBPBdDV4lfuzpUPHGahiyW4dz2v32DrQfpBkLAbJocwQy8l6J2c4VS+XNymiA7qp+
2ZBGS/cJu+7upwdilgrgXsaKCuxTJ5ZAJAa3Psm1RCyiDPiBsJNdiFLtjJwtOnSVC144fTMpj4cE
ttJ+zELGRKWLOAMVJvtpIxMrZRF86876u4IYXGiTbBcjGR0jitOEvot2bn/m5HUug9ckwtXTExR+
E5+O++/NP/n3GjhXsYI4jy4X7LeU8HVtgSDpdITHra51AdFb9/6L6qeXBmrB3IQqnI6oZFyWhj4p
Q2TGxL3+Lud2GNydtegn3N+bd5EKmT4RwgJzAmWXEW+TELAhpMj9+d5kEj9SjApCZRymjTSbAZ/a
IOZBYt2r5GGog2Uk+WsB60IJ8kCJVHDTZ6WwG9/f0qSVcRu6X5bg7xiVdk+p+EKvM6ndzzAxRXki
2bNzgMKNB9Ee+aXyQY8foYkfEDMlBCJuyZjvJi5qnT1uR03ddGXjAUSm5VBJ6xrpe1rG93TOIDHb
kr/K21RZ9aXmZvr6yI4VHerE2GgQ3m+FDLtZaSKaG6vkRuuIIdjyS8YwzhLrgq5KUZoeA4s28IVm
lGcMGEB1TWD88NupJGRZKPsO+2q9LiCsGDkfU9Bj9ZeZKyoO6sZ1XnQUFSrsggvZEjf95p1oNbvG
fIUL40ApCNoPXbDJIkpSI1bVebGjDV2qGc6T0J1X6lETSnwcA0uaR1Vq1kgP3j5mU9DRFEfdFtqR
Lk7X6pSYV7TPso54+IdqHHKOmvYhwyK4KOzo7xfQuyvJ/mfUkX6QwBVNCmTBBsjNHWsr2z+Iu09D
sMDyENYsmb44qD3DSLzAlCJZM5GSfbL+N67ato6skJKVp4dbskxJT2cofGotXtYF0ogUhIHUdW/F
YNeNJoJYBmrDNMCoo7Z78zMaiPyGy3a19gLe0i/cgpq+8Ngladvjr0CjeFxJ10k4oBQj/F9vIcV6
FPa484+VU4M2o2RCHue5lB193DiXWay2dko95R1a6HhOtaFKA3AkA5N2MV+ShvChDG+8ygLzt7U+
GP6nBfggKpIdqQSWqaxfxFI6/Gy4bggUEwr91zzJvH4Ka4oXcXPa9NGvHdbIqYZODNu5rC19Gl95
iiwaOZup2pHO7+Una3SZfgO8VW1sr4PSNEyj92G35Q2tLf32ejzqznEr0UOspi3zJIUY7aylDFYb
9RVBQIyU9gwuMxV36U+UtfRpmpJR/FeKfBOQGeVMKfpIR/DTC/2WhyxCcgW1aj+CL35eWGHrMZud
lNYL2ZPzd4VQIxltdSiTaxKQZ/IkFR3wsj0cQjR3eG1LDKwNl2M9vkuwURkzJHULL0FY0BrsaMGf
MiWGvJK+N1fdAy9AMI9WEwP5/oVKOGUPKgSNyavt/kyeGQ0/KHhLaXLlGz0AqnmYBhZwWR3YyJwZ
bBezWqXBzHI1F1kfMPyQLZwhBMRC8uLiHTjZ/ozDswtXCaW3Ww+PDaQc5DAAgrxpWRre72xqi7Qp
M0MfuF6BoQGM5U2/LWnhZRLsvFz2fopwmb8/hHQnfQN/Qdrkplyvv6D3AhkCQHMnMGQnLCCl84yO
/WMfGmVxvKiNiPTUAtQaAj58xe/ueruuqN4H0XzJ/NksC2oB/exE1itI4MGpNnPqufYPNr0phpWW
nnS/IkPEiI8hzaijHIF8yIlAv+EMsEHJJPXpT33Just/9rrogVJYfRgGFe8jhu1452WAUINLS7D8
InzcP8LhZozJLxkX/qGLpyINMTCD0wThNjneYVwHM8XaGRDSAqCTCx95CkTnWl7A2uy6RdyI3zlY
d8B+3uG9aBPep/fmoSYOvF1mfEPMjCRuo7qKTf3ve0DwZ5vbsf8Ong8y7AlqmtzSXXqP9NfQt8l4
PD6mSv+YEu4l6qQnzDpUyuhMrboDtCwpRNFW8j+d2B863A0Lo1A0//beQLH0wfGqroDvKSHGRxhk
RHA35cMcWprhaFSeyPMil78V/Kc9oONmzeysszDJpm90iQAwz+I94hZI6Qo8f+EmvS9Eldz9j53K
4/4PXkbFrP1ZLFhi6+FgBZFN3ep1W8Tn7IatJk99nPyhdSMGRZesX2CFoPZATgzy91AzK/tXzm6M
MReLreCaoZPYFjOqt6RX1JYKcHC/a0utJTT73ps+GhYvT570WdRSoGGx/W0TRmjtGRlIeKNjxv3l
DiGgfBpV9kzTPR0ETzen7yFPJitpMoYsPSbM3JWv4CFvYZTJJKxNVN+EWqhuhNNd4K2ly2RJjPwg
vhhnOYFEbrPWs2WO3B/kGz/liosowlwt4jVubb1QyFGeByYwFrI24yjgyfS1iMAVBMI/Hk0yFuvW
z/ByMNMskcveIuFJ+bH7YKFSG1Jv9ZICvJBFRXZU8/IVyCLDu6LAG34eEgT5wwFwPSIkw88dY+Iy
I5TueISTK9FcGdDdyLryA3P6lCX58RUdYK+WQKSbTQdp3ndj7s8YIf3ih64spNQxRVPPmc4vULZd
UMYnRafQ7Bv20CDmkc7jA7RhdJvN/ZApxICdmqMf3moKXEzTB5ABAQCDjq8OsQ3rK+9V0n+ixEQ4
zhReRUjH6++wtS6FyNsSN2tzMlLk4LH0G9f/KQYapZ5Ndmm5t2nOQjelX9ELQ3QCxWV67iNPlFYO
gYdvtrzsI7ne6sxcY28kOPWaRJBsIQx8D5fzFUbEXn5eNmZekLFnvqG/JFUqE2VNQ+x9l0Q08uWZ
SsPrqoBb4lZv/v/H1GR9b8cRzjL/WGWvFVcQOKeEpsQl755JNU0CC95/ooX7E8QtMUzvQB2j5EUu
sqOwCVDUpeknT7LkeG6u9UXnzlzAISQwu+4oUvdCqqmyYYgkjYqQ1Xfy9pzJ9P1z7VmZsdIXqMEH
EmIJs/E9Nx+oauef/bZJoJyRFR3UemTIio/3UHSJev5BTh6Ftuqph0qJu0qp1vgQHC36+i5c5Pc6
84j2Jche5PmiSoB9Ip/9Wv2+M/PAgS6J5Z1nI1Q0A5rOmBJY1+fplDBNF87ghdVhfM43gRcte7BO
vRJpHO3a3sCbDDVWYqjhOCXVeuRvUXpQkDOY9QxotLYHeqnqosjE9qyvTuzVaWJTfqPmydl5J5ZW
ug7i/1rmQCZLqhW7twbejVWCczBqbssemvynxE8SUwmYuS9hNVtf82hmBewI8SKsmMsHsRRzlmIJ
JfoQLk2WnXUiARpU1zAJm4bubtylNk4yxGYqPTkOTjWe2H8uFNM4WCCH4QUlPP/qngWR+nBG2D4p
bNIy3Zly7Nd5MPL/vrXfOGj+1fpnw0zQ1p5jUMhh52nvmbSkxx77D2gJE4C9/ouBK0fbytjIBUhm
O1qkYWtIu5V457YyJF1uAoma+ubOzZPlMk4ZxgAqxRTj5vDRdvqb0yMJdU4DobrZhPYJNx3bsTpz
+KprB+e2PNz3lYdsyhiAvG+Bq1ReHYzdPvwPAS+QwDOM1rB1SZQLe9Mb4qLWEgS0HrZrkpFRrmXl
5eDoqGoQKOm9FITfSNfdy5p8sxFOKY7cHet5z0eJgpSHiFIT04l6EStfYb3sAM5dKrQtu/Gk1Lkv
r2iCDWyhAfZM58M2XlOtv57AcNe26XCAG4LaTsTD69VCXkOv64q335OwI6CWtSH0wfLNaxxPckaY
NlvNxOcurj9ov9LhXazCcU7mvzY5EJ9Z1WuAy2W8BvO+Ce9kwk+icfzYVX8fzj1s89nBx9VZfnYC
N32E9I1f4Pu8xXyhHEVx/+U0Zah7mKOl+yrBzIEPW2U5LKytVPWJGvzfOMyrhsfN1+RBn2A9a1Jb
r6wJHM5reLXahWU4bQ8Vjh0I4KsjxVTw/G+Q+C9xTGiTmipcl9LzUJTEZjZm8UbNbObFAHy+wL3x
Q58yEvF9sChLANWlqcxRSSBfK/Wfmuidm7HBZE+Np+l1KZGXzWEzusF4Zl1XoS+xLuoTMjeeZhDi
62Xmm3GiLMiFtvck+1d9uQLHOPg064EE5XIPLyrsNigv2oiPX9FxzJIWH8XFX1NPQLn4eU6Oxz8c
KlWe/UPWgQ9L7H6beUNudAy02TM4VJ6Ad4PH60LSx8gxoMA0MKoVRvvJ/s+rsuOvVOfdHWk6X/Oj
tBH+8CcQtz/v5cvYyQt4anr463dxWRBBcflY+A3wLbESEjp+Zr20N23AbNhFVLrwubBWePrw2bgD
wgnRR0xb/EvM3lP8ZUoyWCrVJCL+gv2SBGJk8s5HHxb7zzz2VMKSbjk9RjqQK/wC+j3gkoLQkK0f
AttWnhdOzQ9o1t0j4KxvZH2ftkdsIZB2IromVEIbExqAYAaNtFS25SoD6kx7Ws8z4wYLaKZeoYPh
1RmnWTlBpIgERjEWDBYcNb36ZyTmg4vlJvYoxiqRnVdSGDIZXw57DVlVEOXWCWvGnc3IyH+rxZkF
SkL30EzI0TmHdqvKGfu8ggLgUQCdsafpdGxwgtuONv1Fyayr7nrnP7szitdA/NOfhbNts2LbFPP3
HoRAmP7GEFOm/bO3J4AjLPsBo1Ho8VhGEerJ/0R6zfAMX+vFJySxD7vzSO51dkKW5MHBG/VUukcF
IrpaGqsRyOov1mCZhHspnVK1NuLKGm4okbfKTy8YcM0gGxGUHa4u2ORugWH5OJhl1J/TDcoDD/0P
rBI2BlW/WFopNEhsY3Dg+shIGZDdg7udHlW/zJTURhgHSaOk48AQ4C0SrBEMDae2sdjt1FLEZ2Pj
6CR7QZHoHkLenVNiTeJFl99XHY5BUVQglZSojdmB/nla4ngrZ+21ZzGBpi3pCf3rsu6ehSRpZgo2
QPbKpF/41a6ag8xFK0pHSAc95n7ZS+BbEBTUHaRR7Z/vdrGpSAxooeiUw4r0Ny0S/PR1qplRKrJ3
3NqufMSu2TfZPfpJ1S8d9cKCwTgAQeuPBtKOhRBzHYgIKbiFAqpFo04j3xLIOPXbNC4sJ6n97pvP
SQNE7+hFFSz9p3y08q0qVDd6L0Ox++zSnQYzLrRwC/lZXizESkuiKBOmvH/Qlvjo2aVGrTHQRax7
k2Wu7684Nb5hq6ySvdDponSFGtdGAc0WmyP3DYyio3bcD8qkyea/VnYCVqgsMt/9IiSTskahVBYK
ISvN62H53SRGH3fCqgMAx+kxp9s+HHZG0P8PPyOCgNUgdL7kjVdrRr9UXnO4+Ri0qbYqpYm1tveN
xzKzUZOHCtX+zpUN3j3FDy7qqHomCDt1f0kHbphHksxAkr8yMxnT0nqsUgWmflwFZx7l8FKVHnll
Yin/dQOVsKmJAJvowqALKeFk2QH5fGnQa2QBuXdE3ouLwYLKAAlqUx19fnUdsWtF76E1n9Yey8GI
pW9GsTGK7ADf8l/6JitOgcxu5F0qv7ET78z3uDvFAoe2wKRmx5RAPNxsWXsCg2w+CB2pNjwFyf+l
VHa9lHkdJ67mieHDvevoxKWBIwnfIaLVS0E60AO4rmNiXj6SSHV1c1YHV0M5h040jU6sfYM9AcPc
2beBxUz2K9Cirv+9/9qGDHpgIr/fu3lL6RvvIS9Sr5UFICylqHsjUOo8fTL4CeEKBRNGMIl/wCVz
jdUWX2arATphlL7f5Ci84FXyvVSo1ZfGlV9adhS00xFLoa/48CgYEpZo/rVd4nqYUycvxb1x7AYc
ZTDfrx9ygSPzzrU/egTnVECxNsWa4ApFYLeN/LctobToN3yqcMFIOdGRhob0/DdNwoj69wkwSrt9
vgpPTSQDZ9CJnBO3CUcv2FtI7phHzE4nS3ng4qfjgWoVvaTZElzVlNu3D/zkMsJe619l+2zQpxcP
Lezy1nEY1+aEJCCy90P9dL25bLcwXef5TcgCsgvJufZL+m4f/RX2zZwoNT3eiwxI/C+vtlMu5Dfx
KzB/jA/5Vwm7qsMMaz0ur/xYTWGKdszTdkwrTR0YyFGrSFWU+Q1c0ZTxLGr0ZtKhqXM5VDNSQBIg
CmxUoevnMNgMuMg9EvE50wI/Aa2yv+z/hpei4StJVG+8TgBHmp+VF50h+CSRZXM4wO6pgG7nNLTb
YpTaqWK6clg1cQUSRRT4prEnKzlWQrVNh0yN2MuI2fOF1T2GZZIzTjhLswRQnv0ZdwcCZDPAJlsC
mW2Z1tlj0b2hMUxPmxx6HLOOwv1+t0uV8MfbWB3wfDaK/EnHngI4gzUQpCzESuKe0dDDjDdSXL9A
SfabRuZN/bmCThpZMqW+7IwstQQjSPRim45rDpUMmcJ+MUJh8B2cgOc53ulKsSLmmuccI5pHuLkU
W1QIm4knLGDlnb9woXAs9mKRosbFrxlbChMewVJ+MYO9Y8Ohx+SSJfygqsj5LzoM05LwiIN8TOfz
v8ksvftefXFoaf3gbbT89D7AFjCNZ8pnIBnFsjsaXBxhWE8tRCOGWbvsI+kgWI986URzrZJ34boS
g2jxwNG4D4aygoupRGNF7qIphSBtFTTHIu5L4w73OoYs8JeuPXXvMLDVaUAc4QkL5DqMNFV31CYr
LM1go0wDEXro5FmaMKGlhA3Vhw9aV6JDaxK00Y5oF+ih5UIidEGi6bZ2UqPHTD6VmfX/RbrNVPdJ
wXpJ1aWhRK2SexSzBZgWkK3LDBnuYSrDEUI5s1yywxqrNLXRHDDamWh7m7wT5TZVCwTqVrEeMMuu
4mA65Ir7Lq1URJPuQADsSARqDTWRg3K00Y6ko8Y7nmPMUXHhREjHrL5w6WLzguGldBe3YXqTY/iH
Pf4Mv6rDsUyEXB3X021sXT9VN6pTIMRkegv+onal+cfVDLsnpQg7f4PDc+2pR/N2XciFHcLguhPd
CGqOa/L8G+Q948wkC1oHeb1AFs1soYrspfOIfD3vTr5qtWQc+cZPlU6dMZ6QSmUXCCNH1yKf5I8v
gfD4YhbujgKFjC3AxugGTeZt+/TRnAe+JUrbFVodTxzGa0+ReBwc2W+QqciY/a0en5cIZhSJEJBf
qJwt5CD4N4aICrempWyaCeK7msVXI6lOrS/ziiMuUX4CPq++FD+Y4Ponqln7dg1fpfsT2XxxesvA
uFS2HSP0tghSX366Yra2f10eKbuODn72o2LI106X+2NZjQziXDZdIJTQifjKhNcqFq2957BoSRUV
cJ/2UHK7g1ALLODUY4YBJFEqUvttNv0nIgMA7XWjsovMfyGK2gg8fmW5I9K9UDgT5WEJobn5NYu5
b1M1PTHy22//9fYz7dKEXddGk3jgWfx4AdY0TQRf5BalKJywYHd1+ejRZlxma8VWemzA/CbfWDGv
YSp8IhihDOcqPX0A8bKQU58gMeE7r049GW6gZ2d52X84UDMOXViaek2fS7Zon5hEQGB1/Zl6whck
haKCmikimJMZXmUe4bXNsKjhWhVoA+/VDokNOFTQOsEZ7iRQn5cj7NHWd4O0gIF31Qg7+1KEcy/C
G47d1VMp4AVAiyL/rGc67CFMEyosR8G/9XtueHTtOU7UPKinnXGFSBZw0LeVXHueSUzAmWdY8Tmt
xgLxigaF0jm2BrWfkw0mXTcbNN0fjvGyvaw0VIXzuW7IE+X0hO5p2OCAXIoAM3nrPuYqBNYQXiiT
WXIIrbBcWBRHjYsrP3ukdOkhLlHkU5Jjbtm5P3Twyb5Kb4X0PniBtE4zN1XzCD/J3DgqWRP9r2JP
2vLISgaONChG0zqygpl9iz2fi6tpCORRQsBaOYh8/b9DIKt6tT2gQUsp6Jg+gtKydS3GMnUiavgr
kv8q5kKSudE1XM1S4HTv7N51SzseRs3Nn2m5YO6y6pT5Yf3Ut1J7xci2ncg9Dz7nrM96ZXkHqs6l
8dzuR0TzE3qLb+ij+79xZS8MJSV5oMcQeVmIk7OHiYacs0hQ5wKXuCPa5WOWGSPMa96jx7TekUln
c0mbhuNiCMEBXz6QkpwVup+87x1D8v7X8BvIxE7A3Eo4HGsn9QiUT6OnaKaB4/Pgcs7Hp0I5hC3Y
5CLW40wsModNjEg6kt4/3oU6C2/aSYlkOCE7y16EOoJGQy2H5/bPFHhUiJOrshuLrUlWTXty+P7I
FvoASOmDp3zSBB59yLyDdWmapG+iy7nXh+fE9td49mlr0gy0L+JK83xHvFbdBAirzDWr2LrRCFz3
IISKZkkzK2vkS/4lb8CN18rtNAS3r+ATKwbgZoW720Rf77H3f4WtHpo/lHfZ6HQfEmvYTM5kVN+K
/Bv+1P3/+xm5nOSLypy1aDA9ML2IFfqSTpbKjv6Uc7QMWU0vtO2bkWsVpcpfdT0GNCd3f+KATqEW
KJDzVj6jOMaWngIfTDCWpIrB2TuId+v/3axNJ80xwaJd92mCl7D0to4ULV7c9zKyP6O2waG3LKk3
kT+cnNy3JeOUiTo8rmc3aVOqJrm1z1YOPYzWK+ozmNgyaV4P/Q/IuMq1pxITTrhDoylh8dr9ocaQ
VsVXU45ULj+Ai3/NL3DQ6ln3ysppLLroIgMopo5+35dl4fYYfLhPFhDYA7uIwG2pDuMy9I0M9b3i
y/D/qT440u6FjRIIChuasbpuz/P2pyjxFk6RuOzsBm7FJCEFgYQmKrrqRFDT/0wmZuohQoi/IcK9
ml9l9SNt9+SwAmxX6oHws/AWKF2OXLt/HIWoIvO7B5cDXuR38C40LvMh9bIqn3yMc10rm3svxNHk
HVhCA5VL2w6EbT3tTVa3AFbEkOie7+9wk/L6yOBWVUaoYlL/BxqtG4uy/SV94xULXrLCn4ZDRj8K
rPw5dFTqJE4oQtlV19rEQrXMb2ZnjwVpqExI0LuLp4HuPH26TRuC+zGKpD5/Y3SUv7Uv7Zspa0Ew
7JOmm7SYW9UPIyl3zGZnKdyZ1wlScYp6fbuxpDsR3ciXqEff+EaPEcEDOFNmqLi7r89VSCA1minQ
+8mibAdmqcRC2vtFYXrDhHExWcw0MxHeYTmfQhiXwjQ4OEurybZ/64K66iY3k9eEN0B1S/toSl44
Yyixl5EmI+dRXQzgkFpjE3oG5ikAuFgw9/A9QpbQZeshBZTZ68oRJkYIzh1/kbUT6dyy3rdxruvr
a9bwpBPo1BTMAtfLLg6HwTfv4ORZuQ0e/AUdAF7kEU3MHhBCBOayqIUD7V6qw4pJD0ZexWI4GZZi
jy8CGV8mOkvPYYtrg2KUKDmyGBAiLrK+BnguhKx4V2/Z87vRcETQ/NqEoofsmzweygWsk+ey1My0
3tfrZR3B6KbOnQ2ZkupClJAeYzrnxOI3DA+5sM/XvfnzNJwpmx/bPg1K0ax90BQ+1urNG7SJ1N8A
BjxlCJaNL2QgMkiZYj+lSVK/CnmmrqEugzptoymj9yRGFkd0NjWHh/JRq4IH57xZgJJCca01ds4o
lJXZczznSbmVe0d6TGZdVq3ALhToLWQCuZOvMNYmYf+8QsIZOiDwwajPyW3tLgWvQpD9GAFFcoQK
m9/gkFflrNzszgbAmhHji9r6sTujSUj1C2dvK7bbPr5ELNX7tTQRebvLD9O95LXnf3q7RH5qA2v1
n4YmAEZoe1w7O5a4iYcE3hfQ6PnkhbuioEI49t8Q6H8/jl1TrIsnHsjI16DP0K88vSH4rq1/pZ1S
gGJTM8kNOUE90LzMq6j4X3GtwWOaMLhP5DwO0ZBlf31Uk5iL6CxsHfKwaqfs6nOGy40skPlzUb0s
qd40RbkgaezCEtLkoMOwt38qsFfvhtvl38DsSFEvnrkhP2Y9q1EG86Qe+AyaI0kjqQk8Td8RmXtx
/qzJJvqoZju0e6SaBaaeE+TPxGjG5r5Y8BGuDFDvGmcpDrrmtOcyVyxUnRjWcg2n/7vPoeA4Wg31
vCDtfh7irxz03zAAu/WnMyJZCWOaF2vWuBuLRDebr3I48fd1pglXq+29kzgz9FxkT4PH06FqQcSn
VjjBo5wULBTMOaci2GWnBzcRECwxmTyAWDjpRn7PpmSWiz1GHgEIpezfQrAxNhaay0/RT4mVtCHe
CmTPPPTGm4fyTyBgy5jUiZuPKLDuXLi7yTpW0wYpOGKGC9vFoZvrduGSYyXzWag5+xINN+FmGv7z
u8RRZ9RHpeGzPj5qteFidMDQhl2kPTtpcxw9Ou40eeDpgXy1zqPE82NOEhQOYWMDlnjECrok+wqO
qr1+qHG+nwyl6FG7YmzHWsGpH6Qxl2XHQTSkp6/BFtdyX/TU9wuieE3mg5iWSUTqOqoVNtlgASr3
NIyUMLWovhmdLXmQJJUdcFAYaJF4IAVeXdzdeXVmvkpabHgUxIbKteAY5mHiFrLGKWzq7G3SjGtr
87lGd+qILHmhFvaPqysW73QG2EVM8Xyb4hLXEKGqdiQTC5ZHq9WivxEa+BuCwjsgbC9yd4KRze43
fOOAPGkm1lpuKCzAGZkIHWf8VZrPVeMwpoYaPycrHUTwBtovGhBNQjcdGxHcyjDcMTf9KTMxKuIR
Ug3frUI+Uq93zm7GjFSf0RCenCV4Zj76Cd+E8eVR0r37vDhOfp3aAWFb5Px6HwEBjmPgtdCU6H3B
MeSHG3YIcoScbFjo6Ts0LlTiXl+KyMR8UlFfn5/duZHNNHuOSYZPFweNf/lZLTsbYM3MoOhSyJTP
JKqAOTa/ralJqmH57urhuj9ocW9thNf1zXNbqr4oB8GBsLEpU/EuHdtO/eVSZBDSyTxWG+9/9VUV
4oUC1feq4e5JM4lNx2O1KJWu8AysYtD3JvzsS8zZ3kJ3TfJ2jjgFU/FH+C+WLroQwxmVLPc3IgMt
F5hDNwIqsoU/TK8QViNdUH8F8v93RHmGTpxH5olwTSQOBocE1CFGh8QG8wPHMZR3o0lPZQaU8A1C
NwTIoXas28wTGHbxINIdARn3LZ4T9/BtezeEk1Qu703z2xxT/4aB32Cl/Z7/PEob2v1T0KNbBWfD
CX/1DRdCd5QwtkHJGSkgEVe3S08jxUyjQ7A+/vnr4MJEO1j97SNA6qJENSjIxAPPKcky4feL2G1W
swRUUJHlYRATkZDEhV1zAkbdXRofTzAYfT6j6zdX0mgW5konDpqAsovv48oeRQ11v8NUGgx+9HBC
VKdfNl6bucscLl/c16VDQpAbfqj8FZLx2712MTZ2vgHfUamZGGSGDXN1YWDnKnAl75eG/LqCcr+t
3e+Ys+njTRgWO4XXZ2JfnLrOA2AsC2OzwQp8lyDFqc9BE2wGQGiGBHwLP33CxG8TibTsA0GLZuqB
o4Wf/Fv+af2cNMe4F/6L25LkEl2QhC3T61VTAShczFuXa20jOf5AXMgJKJjV4PyZlf839g28UZs2
P2V5ImG061XxWC4gZkhgD9zUnmByUAED+vkxqZc3uZYXJjFm3KDvLB4Gg1wrhKW7cQlFI0BcYCqx
GJGtYPXKcme/jo+gy08CW2gsE1HBsXEC5nsd7vR4/N/Mi4QGll5aQm+hnfglk6d76RMW5zB4rhm5
G2ZuqflFA5n91kxZLjCXvh8eAAwMavx0bQs1UJY91sfyUNlHB2K7V4hI8/BtQR8n40hMKwDT6I4U
JXsG2xVbLoOlgU5i0yjO46u2e5DGkcxKNplyhAsBJPVFamt5DOhqzbji3/3/GgbcwZcCJkcDwMFW
ZJdnRMNJ72AZ1D/0Pew9TNHTEvNtu5f5WQ4o7WbE1xP6xm8A71sn0X1NPEcpJ7y+bjhYj5fP1b9F
eADeHIgBbO2opMTBnjtZI1oZzfN0XE0imjMdbAVTodaNULNPbfEC9G8lkpsyF2NkF3kFAMW1cM4h
400U61ka3AstpzeAqa5+1qunqxwgkXVP3Zwd4IpWMce4scTBR6gpBGCipR52cdOKa/zhFRCYzy/8
bjaFbjEmtGJdnWPTP6opHVS/thls5Rkt91rbDqyk0rhWoqybX/cyfnqZu5eqplw+pnZjH/r7SCVJ
rk8S8FKog6FD0STqwW8YYcgvito9DL1N4K/NfuO0aUG92F4gJypjZpQRk/ssz7Op1C8b4Be4yLKz
/Xla+VLsri9y8pv98IdNvlRt7KUy39H5V95QChgRSPar0/hhESZ4+8ggeK11CZy4W0MdiNTmiBO4
kWa4kopBwYBXcFqnWzGk6F+oLX+IpwNHwX2yV8aW11M5fVcU8tOgRWQKKgz4zsQ+1btyIX4iVlH7
FafhrWuy/XIEbSUwE3FWw1AVlWorNbH67JGHmAMnxEmYDPTWBckOUv8hj19nX61E4rBn5SWGu6Ws
jK8gwaL8KEW6oEfo8CA5LfyDRfnmFIjmCAW9vDXkKojcNbd86ACBOD+2z71qG9TpgfvlpgxUh6OP
81MwoNC4x+Vr2JXCkYB9ggH+ylPwydgZzSs7c9wJe88k+e+vXvabv8KBmeb/Uaq9U75vfzkk+rRn
FoM8t5tx7l5BNewpWjprg1RQfbSvd9UZkQj45+/mzeX2O93ePwhRdG9U+uBugOGdryG3m5aNXci1
4mWrbMpXk/7F0hakIv6w+0e0nuWduMbajF6CVp8CVViechFDyU/Wv/zP1zFVN7F0AcRD/rpJp8O4
8OGG7Xr2TFm3ZS7F1RzkZL3Wtuk3SQHb9QwqiRbtq0UnFaUua/FwkRU8C8DGHJmj40H/TAEAoXLi
LzsfG4UjQRMcWvP854LP9DElZ5gdi6Oc+OpTfpicMS1Hhs8UZCv8rB41GowRoE71IsdVoCjAF/vl
yyfVsdVVG9gfhpjOI+ovFgjL6MGM9qF/bEKqUVNlYG94HP5pxuIYBhXP6OB9iKHzLQOFbfnb7Rz2
/Zyvog6P5W9ng1Agsp/5GrcJImmhEFt2hGpjvJe6rLYVCJMWBHGH+iTcgJdCypC7u5PziW6WqLhH
v/FV8Nqz5q7q+eZrJ20yUy9fP2WoliqHj3MgJDM566R/CFOSAfuVD9Wb28bkKM4iikL3SUlYS1p/
lyangR4AdVBeObmANVRHjWJMqtVgJtegCn+QG82vQsYrj57bai0XDcPIG/vntQxOqPQnfMHlvNrd
NaiWU/zFfCWnS3IGgJrUmvGAGmePjhE3AH/dqcGlS8FdnzmBqVgNGY6OmI01i9CZ7WaKJQ+ZgjSw
vlxWK38ZW/vwgFyhoc7u5RGfvnbJ62kSa/6zZMQonxt0+KhhWrsWcHkkMOY8J4CXeJTPD4eM4DYW
m0R2wUN+aGbPhF66+YW6Yx/If/lh568AoMOiMebeX9DqowYgj4s5vTYSGJoYaZsnV7uKvHJfHYIV
fyjsw/zyjEDADOlrd8Jmt382+r2fzStyLrAJzETcnxoRDqGcUKEuHfbzVDdojx6agS348viwsWCi
mjlonD+ojXXRzv47LfRx+ruDgg75id8ein1WBYgurKmuwl5z3b5jhIu7tWw5wclpB1iwLDOot4ZE
gUggrsMJGVt0QkvzgGvvsf/BPM4pvTKXMeE8aitt9eV5swK849Zt2BVWrhe4CPPmuQm4CwhWw5+Q
Sdbb8f3NakwQxfQMxgHu89Gva8TkxuY+C8LiwZIyYKWcz34NNgnv8KmcFr4RPAvPSIG4N0WuWXCD
KazYhJMyTTIwh8DpL3a2xYjGlZQtTCQUiNC37sVUIYf/oXV2/HLySIvq9O5S+3/h3nAxdb61Nnfi
UsHqgRHT4Ji4yuGJzJIwamrX7p+qVOpvnfI3gUwDhVJ+pKhi8d8qFE13pbS2DCO34ZDXytlVCcQt
oju0ziMJa8xv+MSM9pTzk9YycCwQMNrGugqN0wVykoD/FN7p2761Fo3YOIjmlX+1Np/QGaPVVgks
MRyfdRd4VOqkFBKk26yMVB5nXPuqNpzjUBikIZS4UD2DExyTM+8fqEyMWdHk9Lc9qPqIzgnaLoVM
2YqW93unIz8wKwygg0c7lYU4kuR6GP+gbaorL/q0AjdigUnhpr5D++lUo5menf1H9OsHT6Fc6SNU
+D6zkp2YErBRt4Kmd4OFbt510kKLGsnJErTq9DUUOZ4qWjeC9PrvY2YEmC2mMnzxqDri6+3V6ITl
TrDn9d7Uxm5PYH+VXp9/1L024S+Cn6dRZnrvBEiR9NOXlwoJEROp31kiYwK0rqRVIq76BQ/O+HKI
/kviyxGk4qMQYuun0Hj8bA054QcHguBiDxM0brLjEZOu/mpRaqpuCV2kjWm2Dmtn/8qWSR5jGLfJ
ofVjZxedSxUNewdb/qifzuIYmL7tVMGh15OJE/KJNNaHhXuK//NvIVxjipuN+yLBu/Ch3TMW/VJ8
BgBxJkOFDRcS3gBtspVH9pWwsy0cM53yfmDSDBABGpd8AEcWxI++8EIwzf93wDJLtJAMhe0nJZUr
U9HiKl3snO6zlJUOR7eznQuqhmbBXzxMDpETQxxSe2thJn0upby98GuTouljjw1TqVqhCvkjK2KQ
Crnua0UHk7x4EkIAAJAipSzvqk74G/uaaypx1V37DP42VBPbETOZHl0aC1bWXEX/ur8NdbiNy1Pl
D+KfApu132u64TxbA0397LIkbGa/pPF9SuigYckKDy0znh/TWKwcqftpsI/jMFydhGhA/szkbMnU
/9Us5VGzbDxT+RuwErcQ2z+vFy1/GBw1GaSmfrC6iJT1r7h3EQvAUtC9/FCSMoYmUdB/88WWfcKY
zTgPIRwpyv9ChizNGwXTJIMkiNNFw8ooZOxsVdyw99xVIr7tXyvxgV4RIdkoQAmYyM0h/zsmSv/3
kRWgHDomhHELzF8BlvLXZ2mYKOCboA7U1p8xuCCusjd7kt+wHqrIhQ5Pp3172A9OlwgTsutzYoxN
nK7o2nzOBpW1pSQ7k1gBv0gzWLLFZTMQjndLz4KO1FdVyDPrbBKeBBr+I5KaJHplDGZ9AAvcXW7B
BFCF9GgPJtAfuIup9S9ljjRAotnZuTVomrXovDuqks2DUjE4ukljGgfgiLMqQIr7PUuh8IF+Uy+N
Qm2dQUFveA0I+ogl1LHlCZ8MP5tS6c38tsoEjkdi5srxSx4Vi5TYmqSziKDe+0T6Gl/8c3HAJ0yh
Yj1hhFcJB+rR/KaXEPE7lIhw9HsLQrFX47Etcw8Crw7xK/9J+fu4Ipq3d9CA00xW1HnwI793Kzvg
Kgk+74zFIS6xzoJypbuuakmscmc/doeNoL8XuMlHhSZAla0mQLkVJ6bjcj1NxBCwGEKFCSw3+gjS
XUDTpFkshjZgBSseK1zlGo86aB1YY8RUBwc9W0RkwoJoaqVXUhOzbVunBcfegZIc6Q6v1xXJE1Gm
gyh7erIFxQjq+DKphTVWw+HX5/FjGncs49M+yDGI1Ih4aPr9b1PnAPlHu926uerBYOEeP/hV6/IO
OrgofeRd3d+VrArK88K9wOxSIS0C8rKC6inlsGJf9hAbot3ewpIqBl1Mxz4usYS4W/AEegdFqzMo
QGRk9fP/cfldPA9VgS4LmG3a+DKLUOJrRZVcMK5hq5vmUJRxh6MY8kDcpToNYOTze/B7zkbIgWZP
nsGeQmyWpJIk8EOVXyocCXTw2dAGcfs0gtspZoSk2+xWm+1rZ3liBqpUN7M3ywl2TxZa37REO1Og
8QZ1p6qNz2L2glXzP427k5mC2OGxyQKOzzjYbeKVNMEFlD4YEkor1tDNJtKBnXHbpmC8SxiQjGqA
rIWTAHVmdM6xT2/7CyJ7NcrijFQwMADVsbybPD/kumTkx3mpHWdQzLs2By+sfgdpmWK9pqzIHRO7
+OFHvvyc8UPiSzdHhiKEMwKbbNOcL2nA88zKgVtTaikE/hQGet+8AxWC5jEEip7CX2I/Uvh93xhb
YGGUIBdcr1t5ZKJk3nUfqVM/RqitG4mzT6b7Oh0GnGjLwweWMndURsDOXJo9POCc308Wp68qGuyU
N9k3HmTEIVh/0T4kGYv4baBvnsyEjUjHngNdtUfD8LQjFMmUd31UcfDcHa+Wna807UqDwxDV2Hax
pA+pG/IlQS0yA0ktXcdOiCagvxgS3iDExKs0KDRVacjVNzHKc5WASft1koxHY2OF1f3JpC7boEi4
GyRpbHsSsRbeVpAJp5mouzDzPDEzy61O1ytkdcPMjdpNOY4LdR3mqo9jWGsJye1bRMJIwaaKKIpJ
psz15KiMLyw79AapYnT0sOgzK0e/8ZUPcW/lDtpRzfLiXY5+wrGrZhcud6FXzoPya67mVbQqXpXN
OLHeYR4iGhtIUHcerXEwPOOoVZUE69llTfok9+CKGJEM4lf8s2iEvsFELyt4JMrWQGd8SvWctJuL
iAhrDqgteF1Mcd5woftpJN9IbSk4ck8Otvs6QhGJ8xby4GLLwwUF2rxshX0NBsSEFMIapjSaIChR
Q7C7l/6xgdRlYg7neEv1YnQlT8pWt/bPjDuZ52GynwFoGbTa3KZS4etSFGDzxMSZDU4N9j2Jmujt
NW37YtElFul7RILFyqabvo7Y73WAxROcx/3vS39lcsd+93jF/UZySem6/zioJ3CrSqzkuHZqsZwK
mf4KrUDkixPMRu2+EMJhyEZKYIrU72WzW8pZcAVulDIL3OgcozY8cSljkZSdbCgjq+4h12gdZR18
WV/no1Xq0gzlU97tX+6IU1oNUH1e1fg5d/97Qzmx9KGIW+Vm0wUYx3q6o1QjE6RvoQtpEupAKOF5
1WJufToqrf7JRq2xe9SWbSzxqnqFksXsYkRYAkYmpLbYzJ8fK/Ni26a7Ij4Uwg1n+/HgBZpKr8i4
leuLhvnG5n7oGfHdlN1dIQwJx/lqrsS+fNOI2pdjq6ujDoXqmorA/jxXo275HUgW+/34XWrgYk3l
liscVyv3/G9TmIVLMS1RIGA6Uv8iPC/HLjamMOkCXS4vQkSzzw3sWEC6JiBFAFFlivz5Pg+bQU9o
mjTbqm+8slS9da7RUAFdLCdvfIZY7oa5ZPs7beWx6+O8/9ngb5rJhOL50zwuJecLf4K2U5oNXEGU
kaswR4BWIi4Mo3mAUuEbKSWZ6ku+0DYMQCIZ/8cdTULCcoVyXw7RkLwHDNDl3rMJt2jt+ss5xoov
Aqdnrl9CS0T1kLA7DJZD5eeuzuhdM4nwa+a1BSTNq9vF/yGLkVcqNLNBF95nR8/6u79E5q2PNuQr
OP19GBk0hxVBZkhzzLgTHsvRzP8OagCY8IJIP3VBx3JNFq5j8K7gZgYjEev7hiL5wYlbWnULHGqh
JA9TCI6vAjY7JgysEDPUvRPTlNhyEYSQUrZ+Ff5LkMKvkL1mDUsh6NVOSu4MtovHRJjDe1LB1FUy
wFjzwk/urPs0+JiCS9urr4rJoMABdrKP4Red5dWp281S9XlhpZHYyNqueo9MNky7sI/98wdf2nId
GX4lzAPwCxdOIV18DJ4VckZDHqBYs0CjgkT8Ppn3aaZkhip/o9WFPTSvA4uWwJWUee8cyBOpBhex
QKnYZ8Z8/yOENzCPacImLKgXL/dZPMfrvz9a8T01/W+HeJEPSH97LO7DL6IfHnrgOpPK6ZEua6nz
hhhYfGIZ+wH8DyYfzOe7Vg6P0RKmQGcMOfLHQZI9TUIxvQj0U4wkdHB5SREP2OHMQNHpM8q4a/h6
++jkeUR8G/gNgzySKpb7Pmey4X+wxduZthdEb6FBItmeLUb5oh1dnCCYkAz058VHPyRcyT0Pkztv
KWVuQsW4C+00c6RDmE/FNu2ozZiGlaLU/4soWJm94V7a9x+wfP0CuV2EvyxT820HrgZw0glV1V0f
3wrx8st8sPPH4tUK9NzOlI4CapabpcpIGirOUlqnAsf5mp4YZmtX5S/t1TcVGlReQfzxF57yI3Oh
zj1AZxjBzImOZr7xYiXKtJwVLi6L99S+WmajDgecYgLOs/++uaPa01qPtiSjN+4DBbOM2saxbjUf
5e5vS70LVRbOGSXLw4jErOtlW/rxpnM5XQFKgfNL68TJXP9ouHPlr5Qxb+q1B79MtuoN4tmbDJcQ
OdJIx5Rsy9pW08z4HFZ79vf01rF8lWSSGjXJN/5kjUZAyHbCSWrKqct2rHzDFpQNdR6vwOkDJndm
MO/Ph9T0aXRtp9OYomNy6hmhAI0zVrv44dd5W+jF1M3MFgla1SjkktEQM24vTVunG+riAUsSyKX+
RkEqjRlKCMNv0j7OTAATF3Jmap63N1L9IP4s8YqhqYqwr0+zbwuSv/vKzMtYHKrLpBvHcNCDGEzk
OMUG2s5iAucSoWUFmWnOClf16/X97NOJ9lrlm3DeWP19Z0I604bM4XKsyV0KlYkPwVdJpES1wejt
EINOg1PZRlK+k9jQJyOPLs0rYcUBptgCkJO/MSkFJaeNjw235kwN9TO8erXeoj4leeFDxTHo3nzP
zQswhvdvKAB22+xFP0Y5Xln1KEuSkCXsQmXRaDv4z1YurAdV/rBUTFOoBcwgEXkXE5COOTlRbCMW
Q07EC6tFDj2fO2HgF2RVm351OoNvb26UQw58h9pnwvnBdWa/xqMzGT9xxgpVvQ7zCkDXRwUBvRyM
oW5fkrFRfeTl0cP3nRRu/vGcsOGzX+Fmh4HbOO7n4cnjZEDvDUg2TvMh/wF1u5WBpm/TCLi7nld5
0G30Cysx2cwE5y3JaClRDknKyF4LZwdgTvhWs0IC61/AFLj2AP8/2kTw19dQFrbnyce0V0xjfP53
b5sIB1Amxa/dS+axA66V0YqdKF+tzpqiO++7bhpCKNgfTU5IK1DU17lvjEZ8Z1pe0XiFyH6GvzQ2
6JLvPmBUXuSq6NdLpF3VB+bKewYL8vj8TXWJZldFTbDa2rNOcMLBLuIwegMRLnjTg7n2NRj9nBDe
i0ieNieyjYPBCfm3nrSm1LKfcEbU8vQc5kW3/m3Z23QfU/o+Q5u+rc51BN5VnTkaDPM5/aqlAq5J
r9dvDdMVxQtDfxgPHZdW3jIFy0i4p9FnL9SbIg0B8VMy9ofgv7e5FGdKAaeZm7CedJWE8awqq2QQ
5F5wnQIuZQfPIc4YyH7luK+5Q84PdkStQ3Fq4W8kupY8ZSTzlhvxJPYalIKUoer1Es1x2Gor2Z4u
hYlymHa4eosn0agQFhjvbId2x8kimUvlCGT5R4UCr4vuxvKqZsPWEqrbiJ+wPiFRWgpjqX++1jd7
uPERMDBVWYl+2HDG1frsZOiQ9mIf4XXILtv7b6iyzovF6mFYpAOMPzIcg3XCiiDQTpWWZDHuz9NP
kRes+gT3CRtI88SY7gq8SiKRUecgqVuRUPONrm7wjaorY0Hli+ooIHGpiZNjx3AWuZQ46e+umldK
IBD7h8l4zOmKTpY2QryIYk2qfCrEQ1RN31BSqF7uw25bNgqed2tQceg3pDyqJn+U6DBgy1YNMS6L
yW2vZ7zv99MtNFjTcIxMMFLSqlkbdutIfe0XNhWfYRrmSg5foWhbHw7DlXhv947Z5ee7CwX8cYmL
X8iuBnR9maUo6T7ZSc6Fry2OPLmk+8UW8PNkygev4pC1f3NkDDiIzyLqFnBrEup7cgEHrfZSmxh1
isxLQGycUr68EoFmip0A1W0gaa6I5tga0CwWcDg58RpCWXWTmA7kBPL8+dmvYCOBHvafbkwucyuy
YzhCucVh2vLg+MvPVupEG095j3ofElW2wqeo9W8TqHWDRiBdVrS/Drq59JwySsIPtXd5V5M+cPBN
DJc/XpJ4ouZIYWh1X0YZfIT7yiIZLjNCrf/jnM2gmVjs8PDb9pDuh8etFBpSe6/pWBb+JGDxgldU
Y3Tjc+m0sHJOiDhdy9CMn51tHytPuTfZDKkpzrsnfWzc5CCZQGeC6xoU4hy5PFztZvZAOYPji6wM
r0SzWXaSo0cCzXOQHLg6+6imp1UpSQPIurdiuGeWl5NvEuOQvRWOj90Gt+Ao6Nijtw9by8AwRt96
W0y7tCcO/sONWklI318DqfWvfHClHy4LQFclg5aeqlJmaDFoAxRMitgGBPuRkxTd4DT1PgWeZFDj
3WLnhWC5v96OvglnHZ0+Mt51Mv1KdVjVD8w59LuW4xJNxCzNsX9C6FhxWe/zh8XmhGX0X7Pn/gTT
aNmK7+rMzhZERKd2cS7oHXHVQfYLVFZDOlP2KLMl0gV9uA4EXUNqRxRXVQo6Jw2bUNSJvBA0vACt
LKM571amBNzX1xM3vixItCxyudTUgHV7T6MWpcrcvqDfO+oBc1KSvWRjo6z5jrYOp6rHxoJPImUx
j1Z8rSzY9eR0SoTNlrooK8+8Shxv9LjcvWJ4wMoh619fk5rN1txY+BLzioZkgtNYQTLNS+pKQZ2a
0ESlt5T3cqOXbzr4Fz27/rF6oe0EuEULOPZmOEt5x6HJ0F4As+ovinSm3MrhB/Y/ljPWX3lkXETg
+w8vVB8g8IGy/gI59Et4ajgNKJQI22xuCnH4OltLL4tu0rX8dYW6k9xEWh6B62yvTWI6gi7Sk2Vi
91ItHrx+I9kZ2hqDuyZvRrSmNPCWhzjvGtWq9hr7jn/FKjbTSmaRMyL1V5OseeC9/aOgGkAPoroW
f4cM+Gu43blReGKdmo7YAsz7OjBtI3yV2KLg9x6CF7gs3Zhn1N9doBcG2gWOKi4US0dlkG7kMLSq
viFZJ1jKvN964sHz0GBe2mX1NKmR2BfgxVVf0xG/3Taa0X7BeDVo5kdpx4rSGZ5Xfk8qYVoIcN4Q
UpWFh6P1Y0WryTxDt6Tq+SeoHauVa6KRZMuOqrp0AgyDC9DiBUfFPo7irw/g0ltDQeUWRv3YkHrI
5O6SY4VmZdGvHQ2mFy4Xvd8/nbdhFpkfQNeFjAdHl3TZeoYhKWPGydmowETWvy6tETsbYkxf70Y3
pQIkNfDIeh5yTVzMyd1QZur5csC7UbkeZqeQB1te5DIpHNdYXZcnCPekT2rIjocCFz/n5vCx60vD
6EVRj6HQl3E51rlkViSbYrxJ9gEzyiJuRE0lBTLgma1uIYiZ9uOIULiP6e64cj2o5V2y7jyRtdpW
jTuY3lSFlXZKTUohIHy5DwM0QWt3eOGMIUXoocZJe9xte2YBOgapxHz96cIcJRB3EoXbVbpU5b5k
vgZtCxpDa7yPLSyLDPieXd+vrnS9PYqjBL3zincUAJAYi+x3T3jsbPhliyBSTI05UM5f1V+pOS07
PpGeCakiEmjeYahYU+GaXkkEQhOdTjUrLBrvyRjU7v8Qs9+F3AkGo5Ob+ZvWoph4cOe5UFyEsCHb
pZp0CFlz/H3YloGvS2uPTShlFM4RiQ/kfpqDvb84vis1fe1XLBOtC9UtW2YI5gfFdgHb8vYC066V
5cdEp7QgiWHmZhjie+CIdgb5u2QT+NGK3+cWh+dy8WSgi9OcyImSATV+TSo0C7GFCzYwzcZh6gAD
SxrLYjJ7gh8XoVwXW5f/fsJatbJtd7u0/gfBOfYZ9d67AwpQlvQPRLYHvs/7aH/zEhnUJVApFSA4
ZjM+j7ON5ehQix85mrmWZ9FG/bYLv3vDtOGUfPN9JPbYNLGGAW11ypbNEoBgpGWHSvEorr8FAbJ4
WKHp1YWBBQHMJBnIDA8yCo49JbACm8cYJ+vNA4bXkIO7Wdzwz7TVhGMcpiDsowtCH6SrweWtZ14P
hc54o4bO/7BopASM46PCSX42xepIde0NpmSBKXKR1upQHMkqsgB1nnXme0L5NeDTcfqE05XDD6W0
PJaK3+NU3EMw+I6CXY3QXiQGHPlQBNgBETK7UL5CguBpxMtltOncwnKKQZ8pGMoCc+X6QvECbZ+9
KiyPe4178K0gHjMt9/BKXoKuk70MjqOY61/u7BUSQFEAKnAvXy2EkSPP55daaR2bidtngQqmqg3t
Xf84CHjLhVEqFq1Sb1KCmmRBmz2ObNYy5IvMEgh9ZB0Ean+5xS5KBM7JxAEe+9U5gCaDXLH+ZW8q
hiadvHBFymNxYY371YRB2sATnFuzNfcy4oR7Hbz7ka3BmIAK2zyQB38m1i+EPuVU4brGpz0VaY4o
eKq+J1zhzWPcDI6g1LsCkDR4Hsn1+VXkDjzrkOSzacvd27mewn6O7GvYBDPDPuLsokQlpUUSuPrF
ZuidcNmRImWyMbk8KeEPGGO1ycn1yGGsMKMEcleMSRPZChGv7kubB+kZd37rNq4+l3+GEX6+pdLO
OZpenrlBOWU/iMsC8UvPwaGYP/oy0IFXNxc0ZtbyyFpCmlJFpsRlozZWJTczIGxbL1ZyR/cVue1h
T6G0jLkIzA76jo85D90hXh3Gz3thAkgrogRRdnctJTpBqXOWlIbfISxRyJamsTl5YD2aVduFIkkv
erHuliXfRBPtbGoI8pk3vZemzaWZUjduWtgNMcKUpATBU+Ej7fhGBOtHIuosrjDx1awPqaPCZDuj
aGWixQ4jdAFMh5L1XFa3k7PYwgDVNtzelzRqHoJpO9yAwYzt5cF8QANZ6gXF+wP/oZgDX5tUjMGA
c5YX/OQuUMuvd4/wfMlB6YaezQVU2qbN3VLoUagrKSFl9hNtl25yoV0aF7pln4IU5NDRXGmruX3h
JBc35eocUvtb1AN84MQSEQT8dH/XaG5V4OJDos9/dJde2T+DfxbJUGd0aY5RaUP8M39OrpSb1Imw
nnTjMx3couMsvPUUn+I4aiTTTEuv8K0y3OF57bCShHE9pKPO+IF6R16sCZcmYJk2XWfDwQl3HP6b
nLlwVxYX3HYPTr6N9QmtcKQf1g8ju37t1QTJ0rY7oiBN88nbYblBNYuJdVhMtco6DG2435NQrIKM
EbKuzn+9seoK7yKCc9h7Vd2pDTwUnn5rgq9rhTTNLLbtHWFZzK/zvoEwMEqSZVcTlBtyVTVqWCmw
DruRthfX1GX1yt2eeU3TsQMqRM3Jq4cqnw0fjOIKlqiFWwRqlBSuaXtxK74db3qTm2mt5S6zJ24N
zNiaxHOq96BeSl5rnTkGGzMToCTC6PHfy3jIdq4YsHFVs1ZyOPU9L6d8a/V0v6LW2UmTBQ5BuGqI
dz9HmUyBIIQSsjwSNwsRHsp4kKEUuWFR2/KDWdRi6TxIUkSnBqsKzA/f/TseR0OYI0Rx7FQPrQTr
JlMlpaMlTHEH5EbpxZ2Rjs4dozUV9aYkR3a/RvQfHNpiBDnKo9MqUqpa/oU3VkXm10debiWLj+CM
UfGjuLEuGtu4/nKBrCWhztB8CrqCIMSCKZ8iFwON6mR+HmYkr4hkUggG3fuN5TkIogup/dLp6eUo
17osey5OUrqFRaJlT+5/3zXPxDSqDVaGhSQfzeNxMS2eCV0zQmHqytpekt/9ieCM6BhSHLaKj95v
m1v7Iwm8ChAn1VMr0rPU4tRvHKitVDX8XvYabHGFs03PwBcXXaSXGgnfpk0aVfvqq0XH/0cDehAl
n6kJHX8e/MDSsDsEUdWQSkf7npGfi8Ma5JJwzf2LCrM9jNiw9/E5DS/VLya8ueTAVnhR9MZ1m9K9
h4g6F8BuL28ZGEjVhUtgjtipjaXwnvYlP7bJNaYvLQ5qOuMhgsUOhJGua33cVmEqUedosGNUvswQ
fsIUJ249tB15ll+MGpLiOzUrFBRoEcH+yxr71jkS81PVjSM8jckyv8I05kD4Y+c2miLo4xEVIkow
QkNxIPFTZ4PO98mbBH/epyB7W88+JGDU+G//8cDcvWXNDaIrjzHINt6l6mdaB2NWgTQ+gnHf+EDL
PoffrHM1qHpiFLufok5jX0vvcUBg6Vqmi+MrFQZqgWvAQhqTBHyYuBEf/lUvv2qPljoq742LvnU+
BC9ZgeeJnVQFQZjx9j2hKLYPB0+uT0J7yxLB2lQH5/N8Z4zUOGGiocWIASnpKPDZI2wj8MKhj8bR
+KXS4PDsAEmwUE8510c1a7XouzdGQolV6Q8ELWFDxhGKsZYQF2gdgX1h6GfMEb4x1qFGqrfunjWt
74WhHIrN1o92XBug9gA1VvDGn8cM5lzC9MudJZVIoCexN6xf4OXzbbrwBgUhx3/mTWP6eJqubnRx
LQ+XMlomMe7jN5/VjDpp9N+QyIrHQhty4gj4x301GPLNy6rHgsqFd71W32TKjlTAvq7oud7oRBjG
mKNxbdFeYNGhcLzTtgt8QsyfYijIZZeFOL745U278xz/PHB3pQL1KXRuBnG6AVMcVhHwKs67aHRO
8e/TSbIIvQVeoe8EmEuFP0aqC/6sO8YmjVEdl3hz4dy33Hb+Xxm9ZpY3SmoaixgmbrouRXDdivG0
oJi82yRrVkGXjtdq2PUAIKbJ3gRg1EjuVmR5t3bmBJQoBBdpaD3O+twKZ0uWy/6QT5imiTsRI/3m
hE45dBxNoTlvI0Y947g4DnAm0BtWR9sAj5+RFSQATA0GYJ3v+YFad5cHORiYFaQBZYpMhxKPWMqJ
heKPoaoHv4kuc/yDNfFiO/Q6oJPahkDmOUNZqHNdzbrSK0zrGGcoR6XfvWjdxOX/XQktenKgFrJB
9XRsSDGcQWdP3wM/7XwjuaoXFYEPoDPV7Twu74NWi0b6ZEUmKTpxyXd4hB+skqgeC8Ua/sc1r7ix
QBVhIAOjWrSRAhFQcZEmz5A4TWjcAGjSwsiZZg04xPs51bxU+Cz4obJ0dUAT6DKjCoyv+5E9MOBT
xtTcmCyIE0bsZSQfjAwJ8u8Bv9P1/Cb2cfPnFDZBqCEoOK//a07dZZMa7PWXUgwLF23bfgYw3yD+
8OLgbDkd+A1OXak5RXYgUWy23drBZQvWcwmEv/9yS3jnJIbKyD9lHKxczq5SsMGSaiC7FLM3C3G3
vrNU6ktLtExqVU8OcTRPczLXxrLT2fVDDO8YcIx+RyBrmt4jv0VJExCLhJNwBl3kc1k8lZKwJk6j
f8QDjxUtGwaH6cFK/e/oJSmlZqkRQJyNsyD1NsiBJLigNOeDModaKBqoEtlwvcAmPlgX+4rIkeg0
50ojyzrTe84GQbGdbDb6OaONzt0t8WCMoH845KLeZLPO3QTcYe3gwlEhVBoKx1ld9esl63Uj9se6
0UZMQKnW61sO/sycYnAJjAFM/PNyeyDTmrTCSUvVaPfNjdcUgNS2Kt+VcgHOIOpH/WjqGjBFrq7x
m8bDvk6jvl4uOdUqpzPkbINuBzDhlDVkQUKH+phzG1SwS4ZyoI9qjsrxaiViJyP1gqH9Ni8uYk0d
0+4ItlksWm+pV3Tf9qSEgewOjsu5oUJfV75zCzrxsttJ714/fuB9BUUW0WcQT94k7NfOI+CuyVNv
7BPmYsD4Lc5qNfi6KaGmUwiqK8zhs0n24JaxcbAA4N2mKlYx2TAewfA3pxmFZr0tnBFlhlFU9zE3
S0DDYpExdEoxzInRGJinSwhH6/98wrcLxlnJ0FK8wjt+LuSvqh0cATo/wMnzY+XF7TDlQ8ytKkid
81eI19PCJaxnTvQQAseO6wL2wwLUuBxLDIwcQhSsb+VSg5mxzPnWf9NXO42y4FRNQM+dBtrXJ5kB
iRqevIgejulIocBLBinwSeEihbP1tpDNkuf41qO+L/gLpbRQLLl/MACXSTyOGTIal2EUZB91maLI
M2fCulrAJ3GT/yojPbKbAadQyVg7qvIUnS+SvX/TKaTRXfGR0VFuhWgXIn8Kh7uQ9SyQQ2FK7cjD
1PHPKVIzP/YnmY0vUCu695XmiHQAfBOgszYYbieFcvD8udNrHFULwr2VxwHyjMVVNOJK/MAYU0V1
tNqUmy/PpzmetpVdHme/BOu0BM0gJBTmUP8Gc49Z0pNGF2Ej96lRjuzs65PfDc5WuBcrclUQWJKk
G4nBMRjRy8j+nLSvniHaDbM57y9Pz1xx4scEq1kVKtjRmqFPRy6V4L/aGKrAEW+pV4tGG1EKE4Fq
xF7ZN5+xgr0UmbCxEKXYQeHZ09BQZuevKcZsnJL8y2ALnJhL7C0i6bU+dIaM1afUXhaPtkbiF/QS
X+dGQBuWhQ5mgon3VSTUp9YJdebfZE4hp6l2gvIA3QxjKoZVlomz1FxpndR8tJ69c7W8MSle2BAn
YYeB3F1q/+HHpKdMgrSz23Yc0Dpl9Vsd0IJQ0NuTNme+ML+lPt6f9BSaBAJDqZOaTArO+nlZ5MpP
BMczZjnV8EVhTUeqUSYT1GG1EWVsGi82AgJrVxOOvOBkli00nL0ZKfmadvALTZNQCBjArM1aER8S
tFd39W/Ykh7SzLAYXEn+UmpNwpTPuUwkM/Zk6of206ZdWd1JmF187a4Uw8EiQehc6RH5vo0pM04+
2Y+tZfXNkRy44GLeLJ90JIz79rc8oozBnzCYGmPHSUAyh4JsnRaB1YFo9oh6dpzr4sH5BL0Bgdlm
pHP0P9krnBCez6z+47d/Zaa7Ks3CxAtPPpetxI+d6ckg6vCVcBuY/AXIUuqINNmU5qG0Y9r4juFb
IQXVkORhVFGs0D0TnsbiBKll+wFXBpf3qhT/ypXn4wtQ5rp9K8hQ8Vo3wSkTSnm2kg3FYtJw5wQv
bn+iWRGqsJoWK3QgDkaljpw0a9cH59LLYuTgzeEbI4TIjByt3YXuPz+9Culgj0uu5Y7S/rxb2/q9
f/iz9PGepZRqrJTkyc9N0+aTvAvlDnsZfLao1dF4FhfacaK0E87xBKkybfUjTv0m3MtjtazUlq62
e1LNNOiHy4UW1NL25V6uQxBiqX/cxw1ypFjInZQUqwbCjvM745DV13HTnuM0JDqxs0bINMIEZSdg
CYzApEovRcaHT4cFzHlz/VWPzc6dlhMnd4Mi3xFe71RT2jxGssWWsh9emjGGYN9ADbVVcXZm3MOI
IheIc6uAq9GCO6d/4JA5AnqupMJUK4IyetgyaCpEwUA+SDR43WFZpuG477RtCTsYp7jTHeRpdVFu
jAYhpP/Nf7USNO5kZcbK2sZl+XR9V31O6wgC3cpY9Gm7ygBUlZp3hQpVRNdnbFxRELnLWFiD1FpE
u/uE5BtcrBgc23o8PbU1mhhpm9GujShsg0eXC3NicCnka1xOO/jFfZaHOZWjo762tiWmHiJIU+ZQ
xo09Vr3odoLSHmS0Vs7KkxCn/qiJb0MsAg3POrchGBSK7Sb1LAwLIkyZwxZ5wt1hbkeSOY97nL3H
fhFTtTuJ9Xwta43laIx60uh4+lF+0SRfhgNbKMXlQE1OBYcZLfBZ0N890NZ08XVFWlu2uijo8BT8
6tQ16+qbHUJJ7Xm1EOUX2j7TMQaw6YKjqFioNWjMVObxTPM4zeXGhqRjtF4azjqZL08HDCUXD802
+BCZZiGlcBNoSJX5CUz26+yGJ4ofdZXEabJ7nxfDWdk+Cd0QjI8dpxOZfZekZDaZe9jpO7KlRRBX
yv4g66QyULshCtGCVR6AtXOAwUtPLQfq/4wXH0PhCWZ7o6sNZyxM4ZMhgqAi0IV1h+n7MfbCoEz6
flVIfvxcJXnK1Rm9vfRDfn7fDqLaDWUwsyf5IS8WDTzfMHudBcwKRHz+e+57pm0kl1y9NRKSMZqX
Z08y2sf9Y93eOH1xvCWzqgK2Bd1qJPfjbBLabsoeT1vnGeGaEi/foqCtfkDL3uv/SvOyEDxYWM+O
m7n8fef+QjCaA2As994nHA+Q7ZdJBt5U+GdjW8wPemOd9thcWIpx9slBz1mkhR/9Dwkbu5RWkGBj
TwMUZV1Paw/HZf/T2y+fX+tztjrw/NdxBLvoReFcTNgDjLOaLITawwKFXJ2Kr8tqC0Ju/3MuifTj
lqKuU7Jq7/3Rj6DBZ0soYRBhSmhwre5dbMTMVrWTxCpTvO012gfOETzLVuN0k1lZj2t14yiXXwiK
mWu6vASJboxZrowUKjdbHU9OTADbDDByDUStutK4sjIgf9RY9D+o7AeOaOETB7apPf78sROmoohP
zYS67WqYanVA4uDHMQ6muqj7AoLS1rCG9U3XQMqGwWiCUvDK3Rnv4Wz/sIpk6khvqbGrFaq129KJ
BEGeSxFU3cuyjJ4EWI/4vXvLwPhz3CaQNkCX/ZWZ0kxpQPnXZUOVsScQDKhrjh/U5eaLARy+eOuw
rap/BPDyxf1LKsB1M02isFo8s093BerADPXl9M7hJeH/NrpRy6IALAa0204Zg3f7r4Gr+Rnm6iIz
BBRHOP70VNrrlevcWWmyc31lpT4fH43UUov+bg3dbS4NuY4CNUIjz7TAtle2brvSoVrDpcpexbm7
OnRkLIyoIUV2II8O/smk5DWzF+ShLdzbwmQEiofSlytYb0dxiCkSnP+py1hh4Yzth0SHSABWf4tN
64L2TLGjEeCHB3MvTNi/TA5o+3tUmtKcQG8kgtrgcY1o9whjnPpA+67AULDDbI2I1kNz7p3c9q0Q
A08BYLjD57sxQeNhalvF406O6jLfFUyBeAxOTQq1E69q7DujywRsoup02UT6QswtPxQfrMetGP9c
otf8KwAA+BzyUYcIScGnZ80bCAez/IKTS5DtOO1AnPHyu2AXasMIJXDV3AcMMRpZPxjvfTUHmC2a
ZV6Rn1TctSorGSqwuj8WznjEGGKf2R1YwxfIyiY2Eb0gqbL/Xqj9J8sYGDZyWaB7LzV0UuYWDKqu
jwwNGF38hvk5BaBPSWBSwZ7rHGAq3Q1x0girBs/YFRMqiTz3XTXkeEPZmXwhx1yepIwKGR0jQIDR
DIHnqLkzWv+KrPiRdlw4wxVC0ishLUjn4FDsizycAFEDsFta601jjC900wY++f5EZf/NjB2U0sMO
lyCCUheQMOVj5L0/xl/a0O7+HAr1B6KwdGfvmwcE4L4MSbG++TbH9F/GosZkK7woE63xbHgKFpSq
UZKeBzpKEOtzFoX2SwHBF+bnd135B9LLvr5EFQRbmDDnrPaTriMPrI0dnxkzi0DcyxQRKa9nJxBx
Scieps3AVIQcMj/KIXBQ9ZjXhMwS8EDo/bb7uf/PUcLz7L7PIxuhENPQuijfL+8EMZzKdu85caa4
g4yyqpv7nz2xkatiNHk+qoSJJA6Kzg2rPkOp+LRviWn1In/ocQMPpmm6crsRdE5XVcWB3TrnLE1a
8tCGfQ16dbUMejGAF/jC8Mi01FrpeRQx1IPVwYVkm9fnS60KQA6ecNJc4N+dcR0xIy1Q9IbbfJ8/
5f7FWg7UbbI8vSCFmVMyRyWJ7p3H31/AIon/9wAz/cC+PHmACmdMCNu2QFK0ZruEFuuKiW+QhJIv
CGpBptg6ZvzeVBzMdEN+v3QM9/B0ySrgCsmKB5SNsIeOBHf/IgWqs8jp8LN6r9yJcyX73IECp1Hh
HBaMY1cVbXkN9sGABGj3O4ETSHvYQjkZOQani1qGO8kj+G1uNAWPmzYJfguThO0rajwwg7mHA5Ix
BrF9sSw5HbEV9m3uvOUJ9b5ls0ejJ2A2y5FGjUwr/pLJCTtz0IE8vK4J1GbTnrFE2YGEmVm2T/0Z
1d90oOeays8MVsPdrWW9FOCbSSuiW/MEy3DAjSiU7YQNUlm8bXdWhHjBDSCnY+s885Hb5yboi1F8
Io1eXzX5uDJvQgWGMYLne60t7kPLiLL8zAdVASAviRDiNucftQ+g9m8wnzAzCpCsY5Bv4o6zxj0f
5RpdgLb3LvxPKLe4DvKLM8o8D//62C3XLbzQPmEn9wypwCxewoCfYoyaYT/LsVH4VHVMa6rooDk5
wGig6jPbTctM9oEG+Hnjy8n5AC8bwf2D/CzUZilNte0mCnBp2PJSe9y0kKoGEV6lYkJF19YmOFxl
IVJ1LOzxky6W646h+AOF1DorMKWC1bK/0k+WkKAPLcfctC1S4YHoEqE7cJxlJFkU+gPUSK13ExPV
y7RWA+qnOxUrFqCOir1qOSffg7HJA86BIH7U5ko9nnuYdV/07JovY08RG5fvxtLNncPQ4yAb3EEH
m2x+OvF4FH9EqO6jPfG2AkTXjf00xHZ49LVBhtLnFuwQlv2kEh670iXs8csQgRyw05XB7Kd98IWM
z2PU+aRH54GUbpHeBp9tJmbtiFcj2qazhtswH8sCZ53haMnFUCrzXnTuN211VcwmUPrSMij62klc
fCr+gEhpoHKlwNbmXpNQctSMk7ia0/3jfF79AU+watYtS+YccFY41dlPsEN9rIp4xOJ6mDF7nKoT
C7+rRvbAQWMs6JVb8i+/RZXVu7rGD76FNt5SDAzagDCSlHrfdLFMZYGLZOLdlu9rJEzpCqXd7HdG
z0yYA0j/CK4Zq7wy1NVEigK5kXsjL/SrTWngj0PLHO/zCnfPUmCQPld3NX1qTVYUpfPWmWRATSoH
7ySUfUWnl4cEzI0G+z4PJv2m2ztDcW0jcPZrY8gIrRqhDMYnjq9FT9qwUtjut6kPkI009k6gRygl
4Fx6zKF46o6cWJGVseOMnAoa4TcGQeGQkR41MiWT7H5gbkJkZA2JfZUb7cRAIJnVXhXZr/js1XYJ
KkhBoqhmtdxrKymLZR926izlicMBDO6e9FE4Fi3U3yeu0fEEdnHvXXb+XQegOCLprwQmljCWRpAK
BRbUwHacODl+wMzlfCziIEw6Jw6hZ40ZudwqTVpKIWxD06EDr+keaxxUqvquOkINe/7dwLm4E7jP
E7GFofBIFDabQAPHj8BqUciAJAv8MrqKxm4BOc7xCg1PI7LR9FZuBL55rKTwfja6Emvv/3Dr/cNC
s4RJQQW8PkCOV/Xa8Yu3UoCvT5DJOjZMsboY7m9xnFybtoVLBHC8pTvxKEPukzS7AtJcStGgWS1L
k6J9dkC2Dp2QY+70Yg0znTlW5VdXyhvkeEL8q+XOw7Vie/JN0gXFaUS1muSdD32nm8LfOnN5sPD4
2Y1UApj0cnBqucf3mt95GyZY9b+PtMlJL0FcMy6yCIJEMgDaAAc8BKpptXMcYSkqNfd2yuX2QHIR
p4WnJEsFz+kznp8qnF27Rhu+JfJKWtAB3YP1Gmg1pxZYeJ6BWaCWxuIct2xlp0sSYFWY4wqHb/YD
pdCfWV4zfj2huNocCbRmkQ13hhnCFnIKfurRMJO1cU6UKGWNqbMmLOtgNqQAPHd59eRQBCj8+6mR
bg+NJfP5VSLQVX5iHK0SCpg62mHJ3N1C4pyBT7YAP84UaeY1ONRpRcRp19lu+ia9m12bjTqDdDFf
miK+NkKy+sv03By6PWa+kY0wsPuX/1XTd5URRhQN/L65PFG182dSZG5Y/SazrQ5N5pYEmMlfDJzH
CI533Y5XdSZRjJd0y7Fh+PExpVydQiXCM1uDAZZmiyihx37c2t+EDnKNbJAX/tmedv6RTGlMKKDo
ReTy0xPL5gtdOeuSHgxM4ZmgcmcDC7UlWelDt+XeAml1uUiyw9O26VKDbANcb2dKUBZXduXYgzcE
LngvX7vvT9hu+mTKpio9c/rKpCjeyuJLpOdxPzXlKhVIkjp4hOopnm5QeyRwYZYBJLE5uHIufpBd
x0SroVAe6gd1ryMxphvHoUpzR5mzGqMF4u1ObA9rIpxOftOCWa2U1f18gVQ4VZ/e4PntMx0EfK8x
v0oabtCNseR3n2GHk7opzqahWBCs8SZkB90KBE7M1yy4NeJ+dUG4+7wXCICQGYi7zfKE2OswnhKF
Kd5uiwnYpYqjRRGrHgK75au7SmfDNTmw+UQynOA+9BXybe+fIR1TpJKPzZlHXdU5wKuTiXbnV79v
Uc7XqithnBk0ZPORr3lhmqUtWxnICOEnKJud3i6C8tRSYoJzSwD860v7zWQcQbF+yWvNDIhnI419
nuvJ21dNvf0XrTvAzkfzadhOQfIymb9jvtEvmICZtFf0nlPPDl2uCAkeIdm9KMvAPev6y60gy0Sm
Y1uKum/epVZPDkj8XpFmGEyz+9NwzTcu+EyBUEc3zCa4TRESWwis8enJgqjblqw/ombTpuxk7bAK
E3iirXrVh1e0fwrq642r0B1YwT/Q/9Ym9Xh5osYSFzeueVyiwJaZgVhJQHLV3LvTs2KCG2ot5NXP
KOBFqKF0+ltPt+8NndQS99SKXKLs1D4KHxxvGlEcDglwUIr67OO447LUwCRrWlHvoUq3fgn9jNCK
Yb2A+twDJqUHx85uZH9scCSR3g0yvcaKYmgY3MXyUYSxf8jmD9urVKhT6Y5xQHe4WWnV/cEyJ6dd
8ylCW9XM1NOBMlNlrF230i0vASbY2/pY9gMZbjnjpAwddodnQTMOUTWdzIBC5QdQ/JL57D4Ou/cu
12yWMta9Fj/nKwdqQQ0oRZWoBI7OeXKhNN5DiT7ZajweSgKekH5Vv2qLtdfV3WTCmqs+pNu7yDBQ
zikhLtez/tKsa3Ddapu5hOi7vH7Jc16xIbFaDlGmq9dKgvHhhQBE7GLs1qVoBqgiA3qVXmamZZDU
otRcgu7rD0/A5jFnnzR6HogfBd9qTUhFZPTxAPsqd1cNwpl7YeAoo4CCvVDlIaqdnWz2x7EGMC8V
ukOJw+YydvlQBb8Tk8bsIDOQeHClKm4A6dNVOA3MeLVKnRwErbkvUkaze/wZCZJH5hFgtkiB5qL4
+Zdh2b7LTwEXdhrWDbN1KoplafodpOnKRw0dtyLiQeS9HNHzyN8YJHK1eFD2gArHdm8ksYTn0BJ6
Vg15NmdKdKdc60eovCF9vu47S03DSFBFI1KO6lMDxEhEPSf94ok7T5c8oLvkZgr1j5HdaKHdvCH4
7qiy9ECYP167rtTMdginUIKZWD5tjp+S+y6gO0+HWJXHs2PMMJaNrj1BVayJ6mnuSU/KcOnwLaK8
7H75q9KZ/Pr8G4PLoXm23cV6tqfzc96jjjIejOYEjqZYlaPMXYbOPySVl6+MoNLIFGol5DcunQ0o
Bmr1aEj1nh3cqdzQVaS0G97TVwR8nkDvKmWqLM+q4c/0y22frATswAJDss3x9/ciNuEKwWoVdl6L
0dNtvj0TCRLkGE5TEKP2VSuTs+3J6K3N94siZvsK+cs+JdsN8TDJMKkefJFC7vHNXSkFF3kMw4SO
3R0zBwvLYGNGVp7N5/YGC+InkF0FpXREgEXBXAgEa17K20pCc/2aoTH1fLckamOMg4pPRdLmd4oA
UVWst7Xbk4Rggl2Q/4oz2nXPiiX5OpK0T//0WunCmNCluWwfoWT8AvyjsGZ9MYy+Xn+0EoFlIqUB
b6fcTVZB0zz3AMke877/nkSYqoXt7NSg5ZaswBeYVhLEiF1CXz5vIYpYXjaWHFtf0eZh2GaccQxt
3OJMBAo36ccLUzTW3Ris8gTMXaOelYben7SpXQPh/VJ2J6SjFRbQq9qENx1A6YU0UuvQSWKjvi9x
wi1jdcTTcNIDBHhHpjEmTL11HogDeCk+G7BiLZL7mkyiinkfv5XQgqi5j8BzQIBK81nNapNxRJwb
ozxTjDBf9XBjRqgQ54RSPct96g8iWjXOTLJDm7Plz0PA2FZbLgHemr5c0q3+6bQ4snYw98QiKSnO
syG8PwX5D1CedmMvBsF+FhIoo6PSeG4vrvT3H59hB/ENayMrbcLJNjIVEna/kLkS2WOXPdRwXu23
mkOJA3lk6bK3PBIhDX8G/6fdSKDpinlfstNcUH3D3LnILUx/6TjUKyF+Do/JxsKaU69ZLnJiBwId
Tm/OuyuC/potg7BoVku4i8EgwokdL0MlN7dYCQQut3rTnk+rlx1fRKscS9jC+CDGU03CNIUUCarm
yspFotp7msnwl/D/Is2Hi6H2wZ1nILDM6fUkwjwEmoGEcM0tIZqq+5LXi9EAYm6qb6Gq7Emqcyuj
FTdR5aeaYWRillpOcEnMpZSEPsT6Ig7EzSP0BZzwxTvFpZB+TXBEM549fstOb8/ysh6rbguRS7Jc
ILHr4R6cY8Ec1Jz03Rg8JqSJ5m/wKjitwd4/Bo8cozv9k+a6ZvsrrUKfrOSHPDKz9NHZlJ+Fa2KJ
QAOlv8hQDmwmJDpv9w/vzC5fUT3cPAwzvVCwGsT1vXaQVvvge5KWRKAfeZE2yBhxlpQKRwupeddX
Rn+hpzq7sPRzSmAQ7hDAUfZd+1GoC2hSTW0KBmCwO0mykS1uV8JyQkPSoojbnd4Z0Ybxs7IfblzV
X5FSDT+5WR9WHsHcbEqiMn7oROlsRc8Nn6c2xVyX0FyAsf47FRK9vvhbk8XSID590eJOtn3f2Z/N
3x1CPHKkFszwnfHDJGKO9O3EwGQCJDItLM3Tjk8SmQnQmdXQWxaQc8U2DvM/g+ibDn3u7VqHD/f7
fG7HViKdY7lR3yfL6oPKuYQOcG/fqHHyqJK3nYKo6D7OtJ23ILTmC8tYUCfSoG/DxaHiszmKyQbQ
6Rs0fzcodzGv0beC//dkfsaGPCaaR4dPj8k7MAdDIK894OSPQ03XTcXJv2LRPHkgjpds4aMtpuCP
eZOYb5QGRR7xdcDEXAHxgywohHZXvhA83QVsKy0FhjTxvolur3FsYOOE1eAjAXQCR6AYiSh8M9u6
VNYGYzdI4nugBtKOpZtCKb3XK2ob7qS3pu0ejGD0TqUca8BzTMtXvacSQ/FqqTjF0A70C+A7uD5E
zIluPt08FIbnh/ai5nWyAFtk4qYGJEyp6LgOCNy/88Eh8woQftv9XsK0tAf41dSUl46hZz7BuzXU
K3tvHYL3nFW+jkDiC7CxLSgjPrvvAsWNftq2WXi89TwE9amugHBWskmeS+ncKNOIkzKXqD+cdhl9
US47LTk+pdDUbD5beLKOmdWWmEBsS14cbY2f0v4xEI4D5w2yECNuCvw8lwvL4umCrmNXO25y8GKE
MaEmLiPrC+P8QAjc2re9Ir5xKyDj3JCO7X+rhwUyjWveukyJL3sZmpoQUWlJ2rN03GwBAuM1hTla
C7CrndudgOMHPDIPezwCnmvsoBRwDctwcDKaxv89HzilAGWiITiYE+xaTYh8mpZDip3AFRo7QEfL
KWCVLHz6zxkMPo9/VkarHQxecvjA8AYkQ/1uW8665ALdeqUyqtKPJUywlW2/JDDrRpkbTq+2rcfm
IoHcr6iam46V1QJ5yge+tkHx8+JsO9YX2xSxl54jQIFHirV0Ucxk8D4fNgRj9qB4Q4CFRGOd3sjH
qq/z3rnHW02qGSmpuV7Zk/p2JWxc3JyGEyqzK4ZTOVFNFfIa+7300x5W0EwQEg7sT8qtBuTSlMJX
QEvwol5SkkLWdEzCL46o8EHDJJEQLEuDhbimwn7VazoSYkuFXErn73IQiGLAgf31qUH5dJ5ZciS9
/qYcKd/GYeuNP+LqCDj3fSXaXJFBZkbMu46sIZRYaRL4EkUXEzfNqxK2KZM6047h1EOWtU0F2K8I
fFMKgLxuYEFNKPZr5Enmd77VZuS8sQiCOveQ5t4LDpJwNZPwuYbyXQAyHnEWOKsTqsyZz+7miQjh
4hobL7V59psSOY80LhEVZ0cEan8MU/l6hNVOpNLpOLPaNonwMngRkxe2+lk7l6WXmhHE0Ob7Zmxs
WuDJpcWwHPXNt1hM5nlgjVGpGjURYQ5wTP03eo64wl0RoLMnVg2HgXl+8buCxY+JOnUk5RkEYajG
lz4sIzYf/ndBVOrWNytUV+UC3wiFmrxzUxLdOG3xeACrNlvx9Z0TXmZ6u41wHZNG+OlM6JeLdU1J
DIf1Wksz1DW/V6H0ceTBTAKL7VLkr0kbFBBVlX7pHP6/uLCqGzVxSpBEEio+5kUIM6+QGcjh6HJu
R5X9mljnHafeaOD0bbDxiZ2xVdBLDWsxnShhej6o0UZiL7EO7grDIdbEE41rfs2dauWQYFp/C3/O
F/9wAhWtozTpm+Xk9TYOIdCbk3QNlO5lcHWoHNc37dpjoYN7SQybABWyBI8UitQFRY8IfZOBzoeg
c0WeWQPGPlF3VL6LkrLXmceB8RVmv4jc1Nu9E1/m/LtTT3ND1ZOQuJv/Ab1FcYe3oaUyWRRp9JvA
TmNkP+sfQURWtciFI6MApRl1WdD0P9WW1jD5Uw19SXCtcqlKe6htehNxNuvICppFAkNgVyfjkSEh
68RvcIWZr0YoP0OGcZuVlF7F/L0bFGnedoIMRTpjQayx7nlSayQC8InDKP6pHJgvVPQ5YlZtlTzf
z66T7loBVMwEW/mmVNDgkDCemPl7wIws6rF+XJHycFflmCPmNLDQc/WLoRjWl99pbrpl4m4g04fI
/aJC1rYh3JBH7cY6UBliCMyJ1JveL3kIWfcmafhSzUGddVzKIvBkwGzsilRqHvGFNl3vZHg8Zmw/
88y+nfWWpOA/sqzejiBfVEmbpz8Pn5/sasC2xSTW/9r75Q067MUjwnFCcuSLNe1/IlaQs2w5iJlP
4snNMEhbEkv1D48czFBVfni/hDPw3W2k16q06dkL864YhDua3K/u3ajNmiQRG5AVMy7uzcFEFgxs
Yr5a3wczAYL6ik4yBgz+hyB88yRFvyMUvT8W88Yi1MITYhdwBBQs5ptzEMynK71prbIbDNJ1hrEs
4vf/VsWqjKV2LeuDeQRmE+5YXHC8ayGWHJkqwKHJGWOPJ+Nd3mK/LJDhz28RJpfU+K0VPlTd/xQO
4EUTk9QeRrmDxTYt1zJqKhREWdfB1w2cGx+eLWhBNvWtNZb21SdNChFewcl7PCiosKyKl3ps0kho
T8x9NtP+2zCCITXJPyDotcULHfHmjR8EUAxBvLVRMRSAv+kbzO3zzKuzusis4Gi9LSrfM1P+GaIY
VQg5C9C1JP+jRl6ik3XF63CkGaRvq+2HHDC18HziLYT+GGGU9ol/EXHxlpN2i66+qGzpIwHyis7E
9qPCuFR9CA53UHf3HjELGblZWw7ZC7CUwHItgnzgMhAOKj9bHm4dC7D9YsNCzU6zROLexp3zGs7/
krXsczgCXp+W6axwzKlDiD1ziuNCHTOt2+fSr9YMi9+yzdv5TqeurePKcxoaEAiilQwvmXEyNGhH
2fFdPR0r4aFqXGZ65uLnE8bYokIquhB2dnPqF8bzJI3FECYmEYh4n4VcTzOZRv5l2G0viXbstYLA
Sqr15u8hytnfo6iUNc6ZlW55fFPQu28IfbiT9IdzfLxeNbTBnuWt6Kk16yhpyFpiEQMl8CgyqGod
+dQ5KUfm4vCD24DzjpfGRrxj/s9/xewd5MKm9clVFDy2ZZXaC2qzBKl1I4FFv//4wb/LN6nDqrGw
5rdVpTo0AEWxbhNnvJUDNN+qYPhumljUggyfsIQ6kY0RTeQ+xWQOgF/pgOdLPKAHcAqAO25aqPOt
6cIUJ8Skh7F0T9evWdlGqxa3tTh9z+lz4Wmmj2/OmBxyIzAsCwKSF9XpijBqbHsuqXxsvsM91va1
TGkRoZPFyycdAt5uspT+MXVZZ6qrn8fvSF0LQaCQ6nJ3RNASN++t38wluPPM11w0Bj2ACGJhrRTS
KYzgC0my+Vq1vQ0XHKoc1G0cBpTqQa6AI3G7ROOF4bzy4w6Jj7k2QhIY9FuRYSJQDXeDq7yB67uq
nMYSdMNI2px5K6t/ns+gfLS5v1EVtRkzBkIALpdtdxdMP4mm88MUEgjF/mXdGNkNWblNGLq5l4hU
GIBcczbw/UYL07uKFuxU63PN/ORQySUDAapC6MzLLyhHYaTbuk5r1oHml/Tq3bAdHF4VXd3JX+bx
ygEIwd5artP7sKgTPzhR9eOxiK9YYsVxz1s19BY1QwOs5+9nKVEWPqozcxYD35EANIaP3vOIWo1F
r+VRBGUetDggjKVDVM1tZJUCTGUoWZec1JvIFSOyfri/q8/4t84XACde1bn/yZTwpDf5ZpCIMRs/
PuMv5a3hdPgfYBPdplIQCZuUnBS+uJWvlYEKEtM0AdF+RQK0BTIMOPiQuOZLPx72Pjs4x0dLfDdP
ADEfPlmq0e+FmJxiaL1ix/EbZf6720j+sbXWqq1ZkHCfgtOXt/UosMX9HwJ7SD5lD6YV891JEbSm
aDqsWbeRTJGdsoxdvPBM7/pkUwUDIh7qwWo9T4XxY0APpn8Lh2S250zOALQbQR9JfBVN3w6Red+O
6nn0gsNO3GDr9t4s9Ng6mX/uvhz6GseHWbndIIEmVyj2Xv/8ZTh4pcbZyXqvgYPUqUWqRQNrErzV
YjIjJG9s5FI5lm0hXx6aMWtC+/9B+H6MyW5Beh/NjbbMR2Xd1WdQoDj+IHDFNHO9IeiLrimbAW7C
JqaIaQxzidaUvVilL0Sx3sO7d2ya1ZgIyN3wXIixBllHbId5vR3cuLHW445LXv6zw2op8OgRZApL
rW4wfWdAfLQmwD9pvDiTCH1o1hpYO+yBczK+c6713wnNWp+jClGZO68iXmUBTYWMt6WrS0l2HrUL
U9zxPAKfnHB2d0D5eu+q3etcltE3BfDxPNykrFYpuxcroCmkDspu6MKvzP/gvyca//EfRgJL/gy/
MTBUHPf5GdxZ0LSypWuDFH+WlVnGucfDJn3VfLiiNok4IrxfNNjkYUdVhegrqdgLYQjt2D61SL1Q
4Y4m1zKfQ0uhLiE87IS+gx6aPtZfy20Yq1SUt0VWVKFlxCVZV94Vt7YKGJIeiEKQgVmdBFnahqHw
/ItdZbgDZwVj08JNaTdUNkYKQLTllN8LeCGMX8jjeLH1NrmT4qHzbN7hwiAImLcbXNT8IsfvG4oF
vOqyOKdkl6oMD2NDkfOZdMbuULup7V75OJTgT7SPyXtSq/a3EfZhNOyt871UPtDrFkSZWkFfLsJH
YB+JqrenoVZBjYSUXoznVFP/qZnO5CdhxeTFPpTVV6E75hYO70cxe+cXnqnHFocG8vIjMS++8ut1
LUmCnOBnWXVL0+Fuxh54j9WnZU2ujRNeU2hJ30xrNuP6FNCwsGhwDt8szHQjzSZdRsvXAAR5UPWr
NH7bFfjHcFsEUKpW/z/z6vAyDcUDStuwM5l2e9hHUS6GWzu8615yf+0lkYbv5CW0Obk2rvamTuL3
q01sym6VvHVDWlKHjMXmchZoQsKbrCHzHuKzsMUD0s/FzUcI9cCGAuWmJvPzUVSXMFLt+J0msqGD
vz69WrjuY8vWEbI3R8AXTgGU35RQyn3e9qud2uYuLOSUPLGRFZDM7KCIjxLn+PrrXD69Jlxvg/6Z
XqUiSuxy7BW0C2nYhvMWjja4YqMknyM5eFkTpw95tWoQGN0DXzzTNv0srga1sO7EVw1RjAuUN8Pi
/r971ksapSY3b2/aAOUVsLyn3VKqyTEo4kezdpzRI0xTsvan0scPnT5tHaZXiXcrTlBpYUAhHHo7
7b5ESGzK/SsKjrrn2OLvOW7RXD3IZOSW3lHPt+qgSeqH/pMhwUFjTH5O97shfYLh4Fgvg/6MvWf1
/KWXayqQg/7Xgj9SfIOxM/QyxTQS1ZjREjYayVg7NUCrg+USKVHCNWejy++kkUwlmRdrZvt1n8Gz
hcn0LE1cayopwm3HEAmDwFGmAHt7pev7L0LWlOUyAM89qSt+hVVQHGZtSTmXEvXlhzJiks51uUQi
6HHXxZvRIDz95anjvbGyUUPY3cOMBtfmEsuMqjQfKFES75GpYXFO89ohxxZh0K/80TYqyFoGna1O
YY5R9iCBjhfgkyFKbNw4E2AEUd/k9bwRtI0AWd0/OEuQEjahfd8VyeZbC8hEtcWJRGKkfZLnSMhG
K2LQGCD36A82rycozqu0WrgL/hamASzioRSGM5DdDlcqouSfVBzUuf6vWgr3umJo16Dx0hsDvyuv
FMlG8lfGHWXA003mE1JUtaRB6jKc69ZJ0zpHmrV+0xPICKbg0EU3jH41tghtKnIQHk3C4iDLnwqk
hX4M07Xl/MEOsG6mem1bhaKQeee2amqcAKg3JGX17udEqoa6oEvd1Wo0esm++wHI3qUfjIMfAzs6
dqnq2hgm9OUEX4eA9YVsx7uaJldHM/ZTUNB2DCx2A7rAcZu7oN8t5Lyt+69PYse5Pc1BoYi3E9SP
qpnbf9sMn7sxVfxSjn/MAGqhuR9rozqv8G3tewN5XhEALg2ha79qYtxn8gua3tj/VuJcqf3gUWxl
GaACgu+tudxHmbBuVRHaRgSg5D7qBzVbT1eOBnuuMo3owQKUyHOFwDo1ziSgCi/zfM4poBn5brM5
s78kDXtdgdTxenhywoParSE/Sny257JyVMhUWSS8QdRFH1NqdS40dpML0Ob13VcSjN4Qi5OYx1WT
37weAoREdD2mBlQHxW8j1e7rTvnc3MhihRLYDEdfJBA9iZBtb4QVQ8OInpbNwf9bYl70Ia+qwMQU
tX9gXhT9zremix2akfiMSiqG355R0fkTr69lptUr/y9uue2Q/V/uQ3WzFIYUqzNrLwnTZh4AatM+
wmDWHp+OhZWzAuX/bnJIWAPRVJDmOh432Zq5e8zyg7f+Qh2JDchf8VefKNBVrTxkDe3ktn89WedL
/56l2y8F0y36I4Eizd3zK/99AKTopEvvi/3ccW46lUuoFyFnGBBz/Zth9xbW0Cv/qMEtWsF5amw/
yENazwD/bZhgw8+AHVL5uMvkF0uxR+THYUQfMN9n64eKezrdqFTpzj8gNBRPn2N+gh9XT5DyHLpZ
ru6r1/RdQohmUcTV1YcCcqZ/5xrs7bV6/V5qYC/IiYaIk5VMJhyF6KoPxYdaje9VdMk9Gxt7hAqo
TmcPayWHvkEsnPOnxDfnxuPGjbOUOOtrDukJgLet4Y3ahMZWXSmcs8SyICqJlz4cg4L2LS3GOTOb
G2ULyZRUjM2O/BCUF7jxBKQoEgdCXwJHobq929Dum8JBuM3qBnEPa8z27u5vjDNXJZ4UIceTODZO
GuWhIIia0UIQK4dWw/2WBHwn64tuxBBWbGyoya4zBuOcwzf/f79AOIjRYK9C3hZaxD5uL0H1C0Yi
Mq3uz4FdrtLKNnR9YyhSu7lLXet+MU+o6EE45lbr07cFaX5DJMiBchTZFmURhBVyjp7O699LXw7W
+pjrmIeBWncorC/CPUxY96ASlnDP2KSF/oXOIQuWEzPZGfPEz0B26vXLg6TdSkx7oXDvydT3lFwb
3WI78YZ21Bv+n/aRqjHbPtAZAR0IUOF1BeE6svurRd5IgKI1Y9XxvQtWQQL4r1RNQpG/+fvKP9Ii
2wUOGADQTFJx3wkHhc73gcX65uGp3nsgv4hRiBuOCYFgohZKTm5P8RLKZbFUlzpcleXZ1cFq22t5
BFERySlp85JbzAEUNOd58XXVGcI7VjK7IhtUCg9e8k0eBffPPWf6YpO9U7dI36dRN6fcp2gRTznG
IQVDVO1de0Oi2k/ZK0OSlEICuBoHGpw8wwiKG9g0H+zFjMhgTGasRp2Fd6kuVWTRR7VkK98h+n9X
Tuzu8MINWXXo4J+7MSSWcTJWl4/FVn/hZHrOxIw2OQ9eawsj/TtbSA3hsmKgHKYXYJu4jIyLAzUK
Qcz1J4fkbu8BTnfH557HgIrXN+m+TJWuE/iF8LI77PkC3wc3c9UzIF57G/9e8DDzbn2fjCof4lO+
xzJBYRu66mq6J0NvJMzJ6ayzW79ENDSfuSK/l55Mtyz9G1vHYiLMnDWvbJrTICOR4AB9tF0Xlals
ZdwNwiR2uRpul38mNuiBBAFkPfhWpQdENKIHLzYps8EDxWd1kMr32NvejogXApe5qYsvuXuS4vfo
xUghdKZLGenad3r8uoJTz7vXwpOGC8ufeKncpIVvSLQNe91PpCwx0Xlcgv2zV8GcZ++QisRFq4Ag
tEzXqsw3S2HxaVlG+rDZ40sQ+QAD/EUGR3g83Du6EcMpamVDjVfSZwi6YQ2+uWPoPx3t5vW7Croj
9SXHg1I8XyJT6v+OILd64tONVlCAZffFePnQLzeefMRx7IX93u05GmAoi1aeM0cP/CSUOM8JeFXJ
kj9BIUdzSFCD6mqurDnhBMnXYStvX5tg02OHca/m/6+nOZTfEMxnq5fO77YdeQ4A41lBrCFu6z1R
UrkPJ8EVNdYtmyes+Ee5bGYs5IJxwcwB6cEXgWjv222UPXCr876gs0sVscYILhw4GIlLIYbyS9kN
QpHHcjBzYuHPWEmBqqufBLQ8MrSrWwRtUuc8g+5K+2th2blcYQgrhu/vrdyC27qb56rJ0d5tSKvh
MiZHyeQ/3BguoAgylLH0jnN5AFj19C5vVZXtTIyfYbK/dEmYpFCAOphpBGTwZvTLMjDeZjSGCdry
Gzi5mlfrjMPkjwxLbDUNKhDU+VTuZX5ui/R9dVpLPO+IbJfTE0utFqJIJ5HIQehgpYxUIZBTkRhL
3NtfVkI1ognW43p8wmFuvX8KvvzTyVePUEtv2vRQ29v6FU7vCdapm/bNKqTNg1t59dA+jcwr8cbG
6u8/oeUs9irMRbYR97ChYlPeVtjmqDPX6SgR468t5YiikZ5OVvHAjuYuz7tyFKNVlRY92wt/J8yi
crVUwH8I0ZEtDV+UyjEEqr/Z06kgIqMMMbHP2IEv1nvW04JXD6W0v45MpchkcFxSu7KF59xFqfFM
dtFx04rAcjGZlM6MFGOecvGyzMtklzhd1eshQ/YeGjWMrQeKYaoi5d1XWiFpv9wj01Ey8jG6/X+O
d1HINoWAJRGrrmnFip4UIE/G6CVXXOtTAiYnTo/eXPT5QpDEiiafnBD3v5csLf7DUNGDgOEM99gf
+n9eJbVi6Vk0u4B1IhOLR0u+uJZRrrsOaFAcjLu3tLAJ4hAP/x/yeLRmY2gf6dwnUjmJ1yUmuhne
EraNFWeaK3toCprR/ONA5PS/MwKUxEGRBgR44JWvbCfIr0vsGgganu2zHqLBvkAw6uBTTW7NErQg
XDV+VDXS9oji4nGPi0vCbJh8abOoAW6vJt3yitSZSZu/ZqrNS9z32uDu6GZF2+jC6yq9k6xRcLXN
Z6n2NUngRnwdMWFBD8FpxrhMl9X/kzZXtzZxCWEqLLrD73npdstRdS8H4OmNvpFcFRbEi/csoV2i
/VPSzBOf11KJ+O3SaCK44oNDiybxR302P9WT6iroWGs1wz2sHqcAiEWSBZiCggVjde0/+cm6TZFO
/DdSaVNkJq8DD7Z1SXorqFavW9pQSjUr+9C0FDpzQFFnGKALFINSr3YKEuc93xxxErNV7L16bCaB
Il8cBnpObM4npezVtC1+F0IrEsYp3ynGzwNWNItDNgYPZdyr8ipsNsThswaWwHxLWi5LP8rsE/LB
Dky4tSqHXmnoXQ449ylKQNjbzWLaurI2koz1KpR/1osrwmbGNduzGQ3UXKtKwMuQEJfDK353TcU4
r8AAOJxIHOR8y/mBsu/pK1ThpKCR0kyjzpivM7DPhdMpEEWnPQbULj2F6efS5tt+Na4HYyMBk/nq
zbj/5SDbIK/x7xQKXdKG75M47WCb7Cr4eEJPQOVzRyIo17kzJoa8L0q/WqC1FoZ1BHhy6X6XHdol
rfL+lHaWFBP4f9ljbbPTy/IjDT32RD3d0Zha4MdHZvI872wYUgS2cPnjJwsaA7k1C5HPmCJqN4uY
7eT6UetsvXb6we7Bcqep/dCmRk8haMbXvctbUrahUFvaRjt/1HDAUPhYlmBsRsRE2apIfGlAcblK
tAEg2CnhALOZ+lpVF284HXgq+M2kymNVMje7QWnURGv7BcIfmytWbAIMleB4v35EpGLzYmSVyH8V
VfFfop8nBicuCl9pCJ8S82HUZGvtijCYFFp99ettUAFkLoMyJB35pQX5TY/d12qdyPKX/kw5yN4r
nWPZotPLt8wnkjdu+/8jZWs1vcpTGZRa/a0L8n1wD8IXxbO0u8aVkISBqRpN7mpp+QJpl7ptLTI2
gVgK8u4jRnDu2G1zm/7bD4mhcDGrEXBMHUQ09PivuIeRjbH6m0BXOkwV2K8MtPNibmHlxcvsZ01O
+S5B22hA14mlpwYiE/FpskkAODUVNDoc8y388rIS8d0sRpERcaQ9oZ+h7xXPaFWBxzai5mfN+7Kj
SP4yU2xW7dNkCVtny97f4vPxTweWNZuM4W2b9li43DzoDICPCa5edxU5jzYjbbSlWJmL0s066Ayp
n4tcSQAlCsFfaU814+53smgXDWAhdIh9nzqLNUItSBVAeZ5WDmeuwiPkIJHC2R4Pcweo8YpDYWA5
Ckd4olixZUUgf33D5k/FO10M+j/1b9Xjm73X5VZx7IdTnsJewB2PL2S2lNuuaBCoexDHAbVSgRKp
GpuX0NUQzENPz140aX66AFWlCLjiTndkQwJfeAHTxei9msWdoB7i0YNtrIgJGeAHH/3Qw8aJS0MK
93FQejnXiLDgX0zvwhfRWaD+KK1c1nP9chUoMERwPaTWXLH7UQanl8J2kyBcg93hope3nDXgJ5dC
yiBKJz4VE+v2+7Qzh67exRbSKLiUmXGVOH1QMuhV7Hy6QPcBU5eMUXCm+aqe/63C9ro6n5yJEIkF
EBeYjeQvhT+uInN6MGnsANd3rhoF+2MPYJ5wqvPlulEG3UKtORdokKwxUHKgDjG8WGAIL176QjZs
w0XMbr0IyvqC/BA/IuHlaK738s+HgcTYNXhuVlj+RjzdPPS1wcZS6dODl7+qm/OwKnyOIA+VMYXn
F48u5+70ZzUs1W+5LDHrIlXPY+Ik6co+v6e3YJL02gr9Jj3+YHyg8YBGa6yOdu8r3VJ27G/ecO9c
PqjGLkMIDP51qw8zYsi1CPf+Y6zU4ERX5w0ZYqAWxUyTRmoYh0YioMgY5DHZWtTkHDqczittPNdQ
c8g0gvqd44n+Cm7BSGck6aYIlk887FZaFfYUHu0tZxSh+Koe3S/ErD+eubVN0JmzyQ6BrxmN1l0e
RHyF+ebcu7eyUQl69/jUJ/Mx9+d+e7HMO7LKkRgNkCjN4dqYNL0hntoN0KhVVGcsdIEl82O18MY7
fZJ1Y5BFenly7rmwbfeNu7GwE8qRFvVT78fGEXWAdC/rVm3Sajc27qKh9p5WBemTMPllQpEV/wpd
FlmVIZNV3QUcZAoALYk1e9XzBw+VWVVxSjAtiXVMMdhSLbGsuuWJGkCaCTA0CxUlU3aKgs212jI9
hF0nXdTI1AOIDC8uyzs3ikLfFb9whitW4dt8kXwv2rjQqvaFIGT4hElhv650H3+zHE03V6optn46
ih5YxJCaEkNnToBlwjAAn7oG7HpnrdRI6t9avszX0BuANCLenSccfp8+hkgiXRWXEy1YVQxA2sMp
uiSPKOYcqDxlDe36bb4d7fJQ1YgVu+SK0K43BECAqi3fHoizLI+Hy3SWsAu/tqsEiKoytQUipygX
bUr5dHh0KqKfKuT4MqZunV23wIfJzeNWuR8AdiJrIbxvLOFGe+39qh0F7+yRFh6vkn891nka1V5E
VpGc4VvKqLguhR+WgIyCJTKe+dXul8+7FDuglpo0UTslPrp0Y5UYZyYUZKrzvi06ADCUaxzkdZ55
ANCFDzOlcdisvgbflaJi/jkuFOUlpg14NwkvJKPGYPRklpnPdjt8oIYG09AXkH3+EQ+K+UYQrv9B
/Hkp3oQybJ00U6RmtHsoizGng7NRGt1zGekxGH+uJRXQBZMsiW8P5DKTVKplqnGLHSSdffwNBgky
6HHrUU/GLzgb6YQV1XzAxpT2P/7DL1itmN60ESCGkuuwg/3CTzaPKMtr1ttP9BEg8oxfQLCIyfIo
W9a/RC4LvYCxsJZo90FtIUnFdlMlpKfYqP4VYL6wI+W++iuvS9flBkk45gzn1G+XniHJo5cS0dZI
Nr85/CG9NRK+v7AtpW73Us3+Xs5QTiEB/H+s/1VXqqzUh0bRWOLcl1b7qd4YkuA9mQnKY3MnLp9M
GOg6lI53tPyxJ5sXqv6Pi2zlcWyR7Ar+14y2dVZFBE3tP9r05z85LR7ZAca7Dr06WwteMHofPs4Z
mutz55pe18PzTEg5OR7gKw0v2zwDrlnVgucLjmUAedkqwGSydwXqXTYgZn1+Ar/wiBaXYpCQpR2p
c9OuZ5dURAOFRs5TOkcVjIJN4YhKhx0BkqXJxDkhZ6sNk1xBbBffJ07vXLzE+tUS4eDk4e3TpKFB
zpaA1DyYHRn+W4fqSag4ekhN+MVE5UHKWLHMA4QOWPxw+gIvWmHRzcHgIlkxw3KSA/II1vnhvlh9
DSLuwWcqrp2ABITNxqei7Eez8vNNEWfT33C9fOe2eH3ur6al2e4QBfAeEzMBdrtGC0g5rBjng9Nu
ScVells9RgC9RFTHWiDpkg25fmCAet3NkmIMTt3hlz6E0AY+QHtI9hkl78Df0r2bpPLIv8ORK6IA
IPfcPAh60ytN15euBzro8/4O/4WuOjEOoy2I6h27CeOdY4CL9G4e+4y1eLCO1u4qp7NfeMmY+Jvz
7D5DKJkFlhwqMK/a+UhVKG4T0ujPrf60BN10kx4607pEAqJNkRrtD9xrxGbFmN/3KdT8JesGmryH
pG7m2H3e7XulNHju3f+k525EvGuj9qFNbTY1ZnqsXOD4/wue+aIp2v0aoZpaUOzrT7ouRHnykOos
vAEYqHd3M9MyKSrCJyXS6mdf91XJKRqqlz+KD1Ka2HU6S4Crt2nPa6+I1Y3TAaBVW1u3orykPZGa
sFaLsTtcRp1alAsNRQ1rg27o/tc3tVYxm2ESpoft8LazNAGRkRQy+ufgsnmg8we/U4pLXSKvojvh
F5r4mFGLggQ1gFrlX5EV1XrA8NKdniSaVHJEunzJgx4tlA/IOwQW+UvU0rjVwgqADbRbU3aWCVOt
6u29ZT+obkYOt5DntT0ldYSOiUa7abokdsPa8R6CZFz9Hn/ArP2uIXwTxNKM1XIymycFtsBrvvqU
yfD+5fjKtIwfGXFYQjcJwVBbjMIw0o5kmy+4hpxhf33GoZvEcvSpcc1k7max0YN0CH3qYdGiOCZ2
vLM6aIP8CEycTB57rIMumQNkXY9GKCBP2PAklxCw3IQ+Eer9GMpSmD6xxyMzm9d9egyQMNlUTuzz
F1XF4+VUgbkcWgB7cnTgGcjs8IU7RwdcGdyeIMcz5rqDZp0NJmSg665cU14bzDfpGm5Z6JyYHTZc
D1nz1BuxfdNdFQv7v5O0d2E2CkFvSPyEiJncTZwireSMmnovjfuh+vw/PUvlIkig9glw3e7qQt2s
07mM/pKGvYqWTfJuU10L9JG9u4Py4gZOvBgCACbK5ONXB4L/GsXDomJ6BJVKOI/DyG7HBJCsjXCm
iW5brbQH0Twgc4Kp/Ew/wOnWzsZgE4HexJrpOSXaOzXtlDMSstJe1g0yPOKWrfm/uFnsPraB3oIa
tp5Y/ckgs0q5loJoS8mt1621wOa0jIyLV3uHLdgwXTdVtobqY7slTuZ52XznutLxMQNbxrB/KDRa
lZvnThdpSFDbPPh0+7agcvka3uSVaEXp3fp72zvy2zVneKqvW4UEZI02a9fdwOU27bO3G1CSoUOW
LnHFBCsjhhffLOZ6SpoA8yk9la+yLXUsOmDbnXG4lqjtoYwTYBwOgoNL1eMpXg+Sd5d43LlBSOt6
WLdU3JNHhyAw8yajrmUEK5PFdA4rSSGmRzWygEQr2RS8Fe7AxhLjpzpFIJXrPGHDnGLRFnrJRJaT
TNnOuKyTQdvRispzMBJZ/ipAXHTR1N1nXfEKok2JWcG349mSSXi74JqUSQl1K4ATGwQSq3KkTXIK
jbu0iHvbU6CxrIkbMfSMtm2+kULoabIFXBVjNb2lsfIRYWXCeLL8YsVCIlEFRhTEezwwWjmKcKZ+
CsqKLWd2hM50r5VOEdITfvedcopt7p7lOZwNZOGPK3CWuUZn/OiaAVlDXEuGaZDC/OQEAyZMwUIv
W6liA/bBS3t/cR7SvcBlFbFtUzf3pZXxpHGUzC8Ug0u5atZjFirh2HXA3vZ2UUOEmxWTLPtQ2nc6
7FDyZ/zksAwvvIDVz8mWAkR+HzrAkpVYtVIHyLmaHzGBJyG//0YTtR8260cvXKskHpuT2Yhg25Aa
Fcf6Y28Ayos4D63d8802XcmwpTafcCF3ANywU68BeUivqw3tr+bTOgL4vbc+qKNZXS9K6pkOJNEL
yrkED0yXHN0TgDfwz4LMw//zVRtKAwxRGmA6BxC+RTql2ifIzgZ9a9r1Et8ud+LCeD+YN5vTTv9Y
UMSlD3VFDS4RlN0Gmq/1H8hTyu9jYfN5oFR1qmm5kAa1HYNN1llfv+ndCM3f2ceC4YZkLrA0VIAG
+ii+rH1yLMyeREn17iL4n2iKc+aUX411t9SL17ShLwZErobzjob4PwkCuRT4fu0+EQUVoI5RM4Ar
hCoouAj0AwZyuBZ7D/7T6O6Z+gUoCusBedP1q+bKS/QcA24Omn2rkCaXG1jTqivlcrB9zKotoCLl
J/xoBcBVx0TmbDRPDr94Gwl/sukOelysh2fLpOZyFrwOGaH5tnQfM/WmYu/cgnObJZIwG/HjW9Jw
oh4rzyvkwSPxvfKEc3UqrirHFQuiG7sWHvaeq6/oJ5WPq778+N/GAGKGxnnpzJbQPJviVm7N9+Ad
J72Cxr2jc/cC5Q6Zqzg8InCUOcVff+t/2jjb87pqKMoBJLLsOl1wS92Gbah/M/fFGHFjkW052fuA
1gei9Va+hYJjXD9gv0GmULFps6YHvaeph8K5Ol6PcA4Eckq5GVoDzWuZHTWDucejEIGbPZPy2ibv
/5dmrgHr4Yy2fsovapCdNIhaR4vTPLt+rGQbASY8TjLpYvVnOJ0BQ+ixTTjQrrb1PTl4O9cyFjTj
t3CCRkVThYE9QmLW5CnHqcLe12OdxhQ/GkLm5KWPdGmZarLe1i+PeVyojdqtFagfLmcExgmVbulI
ZZ0yH/k1SzJhaI573DtbzPio0H0wODxnQXaH2V82sKDBrGXsCpfSpLNt64u00uS7FB45CVfsuTaI
Uy6h++1n8fJCwlyLMrN3X8OZV7Cxnn6M+qs3Pwf6fE9hQQ7lp10epRwO3eEGWPONsGrAREG+Opeq
WAt6sw8raayYMgkF10V0u0gL0CNRBwI1y18mRR+39dbokqRSLMdxNZmDMWxxIQLC9ajQ6Lek1tRN
Hw1GIz3SYIJWPFMAjzIISza7aetHz48cGphGVdrDlV8V1+mSiah8v5aCZr3mWb4omZ6BqiB37pUn
28tj6JWLjDIoF+NTelLphmw8+wI10W+bXS1ZrtFEm9SBsxlL0eRDDoXF2ek0jvhVKLCv1q/Feq3E
JsJQqoNBTcfRwCoROYhyUYzvoar4zVKiD6NIFnzEsG1edVgPBddUdF4jxH9f+ZDOS29RyZkF92MM
3K3PZgf1nPAAqapNKEHN/7r4HokLH3bUNE4aIVDIGkQqwKmYn6KzAjq3gO3zSyW9KDjQzO6Yhtl8
3bR/nMVhzgJyCWT8Nqprg1jpDgFWDLTZpzuV6g9zw7TxvFelosGWgDjF5JTZQ5Trt2/R62cuwjKY
l5m0CmkojKOG3WHhdL4JYDXJbKI+3jI9gaaUzg/1QBa56syZM/r50k166dCMY/y5jqcK0F1J0aKI
vMmWCNrdzqhEQL8vSrYJdDqD/oJFKQ4DRK8s1lVtow6ycvZmUvw3ekO1nw73u64I8kaybNhPoygc
yMLpGwOWpfN3VsXOxAPfFQfn0g0IbmcxaRqDl20DQaaVzhuyw0pP3r/+5oiPvS/2jELnRi9pD8Ts
3kzpS+LG9xWhWnxLwNZYiE+rtlR8pUvkMvOI/ZKh2MJUbZ+8CA5pBb+zFSYf7WHt2OHVv+BfPSnJ
jpestwI5OCGj9FQKBiVETjdxaJ3i+E8L+xCTqpk0xzTzZ6+/1rro2kyKUc93VjTQ/2dPdk5MTGww
mUFEAwOAi2SBw8rmGKAA/XiesTKJ+LHcPOh5tW0Z09b2he1e8eCKNZYOHTPhahac+7OVxqvy51qf
9lc/O1mYDGaqGTBew+iZhEx5O+dY2/73gkggaKLB3TOniktb44D+l18l9Yd47o6AM9QM0RfcPoZh
My+Be3Ncp2b8gD1Pn1f1DaWezkVJZKSSqMrjTMKYd63B4epSq6O1jjCI9Jwt+DpzJ7fxw65fYzDv
Xp/FWfHKvV7UZJGpi1sqvQeTxt9WFmR/mE/WIkO/yywwoNEkeebMBu0uile21df8IEzfCCLnnJT6
JMAQRRiGNb1UBndVYZxJfO03rlnHDYAaRD0RN1GwE5A2pF17Lj9cOiCT67JAK4ovZTrZZmZdNWOF
v9LErcpMUfZxccyEcgK9e0aIH8RLvFhAEbQRmqz1cdviq/kWjz3o91iXmaO4m93KZ9EvnUzLpf6h
6vZbxsgaTKj0dW5jRni78DWiBJ+CDJjZJPYq2o6CvE4wTSTzWJBp6mXG0jipzabIeNpludhVDmpN
uX9tANmZS+1vjJLExhDgw+CJxCIiuio380ao6FowUZV8rhYFzwek+ksW72ziZFFV9M60xh8wnvbz
VssXUcCB3mJEAag6iIR05YrZnyidvml3R+GNUEQoYepipfCcX94f49ovE9lIhOi9syDT5xH20mQE
cmW97LBMDDpPFUvo7zYSFo1GnvYPcfj0BGJLrU2iQ3EmN+ip7Tkmz3P1p1pDhTTF9C/zvUb6U0iY
Wh2lPKG/+5yRp+UScntaLO6Iio84u1ZvYNe2GcieqXJt/3Ih9JEGSIFH5pOuQzpd0iX/n1SyNpJ/
MMu5bntNFKYi8QJw5O2oOenob5JZ0jLzS03ViZXSIVmgoZnVBvkcs9iXeUYbF4CTxxurecDmub2u
KxO29XtIOhXpfLtL5OuMjCB9JuWYB9cMeZxMR1oDtO4QFwXJ0gaP0cjP8P/i/ovlHt1QAi98l31L
h+aC5NNZmYMmgjAKSppcJdljj1VUtCvSx/o5+d/eL9MmvgKojkuY4tFZd+fV9+962cbGEue7PCQF
7dHWdWsN+IOKB1QJ+9U3onxFPBVQQJF6csHhhGjl3Bndn8v7DkdWmNZrjKqIq8W0UnlAvWF4a2iZ
MDl4VcYmabov9Nkkgiuo2jP5NWDOnKEuV68TVLPTw6mha1ED41HcizLAyDUAHL0oB/lc4f504PHU
AuXIhkNNqtRyWnaag7Kq0fKCppiA2UyV5CCcB77/ZLsh4L6YWv1eZj7V0aBESlfCsCPCIqGwAkex
WTKjv1mfMqCvK4Mtg7YaPxFZSPxliXwvhf6lwEuzGOxMVVRoPR/vTSJDD+k1v70KnmLA82u/xypI
vhbjkcsGA77ZgXKnK8VuWq12CoxPBVL5oKc+CgmIGkr6HeYToJxgt2+8+oyAW1RCiedkIjNr+FYO
ZBUGVIYkpQfXzRVFRPXsANOnbm9TZxipi5Oy0VQ08VJI8ROQ7nHAp6fUtYUBmMwdwz8afY5OzB1/
vwflJEbGx2MCiVrXLUycVUvY1Ga8/RxNU9qPXtry112dRRBsLxDmVmSlZLxRMRkgBgDHYV8/JvVu
HHPQhuTHSQCSKuGDEJ0ukZRtj+4jKzbG2ID8KyQ7+Gxown8J23n5rzzqZ6KNfQlE7XfV4xk/Jvr9
1WB1BebcxL8lKwnhQ84sXBVdpnRuWiaqSZfBCGW6H21ncCOZSYgmLukWNhhVaH0vEEbVSGf0chP1
Ajq3yMc1zBMkRjStc/ta7vuMvaLwNum8UTwH5Rttf4YwYMmzhzWkdE5pLddLPcz0yrL+YzU2Q0Gg
bUVWKFBR79KSEYGGP+2XIr4wHtwlULVPFNl75bWVXy3Q0L4G4BMGJ8JFJAT115N1rMauEXOLMrL7
tcAGilgOn77WuyVTWmfuHuQfpi2560/HWUlLkDIgbBJufjr33fLZ57rBdTZRCof/qtuVc1o2BCBf
up091cB8sg4OgPJjbtNIkYrWJ1ZXdrFc/r6+V6bd16OP01/vKxOX9ThF37VCFAe+bq6e90M/p+/b
fxAFFajg59Xx5BpY1dHPGIl8MPjTPrNqIf7ZP8apD5Tx9NUGQ6fhF5WC8mlTYaZEYq30JHqb8de8
0Ly3l1Tzk7ddyXtE39388w1JqgNMKTwENz+Q+rXAE06p/ETgV/g/iWUFG7WVPSyJ4uEZ4j6aUw8t
NUHaaOG01GD+d4PiqaYDKVUOsPHPiVHJZ/k6B7gc3krTWbAJI7QUCXnwGCXq/IaLYyiYvYGTXQID
s0RUjjk1pjwL1zoY/BIJ4ZFof/LAdi9T9v8a6zedOb+XAJlDgbCy6G2iaLg0TK5OrI7p/9X3zsm2
WbMme29XJXE/1k8bWUp1Y/2ulDeA4DxVL9X49UpqLp6LbAi0mN2LEq/IrQI/YMJyBny/xPlpmW5u
WfQMpVbqtOnZgUGhwW/cr2yFDBgpTsJj0j2QPMR8nkLT+bLK083o340psPt9w4YpBX+4NIX6VHIF
dHblWkLljmkLThvXqUZAv8spa/SwC0W+vE+JrKTCSZxAtJfex9PlOfBVOm3Dh/uDs/WqbOh7xhrl
7OBmHpz5cHFoNizC1odlvp1O25ZCwtfbywRi7EQZD5D/IhkW5pavHxoT02SI4k2FNO+AQUdZkyit
mgbtADX0fMg64N8XXFupj1h7DncX/1jp1jtMmZL+wdZ+naQolsEhptueQoSrh3WMrFcrDrTcg/6b
1ZHHg+cmrqb0heQUUDgoxWWNIC9qaXRS3R/8tHI7h3K09zuoK2j8PZWujhO0Kc61mJv0jT4cJ2+l
C1HyNTpxhujAch683hzfv6xuHDIUSKJAq/VpoiVveoJ57JB2WvCxg0Sm1Fv4mJ57I38OIufRZ8H9
Y/HCXBz6od9/0AqV7fAGP+R5zBJEPay87rpZu1vy3DkoTKLT6Uj/r2uMPhbFeX/hsIAMR+kLvEu4
pxvgSn+wQTivHgL4xzz32PY5qmYZp0D9Do3+wXWhzry+hMSE9cVPCHHfQriHwKsTG+6PLGc78k1I
xx0WGrPM2aJ2y90LOAThzdZIjcjQXxQoUv+Mtw9biUr/yjyU5A/DK6g3VPMEoxXVM2f9PoK/m9xV
iO0ARHgvH9jmlkcB2V7H6FOccgv6N4wUjHaXbzPl1kbgQjoOWBmtnNFzlumcAMI5BhU2VVDld1r5
qpAOaeMIwnRF4OKjzUoQigGlWJFbueSoILdz99pXVjwfEmEEgtzgu2PeeB7FPcwaB+9plzXNMUx6
FXy+eXYpKzFbs56xbdrr4LUNITAREanxhFE7MXJYDSnPZbKQl4IHMt0i2F3eJdSUDsce32tGwpCk
ap8SQq1d4AnPZEWbwBKWHZ+tzHW+Ws5FO61eKuggCsUglnVvXq0UgkP75XNccmNQ+TBBQu6aV6Xo
331aTn72p1WzcLgs011QP7AfZFeHZurQlchDC7Ag4PaOpXEed/Z5z6/O5WYKiuOQakySFRk8VeKv
yzeYrTQSMwpRe5F0CwANjrJRy+ff4DXDkboT3gLMuOXaFQPa4Hi80RdKiHtIPhyZcKJ6tnV4NxlV
USwSs/9cc0ggXO1PUkHj5sbWO3J3AdFm+j447D1sac5G8ENGfPUfQfgBJk4pa4I8y1efDBQJfW8I
LdCfJ+MKink5Uqw7VrQRN5SIzZwALQoJTcsLPSfqAmph35+2zS7bhP/TgqxyghVbVj0kdU82WjHg
+vhp0Xk1WvwTsqPsrCpgkPLdNJn0rbod26KfJA7FpmhYR9h51JmqpiLf7UEPdEhuaPMehK0QDtFr
T/btfWQb6wuARiwITdl3BSu8FKa737rBryUkcn7dDXZYeAgzG2ze3qf+qcmkj1zPZW7o7ZWo+vQq
7KhE+75v/LgqqHI1w4VEKHHT1+92PtM9Iu65rMSPjzhyqGAh8GHdBzgyqOpCbJfgnqVIcbyLSDbW
3vFnojC8603PEGmGoSFluuoxHGueUVxZ/0522fJkJZWKpBARIQanyl3YMs2WWst4iWIlp9aTpkOe
O/DUgycmxbnw/3Z+SUEGgcaw6btDcll6lmSCZMI2ewkCx2I+BP9kEBOimekLZX7LTcVo+tAaiO01
OVPUQjugjcgUCXVO4KNEKwjk0ts9p952nvO3avbxAa1V1cnmENn0CO4PRuj+tMCB2s3KmPbVKw8d
ef6GBg2pHuZOxSdXKjbnNdGZkgj7NaJDLqOISTcSV7YXg/ZQLSijm88c0e+n6nnIw4eAG896Pnr0
BebNfZcUbzdJtYeVAAITydwn7Vdas+pFxlcGcgloFNvuwZphxDYPY9qlbCsE2Li40aQWb99lXH/v
6HqAElLzCy6IRVcwT1+XkLuP5H2l6VQ9rd5OKM/15nHhWxXOuVXwie298zis7L1tw1L+Zw1LoQcm
MFezFdyWWtKQOwiqMjWYNzd4ooLFCVcerKHQicP3xNIcDSy7ikGGx6yiJNcHHqqUB0p9tX7QuzpT
iXMxCxuSmyg+YQzOH4cZNNMyzxX72NBMllMt5m9noUnfbBbwXYHYdlFrKjgbtieIGuJJAIr3ayph
0FcYKJlNZpKx6FQeGp+AAWPQkmvAL5geoS0XV+ZwefXKcEpS+YIBE2mDAnaXp/pCikxuK+rEho3j
JiR00IkzsxeiYbR2n6TKXPNNBaLhJR3k4aq6KqLiCUngBQQQLia52lsoE1B1R6mIIg9M8PxqtRao
AEDVGfHCL0fHKpFdEMMsBhSRTn0Dlp8btRPkfy1Mm4xTRSYyCDyKA5WF+6bI+R5xNMn8JfyuYYzT
YqSZp3FRmk1Izyri16dcRbH+9t4i7CQlGPkwOPMGXyLzT2AeVDj1hcOEc16oemH3brfjLaeQVdsQ
d8KV+eY04kGDUUl+ujIFsSYlCLthqeZvLARGr+0kRXbZvfR2IB/vF2eA/VNSb0K/AMzwsp+jf/6R
LllTJj6W4mGkQH7LcJ91/dXjwxuYnmEInDLVKvsnwMF5RE9eAlLJNCf3+737Zy/j+9+G5joaBQZO
fLVlDXM2Fr5OtGTJD7SqFG7RKKQwHpqao6ltMaZpqwD2G1Z4PVLvAfC7CZJnO4ZlDukntmHPtMEV
Mw2ft4djiCmGpCNxuMGX4vg6CvTbHWvhnOaoyRLmSjVhj3/cXgmvwQNd1Svu8+3K41+ELDFw5tU+
XmyFqhYQS869mEafoRDPwVjPbS1EOtdAgTKivos+W2c5B04NabvfZgHlSG1AC1mqL69wF5+nIMjn
rL+dCOmPYPvFivUjGFn+t+ygZ7hXFp2EBc+CNV6m8f/TxigGqGHbg/aSJFLcnNT8g/y7duBGO0pW
RDMNpi/OzpGxEmXSwwfEaKkyQH7SO74m2pAk719Ly22ESz4ZR9hf7VvNXDn9d0aPAyKV8CNk4Ck1
s6/kU2O+kwxefcm0x0jK5z+lFvH8wjNKOdc441H+nzpDkOjQMlvhHmYZmycwazTx7wixl9hY/opR
Rhx/YGDZS1fbl2msB5QEUZ9qB3g3rLUf8y+43kHgz+bf9eOKtKy6xhRMc6E5KHpYgQrvmC5Vdb+A
1Z5pLP+hNROJFSVr9K0BsLr5125PEefO8O8Rx9q0eF1YEdbpJYzAUB/re6fF6Tbyt4Al3JWP+GmZ
O8OxS2auGkNBlgplvIwSnodgtDHhX0tyx54U0gHQinRzxGzeKT/iSR4qqnzmS9RaliNjGLtbmqcC
QPrbL1GlYCpkWrk66Cpor8ZGwbW5WiBL6J9yQ61al31LzRxd0Mqye8aQNjKSGDC5oawrLRCIZVef
rgP5CInGulVRhevzkOoelS5eEifYtz8VVW0OlQDhEVP3citlEygq0pGmS5k6GvIzg9XWp0e18Ybt
9/JGbqHF6rkj9wRiajqd9R9IFT54rJskE8rOdDu8jpr2fV8cExVcoJHkGazm+GDkGu5E2ainmG7j
yrO2PZv3bkVaY2tM/qbkBiAlOHCY/iEjpTT7nkziQFlk4pKN9LjQDMgUW59zaRKybJ9puDJqoqkb
64aFaQZZPL4YaR+JoSaSPorSgr5d3XW1u5DErhQk+D9If+LrAvt5NfWvDs31pOxdWdQdJVY/Nbpa
TAYjxaYPmhtHUMOAXMVUKtXwZ7pC18DitvaIXdTyiJOcA2xaXYQME69eze9+wIbsNosC3YuNXoXV
7x7/5hEE/qUBZJOFsaCHqa5KWhKmYGtMszC8oMGWzOhZrUX9IcqM/+CNY6gbInM5rylUkBMFR5jF
dioVVFV5gEW7N/WhRl2uV7ZQ8EoK08V95IZH/6TDTf43NenF2EyFJm/t3WEv5w92KReqxJL1cQPw
Z3+DSwl1wqJW5ECLNvK/5ILm+1IwMiSevURLyUGlTSh4m1MoN2WWRWPUo1u0ARSgvYuTAZVQkP4o
aizQ18OhbCNr4N1vw8sQnhDCXF9MNwkJVee5m04DexlBXysBV82s9GRb7Vd6USVpvJw5KFdm+KCN
XhVXK/SOwKO8bX6pQoUZ6AySDJsUlnZBOnqzpANJwr3dcC1KAIDKzelepNCI0DB5v6JCbNYWD33u
HM4wCE3XqYSkaL2+aq/jWauRYUMaqCVhySTxGBbtIugT8+4Jb+zJ8+458e3QDy238Vtr5anDGjzb
N/UQ2z1N04EcwkdfP2Lml3tPzDylMVA2T2BrZGFbOaHmWs45/xmIk7KaGcTg/OBXobf/6HKErTqV
E33vb18BVdHOylFf8i2yVw5jTWBj0cMwmjlV2yWD6bv4Mrwn1UlyenXKi8lvZoRAkZSsrcDF5yxr
DtOcKdfGiK5p121UtN2plKR0JyLoTTxutLQbCtDKBLg8BA9+JRJJEHk78cWYOoGCv7ahSfRoWEN4
qO1rlqpqTSJUnHG1+5lN4P5GMf9OwAyseWJA3IOcqO8Fzcv3Zx+NXIWMC/lR4hbcgFpGqMU4xhUC
3ZMhnVlhlhVhVf6VboLkWllQQR9tO+V3/r0hOJlCnRkv26HpDM3/A19xAacCbL2ZYUwecf1Ly3R+
TKJKCuPtip4qHaNJxgjkC6+qPCmajQGtrKotOloD1pE6ln1y1xDy/8rE1EAl4ASdcCj1iL5E+h9d
MQty+1/pG41HEC1AnX4iEmqbwycS9cri5qY5uFI93X6/2fzH0ErDTwq+bSJ+waxq/NDJ5lGsPk0b
y9SyQuf7cUHzSMX5bmSk3FQbB9f8z5TMVHG/yspLK4XdlkLyeqCTSk3P2EmuTc4lQEi8x6zFGn+R
jN76On0Xp1mubkJ1kAneHGzOH3FScSwXrtIMPg7dpC2/ZET47jal9w15J+tALQW7QeAmw35asOvE
V9iQAsqN1VBTIJ4yljzMeqJ2NVaeMxA2W7oqsZ4MvBIo6k9uJjlZFQlT/9HgwL0ArOuzgK5RSFoH
3pWoC8GHNa2d4rP8sIGJyEGE154/m7pNSsvVWNITAgHh6LS42tNEn5hgVujP53aBooMmYCvhp7jN
hmPz9UKoJNEzBGZEsJ38qQTw5HvGtgLAGDiMvERHNUUaXT3m4t1OKHnfu9xyyrv+c3JoNQvbymPm
E9K32JczZTvw+R9RT4gyGP9Cs+csZNQ7+Y9bh12rgY6/6q3SXVAP+MTyPdi6XMW4kE0HKC40+5Z3
uZkHmqXBh6XDdV957Ydgb9Sohcs0K7D5MafFwkyiu/WtFQvIubPAAhVdfulckj6p7NG9cJBDjle+
amdTpHx4HG7sZvMiFe4Mfphpno0GOnxndfIVpcJ5pV+PmhKWbbvugOvfXBtmG7pXGLrsf8J6Q4pY
iY6W2fzJw4xSGKLHWvT+sEssZd+jh6uaaRVN0in/YnJ/vd8MPtUMO/1eWEuPKO+wOZpMPQVLJMH6
nPn5R0IpblmT6qbFhOoSNdGhkppO2nxX316P4/TK4uUrNCZhgB1ZNOyWgK0wTdH919FvH3YpqrK5
SgBxXn20OJfInQGd0XPIFWUiyWXTko7Y5ldNex7qDHqeZeBS05ZMf97Nuqh/fmTNmZH9343HeENN
lQD0CFQtWvOp3vCl29pJHBPbM/Tm3CYLrCYdnP3vCv+RGfwk27h2KJ4cgkxAEIhYYxSGkMEDRnOW
StOg4Hl1K3B1JVDs7sDjOStHMuHuhYQ7YDZYDHECKO94huD7jOdF+zNnZCmBEgiZxwHmM3ZRk45e
+2U+7b7iIolbQzoeHsLKkiL1Ehgo9zlXFHcu4rurWaPzhwzuYGTYb3fn6TeZ+oCM0hjohxIBzwK8
2Wf4BZEyk5bXWFeWmDRI8os70R7tD+0c3BnkxILYSGn1StaRCr/KZz3b6CbhiohLKVxFHGZCdbeV
rDNpKb+cGGcl9GnT1CLi0n+wh0zM99MHptioQPnEbHxi42Uhl4/kaoVFR6zBxNg1ZF6QudR5spxe
dwwogaFpi+00LlPy6/Nqqbalq/CXvAPuqM3OsKZ1V3UHrV/euIjIDdxWNng7BeKCg44TbqHEY58W
edlzxj8QMW79OcspTFW6IfPwjtnTJMeV+gVRwaE/DLE7/F18hkKwV5NRov2Q7wZt6KbUNekb2R42
5S2WgGcC2W2RksWmnthWeF/mhbgvVHJ4IUeZfo/8giT4mptANQN+h62M/yDiC7pWdknFXo4lGVpc
sg4/w3PlKcqNwXWQy6J/wz2WEQzPQs52KjyRp9ejI9N0YLQaI/rC2ujn29GzSdblVai3LfwSBgq8
k3MoEY8oovf1SOgx5/+zXcPXL6ted1koVP3D29wDM2E3zvupx+taMZWxJw4fZ4VFAemhpHne4Vl0
1jaVtp0omBSPtlJjb8kwb7l0rPsyJLKIK9H0P+lD+092knNSHyPilc1RSk8vhZkfFujGraz4xJuY
SBHvG1LWlCvsT9YEB7v3MKiOqbTwl1InPgwcOOunkbMLKlo/5gm8005ghX2LTLLojaqjWwHuzuUH
QxxrkctN+kj2bnmlMpCBLcsajyUDsCKWPu1NxgLG9zbl8L+Z5pBjh9tFXYDbhcrn+/s1zoX3bAP3
tQk7aF0jLHE1aIdzKyWbsNH0rSR7pYGpiL890Y7YlQJWEn4wTDHMSve7bAUU+z6oRk6gVshg4lW+
YkKm/hxvTM3zrtRt2zYBjeM7Q4DP57S/dUzXMuY1CXqqPPebyyqbmZGBzSrSktHQ4VxpOVt4olC9
fTS69Qvvi9um53dKCfTRCyRfNlHewM9vW6y74w/t47xv+62sq6l0Jzn9k2BvcmNriHP7bmp/xQTq
CuGm9R/eO0sxDNw1ZBGB+ZdclyP3WliTLcCr5kmDeSjnU3MYxsAFqRXNVU3+WvouIWfT9vXqLmLr
U9qQC627APpxj6a7Oe2Vt9Ts+Lia0HtCm4Aq8GQLaMsl3pHYgMUMcD+KSsdfSIbi4AQAsCrx6CGC
FxBTzxrrF7z4uZLGbokb8tp9+HZbWWIiLy7eX3rsmh4xD1JEYKIdWJlMMNroJ5sPe/9JXg+advXs
L9EL3HuEPhJaKLtrOsJOXS9O53bwp5ERwrCslb311zpxSrCAjqL3kom0EcdFdH/h0UlfZCDIjA+o
iC8/ypbsh7twL9bsmTYbxuP0FLJhZ5HRe1/oiTYH+k15Ky1CFwldG4mTa1+dZ9xhkgDQoPWP5YDp
JVe2hygnFmHf0haf833tYlF59PQr9B0OtBzn7YphJ035c0jdyHf6APLhWj8GqejoN2AXCI4FZskt
n36vcYhoN4an6RLv7PYrger3RgjTyXk54vTQieIUPjW2qZqsLqsktTtIfR+GlNtHDnYYGfMw+w0G
8MEFYR2xVSKXA4xy5ArP/8/q96qBAg5LEzMZ/oyvP4l16blCKji6qMpB5zfSa9uPTK1pJsgPhe8L
MhxFfnn/rgm1pf5KccyjFq1d01ObxoF2ocSx5SXL79GEiJlxvroAyc+s8TQXGabRUBI8XajmRCBv
aCv2t0T2/3xnwBhbzqXl+Vsjb2BDFpvbKrHrb91DklyoEIv9wKN4fdIZYZWzfJSkHOkV0Lm2NSae
jUkE644UQvPiR+zWrAO3CHf+Ndz87XBfPM9A/scKPaRSmlJXpiwEm+NadFB4nl0Nq9mqZ9PHOQwW
Nnh4drLechmHz9a9+JQ9n3MiVQCIeKm/bqfeSpFVD2PNLJxe99L+8X4i1Y3fS+mXfVdWyyBNexuv
bfH+GCzCfSg4SHYHx6ZQQeu/9QWYxrxZIiJl6tz8V0l+c6QjJQ5StxldVs8vki9xZjpfMfNYTE62
BnG8rKbaV/DA3+q8ko1TwykA5zCXB0+7MLpkKdtXFmP8W7dQrcVHJDFRr67Cb2o8rWLFXGknKivY
LDwBLJKUX7UpzHnmO4D7UW9inelaaMzjC1W2cxGI8qMFE2L4b62BJfJLAXrimiFWOrag1VyyncWe
GQfiZ6zHyAcn2Tzs9KOlnnmIY+IgBymuRhcMbCpIaybH2/dXwDTW/hNR0KeA0zcdsU79g5al4hGz
BFCm+4dc91azggXQvumm+1UVoQobijrSLlTvg0UbzWGh7t7HJrgYPBsvRWIjjaEe8IpunyVXqrqq
hG8xPH1Q7UaFXkM+MOMZ0XRnkMBI71vefVh09y5uVGBxUxfmknNIG7lnKmVCscZZtoRzZnsIGuZU
hp+04KEG/LkfGZ/p8g6E+N9PA5QMrF3Hmh2QIrCSRL2ogxcvlQwc6yDAp7EE7HJ9hm5y1ks8tlDI
MS1x6/TzwV5VTCHEhqDwq4GD5W9qLu4bJU1ciB73uKS1GzKW9KKPFYdhrV16X4fcIasdjZmWEIHy
ukWEGjkJLo/UcGU6NiJdsvYc9mtg7exCWFBffTYbuLQQmuPhI8rUvUqGvuXdOpGrbihsgOeLN2XE
t+24iULDjrbDkpUONGzfCFLXwPaIwurWQD4KCr3ixCH4JxEjs24oA82xFYBohGGRoTW7upM4SYPG
tn1Ko1gPuXiBkyhebhYzqq1kkC0YHufdpxn12bLLAvkt9bt9ZWruI4luPaBGwHc2YCMtd6Zb/vEJ
a6G1Rd+wBQZmz4SqNPWZGH0HWkCWX+K6/UqUubM1HcqMAtWL0jsh1/LsbQ0F2sDbzDRWNjMyMhm9
7gHE9paHrgZmFVeH6/M8ypqUyl9bwUfE61mpJo1Ka9jCrxOYxBUceqE+wjbBUsxLyeOT/ZkeSH5E
YiDGVSL5aqbb8MHGaFjv99k3sCG5PxNWtbtIkPUHbvhIgT4beQxtVZa1ghgwSbBpeQb6OJfuLxK1
nOF212xCpzI1QNT91c4BotgUqTZLaKmheSztrMPJY890cymw4I5Fjkzj2fvLBK4TXJJkYC7CLLm7
TU81WHcHt3TXDMBUoP5cLwIvagzMZBYLao7+feF/ZiDH/syjtjPenOmuevGiUXV/tKLGRRZcE580
5bTe36eYLsdDkmSyGcmcvmipvMfbxteGSL/m59WKx8FSaha74gKqdelHVHXgh0aEr/+sVLzLr4HE
ngAqNIkOzE2EQS3iSvwe8Sz4+sCkY9cC3/5kF3N/qZI+pT6D0HZ1qZROby6KGrtl4B0EI+NTvZvM
xfNnblmT7KRhwDwP4KVBrkN5NyOHuGp5GnqALEpoA4bcn5bohvMp4oLMvWMfxbiGgQuSDHTO0pGZ
SX8sQeTqbHypn/67rwyuipTHMEQmJXF2Cg2kHQ7J4BwGLtqRABewjbXCr9lKhhY4ahQnQycY8mwc
japSKb7gLO0SJN4LtdMBrEIblkVlsDjByAQJ3UHmZJvWP2TfBh9QD4bKNOvjvsuCvRLKIQDdR5wm
YVruYWpcMt/Ip23IuE6zoX4svSEBt/F2pwKnHOZ1ZVbkJ44jXvSg+5dtrXlGrKXWD1P+OZi743zw
uuROSDjFP9PXi3KibmkcxPdsiY6u5pu/hx7sha1CH03I3quYq1+IjXtkgIULDX93mxQOtcslnX7O
2sDx4BRru0bSibb8b5vL4xQF+ibrHRlmjteDOgVverepP5naicT3FEozyXTBbW+jpTu/9gDGTq/A
CX9V9YCIgWd9QypoXfcMH3G1utd6nR933TMKE8fIMLkH+8IPuvw9LVXQU1JE3OJ1cBiOnB4VFm6e
ovcNbhw4G8ztbUNm3E8OgZWCwcpBqPx2MLu5+npZSRZSlsreXYTtpc+Km9+K8PlqIx3okOjPcvp6
GPbEiQz/DuUl58ewGcQCJyUjL3VB9BOeURo1Bnot+4alcfyAtg3hYquLN7zK0qqTWFUPOFFD3fEj
Upqc4fPRRvCJbPaAKytixQae4HOAIAfw1vwyej9/HfVd/SlBQEzOvbfdHa2fO/2OyeLgYcXP+TMG
Yz+pBQkV9WIDQiXBNVZYBkyLRPsXno0/qiFZCJXf8KK+dDU3DWamlDrdonNeXx4m7fn+NztbODKb
XfSfm7Lm5Vczvo9dMxawiDb+T2Ibk/mSWpTgHviA/iilLXaC415CvPkXRYqR1YQ7Enog352YXrOt
Wa6kQF0lYC23MbBveaNkDMJQj7bamtXCKm3cJNd0QN+oJreT+vZfF78X+NE4ZxeEFfeAy1A9iLpt
c5pxq9fivn2XM0HeFmYemeFtnrGZ48912JCkDMo4Azn3nWKxRqDvxl+sE8c4A1GgDZxU3hqzkTDv
5KDdtfii4nhbFnVPz6xgV4PppIlE16nvi2Xt8SBpeX1yR1i+COawfyooyXkALuxDkk9irUNhjldX
wN5ik4O8rZIl6uP96qmI9dPRAKGfimE6vIIa/vEcy3Qdvg/JSCj3yXQCnAtZNPS9yXFBAJasS9Bq
EUq7x94LQyuJ0twVQt0DC8q02ZJhciv7iqzEiwzbXesI1zeHpIdgjyloHJ/bQTnTdsZPZy6sC/27
6H1BF/34spak6f6wcXzrrVCaDea22VFoQhuJpF1oZi6h14nSTHL2w+VvN4ic7ddUqrNIWTB8CDIm
Xvn24PuOD9VXNGy1HxVaUe1CZZbg5hIKABSoUMx1lYpFkajSKO5paU6IGTxtDyDYOgcZ48QaGd+C
i1poKPDoTDmDdkCimLKlbZj3SbgpYwPYXw+eBnzyuyvATrBW5JKZ4lHvpBl6yFqxMqvUTxz+Z9T6
tHCYSy6F0Nkw8fc7EjszMw8P6FgzlsQXvlNuzpG8zDUdIHNu+W8fS6s2s+UvQaMeHcp7rq43BIR7
CMciXiHWtjRyFxEzoENbhH52dao3eN/C5CU38vlfqiD+o02J7eGfMPrzfl29HJU60s2S0e8bHnra
U9JryzK4W8wLZzQCEdGcbuZRt7ZWd3Nkq/5s8mb9rkDSuV0I4aNBSGT4jV7/X+sUNfk17zeEExaR
wBEXW+9FP5xyNev66iBo6TU8pNAQuofLoGqZRWItUfO4BU+6BHP2FpQTdaBgKduZnX2cfzcMKZje
anbqS9XF0IiNYAQWFkWr9DoGYQSr56sGJlpp+KcJ4fOcKFTpW5JdTFnohTsfCE9Eb0/n/UD+gq9T
V9HnbAFMB5DZJkh2Dzh04vFnx1ATZrU06nRmAO9PHM3O7hE+Jk+Ra2cvTOVMH+E17oVfKQ0yUn/k
7dOmslOShp6hGHG5zGKfAWEXEJlpzjQP1BU3HpoLI8P5w6vK6+9swa2ahjgyLDCVr7qotvdevTdo
j9xOZvKHujFwuPo9PPTWNwD1iWAyrWTyyHeTXZ6mAAdBmyjgmmD5sBbuHlOziqjR9cCSfQKREKNJ
2w8w5J7t+T13AJgWhM0qrjcPXse/aSoJwQ2+wVH0gZ1tXSfX0ooRHDqJSk2rwtzqjs4zCtU/NROu
eYLakbfIW1pPBeol3jVfujVjiSE1QWva/7vzc+bC2M4VV6mgAm2aHq763QyhkZjBuBaO5W19tIEa
s7mxrxXPGRHgQfFIlZzxsRNNeDLrEW4vG6T+BZiIBbKjlh5REvGNZSli2cA1zQiL9cWgika9ML8l
9xf/4Z85WF56T6UISHJyWpA6hNJDH4Hybv3Db3G8yb/7kkd3gCWTVu/s2LtbstUQondVMHjiJ+p1
4fZRPX9UOvMHCfM39pXMfKFXPahD7guGMCJMq0GYOY0yZm8pPCGoScY5SycmoVgoZcSJHVcLmHOi
9VG8iJWL7U/8ztDzQhXEfU7j2+0CnOHjfOPAN2QGKq6rmp9GU6dPoALviiC0SHLwQ2Dv7w4IeLdP
fuv4XCMdcpyOLfNp/NwZbW/DG0U5Kesdhs8H+zQWHwte0Aj7phWVcJ9DkO+BX2CbBdJOSnpwxPn9
ni3ASyK7d5J8lPFxY4xNiI1fkpoVuTf/UiO38pYPygSAz0jgpH/07JnWJg/Cln5UNHpNRX6hnLZS
VzvyY5vjyXdDvjJTqGaMPw2VZJritj8K2EeqBKfUPd7sUhJferoz8MT2Z+C8Bm9bIJSBpiVRA/pi
kW3EOgj7DOnwPTY/HpZhMoYOKKWYrHjo7bCXrnvPSp5iDAUKD5e0ny2/jANP2NInQkqo/3nz6d4w
b+iVSmJJD1a2jxq7CrRkzbF3whwjw5f4g33oQGkWu4qTXVnxIJTypNmIwtODaXizyxhpQsh57+AJ
5szfevmAHyXz5hfYQdDzxRYtN5atOqeZKguY5fsBrAFRvY/ioL9JQSA32WoEesgwtyGwffcoGigy
2btCWfIkVZhZgSzudNmUE3jinp9YtjyP41pWKaHc08wrp6lCdQ7n7bF/vGDP2rQDiFjLPeFjUVyU
8Dww8XeADD9j3ITvBoJfxbbBSsoyKyvCKhKMtJVDWaokzY7pVtjAiJUm5k8ycSgjtUf4b9q0NFkw
9J7CgOFF4oFZ9WIZgGhqlHtezcjdhOhKNIZIGYFaxVANoUfrBjNILwIrYYra52JPhSjid5+SZ+Wa
zLtodK82UCuSmr21YFMfqfwcnFChOUxXRtKXftb+9dYOjHqplJKNJhH0qJrgT7jJ2ODg3eLm+bTe
5Ttc+1PYkDKIkgJ1gVysYqCHNv92ChVFsQYjY/Ywj0b1gkFYE7Bp8aT5bUwKuAvo/8rc1MoWQhqa
7bPKS4kG0qa5aAcZbFHa9XM4Al8Vw+gp9Rc2OQBgKtCpl8zoIP2PCdju2n9g7U3OfJimrujGyRYx
8aOxJox0qS5mZG+vvWjBMiWVG3WBMco6dhXmFo9gimszZbDZ4J54v89qHZ4b9rs87vM/y2j6N1t7
v76P3MNzH5rc3qmZibinmJFY4nmYx9DKBZfDEF2wFbenkh5gFj13S3mz++c8ljKHAPB82V9FZ28/
NOsXqPKfOVHCOUol54RH6cULbd8psyLlCLyqTFeFgX4wD8EaNeEDeNZLpnx4wPySFwbRQzbWbHz1
69j1x/zJfb8S0j1SsJoEvVM/YY7YeaHhc9vAwzu8M/oNawnD/NyNrx2Frnmbqjx3Q3zeVRAP/OU0
N00k8FQKPHnudMM4/q8iPvwxVyDrAyqsXCdGFdTdOMQy+JbC8i4TimEcsf/KqVE0gC4CP0SSfX9W
8FM3KbBJkiST6Oc3iF3HQir1RwnEpHXuvAUg0Pkx549pdX1RBzMpXBN30Ixk3uk4LU1Uxe88H9uu
qoJpxKCNvCnFqAqaSjO5PHn7xHg32n7P943rRR2lhGH9d9oE1n4vaxsAr3zQlcjBrNg8kcsoqm4D
abuUHo25pPXbqoQTQz97ftYq9/61Q+PbUKk2UhjVv2hy42zIyGURZfm8qacnnD7z0kAaxcdpYCcL
an6LDcI6xuuYUfDxuB2ikFO0Mf4zqvDYE2YZCnW2x1AtK7xZbedZsY4o151Fcv0SBbZXeJJ0Yv9d
3jkKP8Fa81ExncZbwc6ja/JY2eRbFhhVg4abFEeHx5DHGHkblXjPWCzMaS0uUL5tVMvxlE1dNVr1
82rH/CexXc+Wadm0oQxHFW2O64hisSQZuRrdIH3zCRC6zvhSR5LMOh6I2fWB+nhUJ3K+db3srkZJ
KXsIggwl7MMsDF43pOzsiSOuflhJF7P3JucAAoFJL086wS+Gjj6DHmw6CceZQo4T/w73CEstZuN7
B9zh6zrFhNzGCCwPEBGYW431AMkh+DBdn8D4LTJmsNgo/F/cDQAteBo46qfw7zoGtynnHJBoULZp
babFSNx2Zw5SoJ7u4wpHwUZZI/879GuAPCXWerKeCxV5DpTFmKmbP0xJ7eUU0hlc4ihhaClOmMUg
e695VaUynTqJE5vScfe+aqbd4jLQndlyBLyct9x8aoL/sG2A1nLSWfMVGUvvL5B/3OWu6Haebere
UWcx/sT6AY+7uPVbqs5j7kBOnzNhq574KZWHAa1VITsfheb32DB9vEejjV87+WqTSL4pfRJbztZl
lUPL9OIfM+A4CYa9tgkXhv2tka6GvIQMv07T0NRo5DsZ/8iZyimpXTokVKy1zIFY2GTkIikXo6De
G953iVAfGSA7zwtokzx6+EOt1oa79dbGBbdKPmKvM2uvRTBJ6iB4AxrDx6DPsGmZIyA8bkGoqkW3
aqKB9j2kecgE2VzoaewTZPvNK2E9h74TDE0iW/LIngZwR1dNIJi9QjI/Gqx+tZXD2ezEPmSmJAQ7
6ebwnEgTUIrWBvtMZESiIfPh2XGfwBHQ1R9i34SC1Kd2rJ5TlsCnT67zRwLtni9scauIbLpl4EtR
tVSjkurMILoPNGxp4WvnXSw4LvDAXkZRCZPH+4LLItvjx29UkMTITR7sX32v0VEGqywle26woM0M
mhRR7EXUnmr0juPPpJbByVPyvwRTYdOqKtby5c7IBBKHn15PJaELDff/0sKLQUiyv9XhPs8wiObZ
4/LuQX2uurFXShOQ5SHZvuSLcJ9QCfcxgqlrsfblqdTZbG8ctmNvVL1GigG866rOG+5DeFsPQGiO
eUlmKmDnL460h87pKhdNb/JqPry63taEuZ1gAo+F56pDzypmwEbM+n4lPA+5d7k+tK6YxdY7ANJ9
jGlxLF2xwrpKzKcG3pnVk+fu1erCm4iJUK9VR+2BRUi4OP+32uB3bBp0hgCOgu7H4rf0gyKo/dsY
PHFK0JdedoQrmP2moTPHA0jCb2TTtNMcfqNr1ynj286cYqFlD8CrLrUeok93xpN6H2GE8SEpnPYa
TTxQKNbD+ayF+UAlUaRXUei30As+ThvFlk9AO8/cEh/IAp7VN0C5tHJwWnsTRGrf7xeLH/eKDRwj
6HRVOXM7WQjFs6PzKpiSJBwSMDIf/0OsrBi+2Bq1irb2M7TQAEGZM9iOTa7y2ukCX656AHeK+ggB
/Xc7a+GGQzjG1r2jx1z16Si4Rqbu/LCJsGFXMuWTdvbmJPdpbyUUHurzgVGaW8jbvWRcVuvntLE7
ifwzqYNkVgMIHPfoCdPNrS+Dw7IBl9yDJ74vdPvZu9M+MtV+Oz5821ec7n7ODKglpWD1zdrfFcTn
dEh+a+Aac/o53a9yvoYQSl5LxmPUr1rSOz8TgTo1jATVHqS9c4lpSJYzEqzfinitvp/u0rXVDzjQ
YJ/D11jA1g++bH6Gj8wKOzl/mEO2xzGjNH6gMXWMHNdZsGAPAsiWBuinSrWa6EJwPnLcmJ6o6TCC
qAq6v7tOpxVN5Nt7I1wZJG2czEjFSwCRhLsU7Yy7M4elKmkDW0knSR4sS0/1h9m+dZoOSKslqwR0
NifDK3UY5Mly3CvLUzO6/AZSWH1h4FDfAhLzxI5s4ELQW7VjIcWGLM8UZBrRML6C9IqJVx0GwW0c
+O300aF+7Efym+k9G6E9kw2feSWPTEMTL4LW4/j7/G6XnkWrEbJ7j+u2b5AU/w5fqJ1xMyYoO/bD
vAgDKncoQFg13ij0l19rhImiW1ll+DAHtHEQDHG+eRKXfp1ToZDYh3n+IW//agGGtXIu83fSJhkZ
nUGchLnFkhNyWcC2Cv8RxNw2W2WVcYaFaN1izIhtqCG/42MahJod5dlNEHfiF6SJkP2gfMXKLp30
S058vp56biJs2X50XAsaQO4eRx/H4dPgXkA1IuBGhLFUDuwxvK5COFE1YzqbNOO++aDWsjJN0Col
bOmB9Ivls3Bmmy1juTm8kZyEQP18ROZz/vOz5w2wYlVA1BlVo8DIAN+OYgoCDliphMNB/Xe5YeXV
GtOfxYotl22kEfvSyptJ5QADJ6pUw3ste3C1DJsB5zoKSiLAZXrJ6pvyUAqV3nRhGsZ01LvNJOD9
BwVV3r5ac2LVpLRftYzjPYGh3HPwgRMTvmbXlBMTWNfCG9MTTo9Vqez4ITeBplBEb8DPqPP9pCQd
x9LNFyRFUNbHiDouL38wIYRPc/I6PQILsd7rTtIDOWj2MFlQ6FKWkseV8dyJ+FIg8naOOiG5FRDK
iaZZfykx3Yd1581N93hW1mGCi43jXMA2mxhEOFbhU/60DwuBvTI4fAAeoajD5A2mS8h6fbU+1iME
hb9U9sZIaxtFmashIbwqbm4LnHDNn9U2an6vjM1KG2V++tmPXRw8w9rAyAvfVYzmMUi1B2a/o18B
hCmCqeZYbHJtu+Ocg5Hk+JhyIvkW/Fkzv93zPRZpUWWt4Sb417ztH0H6esPKrHYBonKk9G/ivhUd
VgsabpPckNMFYqGEa/s0gbWaXtqHqPZbc+11FfBPO0RDezdf9eC+Fz+Sf3UTNXBPu6PJgK18070M
5w0a3ACnONCmretjIlVx2Ax9bYPY0HdplZJcLkjilaVNLKkExCwdOXgUBbjlIbOOtLiT0BV3ASed
Gj1EcGM4dktkk4vHJhxRP2AtPpBwIlurZNBLafivSFiS/A8y+PhFEj2zU/2IVg5Yn4m5mmF2s/12
auwlo8nE3b/lou4Yqb1jo1VmocIllVYDpJ9oyP5NQ9hojUL0hpRgQwRs6KRcOmCsZr5mphgWiq3a
66wReeTJ/Ev9P3o41Cn/O2b5xPcUvY/3r6uFNRxuTdr5V+DK1pI5N7Epuk9qOl9igL6H04gjglZP
sdenD5/p+DupKCbFU9n1UVLPGFqDYX/FEZDZttARkBSFYgUCClEUVOZFLd/Xrfa0YPP7/gq+3Otf
sKWmIgi5P6yW7IKLUMEUsYQnqk2f5AonIvIbqWaWfcY5pHp/Q3ZZjmXHbdBk2mG+3+uC0+i4CUIG
9kE2ZK3enSXcHVAzLG0f74w0cEzoYm39NxLp0GPsOOW2jG+ZxnCH+UQdMlscpTpX20NJcptGwB9F
Uch3s+VgTL5Px+/yHj9Po33FQZVl9xbfPCnRuQ0MIk4/dJRr0iCT3GbsopmrSTExyTnorRDeIX6L
85XK23OJf+7qyXHpRhxvbrat1WhEIAQwXHkKRLclPB+KZLLfq8ZorDMI/98uySfX8xCpQnARP2y5
NV188zF3kP6zAAg50kB+WR8GDrl8qI9mup1GMM0pkByJ3ywN5euyLGkOYgHatOUbqKBVXkdwqwKt
J15CYkm4ktiNzdT3F5+fAUlWOhDgYeEteTugtSZpHnqp+5EFPkaf/rwlR379GCmU77XgeHxWxWqn
TxM5075JftYx0ojTXGycZyKG6liA/UzkO8y4RIncLuP9DB2lbxYFkfoHjOhFyhFE1RRpJL7h6JxK
eK6/y22RfuYNmcz/sE9hak9anKbteAQ6aM2M8vDXGPUVF43Bvl5Ok7jFWMsj+p1ZeBBUeBOTbqd9
eX8b9rZsvgyGW4DjZRC78BiyUrhy2EJ10OvOvxWY6xGhB5YMSu9Ndy5XzmzeLHS+iNtRZBALXQHT
ezLH0gn+BKFkbSxPjYFZnJrRSm26aj8wTNEClzMQixs7mAXsUNGjy+DtqIobbqjNMjxWhz+RYhJw
9YjmYKrOPWwEuohfGLNJ5Kow5MtOVTwV1GJ8BN01Qm5tq6Nmf3vxy9N/R1Eck4IrF99dkXA3LDLM
knY+P0YheUfiCJ3/0R2KEgJmEriUbbcpkUX8k+8IiH9h/cFr3Z51H8D8Vix72zRe5ES7+sB8W153
7WpQv9ZVWNUEyjPWCjXLODQSox3PtFDLkaZmKFbEflOG6iEsFP57DCRXJZ554uh0wtyd6pzLOMHh
yfluS8giBbtNntPUUqR9Hq+APFVBcc0hPA0T+aTqcjN4g3u+IkG73QhXtpDXFc6UULvir7ZFbe31
53J6Mm2mvg51wt2VlzX8aNjsrpusdhaViODjz2Hd2tFmIWDSusnc/QRLn+WUfI29qd9XZZSvpqhd
GCKbT8OCBnmYXBsP86L31VGxJEy5pjBD+JBa3l07U0PRI6RptvPH6MxEIDC8v16j/5EIKMFpUtwL
91Ik5ZCrFoNJl8Q60xpVJ4fyBJ0XTdSBQSdHoXQvkXCeaqXPFuoPO6bmSED9Sk53P4iq0F1tZvUS
0vMvxkizIfMTNk77S+8Ia4tbWDR2R8G867dF6XyPl8oqq2voPvfl28EmAZ0TIZwUAwdTpVCocAAV
qZ8h4763gcPeXn+SYF0xBgpd4gA5HzW5OYJySFF/ZaTzGxaCMSJG2acpsdvvtREq2xRgqGa1qO22
fRXQoMBjy/PXWSb0O3E/GWL0ImwFiVh0Ef6aGh+8MP++sd7AtPw+4hjF6b3aVd+8cos84VPW3fsr
RCEkDHWaf8U8QGOF0HEsQUM0MQSN8DmAfBJv2Hvbl/PC373sdsiQ5ZukYSYElO+dQyilw1SGScIH
CxXzIG2RSU0b6zg23qEL2TYbmmwrkUwmjbV7x1VIb/4JUI4wPOBfj4qudoVklrBT5udgAng90q1H
rDPwTTxiRS+hmuWp9/hl5TxSEHaNJzDukl/9U7lNCz8vBNCKZtw/wfP5E0YTK+cULeiTU8iq3zm/
kYNUMe9zXvkf4TONG1cRc41vEwH0+tmaVb7wWWIekvGQS0ZVVi4ePWS5rdrUJDp/PUJ7SfXHmTys
6FWSjXDyvivCVc7sJLEqGgFl9AYWm/iPfE/YAGGTXC4/DC72nRMZ2idTvuOJSPTNUOtEXUmzGh/o
oMpiVJdsd/oBVIRnrOj8F6CypWu16OwmxGekQmRz5Sh8vCeyY+1GA4hbTHx8AAI/g/fwAY7siuys
pJSFtIYuhaApK/nqX42iFDDtMGMSa/IOTR6+Lf3xHLvwEfvn/+MHoQth6R3PocPvUKHlImkJV41P
LBqo6OtUKNjwM/le2u4P2eXvCfVGPi7XMFhTVna0D918mVyr0GT8EqsTnmShAA96GJ/9AHD8y0Ku
SRM6nJVcoHG5+B5f93tItKSjn6fLHgS2vVakczB6raTOO5nCmX1VI7ozGCCunyX2jbSLz2utfyeM
fW0RhrTk/TH5y96IfUP5Lta87W9jTGyPl0fSOZhXqQqy1txBuWeXyu9mZPtRr8H12e5GKFeY1l33
jgYctJzDjPKxgMrSiZbf/2+Xf/nkUUl/qPBapK778Qyuy/es7XEQ4KA8ywD46UyfzviHphOCElQZ
I/r+P0PiXG0jICl/U5e9hWYWUz0IN6Su9eytBkS73cPTfDydSIFCaflB6/q9gCl9Mzv/NpMDIgaa
f68kwDQbTY8PXZjOGs2IW50JR4EvYS6gYBOYe6x3wIg1IRc9jBZQ4zqw7QmKM3TgtPkiQdsJfv8H
pV4K2D4Ha1WyXfugMmY/nAcJoV28l6DhbJWui6BWvNo3tXnzByXdIHzS6ze6wV33CHwcejY0xpD8
sHMHvQjUvVwM11ZidyJsSvu6lwwrnbIu2ZW4HwRxwInf+3+p5LDm9r95f0dJ/ZQjCx6PGdIAY+el
24Xbk1oXdJU+kkEsY6iNDTU4zSDDZYml2lCvl7sMQk6g+cUZ6+CL6yCv2Of3d/PvJPJNiEGVwSJ+
xTwcv1kguvFV/EnYcUCjPWMHOvPOUDWJvdcFd95Ub+kO+GxpjoAsHoguQcdmrlD2P7rXj6vykTkE
/n5s953l3vQ/SfO/CO9lV6+KOVnHd43RK3TystYn5msIGT+eBBkh/xjTz99dUkYu9fbcP+/gk9PB
L0QCokWFTqkUaPiMmn1aOEM42bGsyDCUWdKORfsh2TDmgSEutMn2RelxuZa8ZPf9XRvR/6Hoelb4
S7E0aZJA3Y8SFBZwf/visF/ePD4dwJb/IUxtugZX9RFpwWUGOjRGLdcHmlM/vvI18LU6jQ3jp0FI
KVTmTSOKF9AvIScYax/A+OeiPkZ09iE3kAb2zvSIZC/08eBwRdo1tQUUWwB8p68j2nxmls27o1BV
13S3GaZpfmoOox56v0p30HqU2DEsOUZXVKh0vE34sRvLFgIvgRHP9lc5756hU+ZZ9is2AtVbLM5U
40l4V6kJOnDhta1jbhBi8n74N/qJPze1Kt+rE+neCTBsqH+l4h8kEir8g5s0eCnkoeRw+XSPFP8A
moSvEnOfaJkkA7ndfhtfNmkCkNVT1oXzBFZ4LsuSI0CyG6mwkQt4uYkTy3eId47256KW4CXv9C/L
qSjWjrjLP9jSO+WWngTSGWZCQqn3mA60aFzsE8VoqLi5tuHUs1qZKOwoIKiXW3Kcm0pK77gycngC
k7MVoOsjdqML4MN2NFakdEnyNEhdztAmbFxeLwAk/VjoCD+eiUN4y31fIi+0SPXPnbYcH7HzRdly
eTy9krA/lBGouvheFn7lWT1EBLMZuYMEMjx+1a+F2vU/UqYdP42OH/iRbn/Snr3nL0lpW00UTy4g
SLT9tXMgLRXvRjh0F4xrZsUFG5TINjMi/zyNTQBUbncPLTzSg0kurpfmTEwveu/4YaSldAwzAE7Q
kUqcX1/z2SCpc2l05tJ/3hSgWkBspuIbNWmgdegziUwiHExbIVtObVs5gLZ7jOUpqSXJB+O2ZkTV
IxOOAxPU5n1x2Dj4750gi7DzvzvplWiAbIiX6GUwrRR+9kz8oPJ7olZsCdOVmgm7mYElZMDMnIGs
jIuNDKN8cGEx6X6PP0wFirzGTVrUSHA8P2ZMuAfnPg+o5PkIH862rtsikUfdAEl6O0tpbtxxwQf7
9ardapk1vxY1Hb+z8YBVnt4rTmh1c6iogE84xz77hoOFJ3dbPvXWDt/vvEC0RQH588kAY3ROdY+R
VSEPjrTCByCUcsY1S7PQW5hrodatUMusaY++baF0LSMQ4CxJnflaFS/iGFmMjovIYsPS53ln8tMd
GuPxOCqQnBAyp9+T0rv8CUQqHdDEjKyYP9nBE7OixD+VjG14tpM6YHlv1oTREWCgQX0Q4tjh7dkR
pqCTogGi726II1Hm7M0p4WBBS2kr/YTGWTq1KKuRU3qwFvh/om/1Skx6coM5KpNzggaeAoXXv2li
qNZ5HQo4C9cZwhtf5KU9eJsVD100ru5dibxDXb8VnTvil+Lh86dAad9aeTwbEZGwb0NpJcEvDe6z
A3Qtc5mhRiVQzXhLC1sVkioSrYnKfy40ME93S6qM04SMvc+SGJ/VGwOx7VZim64vJAna2U7mP3b1
aKcCNUCX4NefQ6EpMOqs67wChFTgOTlmqzStyQYJMQSsVRdbeXWBxpaWdZ+AK1JEHfqALAnoMk+x
U/bee5PUlc3tAnA+EnJyYoTOOMkc8cPU5p1mc5DeOCEqfX0KKY4c1SSZmbaNCk7hy+h1uaJWVHT/
ilFZL/h67Vi7KmX7ug8RKrFtrOYMV1hwm2lsS2k0KXO/ZGEPIiTIJzATNi/pBqRfEkCj1j5CG9zd
MpU/DP9zbKjqqTgdpz9nv7pSNS3l0eukKgEGi0X3i88GLiiueMcayuV4HtrnmTqduXee2iYoKnHa
ZbycRW+00j3uAGMuWypAxx8QlD82NcLZDBUR54+veUSNDSXusE1uBCWfid/Po5JIiBjZI4hjaiKp
W3ZAOHNF9kpdNyD2BIescC6CZ5VHuGG/A4esh91tG5JHVXuCIVXr0C4AkWvF0fef6k3wwHdgnGWt
HOBxCbMGLB+QCVvn5dWNGeifb/jWzU2znvF16AVk3eU6/22FUr4o/qxWGXo3sSNfm0DaFR1HUQx4
0j3TZRWtN+BAMn2nVHiYKtjrPDjePR4zvz5ldVTqpnniYcLlG/zYO9DsGNKnd7iP+zYt/pcxFumm
tN2z2eaQ6ZKlG0/zCjhiS+pLYxUpwBj8siB8kfu0moUxep2oxVsPSfUplp6QzcsGnnYkI+oqc8qI
W5JFeTH+zLwoz5aWAFhRpWhWLlptjqeGew5Q14x9q6NfIs1nPrmOHvKUYWpr+wZdI8IcVHjT5QDF
D0ilH7NTcn1VXb4c9sW9JGh30Ol4oXcxybB2c8n58cX74Z6wrzKhuNWkqamL+RpKDwXzXdYGGpXk
nNc5S1oqh6p10EHFihcFn7SR/ojPyXKK5dxqfOdsXkzURV3jQrcf87V6kuMiIDLEl4XCJkrDh0R/
QCbEsDuyiyARcORVakGuBXRUcnIbmZQCOkIcKRdsEC9KLxEZO86NvgsfmVOeKN57Sd8klwRe0xWw
bL9Tkzad0cs1LcmtVSqC83GepykUyK+FqpeZz1aE0t34YMnOiQlsUvYEUvcHlJOlPTzs/tqzmdQz
fbxgmUxS/u1pkCFzQhLinMnKSqMOkYhpTd5hNl4Q17LZG6uKY8S1AsHyvaO1dKVj6AT1ZB/eMqNX
ddwrWfwNGXs6vViTzjOW5XB2CPcAXgwaWyZHDc1nh75UQo57CsADDaiXMlJCBuzAWZMncs/X1AD6
THeuD2VMujEe+ygr2aPpOPRxbkbIQkD+7KZxo6u0fY+PEpYq4/Dwp/dIV1VSmlcm5JgHAmeF1vhM
11thPAP8oEafUUJnOMuG7aril3IM/8K8Ntis6ev4o7GQM8yqKpj+6YFneWMrUwvENk4q++DI9fhu
fFZRGEW8tDQXSClQzAMXRR8kxe2BnOifxJhY26TIdxQ/xRosgTr5khKgvyGFLjuf2oxuz0Yvn/Hf
ENoeKvQ9NdV/0UcTx2xe3C1ex74yvpHybzkXmdxX+5ilVWLLfgvHnabg1XWRBxa0nqY+T5hxP3kH
/QKtaki+yMX7qWrmh81umseL5hKX7s1SrUkRjSXoEhnt3kGXDJauw7cHSoe2KFihncCQrtrZEPyn
VKAYaLrP3ClyYQHKktkkMJxaFO/NOMhq0MbiAw3Q6UUX4VBLW5wKfElka9qjJWxbuRd4rS/epUMB
LX9UHUikbyhOK8y4fIJIbu/o86i9i34PDcl7C3oIlb5BxtwzyWwNqbDTeMnmCRG9WC6e++Pr8dK8
jyIBAzF75zjfvI2LKuwQ4Qn48NA8+kTOoESmhRPQbW/VLoJTgVBjohRk1irfmUNzw/bT+TtTAy6t
CE4Yq1btWKitt3aVsF5Ndf4uJpVU2JBF41D5t2raiHiv0zs/a96i8ppyg3+nczqEME6kYUn5+j7M
C2EnENtj4uya+iBKSOKyosqQaNN8M/Ban6FrxYGXEtZqhWfS9h/u/ufJAFt6mjXXkTN2vNXbFBz0
/+/fouRg+D3krg+4YKq0ANaX69C9AH881HJN7Kt1BqT3zrx0ZIfev7FhWvoOHG0FsijRt/umwkmC
y+lWr6wSIK1+uMfnVsblixANchlgVEoUXS6yoB4MfIKxeI+idsmH8+6xOjBTgUFASHxBVvv/gf56
d+WBm60+iF5uoLWFcXqWE0rYOwKO0Ail3eyOXwFwVP2enf1UmzDz5l5CmWTtaZ4tenT93r3ufrxz
uFOy1L1sjgvHuvwyQiA6JKZijuF305yNKb+urABteLPdjcFfgog1GOtUnMFFJkfCjmqaUT5EG/Hl
rWggl2P92Qg44lVlKiSvBRrW7ipJZfzcnFpNB2CtP+X9sT8gLQAC4RsUOSWKHQkFklvQQzKH7VQS
+1E2OMPsU3jKWzP148CLqdTPHb5AHJ+TzE/9KrfSSBDkn8bouFAWZuiz7l6eYikYlq9mEWtVCLsm
92W8qomazon7CQEOVPw+iv7WmseO2cuiSSFKOCTLPWOuVLfGNaOc2aq94A6h8VDEoQ5TedBagOF2
zLzyB/vTYSugpP6UBFGtpJrmnphCbuth672yNEi+uHEMCQ9RwYFvQkfhXGEIbW6PGKepoA8xm0Tm
PdEjNUZiYpEj0V1OBVY/X3Hqmvi7mmqelmh/JAl8KjQ5CMRLQpauMti0iiVjnAH6Fv//kiJoVeNk
goiKAwePtS6Nd6yWljt5r3sPXW58LjIRPXqI9sx/QHZ8F5Tsoky2sdB8gMh5mKbmfqQCY65ZjZOz
XnGKQDeMPgMOxueSaQM/yQ0dN0o0+K8iEJua/ByQPBPU8X9AB8EFGSMS8G6Z0Prlp/MPl1HLnimb
U6qB/qL+WMbEUqM2EQSVbvpl5ER1aJMMFTTMtD0Vm2qnbM8dPqCCjMr/FWhSF8ogSUDiW3Yu5IUr
d77dYjeSUDH00KrpBJ6BNI83d9V37X9U/hPGFLZ4swGEPWqZ9Q0F1PpVLvdKzAtVp7CjF+mUbqqM
bIfbXWfqpgsmVOwJdmMzoTR3HJf5Z47jZ7N3irytW80qOTVYsQtMbeFsRY68Hjf7+vNfVxEr89HL
YHrR2QkvKnDCWxCFRT22GoFUpr48KUePwyz1PBV/ubfycIvq5e1M5GNFL25ixfo/ew7YssHYKcT2
A8pK/nFX5/ucnMpjBxQz85YRd4yq+N4GkqCkpWdYVUInJwLw02UP08+uhkGOJsYYvKlVkIcKisUJ
7IFKZoe7JdDq+iUyDRvWw2kc19RDt/xyB8cp+AeiBY9do9vo5YslI+aj/d0kwF8EYbS2ju/yvpNF
DlvXrY55Ai8P/B8kmn6XET7zUCqF38oVyU3vA8RM7tHKCuE2ik2woQ8imEajqdDXh9ZLv/EN9SnO
82V7w90AhVCzlsQDy/398PjJwonNuXoZCyeG7IBmtU5kHUSW7NDVmv9rUOW3Onpk1+q8qsWBW+iN
nLAllq4mJiv0sBWAtT0Z6GSo1kR+PS2lmPSGja6vtXcgCOV6FPrzSaRgllegrZr3Btbfyx8BBqUm
fGlr9U+pP6vtG9s7mDxlWeVJ3dMYx/Ik0csB4jiWoblhXesNtS0fE5twXlaHN3LDtlZZ5I8o0i5/
O4zWbM4QdhOPN0/2q/NmkTyxFjrJID0dkIXNtPJHBWsj/NumeDSDRk4ayiaBf6Sw/G3N7ODtTELX
1VYDxs/GssocnQrST1N4baLkCsl4yK+Jon3jQzM17c5vW2O2WEjifXsxcoSIHa+DZ+0ddZHfkUAp
No+8D6JoJzNgb8PM0RyO/AuQhJQb2t2zQVxq2Twgs6+aPPnWi8avLpXG3Q0wG1kubkfvNGfc3RYJ
2+njI0P2mSNgY4TpfSmn8WAMCT9eDO1Cg13nMSdodQK2BBCe8Nwedxqkf/sRTf7dMWJJACcMTys6
0H4usVXlD5Qzk4IfUuUN/1IRd6crN+mXFAuFmPqrvP9IQMyhn5HrJCkFmwMda1lqHiupRMn/yd7Q
QVcXc1b1gBceq/OAD8DwVYMZrUaidclzeiQzZHv0oBnTzNP+kFaMx8ev9hygG2HbU4yiF/DtOGWQ
atx/7jwLNvU75108tk8pA+rLSlgBG2OeVLEM1mzT2Y4JNRr25c9UA7LaD79pLslpagPbj+vQiGWV
dKiDbqrz07MXvabv3s0WMX4MoxrBpy/KKKB8a1Z7HYUYCxrhmXHgQzNqFppv5fM1NLnvzc78o8JA
T6rvxVRSqpFwigHoF9/WKSqwFfDsdVEIOWD9+KXSFAwnkrHBEBCeZVVJYQmmDFghy6xz3itd+sL+
cV7Ru0CJaczACYdWXbrJfV2OIaCPEchQsHm1zqY3NJ9evYjf77pFGhlpqXRLBOlVvVZZTbQyLJmN
zon1oJHtzKFlagiSyGdT3PqAt6vF/GTf6eveBo2OxQgU/X4IumohFEHB7WuUzsycpkNTdJuNTWAY
x17SuQ48FmT3dMmhtIyb4YePhctweAlqZTO4J+dX58nlmtM9e+W6lWvDmQVqh6z3Fk6zhnBXspTa
lRdXxRt3UXKLn/StcKbyNo+6YMrD2r0GqjlMWQr0eD6LzyKeF6iNqfJ+kfF+nYroD/hLnViPg3rw
9DK5TMHD75ufnYSIMGDUH9uHlNpmMcNFE8yrTwqoktXURXIQ0ilZr/XCkfiSzbB4JspczUSv3LQ9
ca07mrunPFzovNPOMuqc2lV6v0xFfd7ftwUU+pBQJ/7Cd+hpWUAl29Pg5gMzH0lD7HBXnRD5Prds
65C9H0K6raJ9jCjcPCMNVLZDDqe1lHADtyIvrnLfuUd0yIbb8IHN5BuCWE3C8J0dhLlPrOTRrd7s
90itUg8biDIXsfQZmk8oRVNRPl08wHbW1uuWAzeY4YBqp0HZemZgwHaFUKQGJZNbkk46Vf2xwddu
8yGIli3qeWPO1M3zEbmQp+GVIkJtVDKvprMCZ0dXUOxH7yOh+OZ1+x/KCKu8SiOwplK31Q6XZ8ak
VInoWhyQ0JVr90tslox82LjNDgQT+NziCGRLWbfJ9jpIRhGkWUWp2Aa5wbNuZ635yMwF+sgbDp69
cbiAzD0Lb2UivPDfHZezkMwY2+cXk1IbEtKDIVBM3p7krQm1/bozL2BU5PjO0hxAe3NDi/BDDbSp
W6xN9l/38lei5dxTU01tAs1Y/lcdhjlI8tcV7gmezHpLMVs72CxPkUUzCvO7FgpAM39tjkmU3GAk
g5Ten9tQEov5+PQX2C6jZ48yTGuK7ptLwqHoEHBpDbkp54uoxltEiqNa3X758ZjBquS+wT3u7lyP
SV/KhAC7IpkCMIXGEWApVkhCu6feOC5KBMhscoV/BQeRXbmTGpgOa8U6BqkXq8qyiDMrUELxryfb
cQtszV9ubOi20R8UJ73RTxskLQ+45yGmf53pp0atIXJAJKsOt9j3bL+emT5UDTQXxqQee4+BUxRI
6q60IRHrzq6WM2n8yIUUErUr6e51dgWacDVeSNsgHDnFoi6bI9FqdIjS5DU34+env87vd+4F++zY
eNqsVV4JqTdzOPs1OgN+/gxMfJdq0ioWcv767Ttx031s+uAgZ5tWmznX2nr90ZQ6+MzrJ3wdcCGg
JOxzWSn2WUaRQw3onBrA5UU5b4bWNRkUsGq0AIVkji7A899yv5goqKaiGtn89pQzmwc/IPuM/btp
Dm80FNeHhG+1DcnqxjtUKbMb0wyixG4SPOUQA0GwyESn6VBDg7qRwVyk8eOeMUzCcBiE4OYJLgzf
3STpImHPcMzOM2RIdrjTEpM+JbSfYIoXt9t1Z8zDoY9eb3R4US4K8wEPznbp5vrQzFGkrAw65/GB
oi9bzi8GNa/8OdxZ4O7a8419skSIyfT0orrC/eQilckdbGLR775VN4AiVFkh/n7Ut7ZUcKGr8SUz
aLSuxcrfYzwUs20LPYBrZdvfsNttzLjHA+Lr3o0xM/gpecMMyRlO2JQH0joLQJ4zPsU3wy4z06FM
17qofKBY0onFe0mKOJDBtIOzpF/hvOTyGRa/2yab0Kclyk58LVLzGMowTyofW2h80P4j1wmD2TPK
qBe2+WJYJWGUfmD6POpdZD7XID1USkS8cuNAdm4OKcB6fMRFazoxcVI7asTy19Xk0w+LbWMgwVXg
fDreS+BGjDVGcZctn3GeKmK0DYK4TEcYDSkNTWuEaFmDRpV8D+anJLrN3BPiBc34n9PBtORDpZtL
c9AGEVsyRJ4FtG26/7ldEJFbbnUByEEq8JOJyjGGJebVB8IOMlP06eaYJHROS2jl1yXLqOAYxhEn
7AN35x52OXBuThcsU+9pdRrqz1WhgQfvRkU6dWKwfb1TzQlQ39fRJPWwsy78NMYsWp5nnT0mOFFh
Nj0SNsuH06W5tTObzTHe7m3xjQLXKijMdCuAZB7VkJ9iQxI/281j/F2rfGpuUezMnvBFV7sd1vmk
NGltQAqexpkaQVVzz2TKXUVLZPSZmRP9h8vd5gQYG4WhMVvbhwaaCEkhjnkldhl3DciSKrN2Lb1o
kR3IYZsnlfxSHp5Xs75uWZw4TAraplVUnoHcyYRaBTO2ygXgsYt5KMDVn6hMKtHwCnUEeRr9eD/v
anFj3LGNw+IzMA3JQUdEevvYQbhZL/d3Iv0ddIkUSQjhTGyfRlnGnuCrZ6+ly5yQflmOLhfWxb89
Ce3wjgDnt5P4B/itPGRyClcTr9vK91yoeXrEhd2kUYYXnKEV0Vs20aKI/omUXkvPTbKip18QMtMt
Nb0BYihnFqKyXQee/rH9LS+78TsElhl0nXVFx24Wup4A7yGlc8RZBu7BmRPEo3/MpwbEz+zfI174
CC4AdlXNORbpeyokxy3ixe5XMD1K6jQ8pcpve3iZakkghRtUWHBY4f7PYnKKGSgv1q5Jcj5nUSTK
f6NZQmrDVQs7yryJhBq+EkALJIC+RLClub8pIjoyAkKFhfiYYDYSxQF4+Y5EFM0HAc6q0segJbvt
FthrEcB999mvVDK+XVp2NdmIaaAHyQ/cwdn8gwJoA0ZriibyGTEX71Dd0M+iSNR6AqWKAFpNSrzL
f6bV5WjA1gg6BmmxUnYh6wa83gZ6iRknkF3ULNVXu+bfQJf7tx9qBjbw4uhGKBvnT6dP7SiYHo/F
sdqLsOseNoX/gAxQ99KcpQqwAnZbS5yJ2O/y99qC3/MPBT4/vnwQOR/Zs+U7Z8IgU+IiNn9yopd/
DfwTYKtXoXeIB39JyXTl/2MBbhwTbfsNZYQP53N5TK8RNPw8cjp4BKicRGRQQx2zE3JYEoXrNWoT
sEFUOSoDW0CQv05UvusJU56y/RrDxKNdVCM94D1hUawKtNQR4qeq7qbKFlI30rw6WtiG+H+izSvD
mx7HI7C8l3wJFnEjLht/3jHYolcHsCGN97Q/Watc3ejAVuayZPAhp3GfwfN2RNlqgCeDqSu/Aw8T
J6om0XzoA8gxFZZi8p33+9pGKzvY7Fsw9IUnbjCAU4RYvXBPfLroxT/5+pVEIpa4nrd2WzWVRJIg
4Gc1QFR+fouZSOIcva7TtlG2RvkuTdqF7u8z8lJrcevzQo3n4jOVhRIPctWVZ9g93cHvXqduJFDQ
CGbkgvXy1tLPUgvLaNC6lN0E368QorFHdC0RZqHFXeWMmtfZvQgDttTeCu8H1N4sdpEuhEkM6Pa/
HYklcCHzYGLVzWohRwzX0LD0EC227m5A/NAm2DwXoc1kdnKqT7mTtWpbsphEjaqMCJsu/syZsapp
dtoJadhCuClkC5+/YPGTyeWysXp/2moyb9TktKpeWPI3sqcwAGxDuktjUqnWOBcGe4wQmzZu0Im7
aWExuhjepqeIuBt/tVuRW1IK+PsSwPc4/RvsYyOZ95O7cHRXso04dhCzrYtm8d3FEeHDElR81Uzw
zohH2WnGQfX+VKPYANWnsDhYz1+dRup75+PplIqU/HHUwP/AvifrwvsT6ma2lq04uuXMyQFBggUD
ZyloJ9oBG23jpyjctCOqlX368ExKp52Lrr45Q2vCpomgC9nrzNdh7KMQ0H9h/1GNFxMIalhFyO+e
7eWMa9AmQsCru9N/nMyRHSl02cApe6vDYtplIODK7NM38y1KIfGdxi2EBvKljKS3dav2coTS2ZI5
sFKxSXcbQ38iBnCLjJac8Ag9vguNrSlGYWEdtovJycscsF16TIYuRZZlgmDzYny8EqjR1FhL4MGn
y84cXntm1dQLhvxeXzzR4zMNCok2c19JGEPLt2V+P6eGSilbPa6+5OkPAPYudRM2UripcOXxy8d9
WBOni7uF9XtOlPsIBC0goJqv+ph3rhCKZiu32zVcjo+T2sUAI0XvAMoRQXzWCpagmbYxH6jkzeor
HeIkaxDLOMtzJkCZB0y2HFSp1xYHb7I5gDrea669m44278ZYwIxj0aENV1x35vLQ0GZnWaWftYdz
dZQ3b6fBWFCcmcyc3dgWSnEGSxq+Lbr7USzpaTECO23eugLMVNhrBPzd4uSKthGl4VKM6Pi40ugu
8ecQTe3RcxDwVR9r7ocXw2CCjTb+l2MnJLQWyXC5YM1e9mBNA5rf4xTkYLMt7dCGd963UHARxJcU
s8m2Pe7g4sL1Mgy/cNykMhXLHGsDdf7R5/cgtnyocjq6eDj7FzYx2Yyajhi2ZfymYJMVhSdTiwHg
QmpKX16GVZWsufUC45DvNOhkyZMHCy379H7CbFSpKFKKTcR2XBXMk+00Np61ZhmoXqTVz6EHfOWR
y7URvD6wa3VcmMb+XMBWI+dSQSKtoXxz6q1i10xgQBhqefe2l48Wj3aXe8RcSxqnz4rfS2oWHMVD
8W0tLTAp99mYee6cWSNE+pkxu8xOOt0NvrT09Etodq3rSXW1jp1ibyIvAy+14rdvVjyJgFqGsMv8
i14W5OjdoPB8BRx3o9WFQpWS54T4c/LFIptWrpqERf4dVBM4QHK8z+oW7MhweYH3XtkULkqYCg1i
GIPJrzzGHNVctOBi43NmLFRvJogC7VP6q1YZlfg5t0IelwnarWMCIMJbLLEV1Og9mZ9GjNL4GZkw
vU35OvLMhBqcbarc/VCHNwLh9nVBdtg0tq0Df8CZPED4Tt90zMDNu4/+BL7VLXFYoMIcPVvTsR8W
k23xvDzCWNtTW9o0eqW3B3n7KOB3ja2H26TzlCHrJV1yINC6xDeAmoxLzp3y3YINj+ZsL8fqLZij
BKXYv7imBRIbNt1TlDssrAay8T2DI8bAcKjovuA9bKBYTSQS2DdIQdUfUCV8V4c/f2E5OaCiBAbP
b7Sg+EApNrV3pcDiRId3AKHFNrHnMXzAHf+8aBJm1U6vUoZeeBclF0BuUYRvyZK0uYH/8SP0nM2V
RTlYYoQaN19Fo5ZGNMIhR5RrieU328jXNy2A9EbOfFnNKzHEbNgJ2e4yBQ0If80rs0rJLcfw3qTK
U0lX3PZD/jaDC4DOpP3YI3ezOTV1DcntvytPDUiTeY+eyPuPv1mDHR+HwY9s/ug4GUBOtBMA0FTy
/tW2OlW/eiq2oKCglH5P1HWOVKXs//TdhJ5/vs4GWMYgmZ4Wh8UK/P9UH32sH3S8LLMmhJAVOAJR
ODRQS71Mb2z9xUVd9SAZs0xAWNXtDBayAV+Tm+DEpPyznrAjVQliVqYu6hHS+XuyJq9V3L45MPTn
vM9g7HxKnd4a2A0SPRXckYLLxWuvjpFKBl9ZQrTMR4NsvrfoSXz/JIm9vmCzKDIHhL9zfq5GgafQ
SsF8SY22hYpF/akIGcO5De7MipTsggVBycR3UiO1kM7oD5brJsGdMJKaMw7JRXz11EfXDz02Nlx+
evzOdWOXFgTEWUOOy92YL4xcpPclkf/iGx2/bHoZVx4SdvNIWMelrfAH5NRd5iu3/bfu2OQtqImF
scdMcaSMkZP6B59sQbDyt6OPsV3IAJ+1bC+Jto/Mn7FTE5aSRAy73opJ6Vl1neB8/Zqv4Lm3ty6a
OndDNH3g6VH6cFjN1M/OhjHK/3UQAOm95wG4syt1l8gemSbOoAneLDY9Eq8NdC3ztyK3jX1Yd6HX
Lz3uglQYwz8YqKHbuaOb3FWLc2G93pAY5p19CYCbRmsL6AHk/zeHKOKQLpHwFSJ15wpi7x9acweZ
gLyfjYxnopt0vIcI2MznMcJaYgvH88grp5id7n+l8Kc1LVtoauVVWyDdwgye0YQt8nnMdUENf6q7
613LEkASLDIUILxFGCP9acus55o+iHZvFUevIdoZd4Ifu3qhtXraRZGFPI3/sPrYeHciblEgg71C
H3ShkAP7sSIz3RdR7kdJmpG/SLvImLndki3QnzezEVS6NmiFELDYk3t8MhHFCYf/eM3f7VtikmET
0ZpdVrgCbT9ssLKQmCIRrQ1SG4OPpxx5bUEHsvTUL6UMCE8vo9W/VeQL6p5yG2dKaMb8U+UmlFUu
I5KTMFMhZvDW+aBPv2yYJnPPhXUfliPXTKK9HA27Uoe8VUG5DAyGDyFXMBZoIdTbW7evsDRJ8uoE
KhvvmzcVeRyOxTILFyGV0TpkMM7ibTuIrbflHQxgljcuPIw9N4p/o/oCobuAoP11IG65khfgITbD
ONJ8W0v+rQ5/4PDt8GqVzxbGpEJEgVDMEu0vtEQntC7OU/PkJtvIhUCA41PfaasydxUY0HfjCSsk
omIfa7k2wlFi0hqrSAfqdwBJjRiqRS3Ql/KnPQeu+0pwvnqlpWz5OAG2K9oJ6/VWkzKKgOMB8jER
dsx71iikR1QaOjaU84FG1ApvAStSKDOm2D15w8ckkZezf5/k42xRqBn+8aVYFwvdkxCX4PBOxBjB
jox996lZ9VAPlIRiULMMUX4TimuRzohSgzNVe+xB6n3bW3xcFfHkvgy7ekujykj9EU5aAUPew87z
s0MxX/DMj5mZtnERZEBgX0poBSd7u+jZG4uC4uME1NS8y9nnpNhUp1UxZd58dRKWA2fEs06dbJpL
31dSwZNx8neesKarKqA3zLaYZyxBgzCyU8somaTIV4Wd1bJnlymJETyIGFJ/CGyMLDckKASzUmiZ
H1gQ3KrfVsJne+GeXk1pasB5RdXhoFRAPdY+YGgPXVQs3QJlHq/2XLdbD1SqL0r1D6iHBVi05Yac
5jfYSJ/dutuS7cbfFnCqa5tEyphuR3c7+zNjqfQ7ZGy1bZslu1IqFhavNDYJdu9yp78yytsREzY0
OfQTRDYgpS5TiCQWGldIcAfGgCdB3dcgkk9DWnVXuF7lAyHV8fjB7LBvcsqTb8vccsmUlxdVokbQ
5Xq8i9u4K8LZUkmmmPiC6JJD2JB6/mcJdR8+yz1Z9dk9y9WxWHeHtmeM6nCjaB7rHOYPGUQKRx1u
7CgIZqwjaOiSJ+oPkW+hMI2Lb9reKBARa159VGrXyVr2yeAQcFcfdYf6lY/LWjeJJsZHPi7r7+U1
tbYBj1bISurjwAckR5E8f005zs0K7X08drwGEZZ8itFA9+zWH4TTEXKUaGjeUHm4P1neEpsHN2Z/
d5Sy9bUItZEddSyIghf6MxCgQPQ0XRxGVhQ7wOHaF19zLZ/xtMCaJ/pGtOa4YeW+bA01VDPUlAiR
IKiB2Id5dcUTWdOl6t6wuHjxL13xT7Z/8FQP+t9u0E7A/+RE+eSgj8vrzAEQI6rbrFPY6IBfLK1O
qYlrEKi4zJEaQmnINi14aTQwnoHroBmpXiGDFPhf3coUavv3jiHffeu8fpL0Yo4OeZg3IwEZ/ahJ
vA+/jjQ9o/4pkRXQcH+atkGGDLl2gr7rWsWVOm73jbP3gHmVmVM1yDjor/Dw5p3gxob/IrZ1Togc
BPor0RiP2q+rxJyKRGIbeNKA+tblDBdOjgz6ePxYkHq/x026VQGXjGw3u6Jd2TMPF7fhe7crnLO/
wnpSHesiAnihSo7zq628glbd8909NuMslTVO+6nyU6WhowVC2/Gp6V8djyJmc0qHjnIYHBU/pLmd
GgExGyV1Zku/xKhK/3LoeD25qVIxrvx1N3zlrQmVhT3DrYEH4VKaekssmbUBXqPQFNFRvgIKRIZl
Bnl64Kg8x8WPnJI9hh5/yRKguXR7neFMylY+bLWNuxrLKS/8Xygvf/pk2LgHNyQjshIK7bsN+Fnw
QxQCS0Hzv8bDcM0Mj9BdYuL0Jbq6dRH8Di0p5rGGW8ZtqFJNjhCBrzhuGH9GME7l4/cXIUXx5fek
XAQfCc6Qgb7/8gQRQ3tSMXf8Po0uNYmxjlChZXe6RaaijA+7V/MJxkSKC83Pw2Codqq97bpGFOKC
fTw3w188tCvzLzZY4U/ZkLd1u+LbUQaPmHne5BbwhyOUn1ePWVRHIx+b+Lz8SiA29DfkjMf+8w8m
qUjxqCTI0Uuy6x2aadgs1Ci6EubMZ319DhajmJzD3oNyx4vnUubQFQqPA535EG6AN0WB2l28IhRk
YXsw1Dcepjl1C0l6pR09j91UnlWgUfOxcTH7HQ8i4GCTiZbP+jT+wVbLh40+YAecY/i5xnTTTsvO
DUeJeD9/X8HrAGy78mckX8shaqWQoqMHREiS96ezOX3ofhbQuZ+tPtCbrOFloWkcjQxFbf09qtQf
WSGl+tMG6jJ9TzC1xFKWUlFW5Rpj0lBOOAnajM6pWShdXs4w1aiyJkfSKwstKu/WYJTavmDua16i
HsLMOhy6fqdi4ZjGaPf9gzfWjSvBCx5vSJKAc4pItjdgmQD1Onf2cjtp4bRbqkMUYfW95vkBMb6M
hf+b/oA8iUT0k8KIeRZkFxMDzNZxbk/rB5JeL38JugSc54aSUppTQc72X4LmPXji3nGUGOcf/63D
21O63q8QsHC20d6/wUdtFLG5Folk0yNa6y2oS2lh368UWBraEH6q1ipBfPsUlk2+MNDVyIfIMxz5
2AK4OPLlfdyplHxeIZbasOI1ZTiQE+hINt95bId3nawb7VshnalzsPLOYlDAbDQoz3zsL6xGWUIV
mqFTc2w/pF/2jXn/Ov1eATg7I911xZGoJDMAq6ROor9ZZeDpMbHv/pohphsZxZYq59pDCCo3oCmu
VKP6bhEn00Sfl9CAE9HIOnJMh2+Kj/Unk8xZxnISKmnS40moS21hg9aVeic+KeIyBRF/6TvsJc7Z
hOUSTi8pCFVxCtxS8hxCDBLE7aUeP751bEdgB+AmO0acBzHRLMzF/ogfX95T5EBSoHYXqhEjg9Pd
8aiS4l97J0jiVZ0G+tBqRzbSqoM2i8/UCPweg56hJ/d9CPm4Nuzermo79Qe9G/cBNGjGmtrr/oNq
FvbvN61NJR0vqfHw0xRSyHjLTXGQ4MjL/lU8qpJ3fOCc2D6bixa1aoiqeAb/OjeqFzrSwAkB6WT9
AXNhIjmQKANBSo3clzBOO8VjYrbdIjdRsr3mKDbiPJ8u69avl0pdbyshG8fiLx/VbSbU21NgzxHp
kERQN5EzKp6tRjHiSBHm7u43N6HOuv87+4G1gOIHaWnB88gRXVeKLhlvDBEe+Wb+aSaGizSppgUj
jKaFYrbZAB7PLeM9Yk4koygDPG+PHXnhT+dlaYQtQPF9FvBDTW5yxZBUEJZCm6140DpEACHLwrqT
LIQ/ADN2wqq/8K5TuTqCda0lZqKr6r5SQYYIEaZeYclkOkDCj8Hid0hS2yaS0qA4S8St5Zmagbe+
RrP4iUmxBexAm1+cfR7mLo1F0AWyVteg+39UYVXIPN31G/AQ04i41+LSegnc/5qaDTp6MceXjk0P
zX5j1wNfYLloVkumlGSZMMApEbhWlPNSlBH4ne7UhrD6Dl8XOVmKXwXpKvC3rNLFvkGe5lcM1L2Q
FuEv9250f0xLhprP4oJKsmjWhU6ZvDuOZeX3ebF8jFm1X32hqhvGhWbUEtkUnCHpMC58LJGk2epJ
yxVEUYyXmZRW7lJ+9exy/wvLOU+32ppdyITW/xvE0i+JeShkWMwcjhRUF12Vhzd3sO0h4srlGYo0
dg1Le9PzybeuWk6lyhdu0O22hGvrpwusBzzrkCjQf1fXBKwTtR7wzBFOPgg7vMiNniJI+n8n7nwp
zt2s7yOPSpFVRrMaZZDUkyFD4Azp0pXKHH7DTIKEFsn/2OyR/c+zJCdYm9rs+2TdvUUcD1RIhSjf
Xus+CgSfOAQ359SYQYZJM4BLSar3pkFhXA+PljA+sh+XnEXEgBrF3lAS1J1+kN9R/k0OFIc2cwps
JweSpntsJUUYT/WAzEVPQ2I2jpTIHOVgWlh3fE/Fb7I4fIjVAqfaz642c49wofVdE4vhXsuNIRRR
VaaagMWHUJSUaCZ5yNQPrejj3m1wokcNsPWeMHiDHOZVYxL1I27VGPxgnLk3GlxuBL8vAR44+b7x
OlzBFvA/UDGw3QC/eZ2G496kiHdBRKUjE3YeE+swnRN/qdBN+VDxJRhHGTfmu+gH180X04I+6mGc
/CivCOyqNNrVD8KUuHNE06gIMdI9ynJkXt5BBT5wOrgNJZ7tDCi91CoE8bz1ePMEMdu8AUPWDipm
v/+ghsKKxIJp1RWmVEByFkFFQ7P2GpWAtjb/TKF6skwBuQUxP3stNfsvGyl8PqgDAksGfEgdbJ2A
mqW+nCVFLAVnWIifshq8tAMSDwzWhrmeE3nlQnPvzg663a2VfjUzX2CqgWpU7UyrehoZhTunbB4f
naKgNL2/BsCzerCBhjLGLU1wRMshleMfEi38cndcN3nQQpQPrmdrcZJScdbRUKuxKk8B1PuWWxX2
O1xOQHRmuIbRXJ4zILm4FKIknbHWyFTORSLOCobBd10hdjTPcTzX6YUFQHlw0iMYPz7/TG4dA+SD
5zvQtnXCbyiSU4N964ujb+dMgG1JNST/0Zy1xpBEETNcGgytNos64BegXzUgkLqgFUP1e17DsK2l
imQ4dBbGoFfuLca4sT4qZpwr+EOEvzVOvEJDgky5MBwp40/5RzipAdebsfTwJCbbBjtVjVrp2Di5
Th/i3eSXeZsx7/V6DzN9XA+5pjOhu3KIy5NEdJmpT71X5x1Szz3M6GwqD4JuDpNrvJKHsMEov6zQ
VTQh4+wUX2J9TaZzJY4F/Ya9pTJLK9+IelaIZohhsoLiDTQw/Hm5lzJ+L/jAHh7/Zvbgm/FSU8Xw
Pym1hb+C1lp0tWDPtnYGi3Te6WWn7Xced3jYNIw2jVQzXqTsh3zzaztkNqN/g0jhGKoWEMmhau1W
izwaOkgQSYcTWxwDPszOOYYqeeGRFeO3kpUNOLO9hS7BIA2c4IZ8fZN6FhH3dTZwvyVP+3b0mcne
RO/xkbHrO8Tin9/CRCVm9oKdixaOn0clN/+Rfx0H0ftPkHBaYKeuJ0PnhxSZdgN09p4qX/Jp8rj7
r752VYjldQXgcLgznN+rnsCIzSqjQhM7QvnD3VTGf2/I07ivRph0Lpy8DABXmkNRXGkeojeQF3J9
IRDZZloGjq0BzJyhV5GCZDLszVea+i+rPZjeVDybkrNb0EihAz2bQocDvR5Q2VeWx2W3TlBbmF7i
eokAk6hjiLYE6n1dl0nh4XnNFkM2Bsn2N7xX5ZXBZHIO78JXX4TuhkxS8yYFvJd9EZSw+EdCqw05
AYbVHtz1s9DWtX42DMuUK90dzacoiEB5XJs2FEduNfVSxCTNMmXpJNWDq5+e/8u+8uBpM+cvVHsx
UpzPoqHY2JlqLCzcrJWOLXa1nnUrYLRpSB+GuCUIyFKrLUzJtcseEDfl7uM1PuZWuQf1nvuk+uK9
7BieCWQX0Fk6uACR8vjJSrBXkOUDoHUHbfwn/riBfSdgl12BjGqZwEgrGTG0UN1ApkdeUeAe/M+9
lR8U7ogCx1+wAzjWfaFomHQzLSzRZ1+t0PKTGxa9NKuUErNFq+DWwru4dXRpYbFNnx+N56HJyKdz
oGMBY4e8I5GjR4/LTD/WPko97wilMfBhNZh8I2PdE0U36xZs0Wi2HY+aBdN3RV9Vpjrgf5ZvqYx3
CJrjlYmBN2DMKIVyojomj5DPmhDT6BVcZJT7kZMTDbTyZn13GgGCIRoQmFHkba+5NKjSexOS/dqo
4R9BqoCt1OxFJa9E6v19FcY0bNt4xYfPTFaiV0zI3EOHe18ZYTAa/Sf48byEcJsyBMUDv863x3nf
sZBqkHuSXOL/1QWWyIa2rSUfdd2xGhskTRxpCOqDZnILWumPMD/9veFSDLT+WSWTrmPnA+gUlBA0
qIkDfMr6lbcZ9MhH3pYMS/4huIewwiD6zudcwnx2j5CNtn+ex0oAHpt2E2vKhYjmlksiA1wpj4Ez
pbeAHYTIEMNe5k/LPu6ak/kEBDskRbxgZvIFIOi5Xo8qYZMqvHCXr109yJzKN//nCPvN1Nq+Pout
gPquFmQBADHPwOqrBHCmKWKOO6l1VG2QPoNe8aa6uIAtnzXj53pJ+N0fmFy+XZ1wXnf27ZMtHHRU
G+dDtRnEFlpmdk77pWzU+eN1Xq+vOPd72PTLpeh//lPR1CpsthubzCn2I7sja6c7FA4Djcu441Ly
2TaSrT8XBTe+3SYh0Obt9RuVlW3iBpiNw8JYU2sZXFa7BvkLmpo3R02RwiWs7FTCe4yZ7HODVGhG
y3e9KTHKbbD/11K5TJrvZ/uZXJCP4PWGcHyLbrdzpcGGMEXd2SKkJ5r57aeXIJALJRxPUgpS/Y0Y
QhhPNQ/mH0kTypXpszfQYj5E0E6sP8qpW9YSNSISikm8nt9JkUE1ODwV1sPQDedZnN8TDfATq6Vg
8kOd+YS0IYHwHW4EIxY8h06aEbLbNEtSpwJY6+q2QvzKDarcLflqdd7K1/aJnf7dKB8W5f0wwtNA
QSF1N1zNLdWZOV4YuUdXhJo8ipwKU6vUy4pR7MhVt8vLPL7hcCFUyr251zN6RdQrvIzA9ZnCNCVL
aOoFMbAYaAuVYsojY/1M8Qoi5+vH/aKcS5ooyEY4Rl5leA0wcQadLIKotjXNijyRi2ynjeMRiVGu
B3ZB9nLAfX58CyNfex7y4vi3amYChDM7BsKd4Wj/qtbmdG3YB0pbZU8D8JiHh2PKdD2K5HYhTFpK
WUgbZGXJPvuoUtz8ZlnBDZuZ/+3L6jg7IamZeyegHOEVopu4zQyI5xb7mUeO1GiJ/h0+09sSNuoV
WxrZQuT+Wug0UHBoGgI0I4PEtuJKLTB6qH/4RgqBUdddiWNbB0uIsRSdxRZC/W7FzSBE/Pe7lSiq
h/9yFOxM5SG4c62cHhAPrzC1Xo6Toyh/NhsG49URunbTbo0faMoH6kFuLHFWM0ZrYwBnAyeZkeMd
fZshv4a5BWSv8xDbxsz0EUQe7mFA8fvOxrY79qzpyxk6shZTe2mAlMTd6HO0r73hrqvPImzzf+gR
j4JffqCvtoMOd6nW702Ot4P2G4OaIiU8HcTVmco6XUF8OM3rkq01TsqbLZCDgXXVZeP8usqL3KH5
f78ilFhvac0xCgM60PgsDo9abln0f66pxMbsJLrOTUaKsRII9hP2pojM6hxxcjm6ARogdqth9jgV
Tc18jkYee49lJlyw5JG9s+16vpmuGFZID2Uhxbf5q/UL1Z81EiOG8QfGozG+sifrleoMMncXzUYM
iqf49vNrtOH1mQ6qWO4ySIMRbQLOoktvQmMhdUpQFPV+vPEss6fbVfh5HxdQsGRRc4j/3uhsdcfM
F47Z/qjxuBSrffH4PtfMY3aK7PNds9W2t0tmQua3Hf9Pkh7pEgCMalgK7D3XZW2hz8FE7uWGMMoF
/shpcsMILSR63oYnEbT3MauVmwewm04bULpPmqmbzSMrelG5WWTbzMIFPyGoxxsHEXDxqnsNHcN7
2sxePE7M0DiWMCe/7gOJ+LW6wLXo9JSosq7HENwDDa44Mz2x+WWbAUZdiyKsmgnyR7HQ3ag9iyxr
0x9iCwnGH8q6odC+fIoqQsUhZvFUXOP+gKwQQC4hNO+B+dxkW/xtzr9kcoEiywb+RCCyamLTQEOy
yToLxuisMv80fsWY318FMYDOYjgi5lyttnjmoWRlMUp1IYWynXEb7fwZQ6S2+CuJh7CjjKJq739X
jNB3ZUsBjx52a2NhxeJwi+ZjBh7X8yxMlMLzczqWkVoUpyp7GScOabCHSyj3imJN3/5FgiPeWVE/
8j7Sz+HTIukyP/y9fV6osnngCJKaMLcIRpycCHUoShmzfnvY/MaF0UTDecm6vXCQViZD0tJiOW53
6Ktz7nPtvfJJVo7jOmpxwqbRbgU9RcdumlC+/W2MqogMQxuDMXFKrYMtO2j13RpHKmFxmb3JwEAk
kj4oPckq/X4FcnoTBca4BiZhsEbv4WrFAHy9NWYVIjPv414B5Saal6l39Uix9FDckY9dV3TNxZT5
716dBwjijAwmndqhJr/JgRJTugEXHsFoHZe0SgNEnWXb228Y+r3zY6st7lklKJ4WX53TkGIqVb/a
DKT6cFfrJZDNCd9MYzJMCRElqfvVB/rZIbTmGfVJg9+BWttBvY5g6Sd0THt6xvNT4CATMcsUq0Kh
QnwZFK7ecVocVVTXFsKSXjEFBOemLrAjFqyYgWizLqA+3ixXPjOXzIY05ELx4xXqorpTAIJuRqPm
+tqUfVQnaPEXYTlOTm+XR5BprrrKH/33gnomnmGGxo0pnAVD01zGRxEnePIDwGjC74TuMHotYCBI
ieMLSDs/EdGByOzpQMvJbtLmHbZ1fZIuKxkOb1uM5ZK3jE7FBBFbWkqpsn2Q/Tx+o13FfMyYdWfF
fF/irlqkOARX7qdiaQlOas9FjiQlnaY3d+ZM9OHh4YTeI3MGFrkmq+uq9B5wTu4Lqrjl7zWWoQ2Y
xRm7cTvJogtKHukaC0ZMztuFKozFLRoTAfsS1cdo5qBickqt7FcgNjWGbmPgv+4U1X8aFoxT+09w
f1ZF7Hl/oxK0rcyk4yIR5g5XSzr6+LduhafOElaZK4X6tIPUXI2QzNnv8Riz9sv0JbGLzYw22Otg
Nbn/s8kqxwPAhIsmw9MTAi8Ct8Ce9La90ipcSs4AvKhdkddSdJGTkwnjv0+78wQ6a2tTpIHxWjna
V4kuBcH+R5c5YW7P/KCUb5EiPHYsYutpccOT62+Zq4FVwOrmhQU0jVUIlQIpu5uAU+sijCekHWmB
y5q3lET1NeF1xjxXH5pdhbAM9vfmqWkMmedHel0knIuFlOAlQ4yiU+nGt+6SblyKqyOHgjYB3Twx
+Tr1WZ/IOlTQOLwl1fJKBZ3M2kW/ujAoGwuuPEkulrd+dHOKGivH6WFSgO8UEpDFSV5dt6NQECF5
ZKv3dzgkc5+L1gBcwRr6Qsn7LFuNFPlUNViSTCVtOYjnW2psl9Cr9VCaZzDGcjfRmJLdc6cPk1vd
bfRCRjW8KQJxhp3ha+cX6JJsPSEK/ZpejmDi7IiCp/o7UL04kcyxQfX0CHKo4e7RG9r8MUg/zYT8
edzp4wIGWLYex3lBohsO11Ux7yXkDTWDuNwbIn1vZ8mL7RUDSI3bgY+s9iBUZ0o+NeJae/KraUEh
SDV2XqS7WINKSLq3CtPMbzYcjg/JRyHn1sIYWk+JpGJHsh5BWZKCyegWQpEZgL+7r/H++d/QKpwV
0wov0GIoz5vi1M1LjC5cZwe1g3goeFnUn7kwKpncvL4eUAboXl469yUmKwjiVZ0od/gQWqgl3yiY
rgOXeKq85xQF/CMy9ay0cIq8ooSYroyDbBGPMyBKgOSEBC1hmdqM+Ij2hIP+uwfwQwVlqh0OR5Jz
l+hpv9ZRz7F2sEiEst1tJR+Uo/4hLTWWaWqcCBXy8kD127teqD1SPfq8eIZ3g42FbINq7vmkGIa2
YJa9XvSh5UPombdocz3DPXli17Ri0vE2zZZtIH55pyzwBRExbC63XeIODv+GhUAls53PivKzNUE+
OT0m16SvT+0enPzOwNjE9ZRzfsi1YeT1dmVXI/4DhlOg6h+/3JWHuS8tBvVBhVquQ+8LlC+JixL0
Ydvx/B8hgQ+z1XOuzpHgYOGtDj0SX5olqHN3KatayeH+alZ1AgeMuQsD6YWxw++612liAmynputZ
VCEeLfI2CHr+hAdwosXkoUpcxos4rFfD5mkVLQtYWFWOvkFZh5o1TzQUtl0NFZfyL7XYG8eQ3fc0
/FKCiCj+ZoNJaOSY6G5a0lhBmcJrbsApOw2mM4CUJkNmHBUe0TdXkdhrlTdtZ/o6XO54blrmJjVp
lqw6EedGIggL0S5JvESOTdXt55/7YrVYHtGM+7YPSKmxnR7oOFnK2EVZFpS0sn6di14UHyx8wyIk
g9mmtLucybOhIzM5WQxzUxQL5B9aFQGfAmBaVHExysIISNG82GpRD3ahf2Egkgrlca3y5aws0QMS
YCcWcWi56NysWwbTMxTQ4kZ/RC9F46FXQzXJ5oooYgsWBqi/Ixrkc7vGiXEVgazRU4YytwzRbiOj
CZ6hO7PgEH2i+r0Z2gXF+coAStdFET2ipTuAE82fapx4qE9zyTVn/1E2P4z4u3l9zBcCLHF4aT/2
jrzN+ACLAsThMfGJck1XaY09AG4SXiVSSRU9st+JnWKjovK1QKH8rkeR7QjujVJjgomZYR6Ri+D8
CtPb+cbvQxOjRqHpY/xF7uCA6WdmtibtWWTDayYzOJb92ccnag0jePLMUfYU5OceLNtG6HNnwG6g
pGmX+vQFNSNtyw40kXZBVzSyOATcajR6a4+kKRezUfc3SkIQwg8DbReiSKK2JsCd5unsru55+s71
kdgbx3kUm2trcXPilgRLdfuYBOnkxWzqmWhBp/jkAhmCW+r/IKoW+u2xT9xgAfdy1cTNdM2t2fak
/yT7euHMhtVs+YH4R9L69JYZp7nfpHRIijf5DDD/BlSM5Qt5ZJ1KKdzYFwMo0EGaqQRJmb3o5/vN
SaO6vwUA5cluN5arIL4wX4mOJyySsLW9q+5aaV0VCeXJuA8CCG6f984dzbV48lFhmVsCxpcnSZp/
rqc6rCAUpUPiz1FK59iF+9SRFzYoaEQ35+wn/Lh8DI5E8JQx/mOCRtub+hNBOQ9ZSuAmXlK62X01
cN1ia9QQYvs5HyqoPK8VMCkZS2DShmqzn2+JDfyy9/wrvXqRzJv5pt+VecxH9Tu8/Tom6MONtPWP
PfmM7VKaTYdZbJ81g/l/NsL0W6JZHLoa1UDF5jvHxkDnm2qOPAeN7qxZFQZz5SX766TCa7spI41Q
beVVhc1n+8Ecn59l3Hy2pjyPGZEDXsRC6TXsNELv3x2yQIX6P0Ypc4GAbEF9TB0ikZRDsuSW/5qC
EK524BpX6ns2r8C8CFahABterkxsTHm0W+hD/jh0k6ciuN1AAzofCEY7pdZ6kHNbxvn0j6NzvUSO
dJh7y3ByIKDynJjIlGG9aNaUmmwXrIszBq3EpjISycTA0XEa7JNM4qmcGUTpekQJYOo5Ac/4grOB
UZ19kZcWTeEdNGEud47Fij3Dtv0W6G/EkH3BOWIOa0LMUvHgNxUh6N2oh9F27FtKv7llWQu/D6Eu
sTXeOvfvOWNVcM8488kpY8vlQ2mun7/yu40TNsFmuUjhMELiWxv7SCt29Lh2I5AUVegkl7iozvl7
cShXNIQuQ142H2JXcnDb+graOAqk1mWhSjjBORlu2hq1JSXYCajLXEJOg9sW0QMySNEGquNapGKI
YXnUaK1BIe/BHFNbanZl/bAwmK98MD4VY0XbFsj8vPr1yGV6Bd7Ye41y06EgS9/0ipArXFtCDcJ3
e6S1C1PHwXDkvxFPKd8aw0x6Ke5eKZlxdlpiAKsxXk0B3iUBjcj1gCn1+MPdHrutWviIUyWNmn5K
dGDi8sTBNaDkk3fbuJbY3KCEao12/qfWPZ5x199Cv7yfATvXuDKG5xHuCDFYg+Mib8ARbk/UEuQ/
xT4zGv64DxwaHlQ9WaMmaxIUqsNyUyOpLvUgYSxGvG9zfkMPgkroyoNH1VgWmYjWhqecgFuVyvKg
K0Qy4ZScAJarARz6dJ/8hp+7KR4lnu0gxMw5RCyafHH7QbX6otZtd+D4cQxCd/PvcvDblVg1JvaG
3OXppFhSmep6U5i3lbD1k/MFhLeeil6p9eme1d4qALVfDMva1XGz0mI/hR/42xAlXTBS65PPYyeZ
KJ3k+a8vuWmaQYls9qlNSO6C9sa3p5IwcmHU9hc+FNPXNJ5ZlkQ09gSRi/GusphzGeoKUhLJXTkA
fCW2e0+BwksY0bP8tk5Ki/Dle2iGhMJ/afDih1IzswD4f73SpL3S4w2ASSA6xxXHUlVTU1WEh9jz
0oscs8cAnftExFWX5HwMK7mS6skFKLvS7/jrbI/DOP06BnkuPoIAv6RKQXerTfDLozgvUAlDaqxA
e82EgMDr3kCDXpnlrX/+z/BSOPw+/cQt6/3Iv5VnN2Sj9jueLcTPRo2RRthJgnC+SWzKyvkvDLja
FqD2VixxUzPIGlVC5MaCu2LYmypSZAJz3vrTYlqr2qYRX28iPf7p4u8/cSGf20JBqQuwcqylmkc5
xh8w/5AggFskaLXEnV8NzCC0k0bdld8LYiNVq/3lv/B7X5C4j7IsIwLtCuLwZemr8d/MNIJ/iumI
whKqfWddec849BfNYNPV5XfgnRx41QsoANpobi2NFEFtnt7onXUDGeYurv/SANbka4FJS/H5uuPR
BlhSdtLXB7ZCfIbY4GqzO3biHjeAXJa9l2l0Jdj2HkR+xTwQxIAYf4qs8kT2FEn90Aqo8+YaN7Kz
fDSF2CODjlFmHg4SklVuUp2ZfOcbNAuRwfziSo9C1kAPBJQ314PCsWb9AfCnOLQ8/FtLedjdodYv
RcWC232UirMCStXbFr6jYcEYjwuy1eh7B4CeaZOeILGRGKszojg2p2AOF9gOAQlHo/Qiu8AHJBQu
bY9HGxuMwt0KGkxaQPCIo7+yEIQZseIB/rZL32SrevUvMlDAY087umXYj/Yn6KdwpolRASajn2EJ
SOpVynWWgPNG4b6d2KC0vMfa04LT+ks+K5pGtNrXA9MUCJ9BUcPvtIz03p4mBK9+jj3EtA3+NhXW
QAaR6MP4OrM0r/vmSawzt8w1R71x4LBojsEAEpR4F8qkt9cKAIW06Q4aqbAaZ9jr5B2DhiXwolPG
GVh9csb011MKf2QxZ77QmbgcememniAQWmD/F9GGNUpvX76TigIYYWtpNH3CEC23s9EojK3HnaBK
qVYHAn1DJiQ4v67QWDzulO7FTcpZC7VDScymp1f0bwqJiI7fk7Vw8UmkXVC6DgJytR+Sze0q0qCy
YELSDFMqiycd1g5BM5I5cAOUjRVgGexaryoEz2RRkF6VetGEyZq46UA1y4XgZAoVbWFrRYX4wm/I
ykpAzhJbG6LceOKKBBTN4e+q2JP8rRs2y6b35wVCr2Z2VYtKE3z80UetJ/wvvUdyyZR7y0X1pwPO
HI98SlZw4l14Iv2psu9HzBT7HptbwyBXa8XoNnzKclAyidMX/BMz7FA2oB8tw08WoSE9GQMRKqjb
bcBgpAmlHKD6GUK1JFkslLP1C5DIc0GqZc/FeQJHOxBSUfW4Womgf6ydJhMz2kouzLjwdEm1bj9j
kApzXpEbjF3gmCpou5iz3a8bW7mJRq0PXAsE6jMm3BGbCPZaz6iQgS49tbTy+bSeFzrJxjViKA2/
U/xrQEtZP/RTPgbsmEDvAuu3HbnyZBjgRQ+Wy6p1Xc2e5nI+Dvi3QQ8yFLaE6RUrNcqzUl7Y4EHj
iidUvlTmAfzwwT+BgcqcE9EqsLOauN8o4TynE53ObXFUdDQzeq1fhQNVsKOs6UpDQ1rAMoWv1h7d
d4YT8nVcxI+2haSKlZI9NHi8e4wlXYS+1CI6S9OhfGkQRlHPvR4GTtZl8r3+U3SU/0DCPvBn+5/w
2o2yoAX8Ru5nyJa3O/vkGc01Oan3sEel6I3PeIVOD1pie8y+i7Z2wtQjE+GkUwJzLIELo7E1S9R+
uZ2UfQFnPBuMVS/JVNqm/U27fxkbbkEPq6Y11r4ZBYkgX7YidamdxxNeUrDITuaCK9tPYMRskovZ
FoyDTANaHBrsdU/T/8gb7l/zQCuE+M33eGeVz9xNFS5vTc9DeyEl4Xe+xxaK2Y2yUNaN/yFJtitn
DwRxzYoomdC3gKblm5bE6c/juvt5YXXx36JFun9/RPxKOpELL/Ed7cRd2Ge9JEFXHBbVZykvWwxp
C3BciG4etx7ssRfeL/Fz0sNHaS1J6sFTnY/DD/jgrTM06m/4Azuiq2KHmDNxKzOFmVjyWnkrIjX0
HkGRKfWcJNMEHm7F248/d2fgzNefVQoWLDJlcVyXPbegTI5HZztSVojjfBcZ78pya5H9RdZxhLMv
6cpBV8wJgZLC3NGtTCWCFdYsE+08b5L/MpRxs4q7U9EUuze9ThHqNI1X4KZzxFiJQEcc1vyLhYz/
ggewAzxQmVZKWCSbSdyFP0+ysETOA1hl/H3Ljt0zbs8Z98y26B+xFRtjSD0eDto3DJucTT3ursgj
lpqbRb9qO6X97d/bFuQMZA2oqwnieC6tiYRytao8SGqgzAyDwWzx6/8Ag3mS7of/cy3WlI2lXPeh
ULm6dHx++FMMl/dJ46yNZDQ20Q+/8mshLnXucAMI0Z4AHlfmIFI/NbTcTNQnVw+18AywteIyQmDA
8Im/zH7wuxUnclG2c8CmuLGT/Jhs7SO+0Mp4ydyhSL79zTQ/IfUQk3lPI/Bqkv9BaV/8okX9JcEg
hMS7vGKwrRBzW8D70NkEhHsFZlhD5B8E7bzqiwlTSk+6+SNAEnLBQXJe/VrgoDRWlfqa/MnENYFr
6mFPkfcMIMg1AYdXYfElgDXhbzbcIF3iHhuOdgQCppvXVttyVywWzWqlHqcl1NgZOgUDCXm7hJ36
M7aylQ49DCQKN/NV5dq5q4Fvk/ksA286ldRoT8wiUSEBEba9VDfkYfXq+CujWFj7iL8sT5cdG2qF
h+OK6vIelgZvCjUVyCRk3s73vqBQ2CrZ4a14zidsIqt7AP3U8W5k1jAf2AnsSyKZHVtgH2nCKAaj
rSfNn8eoMOLaKXijdue7odh3d/uW+0oiHEsw1HCUCjUg0FpNlAvizGXpIcYW3mAQ3VEA77fq3/bS
eiWSbX0KU4GDEIEQK44hFxEpVCzQeJ1yRb3TeEGBYuEyGAsWkxH54nSwc3sj/2hXpzlG1LSVC3nx
My0MDTbLdoyFjnO+o1HyH6eR3kKtcEN5yun7G9iLcdyBRSITy644xDhkeK5RGqJnyFdr9WPSvJDL
XfCVzq5hBnBOkCAddGoklN/3TPj0u438b2/AVjqQTwyGC1J2qs3Klp0Ji32vqTRjGgLcnWfHVbsS
QI2+3qvG4YszqOVvYoX7g8UkyLLGhkimuLeKZhufp37qzk+9B5UIqHwF44FStMBHyZnKsf2qD5gC
p18anJrEsevC54QOJ1t7u8XWrQQKwuisNo6nUUwtk65mVpp7X2+Va59dlQJoUVFKNt1ONTzmgwUx
2PxdcYr03HWvqb8fiArZc/rMu/oElbo8LTnN73cUPFMFoq2jkAORi9edfPzu05DT2nRgAYrPrIR4
3RmWZPIfbC8moRjIW9oh0YrA3q1XImmv9KjX3x87VpCqHH9WdhCsIcMhsdwMpBySPcEIY5Q5C3J/
DiQegpYh200VXTSQToBfklMjdvuXAnPsZbVpa7UxB1Hn8RgbHtpsfX7YIVQosSkd/fU18QOqtBJ6
HInrbRHPEwwocn55S4HE9xlQ+Zj957GKCCwn1zyjCOWVvXsI2ZbHdwspqK/34vfjgKSEhxfpQdwB
LuE0kdx2oBV0URfbk3YhtcVep+ELDSgzrPmyVfQ/j7GQ7NPjqFPx9SJ7bKDPyl27djRHnn+QBf+f
Nkzt4RzVHfVNfDh4FNFuFqA50Ka2asiF+3M7fGZE0JMyjU0a5TcNKlMH7wvgQKvC6q/09ZyBOCnc
CpiLfPNTFzxDuHYywh0WfzYR7JmYzmHium2QJssDR4yQUb5wM7i7xtUUymxwN2aDhf/9z9px/KyM
yAj0/cZXEX7OnUlfhCqNfHWnQCi/bRcjY6N10yjcWn1H3v3IuhqqA2CdXwjiRJwBir2pP7loi7lN
7hPCigaM9159fOhLDP3Qhcvqt+jhcfud8TAxvZuF0VuPEgl5nARUsiFlj0c/s0srfI8sXWkGBpxt
vHupdg5LBNVsskMS/V3VlbfBU7dmofEpp94Eqb/vxcr/Yzwb1IPxgOfynvcQwE9JmGdXsnhi723g
UAjEk2pOF5BuNAIYPY1W2T/MkIYXB6+Whls5yA4fwskTZbFGj0CzDvyX+BlrvUHsLrdFH1bzZlzx
m/G2D3zPdBbMubjnYyU9wUOUOusScPPiWQiPIKeRuiH2SwO7aXOQbaL3o7/iG3k3Y4amiAqoqC/l
UKjdw/daPK55UuqQsHVxjZgKxMxLUSUWjSJKCoPlRec2uG0jAKBn7Pl1hAz2PQvDtI/BhC5iGE8l
zeJIvu4kSWWFeVmvuBaky4qn+iP8x3Q6lDq4UWsYSk6SwogwOpQXl6t5oS1gtmK1J7lblZWs3cvT
ahK4yJWVC+yfS4kN5un5Vs4XB8OK5JANC4dRdUxYgztmhWLPnFvMRG6M+D7QccaXO/MIqgNrt80t
9GNVjU9zi9oSqJrFNbwWKwdLDq27HGl0nV6yTw5PR4hzvWvpvn2BrwhOHlKRK5lrDbxnfBdeEjsZ
6alJIGjDZwcAtP0Rs/KGcHhtknG4oMBK6YUMUlZQx6LITcIHZxbeX1raWV5yhh+PcGDABkifSG4b
rjJSg/O5M/Y+BgI+vqidace3zJG49kFx3cVMCqJQVBLUGjwc/K+KfLbUS3eKHG45CjiYZzz6mVAx
ryJd00zedmxmqbd2sNX5qU4gCzLvhmnstpTRctdjU9ccZ4uE1YJJP7g+iB+W6EM/4JI9JQw+z2Tt
VdnsajEhQy2zQV1/S8wPWLzOfuSPGjLguK+ESHPngkOicQrJlQWdG77qsWWgPLtA+oOITn+w/afy
WitB4SCdf1CAbO7kjB7miwy5WSZGLptSA0p7ZrSh69tek7ggyAKf0H4UPYNfSgxzYdpaB4J1Egls
T7jc1WPo3RsZedSTUYsgtw9Xwl/1vpH9DgvgMhy17qSQAton76OMagjd440nDCz3scix7hHCOSsJ
utaEjv6kYqRRYfTPKoEVGsZBNCkxNYSale9YOFIYMqUQZucpyMJQ8FD1TBo6MNQbWtz+EwJu2vo2
baydR+vS1Bjg8IjhK7XJrwMt0dw7wu8qLqpOaRN6B5e9rlydrok4j54SG+5qBmXIAfVNOMxM9fMs
wzMGIye5cDU5jK1c+ENhskh51qt/sDLVI5J+EO5y3Hjka/igMkrI9J/BfoTTPzI63bpdiaQ72hb6
4C2ukIb/kMprR8OYnY8iejD/icZY2vQGScaM2nQepMqHktU9RG7nJABc/KFmESAye0WzWZW8a65t
DBG3uOnyoaFLYV2pVBCgxbCKuBxviZ1bbFDkH9ka0JAdPVlzcuHPQmMHTrH4lqpZelgnyip+F1cw
2/xGs6hq40w+Fpvwwb0tsoRfCM5rGQGwfe5CYGTavUng/GXZpXrloGSJMeV9aCbwDiFAkMPigmQ2
e8D5NcwVBCWJIupTyYr7nZkrY42gqQZPQdDt19VUatzq9DQILwLdZ2dqgOWEcKGiu1QBq7lK08qi
gU/stcM19+VNQNWGXt1gm0ecc82cmvWsG3MgmCflWjTjxotxpBVIOh9tBFmP5rgifI0FYHH9XUtO
j/rv0T1bXcqfHGedmquoNa5zetoTQM/DjOUzpqSnYvpBL4LYjNtfrLgSyDK8TN9Vj8fta2dX88yD
ZQDDHyeNzPIV104Ds3JAE8R4I14AYOwJB9z7g1ZACoyO6k6NI9ecZNiHz9HDyBfUn2f5UjQhhCeN
L7ZMzaOw8vsW9zz7mpDV0uUXaWTs/SseRgVD8uhHt0Shc5pePuQIlsAwcWDK22MTsOZySdy7f/sx
OAJfRl7F7OkRL/w38f6GnzYL2vNP0leS57MbomfTRHPW52c0lngYwHCmD/Jgpzc8zByjcX4A1Eit
CrOSrTe9i6cTfy+Faa932FaurmAI9uDVWSgC97TomKy+qI3jiPH7BRNRkcgMkAIM3NShfc6KFr/g
z7nrrknstHvehycwwmdnfyrIgMKRe8Du8z1ahqfrriYdpWaBhizLabjsvm0HiMNTEHRT8EGrlyLX
geMx4l6KWqhCxl7VB8dbCABMyvalHv5SpJqS+SG3B23TbB1XTKY+rHKNNSdXT7qdc7QhcVVCpdpp
o/FJtSvCyMJ/VCPnT+DKEsyvF4G5KC3u1L5qj42KsvZRvgfKi6r7vWrB6RDMUx5482h4MsvvEV74
71ND3pOpRB1ej1CQgGh7UCx15v8gB7MAZncW2cubrBxoOjeKyPtf0khwPzCjV0qD4p0+y2aqULy7
qzi/dnjr65QTug7o4MRbJoHpsA/phrNjt/EpmEeL7Fgap5c16j0TFxkcwwW/V/vCMPsP99Wl1KRs
AgxJxkYksxa2UTIFUQ1GJp/cu0wCLPDYWgdAiNWKjP9VlM1KExYCn55xgM4/aixRTjStPJKUjj7F
R3vZKcMbVY59qkpKK7LkuevrY+R+xmbhFEfI+Ho9UgqzsLIfCH8JBJyv0qJwY86veNOPusf+twAG
0mYvmn6Q9c4TDezTHhtkqP744DCeWX6MKTWmw0BlgEeAFim4jLJni8Kv2n/BlxWejXlBiC5/N0KI
qqpV5rvc5gfIFH3d9TQCbR2BjyN8Ys58AEO3WLhgTmz7+ZIEoSNUaF0/qRn9eMBKE5OafMPfamaM
YKvK4DKMWEUOlROVDT12hlcN05cOCyUHElPOqcTNxO5vb6L7HV5Rzr6nfkov5yJnJI3AR+Z2AniC
Uz9B9FPz+LO9OanDpbdOAzxP179f91/T45v05Z7w1A6cYJsw7yYk/DcBeqOIDBYOQ0BJavVkcRFR
nkTnSJ6EcqxM9VuLV9D6LbU8v7mAVSttCDvbsw8IY0TwGw6iX6unwqUL4mTQBPON3nPXLjYG40pV
zsJ7EvEy4kTlGRs30HDm+YcuwbhDwVNxWKiCesZzmSf/xJny5yvltq2nsRGWsya/pqIW5PZxep8y
G4mgeV3+5feU6HFY1WlOII/5pIvHLO/CoZEKHKb5+Yo7mp/iCIUz+pUMgkODc12xM1vsVRueUsws
4YrFxD13bxGonS7kBQrk75Zs5wcsZIHg1fst4tn8XfF8R9aihumC/B88i2qR22Ew5+Q8v60FlJsP
2cgwFB+n4NYHUAxrUPQHxU4/TjGgwMcsEToIcvPt3QtG2IbTGlAsyeleJrP+swFjlXqVs2nnA2TM
TRLseiscfd2yDIdBFjPeaedz2aiw4ODers6Lqy1Q9pZlRni6EZ6CaBBfJAFH3hklzaCoHZn8X3E5
41jTBi8V9FpPPMrFrA5QVmH9bcaFqeiZxaqYekmZ/DBo6Jfua4oZkSRsJCPfzecQmc8bleRj4adw
VkHC1N8PFRgC0/9DxKmd5n21Jj50tUjPYxkduqzG8hROE4k6yw2ESqMqu+FD7R6IWS0poTr37FvW
tOB/Fhj8PK7wzLNOYlPG2aROf8H3wcL+m+CJ+ff7NAIGnwVoxBQVzCfY65exMic6rLQt/j0A97i9
Hus9loHZxKk35lLPEObwcoTGUyX/O7k6rwPH0z5FCJEJijP5yjkD01ZdsnkKPojWfVlcGoOPCMdc
phnDdShvhCK+tXljfxqJ54YuHiRaNjKpsyNTu1taGRdZrsXaVu+Zyfd77HKxGYQAVBnq0ssQaUGK
YcPWEMlYNPI+lw/ziZnnPq1r8LqFF8c9ptnTogyML93IN8SAiFAcsAWxgW1OURNNNQFEW29UjQ+z
dlIM0LHoWqctpHo2HbVKRyuw3c6tG7HXmvVtTAK2gIC5UVgAaTsTtEf69BGCVMpgsPoa82popS8A
8C7hS81ER9kcIBqdNbnkZchjnMBHNyS4E9wsOs30zs+b6Nv9UApxC/i90C8SDAa5l4cse+/xJFjg
s/Mj58uhfUxwFbcVL+dLOlgrKMYkHwJ5UXg4zWRjpEzhxq7HeaGItLt98j1rzNFtT/8qcTmWvhyW
eDrr/W6+2QJdENhAh4Vm1tFIEMuP6P+yUIN5Pj2SK/q5w4EwDfbICP7QSkxGmv6pLJ4ViHzPE9fa
o2CQTMTC7YlznolbpFoUXjIhu7Sz3I3wMD3qkHjPDsnneoa3O5qOKhFAsReh34mrV6d374jETiwW
B7Nr3X5ZqwyUaK851S0GEX6cd+DeMBAJV9trf+6/XBsrQCJbRfDFRo21ARPG3DYNsBjZz3XV3pJJ
QTvOXwOVgXehiby+PdOjqW5qano77qN8pXg3KLwsfgQadfBWVvGsQpOLyMYuo0BiON1es9+FRVB4
yqCKPA4TRvtYhi1WJUiSGd9eYjpVw1az5bGPHMmDbqP0DZJ0sZsbUhqIsZKq3Q0VHx33LFKyM3a2
eKxuCfoW1TFfcKMJcm1MWG1g3dg5Rwh4dYWvQkJXh3mh5ep3qB2Vbj6XVATpH27rd/KpY5B6BW/C
nsEAQSba15DrqKGiPeBxuZvUhU9+r6FefUHONjpWiz6m4ulwZbi2KQB3yhogCtVJV9PFP/wBg/bz
v/TbWUhGiewDaD7TG/YWoddtabHAmvK2N2Bp3cjcetE/OjQaxHkJT3A3pDiU19ynEAYs/ejjxwh4
FoREXE9BcpDHqQwnnlgeTt+AsWz/2KYjcgjA7udEfmom4NROFP8D+GiShEhIf9eXivVChQzHkoO7
bj5xcvhKqa++CNfOQeSoazQjc4+eFV2tSEjRe9jXOqYdzVVCgod2y8jRdUw5JhbspTA9Usgfy4ux
IwWVd6sYvRp8EnlcoVzMhq1XLDXcuPhJrc/+6PwERQiMfT88SCmOeTBmw6MN7vbAYHlIl1RUeRsg
QhHQxTQ33FaJWYNthL2vUERMclqwDY3s35EeiOK0Gu3Ojm2D2peKJKUSdB90xfQxrk+AdXY0Wcp+
QYtSjaUkofxhHVGegx/C2wpUP2ECrsUG344VbJPw0Mh9FVph7Wl39m2tGsc5BjvQIfbZNaq7H/Lb
ZA96kNIZ8tHZYsydUR3H/Ha2Sx7gUBw458POsG7kkO0kRJDnImSlZlv3dS2+giqdk+uvNm0/pky8
R2xV5k6yI4qhQivyJMZrOGvmtB7InPgOi+flPvKn9wMYzvv/V7aKV33R+sL6x3dASlf+WS7gx6CY
0m4fQwMhnYv0B2WCRxetlUAl8WTM4dibgMbYkDvMsysium+iOl9gbzmvJlVsWH5nJX2vntLuGFcX
b01zyJC/vnjZECosxtoiu+HACuVgtuYHh6Sosdb6IdOCmYQGI9W48+a4eYsIothl6VJo7ik8Nlym
r3e7Z7Y1ehirlP/NK6IVWBrI1wqj59GjXEjzE7k+1HzmHLdC/dMuVvC69G/FyiBlYlw8dJeqYHPo
St6BMEgv42tuKdWOF/02g7PwImVUN7z18tqw3ei72yqhsNCS0oFzTmagBV4T5XurT6/C8WGzPnj9
Wh+g7VSu8KB7iCMVw5AOxMjEnYxBmreOtidBNvLntEETJXQUlBoC8qRPgFwMtu7RzOm9ilSYBcZf
gk4Swqn02IELj8H/kO4VVFnhhmT5emps2sRZvjnwgnKMv1j7KvzmSP15+Q5iXDrjMBu8dbYQL4eV
qjllQruGIxe9OWmM2eIUAAnQ3hS6fS9RGg9bjeAxfBZr6HWzMWE4ZiRqhxKlAALZmYygRT6M0g5e
+q2rmBOxIP2RtYNkztZINW36Z7umHoC8wlJgbKZqmvOER9iTn7Qzkg7v7ktgGVf8hVtImyH/mMQI
uGhZ60SdmhKjWtqxtDY9+0P/u04CPGOy29pFsMBn68RsJpX3trdEXYI1fhnFo6YSMZn8DcV5PhaH
I4r03f0ApJfSNLB1vlJLvGcXmOBOnxk3+a7siiwTJHgObmGfpQfYbe9UMN1uLJPxuLoOB4Y6rk/h
lx2ZOoZaJrr+NxSf5+wwI8cbEUMbseN/kn0nNzovNSH8RwZHQkpnJ/uvNNPqIigm2bkG//Mbt2K+
J5hcQ8I/wFl6+Im2FqBDQ6l+Qzp77nKy0NnmyTBOR5nabKBx1AcW8EjL+G2s2oK7QvpKvqKQ1gaC
Oo/PQh8RqKak7+Zqtr4pL8j04WS2xu+BxgF2UyhQzoAD7V+8X9HIXIGCMpaE/v0OXdGSmRgnAsSE
nJ7Bgaz5UHxX//9OPSH57qdWyuqYuGvyZH9Vq7yJCnk71mDu8tTYA84sBPqHjuQFZ3x+x80HdLOb
cagp1AhqCNc2PJZElPAHEDJIOmzq3RhiDgW6VTkS/opi9+zzfaBbxL5wbt0DeCVEjO27t0W7EEdr
Hy0NGn2RAcHLT6YfznT/dPcnRfH6MIa9N7oWHNZc0T1Oe73BYUntm5/sJ7gwpc/TG86UNZ7Y/QlD
Mq6yG+0hdb57sJZiWovFlCmI0/1Jwr7D7azKjQEICkyeSPwySnB6gYY+MXe2++vabORJsAl6fiS5
ilAyBJ0vdhk+qu24IuJFHfCtn4BNzfJOAXSIHSkEN2dAaNhN0b5g7iDB2E4amghkvxJnXPlRKIYd
MLI+MamyqbruY+Srj6DN7xobuoD2bkRhTzBRPwsVX9NSsvdm+QM8CAwUCYWqGhu9DeEFxoYK0a9V
OJ8BxFJ/OkHMJJOamUPZiTXE/Q6m9D4Z8x1CAhLbyydwM3siAbxS1yy7zIsGGqVyzdm+Z7iJdZk2
iC5+U3CelF5/TxECFUZDhMh4zzrV6tdfK66G8ZD0TZYlZ8pGif8g0RCHumfx5XrXOFaAAmKHyC6K
qtlfdTQdpN3MrRpsdP99OG//izwv7B+vAv9c3nZU6en5papJWyJOd4eU3CIyOELysXzxP2FgFqv/
M4O7+cAzLwB6obWy4iA5BEMCch6/DtDPpDDqwmlCqWHyR+XV+zW8bfOzfpeLbeagJKa5Z/52nGbK
6OYnJOjAnhuAaYlbpHovovusXG4hNb2dC4k4W/kByPRnpaRbt5qkDZUJjEiILEFkcuYeM8pwAmMG
UjT3pALYEw1jnP9mjyjO6Gj3Zf4I5pvFwG9RopXWMPkMsWqbwfJSG61jWuERxQLA/YUD+9CrtqMc
s20RtlNB7twh9r86QWVx065LY4W/WJak7JV2/QttTr6EQ5ie9Ig9aNXvgSQqcYaOjlAVjPONG1UN
2GzzzqbVIIfvKPQo+qlKdGELM41noCX6pA8V6ZSX9qspynQln6zZe3BAfLK0B1zxVK1VOgvst8dd
Ev2Tmhj3uYmBnVkVX1FeeENnCFOOVoopvKc6ezAnxKxW/1JbqHS0/Y45C8LthJOTahgricdFFW61
hk8AIxvTLymfyoX9ShmQWxDqhytupeazSlQ/mUcaVA2yZsrlQlIleQ9XQdf5vWjC+HcHkFWFksuI
tQneW05x+CIzZK+jWUQxW8uYNjGD86GmTDKb4VmCCqQ9cIe1ReIy+6zwXyrAvwQg7S1p2QFq59sp
HemBoRe8tvM29zGINPEvc2M9DoX0zrqWIrHJcnBLhIJ4TXg+SLwxGNinwsaXVVEiyjiVXjrH8vdW
aVURLWtwe7PGzoNbmJcnAK6RdkxzYtwpu15Nng5Co1vthKvwownWg898JxhlHJHqH8YvSuGtTVA6
t6gHPxTrUSwLIh5PR0LfbChbK10dki3S3DlQufNWPQv3OFjmak2bHSmrB41e2gOW0sNgwNaOu4TD
frRq9DRwOmFdilN+LXWlLyMVxC32/5EwyBkwxJ/u+gBW9qeRwyGO6yTRmt6+lNJDR/WwhiKJSWrY
++twNun/wuItvrQDF9gawKr23TnybGHMVL+j+Bwn9/pHt3G1VEb2ZQnWKflMXyK8HuYX+UMFdyXd
FzgynB6p2jWGTQgTuKezlxaOeh2O9YE7JSTEKUtx2qNzG9jEIg2TpZ2PCikpdjULaOJs10Qz2mtv
4T39ZaOvDlHmdLm0t1a9wDELNiyw0xVoRsNV8Mf/gQSW5pSNY9OR+P3pEd5exjazLAvYSdXRoqGb
9KAbfcdWuKbVo/MKPryz/33q4Bd4WJHLJdOUKIn0lItu3LegK34m2/qnVe0x5/c0dQ9fjOxPm33C
wrX7TutaipaXHuwxp35xO1OtDejND5hoEhWZbnIm1B71KnZ90abUoBtUG7p15eRf0eh97LddvP0l
T/FkFu21+3dB8IHPuB963ikw7HTwo8UTtDG+wzGIaryB4ZuF6jM63qiYp0ewda5x6qxRaXX07veP
DCyiSJVJdS4zC9oMTP/+m2nns3JkxMUvpxxDPQUBy/7ZkSkIQvEfSgDip2HA1uRVOUS8N7BHc5Dc
3PKmRKShfc8TabcvekN1blRBvI0bkWSc7jqGnKNmTGtC/yfL0UtBBvNKfoWVOQv+WmRqNLgQ6D7v
fK0jwZoXphzkBAe8SxQVLqx5lASo8u22/ZGyJ44UYv/GFrOZ4tz+4BwHOreQnkZlKsAoKkUgybu2
E09lalRwDSKUK99gWHCagngPFO5t3HdVfOKHftYpQoW4V1bQfvpSNVi8ZCZs+s6o9F3+XiUmCEvV
gb99q4b3CE/CZWF1qelC3qVNtzi4ueUkY8CxqQDRKpcDLICGOO6baZHTlc9TlFO/o/vozduhLMsM
fuH7f7fbGeY/zJ7eQAp+4S0mU4EHY8Kt1HNgWI+1JR6xmfBvQejl17lc4k9E/PTXHCdNddHbj3dw
nQplJGHpHpbr7cUJILNppMZBXqd19Q43yproV1CG3xuAgs6CujRC0J/9MSCAB6w13/2cUNP5SX8s
pMHYR2hIjsSx3kW1i2DVod5S8T9uEhli4gck0iv68F/6pzdolMGO2sS1yuUIzg6QxSdp3IobzaWO
QiQoQzo12UI3TSHLc27H6c/sOqzV+rgAunokU7tE5u15P+PWII52Uy9KSn3ahzh6ArNz+fJY2NzB
BGWKN+Q7X5Dyfek9RTA0WWaqOjz+0LdT9/ttwDqqpEP4j4/bsCOyNBt21pev/X544XlZkGFDheSu
YT6PSNN8RSdvaILN8CTB13sSXSsKuFP9fpXqcbbA1TunBfYLv+qzj6orH6tbZw6mB0FMlNH901Iz
g1HZ5aBSEDgDd/L2DBT9ggrw+nUcCBXxtTHbVrrriCqz/9VS5QVnhZAdcUH56lUc1fpQPWmeVRT0
U/oFSe/jMAY8+pJCxe+/nHg0SrJ7p5mMBk0/gd1/MAWg0jO2kvY6zuZ9nWua7RDqrQKsQs4LrGG3
3OoJHIugKAZLlMFoUb1SalJdENHrzUbd2qGVOyA0osdHlJ/MYu6eUmyjeVbijtuHcAwyMNimVqmN
GQ60/uIoeRYV3+FFfiq7MI8J3WBNTbD1bdfYY4oEaU3zE7ur2MhYPqxPUlGNTXxbBxatxrodO+kA
7PUiFugAlxde/7lLiE0PLCcGVjoWICteC/OaJYd94LLfypmdb35lc/ieS9YJWDvKfbcuVAPSB8tR
bxlj6zT2sCbwJvhnybjBxJephGDXoxIbjtcN9txUCnXBVNExRn2XhZ4lZjzvRcmrlOt+EkoPQk7c
zQ6g+jmAhU5RpB6oED1SCrkO2pcn9ydyrkEyM1V/TY/otafhyKv7mzp2A5G8ng04Z/FI3Z88+pIo
p3FKcw7fgQP+iWkz50wzzJT3MKMabxAWyQxCtYSBdHjHr0ow2Tjwb7WVwIWgN/zCmWL+zrKM/LbL
A3KBzEeFeH5KGh1TMHbTgeUWM9Ac2zqHn5A7FbCa4oiRq2qkZDaJaGqp5JWq4F1Jz/FInwUW/5D3
XpBRirRjttsY5QMQHJAMV15g30V77/RBNY/idGnMrzwBP+lmiZPJwsdtP5KWPmQ1PG2+9FEoaQ8R
JI0hdczoDqOrIYwBKT3O4HQ7zjLIb1ckkkU0AODJZnx+fWkEeTaXd1D1IQaL67qIzAYhMamsfwbf
/yRhgvC8LZ/OtuJQ8+D6lRIKQcMZk5/BwNn1ZSFDbGAc5W3tcp5IN3WIHj5RDjQDCLEQj14I5Qqc
y2sbORsSt41YADM8kyBLT7gN0r6VB9jFd0+icvNYSbuU5Vl2gBIfQ5+Feb4lTKmKec9FrxwiusTJ
AVv41GfnMr2hnifae7I2L5pSMt8gfXD6RnkCasow2HTosMx0TTBdAaVNZvqdBS3RIbLJ+eiVojSi
y85IaGvCrG0OlWA9NMbFt1L1pbT6LATVzIe89ntQim9Sk5/vycgg4zosW4/Xb+sE42VMTvBJCpE2
78SfzTTORfq/llIDdQVWos94NZ+4wrab/JITlvYHUG0sSIQC4dKr0MGr7fniS/71bukEZTKZAYEM
XOUteT/UAbpqPJnfjy6PrdBsn0dBncO5jcCENdU0aCAUo3kMqG5Q/o1FAnpbQu3rWmktWnQv7QBE
BlkptrzA2lKXCtcExsIaKQCEkcXz0jn61YKzNddz4ZDKiNPhh0an5fd3wyaA921R9wAce0qxRn5k
fNewb2B+uliiAKV0O0AJJWqM6EcOiy5i8GkCth1TvvtQUqcb2OrtJ5d42tcijmtyo1IQGHZws/Op
pTPjXOzMmHf7Hvt15nDTFKe02MVKVBEr4CRXq5Ig93JzvIuzD/QtnAjbOeO8YDEE42MApChGB0dp
+cGRQnpVBScTbd8haie6KSARPu1OKLOhYe058f3IlJUCVRUphNFlkHDG/ZTwvrUi1UyTpJejKjp1
mENuJWX5XSSrhiPm7UbOgu+kV16Ae/AXOXnTwNTCJ/rrLT108TAKb3AlI9HaABNha145A7IBLqDF
6Ujss7yF8TQeWkchGD83W3OehWowAJg6XCRIgc+CCTWBj4p8IdLEqnjgfEgAG2fSc9qPU14gHR55
ugFrEV3OMHVzt6rKYzWqNxHGxQQmr9gdqRKZggqQz+LRc7SN95O6/UyXrdQYp6XC2uamqJLlpwPh
6AMlr7+dFbUoNdW33lD2ZyWcK2/1tOtdVRFqorowCpudYcxOHESG/WDa0lLo+OhjdGxTiQvhMhvm
HuPDMUP9HMXiDSUf3kYkTgif7arKD0FZghzmlnhL+j+juIbvGGRIMUKYX5QEQXaEfpJZX8KWc59f
p401rAlJg0U0fwJi1c+GyDT3e42/7u4MDA4WguvS8MpYtkLlMs4eM3Bz8dY2fnyiknWrWVlOAle3
uHkYT/g7g4KBAF3l+zNlKDGjN6vQ4mmr05/jE5UJGQA59NAggonQQssQt/c/mfUGTKSF0jJwTYFp
L1cmU5kXFjmqNg6KFBUh5KGEkVUBpluma1kZnEQh8WbXCDOQvHEKyB6MnHiKQGiC0oWmXFKcEgRF
sp4QCZEk4YQEaKR8bUrTeXmYe7kzMReN9sWspP8483UJ7XrvfPDooWgKY0FuEp4Ka2bKKmNVY9zZ
AGgBn8I8UTr/ffyDlS2z34w/xlH0WxoRfzKR2uDD4kIbvUJG/PXdmuTgyrS8CYl45N3gYWPXWvh2
NAl87QvnlnrQvgSxZIX5QY2CiYUgPO4J66xYscx3Ie2GrGUtGUbcnwYcG0TT45jRM3nMkVOfwPAW
UOeuExqlbXfqasyC7bSjhCZHhz7Ob+0AacxtViSJheN+98t/gQjkCuNJZ6vRgxouPlIixWnNC6Ic
7O/dttofCSzBBgN6mFfSC6cOJvFOvQ4UMFCc7qgyqMdgJt0ZwnWayzJJ9MGX/Ub5kBDwyyL/WtR/
jFWtl69iP8G3+8RWAIrzXWLo0aO67Zbx8/y3aLKJUZmb55iLD8yRxd/6hL915OReNhX8Vn3OP5qu
NtfX6qlGc7ipGLSGWcyQfLkH+2HTRj1XKhhR+wIxYR3w8dPJZtZRVBygz+MWjD2KsaFwrajq2Bhe
rfPX1E6MphuR1CC4tLbzyV9wnme1FCEoUryZB051JQhkF08mTXwsl0G69e1CiWFXLNA347e2TH1g
UWcc8Eax2MU8UM2yb6iWwqsOEL52JFEV6k3U0mmOa+pcPTCmAEOuJ7KvipWDXzYXHaPgbjKgdPDa
aq+ifyiVnsQaC59Qkhb1Q681IhLyneRXvjMkXVJsa71A6IBuQ8EqJsz69ZlUs4R7VuNa7j42Mg1L
jXUF5xualHjbjH+5/XszDzR0AKMQZ1oclBdKuqC31oQrqYrIeEVkXVMSou7jVGL+/oOwLXmiXrDv
a/rHtBN8SKWSui6SKwjMdXnSLRtAP5Hz3U5MfbUoxgXiYPTN9YRCNfUbQjrDZhTZYP2VY3Rs16QF
HSQ3otHe/Wzs1DFkB5cXZ60K7ThaBABpNv/jyREh/TsGmL+xf5T6fcn33/uYMSlDPtdsN1n28RlO
4hsUB8DoMZZHLx7Pv4FKasRLIVJBy7jrjPbAOC3sZ0zHNw5Qp2hp/RqSJRH5uKxENTWPMsEjZY3z
Wq+gHj8YPnjbBzSNXkR0yUin3u7Y5ngkEJSRjH5rPwrS/i3YQgffiRlOPoEgt3E/vLsY0RkXpGTy
XcxOJJOxTXfk/hX7W4cOKZltcQlTomyBvjs7Sc+N8s/p9i68FRl/G6GLAaRwZtqt/uV1I/80iZkU
2z1iOAVLuX6sOvU0575rZ9Nhz0lXbOE4ghRNLoOfNuvxI3DSVQOFrNPqM9N9gcY5BdtPCCpa2iSs
6W/F/pQX8cvPqzsgP3jZJ5rfe3vE2/08YTIKs8ibHpGTONfXKs5BL7nFMBPY6eNl7f0q9WxiwZPD
W+2pJ97V70hC7gRM8DdWe8HoiW2h/ATTD0625tvo3o5p9vAwfjwmj2hRlyr2vqNTcVIvwKc2LuuN
pwe38EFXJjie0lJhGG6wUo0/zeQuKuZeA3pNmn5sMy5N8m5nJ/4r89x0Dd9T/cY2abvZ8tHN6+Ub
w3t3yRMT0Teak1c12ExQnd0Iiui+PLu+dwQqYOSjMyGl0P8ADVVIi/lnSSw3bJvyIa4C2dbR7hJa
H1ByoliiquwiFgd5FBbLx+BLWEwh2jHt2nu7/GBf06ZfKhIDTrTmJyszr9Kxtg2LmTILPLMV08eS
Ws/Oe/BLY1rckUWcST7dujTXv0xVm2v/RXMTVmox//ZlscEfuSpwMzCRuAAohfduBRgGkH8bjTT1
cr3vYQvCTj6ed1hcmpxANEZTDcL8aErvY8x5VqdK4xlzAXAGEA0JXQ9z5wXVnV+fNbv+aNm3jGsR
2qqhXzWfP6KbibOPJWnbH2z3iuzkxOmIkVqUd6dYzD+KHSJNI9+Sl+GGQGeHXX7McQKPQcqQuHLE
rQN8lgVDhoiGlu+Y0tcjekLdQ8hHBM1SZhtvmfqezzDofVtho4SzLdXcG1PYKRHUvJPbzilcm/ql
9LxBTdzBP1Lj6pZYE9Yc3As5hXX/+F2KOF7L9ZSCewFvT0qfVo86flx+CU3BWL/M+6446pf2t6a3
Slk9ZUuedj0ZYixQ3TIcsq8tvXE6OqgTfg2ZKXEev9f29F936cSEt9qtw8kC3ynr/MOn/MgvBw/9
NrNrDqdAascm2PIOJwxnoVRiEnRE9SG/sH6tw2T/Hdm4CrfnqD/eVKDnWgC0DKjvOaVLQpXTciB0
LWSoTtYzZYC70Ow6tRQdkLOKhq+6pL/pAVIh59sfQsGzuNjcr7/wOehnfdU5b71z/ndhJibma7ao
e/qLX53chYVyYfSyRL54R9DtZyqfTr45EsdhZkt1pv+UuNCucsoYr06TVvO+Wtpx1WYoz7qr15P4
I2beS3vOguO8JsKoQvMl5Hqs79FuMM9Zo8BfRbuH32CDNeCQrb34wbyhHl9XLovYvOPd6/CSpCVs
dqUOj+0/gPSKHobsuvFjv9/ibrDsAQsfsds3jR+CAiIkwsiFdI5LV1yiXFxnVbSxdFx3yCyl06uG
23aJDtEu6JW2x8xphsBygSxeiERA7HBxbhwotaPC1t+Xo4pOcaZJcDylGwJVJcz1UgXx3Q8WCsoa
QomJVQH2YaY1Hg9lB98cy75eYNp1MM+VYW8rLMlny1hmQxvsOZWBar7b1FY7ZzGGiNX+mPTNX3h9
LibV0Ya+LCbf34BeMjkwQJWK/7hT0EC8aYccMSSiDJKw0iuswSzHjRvvgU5fHXhsEzN510ZyAfAY
FJRH1ahJZTI3//NOtygpVXWglGiqk7UO2u7vPR3iksUFhU3xVG+D+pv+h54GgqA3iK3ZlYCoJ3gN
e05YzMqhDaEyHxTmJob7NaTkkXCaz4AMejpwDXK9Ra5kfh7WlJW9+y6DL8Ac+ZiaTRFhPRBIQ+LS
33YYzcivHTPZpZTH7x5wWI+Mb7QqIIXvU8RRQB1dIkHSCdIQtV4LkFFheDClD7HPhdZGKI7HlYI6
zdSwkph0w5h994Nvz3ASYPZMsNonp1pREJqdGLlb7yGT/IyTWBZS9U9nvZPnX7DFvDrgNizjzprh
zvG1B0uscWUaUetY9Pl/lcSxWu3X/heWF1yVF/zMiTySwYlNOGPnDa/ln9Gkhp3VeJIdM9NuSuSs
hUwNe4xH2FqTeFXwwomZjbc0qZGUB7Arsyz/2RksabtX24W0cB5Hi16JfuChcNd2yToAUHFGBnIy
9uv2wkqnaJwx/HbKODM6ouGnY1RQ8qCBOI6LPChICAYKeP+odKXGr+9LYf1rbI7GVV3qNMHSjCk4
xGWJJ+bWhPM1U+sBZKe/MQyJ2HDVihHxY/zCOHoOFfFbz3JwWeWCHd4nUb3TU1nKmkmWPPqGtgc+
qk3gah5Qwl1ovU7+qnd0N5yD9HKQrIoaifqHCpOJzAHMC5oczhlfxf4Xe3d3Kj6x0Ok+NleE7odP
ndz5ZmcpIuvYpMBnHf9qzjjzqC5tjIZyDO8SZXVp90FxBqhKBehA5eNVjowfoCXdNngbkPahc1PV
q0LZy6DxDF0iAskvKdpRZ6HqVqR9ZYBB76zZRx5Ynm41ct8LCP3xuhus5+6G/XoWtRI8WyuiaHy3
TaU2Ji3Iq1Mqxz03BI7wVa9s6PpFC2mputO/FPSuw8QWQLqcWWz75Ll5qp3CgxfMspo8blGmPAtd
vUdevChPFNdjtMUHadEpsmZitCvUFWyILLKh2Q4tLntdLJZkYbPpJu167A1KjsAVM3UqE4Qk9ESz
GLenVXiY2S6jeUwFuB1FptIQkMG7oWxQWOITmzAkCuHwWQ9i7cYzQD1SqkpTyMT41uyWiAMQQFGx
qfEozt1P8mWFKmC+j4tUSSVqX8OfjJliMqFFJPNbMOjUiBAva/z+KJ0HxfCXkRefhY8MmExIZIBw
IStNc0tx+7awf/q2S1VwzUO2zvk4NJhLnZ2EcF49jdnbMrXw3lRFhgdcLqF6kLMvoz8j/t1j1IYV
Dl2B2PvDaw6OeMc0axHUITXVsquZMdTwGR4FVtEivwFG9R4ASnkvdH/eJJ/tnE/Wug0IWKFYsASj
ikecWUX3i684smcsZCgdbWGFEzHil0s5A3AVjro8/jgFn0/GmMPIwdUe93b2nrrLWGdxcnRLHq+o
QKHvXwrj6K+FEIz96dTm5WbBsqnEoUbM0cGVLH9ocoAcGuGTq2da15OwcxsdCMLmF26pkud+oklW
vJ8J3uwNcDjy7pmtSn2nyOsuU1HqQcMEPl/2YSYZdC4EfeU4bNtSYBAQkyYxn8076z9DsKdZqFkt
vXWOcQqn4OiuR8818NhhHD/E0UXAb/7x4/uDhjYz4Qd79SEXIqSVKykZPcTw8RFq6cB2C6QDsw+U
hJv5IlIGW+6VVI+yHoSQGjTc+BOQOZna6eAmnoindc6z6EQKUNW8RvgwvzBBe4bAYcvOqCG4TRCB
/Id9tn7o8ztQNUrIZJcLPuoIFXyBTkXI3VhzccCp/QhaeJvR+fwnOKMhxyrLZwF7gbkFcOcGkqRE
TcfbYfNP+8VrjBKSOjcQdU9CCX7T6N3I+N9V4PtdkPUzeUa0A//8HPiQGnYqtdZCTLfFRORhCftb
PLSSgiAIrt2dyoDPGiYD1aKwDZgCYjkwT3G40YDfGF48XVGAu//I4/WPsWV6pcBE5sPcGDfl6VWR
JRzEgbktMmiBRQwe+OCbDDSHbFgNjoZ1WtE1jNla1MajB1ADyN7rv0yRwUou7OMAKTKKEWew528h
05qN1ccpayErlg+Ggd3G2JyD+XKXTCboez5T7N43gkCny8CsfiGhPnsI2ZLecHN/B55iB90byj71
q5EUzbxWyCF996XRTEESCMPXkVmENpE7LvL5pYzQVqZNmULS1NkgTnl6KYGYKn5xyh/nsAoe3lf6
E1E/rq8WZl+tr3VK8TV0wlVt94GXzaouGEl/wAGA4qOJ2zjSa1gAEK4+Bwq254muk8oRxhAOcljT
rp3jpy7q6uptNet/JVVkkuhoayqwirlV4YZ3iIM+B5ffcBrkBZ+jpu1VaK1wD97QUs3IqmKu8hFG
bOrH8PsjTaaArzVA2FrpWArm5VxjRKE49jsvwyJv/lDndhYS8LbhQtIGhkNKxJs+SG5xWE4Cjuju
ZkLcTiYHXMJCHP/ADY+lFeSMJMWQVchf0bZMOQQPX6B1RcFNqT2fyVq/R6Hr5zhYcVCK4InA2WfJ
6qcx0l3aqqyVdAOyMqnMUCvvNXua8vLDbo96ZQ4QrmITHniamx4v666oXEKd0mzLoMbZ66GJ0ydn
Zu6trQhSGbjqqJTRsn1IGXmxLXHHZb1vQHt0Ja6/TvBj4Fpuu5XttETvkvRkyhc+fzMjI0aByNdN
iz/7tcx2P1FPjOrOBhA2dvWtm6yA/E9Bbx0pEHAxx+xZpUx9ia2y+010yqrqccbAOtFwXBJiDfgQ
Q8tGA2muhcO3x2mubHNE2u80K1cznn8anhdPlmehPlVBpUKkLkQj1xibZ3lVIyGIrvyd3QtEOr/l
zQiB4f4z3Zp3H5kQD7v/iEkq0TD1jHT6AgpmDQeMMzIZMusZh/GL0xPnpppbyWZyXcEIdzjlHhxl
aAKu2spphdo56+Q18QKesIpg70R2kk93Uc84ZRXPuZbR5fYT4h5o8zSLWq0Wf7mCAor9ZGs0Edm5
RQ4yUJlYT0wA7jojr6C7VSQdJgzff5h7P3NvoFHZYw8EaQlL+Dii/ReWenSDTEPdm2CwLw73rXR3
3jEHuxLotwREpKK/cskn1nsPUTSCfYTN3M5DJSFUO51zUCCWfDblFumjL+qNESVt5r7ZN0kGoLWr
OxO+vE10sI3Y8mAPl4Pamh9sLTB3T3dxQwIC3XsBVY3TqHu3e5rwUlPV6usnu69cUzcVLMhO0NzJ
WFqsX00LD15nEWqV40zlN0x5IH15cBrAfWRr9mEi2Tpr1p2y2BCrELulJvBy25s7YuDkjfKs/Aaz
elFoaks/kqiSv6vF+A4l5ye21ulIL9rikJzKX/PmCNiy84vCn5fh1OYUSt+RsHIQlmNmz5+JwraO
InE4Ku5bZiWHO8PZGsSKc128U1DEDSY+C84Auh+CevFOCQO4qV1ZOSTc71THjOMI8r0AMgz2MGq3
NuCQBnz0JiNNcycFaP9jH+e5xaNg/sjqCamUJr1sbDZlZOCzp7lqIT4bqrRW1eNWkbDaKT070bzf
3ljkHM4SDM+PhkwlYCUboClPoONIqshrXijbpvaI5BvNRG4l0cyVzHsc1l+d9ljKVdM+QQoyxLYl
sYXmAfXShi9IIf49bwajO/Wdz/xpkni3p8saHcowJdncK1u7kdPUQJXkHHI4NQDHy8lDxfTi+O3J
J/pdPL3OKSlG4oaFB2IHg5Sj+cKsYAOcCnMCGZsNw/mxulxW0pFkQEZfXK9+yHitPzgIVMyvnCnx
v16B84i6ksxe2f2Xk3MNMp4RKl+goeANqz1v4O5Tamff6bOFf0N0+nF818TJdmug26EF1nofXdTk
njfm9JTVgcdhyOSoG0vrTrCuInDVGcnlLwyIkg6hNRGQp8iZxHbGV2KbsvDpl9tHjm9NQYqfzIwn
4wZd1Br6CicRB2IEfY+E8ZV5eLSH3heeFWzW2bDBmTDBOVRYGNylA6oVUEmQOL6ME9huKjil0kpz
LSqDWoh8GskYC1b/uusSSS0Lygbb5y7syCzmvs8ekchSGekSSG0wuXvzP7lbFBBhTTkVr8cGNlVq
eGNB0g0+2yNMaz+OSYFE+dG2dFwThyL7FaPneXR+xyBpb/tKBTdTZpxpmYVhNgCRGe9w8Ync2BzE
mU9qD+X2YOk4s4DAoiiDgj/vsWUQUXS5V0Xo3Vo6ZYgSnpTnndvCL13doTnHtNL4vskzPOHIG2D7
SEMsd+gD9ZT5xCvlDmHzZBzJVABSsKHh9L03Ozd0tSUCeNPvCe+fcQM7U1RG46twzV6TD/9iBsDI
ZnY1fLwb1UiPzq3BZdcXVxSTRQCE4K4QIVm2+r7xOJe6b2UNNnQt3E11XRNhE/nEyuJJE11pVAjW
+6YRc2KVwtFxVrkooHwhMxiRqvGwg0OZ+aYBDsvkJbKxJarbqcDGZPYHpKbKb9f/rOL90GwhVQgU
Uxj/XnJ9T2p4LX2YjAKRpgAP+CVpR8/0QsLnzVUN5Rxvnl64IOABbp+63nT/POI6ohAuL+Qj540C
3ZzN/SGjOPbCffXi9SnzU9w6/SmyXggU2Br42dQzC2sOAcCMz746PVAsho6waPBSrE15z7NbxKd8
xRJ4wDsriIbojSkaY7DOoT0Whw7IbZerlCCEsx+JOwfueOoBAJ2o1QhxwzHhHwI4LfwTWiz295+K
sstXmqR2Pcm/qHXUw8f1VuJKertNDJmsoddYZDErEipV2g+M4Aifm32IW9pRWSpiG1QFBATCl4BM
S78Fel8mE38UcGQw6IAf7y2+jAbHvMrsIXnijN/kMJZDzXfzSzGwNY0qCUTUCFcuH4ul5+LXE7MF
1zcdkZJ9/Rex2Q0UbWFc0u+Y+2ZozKslRSSxA9X9XFbTaB1MoDS6siENoR+u+OPGFc2P6fb+h3dK
MGt8raY9BhJymVSAQhe3JtIc6KOa62E0aPd1A+z7DTnYnLIGGOj+kmmyryL1ECzSNEEIDRKQdI17
BqngAzqRbCipdToBujtV0VmS10gLVViQclpZVWscnwjRWV7HeCB77Rf+GBtnthdFIb7bEC583p1l
qQVpJFUE+2O1ccPFD8uYN/LckzNTLdqdBvUHjU/S+8+rTjjM5Jo50Bdy3up3QzFMsY3K0cuc2oWB
xi/2fJVtcQhxreGcgJ/6+xRMtlGqKeMpL8rDkVAsnWaSnVrCARA4/TnQ0BkOi1vHU9RxNaFsjDkr
IxKI3AQdU2YKF+5JcTIqvxM+qzC9N71cv1srwPpd8RHNjWkjwGBnE7SkUytXZhNeLetAZYKIVBg3
El9J0RpXD5myOJZbt/3xwnbNtEDll+ExMc52IoijdNFBH6gz/DFum/lhMFF3bbq4e1ACbR6FWeZa
PNdnYWREOe1vlUv2CSCyWBwa01WNmtTg2sWIZPudx6IcYDKm04/jbUzkE3uiDdurtyuKs+p3JuMU
IZI+TtBvS3lK/JCi1bztE0PxUaoDTjZgAdp5dFnObb6fFsI60iT2gBcTv7dI/mfnI/jvBRtr3aor
uO47qsejYZnxucZeAvvuG6fQJmPtC9W4rjUsQUoRs1G+PshrdlHsQZcRuJsbDOWentqCD8PugpSX
MUohcJO8p8aH72i5tuQxhRdYCBMIbBfBzMVKpP94PVcKPTBgZPt6E4vHhqybQGPx5Hfb57iX2xBY
Frbf/0OfUEXlaMD2Hc6Hsu+AsladFMTJ/MtzdLVGoJelk59OJaGnrKnk1pw1V8RLeStKxTiJQL/8
eWyf18QVcm1TWu6nh/vxnJjGs0Xz4b4MaJH1m2S2R7EQ9C1ryueUCuPIHN7RA+YOTRX9wGUT6JGC
aPqNG3iW5U5XIQEpdInHAQX8PvqECpDcck+l9UeYK8uXtYOXCo+qFg5D+Xox9PeRfenmJwvpIVgn
IhbuDc1H06CdyexJxwaSKBH0y4cHm8rNQ5Pa8ja/PWqJ4LLFkht5j1ohlxxOsHvSAJ4hOIv6DpQG
bR6t9P58KxMht9Q0U/pgFKYJNoe/83JlBtFjJ005HzMhuB14UAPn8o6DqA2twybcR8D3oaOl+Mfn
hMSm9miN0OefmCkWxGW9DXYLq6mZu92AOb5mIsgqhcjpUOJK9tCo0GbAaeF9R1duFIt5HRtgNEyS
TN7ZnWM2j+DrVLAgAlEEJoJRPEZGSOl+XXKvLI83SDjoTZMfHKghJjlhvNcduGOYApXPHL2bNcyG
RDniyCOA8+pckAwkXnFSMW/ZmvRI2BtkVxvt87BfYScrdQhmDjiLAKjuv7iDEj7YFxReJFY/+m7U
zYbPA/UXhjTz4CQreDGftWxqm3OtS9zpUSfh9m15xu3XGXq0LAtvblgTLifz6LcaDajo2Vt2HBnF
9VprYIUBcm9u/VyjqE82OMCwa2I+++OXlvN7eTM37/lRtXCHKfu1l4ehnvLaaOGhTECVmOtLj4Ke
QL4jrHQnsIO6i7YhVB3sMJvoPJG9Ss6niK7/GBWfuK9POdNJXlccrQ0UILKpICfzcFyXdf06Lajr
a/27dkzGWrIxyv1StbcXcfwG7G40Pzfsk8VdFr5gYQto/2QfZGzmDbb3WOJq0Jrkf8AuQceqT57k
V99kxM2RzLP/3cS5onD8y7gR4qSWprep8uNLgP7l8RikI6n5MfQkjqGzioExBHR9K+h1P0h53DMI
y00LSCTZLR0hnqgjzPzeZUcAkrq6WpvkVAx3sNQzUOZ8Ijk2niuclgSV1xlyW51MGgdZczS020Vt
QJptynY+9RAtN3MeeKvQCBQSph9Oxord3Zmdoqz/hOZDBVHMRKTYaaKYfj9PEKA8WzyCNbwbQ4Y3
uQK7QMCm68+LRa0UQUhBGhaB075fNyVFHMfm6Cf4v2QI7Otss0M9jcNa2oooj+zJ9yF3XTVuL1eR
KWusn4aBERYutlyubaHeFJozjVjSWpod1sAaVEbxS3iXstRi0Jpqb1MSBTllWk/VwR9bTuX7pWVk
Cz9WpKWGtzsUESW0jS/SJf+C9VSLnZxbVskCEIwBeTpSfi5Si6mceUgKkPuh0MWQNXdzPuKMqrga
6DSoUCV428GFD+gnx2FOrMAtgN7c8xa0nMMNfmCXvXS+TOjs8ZCJGsYyRoHNXh0Kf/+05y287ok7
XfBVLrDo2dFO92GDgXcj7vZWyae92C09K1CEIFA2SbiwrsVJQqDOlAj3uMqIg7jlooRi9jdvYe8y
RTJbry4yIDnw+irpZH2tVxpmOiymtpZzKw5ayeFIhGSfBSJM+6sxAIl/htw6FOzAMaizGswxLUNB
E3n5mlgKvGe2koIun05pXNHcgdH8eO8rntFAuCoZutDSn3jpB2c2ZXyWJ04BQlUacbSWMabI1B+r
p9m/Q2NI8j+ja+v8gCCGMqxgM2AyVj+NzfKvl0i47LF7GATg8dihKHKOyNdefEhn2F87SRZ64ay2
ClNR3pljjHM8ruiwzHbYlXv5KyJQhjytRCon+TVT1lCh2cROQRmanfxqxDE6e6A2Vf2jyYCdhCrU
+C5WzRELj1KAI/eZYssVHyaZ0U6W42BDwxnoDE4NjtozYLMtPEElJ8bwRW/2ODKjFwoZrKWbLJIO
gFBKhkIaIjp/g5dUBUqSxmL3V3KLj0V2OtFfD4dWEb6Z7Tkexo+gMi/QCEHi0iAqA0bRJFj1bmie
4cFEPOFr2GH1lt1d6sPOPstK0Jv9OE9yS33hoEawRNrp5RH/jWMq7UcGqNwp4b7nzl5dbR46w0Xo
zRi7siDh/pwHpZ31Yn2sDmigFrX7qUYp0vfYh7+JYqwbu4FLcimTcdSb/XyG9UYlTcGJFfKga4qa
IoZNq0cNooCpoG6ShnNoMi6re3HDEVCLj5FWTkQ4mcmzkzgel+c4vPeTSI3ShaoQihVo7H76EV3V
+g8UBch6yZoSz1DtOydddy79Kyj7Off9ScIn77Z9TzDSwkEltjskikKxomz7lC69HMIta1oXK62n
rtctD6v+Su5braqRsNPT+r8cm905YU7KDz2kCW7C7LRGPbSHEdU58XSoOCBNA5WGzerVXpdX1E2+
ip1R8VZ2s1VXl28oAxl11R+U2ry6OzoBrLs/LCcL63Fg87WPHMwC5qE7RD0+75b3MhHq52Rb2d50
6A8c4j0d9KTaR04tvrHEdtRQin7nL2WOgLz8/aQ38+aJwPA7LRHGf/RPeb9d1kKDG0k7b6b7cKIG
QYDR0iJIh0Exixkr5noLEa8Ta4IKDbm0qNSFFxiVH8iGj7hZkUDP/FY2RYq17Ao1ZiAtdHTdc1Ek
0GvQ9fk4dTpSe+gI9Wsv/5R/9pLqc4N6S6cpTl/Kp1T9mMpIdGqOscXpnZRL6VARCgnVbiTN5Aij
c5PPdgF4BkPaSwMxRxhAbJIfZ74W59ZDI0uPQB7B9EeUqTlK0qFV3SRRKHRIlnuARUtIp9etJjEp
47lWR1maZv52JqbbHjpOtQEWWZf9hXCroL79zCMka5ykvQ9Gx3+fY0HFsTYilyH30csXgXmeY7nw
0/aciIlNNjMDUhE9JKyM2MNcB2fYMvJS9ZuDbu0lk/N/6ot7rNKEj93X838wcHxNRnsc1kdJAK4T
B9sEoUCmfRrXCuTP8ff1cDcsi7u/m/nOn78VkgXJZvbS1te/0mQHNqm7zGgd0PgjDhjEzhvYvS3t
OD63QoUi2RuYUoah0KCjJektxNvWNuyUIEtchkKqlTuaWeazMuGHJUSFknqRgoXgijGPh696Mb/W
3LIOxTqlRspSLHKCoPia0j7WnISoBp1eJ7slYg3xyDSTW5f4k++GDRuaITdjIRHpddJsSU9rUKCJ
GWNWyv6BbqNkxfMn/gRFVB3gGncGbAXMyecy1pVaK4miTroX5pjOR/TIUeNlbGewGPSyC+xtI0Y8
u+KxaAJyuVsbiG1fNRoP7J+T/w6lKbtrX6R9aZ2xpGJRY2tx0hy9Rjh50y5R6wHgDpRu7R2RgAPi
mooxP1vXk7iFqqNr5A0tmC6N1mhOgewO38oYAWLUpTcE6boYemN4nbSMQx5vmAsMj3ZzoU5+8NoW
Lh9zuVTfUxqyvo07dhllC/iZOPhpCm0hR3Ikkgd/rHsg7QC8BzJhklN5Gyg45X12grRcJqVCjYK6
hSs9YEAFIagy3kREivJ9avfEd5dyDXOFwO/qE/qDRcgrs7FJoFl5pk9zGDGfFhPVGJYfWo+rpTEW
bQk/XayjcXxsd14V/hKwDUXAh9BU+ymnGVePxzSGWnYbzKQs7fqWSgc1Tn1UfybRKQNFwAcVhkeW
MzOglg0NEA2fHOcgrZydrQ93gXxGHWdjbY3q8fRcipaxYhVWN1dEfAIg2aRu5F00Z47REPJwil2O
NNfeQK1PwSQgdsgxb9+zffW69LQ2+VrZFCATUCXGhrk+qNy0Ur5wE3m5h7zQkgHlvYXTZ+12EZ8e
ldj2bKnXScvRPeuQ5jhCe1L0kxQ+Ra1FPOwCz8hhe6sa948jU80zbP2UBogSkyQMESfgf611mbTi
J0UPYCFclhv12pdDllrwnR9BmpJfW2A67HXZjnx0u3uu4fNF8xfFFA3BMdHToI82y9cSoWtrh/Eb
o/fJdtPrUIxgCqGEdCwVrtTX4jUGO9oFVX+0mREiEf+69AkHarICWCrP3xOUdzZySvsr4yXPa6P+
UE/LYGQxRQfDv4jd6oBjTahryKeviQBoWiXRPgIoACS2yYM419OrdYSF2D64ssn6YcutwTmrebPg
iKowpolgjlN3B7f4xFVj2g0aLRSzUQu0CImYv8S+h43MJkZICf3a4n1w6oATlUTmSKj76t17GU1w
td7vI9nnYLIM9lPIFFSRq0XduTrpsZ429/lafVfQ+IQ8/QmrTDEHhtmgNXtM0XbAPDV6Ox4yIXV3
Ko9Hjf2cDCDQv2Ja2plg6MHvU06rPs9N3Y9iQK9oTke6cqAyJX/tliNUsBMPhIMhDS63Lc8+S01K
dX+dfF7l5G7iXLP2WOwUdUWpFGLL+yjOMymPxIxPdpI0IZLRemGtPNuWPOYFQa9pS96IsLH0dVJQ
CqPhwk+dSqkyEmQFTxZDbOcwAOe1rhk05TgX+R2Ue+moLv/46xT427qhonsNZdTdOqfvB6k236VR
Y2ACmPRC82YlZAS8MamygminRwNi/5AcDdWorBBNheEYarw0Zcj9gIA9t505VgqJ8vjNZCIgfkcQ
hpRy5VtTpFINbA9egg1ZFDU4VlRX0BIKaZwKnabXb25Z833YnMxCwzts6El2tSaw3wHgqRywHVlZ
6G2II6Bn42071kWMxsqzcQIFyl26timOKeRZhR47KpaZoblDTNgu7Ij8PT7GCAAMSpRt7dx4mYQw
Rx8RaMUcRYfONtcypLWCDqUYjzzAYz6MuQf+H5OYcYtSsSEa8cxKlbMj76qNow+2ELwh6keDPVVN
VpAgMjVpbvK72hPQoWMvUGozzWaWQcXS8RrIiNlpsESP9BzqAlo/ALFjXi8SX1aOflzy3sjN53DL
ApGg4Wg7QoYKEsJGio3BZKs1zXAqwYIANk8ZbmiHboGx+sARE7ebRHLG6gzE8kGdYgaAuGPwS9x4
/mVXxoaGFummx/L5pz+rWkVOKDIOumWfC7LOlsTH2o5nZ9NXvYzdbFyvZA+8QuuXlDpigHW0w9DS
KRFlJKVgfkXHa6TChbXaVEME/2C7mPTKoK4T7izPh9fgEQnWrj5b2BWiqRlboCBGpH2TyswtCvjS
FcsYyVdyHznCG8QEKGuxOb2uYPqRS5BMGenD4Jp/69Unj+I3G28OazHHm7Y6xz6VA+NkRudb2WQW
SqIvj7rs+v9E8tXaoccBoWYeakoHWVXIQUtblWp3F0R/bTIwKR6TcQXH4q+nLYqeJ9VKDc7apWJN
rQOumIxrIpnl2gGD2qXrXgB2Vvad9xzAyY5vtX09iQ/uASxvcZQV5CxRtYR+c1FiQzb5UoKKQS6X
WZ4xGGb2ggvO1QZ8sWz69aQ+YNoBb5l/AzhqMEzw92o8AKCI8U+WZzX+0GzVmfnX2GErkdt41fkt
uZk+kp+1gopVlqCbrdphE95TMiobIl/P79dvrC207oUpnUHJSonjOSmPTxMt4uXUv6daWHvGQlc+
ZRaJupYizfYNt+rddku1nhXJuhZ+ROCFBvjxtnXi044zYxzQOIO+OQ5deL79qlH0wcy2y2XBb9p2
ThX6nUL2JmAhR2n2nClYOcocc+W75yLjTj0X5e2KkjvDqo8IZrnrozWAKv1vH+JKBrwEZlMZQUxb
Y2/mDdkjTYaHS4Q7nP0d0yY2hpH6/JogffYTm4RNokyXjikwd2zL/s5f9Xhx0QFtjMIio4aspgdF
yvSrmfH4YjsjHw0CNsXoT7um6BZq+M1GlFIDPkZ/pEIzVJUE0Tvczqc5jHFD81gSya7MhDW5vrwP
+DmFZL4jQQQdqUL5j/4EMeA5pw90Z/JqqgtxllnhTEImJsCRfkTaqkXdKA1/hFhHJjU4oXhjgoiJ
yNL6BLl2I4IKm/gGnFEQXt/3kKlwbNrQupdAaQ+ST/f1Hh6eV+TY0P2dgERl6twOujbyOLadJIYk
ZfKnG762CI7EyqlubApCe4axdGd+fgusu4MNXSeybRj6x+X21RLapZlB+KvWdxvvPY5E4LQN30Dh
J1Pv9UnY1Iyqkr+WKepSrqoefgR//1JLUc2me1jkOkEliYICD5d7x2JDuIpC4jfJz+aQYhcUuMkd
l0gcFWmerar+pBMZcHxhcWlrW7mvfB7iFVq45BHIIFkkudScUdm5wJ37YuxetflOWdLKpOGmIfHq
MXfKyl5/1H7rCFs3I5DenQvue82d7pgkc5UVcsCiSLoeH3N7p8dA0fvwcVZEMxP2QK4Y3l04pjFA
VlmOlM9/BZROthyBYvruwQe1VOZHeXNUppzEcoVgBaq2zwfTM/VF5SGG1X2+HTuy2iVxdgTmP77P
3C2jhGxI0e5ZSQNgQ4ECWzSSJzmsSGliFk6QXsI1Y5PSTJZyqZdVR941QYl52iwZSSiZRHrayhsh
Jl8Ev1qAp7Xxp5X+VAXHW1RxCpgwqDJjXgqyXfEKo9yLqJNewnGdzx4oHL1wsl22mFRoL4IcZRvm
8KpwMt1JQBSAyFmBGUmTuw9fbFzyVPzsq2abN0RZsGgluxeF4pPwX1UrnukGK7kFfxfMPZX37abZ
Lx6MEPfS23h7kUyC1fl/ZwIxqqsDw1Na+Z1/ZHND5fer5xxcYxP5YlkbFi7EHCag5JnmVPkfxkz8
2DqMFhRPlofAYdHrgIhAxEYmCF3UddE5XEnnMFvW3ZOjmmpSsg8tuTzNFB1d9jlY9/m4v95hr6vE
gCnz3K0DHUVA/0rImJ1pUwiJ3HUTo7opis5iHT82rm6eB5WrjVjlWhROTDZOSb4B1R6oglUa8XAg
w4U728QflhiAQzYxqSQBsM7kjs83Mrxq0PooLK37YMBtQZOqtwVMAye7BJgNvEV9XTloAjzLpVjT
ajfcxyAifeC5rGhE5iZXdy5wvX8A+WA2kPlJtPt5iLQAunkHk+pxzmHME4msWjW1TTyHoKzgeKax
DO4LqHOHK9juA/oLrdBKnx0rQEkGW9J66KDQ8hoUKIVRo2z3sNHi5fuzuSyWzEi6R9+h23I3Kcks
JL6uPKuiVMsdYiUx7EDwd22KNs36hyaGszh4RYVGoiKZE0CSLovHtSfG/KBArJz0Z152dOTRHLn6
ymDRAefcsXSbTBJOdxUB/uMgI7VKXQhbNpcfknqquqpEBfU/EPad6n+i+6d27uM4FrE9G6VwjIGc
hnBkGW9M5GtW41GA8rBOCAk3aZfDrHTunNgnerZq+qC2PoS/BWSkw0EYIvaJQRL3WFsf/SAtbtKu
Ij+iEpLR7JrBl4EIDuZSm9yb9D6b4ASfOiB8bRm+82I8s1bgJQMA+KJm4i/+fhd/0/rPL/G2D+UB
4Lm8WkbVhj9pOFpzZ+pBCXOFJZbKrcjGQQQMT0pECUqbd/EdSpot1G4ZwumqItY0MX6HTytGQ3rt
5ohO3NHiQuBRfH1Oxi9Y3llnWI1GkmZdrIevgjZnePk+pJdNMMm4B2dRxxAlMZppa6rufPpKPVFB
19DwTHvFoNV1Dzy2zwr48y93Mi2w1AaBEAtOwCZuVv3aDCuZCCwJfj5WCXfI8OdCpT+2958MZNbC
1QWdE4mnvzZa9nxKRQd3i5lkJ0/tCfQ7xsmCvRWc8HZ7wMpphE/RP+i6+Uoq5aVNu0o8r6OnkIq+
facnWHTcTF9kCd4edpvDjlgzwJG2e2UxhA78Aflsa6w3Foqf7hO1/JwWFFJxWM9Ap7au9Xwj8i/5
TKVltuBE1/8W+iizM0VvNHzgSR/P7teohc40DOK+gCSCmQQXTz2t7DgNgS+OdhhQlsyvne06UH+v
WAlFlXv+kmQWXWeCExzCBW3UP6HNOMs6EBprzZnebxTc3mH3md+pJYp3GeKIS7hNe0ZsR/TeZI7n
OYqVGP5HizfS3xwv6lU6z2WzbPpNJm/peEnCiat14tgH5ysnAk5BGiDhn/mW9O3YKRNPxrhm+32k
shMyo/WXleRNMEqYUdV5OX+0su0dpf61TH0UBK1ThXdSy6RAwt4IUnFgkgFvB7V4JHplnQaiiw3k
BVd1Mmv9UqluZcPFKXHMLPNuiklOdVLkQNSjXIODW8WlHMrgraungKRGsDsVNHxAQzI6DA7OroLH
JRFKf418GbIUC7OYxXP+6sjjcfl8oIquvGQW6GGiEcxjGXbsO22jBk4EvGrUwpf800rvu4mdLTns
L+GsHoeWJIESYmDpyb6ZRlGuSNpqceCWTMFSPKbitLlPuy1DScZtsSOQgQrvoi38du9o8kStfEPX
4Lb/sHGVXBwI5pFj4NDBilCT4b40tN4g/Qo4rMJE36B4W0WBhVX+5dJVtTD+dqE672fJb+mSu0a0
ziTgHl1OJA7MFllJg6J5wMaDUJ9nuxLg9jMg+kTrioY7Tq05iQqHhXTp/eIjGOuhohQFlq5+BAk3
Y172ofOgvU+Di+xD/c9I8mF9h8i0sPq1zjnwBiOSY8ZkBIZbMgWgQ7eDA8cjLqdJoUm2Rw3hBTQh
x5wekMVGivHj+upDYdMyQ1B48oBpeZi1mQdeg6B2sSYSwuTX+eMIqaeBWr9My9P0A6w5h36xHBL/
PzvK1YzRFpYKDRm1TCxVmzzPq704xSSzWsgkm7IkOURr/5Ww3YFIp0H4tNJLdMIYVd7R8Wixh2oM
RrJOQcGWb06GuQQSyPCcrg1gypMfZTkqyISNR0+jyCHzl1KiM3g3ROFBCVgS63zqAVhybR9sb/Yt
03oNYSbQUuKfgHpoLSCAsDa+fEp7hsZ/dLxJ6oa39ZS0BrB40aFIZI3nbD1bgBhiBTcHNQL6Frt2
9UQ5XkfU7030659R8JjwqNmky42QPEZEaMIp3yvelXtAfTMDHA+2AvrjP50zeFBH8w2ePolpjBKA
k6PMFsW5Q0m4qgboYH/boccF+pXh/VXCap3AQIxufxiLzK5LEUVE44T+h8MgucB98H7iRHHlJz/y
S/0AnKCPn2i3YluCAURv+XgZ1W0y8FNtkm9+Yp4gdBTKraMw/BFqYumQ6wU9gjbbIv6yA2WV6bqb
SruNQtvfffYy25gX9iGJJoH+IEVG+wl0DNKvKPrO/DJPxevglNURsfAVU5dC/NuU/dVUU0dElSmp
FOwOdsGEmXZys82RpT8N5pG030HXWSF1jpgjLPloO1vyuMuqUDVOBF+4cL74KHS6M9aqV/RbmL07
cBjDyWGHhsqXC0Da7O/AJ1370PHEI+YV2LY0/1VIFS7VZMc0X4tDye+wehhVSbiksmP/MTcc+VVQ
rs9MEym+JcoZN6Jhb2Tljv0Qg2Do3u9lxseUzPRLriGzGHHQCGKYWipdvjW8axRfys79Dai1URPo
H3HyKrYCU8MhRJr7JBb0JtT/MtKZYxJ4FK7EhMywfUHfM0y+ItpLuL1ue6kQSCtvQ5w51YWXEbCH
UAX7Nwn6tzI457VnCP8TJ5RtKHCwQySIhtwLe+zFZSXXkedKPWVEujMpIxH5BjiuKp83BAOKncmh
Jt8EDijhbd8nOHCOZMpxiiiVcngfXccTH8R5Lew2oBonTHVQLAXic3q0wbrEF1bAzUyXiOsAOjsv
BcscdSVQ0OJx+k3WATZDm7ooX7hPXc+RHB6uexGXS6fq164by0ZzEMZQWk+nFdDdZarbqLBBEub8
DadQX/AI7NNHJ63Gmhw34OQJQiV3amM/7PZoFKl+txiNyBe2RCyX0RNFp/dw7+duAjqu2MZ3SrNq
JK+TxmteFaRrIV+fZNej2AH69jhP8Jr413WetyS7W2Vy41z0XCxKN/8z/dTVbe0moX8/zqQZcDZX
o80dgvr4nh4dgxEdwWdjrJRxKKKOXYTupXSDD4JBcM2NyhpzbBD2m0IBYh/Z29GaRv/q6R9wgbWX
zGdhJZuNMcD4SSEShge2y9gyGVII0Wwcod63QdI69nXgX1+Ul/qWEJshQ5swoAxPzY90g/CJG6wi
iR26ym9yALuXrrGYkDmu9TKxw3t4a+8UTD16hpwojYDEcJU1cKIBe/EoTVxKEF4MqPmbwfFaAwp0
0l9AjnV5Uo8hkzQmhwFV2O8UGJLyHKslh0zsaJJkvdiS+V8v9rl/f4NsOvhJdXqCZjuvpB2bXvbc
LcdxFnOjVfi+4sQEAKvjVbAibt57+lO91I05vU0obu28VO4UAmlRN+0v+ZQDcgMNQyFpvRgIOOYf
/CPxROC2/752SaJcBdEK1+/0TFDWMkzX8Io1TdSXR/7E5msnBIGee9sIvvoGaLyb7As+Yi2aP4Ei
98otnPUDkkn4dciLGIlRXSoXmghlzJTK827CGdgG9fjvMxn1VcHO3EFgjPyy4R8tGXBDi24BuUJE
spn711vvximgTgZfuaUCLk1LKverdsnXEmL58jQZUU2X1WNlQqaB6ejf36jnnkG3Hu2MT1ntSdAk
RKUrgjCXfgwr2Le1Kjklcgs4aMVXF7mxIZP8Kol8/aUg1hdsjwbsbMEjGrO3608AGAbz7HQm+sl8
ea8MW7StIEFRVyson/V6tf5vkSsNseKui8mi1cAdLi1XSkUF0z/Z+bKzu8YOt1X1aSkdqtGCimdJ
7RUt0DtUb8VyTBLSnmxWpmrjeR6MJGJjUrWmVZS9xJRAd/Zewznrg0ygH1UR8urYBmVZCVVTgdvJ
Q/VgSLuijiYh6O+T7XYsMw2JPfhY2NmLS5Na+zgTElzMta2f3GzUfQhFPA0AkAZ7ANytOhhtSDNZ
BUpnRDD8crBwCoCl96fAAItk1DGHGcRzTCXcpItCXDGmZyUJ6JlrCYmzYg3169qYRkLR6ee6Vu/2
q9MnGH9HeVqivnZsO/Cn9TCqksvqbtWt88gpZYg1sI6cxZ3BeVSFvpm1qj8+HCiiJXoOz2uCL7Wp
TQNCtOaCaL8WWogPT6aeeCBFtGLCnZQHFpuO5vWHKAL0ozhOxwCYPH5MOsBK4G3ZBOavLlMh807f
8GjCDXL1QLRsa3o5A1aLb/cmTp1tqFp9aFwzTOO07IHadgBC6VjjSYST6f8HeSb/6LN4Vt+rkV0N
TykpMTTHh4CVNDJGxGh715mNRjTr4YnfvmUhzcpAMD0f9yJs02vPXhE2PeiQfGmMM6jK7CrZp6ro
Wq5S/nXy1wDS61qsZRaPRj6aDKvx52xGVS7qvGw9fqYu6Y21g2VjHUjU2EurvY6DCTuQnt3lR/5k
ua73vUKpfFgQmujcmGTgLPEilC9Z49ZNqwFpUnQiMj9LXRyBB5p10Xiw23uqD+oa4QLT2+oacvNf
46JyqhvVHsqfXRL+CWoOX77fjf2UKLx0MJk2AgRWJ8RCger9rH/3j+MWhK6uVwcPLwWQaWoqu5G+
NW7DLaxKLU2l6EQG80yeJfMhlQUTjkT0KFJ4Oogkf9WcNbrI7tTK5/u3s9BTJfH4OtYS8WRc7S2I
SzZWvlCA9UepGgJlrAKCY5FdgJUxYztzoQB3DJbRw0V/HO5ZivLfTE0T7S5V18T0UjSX+YS6uVTV
LbnKkQvg0orjak6ekYrgNfNb8Eqjz2V9hpBOntGGW0vwh/4LwDyUpDcF/TBr6lt2Luwh3PvoNToo
pNwfbB3f3QChO7L5b1qyLS3wExTjTjw24Li2xOA40dnr5vE9PR0ZNpG4NuURiSEkwqTcFnNYS6nH
0VW9bUijVnDOlHk81weud9ViOFQKPAaQUE8Bn0iM7yt6QIqRHgB1eai+nyBV7XQfXn2xAi6NzHte
Ze7rbFabM/oF5eFuFer4rgWTt42iQ7LOox8ffovg0Wx3Q8+xkl34yhIQaZ6LCiVLsn3z6vbj0s1N
HgiKnevrKDPl+8hRaSZgup7yrcjZzZps/pCw4//iSjstmdUpyY6SnsKTsRmqfhWd05SkJhRIgjdX
XQvVGcjl0mhuNLbUqTKmlSJijPy56SSfC6FvE6+ZgrV/zlE6n/PijVekPN29TypdRJKBwdnq+KNs
vRqdBLQC5qaqCMuHPlJm5bZaFTYN7SP/GwVPI3H/BGg57SOMgrN6yrwqhGpiFYO95j9eGsL5D+MM
ee+KzRtRuoy2jRQ4R4oWlYtYL4E5hmEEUaaRJiyLalbapGwBCSEGiCZ83Xwp8M4LsK4CfTC7KCgX
kmGAD5FzlvaXsf0PzjgVq5sNTenTxxCWP/bCjuHT8d6f2Eusm2Ez3ynlGtkkrIVfFxQQBzDhKnWS
hdJI5/Lr8I/vReb7tvuKceYm48515hnHrit9RKokqXRiQP/p1eeb9utpZY7zUXe1YW1QH7nWLyT6
LgQzywLyc0QoWWwSNQ0BHwC0De8oT321ntXU5Wx1IU3jRK7WhJye1kPcSWuJ+9t8Az3TtaIR5gQj
vmRL/5vh7/WBrJRNMH1SAQmqjULU/+W01YSqnbtHJMOPL3U8E/yjssr+TN4h8if10shpAvqS4saC
AIKXcFsyozliMwMwSWWxsnvygDxrDtvxF9CRNJEL432u1fNe8+Cwe1+JtHA6Hl1wrzBptUCs2/rH
rDt1Vkn+5OyX2qjYWsSqdkcTpQkoaQ1c+8UH2KrtthEzGK+lGGQiCoAyvKsBNNTCz6gmREMSRGGU
qVqXmMaUw2w9OJfoauJ7U08gb7hwWgBl7Aa3Q24YMWWPkvfXlIzb40turJPUMljHDPYuSEJC9T0q
yJfzJYAA+BzvDYU7RuLsYsdz+ziVdEY0EmP1TQKiHFmeD59eZf76RJIp7bUuvUc2ftdPJAChUlxA
Sc3aZ8I2mdyaXGm0zXADUoHLFQLbNjD+92CRoM+LZ/CQ4q3nAwO5uyGj8ryYfe8WUKGTlDYtAMY7
F0P+myEaEZG2nDPVVmm1h08bioB8NCv6/r4w3r5T0ZUmxnjNJqTUU84aP8+0sfbD2PJSvy9r4pub
cK8C53RyrZnbB3R14AvjVsJ3iq9lNo+ioHzbnMno54sdp45t/DMIN0PX2oOyzWX9qUdnST+dHyk2
OOC5gASWCLNs/MQX/VtX9LEiBZVN1gbIWpcyiyDgJEIw+cxVbRRfH04H4zOFjWpPgFw/Yz5y1evL
biKi32UTI+rZi2sspzv4D61BE9H27j/wKdjmkiGyHGY/wg2nO45VdWm3SUxC7bfKj6alYp7DNv2p
h4jP3RC8DNAc+nuTzGwUhL26UM5yLzVr1RzB5l0VbkmlogO2JqQIsaqRaOssSuHlw9Z1/Kcxtyzy
Cun0z1ZkL0qZKB2zYb5zFQu98woVt3RVouCFMqq6JOwwbtRjozHOGH8RCfDia3uWOcrctACBwpeU
THmznoSPC8lc/y4gcd5/JviHdj+CnRLtBD/rksMj1n9TavZIpr3wlgFVyqkMlwrYyHl35QuL6b2j
hZAbhkR0lIrSyOTOIVXw1DankCUs0Qh8tppjctBiSZawdzjjez7WVcuDtSCWckPF+zTDtLN1MfX7
gvCQg2hTd2XvK5ZpqlNaHwDWgyBiLlSUANtS6gN1PRKprBgLPzog7Fk/nj+ysSBDJnrS5VjXiJ0V
hh+ozRnAWU0iBUMzrni/i0osz2VTuhiLpmKyKu4G25uGqtdarBwHeFgLFVO/k9SErNBbTZHM0Rt7
I515prutLOD1Nuz/ngRUcLHFir4sVYTIH6WjfgERXA6lwLWNuRYdubdZpEkqnJxYd7PrqlbFdzcz
hNGGB424XaO3IwpwjgqEWmeF4RF9r0WNUNPYflh90SzjWJTl+sVYO4McPvlGLbt060hAK4/nxq7t
aCSw31OtlLikKJssSN2R425aYyFxDVchdmF1Coeu5pxJ+6gAvQOspgi3M796GY4UxYQfBptafvpP
z9l3eCjZNPwdROdwKCP6JHOOzoy9ATSIqQxGUluprnEnUHlBNZJM+4KgrCwccxWAUoICYV8+aK10
NbsWzoroQ4rL0AYhn/aHQD4Mip6Zc3k3vcMfhXcWsgcz8AHDt1YU/mdJQ2dA+8fhSdd5d42xjC2/
mxrZY6gOEg9SKYE1ojBE7cPVhVJH/KxfmppTLznMqryHAefTjYdzpSSW6iEbVW2U5J3VmY5jn+PZ
QNmCcICJmP8w1vLxM446YVEHy+pJZIrtRkjj+W6pjLL8NQWm5072OqFp2p6QQP40/117kfXfkDM2
o+LcItM1pKGTE1WLM87YvZ24PsU84IuxSOhxB8214VCRyygcxLvTh7S2oczoHGEAeG3JPTQxSm9F
OhAqdGRV9obQQOVW+gIAtar7ZC9mDQ/fDf7RPKxeITwFqrv/9lulX2kasP3jYtaZ1MHSrinkXmgO
wP2iF3ydPIszhuOXbrzGAFPfbzmRva9o12oYWD3UluZnZslqE/0V3024JuHmf07SM6Kv4pPdt1PG
FkyaXft4ms8P099RY9U9Fb2dqPLu/VwSOxvs2rcXD4NH0qtbPTLzkd45+MSfCPI0u0Xp5I0OojfM
8v7rzG+pYRcB8edYxib5hza3l+mMMLbySjPVcjtv2N2lfk0bVVmDfC7MLlBC/ZRhtReqTiqnQs/b
Rc1ZHaBVgiwnTVTuIYVohJyISDc4eO/331Hy/AHjK4HWq0ZUVN4g9Vc5wYsibARz8LizG8kd6yL8
WrByPCYypxI5OikIxfEVrbf+dQNZWmrX7qFwm+7w5znYP9WKSHbQVD7AXMa/o24sHOGQU9601sVW
+hSyydP1ivAjGB+ZL/PzX4KlsxKogygKXd5zwwyOIo2lCaUKXhLCOM4iHpj3Cn2iGw/CnSYGv5tD
8P3d4H9eeW4DBJdU9S4UEezstWXdkFvuVq7RJEZ3xEq7ETw5C9c2bg1TgM0A9+y740HqfenpDi82
rlc/IW3j2dK7C6wyhoW12QVGKGkD/DDT1tEMj1U99HgmCFKNEreL/ezwmYyBilCYaugy3GXLa2fQ
7YiBb/LKyFCZ7z8oqK104yB8JLzSfVRCNKU38Qzo1G+A15VRxbBWsNaI7kbVsjs1FVm3GAcT5ZYV
ohwDQEUBucbD6zCYD/kgFNEaB11rOcBv+jM3eAOy82wB2rptjvzgiCy2jpjJp48rPi9w0o/U8zLO
tB9GXGeent946b+ycfwnMZZeD0+drnNWUdAkU0qoekUbhX+GdgfktEsW4nU73J4dVZTmYUaq84NQ
1r90b3BZqoV8Xtf+sHkjVLlI1haHC63XGCJrN7RZiqGB+6n+wlRAE+TDBX2Mzh/HLdbYWhW38nNu
1wqNLydDkGdXApu4G8sjtw57+5EVu7nrgN9mqTpfjwfBspLScRrUTRV6cUEU7K5DZeKT/n2DprJW
h/H5nPzBEFLTrtts8nSxr9hQ9kDtK0jQkFfarrrQP9k6k1yR9fJkdGcV2F9mFC7HCtx6u1wcBfd8
y8BTp0Y2UyTHmG4VpCvB4xDdQ/bDZ/uXsctph/Y55kAOAFl29vT5IwOYo2VyvvltauyEQtk2/EPk
eNAUFhmsyCKRd8SW3TalqJwDObNayOE4+Jr9AtwqM/XrG7BXVC18F/tG/7SUmpI5yaYhapmB5N/f
k1iXBpUL3iIpffyhfMG9H6HYPdy+R+yU2lWGO3cerdOtnIorVFraObH0TLGJ+7/P7WKZDSWEuvjw
H6d6a4UNJXv2dxAus6nnMgjx+nymCQkfrKCYPghLf19Lf8zPifzeNZdIxqvsjlqVNrD+LdachURg
XvaiG4mN1TfP/Akrnk2XtXKkVD1JEDZCm/5g/GYzXRvfiOjuG5TLUaZqVBOm6PZPYs2ZfA6SkM38
cR7oqKBOguaxE4EBXH9L3zvdT2AYRvrUqMar7ekY4a2eX9a+NULXiksd5jzLGZkjHFO1//kJqGMq
oYd8SSoApseuI9z1RH/ix9qBsNKay0PogjgMAbAMy/xloG82GSPJe3wyTtCyee8syzXRTJtwWOIo
Gz75YxwMBaKxK5sKoAp4FVwVk1w4QYeOG0E1n+WSNXyhmswD2EHvQoKCAimm5srpLPsKjJFYA7jw
OlbSZ6oVd7v0hG+K+CXxoi8vrPFdssfacWavIBdNj0gDbmcrgYMpVuloiM8jZg4uVccJzN8F3yAu
cnqZGRRltrDwVENdkkIO9HQ2Z7MSD424t9l2DBTIE6Eal0kGCReW6ApLfXrGnrX/gQ/sWQal0g8o
KyVqnWjq2itt6R6gPWfIWRxjiU0q/Ft4+5r8lCXXEF2F9BUBPyF9bS/x7jL5qqzZ2XkzTnBfI3TX
VvLU20g84a2Lr7CpIgYOBOEew4dIr0lJvrlBNXWNEFilqqvv+cIfbGCey7LyoY2sZVOgLiw9/v8j
m9Lt/foe1LHuWIUHjJFM6V0nI1xwBIHl5CLLzk6Id4Jxi0yMmWxQ9oD6lNDjdd8CrLwOY5aUSHvw
EDfL++SsAatwxjsW8b/YorLrChmsnHiB2CGexmgwKDSmFjCXQIdsDt5kTxEzRm3Xa3WAZXDXe9Bq
Y9tJSlGLtT9sVr+koqlXAa0vm8jAMD2iGLCjOQl2YkK8OwFFySSVvlDHDA6f0mtqOuvJIM1yDGMa
9VrI8TK440AmvwrHmC4GToCFvUbcSmVb2z7j0Gc9DcWSuGsid8MBvj6KYVe50M3Pj6jwwOcQ/rHO
OM0LVjQEZ3He9AHaWdYdETQOsLec/4ym2nfF3nUEFkGeFaEkf1P8brF3u2xZhvhZM0EgyUCm8Kja
THCc4+pOtrp6ih8C+yVJOaVFOb2dEszSneKEtLuiJRlbaNUCduorh+zUwJPTiWYe/O9xVAS4sbpY
hUdpvAnN49GRQpVLMkqb5vQ1ADMwbrhirX1ml0manwljGYgZNuTsLRLYlYG7wBE08azgUn+BFuXV
AopIkez22Q7JKcv7xVdXiNmg5sRIJHPApv51W20b11sKtq5LodLROMUpLhhiR1b7AonprrVGlVZ0
9kblT9Q3eGf9CF/sz8s292Ge6miR+eXcD3vtQydJ0vA+ird2wdOTPiHFVTMpYNrEzh2rq4kE7Paa
dcdvm4PcFfSdh+aq399oQXC6lm60tU6C5heuLCp+FMtVrxXhcULH7u0LBcORhmdDdP2f/oU8aqqA
tA2a2DIrV2hAeExlLxjd577ThE4mfNGWCpm5VeT75GcKnpO3eHdCW1P5ZGfs8wad2S9nXAf7SYaT
bRp4ylZwIIbbWVXSqqIoeN5et4TO5umVqCkLdqKnThur9aKsJBrZdGChPwvSYAR0CyJG4ePox57z
vWEKmOVYQMOTOaxKce5+uqlGNY8hmvhkEXBbdwgktFnbpUHxLHevmZjhUb+9Wzh9SegCkrGvr1Ui
pXvRiZjPDkV4kTP+LY3h1XsxRYvK5YTI3lsqvFFxpGgJZywLLq+fMMg7X7cDs+9YIM8jBvB2qwZM
1QONhpYc/wu6188Au7h4uu8bMIJxdtj5/f21D2fCXA/uVA5DI2X/yIKuwy1SXarveu7HAuZGFxQ7
L2ztRS37QkdA2xu0IqP7VqUwmZYIg4RaRwoM8UR33441a00FNW20p66w+QpYGCZa9hBA9KQtqupJ
lSSu/T93t0EIPTLhdclNCZIDs4SBVytTU1CtRRDNo4sBmwZwLdNilw22Bbaj6ykYbVlgs2d0oj1I
HLsH+xL1hFbn4a0myr3KMct447HGm2WhA0wlcT3YTMBfCWS5kH1Keh4xw1B3O2OTWC8xec8e67I2
E5CULv6geN1z5Jtbhwhqf6tRq3omq2+gbOO2+yD2LgtW8WrEVs9Iq+dXCzGhXuuCQYCDClRDSunF
pRqrpGTfr4dKVhHitHYMs6mL3Y9wpYDB1l29JdlDUClIM9G7KMhZKCnHix6mBdANu7j4yc/bSAT8
dIpN/G6cNT2SLAczMTQilmiZarJ2BAij3AY499vHxvVDzz59jpF9rp9jttDpQdSgHBspgwQMjLH4
DpEGsjMbhQ91RsroG0GUzXENUS1BWwgy9KWGIYsBVR6kuA+hBnzWmYq1F3oqWSRAOvlBWuW4fGkG
y8Yra1E4X7wIlUkxN3VOh+z1zwemCFEnoejq4Y42O32rVTQ2X4BTdoDgNS4xLhQpCz4EM2t6rmVS
nAKuxXHIKqPfdECywMR/POt2WXRjrfPh5FSuMVJQ5bu3nnK2cn+2nqNcrPI1RDNbKWoJrw0DuoRf
eyIou1baEi2/jK5leqF50fTwjR1rwFxKREBf/oU8aLbOmUU+hV/E3ElYH1IGbcxJWynYPPD9LjF3
cZTT46DVa0RS0WfoIeeG7yEEbjnFhOgcfDG6hUhkk3HfUsTD5mn+zcGdDefuiVklwbbnQdeoxyA7
YcV4RbkSwy1BSS7la1R+1KFLPEjSb2o8dqmfUrvvy3tsU62eNVmJtLiYoQQb/bJcHDU4ap4oFsbR
ODim50oGrBOL9sS2Q4b3vddo1XSyo+hAfP1RNaDDBAMqW1i95+CjoOciBDCtQwa7iWaa9RRYY++F
WQEID77kb8BszyN1Z2Ev7hgmihByrhcp5UhGcUxNvVlJWrQnK3Vh2U4VlSy6eokVXKSOm0zlvDnO
Qh4Ice3hitwVt+uKMF2E3p4gJ5PWIjtuCjpoSaXPQnPm5bvQ0R3LkKj/s2UUbUd3Ac0aHaGzV4qp
RG3LM8Zk+N6ngxtSs4zXhfT8nCSe6SHvnofzE1UL31DdnVjHbln5zHocxGj0W93oY58FFlceEOZb
j7OS1ZDhf+eGS7qtHjzhUZmvBMeYCnWqtYZ564U1JKcVLfR1h9yv9g0OvfnbxRAna+AD6G1NhMnc
nvp7svl2PLe/XS4LaovspvPAIcUQ3e9F/I9u/U01z5b043UPOW1gm0Y1niz20bD2cXrP5LmzWZ29
s9eAq7oVEVO28MzyFeK2ragIJtatIFvUaoVNdfXdGNH0yH3vYoMuyIXvipxVmFtwEbesE3HmTj7l
wFtsjxhLyew2IfRmi6EhhlxR86uu/CsyOdYh60kmhrYLlpd12bwbZBUq0aR6kjlRbj6w8hleb+Xf
X69pD02PCrbTCkH/piN2j6SFiM3+9iHimYH8lNN6QZQ3EE52GuJz9W7bfP7X0lDvz2AZvPs9mBxl
XqrNcuKcdNnafjsOg+GTsQ62JIwGgmAlJg47dmUKpeVK51gsSSwYMOWTXz7W6+z5kdlUgJUeKKxv
Ckg40bD+QZnCo3Ks3DBjJKAdetmZIfmRN2GlIh2oBXYX1X4ws/ff1T1vKNrOabIAd+NPGI+M4jjn
kLEQx4uqFVzK/ZDv16qREREWMZr/2bjabI4kT4K00w308Sczr13ATthraPe0D++T9fUTm7G4sl5z
7Tz4bj3DfjyuE5128VEjdAA+cw4AD8+Ddv7G+biCPTueS/hc6HuxlS2HFipeygfg8BsXovAQt6uK
eCQHLRTio6MshzWT3Dammsb3SJrVsyTw1DkmEbmF+YWb+5/jeTvJNncMV5+APg7Se6AJqSc94GQu
FW/31wC+pSOzYlF2VnLc3uiJT3pgqGeoyEEmOqwCFg714/8fZqB/GS3YnzO3EOYjcRCOfOVg3aX1
uIfJ94DXeFJSyvnTC5j5UNqGJE4KlnWjbdMm2NaR9XVbhtcAR6axjLCZlFDCKVzGgdsH5Al45O2N
5xvPA8wDXspgPHt3gEmcjp7RvRiTE3/tMnH01KfOw+Wy68qDdbV/2X9ulYm/Cilu+RJ6lY6P/xFp
7/0JBGLumMb4hrkuItqsXlRX/k/sq+djwStwU/gCRjk1c6qp9gA8KeEiMGcyw2Y76lRc28Xm3n7E
90QlJwpFyYdNZOr6XAvuScFsqYhOQ3spzuURYz5roxamie7bWViWqEYIyUXqWzhApgpAJZORLg05
f7nTJecxbgNJHZN2UVIr/3G9Ya4+AQxEvH/DXDtRv7DjEEZmpF0xK4KUulnKTHpZPSFGw7Sb9tHH
d8eA2t519FZrArwa9g1jUKZU4yYFnh9ZKlJcQvbo7J6m2a/U82tm0BSbTSznRhsHyzcFTD3xSyLY
3WCx0hTpn2nIEi4bcUDHVnJ4JpQmdVmGAx46Uj1vWSWboUI58vr0DRlO7W0Gxex1Lc/xPNZ8AW/+
hVATZ+x1HMunnKuCelKYSkLbK+jVhj8i8Npf0mvNGWLoKgEWGJv6vLjvpjdp439/K5Ik8udsHKfd
Xl0mNrdw+9aJKm3WKrCTzg+o8eRj6XqLLRtYiGNRh11pb4tvgCez1EkzXdN3o1MJ/92iWy/Wkyyy
r7fiuMUIHSYQwux96HVT0cS/F9QqfiKMhxXEYDPTJBrooYJ7wSF8Urqsiofoavk3UvoC/1t8N4mP
ms+5mg7Mp2rE4OKhJVD209gnkBpaQ8Z7s9/FCjQl5e6KC5JrLBB7C+inWxg+0qtqzP895d40i4Eh
shcPMBS1N8xtH73jh+1os0kjeKL5siyGw29nlmJ1G0bhiRHVjyrboxQKeT8lCgI76zn/Ft2+QKuJ
uLI0JEtI73hnd5YvQurPeXNmYV2PlqkfQWypZS1zx2GcIBMyvbWVkX7v5ueaxzDifD3gcrc3Mamd
FbE3GFKtjALNOKP/LrXtt9DPZP7wFVU9ScU6ZK0cPIlSQ4+l6ajyFJcim5/gBD1okZ6Xg2XGW6Pj
UUuh0GJ628PGAtC4cPp05xjprUffpi6rPKBhJgVXP9Vj76wZ5nrngs4NiKGZusJWs+f8vQjc4SMn
ejilGV/ronOME42R0VuE4snSf5wS7yF/5f7RizykxDVN3U2FeCCkAV2oZDThCB1BKbCOjmoHzI4L
iah1TuCV3JP9rLFRTpDFBIfgmRdDSJW13pUorHi/aeE3Z+X8j60eTIHzG6FNirrfuqZ2bU3K+vq/
VDSjN/CkaryPo3hYrjbQob9MY8bYbBytbF4mY8QuHcTFACQoFAKo7YMvjCT1Juybh8D6BZPA9wMG
g2FeEZ4J4OMkLAi7LftCn8vhpAUFptBAbqdeV2tZV4bpWaFKDWFUxCDmKBFcamF4wIcXGPtNuh1h
JldYrPZhYBef67teO00T+cmtzVb9DTPye/BsNXgGvDAqKDOPVTd2tX6VYcp0/cxSeMSgB2YTaxln
dzf/kd/rrn9YE9TtK6dnE8nF76zuqMoZrBBRV7mLcYKKVZJJzcXc42ztujbhle97Rd/7AbekzHqu
XS81T8DJe2GlHwU2QmHpXhzMsb6jDkWgy2wB1dHQZgBSCVffsSPgrgjp7gOhlN0PKRoOUPNN2jc7
imxl7ERerb6WcJQIE/8eMTb/yv7oPLdHzUw3NziqtQVK4TuNcQ0adpZKP94vSLvaA9d0Qha2Ad/o
M+zHLjQ49aAFU0uAMr7WPAVl6lmTDNX5FXjHfG/NHGlgqaWU/sF49gaYAmEuIAlJIYjIlaDA1fPC
Mc1Dyo9phnL/HgrG9I1dlqz5RAvxQFDxvRbDFhXQtfLpxxvxNDBZdnxpsBLdJ8NV04IJukEEj7cX
jK34fIbxeF/xU8VnFVg/GiHBsB9P0XAgzB46vjUvYN+lIH93+Phzw/iDnHsGlIF8qYp4dEnrzhDr
ekOnRDzom3sJ7S7UXZ69ucTSZakoF247OI3SW5f+u87mTGz96nYUvNEiZXjaxynn+i5VvaTfj72k
QgWZMCKmRZ1pLYrK7uAW4FvnyfFN8UM9AAR+TcK2k7dv0zd6aloSE3VuEk6PDONR1m32P2iaIa3Z
qZbZUwjBiavniqXZjjGtZuOBg/eMIOCWeG5J1GoREdYCKYMk2/ATHopcWMUVUAlEoGU/ytyV5OsQ
myiMhrWeJF5JkCws6WOkDHPLqN943tSlwOoT7o4JNbUD+7yv1RB96BgYh72A+41vJ6za1gdVkA1O
K5MninTaZyD+apxqDbkSAWtgNsKVCIJE4v+M3ehAcZBRBeB1N48Z5ypJWZUw/o8Mc4gg0l6BS/Qt
tG86fTd5HeffsWrEB+vCbWzF/y/Nh5mQXA4/RADOrH0toK/YKDrS9gyrWJLNm6EP8XaQBHfA5P+h
wUF7pxflPF5bhusPcfUnxGUTum9eznduCxTHKazcX7wO10VQ0xpre0Hx3kX+2FybKJ5olr/7mp8m
/sPa163VZ0HqPu9Oow7SXTpG9fkl0dVRdPkTmIEWAGqEtf5dzZT0NOacZnICmx/d3pRYXSQarV7Q
nc4b7o3cDJQZIzrr7J/6MbjhrObhvZgZTCjXf2XQ8OwBTGXkPQfUFVITMYHKUhMnB0qkRPYIj3EX
2hoNng3mdJbHT+2/hokT3cTF/BYy92aSTuxSWpbgRywEyWsrvK2B1Jp3RIYvRSQFJ/dghVJ80rw3
sAWMyD48/nseaobei5btQ1EgH4bNlf5iN2X3Q8lOK1SJ4eeXBy0rnEzDiI3vCeawF1A7IGXyP7Kt
x1I3WWBc5Y5MK25TkXD/F9n4EQZSkiZO4y+drNfYLQxmjirMt4CRRTt/f+wWcrlzKtSEQqJw5HAH
x2kWwcfT+A2Mig8MjPOmdA3zu8kQ66zD8zQEOzhdbkwBIP6lSJHl1ChveO5oaqFNgeKyVz9vD3B7
gNmHXkqCnY+Zr2mQKS2A3YW98sA9Dq0T9e9clVcZHm7RRg6wIyrDW4G4x90z1lKM5R5qubCDMA9X
lMC5dFuqAfHzfkhDOb3mT15wv4Udc4FIVblumWrF0xrB56BNqLvzzfmnFDSFufX+tsJmVMGT9lJM
hTVpOyPdNIYDyklvclCMftL9Irw12kB+vC5Hq0kSSKa+jV/1JboVo8e1R2TKD5A1WkpDAqLRSxh8
CcN3g1Du22rXSieM37j0IPrguUj6pjPIHMQgOJU7/5qxFmR7WgSDLXlPzaZPB8iPMUJ3rD+Va5Aw
AJ7bQvsnKDxqRE0X8dN0Kp2p+ASBrog+I/lQItb+zIf7Zn10CnjIaS1DDJZ24fEXscfNMHzCLK4P
23HGwygn8q55GFmV1nwbbqc5TOfjC6UqPo60PRdFYAJIJqArvJUtR4lNCwZi060JlEBDuwGCTh0T
A80jnoO4ff10kV+Xe4v60Ux2c+uhKWv8xwHz3jfXGpsmXFJ26wgRasEWlMTKKG7EO9rIc4F+uVVL
olbmCCzRA6703OfVFjnWSjKcv+lIWqeFoTfOLNYMwQXQWvD08PakNAa8MQc7Y3RTAAaO4/tW7gwj
O2QV6aJBSTIKhcNmZVDbcaV3+k6WBxDuDOsREPnUw1154h5OUv+E/FquWzuLgmfO6xVKqCbw3n60
DWrxBIRzZrZInVsan0hD6qFjhnYA0AdSrjpCNFcvud6l/PCXnQcxeqT5A1M9DQPCQ6hwMggo23q0
E2ZxXLUlTuSHCJHt1jRRKSAQyXBf8CgJ+VBm9J28G0ay9B6P1cS4Fves71+mP7eytpCXk8CKLaRW
AvCmDdDzqrPgc8y5SCkHgqHYaeMXUx++1yV+5dGsVIB7sdynCiRCqyS7BtuFNPNWKESfZD9t+hZ/
7gOtp8HxxPsZ7WZvzIWg9pcXUbSe9FuGPaEN1rGNvre3XIUDsEP9rirXw/kSrn/bfiAG9XYa+jAi
tqwDbq1L6GtZSBB7fYq5nJCJiMJ7SlBQvleU5zNFDb8y0PqCyspRGapIRY9SQ14ZeHsJJgpX/7zu
nQCEe70WDXvos3ZltP3VsOEokWUQ0AmdrFnzoI8iEJrDfwSd36CgEGDdQpdghkIswQ/lvozwxRXh
i4dpzExJGLeo8HALkgSNCsRcpnTq0pilr8G2RiW2UhANsNHbn1G5saDdXSadGw81McDLDvm5MM5e
0MmXG7L13LGEzTUfYZlgL6lmApyM443+0IvsLiJlV4pUxO+2xYbBAtPvq7Kx7sIvpUrRdHY9TMrz
mY/aRjL3L+Yz8F6E/YaG7hCA288+bda3+PQcszMFHukS8ChYQVmgBqjp1lpdPwuAsjURugbpi+oy
RZMC3QrDo35JNMWWFIDksHXdqTBtxMpKEsEP8IyeE5d7PtY01t9dfOkPzE9WBkqU9PMaIbWJg1A9
uuhWxm2RI8H7TXeyHm8UtoxYfUXXjlwh6KF55ECA2E7gVpXO3orIK/RBhaM69TE+m+qzXcci6g1S
+FAcL6fUwJoFpGJfle6heWVaQiHzkOPxvzOj2nBNNrObMuFxbpDMkRDtQm+kR0Dh9xFkay+7c2QS
yVsjGvneNtH/EyQqbyJP+EIdsDnyYEj1tYiB5vHI3wkX79r+AAixljmcRb5r3LOhE3RVZcpcNmYt
AchYKMVa4Qx2n9eWy7OSVPQd/N210hhozMT1hZEuKcVPSrHppBuYkatXNVTA4jxKiYjctethCuJd
5QK6GgD6roJjIX0rwPj/1py6KWzSbBeBlmXkDNYwer0aGmGYbMzEmMmTqgXP2yJ6I9CHxxZOvrgq
rekQRLQyWE7TrlHE/jEzuJhRbxbKywFXybuxf9rLCcp8HRqVqO5cf+Ekj4mRJUrrgNm1k/mQJQmO
sPZUgnbl6Lj1bvQ5ZOcL/2pb1CdLUKVH2GVd4Up+Jtv1PrvUWVX7+iBGHmFwzJAE6crxE7bew3wR
kLcZnCECCAmKU/3pyq/gL4tdhsk3JEYhavEAp2wHamUyAKIymJYSLRPSud9u/K1p+CiW1z/a7VFw
2PqGLw5VZuGre4lJ9IPtn/R1u63pnB9OoECFGeMYjNGOAgVrtb2UaPCJJLbyiPTgz29T6yY7BaIw
RyXjr/ed9tJRHWlr44Y3VKyjNkj76dv33H68NLUMZdhctCZA5EFHOLNSaKejOAkiMCZctS5rEjik
b0l4UaVXjeAFLl59Esu0COAl+oC8Uy6Ugu1Y8po7S4mMFU4Uj3h48pnzyf2N+uQyyAcwnS277qJM
nevqqRbNFQBkq2w9jzclhuVCtQpEewhpYQKamHnp/Ky9/A0gLIhWIejqYRGTZUmjlPl8vPo2iIoI
CZseKnel3y4zALCQZLFptSkr655vrY6NjejOKjUd7Uq7lAwUie0aEfln5Pr42xES6JOE6daWFyG+
QZAGxh5wMyT7H7RoUhj4+SvYhcmMuXOHU3t2AsYgL8NAkgYr4XRAjndqxKIroRZFviaq7Opz84hA
KMIXjSv9RDYmqKXfaJJi8F0H17mCsxQH93m5fTXsfEWwo8r9qJivUTvtRe4s7bV9GN83Prctoicw
EbgRpalno29PyIjgI6EiDhCpYm0ZkaX8BLfwBWEVCc1BF31ls3AQ+1VWNorprAMPi9GVv9LQpML1
QhIj/ONumyuOl0mUAHXvVe70dgnBzFKN2/yrnbM9jQSZwHHqmDYLHd59LIyL/lXfBtvB2pz47qak
sJ17gwxsGARlPkbVBQjWUEXeY0ZAO2U8E8T3bF7cpIYCBVE+JgnFiD/ES4FsZDKu160HtPHOJSXw
rcaDYp6CVSZ+h6eI1qf6zL0BBIgqxi4eULQuBDaJ9dmVOGg78fNXNBqDf/VepC38iNcTYMyGK4jn
WQtcCuMQwtzDoKBElHc3qBJAt0Hlu+LQ/h70zWD4p0kPlxD7JHqFx6b3J8ur9/zDPC3H1Uaq9GUh
rUknMChTwXvSYiRjbh78fsLt8jk79/JVIGRtrmODhiF7ePBjqmqt1FgEyuW+Ah8sJkvc3HRslkRM
yim/CSVLww7eO/9Af6RbFZRVq4Cp4d0dwc7RaeNLLZt10Uklkca0cLFIvvlVD2fUptIHyaXoARHt
SD8L7w3MI4HurJqtYqt5uUBJlXP773DSW7jCgp8rx/742dOKm+tGagajrDRHHbyCtR6KFXMIMCdJ
7f2DDrAJ4fBjPrJtT81P1XtNusXwNx7kCPmw/dXifU3ZnL7AwAf3uzFDsOh2gMvSEnJ62M9AlGOZ
hZ3GkS42BWrR+dW6A1sQm5yaUAH1raAPOPTGNyvF3THfPc076ROGTCyCtF1H+KlZtIzwl3zyfPsf
eT1lcX1AacQDEU7caKN+PE5FRb2mPbvYgeGo0f7UfjBRydtv2ehMNFQ2RM3byU2+Lc3MXqjobeLF
tQL4N2GCa55v6LenelGNbYd8Hi9LEBIVoGoIYKTtFb2xdJ8kub9h4WCB/r/SC2CX91hEreXZrCXh
hpiT75wtCKOL9s4qMktpeakkf06T7eBUDFI/mLgdh63m8UBtE52Uiso6H0blM2sJHRY5wniGw4lb
4vWpPmwP0HvMMENJ2AxlUB/D88+5scCJYtvsUEfqx2oR+UkMI3wie74tvAO8rEKVDdbvJj7eWOX5
yOBTduoWx5cJrg0wUjVVgLOoseUek89cjgA5iNydkxyedW4To7YBdBsMXpKAx7iDvww0lOrIjcY/
BRzoByaCXCp8cW+IA5JHnuNFCCAZmRADLuh4XLEpuyKDBCy33efd0J2h8O+FgtzH/nt7V99zyXA/
vBLM8zYJ0ZxBqfIVBtbveiz5ICV1/vD6mExafeI0UqGhLGcJJKEt1a4V4t+dmUwIm12CYth+m7M2
ziDphqSw7MIqSHy28FImr+6WLuRqbCgwiWywVGuz5Zk3j4DeojqL3TBvBLrrjpmRRMiijamYga1A
sZvW4jRlTCF95NxImTtQhmWweJgstYHoHu6MgtMQAqlhtQJktf4WQmUjOTfg0e5HA3UNaYc9d1wY
PhNPzBW95wZGPGQOM8AzPghWnwlHp10y2Goz/YamdwavbDiZNhXit1H4UIHn5grWaM9afyxTPh82
K9a8bb90FwtEDDEXE4qke8AVfT9f14xSY8GcjeqPN5wsSFbqHbqKo0P85YtXjgMNi4SHG2sMhPxk
YLnkApnH4FBwov72mBkHlpens0R6Dmfjcw/j7ue6zKANd3NHe1U9vFMQfqi+OBfsFPp5lhgCVuMj
T8+O51zCswgFPns7MYFbSSRDYbdV1sNC1aBK0kR2reDPzUY3JH05mErkdSZ45Wn9JXzX0Enn0Ml0
BiMHvsjmn8zJu3//c5FVsmzZGLl7v+qjSpSiRW1azw2m7VAfKpaFmvo1lsrtWYpLc+/mBN87jVHC
sosZI5iceOPc9+SCsdUQYFUnhSKsfGu8KVDB/1Igi38n2Gxhbc6Fu5aFuawbMSqeJK/qR5ZsmIHE
N65o9qS9V8EleYDpFWPdQF6ipTwu0sGynfTa0CqWhw6D/O53jTa1+Ph+KAYGST4vaN1nTlb7M+wB
J01G0rx65R9dI9Lu4JDgKHxj9CVt1ZUoq/j3dKGfyNjaHEgofDYvj26z5/MkM3mNP+7U22J9R79o
SPf4Vd6n7HAWjXAN3Ch7B2I1SallQXoJkOZ/MLE8T14be1qAkddD3dzpAeqK4bqCyj4dZcd0Lm3c
W0izhLg81Q2uWTHK4E5+RLSHNbq9qSk70MIwuJOvaQ+Fg0010LqBf8tDvh6H6Z///5R51SM7+IdY
02plGcwNEHfoenFdz/wFN6AZB1CRVnINBoAXTpHUGs9nZ8QYS1IeqWB3p2re6NUXJqz6A1e+urFY
OQWDBeKKBrMs6HX1nIWvgZGt+V1naKMhChOn5baM/cO7mFCg4aXrZcvnXmMWd5SgFh091bCYTm0x
nV9Am/wi5dLu5d/XThKrst12yodz5705t/WsvJev/QyduARdFf+uoqVN5kuSWTXPlB2npxEGzDxF
QHS9TRFlx1AiCs6LJ6m+2wxiGtAswgpYZQU7xjtNjuAXBK2fNMaw2MHiTIaNUO1W/OfMsorv7MJL
H9w2HIPia4Pjx6bJrB28bI1NrYMkxzrXslj/+l1Wh3nvtOS2/ownCrNK2E/SLL8CtYv+QzjaspVt
5XUOakMJmBjfWMU3JwubBSajgZyA40yX4qX0HqA8yrI0UrHd/Bn33uSD3QwBxkSFqOuuyKt814U7
grWFBqFG3LqO87Q/9A8IDREQktCRHt8yQQ0iOTf6PFMSiHFeYGa5imZly/O8Xryy4JesF6+Eswfb
G+wrRWhkhs8koSYQNPQwOpuF/I3J+JUx6dX0bLCcb3oWJhy8WBA+E+cjL+UnAVI+ZTzZc1nZrFst
nOQJSqdCzyL342lFdkcLsDgb54zkr9e/elfm+mtp13ykvRXKwKh5F9mlt8tAJAAANpQ8J/Lhi14s
MOyvYimbxettxX++J5j4FBfS0sm5W+7w5+4MAJfRHkucTs+Mt7m7RdBfHuSVr3520+xh+YD7Lqbj
ri1gI3GVZGi8DmyTT7vnFnnsx1PFcpgUBU353tZmWrzc16GKjbwKq5KzukiOcIqiUiZ2w+Fd5w5u
HkplsbNsedXw3oYL+mX5hguli1mFY+7bGxgHEvkKYYq4wLHyDg4Xe/2i85bNP3ht9sKQjlVzfw3Q
7EXZBpEWXaYu0IgnR2CArCcZj832oxCm+QquGz4Nvy1u97JPCzlpZb1ST+d7/b03uSDA+o+SrOUV
aCb9knWIJjzdR/wFPKytcHauAtlAaHjK4d6jJ5m2DdulK5qvPx31Rpfb+ebjwVZf6aALH3+auQDb
nmcKdyu18LdRnsk8E8tvcyu0mGPE0vwBGB0f2QQ3OfR+jGAOoPl6IXJ4PQUFBNd/BZJ8EOloVjcB
UJDKvIIkaP8wD6DnsPsVri4sFlyTU/G5AkxGhragy32TEDu2ru9YI/WEsz+w1dTU7BFSGWd8B9Jp
fhkPSQ77DyPl9tGW/DVFaC2p7cuqEvhoJ2wrqnvvlf5rwNsvLa5mMCaQ2ByiM+smeWPuv7DqvQtH
zdFonXvbF8VrhLml/5E/G4ao2BYjiHViitKqsci1YyLGeQqO2maQuPrcocWBflzrll1soSdxGleU
9Q5g55fQY2kBr6XYHj0Y9GLRhWG/rbJGL/xAmG13T3dGEPGGkPEj0h0dksl4ttvjpyWLTBadBqWL
S88maFj/joQy4hu5EgP67z3p/abu9WEam2O3tI3FHOJZKs57bhVCbifj8/PkiUNx5D19qyaxxLj7
h8zh6EN3V29gpRz/VKzQdyQ+sVvKlnE1dVbaUyH/WGOn/aDZT7mzf3e5HmTpaSzZLsfw+/XYp1cc
l8iZbUjmaiQ0neRvCPShAi0Pl+gzllbZMxFzQDNBiLh67Qa2d/BWYpG0dJCTHrJTtyrn/6J1j1kA
d1XIsuHtGUcEhAW2jSby0Rg31V+cL8ytwgcVKyluv4zN8j3GSw3tpBGNW8gSj+xYMTwrCritqlPv
okByaIZCiTOW7C5JJA998D2sXN2982h0miTABu58jRZPj/b397sQV/p3BLDiDFemWn460sKac0RY
GiX7DOHn4Wjt4aDusPexxDdtWNRqUJzPwUMyJvRAs7hbHfVpYYN4jWCqB3L/PkTKDgH8/Gmz0g/I
+9MSTPU4/EvzxVHiU5nJ0IifeSqhfYoBMi/rsBAr9UHcpASp8HKFbLy+ELtkPTcXTVFJ7a/B33fm
79/cy1FmsG+SSdxKimEh5otqMH8teMgdaWQ7RFGDVrzXXt09JyuR0qYw9Hbf54Wopw8fUzWP5EzB
i5RtMk05xTIyZUMooeODXbSILldpRDKQsKKs9cZv4/Tmb8Vl5FTLKsFUEvrk/eCwT3JjslTy/xoD
RksQN1BH1ZdsOC2I7Y16OhsnqRzgkYHAtDE9vLyME51uuW/BIzSbQX562+nirQcls8VFZ4htXa3G
Y83tyqPBSJLPC7e0qi5v+FJUp4OmEwgIyyNb5vECaVsFx4UoadbVu71oc2iJmPmRCPezDcUb2URe
wyo6c4CCKPF7RB488RYB4bpM7Z+m8m3X9bHKxoSZWoUxPVZ7Ts1PT2NlfugSnH+2oNiLEW9KzD50
XhFMIyGEVl7GH6p0vBkshu3z1e4dwCC1ujrFqcQstMgGuN5QpGTyHGl5V+PIDG2pmsRdLTEtI05t
goZiN6/88NE+dnVfknhRliQHN4Hz8rOZcCARxojPe7qa3M2blYhoBKw1nwIByj7MxfXAD2hLdLA9
8ZpRzkJpsXCEeO8ojrVJvtISBPGiHzTucJChh4GYFO+rI547ez/4cgPYhV3gpZHeRpGOJzR2u2Nq
wnPIFcwvrgKPARE85eDNhwAFLPiRUCE6G2LReGmczgd0VW3cRmdCo++p/Yra059w8e1To8mbL95g
FMMLDDxRbcub/O7lbkIty9EAXgc/sg13wxMLTcy6a4Y6kOqqXHWb3bHe/+CqDjYgi6N4GVn83+xo
JsNicEOPOHnOAqtXeBYZcS+N/xwE1oyHXG7gj3bZB08X/a2hVsDJVCuLPdp+NrbQsuNxzN+IotKG
6rMQFFtZB2O/SItI5fqfvJWuiVgWA+GjJPr0qoz0BKEzm6cHdu9ZT/TvcquHEY5dqLEkZtDcUBHS
9IXgmuf3S4jUiAAJ+mHx8GobiU4qJLl2i5srlgNhx7oiOVPf78R9hj1YepYgdKpdW4RDb23IEokh
RcU5tNt49EE5QvMzIeOJ6jrgU/eOoFVoav19BXZoVxDZZJpUDBGI0LgVBLDddeonsSO+tWSp/W7Y
UqR/QS/2eqYWBzCeeBTE/oPx36GAs1I7ehIVxArBb7kkLnDhIM/CJ2XDJpGa3iexPUHHagG1qcRE
HjvhQ4q3onZEKCMRzmhxhE9FBENry2M+FCxUwaeliPkwk6wtVXaiatlrXLjvkTmSwX8XV1PlE+r4
Oid9jzmPxFtkg0xTQodOs1OA36fuo595jYVo5fcdYqNcrS16nKOE/hY4R/GPp9eJvIMfhWB8SxKJ
WO5ahDWCJ2Zs0PGMsHhB057/Neph9qkvGXwnJNPC2Biqu8cC8vX0Sg6zatgzeqIc4w10J6TaZiL+
y1R5mcpLkOJFA3+1ZJMROqnhMd95JfUip1fNbOpqOZTnLEXfIETN4n9/UIVvEZy+HWyctMrgwP0F
mH4Ft1tuqzEsF/VY+iS0V6UA11ilUjJq1nC/8c5pxuxx5Y5sAy0emLuKIzu7vQr/gCN8egQnVSlK
VIS4rVT3uqyqS1FDq8SvtQxrIdZzcOWowzM4c17IeXf0WoXbBjFDSA/nRIRh/drX2e1r/4QOub82
v/CivT6Wo3evTxtNzW0H3X/EXZxWX7w2mKQXawJmAE6hTjHTvTlWprmuatDbuderSRfCdWaeQ9Fy
4piWx39GMHskIgtY/F+TJnTQOOzNfbdGd4koMohzXymYR6LE8u4AFADrh6dqaBI1MxEAeSIbmRn2
Znf/Rsu91mow0rVfMnQyRsX+vqkR3w7WJAjutKcgwu02Jrm3IP3badUuq26TIFTfZfUAks1P55T6
N+llc1hvalecrpU3mk7BsqWbKYOC38EqzcQjpAcJwCBXgV1RZw+aeccpqB0ehikSD07ggPvxgNxA
fBDR/hSRf29AMz+MbAApR9kRaJ54yXTQC5D8Ec9e9GwAhH+kp5bN4UoA8nBjO+Xa3VHCjFE3Gm6w
JaiTY8QgGq8N0tqpmZDgr8m9ZaMV2FxeoG1Ls5KHHpGBvdYBybv3iif1VTW6Nd83CZOvL3SkxP+L
zGyDS46jLQOWkds6TKuDWS4E5UyoLMm6Bf9KFGUVQMZCdPHFZec5Yqxu6DtqXfdJk/3kqC0FV0tI
Ibkq7OqF6QepkpfC0KqR2+e6cA6hOc72ryPxKGDFZ4YzGbxglMotYWyU0ovWozF8adBnNdoC9CBY
HKnrfewfe7/FjPaPY8LZeS5wE/33IPeZ/WMRxYy0tCM/NapIaoXcGsmSs/qV4tns6cr5RKkq7LUw
Q5gR5SA9A08uGsqgze9c4n3APyJF7TgCM/A+nQNCYJ//mAm55RGDJIGrH+SHvL5ByA1ywfp4fv6X
YfZQkDtLYtOxj+qKcqpHyhnfhvR9N++3nqm7hm2A+i7/R06JIfe0a9Iar+oUznWBshunenrG7QB2
MIAZMPd9665MN/yVqrIGQ8wrm7b52lI+CDNeWDQp3eDX5iMI+RQU39X6xSUL4hVJ0PTEegnCNvW9
n3TzZ3SB51+v3nY1u4IVJjJHUk5Be2XweCXARTZbTkys4xgLEX3ogoTCtYEh1Sh60NKOitckLEio
8pU9rCEN5yGtb2cgjfj1EF5ohOd7p9k4es2XcmKGoX8M2z6uQgk2uli5osMINYeBxBgjOYJi2HQb
+nYQQ9Sw8I1dyGWDndW+lc4Y/tN3ns65EcIy1gt3/0kVui8bGXGA8gejd6W4IQ9NtJDwmVJBUyR8
/GBQJ6lD3KXaTeaWyQpuJIOPLE0+MlMVbDqelA/3FxP0OcmUOesTeIiQlDh5Ung3XgeM8Viv/bFW
qBOj8tDXdEyRL+iQJv4/VXCkXkkT/FYkvcK+qedCP6W6qH1s4DQ+rC/MStswUlITHPYw3HeP69SM
wOrmPK+WZ7imU898hf66EVDA5aFnxJGHw9ERvbPrWZpBdzdKCk00uZYLsJ/6nVb1mcbJd+NLLvOb
1lMT1DehnhhNGPX6mwoLjmGC73hKg6yRGfJ0uaS3YnxWpVayMXPUH7GLVR6aYC/ROv7LskYsgloT
T0DHTv/XdZH/AtwT0sYq3zBsKm+8qEMDg0rn9srt/wzAZsZsXOzOIuamAYfW17J/PVPNalVJuFnb
nc6xIvNlj2SXFUdf/rmKOSnS4povvRpvXcPTwEXB9LExFKzX5hZtX38dmHntsAqm4w8gFaZw1hVy
ZOdinc3jZEUi2FQ9RiOMLH95DP49f0R5IOi8Kjx+RxVerJ3S/LEcUd9zAt50U/qq3PYPIg4mWmf5
IbKthafSB3yylW4xJAgO4JG0eICwcMy8iknsxJAHgzcuSiol92+Y1BhHqdcFlHEttpDVoyf6TRJR
BbZVkhNApx2J7IVFhQyUUCOllFFyfFmo8G/nwAPNOs7FXvYDEkX01Pzki1BdOxWMtxFcuCbyD2Wg
v1cjdOVxbAM3Hx6v1jBILS3wGfeZZ7PA9xYLhGNI1nsA2xMU0mJWDx+rQ6CYS1MGo8vdlc3xmFLo
gxnOk+qmvmot3n/Af5hI9+2hVxuH0yY1c7abYAkfSse4fR56Cpfys3E+1YivaU3LVsY4EOwHqNwL
w7SUBRkKSXNPz3ge2vDnCRftb/ANvHIKVpGyD5/rEsECmWQBFteO9QCbY9hzTcQ/6BjKetH7o4wo
JP0LTSw40qx0Z1YHXVTVByvS1z1aXRBuqIdDi7DeEICHD6nQhbUAg9ONxqaRIevjkpSHZTSfKV9Y
VK3pU3gyrHvZ9bVslQ771bquvLCOzJiGfTUSbmcKpE+wB7vQN3dyfOt5E3eQM7U3StYkyG3/uzNd
4M/xizvnit0Uj0m+QucDLv82dhG1AMtGvjshkwW5BKbpWmgBYQ2DaU37VeGII1zBuulGyO/TnGlM
es9hc+7tARwNdEVNZqMKdzOnDOOZsr7wv3Ys1b0yG+NjsJxbLPcltBvBbvFWnecHYGHgi0wFzvX9
3FQgAVcSBkW3lw20xgHiZEaQ0E48+tDROZpwmNseccxN2zlWPNOY9w/JwAaoIB6vDGtDNApxSehL
Nri+NUpJk+Hda0niMYvmW2rujt2cQT3JHG0rog73XXXDZxWnZN7EY3id5koFgQd8mX2XKSKQqz5N
MHZHS1YEXX7CoBz4b+6JLHNNUwvXCbSi7utO9vsPimM7uVouWZI6C+fiIyOqfq00/kN0jQGC9xzn
YhQuB1kauD3pqDWmNRaKRs/cM1ROBQshnZ1N5qfv+OLbm1CkToF+Yg9aBE5U9sP2XApGPI/GcmCt
5BwRiAqVJ6s6CrSR+7mfPq59mMHsXfWs0S6N/Hx9n/rjZxsrB7awh5aSbqTt2zikO7TwB7qQMsJP
2dfgcCs9uFBVtoJp+TdyFO8mgMyEffM5XCkbmdAbKa1BWuliPtKzr9OoZ/Fdy9fnTsPmq45bSXRo
o7UncxOoYgxXKSbzSTjDr7EfrCeASz0mqYCtcHf86AaJ9I5gM+5j4zlbFSHZzMA0bdw+aa6zliqm
fE+rAEqN7qZnvAdRjRJh2XUhh1Y3rrW4ZP4S7hV+4ablzYB7TMiapusInZ85A18emh5VdqMgYapc
RTdzK23p2jy4dtywZJVsxdOD8fHKV4MH4SkUNNdi5DgmUg3aRii8U58/xl862f8hYs9zCRnWXyuR
WR/WaxCbc9zljL3bC6snkm6up2nySBlKmAqSRNJDI2a86GH5lBf0zaEj3Uw/tfIJodZJm+OdGbWg
x2P6D3CZ2b/hfgdc1UXErXOtyTkJy5ck2ofpzwIVkdH9UkT2Q4baW8069lEsH6xgHFJaA3d8JsHH
LlCLdLkn4mfY8KgMeWzGk6G+yIWIUv06rIXlPfvYfNLVnUoLzEGiTkhdprAwcb9n77Go/yviryCY
A5ynkH/oc5WAUh9p4rNkqqn+V1E7R/f+SyWqTI4FO+GCdJ8wLpxxgsJYbGQw6grSuJzoXOnNfYWC
cdCfAjTpSv3OdzBiuex05p05g/of1HPNj1+lR+jYj/YEm6jxXrU16cAblhQ8BBxXfbpkX5XTxUuF
YtTBHRXP84GMklMBLBxCevUaR6Ics1LlyLUJ0o6jQINA5ji1ryTKz2+P5txNmT9NY5YU23zbS2px
onMm4Y4m9/cIPyboiGUJYVXSzbVTDUx3TGyWqfe22S420Zp79/w6oMHogUXUS5E29BroIdRxxpPK
aEHIXXgY1mHo57xaB6JUP7EOyopxEQECkDiLy5pxNVie3w+r3OZrpu4emh7K7sxTs/CL7vIzTXmC
7+9zMvrlL7HVgJCVNqV6GsvaZtssAHKDFzXhCn3vGltnqktmtTFGfitcy7fVmHipLtp7WMaRZq5x
5tKEZFjQ/3bMT065b76VvIKbDh2M5gc/WP1CnbVGCdqTpuHJ3vlfU27vSEud45zt9TLtzYoNZnIY
5jeDlbRtqY6uOGrHTYxwOB30PG7QffNcXBqCYv5gSGf8HQrJI5q+nFtfqdWc6j9jeI6qYf+8+rp+
ZlZ+cJe65H3pRnuL1e6g4NqdpyQy0plQ4+E+5b8aGYLt2NvEYKPbWqbtjZHxsCbHPuWcJXZq+4xz
gi1/tYhXXKwa1OxeiJVjtqqEtYBlr8opi+cFdtpUaKvGBxdeOsGGMTBGHWOsefbiBZ//BmgSQeBs
sTTNNJTtWLbiNdFZ/HbJ1kbUGv+fPvVxGZeG27YBzLnTFiKDmTx+HSiJqe4qbDNZDnzSuP+MzSaI
DfTrAT0wVqp86ZZAt3pbrocY42fj0TeLi59mrv7CitoKmpKn6Mg/byU7kCoogLcdvjz7vQO8xu+s
IA73uTmXPJeqisz+EI0xsZo0HDQkwvd/h3H/wtALsqCZIampsHuGKrDzYol99PoKc5+XoYzfyZtD
M/huOcbR2OAz4IOj0hQGbYCQg+OzecyTjhsciG5IfC/OXge3vz+KZyB1ne2SImjsV5tddpcxoG7V
aKgntEbNEn26PWqCPb4duOfGeVls7JER6Zinxp5O557GYMPlblzztcbVQw35NIw4ZeFpbdaD+FHk
jyMlOS0lkIWUpoeVpvsaxI2pl0esH5bLZ6fxS4BPzdJ5TWTF+wMdqC8LV6OgBwW/ddi2kNWbab84
j6nZl3bN9/H2jaA8wlxYwtoyXx4hWVGUxUB/zFebLdVctFVpSQaBcc0Up0Qa8WMrGmeVCEC5z8AP
SVE2STaEZ5IZk+F4j91uj6Wh0peymYgQkCFOjYBnx/ReftCnyVrNl+bXt51joXOG+GtQhqFrzKiB
wwCoXgaGs+hiNYWC6vxwjE1Vn0Abc54C/9xJbFSeZSLl/rNKW6NzU0P4OEbgswtjfmiemReJv4t0
AVMWrXJqBYaXB3JsypuQBSYY+LLgo6u052VTlIh/QAH78k9aTMtCctjaH07/cBunSuBxXZ1yeujR
0uhp/zvgrFtN9hU2BSIRogity1qTw9A9JvzxZMe/bloiwT81bjtFft9v+ZPwzqtDNg4U2cvrwHEe
UTxo//fZhw+KPP3WiK5rIvdbjRKqpkCC+O6IjVaCesv9hdFWvabuLu95Dr0X3tBrTr4dDSrJnu4V
IlhfeU9jtGAUovM5iWU/J5Q9gL0Jsr+tJgofjn1bL2/qQNNQehxodLklmTMyjCK3/DhH7BObr/cL
TluHZ4v8UltfKdpss15ZkUQD8Dq/Oqp9FTyVvFkhKPB/OVke3k/SOnMvKGUfddRDPanYbnurHOQr
HTEoPmmZlheEWmCAGKfelVC+cX9Mq0uu/pUy2DCBiN0tHXivM9xtE6iMxuQ99bvM9F0AbC02ZDCr
p+vsbe/42hVrf9JgfQyrxzN+p1ycaCkPM9qm7N7qoTriVYekr3eNmZnCVVjvjlCO7Ay98YpWHKpe
pQ+B0t41XLOS4YxN9bHijwEkhc8Q3FFriiMxc9Vmh4IjhH9ODh/sRDRwBs6itsvdFcqtVFzaNxrm
WnoNfgpSuqEx+UVZQ0nyVKI3EDRXBeA5VbEw52zsoHXJDUXEx8hpiLVel/uohpxLf5JGlX2CwnM9
c6BOknqDxl5wAkgWAyWkxMI37Yk3vF1IDk5z6r4QAsMwBwnFtYFiBomhTIv//plHLwbdFpiC9BKn
gLaKldg6BBEPfP3KnlLDvY5KVA9uIFXNsdn3BgBmZLizcE8AkSIkz5Y5jMlue+fPMRD86a8IFPtd
+/SFa2SWXhv5WBLrH9r0S+3ReDUNbogJ653f+9VRCvK5BU5cUeq10CJuMSWpE+Vqxty2PzoZYMvL
/y+tPCGLxlUwQ9vqApm+IX56i84yPmcP8a7nBbzQhv+im6XXvWT2N/j6GM9dovMqFND3/0A1xuEL
0VMFFb2ZjOCUcTmHRg0gm4ZDltBiZFsrO/eJC877UayNjmbng09Nr3G0Mp8IR3BEKphgxNlWAq7t
Tf1J3fNjQjxg/OlbB43funQmC/AXtUKuKUY+PAw3iPeWcAUEthAksFUf+rVoPGZEosnfZ27t14LQ
tYwTB+wYjgZnLU/DcuJgrkdpWhZc5hhf1GA8KD4OV4gvlnIDkaJClA0svNPH1HXHYCuAZr1Q6vCc
xhpnXSOhDcOW/M2IAqEQIxGaEqWAEBSgv26VAY/slpDxI/EkuY9SbZ9PMW5gijLDhy8PkovfFl+e
FqjDcgbDO0JcaQ8M8hI8SW3MoAcQz/N1iZSc8bxdzFybOqj6ft52WCoyKr+A2IwjYlGr/R8nJRKR
mXCVnOMOHJkcqDpiZZfHm/9wwPKSsnO3xFvOl92IBo3mUGj3mzj9gLoFc3T5QfZ0X5DyrmQLcHCJ
vYOWH65j+hFKsp3UvNg/qENu859tv/eITYG8Yye4P1JRrtyHo1yAg++U2z4nVEQXtNTySw14NT36
6c9T0dd7ghiK1RSCFyA7AYgK9MRfemhKLmO6ocSCn3MPc8hVBF/YXoVNheyiQtfMdo5CpGC7gtU+
Clrqrn9zLlD3YSfDIB/fxl95Gh+435fqaNL7AztkY7miYpM4uwTCF6b7cb1vqvM0woQtMPrH1wOc
DTyNf5YOM575abAeI5KXpJKqhhtw2mvaHlYWZrWhzKBkT1iBGt1X9/OnFET8lEbZd+r71KB2WqAD
toIcGeldlwTSkICju1/ZEBDzfGEzhtgH3GXNVPN1UH6n5bOcp0yHt5ipsnIgWi1G70SeE2nPy0/z
ncp830ecB1rWdFiZ+GTjT9o7rQYewhFwY38cWGJsLgCETTDq9gO4pPKE5A2rtVBhOcyUVjtN+iot
GEdCaHynLBDrs+FaZBSYwclco507RuFEA34o/grhzdZc+o/7Puk4QSP8fju6px2r+fagIfEoxjAi
sgoY+CYziNtktMvWhphjmBsPGrB6DS1SfzKjqe6/atlyTdAJ1zIz1sKlj7A96XRsI/CSPUHm2OS8
Kb5xRF6ic9Wk/kGtfUZ1YQ6W0wPYJTY5LpknQ281rb9PiZKHYrp7QCe4qu7ldX1QaZ07RR/4wGWV
S94IuYKOBNZacBgYKS3zQTqQPBEwCcL9TeKYr4m6F83MP2iBdkHByFlKpvROi9DLU5MkJDMLsMH+
+AJ8isvu9/MCLQsr8DWrIgz/q3BpsHIponIj3aPwuy2cfNPqP1SPSFIFga+1VoWtI2GFGHUYqNgQ
FJZPNJTEFt1DOfAcMHKwHxvtwJR5gB5PAkhBJorrPS3dObd2HP66N0k4t81jX9+/dT5g7YlTmQBF
mz7/KdFgNVhJl/Gqr6ENzCAXRh6fVb7AdmBQ3N2273+uyMJugG6yT/z7z/UtXUfSIcxT9MCvBBEX
KPY0uHjaig9xO7ehGWsMeEIA/Zg6CUXwr5vAzfeD0N8Wh/AJMlQTlUEdWUsGIRyuZtr7HSTt8s/1
ZsC+ViiciGCv/s/b3GpVYdCRwM7cT2vXY53H+WwWK4Lv6wA5yBiyLyKH2PcOeqBci7ohrx2hp1PO
4iNiXC11qS+VGilLpgX/UoU5K4w+RhqhxP3n8Ry0IcCDflNy5MEMi/LeBYy3JkszqBeWuqPHNAzx
57totY5+rN1Q+MnYX0a6wn6awLoQHzXfNsZWLLQqQKBZ5QtYnfr96BL7BgmEPbJzTOxfFF/CfnYl
zzohDN3JNpbFnafGMM9ZKWium5v36ajUrQMW84ugXYRB86XLdZzKKaoKdd2edMortK20YRdSA2tj
uCh+OZNZ7HN+OKiGR+ziW/E5mvrGUMrM5HT5oLZnJzaW142CBlkQT+4KH/hgA+DjfYedQAsz7Q7u
Q9Hu1UIUGSHI1QmV7/NBlEwbIBRLz/T0NfpyGpQK16n8LtTQghZpii9uPvZdzIbV9ON8zyBDj+ZA
5yNDxtCqOo5gGcpvhkLEeh5BKhH3nXgVINs/moLo5DfKy+DL6nY2BCPTylB+7WNnv3MWM78+500+
rp9bnxHHqPPFpp7xJmmbikEYhCpapQDUzhY+DCWoByyTOci+w7FPPMQ8vKCgFwdYqLr9dqkTCNxb
ryjeAEc1EC4oXgSdaNh5Fx7oDUhpoa+4IdQVa3vtUiUhZfyWR6IzMwNog6hl1n9LLcuP0LfrxrX+
EL29DchY1t7tkkcc/cDmVutr3pUTx4PB0xY3yG5n08pzZ/tXfy5lPXDzBmnW/zwrssXcULll6Seh
5fZFsS4sVZCtpdgat2BYQRaej1zWp/4Sc/yaGrkb+F2bCLpJDGgNFYVD2aZCVGCIdz4Gl87NEV6l
mGso1IecSmEkZ+AygjI39LDDF+2YA5Cb0duQHAjy6R/PMsEcvd33Dn7CpcT5Jsssxzq5DV3g53Ez
8OdMx31N5cIVx1tMIxugNDVelOY79mbssuAAQdq5AqRViuR4RTkko/yoW47oQkgIbZdNv4+HKHsJ
VzZ2vE39hdf50QyuUbaN09NyuvIqjYnCQthg0rfMnDRa1VsVuZmvgrO5MnnNKXtcx8/S56rs1KTT
cUAbvTKAi8LhhEw3J4UZ1Vihm1CUCKRNwVJ7uMpTiKYKtaLTj8mzkuBJCQ2NXX0Gzzmcbf1WwUIN
qslWJO9Ez3oS2FICBhmx4trfDGqZqC5+jVyXnA7XwgXilPVl6uAVjNtqLPVwUT7ne/slyG3SfuPZ
CxRyIOxMBAJXXO32PaGm7lXwnqmszunK7T9ydxfn8ZHWqwfJjFWKg8/982nVA0SbwLJGVD6TMJFR
ubjhWj/iCM2rZ6fFke93DBDfDsMCVM/PittZU5a6ksg8PX9szfYy5nZcF7hgjg2sJShM/3CDtvJz
JJStTQYFbAqjZhAErBDPuvP5xSkBR69OqsfYNR2ge2w/2Kmn8Q9PMgnZG/meX3j2+OudU9yJPbjA
0aFTs84DZEKbW03M2k+bPY1huTdl5myGxzh6UjRQ9xxMQ4VcS3PNMKAkvuKnW80GfPs4FFsyi+3h
ko3r+RTnV6jRXm5b3ttv1lJWnS2FTqYvo3XUilXu8NdsbVsbehX5vjR4ooO9IIRr2jXi8osZVLRf
1ftC2TnACw6iGb99+9AZkJNzuuPyp9ipn79Bd8fDwuoyJDZImcnQb6NjcECwdM4qNCyls1IDomZt
xW3HSGe1Oi9emrAN2PkyvoYiFMJnq/SlrRv919zdwtUpRrs1Sus4Riy6505Cz9GKhdzrttxvqGKj
A7WkJf6Q1j4WSRExSPhiHhO7MugFAKw3xOmnJcafcSwiezMgoExhQoEBNvp5LXSgO2y2IE8qnyNO
LTlTAP2s1sgYrfz4aMC51W6VIUsIW4kl4jR3bDJpiKhj1CfdSXB8143cNbfxFfOKq+GB710PSlty
+uf3zaV3UX0dnL0cfQByhRYKtYqqPtYBc4rc9wtu8U+IQkzfg0pwPA1tNctPL1jxueX542IAhuqu
hNNtpdoHmm8mAxDS1+QEbZaoqXlBa93n5yqc0DboKd1FbMc271w7q2fYFxuXjJvov5BQN+4wpRqJ
y0mJYIK2gHTwF/GEiHykECIUIjzPAlnZMnZQNh8QHXi2YJmD/j4j17HzK3cLuUWHa2aWn1NyFLJC
D2pMCsYri7ewlpdgMxvX8SApUuc4YP8aqzdRQNZx/NshLK6Sztl8y8wqW6CBn32Ve+fMgnfipGHV
2jUuB7wbapyMnDhu02MLr+VYxaU2THYVmVb0N3PSOLpaOMJz9N40gtI2YV0K6/iG1kH67Pq/HPt9
mATmPCYvrRqPmh4IQ+eB0achE6V6JaUTh1pguORqjMeMWmp+cEMF1GPsUKyTXWNSAf1hFPM7hjHZ
l6EBsWnEg1tNTqUYoNGYu/gswAha4XIbb3noEzPSyv8tuF6KFxI2vqd4EN/rPT5Xjr/FUJgksLHH
oTDCEuoGE/Y+ap+OBe6nCCgNJLH2A3AwxHZ/uCRzad+g8zbLFAdABZBON3+gPXpCc5jbZFAByy4Y
xILk/q6GphaTVfm9h5NXpeHHVPbvAVqmn6Sj1gQzaYej7xXfksJH+EJxaKj5FVQVl66E1CFeasz9
hsjm+b4XIU13bXp2ATAyeI25/XKYtJiHjgJ3luWfWDWRLFPhY8uCG4TRxXSw/cMtAs76kYJd4/b/
DSTWrLCNaLIMtSNiuU7RzeZeYlarUzcajU4GPF0HUnMjqMlJ+bdNAq0Iz/cJBzJD+X7ogViuaPBo
uLuRGDqloIGjNTV06bPmpu0oA7hasTHjoH10JvxnwXLaDwPXFmGoxmdZUThZXD49+gLC9L0wgwN6
ZrHy/6W4+giZYhkQAeqhpT2PP60uhY0cO0Sp9R3rVs2njIq8K88mUC5aLUmXgnXANSFriWO6IyQX
RIIyAkQSeWBoMZ+XK6qsypx6+nO2R08rKkvRGLehNkBZBVtSGOHZAETA6M7w4B8uGXMK8W3ocphP
J34zrVG5KCX6MO8CVc8RVPDUxf8jdTkEYWRd8gUYmw0fw8KHI/CRvWTmIvBrqno9ln/ihs4GyPNd
DGbIqFphm0/juJtibsPA4CXfaA6GzVG5gxzGwNRC1QAjNBIIVHUyrmE6aq+P7H/PpMHlSaNqk3Wh
BT4tFAQTuwWEMg9dfJg7WuK7sxhS9VnjyCilUCVvyVra3g7oyeIp8Exa1t4vIo81WdRFKuiO3ktz
ZZdz/EukMnvMcd3j74x9Eq3AN41LtquNW5Lqw+6L05HAY2Efymghki0I7xWC0YsaEX8Xq+YnXyjH
xYq0vqj4joAkIY0WkEc4CK0p5972ynoY8vWvuB1cmS8aKGL18OMkiB7g/I9Cyb8JOQfF5OuenSvx
SyB55VvxyzfyslmISLTy1cGD57GcbKgO/MxbvVCqgV9zB4blmDl513JFCcVX5jLnF7eskCA8mkMS
HE1l8ZCFcWtxLWDTX6kWDtqmiDFn6CCdVSu9X4W7NINW1OjrwkgSYeuGmpEgJuL9OdXLSYNOF1s+
p2NYgFXEjwPUjEJmWpZ1/rP8CV0eXSe/nUihxaLIpZ3sRtFeTo+HOq0RTdOemYMlrLjXpUhtI5A0
a8KeN5pDtpMvEPFi9nVh6nmHQgEkInOBibwnXP3VNCiOW3dWGIQRsfU1rxr4CR6icF4nRb1/zex7
4n4+6IF4uwSY+hi3ikx1Kkj5i3ZntgXO+4wGRtyoPLBXYQBdZUeulMNFeAMNcYQuXKGXoexY4VCz
DZ4IVAAZKZPdee475PSytxjn+nQWfTs4Y+/aJjVyB70NEk+NZBbeqVYepyGku82D9FA/zvsuTct7
UBlF7KafUL542Wurbgqq54d1MFR/tFLnTw1gENt29BbIL1sl9P5i68wEfgGOl9S1Sg0yynnF5MNt
e08CpcCaRaczoKgLodfCwZnzIKzgR97Qbgm5oO/qE6+JkWR594tYDI+NsCuOKumJix4HnO/unC22
k4K8g7xW0Px+CZgUMA1MLB3yNKhhUzcA1OT+L/5SzDziKKNRGmWR/nUN9hLrcJUoEtXe2X6BDhZX
G9jl+ZNmsdn286Gvktzta057qn6XmXJTesJMdaH9wT1LgJBh9Uy0KWuA1Z6vZ7Nurx3NnRH597Nw
EQE4eoGK6svnMZ4ncWbE71tUD6gRkGHIkhCr3ppthCpvgpCxCy7BYscV1MeIgLgmw2yhGV5tbsuC
Kola9c0TrZVryuU4XhLfYOqDLXk0fNmaG5vRp1YSjeRrADB4aLawVrHuZRH6GZQkylgtJtNWSTUE
+9BJkuvnWlhtDeFb6uSVgJo6wNEopeWzKTnBqk/gxgCYiG/JuKERZQSfqEW7Blt5Vo0ZSMj7b/FJ
gfQ8UsTWs9UGKEF8Y8HYhwrcbL1PT6dZbmrmO+DzrW/V2KeF5+jcrQUYr188idl3uu+2nCzbXlBa
HOOfaxfK9cLjOL30TgNqxXjqLg9fHbJsLHrEIEfpYd+EM4ryug7nl2pltC+rSw8iMzpdDBbuHvym
f+LMUmiNA4DkJwUY8GrJd+7Kp3GtScMszfHsqtdG2l2TtnomvJbpENEx2Br5EgZstbIcny7QKc8+
ZmQePjTBxkaF/HwH1Syec/oBZb7Y72xHYI3q0DXLCcnAk0cIXvfnxacXq6HGXXSpuLCHSB5/b5ye
NB39M0YzrsSILKbpS8ZYES3ZgCcSL7sLp9himcqWz5r3k00ZcTACjJsClPfZujBQTkCfUz97cLra
SKsn8IcUVTMbp/wpGu071gVO7HMgOAvroi4pOwnPDlsE/QoDimzGuzpmvnNpq16HyvXRp6/kChBv
ga3WU48SD/vlf+R0zWeHEe0MxOH2iDFlfAQAvJksXWjsMXzc97cLu/9j5YqPruuj12GBtbPTpWcW
18vnmHRw9q2WUU9CrisZ4L8cS69DwsDoo5HajXeR9cN5lHc++c9QDE8v52b5+bYMjE/SC8pZ5nCM
E3kiDNfsgNyppIlSN3A2Qgjg8Jhg7WWWxrv/PfIeeq+0XUM4xA7pqpgaMwpzJYPEIAdAUMmTkUE1
yjbgDuy+XpHAeeIGeKSVTTqQvysEdO+IySvycaEAmr1TiP8Bbe8yGSgRsQv57u8yVnXpwSOrfH0f
3ru3SrWeb5c5dRm4VZzuqB9//6Q4R2FHCrihuwPv7fomke62lPezmme+LJyDuCwCshz5tq734GMN
uwCUTvsF5zL1rl63KUscCl8AJUHExQGGtZ40RgnFmJ7n2Qtk8iCNwku0MUBZkdjZLJ1nqo3DFTfj
VaTBIEVLZGqhmoNt7kEqzUAURld2Q8E7pe1HSHqFbhudU84Ms2xmViaYAUdtOisQD8FHlkLCh0BP
h8W+5itFEXqp/69jB29oRCTHxNbBXdbmiE3xXYTuJKuL8C6DdNbaBCPNp+0ubiR7rm+YMcpQ/tx3
C4HHgFfzagJg8daUuS9F9Ee1T8f5SIIgGzXy9VgxGXDwJFFY6sF9w+x787S7+3ESy/ncSWvryI8m
bHgPxNU2VJIt82Ce8+Ztfaq0z3JOZlrJmfAOIBkA5cQUOLtcYUmblpljUTWMHGfZQi2DJORkju51
JvJQcGX/+nV0EWj2fx35/r/82AuwhHTcUacEfZdjBzu3MNErnJYBdJLr18AfdnqwrNWWOQyscxGM
jSx4RvEeLgq79yw271UFkukhlc2WgmQQeRy2q8n3dAXjGGk+yG0amPWqhaDzhnBzqBvzPi88xrrQ
JoOQGj/C8do1V32+uonJcBHtVXa1xlGwksoUo0hSestYfOz8+iafkTbdpS1I6DtqrXI+z4d327eA
cQHJKGU7mkH133FP42LZTgiZY8BXqoK+Z00qNTqNPGyhfAqiaPCeq1p+ZKtqEIz80JuuF2ThG/8v
YPjIw1a7PYYTZUyBgrvsCEm7hFoWC7lJP3koYQJGXjAxoIPGMa/VPrQ0vYeuHrq0b4OzE5GeJ0+V
nujYxN0VeD28s4bCF25COwN6WiBFr4T+9M+nZmnG67j387F9Pb8OlSEHVnyLUDYVQy5X7o7mzKGo
ZwzlDXCx7vzJD4Im3Ws9PwhW3jdWYfARFJ7X1ytAO5l2bYLD1o8EfyTUCuHcsEC3C7ezhQKgD9+D
BhnAnuHD5LLnGHzFkquBicVCU3Gyh6kezap3p6b5D2FS22v2Xum81NX5iTYucz8XucspDT6FZzXV
jH8/tkea2ajisVh/H2KFTDtR4HlJB3g5JON6gx9FfOa2Ff7rv1+XN4//mX8VNSH2DwaVaYNZlBPn
ODa2iWjKfX2g7ACtUaCzxEsYuSIhts4nmdcV0xXdf07FlRSjE5jUP/42BXqFScMttlj6IWQ0EeA3
w8nOlJzsPnVxpIOmWvL1L+vlOL5d2Mao9TzjGwhu2iS3omdwXUVVEpmLaAobo20ttCJcZBDIZSvb
cb7EsPsVuvLD7hNWV9nv3nD8DYICCnSqWdA2nAG4GoCVLkzzqRIdh8HX1oIooK1kELz13pLmhIwD
WNXERqTYAX5YHcuyNo3PyISdEUGoWay+cX5TGLXcdo8RhY3ni0nOQjxto3HAq9jqJZK4e7hmDRCD
BXeGFsq0msSroxvkHvEt1Ouy2yF0v3Zsq2OWDG9tTepdfPJfjex2lstB4xthjuhmXolsJUnSmyF+
t/Y94rHyr6Okos7VHUwR4UZsd/TqEIR+T+YB7JmYSlZ2LmdesB6jpYldgmF0GFrv+fz6+Y6JhOb7
2FUtwozlr1Ch4xpi2D6hSK6QFTjCpTzHK+08muqpSPligLdIy6jX0hQMCv9qvGHwynbvwzvmSLWn
wyn+mtG4c9PwOHXpCk8Nh3Tr7Brfwi/httoo0GyoZ4XdFXf5N5qHnzmXOHhP+k/brX4GlsCIORsy
8aVsM0pJCzsQt6AhFYuHpEAM2xyDW0abOUFGagxFY7AQIGBcsYyzrbgFnvJpiTyEFQzvGTX3O+eB
Grxg+ZyFYIMMk+F9MzUrhgFfx2HzwT3UCD57OLRvdPEK+mWm3IvFjqrbE6h3j+wAz30p8i7QLdLN
qYho4RQKsdKjwpObufVOTsBfSJidXnJntjmsYSAb7KOSCjX3zjBYlQOeie4WAjzc2Mco2fhrATB4
Bk6e1TK/BUMooGBrnhZmHJOuv45Njv9aOGH3Ev0Fcp1P0c3264EBe8q1evg5XcSA8oO1IAhfeP0y
jYyiHV2mK2pev+4lwi1B2zOlB49UGyKUYOIHTBtQ3r/TZdk7jA7RvDPVpa9kknToMZS0saXp0yPs
iEY9JPvNA9/Szrsmd8NRaWrs7FgUG0jjgqWgArEijzhmnFcVHRz44iXmVXza9s1aaHxCrIdVzS4k
6AmsTIiJaPgKAuUG31fyyiZ6tIX80b9XaI+QKb9vUtVHDyabvaX0C1yedD/oGW6fJFwPsC3fRTDL
eamvHx5uW6ZVNesNQEZBX+NEXAfey3wYguhjq++uoKJJyra+wasAu/DLJ1cnXW6NDicFGNsBNFDX
NT9UEDzm67vWbQsFUtxsbSGwKj4oeFF8WHrPv0l6XLW89GJ54eQ/btcDMtlFWurCD2DVqsqwfzkh
5uCWgR7ewGfDtunUBkBlZxIFaAAENO9NAaJe1UoglWHhPWDPWrlqZ0lkDapnCDvdRMmiNXtkffVi
VcPukmRGvQZb8IrAOpmRdpovtbaR3M8pA6pTEcL5O4wN1Uw8aT+Eo/ht85gxZEe6MZ0Z2bbjdUTg
J5rhP6zZoFPLPF2ZXAiSU30FmcudSMt/2LE0x3ToiGASLonTngaElrZF11imkwgtONxn8wNpNqqb
5lrBOlJCvmUwha8fSUFZIx+OVxVnijYZsCnhg8FhbzaY+FA0VSZWFCfRT7l8IaQglIc7fV2qnym7
iAXLHVaswyANbx2HmYmGUt266yyWBbfQPwlF++yESiE6F7QEzEkj8/Xci0PKVhofjXkgP7lo3ZP6
cIHB2RkJYLFnf9lAlCBdShKaMCwH/FPQW6Bdy9wp80zEoKt7Sw/VXAxR/eitzL2BWZpSxVxEMTa2
MPXJVvRL2NqFhR9WwwL2SUZL+A/JKP5prV/oWuBx/F7CpbzzHqZoi2502yLJKdzaqoKsJsHPgJ96
mlBxEaEUNecq7phU95cv6e/nWHfja2+FsdTnd6qtUj5g/J7LLUqNvChTuqGPqQWKOXcFXdHB6hsZ
RbdnprjzMXRsNaEyHFu9qedy5NfLf99Q1tgxfffclbfhzXZPG6bIt7N3xQ5RFtzz7l0FnsrhBSj5
U4Rz5ybJt1ZaC3zcnV97fLO+1fXJWh5LQief4fxxPFuh5EfWnko8/3j17Wj2dEfCh0Cec2v5cM5f
k2ns3Dqgmxgy006TvCW2l1ErVcSJGYwG6yWRL+YHIW12H0WuJ3Jo7i9QV2JnirBYCXbOs/ZNYsLm
sFF7Utxxv+daHdSCrzJWPyHcsaLhaQ+TDCXmfYSiu4adkTwddgt9qZtdfScPpkEtoy5iYWSqqYiD
/8THDndx2otBNcsRKoFwUacD4FAKe3eO+D/Wmiff4sTsgDktHGYjOJZPbTNF2kDdHMsHMgFXBc9r
VhSKglqF+LXbpHMKaql/1bpiD1DxY7yUuKvbgbSoL8Y0B4DCaec9RNZrYf6rifMXfCeQ0kiW2c5J
P0XzO1ny5CBoIjnNtda4O0i7blIob+W4n64CrK1vL8f9/88UxeRN/VlyislOiqtetLKrr8pdOwwf
tdDCgEWhqIKqg7vgO1Z2N3+mVd764ydTCxoo52wYzQRoeKgHv0besZntG1S8pMnkJkbkLslFxYEC
N3YAGagC+Oy+nokKtIBWBb9EgZ7rkXsENr0zYojpEATW4T2JHXTzKm+nxsZJp7JvzdOZrhh+kbKj
Smv9TBcf3D/b8ZdeHRacApogsbCF11IqHjUhTlPL7ljBo+ZPMxxoF3uvP1kMclG9AQOOap8awGLM
CchbeRsaOebaxOFJUCJoafrYngZ2L9qlgeamryLasMeH55EIT4CGVvZUWkuWKV2g1CNSxf3anATx
55EZEVvZBS0CinL6UhIlSOURgdXrvaWuwgDKOkHxz8dfhEZ/eywnDFdzqY8hzegWFxg51vP/w95S
0Jg7+ose8PwHFVfZjmnpMjEzmBk2WftGjAMkYfey33QYwxk3rgZVhD10UMwrwh+z3VEkHjHZTFag
yip92IQ6/+N0xGZ0HCGxJWOgBmN3DDN2QUbKUPTzPThe+zHXctpwD8nDyJ4d3L21Rd58DG2XvyRo
f3MK9OhvK/prA9r6x1Od7dbGhS9lT3CLHkOkfS+VqBVpZp7+wqs7heZozwtix8zvrC/PfIe72F8A
N1Ru1zF+UOdpefAr0NpGHHsZLRWC70rI7JqxGCssot9shwfGEM+5sH/hNRpvxRkOAEIwz7WDqJu1
PacP2nJ25srOaj1RP3RV19bb8yPn6dU5sstAhStSejiYPBNAlY+87qNO5I5YKkN3fY5cu4XbtUb5
L0ph08wFbStS6VWJBz2qQc1KYI5oJ8EfqpOEnNHurj/i5BvPIKx21mQN6P1Op1euZ9IKkInXYGHr
H8ajhmIl4LffGQe13GCsxfzRRDHssVmhyKGvUv8i7vD1QXfged/WXyklz4vJxnW7xT02xJVP6s49
/aAgJKuYKuOpnpM0s0bysh7WQiEhte7fjvR9i5/smbEqFy1C6PNkO5JMvFcuzocRrA9GY2B4A9Hm
QIrvzwrVT3V14gjtjhrO4i5cbaE0693QgBERzcQyjYZOzIKb9t+6+faNLCNdUDN28V81YXDDAjKE
TmgBiPgLfyXc7QFBkQfxrZjyaLV1SMZLA4eSbofyws10++zryuw/V44oGMiSWXnQvFvRFLabLYO3
Kd/+II3Mj03pg95U87Co7SPqJFXyvMH2j2CviTwGcOoJChEctx1KM2UXJ6hoKNt25R0BGMF8atfT
GtVun3of2GB4jfqE/fFE1QIz51jI66JL29Vj4gRfjjfjCAaJ6hCkmlhIDl+JMryUsRXGaLIAG4eN
9Q0EKy9ALXcM8IlpDBFd+2WPSeqkivOmpHYVyTSq/J694cG7Bbd//73N99Uwj//Z3d8qi+9GwDZT
cKE15Jax8ywRx3s1kFrlLq6/oz5JOelBrQMJEeR6yaQjTdizYgDhPqdenRxRvVSQpmO4z9rhlOZX
PO5nkLhP2AD0AjXe7guW7YF84kfTwSIWPmgemNg3RFKTxw0w9rRTfcWcVXNajCzfMDhHM1Wcj48E
UdC5ozojmxG8BpAR1+DEfBl8YF0ol23QB04qJbVQtBNnO9sgek+4lK/rkhwwqUeueXaX3Ail+Fun
1GjTU+pAtQ15MQ7KsHGgm3c630Z1W0SSbApV9cYjbfL3KNwCebfLw1yNeKD5G+tXzIFQDhUjAVmW
/foetKYIqQys2XA0Vr5EEglUyuY2IETkjsQEXbEq1bQE9xWVXM1rwFGrndWPhQpEPdgNMKddUX/e
ixkCRaaBQp+h8JnmwJpndili7Vthtk9uIhsg8fWZMxWcTsUuoNg5GLJh7GPftxLWBchvT2/tLP3P
tsO79h5DUikkn1By+b+lKWmxwxzNC4jYCPXbvbSkf2GVdcTwfFtl+lxNi7CHOf+2h6Ceq5cl8sbl
j6pyUCmBbOkuWKg6Um0hw4qcQoPbhAPDuuFLVP1H8k3ew9Ie/O0x+9oIsN5gz8RPio19Ejyuwq+Z
mV+nDJzQLypXKshFdlqDxdfxJcC19QiJSvmmN+tZCv7yPRDN1l4O550jX+JnKeX+IagdG0ryY/HZ
0owjfHL6YKu1K90fpVWPsAicgqBsrJaCOxeTvT9ktrla//LwrwEVhKnIYhGuTxkMemrx3VMX7BIk
Zyfs1cshfnKahslO8PW3EDDWmZ3TFP7QCzg6xuwFeIhOo2T304UhekPBuPqen3rVZjuSOPtmv/jG
zdgYZPC2tccYWtknqEOsxQghnxj/8hQpY4IoesZ0JHWCzsk3IEanaLxvKfwF6lG/vMZN52ZCfzIp
nHCqFhxe4Ys6n34WThTnvU4xH2HRwqGpiiJReft9FDQ37Zy+Z4p5UJ33qPfBeKgLFNDs3HZrrX7s
8nJPf7KZsvhRxnIwnDNl7HMk7Zec3mfmqnlAxiboP1L+4hMohXcEccX6UCPbjGZeWlzvwPoNIR4I
GkFVNhY9BlQH++U/4cQMFio1Q+eXB47xtSlWjdYiJdf0U8jrEs4vhL1iB43/G+IjE+ioYmN2n7dK
60lnfoY1v4TDB4Kno9jSAR5QcHQPYq0rpb/yLllUePgjSiP1RB/VUIa9B3M+PTQUdmyid/6GABW1
kalGRNoyJe/JEBMkauXLSTipvr1X55h1DElkNOE/rMni8qXBP6xq4qD7cofkVTvXn0hxr9FMJIvV
fFAN9bB8NBesvn+awqjpn1JjXtQtPh3ojzXhTAjBrkEDModK77I38At70OnJkqRQBWnSttuMJTr1
3TKAlbhTvvActc1j7qFODQBcQhjUy2vP9XZ1A0STdR+EmOaSjrGuDnQNthVJU7yGTwIrnpyPngPE
zkM1/mAHRAy8J5PNQnqCieOXH7OCfCIe+O2SydBkLSQfdleI3KyAAqXWRd7fJoHJWE9BzwoqQcqK
BP0RbY1/MaLoEs0Ue+lXxLZA4Xe9m3jk+Mnu1lbLQs5+i2CCBP1JkzoSzvgR2LeWPR2Hb4nAESBa
SAzng7fJV0G+MKBUaH6ZX52L2XEjHoiqhiIPIc5QFNoDf6s/HPSFdtgJOxZUFhNRPeAJqt0YuJrt
Z6mIV0gDQ4S08kEu2AjE7un5ds4IC/iBo5Nh7Ulc8cPfOifT0f2jPoc5v6bTV69jpnvOpF2IP5FI
fjrB08I8CfRJDgTtinU1dP/hdhKT2PmOmopIM7GRDcF0jOwPltmeIqegxdLAJZ8a/I9QMq38X1wL
LG0HroY4tXJRgsMgW5DdLSs9PFWPgcba2ZaQGD0zJW2TqW8+JSZRQDQ8ZWNhDW5kQMBL4x3eZGbc
hU7/NUVBX33LM6DJ7pJAp2ZHvsphBDTGoAR31BO5xRxUDs9Qdv93tfFaYIJbqTBhf27zFnAorE6b
CJDsE/hcC+tqgmjqon8Y6JTZyA6aGhci1odB0klxovd9GjkOr6G56kjE1M3EPduJ4MdOvXWRiX+G
UO0YnbjviEP8GTg9dc6nlGYmqyz6R5q4WAMLURZxy00DYU+zhUuemL6yRvnTtSOrilF2TrR9pe9m
PzB2fIIWSWoNw3x+PbjGNUiAJxEqwzeCFrXzhC1ukcnO04Rk0iai1VDdSXSYxREroI04n3QOHuyT
fX4yRd+S8x0lkum+FeyzztLcQs2NSwtILL8c5SnXpKCro+fVLFG6N2SorWW0hyPHDHyzMysuVBL5
pbU8VyggQ39QHx5xIlpXZiODxuH3qY3tOiHb85IiDzu7hBRvxQPiD9PFocWRvCqS9e68cZJ4zVYf
vTx78/IG0oZ13Kxp/vdRNXe1zYylYzV68emhNGtEa1dE1YP0WevkaQM9b3Z0h/vOacIX6ZalGUeT
3mTu1ShK4noSxOd61FWlSZiBpCWBvT/Lior1cr3XJMJ5PtFshDNTNQUlHg5L4eZVtUGE4EU7JJMY
O+XX6TStlmXiqApDC0vHnOgNuvSGrC9a2GH+REDLraKTIGuHyuSG4E1zLqrGMWpleUyP+M/hBC1o
SlCROYs8qiY7S+nuTdrqqyExBkEb/p+FsZo8QAKQI5gYxvziE0AVgiagb3BfRcMhEZAZvary6OY2
HM+LO04GobuyDbNXfX7SfT3A3d15eQVqNG8TVogJvR9Isqz19Z6zcSY2hjgy9ScJ6k2YF1VFwckK
axyM+neJCP/wQgxXxcBsQi7iM2SreSTLikJmLMJvvaa2GAN3p/LZFwTbH6i/+jYfOwc8Ko4LgBvG
bfDH3G3LSLWK5LJogdJgVbpTvjFXU9GVa9q5a1YpB5An737euRQCMcjZl05u7zIU/DH/p6kV5wQv
4lyTpty8bve5cA33Mq1oJZFMAikWNlzaC2y68Z0m7hOkFkAacWw4ztkmji4P3aefoZgwX1Ze8ibP
IgZVQTr6LLOMyqYVJBibjCPng1VVkGWWJ4Ai4YpdRJzLoEj7rW7CTiYqqrFMjupAbZfmHQ6OqGlM
sAK+tuYXqdbz75UKPMiNY0HVhFgLPwdUMSa8YEyjtVLkWYkwtNooQ2qt0e1MvU2f/rg0g3/HR9eE
Ps0gQdBo/nd2XaBcGYERhcGHiIfa/DCmStyYHWZGeOWFMQhqJOwiMYczei0JPz/zNFAvqpHuS6TO
GmvZkaKsILK9OoXGhO3zYlA3bV25BvOLWAdccNZJX+9oB9mI82ZVITS7ohAn9TanAvL5ucv5xm21
c1K+n9p7FDB+4KIA7Y9LAG61vYPzU2UShKwAi2aXc6Ut5iRgZpbJvPDSSAA2Vl6STfCf6Rw5ua84
4tAaNUZXzVcYRjlNWNfzia515I4Oy6YH5CRIRphN7MyPC1/Hli+U8UYEjI6nkmKbm6y/7AtCZyMA
83M6Mn9Wf/9l00vQNNZwdGzUioKjiQHGTPxHoFsX9eWYo6EnvBwASI+iseeuQC6cf0ca+Z5QKtxj
HMrU59rFteCsfV63nRILhXeyZdVBdMS/P9GSzR/nw20ked3ti6J2QAAzIA63lzoW1aDOqphh/KVE
V2d/fA06+aFtH/fdq3K0KrQByfvw1T0DTKb5yaSENNTkIUUiiFS08K5asNJHmLclHTXzdInKmufC
iLLBBGGr3R7/iSyJ0GhHh8s2NaWV/fhLNjZkDOKIvrnTvs/RaDiwbGP4ZvBuIyVO+cMi6aLM1xmg
TGJbFIt9qNkKtZUHVPXp/iAG/M/SmUynwEB+K08EpAbQmT+04Cvyw+F9zGK5KZ54k5rKznMDpCwY
AD2Tia0MrqQWtO3Gu7VjnFbfX6xkpIzzh7cBxLfCymVFuETQKSoCSMM51ifvUBxbdj+NK6hczNhM
6N6Z4klT2/3rmPfX8yzapMqYhw8RhPFgR/AAqOC/wEcn3dHr2doEEqOxyZreZWzCZVYS3Z4asnCP
DUOH7bK69nDSrCw6B4MmBDouVhHuyZsb68IuYHLrNsDYmmxkYGxMpex66Oc1aXdftlKilL9MoBRW
2pyAQbUO45jF4x4NDE/rkANKEJ9+zQKrb+8M2tP9ZrZ/cruhgdy8gdvschdEijS+aBkQc7S6CC5v
DNQy/hZyov+qfKkeXWHKvgt7BZkjTNryoxH0jI7ouVLv87kzvgo8GpNYcAp/6BnVaXJ77HY4aQ/o
gvsPU+Gt2fb22yjjgL0DOnMDhmrQu0GfQVFQzpZ1OhAnLQy8mEpPgPpV0+6F7h+NfJMeKBEW9rbZ
MOSFAcfuEaLjVz+gN3xe1iC/EgJYWOXx8rpx1/DDDGiFCNJaOuXEI8YkFRa39npUAJR8/FYxVOKa
oWlRK9F+9kepQRlOxyt2khyMiCdMviobdYfj2ixj/OwtLkwxShmgv4xaDrkyMsb0xfJtPWFTCSy6
A3SBR4mDDPNICmzdIyUsorySuuJTOn7eCygiTBPXDnsSzf7H237unmjhCi+cRR/rmAGNWz6lBVPI
PFdX9O44VhZUY9qz+IzsyGo8/FRlrblJPFvbxeEnfrIipEbPsNMlpR/emrZ+440CyBpRHpqDchI/
h7FOLLIKvMLZ4Ghb/xdgY+Y9OSBVKg0r5ecsBpqhQhZoiXxAUlGuDfIAA0F5Oh8dFInNoI1U5QGV
GqAjqIM7vO/s7HT6fVzKKCXaKAryuQgCULGM+X9+rmy53mBG/zqkjFaxH6sL/XGdawB3jvzHKnQl
OJ1IoY2HsTzjhGt8tpl+pSUT/egHBiM/Rmny2GQgZR0y42THm0Mgf7gxvgJjchqESQYoetdR/GpI
TEZa0ED+uDuvaQUFAHj/UAc1qBoaE+p8k0zBiXEFpswgBBX1Leww7YNmFslBxidwTZWWcy8ipSmR
/GC3w8hWrBej56MhZS9PWOqBaw5wwFTe9gHU1DWhgxrFh8z4ESP7LffmjJLQbAfPdeQ1QX16fDx9
WDGM8fK6VkMHhnvQpi+yCaJdd5oXiothsJ/yr4tXGzMaHvoksK7rcu4RGSSYpa0XJI/SzdI+0EHM
i+yCHCLVKsVCtHLqpwOnCpDZ0bZzjBp1Cdhpeq88kw8xb84FItemdKc8fK8AlD7b7Hxm3vZfynox
LFA21bYsFFT9Yy1IIpuZ4IRQy9+RyWVHpUVTI2gQOyOo6sbEdIY9UIb4qJqziNu/clJgFEmEA8PJ
hMv+2WKQZLAq0yt7Bj1W0iOWhgNcao8DarUoPKudktMp+gkcqBkddMbE0Gad3yUHIAwcrOnsYyvH
4SR9bV5yywxdmkrotEDHj7g2ZtUBhfieAYN7/Z+xxcggN31N9tAXiorVqRVR73th++3EQPeBZxXQ
ZhD1Kk0lLrkrQLFZg+by2TruvsJ/TKMVOdbmciK+Oy2ztNqvO8NhXBcpuiNhCa8+rNfm7/X8/bOq
e9qzINGfEqESTDI9WXQDneqTvGRvg8ccOtHvF43SAhj7IpRhPvZ/4wlIKhTEGDH4TjVruN4JWgTH
huW/0kR2OATuHl5g/VVKmJxCRZjZu7ThN8l1HxNZ1RswoduElaUc2rXilGxa20roNxImTAKPQi4t
C3INHu3ectL0J9YlhH9Ck1q+Fkk4lsxadErnTx9SaRx48xkw8+26IrvfQLiM3gsRCMbiYgkggX1R
zmf3EizkJ7v82yHSQMlpxyk15JyifdeHhcT/wXwFg5mltAytFQKuW7fs6xDVJfCcVdXtLC2BGiD5
ajIdBIr4o831bVzci/qpmwKbcW4GddX/VuzkOeX3H4J0eocifGbiYmeRI0aofVakQNvpNb/BtqC4
MceuCCdom/XAy++dEEH49Ioxd7YNTaCHoQswZ9fFH00KYriADvmyZZ/CDZAMCkfjgiVmUDOLxqbN
nJwKqDo1MSMqa+6y4q3/VZidhrwe2GpJlaITprNdHoTMlqOF47lzcwuyxkVGhYdPh730W2TRLV+2
5iP10U0S66i0l9KOKrJsk3p3cwZFfcGxE1UwcGIEDO2I9iS2f+ZkjgWBWiE8fH7T0z4U1ocxvCY/
i6+XD/nzqQVJDmZgJK8ebn+j0LcuGgf+cetJ+P5JzkW8sUurYC9/FS17msQK7ld2W2UJ2gLwoeDZ
YmiU+kvwLScRiYwlZz2sDwEF2WOiF6SMDwh1EsYDmxbyoXa2hD2PnbJJa3dFp0U8bZ8lTD7UMvEG
oh2grc/6xQyfeL+vpsNgTiw4ybV9d+oAAgY/WM/rmRPI16HZrRmPDpfwaV6vSMJsI0tzKJ72wC8d
OMD8FLHWVFNjRT6+91qJCvsfouWFXdVovGesCeEs3tsJurcWRBidW9uLetrc2hm6GpCzUZS1jrbM
GztsUxRh2yshp6TzbFlBDMolaWJOBf6G9pPTIF2cGEjEhp+4tu0dk8mt8NdkSqcWXDjgDEcz2MSh
/MVyZBTkdOc3qF4qfZohzTEGlkFtxRbjmBm2KaPVzg6hXY/OkBUOK7/yyZuppfTzZo5BVz7WbGng
yequQ3UI8sDUmEWNKZhBXbCd48LvCLcNa1FEfp2imeLfpe18RoMK4NUnwhJsNhpo2hqqTucGzHZV
Dv1C4EDXykk88ESDwRfLciRVuKxXb7EVs7Pmh8a/Fy0WTu1j6ruLhdlOFUhQZyAcn3KdMbRN9LmO
B5SGPX7V4FY6q6/QsJKwaQ5G9vAmwzb3ByTUzDkPnwvz/PW27ortd46NDTBcYyjrhyhRSERWhUUt
UzdOObSvkq1S+ziIk9TM6oKTRlaf+dhQYP/wKmwAE7bblIgucvgfuwcmvEWRbXzc1VLk9yGGPloX
NQBNBmZXGSJUWCOL+TJ6YcpKOFl0U7U/WUaZeHIBa+1XLRfwF0zUXBQBb1UVrtpn3d9wlz5q3QnC
3QIC75Bjc7ZbyAUJTXgxGOpSOx7B0oBIUzR/jRVLvTRgW2C/sA6xlUAcLpd3OPYWUGFgoKIoBGk0
izwLxhfblPecMQnIs6hEOMn4aGDNtBtZ1W73uJmdJe4+NcJz9glW+eUl9wrNIVLX0O6B6cdHsQwG
LUGPcD2Cn6G95RM0wv69chWBBngJpYSjfYsy1Gl2zKkXNCsf9EN4WAA2mGyZ8b0NVej9fZbt4BQb
OuVsgTRXCLRsHsHyESF/ikJxX478W0vjxDRmkvVWejn7hn/kT2ls8YQp8h7wBSTxGxsFclejLygU
ZLkCKHG3Awql+HPUMpQjk0piv2mCdEEYfUYNjPyIXjaJizHECNG/KqlDdDkLmpjNpq5YsG+eimjt
sZq4AzLJI3k/3YXUhu+lVu+1sZbp/1Qr3a8KUp4+7Ldqot2Wz8IvCUlzTfvur6ABqjxk1QdwlShp
h2DsOE/P7EeatReF7sdinvVREHrNC/KDBpOPZnlM/i11pCe0cRGLBY+2LiEBmCGeI95gwJPIqO9A
YZfSxPnPYWZiymLh4RxWempYEXtJtQKaP+UQ0aRGuUXquetBVJiHtCJ5MPcnYu+IIBPuPLEKX8bn
pjNTa/ITvw9nYQ3noZWi13Toe2RTH3Fln5+VIQTYzugCbRscnPra952xNODTWd1bax+yu1v48lwi
9pfTWY43Qf2x0MepYRf38nXPmp3Iv2pp2jbMWybv4EacJw06dOfICDmW6chvmGI73Dz4e8Q5Dh+7
J7IhaJTuxXNq8GMn5xoMSw4H1DvbBKWX0nFz5cKuXlAkUej6dBGkDupWHT1Fi6Hc7v4pRBw+nEBk
l6oJpI8L4yz8SKnXFrXgAe7fNKuSNPhUdhvWzK9tal20C+50PGwChe2CcfpEgXjPt4vn2kxzU/xw
vGnxHYNmk4baO+lLHcoC67TQzjwls/PlKggHlIz64Ba85lnaX7C/94px0wLFM4UPQE5o4aqEfGDC
EYFwZMz83LkpFcne7jmuqLYxk/9q3goGO+9zgpSfNcrKDQu7SH+Ou8or4AjhuoYS7tJYoBIpjVmN
odgKDFSwKa8nBBVpZJY+muh5g8xZsDqzUt0kCBjPYp/wANsp5c1JgqaXvA/NFdVGo4CuGGFmLBH+
MFchmMfiQIaEJjmfVeplt50NOt5Tp8fhqoD1F2YWhM2yyQhionBpchSSaATw05Mie++3dAljNi+J
iYeXAVcBMXi4nlJAKd1IU66KrBMQZF/s7dHVcbF8vFnklhIP7O18ea9inc2ZJu9cxnAhhHKcBcN3
QstdyuVtZXbd+gCzzx6/jzJwNKP5hWTZoULM4l/xxO+9AA+KzSLKRmBt/S61F6NEQyOpMh+OVZiv
nrprY/4X+qWbrIhnQM7IzW5BruXWdOxRdKjDkzR7Z+h2lKYBFYBX8D9utm3ZTL6bcUgSGuanbfJ8
bfNbCiyOIdTq0TX/FjjBnnjnR+oqJ4vpuW2MqPa9NUjVQAYkxhTvJIuZQU9Hc+ZCm6NVrYxVzDDo
2x2taH04NA/0+TKlfcgETO/fJT950COqQ6GZykHwCkTOU5lgW7OVSHJV5QSMmBK6VfcMsIPtDGVv
R/AiBXXhmfK7f1jmb9c7j47Ahs3NNUUFQj3JAzPUWvs352Dos138NLF92/pEM4TufDOiy/zHsLjD
pXikRNClfwOdF2lP02abcmxz5uWUydNHEa63TERBgKRtkFcyJP3V62FN54MGPufHEsg3wfPLi7Pd
SxdTHS9zpwqkJ/OeemTUpO5Dzqo2zJQAXXaMyLD8BVDySpOrwCyp+Ak91rdLPG7MeN5/k3iBy0aK
klYFBBX0M2iCNzjFGpHAZUknhKmKrhBBUv1fZLtxcg5Carg0SHUXWUXOvUUeroBhNSyYi3aJb6k4
0rwNRz18P4UWxUOFLj4flJHns+Ydblde6pLuf4NIJJodL0AkBEDPOGIlz78Tv9PpEEjpzolJLOsI
Q3bEQwK7zT3GNoop68K5+T1bfVzHz0VQpKvpBGU4i/72lKbnj17V9ikuJPS/zFZw9en3GUyjylPX
j0073xNNsgt6jyPiur5eF35uuFQZUeCQQncL/p88NWpFY4aEHr/7nmD7Muy8KwNTu+4ORTPoTHfP
fNxMyXIvEkNOEtznx3uJRsAhkqZaTeVrNnBxy7l3J2VtJY6AmE+erJKhCezxVfqjwS+bvxJrmI3I
oY9tBjCaBKRsPrki4X6tqsNkseO/thJUyWMe26h5NOXOvewdACzx8OQbK2aB7RPDGABcqXtnI0ck
lmQy2CbMkF6PX+aPBtUzM2k37j0fy/XYSPfXUi0UGTYF1gNIYdhUoeHrvLMthD4K+fOj/s83taH9
H378Y0SL1hHmiPqdQIhmAIhER6zcOeD1/SrRi7M10HWi891OPpIZfcr1AVTgVmTlBUOlyKkyMQlo
Rc/tUjY/FJDtVewdW4z6/z7cCgJ/j4fUsDumO+Gbgfj5vWIYNThm91tVRXLWE3XIi+BkXDh7c7wq
PUmjNJlNws2McRTntigsV3LNxNZ1vwbUBnVZMKGf4pAglvoe2vWuYr1XFX92eFgxwgGOw4O8y6fc
Mzief3vsbqh7CeJ7Co/82JhO7vhsMleYsIL0b6SE809NzZgHQTPovX8G/23eYwJPhIvcxI1byEvX
AhPWllo9O3cTxtoim/qVVh4qf45Y2MZK87UuCEsGOaUIlORKgEmZbJuzxw0BdkSe3ni7imqMl3JB
LyDkPkqTfNpUBviwEuL5JITuihuuO5+P02796HOsMH8wyhwEyl5YmSLSXItGvuTHO+t/f60JlZNQ
QsrXhzNHrEJvV5QZnN1/ZMJpaTfcYG+0PFX9gP+vj7dbx0lqGzHO+vBjicehBjadYz+1kD15We4w
UJCuAt3cBo9r/1iFUlfccQKf9zZnCiocinHHoM5XaCZFlZAy/CgPcoY6QvSOhZif9AwkSLScLDLK
tTbgB4RCA8+PMydFJHQPr1449CW0heYWT37eAOheGzilah0+MmN843ey41g1LLR0mBZGQ0YjrTGx
49B6AHe6HmG0LceXwrgy2o08m87xC42kCUsLNhI+fg6sx8f8gWMv16nG3v04JgDMpxfRk421J4Lq
pGYnpVUzWB1tcaJwpIZlcX3HJg6lpDba7HON8AgVIzHzh5GUHaFs/34LP+jmcD4r9AOCb6O+Hxdk
dr41gN9K+FV/B8Os64tDVgu9gEKsl5ZxKgYnpend0c0+0egyjxWtV7smF/y4WYRORH6WYOQCIU2i
th/EQeO9wX8U+rJNtqZ+l+dVviFZW1DiA0tnoD7Fi/AqrOK2CO+KLXJhE2OnroQGhgY974STewYx
FOfRNoq4qMu12naAWrqGv4OUwwj/eDUcsjx+YhbCPi4rPLCRuwswQsj1+1wO6PclD71K6ffVVRBQ
GOWoZv1G6sY+wEUC0y8oM6XSaUmbVL4DNJ/aqHCYBnp+kJnkpx5XjQQBardMe0XuxbqPzZ+DENDc
m4wF37eadlMz3KcPMATO2yhlumwHbpZopS0H28gQR9icqWU0Ha74LKUy+zpkO2ELzYMshFioJgoA
W5uc13XHTlpuRDBC6Ux+JbEIFK3/CovdqWZmfdYnnEKU8HcV7tTJmmPnMhOgV4iZypqNBGFM8vHu
tiVJKrqmNCGcLHtQiaQcpnB/zDpCVHxzrg9aptMZ2SXGE+IXKWBQUq5oABuXSza/+R44LcLVJpsj
+6p4SakuuRudl6xrsgS7DxIJFX34lAYjXgWn/pvxCEL3ZqRuxha7kV3Fj6huCMKxB9dip0AxORGx
vjHworEoAX40lEDpYbiKcNd/LMr3+0FJmd7BGhkGVlN3W5Uttca7uERyOft6AKnHqL099n1w+TQf
XdrsZEqkasvCTPm0oQLxOs5LsNAGFHn6OeGb94aPRbsY9j3hrHrEs0B1b+WZlGMVSlLFscQIegf/
g3NUTeDZPAIlgdsVDKNFatn16jHPvRPYJ4Gac8suuM9lMLGcjfR4+9gZADZWaa2/PeJ9IuULt98U
1t3t+HEpLr+sMG1xOmQoIQRr9J7Q4/zLUoMy98AOvqITDpgcjFiUHr5U5XuMEekXCRzu48CfQ82m
wwrvJN+IO9Vs+WdJ2NEyK8ICTu5EtGuAuwURqnSLGtNwy3prhTLRigtrd3J1IS7qf0cNH95K3asD
lmk+mVZ7XFKYbv+fQtbR37UbqD+qz0tkwoksTBSP0WDdP1Cj1uqVyeOQM4BYv+Mz8M6aIS249Vzw
ewYjEAXTomrwqDNEsFmlQKgkzu947SslT/GNPX9caWodEykWewwKLTDPXbJg4MSptEQF3amaKoDp
k/cHUZ2u5/5eT7FvxFAJjb89AKm63q6JkGQTL5rYQ5pKKfZTLROZ95X+m4ZLhnaFja4vy74su33p
XhEInQlLVntjBgxHQ4j5ntElpNO9ST4KbmwgWULtyEc4dlPQcGtrscrXBZYfcew2z7qE2jdV9sUk
n2oXLf1wNTliCHoyqjYSgL5nB+xH92kxjsdNBHb2Joi0G14gWeSUflQXV2PRU15jpHDogaIWRG5M
0QXe/0S95JjJrS02JDopvPwMqFWnZBzBEh19+aRX8NT0Jsofb843gLtvSjzcQvWAelA2bL65fVUK
m4bhUoGdEn0QQ0d8x8K9kvbDEjHpTgcqvFfh1e18qj3vOMZJ4J3mhE8KqFuPwrNn9Llx2r6ZKoT8
YOu7g1yhlYsvXuPXWAw/CQe8pCc79S96yqSlT3Senp8gKOE+sR6a9+InoF2+4Azs5v4T7Eqeof/r
j2zuLc0yHXoQDB4Tvd2fuuYs2Lb4jbNltRsbpmo8i7Ic+aAwiOWm2slrhAVOPMaIQs0EJaVPndzc
zRuBwZvUhPJfLSVG19Wtt0bUm/KZ5PnnVIjw0IVD1gzv/0lnXqkHAJhO4acTMjNK9ZoS9cxfKLB4
onYXXEcrM0KJ7iyn613doZO/Rz0NdDYqw4tQo+9XSSbX52oPuZ5zXEz2oJ67CN68vPf7Zxbyh8ll
KOApsKRlmNB/WFFL2s1debptEAqaDw4f9+8zh4nJflc6SYRg+/TDSwF8Dsaw7yKDfLCXazl0d9QL
mSHUJxBY9B0+S+YD8sIHwovM+iyTIpjIhc2t2ZFkSyW/kvzN+drUfPqNmZ0bGf0ipUGhr/D2CqBz
7Bn+SS2w+N3v+YW0n1ZigejnLQZz49djCjQypDxT9XwAmaDKwjTqbj9NoNmUlODElA4juYHnn+8a
fDqacYOLuzDGJ784xUkv5tt3s/JiiICotP+w4LFMgh/NTfWoHX6fAEAWrWlg27Uv7YJ0jXU7TZ7f
BkbM78YhXdk/q+fDo1Q4CjINA5I7suAsnAeSFqyuDWdMf0U1PgLsFc1WDWh/3JAT0gEGkK3Ljvuc
Uncji7h8TsVPfkHJxTAxNSTtEg9enS1c12XNoa/ieiVP8+Q+GJDAJVqk1gAuqtVJ7P7xBXSkLwq8
FqG9avWwUDJCYgzf9u56F/4UJl+bbPUb9haNg5CzmAqypcXSG5mqMMxUcwOOxrfgvLXa38nygkuz
2y76qRzeaqbJOs/e2T54sbnu9QH/vO8IZQ4lSPvh/Nu2zuCIzLDjZdlcxOLByHaB3djYHCSgiU9N
QXqHa37mvZlMdeSfCUXdoaKQQ8/6Jr3ahIVZhtuuRywvj+eBstMvy0johAPwWfHLvGz8z0cdd3zs
A4rqBot6OfqQ1SM4uJ5sx6TpsrsUQwt/DjR4bETDosx3YXV3+PoWlLh0IhrRBDUkeDWnroKTMwkX
+bP0sUClALCj6JoEKGm+in6a6UBV8Zmi1pwK0prZQ1Fd3/JzK8M1UH5H7ZpVtnhXlBa+HKvZd1Gl
VHKUKc61XCkG/CnTPll2r5RyzdtMGC6zn1nyyqqR4Ci1tgZMApwpvY6swcgAoH897P88e2QW/1pI
Rd5o42mPQypLDgeu8D7Lo2hfQ1p/jxqv7/zw7PYNmrdX2RekSWWYwuqicC5+HPam5pclQS8W6bpq
RxTrCu48CzHm0+GQOQDidz+F0PI3R9ZWKEn3iD0U5WBjofVuBj2ifOjbShqBv4756321rU8j77PY
nzOc9TaMp/2WW9gTlNC4//C3YsEMwMG+AcQ45xfU58z9+Kz2V8S3JEskv2gD51Z4nY02z5NbgbOZ
KxGSeuSh25H/0+QmEstCCcmmGLIoyBMCMgObrXsxQKcQgVxV90zZqiiwi3HFB29bCHebDEzV0m8p
XnEHUGtDDoryFiayrk9ShNJKSBnUazh6c10qLq+h+97JvkXaG912z+YJjeWpRChN3pwr6aGhszRy
friSRJ3cpdgM8XRO/7LNPImpbtS03FyrygWPWTldPVdb5bqHZ6uqPWqKcRicFkaKlB9cYGW1yV5S
ygbsVsmEWuetsdXewu9WbwuY6GLmZW3RFo8jrLCjFYnN8szmM0CyBGy/s64I6ym34tlOIsaYEMlR
UNKlzWlhS7euh6nJVIDUfH5NafwCMBtQQWovMt2phNZeiNQ8Tpe+kXpl0RY9bNhV9wKffkHEgOjU
+2CilEnUMTLy7+t8BhGZ1s4KNmFCSC1Aixd/X4UtwhtwH9F9982c5tU3z7ETBQ7qEDHm8vA/eMkk
7Tylvc1gl/fxWaoB0hZDd7QNXS5r2vqT9yQbM6pnSA4uPqwktm21IJ7fpz2b6wB3/BJKx9vY79jO
Wc1EvxmPbv71vETEP7MU95WsmEOe7U15h6Wzq0DcJY/eC83iVAoqLePjSDj+cgUIZBKLawsaNXF/
mMzQQ/jLKkiM8VRpSiX408LU2gO0kLYFMw3bIqXzK5S4FOHVH+jKUvEq6Ik+oZR9zFZoPcOV239v
YEL6X5HuloOjc2ZfBoxnRFLWRQmywOotVZOWSHLelbWLqTMGAxHITkqHGav0b6OdQSnI5n/Vprpv
hwjpkBTpUHha05kWq/WfVelKnHFjQviO3EYbj82O0ERqHe0v4KKZKFctKaz0azkTf4EXKo3hTV/a
tUKd/ihm9h00LSY/Z14n0yfAuwhpUzIZ3anG9x1QSklKmK00UU+8mMv8rI2rrKH9FqgLhXa6TTUV
U1DuAV3w1gm1MCdz1RBh6bDoLbn/N1tkm4qpVNyDc2rRSGPcXQTIJmY2LN6ngG66KrHVCbsc+KJx
ohUAJhH1m+13Xv5OSnm4RuxwovenF7p7ZHbiFtNG65WAZ809iKxfKPQkKc42A7IQNfr+98P5/K84
eRg6qFSH7/myVwlaJno5TBgx5V4PCVd7uWetgSBDqZqvyfkKTqhPP1e0m1O+EG+l57k99vbqyNBy
yOunhhFFuB2NvM5F4UhZwdKfcEFS35OMRtohKtp8eJZOGn3vGjkVZVYiOOhXzFI8aX/qHbfMyIfU
iLfqHM4bmk6bG8stUCRjoLQ4Kmsq17AcLTvxBsA8FX6ei+bt1fyDJJCmzxtOoNeLDAJmLLm+GZht
0CzyPpyPvqfpK9ES2htAv/S2oJNE80vD4KX/attmjTzK2/qbxg1ampcaHIBK9YjXtLax5b223H5N
Ue7ccwmFbJjsWUmqEiB4LFXQddNW++lTUGoJIShENpOxQlN6SkrxQZEjKSh2mqVSnl/WZcf1EiB6
c431sDGgHM7jNk0UE56csKrexKEJDLwjyVokLJ6NabZKAfqdn/xbT6chvytrzCFUd68Fw/I29JaW
WGe288I5PXeLW2nUF4eboMqFTXmlVUr6cA609XFtiSElJzJ7rsQK+o6LYMP9Ou1Gub2Um0nyAOLc
TUC+UNK3MoGt2qo2r0T8fB0NJ4yCqCPLlmhFfTnELGKtpKUBbJ8+Sgr37QMsRf81MBifvYif3+s6
uC7WbUCnesickG1c4s5rvJ2gwahJnp/7RT+eEUGZApNF2Ujil/qkSGP9DcRj877pmU37mGwxAtc8
WBgulWP332E/U0a+tN2naJsAAMwHfF0kbw1vYTeWrHoHT8yaSdKpUlgPeApJthm0TTsCznA3Q19P
CKQXX4Om9nnLndFsUAcRNK6sXteuozQCHRtqCyfWQkSzDLuZ52oTPAwfsPtWsZjqC2z8kGJ0jqlB
/+ZJYDZVThHX+oRz8yHnXFVGDT4GBZBpe/2Q8C+wTx9RybsLERi0OTaelu2fphUaZ4CJENSsq29z
0zVPAN8rt7+/9sKwqBpWD0pT2JyKTQ+2m5gCTRUUcmRhsHSKvmvBnVCObqM3RWY2aCl8egDHmxiM
Q9deDmfjPgvrCiGfnIjMr/K+cBF8zv5sr0PiFSnw9L9SmfAZ1Sh92hSsW0mHmlRzyPPKHz4PTuCH
AXqEI0OxNh8ATHWnhPS7wyQyIFWW7SUM+5fisaXhZydjpBTnybA8uhhOtZjDUQsBpcX9oVWSRMkr
w9crVIrHEmmWBdCtD4xgTGnhCTtvWZRPSfkah41dZZmvQeS/NL+MyeBYXkUw4MPnTX8IOm0KajS2
nV97yLpevCWC8jxPx1moVK6YWCsuW3FA9Y/1qj4E3TLO4PzeqC4H/DryJgMMJCJ5zrrsBBL4sKOF
2D0vy4TG9VK+R2H6QBSz/QOEp5w0UD5C7cZ+ffq9CBR/D2DRWN9vxt6+qca/2KromAzcpkEFwdBl
sBqW3ht+C3sVnAW84dff9QSLgCFITdJni4nS3hccwyEsCYP9BOXxZQxc8Nc+FNpSh1faJAYR5VXh
Rq8OE54emt17Otsrt5swKjSrrbJTobjuq2fL4+14kHhdiqjQu21HzLsi8E/mbfFLI0lIkZwHpuJs
Kcp4oWGeY9Sl7akryznKKsZCXpLMHg5DtM3WShezxg3YE2mTWxDiXKbpyxrlabut66CDvUi4tvMP
X4fZSNa7HzueSUkUmsxoum6PwXwN+cmEcgTXKL3j0dJnlNYQ5PWmNU5XbJwBIJwTGsOfaKNMPpub
rnd1SC58sZ7rYbHtuH9sF97thRfjHWDptCN6cVVP8tM9bai399trdYKGQZVlJWTvqFYabfHGHSVZ
GS0Fjarc5QHsfWbEKy10tMx5AoWnneNfVv07aVuHr6jcqWpPwWyl4t8htw8L95aQqnY6WwWl45aI
Q4dGzgiXHMFEFSPe0Z4D0t7BVftQJ+Z6hyIl5mFlA4+g5A15Y7RM+f0FskTXVoh+nALDASJWmLYg
AdY9xzBcvXsZ88Gamw2PkNb48ymuD25n8JtzwDZFmiQ+rrXqu/+WZoswoxIizC/4h99HSMfnzyCw
DAJYBbrj/2HzGcTbdDnbZ4KwOzeaG9a8g4f0gDrv6m9/+Pfjq0OkbnBxTG4HF3NFsqpABiEus4iY
d9v1H/Wa2NP2fZRhAST+4Pf7S2Q+uHczuddE1inU47vsbqFbPytpw+npbnisJkbavHLGKzs99VSt
8otAnwtcWY/BJMKwjo8I5VRNBpfSbtToN5WewBeDKz8wRXHmfMVpJdSsFUd4eA3GSBUDcJ4mbAZU
4tj3jj7cdKw3e3cEBt2uV7bKEW3g8NzLCH1uOAe8NG6AT5DNrfuqIgdDEW5wStUy7O1fa0LceZjK
sOUgP+rZY02A9kWwSYAhkVvmNxxU1TagwCNVakyCUSSvN+NNRIveKOG+srLkjfQJkDH592SAs++8
HZjvJ4dsLiwAmXIym7ZqF+dI66c/ed1w2JdRcbnbqV/DOaSiBIJqBXf+YS+GOJKxSB1zmVVPGZY1
AEU9Qx9DkqWsw+kRiF1Sb5IROSPWg//wkzXqWuA1PPwWgj6Romfy31+amIDq7amvVRdkAl8gcMPS
hzADR8l1eNMJS4nlY/52GZkRiuxzp4a5Jug7xqUi51Vx9Tn9uxTiE9h9jUELCa/PyyMTfDmH9oLj
pJKeAYFK10ySpRkRoEsqqPSJJoxvBQQbIR+9QBRscGUUPlSIXTd+DfSnRfANu57WE+vCZYDQWQKC
vfQW09Ni2WsPa5D7/ZPhNfBmG3GfI5brApyXBg5GSpoSAydT2qMiMXXOyjos5tLKhRPJ3n4GrmFC
dVsZCHxCBOwnYMtM9bfr+AGAVMFtvLBMpq8tLSHVB5foQlhnsgAiYWto+vwf78OA5U8pz7bdZoil
elzGmsuWH5eFh6SpcPS7wf/+cw5Zh0xdkjW6Lof1LrorBsQPwkbGs7LpHBnH6/taqeKD2R1dwWn8
jao3wx+toL6wKTykQHS5iEjflNiZx5sWuZAprLjJ2MJL7Wq5i73hK48qUi1cjycLlst5NQYx7HlJ
D+XBrc3sse0avsBunSJ6czFkRSvBQ9/p/9sxdhucPXn74PPCNebEFmO4fRxY/Uh0KMaZIhm2aY9L
JhVddCKG5TNRl355RGEzRprJAe/FXo6UEXdq5mNUOAra/irZDpZKGAaeyXzxs2Hn1xk1rRFw6PBR
oxmeHLEatJFm3eLrKFHAWbcITt/L1qLR0x0wTqE0flecOT7uEh7rAfj/M8VVfXhrNkSYzF8qxAl7
Hh3ICsUcL/Wtt55qXACZVne/Aftdkzrgw/kZjJlGKpdvJvSvTvifwZw9LGYcYcx474oOueLWsCA2
77ePJWzAu8A/VpPVX2ZTaaFYTXve3VIQl5qe1E+2NOLwEcKwdUSi6eNAjj6HWErMHqMO1yk2PV6V
gw5ffoh53bpLbl4ed6hpEKm+amgvCo2HSzBBG5N73aDZahY0ZqLKc7VkaTJExSZDR2VfXjH0OuRW
BwR6P+1+Q7saAb5+74y0sJCX+rQ7kamwbYNSBLHd+P6mZoPYApOlcUoCvIAhrMXZXW3hwlwuVyxu
MYkhNWAgRA+cy2wX/sea6TcL2wCr6//zhRZwAMa0Ut9AgGyJfQ35OIorwdksFJVP3Iimj9BOXMLI
IDzNA4KvIUbiuLTsbSXVP+9jSLMFrR9Jc1FT5+qeC1LndKSnxSfsedZIpMtBWeljVApTkh+tic4u
ZE0guocnuGeRtOKpim/54DR++fKmEmjxCw6ROwBGbXN8fSbKKgwQriKA6AkZpizZYHLKNF5E02Cw
JzXBz4iknTun/tcZI/9zLk5kAjo6nqyk7rwgcnUgbKzaZb33T1Qlmardf625NChdOyCF0EecFlUQ
Mdad+8Y7imi10zsT2rCLnkRMbP4sIYF5eWkYpGn5mYK7V2Ff2/OJgzq7RWWB6GkASuT5JU16zc5X
ra2zmsWlGWEE7Rj2xoSPaF1OJP0WxTSkPXn2YvbihzIJdtmGl5QO483hYHT1VHSSfJ1CVQWlDxlm
Q1ZIbtoTnvhRg6ldMfxlDuF9qZx74Cab1ydYz2wdyBn+IlB2uU9VOvAv4F3UKX5Eh2q9jrbVgpHh
FA/+uCd7V6f01gda9Ojdcqg3sFz+B3xNPn30sf8X8kp6mR3/tJGXD7TTm2C0n60PMWQeVkc8iMZo
93IZRgnXVIN7Us/dJl1rURGJULS09/atah992N8F3qCWIbB9hWUhdJENeIayDqB2YmLUAdxg+tNG
K8xk9HkskPdEAgCLY8wZDn6x15YH5le4s6jgANmP4ajg9wq/5T05gbg13fbz2gmn8pluaJOv/xvt
8LG5OC7iqW+5i7HvGjla2ZADfMVpILVpRX5ALHh7xiKv7JMdfS/+8hREJAKUC3lyeRpEpGlkT8Jj
qC3aRYVA07de5HRJ+9ikuotMgUGvaoC4lhX0w9vIHL1J+UPcNe0oJqv5CW+ro6K12R6TUkb9CfXu
yupCjC5QuSCXVzNSITHkC0PilSClqb7DNWczhMB2tLMHd5GGG5OQ3Xosz+LWWSU3KlmV2sRoTM2i
2zK/5MGYEBdIvQ8AdW62O5JOz0iwHWksoaEZfaBO19OH1flpnI88YNy0wMvXW7x+BKsGk9Yc+b10
3ePtSd1+/0EHBpWxbWz9Q017mujzOf+JQKhyQhzipqEYO0si4IleBb4DnK9jJh0Pgjx8foxteLGr
SlZv06hET3iTzDiYcJ5e5koXI+6VAALl3SlTZZIdb8XPdhQNIcrG+nPrikqPZJVWUNtUNbuRfhd/
omRsQMgjicdRLGhltqrz4j55Cb6hplg4g3OktkDu/ZtllLwRfHo3ERTYo17k0TZUKVTitzc0D9//
/X6L3hIhIhIeXAe1XEYbIE+cUgnmM+LppupJ3Q/P0DENU5oo/CUbcg6OrRHFE69UCtS567p/1ChR
W7TOqFO4g45MTqp5T+7WxcwYz+rxUC/kobavKTlyD/VDhawWBG++245X1b/1gbicje7BlOEsTSf2
pu4biYE8wYENgLreV+v53iqrbUFzi3jXZ/yShugeqFSEeQZkUM65hwbGHK8rBs/MIbnw2Wt0ED3O
Hle8MAg+trrgBVSx72xgXuY8HS5Tz2c3bVp+3SCGY8VCMabtJL5VjvGnek7jnzVN1k89FdgL8grm
8On1oFvpCBEMjhPzsFNGwvktLoCdo/BlrDh4JLqo6/7GTjLkuHQi0kNuD1dHZW1v+MX1kZkYHVgN
T3woY6ToN8j010E6vmDSKYaC55uWznp0+5VDa36+xxOk9q8/e7cIB6vhAkHT3hMfHIIwK9DesX1y
6lXgRkvzRZ/nK5Zl83kvQMWOJsWDUQPTlmQZNRfa3+44Goie0PcZfkYQ23tplNWvDZJqacTTTFRf
kLXU1cHwD5bDpzPj2x0SEKEAS3FTKVrD1lZMSel8snBO07K6W9AFQI/aiFQpbyan2p6JEu3V7iu8
h6wrByJqQvgU7fmaT3RkdnxeKnm72US3R6+RPMtjqBs2v/SfNr+4k9tM7ylgxUt3hKB7AzP70sou
aw4uE1TG5Gy2rDfKkWzLV+j/CyA+dotq+JALISvkVHbudd/eSC0gZVd4HjWQUU38746UqvKRT9i/
Ydm9N9fneGU6kMg1DmeG6ifJ4Gol/forGyR4o2mQSs9W1QpKTtgPtFENE2J7wP+ztro54c/m2yaO
wQ8qkqN6l5ZY0ziUh2Xr3eLjt5UwVNtvxSk9m0Yc7uGQx09wRimKtoOjtD8oFU3nJlKYFUJE7Kti
tWNwtCn2Hmz9iTRgThrblANY4khlEjZDNVVftiWyYbj+UIoU3xyfFmF/k/+WjxFe/a61J5bSCzXB
tqfmwZ8WyQ3D/nwv6OGeiea2sD2pFvlt9/xfdDX421vUo0cCmHIaSufukQJHAXzR/hgT1jyI7sZi
RyNZ8NdUG95nKYeyP3NW5o2xe4EYd0IjaQD5qZqtgVbkvAilNtYVHtJqGiYgKqpIcnOXeNrIUQ8o
kRamPAiKewUV69cqJ4kWOB6bQacyJzQjf0N+UVJHfvUUjuKzzrtzG/VzJovphzdQ3G+dmlevRtDt
NHJHQ2AbiU7c41gZeehuOXfAB+QwCExoXuC+QZP2TFW8R5bvT78q6K4nzgtgKNdyxIz+42M4L2by
2LI80E3MJpBqdYMurobPSkUnRKFghK5LcpeTjBfF57UF4sIh9AzTK0Cxw0AgXETbHMZnNJRrtM98
bHLCRJMnjKdHroMsKbph/hWcaTts1YZC3ASjDXSCnMTNuTv3LBct3g1WUTP+PuKUa8F3qNIHjqXr
sJ5NtygQjz1ktMu68nPKw9WTJs5H7L5tJZmkqvnhBK+YN0r1S60GtGjn4VGi5cixYGuKpuAsXtri
YrMjGysPe5c6KywyUGfp7eVT+OzBZDH+Qh+gR/i6yPQBUFOvH0V6HpZSEgoEhRRyV/nwJYml50v4
ApZ6Evp9txkLoovQ54R4AKBRb8En3BzIW+U/6ejiijxcSHGyHHHSFS59nMhTVle17KKaU7tHAFHV
8sBCMS2VkYQSZ3Kzo0PosNdwEeciMBvQAE+YmpUXGEfLTK7RfrY7caSDbsP9KY1eHPaWiJ2QAweV
yugThtIJQV5/FPh+D35RRFg2HLXMSatUq+q8J2yWM7uUeTkIdfPrmkq9QyZsVT7pFJ22qxtYF32f
cYO2W+BgBJVjH/rqc0Fmxk0EzS5k7qEmV78aOa9xEAQaq1GyBf21KqjO/179pUKG0dvxR6w4Nh6m
LrMzGbVjaGjPEEi8uKxYe+gA4uXZGr9guVMvUlR3u3fPfGUP5oohfYnmTmf92ivCZSTQMassLAz2
8d74/KXdalN+pBNXi/W1+GbgMNTpte3uhgIEeF1bacycbFth3LomJaklzPToi5ThiWmHGAz26Ex8
LvmtEFc2AX3fCgOtWX+tDverl44ASFMfaqb57MSlSCstZe2IRK4HnSXY620A1scmW1fLQ7K3KGXn
+rW2U9aFLt05Ja2pV9rEZ2bxS7rcDHaSsyzfyi3/gqhSPW+4beSO5/tC3ErxT1qQ2Mh2tazKqhfB
kfS69URE8iKCvRrSGwAYjiiRgISCMl411vtcNZ/XDGdb34gCASCA7ffkPiBdtmWAEV9RQExXkq42
e3d/T363E0/7jKesanaocTXM/UaJxD5DaW34k47HMAMPZUhCr0yW6zXx6mN5Zg9jkN6kRyhGv92C
JVc0qR3pkQp2ZxV05gEknvhtXCV77OYEzdmBVIbpEfuHHG6aQ3fQNayRmVqKYn+SAtWHZdf53YCs
i65g8rF8juCYPCCpAwqsrxFihYcgPmm75eFRj4Cxv29rqPGomTWFllrAYEcsS8ycdypSaFOOGOkH
TOcogXWOJTGVXlRcR+W9ioZ3WKXSqkSaeDXoR+VM2yAWg4fiq7M45lAGby2F4gu2Zge9TEpUZtTf
X0ANCih3nFFQNer2kADVdI5aTCfzTGs3T91lM7PACnAf6fAFoNdhEhexjitP4R4URKd88YRO4IAP
Q7CJQ8SucN3Hql21Fl90FY9E9Gm7sx3BbkbQgS/QcZdFLu054Vd3Taft8Y0Y76hH7muI+JEQtXqE
JJH0j4cnO09iDInrbCQT11jffBxV/W5h/yt5NsZlyz/OvtMufyylxnXqkiy/iWYtjRQn07eBqALI
UiztRgf02pLq+Z8O+cz3v82EQQvXD0cgIHuyYcie+6+Y4st8eEC/D3Y5V89hN5SLkyrUmJZ4boYy
LpFqfUjHUuFq2NK7+jr0D4swWqbGWFO5MypDxAnm69/2tML/HkDIzJ6INjrY2CHDH45l4AGm6of2
eTrZdUptRMhXsC8Jqo8LTD5xcBRGAkongqEvLbsiHjfbrtHPQATnBph3TjPhhky53G8NZVUdqGfG
mcFoFRASLfVBr5AX6a+xYD588dOGz/kGG5ngceJhmKdk6gBbHEG/SFfFinxMG6SMUB3MLoi8yU0t
W8zfpYfbVYi3vVXlbHR9hzZU3htrYb3InVE/7mWrOcGX5s10UzVntHsNzD2XllxgP+UMcEb7vbCP
vztmC/o8/n+xDRIRMXw3CBW4kLDIXcKdDxcscBW5oJUQtpyGSTzF6ma5Su2LENSj/gaqotv9QlfL
BlM4EAl7d1UKnluPkjY0EDe3xjc3e/HZBoEH0fBWG5LX1mBPzJlLMCXAsLo/kHP+yfiEfCPnA5IM
qyWhFzhHDck5YR9P/7cYYjkSaLIJmOAX0pXu7uhus3L+mN2r9o9ZsLg55COKiOg8qhqNTMK3cUC2
BTD7XxiEz4hY0ZCwN1jaCXghGqSX5MWVIpYN/cA2e33ifIOUFQoBrJKgJSqyh9RFv0HILojtBu99
D3v+13rBfMgjxptLxrQp1NHRhCohqtrvasziXR+YuU3LkU3FlpDOhHcq8zUZmaZdxsieROHgLYR1
WmjZLjXVDHpWxFb+fOJA7iVc4bcx1SkYibl2H5OGKRTnvXpE341yXw5rwbd05/3SGD8zXGcgviVs
62L2cESch8nENB0ihOE9LAVHCRhX5tdj6bj/0kUe3GBCWpRHI/PjYtrGPeB86a2K6CFkV9V8jq96
PUuJTkeZJ44SfyCMYxY4eM7lJe/7+cxPEUU5T5gMDbDP/qE+xhPeuuWkPezMJ1AIu2NtlUCGovKc
zL7ozoUjT6I5QViARJxUr8GEf5e2cnAyxvxrXYg3ZTO5KpMhmAHV/X+H82vDwoISHBBjpDeyt7+B
f8dV1AQ9xiM+UbzZCB1z1DzK71LFkbeViNd9uN1AkOnvSKvpZBt597uW1mLQeOsCmz14xv+AQvZJ
Xh0qFKyigBLcjeMKPvR2uhvu8gjpyYgqnP9iOzoSLxD8zHqs3YP7k6ulIhM5TCIlVIDtG2GKNzE1
Lrnc5SyibqF5y+KOiP0H45/Vp0f268EODubjWj7OoV1S6YV5aa8aBwcXi61k9HQ4G6RFVHOd5WrX
EMFy/vfMqDNFMHwRgf18LE/lxKYCCyMofEiLHgOMhxeKI4aLgJYTb9YJ1SfgjNi0aBZfEHNiEYM5
p+8V7KtPffmNxGxa8R7CK3T2kxrrCzA3AH9ZD/XjoYSvjvZRJPmh+ucqTkEFA8weUKnHiOCvyOq0
w2YHhr3ixM1IE1XKojbLzSZEIdv+hDlVgC5L26kz7r640U4xHHO4Bz9Nu/8yGF7ltrYXMqF0gYEx
MBLUKTw2jbannxI5TZsc5JTBxDSAbjpLv4QkiRCgt/lx6yqCFe0SA9opO6AuOGTe6jtY0HdVoop5
mpwQCpBwC81TvendO8cgyZwtg635iCczeTuhMmOcUU2U4T0O9DKO+yTHyhDdG6ZUze1ks9a3j2yl
FQbOWDhKJJ8Amf2t7FwGfKPeyPJ/b0NKgD9XxbhZeoR4i5zw+VJ0tU08sQSanDvHT2qK04oRzJs6
ctlRxCopLF6h9v56EJoBboSVToANNg+/elRA7LviAADpACfjIeneHDH11m7xj7uo2l5rrAENtga9
WssOnkW4uIPZeHExJ6KotYuIBr6oX6JQT2TFyfgAQPqtsNAfKXO4qaBQT4fIrCkyLsl9QoP487Zb
ijHkJks3A1QKDZobViFinAyyyEoVzRpSPI7pWlX3A0UlZfVoHsrS67jmCckhN0Cp/KIyacAdO30v
Vsfu1D5TsaAeIAfgha69UqRfNrETEvqp4pTVy0xWmG6aNtGbtdYZEDSJAZxaZ4vkMUzuIk0TARM5
0W/AM4K3EpG8KxuUuwjwRci62J7X6D9sGMtR5IbB9VsH09S3GRtP01RNoenaQFDw8nmTJzqz3/JN
ONongieWB6FekyIR08SQmacPQr7vc/boDUQYUUyROorSyARVag09wLHn8INXOiUTw5vs/w8wH6YV
frJHPl1gFW/BxLHJ79ONjJpZYb70SjjbKEvtcrxmdyjgmX7lvGr67Tj+ETJ34IvntB1RMPCm99KB
4f/GZO1/mqpb1QT9hEpa2wiC8rxiJLrxK0fE1InQZGjkSShKxDB3EN7DKCIDYR74bc4pKM1Nro5Z
fr74wb2PVlSsEwAHz3VnMYDbrVNQX2JaB4BB9ax5dR1hzwbM3xiGnuNBLFlJiXhYpMRB8PxBHTqe
1/8Gi+azy00U6iu2JVelq3g2HxqnuhuJkF/8eqJeJ1qUOaCetjiAPxCtbYKISDRf2ZeoMJj2wZWf
dydRMHBh5t+jcLq5eqUtf75l3lx8Y+8fE74K6b1VffLT/rrrxXRpipaIptSCRkLYpeeJ9M77qPF7
C9mJ33Ro0H15q3mB+ZqWtdWC/sEEfG5OTmu53VA7EmEDm4aXf+tqCC1NIbex3sc5gbE05c7gBzGU
noZbsIWdmuIkh3j476v5spvOHv0YrMV1SP7EKcv/lriFYRGCj67E4lSe0uwyx7hvWA6XtfYFX7aw
Hxk/oCOXMd3UPOiZjzrEu7+qS19Karq7bR/f9TxwaCLun0bQ3tauaFslTJQJ7GjXOKQDm0TAvUAm
Vih9HW29Ffb7otu3XA+Zb4wbzu8wwJX1agBsXMq1Feadz02m87un+qu4+KgrHSFkR08o/Wa6cT7E
WcnGUiwr3BMlJmv9kWpmc5uQXIvQhSheKktuSHPkzabfe/zFppCw7eSKqQ08FG7RmyqYRmlUqowC
+I2O+wnTj/fRAvM5K34I4Huoslh188kGfEjW8Ef8snEQVwhDnVY4b0mnqQeFgT1XYpK6ErCPnAv1
Ft7nU9+gGXNbYspbzjGi6Bp/2E8vExkFv6f4EXuIBQ9fo5Kf3Zi8uKhM+RI0lBd6IAlLK9CfkTtx
lrkJkZL8YUSHOzSj0pCyo1xhzeqjnsm/pEHP/6hs/nwg9UeThVcN2kGGWxn/ltoGsuciyx7LsJy2
21EaiugrTAHyic0cI6fa2VXAn0J9OrkYCBLvfZ45mtVzzlqL+Qj0Kbzg8g0PIefg0CERQ+seAwJ8
GIVp987CmOKjfcELBO8lUnke7e5RKH1Sfk67UILNHjHRDicNn/tWIctYhUBWc0DO2+o3ryio88m5
gEIJG65AgAFPyugKtiKj7xJS2doBWdCAoHwmpc3sjXHrzKBpbbEVjHyhvVVwPEZQCUAR/8qBQNjO
Xv39p2KWHYRnllaXJ924JjQ217APRn5W/BuEPrHQlOElwfEcRddXw0wz2LtNjGG6eVckCPTz1sgg
Myy0MFQhYLdXkoliAGKBBW+7Krb6jn1d1iiOE2KeBFzoFoPNGbZv2ADzJqR2mBfWvSErnBHJzY+3
qiMgiEzu/7VQO09cvIxZf/B3q1qVSoEvlLf4XTEeSEFYtkALbS9cazJcjyp1JpEeWHqr/y7ckJ2e
CCZK8NC78nWmcXI/5lw8nvjSmsz0QQMQ4cqmFoIOzl55CXX9giymcI5Qayg6631St8bBE3uSqycp
AVSHtgexP9bEmeaa3Gijfl5FHw95r/Y3N6A5mZ/D2/fP8uv2Gyd1KdXSp2OGLjC675ZSuGv2cQ0V
PYGOuownm2x9vAisu6oeyd1Ic/zjXZFn7SAu0CmMyc8BSALoahveW8xEgwN7n3qUK4pxdsaBwkuI
c9bVC5vbDN/dQuluuKWlOy+N8joAhQbSalQjIelrI19OJsNnMYndBhAO+4DWFruoP8YZn4sxMz2C
Dir2V7nujxA7kpB/uKZ8pURj302HM3Eh5qz5y+5vhqQ5IaqykgCLI8EiUlFU0qrsVs/uOfM3ribK
KlX/fMFI29yY4GEawLoYrI/cef8Jkxj8gFVECVnbP/0hTv+NVw+OL3rgAB4YNO1aI0bcLPuibikr
a9GPI3ndrl4RzBZDGouyodVfhAAToIxVjCz3RabpCkvbCCUj04aPuj73fwLEq1ffDOSLtg2/hg5u
smQ6Kuty0P1l+IVYe/zMDoc4/NfpoErLj9cNEV/oo7uW+AORuVPe+vw3LwC5OJMRM+/uhFvAbEYK
4MDZJy0OOV9gSCwYqZvT+IfJ8jswSrQn/3zzqt1YXgBF820AgAE5YmfPEsjJdk9UNtnN1XBcfkTz
saoGXPM8B7m4/ROHAGNCQXjp+rjChSIRlTApOt9uAi2509JKmfu+1/sM/M3pOuO1VnejPow1xRO3
WRcMU124Q0MqGVu1h3AkL3mZ8VRV6xIVspKlyCxhwdnnwOLxG9tF+kUrynGFXo1UeEej6o2I/c8N
nB7Wf0a0qhiFaKaOoWeXaDg2oKYmKT3N5a6wxSHzTGrVcPiNWRhiHl+4RcFeG4z31WiS0PVwIFxH
9ahe+OYWgxCGn0hP7ad+z+JqbG6R0ApRlSspjhHOdqdke6zI1uO4XWabLzjD5zIp6vRw6zUU/fRQ
gjnbl9Bl/+HQr6apCU5XiZBGIkORsVk2GWDteAbhBxo7anLUWxV5KsRA5CVHtotIzvjYKHehdUkQ
Ksv99IO76QD+MvzC7CJBYsa05WbaII4zSsC3HkPuhyVjMfE2iEVOsZaY1ZhAQbS/RgZgB55zAON1
CmXUxbI14e2o7qUxVk2ieTofIsQR+qqoo6Mz3TqIv84/HwkJfN7z88mwrZNagxiiSWi8JE7viYMh
u7kJZQnM5JOl7+mp+3CE7dB8rQJgL+/SVXxnreT2Pk2od3FmG5egYIAyMDrba2NL5qjkCYfNVKwC
VTxGIGw4JNkQGXx/Y0sJhAluAMN/HcGffpjsz/shMPD84TcgWfdmq5GO0PRw/uy8mUfc+VjuEjxX
GbXwNRTUUtvzHQ4uD+TjMmoJcXOh1kvho7Ps/Lw6f9QYhvbGtRXUud4/FhozzKmNo0RC4/Nqg8V5
v1ZQ3fUqUjNBh/U240vy2AmPc8xmxA/hA5invpPigQof329Cucuo1E8Oj8wV4nRyhWQQhWRni9dr
7z0hguEgetFLSDtl0Eaq8aqI+ivTNDx0CrW3IQ2Vw9iyIQQ3f2aNMX3UcGwuLbEUeGTsGYT1ZCOf
Qk/566MDuLkEytVCWSYZDoC7OuUwTvGI9tndzjkCqBzfjZsqQo1PywYQhmX/cYQ+fkLqaexdqF4B
iywk0f+GV/nQzwPGQHhC5xAQqzFhMs2VBFOSvB/j8VkffZ9ZOaGk0Ip0BFgIOLZ2JcTynQk5TzZJ
LWeBAaEHFKuIqATb4zuzpGwfeKjvbGQpoJqpn4hQabbGY5D0WxUk6xXw++bkO9Q2ebnCAAVdIBiX
nsRjMikb3+X3Ojl3LFgSMFf2jQqwNFDpIt/DotYDNO7QQoC1oG51wItrcrqh+VBANAqxJj15+IGe
Ovb0iSZ3AIXlKj3bytTU64Emf/5LzYO/RhNAr7o62gl7QHH5EyWia0yZ7nejF2AbkN5Rn2KCUsLC
aSXb4MvfWzxOOEldhjJQNgrT34V/JT1/1XPVMKT9Q94w143fZOzHDuSd2RBSBHnH4bKUhRswI0EQ
/V+EoXjzGzEZEs8I0juTZcmo+2u/bH88GLS0uWiXCu8TJBc8RCdmso8ubS2035jrKcrkTflGaV++
BzjAiapqKpKjRCIBuzFfdlFcUU13bOQ39WHGzKpz+5Jqxgks7/b44y06fHLn7fdATDLBq3gX5ORT
dbvGxFzFGMYam09wLOxbzM/ykWV7XWen+fdQxlyC/+jzRc2Ywk0hleKDqjYUjgt62wWsscvOHBEx
8XZ7ywph6rGaNR+QOiY/KictRlbfpMIZ8/G5PKge2oLAi2Nd5trSRcgyU1QgAal6fR2LgSj7Lh1p
LmWlAHwYLMHRWxjP0OlGcSwOs/nDGuv6SD7zF62QbPWP3yH+SObRJpgfh+aQhRI4cvCqxUVKiPYi
KhBYGtBKXo6Zmwhyyspe3zikzXxn10LJOC/8xbGA8jTfl8YXamSeoenCZqn6YVZnuqWHP7c9FRye
/iwjSK+IAGobsYXBrUJQRiPG/m3wukAETBRfpiHexHxU6fk8XxcUBq/5XgdxVnOgWOtt/VioWYIo
Vdbe9jutQ+/2p9P9gWSOJee+oqOGqG4J94kg+vFGGQch5r/A9lMm/dEwuCtO4ayoGGhoHjVRZUhh
TGK0dJ/ETcQtSiGVy/dzgHsUnYCIlj26kE1FD5TwvgUsbpZEAlX+cml17Fmzdye5LDcJJWtS5net
09VQ+Jg4viyBeMEOMkXIVsMyRqF1/azv1Q1es1RRbJvvlcYP9ln8TVmKJ/f0Guj/1s/0WcVqjOtU
ASOTdCvd3h+XYKbAac6nWyljf/V+yV/+IlZuZph9zgtKHX7zXzTejG5kBolRh0nljI/NPt3ykvgn
yh+NWk4apFbC2IIJoW+HSC2S0HqLMWwbo4XKE98dVhyD9YEsXXkZf6xBzazfgF7LWDtAl4TIZcVz
l0zT7xJVPrPqS18ClkrVoT+8b6in+IevDklzi8+F3aZ55ggNH2vvbDp2bnsRGmtS0s3Oq2wvIaPI
a3zIgty60LIgaW41fq1loxMbdJvUvfyeICKaWgGyvhnHN8EEuyr3aVD0jXHrWG6k3QZOwiSkVx0x
NK6lw2mzYygfzCpyw8z1S43nMw+ELcs2Zv9WPLJ4uOu7Eu0udsmv8yjYNfWhySqGtszW7Uc2OQ/R
r0A56ZSeajfU6mRbmdkajcZLYHgwSOrxvbc/9GUhl7TU1pSt9f1IKbNUgVXcI4f6Q0fKINeJiihq
zCF+WMoDCIueuekHsuojPwfOXTWIC1a2ry7vlTEYwcMhssEZ6t52E08vYFywNFp9gyv6x1zyQ99u
vjsCoO5QnNI/vy74Uyz9Kddei8IReBhLriHRwAeJ+pSA71AVpc7ygKIjcoVcbegFXFi9uwj9c8jL
srhJEW/x5LmIARm3pvK0EJ9CVZt2qVyJ317RzXbnnWqzqFgck6r3RrE+5hRF7GGmGUcUpv+l6AHV
L/TVGbKE3mWQwAP+98lOSeukt1xR60/vHoHl6GYqtSiGqsOGaJyWWIAfiUWrD7XqhsO3WkOtsQXZ
zBN4rsnnKMY5mS2nO9wx7JjChGVP6ofVbSkgILjN461jIsSzSmyCxQ1hWt5KiFPVBo56Mu3TKL8L
Wi9mcuxddQVmc2LNbNFsB87cDVrH5PdEMlrAxFGfHhaxMdpBVzan4xjNN7fOeMrsQgEaIASLFAmq
RHYJkGgWKNJWan6rz9pwBAfpbtXeTHdZHZ26RkjPSRijpP6+McTF50OXspgfBR5PNiXlqp1Jody/
zgxud4PcIB042Ktx97HsD9P5/bw8oF/fRcZVHh2nIMbEhv/0bCt1RSv6BNl6XOl3gXbQJOkUYLrc
/sMcm3c6uMncUqjLW8speSsMStPj8sDyDn+wB2fKnx5E5rNQZDeVknsMjzd2imyfkPsbUFWjxc4I
dbB1yabIaGNwNfSrfCtgtfb6tbv9IgfJp+aO7SeKD/0sDl3pYWlnQgLx6HFl7S8X1e89HxIXSbfC
BjHy723GYIBBRwlz+FRFLowYjX3FkRsMTJnHufKEcLsnAqQZ+ZcSNYxhWIYEYw+0+2yD8s1lXMr7
fdETN7YjkhesUlqW1B1zT1vvQypl/UUp2mi2ZmEe2thRVJxLY561lH1DArl2EncvAtwNzR0iJKAT
Pm6mCzpNs568X28QpQi5/wy14+AeZN8pOe8CxKMnGDGVUZwlhurGKjB02S4TLLbaDUUJsKmJjxeh
A0iTprvmwiveCJJkoOMrvKN9Od778MfZU2ROFokVgtkcQvIVuJdnWyU/CI831dwgqusomVJEiQNl
bchXC5AsYADphdufPFzE/8jRBY4FLIVYvUzW+ZI0t/gv5wMOLqcBKO1jX5omwKa1Fj21fLnnGYfW
Kb0aMmENwxj37K/MXWCY20bRND5taZ1uVoB6z4tiWRcWmyVAgN4/4si0bEaebUvx3TE5xZlz1PHY
AHsy4gZxTTUL/gagid2Cp8mN1mDGeCmDQyxaq5b+fSQaNcMJw9wySJ6maCDlDbDJf07TuMIK2cPY
ehIt+FweLj+HdJNRNoT+sPeehQeMmqi3/Zuoja01T/B0hOGoo+378Pk0YwrikLeUiHVyNb00N1kd
wloQsCv1Tw31sSS/1mjfmHe851v3UpeFGnfMqdISN4Uxjq/dtOwZeAQY4F77RsW8R5DOoDfMpCCE
9T0/DRYgNOP9fG2+RFUHz2VivDqa8z4ygOQkSwJiRQ/2TsFyZErnCUFW0XmrFvBJSxKSvryCUXA9
vcOBIvVOgrr5RyUUoQ3IKYZLrrMpB/KIdrBVDTbxakKb5SgWCSrdEWbdyZY0mMqgMg3ro0RvkdGt
gpI2J010cfUBC5p/pmD1AePkOEG4OM84NUSPbKXZMong8V/XW4ppSsqrTp8m3/hAenU1/j7Mz4rm
LJfixU//eZqyRzGuHCIEiveiRK51eFIe1SIZrZI6YY5rqbhm4QkwZQCfdE6e/bUR/w61r6NufVQ2
cd3iSvvWKXodCSOTcxayZcjx7uTlSLDEQvYp4kBFEIzRmscKUhsll2iRv581ZZe610uXxShnfui6
dChak4mGbOchcRBCQ91QZRwWb8YfOWrby9E0xak/va3kXfrC6oeYAZqPTh8lNOsiHsYzCrC6UT0t
7NwDrQ9hePJj6i7g42zw7kiCfxdeoOcsolMJh4dMW5K1ydIjMp05mFow94axbdylV+76Z/d9kvHy
8BLVOOcG/0+Dz9J1cOUVeBKfDCTpyjHTU5Q48loRn8KNkwawINV1pujEy4qZgH/Tx0+p0/HpDQiY
ev0lQwlNCi1xqD4spMMimLzOXvy1BsYsRFlSk9x/JJHnLW6bcv0g9XtrCe0yw2LZc+zrjdVt/CMj
ji2RvHjxeGkh0cL3AmBn/w2vAt2lFUqlEqaw+CuPa/wUtQCjWonpbDvt0zF3/Bd7JE5eZnryr1rU
jDfVXAYIRA8fw8zmfxAbTwn2P3y2HLfhASrxfWVGqC2etBmxussQf3yqJ9blw/M8NKT3jVNZQpPW
3521i5wobKCOohZ1oX+kqLvTXhdsglM03iHOZRNFdIRAgCW3dox731VivfgLTfO5IJKrjX+PRiUR
e4pniLjzGHg2u/MaAg7GkPBHb58iDU5PtMjDrc5yfhTYv18q5T6vjjwAV9glVIRdtesfYyJKneK8
lczl9jYMiM7/ardlt/2bxaao8mD3AzFfhn9BBGen+n4bZaxUCLIXGqCIPtK6R87g3bJZwNaF3rY5
gSlg7uTujQ++6oFBMoL9iLqQQMfeJiQD/GuFMAzbk5bxDW0q5Mjo5HaLagVD7lplJuVnrwRU1Ikx
DMOmu14cW617StMuelbuuiL+WK933Tt9Na40GDIYWplpYefSGV+APMN6hcgmOip/FQBTwL6ChCKf
09WSGVicLokM75r4So+w0mpnbaAEps27xCU2O405GIxtAZlY1VyT2+goOQCr3qAI5hQ3rfPnQ9Hb
PPh4WgZsMwsD3ErdohRhXKU2CGWEDpQPaCofOHRWNEMRu2WhthHii/CUb4wXyqy0RKCyCXrRFcuG
cksIiQdJcIynIrPUqyQe72op3AmM4arR+mlq9uPA1GT88VUgYy3Q18scUG2+75/qoXy2/gSf9y6S
XYoMiDHIqVKaqBOMU6rmPVt5/js+sDUVmo+v0Svf850zphPD77gTICOufLTNPUstAGrV+Zp8S2RL
3ByvOa7lXywHyf2L10Binufy638c+hw1Gh+rf9QVFWkQ7jMt933AlLclZ2o5j/F2bZkboZgxpe1l
pkQRTDHVGwcJ70QGn7YaKuRqhO94zSl6fVHfasSGmkJH0rhhOJ5tmaabj2nB74Pvk3FU6h5LFTwH
Hy5IOk7/qJormwFyHZ1Rs+uOU3S2nlcDj3Wk5Ny7aWlqdDTaDqDP4SQdU0lWtGyV+iJhrj9UtGRr
Vm1XhdV+d2385ES9V6c1QoaZ38X0mvKkOPodg/RWY8dPOy9QYqjTDaYQG1pQj5A6A8VTvrt710W8
fapVrFczpoGuJNq7ByumZjSSDL5K/kVD668Ig1RSzFzSfLfT1xzkw92O/Eg1hcO/VyKV8CKZxpJm
zVeDMUDkuSFs7DT0EQVIlnLHYV7KDA8E6hToPJ6zQGVeUSr2p3kNZAW7KjY1d4wtuxfrLWSjYMUU
9qPfKSFfZgx0XkOKsnDl9NZs/009mLiVwdCC5XSYB4/12cKkB7TICo7Rmqvx3ZvB80BNrL8PRfgH
zE11VbzLR41B1OVyP6JP9fvGaxxK7FAFXNFlDbAOa5VwQLa644s9Ctpts1XudXQCzU5/BJjSaqyN
L9C6tTe8RajXPEXCcwa7bxI6RwkkkYwrUjZbL9nTKKLtzf67ZCUZ4ItdUgLyFuQMI9zYdWkCb6WY
UM53SJwdOBKNoosh7XkePnoAR38sbrbNJrjyIaQglyJjFmS+xyaqzCZj0PCvWkYxwxm36dzIWbp/
o8NCJexi6ZR7NNSKuHnUgRjXekpivGuHLoOSzdshCKeUry0HjyItu2RnP7vP7i1Fp55b1HLY2d4z
pak2mcw3fnHJq/LwU/QDJTT8l2G1ZqkOaAIjB+2jaZYjak+wqGhOhqiB5s6o79c7F32+NVy6Ze+m
uM4zUP2/TjYv38a+i02tUMBzt/QMjsqH+aHYmoPYZvBcB+ekH1lxEj5uKlV/bbueWsKdjc5PCRL+
er5gmb+H6PJY+8kfywkbJBWRfedARgq7qhiYcUorNHZiXgrl50k1Uq5gzsXP7o9tuPsKyKb1LRzA
e6lWSYVVo8eFv2E4rb1Hz68H0DACTSWFnUOF1hQQ0hRgJWROd5GR5wcd0G6DhIplN7Pi+gvcPZYq
lkweZBLTkv6hSNHREBcxjvwa7yaHbzmoa5kJopHHYqRWtaJ3vzryJvkhGSjk1FqBdDi1zCcOECf/
Vf7SeimbS53yuCZxhXsFAELCqxaJefbEDpaApSOEMzvcctN48qxY8c691GMZZ5QWT2Zodr55+XRd
JLqrA4jBuRENJBMaEduiarRqEbRlGt/G3xj7kxcbd7UJk/73d2BiRf+c7CqFuFqwkCoQaOBg9apo
OgMikV5D9SowvsxjuzNYiWhtQxVcOh+Ds9rTVbhdvhYPolC/jIoDXHxbqHRfMykuLm3pgoyV9qAW
z+L6aApGS1phnPnqd/jiijfkPHoRd8k+dGWtJhaDJPm3j3mEvY16kNDUBJZ09cPkaFWyYh12gVSQ
y8FgGVusA49oczJvFz2q4C4cKZUCpr2n3T1L5bbilJ2d6Ai/zQMfp4orTHScyAb/ASzdR3B/dWQM
D4GgGWtT6GlXKvUCAVB9+UNR9lgVG/WrtdyEEGeuUwpmCpFx4Bu79/zCHtjmq8RrHkoYamC/Io4m
Gi+I74nB1gBipWvwx2jDTdUaPkyKWhFNDugapFATYaC/7RcSmPTXs4iMoXM7JxSomqv0pJYYDD94
+qZVwgfZJi2/y16JYibcjm+3ZTM/mJqQ5DAUjGa02koVPPKIrulgp5QwYy9mnEnctkSouqO/dOU/
Rxvqe+ix2wWItdAQpa50sqCD8V0Uar6u31+NpXAOXjrB+L7+oi2bgi3V50AxarXbC9MkavziYzXD
xIOOZ8n7nvLyRyfs9ZZtR7Lxq9B7e2sjT+2q/ks5UEeNoBrVx7wFuBTJMVy5h+utSq3JMFzzm1wl
jMseYLDkSAWWo4xTpX+tgX0lcjVgVlcUTXZFOiQM4HECATeLLHRobSWUq2pOJDklGqLQUoh5dcHX
9fR0Y9MLKb53CNZ3JDOBbVj1NBkHTpwQLtjirHvNfai42aQVo+gcxBZL/Xw9RHxm0hxNf3B3CvvK
rlWx+GHI0jV8GwqDRFdL/zJ4/NC5Hixp/lJ/P4FNYglahWkYtNZrZGDbsx8hINquQJrzqW9IWKCf
h8+wzaBLLd9bCgOf1wddyXo5snk+3DFNekp+3jOYilgh0YpGxzBD0kn/hCihRky1CIfvyILe2dzw
rvJ38wAB+hTdbtoqN0oAya0ucsbOofEu9DgNBZtA6gM9G9vgXhdU6T+rZialIdwmAwgooaltbNWO
HUWaP8gJE7faue5qkvU3nqlzegpZmKvFVi77kvxIXg7bgCqm8X4vXjlz5C4FeB2Ema8yaD2uGYFG
1hcDv9cC6yyOFjtm2yGZH5KT4LUX0iB1ukyvzFhPK2SoVwSoQOa7m/36XlMiAWlrCtYzdwpc1dk2
L2O3KSSyO5LMyN0SPAxMGIUcXd58BepOL4kYgf+cYcFolyuAHWjPslcoUxB1fCDJIRbezHyVxV0E
wjW2I/64Yr5xvnLaXuVIZCW15uwzXpdfV8WWG64uv5pjNdcl+FjNdsSc6rqsNkLJhmqFnB8GfVhw
bBhtIC163T85z1HDyWKTBW6IJRuPGTc6Jv10w8rs/Gxqxfpk7m+chC8IJRGArIVUTax3CDZQy+CY
kxT5EaZ95BHKFD1X99XWM1D2i1jNhbF/iISKKmmlUJkqZXHddsv2hnMNv7sxWPcrXGzUYhYJiSJT
gxKGtRNiHygdV9nSMRIDO6nEWMnjBeUa4juJFj3lKkxJ5KwwJuKWD4JvF/MlfoooBC3djA5ANzBf
YWcNfBXVK+hgbAz2Jxe8kOIcI9GwzlDffjbDUvWFnp2q7ljc99bTsebQqsvHt41AuHVSsPKWz7tI
48Hih9UDjRhuAmSI9xzWuNSJ0oIuz4ZFfstFoYUTQ8eNDqmRftj6DnCN1qUq3DoxIDAFR4qTYMFe
UhZY3wnXBu8MrS71ODRlNoeH4ri/ek4IN2Lmxmeyjl0IkazAd+dpqj01XA2s9VIUY+Vj+XeHe2ib
DusyLNAC3cHtp+PWj0u+zS7Xe8I1depPKZCCXnPjM5ID+JMA0CWMeQ5+zx5dXHIY/r45NXQRBfSm
xImXGf1JPFpynxfNCudJj0CFCco1HW8GpZWhgfKDsYrAjdHvxM9JX06qF/1gJPGNnhF8jg71Gv3d
yY4P7copAvkvCsG0uCWJ5M1ve7GuSPDlVRFmdeGCnRO5Vk4z1UKhl/9lAD+vuvN8OZKw7qWCnuua
yRk8xa7bVFb2y64KDtW+zZJq/Z44H1+Aca2O+c6aa6fS14jLhr4j18TKlLalPB7QG6NpNhut6EE3
rSYbMS73BS+PZYiicPMEU6NcH3RHi2RFqRdP3IUFotysw5RtktJrHaCQqyZ8YRLIyPAq2cqFgDAe
ii2nqgGCLbNCbm6N9qc88WZp24Sdv4UwbEKL67ZCQhEg4W2f/OAk26FqJv/GIu7TSCpI/e6N0dgO
Z+4X+LaS8NunaCCnvyvJDtf2rmZpN05eQmPFVmhhacItN4e7ljhPh8oC/SCfh8JMGkGJCeWng34W
AAJ9VrcyWm0WUrdHyuanoc5grnR5INdUI21w8UlIGiro4bXORYqL7ZZqOmgeSfEEg7224o4SQtnB
SYUXmaP74KUEK1WtslojPCWvqpDn72RePwS8SiWplmzd3Wk5YfISZCBsrAwYCDH9dC+UoRcL1mEB
JbgQCBQudN1bEiRcrWukaGmy84pf34kQXMTc65zxJvY0wCRlSRdlcFSU38B5i0fUZ14OWDsh1X9M
Y3HwbiHsLuHdxDqZ3Y+88NXoNi9VzfeDQN2NA1cYo9nFw5zn0dg8jFW+TVZyIiD5wx6toKLs4RVp
a93LT5rgsvJLJauxmyPqxxOPBZMa57980SJonu28VpNs0T8B50cJPyY0qN2ix942U7FJAZjTRP21
6vyBt6lfzWMXUEN+wjiSyRBrEs5kBLw44zKovhiq4hhvfGQnWDwIqwbJ8cHP8FAs08Bn7FIX+Vrm
cVZJz54+qHn15PgFFbMBnLxu3kYLxxCu9I5wXf7g4yl5FoHa6VkfBi45JKbxrSt5Vlv1D+bChyPy
DM9rSB97C2Z50kP3kmt+nfFI8Kckxdy++y2TkrmWcby/u98WwV9e9fPY4Uz4zq0e6nos56CUMX5L
vm1YwCBJL6/tlAmoSp+IjLv9rgQ1k25sn/Z5WIJba5lKBNzvs7jegvB+afXi2gPSxgVBrgmwfQc/
eDGytcGIyH2tSaxZZH+ju0CVnyUKx+M9PxTWNBIsPi37SYUYdK3HLBNilz1yRIOK8X7i54duE3Be
Crz2vyc+26m2zx7/4sLv7cpPs0lQ4mQt8wFbyuyV8SUbm0FsreEwSTocZ2Ys43ktMmfiOsSe3M9m
JTzFUSbymTFP1vz6fPktUQ4oplFDGJ0ntRWuUgQM6rzg2E46xJ+F+rQP3oEuoWCY/FtgELwIeLiC
fz2cSUq+B77zRMRE+50kXDA4M6XnIBy1p9Vydo4iLzUSHnQEwgDsbs7FlkBPoPBJat5yiU1KInII
n4PIVPnMXaSBvf3u94xfz4M/S8iIoLu9pOl7tt1bX0TmOq13Nl7UY1I45aKxWIYFvhsB4QwKqNyS
aGFOYIE8cIOzERAjFup3FzzMZBYgm8zo607dt6de5Aw9sYYpAwn+HPBqtPF4q/nrExptTEAwmee6
fN4AlKIHbg08z6DIDeh/j2dfwmyCColgNjiZoVUzPZ8W0o0O6K9Zxyj9xbfsuKn91FQFxiwlaDlM
A9VvWjMUla+CB+KB8KxcMkRerih0ogQde2iIce5UaJBE4OhQMOngVQRXhdrqg1KyAMed6YDbcEaB
dtDlFTldsILtXir9I+1thkUFtIFpJwJUnN1zpPTUQFcOx8R323Rb69u0eVpxO+PGSBzVX5FStnqM
jv285dUqpdKW7jsr58Fot/1jLhJAu5Jt0TXOFrSyhxPfRCuKrr32YWjPr5OiXU+Kohd/PsdAPSkz
r/yraO99ZKtEsp2qnn0tVyKaOJiwN3/M9xMtmpm1GUXCYeR3L2Qz9N4GuZXgJ5jCvFW2hKRoSS+L
FyFFOIs87Sb1r6C/UBo2dW5T/7C5dQMmXJdIxXPW4Af9W2CmviKqfk1pcm2LZMJxlf6A/f6shpzq
ZTvFgLRvHqwCz3zbsd3/wU7s/F/6rujWuqAk9zmmVVXDsbEgKbDEsve+cEf/lgfnBZscBSh+brwT
bGUHIL95xpTqzU+lOvKgZq1/oyUaGfylkFoRQvarRZobOQD6g3puPKonvdUdsPkBJSR5G5eWO6lJ
j+EbR59t7pd8ff+Bt3d32dkmSTbDZZpdRVbGKsnOTG0f5a1h6eCyhGYuOGaYMBrsPipieHLMsVaU
6yx9nR2noluKbAHOuIBMlQIf0Ne2i//MdMC8eSfwWFqiTkCobjrqthU33GD30hL4+mqlgz89ZXPA
CrcHXOFGNzZOkshpkkbGVvoNtD42Lm9K2J5SFkYvGyB75msQc9XgVDzyqdJbx66Qm8cNYNmWEfzl
CZZokxeGEBhe97/mTX2QdStVfQXObHVQ1816vAp5rwJDh7h9O8wTdOk6Zh+loEu7JPyT45hG7/4P
ykzkgpruaiCwrf5sYr1HsY90FbmJYh0maFNN10lWY2Jexm0Zq5APWO0Wrve73cEO6Cpr1oUdkozT
9CyazBJiC9M0Q2fTaIFG/fRsSHjzF2/G4V2fDv5bPj+SywleHCVl6gWvBrD+uTuBAFoPdIGLauh1
U8+/TKmEXKoPYBb0n0JvsMR2hNK2CAlDfnNJmmj3hDmX19KLLpwKHIw5zt7vtY6JAlvyZO9/Ehd5
EvBloEhnOhJX1YPx2EJ7f/60e1n/cD2tDIH1nYLD2YE8gew1FpBMeLikwNxkd8X/I9gRJjj2odXk
NExlqXtooBIwslmmW18/m9L0j/rmAfsFOvm1LGGqyWU4YSEPTO64YZiOx/vAvFMiznXCw+zscS/u
vgUzJjo3I+dpSjJ/h9yA+UJzsU9eKhkALynp5SnKomEbs6P/j3wGAgedRCV9yo47p1Yo9Q3NuprT
UvGte5qZG5158Y/cIvDRYbv/5DCYBod6h0wrshaXoKa/yyCqNk9PJqVucXvNt3MDp82C/aGaJM95
Uz57st0pXWo1xUBpbEzUIqMp5X4+0DtCQyHpchd/noU25tzbGNNKEQTW9bbWvmPaFke8zBHVmK73
BPma5VYVJoit0DzxXSfx6thMNS61W6KsnXqS74xjo0sXHRSkY/tfR2EWATQ53HgUqtndbmjCGkAk
LLb8H8c9PIi9z8ie/JYpjI1nYA7nK22zPuVfqG7LZ1lQMIrgI/HNsy2ygodmWfRKtgf9PHu4utiY
/kPZSKqVwex2Va1ZMIW9KBlxNBC/6oQvOBOhgZu3VdL9ye/IKhVU6jmmlLOgK7k8Z0MqCLn7WYu3
b1QHbY6v/PsahLtDCwBDWdBQJj2RYM2CEfnAb3KDxDkThscbJ/Z9VhAWbFwwM2HdDzPlGYsx11Qz
1WxhJd1c4xbb9Zteuw9gEXzSt5mPoxGhOAHGFeUiUa5MhJ5maGbSRa0Qx+e5jA+RB44lOjt7RRPZ
qC2u2Uxqa18fTRCs1BgjpfijkMUZuimnBw/CzqC/cJckK7q9bpo/sLWFCJ2FUxz8jzCxWUILzAOc
/YzDJajetWdFhu4IkW9uZxdteZ6DRlRNsHRTXEpBhwalc6f+wtceBCLipvjEWPOWGFitDBIocXOi
2cn5OXyIraOuM5bIrEsjFWbQvOIc0Jc8JLJWp5rVUu6AYW7jJW7EkxALf2gldOiWM7hnjG0CuMo3
TkNOYgqdv4PUIDpDPqVa0+Q4lDCQ4Z3jgCe4i1shjoWRESx5fR1HcIIOE3lWYWwVqJCw5OnRMWL+
g4EudXWxKDn00PQHE5w06SgUpgZIpzWvXOPQftjAxZwM+yKfrOUeMP91BplxyOTEqvwrDbLn2e5D
UXtiEWyiZrnM5Ct7BDmaKoObcQTsjlu7F59OnINEnF3FEmChktbVG/+9EeqY7EtO1Ou9/RtKCCHR
RIVHq+BxO4twH7hA6bQxLRhz2/w+1ZcaCqnAv8WrMtunMQcOUcvUqWzlatf6maxJqO4gbpMQcGMH
I1OPTfpYPU4bwEU/m8Nw6aOBwJw1xTqWCCVG2QPBezsMOB8DWof8nyBzxXPGZcZGd+UgAl13NDg2
TrL8VtINIckS0+WOo2b7g+IUeluN9l2Om0VPysKosqGmrdv1ggz3l8tPu/Sp4TK4BouJynwi5OMx
eLGMAXu7XtEIpSpE4ny882++x/qK7XcqohJcjKWHIPN2Yg1w3ng5mMYUVgV/VJOSLQheOUZIkLYU
swik2ilXrIOWenk3bFkldY01Tyv4U/Q+eAkgy+V0dnf1Ov8xEAbmwyAR6bLpSxlwj24MLKfCwkVs
JVeJjyP1LhNW/PRXEJH08J8kjF5wvstNrmAE8Afr8F7JUqQFx42vGUaMB7AoDofnUOvWtrlgjJ8h
96UyKFvxQisELA/nnFKlYnhBy5Vv66LV0YkGkr5FxEgRUPFgaUHymHY5uji7lSEC4uSRVW3wvi5M
La0RT/M3l3mHzj6brtJQQIeIPDYHeORHn5RxJDLVcdefi3NEQWmyDW4p0GEi/P5k4zt3IY04QfcT
+9/Qr3cxVbNJnPjH5kt38QouJ5HdvY76G8mW9gniKuJQPSy0uwddjob5nEZSM5hLS1h+gWqOpdVZ
pBY4+vAnPKAyI2MWHcfnfw+EbUgyWdYtLaNrD+h459vIaVyLvGGTcEq58WqfkV67rFtrnqUIdJUM
ALe5Rgd5SFWk3PxwziwKp0HCfzOOi1j+tHcXz/Vv20yhBhfHgq3s2a9peqplCrpbzglZ/qAN0R2c
w+9Y/QR/jB5Xee0Isl4CfeEYpaztao1XSzgwA3qz4jBUY2XLgHc6V3ktp19wIuTx2W2Dft05Jw8g
bXRDa4368ir9e+xjsmZzNsFj3Vgp25qWapA4LZr/FjN1mRNCOigKtM247/MFEJd5sfIC6Xk9C3CW
Np3ayWzz5sFHJcMRbc0HC3NaPCjabXTJuf2TsJbDVvUil4ipTSrAw9f9hXNCIGUqB3fHNY4pVbWw
wIR+wZK2dU2R2piuyFBMdPdPaZYKf489IvWGzeE2efVdUXd7LFdGe3ZOAIbCq3WOszllHx5lrYeR
XTfI4XlmA+6TSkA5deBBVI9D/evuM7hL06hGtDN+8iCBsqRcp3nLoYbJ7zN3lT0PafG1L4ODsaGJ
dIV+HC/i+4fCpvtcextrCq9PKQY9t9i9iFqPReojNX2eWtEYiRzlerB8rGJdbGBkLpr0xosDrvgq
cqeTUiYpoeZgwiC6jaYyWwi5JoqaT6LaXKgNB4x+2LZe84Nc6MLrYlc82x67U3gLjQmK7z5WWw06
AbfH2Vwd2br9EKfjeSjIQzTFzIuRXz9xqR+csjhM5XTHNMPbShYy9I59e3uPup7b9fxY0hEWi6aX
8kesqOj9C6JlSPIhGDfyS3T7Arzp6AOEN1C+QkDQ327XcJU+bgqhmp6njzwZnyaN15AABvdUrVBS
2HExg6Q7S9J/WTDAeMlAjHCrZm1VQTGdNujgSFz3DkaIjDrMLtqRGRc3Ur/6S2z0ey4iofHQ8ovS
bovDV2L0vytEU4WtfCWUBng47zxJ1L+fDhfizmSZyxz6LlGdHfU96wSy9cjAZNc9tCJoxdpSI+Qc
QBVO5233R3Wpl9t+cTfRkZVfji1wAfdzHbWjTaPL+aYHJdtgaHqAjB2B3Kd/WJBS+uSvSK4EIH4p
2TE/tQ7WkmczqYG03Yv+0kBaZb8tE6Q32jJXueEqfPyrvfB1RT6Ab/jkqjbUFmOurrdrmW0GgRBQ
5PL8W+e7knSi+xaYevFMqyZDDfJ0KilgPmFNKoc/kb+2KeqqdBNpAa/Vw5Wk84MsuwbmvC+/5x4e
GtxSfBNsUytJjIUvJafX2BojV9jIj4hqHZD+b1zI+++rycI6/TbTfN0g8/nokJ9m8Gt37rg9zTn0
7zxapvJQSZ2A2mTyakss9JwZXBkgqhcz70NQDOW5BoEU7K7WDwWMy+9ADxEJHHDQP5mjbU6cOnUi
lPtJ2dTU1M3d4t2d2beN8yVH0tI0bcQZOUauFotqhF7I+f6uJ6jKsYIDVsqy852ecO/GVGkvBEnl
E9CC4p4evPluLHri/ryDxefW2L5mlIH5mdsOL/njPG+OxrO8ifjRc4b6QSx26Lhd1mfFRsoDcBmm
thbezL5zHLNb2GWvIpjzAXrZFZBKQzdn9EA7Bz3LAtulbknNYtAL0OCyNvaS9cU6SQMCUNqakqBM
HOA8U7FCB67pryz2yY5F3BTcRjYEO6snafZrFlQfrV1o3tvdI3NyeuNOCwSFtEOIFhzei7KWh0Di
Z4mFUYCkomHWCppiEgs6DIrhWoyFzzuUU1puQUdvBcHpslkzzcyygn5Eocnla7JUw9zCjnxTnp8Q
ctoPoKqyHMjR+Pwxngj0vly2yzQLFtrPNDwstPP/wrCLHkbYJ8JqSoaQrXu15kcJ026M4KtMcMWv
YqrOax5DOH42re3WPG7TyBoqz3p8RUQjqjcGmcqD5PWwcKQDYuXOD6RVAoloHKwksNE2ibUEGA+w
/tpThwAKp0CA17iDGor5W0tm3UG+gFRulh+wpDhWUwygR8WG6JLOByCNoktGOvEcZDAi1ygZmBCx
GJQ7qc4uYYuFNebIpdfsZLmlwyjRi/rrIXjW9XPNAf4No6z6RJvd1OEr4QpEvYpLU92x3WEoSZpF
bNDKXARtVefp/XHHn/RdEQfgBJMeXlRWxXi99XacFjbjLY3p/OTz3bnXWIdQk6B5vp7yvtPlcMo0
4/PlUJsDRvP23FnOvqA6UagDqHS2G8uOghP8E1JY+V3bE6Hed35uKrFd6R0S0mV5hFW7FM4sdFRH
9ZxlVs1BfoCCRUnnSsfsXDu33T4Jm6iYGn3NsbOz4X8ABbaBm1p+Zp/GDhZChfB1OTunCkd1cpb9
7Ws35zuO6PYRaIcuxitiBPo6jji10AsSfEmHYEFDQ9Ojv/vgDNIkUA38hYuhLqoqhrsmjPy9yaCe
RmTaiv/ml/jUL0U7Pif2DdlrYnWeaLP22ISjpC8oe+kDi5Xd/XrBNR1GDcfmN8T6Zv77o9wbHdBT
YIDFBq+0RgKCdH94h4XgtR0dVUmMpPxYI8c6j8tF0wcf8xgkJ1+2LSLMyW/7FMAfmruKFaR2dm8x
A6qtsTaeOZWE7GwI8JqJWNtG9Nml7ZoJJcLByWVsxUsNfdNrjNK1UrIlFUTr5c7baMnumBQaLSO8
4fFk723zlV3bPFiTE6MgqpMKfKpki4o6UlJuxaKNpood3MafWK8eB0c9i/WRRPnoVBdmB8+ZOYec
i6puphMYuZ+9o/dYY7ozshKZthaMftczyzyIIVWk+aAWSPIC2RzI4Qg3l4QxJ8aor2rs16KquHPp
/T/Tvhv4gZ8L9NoRmMcIS3YoA82b9nw2UjbHY8HkSJWQPt4TKy8nBLiZ5AI+ci/7R7TCwlUgsNfT
UMuPdQ0h5KHwevH5hu43MEitbh7gIUg0NAXO7aHBnP/xdaOfmysNBdvA+zcdmrlsYRDPOGD+4bJO
RYfcCkZ7qRs/c2ivClBL7EZYZHP9yvqipvoFjLkAjNNGpkao9OD0FnjfPdeDVubRAMqjERCfDxqO
CNbWDX07Ic+ZMYVQMQJZPoVWKrJFHPn7yZlaue9H7hOHAgCGg2M8hHdmooTo2DdMu2N5NGrsHe7E
EXfdlI5x70nCZGPKmHCTXNltN5znpHDCBD4RArtfXtvF/BGl2wr+ktYRLw5TYvhcESOzOSV7/kPN
N1U9hNxeDDX+qbD0+64Ax4Fgs6iheoNNm/4zSuT5Nsta8B74+/6U2vAq0zMvgkVbibExkc5ad8Xx
FwH6HJV2kx6q1n5i5rukq9Tl7rZW8WJfTsZTFOdakk/HgHylNM6MHrZ4IlnZCXi8tVolxxrU/CsP
/4NNpgChwQXMNNbG8WIyj+mGnq6/wLml9eX/3VP0yEAK9UBlhO3OBVvgjDkIEfGAIyBwcUowMgsA
oAYKyFZBgcrK65sOvFWvEAPp74Es5LDCNk82XcnhAIzbsjxxibOAaybxmg4uMS8Q5LJjiOKnZlZk
ud4Qz5N+jg1ffhxZD8t9uOSEpsTYwluMNaDyHFeBww9/ig/6ht0gb1gyG6H5KHJpGKMeXXUOojfX
rhD/Y7o5C43qxWxf61S/yL5vCTME3PNl7DkbcPH15sX95PmWYkFb3ArPqPn1L0LrIC4O8p8+4oIB
irCTmTmCkRhfqVeb0PxzjUWfqsaMRQZTcsTN4uBNxcWPpz2kFFRB3yxvx2k1gkjDMtc3zgSrcskg
uyVi0bEYZqAnfarWOpqTHWWSU/aUJftea6R4PSzBqMuXwVa0jli2oxekQ2G8zvSGorQ09Y1shFKw
cfS6GcY36WlLq1pCPSepDu+NfDfJxmle1AODhVR0jWUa4C79RVGdsFHUaaAApnrUK4Sfb8jvF7X0
aueiH90j+78hV/7stprPL9e+sVhvpUPyxM0vuMs1Wz2X4hWJZekFr2VQcOmpjmOMqTOWJk69m0rf
mHKt8FrH/BT3U1Yjss+aLDnYRVnv/OG9pdEaFevPkyA7Ut0PzaTj/OrGILcl9WjXEMK8EXkIGNny
xkxR79m0VxllMf0u7QI2KQXkyKMzyZqS6LAnw8ePyDyVzcZGHBK3DmU3z1O82thrtQbX1gwNUrnb
dmJpCFMj5QlArdYYobvqXiNARqepSZurMbAhjMece8xQe6IG52WGu594DqIyaQ0lsD/rhzDHW+m9
nndLAkqkSYirtGJNERVbuzBYHhitKWVYol+XfgRhBnO557cv/f4/U2QuenwMqlI3moz3lQkMI/QU
aaFzZC4u7+eFWRRevhl0iBDzYnExeM/u3UlbiQhRBj/ive/e09f/VYC9tF3AvRSBWY1Jc9IGACLQ
po5qDw+G6YZpCxsxYW4twI1ZgjB1D20fphCkct7VXepYWhTJjTKCM7HDr7Osi2LyiNPasmy/Ij1y
2N91WZkEPMMUHjck+G8uE3IVuUEdN3PcdOvG6veo6YPuzcD6/27ToxVTpRh2nsDnZl03zqddNEoz
J4HJonm3bxjLLWoxz/pJYRW4517mLgFA7jL1zXH9XfIF+XrCOJ+s/xcL5lLVsm/vCCGoILNJxUVI
nOXFj9O4vKi0tbAk77gE8NaBInZ3v90mM3e6webx32TWrxedFyEHj7F4moYXmgOe7pCeazHwUOfC
apYgJZI6oL91wgUbhBvYY6y/8cq2Ky1LS/OAttFNQgmeY1Hd6uGUIaKQXUb8JXj4ZLiA42v/PkAF
FxXEObl8HWsrpXFU62+I1o01+bzMh7LH5/D8XWVVQctJnkxywKoAFURQg0pSNMCjuvEZCb3gQ4xT
NQjLM6fBOS9sdDWNcPeBQozrq2vhciRYRGKM4VCCy1KgT6989ERKELgK4fgAM8HMhyzgf6r6ts45
D3oWXPG2cPMkYANUGEsdFu3w1JxjIVpUMl+qaynXvv6vU4HI30nvX8QQ8ChmKLy/1SXGg/KiY9nL
7ohNNEUhaVdje+uYFeMRrQGsSwXwHIj9JlFGmWX9E6y1oO68EN5N/FDywA2J6NpxjcTWSf0E53p8
9NNPgt+Pf19w7PvBG/konNO5puQysAfD2xJiJ7IrRhYrb76bwY8jZodvPzr13ZNKpi8AOTp/7kqG
hK+xIjdYzfGm8OrhxtVVPrcJ2aC6yrlnlAJZJnApExrvMNOiyUMXJkurd5pPHQegTbN7sA//tz1G
cayoj1fZiXpWf8bUuZOqKNHe59Hqsr8CvVFNQBJgtgOlrVLM3c4hivimiMoGmfX1PaLR6msLGOvF
E8x8inXpeAkJ6iIRbkyvT+heW14j2RMZ7aQnYGTcNx6LTBCPj+Ll5Ssl/IVIljGhm1XBfuqFZh/U
PNa3EaXNFG3cb+nWcYb1FLk+sYEfY9Z9R2xscGrf92TWktKChtI+Ni7r+i3MWIA77xlRTFwPeP0w
CYyldMvVV2IvVB56xn0zsEx5V3kfsyRX4py2MMjmjxmN9MnDrN7O3A0m14ydfUu1oKKY4+AwK9TQ
F3PtXX1sGevdo9heU3BYiODT9LK85J0jTwZHb9nmS+LyXYPHTJ/iTgtOVwhuIGkRzuHswwmpk9bi
NZ4t5oehywbkfbokO2ap5dg01ljoE8z2M1UUU0id7Kie/qDTkKe89wshqJ6FMulFxFxdLPoMdpLJ
6OCOOflGBFExTdYPN8hjPpnKViuMSJ8xTWa4Q1kY/5/i95cqDuc81nIygFMsd75u8yYP2uzkslkI
i3tV9nJ7ugNBWd5o25gGSe0eHLRVfuJEmNajvzYJYS7z05ltUwKb5tmYt38yL9bs8Ba8XihmaQ6M
qxniOMbOTqHt8OxZ+x8W9XSxPRno4gIb4deWyw/bQ4WyGXlwdFal0eH7TZa+hL51Z3wGg1lzlCx+
Aj78I/l26MlujW4cQ4n4zzW8fs74v7Gw+RsxOHi4Dm9PNltyme1IBdtlMW4WAl7i179Rr+KnoSjR
whMTrSm8mOBytTt6vRqcdUkKDL8CIOeSoWn9A56tDsJF0CdyUnEeGMO99sqRrSuOBgpVumaNnyvB
XnmVUcCGzASqDnpghQe6eyN3xHQyh3tWV3Qu5J/39vev3PlaxRlgEECf6YBk8r+i3OZfsCZoHsQY
OR0PNgAMj2Ce/qNoVcp7vh/7KcSLFiYW5gNnWlHevDuj/f6GDQhHC/QiH60o/rESAMz6esBZsiG1
Llqf0ax9EAhPl4KpSBhVAopnWP6QdJKqZ9OY9a29tSgk73kN3IMX6780hW+pJV7+lW+Mc7lxVhBv
YJWpCt0lnmJtUohodNfKuQUB+WXiFfyg2oBGoyOkWKAJmMa0BEVur7pvGWk02xrEZuRNWk+nOC8V
VBWyBHLffmQZbVT66tthhRmB1SNqm+2oJ3uFus4LefVsjDuTljaS3/y4RqARL1/D5TfdlsC0/Fl+
T1K61NhsYd79z+TDjvhoUVxGoP249b3pT3NEGbyR5s3f+t+WweYkCs8eDGQyfFN7v4xNf3nAqWI2
ZAD28/PGfK7J2MzBdIpso+DY4Rk48WB7h41+4Oa7E1obqZgxFO+gfnpeP8kYO0lrWjP3Nf5jrlub
7v2jfXG41NDxCUFvR9mAkps4GCkBLq3hEohKLwTUV+DhKCyCbV3MpkmI1Uo2cE9Qqpvx5QDOonP4
RD5fpOvzAxcDfPpsf+D/lN2B5ODvKe0KzeDOH5Ip+7Oaba5u8Y7qN249DQxtr1NOBXU8vrD6kMqp
rjhO/RAXbW4PavjCGmWD7Ijc8onrN687gsF/LKkstv/US+fGKfFGfSoYL4U6Sv3vrlDXqBMOK/+z
gFRb6eUHL4ZGBeuCuaxEn2pMxzPXrZeTBmYRvRgTp3tcs7IxFUwBS7SQMr+XCPcaJ2Mj4nSk2uBp
DdqaY+hqjnJMcfiilzOj5lHZTKxY5yX84r0SFWbbo4qaBFxZZCVZ4gv9bUFGIGS3cA3fsOfWoLvP
r4/1AuYWa6a7sHN+LOKJsZBXy8Ldug5AGddOBafCZ9thtEr3OGqybTjZWax7DOOXmYoLZXtj92Nv
680dpq3nPHMdAn3iz00zr6hoYCEmzHj2NiNPlhIb+02eo/qCHuqj8Uxx5kzA3y1cnC+xX0PaUTVz
lrYcvGKQhGHXtA0vSFoMkZkGjzFSmN4ZTvFFvgr5psbwD1faESy9YkqoDUXJlA/stpFYeTA5S98J
jvbneKuY2dYYOtu5B9RgwPaGkn+Uu5xsAY7OzuUPzFPsQB759jV8vf1APafZQ8guYPRUOREDkZbU
S7/mSdEvG60if48U+oggkHu0pOntHcrj+Vf+LmDjvEAhd1sgVd7809p4dOKv609OqiyjusqSZff8
yqqmHWvsGysya5sEgvbYVbxoA2PejCSuoohZ7IEuXvtPLQ2lcm920qmbhCtgdvC/pPwSPOQzrHoV
UcfZ2Vx3vgUCCeigTsIB0OmbItX/J/jbPRfgcfQruPZk9BbiwTeZMbYIB+L04A1GvCD45kSZriMW
T64aRAuD4QlywgtKKZGJ6cyNucuu7aWKL0TONIlfuTfl+vfToCWS7II0MYXJOWVcHs6BCmpHxJVF
gyZT/A9x0N2I5pPl1a9uNt7nS8e7+C8QOqaqLQX4fCyVnk69hhHVflKy0MDsZjp6pa+j2GzAxJxL
0wCW/Gb+jhztVIOp7hXn17uC/xbaYZzx2JXmCewI4tf1wF3pmSE4u13Ytqxg+dXnYpu8NpAwz4gS
XttpuGNyRBXYUUCGoBulHhBMMKlpUzIPSx7SINNb96tsD3+R8QPNHqOecbf1QpEYVZzwczawslBl
34gE7qTSVNBx5Zyya0iVraazjH50WG7/w+zl6I+91wRD4fChCQdNgqIro7JTk1Rv+T4TwK7VoI5s
d9VR515mtZILF/ojm8mB1UwKe7nVliIscb2ri/dmbEkBpsgYZ5t0jri6DqEG0d0R281pA3qr4qpY
F5qDlvNCohJ6I6JkbJfieX9GqoQPukpl9tXXhIs7Iwd2bbV01m4BqOeRT09K4KXJJX6RvEMa+b0t
Uy7dEIhDPakicPD2m2G78LEGNqU12D+dAg7lzqwHURtWmy8EW9VmHY3DG4+Vh1af9uvuqblnro1H
5NpiGHmspIu6oNTko62d8ldTX0mH01gmBhwzue8HS2rtVu007Lgdg/MsvZ3ERoNOAlOCfSxjdngo
Zlab8VDc3l+u2fCF7W6LMwLtvenkWs9wMPoYt5ggZhwoXvg1AH40ZJl6O7H/t85vYUK9ZUZe453T
kH6UReufUcDHuSjl01tCenN5smxFHz0DPbQQAENpcUPW0Rg3KjKyG8I+ZhIhQTZlVyGu2GM9AZKW
zkLaqJSbwgDzbay8UF5b3Z+6/2Axn4Ex2IK8OWnENJ3hAIjy/s/AQXlxGiHmp6yZNnZNiSEU/F5/
syW++KinhlO4yc3wEU2WcrA0JzayvEOwUU4XenEA/6idWs3Bnxe+Z8dP9IoodgLz47Fcl4qfmIEY
5AV0ka/nQfTGUWFkJAjDj2upzv9SHD323y9JqjBIU1ZdFxIFvicvHWOXx92RmH0jcXOAuZoDxSbO
QiL9U/8D1qWjAh4OI9hFwcIpbfzjUkSmxRV50rcSDDEz6EY3QEjfigAtaqrqlrnAv/5qklKI8tYB
UC7DCkwwf6eamLoCvJLrIfEON7V9yLeUR3OYdWdYLD3xbYdT2xnBtVkOXI94tS4i24FKEzhxsgRb
a4MX+jc64S33W1kElT4aoUmYBXiXpuxJyyIxdpqgRWDKd7+I4QG25hruTmrI3BqauVd20/PQ37jK
VbTVgTsVWjHwUKlx/uJdaWeNf5zWdFHKiI8fY2SpXx7ID8aoNp6mlTnYQf/S4RWHE9BGu5UTbayV
kLb7iGmRwzJ3KXHlB2kLA9uAtp7Pn/JEq6OBgWzAZGNRRNiefbu5j04HYffRMXcobNfoaoFjcAQQ
03pJgf5Yk0HjQwOg0i/FJ6woMynh2aa5VdpAsANdzyTDGTiz2Nj3TsM0A4gLO7K+4I/BctKUP91K
ZjUI2/ZcWyFrorkqrNvOH2J7u9jOqORRH/hEf4oono6xAMMMrfRpPibr5fhBkwvoZFLS2Rsu2qTw
3v9sXdHTH/ahVydlrDvW2Q0hE9IZoVhGVL7NlHFH79UNcTcqltg6DB8Mw1pHoPU7xAfpXrLH3EUa
tWekmbFJYQSzmS0nSMbtnH9xzzSOL75zPIwp6swWYtbdziuKu+AAoym3ylCOcNguCzFrIepfKzHI
vibdqEe51H8rSFqtCW9tH8awpHc0eZUEgkA0PumA7q+mJ2Rjc78ReM/kJVN+Qg/XwjO9pwwfHVy/
+9ARaMmluWOxnjcKHB7TPlzsV+swCpvNeP0kJbt0M2WhIPrEC7vtVzzxx/ooPCYFuXQGlzxCnU+W
6K5mby4Zboj6oitrvUmFhqpk51/q+8pK0nN48UmMRuT/dX1iXo8Ceze+J2J4qMtiUduMQC8Nodfa
tC8MpNeHbGQE+KtbrXOK+tsuw9XjfngY+XfL4zP4mfccaNBdbDh7UMCzYKlYOH8/5au37F61AYIZ
3QRj2a7VkELIc13SwVCNM3Gi/HvsmOpq96W4nyhyhf7U+k26sRQazViZrtD7NVl0uf2B1KdwytVt
s9xHuD+a04ZdLelGYmB2hcbP+YaioM10ITy3f7kqjxXAh1ttUJDMzxAPixZ9IVjL+ghtowkL3adL
flW+z1DKSP3DXRwerlFhsKXCx0dcehecHkMoKjvadBBARgh/WXrcCPKAbyIPPFUZ7qiBFMS0rZBA
hoLMkCmmbN5Xal4jcvT7jL63pmgKOe2ed0VEOzIp+av7Jo8CjkmFw4kPOOHCx4bNLs0YP4Nmi910
ufLvvvkDVgvQse6DX4hJR8mBSjW6yUpzMl+f2pBdQKzHe8wslVBHip5oI/+WiTULGYn4RArj3rta
z/uq0Ii9syaBt+eec9uJRI+qIyWvyCVir8F4gk9TrOJBavO8cNHjbV6/FZJTciElVPX5sLjKdB6n
LSP1kU+W2Ol2qU/lN7NZ4hQMfH6d9PWpWkbauhlmfY+9eWTBBirjsrEglxUW+a47OxlmYv5S3Oql
iIAPy5iMhmg9BU0bCcycEXpdyxTpb9TxskJtFo49htc2mJ0Ihf0EMKCxZg8oa3rlqhC/bKomQ7Fb
aCc2Sz6ty+7xwgI3tVKdqrbKMegjH6hLVmtn/Rl3AdvdQWVsjX0Z8Asr3mDvDJiu717t9AdCAyW5
K3uJqNY3oQBh1pt5acUeE9Pp6LcTU6rkIBSDdGRh0nnDB6LYygLbgOXA3qzqnHGeM/H6tBz2bjBn
9rYvq2rdfXfkFvS3mScVOOQLmVeBP+4/wM7V8e+0Y0WNNg61rp9ot2xJ1ASkV3Ruy1aKWiw2wATB
G9RUD+Abo4sBV6DM3HUocak60sgtOhYPNK7A/dsTI7yCmuS8vXLeQsB893UA3b7yLIwq9uF3NzLR
0bgk0PQlbZwJDXB3f+SsED66kEUe7wXUYRB/HUwzpd7ChBmVwvLi70cylESMuXdTY+pQ8aQmUYuo
Rqb7XSJA2r7mujqJQbtaadec5GFHhCsF5U1+TescFnrR2GStX2N5CxQHAnFmlCFBfta9vZfjioAF
EWJzit32uLckrTNGtG0Usu59HBHyZZjrHR3GW3iU4qZm9EOmKp4PBbEWYYV+oyq7iUTPXxTSTlHU
Zok8tovUVJZdHE89zAMw85/AvTt9wfHPXT0wXEM40S+94WheGz34TaIhfpILSE+w01xj+i1uNO5a
obkzecvzzmcjY+Lw+FRGeoLItkn0PdOfF7bLQMOlC7EztHrAjGYaDywB1yupyTthIQvhr024rAaV
S8Pp3usxRcwkUln4k36zPhn1Td92yCI/7OCJGP/SM3xKIVPEBQPnPMWgzqEpLgl56EKLz4OhSo9P
N/Ck5CrcMIyzabU78uuWdwAFjskCGCGrX5t7Xvs1pwJUg6sYQDkVQ8OKnNVhDrswbV2fWGLuNVSx
Mk2xvvo+P6IVLJo9Jh8YJbFwCnHYgtQnNaYV0rFrK/C1CsiWudOPWs+11sACowkcaU9KAoLJYQdB
GQ+L0nMKKBX22H/31tspjRwX5gDJMTLzIYuoeqIS+L8r8exc03BiRn19Lmd+xlTTdoHUhkCAELZI
wtB3ioJTXo+rdQOPJDM43cClz4KDUwhvhjjJyA48xut6481PUwI+JD58PE218yoeOicjIj6jC64A
hPgtfiZDQPMS9VVY6wV11F1LR6sVkKQnQ1ZpWEz5D2Lht4fzf+FAuBe04Wjn9mOhxx6m2XvrVSNi
iZeP0cCL2NYT5h9xo7Dq9g4scdc4qsRTpfvGbapVPhHyn1VEDPfXWQfPLOSShmSJh6g98jGmVJ9Z
6MrLJ0PC28cmEytE5VP7vqCoKU8s+y7+JJEvJMIqX2sZo78P0k9M687XJKETbwr9qtOyTKjS5oiQ
zRlBFTVikU4bQlGUgRVHllacBCiLLHmC6pDlq2q2jpXjewv9+VqSVxUcYCvhn2PsYtXWC7/A+qS1
nPVYMKCMIFv/cOBpMAdLERefT2muku3vrN/JPxqVN9RCwsUVv+5UoRD/pRk4WijYrcULTG3OfW33
lyG+L5h8nDTa625IHObgAXV0Z+bLUaSL2Ral1T9tqzSzJ7Yjl9q01DzHKCbYShGx1aF6Ebp9QRZf
Skk3uy5ZXciOM7lz/zeiEhLu3kLsqHZEEEdPumlCwnq7DTDz/XvkTly/CedHKsOiwqMRM09ZEWC7
JcEt4mXhPladMAHAsahYgWo26sISmMqvTkZjldekPMZJmBrKPvz3qGKVV/Ig6BBXa3/YKJYNi8L2
qvpKYMd4DSJPhiMIPjzhl42LmurzC1PDIDg7LvBCKww/4PVfi6kTwoPRMLoq3h6xItsFK+BYyyqp
wjZarHflxkg6drIlMks2a93lZnPFi0JDYeL9MZNkPm34q9ljiMlqNYZhl6y+pmSTDENsCFfhd2RN
DMdVJAMBMSSXTn717IsD40tyWNWDHn31mzeE9iLL+/Kw7QRSNURLLYnbOoJg9Q1/xK/bk1rHDUq5
AbT97RAbUEe0ZFYa99Q01hPrer/1lhz8rtT5pYJCZvcACTOyxnB2k2MHntBYgjxgkpW9NAAFO29V
XWo+GIkd5pT9/uppYeagGszBWywrvaTQq9SVy8m5NT/GWVPohFfEyULsSrQNJ+fRW1t7UYHdhr/q
CyYZdCaDwmQEIEKlniVrCx+RWE+zbc9WgB3osUClDxCRK2s/3C2+Tqee8E/sG1RoJCmnA0KVLKL6
S9gQLyDY0bRTU6h2EetpckdJvOPKaeQ+MYu2YTtMJ4hjPpRFEGjG5sDgb88R2gArGFqlMQcQXC59
job2VTzXpiyRmbfxLY/08mlyBMsx9Ia/8Nx66EWnVMObMwHUIewrrujQRXuNMuJgJRJPvXTqreGU
WDay1ox80l6W0jjyYoJixJyPKClLIyOop7GeXBGMhYAD9/A10bEBIxHpck1WIlrDu1sCOwbYVgwT
HwEHLrvFcjS/fnP7zBeBrHllQz/WeqJtIEtax3ktklSHDjtxEVKPxK8KWuSTYQVr7vsOayFUf/rA
e/q6whnHUi2yHxKoo1fkANOS4WmFC6icVJZmV5Ny4fdH49pmr1b7NdmoQFCjOZPhJiAXkSFU1+Hr
eCcGBDAOYu41lVHk9JECtKrzzeCX+rEVgES4LtGIKJCubsieSUDo4qMshKUOSfWpBiUTGJUjKLP/
1lmraMEjkmfRDPR4RgD9jYVP/Ke3eqR4edqCGOJ5bEiOBBhV1U0JzHFn4PEmW+/DSaiZinFKDfAb
rLi/UpvAYKuamZCknFZ8WMqFa/fh7nKxu4w1NJ/xwsaU7XRBGmSTiM5xRmQV2P5ukzmtyMenGHr8
dnZopYel5ta+xSftiO4gnAHXaxmi+jFlxcrR+jwaK27WIWeG2JvCh+Q3KSJ1OFjYArltR72QfRNj
KcAO9aDQicE5ZqnJqCjJA3mmphFW25/nen+KuS3NYezsSRPjdkPkik8AqVIKZai/oM+nRds58tQ4
AfDTUlORr9JZY8hELozbVzmJJIeqNBorpMVOPRisJuWzKxDnh+JrJxmZGxlhBxYjyqsQAKH12SFm
Ekh+9MmJJl+i7sfMbw+htzQ2qhyv6ib6jont3pJZWLXxeF5VhdIRabvliolUFXgzTL6HPV3kDFXN
PyuMZ0mmeqVrTPEuzAGPdoE43qa9dFbgY5uHs2V3r7e3D/T1hCEcK1znQV96FFecf4yDM+Z90osu
dyaeVKkrJPSO3dDBYwOlMA6govQObsu4ZuMaCie2FjzD5r5LsqW6VpmUZmGlivVHox3Ud7w/90vi
sII5S8zR1C/1NmoPpbmKnUpHd44eQPzZLbaCsaXJYA7D3+ylI6BnWD66EkR0AmMFVHBY3Rsnd1gp
nAMKpCLrs+elw7EhkLPifj/Bx4OERqQxsNyBpBW4W1RqdP5uHsHnHWadj31sHR9ItthFkfw3ntby
tAtTylwNBkFluK1VPhGd/DF9WXWCJH8UwASzUrhyVQRP6ID+uLoCHTvagQkv0mvmtqnB5vEucw4x
TQX4eg5e5F7puv8FJHuE6r5S8vTvtjQajl3nse04g//rLqWMLT4Fb7P/fW+0fvzdPbb0mE2/vJsO
lPzkIMOt7C9FdK0b0HYP5bxzQhG5s46xfa1N8gHYOfuAgPKZwHbMgTHsOZSxe4q5rMuyzU65V0Wj
Hvbs8z33b8KPQ5a4Gqbs5wvVka2zXKQpoqA+n3DlEyYsvuiYzJPuz3aO6uBXyumXrceteWAiTHRY
2rvVeHujBxXTKhL4iiJkn0RAE+47lyvLgZwYuqN5FNHRwIqxuRaFzaKluDX9xbqo2a9O3h4r2d7C
UpywyZGzHPS2G3r5cOjqlEGMU4Krfx7b08c49Tjhl7Ji45CxMn1mwZB/C5IUKS6wLRF1vfOLZvBz
UnNFkYRiM9L9VIx/wyAnLEJEo5GEk7spSYh2BcexX5AEC1XJJeK2JEq6dVQ9U6jGqUuTKRTcalVf
Epi6kWcY8ZbiAtvcwirzaobIDHeoNjTOVb3q3kUaLEzhkYwLReisWqT+m/15eKMm/D3LTqPVS2wJ
2lKCf831kIm58+rnF4+aYqVK9g3IztCz89D2lU7qpCo6ePssSK8gVEG2BOIbuckfY47UZiAFKplM
rKXIz7r/GejAyDJNDJtnk8nqFLhYz5hbNLZhmNsqHmQrKUS5AYTWJH0Kuq7pL0sicK8fW+Hbh0yk
kKPcXzKqDgOZaZ6w8G0RgWL1f3gTyKPRp/awa47vUV0D3/2GTeAE1dIpCbUK0c998XuvXR3J6DO5
B4ieXZfArS8Rmb7hDZ/2Sg9eJAh01aL4BKRxc24AgIdf2xIKuvwjpGP/5/jMxBYtituofrvyQLGw
1YQjqR1dDaIinhYE7vWcj2uWMcO/EEVkoiH1yJFJT9JYcz/Wa/E7WLywVPhTo95X46zmedUS5S64
irWcffVpt9KpBFj4719VYNiHk0PAIoRdBfVRzUP5WOtnq+k34kZb9uMUdUCiqRygcWgYgblaOJ6j
gflY+EbyYOWpy7YDq2BE0iS/+Iw90/6b8ok4a3uSAZnAnVtsalm5dZvYqLi/FCJpLA9s4ENngy8w
SjCveW4x4YNodsi4TVfaYUVcXAFw6gE8Y94lpcNu9t9wYReb9RYnHf9pa0HJ8qjGSvmO110ud1kl
zRRqyZWAoSz76q/tObKmHaXdueGot0xL61YIkpYpbpMGazpv+VWRxKVGsg1wSI+6ad/pT93fz+/7
s8gP/TOIrudEXYntIcxRcg90SbF9s/fidOS/ymgH7Mp+iCNOC0wiua+jQa7GB9wmtHc/ErvwuEtH
fv25n0CictTCmpEcWPPu8LESSQv4E+Avvs4mJImTfITJzQ6zEcydfofYdNmQCVrgqgWnM8auC8h2
4/b3Z5sgnZsYSpPMvw7jA+NQzw4g8ZaFnuUw38qHf2qRYMDDwLCcFouYUwXT2Nk5HE6gmA88CPgl
DRO0OrEgFORSvI1lKXSq/dy4sFP7UbcP121kXyliHboeG0FBCvshtDQPJVAy4qeBP0YrCeu5hokg
xz2aWKhoNYc13EdhXKVFaQ+5Kv0t7VFiz40Bvvhz3N9w64Kn7gNfkpVbGeXCpQqQE/jCa+nCR39I
O7CBj5uETtJjN74hWXy3tpNtz+mTj7TUNQU5uXKJHFd/wH5mqNUHjSpgDzpijXwuWSbFSoG+qGS5
e9sQHwJUSO7vOvQO8DuDSvWJvKsXRzty3k5F4EedvnMDeWAjbG7mpCJRP3aHS764l/OJ45xJoS7A
Id8l4AHRDx06aLmMHwsayAPvOULhF8FoQMw4p155sMjI7/YpJg4vGkt61sQnl8syRPlOv4g/78zL
0nqDwpq3Wc+BYwEABVEo4ryJM9/0+u6mWpHF0e+TSomnjC0ilJIjO8EBIJ67gD4ZwO2eaPf/vv3N
TsuA5SxleR4aiMrt2M/1s1F4IZJZE8sBdU0oCxoU5OWAFzgc3c0OxZiSBAL+CqXVkFKCAG7WdmK8
IOtDNx9rIIdjrPkIXe5BZu142nvKIQNhYfsIs+MkJGW/BePkhrcvqx/ivvR2GIVwG/b05SEtn4T6
5A8L9PVqf+492qA+0KAJ8s7pZ2bLiyhdsi979Yg67dcI3nsXIS7hCSmN6nqbyHRucVsILwtygxKe
QqufGgPnAiQjAVUqIB7xajRDS0WtFabDZwpW4bpZhzoT0g1erUAn/70NHJT65QZd2eK3r3gStdd+
TkzBGqarQmm99zqWHl6Gz6/FkSQw4KKTb2C3/v/sld58/v30KPhN9P7XWC3b1g8OL5x/6ecJifbO
uzn487LFktnXQcRrYH3AUZtR12J5gwoRzPCvAen7PPwffgy4OsXW3gBpUdFIkWo4uxFMIgskK/Ns
ftv0t+CmOxqCxwYnHAqRlgj6ha6l6maB6p+lhLZhOUkBdY6MPz0HYDmOClXH07gtm3Fex9DL3e9a
uVEq2HrYNB9aisLFg1OmJA81o1vvjvPOFRcZJY5IAruZBGX4iBZ1SBflzPHlggCTs2v26lHavg5y
Uwvs1SFo/8Enuoe+el+SvbRlAFlzmUbPikQGw1+l4mQMNx+L52ihot99j8AOpjo8Z3g+Zi90PQ2z
UmZpTCufYmN8+qAijWsF4UpArHKTsi/A+/YW/NbnC4R8w1JoBfo6NNjhzJvZrlUWMC4utSXankrq
+d72yCu/6sGmyqXqnt0Mxhk0GP/8KpniPMRAAD5oGrS1G5rohnSHRPpmCRh+gsrePI+0icV7WRdr
nU2k+6ZpzeAVdjkO5bwbv08IH+SPpJ5MlF3FGQxSPqPf3uXsb7yClcYV76cN/KxhMwkjP1rLotL7
xUg+VjHEUXqU4BGi8oibE/bv+Rk+huE1fww+4Gd1KImPfbhyYaZrqX1xL9n4o3gMpQb/c6EasiyD
T1YWE8ECkIrakkM39ObCaeEyf/FUlWd1B8OoFKQ2BPf2We+WdjqrmzARZnZ667By6OhBI7yz9OfQ
0ucBJbZp6av1brOUBgskQj1yq5zizyKYDCIbX0ojLr+S5qPqTBVCgk9pWcAOUXuofavHky9XJ9vw
Cih6UJKVxCvEd5To6ymuNZvdXFzcKuryRyGZdbCjoS6f635ksHUIvQu7UJpEQ2rFFoxW3pSFW8Vz
Mu2Zgonpu8+0wz4pfrbtC6y1UD+Inf/Cb8A4Br1Ddb9/zb7YKRxP5JOXYrU/oTSq66s78qgZt477
3AYu0hBhoRHsC8tRWXTw3TV/Amh9Bcey2hGlgqSx8sKQo+8UWODcHzvBlX9pmmXphYohCqwTXcV2
xUeK327GMU3feD0wIB+qWZQ7bmjtDzVDtx/5V/jursvJeLoJGRU+x3zGcQR5IvU0ixmJWY7kDJR2
o5U2WHxj65xUKYgunJcHIOX37YFf4PwjlSmJ2EcWyCHfq0pNiAcNI7z8stV5O/oYWcU6yeQuUcw1
FHyUy44Y3uk+HLrI3ZH4QmyDLKDrvCiEwAaY/JW+tcBdQSBV4u9mMrOVIONpyFRPYnI2ifU5v2Lo
4y+8HHY/2eMynYFf/52fgOKz2YT89ClUPfsZH9EQPfxiIy3FqEAANPNU2vD6iMjQWCHeQic2LuWT
vDrNX6tfsug+1Y+/fguTjiP1E/ZgjdATVrkBuE1QT1L5n78kq/fsML2QJ7YwC+utUbr5zOFwXmct
kIG+RT6ynGiLQtt29WGOK0xR7sIjS3ElWxR0VUhAtiJ5zQCScbtcXIZuXKsfSgzPFyC0FjhERS9p
tbqrq/nflNdrAKF8laqKwKQtz24B1cgaja3mbze7ZXfTiOEuiO7vVxUPRY87d0r1tpULIzxog8+2
FlliOpcfZ7L0J50S3SJDF/4m1gvHxxmqthhDWT7ZxkIP8n1YZuZJH7b3+rJAMaEcI/w3fBQO4SBc
J1kNloqn9n0P/CHcKa2vx3MjS0HgpKvurDZr8Ou02+6RSX6pC2d0Qk7XwaqTw73ZbDbu/6ochIAy
ozqW+qIrUptwtVVc6fa2/sJkUjQ0dJiXqMcd71RVONC56b5C9K7u8QHOiG/DHdolSbb2IqOShNj9
XzWiK26Kp1bgg9QtWupDqX6mJwvnI2FDi49XnjrIS03VpLh8WWlXIJtZiYI3LjNT+LcQgN5G8uLg
8GCBI4ib/SOi8L4fPplZbsRZoe5C72A3kZRYUbhqiDiTpgK8ovQuVMD1UvWMN10NX7FICmovMd+m
MIGM/on4qQgJY3OQBggNgcvVbVUFgCMmHwmEGiz5am2WCCOHZrxfXm1tmu5l77O69k7E39rS1ccb
PDlpbHPhv7gPsYs+TAN9fky877/mrIb1hkvZldgNvc5qjRFYOgWdEVcUccujmRGLJ9ly3uPPLXKu
MWYVeOMiNU6yi3CS0u+orkOgf3BO4Mv1NYjJHY0utyrV/ewQKNYHmpmhzBptBaSq0FU8bjY5Ufx6
hHLtl7tjZfsgYUI4NJstJSAvxY4zZ6LnHE5BvSbnYtoDx/SkU/f1mGNGt+ZkwzKfBGxxOz0SIBK9
H6VHBczXIprb1Mv4NvbiLLjWtRbqfRxUiOpDy/GE6/ljvupUUK1bozq+e8odseKwBynXIaJaIitp
FCJsbjKMlrm/+N65bsv5pBY+HMzVA9yM+eK/wdBNepURvTQ2KcokdFXQADN4cjY5ixAWA1qfS26f
cRlh8yeO8smDAdTvxVM7KT3swP8fzpKEmuoghq3KKA1+O5sBnVGxGlVQnF3sqDFseev4LTTuVBM9
kHWTe1beuRnSl9XHObYsXui0LTJG/oTuAYs0Sz6Pto3NlB5BV+QzyQEouKFaVDIHGiuEb67OQyHn
QUhAzxVoEUoA0fGKaAoHrJ0TrgVBv6Sv+4IgcXoGJag2yFZfb+r56o0eXQ8I4SjV7M1CsRYuBHse
mG/b6PHhTcC2N8xZjE0wKAUQA4kXtZnZOoZKmAWNyRDsqq33B/FlXd3SIBXp8IB7b/TNV+YmT2z/
eIzyXCEkLfKZ5yy3isohxJc36Zh1/vXSD0i1FgT3JBo5eKq8O6lKhFOkFoSeeT3Ez5MXFj46hmOF
RKqX9U8ag+9CQxRaQ/t17PayZnnNhrAonBZjAPTF0YaEJbFmkr45DnJ7fd+q+INVHNH/vtkD3j7L
+xXHTCbI5NuGKREoKiJLLu4ujMOYC8L361iya5FYjZbhfsCUe84gp2YEodvGOLYUMbS8igeNlbSn
Kt/n9pMDCg260h2OGjTeMIlqr9qvr4IOtTpxtsHMT/UhNNB5tT/VP+eJHA6py+37rPDmVOQWqzS8
+cEDyATubLf80ocUNJx45jn6osRR6jAhCkkZ7hyzOOjvbN6r3KICq7CwDzROAkYIvboQv94vkMh2
VS8dZqWeQNsEklVYuoQXVm3RxwAZAzOQznEqXg2G0F2ZA9cmwo4pwtrzDFcpW6McIyUqNVzAqho6
w/ENLs0Sk/x4qafyyF6eG9f3f4fiUnMSKSI84aMzkg9io7QcDLZJ/3TSlboodCVEyxSZAH4bTyqw
iXgfMEJVBnGnqZx11hh+OZbnplKJWxN6MWZjU4icy46FaEUXk8bfQVpuXwld0Lqtd0gr8PbJvid2
bRhnnbOuhcA+abGt1qxHUJtrlbH9xdj35GmgKiWq8r/ltduETu6dkatTB7ZwR5UmMfJ2uqcbz1dq
6queBB99OfFUXjIa6RJI9ixtKY4jD7h/ICxZWfCSzh4vqu6y30PhXWP+a44DF/ACJJCSsHkdy11a
ByYAbAtbaDl9sAbx5xpMRcegHmNrTbr2j65TPPRRrlJJ7egwP5wY10Tz78YH4V8tBlbRcQBaZK+D
PxRdRtwUp8DjRK4zhp3HFGA4GrzRMkYVRMe7GU1L9+NoIy2fg6OLL5otR9uLiyEzjwwwdA96Cecp
Ibi+EhIrUddRay8p41SA6yXDmg733JrBPtAycOa8SYIXL3So2ya9ERs0lYn+gfd+Jabw7SzR8k6G
cYHiYli98yQOIu/TiHF/tIKi5YABCdqqAbHY86I/X7QU3KjoUResiuAZ205zKq49fbIVfjnvNd/R
YPOhnFiVmAqoFXT1s7lGozkUKYT2b4E8OIFIp1U+s+tTlqzbSPgm4m787zK9BBk4ThkkMn2oG4Ep
NTiHiSU/13RwNnsD31mXDcpcpcBeGLCIuC14sjp79xxHveqa7uTb1nzBbybMdKSP8SGS/oA/EE+c
PMpd7CcWGsPC3v6+9yT9t+KtK6RM5fgYS6dmAhEaVcZNNqItlSLQG9895/LUvwg5Qcfvw80+T651
T6xMP8iS8Sqr1bb1uhrHXIhHQCK27fe77pgOnFHs9HTPLEpQQ2G2dSTYV3s0n0N9Sqk7qPVsEQiZ
TYkUpCS6D+dBKS/qFK5MqERMDRpb5QTOQheNSIpu6JHPPup61I5pz6BJiWxkYis8UHJ2q+7lJHbo
OrKrzLoc6hXvLqeyOkDFWj4VDqo6d1Uj3N0JefbvH3/7W/MTvZJhp2dMdWAkPydSOujQhu53sQ+w
Bi4J0ciBh9GeXSKuSZw/wGojpmUkE2Pc0FNP10Fojp/2fPhTn1v2obAsc3fA6G4BKK/dTJEwaB1z
ETRo3VAFPWLkUOXwyPGbXh63yxsIq7bQ6w5x5ZalBTL+FgSV0B1E/PWhjXY+2YwAZoyb3j2J6VbM
iaLPko53MjkyKWhpX4vFwYlu+nM5xt7bSMgZTTCrcDkqZCgvWPvV+zab78iwzik9o+zMMSp3NMgu
yf6yTcblna5zPNOy2481EMkfwzIXauNiedie+EAPy0MC7bw82WG9J+YX2LQXOA1V6bylSP44novG
oN6AEoGC1Sbi9DLPTOn2KU5E1aoN0O1j/nclrltLH/3XVMrArkDvKZu6diOPmfKLP6NLpKNKAl4M
yMP5jfSDBdkI8dCLgB0w4dsm8GeQ3xbdFNzuxpyjFQY8uOTCEzxxJVX37jpxB1wSgrv9UH/ThGqx
yy5epRnvRjmMmRYOMVNL7lH06hY5VEU5DdRtRQXMC3ndCTH5AlvogVV4JdMEYeyRD5FP2FQ5ySvK
SJbx1w9TlB4YdS9iiEpzoq/oy//cwuqjGbW20xWLNXNn3z/YP0r//x0IaeQVcOA96TdbCX9aotMS
Cw/eet7f+6YNsVgFHYCd3AzrDqYWgyugzBEVG873+VuilnKDVIquztyV4h41Su0fUO6SSvuRXF4+
cc07oDxjCbCH4DZ1B8McM7K4h3VXUne5S5trVJZ807fWrEcJHRLnPen5ZkPzPZNz9H/XI3jaqZCo
iGjsdTXKDB6z4ZCSqN2QNYZNIFeKKEnljc+5XLnA9jHYowdgopsg3wOD2hjDVfPanzKPdpN08hkw
ivgMZ0RxDDD73erZoeC/+wfPHNn6HgupUd+I+Qj4xv1V7z3Dym+em4kHJXvdfmGYMSqrVqKkvouW
NUuUdx/zSbZ5Q+MQ685MkWum5BXezxu3g3kfPZPaqdcWG/WO1Rt2qMA0rr4/VuLAGdXryXOQJmgh
B1n65freNfI2LIp3nqb1R+F8AE/eQItdAstP4v0RimWQ2e5LxANA5F3OzcJuKJPsMvvBwXXkuj9S
7kVI7puxhZbmPSYyN+Qzf8FgR7Vl/ooOP+i9qB3NHeN+xvxpXnWHNBPRixANKVzDWUGno+FiIiO9
y3oeARTyPXTa3/2oHCMBypTD0RMv4mCEcwnxIbu3S6etD3Ii/HrIyz4uCNtUVdu3WACGfxGAEIb8
Ghpk+GJRhTo6jGAcqb9cuIHFI3Heh92I7fyYUiDLGEhfOgz3fuqO64AkatUPoo+a7NK/pCfBbmdL
0i9SphepD2iMgTAbrVu6xaokcd5AOkpcFgBIeKacMz2ZwkY8beiAHJyf29xrfKVuYPOaXUnxV1v/
79NZR8FkV5Fb6NCuEawT6iIXMQ/wUToQhZ6W2basEbCB4U8941p6/BCGkNLGbUzwnlItMOVuPHOo
D4m6cfktptYXg+NaYA/squ+BR6yZngUUW7bTx6LKMWnH2tPSZ1y/V0PFJ6TD0t8MQuyAsyGEhHlU
pGPSP/PO0EKwCUh3V6kklhDwyzIPdBkmW1+cbrMXLdvFonYNDvSK9LcMCXBEYRayjp0QsHrjikf1
L/CqWIJTFL9Oia4EYPgH3Z9KDSGpNvheNfxrDdgHcLY5uqnQLhx73DOOxsID1RVeO6+t/JhVZYek
0m+1QcfdAbT/PKXdDQYkVcBfscCsizjhOE9m9mWXmURi1a23rJ17P5iOTQvL0nfwPQgnSQ9AAQVt
/f8xNb8ya4wAGOv3WU7McHrwWfpKSR2zrKh3wZUl1DqhEz4gopk70/2npm936zeyGn5567v4UmnG
zHdm5Ds2iNblTZDXtwjjFIemdAxz1WE3zBofHWqsDcDnu1Kc6IFLuVzA6D2JuibOktznKYNc6CeB
frchvdKFUEoXIE9BnNdYRy6Ld976AhSappx1I4iEQovkH/Hc1TudLO+cuivnWzVzdEpU/2QY4W9v
mhLsYOXjk32kxxtMC+I2kL4JeZVNTJdKUUZBRxstx1ZbrOu4W6lzM6Ez20o/T3/30Iu+dq6TAtw0
CpdYAGZLZbYINXYAI4MXqXc5elAzAKLCjR8yrihNYBJp6FPVhXjyCHPdu4NvdB7fJ6bLgETnjN9q
8CxKE83NJX+dwnQaoxw21uM8DMT3c41VKAtOf0oULFrgshdl0WHbFiYmJ9eHr8nH1owTRFV9SufA
8JzpeN594f2gNm1TWUStCOSiIcTrY8nK1utm3zlKzUp25+fAIq4vSOdth014tIvDdUIzu96ob1rH
W8MV6IFq33RkN96J65Um+WuIx0fj07+FroIUTqExo48WovNt+7k9byvp92t5SD4D3Oti4XaZuKtO
VnUgSBjoVqF+xeVjH3iNFaqcdotNFjA5fl2F65lLXoZldaM7I7jHjUtJEeo0bXlITzMAZiD1Hy8Y
v0H/YZMxoRmXOyBxsi4OEOwkPmeeNHfb1W6Pd6g2Kk9sM0ATBroV+83rRtlOAq7sRfaTcYJSroBK
Fq/O35uFEa+dM83aA5PIBOdl3DpdOB1y3awl4uGpmYy/LRxOPkw9JC3Sx7U8n9PZ21IbtfnLjMd3
Zuz9vfVmhJL7cn5hw/wc7crHJ7dP8mU7CxI3tEtdd8+cmEI9myekTv1hKAjEUmORd0u7Zu/gP8Bh
dH7CMO8jHoRsRMlrAlSW25nZYacSiZF2AKGbR2oD/uJs/8mYwPdgudpfwqALTy5ZGnrIAePSVowH
I1mIUggotnyPvXjjqwwoZcSCWYJkXbt1Q8EguowdWtGMOKLVgUM53mHtLB5uP6tTM4T9mp1xQz1M
L1WH9g3taCJUUwo2jUz8geuGIHB43/eulRIwlyewMwBmHr/uTsHXFxTdRx8hsLsR2TfE0iWdO93m
/cLBZ49nydN5/3aHbdp9tl3l+VuPdWY5Acw2UK8+N7RR4dwG0BSe5+1UI8CjwU15QJ3yGCJDuwTL
I44Fs4xBVsrL3qcJK3XEdfhVB2H70yq/ORCW00eTO36wRtPjAMCuyUCnqVxjmyMgtDjTB4GjGLNJ
wDS6zx1TxEajaogNAdOJLI3OcG364ATjeq4arNJ91VN88bIL9WVKdJIoOpFTWuvG021WZQ4VadvZ
RQ72jrh0K8KOKI35JoydK5Qdn5NSJg0ZbDGJyCnfbnADQKd7DOCXGnuxobqA1KEsacocOcMMXjPj
IiYxgnlSvoS/CF1oE1n9kxjJN+690yOaStIlaPBsyt66v/xnSJDEU5oFmaArsc3+odB9hk5FcQBc
f13+OG9caKZv8B5S48QZZuQhWNfONHvIuk2bPgNAsnrGYm3VEvHTA5GoyFEgwuTE//RAk7hTlCG4
UCcKsyIoncpCnOuioyEOdlxySW0SxIqnFy6wrXBF2/W7qx5oRyptvJ6fCQC+z/Lt6jDloujMoQf9
3yFQfSJyeszq+HZUpDcCwWPhVwmFt2as2UZ5p3XBci2ShB3BYS4PMyE2Nq+bWzv2WOISK/3XYPYL
6Bak2/PtyYXSdxX6Rov4WONYUQVRwRQiWNkxD+vL97auj5jJNxFZHyBBWetA5zAMd/+KVqbARYIC
z68I1fB6IhN6UXjss6sr8syJsGC4zTC4cdXA4GSsH/E2mP+k9h7D5z+JGUMco/WBFLV1XmHMuCxm
2p2B4WbGIwAbZvsiNi9dDA8RXgrx4pkDdL4skm1n9/FrOkm0idN/OShNq5h/ywnsrIin94mo7W0A
s0mbiCfr6Fhsp27lX3GbxD5JywelEnhe49QDCGURJrDVpkc5LONTqyNf3uqYykr2IDnPGsOiBhwX
ahS2xAd6AOjU+YypLBZjH1zOYBUsqRqoPy5lpzanNkWydl5VGIOQAV19sU+j/3z44etklAg32l5f
UfV4Sj73u8lghPiuBKy8YOjBjl6KmKCWkzUazcOKKj6SVftwJEiGPKSTws2RSuXD+6tHTNEsXxo/
NggzFUhtqZaUKVDb8BjwJvnoPrcdS4dlc5ZiCYddEVruxAZ+Fhgky4u3k9B+y9qL74YPJ2TAPWoq
lBwy8Ev1PaTrK5j0FPMT9h8vuFhVG0EjPWiYob5H1X657+rsjdwS2TKESKMGMBgr7KpDmbL7x5MU
TX248KWahFEs4R4AwJaqMTOTztKeJed+eOPBx5FkBQW2B0qRk1wcR/jTL4+aqElyurkae30EzYgq
QWODYKIzEJyesJsD1K7IT8O07X3oOMGRE98p0sdiqRU6WbOIg7NfSAAit/veNaPrR6Ku/7VcF7qz
tham9XzU+Empba0spQf1leNMiO0ei6SUHk93xef7oO1o7jUpYhliLCaPh42fLteCYyI1bUOZt0rz
KxTSqDarqKM1GEAXVRrFoWv+d41VTuAs0EGuUYDdUj3OGQ0ySuJWWn6HlTHphAJ7uet0D5U4tr7B
a7dHQsqdw1z/2A4LxxiNlxpkVlXQLNBVvQH5kem/Hvu99p6ZQ46ubLuZGQJFlzEXJg2mbBeIz4fs
QgUpYxkLJnqG5z+5hJGiFmp607MXMT5/m4wleMCLneJsXWUA9RzscVwMGxXK0wpmFdZTb1YrwER9
rVW6du+ELbx/CKK2GHPTkVhFOK+uUohhsolObcfYZGKN75OlXH5zR0gyY+0sQ7GZVPJ1CCL4R7G4
5xA3J1f8AVMPu2q68ihe6FSqY72pkd2Di4/DqIeja95PtAPnTpIjMnkxnGDCQSZGh6B1eupqJD3r
cjKZ7VrhKQvOXyygjcscZFzmMudIqVDMoIrzOlSkMbP04dreNUt9Fh8Qc+8xCc3ESt7VFUNKxr/1
G8g70RAsabxqzUlqqv8NXrNgBsqcpEPspET7UQgxvGxxxm9xeEX2Qom0G7hp8e0KdfMFTNql833t
w6iRQ3uk1csiXB8L5BLeuclzl+a1PO8KHqwtIYq/lqSkhsmOVrQPJQO8jxQJpbDAHvVAUFYXLwjJ
QGIZlBL4EPHSkwu4NY77BfjCnPWI2/MEws7DqY3Qw0G0qc/6xEmf0CdssFrWOjkb5D6L5W0t2GSs
YK/VHx6hbS583LIAk4TVmjUwK1MZRNqLET8lOImgO/OaZahIVtSGXB535p0Ie1797nNPbpopZ4jY
Fb1PFeIXcH6oZx1jRhtrDdJJDne8PSme/gNR77Rjsllw7v8/dQECFO6fbOPjEJcKBAZ4VBqXqYes
djlLCJ2evyLBmp7aDSUUvSRJin0WB0BPugoJYiJHMwC208Wd5n8Sex35xhGBbBBO25xtvpOBUxhF
+XBVxzO8I2j+TVSROUOOWbmpwO4tDTRcyb8JH8KE3zMCMBcFFuqWTQWUXEsh4FR6DbdQ+JXpAKr5
Ozls/FiLs+tOsVAIiEsY52poS2XV2VG69rsYfqwLtXuhpRQfRAjul784oiO1vo9u0wdrdG9wkrwS
S9k3Lj9RAu0fxojq2xNL4oT6sWdtIITHrKV0ZnPIJRTsBJSdzh3PAR7fp0aHq067XZSAh9CRDD1k
5PXekO7JTsg99tGDKRAEjvjx/eegIJY5m/Q8ctl+iCo8fm1hW7L98zK9BZ0iSwZd5ZkMgV7W8Lwq
rbC5Mm8ZSRnSxCxp1DVKWt4Zx0OcTYb5lBC38K5SBvX4gu94DGoGEFBzLSfoR4HOKZobfFELVCK/
QrBAT/UjbtnTLWVcx06fdw9/tHphQ1auLf74gbDe7X9d40Bi+i+D6B0ayENVz9es+CCBHxqt19bk
j6n+T2qm6qBjYSvv2FO08YA06Ie47d6JWBZ/xuN5fT4DxRXS2hiEfVIUrtxC4Ysumy/y93PH3ffv
wUaad/naERnKWbMFNfUbml068vHvKW6APArDQkTE+Htkb5giKLLvW+D3Y2YbGkZwlZpwDha2sJeO
Q5fCUhfJ9YSL3m9c+xAkoMaWenNWeWbNoHYkfH1ELvTKJReS27wjxZ+nyr94AOeSH1TYUeomqJHa
YITws25yS4u8NgfYluJsfdj0tzItVeyVzJwh/WEC89oJmmYZPk75LXi6O+j2+81ZqC9K450OZYnh
20uXXnkj7kygBe9C3gaE8M83sxOrkOzJNf4b1yY5z2isxRXWTO/rQ5Tu6oE+58pP5YHJYlmwxC6m
q+vTNrP6XDi/x4t9yUTTCUKUyipofukz9veXyuk5xyuDwaZWa2UcQZgvRtYGqr3hvx0Fn69Fu8pt
VHeG8QjGMFLpqpYKPgnfDkkEKeSg9/QMrpnxBc+fhsAjXZyuQU4R3Nsj6T1xN46Mw3ID1QyrHN64
Gw2DXy9TL6NyJbWh4L/5SsIHwwBd9joxwUaA1hflXUTPNoqHfAfOAQPZw33KtDU10lRG4EPYdGH3
na6dbAHLQQvFlimpb1N002QOYMGJ8r9lRnE71S9s5sihPT6576sZdKl1Xka1Oy97SiZYWBRoNE4E
LHfC/N7ydWmAMiIcpSBmwAg5AN5THJqOuktot6Rfcy5cLzr4G64Af/YbE90Zfo0bIBOPBNraoIzq
spQbLLxRuVhm7i+bFN8k+X+NEarnddtL/7EjgIy6Iak9x0FmqYPEXOQGDiXhh4MD7c2K3bbkdMyc
7VUaeZBiAsIBVGkeLrqkIqLZlcPMq5OHD5Ur0wjmpVSQvK+mQaEUBkyPu1XMA5kDYgCbC2N2Qf5O
Ex3OKoIkq5uvkJPyPqjuWYH0z3ZId68hd0O8wmmjWiYPH+BnadlpBKoop7WyoOjPIyY8qXb9yv/P
qCkHak3J0Lwt0HXMDIO387SmLS0ZEQ031iIsg0tWfLfwRRILCGGfYCCfBvJAEkcBBP7OpQ+L6ZyO
oYhIMZCgxWgiOL4XCaOcMwN1AJrR0XF2KEfp4nwZq4U4hszHBcmZqGQMs0r5S1Fn9VxUCJ7gr7NJ
nAfF+J4Y9gVZoArMLfiXNElZl1hJIhIFL9g3XJrBY6Dv++dHO7Hqg5gHlpe3Q/nlzbe4l7yVxhDo
Nl4oyVsBFaWg+qtEQYZrRJ5fTOL8w0ssOZr2ti4kApnkhlOeCg2LqiHYZOUIQKek2c26NVYxQ6Pi
pTqsx8jvhP1etEwRGghu8Y3HXTTR8u/NpV9IKnggQGQduAnYPqJEw2inmEzfJTnHRnNHJZd+IRs8
TdSx1xH9rRtwmOyMqZ1h3na59kn/ME0wEW7kTPcwkJ07ayV868Gs9Sbp4eH3pu4wYoMl1ZZ6TkBT
NmfXibDZrDzCHq/2qZ5li96/5n6TmF3wqurRHpBHQUQ/nK6Toew9UulV0BEoHduxARrTK8GI9+XN
2yxEZKprOPvzoU3g7SnHmaLbMJoaoEg7WUEfXiaU97rHRTQNvFMk/Ma1wDl/hdL4EEeGFt3Wipmp
78kFbxJ+WCag73PYtRzQPdEBqGKXlzranHRMcURAtKPqLk9KQl3Rm/lPmKEQDvbNW5IDfb4BQ/Rg
iIIliMCvNYtyCXM3klgYJJqiicIPVODVBhPC5pFZlEv0lDqwRXPpvvz1jhiiHum+o+x4HhzqxKGP
NUNej4YuXPoyby1iF+6UKxBulc0Ueyd3y/5rG711Wo7Ivs09U6ciDISnRCDcjpT+iEUk6QIYAeii
V7kpBcyvX14FaMceJiZnu8DQAvYS3o2etGDeE9W1yOzWPSSdsasfCPH5LOIw1omIXpO3sfnOT5Bs
wlEm2J2x2Mwj6fNbYke1uATtYT69OBWda4fNGlW5VhO5ilhqDNU/FMxPyCQfIUd95UJe9yt3+IeN
7hmBsrCY5d1q9DxK8XxTXgNKZUEalSH1dVaf/v9Y5856PO1SfZ6HHr4tIZYUtKWhigng9VR/L1Oy
ko6NHgcYKWqG6pEwBWENIBcIezFkU2JY3yoUOjaggxL/8dDvn9kI3O+oNIt/drdyFVeKSAgHgOnQ
qKg0wIWKqYE6aLmtQdi2xbA6DoWXLStIHuZ3TLHCovWK1de2NFZlBzHMdjg4ApR1znQewHrBmuKr
QTgZZ0QtJ8SbDv2d+8vtXz/BInMyAURjJaYz3sdMtYvT7KlL+/Z5W36u7T3kwbu77wb+k3EZ7Pe6
+C3tiGE3fOEDZWy9c2iduJmtQWFUoI7nCFNc6PeKvcpnFypnbJCZ1t53op9aaWhUP0HJIkVrWBNK
tkJ/kVrFWrM2h6yveazJi/4OBp9OJxO5z8xjDgqmxNoLFqTh6TEZKT8b1ZvFcvBRFeEGFm7c0KHj
31UV9HpZs+Z+D6uhXrK5m0Fk+L4aCNoV0nuv88EonsEwyopzsLYgdSOaDHKlK+vPPdKJr478gUM6
/z5kovwuKAzc8/hxLa90gKLETiCMbbRG9GPTJmzLuc7GGfJaw8LHox/3ItR8IZjRZM4q4iITnUDZ
1fADpkSbrDBkHxJH5PzvoIkG6mEd64DadlOgosSJknRjS7UOgovLbzaUB2dVAM2vOMIg8vCzfKrz
B/ZNMTJ8J6mklhj1PbeJYU8PX1XLrCmjd4QQpVa812kCXTRI8B5YwPkeg6TEAbLstr7kBwLnoV8F
t8xVUi26McJgGM65xB17iyDkAIs4w+2+GJF/8G8EI1fERoH3YI8eoi+Ykjz40OeWarkK0YLCUQVx
4GB8GalijvnVjbUYIfSwl0iJInrpUnuf7Qn/fuHhVFX0P0RvPZgxJuwwi1/tKVP7HEUT6uBVL78u
Oa5xd7XhzUkc2FrFztp0a7lIQUTzYunMFIttoZeS1gUpEMEzC1PnQaV6lps/EOXynsreNaTR66WT
1M6vBBP3Tc7xyfnnmnvXVEjWWClyq3lZo6VKHEdk4LgJvWcVm1LDTMIWpCDXJJVGS1dPRkLZbpQ3
oYmhJIYAEicUv3vPdPUjrEbEg/EFvPcouTSjHtqeBylQZbkBeGzEhS0d8ZHzJl7vBFoo6gx8Zy+s
j5OkrQrOT86xxeY0sePj0eT2+Cq83S1EQxqaaWEa25tenNWCppLzKEKS8xon6lkYzVIkkZVoOdYB
VrYjXWvlJx7yTbDIVrY/DFJKMRNRYCJknngE2LRkGjUgUfnBu8UfmazPx05Pub9mHtdbtKPxcoeg
YZa/CCBLb2ODKXvIru6g+F2qmb9i/cfvT2egHBA6u5ORhR4Guac7noTnR+Mq7ZIZOil1UGcutGjV
98o34A/mNS0uS2W3lUFsLemAosmdxn6YgpzbDKJCthl9iH0mHueZE+rolKNsXLyNe28rDBGkccBq
ulqjZsBvtmbM9++AlVAZXRlNaHkEaRmWQ/F38VKSLS7qrkFwWSMR83NIHalC6iEJHjdndlUqT2a7
HYPdAs29J9TnVEqTQH1POz8/aSb2Bz3IcQQYEKnvVcj5ZyDH9TblVlJsbaHDMHE2NruQnMfIlAHQ
oGCfiNcdy9+X2WmMxkUSmqWQm3TdTW6Dq8FnE0KmP1mt4wQdJh4JW5GvMwZ76t4ygCS84asrpntV
nhzwW1Ml+1XrvLTUPdoUyup2YtIFVIzqCBbYVNL6+4k9/TOx+/nmnBK4oz0tFRTWjGt6lobqrepa
1D33WKWQryp/ojGWU8DoW2xSzD/kaMZeH1YIWerahNjwzY5jdg9LBr2LzacuI/zF3V/e3M4rR4cn
/thq57HkYc4i/w0G/JudYkpkNn60t39CNKERN0+u7p76ZRh+nR6gCbFGmCut5IU04YJMb1fMYz2G
zZXLDjNzf075KyUT0H4pBgP3+4k/E54viJdKFOaYTyDv3w6nBsyilinMpUHpXHY5hCuP5r3FqYQF
WnDPzpIxbQ3ISYeslhHXXG+j1r+jDnZJcrRGYV1P7eaydPs7YUVRPWs9ZRzH6mqAlD/D0TpP4ioU
lMtmtUEefsgaqmTegBKsYamni6nSKt5X6TnBPG7JZCkQZ2Jrn01grwP0Y3o0FTRxwrozQ1ZHJr44
BPVTnpxO9HLAQ/Y3iwqT+Hm3bbgmcVFJUmu9VRsjO4iuVTAcasSTT2kfV9UrH3LkMSI6czspkzTt
sSTyWEucsSm1LCfg3Is/KBrkNBYqsg1LiH3onYyKGtX1I4Qt1YZn8J3p9oL3v8DBLwHiQaDVZbGX
fEbNSkG5bvbHRw2STyeJrRVWmlKxpfLOFpuNae0allQD5tPsJnaQUQIBavKLU2yhGoVuOOs4Utc+
dQg3vebtMV3UbvsKNOcIqkhwUP5wtobNUA6q/wy5Knwb8j5s0yYeRQ88z0BHMu4/aPNuXpYgQ3Tu
EbWQ1Hz3fYOa++sMGTmu0GgXkWB9iHJ2bgECIy3/LXbyyuSYhwbrBM/HMeGaD3PJL2FIoVPTontK
IjgaSwcEPG6Pulbkqeafo8d4MNqV0RrZvOVLl3WI3683/idhq1H59JFpXqwW0jgWr3cXkryo273B
JQ34tZSUTakpCfNf7bjJz1Mar5nH5+e3tHFy8eCFI8vmV5pmyDojEvcJdMPQRFoYIQoSZHkelbG6
OfI8WETk3l1hsDbDiBFyppXst1xEEyL6E9TgDTu715RFBO/Kot/yF4UEqUn5gOpHYUJSTu7Uh/ri
txzs9jD9fecCBkgFsly+xR4+Mga2latkQdbjQA3u05OewS5ywjpS+YWOq5afaxYvqQhFA1GoC7ND
1xKC3MBE5dw7+7v6JgC0oa2/1xImPpJKXDZlvv0baUPQPCheRHecu52yfwRPXT2WH0C73QFixgWC
p7FRn0plWPUgA74Y/gs61BAX01z8oUTQLcrbd141+fVr+f77Igcy/HQbMdnIzZKaTAkY+z99sXaX
jj9Mr0OV3nAUQoLNv2UKbALSWOW1NOJnyuieFZ0U8hoeWNRDQ3WtIhVcGxrz8JKec80Rfued2r9q
8Zt5hCYupqW/NL6nPf4s3e908y/Eng3rui76f+EBSKLet+RuDOiL6/PJNH7eHXzO43eVqtH0dpvY
MVh3k6gisAUdlBShbyFrvsUfR77btwXpeaE/m7tJdEBXEBqReoNN17W0cJT1jJfFhwbpUiJRrjEY
wIzG1lVtFHcFtGirZiGTOeRaY+ZsCJaSl58ydOD9tSKpOiYDqm8eZAHLWsWtgbupYkA+II2agyXe
/0qEnWXKvtvDJmw2/oGMqXPTMJOil2RUWb/mhpPpvnPSTohMRBkn9/lrFNabVkPo9tN4YxTVToYP
/j9rE48bZQNRA4dI6zb+sdi8vBuBTOBSZAkm2cbBWLcLTP7STxuer2ODPusXRy7uT77bG4CaoYDx
J/q8hBV47IImACJ25Uzt4mQOupLEWl8kl5IciCn4yLR0wCErGMheQDAw4VyaflPytQI68oGi1dlt
jvCBL0jb/Vn1lsjQb2H84Kl7lAkClOHH4h82HlFW16bxeqTJCtqxinDwoBvmmGjEteXQLlJZSc0W
n2kmIVUHDhRDJ8CeqhS58kni78XsaCP0cLtyofdURO5TJcYUcFLl3f+gnd2WGT2pC65foJy87wBy
Ou/GySTkJ+ouPyvcOMGOJ9YmROeDDKZXxPDTYC9pj0S9pulraiBBaoU+Ln8yIMoffUvTJOYuphcP
AainPFOs215kpBVzGRs49GyIS/r8iGVyRSJy4PllySIEXx1dfETZhOW7uFiC2Sn90sx2Z0IthJJo
akEvBJ8jaSKA+2ufI7+uN4Nr8UkjkxROjeu/k9kBiliS+51W02skMP4yvPuDGPxXJf7OxuwgkvMY
v3VNqffEXkE28svMJQFMvif3Xxc+ll/nl0aWJIfHC62K4wz/F9rWreJ6jhBm5LA3dqwlzTGjz/s4
oq8LVW9VsniEbDU+RIDrs38UZvcfH6lPPPrn4HxcZqLI8Df9yrctn8sB/kkHvSHY8w2kSC9iTs3B
EH37/unEWJu5zwz6CjqdSdR4jjShKOtjPKpdYL0tLHXZ1thXNIcwgNRfVj81eGCYbaxLxI9se487
6NyEnP4wSUUIXPTUXjV6eW0bsizJ/yXnfi0u4Mrom52SubO3FrA21KZs4wK2QUoB2mDvWFPsB1yu
Jan0KnvnJGo+Ek4TNSXlkXxuLAeeMFQKre9o1POk32m0wmgWJNsBiO08P8fyeeK/iizDP/fU4O1h
EGwudiv0ss5yVfKbMfJqE8g0AFWvUKwiTmE7Lt+inoM0If6LRkXqOawktmmHogvOrBWSVr0LLszi
U7xJy9QoHORE5eIr3Fow6FukdVbDgJQYOqqFAmLazECpbRbb+KrRAHWbTKkmaPat8noudKzpfQz/
RYjSS09EXPyCMDsZCkwPIaurNN7GgGSdvWQsx2BknUC5qRUSgq446jX2M72+mqeSxH+xyXCE3Wx+
mbi9KraUTTv4usJRa45aIoZLYr7OOuHzVWCAe+oWxFN1KTc+oKEVGH5IkOZpdcfic+wSnNHVLC03
KagMXGpHnLNr3qPK60uiJJMUeUD0E39DsRCL2PYXHikAd0FGWWHhtFfhYtdrWS0C9k4AtMZrDKIi
yLO+G3jvRiHU4aWHptTQcOHx0/MWAlWXMuysHJjp80hDVwHOyS+ipOG2TRvT1xsle+3tr0zOs30e
tFDcbWB1TGwIaC6zG9t3hFDClQPsuABTIb8nokypGas/iYCrNBsVuO/UFXBRJ0Ad4jynTTKRR8AW
x+PQT6IYrMuBN7QuRp31pcGmi6jrSAGC3iTCRTQ/6QhdbbAoel5DjY8UJWjWfsfYPQ+kwcWy2z6/
5Uq5cC3WouEZGoF8wC8oXyK/jCOozlH2jAiCW58Nudvaax9WA6LSZJRxWe+wQ/FjSoK16HoUF1Lw
xApA10tgV9+seBiRb1oPkpTM68HRDmMNZd+FHivrLaZWkQYJMSZ2AZm6p+W6wxufFRypcrubskD4
xB+/fL0ARpxHqFamdGulsS4tTqXbdESSzzTh3iXPja/lQS8z93beHlyF6hol1R+SXnStoU25hTCu
xpVqN7VNMfQGOM3fBaDCY0KcTrhlYuOGB5QWxVIg/Ywd6E7H8pxCTlaxGyQOYQvpY69Bb0tXTntz
rC3ihlAh3ls2QxZrMyqLC6nPfqNR/7Mi9yyGt4nxibM3Eg8y4qe1MMA6SGQP3ITZFvInwNuPhTp2
OHIaM8QPhKsQTZgm7NZML07LBog49U6RcolKAwO8B3qld4ymuUkuXOCNB9fFAs5DJIdWCWfxVrIH
HNXtsYI8Ukq754Z63S+6Wtny67+DJbkB4woxJYbdkVf0vC8ABpH97q72ss6EYf5ZqcoK2PMN/gR8
ulPi9+STg5e76qpT2ZeFZRlTAFQWaeaTTlvg7XB3pMKz5+Q4IIYwcMd3afIvQeZIh+PxIXw6Uy+r
uUZtvRfNNtUTDfNEwErg8um0goku9ecSlFQklxqNP/kAFZ25uFoyrNVkkKkWkj+ntBZkvztCY3/V
FWq3WojF0SHgF0ZzxfGruRTWhwaaXNccpAQM1HchdSSBVJBq5LFlZKgvsEBHJCpMVuU9vHU3phVQ
aZ7WHF5cekIU7otFwYssV7EfehJJOijuLkMzUDa+fO0/zvx0hV06WysVaycOTaGSk/ecAcPIHJ6z
U2gpAfB86beMANYrSEgrY+1U3F9akW1KBOrDUnbEbRP7XbQXhTD39tYTU7ZvyE4Q0Ja8nKdDauMj
B9BrL9yv6o2M9r374NqHVUVFcpkBOddzzLDeQ60JqzSA6Ppi9LamBOWy34KYi9XPwKTXxKxT0tWr
UNdlvV8mCGaGLQ8u43r08wNuvKC04720O6iObZvyz0JYL6eca9ebZP/xE11BMId3auwCLnW0JswK
/lE+4CIaX/BDvVyAJSBV0f1VvQaPNQKwVtcUoq6qepLz3sANEdmdb5hxZhGk13hHZQX5w2wevlua
PSKca8aoOqpV87DBDEigqUYCY8KWlPXMHNGHZbBZFnSmu4e0X/e6D3vb7zhXitCObDDRS74iL2Ua
s0WH8OhRvAXlRTm+4PE5SqK/U+PXUgw0K5s6IGNe7FYXFeKgmHxKAMcRnYVZu7VJjII4D39DliL+
maMvpiWHtUigVjg8BO4zyGE3Wwwt+zeGrT31hMVeaHQO93/t77z7EGko7UeE+cLGtiYthsNJ81qa
HLmIu+oiVrxVUei14BfUxIJFb/2gT6iJ0RQaR7xMZphvReZ+jpOHtdoVJO4caQgbFLmk2lxk9G/y
Z9H6C21pkzRjlTcwuG9VvQSME/0Xp6XK1u8Vzk6HhCgwBMep4xYE4QDivjNsJIIJfsE+x0xWerxe
waRY4d6wub/liOK6jmFNs9YoJ/ZxQpabo1L7/0mpepeMV7uhaDv3ftcbedZi/FihOSMfbaJc5pJc
/pBpiVXPxDuFLLuoZiSI0qA5hV/ZlXwUuno7T/RBnx5rVzDQo+tgbEr5M4L1kTgYzFQ7dM7zoc6Y
u495jSQOBGcZF5Dk2QqzVTwIy4sPLPHc2Fzw04jPqb5u+nWk/yu5k3K5+xvG38iqiAfeeEP+Yy6w
aI9Yxn7F5i+dM1UTQBVyjpxkigx0CEc2C4tZKF2nUqYk5Dc8YvaPgtRmQYM/rNAXJXqbDcDkUjLF
RGBE7aCQEwCaRi1a9FbzS8iFCdhViQuHA6Do/QZs/IlLZ+javs3dNOteKY59uUZz3UqzfZSoiTPq
jD3D/8oOBZ7rJGQKrlzpqHiWXvwWOAARu9eOCF6DFt49oE0pNjGnjs/xyFw/4AobQjCFMlBcVbvE
8BzUXcA2xC20pHfxX47QXptFgFS2VNPp60hJFfeqIUCoAXj0yjvlIMmDdgs+6WUvfmp+jIbzXQJH
LziXQNep7x3I11Yqv/j7kX2QklkAUMgLu/pmFaLL4bzv4xKLkDIUW23tyTvX6KwVJYZ+bEeiUYaV
Drb5GF5QCBrstqpOI7KnEHssdDX82AAlhyvXWNj3vrrFwPJlV3inB4j4KB+tB+EJjCAeP2TAtIDY
4tUBBIYLDeBnH5r/8t2SC9HLlxF7D4D+slAY92Mb880uQOWBoXeYbi/et7VGCLSV5k5diTGaRLaf
kwMK25usFM7MFQj6D/+ra4SfxlniP7M/6Voypn3FWHrAamwmd/UR0SfrrwxA0kCrHVXcoEX3zLGE
A0pDzNrZ7Yyd4U4lRpIsG2+6Xu4W55JCSyqm0sKSoP3tL48YggKlsK9iCUyKTJdipHHesBAqAcJ1
WFGBTROTn70AQPoALgJOnAszsYgrWBBXNkok4Dxj5Kdcz+2+iBttZ5pdc89yiq4bid1Ku4bWreid
7cxjYlL82PR2BH0NRcFPHigvcx30f5VwbUFkdLnatqOLG6aCRMp1TAnLgLZHeGFHJJ5xyopI+BUc
3/73KHC/Qcnn4oCdZkyyWjt8LXYNRk4y14xQkY+Uc2h3jSkMG1BQjRNvy3wkLigRPOLgmZga9K9F
6qzedaaaTl5qwOT2HkdnMry6QNwc8rAwFTklpGZze90haMlKoqGKf5Lt2bSYeyYKw1wCQyVZNM5E
tRJjKR4ukZCSWm6XJehCQygpIuAmAbaL7fewipjgoEgfsVny7zvy3wNwn0ACjj3OfkAx/hmNtqQB
f6/SLsOErLzxEK+obN5h2qcIHsVVblKCgpD5C6XkXjGx04i+yxItwqQKcElfkguW0XHOFzD6A6Y7
NZYrAdNTYIMSBrZyxGTMWTAzwMj79D+UqoFBWwPIZyNMeb4y2xz3z5ItznCp99c0yDsbxzXktwr+
MwdD3bTZceyuDIV0ODkVuV70zZfQ6k5BFQ+oXzFdJrGJsMEJ8/5MFNx7DmGeD4/MMCzn4waS3ZHf
dWai908KIne4us7jR80PvZKo+q3eNQjPElr91UeLDjh90bGHe66vWx9TmjOTst3kvE62xfWYexkt
6fThvE0lZ5EKtpA+wdKGjKTN5MRpGMYHfvoeGgLqGmpMoYzFBtPXSrxVUrKTblAVOEnPJsGEd2lj
U9Sq3e72jsS76xMzMsleWBzFZlSSmhhTB/7o3sW/mrxtkSZ8CQbn+BJgY8nn5+GzBMmhasicevV6
iI8dusCnGw73M+cGXKHZuRBt+pWp/O/kQ34llL9N8drK72KlFAojYID10x3F/YRv0+i6KB+k3fTl
a/ZTVKb8ZPPMzW7KPLXPPgx4TS8jvSvGQlrZRCiUqlCgYyzMNpvXXWs8HDbIal3Kpu3iyaMC1vl3
FpnMmmRQCtqzHXgHIfgzXgBZuS6ZuFRsybss08dP/iWUKjL6/gT6ipu/Pn8ce4wOfAt+O+QDq+2y
LjdwFqLXp0uGaNTN0W+w1nGAqOgFetcBz9xgD7vslK8IYBP+O9GYhAbdbeolCMheuulxSNx9W317
9EJPCrnUETTIHL+Q3UVPfQv7zz6DNvUgaqfoPYX3XB+lex4oOVsqVxE/1SiHDpF9fdOBQL6rlM/l
+0C/0ExEfSPPbj0hyv3734Is8bFBkEQ3tGzaKXDowY8wnEBw3K8E1YkfgvXUZ8mHK7nga2/ni3hq
/fl/fjwYvThWyzwIci5szNhrtVdLyEwQ8B7AOn5q/qStVB6ZHNMxd4oumGEmp08KJyHf/tSwQspd
1zjBSq9kks7ZsCn4JqWt8hIpPvHzORoy/GZd0awxILJ4lokxUVlyG4B4mKn8n3eWU+sfLIGPO7oE
5kHBn36DQ/Add4a5aZgtAVVCsSmnRtB7wD/iHNdeDTYjiiTOhkJGwhhcdb7WqAES+OCjTCj03ICB
86bszajYsjMFlqHg8jjtJcNOuD0darcj5QaBG674OreCrU4POLA3zzbbGISDI8zk0flboRXXc51g
op58pB9GGjkr5RFEngma2+af8oUd7GiPG64II55p7+xENE7jv234C4jS+qRAe6FEYMeLbIjVa4li
w5JWyGSjbZSyPrgDASsdcqH8yt0YEo02dI2c2sWszZ2eTF9XV1gRWYMyQwVvGEQTKjJ8fif/1qzE
srvYdTvFbnfSqzfLFBgDkNVh4tgAdcNO4qWPAJBk7nXgjmRmXL5CRTyq1W3vHBcfML3uFMbAWB9N
fLMas8dS6+fuyCnZl6V0tWgzbwaFd2CB0q5GxIf66UObkfsBVoQfXZZ64RtXqe5rsjxPo/5XyOhj
6co9/hG3niTJT9IgJ/bB3kqzcZ4Gv+yR2VQOyRjFGseXW/exz4NmhEskh+yCaQY+cJFZZpSJuhEC
YptW9SRvyL0XEge125UTQfh0GtlghmERW+KUIxohgGaROUFJfC+deUP7exQD1uNS3nBIZkNKDO6f
WZmYN2OLJ4eRp36gcdfoSIf6hmWOW2UpbBEUwgAr+mvTRGHOKxf2GOHUfX6sgvLP8vQlsUoN3ysP
jgboHS+Zn9ZZJyWJcOKnpq87xOvhrRFz6Y2dpXqztrf7lmV5BQBdRdGCQIB0lQqclPp/tWWQPL2f
dkwtjv/8aEz5rZqIBeqzR0Nqgv6oX0RR1vqwRpeNS8RHLnRtRaPnUwdaQF+QDnFEFVVqHoEbiehW
724gqMn5sLzAALwWV2EgHUhsfGavqDjwZDWKe/LHzxvotK4VcaElF5vP2EdfBpTVKl5AqzJJDA/U
zBHwfRLPIp/FZfXWnFnZYyoSyDkuTcQ6cp04vYSwMnHbXoobegEknSTu6uWSB/GjJ3cAf9mNsHcW
sBN0z3tpv0QgIua3q93FOzb+wcNW/UOejOY4W9prZKmx4EvfPHINRkBZRj/Ry+mGzspBIPfCfHTN
52pdfAydSelU9PjJx0r3e6xwqmWjZlepn/GENje+4ZibVsS8jUZQAyaZtmTsbAbSc4GQjKmW9B1Z
zQBgVKpbzspaLqeuSl5LPViJizA4b3xVERV3X7u19ilH0iaxGQtbZJRovhSDdxf4a5fFv3SPqHwu
3V/NIcH0m2dx2rIDOJ0OGExD9kpLLwpY6gIS9yW54uoBvBcCvi4yK7tdU4xrY7NJT+0ExkKEDee0
HF7XKsNrUCwJrz4nHNPx+pzLv92enlKnY67TkN2PhZ9iyppf2kJ6oIHtnMQykg8n5sM2BNMdBbIy
+ZUstFt2kaATnI18jPFavaXwUDs2W2Yyd851Elkms/zXX54uxP3I/yLR4WL07USRP6czJkpXAuiq
i4tZ68X7EmFXarJgSANVtRfZai+2LxjryM9hMW6bR40GoGJ49aR7r3zNCKg/uo/d9sFxfL8F6fmB
9ndFBZ9a29xgd+ahcMEMN2r+axAodtgKyOJt/OmVyHyhJyRbMw7desGstZldD0o3pZj7hEZlqbUl
LZ80O8Jor7TCnHik0xfsGCPHKLGBFfS+RYXrU5SgIbHGBE5obtDZp0sbmChOxcBhnNRR6HoCT7oI
GA1k7RP9tFMp151Dw1XGqvG7lVRs/jxg/3ynVW/6nqopg6jPaV8GgZL4+3d+67oHGhrDQS8MFo1O
0idWvLcL9LbQLi0vgX/CxAkJx6tWd8GNdH59szJRjQNOPfaj29EGQ/cOwObscOR/HRcPd6CHdPz1
DjN9XYyjXsKkWgS+nCM4tDPPaIAx5ff/PUS70eZsGWB8/7GnsBs0AaB8vB+YqBv68HLlzWQsMP3P
Ior7us7sV8KUeoVMsrOil+9Ojp6Meif4G+J2RzXEm/0GPrd6+IBPyF/0Zmykwc51ZFs2WNFo3tx0
IVGMXLl5Om8NDFUv+PaVxPTs9jVgSS6hcUvwrblR8Ad+aV8N0Y9yO7DBO8L/kIWXFK3QsENB0gu1
0a4kXnTF/V7VrsbeINmrkM4/Tr9ktFxQpjO1SmvZDxBSsLJXVL9Bl6Tz15o3P4Fulc7ODV3Fg1d9
x9Jr/ApBpe5eLjhaCUUCnXEmnvojCS6BXkYD0xSxA3GksivYJHaG0IC1mqWCBBowiJRmzonbJpd3
bCAquy21SDTb1G18HlgXaQ2om8tvnDrhQYK0znmDZq/8eNeSBkK4EBf68mbaWZhdJz1qoNBpR1Pd
p2AufMw28FN+mH4Z+Es2rHvBVL7w0TCq3HWhoC1g4pUu5m3G+KAKJPSSSf6JGSIfPZUcoepZz0jD
O3XtOsIYf49G6yJ0T1LopiXPya0Bei6LVxH30Iq+NGUyuFVerGyqq11N896e4q18+jr+rMKozUfe
yLuLsFpxmkDz8pXV+vuFXGAz7XJwPhORhTZg+TuMQmBNFSHTSJt+OOCFMNcV9EXVmhHp5M4BontV
FhJ0IKYXT9HjBp6+DXQlnG5tcrjqx0n5qcQJ/v1XIWsKANl76SvmedgkRruFDGpIv9DMo1dqqve3
eD4+BeNmkdt5YDchPolam1GN6v+4DXRmTNs2mHA6tLbOKgUiGob5gl7JKV8O6pmtGlrRHHdbjR7y
Ut+L6WQbrRlIXnknRmnGe6M0S8+rwRtGp0kxWvoLHvvYZF9YSYwineo6lxUvY2elzTIz2dSrANDJ
LRqXCXNn0q+uo6FRd5E+NBkEKQBzzdcf5y5SBv2px0GFdOUeJjbjvHMoY9iQF5ciUR7AA/pkELK+
219TZEXb4sv9tw3Wocz1d1dOawFTu+8WkmtHcT9Wt4yFYHcx/07L1Ici2mxpCizjsQk9lojHwFRI
AtQJe6Zqxfw9/u96ucLwurRvT/Z58J5pTS/2pj4oxTB7Aq0GS+nv55dh+Z/LKAg/4UtnwKs3gJLv
5D7dgarU+8Fbhyg7Wt1T1TiUCAgEJ0JTKKz8tc04d+/hC4aPsT9lc/7uhEuroilk02Dl39vuAg8c
ygjbL6PwNKpFEGty8QXa8I9jR3KoeCp/JZBf0geI+NazDkxxGtpqvZP5o3yuM+HFQg5hNasCgYnn
fVGIuXxI+z1Ym6sOEHuWw2zxnk/3TFV+/EyKwo6qqoe91aNhzMMQh/OC/gkpw3OQWZoRrLf0QtEk
URpxv7GszsBtMNk78dAB3B0dMYqPb3xS0GC7kj2uG6EZGRE1VwFHcLZ0e2I68bW+GJN/ruGkjNg/
pXAwcTz1lkGKf4vmvK7BUc1rML3lDNtOrNSJViyMRD3Ih+VdTo3+C2hinycWC2KrtHeYAGgm1ZSV
1nfbI/v98mM/YG8v/mLN8qFQ0EXn2tIewPn2m5WyQXTDqcXb2w2p/HftTqbghNRxTQJG6jtZsMyH
S4cC5zhrCH1nfNz9i6mok4Y3vjNDzGttj87EpQ5vWLTWTnLy2FasWw2olxBe4Kvu950iqVgpfJFq
moLK1lpe7l8Br6n1MVuEA9ZeY/Mig4GBd64OCk23coYW/cqdrsDVSU9zVpd7QoqpEhP4zMTeEQzF
vGp4QHEVfZFo1jSotuAMHIBTMSmY1FnnPTZ3X9kQ3sDCOgVmToOyVnb9/+MM0ZcUH/WHIHlk4fMO
VMQGayszHqYqe+HTC6aagD/c3Pb0Ef5hl8eLFrYbHzvamhko7TbnZCwDnBTMTUkseE1gpcdgxf3N
vyi8ZCrEuBJtBSN2KVMD8uEJrA/ZahUy0vKywW/WUw1qXQwIhPcSuHcgA92PBc6VESjyotbsgwib
1mhAIwPKF+R3Cq4/Mg4QBAE2wnErj79x6DQ4GF6HjL+2/Y6Tme6Z6BNcGDs2RQjvm8IT+0b1nJOz
AcHkFtsFrE3z9N4T07hAgKttz+ccy69kwBG6cdyo79nYBfSan4/4BJ0OvBouIGGPcL+QVdP7qqsX
ArT88j48srE+AoqZwmOWBPK2xy4cY+Vq7g/whcq2YLCphjApiwq9Hx18Bs655W7RbWA0yEjLy8F+
97xFWFaHRynb5lXHz4zL5yThnPImGY9LM/kVx7S4GHqQhycHZSq22wE+/eMl32p9XEegleo9a9oV
a+BoAtFUorGpos04SLCT7G1kzZeoFcbP0nkl/QyxL3wv6WWSTsDACWqo55Bhea6Oon+yB3wJDHpE
HidyRIYmzAqgt/dnUoOOXLzEDymzn93JFE++o6n8BgmosJwU0EQd2tbDRLU5mtds6bh+0vDgUuL9
xwBzoC1W90BWlro3bXGRCJk9qBZpjs8s3Jh61LK2tdKXcjpLzk8Im2N2iqRc9xGkO1BBaVAHe+K3
hZpY89AlytlKDjWvHD7mLA9H5W7KgqBpi86jqt7u1IiB2+50bcdCq0KgoQlG3Q4C0t8p8371d0B1
40KOF0RZYf+mWamycVvmS/bKJR2MYtFbIGDbCPMc2ek779QDk9BdgamAGFAu47qbEnQdyWGsNIaj
0aQVxEDt0sZz6TyqRiUXb3ApVsvSKMm9SeBhlG+5bxBPorgWKCBqL81aNIP/5192zGNxTijmHyfw
n3a9VOrdTqhM47ix/69+8ayMZyTUz78cOiuxijrffOeePKFrTmyXUBi9S41M9WLUgradzWWwII72
WeFcrtE8n/r4qk43E4isZSOibn/xHwkUcqOMtbq1XXx7ey8TnPElCq+OueSYCZ9mAaCyNuXzCHeY
l11XS2XUhMStydndWO2KRQPizXpLgG+tm/4L3umG1YRYQfAFlhXUBksVgchzNeXOkDLHlUY2ABKw
dDtEr5nIbpJIv9dl1JFsfEjuM8pABjODSlENb9j6kh5chHm0rWSEU60aZ5Tcz4YQTZO6+5lW8Q5v
cR9yse7PH+RNaafQHPSnRHC+aw1ex0IbIEBv8UfyAgOaOCZOMuVzztOzbjY125ewKBBLchCFJ7eq
A3cZwoyfGzmh9C/j612UMvA/SPzNZXmt5g0/nV3rXB1836esIMBxo92SEyyk+GZv5cqIpUiMIqTZ
dxjSHSDNYucBlWCl6jRfTiymIsIG2hE3lepmY63XqwkqidgbjAnvlLl1tfyVmyC5J2XMKd1WNyZx
OFS9UmtigmmjrLg3ErtVaqB1IyF6YWwzu5bMvhYkJ8tKy3VadyzOIQFkMTjYkMi4NIsQpEuqjx2O
cQyFalTgBQiFQBgMKQ19+BKjuksfaZYFMSdMcCpMOj9C9/ehSzyk+fxooOhl80n9NL/cFY42urye
TkDbSjpfGo6yrbIXuW52JePcF8wj1iWVXbiANlXiL5BazIMYBHpHA5aWziv2i2AbxGv66Q+xQ/s6
ZjHU2YoS2ggy5IQ7qNfCfCfx46jMNjozUBsp3XpYtTOkaQjYVt1MHpyYwt/aohE121XLMNwEFu9H
vy0aINr8yn/3M7Qi4lCR9CKe8FOgkMLKq5xAaEypDXLks+J6bO8gdE1aep+8/gaqjkGu9nYuOeBz
lCIEJRYPm24mzry0I5+ogeh8Fo+OgvQ94oF8t+CxbBusWcmPYYBCIu7Lc5rfg8ALg6BYsCFX6TFJ
NZ5eaaY+gdE/M2g2Yg4eS+QiSbhDcgEBi152dKE2v+mTd8nzFiu3OBBdjdab3H6A+yOJN7t4Jexj
iUdcsJmKsQ1Rx+2HAw2p3R9uWwGhuLP+OS2Kj38oBt+7ul/HYQhtr4Ms1/jnwXL1bzz2/NeuYMwZ
fNo+D9ClTiyMlF/GX3VHpNe6IBIh9ei0s5z5DGwd2/ojTvLycYV4pG3xZ1oZfzQQ8uhr4iIzJ30r
ZuV5pQuoHICHER0o89U4TFCz3ioYcaXadDlBp/dnd2tv2+eSwTU9fqoxUlrhTKsgXdeyCpuAj7mm
Y+qtdQWTkAdvlUteB4KIi0d1w0BNENuDQd+m8vHwU0g2PFH2zcBip1y0MejTMjDtzD8O3nOe842t
g76io+MxNkrU+qOx7nmKvQXbapo9YR4ASoQn0sF87pQsoa84NfoBQUYvX/sR7HGjxlaObGvuQHSR
E1Sb7bsiciYliygDutgLbafi135Bn26yQZukd3nR9TiS3NeAW5Dx5jimBnxhBihYAWBMf7l7cq3G
+M3gZPENmrJWwEbEyskMSYQqqit6CmjJO5vWpvBd26lnF22EOTB86q/eW9FZsiQtD3Y+1+HWi6hV
KfHgiSUYwGmYT98RJvWveebRrS1TK1KI6xlk7kxesKfXmaCBR9z3S1cZxduIfOdJiVgpLAg+O2pm
6qub1/Wp4zvLPK8P9ZanviWOTJKbLKWrWelRLUtIczOo0slxYT3QZVAsG7TNHZlXc2b/q2lxkHZ+
C0xq2nucQUraPcAD0CCibpQnIgZFpCmchY3HO4IEWP5ELQcJ88F0mC7n5ajSnSmLfWsuPRX+kDxt
2f1jR6H1p/7yCy+zH5ds9YLzMR9WT93i6KUj7ydON54h2QHEluQpS+lYl0VGhxuFdT/sotvsQuBG
xwiklpsOkHqvYID9N+izudjckmaCFTt2E4hpZB8OpSKh71X9lHro1255igNBEiFozfFJNh6TAH1E
Wn8qkbjA8XC0N+y+Ajsq43XyZhHG92xDe6nykq5SomANJw/LAlxjSv24rbYCOCxBZNw8DM0omNgI
/oznby60HqsIFuj6zNPNba5BMrx7sK5WxEc5eMcvON3KBA21mCxbisrNm210pN7YxO3/hJ1rtHJT
9T70fSFliJfaBDsSp7f9/aXGgf0HGbT6C5BxT0a9GzWl1Wthe0ESwrLOlVwbFueod8LJIpcckWyh
mmEv8nvqKoWkP3P9qXh2MGcuMrOYS7NzGz4CJ3QG7XWs+3yRIh9k5GZcCNs+li8M7k3oL8J/mLjB
TgrcrxpIhl5v0r5crlGaH8lV1O8PGqoOXJ4ncFqo9seHdtluZSLjjV0lRspW7l1mV62fFHG4sM8E
bkEjvWZUaGR9xdhLkDd8gb/+pzqXFFEmw/9N2ZbgNDwCNccZygUjC4E9cAGLrqU3MirLR+/Zq8mZ
P7Y2jEQmIACcZRmaRNQKbmKnPFLUaNySnoLmdyAfL9j+h3VEZ8hpUXK33eFRwcdp2cYL5cnHX1bh
FBG0Itg5O7KFkBKCD8YcTTlOKtdMvJULHuFK5XZC1sPbtn39r6aI4Wj/UigJzW6ZhhvU1q+5EXhW
q67MfgVjQSKYwQWigoARw1BeHdi7caC9SovaNZYzHneqIM40Ba57EQOCo/4CF9Dym4sIt8EOoKeK
uUeYkhUqsozg7U144HDbI9d+MN2kBlHUHt2PJYF0zIUZ0cral+9WM/hmwfu6sf+FVO536YiCboBv
yNCE+mVthAtPZejEGz1q24FbKlCR91DQ32iT3yWNlGIImYgrMBoF0zC7yFOubst0zNpuuMN5Bw8A
+/wCRwljEVtan+L+F/jgBS/OeMlCwX5MR3wwuDB6k/LfJSO4Arx2gtUG6tvLzh18Gt387l1KX6Td
tCbRkieG9/C80MsZj0DbasvDSt7O+O9nBXVTLvKJHxCJfLmdzZy8mHP+zekWSxprjRIhOPfPGD1W
YN99fQLSY7ZjxAXGHn+NrTbeKF7sMU/zoRROnPi68TgVlkf6PFuSTpSRk4VfJeZO+IrhCGUK3QBo
ZItPivCD2gh+TNmI7QWB6qCAhU9ZwCgE2WywdY65J8A95GMMZ9qADg3fhVsqWxAcZINDx/d0M9Di
OdLIw1oDLD+ce3EaWe7X6zIhkQk2vd1dT4ItIVHRR9nFXYmlQ2X4TVN/j70pkoUsQppAIRS/8YHr
96Ch8KeVxpwKtm8Uc29j7wrqjMGnNtmjRnvsJCatvijh1Z3RIetbpNMbUddmgsnn1emKEd4Mf3ng
xZxD9NuQ/zdlWs3N9xqV6nWickS0opXTuwIA5AyHaK4m2oPMSSO/p1FJGTDCy1CxV/oxpyXokktw
P2mTimRONKXl8dVz5AdVup69prp05hmM5eAARvwx6A1toljBcKNHtgJ8IMzF1cOieQaovWu773/z
vxWrL1H2AyGbfU0cAxn5m4+RfitIDKIc2k2Z4FDE9ZC5ELvPiRICm1qIMPLaFFpXlMqmAsb/kXQu
4ZS9vqJ7VS8DYK6gbOdxx2xx5mCTGYnwYaFEc7G63iD+jBy7nu7TMsMXepyWFuWLrnTvvTYAFCCC
FFU6ZCWFeHZYa+0HOfqUPII6aYvI3ow+BNrEvXey4ABzz23tYM7wcdnn4VSnrFrkCj6JsQQ+uSai
ygIzhdtSbgFqih8EvXgoRycO3BEG6s2NOH7cnq7h/gz7H0cdANhuTwWobQ2bZREqvytu5k3QTs1I
gQw6lSP1plmEOhS/wxbOMb89KIgE7YyOi2mi+iIk/mXTqLASxTg/Q1rMR0svGZuLZ/8BqKhgb/0k
+RvyyBhAnrxTsiumXSA5cwiTsTw1MUh9xeutN8zV6ZK5P9u9287X4Uwy0xDy312C4X7SWSRyUvuB
PzgRDnyCA8GGMCtLoTOlGBwKZG+2LOc6h/Rds863j7GCAmBaC06ROKDfQ1f0Gd31J91TKDHkjUM0
7MPvjN38O9bOTPEvRzHwWR4l/SZAliXS3e8wo4Gu08WdHZskGET9+DhckAPkbBldGYqOErm5nxyc
G/jZKs1nGd55VFJXezbscErNQETU25MURUDqokYzxWqBnNMROpoKRRwkInV3TsuN7NMJNkoK1eso
Sy9MAbW98N1b9akFV/svKDOTNPMQngmmi1aO1LC9waVT2Nj2/t6CKs6PNDsMv2TdyXnZ5U0M9OSw
1EtOdUEoNcny2HX2Uzt0jrkcu6DVHTXh7MnXKvowK6WXVZTtwLz8DFVYt6mGIj44o5oxwS2EF/9D
3++JXcDVScUKqteBgos9W6v6Z3dD7eCdjlURKDmPEB+f2hJYpPdfITrm08UpGVp2fnNekdgDWc2l
CIYAhn4pTwlrfI1q44M1UyCrR8W4Y8jiIRlWBU3rA/JXseMuYG8G2/qox6BTpwm3INYgzs3YJY63
njbKgwSvVJJY225eVFs4UjTwht/PMkqxyu5TK/GzIqkNG57jqIIW64/nzSjthHrstY9UJbs4NNIm
vbD7Gb4zdRJ9K9Mxd/jGqQo+hT0UvYgR0LeddTxN/SLb2Vp8gmmH8+RMcM47kl0ddSKoFEhjrGs/
Smws2nw6UI20ccYpSoB/UHWftE9qwC0aHKYLyjadayQjEvuyr7EaQDQG0CLLToz1CzabyVvPN3bO
zk92pxypxBixv3LKBn6nXuXQqVbyE5/J0fKpoQiWU5ZpSxOGEdmQFft0TR0bNvO9yoWP/nWtkG/D
2HXSNDXVd3+FqvaRRY2GRr9r7BxpA4ehE5567Wn3Iuwvb1Dvf/rQnHJNYmd5cmnksgLXKesh5WcT
Zgwpv1NneD0vOXZ9iTpWYLDT3ha/+5LiL2YsnwPesVBDwjK5DXYmS4gJ30UU7coRsjl8Jgvx58eV
hpzjsbox2jiRvEErGkMQnaEd6jfEqswCrFFb0pgqgBhnlopm7R01Mj17Vc+MW7ScRZXxvUYtCOq3
WEyqY5EwrkKuMbX1eoYDTN/J2u1lmP4fvY5raEeLcpbCyDotF4y2zxviIkdn1m5v9Gz5LKajNGxY
tiDcyel2NkijI1eCDkxV+RJnHn06o6qR3RSkaTLBZ6jO6XgHUC9Pbez2Vt47SNR1Q1+oI7A4oujS
PHIS2YvG91m2i1hnLFUgvGYjSdjLALSKx/02fQ1wHzG0B1t3iwsjvpR2I1I5IMPfXUAO3kZjOgOO
i9tJju0d3FV2ECcY3RuYhHpW9l+ucj6YJFFQ8Ro/OdaHKleT0WrgKpvKtnTE37s5vDtQ6b7Uda9A
HrQsu1dofKoQazoVIs852U4pdGOeQilec8c7KRj1XnIqrxpyx/icDC1pt5CINJUCAZejPeim4ZHe
OhEjIzmk1hbu9jl9I6tmpr0NNkFRWPzieSEtN4H278c9o4f/izu9aCRu3/sDfInKT1XvykKPkhsY
dKVBCRGv4/LCLQWZUM3WUadmJbI6/IgJCs7X1ZSZRKLy7MfMPcFO3k6xjUTPPbq1JcQon/JC+OpT
CaxFnkrY7jlLgcgKJY0btx74MoVp/CwxcHQ6DZlFhNI/qaUi3BPzGNamPCvjvBe86jta3yt2ZpsJ
m8f9qFPFwzrl7Jlr5QEpJLUQIER+WN+ZGhbgaKm2fgGMq2KSoblOFAokeEaFYNX8a5PGNst+gZHL
X7GyJMhxlAflJJRwCAZCEch3kw/9+xL4u78GPxutu7vfuJAB7fFB4s5Tv5aCXwB0hbJlW1oRKBwW
jCKR8WII5cyCdC4AqYhzp72dVUP3RXdqoP0qDl4pua3ruzq11Cg//A3skhXwl+saGbPnKxFt8H3g
26iMPYi5qeU1/dxiAK12ZyGTy+nkS6zwWSTUq30vpptQwP+I5opQ+mWQg4OMNBfAVzJojAmS1blm
+DozSUsxByjpXuSYdH9CDNNEANB3+YfHrYQBIFTzKnzZX53v8Jxgms933tplqx36jayQcE9e3Mvr
RL9n6qUMav/SHHexytuQyL3U7RSLWwxSHESyK7Egb5B7P3N1JkUJ2+5zSAu0qtpVeDW6i9166QkK
/tmqDYNkDbA36yZ6ZoDcOlg0j6qFr9KrxcjsImZd3OT5MpaHy/yXBxP68QJjU1odyeTnWf8yvg5F
tXM/dausgwEB4AmMAigOIlb2oW1gclFLIzcJvq4wb1hXtCUZCL2xb8lVVy2yxi1hCQVc1VGeVoIV
iN14inTHE3oJg+dTB1nzHEZBCWvAHBeoOgj6QKwWTITe7JXveMKi36jSYhVEIVF7FUqw/0dtKkfs
sLMFrsuYiF0FjTXbFwFow9DoqFXHYN39lPVd2k7h0d22qtHbmPcyq9NcSjOr1PAjBwk/AuQEUCEa
O6bgbiRAYRpNGm2Dw5LppVdi16rA8MDugtmHJTKGNeHcL84Ujaka4ALIjGWOaMw5CXWYMX0LuK01
PNIbyZYw7EO4q68p8LvT+qS21j2m3tzNnbE4SaSh3U1aKM2WUtCa32YvGHFBBk8icsHrh/Q39B2Z
Bf7yiVuUKINw0tFEc1sgwnNh/8yF/IwA2/2FaR+p1QH3AheRf8HIiy3Ief9m3uNgWuwo6nhBWJuX
Kila4TkGxU1lPJcfPdkAwDottli2QwZeX1XqJ27qtOC/qWoJMZKbCKZ8PmxnJNgAlpfGA0mJ3Szo
MtM47T9I4EdVmqnMsvvwAw5FcFotmEakscR124TZ+/OCMlICV4qlDK5Ft8fkPTL8s18QJKhYzfpO
aqIN+9zUDdyCx2gPLAkPw2qDO+BBdnYtCANUCkLZ1CxufIEGCaht4foKFtAIRyIC9kbW8K6vubKs
rOmBdEKoEc4+6OM9S6nbY1stDtU7ZdIDctjM/Lczuo3nNzAOr5vryjlaQG3PufGLvxqxIiCLVQZr
0NoQYtLmoUb/4XWgU6ztjujRnyW/1wlTznes4YH3udDCDNfOcLLR+XTJ82LfO/RYRVXIItvkmyCM
5yLjZQRFWwKGmGlltFZHi0oZ0oLrLXeC/P4xGWsa2mYjj8tvpXKU8e7YueQkLZtVKd0xtiMTLNgS
dDd3hm9R6f/mGI5yY96o+FyaGVeBL4kUHByLZLDdy7xu9CyfK1I+OKQe781Qdjpx1kTBZe1ZfJzs
ZwH8IoCOvner1c1YtN7Wx9YdxDHSJ8oHLgsPvvBU8OWp3wgn7bQw9CMTjgCW6/nKHtDKVSFsVMP0
B7BjxP9AnMDrkOfJF/CAiooq3NnrFKXQ17mSM9PGFK7LBvNcPZs07nVPDBTfwV0+PjZFben6MWOa
S6RsgS/eAhZM8XHgfNy9UYKzQgVacJt6YVPNYOftBONzIHL71GVMcGLsSA0vP5DKFuV2d2NCNtVg
9ehSWsQX1GhD/r26xmDznVGqKep1UKaE5hjJJTdrHuIiqWfNlzJ/y94ACC42uqYEx/WbMhCUElUM
UrMPNeQqshEBju9W0kP3oA4kBHEaIpBEK+k9tEfBq8Sd/6l87H5eZA+FUGjVIrF8uVNg+HjPrNoY
/qEjRShaULYGuCITHWTpoPH3EgcUMZyNK+sFcbtVcV21xCygfgoYVZkpDQAtYVv41tFJncJ/1zLz
vjxZBYNifugIWN0G647RhZpocnkrS+mOMZIz6tDn7y130LJWn95JWtYFAyhYilEG+BtYKXxaDNOp
/1WMqQWMmWPZJUT3twbLCDcvCokUHR3dCaoF6dfiT7QhGFTHd1rUOx3M8Hh9X9sNKkzpqvOTRZ/F
c3VcnO+qe2/+ze30z1FEFMv74a2VLlSijjcYDzTVP2a1BupAOZMkzMQ7LTvEM151Waj18ElP1XN6
s/5T0SJSJe7XRhPgzLxHOU5mfq+UDH7mqjeTdhaN43m5hnHFjBKSYq71C9dewRxTxPp0ZXWYp9eF
hGXXP8AoMa0oXaE1Jt/m27aRIwfSudVJ6Bbwn+y+pAXx8gfaQZ5fhCJQbtNQsWTsvrPiitl22aQx
69Gpo8zE+TlD549/sc9VfFNvExAO2IB6ebRmPLuPpQfAW5+HDN/8ScLmY+ZfEgfhsX/0lPdh7SDl
SbY2nKXii+zUnPHdRLGTLClQBPbKfoeACj1HUMNH0xvEH/ypu0OyeZs0ejwK+XGttT9tNIi7Weyi
t6tHGtiKK2t/5DH5Q8dLUfoFDIvo5GnZzWhoCduLIZmon39XsdhBvk/oKS+xR2vfSoFxLiEK7JqM
PGdGey7oUqyvPWpx8oq8wW74/d0bPPmuYui+6PEOJoCupXDoCSkajMLPHK+Iktkm6MoS+MyH32nM
tkBfX2UhRK/WTxgRZo/kCaVWSABbYlZixsE2tyLcRVw/qLQ9HCL8dD5z7hrK6Q9GzII4lJifYsiO
IzV0zMNuqv5bc7rssGdmbKqPfaKBN/r0qx2oH/zVWAYvu+F5U5w2UL/qmn5Jvd3ppQrfcNAq5N+9
yCam0pXIg37DWP+3ittNxeQQN3TiMfy7YGLh5My9MzvrmFKvicUsHQv5AiTLk7J6PruT0tXKmJMD
+EgOePdoOFeNYnJnoZFIe0yCWMiLnjLKq5UuNm1+XtgFLVcmDMSJhFZF6i2bWyZu89J2c8vrtQoQ
FonkmupULutL4cTnKbm8RdPCLJtYuHPVquLKGzUTiwFPitIUqfHs/UDNDBMkvY3rV4A47L8kOKyk
0Krdp++PL2zLmQa7TSTpXbXIYN5d2w/CP6zr+jX7wEoTwTFwVGH1NhpBHtYBd8qkUMj2V9rpd271
EKrX9BZECCIlGm5J4xDexypgQorW/hdlG9l6LaE/5suwzB/ASSNFFSp7IiieLMXjiuiFmflKYhLi
cp22Q8S3tB5zBHCrE5yK1PcGCqBfeCcfKu9Cs6PzJXiI3rdrc6gQM1Bon/3/ADm2v9Ew2Gn/co2S
KILi3EqM2N0zTbfQeJQLW/+DQNgb/6hv+3O4Y9unjbYDDtvWhWZKqOHJ+9CECOoOfO9fpPKgNfj6
1fWuaM8ZCBFqbs3DNSHtuDxlhRiNs/+veYiPyN22H9ERewE/wq4+L89nHIbIrURYFq3wUbunh/4p
a+HQMwqJKqj3awVvMwtHNuPq+cjbEaW9MMx3SBjPAWzqRbpfaPzu8Z6451FNPwg+N2tX5RLeZiq5
PUpzMy//lhnDUX+ncQ2z29gSab0fxPvr77yVYtPqB3nJLImn8OCe6joCE9IQw7F8AgZpSiLn1GBK
aAHcO71lyCEomoyvv7fqKkTmXc3Jkv0UcPi5zCYwCRMIFIIEl4FmlGxasR+RVDEBAJZFBduLBIzY
0cBElLc6jXKXjoWIE83QH4zgh1Zej7+Rr/11yeTEb99mzkqMWVNW0ppsB9aWjXLsjhayObvQbqU8
GSx1VgHea+TnHSWiGEXgTKeftg2DaGYAf+OlefZj5JMCEANVYdDLwK3PnwwNYzmxQJv2dMKEx93f
0k/KiBvKehzbNoH0RrJ3R4ngVoigqhg6goPzguq0CrkeEuJ8qwJD9lCQsyOPgB+oaW9A3C3th73v
9D5M9jCvKdgSPp24ls60B7oMedPlljK14F4/GWMlpOsXBsipn9o09ERm7822Be0stdGMfg+vQ+Qb
nLc+fGM3qhLsbmoPoXAUkWVRrh3XU6dsD/HFyfgmE5A/8yjToWi6026ddVOM2n4DKqv+t7SHybpw
Hf+CAMlb3tSpPO9cVK0sBjElo2+OZM9hY01Ludy33ZeW7KWSIcIDEjoTTth1Iw6SPkm6YkTeFzX3
D+SjpV9hn+YgtSi1voAnePUhYOkC5d3/tXjoZGDg9LG20csnukR4t0MftG21d6hGuRpZw4FgNRe/
vy+OJzvLwODoFnUNvjGjKeVmQW5MNgK/ZS+0cuybtKU2PiezNeTHBWsDnMCHlugpM8N3KG/m5YyD
rH1G4ftLVuJyqNBJKNhxJ5FAge/FCphWVms+q2/wIw+y1bmuP1SPnM6jGstZX0IbFYHO8PW0rq/D
Vc+L2+Oy0HxrNQ1UskOViwnCohZYOUt1PXNQsFImlP1YcO1in5ujcRpArAjhQhqK3JTBVM+kmbgA
6Hh3rSMzkGgJ8MfCrCdPY4bkQIgSC7AFjOGk4AADgzAYKCN3gDhGoMYS5Q34ZeCbKiaYAkZG0FDs
X/Hm1Rg9CWaH06ERvx9bzUBA2oGnW68VgyI6+zM4MheewyUkVEH86obG5Im+J/6CvZPIR5sfMQc4
lUG5GkfDAp5YsSw/scY7XWku1Ah7SimGxzg8eGjYu2NUk8333TQL+3NdIoa0B9nLD0p40xWge+zz
59AKzgNbzrOag6J9Livhw9cC3v2RbOGW0r5PAxIFq53h0VgZytv/VuIQhCitFzVlC20mCLHMxA/t
OOM3JF+tR/jHNgXlV1ntODqmuEB+zIsF8oDNOwIBawBDJTxHQkfa/8ynF9w+y/y+zImusPBCwT22
w0EselISSeh0ReWzr1jtjb53OdvyqrdbJVON5MWRIHQbDT190hQnFXD5Euurs/dNY174sFvsB+zH
W6zSXJbc0RT+IEehEfAMAb/s3lP5wuSPxifNw+63WLmyXDR757Zznsxy3PgNGXJNW1Q7GrnLiszq
CG8VQN7H3HYAS3M54HKU1jvJG/HOL18f6NKjMnhMUqVVsXXyahz+FyuBuJnimsK4xUlAWOf4GAn/
cDSRcXK47gW6H9XzQ9naMFEI2IReXgpxO3E21A9MN47ogtKknWoOh0V74RqcRtGuXzNcSMTQUBLH
nQ4mDfNedikDazM30lCM70trdJ7xQ/tgVirCjmomCvrW1ajgELI2fw3E8tbSWoJ2aJOOLMftCIkr
9dbIpXroYRDMMUIoDDQLrlvRNlMj3qs5UV2169Ljyff4fg4EIXin1H5rjdFIc8gh2lsDNWMyeGSu
WXw7OkXOItvHgo+EEX1GVwq0AUCSdwTmbJ6SHTbRgWMZliJwYbvwON7JfAyhUE97V+WqfCIwQPP/
Stq2Ay1U6xLhNgmXyQOCEgO0ECES+NTx0NuDeGFNyAjHQy3J9PnSVKQMZkF/H+84HSAP4l4ptPyN
87FJjSKGVcSn6YUnL719P+w/FPfVzIQp7oD10S/xZy9G5hnnNfU4WXF1pEZ2dI9clMXN3XjM9F4L
em+czoNNMhMVBnhKUTup51e1BoUva9okcw47pcIM48JwNhQeqBEJxb+Bl/CaFDtA5vQ0kPvb/BIO
DwlzlsvFrJVPNmPwWX9rzjYsGgKozhJ8Y0Lq1MGdHypZTy1RVmXPPHKKOAa9SDFFlKYlXil+5OTg
gMwOWNhDOv5Srn9jmCyiuOeeZ2kAuNp5yavjQNyPst0ZLX4RonKfTLCo8GRV6zk9lab02CsKVFpP
Qa/9nk6tOeDZizr1UsBejObSNasgSAsjDpmENnnyKQCWRhfbsuSGrdCrxEFbSbGiuWPo+NoVyyQH
Gxrhvw+I8n9zM2eU0I02bTvTNGcESrjXe8zzDcgywCwvz41UqntoinIa0mswqxWGfLPA7Ut4kDbb
CsrWDgsWhZzphTzmZedmI9G2b0CBc2CQg6X3mANeelWqUqqZgH+95b0TZkUe7sbjqenbl3w6C0CJ
Yow/auVrdT/mkSUl1dqwRcfttpBTzQ2LvUM2MeY3/qwkc//+DKSkGCX1XFShQYX9YP+/YwaHWsre
VCpXB9dDIYbjR5bIkfhmLU+yYIUxDM+puG5AOr7/dpzcknIGKyCGYP71Xz6qVnmtnkJpF1MJdq/z
GQufGL+4qKnKUVXADvEQy0lVemMwQJ8rvrHSTgLOm4g0MliJ9wCF1DmhXc2qzp8KU5CBwwQ192kz
d3vChwtgAon97Qaxff/EbjyuyKNP8V12vxPDY/x+RhKN/l+DkwhBFOVbWzmpHTok5a6NFUL2rhUF
qt9yQGMZAebbKcRQbSWU2HHVsJSNJtVreq6sTumWDl71AsdhIJmYTn0gXGFiN6/VRRGKofQVXmc6
uPanTTLuJWxTes4r2+kmuTdxc/hAmvZ9Cf5YjdTkUqZ2OUiaqBBbuWmDDFZzWzyxY8ZxEFaFaWs9
R/10rR8WVNbWVTknYTZ82+FApJCIMOg/O/RxXUQkQXDaaxXPx8NbuorbkKAjFaDaiPpK7jUb1lXt
zozVtakUnmunc98n88FX9CWKd4xnnqucEXTBCdm+6h1JoZbu+l36AVemk5FjoJfTjsy6IHQnIMae
71mhuymtUIyBFzFq0GUZ7X1KobpN595VCeJQztgk5BOeUDiZVFfuvz8Bc/0O3HM0g8mhOprWnr2f
1YhyBXRAM4w7V9fOA3VYhLNKcL0PB491aHpl+4ECA22zPCyR30Bn3x3pyMA+uchh7oAB9toZY4Yd
qISO4TYlv08UaIKYxm8C3r3D6XUU3y7y3QSEP9RsgaJgunQYs9+csTBu2d7//+cbhwTRrWwJcyle
13e0/8RVpEsrtxrm/PVnzHB3QBn2Ee+kkg3SVJloUBE1+0iwk428E6hzZ93xrGQ2B7ysbhZ1tV/U
ZTTKKH+mqIXmvY0yKt/U/xW6Q38lFsLNqQKSAePkZlHpsBx2d6JMz0mLU4Z86klcA2mibt3RBO8Z
zzCMVvU+k+fODQEENmEfDCyt8vW+97yzjPCNhrS7cedFOyrwPXqgEIfavwTbvIv/Bf9atQ9nI8Lk
l/OGu++CadxK8SLmsr0pLi/lhzRSIXFErG+6Az1UsbCP8T2mC8PP7LjkYHczrizjZaXmnLF1cEYd
9ErZrYmkX7uilVZBmdeCYLowXCs9O1Bcp9Flry5TWt93ClLW/sbqlYLyLWX9Yayy5A4FlogsMdqf
mViQnTF7h80PoLeO9WY/oyOmmnkRmcIKJpbxLB+0HOdtTrVvp/MmrHOW8itB523TW9lyFibDZwZn
YaBp1QVXTVLpALfaBQF+fILb+p1sRcM2+BJ0SSaaFfMDLHh7foucwwyycesOwHvk3ScZDKLnOmqe
fYpehAqMlMplIsiZ7SmJF7gE9anon34BHbATRgOd/XJEYp6Tv+SSe7yXo/h7i2V1L3TXwqOAW23q
LbpYqPkwMiqUqt/JCVB1dBWvrnIgPZwfD6BjsW7myxu6LgK3i42WPg4TqDaxwlKZ4u/FD3yg+NRj
e1ZkdS/w5hnIGqBFaw1XtBfrVrYRUbwZHTo53L0XIXxkz/Y6pSWvwOhmrCLRz+NTHLCTThSCJwpe
/JhkN8dysdprUThglayOraUhErU4vSi+rDNqCSgOSvIuDmbDvePooqdnBdjUMuGLy7DxGNjV+n6/
7TEwX7N4V6a8vZC/dYNNDuF9bIe6mwH/TiPcRxpCMNAviPMF2rYo5Eq6t4CvabnaqtRsuWHQXzZK
7tgtci7qNWaugjgh0gaXfMpDF3LFn9PJwkCmwHkKNb3Rw+b1w6WvFB72wKusF5/zEUuSfMXWqqsL
pE9Ac88sMA2F0tt30VclTuznDnF+Yv/3KWzui8Qr1lhSWmlDxEZUP6mtEH/3FucO6NHSnZ9/xo81
DoucoH+L8A9dFT/5CVs4B8nxjLTNkoMyWWjBco14/hiUUhDosMIMrbL9f6nt9thdje4nINBOGuLJ
z58eii+9MBIEfwjEMYM8eO4HxM2Z5+npqclbnWvCe7La0aozBy51nwNu8PsNufokfMLc5ojhywPZ
FeDF6gtqt2AWFUV8vpaXlee2HhUBbYj3a40YDtgzlvPzae0XanZ93FBdQW8qSzem/Ar5P24gRoFO
9b1Ak7RMtXslx4KblS+4C6LlWRB5z612v45n+EETeWV28CYgInlFeXo6RAkvOdZM2fOgnwti0jdo
NafT2uzCe/N6yd83Sdx79AgFco5MCYIoM8sBMKkGzvfXR7Si+ALEv5JDBOJY6xSUza2AWzehZ6i/
O9Lmat9ZkbTlfhRGWuRDYq1bjbszCpDS6z2bEMgDjNmsJePIr7GKgF9fQBUSK1Fw1nkRa4z3w3tT
4XMqEL/Go8rfnqrbe8tM48XkVuz79UBB71ee7ri+BVxj/R852WtD+kAywtWnjaxWMbRjVhhQMpkw
QEbQSv6ZtcWEOb19gPgHkt6HXqQfbIOB2STlO9YP+leG7gnvtOt3FWdXSy3QtOLbMOK4uoJqrxoH
7f3PjQIDxUbwsSLedaiYWMpc3leN7NjwmUco8wSciNPngIjBTXX/xHaWRf9JQyOIsOgfK7jGL9/T
lKE/gZhStao6Btwjn14M7JT21ZRYc2uxjALzavKpE5W74peW/yhkrZQODx3pvds4YzC4UszfiLNN
O+6V0BGpMer3sdBFjS99k32DLWvIGuWsU1SQqC/KEXUPpmCjqsNiX6+Ja0zf5LNrC1pbUPSZOUJy
eD2slKAg9OsMOrUHyY01ipWW8XTYngxlkGHwbSbxzrVGF9oWODTN81w34RTJUwCKljRqkUJLM26D
UIIpCJSeBj/hcaHNfFq6t11D1qD5nb+EUvt2D4IdzYwh8gWJTwS29XBDNmxSLDgga9c/N/UPSOH8
dQ3A+GKrAB9Zy9sVUzrXJ57HWQfGr6xhyi4LaDw0eU+jrAUxxG/rgR0y+nkzhJc56MAfoMtYz7lw
HaHtT5j4kg5rKSyiIw3JEPWax9xa1tTTYWv8qZb6MhEUu4DnARbCJcWyG+ie/WkVLd3vetLNpeGz
n5g1c8nJupyrKOOnFPJqHmwT0Jy3P8CHIOL+YVQPWr64Xb4xkhrxE2l11e1yLOdf5r14XoeD1yWE
D2zffA7xOr41jNj1KAkrflwHGP/ebur2dJEC6lYU5xMUBZ+pTWwZ59lmNrkZUELprmeJcqnNgrMn
GFeqAOhV7OavWUc25qTibU+JEfo1u9aMjERcQG4yqmGZy+e4M8V+ReDpEhStCUlR0ODLaZVi77dV
eO6N1y0f49wdGan+Zk37qZZlCGsPfRPfxrKDwFcBVWQlLXbzQtlaJJKBQOzGIVOTr5XcV5rui1dX
3VgkVkcAtfKA6dzpE8LRhVf8FSgOIqgJhyNQlo+lUj3OHpwOMYB6JS1tXz4yi/87LNHU8ZwDIfBV
0tGI+SamJo1VFs6NE2oej+4yWQn+1B5vcJ3nI8T/NQ4W4owZTvjwDOzr9j4XATlrvHyjCN94vwb7
ec1RXWo1qUVaIi120oDdNdU2yXQuF9eK98edUBhJbo+W3Iuzb1ycj/6zYCzMvrqD+jlkXUxFVc3h
2PtAIH/6dO99V8n09J6ExJc6K9Ahb1A0M1d5ghO9IBtJIWCCRYJVbiA8utooVUTiOfvlX1HjFQLt
jvu5HNzF8EGhAV7K6rhPfhfWZmKrwiVHeC5PYJh3dMFq+YHoIhI9H0PP2BipYS+cs0+owG2I+Jkb
Myav/pZDmchdJjpZSlf5L9Q+H1Ro1tFLeTblpHPChwnuBWq3RX6nnN5qDnshENpRbudL6oDjcH0W
ZyfwMiSAipLQ7iIA2Z/ShsrEhlDd/rMBPKLYKyCywK7/BPsM8KxmvFOed6UQFSdQkF39g5w1UAAW
ZMgK5nWl5nl9BWQ/fzUnJUmzZxG86DfNubzzLPhYr/q+axoJhw830T2Kc6hte6pkgou2MwtkuAIq
+ReqCSC48FHGAUfTn08uDV2OxU0eIV/w2Y8VW0O70IIh9BzDm0aeRHwNip5CY4qo67I3FhnKrXFK
2c2Kdz3v0t+52M0x73acfinZ2hs3J79/0BsQCNpuiZTOgMZq9AKJaI1jJeBa3XNLcRKNtyU6nwje
wozw7kiMTiYGaA6mYuY25VAzOPnjAQITN5R5ONOanSJgbxvmSpuYyVcuAOPPO2FyEZk3Sxgcp5OW
azAw09ljdvbAm4LDCRFkhcWIsGt9CHwKzA6mV41YPFMaDmG9mDdOXWF87DEkcSsn2uHAdC5DleQX
1JRppcSzbHmMnu7j5XXwETKa++55n5t7YNo0T0+CoS7qM+TXRDoXCtDJVqItF9RamncoNXUiQ1KL
Yd05dx0Df8g6+X785oHsWNO8wX3VpzLgP/DPz7HyodmphXF9gQiJdGIbSXUXaepeaFk732gb5DSi
KofW7DB5HDGM1+rsFL1+wulsOdh8v3zwoqlwa9d1fw6TF8RdIDQ+65DPIdKefYMXPwUBP02XFaqn
WwIWMKm6yl/ZP/ljUpNn8ALDvWlpq1+59CCPg8fw177YuUOh83Kg2S+wTzIZnfLWwwR2gxcVhU0v
aIK/GU18fK7H89GXeymdrjKWJMSLNOmJ6U4dbC/fOLmUy2xFOBVaZqtGEV0mc2fQhoi4CoP5MUj+
J5+k5NC7cRUo08ZZGH4dNVGOzrz+yhrnbDh523lf65AvbBdLUw6rWj1QIO8AiGJP9rp2bAx8WzW9
4+PV6Hf8Oe+cpG68ILdk58O/10DpTZQbDpnBp9eltuMz+2nqUJAIvjM7C+q+s+w5GrUh9eoxtrWl
RE+42UyrwHZt2018TwMCT1VtYaMg2mJF9AHWlGhrA4OVVJSeiYkLUQJI5VQPM9uHsM4ioC2F3oIV
/ab6h1th9EIUzqHx/fEnhOseE//RPmuKLW3ZqH9GCTPd0RHe0GzhKUmVH+JPNs+5JXcvwCw+UJEi
9aECmyeGRv3lBLCNQ+VGWkFneztxTQetVbFdebAkAOLILK2IWwzKQJ0OOiyqAhWsF1J2K3t8q5a+
X+oXZeWGmdS62rGv8o0q9YLMR8lEj3BlGSnUDciKfOXvgaxQ4m8fc1YPWSMhiwK+OlC0DhSFp2L6
gVnePwbzWlyrHc1mBIuSHfx0iXq4d8BSPd75DdYcvKdkihkGD6xJN8XDzMw6sdm6BaRTdsd5tCcZ
CiO4jJP1BsM2MjHSCRbUQe5qwvjNDQ8bvXdUBVf5eztsQGP9aKaPvZIZi+63tN7hNoCKK3dSaNfd
8mLIfRDJnHVTKS3md7INvOB9p3lUJj68uzBaLp34pP8SwU8FTJAm/S2n22n3+UGDM414r8mtvkNO
x7xbk+j2va1PjMibLMlfiCAYJYL7nX2MEExpSiTF1say8oTMO3bIUDT7G+Dn9Pm4X6/Ahd4eL8gf
9Oy1pBt8MnK6cJfkvxRvKtmRqxfvBprl/liuqL5QfIL2G7+ytj98MF7fUijaMJAgFaRHocqzIteb
VbQTD3k3PqxFR/TliPsE7LlbDO/+29KFgtSbqMcDvYWr6+OSTYSDQU3C6GUXN65VZ7zGk7L67bvN
6jMZQCqEsOF7FM+QMp+oijfaTr1Ix5kZW3l1X4EyZlx0fJcvYU57WftkxRYhV8e8oSmwYgZohFsH
ejEf+nWR+Rfv8B/4J+JDs2J9VSjUKOBMmIEMm4CApXx4707Ucz9gRUdowzyGshZf16rWt3+rQQjU
ujiRNJRDdzmbAmeRD651EFzuIx0+lCsZ2p5mtBp0te+MmHN/FVW71O+Eqzos2ebcIRa2HmFfK3s4
FlIioPHiT+gwWciM54U0944MTxddCrXC/BDROuRHcOKHndhHvdcFqbhB8/gj9Bi1gj2vgPi8i34m
zNouNVv3wryEXHYkMFFw7TV17Ewmb0oTaRDxUkjcDwRw2YjFq6iZvtY+qbVVBCQM27fHW6hzuu9q
tusfF0leL5BtJVwl3LsChfvtYTRB7etvw4FvDZAM8k8ivMyPBpJxjobqIT+S1TpPAX+5mnGyXrkI
lB0WILrg8nh4VJ6TznbW6zqw2jLEFecKa/LJ7fpLHhZTXIK5Lv9U1CLHIUMEZfy1Oq5hyaRVfiml
TTKigQQwGJ0+TxQRbtUN8MWINgcc6b/x5wqgO0l/YSQ0MZdqI5EUVihTu0BBKfoPVCdxuG+y1lAw
lWjzb33I9hAujpHfnyBxph3BR5e6oJ7taZBOc81gfN46zfEkaMeHqqhcoogyj7Fi+RYd5l4y4RWl
MmM6183YdCpSNeyqKeFAhBiAlaUu5X7GPP1yPQGe9yeQO/7d8cblkI12tPdMs7kxuk8ybmlK14vI
jzzTF2XvTeJJGTPO9j4ba86JShQPHewW+nC6Q29Brcr+RHLqj0nkwLdOxoHiVA0Dze6sBwnoFlcl
5IGih/BS27MQuE2y+fPSB51Hz3+zoOGoujvrqcsff+eo5WlIjZ6WlxBwG6ZqCyow7c/R0pC8T85g
ARevsVFCYlsh0yl6zQCvy0vAMTUUL3o06froIxakSsdK/qB7iFtE4VYA5+ktMRqVLgaPqX5rh3+5
KdFWa6+lV5o61PJ9KErgJnoeUjdoS2FyXDeVG2RGkP6PoEKQq/E8vFvBIFa9mVdHVcdq4spNtZ1J
buoDfl2Zg2BmbitzyeSiVbf8G3QwuZSZVeH+mGsZN6pEcWC2E/USBVfrmqTpmFiiFeV5MtUAEUqf
W+K5Zm76PyazqgpnsbMPJMnyQ9/GmWriT03yp8F/1ekf2pVc2I3x4CBBuG1mmUnTPQGOrk9CHIgY
Iw3OugDYDx2JnnVCuaNPp8aLDiLaJ+mNjSSpbYpVAbw4N10VLDS7n6gHwplr1c6q3azLRebkyhOW
LONlaDza+PiQKWsjC8Un2E4f1TtF3D9UMrYL5yhNYhm1vjMzTVGSjSnmkz0DXM6/NtanBbqEe7Yf
YBz4AwATqBPDRJX+1Qk2yub+iJEaK5mK7fiJ0crdjd/R3J3mLt8rHObK5RgE5y6tcm4NhNrdWwfb
fuO8Yyt2oa/SVZ+yWt50CIRruSLmViS3jrHo01Lkmzc3YpkvsI+N2dO2VrsPP3lPwJfIpoPLac5X
chVkNxYF3cr12eyeM3RK/NzpLwsv8DrZvflior0o3kLXPemGE7WRC89gaUl7DqtBm0oFfQ4bMs3N
fKt3dyqXWpAMzWPzP1d2PRln6xMyK+xh/Ec2MjMBM9rDnQNgspiBsh9ukRk3I4mPjZ/uipzbo1tV
YB57Ca7vj8VNEpG7aHedGx6kfoGdqEZltIazgFZjvoBujjcy665ZV4mkKahko+swYrHjVNXQXjrD
WEzNPs2p+y34em7gU0V0GVpHpewvNoS7N4pElfZTI9uVZ94/GFNMBrovEN+b4kT5ApsFR3fquzAM
IW88bH238quupnOZi4MHcPsqIIxXbPjX7bkQ/ey5+G8rkdeFNqQtkSCpZkp1MKEt7SPrAxw+GU+I
1rDEBNGdRq4r5YNJNkGclGAkTIGJj3jLbyKYlIG86WY1r9aInRLLnSo08BQ61DdIQ7p0VGwEzF1V
McVO34seHLxNQps/EpxOCoBtNQqiqs8zOCRdYvkugaJqnB5bT3at/wqtPQ/VSptYSHktOM9MgWke
SVi4TgXrH17lqP785aZQfMa6pHeHgh2ohtI2dTogYgOF2uM7C9zD2sZhZMyhxXZyh2LKObdsZHD+
SxzJTkmzbCImznOE8hlmmKiGujH4MLh8OgFp2ZJqNUoLJ02HflsMkdB9DcwjnmSsuRFe6UT8iEhh
rC7KHaf8Bw5/MTB//OncLxUzG9eoXZbjQyfhEnm8AU1o3i73u8Sc0oOY+b1ySx+vd1rsamTf+Uwv
HmwHGxK4wg7TAhHepWhIS1DoFtdXMr7lAc8KkOJkSilItjw9jXUqlraEfOBNaiQWh6gqOc+VsBCs
VEuQ+4aj0oHXry3iRrPve7y/rfxg3cjvwEfBJMmnLtwJGCuxIhWNeYaJJqEyig1oLfFfYsWlKVCF
Z4YU4Ztse0W/FYUsZ3UZSvqaAMMsClhqDw9cdQlTzn6v55cvxUAIbylW98hZQRNQvO64g3YmHtjQ
uqTfI8Hl7CilamBu4vG8pnMm9XwIDN8lrmyhPjlWumNoTw3NbhTrX+DDgGFfyEIWEoX8F/3NmylX
Dq+9K7krn8UIAhq74RTyQgBEf0BJOko0DXMCZf85N3w577Tq5x2sTshu/5t1xbqLDSSNgY8q0c4M
1lE6K2Cdb6IDCPAUHMUDRA3v2uMjBuhrR/VhL2DI415tPzvwmjCjRSDl7S9cDc6OetYDp1lnNMh+
HsGq69/XboDsVf0665C4KyzSo9MzfJhn0+DyNCdMD5aSR9jwnZBsGHLaYMKh5L+Bg3bgLJ3Bqvkp
nsxwVNFczkmqk8rAN/2loaHo78D/bOXeSkQAxXbEPrw6xv+mkdqRwe6pXuQRSu/xJLYY3tW7p9EN
WAGH5taTtoNqbmiaE/U70FjjiS7S8J9XPrbkNgNYU0MtWnqOaTVGx39Czn4L0gMIdl18ROlLMglp
I+7020M3vX+6GRjQGCc/VT29RglJxUgH9Y6gLWsfhlv/4p/raLM/03z3465xJcFK3k+lS5G+9xYN
643xI5+yJAYoAu8sbCQ7Ep3p5gj/I4x+8Q24DcwUDXqeFqKJ+l9eyuRzarIpwLcgAR6eIIl/W7yx
dpqK3d5FhX8aXbivv+f1VQXOHrdQffm0ZIrzuVI4F8o1+IRUf9q8KuB0r3n+kbFH4ijRfg4AEMaM
es7CLVpWM3HBNnD2XC5wMjkjJVrG/h/xp2Ah/aZ0NHMFVlSDjsa32W9zDmy9dk//Ubu0CvWNn+FP
5FFp/tIB1Ug4djqUOaQgcpNZQUe2LWyL4heldFOHNoKcqO7+Et+OE6ocYs95yoKrc2sEa8Vdm+fn
1J8uJnu06SYXEWEhX8BOJeZlcMR89wL7SYfoEv6RWv2y8LvTkVGfrvA8kHnb6A4eBu/GvYe4f7gv
TqNTGofghE9oel21/Fq6Eih0YzZQvZNBFb+o3Aa9rssqLo6QvNYU9//+MA9DahWICFW5svUh6HPq
idaY5Wb7hEiDbqijaoFf2iRb9NJTKOn68avQlmcx9wDRYe/Qp8kX2f73Q5GFqIOyTxkv80hYeUd2
KfEH5BCysIIkb2AzZYcayu9VAZIUW/KSp2rRq58neKpAIGDKIFb+ei4g4tioRnlzkXPCwPLOa5PO
HPeYF7pEZ7M8htCFqIpOqwRgI4GMAAv5k29+uQU99CRXCisoypiBAejZwvJAo/cokJs0Y5K21nL6
iH2r5k4Ui4YpXm02pOQ3gj0+1dNAaSn4dYvNvX8e0mvXkKzIvgnGSNORgrl5ONTQd56rroK80kvX
SGNRmSMV7bQxqxf8PLGXBYSfkq2AEUswMzEJ+VkqwJfmFf2OAj5h3LtapcKkrck5N20corzs0h51
F2XJGfA8o2sSYmoopr+XCK6aaCsyfoyA051n3uyEg1JJkNfkVR0wF4vpOCKrbPrN7/3KX1jUPcRf
L0Gie6hNbS3bbeU5jXe39Zre35F77bnRwPEglCntqzj6pvoXLy0HhvZpSYTlXwqaeBKgDcvLVIzk
u1el8mJAbHZQ3KkDtnWNGpmYeMD+893bjwr5XuRvKny1KJPopPbyBU2kvLnZ3xqV5GYsu4x6meUp
gMOJxcBHnQOPSX9EdmMFKDmHJnlPGTd7Kq1JLkgjVFbqhCiGtjLSPG5lhk70IimeSZEHJR4ZF9vl
QwHvblNc52WaIj5cqRxb7p5XkREFVVon6/E/Pp/7ZFOAt4PVOlW5vF5wlVWVhomq9bxSgBOPZkvq
BTgpAUpcXujGnDedas0P8pZsL1qRoPpeGytJl+/B09eyZGsM3HHnFHgIpxUNlT5wDk7VobEPgInY
cpBWVkXnto1YHh2j6wsQFf/Uz2aHhqGBspCdxzPmW8B03w/A71VlnRCI10Z7Ceb4l9vDMOjmZtoq
EoAj27zflq+9VgP+OjUKhv74cSNGgttF5bT0FMMTLY37BLnkxjOxxajpl27WQW7/eGy+2WlFOJ/W
mo3r8QMqERLz5i1yLizSLBu9WMzemjjvdbL9xXVpSYcUtbGnOT4ks+TSk9Tz39SPQ+MvP583ucOd
B9K7VMTwuDWBX5Mi+v54zfWpTBVj0I5tAv2w0gUcHYqioykAFntRgU7sVT6Ga2/YdIWxw2Enx3zY
OMsLmHtoSI2m3tVTFN8r/n6jjoIU5jmvBIf4hI4n2LnRMj8nrDlQnYHk4+XaOLNRcUcROnVGobQM
JeH7lEX1moNBcK/ld71R8YXdQAQ7bEAYYQZ7w8durSgQDcLS7VJ5CkidgniLVn4yMh1MLfO7v/IN
1J/3kLD6SnjTIfh1jozUnTFfEGuLtahNf69Bz8n+gZtnq3qdryMKwT0YsYJs2J7hNzfPEfrnd1a/
MtSc+2QszuZRkwZhywj57Yb/KZpvGjpRxF2/qdYmbixKukwU9H6XqiWkmjPhpdefWBJMpPizqP2b
Bh3US8SzPiQsMMh7zoqaQTw3vJyfC44hRymDc47lhK3C4RQIms4j03oqI/rwRyDCBW57dyWgrfxR
bI4erL1V3Jce4mpc+1cmfwB8M7vakeniJw5/hWzcrOW3k6OfRJ0jb9fGuVapW09bLfcC6M/o3Ku3
DfdlCfazXZyzQFDKhRtOsSXEcbd0QKjCU4zE1IVeZbcuOVRUWMWCRJLBSyvZw3Jl4LtFh8LwxQEb
1uUHgURLKNZ7j2GC0IDDwvTovQVWH34bOn3CJY3AcHHtV94mwfKF/zddpv4p0LFnxZxvnd+WnABq
HlDWJuPXC/YOjdRNKfNkGu/fUp+BR2WhI8qvneciaTa7jrKVtqrEFwTKeiSd2yF6Hmzxpcsmp1a8
/s4l362+LfG4mfNhBaJOiijmmsiAgDHVd9LKYZZMDK+LZlf18gpEPAvT38vLLQ688EyHE1fOHe36
qlo5Dfwhqcv2GzDTaCfgn63PGnJneloNritOpp2xBp6FadzgTG4+FvUSlfRrQuKx069uCI98a/mO
53FFqXV2mnMsKGTCdPTHByNXg0MOMiG4zmzcnyW1oDtOgJm10VDkqnKb9Nk9KaUyVahdgOhf07sv
Ve4xHqbnKx1j+fRUuCauJLyrBKd7u7/QjJAOjJ+OjmW0hp8iRJSt9ru7xsY71RUn1GRhoNGAC25W
qxJ2BNO88WuuT8YENUvqwpBxlEmmnfIfUBu/s8lhSWDEx0zvGcxB9/AUsCdNPQYNKQ5gdZHpLV8Y
M3PoGK0iTeKWViuZO+qdob0xilcroJVFuBTUtOTHJw2axDz/7WjmMM1TffcWW9b1GzMByolPHGSG
uxO8sauagI9eyweWMxBcMr8Fvol8Avjr0VXaRPvjZTK33bOG8mvII/xNSrCmRXWD61i5gZGT7Rp2
29b4cHiuqLu6fJgTSt9Tt3+9LDg7cusmnL0+wJsN1BCjzMR2cCrF38xK35rm0t7B0IJtEUUXl38j
iCK4/TTAFQ6lmJ2mSMLaSG8IzhvdIzPLtaZKMG209kFiZuz94VXhq46+jgOp3g/IfbC0mia7ok7s
MrvVhiq4eIKlIxBa1sr7XeDhn4TMbyHSl17K+ioMBGOOnXukSNQR9BxwG4HzUyRPLJKtHPYADXyM
5CLRB9KHZh5OpQY6ZQBHTxtOtOMP44yyMKtIwHD42FVw1x+yHfdT6iSFdHce3NNsLTG67yz0APH/
S3UlPJ7er5hTMcMqqPeCCU1UbbAL4bB3hvSZ7SSr7vAtZdTc+kTzcWUKu0J6LrtseN+M/FCUwQy7
GcCh0xGnzzLG/mlsD5M+Lv7Q/8skaTg38HH1+KQuHUPGwxXxqGGo38jHsDfETgPauNRQYRB0z2uY
NnAS7gFUEWL30rd9lScVf1fe5g6GgHdO8g8fIX9soRxbcRf2B8N1d7S/o7hMKfGST7i2pexTDybm
KBrPq24WwLINHdgszwQmN5K9nzw1X/rbT9Kg8GLVsBCakJtNjVaUctAkXAv0xadsdBG6EgjiEHgm
O1wiJin3gCYbGI2aErySpkWa9nT1bQoV/LYcm87CnlMYU/8nDzOhbAwNK4EP5KMbvlz6vjJuzmYF
zk7hyiohILXjTbAyLxuDag5P+0r3hcwRIpsFQiC9eY2H0yFEdNzumz7GKD86554SCjrAHfoqpIFl
MALtUmd3bgNFVQtOJnQMyznWgFEqOfZSLJ3nJIfIylKkC0If6dY3d1t8uNXC9aVrR87daNkdHZWQ
iKb66whA6EDxHm1yqUNQAAxtlNg320D3HB4novkX7KWfbOe+WyRbjJffbsQ2/VJs2I8Q1HUs7rev
ngbEacr2AQJ6yqs/edQ6bmj26SN6cbjQLqaPrzigtK302UnANKrLDGln0KthDGCELzO2XHtpFYWZ
fglKskCqfPuHmS8kwUVAQrTlifzLyInN9j7Y4adb53ukXYfOcBnb2/+DzWDPQ3YYTIg603z7L56A
+g05E56unrQ7sA7leON/fD//+yvFTJyoAyEJVdmwq3kzG3VA3DaziGG6ZlJK7HbHgS3GOlnhL3jX
SoCi35RTkc7QjLU5XyhogTprIAwbCILgV4/59pB0f1Y6ZWyCL5J3Rzwy2r137Qs0OhE0ZuJkG8MA
VyidHVHeMewELHVlsBBNGP+XEKGewwbMueFI/6+JH3eZndQvdEvCPWm0CG4JGdwJuCUNK+iPIs1E
e9632pDncfSp4guoYNe2nKXk9u8k/VObFfyKAYmg7Ph0lBXec9NkGwif5eK56FrzHV9sqjyCmFoN
+78caNQH10ik4/fk04s1TRzpoSCyGDjTsOzIc/3eYoDKXotS94+vBcpNALrKbaDXpxd2RWGJ6xiH
L1X+jPRPsg5bGuSuhX7AhOoA4O3f6i8t5jr/XS5MFK36c3NAs7uPkrO313DhcJ3v7EEDyUB71dZ8
AD08JxlFRIgsq7uQXzpYThWFJ5foyGt0Bez/NsIJnDU+0P+zuIFQkySaCKdWSbzryM/OOVtOsF5b
UC5fgaRZWLK/KrB0xICy4FTuRG8AHlIJy5UEJaYXmvoBSXLMB03yVV/MBwl4Bj3S5OGsrxAsoZjj
XrBUfELx4asO1J13JTSalZNzgL4JMfuA4VumjzB7FQWBhYCMgsrFOgzBXQgBUSwpIn4aR1Vfn/Cr
7utXPcg/nd4RggMYcQqdQ29t8chbZ8P58ghZL1Qk9olntme1wIPSOzgaZjq3oCzx/HLXzWwbNO6I
L45RWH+Vpk+X4QfwiO+ELrtNLoKcKncxXYJxY8AoKujzM9943Bd/r4WZVPkwEdEciTmXPShTjDGH
CgAdc4KEj6dbZbnbk9kwhRN4A6UZy30NPH62EFGJaG6SM6UkvA5Xf7I1IogmnY8H4702E5PIVPXp
cmscTUaGg0MRbQBZp1ClT4vpTbwYG15j7gVvsS5o5PuxxNFSJH7RpOm4E9EMwQ0WFlsN6YGz5/Lv
2l5xbF0QpU2R/wwlX7uQwVCpp/vjlPV5lxd3sOmdLYEe5fQu6L3aH9iB/xd5bkIWxUQfLtii5QYZ
tWuLWutJEnrp+YzYReOWlcvDvnh0vn7t9egdRQrmIs5RXM2yUi5NxhvFdw0LraRYG9Ws3WUeDB7X
PsZ1nrKXm/cHAtZT2m0GCM8Hq5W0d9h/IrkZgsjI9A3EWXj7cHegr4FwDktyRYXh7MQ5mq8ZYTq8
537kxVuS77vw09yY8uSEpq9a8b+vw1FfWlUTt6CywH0RQVISfufRnEQh631B3LtkWPR6h/RVu5qr
9wr39ovfwp3Sm1sJHkekhcSo0qUcKO5HSdDr6LHnCFxd+hQnUq9vX+YQGtHD6xEy6vb035qA2WWm
/s/VFrVci39P1BFiP7XBvkBmctpK2F21DD+aMWiJqmoGZ2DoI8VDzT6ArSBcfPVAFZmgz/15+zDt
EG5nAZKSUOvpFJIJsl51MfyCZH9R3VjY4UVw1NWRnh9YW8JC8T8b6bMb1Hog/6UDnEaDxf+V9qg9
CpTQJM6ogs1R7jFeHvlaAoPKESMz5s1+X0dJFWCEVlwBoBFAGIozax7zseQ9WLCyYOMiqJtgwnox
cCIusFNdQ0IAhmF35D1e8Bf2MNNvgCMZyv9DK/s+8L7b/T4p6WijgUCszvvhSHtc086P/hf66K41
Me+N1GbmX0YNuh9tKyOAbvh/m/rCQJsSX0HnzXqcwv3JcmeC6X+gFOQtlzga/jVTXBMtbhIplkEu
fP0Hw/R6GF+5RuN8355afmNxx7FDllO7HuRnXBF0pciCFyjlpJucycVBO/jEGW8ceYhcFrqbRPa9
BeRLQ3F3ESDwFCW7Mf5i9RptcJkZzyXdAWsrh16nFfxyM0UQQMEws9gmsNlx4x6cZ6H7raOhI2Fk
HYpQoUOC4QfMMJT+Ohi+NWdbQ9+8k8Mn34OOtymsin6AD/T6yq80jti/lJkkHgRE3xGz8PKe41TP
OBqt7P+ZIXubVRl+PqupSV2vLcKJhqpDuGmnA5I/NHxBpuWFuvK9qNNHN91cBkhvbcQAlXZ6uLjR
XeHw/nYSmAdUvy1UCkCrwowaBGaGwiU6qN3lYng2xYDAa70hAgz79NQLSXtFZOFhoT0mYbzUt/g0
KGziMn1h9rQgxY2YgKSUpGoTQm1cY/JvIpjFFh5ckXAkHMNXgZDJmGjhs0p9/e60IuRfkXstNvob
0rBXpC5M01N9OHKaWZHSlCeCztw4O7AeudF0P5d510HI9TsnsHYDiTHWD/CfcTqNIbZZVS2kvxSc
AZ0ykpuQq1SYewXWGci6aM8Qq+EErxNu6K77o1/0hXIQ1pV4fmB6xibpFlAU8/w7u0RzjXgHQNzx
woLinPFhc5FPRK56t+Jponj/qeEyZ5vmvRUdVvk/uDssRyrJPC73+eXyZ0TLp6zZducY6VwR27P/
8piyTbLQT6Bz0+E5b9jEhjilYF4T+1vDT/yhVYzePXf8fgNQNk9+QTWcbicxb02kBuuNBVNj87F0
Qyc7QP/7HvEmW4L88Wp3VCUH2Vzjm3oExi3g/b9GjA6GwK2Oy9hXaajB/yZwYmW+btwGc4J1fRUZ
yBFfueejdpfZDi+p9eHfALdpoI6aKPWXA9IWunn/qvPv83zKZloQjbEt9N2Bx4xo+32K9HekWpVI
jqtFSzY5nAbKQLjYCQzD3dOBe0Yh2MBdI+XKV7O5OOQM5gMnNCRDBrvFpmr0pgEpbFQGKIRGKKD4
4GnE7EfNrA7b64KpOUGmu4tyUFndW5LbsZ7pAvbjZCNZR+3P0scftBvTs0c+T4/MrZOmAnYURmhH
GmJdEUQ5Jlq9mHGwelTcDK4K/uDB7iBZJLgVLrFswnphbow58GwatHrD7IvfL+vTtsPiVDb0wNiT
ynyNFO23P2WWbp7+eq2gzpKBW6OSrizXNZAQMCAcnoWOftlp7ZvogwKTvop73i2omwCMOzafsJXi
KDBcBReE5GQgTyWbNGVHkZ2Xb1wJwbrVJiNNVaEUMatRHiOMh+X+9qlk+R46/yr3pF6f8P4AUrug
KGX5ivjFdgdtGpuuIKYGmYWvvS3KpPkc7pfc2G+9EtPpVEl/hnXo5vbjlMtq/pP930SGgRxK0jWA
rKKehUktowI3xRuPkJa83PfIk/P+4TEsn2m334QTNFf4rIsARllFgS/DF8MbetROqY96P6Vj8m9t
TyV+R93/f/TbdCILtZwFbMGRsdw2hNlj1S9xQK8QUeeVQNBFtNMWrmhG3YMzPPs+DGGu9tRAYVFF
kUrConXvWM6KRLufJbTAXqBGJKocxymJ14DB+0xE6I4KA7TPpujYYGBjabF/vyJ9ksq/DHHxmiv9
mupdDeS50XO4a2/QhkWzkW+nQvvZz7gdzHm+zrxYeq1bPcF/fRDLlqbvKVhznXm518qVnVGBc9H/
wMHCIZCLMM39X8sNQxd7rYS0ps3p+sIqA+DfEu7QccRtIiSWwSjIyfY7/24kyOQQKQqIUUFnMHXM
/Jlw7dBigYUdzgnAaiapaJuwP2zLUH7qchkIHk4AuA7N/ZfW6WY0jWAzp4YRzle6eyXsGRg4ZfYa
PQPyoRiRAUoCDEt0mz7Q+EZ7gPRoMh64tNwx2g1zU1MBpsoyv7+v2LwrR2t+U8t6EYibbWheBiU4
Ulqbhkspo3GQHgl+3fwZ4Z55559upJLNgbue/5d2cRVsUCEFgk8DxrlQvYNHFbTpftP/ZEbcpY0R
/wLDEFmlU6uM8Cw8jCvcuQnhdEMoiIFngT5d0qzbVSyljXMYYJvGj/prPgVGOtc4h31JJv+2ul5N
GoF5+paW8+c0Q3SCC7+r7csGcS144AycFF9y5eUbOYfbZ8tHVG8eYphbWjAtTsM87N0bOCs2sZfz
iQf6bREx0JMzxv2/V5zxbRGi99XvZie8/bADsIJPsyBPr0Cf1j+9gRgD5+gw4piGf2X95zp/hjuY
4gApXYnrPG2qiLKmERqyYAW4uWXVNFfZsrFEdFxyAKJ1RhSnU8QEQ03Nf10c63uzapWkNtgHZZV/
nOr/DNoP5L0HbJuXc8phlbyfSDtq2W88U59fG8ByDZ9hUgX59ikv+jYl2FcWZ2fM4Rf7Y+K32xEF
EgqDXkobf/BXuMrsoLOuw+byLuXvcoGVidBL0HHLByPZs1DTkC6CQdj0MPD4EWLJ2Vl4McEzyIK0
HUppJEgRv+Cqy2P5AZXt+tDlhm9oFEOn+aRgwI0/sjyff1vRFQurqRT/bxLUVlQDK2J8agRX8bxM
JwhTwaC/IHOZgrPqtbrJAmOd14lXZuQ3o+Tzym60uJG9z8zVDsCSenGe14IUP7kpwl14h9EOaSlo
11qmC+Tnsjz5KpDDo4apiEhDAI7GGEK7tagPHjnRGR7svQjEg4gMUB7/XV6vAvzve8RPWj8eTp3B
9YmE0yi/GYpWlHdxMDlTRD8/AT1JMwLLdlQmYZhuiZHo6kavJ4LIOGAaNGlNZdB/0FuDLEU/7VVd
n14Ta5bY3ZgPyWDcGnBXkCp6UuXMwFBw5Gf6DWFwm3pYE8Egp88LR/lWlpp49zDnhBCT3ryRjOdj
6vuZfsn9IFW8IUwiEZqv3aTqBIbIg60kFM9Z6xpmyVqKuTEz2+eZzJOJxfbanO+hO4fZAky+ikQc
EHSKWjJQB3lxeOkU/U+8NxI83FoPrfgKH1sSYy5b20QxJQbgH8FvhWh55wn3chROI6TET/FZ/dY3
zvlZDtFbH2v4NnWDcspjNtPPC+yDtTeOfY4i0XFggVhtQa4T9cBGRji1I38mdyGBFrVHbO1NDhb8
HT60zMUy92F9t5tyuZKSYWMB/CU8Az/HeFZ9sbaEb/EUvrfLu0EkxlTRnUYRNJHcOgeSq3Wq8KSs
rQwb8Wax3hwqORji4xDIVa2Eb3l2cztm9YMGe6bnHQ93LbN+9YzVFnq2NKFTQY3G9OFR1iC6KH2F
WYVunfXD6rG9YB8wYE4RVXmBoWU0mH5ukm0zjXB8uZzL+87zpp7bdv79hQ2GGxQvh2xLsb05BJiA
upo1JimYWyv4ui6l3fyJXuC085Au/g2dfYoXrx0W8cxkPocmlerIfglHK3MBs4oPjFTMsTU2MTk8
/08LKKUHyKZNKJ6WCqE9W+9h2m1Nl9kdIUWW7NnyW5be6amZA6+bjyeyWvLWX55zvR+54ZW9hB+A
+kVMePh+YLrUPlVq34r5JBmxRraBZFSlKacpoqkbmQDqSzvQymQMeW/vcTUQnC+8MWURrw14z/CX
KEwBXBeQr0FK+QBJvoAoAqQK/tL7t0tFoxf9V/xa8eRVv6DBiPxwcs9FXKH5MpDpUUk6i1ejHbWN
S09zvGngTJi+9S2JVm1ZORwf1/DPss6ngwkkxuTKMofjLPt1YpWX60ftC3T6hUCylGC6OvKxSrZ7
/Hk2eCNfEA+athkDbF3V3h5oOgWxaTfPwUkQQe2OtcnNK2m5c9/R++K66kqQbhhW+pOS+bu0XONH
KSpPGFbFKLiQteb5ve9alC7ZbxqdXFYNxAJUiEv0sLsfsopOhy4kyh3NcH4vrU/t797wLb02bOEB
FSG0qxsSHytOacYb8TSw3PhgHdK+F9F6YGWXdCGRCN4AAgCX2e7PHLaY1i6wuvKnFeevjrm0Xvsr
LuGEeUYhzyRCFjL91+f7R6p6VQppSCs+LSql3C+tQmgtGGcAzV8r/SbvAIIV4cjdt7fFK+yfrKSB
RS/3ON8i7Z4ZRCwhXaAq9QqIPTdT4++6gHVppBg9BSloNvQ+oN/SVQV4ub93bv9kSii/rJYrnr8p
XyexfFsEs8fQFwEkcpkIJU/X5l2FIOZdG2y7jq2Tgwz4g+s/7G8zxYTUfYhIgEb+zJsuBeuzKQX/
iUojrkQarWnjWMgpAKL/WK1CVOR5SB5oY5YoV4irlUM7QTwImOibM0OcdbNWeHeAwuIIXSB6zQt9
VRMJGMnzgBIvJqXXQxndNlMTizhI39TWDFHb4xdAh4IzbMpnUOBHk45jtcBtGw1My6KW9jEL/Wqo
g0H9EuANuMbEgasq8W3UfEoEiqQH9lTEBTNbs2DLI3RXhNRUfpIi8IEj7i+IU9p616BUAblm5Rbe
wxosyrQcrHY4ApEQN4IvmYWWN83Dkb9ZyStzRX/6gNfg4A9JnZiDRGhtd804iDBag+AijxK6nq7C
EqI2jjm20d5oe+pcZT3ooDIY14nt7kMh2MqUYH51MylFpQx4A4NgId1OZ6iZ04Txc2Ax7M+X1oUH
pparu+dhHK3t+xMKIVRSbf//CTNKaf0ZgAAtwLhRUc3U4/dKVIA+JPEdIjBdzRDxL5fBJ4plMNIa
kA6lbg0Qq4ayVeAI6SPUYTmZPz1ICuo7mE30zEXi+924rIyZpZohgZfHwV/BMVZEzD53aWfh5Yam
tM/fn2GqzQz/7zbzVjJYr5dZIcTxT+GBdRPKpU2TbHMnMU/s5z5WnuP02CJ8GbstffA5XXjbn+4m
ZGgZ8MrIbG5vleuExyT/FIGx7W75PZ4P6gp3Y3Y17U3FrtukvG//24Y3TtgPcUezYREbQV/WVCph
pxGiG2MGIXyQz/jzdTfXy1aNLKN4NgT/EFZ7G5hHjs0LYcuC2ksgJ6tSAvD06pP9gzuKQ8q6rUZq
zrGWMO5WQNu/J0SCZniyBg9aivnFMsbL2DUoSMQMTI13k/+UESW2sSGVCWCw6edewxNyx+ramExZ
+yRSRMlpIxX6fVNgAVjezaYlzUUCw2e+zp/bTkl3CPDYSKAJvkEHOdya8hmj7652h4yJ0TB7JHor
EW3HBr8WG+xtPxksivDF+apKvNZLKsoFrla8eYmZwn76aesGI/ZNfYUimTiEt1u7P5QGLy/21QFZ
ya2UWC0kbDpwIKiTefZavGJNRcDStIcCvum0hoIppjLyHHRhJoXTTQ8tRxoBMZP1cFe641/ZeHOk
1iuzKLeY/Er3y6tNJOJI2HOxSjLkIriIQW5fW9zppXWbMS9bVP2C1KTl5EexLHkrLOCyMWq71aOH
juAfNFJ25Crdvgh5FQMiPTX0K3XuUFSutlsZ9FBMUsW+mkxW02xGRWGJGezdXuypROsUg0dVfLBe
5yzGwFxyGom5Is/IRIqGIR260bexHgx5mOd1bG18HepOkEf4jIW1kTbHPq1eIyiy5407kmWAESIR
nc+pz2yLdmiY084aKtlAc6Lx0cbN7rvWFxL3ENI/hKUNkvt1zI/4a+rMRyoB4MJ26OEfJkeIVNy7
Z4KZgoNPvzrzczwNsc10C3MZnmVhSZX4DSJSnCluubRvv+D6xvxr+Gzy4BYMo26aaPm8yxx9pKAR
9qOFAMw+o7Pfc5dGh+sTi+b4Ypy5jqLrklk97Bjag8DbaiA0HwF/NMCw85hN/coFOtlOPsq+Ocrr
Drenx2lQhcBnvGwU4++Lrt9jRXcSILijl34Se73lC+3RGqbVEpWPiShLsHn/btKLByus2mbf8Exx
17W+a0QrK+kZMUb408HENISXSoKEUCn1xxEGCJbxm8DLeZBWqvpJgjtjq04pjDYh5Ls8wdjpDKE/
B0BVxXFBAROCh4hngoTL20tVkXQYSTv3BWLHXCHYkDYRCyYWNZwMDL8NZ5mgq9DceJGJ2La+BitN
hzd4rH/n5cYefFSQnLY3JVip45DW+C/r8HkB6DlYap/3PmWGS1VEFms5FaKzN6rDLflzxdma2mt/
0XvU2Wc0hlx+LRe2CfO88iPxSvlk41zkuhpycd6g722DpC1zFk4hwqoiLLfQpnaOlQtPIRWMlCmo
qbNt6L8wdGpSBou3zeiQlarQ6aqqO9mI2vgrnNd4Ct3cIzenhceHZ7ylsvecIaGnpv3OSrgbSlL1
/2erR3nwZrB134hQB1byPJty0vub/JoEGrokm7lAZypnadxOscc50sYF4WGWsR7Wv820jGSzo27M
CL6veTVU2Y83R0Tnzc4oF5exA7Gk6wAyXQK6vF0nPclkOncbXZTpS1GJyNuCT8/yyV5Xwb4jqgWm
w6fFpeLFnCbg8fnoAYMH3NXGaFmqeBZvhSU9lNqyAfRgEuNyP6S5qS/nyv3EEZMmZ+4jfeFAPVAd
abKRn+JDj56u4Q6jSdV4EOiZrclsc+/Xw8mPef3dri3uPu1KcTLIU2OpX0j7GwxMh4yQC/+M379c
B9PYc4MAhHorydrT68KniO/phROSbohU1Emq1KjG2mfXF2tmn3YXm10OsNyzfa8VylWGfGQz+qiV
YjtgwTtzJOOtdXL+c9IzyRAPr5tkOIqpr73haiHS08vCT7v+3cYzvlpcA30Bja7xjh7e4rMutGSj
Qr+PlaG/QlnAgUfajqUfZmrSs8z/S+zgX+9yd7vBpa3lPi1halyfRY+HHMDOPu5E/PT6lUWbM5lK
QwlyFVjnBh22nQJbhSnQLlUt6R/umxJb3OJVpcrbbA2xKES3HNPEw7SOGyRW+kbXYf850Nzs2Ohy
scGifpwkvcRwcNyxXpBn6Gh9hr5A4jG6I9HR91NUaEnhUmjeN2PxqZXkvkLWDYHi9O3bZaAt0PTk
WN/Lkg0RmY8gVjFWl17F5TN2cQv80BrotW1IVz6EX3OVl4S1qyWQzr9sKNvFRDLc966toKmSGFgt
sNByNMMRWnyAe0sVFSpjTuwH1IMCKdtaEQ8QCWGmfQ65JW3CKKdc96l5i+kQcYCu/b74tEFr2OyK
RbnrLoH7Twlw4LZaf18iom4CIJ0a/hbjB2VsvMHcXmCx/3lUV9UzCi8OXDFGlEd2dsk4V1GeKMIJ
MC3oF7vzyd7HzoB7ThmvDqRx23HDUgsCHv7fBEpqHYLuwmMyd58w3yJ3OCp5bHh/v4ghAIZhwStm
OawLEhKEV+dSy+TOiD+VD/8K0dwCJDbgFPK8H+W/QizLy4zhsY4j7H/OwkTwUrNn9g5BVrhcJjXi
opgoEZy36J323bdWdTjO8pE1ULb523B1OHHoe/pUNdIMoEnJOGUNPLDtqGrQWJtu/HWKo8xA8jlX
CIUJU0vQBWjBUAGq97DwFs7qgy8a2dvTRenmq+qCkr66j+fuGpo0KdZ+kkjc/MpSkWoI32dYlBFN
PzGj0woMge3vtem5gZW/QHqSUkYoreP9DSUWqPS2hiKav+ZcammH0JqoRQCZ5Yw0dZFKO6jCdTWA
fHWR+MqMPlIwQLDYeZwoLesViueu28T0qLGcNpTvh5EYj186PKc1P6yLbnNmp9ROz0TxUmGGw4uf
dEVQRefJCamvR/xeykVESCJtJxlHDKPPI8WnaXrey2H96SVhChRw+89fPJXxbUovMuUdjgrFLPh3
h5pz/scw4ikV4l5tAuFSQqT3+haTxTclSAxFTFEcAGvCE1wUyyb5Sw9wpdhCE5NvJ5ujYRVNs66W
REZhQvzZQX72nf2s3A8tCkwVp0CDXMAcF60b3itIwR9uHb0RXFlMX/2ylYWBjDo+mtwM25bdAmmP
nH1s3oZ/3DUyZx/hDCykbU+/1Xi+r9tsAiUy9GWA1XP0xd8o+/oT/e+CBtoHKuN259UNOqT4AscO
aC6kseczNoqDs6sNSqptucrtLcFJExcXzkjbcMOJL9DnV8SjE+UeRKnnHxDIhF/AVVypn+F6aeNA
f249dGt9picQ5n9PxXCsOLTpAjRNdUfWC5EEOCnlrAe0duWITzFtw0akfDdCSl1Z/ZmnLzYoXHKz
TRV4k98uL5CrcA1ejsj9VWUnLsqgONsCeJzRul5+p24aymgG+40gWcXmIoii1YkjidgqM28XSeQ3
H1KWkjmSbS/umCnL+Pz8NcJMZimk+8z48YNNQSVqBvXUwNPf+g+jwtrtw9wnC9gHccIIMB+BjpGL
2jQ+JcOjF/vVW1lDev+0rtnBo4pGQmiQq7Vxd+S/TEKtk+ABlTRFnZ16UiEHhkokPBrdgxUndedy
lPBO2cOt/XfSFL0Co7NuPfDZ3GmBCsvUCV4lO6VLflbW88PZ1M1z6h3kpVYhkMftll6l/3o7884C
JMqfsUzLNDiNLP79f8SMe5uXHo9IzUHYx+egY8PcY9/j3IsVPj0Evz/FnpqBegeRKzQUnegMI/57
BCLGPIvJLGkisConhIqXUlvndcalqplKqwoLKtbj0I4g3s6vT/VlYaXxW+Gx/Sb1KAH7rlV8Pyu4
Rrcoim/tXQNeqSXzw/RkS34voJAHMYNnkEWOWEZKRUbWtan5eHJxuvbSIYT7Fq25ZFOM1CBO2JqW
Hd/2pkZY62MeVsGa3pA3Q2ZSvmpS5ppSBwxoF+txh5tjLT2K+9esnSopDUs2QSCeLG4Obcpu3HkF
jbPn6A5uMQruHJ2uhvyznHva3k0JnWhOkR1b03MzmQIiwlUEbjDTRxqWmAvb+wsMG9y5jygo+RWq
p5IhvBLPZNe5GRk15svThiq8hNAagGcMnupCHTALUx3UrmjLcm5dA4NXdl1Jh4gsQ81cAEvxBjVv
/c4zz/xQmz+bjWcai7THNzayp5vXf1km598JJleynJwVDvY2g+zgzkeiRIJ7eQPuosVv/WoT25Mn
Hk41rfszYy7xRLzmqL0yv4nY2Pn49u252HJ6ze7MM61Aa6inSu33T0zlM7eLbjFg8tnh76uBqCa5
2VYgfZSw3qoF2yohkGISSZeDqymkAhiN4Fku8562KrtbMywDSw1JITdRoywgvEE7L6+uttaJuhRz
NH6FDTKjh+ALykhncHGMZWrOM5y3ITV2O2Obn0QsZOHa8BFqVXORp8z8GL79rxQM1OxPronlr1qq
RRDX4Jiexxkwu/IaZrMQ+5ULO0jFc7IUNGHhUF+DWUIjDobBBY00fZpTrs4STzShYXbP1K8s1DVu
qjGPQkmBKbE4GVsj8wYyDoO1i+U/wiM0sIGJPJ1KVqLu7PFDyTh2E9CsZb0db+2ElOYaKmQT9scl
vE1xLa1RTtqXSNTfeHuvaDIZU1GBKlB/wHkNkJ7H87djLuCs4B8rgYFWVLOfsbpIEw0qDo3LaBcO
3a/jnq+x0vn071vXVYf0ySD0DdafsHHRIlgYtwcol+A64JpjxVMVD7lIsdy9yi7vyzDOw5QVxEcf
8zLFZmU1yPPBxvh6dPi23jlVkOamVbE0SP2A71mh4R7Tw7dmP6a7OIo4b3WKI5aIj80VynXJ3min
iHrRUvd23KT6LYGJ3CkBZU6aSAx3GHxYqhqq+mXYUwT8EMRpIkwZ/csxO9hzOLl3XhfD8OGTRKSM
vQ8MBoCKV/3Q9GImsRyb9bR342W+NtfpDCFhyrCTbYTwRHk9qoiUi4AaJPzJ6RdQAIuw0cF1kX9C
cZoXojPo72fkpYtXO82NgJfSpaUikgYkg+RlWUQZhFQQAIawhhcZGrdRIsY3GEzEjm8fEghu3RWN
1ucNKnaCmyiVSSABEzEb9B5Vt8daGfEO+D0krT284v4tInv7OOQycu2WDJoXSSTB5JD6vPeU2mHA
FUMdF/OqLcAaM84yEbo3QPTf2LxD7BWzbxKuTckHOtK04lTZdzAgeGO+AuR/IMX92td5q1hgVx70
2rkmfJMlpeq0xFuEAmHmje8DQXQ3qdvF0o8tTO6Zd6HA2YQXf2hDOz0miC4NCWWURq/nrTECVVTc
CzN248dZIdS8w45/Rg2iHUWkYQ8DVVgQgok00sTuQSzsWzCNBe92WzUCo02pTl/Y1esx4BlM5FTp
VuOPyQ1b/5poQuVU+EDZcm1LgblX/E/7buoieZWS9z612bg9VGbcq0yHdyvef4RHe3/vT65jWGKr
ImUMGCF7/eTwXiP4YeP+UoLHaiISha7ph3u/Avo3ZUrbX4OqawoH1++e55nlF/NktWVT9baKI/Rd
6vaXlG9SnHHk2X82r64QtIEYCSCO4CgBVjjEBxGsF679rtm029hnje3eZ7TQfAtlaHv2HT9nxKIE
tQ+cdzXwpdG7ONUWwR6Yk5YvZq0Rnvi8/Ky9JUWYWVTJA/IcbCIGYo4lkfjmqviOiDaIXmRVGWrp
zQ2j1K6joEgWoT+Kd5g/pJqHKaQUF3rN9v+D6HjwGC0Wb8F1p02al7Ee9NZ6s45qOXrzuoGyRi8V
C3YTcgZ/vVe/nxFhoeCP2dDQQRqT4CItzRa24PPxJi1ep46SJ2NTRdCGOiHKn04OXshP6MrSlqQ7
PynY7Ubzf6sjXa4xytSVc4jMyki2Ug/4UhFshRRrDqdX4bpM/K1W1Ym8j/3ouus3ZLkMuXzCNNgj
jrqpS3VH2OAW9+sWsYNsMeSPRUkSFpkQORbQuQaVV7+Hg582/z1wR0lBnmCC82VuETQ0qnvLRVMC
HEGMYAk5+CcLaAcP7MiwnwZIA7dWgiHP5CzzfOMLWIV+OIu47k1D0h5OzTs4qph5iCr4xRYha2Ev
biWs6IYa6rQQp1qKEn8eoByL0O8hrDKHhee2FoCinPd15H6yqlEwN8zj491DB+/Q+nhbXKc6ZwBL
AikcGfwhgdykT2Y9/eaHw/PkT1kFg34NOcaZrlfGsfrManA1PIjuflsym+9Jxdd1vXuMDAYTbGjA
092orpr9cyH9Vv/DZc4Y/dHCme2qONW8NA/wjXCUjOnXWM1r3QTQqodHK1kVvBKgGNQ85n87WNGa
jZ0JTigakdcElrQz1dmCUfTa1ZxCy9ZF8cucYDygPiJLk+c2Dr/RI9DaVL8kbg3fAot3ezL9ivOp
5i2N/Rkc2qVcAFwTmGpHGADh+fr5tqXG42K6DlxbSGd3IkA7VLvehrA37bhyyo2BRfHtOXQoZk51
PxxQ0GuOVXBdfTk9824T1LPHRlEM7tgYDWsVtcA9byoEsxx77a8B9ZuGCwfSI8xL58vit/gcu1iq
g3gADThWA61keDFRv4J2zS8QCBNiI4G7UjjAVlPUffcyOBfcJYpw6/0T2SwihpovrB8Z5Ox3j4xP
8CV1fRbnuJ5TnT/pfByQFdIopdi079L/W4/3yKUqftWYA4GdXHaFj/FxRsi/SYKK+RrCTWkQDGK+
NNcmg1bIZWiQxz0L8XwNCLUw70L3srGOGXupzL8g8fXClmuI3MjB7AFF84BzEoOitIurExlNL6Hj
wAC7/32wfLJJzUBF2+JCLGWoibhHH9Xqsv0e7Cp0RHGy9Evp1Suy6SluFqIk9JdzKJ/EriHNpIrO
I9ScftPhdYDulS1k01nNkrbEs7HudbK1q2LTuFSDmZioEJC9w4VZxVXCCT7BEDsEJLNRqko6VCPl
/HMlAURFFrZhPakKz/ECVPgdHOCBpIOx4D4J9neNTtuDi3+qlXXHYA50dC62rL2uKF2T6btqS2wY
qPS+juXK9sEGtxeAJHBZQS52zJwtwK3QLvqtRkxy94FgdMGk3oHHRF5SjWkhFme9bEQ+f/Dr4Ay5
v7qWH7jAZBMr8Y71i7L6k+6fhZ61iuUFxhoHtlR5ad8ag5vWwIRswP1TdjpB26LSH6GSVzGMbgV3
KFilvuDmxxKySo5W0yNo/XoJzAb0L06k598XI3+LvTRrPSreve7HqjWH5gLVBRe3rHMPXBldPzOj
+NdL9Zpab8gwHABSdkprlOX9oGC8Vu+wgq29aVMchMuFWrP3MWO07JT9fFmp4QDS9uUN56VXm6T7
zCcmyotKFjYDmkf9+lfqrH4OLa4Z/lJ2odqlyEw6+nycE8e1IW/vjwnr3KJxdfoxoVNr7IjpgKBH
sYzqWsNnwSDSaO6NlGJb2AhdP6VecnGjpxtH5tkauc6o+SklVeOiS5tqnZW2oMWh3PB1vJxJz3Qj
ddUkC97FLgSoBYYPQjv+fXt+nmJoUnVwqfcyUQ38UqmDS4GnUKNCjA45oxLvxWLTr4bIVn1h538m
vicpW9dOtoIbZlH7Deorx+5mlcarhXJeE7bScjNzoYSsAS3Pj9uaanxYJvjJIQji3g9PiUTw9hfw
MeS4T0HPC6zMecVCD7LKR3YShCTxfOi2rHqgWDftoff+GUyIVi7XuzFQp295HXjog2Z4j8PcEobh
LHT4xzVy9ui1SLFc36RTw1cPOf64jLSxYgTLwaUl/25vR1Ed0TJBNyo/AAyOpObUNZ6yVDXiwY8/
jN+WQnGMBBgKnLSf90QD30nN5tKN5ggJsRjvrd6y4xv1tRC2ZJwOaVHkZE/TjcNvDNITWxg3HFKB
JR69TV+qfGK38NiJzI4XzWorenK5IokA1Zox2JI+vuODWmIaMmd4Uc+4zsiuLvmW2KKnko3Zaixa
6cMgwOApn5TKCDcpV6Svcp43xJUwDQI3kFIIStkvMMu3SC1bbFmy2dFhppp2Nnp0FAfUrXQJTPxo
igdB7e5b8d4ufy8vpBgrDeZ7hC+J7OgG53UWaE08Ct8rb7PxsemOACQv9f00D5khVCF5Ank073IU
RhdYUKRZ5LxJ1G+K00dVhFz9xLUZ8kSP3dUmA/OJEIokLWUCUOiUyn0zl0ROUfkeLPpCCoUOknR2
mA9uhErAAuphps4Du2UOLAxf5FDIrCZJrbxgifsVafFloSEu82iR0Xum9JNmeO+HWREESGuuqaGf
uYRV6sMI/d/yAVsUGbw1Mncm5QIud3kpGb1Yw6WyM8EJXSzjhkXioeMu4suT7VsHxUsUHFOAdRX6
y6yafF9tLw373m3TaAcCK7mzoEwP6ZD1STJQbi6sLzR21dVHVkjNIcxiphGbxYa3lm/BuNYJ8bc/
BYGuFCvp/6m1x0n2aid5JAa4/Yhzeey4oSv1Qy9EGmfphR3+Wz27QfsphsE8Oqsh1/fUT8vcPbJB
EInW3j2KdiT6jNsa+EgF51GFKvoULL0BXR/Og88OLuk9zrq+Tru9eiZqr1I+1DRCy/8nxSjB6z7y
/B0q2DBC1ZvAsll7Ydem/HsbRkKZYPUAwETQZH3vL9UnVv9IIZVjpXC8SaFeJIQ14PpZa/6sx6PT
CFQtpZyBo6oXASViMbuxXpRMB+hBfKurg59X6TKoE2tOsAwsPBc28kMIAhWnhdK2Dl8DLbwa07Dd
YZN7Jd0QZE93wIMVshHXXDPhZy2khGXvGrE26Uek4ujEKhWRzjXVE1J9QFeAajPqq9UYkEeM0r+I
7JjIC/qw4eEYocU4sS8TG0XfO9+UC9fmOPWS8pvv9HIOxuhdzYMpKtoHNspk6w+DaGaZptSuPYOs
+g2tbPr3YBXAcOwNkAZHnHWaap/UaJlnglPrZ9OedllX+N+PhNbNYWlWesEsyc4xcVELcxEBY+5Z
OZHwbe/DuKWdnA4O0qcWhBtgM1aImWunrr3olLvGhjyJOGmJGUuCGy1WiSzVtmoTs0GxhC4Pa4ZQ
fUxasZ6440D/oNNXC4Y9XTykPsU3G4YxsWfTehxJyR8MSpY76ixqFnIj4tf3zm2m4UGRDMSPA6dx
tDPlo7SqozDbv7BFSA9ZWU+kYZK1Vnv6HYrsLlkX4yi7yll8Tkyupg5eDEsmiS8mDTaF2H50kITq
UwU63A0WwUaCE9A3mOho44jsK9lC7vQ5ccXHYpVORr5LEGMFrawNOViwm86p7rGsDhWrMJCue9Lp
sc6Xbhq1uqFojnUOEcJmof9SMKAh04bH3HXyaBDLH/oumU/lTfNb/NwdlY5RwhcnqtUondxc1NQi
2UDXdiOA3hLVBARhrYXaHbLUoItf2fuSUFW7SqNwqIlxInLthb8aWp5DDXJ5FA+AzHmziJU9qj4m
81A0JORsjkW+4EC/WvACTKsyBcjvFELKStU+Fr6AgCW/RY40weT9ez2MZqBdPqi5Jynld5qkYyBe
JnKAEwFM1vyLbrrndJ1dNuynFfNRRiWyJ8cfOfBdndW6SXAkwlHB091hn6TtL93oSeGfFKtfpzMC
Hfx9WgjbxM7fMfhYdbM9ZUzGwx6lhiYE9eV+f6yWP9VgYBmkeNdqZAAv+SBihl4ejKRupfWZW3CM
p47TtKEvbSy3Z8hgUT1U4QeDBdLNQQ2sTkgGgDNZyyvPvzEIOinnMehCg/EKK1TCQKn/bityjSC0
KM4sQucD3XX2OyJV2lURUnQYq880cHmv2eJ79VSFNULoyg6RTQhUA3gaAVQYhO9kpSS8+2ixGJKC
2rLTtzkPYv6Rw6a0v9OjjWieifWAw1kBFAsKZOADBkFPA+SnCdiIan3Bb0+kw0GGAufWazgFig2c
mXO6IGUHz/TR3cueTGBdiKR6cVcugA2lrv3YSMmkrUjn2wXf0bUiJrKDlShBH4HD1YTh2NR6Qu6t
zz/heEGTUlW8IGc3pxGfWy8AA9d9B2n82t/0+bzAVfJUvwUWIkHceFtjxd/2w3qzyyJz+FliGuLD
uP2FXgfF27wd0du+fESakrWQhzT9j68iVm0KRYA+cpP+acJ7uk02A1P4Pske9Cv1Nr1k36LqkXYU
jR+EHUGiZ8ZwYCqdW7HDVgr2bcm7yYhOdqBiPrrhFi9CzC9AR9Lwz+A+8p3rMUCVqvTlraKvnA7f
pzPcmQ+jYcKkr9IWp1hqh1vNgOuuwJSEtNs5AOB7fFXFWAo4PoS9vGea+cSzqLXI9IC4nAxJz3B6
emONvXUcAPNVxOOwrjR6GcV6CppqCLG2hIy3wW85OBQK8UbaaJByTyKc/o3Cyt9G/sLt+gxhW4Cp
06P8/ifij9xKEGvbvQlpoHT+70cscQUA6IGbIAQaxXIAjV/cLVRWyArgviU9nVpYox9XsrrmjDQs
x6XoPaXM7V0pfICW5WhvqndN56agXc/Qhij3uz7qtOHkhr3xsPM3hKXeHEJ8LE0QXUOKjZ/ndb7D
nsR0tFZSzpDxrr9/79zBvlfzsjklGZ3qR1Gaao+ede0JiVzjajnBkFwrpk+tFTHhpgVDbovf96KR
VCC/o7SVM7+0y6mMYnfpcrLsRDY3s6XTmpzZ9qMznDHsAVAA2XzRXnYbptelLj2bNGVNl4Bv3khX
YQBGPiOB4hrXFtlGbaadvPjAYQ2hzRfHcsDJpPes/9syqws7TUP17okGNMCcP2PPY2fjDv0m6tdd
aVeNBE7RgA1YAlG5GM21MqeOWll/Rp0aKh7nhFtpkuhXwr2pcuPdZ8c5g3CjR4svZq/dEKCGI9Hy
O1lhCDmi/HZ17HeFD5xZJVVq5jr4u3F7sz10BDN7Qs0LLRxPLGcQXfdP+jPt+hCR18CMDoTfa5Mi
uSPndjQARuJ0sr/2l/3OFv9fbEs2T1pTFbspoK6r45+31DHxySbkq8BmoUh53lVV+XaMS8yzarqE
z5O5mqq1x1RWmQkaRJsGZ7EFM/txPtvLM+ZiPcv/wuoNMXbKmXbUCniEp/Bn+s2ZrsyJKQAOHlQE
N3QnkmbGmalpDU+UiMOOQrZN8bu/Zh/Q0JDpPWkGOIHfxHUAwHkX5aQXI+uxt+cp7wA2Yvwc54vf
ha+gi+VuzKwzjW/dLWOCgaYrD7+s9JdzZv3YWrOG/j3GpNwN+WKCA7p1dJRyzFU9CYTs4FAHBfFl
lzyXvC8zBf8l0xaFOFId6slV8feb/3gwqF2F7j9tL+mFAkw+xUKhsSFBRgZVXdK8pVpTFdzmoCkM
eovo5IjYAuNacCohPGpanmWIEddWUJeaxGRAxL5mwforBUh6MeX475EmvIme/Y3atZcv2hgEBqb4
H3Xxi3ZDk2LAh5SMfVoWO2oqCPqbjxjCPvc+UEL9tIQaNPBRsi5JEHS9RBDSEHOuNfGSHSgUn4qG
ISry74RUzPSnS5bq6+XErzD3Zy2KJsL82ZqvSEYQScqem38+i0ggOTZ78aDhB2iF5aQy+lpGV6oe
+nSvCG4+AH21xHUgoQ9JMYffFWOee5afxiAdXI0bQ0Wz5i3/nAcTo0JAITrN0j2PFd4myc3AK3gJ
SH6nI+kbCz4oerqX4+ng+N0kcWVXLllozVoJEZZoJoJluxry2Hzj6Cymxuzc9r62WD/HO24WPZVs
LvrK5fjbTx7jw/8liYwzU3hIo0dSZeDBy6beljayLuJ2u/tod2Du3huQ220VROcRCKrmppH1mJ0l
0tBv8yVq3KgKqq86D7QHXUxXAzduWkHJ2t3Lonv+zhfOQEpfNAHDXK0Dv3F87U8q7yeQbGMAcoV/
Pcmoik+zzqPbWj/LVBsCfvCllqBEz80neaIWvzrmpdyQTiDCc3VKEq8yTU9yDkZiGWhvVfk41RbR
78HQuIIZGERH4whhzmAYnkQSrFbAh5QYVmXmWRZF3OgTdiIdmW6zzBFYI2dDIkhhC2uMBbMyjLRe
GmYqzpfpgJSrmgn0iBmcU+XmbaO78svzZOdAhy2L7c62v8MLwGHH86PznLor27tnH0PG2bTV/npF
MXSPd5faMFy6KaSzgCvQNr1dW/5OeE8NgrQfediu0IdE20gwStCMH8Lfl4bLkyF7mmQpX7UO4F4V
5+Bcy4128pU9JUu2imHodEvAPsB9fNPA/67i8uRahQxstyZSVWnf16F7oQ85fCukc5280o1vBPLa
SLxhwxL4+rZfFNF44ssWjw8+ygeU5dcIpPTFr7XF/3YsKhVjCVkpYNn5w2qP4vKCWHC7Qun++FEw
EVkCTBuP08KhVAdb/eHMtR0kMCopKp9gCt4r4Alkx1cplBFjyrvGIycsG2/JdVoCeCB0sYCEgyLs
HhhEAE/JskbkwgVxJqNvI4E1sfFmlVMp+1U8z9F4iHupg9qd0rIbViza6dxAGMRx+QW7Xnn/tJHc
O1oDmrMGo8/cyOZFzUyyjjJ8hNk/NCZLJ20ywIo10C+Yy5Hjhk5xT3Fmca2ysz6OYDzUX/PBN7ww
EThy6pZPcPa9B2ymgFefwMcKcmNlVPY5yO/ALhzoFcWR9qFRrv0gU6cqWdd9IhPBNtZdxwfWFe63
JHi2GWz7oh7Oj5JeGFeoksxx0VRSQCIjbMkHEHizE4f3R5rjicL6Lrpx6Of85oGQSWAWNfidOjoi
zw7Zhz12aceujEXNOwcMQuCobo1JInkRhstXHDrvCpxRV5cAbklcBnrZ/jjFSRivW+ubqCxWXWa1
tFSfDzo55E9swoO7vv9GSPByT+mtqwSL/NyGS7h4WP1w2LjMCxApCHWZqPBCMEZhWVzGgWQzkPnf
cesrgA0SHpNCscQSgR2XSs7USHZ55GJDeqdB7+ercOfx7/svT8ZYdDpD1IopvuIWrxuwzf9dAngJ
WV37n2cd1PXH5AbLWt1lwZZy+AEYvJ2EH1Gw0ddOMX8tfGl+sKcxaHGwsb2UDs+eVOSt/6xhOloh
8DjjTP1gQUFQjRVuM4/NNjdpoe30Rzr+jgXzjchQMkpL6VOHO/GqGU44uN2z2xJcwF6SqzvKwkTp
sDjVJGPloty+TOVaikx+Tw78oy83MRPbLs0m3S188RTMIrF0aZ6rMauofevaZQt609f3nGmcD2DT
m0ODFhWh70zJSps9swQeP/naA11g6HES7Dt6SwDCXTdXcuebPXbcqbBR6nskgy4yeJY58f2htDjK
Yxgp30/Dw7x+Xez+l+HEp40mRgkOyiP8RNz5uMplRg1B88FFFabVJhoVSIQGOBsCyq6fwhPovddh
6/dHMuZTL6t0+lvBFMwGU8tWllyAWYVMPaPla5GfweQ6s2+9ZVb+SBHHriKv26WCbzTrIeN1+Oml
MRSc5qglu7FlP9tfzOaktSI/NLXEosVL/WncGhCEkGwcCBGXOE+OOFpYq14POQL5xavdI++cVYkq
m9aYWf3E9DuAEcAakK8dGWUQuFZP5F+rWh+vs1+wA11V1p19Zyqib0rD3bfrDN9NtXx3ZfDXg275
U4/vQs+Z8G5rwXMIRcJmYXmHC1VQut0q3gvyHGjWv58kTG99eOUBJJO08M8WeX4UKK9I4bbvpXC1
Ay5XfBUUtCo7QbswgmA1xYVIpdf6a9Li+/Zj6viHU1Bhi+7csiujeH+pyp7DV4fW1WTcY8rAcsz5
z1bJmeFq8t2JBjBQalYRBVNmXUyY+NaR7RfCR+rzhdk8x1GIiQoc0ACp1REEyA/YRLuRJdTBAM7x
VFnp1t71DFIJPW9pT2tLeyEueN2T1PYsMDU4uuWCO9RLY2MxPumO71MCU/r4eAo8rzotEjgbnqj9
wFzQAGBiIwUK7QRIDzNHKTZZd0m1hciM+G+TDbgQeYakhi2xFSJqxS14EVCNLqlZsQp+9zzZhLPE
GbpYlQNS8LsWvVg5nuPSMOXgyPBYiC7FEkdY+Cp/4goBGwhFW+Cr2J1F6TMqcdFyMYj8yqgiNwbW
WGB5UYp4evL+pj+50A0Ap/ygoKs2OmRPgs3RO7P8diA66BvIkMmDjmgOr1v6DDKSh2pvgCni1dez
HGiK8/5Ezg7pMskKWQGhESD55k6iIEhEsjaYW3PIxQz3QE50DiQ7kAcW3eWRA61cRgJAtXnZOXr+
Qfa2+F9G9rKhRDQXxc40TUk8pd5jdTtcd1yVEzLd/pC1lBrVFkqsSOQE6X0dCFhSDaWcaWEDALj2
v3mn5C7hjgZQNfrnVnqXXPK/+rJSdy7m1291sZuHj0bdc5b3Dyf4XoZ9MGmeOFWHISzdrG1XI/dV
vIiQYiJnq92NSOwM3YT11Ojd1q5yXXlAG4O9EyVtnB7Y3DzbynjxYWUPsdOiLBWncqTMCcP5qKMo
YKxlnm7WU68a9koBky0TiHByf6agD4e1krDCgCWNWOurCU/aqMJ8NGGnpnL7VTcJVS/zpIwLJMXq
a0Vk2mT+qs89Hs7PvuZkt22CPdAWCiQ8rm1mwtJhoXFTVweXhjkfwCiav52BY6uNGY2xzeRpK8q9
iUg5s+syGqBGnuBQTQwk4+PjFWEBr7igRaE885LbhetMw2Sq1PRyKg35NsKGRwjZEARRoB+Kh9Sp
tbyU0SUDw9MYfJzmC3vXYS9UmsiXjfjhv1e1dfsp1gq1vOwgky/i8UrkANkO/q1O3MH1VQAMDOL/
YIJgOLsNSLCC6t52t35dp9Z0kj7+tnjfhnuH64S5Zt+T7+GpQpkuqOeSYsTw/1U8BBrPO/I6HRPU
T1+14NmGB8QO5j6oEByUvasoF3eQga5vyTjTY4/ZIvqwlU2V5cSTRoEMTPeKp5pqHJ3ecWbWZL5y
SbtRodKCZ+w4mbWuHMl8ktbdEbXnDyDmA9I7jW3F5nWODb6LGeUGsB1uz/1A4NMnDEUBgUlp6xYK
Oh8rHecU/tI9mmyG5IvQAvrScVdlmaraKcWPJh0SmH7SE+/5zV7w9J2LYwG/UBr48JkCxQbJBYkM
KuC1oDf7IwxI7ofcSLmRGAzx7IGpNUFIhYx/Vwt0ct/KkWQdtPphDeKrukP2uffEozLvNso9/dYP
hQxyfyov1OrMf7feqbpC3f62wYwX65qgQDNH+mk9PyFx865/mp2whVZVcFNkHuLEbeCRCWBhluwi
2xzIQneLC5kolQHesDVnH20+lfNgtGlbnqmGLlDKYYBsEkS3B01Zku5wQj3LOfwUm76O2CDfphZv
sDuWf6mZOH61GmZmgQPFPY5VUsMtuaW3cbCTv/NrcM2ePt1ZwWlbdtGTtK/UgrDhptRaQDttnpdN
ZDfAiczUymF257O2oR1rd3ILYer88kISbxRdQh4VUBxPLcDPm5M/TGCHlnSL/p5xCE76kNt/adz5
O0boNvqoiddwXrvUmtjbScMehkzkjz5Qh+7FBbcZ1A2zPyyvuraE8sll+oG/mnWXdMcuNLrj08ma
j1m3RO7R1SWtIDqTan9oFZ7WJttDNOWM/4d63gAkjF/JyM+GnQXpZhta5fklYldZii+ssbuIhHN/
OneLl+BpVwq3z/LxdklN9YmSmu+tljCWaE50uKeal8HhDXrbfIV/0qWMMiHYo9TjUJ4D+KOkil01
gpdctPl0YbaEoVUaqlqptU6G4gmnrW4f4tSBC6Vr4AoiZ5OKOg9yzMnb506R/XH6JnwJyTitTHo+
SLKEnK7mZjWxdQqpH16cYrLbV8DKN2swsja46b6654xvvGtBQVxRxb3sEODgM/kmFCB9YeZtIEgl
R90ZGSo3f5f7b69cvZU74lnc1DYX66IS6yptOVMIHTZCfmU8s2Polgo32hFTAZoOmWzk/or/O2i9
VpOZaj7cgdE0JH8qewnKMV25q9MMlt8jFemEjNhacbGdBQXKazWe6TinPoLSnYlsA7qdXalgFOfJ
6m/2COB0FSLdhd9yJl5rVCuXSvuK7MwKd5cCiEt943ddJ05S7Ppo9UobdliQled0x7FfZ64l9cT3
8gYwUizVq9pbtx2Bv2DmoPSx/245z7z4r0YJuJMrpnsOtGszvdlTq9Y5MoIXsc7amYnrzUiu3qCe
bVFwFETnt6YfOwS14TiTmB/lMJo0XKPR7Rd58xuHhBgWYD0VsDuKVJ+vlbA3ZkXtBzYaYIBytHaW
aJ2azkR8+estIJnzzY3xtjU5NJea9Lfex2SvxeA87oY6Cikm5iV2PTvQQ4tAgFtE8t07qx86rs6t
hf08uoXDr7MOXmy84Ag9pB+Pi6cLEejkKMkARG/Cfm6X6eNIyFsf8G9czQaOfNXmX3ylXW5XaDQd
nCvn99rPbo2Er/vVQZ9YYqb/mhEr01kxdOXEfJBK8loriSI7dbEcqVgGTElr20+edaPFjYPUWCHd
XJKCptG7TcQ66m1jooOmcqu5DrFT9e6itQjbvBuE8gNR6ca2bI+zSessrcEGvr3HcABoEXXUpn1a
MrjaqORLxBi705TgXDfl+1cwVdmaWUV0DXQYqVPSFnHg4+rHEhhIrtXNf0awCC6+vUmX2bvD5CEU
gAApz6lA2kcpLaa+PBRLuHk32AovESKrkjB+kwMpYA7KV7/RQKxXGvPM0ABuz1w7qtOV9Hd8HR4y
wyikMzjyM+Ssh1Lg6+PupwUaSfDT9DU0byvPRyHAVoU7LGCdZncr8kterfwHpYCQCeudwMpTHK9W
zEqclc4OVtkYJoSPKljGCVU59qhkEv9Jl6Dh01MotsAsNGynm6cjRv4+m3dM62brL7p8Oy2tXuVL
FgS4Em3ZU0+5Lm/X8rH/NPMK2uY+NapCT84KBoV58etZyJoS0ai1dHN01aQH1Dn+NkaYVxo7a2h+
5j4/5kcuQuwL3zD1jyojgDp8m+Dbq5a9e2rtKsh3ehOEnLay6Dg6TyHSJyZdw/9WYp8u57TwQAoK
4xgRKNbX8r+XPmmu9NCk/Erd5AUvtpecmx8GR+KbKN/6G672SXj8SyFfkenQ0DPjm7y+ukY2Tg/n
8+vZhgheovMEeY/w0HCQJ6ktUOMIma2ejXG1Mk3zKrIpLvbqpGJWIn7nIk9LO0cAyPtEHgqGLxS3
N/qy9y7RDf872/QQRjtD3C/Qe4u2PvVXE/f3XLPmSRDdgagWS9rS4n8YAZHdOwUN+ndyaMw/nb+j
cDGqdHS7vej7RVMTDdlqY38eVvlgTOV+TI6tYVXEEO6+qhBqU/3+yNxDZRlPJdnz8wSB9MbLacnC
dgD+U6j4oF/6WXbLjXouK5j9fduIOQHZs5a9phs27BlWLAGrYTNgsd7+GGJ4sho9xdcACIH//y73
+EbfLzDu9SRTR142ssidrkiBhNAnaEagrl2T2sNA4ujDuBcIPmpvx2udwYGCU00DcW/3QYCYxm1o
t3O3JfPG/iUR9N76oRhJpX02DkaoJKlaO0u61fb/wfjsZNc04EGxg8hkMLYXmug2hUF4i20P0NnI
5LuQWZqSTyvwSZzRopckWmHAB6Ow6asf5zLO/OEORjn1FJts+fsdWhGbm5likK4AHiRyzLYs+lMD
U3ULelG2AcDeymutpNxpOTZdjBIc1c0wjbuaOLJKGNnpnecVbIIVoV8hW5HNLj66ScCENKvLBLKg
QO86WQgKPWa09dP8ZLPIj0OGp7tZJ6YcZrAwq2v7tt8De4e80kVNTxEEvuDZaVa8/IyuvBh6pfst
miVhBrGkL0TvuWP0pzwT9IB/uL3oMvYB+OTHYp2yu8I9qeDOinGF85Mhgyj0FYy4fGd0LdIT7ffR
eMxLuiPJV9jTHPFpQW5XQHS5P7nQKrws8BRc9Kt+cV0B+GsqsiiygBFhTc2m20BgdVGxNr83AUOf
KTpikU1ZbIF93Om5+FqFiSpq2YQF1i90nsNJc9DjI/t3ZXOgGUw4DPFmCNO68tR0SMMTc1akTsl1
Xke6TEshMSFaEnnUghVoaVU+UY6/JP2Sn29/OolqJWsBs1qXxCxJmoKZxObngcKxKuZvOFZ4eO1d
o/JHRYNiKO1xy0f9swAj1SP3U5qeLlaCr388st3YDD373XZvTKpQAuRTEhYLeVrXpGFFEaKlrepT
V1jdVPGOkCm9ZCAgdnIraTCMyuIqIZGrd29z177CJaoAUL+qxxJJVctZSz8SG9W7ctfh5ZurZpmt
N0Qe0qgx8anDU7KQjM+6UKObyZMPf+EkVKFmTdOkiCAMZKDzHAl07Gab1nBNerdCPxp0A0UZGzlz
yeDYi+5QpV/9GpLLoCeM2NP3l6MFkOmnRnkujRigX5xVpt6EMqxdNFI6v8dHsVoT/kOGZLq4s1wB
95gzZw5Lbzw8lUVgW+dQ/4RQG5yf0w3YaNnZJ2NEkCxRndABg6NTCS9ZjHlcjUTuxRbA7ZcRqA6C
48LspA/ne2z4tfs6YABHPdv37LafVe1kpCuozoopqGe8q36MJCGAtQ8glm3XNgVgU1I5IKE5+tbR
SkyvjRlVlc3glP9u+HrPjPtmYiKNQMatGARwcLNTLTQAdiBqm4B28uTN1Y9mLNbe4ZIHDXtS7qKF
K6e4O1/XE+0Bf3twgwD5Lbauv2pREK0BL+FxujA49Q+JgOFrvB7H5pOpXIYMl7/9rlCi4FmiICMh
L8TT4t3nbz2jP1x4LExA1pr4atMlYAEypoA2v75ct6hFF04pEuJ4RyyOT856OuZTCdsCsoTwVI2A
X+98Qy9YCvFBua9/0oVn9Eh62qJ+4oBmUBGJX4IkNqm67fTBPGR//Q46Wu/ltU/bO3gs2iMLA0OA
yOJnjKznZB0cg11e/YFCwSPIAc4j6ccCeOlWqXJVhG5GitSx4jUGX21AigzRi4lAWueAS+LE73xY
TY6+L51wkezIJrPN+JhZaUX7pQvNf0Ir0faqYwDkeF0HQLXTyRuGtWkUyB34egljk7h43GeMd5bm
CQYAmsSQIMozP67+GKwEYZ2wjdo/HzQXH7uOwKyCyN6z4tnZrAA22No3CMwziKwvAy6e6AgPEzFt
tlNot5Qq9LgycYa2jy4B2qewbMiDjkByXLMR3ET52pVsm3zQzqiUqe5LqhxxcZcqjgFilZKczPaC
tcMKOOMwzo0ZpCfyIqBllN3cx+dFQXXjU/g5MjgZEsm+M5foWLY6dW0N8IPniOPkA/3fbV4787sw
d40cfdhPhvgnIWRt7sQlBBzXpdSB7AAD0NgdbgowBjkdkPy5cXjob11GkGu84IVYp6zoYxKQQUUr
xwIh7CH2U3UwZ4ZIXnXaYJYPLHGkag+wJnvyAumAHNVruW9FLtECMDlSNKwjgN9NJwY9XFVXnZsC
uT1hQ4v6S8yVciJVtBsQnCeZZLF1+r+8QPTF2XzVKtPFuQT3D1mFjrfYRzV4mDdq6gMiDm4+Isc0
I02HCAOKhGR5OV9TVvj4MiSDBBYIcby59cyY/mzhquOHTJJnmqxPWfmCNzJ+c3u/5jm3VZtH/13K
qcSn9RsaTRt+tWb93SsV9D4pbpQw/AsNI2OYv7sdf35tGviHFVhnRb3HUDtPRK+UwdHUhOuhWq8n
ylF3i67hAIIbb+9V/tStdvJxcrTGWb2L0XD1xJylagp+vedMhSH6ZnfvqCdPMUJVP7dvafhq6szK
Ci4tAisXK60hV4DZ7bZQ8Azc8paZz6xOvOB8qcq4th/MV3uO3fE0qt8UdGQn9A9W+xkfLdqFH0cl
YWAMhOOtL337y+2L0S3vo64Bky/+HmZBWnJC4pAj3YbBAj25uHyQD6CszazJHcwhWn/bQfcyzT9M
iofUElrjDwDh1gCKU53jI8PGE9Q1mI4NBTEH1oZ8RnVFfwQlKGP571dyFegio2DkRwfFxUG/Iq0M
4tV2qZrGprZ4tNp7AInRNC0ysAp+2q48q4lFqJG5nZ4waXGdYOnDOpbwuvodxFhjVHa9kVtotujq
vEl61+aEFLG826X06gc1Ib9niVIE8XQJtDw7ap9tv5/T8P2ePVpivv06OrWU/TOTtiOg3V8AS0yP
JioF9LJALCz+rSPX9LDw990yqiLZnEcusnw93afgxj33SsGbCHlq7Z6rb/7xPzGdgZ0djyNA6HBA
+CT2v9y/oANVKt0TkhWfqcH7IEBGA+LMrS99XqXZH+MKg1xmfx7ftGLs09FFCodyg2toO+KEXCI2
nKhbDvsCfEWtRjTa9tYPp4TYXAvghSLQsq/k2sjFF3AQ2XWfVrO7Ug8RMp8xLm8MtxZbtvNp5dwD
+/wTRGGIVLzBE5V3xqR6JjeJhqGjbK0oyS9TDvpHSqi/tnUW0dw37N2qJc7qWNue7JLZwSbHzazh
aF8q0+fvYRwBHGU+AecL0Wk1ffZTi3CLXDph+QpNuW+ZBMc0e7FFh1VQulvKggF6FFqW+hj0Xvkg
3JZWG3mxgTjeN4jYr61Kz5TSrlDxumwPEmEbjz1Q3HI5XEUu5fSQ13iLM7H5iCvPSqjZyuMXusR7
w+O038zLC7SO9VsYUn3wI9GDKLQ4q23T618rpaGTHxYJv3HjNpQFSC1tMgtcspXS7Nvexd3Bqv+5
VtnNM/IUGvwSnx39kPldYwl30FwNju+ywVKBR3xKNALHNz44qxOgdtb9BRJRDUzBUvUDo60jdavs
e8B7F/J6+wE9FWI9MfBT4ExHRqHJTQVkEuzBLny4F9wK4aO1uHW+lDANAm4EYq4GGCdcMKkmUl3Z
g90gAIAEkFlUn8Ng5HpBrayt5sC7fSC5z3RcU7Cj42TvR1lefGx2HwlikcULabXzXSykVpP14KTc
ZpxNk2nftMMlNQ3ylkzoH9xi1iJHRqullu8gaFmGBCIUA+sDuYfdPMXFHGA81hyGBXtz+N34qvKO
lG0hyP225jq0lSl0QZ1BR7Z1pDF64Nl91gMXUUTkOJYDXhCxzaJLq6Yw7ThdAGKO9s0CMPsUQk4n
or1omseHMdRB9FgTNwqzCgbbZeaqHmXOY0VQ78tFsmkDhdrYgThMS1awAABLf4AsQ8XWUqFyO4K8
XRBcVohOnTyLRuviPDsbDWTlGq4RH9Ogu/joBx2itprwsrmyEprfs2V82nUQbtYzXO6U0boclWfO
uyWNywtYIn3j+3x5CRe+YC7jxsFRddciCV92buttdtkpZaSIufyaAf2hRzapsgesNrj8w6aeHtOo
B5VGe59PEOkVJdhQmjwUPzCYs16ya96haPIhtX2iw3OUXUg4RgGbe0LNMjFlCmmK5uWCG043dmxO
1kYyYOAgVqgDrysRT8MlApZFa8CnStOp4MMFcCoDTi+Q/CKe/s90mdRZn+jBiZCnOPX1bIRH0eq5
OYyxVv6WzzQGW1W60BgjaVp7hykWcN9PMAG4XTlxnziRoFu7vuauHOT4BSMGc8bpn1jG0Sjve7wr
JbDSIfWQqUBBBhEtZRCx+mQ4aHEMgi34fKkGUTjpUDjeLm78slKl4CVPyOTHqhebtBQJWMp0J6VQ
/gMJuqguWOeuB3tDEhGlurDlAp/+DNHDxpjO5YwDfB65YRj0W6n05hpq+rdpzvwhZU3I0+hqPYPW
i53dlKyOQUrUbeZpqh7odaGz3xFclB1i9vUXXQ6mrbKZeEj9xr7pqLUeXrCFf9Bargy3WTKi+OWU
NC8Zgb9BzzJayhLQ2VQIfOiirjjT2nL8rPUPjbu+Rf1c788x+QwdvjWI8sTJAmhTIaIYXmTh3VtA
dyQWcST5xjzk5lKNfgkIsCU+MXzh/OnoBsqiLjrWznuyDoV2SZYL2TE9CfU4GZSlEo7uqMEg7u3h
nmd21JiMgtChI3q5QZlfS2So18KMgoxAAgYVXTv6VuIB7ME7SE7pgRoL/o1db/iFF7/ozNePJmhN
kJjEzPllFFIG0HpJ2lA/AXPNqXZXB8gkV2V7arV5o5pqsHaARRv+J86NlNkySEUfzHqQUmPljDkU
BYkTjtBP+zjg3PF9ebeb1BpxVQJPZK2oHNk2ZlLtixtHXSXKpMDHGV374qawjbZHlt6kthGD9C0H
IxYThzf9s2Ryrb/u+Iev3H4AdTXdUM/rf7DNT8uCT4ajzyHfqpwpL2XQyj8wuicyKhfRQ0fu2Ldp
7WDuBEK/Cok0kyLeOHrjthlCRYsua8tc1Sb8napEyfOgjVzSsDoePEpXrfqIP4ctb3GwT+mAEofb
wGr/POr2hk54S3ZWFlfDcmWjYjw2VBurGnGInPTrI0X59uAKjj6YH73TJYHgGq21/NOeedVrd2oN
EGLfzsRp1sC7JKnp3/epSuy7eGlvEafipNsTWg7YFdHoUoVdASqwk992SsWPoKMLYjdmUO084yrs
9AbXtgR56fMJKJlCfOSpy6HThoQZqZ6XkSYYh0bBOX8YrZZIyVNgv0jR79nSXXYXHphMQ2asoEcg
sPq/ssGB+hgzdt+/LV6W9EXty6n5TSWlQkQ2d01o4SPkTXtkb/CUNE8VLodSK0xUVek4d9fyvIp7
ELul4wOnJoD+7E05ZlwVCchuh1eTnp0IlTsGbrdAtlT3Ia7o+OdgMT2HFVL2s5p/lpTRVs3tcW9Y
ygFyr2kww+7e61V89XYqckW0cz/86KNWF6tl/qSBlFhsRu3MWoS45AxrbleMI8pSncOnXxXOajPK
blPSyAvPLxhC52OtMLCUbPEVqzEVH+zp/c9HufLW6tPhdNtzcpFylMdQBhHc2ZSDL90eQ44TjnCq
weNurRg+MqGavWcm79AGAC25bfM/90PDWogBzwzVpQN9HiqF8Ppr6SjklWvbEVNaDESIkcJORT4t
O+2GhPJFuH+iNKSuMuUXGIad0cTdaHinjktOde0YK4sMRIMuK7xzeldjO/5bznSinoZ0qU64akkU
zVeiJjtwYVwocWi6jbjNmF43H32tiOImGGrjgYLa0+E6XyrcmPjXNA5vB+T5A+vBVoFUfg7frm+8
OYqiz7kP7cQH0bdaAHYRREVrU6bZef9xhnacMXfky2WOYXlmXsh3Ge9Fut+CHuKx2TW0Y17ET5DZ
XKl7HqaVgUaqyTaEdpz5qr45NWRD/mZw0cDKLzFLQty/97OYhOKHqnYgPDuKlkw/W10k7eY8PzqS
ousYuopIr2NDqs82PgaTV2DpBL0Cd8/ywmwE3GrSwAAfo22pS0ANrywwYgK3dbF/JOvIYL73dPs2
JXgQrjasxUOYjdgqPu6QYU/GvunLS5kzD61VjXafKWbiG1cjw2k2OSeBZ05M4x0HwGV6lpb+3JZ2
ehZW/YXYynHzJZ+tkhIXtHVNBhto3QQPolP0rTs0tBsUp6/2+GfH++Y1PgdyrYz6GCHZl43mSFf3
ZYWphoOemIqbRUH8p70/Fa4P/WZaf92pdZJ+H3LL+zYEOo3kmeGOhEEn0Lny8fcmouQW9NVFFgKB
YZ3gmJaupJq23MYqx4c11j0B3IObQfl2eTGuUCfvEY107sYQfkcUoej2RJAfJ9qiu52UJbnHlcvg
0cD+Vph2BQpSsVo1rqd9bKrDiojEcGDw8BuYW62fVPW/OKswCgPFLzDbNn9eCriXoaEF3nzO+s38
Gcpb4K14wmkVzIvJb+z85hQlWXIEHuNAAEjfS9Vg2KFQU+6EYqvcj2pQiQtpVGvfCW0hJ4peXaAc
Nx5sh2zMJ7Sc4Tkl1tTieYPavvCwj1LjTz5D4SOTRD1BYmG+PdWooy+lmav5ihTS88/xfPEmoCxZ
XoHfTl+BKUp0aML7H87iZw8Cb3Cad+c9iHfN7csHmh48ny46ZD5fuB4XB2UJ4CAn3gI7CNmYLLPC
w2Aoijc+5thGdH/jRwpx1v/2hTuGY2iNQcNSkIS+OSREc+ngqkv8yz0UhabQ3RK8KTGEuURdNP7w
w+l/kjrI4Q/hdcwtlVMgwHu+W4SBKIbyIP6PU+NQQK5UK9snYuEt2PTUBasf/ECkSvudz6ukoRZm
pigZizMQPnwulXg40WxLz6kfQRJmsYRMxX2ACcY38pyliRwfh22gZcopZ77RNciBzEaJLJhzYmDL
Y9aQmRNrkFuMP8bEGJFdMUk3ufCJRIWNzN/p4D5P+gNX2MPV7lHqXsbCP3ggBJ1UeRUxI374bu6y
jm5+MQSurruVTAJxhcwLXtdROusJGS+yMNx8NjQXd437j9MJf64Bp3iU8M4ii82kN6h9KlRpWfdT
ffX11WTcY8kWzpMQy3oY5/xnYyupM4RYbHdn57hVMKHJTFZVmauH6ppA8eYvUVcJopkfGzuxxWOg
SpzPWTj/aR5ISHebB//t7cu7C/j3ET0+SMfPuNjnMMvvno8Oc62/tW7vDTcY+tq6VRifUc3VKYTT
4yHtaMHlFZaCyLyjLAEfVeWNGGtUzeP7u78P1/5XkOzfePgznb+rZch71ONm4UWANxUWKK5b3cpr
99lBXX0OTJKt47hYTE2c7aF6FY9Kk10CXP/ikLvmhaW4JSXRGggIw0pVBXaQ4npfvBJ7aqsPcsYc
DStTnLk9E226K4VoKvGdPAGYERAYeWKFAHTtyO2D7YV6/pjLIwxj34YYpPAmCX5lpLLXLiThHd9h
gV4EubltIk/jw0vOABfTx1fSuoDnOO6gESBWQD/eQMchP3oRMx4ZONxSGTJp4K8jpTq+jzfIegZb
ywok9VAOUDIOMA2kndxjYthU4pOxPArbHVPObfPpEI9KTLDJ9o7LO71oQCPjOifbrI02x+SvYdtj
A5ddiuePQ7CLyU0e9hgl62vZSEGc7LeBGDj1Q4JsnO/6BpgTEtcixY6KdKWddcSAuWRVugohNT7T
wmxOQuxxZ9Gtm6COzNPrMWfMHBnm7v0vl6rZt4pZwbr8iTdq9ghiaDlnIze0uezXZlr1yNThBQzm
SOQuuziaHniJM0kh+3kUsWjPCZoY7RzyTZrzTXAPI7p25HdFRhLCtZ/+vPFtTcqTe3xnrVkl7aVu
pDEPT8mliY9Go7SoTtY+kGeaPuO4P+sLI2xHZ301Yyc7PNh5/eU8dEEnbqAj1VYZlnglN07+6BHk
Joxp+ERH1jGdljAKNtBKV/CDA3V+fBEx7f48aGn8Wr3M+IA0zbYWP7mHyiIvM7nNo/hnl0osGndn
TN1kK46j7DDKErU+VdTSkrn57j4inu4XvsIEpwf3Nd5LlIz7+F4zRv4RhtdBav9gM4xlwpR2Oc2g
Z8flClYXe2HyBQTv83RnrDbGwzLNBEsJJvjVYn+4zy/cpaG5ZhAq/vJAkXejtYdFuh9P9cS8wm1z
TTDDPKmvKzWz9IIRao6ZgAEHpDj9ncDl+sKcSmDmCuffVHBTGbAkTexsby5XnWVl5KAstVAhH48X
fVa7UqvHLe7CFiCn5sk0Y8K55ZCO1lBVqg3+1oe7Dg9Ac1gsiYn5HkeOpvblNTIQmQPYez3bqXBZ
FKN103bVutjc0zk6N8sdUmWrcGQnaPYeP1dhMuVz1nOAGMZeA43RBLy0OtRuUnF4jzGYm7SQOqNd
oCXA6TXsRYQ853l1OQXwR7YA+ujzDvioO/wfAdOjXI6z7vln0gYbpMDBFaWvYeCXa7Y4EuTsRFEH
ZICrHHqT9zj4TNw+SBeoB8y8zH2H0uiJE846sjgVvelWZ60F+T1T5eakU2Pbt0HsqxKIkiVlpAOg
7omWoLey4bf6uouapHnpOAPobznxaWsg/9ccK9qRMHJTwGWZDQV0YHr6XZNb+/uO6+AUkcZTkHAN
2nTHAE0sWH1U+H1CWRc564JXsGVj6bAyTZ7bur7Lkxjx0ARSzeJV/8QAOvHJZ7fGVseAAZZeo1wZ
Jsk10zQBhGu8VlymNh8LjBSmqyJbDOuK3zDiQvMBI2hO13AM7JIPQCiPWT2x9wU3/33NXebwih0c
/dxv1+72AcG+Re3X15VZHXOmvOC6t5Y5A6PvEsAowrKedgs7ybVTPlAHTTG3lIyvM/pkpkUihJ2p
FQ+K5Kj/IR/tX8Z7SEDOLMi9zkrcd+6b1CMrmjt83VBu+HtY2N19nmIotX7x882RjNKlVBhhAd1K
3ToHNCqLv94tzz6niD+okGiljXv9DsOzmZPPEqIRYKudQ9g36zpIpQy/JOnElNDgHQEWsWSdb8Yv
3FiiKNYsniFwbtvtyUFcPWN95x6YqWbi2+XoLGlsrqlJErAhxpS24YU0tT13HJkwKnZxF2BN+CUj
PIWs5Wd8C3AsQNrH117H0OapHnRkAaSujWWjvMDTg2WHPPVKHniQuKbnwuZrmMAj1lnqZsR8qmKm
q/mLKh0p6hN/tA7WTRAVw26f2UP1DZzAl7lI9+4gVURCPZnUyMh8nhw5IaDrOHHLfGSTmheJ34JH
56ihJbuYKbtx5/noECNzoD2s73YXyfFiku4Xzl8bLiyGuvxh/9G37HAnu2Sq0XJADTA+wt3dnEN+
ivQvZUiItLBRpO8E7T/n93vm0a7POvfgA249GSUB8Nqf29ckOmYXJWbbhyS1UVx/PV6RoRpoon3z
epgBD6eZrzTiSbq5xdHfC5LGcXqxIae5kN4NVpIoN67v9VB//bDKwidiJODlM6ma2ncttz9IRtRd
KyCizHUuOFnOg5hp2ILicH+0NU2RGaTxW/BNNS7pgd5n/BPMpc0yNQKAwL9pSF+iT2/pvQbUkwjM
iklz580kZnh0T+6v4i4nQ1E4AtAMeiUpG6BfY5TEsW7/B13Idu1tcCqaA4pEJoF0NxCrD5d6//ZU
G3KczENA/5WUKsd2seHCjMH5xUAll1BGE6t4dU5aH9ZtnhsOYTJWHXBnHK14666m9T0CKwi9rAPr
Xm7SP8XAleplXQkdv8h5J+0cD0rnxIlILAHQyjkk+MXAwEwxfaKpI6RODaybwGeFbk4eMoG17pYn
k9ykw2IOGIUfr5+mi4mgXXnx9mriXQe9IdH+GU88kwXYbsXcxID3IAaJ4g12p6Xkm/0VV+T3h5bs
HbsK06cMC7gUHi3dscjUFdZUoJbf5NBzCC/m5Z91+pMqZmMLNoa6R315u0NT3p5FPnfM7WAXWaWC
8t6segOoUtOOSI0xGn+Z9AdjAmXQsM8wBAl12nIZ7YX3Xltpz8e8AIdrEpRKIdE8gkhMYCubJjpN
ah7meJJ7CPdksCcBlI3w9Eugxkbe9R9fJ4R4SPxFUgZkK8Cf1YCrspoMw1thJqoRnlmcuD5GxAdX
TYrnYdv5QrQMi3rwlveXBQix43IYKLQNB7ZyXQ3elCi0eNAqELm8emN3S+6YW1chKS3+k96/iHix
4JV0pyeAD5/XuZxzyBWewQLuIHyS7qH8VKIliNClB5uhtgC1ZL5DMGEVVho0tcckJLr6xJ+aO5Xi
LfWq8cbT6DNu3i6Nw/r9926kQq0HXyMrwI6Oc1GFrSnwnRNamzcGo/yAJyYsh0USmR4f28XXOybo
Lq1dzVR1954Wj2uT+Z5pFOMRHzUPGbbH2m/PQPOYkKPtVcNUcovjWXoJADlXAxFLamHrFuv12mFv
+1eS0fwiBFCx4hqTZxkxHC10SvArrb5UuM6KAZh/ZTSI1KgUQSLKn1ASbONLSBOa3UW1G07+s+9c
BC5QDnsD0dpWJsmtwGoo8yMzsW3wnecZ/Bt9Z/JOLquhOaXtfagFHO9/h9CB8e2/LRuQ+84ls6OV
6kG4Louwh6E2jUj9hOYi7vuVd1fBbLaPBl0zL5KHLJD8MnxHViJjulJncHREfahgfz2Mq+Dz/Fl7
KLbJlabvmjRDhQpkQuzDb9kE8Ys00L2AfyXXFv1VLSlLXhUlHZ3OluSINFRbxI3JGxbHMPwv28Lq
XdSRLCgNK+IzanqgAqzh1XD5muo6Hq58QkU91sQ34M7O7U3xZrAQFkC7i2vgA15j2WF6F79fa9vz
yEX0aEQxn2utXhWs6g4YIC6Y6rGkCU8ektPl89gy9Yv/GKOO6il+p0Dl9lJjemY1ARResLthYGDg
K+9LDVtWtzZU79cw6k6p5R2gCRf+0qpnsC14Li9yoMtRJp3pRxZmxsPoL3RK/JXNSLdMh5MK+BMD
fY/Rj/nZiAuecwqzuA2j7HBM+FlLzF1s4Z2PcuCxihSpFbGlWWthsC6CtzXLhpF9FRebyJeIX1eR
vNYUTaNxlkeBdKisvMdo05pPgPVVdXFwOdEpmCbrdfXy5I14+1dN6O5UGTZbem+sum7I5I9ThX1f
3TMEXr4u+75iM7t0l4CSoLhdS/g3YyBMAYyNXtr1MMhn+NmRed7lMkv9M/s2XP4Z59B4VMSLl0zN
k++ynZWI2yukA9Gg02gXi45wrV+8vdetC55h3x6ooDgV0OU27x4YRX6zIJbzxeev2p+1+Zvbn4+b
rAAV3FQPDqLmXoAcjux7JxR/7KyBEXN3GasNrghbxfBaTmt3alDNb/Ezyfh7AAuO6d5bFYvXzGh2
zUIPX+ngd17X3qXfwCPvKI4IxtICAwiVMrodpKH+SXK0nZcmffTryPJZbNG3M2nuGVGw/i/R5xep
jpou4HVHa8rmtG0fEJkutgWzxfXVwUQxtqinot1uPh6l+/D0cz0dfYT+LLn0BrcYx6Go/AWLMtaH
/ktLteK8Prfa9Xra5IP6gXotblgTuJ3Q+t2ryExv88lODG2tOo3BBxgVcA0gnvQdbgBYoEkTD+8n
a3DcHTiwop8qVGIy5clCGcfyCLvnl6mlM89VsI7b0Nlf0LSdo6V5bkVXwKOEEL3t5dVHJ7hxMX5Y
atOXWBgph0XDJo11vJIIzT6gJB9C24dRSQoyZjhhjBQygmzv7XGFdtLiZlXsi80vNvDawB656Y9x
slvcA90/M9Xs/s0IeCVKLpbEE5KXcFAIi937WH7DWaJfHM9hCEXfuDan46i0cJhDaw2iwdbxugS0
9dv8C+h+a8q8d9cU3m3hGCM+WmVY317c/oR6EWiPhzAfnyTxCsdUToFr7eQvrASE1MVTdiltzI/p
iithP4voU9pVEPc7LkbJoW8JGOoJhz8EAQN6n1wG5jRu1xGpQoSAf0isTHz2Iw0I+uE13vLkhUFB
S93PZGEyNJo7+qyomtsov2o25tzAJE7KR2BMZmWS0ybCfojUmeqrExz6OeR4nwCYvRH8K5yK61Kj
i3YrJzzAbQiJq8AVg0/SYIhoVDprhTX0AG1SaPLXNhvZV44CaSal+8ZhMBQ44/LyWgPrDBZT6sRR
5RjHEURpfAWXc+6D32OOdJ3lKt/kCknV6ie6MIWkdAKRmhHDkT1L+KFXeE/xA0QOcvn+0RuF3T9R
kq51c0aa3jK0Kpc23aEx2SwUJZP2q0/i/Gu85WI+GmMnE7m1t4KftCfwIblDc6EY1Kul/MflEFmq
BiqZYqlCe+lhxa/tPZTjG8IUprLeqJcvA+iSv5M51ouqo/lefDcvOcSAKSjIgfCoNMoMWPJmY3Au
k9jIAqqg4qUjiPMyRNUT3SyubnPPmZjNUTGRKWxo9H5tYX4z1VGkatsuzSO8/VhjjgpNGhJ8gjYX
6ZKmTQ6q2fy0jprhFAVpg29TcDRJNMKRCPRpbiL4KkfRX6pciycJpq6vybQDY9GOIGkhIlYoBAMF
266XftA0qx/KlNoj9+Ot3ttraz3v19ZTcwNOBiVv8VVVDpWjLosKaUbJhN8lQCRrHa1mjin/Snx8
cg7Dh9EiTdJ0BHqjElf/09777UGXK2WKpcyesaGPyygudbNeLqxuOxsfdPeG39myPGgGf7VXqJrJ
v7cvJREobFWyMBPdu2dz6xAZVMSAFr6RgNtFYEauTQNeE/0Lj7OIskVdDtKvzK71zrnyOX2KJ6es
IhMqWc0lTju/PH0RSbA/4id2txkw+izjDdC5kRDTLk5So3wk9KVnT8EouUMGHV0KFQg73kjt3EPB
m8uYM1gycjWsmG32uXClPz5hLZYDtI6YL2zki90x2wir+Z3mon0r0O1QQiD5IgQIW3TNrmTme/EA
lj5/pK8FCq4Xu3rslOFpQVj7ueDqPsIa1TDqnKgKn2zGBi77We6MiMwkewtXKfg4jZ3vCvh0V117
gX6AXGWInvYZomDNvq2WGIqmDj/wer/tjklanGpX5PKIzc3hCHZXtqrIfS6RqBlQN230dBmHUIDK
V8rAasnXxtsnjUZGgj1AFeW/CN2kjumOCbu8I2aqo5pt7FnU6CBvAJIrFsw+ODHgLZL/cqSxg1vX
jkthcBp6IW60Qo3HRtJ7VLLlJ/KVYMsuOZyxJTSfeAx2FZKjyu/K8KOg+9EeM1K9XDIYcBtfORRn
A7/DmaJ4ah+yr0xfrsR3GxASj2pHpoA4MPWk1svHJyIZS7NMCNURObjM4j/gZ+b3XmRXDdDM0Wsi
5UyfSv5wGmVfz35gbutvrAG4WaKUn7tmfVRxsQEH+YrrH27pTm4V0ng2e0rZXlHWig8ztcm0B9u6
vJB4wBjJTgB8Hn7rLZW/vr2aQ8kDcvR2g3OWLHQDMnVaNq3wDayqH7rMLTwxrGGWmZdqXnwIFfr+
qvHKbYn8Dtuq6Q3in/DqjfqHHKT7CkVy8yeesklr5hMMaCpWeM5Ur90FldKSOZn8/5bT13ZJ0IVv
hCQ8OD1T/3pbSsETUX6CxOZ6DPVUU3DgysHLHr9UkyV7lOoOhNswzJvmDXYFxV+FtwkzLTe1vBuj
KNzbrk6wWeOe02od4R5pmKgYW+RuL1LxDK7A/TqjL/Y6/5QeZfKTVHYQ1jnOP4kFJ0Qq5RGoXqIe
jVFagFHGUkUKYprWjTZeF644ZwXdX4nL06xYLb9jB6/jEQLPV/LQOYeKDheYZutcbDph6CfLTyDK
/XJmcdVpkXl7wmGiJB6F/GPXg+rrZJ3B3q+OoQbye/AEfQO3H7Wh55ZI63xGIwysrfHYm9f4Hdpm
f8G3zpgTHP7Xu7tPzxjV6cT41e/z625R68R7DM/WiQZfU+9VUDopt+GQhC3IRJb1yLH6hS8LH5dN
2/kllVuAFsV9F0SRm55fHhf18lVNT7K3khSK1qRWShWpvxDXH/uzEI7EKYUucq1dxRaKaoomeH0V
yc9DjlZXtNInYMdJjKgUeXYlYMYJHo3n7vs8ugmksz25js0UCQGpDX+LEjABFn3gZ2NQde8HmaKI
7mymEmyG/8sVABxfYrgcl1E7fyojUsxScK7a7yKV9mB3z7hK2hcMzPCs8VzReRkzSSAKXUcHv5kM
mFO9V5jTWoRomsgsG+cnFe7BE9uoFj1VkZlfdEiu7TWCr8SHFJ289Yi6VoQKbUDy0L/mUdoz5cr6
HX8zgib9ZCWpoBK0036Th1KuXBlgH7fWyYGUMmnx+Rx/q9TYXYGFzcz3pJ1QT2haQplNYUIJiyUr
u/Fg9swH6mChhR9z6MWG+HKfEMCEJsEZJSa8hloPMx+XhdMz8cLoRsoif5cS36PfnfbWw+JsmLSg
wO7Okhoo4+NDgSFjfjSZZlu1xn6y9g1XXDyxqX2mESyc0pJQamhK1HE1OLFg+5cpWTWpqjjWep8q
QIy0ZCb8YL/Os1bgVa21qMDLY7GnVc654HpBp2PEk1CMX+xfQIjbZIu3bkkR28Eyx1/ExRKa6uvE
KKxzlmL0DhQjlFIBsDH3xhPuUkcOr5gEgz34z5WBu8i/1q80WgBS5DN4XxgT7sK9A9dfH63k5ENj
63vfvnqYqXFq9QJ2t2Z6bASUPUWgz/1eQRBxj19I7XVTU54i4kLnRQf3AjFg7Se9q6ik2FoGgKwX
T9isvUJm1zTUFeekGDN/7NEdI91z6naQC3vSqfuLN4wIM3lI5GBrS8NQ1K6t5CYqIorK4vM0VZfL
MYSln9PC7qiek+7xRPfL8PaKWOm5n00lebrmpOi9xLGTdnf3YLR1NBK2gGFzRVUe9bzPu5mwaGEq
HcvRZVGWUh48CvZT1QWO0joAoPRZjEvRlD2qHZEnNN20kWkj9WD43UQAkPu/MmjzIVumBUB7Z0PU
v3yGOE70VJ3jO70gFQv/knv88uQnb4dcnSKOVWY5SngJimAWaqz5azUM2lwtyiw5E7Igh9aAOGbj
QxxSfuIKY7d4Nej9msInLkgG8pef7IAX938IVeUWotSeMC+GbD+bu3bDj7R55PizONgXX0CxgfFt
t6O9r8qQapnzZb7beiheTWRZwvvXuqBYSWYaZiK2OYCV7Pp+Fx2zsMqgFj7tKqUIa1Vyu5Ngwv05
HQIBJTEWzcbuJMw7R69If6IT+JLxGCtM08e95JUgItlqZhS8934HkbUw3AAsAJkPp2VYgumRqmFS
NKpA4Hws890654IgKvPsRwwUVVXrrw+vQl29yXGsVajFnhjiwTDw+aKlzlV5d+6vzwv47RQwrueF
gb/XuWGeTXYQ4VQg5cZrUyOgP2Rrwe2ou8qSDINIGK9IKo0IcopSlGcrhaE5A2r7gpN/3Tjuearw
cq7D7M0+dRM+Kf2geP/6Gah2CnngLTvkDsbSM8ZhjLMMv9MEONd9c7mfRrs+YZFPx7XnURabjgyM
7FMnmQ6d56lHWZiteUyL1aMfLXZq2nY1wCwgvOiGRkyhIsI5palLfGCyCWuIwB3sKFTDeQp8uLGI
CHe0Pn3wuYmE1h/9wFa2y3VXKRIKzntNc0lD+CKqWoIm00jHgVv/LC3X+v+9BcsLe3b4tNr/kAi4
UeSkh18x5cvqKf3qU3AAsHd5mMx8OKkOJ1uZqjnx46ySHktxjeww/YSSDs1dNS0bY5Co1poiC1m0
kQ1IJf1RxtgNfbYUJDWD6YNQt2/sqNhy7+6T1Vyt+dao9/+8UsrJJ+USibyhLwNspLlS3LgdWF0a
eUmE8A+8UkC5YabrZvGdJYFCCQokDqdLvfgpLS9SZFMIVAWi1heXYjO2vE9Jw5hxDXfTEsvloidG
7nd6wXn0MwGdhQAoVWMIYpGOgBVqL1CJ9f9x87jnGtb7iPxJ7REcCY6bIzlqoWW/dJ+l9itDLs4u
rT+FfsIgb5+m4THTifWQuCDdCIRxsDnm1xSqKnfNXjgbSrZeusHtlD9R9nwfjDDUUel7+oWH6fnA
b60upLCQa+67w5s3GDSV+TlXTzNimvAmf/0uHKP6sc2SkX6R9YsBnwvn0j6YYNjVGCxVz4N2SbEw
YDmgU7wHeZJo199zU2QDMDHdjupZJMJTU7hUOnUclzUHoH7+eqdWsbW1S3a9D0izero3yu/G45dz
Z6DsXqY2VakM/qMUgx+f2jFmd5SvnrfyjTAe+l1ezcyHXyFi86EMxD8fq70LZc5H5nYQh79i0frk
4lArWDr7AVwN8uPaEQlhOpzNBC1BBHsOUc/TLIf+koWsCpZ2fkptb2KpvBjHEtUhSWBrDdVc+h5I
ElrInD2s19wLalBU+HK44cTa7ZvDaYZ/tND4A1UlFwKDF6DILispTrmkeioZF9iVKpy4qGuENSy7
yYdFPMpzLMDjGE+y/gFy5GVneN+noBIKN5xeon1issC9Ur+llCtABFpXCOrMZD5AmbV2u1l7iGeN
kjNuZFZGKRIKAaunV7kORONEnw1twTSZ0CjOfHBWqd4WP53LcaTkq8A9fcuK3MNS3dAtYkr32Zeb
qPo+59pIIfFkaoDW9k3ai/9GqIvfoqU5SAtnPdlc526RwjwnqrjOa6seftVEndThoKLTqxG5FZ/R
xbabtuRKKQ1UOHTFSywheK9zo3JGZuKj9a0Lrf+TcaC0svfX7Msbri0oywzJefGrASMnqnVCfS+j
mwS/nY84J7ViA2oOGkmLjVfJf3oBMuCr/rJef+sFFfpL/5Nlvv9XbPiat8PIx15VMxr+ih12h43a
idU0Y3dZAIEW7rKImfaKOT082zZoKJ/UVuzKS3uSMN39UAPr6TuhwL/qQYj15O+Q+Kpv3k6VHtCh
ORoJEv08nsp+l66Lua4re7RrEFzalDb3qWBb+wGb3iPSkliE283l9tATMbvw7A+VikdAXCZHBsaZ
M9hMaSvXxSwwbnBNE2Or5bhQaD7cFxtxuI/dleV88/twcKernpmIgPbg+0XNbdP3ybwDUjGKyDBX
ClJAVmNjTPk/rnhAOVCTIpSj37cNBSfA5FBych8ig0JmEbRng0zgRPQ7bCGygZ7Eq9eb49BwmogK
kVlBQIDYNwIHwr88iuc2YspId5+Zv6k1HM3tb47OH1VSmssWJmZGjoXhVG9Zxe5VO3u83gKb+G32
KjT/JpsY/DaUuyUqjKQQ5YrCCoLP7l+QS7CQ/aF4JZAhWcKzt2VZT0J6B6CmsUtyLs0O++brh8sf
fWJCsNlQmcA8ZDc9pqXVKAvIlkL8y9JJgVJW5nQpN13VwakeB5WzvPHbL2bVG5plC1QDcyTlc7SC
E15/oGzMb238nLmt0JOrvGY6ZUWmhPIgvAWBWC6nVVhkGn02JdGStc22cZddFr6DA7N2kgIgkHXq
/Cwsxjg38dIrkIBnBCI5YGG9giMfqfShHhCvILkS20yogERekuGlE7WKXFzWljObiARahakyYh4t
69N3lOSz0GSkSoo05gyYi3l9qRVeVONc7sEkImKZ8RPpR5ar8l8MP+MUCdQKUfs7k1uS+08Nox2d
IWgqkT7DHULhJ4+OcjoZH6w/vlbm7FmNldnWJUsc/e8XEW8bkLqoN3nGWU1w+OXwLjZkHt7ujo4q
6eqHfbcIp9BynkD4HFLZSJJuQ4mrJFyLugGKL3mRKW0PSbURXYu/pVvwq0iYtmtNLYGX0mzSHHmJ
YpJIg/EdLqfmAZzQ1aiMcZgw64Js19tNvAAWMzGos6Rx8dcjkvriYScYMoedoy0yMjLYSVLYbOKc
jJmV/r+208JhuT7NLicj7XMRZBiHfzJ8VsejcoXVL0WCAwStI4tMsQ0MfhMSgpQ+42706uTWbEha
Fgamt3Som+PHrvvZ0XArrHjkT0gLswmVU6iH8ReQ1nmh9Sy3ik7VjsZbJhbpsi0GAScsLG4K4i5+
cXvvpa4o9BAnmtewOd0kkGm63rUiuz0nINSjtcuBPo9MNvrIaNsv3fJqXCqTzIuYCEzrtMRVRoyK
n1mdfWKUPZIKa2JohA0Mzpd3ksTbeHACiPKpVoTpCiaX4bXOgLYBTgR0w/XGMNaX01cG/Dy50vCx
1zfMA9cpUJDJRHnRV+nbWs5uIJv4i+OwxBC14Yk20+Er0rexKyDps1O+dKTEbo7MBLMPO5X7PomN
BAyjzVWDBBo4DtqWdpKIF/Ayn+jTRKvsT6AHOs2ljjGvON576TiOw4FVYldxLaYnYTE8tgAkalIE
KpdS2WVtU+2kNblMSFdjCyUpUgO+EK7Mt5NxK2LfrSQOhsu7b7vyhvi3RtPHfysuAtMlvZsNmVOm
B3gSE8IDvvBN4p9SmifH6ooZF86NLdym/0mH098L+nLAJgUVCJ+T3npJPnnGoQga7aSdg3+ZksUE
7BbBOvCDJeYcEC+TsgocMoe9q3rkn809G9plJu57StoqB0jJoiN9Kcbe2MeoVcIMf7Mfg4vQ9AbV
uIdFDj/+5eOYRmaugB/LmprNHdASg/yqjg9bWEIonHXd8zx6vL3biaQxPnlKk6b1pjqHjpeVeqko
zaoIXveWODP5xC0gs0k/fGaiXi/X3BLiZyKrIxNW86W/ykaG+miGt3cPZh1ilhuXwLx0d69iLCMj
lHZPq5XnR5aTmVZ2NaBXe2i1B06qDBgrghNAC/15iB6Or2EKRKLnkbGS2AjrWy86eKb9AtCQC+cw
MPqnKbpwf/DK02PauwJ7JK0v8JDF36+YT1rnpIli5UxZ05XXDsdmNgkLRqSC2DzDbUJCWIJY2WLT
PHEARjpwkWrbGdJwba97qdXxdaDXSf622aLCPvlXdbEQydxFkihJy/1h/0aezgFrjfEtS21UVd1S
LMWMFnk+S0c1CGUyfgqWIDX2mDfGnEl8Dzlo6VY/Ww4DZxNQPthyZ/VqM7eMb6fK3HT4HopH6sT0
q6LFP4G6BCoh+O/11DGzUVi37yP063dIJd4FfjxEU9cWUTmRVYZ+eviYzy0RDZb9DLMkQfMuNaqe
JBmxRDWFF0GiYEMxpYEUb1ln/HYGuqElDJVnIkM0sICwm4ZPNp3mE3spCSPMVQuCYFf5KQ8lUc6+
ZGUzJss2H/ve+PY8RXD0pn9rWkuoFMOA6OWXNezKvhxyfN9lKUp5MH93f6mrBh8v+U/R7M4y8ViY
DJ9zH3hbuzIUho/pcXxX9PU4WSbSptiSidSD2k41W3u/4PrxroCsDcmEJi6ELVWDX8/AWxtYfMdd
r2LOHRKd9LRoR0jmwKW8a+VKfM+ex8KBVXWBfgiMObUZCksIXblMu8LcbeEh2fkJR+U6L5f0hNic
Oo9VIGv/gxTgBJSWpnfeHg3MTGaHe02c0Gb8NXgQjuvEGG6Zvj0Hi4TRYz8ZLiSsEOR1GjYOJQsS
dQeNN2LDaU1CFh10XqoBkBz4IYISYFM5+2sVWyOldSa6kNJto96JBNItZd1+acVMKJzUsx9cOWNH
f0rOPCuD/W45a454kFa9MacGjRgyen3s/aopur+jgDm6qU4ldATxN3MEHDuk89qmC5muv9w34DPo
Pd8PkJGThietAza/TZpcUef4hlsmp2n7JVTCOJ/PK90zgwlJRjSWvG8JMJJSme0gRzvphXViJ8Y+
YhDzYJ6BfIgdPdyRbahob/xPGHLfckKgP8F7YTemup4f837iuNKs+LXU4K8qEcJJot6bWWxMQxop
ewj5S+TfMhmaZQnWYApCnyPiDghvxrg3OuS9/NkBMe+z2TuYdabYWscIbtJc0+3PusW43+0DHLVw
7fZ1sAksEp3MBC0F4najKI4xrbKSoNY86zQnHVs1FE4zJnBE1YBmxfaTEE6nx+RvAaGOpVg1hQsk
/1henLQO6DNxKMnDVFUtRrr8LHIzIqTKJ45mY7jm2TzoVEnp2ww4QPA2xTTsSfqsWKlw6k45la+W
Dw8WNVgVW3QmAZzdXuMOxAf/2wBRr0wX3vr+tBM1PlCMtVt1IeT23FU4yYnTQ6Edgyrzwf0PkMvF
HG+BLQKUv7LBik5a2w6kKqZEky6tJV9KAB36thnQ92i+JK0IfOmisvjNanNFazzSau2sqw8MCPq1
1+L6Wu9jgjBLJnS2b9jYSEE83xeRlfgAiHuUhX1kBHJKSa8QLpJj4i6+wRHnsg0lKopjz3ik+srQ
vES41XbDaaznoUG69/4LUpG/NO09JFweVwS0/DiEh3PmVniQye7RqYYpcT/O5EoueIiBdmLTTlX6
3N2Fpwszd3PwZjucUq3w4g8ZrGpF3e9ncQGyazzZdPRxRO+wJzVKRTkdK1R5AUuxSZRrBwiMm8RE
ku1cIAvvSFS50uvTOqNmxEaz6h+LTwvo8S+kpQ4NtsELFo120kyw0CUodrScl+DVqk+8hymO02/S
NXVhA9IobgLQ3rwCaOpfClYx7DgGymy2hUy8+unsVYyhVFlHQxVnciO2qPg8i6fnwi7nCM34Jud6
gj/4j5Wd5d0bw3qsgcy6Td+OwhS37a+BDCZHQcYBbKE4w5HCP40Or0A+nrSIC4W86Vxag/JrwJMe
ZSFr4o3A/JxqNG2GAy/QxkVkNkCIPvsWV6bk3aAXSSBtFLRBCmqjXrvhwy1/foObvFgAXevuHTbi
FpO9SntBWuL2UoQ6Z3z+sSFuvZuzRvCgE/YRDyqEsokInWn+GjZ2J/ojvBng8AkerHbQ0rHi2ian
q3TgFceFdU4nXNG9mjs91o47Z9xQ2akH9yI6lOxIu1hbfUVnTxLPTLKwxztERhVVmbCLYr5txbb3
5r3Y+RmI6gUcAd+EWnfGjjdjCdkZ4sqOr7Gszua1wd3ssJPAqTM3OY0sSL9zoEBghLe4mCJ4uuIp
qmDIp1V8E3upTlZt7FgN2j7uz7DotwiRo1Vv81CNxdR1Kze62OkXfu2Qqr8ynINIj+nXYN7jEEe0
FYbUZ9Hi3t1Ke/3yQVkY8cQpvxAH3gLkwOl2SeFMs0bXVErWbI+WUV7hKoW/udy0OhB/1RxtRWOp
ZKuBxR/rVkXc8MoPnrocCJMAqh5xRckh+OmULwaLYDBc1xQ7uXzv27UcyrhxS2dH+/4FHg9kVAxr
UcXXofcrfR8gkq3Y5TlwA9QIyGw6XaSg4Q8E9+EzYEIU+Pm2tIKZcWxAdwWRirSdifD6o+EqgsBg
nO8YuJB8fbV1YGbguVItx+piPQ/Ruz5/uMMfvo73MfEs9YyCwTHsSPZ81pg7ronrNlN6D2bPWOOB
VkMEXYR/UmSzwSahIq4jn8pO330+UN+0Mq5l9e2CPXPHES4euvyen6BNpL2f1PzH2InVhvXQcDCM
F+ZDEh69/TW2FJTive2e6XzwR7Qm5jWOUQNfGcNHy+CbO7Mi730lgStDVo1DBws3XdHjMt3Kmp9K
vDNBqmx27LIBGy/y2tV8sMcVpujoNA7oytm1s8ubDiyMdP2UoFs+dedGSHTy+j09OuYgJZpdbXsN
cAgX2Dyr8LQJQHIJfiX0ANQMeYokKzWTw0bRU3yrwjyY+x13bfFqfqPkLE1lA1NKjfQrXcJYkNMd
wLScb9qCHQvJPqGSZoAqUGy9M9W4zgVZy2CyKdQi3BrhSVUL6n9icihs7hj4i0hgs6H1tywngeCu
+7GBWhix8p0+sfZzBXeNyapkPqsrZbJs5tL4fx3GhdRDE7dcaoIOfcsJbRdSwM5FbJX2gNBwTRFr
66WqX1PRFcg8dSxqRJG1utHAhg5t99/U1beJVW8AIN+Cn5V/UQWKh9ozTh1GMx1viizFAAoji/XK
Tzqltcmuml/w3WGcyDOzgBKWQRKxiOuEEuJ6nF8MAO5QtX4xjnzn0FHvY1PAbxzRCvvRxzp4fv1W
74yfIWcoxAITRU0No0bSYaek67hF4P3QaCxrLzjDZ+EushC9ngFoBJrLFtkXtTTzfOpQPCMxoZbt
z1InCjTI4gOW86oYTE/raYWaRCXUxBUpJ1nK43lEQkk+IqLoQQpDHvQcX3yqSrZHEXYkiZJlo7Na
Anb6nZAW+S169AAsHqsGTS0fritp6I3TCnD6FuFewMDmZdBQR3jTPhGxKPgkO7ae5vqJRW7v33Oh
abQyCfQJGDqmjt06Xpiy+FV1xTWlY8hP1WCj/YJidWs6VCPpI5d/p+ZTN2GskPh2shlDaH5yneOK
BR9wxsQS4grFoh0rp5KKmZbA/h+BYhq/IYrPq9+ZtEP9Mr/2f3MsSZmB7vxczmOYYoe2yHrTLOqD
GfJUCb+quBImjnanTq5YCm6hdOZ30HSDlcHgspQ1zyRPX9RMCUS5KGRNs15m53sybuzlu2yCrOZg
oQQHdQOLX5zdOZ1mzf+zfVzcBUspV/xWz7YN4gOC/VXsVJSbHMiG7F3/M/MpfaOBGDbPlFa22icu
p5utQsIonS9nkfVNBUaYQ56AARUh22HVwkHXtgWnzlJAzNuB5zJb9k52Czfbm44FOzPLH2E3WCw7
5t6hV77Ewb8PY56HDH5Ggo/ZKrn4Ll/7Gxc05HMdK4vTwyp8DCoGPTJwyqBSlO/2blVx8kDgObBc
tKqs1kbgNBBKZQVvbbod1VWp4Ng/ShxeK7Uu6iXmsqv8CFq90dMyI1gZhleWamL39QsARwjslChN
SirjWZJ2cZ9QQyJu2u43Gvmi43ODJtMWqFPQHz8URNaVCF/VCcSe4M4/KdDP3ajYU6lCHCsDTd3w
32mdJQq0MBb1XQJInVDp8QHak8eixstbqxqC4eg4QM7G9snAw33ts6n8RP48fWrBzph6A2j7Fz2U
IQ8z4Y4Ng0E4rni6jMSQ5W0B2seAQFB1z/21NnNSWb8cqGbs+zh9vweenCqsN7fexiZsW81sQJvo
cizWwI0dQaqG2kv5HQsSCoE4hrBwBvauhUr+z2CRxvchOTaXJiaR2xHkpIIRNXz1ZGDh7gWkZ78E
Rkl/al067dbUXxZ02DrSJ8vUsNebQsolZkxeP61gEzrMW5KrqvoZMOPa/BT/GHzH42oxbFDU7HkE
TDQO189UydBLD/lTMJTOH7Rp0iXLW4vr0azk8+P+DHiXq/C+jL4mH8DIfndam3vYaB5l7f5/9g+6
zLtFXpDc3ooAC0mnh/kA5p6RgTDmp8XW0p5qNZgYi6KZfg9MOs51JjsgCXpKAIpMTRAbTLagM2Rw
tfxnoNXksUNmcUNgxxOzJDP1qGqtNsrB6BbqCCabpMcw8cmOjyjC6H1CeiU9Nhd7hbLdfgZsuj/E
QgE1Rk4iWjB0+4Xk5rvIEQt/mWkVBhg7qXyce/ewCP64CBKcqRTBOjX3+jvUVehaft6IZCGZuAAA
XIzvbftCC3fc0CfXudByKWLfB0Qr4PM2sQv561VDi9agQgQbi41ajHUwPChWtSXobnuFgJZ16G6c
jiGiQee4H+MvoYaNCa7+R8CVqBa7OtnFDO2VJZrAMwIenD+B2feE+QU7V0OgTGUus0731STaIS9l
T+gTz269+78f2NENn607EIwlb9mo4AN7rskNXb9HEKSSyjvi2Pm7kw4mBklCzzMYcFTxmRlUlqEF
IWkxGjkYi6jgINPOS4+gWeqqZ48emDrhh8kLQkKrOHYcpJ1nbHNG2HmHNvvg7zlwhiX2nJZqToU4
n480XbcxHvTtbFE8mmkhioYjZnV0+IkB3vW8hgiQwEV26SH9NPGFG1gBO3NBegEKn7/Z3DAzEs3W
eW71jk8tyvE/bKyU/TTqvs/YLWBiqzYneXEaNJA0H8q2rAcr1nJ4q6Bdfgi9CMKAwQvydnxHxfK2
RVx4kjEz1eX64lkASH9ZxNrBgp8gPibjPQumyaQLdLhCz0L4EA8RHGIWwxjyYNbI/NfSVL1f+VKy
EgjDGUkyLmRG3PbbU5qZI3yZfDlFAKlcyS9CFPtylLcBxBnN3pROKR3/gKs8ivoWEnzNw5pPzZil
IMgecPuo50QTeiCuTJWbbpLkidJFFMKD3Ww/hcWAXMPGnwPxGP75w/j0fm/zbfs1IIqx2qCDKo5X
yF6Kfl1BYmFqzR/mDwbRmE1b76L6bAPNrIyl4z/5qSBmzLPqbISEjYWiLROi01kQ+msuhyjeXd/D
zZquqxRhoN6ZSG0/OzPC03TZTnXKk1L0BY6E8lie9jpIQzXP9EHsNXeKU00GT7IcG0WM43odBULH
8uKz39Ofy/qIzSaukUpXNNvXNE6SP9Mw29Pm+8ySzp8FE9Pe8bBzP5PDzA4tfBgzSfOcmUO3I0ti
8eR/9bEY9gVD6FzjCYkAQN11Extu27Bj6na1KHUifDCmC6lEbSYrDVTtjiBt5IVL4dn8sw9uKn7l
2zsz7Qb9Py22nvfp09i1IdC3rBQMiUjITAqWgcXa1tdweOAOu5wIJoZ/f6VaFPAhflOnfaUJ1Da7
Xu1baF7/ppu8Q1o5NtwZopsjlcYhjjCqu38YeVmZmJdt9n6ADy+6SyO2klaK3StoHmsJvoy727w1
s+hSrrjj8k5BypyVe0FfcW1ol1siYvfqDEIr1eg1Cp1vntQUU3DidsA3MpQKLGhC/uAxCZSLLCFF
/iXo2j5CnN8TgW/ptd+ufVbePoJXBCKfqegC0rZhnoajoKEteWaBcPUedMkuPiSv+0hlKth8+ksX
L4g5ildBVu89cC+0y7//hMlJvR0dxQkMz4+TtoKc35gjp5jDSm7ReCFX7m9guU5xUzhtKzoKzXTL
8oeNQqaCtdSCHPraMY2iRqZqfeP3kRRzyUaoGhJN78x2h7aPMGtipSsdW/rKrbGpsF/k0a1rLUYh
J+3LtA1bb/wKo2p0GWkWg2uVIDaSH0sLv7CgcqfE0lxyaPqljlRkpklGF/PyQfxNKtmtkfwBgs/5
DpU5UY8hnhIGkegVN+EjnOsXCcNPz4MNXAZ7x9c61bxVH8konhtFQ9/OJopPipk7ylsU8SwcurXO
2YSpij/5Qy20zr3gz+vO3Azvqp4pm6uPVUS8zVReFLiEKc+RWpDmADaGmJR3xLLEoNxiFTT1GiZM
x9nXuJM1F/4Q7qKgIzTAG1gwyElVFzrrDdwrLguUxnPVs0caHKIowVO2TM+63sWH7hZ9pWVdeMZR
AVR0a1AQFUWbU3oPkr3CeWMpCHPaE5MWVg34FkG93xHBeeOL9bLDkxM9v0w9ipo56fo4UxcrnhSj
N77nv8ceyL4QxPlmjlyTsvj1OQ5OSzLC50zt1qBozj/i/sE5LefLUR93ORr/eYiKCdlZCYhMTeRD
6QfQWpG64nP1p6uwkjxuTFS2cHhVQdVJbASSdG5YxybeFrpawYsQgqdCMJgow5dAlLNVStg9xoPO
v5MwXey8o/V4xWwNOL1+1g/ZMVy/577Hvw0FPS1pq7zptJy4O2fFjRcbziSYT1qWXrDbcc3x1Iwb
TIEZA5TPLcKOk9m6Ar5Q1QUXpjOdVJ7JHBMSe67Qr+rCncUiNMGC/21Dq4BwSTyVjJxQndBQLWpM
uVmL2dyEds5QaEGIfERLjMR8NVQXC6el4O27BFWKKtZGDP8qzCx+2I4tGiZBiS7btwkvkJlFeZoB
EkZ6vCngYalReIxoH90BjaFkJXC2YdhV46GkyiasVef9yrgn65/tKYLW6/8ADzHHSKlKhuT1pNep
x+cJHAeJ8Vvhj2a7SibeI6PDd0PV2+cpSYOALcAAZZy0VAoUsFek5WzXbL7g6diYRGuXJCB9tieH
LlSSGsLnUlDR4NUqrfbFz/Nks/KN73l2vfXJBitqEFZWtEJX/UNni3Dv3EtWI38IPsw3xl56qt9I
9wsOQUqakf+234oHlfgvZMHGHuLQDcWKRSQw40ZzsxJDw9nYo8jw1voxdcX9/wo0INewQFZQ4yH/
XHmpC0+15lfPPj4FK/PIRu1zf4xaV6xOlxW7rW0MyW6gAyWGgjfzwa08Qv18dFcUuXAIJqakXZ9b
pMWsfZda4HhAFyZ/qV/JvDQ3kML0HIl0GvKsC+beWRNWb68WmoFzBpbbRhsGc3KImi3apqtyz/iX
pfhYcj0lqj0/Zm2S0D/ldGuLmDVTDFBTmZOQDAGfNjat/yX3otHymtPfXrs5C22tAp35pTBOKNMR
xYN3RBwOsjr/C+HUEFGeZ0e6Rd+9Ysy7aHAmQCS1cg84f9+FoFH8ol6Sw4NmcunrmZHrMEG9/VYG
XqufI3OHah7cGlyLZNZs51If17W+khEF+i8KBqsRoQWW+uYyONyNITOlmJFQQzAK+Jl3jpOmbmqe
g8hGyx3NnuJCsiLS43fRX3tzHWjLwongTrptQcYWdLG9aXYaImhjZUjONLfGAbEk10fXpziJerGv
2PkslSEVu7uy0PtjFjSGIEY3tGqRcaelHEB9AUntus1YXCZHeIK2IiZ9/DGqKOUKApaeJVolFTV0
RS/xB7hCccRPPU0vE4qhfX+tDX7pNCeMvj0ZdyCAl1h+2MzQMTrAMSTNbc+wD996CNrq2Ci0CeE2
2tCDGqCcAJmO6SMBGrmiqWHyH1SBRC7/HTX/HabecL3O8H/pz3YzhPdsIaQA24ulLhNEJWm6cCvQ
1iidXL4F48NCB8tRoG7CqKiftOk0XMUZLdD0apW/j5zDMg/XdK72y7+2fDeg8a8bJjryTAdETK20
OJzDO+1pwyl2KFwL8IE0yWt7zdYrsTeBtnX2r6+ompiw8VgTyIHbCVkK/XVXFmzYXztZEmMOFdkA
KOyvSxoWF0XKW90AJEXF6YmWpOLD/rV0QmdxkFk/6irww3doGYaTS5mIxFPs/EeL8ZVwAcJnXOuv
4/NyLYkoTrMrZdA21xal/Yl6qFYhOs0NJJRQNGm6wWb7mWTC71ovzS61vX5nsgOM72BidYtggSqi
Kr8IFpnzvxLSvRa9LgFNKXPD8R8M7IbTl5ugdmIPXGF/LdDZC0H8l6mMsYjj8NwAT+ZBrNtCLPza
PHE/TX0QHB0Y0zTfN6NuTxCXBw09OddqMkdoj8nnrseIaPK49sPJP1XgJqs8lFNkiZCqAOtwLb0g
t8xuwJ6wHcHQScxLVMu6TdwoCQd/S0Qf3065DTl9sTgXUKmpGQnqOgwBoRv7eLaP2dUxwCVoM7QP
8kvnbqzJwHN2XXOQlmNsxpNV8A8DqdSzwhyiUkJGY+4dTcw1ydq9pa3KyGO7JxqqSqikU89/jFnO
cBxqNICIgAm3IoMQkleep1x7oeDFY4c0T8kq7n9pryap3iEWDSVMBqaTIekzVQSMOGbWdGsIUd+8
Zlfb9dbwi2MglFAaIpeCgpJZYFCvdmdGC32HqBiCeHSL9dTbnmvTjiaZy79xEf34P3g6iXDoallB
8aok8UkUxrqQRQ9rpEFoZ84o3FZZ4DfN3cTQC/GKPME4+XKOelx3DAwT8ES0cBFyNqPaHtfNmQGp
zNrtq+ZFiNJvaeFG3YyOiOUWikxLkejot1oeAHf45Ffy323Bc8vdPNp2LjVyfOoe9qXsKQ+YzIt1
JnPRAcSf3aVu/z3/iDUbFRQxKbZpltgg2h4wJjFnnrwDKPOnsolyOm+BwSfupSJZnmbeyB06qUok
P00SLvrrX2y4/37SwIACZ4CW3G/3+f+RoWUYtdcS2YLqKWXPMkr4kaSrUhmkyssSJQzE6N+5GtBJ
lKuFGdX4kOpI+Frhv+w/ZRmBSdj4WwAyECM875CjzkYwPw5kcz3oGwf7RAhUDH7iDxvQZivJGI1O
/nPCdW2d5RQXO7QAsfHoyUbUs5UFFcZ3kOj4bza8ReNswqhoGKk6exCQbqvQSwV8zqS56oYeiGSf
b8FXZKRDIMvp/n8PsCwED2lF1vVvDQxENWx7EUZZu61Zk9clEYJRFWQGeXYxNzWqmi/q7zC6niHq
2e+agwc4WuqlPe/wM0ZH/ghf8SYuL9qlVCuXxaj66sArVeXmoRNJ9SccIWaSC54psLLcAjLckklq
EYWs2iU9c/W+7XkrGSyeIfkCv9mWNUXDg1sSxro6/8hCcIypsiEQ4BkIEDgP2KlM8QnSyqAetD8w
1EjL0lHmZWuawE1ro61wLcvplfVQZ39vmlVzZ86XPU6Rc0CLQ/s5kaVI25KqxUKqf97YlLJ+KHom
8oN7UFAkYhycG2RmkdkgJ6MVng66IjaMXHbyiIWOORXUyAHWS2DTOonkWu86GHllt5QQWKhT1TCs
VX5q3zE8o5DA7A8h+93ZNkfNwGpiO7bfZmvyiWJB53RinDzR3yqSHt9stRDJi6dLsYDsMydHDRHX
Cq3vEpwYKKXVNxHaBOpafPi3dBc7oz/fAzHDEqdejAjs2l0a/4zNvyXI+K7QYMCH0cgRLzfuG2ox
3PhmiQwgr2LK9sPwNeUVuMKqN/yppihwUX/fIrd20R6IBJ7wDL+sHE+KTPU8qEqFVibr2+AbhLl2
poNlqNewY0G6DRMIl7LN8XIj7r0j5Z6LK7RVXVRqa1cZ6pLJVQgCwytS0ZHbeutN3U7Z/rK7AwBy
VCaGQgp79Y5fg5JD74ekXhKx7VfIRyVUM1qAsvePjk/HpwgkkxMFmcvtKKOjtiC4NyZrA5ary7v/
fHO8LdPr0TkUhmFhb/8zg2mMS23HGe/O2CcurKQN0GMZPwDGcsaEF7p56UYaqWs+bsHnfdAyaJPc
RdSx+MgXgjWYfeMejHfySnyPm5Rrmouf49wWivw6kWP2+G/kP7dPIF5IpdCW5JKUsY+6mh6j0HmN
CGdfu1mufHZbb2Zf65Ysil3DRpnq1f9YKl6MRw1wWXOf410pkvmO+GmMR/8UDVZy500Rw3/9jzZX
6ReLm1Kf2nqsLmWcEIuYmvhBw6rC2+/Kn5mfy8jIjRBTOc/s65NLh6fYQoU26XvJcHrCy0q2GRrI
hONWte1HmE4PfWh+0dV5TwxCqGouaFZIEKwcNholOv7zyC1h652Aufzafz8wD9J1kimKfDj5eJZv
NkVlDZL3QukZDUvRnuA6FdO4DrPQJZH39NG9d214sy2PUMilJPieafRRkLUZoKkSLt4Icsk95EMc
10ejs5q/MfnJVpOiXfPqaqgrBAvz8mjVZZqxX0bnIdbye4CqM+ws8uORWCoe5ZMVxD575S50Encz
J1vEThIQULyuTvk37bbKbSXV1mVRBJHn6fU83x2oM6Yy1i2y6z7goPsMZeriToq3nPI7X7M/H17+
LwDZkA7+pj5RQVP8vVO389MKmOHdxhaYbNd4jWgVQpjDGzSwZUXbWCoEOHX0ojOyDspPD87wK8YF
Y32tnfn80juEIfvHR/2I30arxiHqmuj9RdO2jzXXVSV/8tPDkUnPylujIXNDB2p2V55+6aCQuT+0
TVXXKtKjNCYANl99OELOhcybDKAvmVidkgo0SMLLqe+kPsuxdYgdDIr0fjfXvMYBL1U/adf8shcd
5MTlmwLzrVoD5ZM6ANGMcRiJ//aNikGMAJ8r0Km+9JLVFASBjZ9t7pGpzOFfU6jq/b0hj4P847vq
ZM6rcL9IvX1ujolEj1/u+L8hcir7fZQd06dZbxCxpY8u5BRwpQKxY+hB4qUPv6d4iztH9srfLPIz
Yda+UeiLSsKu5tYIh2Rxxz1VZTJaivzmjJSLrAN//ZQQHsHLlqjPys/ZY5muS9lHrM6kyAvZ+QCW
VirWkWoosMYHCOTGcWwLIw2JeGMuWUXzLef3bI7QHLDirFpHiSc48e0k6URUFGTx+TrvbR/UKY1l
t7VjMethF8B3l6Eb49GOthFoEDWFBPzBLCwT5tKkAFxAqcqCimlKR3WYEYeSQbgyOUQud1THqGV1
7BTj/wDvAf8WskPaqqpoRGGdQvZKcYzetWu7lsjehGk7D3WuBFgGhLasUITKA04n+i1vAqUfYNDw
T0PPPydYtwkXhMiTNd9nfL0souvppgpWlDTUc2uAH8JzcUTrrzB3dQQnqzzt22q2NRBHgFGSgUJH
AhvCIBE4NiZ1mE8iRWns66uZZT0fEcjuo8jCyQYE1Sxw2FAPCqodzNOtv49CtkfZFfFSLpNK2j/+
cM01ILVQgt2v/P/HhVwUUeBTf2WseV+7DY8SEzH+K9M671g87KV7di+dR3Q+5NrWWhGMIfsSoVg0
rtA6QWWT6m+DlAYi+bjEl8eyrZ/GjP8hMdSVVwFSkRhyStnaHMCIKC5TdVgIkD7U4D2AhaqjEwHe
4rmH+7U+jO10wAwZvzxgXEgPaYFkfmXcDoOwP3fdACIubcH8GvjeMAWhZ3NkvKw85WtrzLHY2FpF
B+uTi82a6uZ01d1ZcU9p7nW359FDPn3+mtvdvNzVRHnVD1oH/qKtLcDkpllmqPo6ZKJlSeaWpXlW
UQFOpOjNjIf6Oy35YqusqpvP6KmhjQP7kObgeZNG71aR5rOqcHEBzUym3WWzWbH/rWVDmAQPYRZt
uYyrW7kbNu/LwIWiMuRPknwOyKADFHbmjZWXG4XTE/9PpbzoKns9sPikC2I+5fzY/ws+x+E9bXvO
PjfoZL5jUF8gfp4aDWmlUVARxVs/B6I5QJLnuT+jg8370MMDZq7hRZIrxWrPLG6bauuMVN/ym+QY
Da0R6vZSiM3s8NSi/UcFtwBp1/aKfW916jyIPmvr3Cu+pwiq1Ydeut+NMGFkjYMHkxDJsiZVtsN/
UN8LHz8Kj0nu1bzfnGI6UKUWd0tfWDoUdbYB3aBmeJHnVnWSHKn8/owaAqwNSBgQQ0swwFGWcD2j
alCnYjlwadlM5FmRTSfSl9VWVifVb+W2lZF8yN0p+P0i98NpL7rnM8AdzxszrbrIMMcvqG6lx/xQ
IU5b0ijdz7XKGaPb2+SssFrNo0KY+ymHNKM5U9m+C3haURpeLbDQKlFScj1CB4mU4LBZk9Lb5ira
4oyrjMVACNu6P34P5szXyvovDGty1cO2Ju4ePwmJd0V6HN5VSr+Q+OpCv5MZwaaAC9YVhgZqbpw7
jhMC+Sz2LTwDWUGg5kgb4DgJhde7w92umG3+3CqvYY9BngXGUhcf5+QSuRa7LYh3L3XxizzxXpvg
6V9a1YLNTRMz6o3SM/TBnVh+AYk26PU+Gl9Dh4VgdFeVgNbem07M5ueh8q9KCpFc0DOWF/jgKGi1
H39ANdcVJLgSiZL4WiCB+zusBC4C36/SyQw2tKm6c+IaMqv7LFJhbzDA5FuYKR6ihDpBqDeFbYVD
/VaCAaRYWP8OX0bB5FOnSY5Fqb++rLZMPcV6HTRqwQmvKMIj3DhRJ4uBf9lV4iqaOk22RSyW33lR
jspG/yX12g+9DIbA7vTkV1iIvsyOORSx0l6XB6TyYkZmT5aXIL12pY81hASrW8w/Pe89hB0fR//6
8Edrm5O5OxumvHHQkL+uUxQ5da3bXNk6GfEQmtADL2gnnbT8ddwudionRZ/5UdZz3nNn2oER69pN
vI/Pa+4bDzPLhpBQtKOxiSrDomHYY1nWnn38gEzH8S7YLcUuZ8MkWQ+yXUJ2g2fBi3+c6fXW4Tdr
fLkyyLdwqhARR17S/KWE1ZWiPTFpw2RfJq1gCOw8kJaKXgnygbc1mfoM9eGTodU8ZdPqqDLy+91O
rbzB8+mfvHkWdQxHErMFTVZ64fvkXHuZGDg9iAc84hExc4HevxKzMHno60Pjqdwmz+r+2IoioizM
wv2fL0iQ5OJl7g5/L4dviN2yywP/RWabrpvR6k/TE7lx4MthwoSb6Ir1Yea4FFkQhSBEIN0lo/pA
txiOBHX5OBwxci7necu16Ox1MKgw0duZzvqedzC/olHUhAtCEJuQ/Wb5+qeOUBy2ah4lvf7HlT0M
BCXBfQoBwZzd+HEp71441ymC+mQaUKTEFiBoeERGdNGZ4l6RO/77NOTxosa6I/mU1WKZEGOxGNd4
uJ5Gz+9GtWXcFCncerRhhj/UfnuRbzj+O087NqgKNNNnrAPjb+q5OEEtS14hzVVFlbuOViOe+B8m
Vl6LbfNGw1QFoCgtozvReExfwza9kOo5MfvACUODoH7o/Ws9tglXeMvGsZqBV71ZnvxLPfzyItuV
7eqrokWFU8lDShVmeLgEIyYz2+pyJkJo6wqRroZvr7hyuA+tiR547f2gElhDAhyUSO0pIeGrI1di
Nhnr568TzBjlMdxVVv22PUMFuFcSodwqo/iVXWeaYxl5xEoaxV6hRvuG1t4x9j1bBRxXY9WWr2qf
nSSLVlsu9i3XW3KTjjRSyxvOoPSzcJ2+NX6Doj4wDLEndVwZSaFi8MXaV9r3jgJlyHCR7tPKVGWX
BLneQUmLIak6DZwNfpMpx1WHaSdux3efeTBVHBa3Lbs+tlRIon+T/sVCiitXBSXBEsLtbRLURTxr
33KxKoLyoJJj/jas9kg7i3qN9VCVOGhMJW+pheYCYrR3ujHmdAisVnZI47zFHICW88ZYspzRyNbo
5IhzJfdmguGoIyDSqsETj8rpXk7thWw25KARRv3DweqTA+Gv90iD3eayIqrEs1xETjBuvGipj20s
BiqOC3aN4LV1AO81RsMwe+lSl1RRHnYfYFoGlvxGTTNOzUOUghN/Flyu+1fP0eZXRw3tBzXU8mwm
ci1sNKJDVumj6g5UBBv/l/5IoPQU/JTz7ONgALr45PeAEU2scg0zVaBZcRGXSbFKFL3evMa1w1lP
R78h+tgj1y5ZO5az9PshkuNneK3eQtIHQiOvXd0lmeHScLDd/xIe3f5eEcYT5zAL6rB6SvLAL01j
EyKody2saPE1XDCkFkUwSik25ujp4JkLYCw7SbEWAUbuR6dQT96byodPcClx142Rkj7MDEX3fF/p
4tnklqMuq9rAsrrcIINpuz5fWShvB1RIvySFkzRch7D7L3FJY3MRiqN7zwpUVLUJeT/1SPe0n1A8
gureSVNKCqzThczk1AMvPxPkFFLTRKfDZ4K5dl8hiQZ6DrSHhvs14JvP8f4805T3/XAU/BHBnLyJ
M7z7w498UCmgyIc01HnBDbhRR3TMV4ud4kbULAxQoVun+KKarQHt8E4e4sEuKSkAXynOIPdFNBcM
9GtOZJ7ysZjP1IoV0S5IVCHT4aFYW8VvnphLW1CkXZIpoP/omsd4/uGQwfqdSqeEO+OYu4Uhg282
g8lBLOGywZS92ate1Epi2nMBmVO32P2A3qLm7zeOjlCuxVTw8x2uAzlp7QKEtHnz55bw2AgyADoj
H4G0oBCAH+9hRe5Bb0Tz5/V2P6ayYrRJM6PDDfJCzBd1KTJG92+MALrl5pFHxEoeGHMT1iGaYMmG
PUg6lFX/yojVnHb8hMBVBzd7M32VQY1QyVQo0KfHIfmeZPMBG+5d3SfF1noDRPugMDUI/dcXmDXk
fmIoridu0LIVFYm8nAHQrbXsjvKK5XAZmwK6ZJVXTXZU2rpRLGdyvE2wU5cZi226b561lVwpuZl/
E8wtoK2UdPl/AGA26H0eKIufTHZPKw2k2TITkDGQgQQ6+mwUE+WXGiIXPqP37z02TxpjazehHIOj
evc6iHqJJU7jJnRplF32Rl0xOxI+5/JO1tY44RFUAbOeQsD4iCrOCAmM9jkqTqWv5yffZ6M4HONC
/nnRqdttpX/HeCiQ5m6K5IGrU7oT4Q0f1eCJtW3/km/0s0dVgJelTWFFwsNjhyoUya2jo69oiKVK
gDIaIpGi78vltHxy4y7223dZuoe8bCJciWVoNdUxwt3AOscfpeCHNzegxkQBeX5jUDiZugDfKWqX
ITXtKtp3Eyz2PQo8UehJJKD+BC1uAREkbDJ8waV3rmz7hUqNm8tHxPEB9N/rtcn/2VIedys52c8s
x64nv5vB8b9+uSPbHgTEbFRBtzW9YJpEwUaQJXALf6ISp2mVPZfIHo0OkNxF3kFr9VAG/fRXtKVi
Xv+6gqX8wAZ0xY4g91264pVFLNu6L3kSEFK/TZNJVAeQv036da3LL9ARu8WxESDhb1TmibiiGjzb
Lkr+Gw/A0rXaE4hHXWFDZez9wYK9+uvG9wjtvsYTr71Ba/VHY75PKxpt0hLW2SFeodYp8qeQ9f2p
ycSKNCT2gKVYGY+72Jhy3cFm3Ij4OHfanZT5gV6zoXNy/mMqsYoH+hznN6ZwqDNg5++37M4CmEKr
NbRSxvXpAb2g7c6g+xUDMBuY2eCFGvnLcLYjkJInyxFQLJzEANzAH/wrerEMIMXWYptIExB1Dlwi
zz81cdfIobpSisImdKRTKVdLDv2d89bujKw9qSGOf0Ns8B6aZkU55ewLNp/IMvofFTgbBybi606N
sSjLW1iceFdDrokpbolFZUbOHn7QHYhoYEQxfwilwTiJpALNEWaixJZ4FaHEooAnKe5PxDx5icAq
YM4bLORfGQ9ooHg3h5AjxpC+e8G88ny/CkNizndxLZgBaGMXgyIoXYKcUs0NNVWBDFKxCfCcRed4
wTBlG+C0+7OhVi8mXaMjKS9wG+k3QABHDo7Cp5UmIM40lvjuwmGNEzeMjmnkVRAAQGP2kMHVDIhg
iAucuiGS+WInfJvyChbW+Ha+cqc/nsti68SYUPVzH89HkLFWR3YAvYXDRFstsLIpHLwXacGgJvip
V0AExq40eY1t7NVc8M3rD1mEYcPGw4qGKmxPx9Yf19R9W6Ut9V42FdZJfg9bFqW2sxGM2sM6bhJK
Ag7sCxM4gJl0XPw1Fvc8I6K4j0X4kq6MPodZTzT4P+Wb75v1ER+FnCQhTabLzjjDuEuwaYYVpZxn
MVx8uOYp+wN0NTfYBi26XK2aiyEnDakJEEaUOBFn4GztMfl9LBgb7KIPBtEr1pGAyZMssbBi0ZC7
MxPCKHcYYBGf8yJmumkSBraGxj2KP3a9sUPRdowNFIBbaWDuGfLdxd3n/XX7+ZogJKHZmSwGw0Cp
+jq9Z2AWyLSSxB4haB2PpDbNvzrzjqMDfX04Z7NoLR17uprH4gtojmFboo8wRH78gW9lCGplj9vH
HDUjuAyzwiApHZZj0xi0S3HVUifOmmaOqywa2OC574fJNa3MYGp33cgpc4qHE8uDcr1Qc0dmkHNv
CCDuRmkn0XapKvO2O7ipXT62VZegGv9pZTTLLQetyk8gI8asnaM+6z8cP9FAkIyDIOykIJqrvoam
Fe6/mhwAipxxBS8I5kkVP83CDou8piUEOilfdV5mksf5r7TvN9zv/AmQJtzqWR2p0zK4P5JnN9ka
DmkUUWpvJTSa14AyB4cx8phKx3QfxPR+mgZTXSk27hISO29WN9ZL4/8kKOzVNkUO4+9iKPFpxOph
kCIgErn/uVH4C3k3+HdD1nLzzdT2NbDM28v7mnYMBjwLEqdGSX6nrfklZZkcTTl55zuUxaFBnLL/
ZjAjvMh+VqJJ/JQTq8PYiDcEbh4XmXPLQsqrQdQc7/ev9D6gSOgjCjnKwuto32CbjISKdnbg5Npa
BPzd7JCVlNsqpEZ6V2ByTDT9smKmWmR/4Rh6TsgY7jN41fsYf1JkAABg+jZhOO1jhpM10W52ky5x
EjRlm8y0nDm+rmBjQtuYNAX6+A+Cjw+dIv+Slzmx5bz+Pq4T0pg8OcTmGCOSAMv1+8jN9vtNA3hS
qSQ5YOOSXmubSgAmfJ5mTmI4urOUEhy199LIvmNVPDRjT/gNv9AVlPdZ+SgOKZookwujZ2T0in7y
2iriHEvIoV3N7/d0EZo5QsQC+8t9kxQaZBgrbAo5qFgM7oLbrG8m/Wio/H83WKpdQfqniWsrTr8T
RVYnLKGq6Xy3kTlks+hcfCYFqMHQQcfubxREXZ9RwgqskvaecQg5+hcpGng7B4eAosTvLvJsajTC
0IUOj75V85MfHvr1v9Ro+o5ZeI/UDTSe7c1czK1aTcRWP9NzbAt6yXJ0fyBuyVS9IA8ZqIgcKv+F
KjTaj0oDTUX2gMmtuYcUmOVJGM+OLHiCSqHEt+eSSO6IAUmou1b2nAVwKIFaZVqz8LeOJ5/CyX+I
cVLyvtCOt4L6d8UtqYIXudEyosL6AAD/MfKMyGKI9n39W1r6PBJnYm8BzJ8meRuOmrIXBWTNdN/c
YUL9DJmcumv00gRXqGoRBO3bjW8JiR5p68cqDN419fkNDDU9Cqub8S5rPFKZKfa2wJ+TlWCBMg4C
YFapyOItGCQ49XC2ch9Se4A2CJttz0x85glT+pnAWTyYvJ2PmBWFG+a6vwpW51PKwjO0ZTK8DJ1l
p/otc0LIWI4Yc8piuQ//hi7lxgaXXmYe8HT5Gh/mXvRAxhL2LmQi4W48odlU54Vf1qaABagYGj/7
WHmhU34TTaNPD9sFKGg9nKBN8pythD8C2l6rFDn6k3eIzBl+IJaq7o0XTZH5eP5kukA+aJ5X2mxp
uDseLQwifQrakMVAMN5XXicJlyDs98b47hnUVECa729LTntEHykYENPe/MYYPSW7TdvcRbrjStVL
AoJQ0mc4cUCIZ5Y+bWdJ5HKGpyTIpVJIaTefgAaaUv+XQiz83v8YCjTkR20WFaelhytVl4KMrpM2
duQ8Kivsc0E2iXi6ZoEt2KkRiHe0kb8mu5Thy4AJz+WzXXivvFd0j1n/TchRzeM6r1D6WpuT9J6B
dl2BbwCZjhXZBFon3C8hboLXNDFIIexaCeW6rsGUU8iapMtfY3VQO0tscoOgwrzL2nSxL9Wwbb57
+ndknoxd6/fCrno+0e8eIsU2xvAHXLxgH15qdyi6RXOxhtJr1uHK+nMDgt3K82UOQkhHaoVl2RIC
CgoH+cAO4UuCsBIwx+37v1U7DYYcTPJKtj1xVubRkCVMt21hIP8ouo8fM+SXPdzuubLc/9AxmnEp
9NOpamOOaIh3ctWr0XEaZeU6t+wwsBbhLwMV/oyiC1mt9phhNvXvIq04ar0uNd6XgpDL8cfKAR/g
Meteuw1wXMrHwE0uU1QbeHP7OOG90B2FLOZf21kkQrxdwSINQyRIsIwYs3V27ndfWnBHUzs64/qG
LzGkq9O/1KKhfjXwC6d3+KzDA0KsgQoa/TCyilK1eQJiPwwh7/r4UjuYL1zfgZwaPb88jLbNLINZ
YcvbwLXxJzhb1Q9wO0/7dlenmzHGLsZsDhUl3TLmq0H7/S5saCL8W6FczzqK7nGC+LIVc83D1SkE
YwWTkXIupvAhMvTEcXoHIrSHZpM+3sz0zRZ0F0l9+zbnjnFRVkKkCQVJFKID9oLk+BhPZvTmhhYc
u+4lOZW7nLst21tBm4Z/SLLSzz1+ZVN1DXD2xgdm7oT8r02UUDkBLnulkgBq+sDs2kMn83sUpMSq
QAg23GonoyfDnxWSUT+u2onIuv0MkYlD9GS9tTZ88VgSw0tfi/Hs5wVpHlFEqpRSO8UW8+LH7h7q
pR1IEgdMnbA5XAmJcosqvZqMVs+/3E0JM0E8PrH2uhgfdzQMOgZJZLJQhpSl2AYgOphskiaSRF2k
fmEwXAcTHpPZfuoFfed8GLoNbDZQQegzVNSIzmo1PVMrmzCK6OcRVFwsFSYwN1vsdZfnpSSHS7vA
Evj3PIKnni+SlNkrbtuUH7VZd+rsFKl5U+OrpYPkEvX8aCjZgjmN3NRGA3R+Ons8dk4D7bb2/6gr
8P+p9aP4M0yoHIOJdyUoYysQEx6UH/8ps2mMoVmhvFzGdp47mX2+wRIjQ0bD164+fmB09Tt+3epP
9D4oV7LyspO8tMTaI1odJd+y7ZCAGLPcMxVURIZvafNQUDkOjMwmcLYpZ9qvMSrTM7T43m1gZrnD
Axm1d6FIfKpI6SjRcun/7NXaypU9OR6euox2N9ceJ375pKOTfNV0+yrStBDMUPT9FkJg5d84+b7L
qlhqPFcJDKg74pKW1IZc8VP1KT3uStRelwUymPuvcKt6vsupXCkT0VdW4eXZxym/xyNa5kBQ1wJs
P5Zn9aj0hib5cJxx6YNBRBy2Y5aJTM71kUFCj/KHiJ7e5kR8n6t1mnPfwvCF3o+L7RMYKqOtjy5D
d1cn4cevHmFVCGjRGGYF7t/TH0Zm7OqmG8Ltb9s7u+qoX0E5zAjBZVwHnot9+RtL8Mp3p8b3z/hE
+l61gO9mkuTJM+zJ1xw0fBilQJFA61QnKUROCyhufBnrZcVQzT/LMr6zsySbgJZ5rmpdpbC9y3Fl
hy8ZPgmbF4J2GFA+N89n8Tm3XgMMbS1iMEPs/8SZVoxWDIpWx3arECdt2ASlg3aoa46H9F4+rOIJ
KwBUHN9sSBbZIO9+yoqP4mmMjkkqix42IkneILs3oOYXY42gH7zQLJm+UWPSzaJT2xw0Gaioj4v2
Tdv+lZtcCgECCwniuG/Cc8S7T9k/zv0JYg/xTvCFQf4Zw6Tf8U4DNsI0DwHFFJXN9VPQ7mmleN9o
9J9wDgR2+dBSHh8ayca184+DVNVo1l26aTqDmGhp3pRNnwkE9TExEwRmt742PDweABRLuYeamLNA
U9v9WrR0uPoa5Y2x+XN99V60jNUEFZ8fjHI8zVFMs2TW9KU1mlzN5BkQ3bJ45bpVXrEeIqNyg1BY
Sf2UJRtMYUje42k3BKdNCpLeAjPeN4n5jypMa8YrIdFV9QvDX4YZyL3bEgqbVszhX/2boKx3xV3M
AGeRWy6NXYlrd7JFrciqIA7c5FFTIW4Wme3LZNr763WnLBVNo8YtJlXsXh7ve4+qa+UKmZ1URCJK
KU7/wAn8HUpQjtKiv/3SYBdz8OVOicoyrA059XlLRC9oT7X2oTMga91TqgA8U2cvgN83wF25uxew
EKlZz2Jkz1EXLaUhk35VdX+01kisTx6mBzcGqesokbHzAxbQy0tnf7ehJFNYqEBOO5WIa5FgZzUe
1E+Xh8FroGgvRzUVgnxMK49iHCumUJYg6Fyi5GqKUVKNY4g7cvExVM/zjswtGPJKPfEE312Nmo/B
HFAuK+gaieCkK28uisd5VGRLIiZThYs54YFh9mfIKoLH1/gcLB1o+tauCJIfxlIcaJai0s8Lntx/
zvNLscKOBZa2T+D5bEpfKc2LvguaYNrwjzB4EN5jTNeIchdevS6Mg+DEeNPHyFaUnFhKPaTTD15v
B/KBOFagOxLGKeT0bp37uUXBP7utdUOUclMqTjINCMXnHrg+psBFWCju768A+UfeSSmfB8Z+JuO6
LIoxgECO7jjQsJcVwuicMU8GpVdezSh+GZwfuKk/b+o+FcezUNgjceO2Xd9qCqfb1ckagGmFdUmr
Tddo1ZKc6aHL0xpJyBO0/bJ2+lzGb/ALiUp1iVFQ2UZ8fHvW6dzyoC3qumDyS1fSoTFp8VituVYh
SIyWgszEklx8MROKZ3342jnAeqDw1STDoDZY/j3Aj4ZQtiJVd2KGkKviCbQJOQXMoUCxl5zl+fDM
g70nrNtk8K7RFhKPQ2HFeN/iD1bN/46QEMkc2f7EgrajHaWJwTsCKVXq3Dim7PdxLVU78pjxqwtW
mj/XZi34pjlYo9qxDU9c/M0cj6Cw0zmHM6ILJlJxFjowb+jGgCVuo/UTTbl/FB1ntnthLphO1Jy0
NR2SIao9FoQcekf5sOH1Uv9TsL+mfaTIrh3I3eiKfLCG0JpDV46qUvdnqXzQTGNaAcagZviyiJM5
LuAlQu9/nlexIqxX9a3SkQymYyASdvCENyvYeP9/SNatJ8qPHG6h7pcaa7SgrK3ze8ZcbdWjcMmk
MkTKxCyz8kcePejjTiGCklaNiHa11DzA7w6IK5ZRHUhTsNfnw5/q5Ay7TCLQt+jEG60+V8kiEQUh
4MHJGi2B83YhDe59yMmHqL502IgvqFYIiSRVyiF7J8V13LSSLVELzu0oFJKDBhmeRka8NoQHLypG
JS4QS7Itc8eCi/IKrCWzB37s5lheAQeQU545BJ16bH2JHulNCNnIM5gepaOrLK3ZjkQZ7xKzPZwh
wxHMiVOMs02DotOeGtfc4ryhnEcXQPnppEaP81xrt2Xu3Xxt272LOIPeJ0gzLFqFsYAnW+Be9izU
C4uFiTTbnzYdeKMhYBTHCOTGAA+TU4xP1af5ewQBUdrgbwdMbtRZZ93jJwWj+PZktgMgfCE50dao
zlPs0jkd23kA6/f5U7HC8Ij7WIRQBH8I62LIK2H679PMStX7LNA7l1XrNepzHTSVunxhIw14T0yY
S/DSHya4IQhsxKA9irPOl1nnfoZT6duh92P7NLpgIVGW30xjjgK03e/6jd3ZWBqEWFCx+140/1P2
fb8vP06ZlorDEvItOSSr8L9jbnOF1G7Is31C+0mS24HaFDVpIBSIn6y3kD1972TDDoHSY+xsJe3D
SkC20RFTMo+P0PkUZkOoo2/J5CFk2i+m2xg+1lhWbd/a0FD0u38U0Qy3yfoNzQyLH5cBfIHlo513
/57S5zZRsf3o4cRHHZCIxsASenLlvZ9jKhE7u2w/k3i0NdmQnucqB2jSXsXx3acM5VoSlNdzG123
OcZBSVdXyKuFCE6/BZ3lFHCsFIkRfkSX8IPdaVpDRBJ5r9T/tTKsj5bZHdM9lr0xcpvMFTYbws4I
ZLK2eGZ41pBNqa0h8PVPoYWJVAQMn9idQPWD+L48KFlpa2caKmsxR61V8JayWEfWEzxNMj28lUaq
Asn6JcUS52vlLEjeGhzA0gApr4iA8lUt6mnd9Iu1nvvMNbdgw3BDcrOUE02CgpfSF0dOI7crnLu/
dys9vC86i/l90JAJNnCT6UdAw0I/rHp0QQJGzDfWb+worL7nRdi3g2M8PrQfRsnl9w0i2Gpy9xmm
R8soir1syVUlxA9zmWIi+Qb6oCL7z6QsoWvEhMD10eA5e5bzpwDudHepMXxJrJwtdOVH07jlLrNS
r1yidlPZjOOXazguQjD0xh+exCAZF+53FET32HfI/78H+BI2F16Ad46ihz3HpzeOx+ZsyOFR0nMy
1VPoWICZGN2ZfW31r/MEy/CCBF53prsCIwtf3HplCxjud8POSi5nbCcjKNbeM1LBWYQaVuZGmpJj
34nlaBk9VWEqgNZuXVR7AnYA74mgDyfTvdM1jm6759Vm8V+v/oijZd5VGTD5gfLSHSPTG5twyVhu
ldfsdLiQy8bO8oULLVsCRAcuNNFsyoMiQgYkFfapEEepWjQMp6Q6Ycp5ZPfHmRm88/F7hn9Ev2S8
29w4rYev4Vf7UEenGasvG3EhlXP61h9QG8WXiVF4MO5N9KnNUzafLA6uy3qxP+xw7uOAOQlXiu1o
DkF9sS6Lt9FC7GNO/BddWagrOdORni5Oz8a3dfnmOx48+Tl/TbNp7oo10c2d4O5fR6pzh85BKLLe
y+JhjWjIQi9MaC4baxuysxZilhx6xazW9qMTm3+sOggTcl9Af6f/QfSGTRdZnZ0RDoW2MF4DJI26
tO1E/0H6k1qezV7ypANnQTQLlZk7OaJZLddhsWzgzOlN3WL7zLqgGZ0Qyf7TeG7uEpPe+7Z7ioFW
WLnY3DyFN59AitAEhoyoNIhnLBj7acPMHAaJCKr7lFMHhmU9nd4HU5MMCrb1jVOtMZrEQp6JldVH
kST1ZJ1wG1dwH/4TWdbXDCkobYh6sHS5xHDfxn8fRZVsPox0xWIjfPHty7w6z8sviBo2JDkCmuw4
n4BNgvbP8mrM1c7tiLUBSrdGAK3Lq/uFL4MPd2rjbvxCgybBD5z/EkNwpeS/r+hshAM0RYaUIAzc
V0VWy6hN1Id6Equ0KzLILIJGs6JkO9de15z2rPxQ/Ihg8cj431TmDJh2zvFyLtqW0Yn9Ddb8sMnR
LNJv0Yhm38lhgnRHgowRGqUk/UfP2ZSKWFPvvkW0Es1sEhR73b4PKNv2QsC8Ixd1s1TztbDC/f7K
pp0glZGBUIzaFgN5yAoccLLUPnd/HXe9oDs36Hd2MmyGJXVUT7T/ayyJZ7D8gOT5EBVOoLcRT4cL
TbfX0i7/rDRM8RKM0cHN3sD1GvLP++T9M4dA30/URVqMTwfL3fWMTejO5G+a07/9Ag+f6BY7E3rP
p1S74qedjCrHE6qLJK/80B4bOPDjZcUY3BFr+ktEwj2mYN/ZC9BseRy8EeuB+bpUlPA2h6ECgTIZ
pJnJNCpS8MGmeCGSKZ7x0ffQJe7Z2klXyevKC0usQN28QLH3I4IK7zlJv/5sI+wXb0vXRy480Jc2
RXVov34s9N77nzTvKKSCl/MZgYmZeIf9hZfx1AqNa90i1pRxFsLt4+9tYATAE0oWiEUX0CpVxAoH
YxsLJdIfGFpQlU92TXssKMe5Iw6msH+UWNkpSnneQAT9ghyEJJ/IskjqAXzI7At0I/kSZHR8ymsr
BrAFcQX+azuuzkN14AHoMHBjJZ4Es7t5ILrpTuEq6vExQq+6JP2ALyNpkKHr1Uv8Ty3HgluZICnb
LEnzc6Y5tZubyqp16vyCZD1/beVYXECSFdjY6ts3D6iiDJ5IeOgZfplpsF0Rky6lOmj35OaRi7Ps
MDh+movkhVJ2EYiuWoHoIY6u9mZA4zdddN7d88JvPkxh3bsNaE4meVwbHKwLrrtMOHa7bQg6focH
JZFoir2oryf/zQecKrrV0t4GHlIEQMF9C9DzviUdLFU3PqWk0+EADwqWSRcq6NC79+bGRGz2jpgg
JSkARrJcm8MgOI83pAz+oD3VBMpDQ1cN6KFyDc39VBPPivT0HYunzEsI8SsD2EX9dxaRW5LcGFWM
ufeg3aXEx7C6KKd5MCIc2zJRzojXwoHwS/olBvH+e6vjZ5EpqKBHpdB60IY69kwKNE80bvNlajyl
QUWSrHvAv1Z4P8XvRV3M9ry8Y7iBaagKKCpCsVvptUpmBY+tMYQ+v/VH7iSbK9hGmTv/PhXSQ66m
oDYX7EoyzgiaTrVRv3dXOKWKjzn6aD6fhaACg9ZanvncFKRVpJ3EUzD2jyJ1SZbATtcetepmsNtb
lkzaCfxOISYQZC0auIATQtR3p5Ybh472lDvzhMCwKCurhlwIR+BS/keBHw3ndm5E70k28qNNQzDu
fWu6PO3t47lUugaoEMJpLKYbasvVp/1Ks5TlrQqHekQ29ukNEIBA48mbesjLtSM9d9zZOv9lF/dO
9dhiDssDt/05JuxgR4LwkwcV040J2AV4vPBFN+g7Qa4jz/Asnrr98A6D8lw2Wz6Z/78KxqtCTGIn
4yaSM2MQSyzMDd0KJBJN8n/Sl32vkBOqP2c10aWe5X5ZgjjzSUy9fZPnKpvG7pf1C12ADwJFi0nv
J/MoYb+MH91H/2uQIkfzi6oqpgljqnGZ+1ZjU5BaaSeyd+bc6EaFYZygMk5tCL+36mzmmbER7o2N
W4qPceaPMw71c4G6RlcCBBJzrS68DNnnDw3ZDYriY+aZG+WDnTYiZZDk6zxYAXYHWNZ8Xv4hWxCk
VYUWfHQ2/X2KmRyNyaSef/l9KvseJrsNuLesxMx6uP1yMNQyexqDhp3iqITgSdFzWmaj0UnOKVT6
EeNmxbv9dXO7G5Bxprlxi74UBtI9cIbHHKX9WFdpHVMKfEjyKEuJvCNeqUHWJdoafP6fKK/ANEiK
KT6Qvxn7OHtQSXubHeLcpVADf6xkX1vCD0MDkAyBXpkqmfn4Q1qZJexNGkNGM8/4rfLaVzBy5+ec
Jqgbk9BjEO2lSlwbyeDtoOnoj4RndzXSg77ZrBSYEIbMXv27uOTgy4xWRA3wbPjndiEU3t9e/odD
TPWON7pBa5Al2P83qHVLkapx20lyK5xfy2d6iP+pWdCetK/870dvLpfu6W8+wwi0Bgl65z6gN8bD
ES9uOkltfkxXAl3/e9BZjbFKpdCHyboHYexL64XpqvX/iTlPHLVFGezKR6RNpDEZcB0GwNSOkPJf
8340Q10k/NIqr0IN0u7pe2he8P5myajy1lUhEKkzNl1r0W33sUhwTa1ITLfL8LiO8QscBCq2maj7
IhuPvcVABIVL1QNGoP2O/CcBmOEQHgRaXt//AylzLDImGACMdLv82O7NuBXZs50ljHHFbUGsrgo2
zG6GnDoK1AMW0OHUgLVWpUaYYoEuw5BG5C7ScHz5yJM2hJnR17ekNG0nzZe2wKBOv6NONTKaNElh
uNBoyQ4+dwLHDg/3Dl0wtzhIfS/SBt9BtKZJzbjs7QK+6XOJlkRv/gfD7kt7fU1ppJRfYQqBCOgG
L86T2LIk+KhS3V3YSoUgqozgjK3gbC4dC9s9BzK1XTRR7IUhZmivVFvr5JCfV/gQ+3MpZXHHAVen
TyOCEL37QsgE82ZQQFMqu/RrcNAK8gCflA/0XOBo9vKpmO01QpKopX45DrUe6CyOpTsrD46OCu1a
6ZRcnb/JVrvj3OPXjl6f0V0GSARTbhcUYqLFc34XJ3GOvPaJBN2yuUXgCaXP7SOrUXP10mJKkm3K
xgJzyxZQYwbP2ksdyQm+cTWvMiLu3+K+PIoQ7TeK9P1QS7wwFqIEqNz5EsffM8S1pIKcTh8Y6rQk
rJqoL7Pb8M39c2LyL7tqd/bfs3eOg+KRMEDCeg63FqpZvXn0PZuYVupUJvUWmcrQV13nCYsd0/k3
aGYpioLe4W8D0Vgz70RcsQAHOm9qrX+PrKw714cdQ44xISF1amlu5sjdDNKXiXoaXHiNkgiMubaD
rg4FHMchW0Va6uHd7lfPQqmd7FruNY+ubrfxBaOCDI/dou3MySja22bUK0vKVvt0QtEM7y9rNMpr
78DNzLxF/a5kbKhH7wizwa3JbhdqWQ9LDywfkTh+e9FxEeiyS0G2/xC2GmrAZ/6i8JeOAYgnAnt2
9AwUu+UjehlZAOf4ar9Z1kiaJwgFqy6vlC5xylryF28nn3ozHMrmkqeSZboMNW6E1f+eSSMCiZSU
ufrUm2E4+kHSQ8AlFxuTf0H1ERChnevLyNuUWAtAJGpvzxzCA+KAFioD1e+emQIH6VABuPOW2dxN
WCF2M3Git3r0oy4Gjgr0IwcPXZ1b1nKooLUoLuYbZSDzCh1Jys+iCGBNNjKDscglyOSmNrMA3t8W
gUmntK/NRYP5BqYi4s+X5CSfmvM/vvFHL+jPUc+a1UFt8QecasxVBYqXuNzlVgIwox8TDwFRKGVz
5LjP2FvcJrX035x29t/POeUKsGhsh5vlXNdIs4NVsE24xGOJ94Tto4PUhOiWaDEn039WBbD9Co5Q
KllztGOa+morlYtZVKW7OnVMXEqEKepcj2sCQ1NeYjfUh4JPYZUliX75QUGXewntogmRulMihExc
mWBzjtqisI9WpCbztg5IObpG0ADFDOH3XuD7popXmhO9htNQkwUmzejQE22WneDDV41MglFzVGaC
bdYDPcybQJ0IugI5XlCTyru5Xyjq6YOvMK9I3e3S0CvXAFe9bf8K+cSxEhBiQ5dgpDUGX9AvnZg/
n56RFjTL5RrNaz4OMHQjCWm/Vwt5Xx4l5LNXUQPjEOG7Lvg4z2gG0ghHmQgjqdAIfy4HHguuHx0f
gmYMrauUPPAkbSsxSphMH2yaWnVBvynqG4uVOvTRPo/+bRNZmGoHodOICslOXWdccOu/QKYefhxE
myEmmkvidTaxuU1/mr+dxJulnuhJPNr7+VdWJIwLG6QrpCvMG+u0qx21iW4tD5C4KKiro6yNThDd
+2xG0sego79SRKWvDe59gptfzKjLa4qFrLUZ9stpcHQDsXQ2tpDvfBTKjzjMP3zG6dNpgQThmbuF
RNxYdxyTSxpBvkfVmGunJYeMll8XJdxqCvHcFg0oQ40bMgdTM23LOIsF/7LhqPO4zBb0fILaIsZ1
DqQm2g2RtIP193omYAnTd7KsQB8J9Oy7Q2n2nRk3D4SI9uo60iszwjCajmlKcyJdBCfVzir9qgEN
tdE4UsdArFwr/xvU1mSRaoRQIw7dh1y7IAspswVIosoXe+1CTglnW35nhSWLSXpy6ZSLue1vISEN
0kerHwhW5uWens6gIcvgbeI/qiHpTOkLDmeM9zbe+s7HVkTvnnSTaEq+c1jnJr9aldKcA84XxiVY
jrKPkyZ6IAu8ipnd7AJ0Be/DTNb7gQz5CP431OPrVvGyBjVruCAb5p43AhsGxJumZF8iCsHP2T1u
GhDSBQCr6Wd7Soo2Mx5k0RRlZpmStCJmht9T4p0+Lm+s1smeQAaT0rop8Cmiv7y4cccggJGE5I5m
AKd3PptF1S5S/7tuvL1Yqj+SDN7+qv1SarSCHntPu1i5D7cuYyeJKEsK5FC+TS0aBTkxl+jvDaN9
Tr2A631aWyYo849GIpSz1t1k/jO6Lx1CcvkMzf8X/MtVYGAqtEdVbxUkkMW2azI6CuA8z4BkGhyB
efo2Poem3ofYxNh+z5pbZ5qDoVF1440p6SDV7J5NV8kYbXI2OBUJRfxdE+r5mXtZpV3u9FcTCdLd
aMOdBeMs4DeB8Fb/CkzaCgRPlmu5xI2AnsAtbPsBNRIIiMpbZEHpT3aCfnfWJfmWA7CJ0ctvs7yL
/jEPCgEob3fjmlrS7Q5PdPW6Vqpu109QHXIgPsvYELvkq4uSPp20PEdMDquITrGK3L2h0/qfLS4v
9YFbnXMIgxeTgEUuZ5etTeBMsmb46PBhpqHxTwthknPwZxkEqy07oP0ycYPfjuYb0yBd9OJCWn3u
A3xfoHlYN2QCCtnxM+RgA8GEireIh+iSVL7laD+b1x/r6TxJNIQV97+tzC/vPN4tXiqFNHvaaL2+
C5NvnpPQbkchB303pcdDfag5NH7O5/WoDimSqazVEF2Favvi/r5iIiV7mar/bu52u/hzUZ7uZPJa
C9L/eT60F9Hh84l5/5pt0fTm56mDLhy0d0YM1WRsSIJCzNoeEQlvKbLdvMKGJjYO4YpjlXsrsXDY
+HkVj+89C838s0pcQCWHiis5UyQlB6mL64ZFfulRzR4r2TP5ACN2v1bTNlMVjLmwvwuSAFGGt3uv
DyapRuEl2gGeQqdlK5AiC/U8zOtAq5U1X+QcZpVeVMp1nQmIP1LtT3T2IkWQFs1J09ygXn/cN9NW
8HgtdfAELTZAXY8IXX50IqLRrDay+NRrKa7kfaxCQZsekA+QRTjCKj0Vf8SR0bgQddBOnSfKl+IU
hqQ3V3FjJ0LCaBygPEi8NKy9zv0MX+32TQyFD9GSVhHZrjwoVIWqO+0HtmK4Qg7DU/Yx0LwEK4mD
EiQIdaMZY2KkiihbJsxA4fNWFybT7UGuSwKXyoWZcuR3aTHVtE6NB99efMl3jntqCW3iKmW26nhu
EuyBq9scF7XaMK6Mzo8n+PnTYUaSYeUB8+eHN6GL1OTGd0WKu5EspL+AHGXlrYg1CcLJHh3vSMrk
ryPX3ox4m2G989IBGleUeN/Jej1vcHk0rqnB1YQYGZn9UJ6nbCTo/k5DUMfUKS6DJyXa8oB/xPsD
pWMgolfXgmYo30bxHsm4q7udu5Ox0WTj2tHOUcroG9ivMlMyC4WOgzD1pCwRsE4pymcooPT7DpGo
PdFRWeb7a4rmXZoda0pbFStPpwChqGwJkkZlhEASfc569y3SVSjARHUpZajY9cVqzCjpGKn27Osm
Cj35XfRmRF/JstOFMS6BRuyJVyvjgFLh40eTSaUA8/+eiWZWWOgqXOKz2DU6bxsa3DoqQpFY3PVX
4Q9woVInR+hucc4Wp0aNcT8do+ZVJjz6iF4K3kZ7Uks8EgFVF41Ju26K8Envs8qds9EUjhvq08Ma
HcPwf1QcBdcK9bd6UtjwEv+bC60QcWgUFn2BsAGszyqTOnEsG3209IkJrQQ7mjnpz0JLwNscqZ/7
bf6D2P6PUJ2A/mvOljvaYH6BbPOTqiYyL3RZzdU26ir35YFYjN2MLMHL5NRDbzEYf35qp+umJ1Vg
ZyjnAKmK0CvCna7zSXm6cA16I5evSwYp3Y1TshEJZazwWeBQ8SjoN9nQSXgsnlLsKKXQIuSlsWwU
StsydmusKqxo9yHuLhYDPqpYoqIU/gD3nwDxDOC53eqGVWB/RAyfMgcMzi1unQ6rynBbfHiMMTTV
V0Cw2ipNQYcc152SB25YprneYJN6pN56JK5vb84CHPATzOieTkcdz5H6iW6KXNOW67TSIs6Wq0dy
gZ38tKouxOwLnFIGWDvVqxl/TopuiKun8x0kbz4BkBZeiHhDWdpQwwfS4L/iw5HtLPN0gZxinM3q
c8rbdVYfKIkqjD0OaM9lCpdQ/3uojzlgbmF1ISxt8fyvcq3wMyMsrPnCowkhMpclMtlpllFHvCkt
1QLQ3iMbDqv550fDFPJwMzm7aWv2ynS3NbO5zmNaHWpLWQjrCjSR7012DLi7s8IhdNGPHec12doQ
Nc5HpmOLsLNrX3mHeRnAbvVV/s+OGbOirtDE7UTzicSEnaRIhpeTQ59eFKcvm41SzMCXw5v/7gNZ
jDUKMjK11eNFaZ/1dg0IfuWI4L3mK0ix1RbNzdDYKyX8vKQEY0hd7hqRILHdvNXyhaUf0+8f8xpg
l4EPU4sB9vqapV4BwpcizsqQl52A6Q3okbooEh+wGV3NPobvSDymo/6nUlo6TSJuyc8kEYPXdohh
ZXzmOvUwnqoIpPm/GVCCLCG79j+d8x5BPMG+Vke/QhqY1xJ8ZRlpHNUEa4/BAmPeiDp5Xx4UMKgY
0USj+c8twA11UUKvkLCpVmVKKqmFxz/tJKeTaw2QSp5JB5Ogsfed9amnwUFW5S0JWJX0kQ8zDhqv
0dosps1WvELFw+OyVdh/2e4jF/2S6aRxFhcXwSrzZshOeo2bOQRyqXx8LF5nnO7d8GSA90MkwFzo
BuVdFZ0Hh7pT2cj18yeZ249BFEcgiYY94WZ7M10QgEMyjwGEmeDsiChf/R2WUG01BscsYjqDjtqv
xTMceudbZ0h8Qf4kxzhPE5yggLlH+m6O6W9z0R5VWLbvjzSwdpvMQ6028pH6hPb7FAMD4h+B5QfI
/MSY7BRjAuGn3wUv01zrLikQ3oDTgT9n3Y5YsdDM1JPI1fkzGb5n3KZHXbdkIJmcpe2IedMbXMfo
RI69IcztIq69d17NpHcpZQT+S/av5tg+yNApYyKL9YQeXDw57WxW7sBERLk7tcm+Y8PzoHFltPPy
764gaT3Gu/QWwqwNBbIkDSSgie4erTXzjfrb3MjfbDRbwQCEyp8Fbie0RPqWgidVJ8Q3P4VWg/V6
Ai7evRnq+igLi7bE3cLm4YfCOMKyiE0g2sNXvTeP+WwN5tmM31Kg6JQnbIQZn1aQ/s7vaTK1fuPP
4AYUx/TsBGsMRKxrcN68zc8oEU4NsWHo+x+peOz0KbxDukXzGOYahjgK4fJOteIPi0QoLLO7gsO6
8gzwApyumxqST3cSqR1N0orpGBGoJZ8W+uvhI0W0FnQTWDyn37R3Ld6wNaX9DTLqRGB3SVg1f7K4
8Y0/MMufpiQ9ZcL2q7I23kXxu/fnVDGBro2KF2KtPxet7KjHmuHq8FHo2Z7M/WlcRsOuS3NLsITf
3+zLdFlqyH8gKj4wr4QsvAkXcsJGCPU8mYBf+HWKtenKZhpEYzPQy+87E3nXnM1ZWddllW22gcYO
hCthUUVf9nxfhJtzsBUndbeQo1iaM7S+enoWWjGQ0f3/IKdJK4Xe9lgDKXtaGYH8XWC5a0pzA2Mv
PnnzQdOn20zP4r2quA1cvFz5+5e0rl7EEelgEDI/K4ycZZt0CggRsNG+l0raBCdKmeTryDlSAwwS
Leo97yjoo9EB1z4+zNDUm/3eB0IqmI4B+wiGIX0HITdYaoZ6Ry9JN7UEjsCNRs+KI0Pt81eiBMLk
OINKOqDtpQzPs4KifIfyf9PSnJSNhw+tnP1yup5Y7hnhWxQLTrDOCOfOiR/mhZ6xQibr31kV6/u9
EFw4/Iu3YphbGDDYaiZO84HN70m7eBnGqzIyjSnZRC/4gSHiqGY8iRVuV72STPc0lo8swwmEmMfT
ONlBRPF2fvW7H4SU40mAY0HctoL6cntl8L2lD9f03IWUP0pJGB+HQAu9Z4E2Bseykt29yGO/gt+y
znlfr8xwN9kgfBQjHx6u6x0YWVsZsXDu6nARq8GTUMwCbG2XWOhYmcFgtcIaRockSzoJSG+sRMkb
yoKG3iIz2AFZJcj6IJ9t3IlRInSxLT/IOlRpZO3u2YVs9jZ3atWpG4dm+7Tlhg3OA84mcyYEwFag
1zfTfNrgTzOGiFr9UcSMeOtk8jab/iQvlh8y0tvXknOlUsqhV4tEgYyhilRDN7aPXNGURbK5pW4n
XThl2qUtFKz+c5hq+GzkQNOKw1EbyK+rnwigBpSfW78XVE42X7GsrO/J4LgJJoPlCfm1Cd8aEISk
6eqeuuIRNZLRIOwa6YkKWu3PoxW8sFUilPNJTLx+5J1316lP57zrxyeR3puixpvWeZJEsnW2U9Fk
JixT0ZT3pF43FTRSTfmOpoY8qN88r5cWc2dV4uYkm7mSeu0OVngozNAjgWWODaD/0AhrQJpvNB2a
uRIiBb2JCCEdq7yz00knW671HBTMAOLJG4kPxj6qyY6KbJANzQEY7KtfOghRREVtSsaIW8f4fnWD
B7EVphiOKU5ABBo1r1d3Jj3W+xn79PFMIadQKczAtThI8H+eHMThXNmplOSOlz/NyEPOI6nppzh4
gt6fFyLMnozQIiko8Tp9BQQbtrmApViXC4vVV2OPx+cwUNboBgYEeauKoxLzXVb1/Dr38jEa1aN6
aYl9mVsJ0VYHuuNPMdbI5EvunvZikY479ZFTyreuPQ38fV/yeVoPoT8/XVIv07+RtkTTsmCttFPz
gYgmO95eaMPim7w8MOuQ6V8jxVD2j3mA3J8yP7pzTWP5aIT8DmeNyNRsd3OV93Nd2wFbBi8eiblc
LYBeasuByGeQfzSAyiLOCXRUgpLtoZ6ouX4Qwgze+Tgt7egjkQ0AXjhv5Q8ezM6AQmggbwiLH6Mw
UdYhV1mNINWnzbP+F8srlhmMWelmff8wJGMLESgtZ5UV4wm6J/C/Ss/nXQFEimP67plZ5ISYgoVa
rrVplBGlOvaHLpT79POKzCfLcJX0EGvybFBjMaAUmQNcD38fSEvaJmqz2lnhxiNW3D0pdLhOplvs
v1s/tqD6RRKpd2jOyFy+/mT4jGkgqTlTuiyr9VpZogxQxXqAobJJwBzGtjA459N4TsOeJYK1TU2z
12XbM8FzihPfsAvClcQOQlimX1Qvua5LA8+dXqgqKM2YoCFhvwzXlGwLsxaCEbQDV+BrtksQ5U+U
+du7YZvT2BRp6czTma3f4ldqc8o/LSRlDqrb2QqzL9iZ1ZpFbkUGUYOrrL7eOzmjgkgCgfOA9RFa
QlL+y2221kxlH+rW4gh+F11s9tw5x1+syeJx0WP0WciE4SN03i5WIN1yZt/Ud6mxKmP7M7PNbHkM
ofp9fKXS46gOdo0HVr7q5xAYSO6rxEu5PvOLFB5GlOpeLDNEV3LDzpgU86IKgsNusmFe6oGUIhm9
dnzRfeq6lg1tvHcRR2kNNm5NQvlwVLHs5qROrSjqUHj0wpsyGT28ocpRWaTa37QjJV/IKNspP23d
Gh8W2m8NmtM4cjga6yWZvRf98bgj+AIkIh4yJFa7K7vXHweg6EvIg/7f4B1y3l3L22RzT1+nUvAF
GqJVQhWiBYEEtFXhRURyu35bcuJny6c0lrIl/6fYtnAfkq+nvGatTSu/Msb4KBf39hWeFlcMTPmp
qJTzwWY6KyJLLngFwv6vwLxTDtb7PvWdzn4vnKwNpl1wVW5PdaaiIwP7mi4n/pQv42WePY6ZAEoA
qI2JIVNILyKvXtE5o6VRAQugTDoyzGVcXIYJrZIPqVcC+grx0TrAI4VLCdVvfac0g0N/wGpq1bqL
jCBwiR6z0Q5axdnb3jJb8eBrgCTHquR2t0x5DQdsQWQD56qgdUWSKxjRZvoR9NBSrWPhEDJYhvB1
31K50cMFKJMcsXaQvVjH+TzUSPlviaQ3VgWIdqqDKsVu+cVLZr/t4oZlYBX2CAOtd3+Ic22CD4jH
cRqdJ4v0h2XTRlCsam09koruhJq/Y96oFN7B52YaFcaQqn+d9tgUyomLN6y7VCajsqvOzg4DsxLR
+fN/Jcogckn9tTZrMs2kQqpLQOZnLaXgV/CmD36LlHqppBTOOXgXpkaZCbpq71DGSek/f6iWkbLZ
KDNiP7YAljb85vds7Z51cNl0ubwabwCWy5xbaA6wmMIfXGGHQGhAU4elgPRYo3Xc2AZMaynnrUdw
TbA3zjLBH5l0KRz4RKzcVYPC6y1NPvJ2mSE9OycKEBt4nhNEZiUPKJELec1pyBBGsiNmKbvl/koh
EyeK/Cq6zUqd0m0cu9ORB8MHeL/tzgMZoahVDPma6bFFTye9M/KInd2hl7DQgaBO6JWaynl8V6BK
QRyxFvr2akYOl5Qx6lRt8xsHHpcISHW7ygI4h6UK5YD+ePu11cMarltqEjYgQkSnGyc/VHsRqgXS
DLczzgcLCRwObgCr96wY1aiAQ+J7OMFxrBNNisZ6psJGE7Y4SoAeLTxmq5cG4av6s+/hylMUMXAS
GacCfi/QTFTbo4TGJCV0nJYOr+yHVmQO/a0ZjI3vyT6JMe2KRs9x+E7izxhrsF//flQvbKnlzCgO
dF0AxKrUYFPmkrRdpupZtEkCpJ1fVA6QneAXlPvhSElL1qOmiUn+xgquS2IbAqNf9yM2K4nqGcrV
fopEVwHYCE7c+24uHqyQoYMlAORLhQSa2zX1XToNrc7XPmTvG8RoLzpxMb+CuTaEChsjaz0zXTXX
9BAaZ4A3kC32OUf1GNhj6iU1nmckE/g3F4n1J08/5aoopj8BndJqAVgBNCZoaa94FqNw09PSetCT
2baGIUZGfRb90M1h7jU3Kvhvynpu5Fo9olvBAPMKx+qmG4q1QWZRw92skCWq8jIy2NEEkuhIu8he
jg3CZ8voc8PtdRX6fW79//OfEkOnCQ3+hx63yc4hUmUBM7EoP+DccauD6Utx0chluImLUm+qrEWn
mo4Qp4YYnAjYIIxJYdVZ+Jo2SkvO6IPNolhDPUkcTeaYgPnBrR67iVY8GWScQk1E/8eGgRkdoSvC
foLGq9WiJWDpM3Ymw/WOPUtO84OQ19kYfQDHHZSkB9vgU0GajYayF7/1YtKt/eL17+W8IBeFCwp+
Izcmq2GPx8OtyPZHZPHF5rDdQhzPQ2M1CQghykG9r0el+GrReRvTy3pMjpo3qgTPZdri10Au4KfX
Doe+n+pt241mP1mMgo5me7nCdluy7eUAkSdKRFcV0p7my0ia9nY6kFHar1vasUcGpKeoQcMH1E4q
2TAXaB/EnlrQMd3I8b+crm/oVRXg2q3lSi7PO2m0mjKdFT4fiayO727F5ZjSZK7n3K/hSy2q+H6O
TqDnH6jt7iJJfhpuNGLbTRQvuDczh/vXLuKXoSZVBEUgC/RZP3tMWJ0HL/PQLl1srI69k/7LEPuS
0ROFjOASdj4W/l49tllOLYfUf1ggpljnsmS3u4Th659lRuWTFBZzNEXzwGpaiJGktnPTNTAOzNfT
G0ae1LEHWWbr5qcLF+fmxSEt7pKjo8Dc/13e18Nj/CYgdgbukVXreGl5iooYC0I6utyzCRltA6EG
8bJGuMuLi0kjnLay125T/Kvgj6tu2acnw8jMpD/26q6fExDL41a55a2XFIuCF9DgTMhOj3Dm0gI9
XmUqF+XoxnLgRpv5xhfmxia/HSGX3kTeee2GaFn8CSINAZVIEfVFnkhQwzAodzl1bU+DeaQVaW4/
/DiNpN87OOQUIzgGrSVGn5444EZTZwDvB/u51DMmbPhQf/jSCOg53r8vNzZuE1KqLWYh062SFUJY
CSbinlnh5uwS3GZEqggb7y9Eq8nZR4gaiIogsadm3s7ub0zimI6Ik/mHipPhbOC725YAmFLjxJSE
PjT3xhuujKw6cwJOzJHeUWC6N1I25V0DN8HxB/Jh8tDeLq5f2prcWunsT0j+jbSUXks4/BEPa8ju
KRBNBu4rutRlIM3bLzjlnxC0mOATraTZMy6kSiJqdzF3ctUwOYo30+gOFB7nwsqpa5Ccm6New4uU
ZsFHWas9s4XGQ9SJ32Xp1ulwv1OcxVJ/sj9ieUNbLGA75mOKuLmrBzsX8+3sys71she0uClMMDQn
NDTBcSflAMskLncjupBQ/KkGxmWEz8VAbagigkgz1ofRM7W1FoWClG4qYeTxld8L2/R74IGqCvTO
fgdDtGS7SpsgHxRYxAobLUqLwFfezEDJNAb6gNnoh5j3rNGzgqcMmd196d3jD6VWKEaEsqo0KJFm
cvqvowmMZ4gqze8B/rxOGrVLjUhHUp1bDMEuvEbyaD8NIZBqq4LoUcsQz9OSoZoE3taEuhYZuq7E
RFV9sZJE4A1WTza7kiLRT1ytRndQlhHO/nXT5hHmtM8vJPqot4acnlbBI4JxZNSjao63Aw1qMHWu
BLQ/133BndYSjWGv02AXka/YppL+6bNP5jhyyoowujQQQlJBVuXq0L+smmoN+gI1bryoozDvfazX
ryK+y9lDRqLtP7Antzpp9/uZaVTmZSuC26sST+KZP7b8UvD/UnYuEysCQBGe1kihpUCsn704YnlC
Gh6tFjHugm3h3IvgWkxdREpbom7qSNQUUekmw+dMNYkGUBIQF6Vu3zN5VMrz+1UUEEu1huHcW4E1
Q2R7QjGcdme7/8YY8g42pc9rrKlGJwgY3KpW6YM28qd8bLc579aPs3xAwjwXK71G+ZKyr2GrnUZl
kt8GO4fURjUwGln3hs1s+vXiNm5PQybWfL420U51+4uEJW12uua61aBGJSh1WJn8E0GvbjfeY5zt
MY174wyHM7pXgQaS1/13UNhNi6q0iH2vAqrYLlbHgfOlFlOMfNtpjKDbfq5KAGhcblKH/EjvbqaS
VgPjRwmhANwem1oCnTwf7TSSN2OElyAl3kIFZmDMkb3/gcDy4U/HrGjI4Ncg+1q1dZ9TwwFC/+aX
N8HO6rCXuPiRZfJFAoavQr4nqYUV2nejXR42L0JawP9WaKfdd2/ckyV3+U91ro+gR/YDZEnSqo7w
AKWg7PN0Bhb/uICwXA75llnqx02AeMYR07qQiArEv8po/DXYd5M3EWhy57YLEQJN9yXXH2f+ts0S
8A7UPwX8uzy3YMmFEN1IuCO84aQ0LPDzxHwezoyO3aKeJ+03RQucdsbmB26GAoX6ogv7LwoDh3vu
b4Nz7XU12NEzG9wjn4r6k3mYdlSx0ZPH06ZzsL1uMax8qdf3PgDX9ADljgETsKsEi7feoaW66THV
bq6dhgz3RCcRdCd6aE1vniunMTNR1DirIXJsUdVF8D8IiMgZvcabC5J3mdpSfD1l5jwkPreYZCeL
Q1b/LkjEI5+Yy4Yw+Wg2WMAO5iBf4rr2yZdJ204enXF6LTPjSGaAcyY88g2nR//aE6P3F2ggwIh6
bYaUStRUMADSf5Ry0a+u60ooJmfP+PbzBXMXBXcjkxbDxnBqpOIgVMhuUgxFsSz61TLX6XjUvS1R
rDCD/EbMRLusLq5m55PGqlyxFLE5hhtejKv7zMNr5jBMxBLgRuJpnR7InqS4NFibPMV1dNH1dgt+
TKidkQWLor7hxZZx2cKdlZEunn3hj9WKfC3aXVZGAtxeqFmOoAzWW3cLQjIRxjLUdLfJqS/1mRIs
HM+krs1yGpKZUSyYGa/0pqo/f0vj0NPNTEpGJxHP0OxO2IGBDW2lnTHvX4F1jlG4opU/nP65Ufhd
j129tMhMPI39PXW3n3aowPBxPewKj5fFsWQ0qfeX8hFceUFtlsNBeCq3T1IbbrCtYxtP2HVTxDos
dDABfVynaZA6dhjT2pP2LwqhflPaCjG3e0G2vh3wVlS2+kIBfk9pDKrszdzP5y0zHDsgNlWtHlMR
EHxIT5iZqmShT/Gb9cFCIqvcTtYy3fz+KPYTtvtMdnnTLNXyi7YnUeGNqRX98hNTr56DBFKgcaNE
Upqmmr6cyYlIpY/Z1moJ4sAdV3CVwuHm9+83AMIjvR2JLMjeVG6hXDzuc+WfOpus7daoa9hcmmye
pTXXeEGHfNUgn/5yj12PBdGJy5Ub0rcIKp4RmdLG6J50gsm0Bm1rcF6+fOpRpP6u98jLtoaQwTkc
dHG+MtXbtyJBOLHVlW8Oy25Lg+ZFEr/VVrMamSLpQct5BRLNAzrY0UCSUaBwe8MddRO0ZpKJlwas
To1HjhUI9d3Ynn1ylJUrIy795ye+3XA0vsQe745RFDNDGslYJ4F6Ze4ITSJKYsocqWLwO7bE0qSt
SPokQ87IIqBrk+0BIPF7xZ05OFWYHZfP4ElDcxI2vyz7wjngcTeqIYY/S3eTO4Mde5nv9CunfwE7
uk5uJyTEx7oNMYgF3G8kp/082zeBUxyJ6+XBvVhR85AondMPnWS2UVX+nVHSVAInD4FRDiAaIIcr
NG1XZ2R2NhCeDXRsDctOJi/A/+U+1YMRrydIzv1inZGyMfg0TvYo3d+1ERC9EQHodwk/2Jim98HR
sMJcBrayFUQzhL3C3ez7CuTMIbvgTz4masQcQwCrfeNth7+o2sqluIo0pCR4QS1aGzMQM1Nm3NQ9
DpsSBEzUp4pHvMXGYOwgyYs6WyAzeNOtkUgKQ21UqvCHmW8dVWyy3RGT1lihwfYWlWTQ0UMm1rWD
kTR7S5DSTc6kvbxEWVQOc68yN/muhaHQK9VcudZJ6Wkmr2jFmpsr62SvWOZYWmQhdveKigbnCrvP
IVN9VgACrtSe/pc6UwI2xOTGxmPT3/iIKMYk/YdYrMn8VrCc7uDnIAyTH1TxQS5CqR/fQG9SZtJb
P+bLR45xMTyrANrmxL180Ms4HNSgVoXFYV6bM8UazwbP+RzEyJ3mhBLTstUWB+iG4IH3FOcqRPlr
zx+8/1Wb1jIvstBr/t3SyZ2YZTWxOldFBPvnt4kIUgDPoDNCzPznjGRrXFAKKAPF5vVCDr6i0YZW
foFwZbwXzm91keXWkeQNRUhWf5bNt/YEKyH+aApnaRCo7xcJZfRK92ZqdnK7m+Q7Vnxx0lYE1k44
yvR9AElxW+i7isA6Hb/zGSOek6JQLZ2soN9xQc/QG4xuuJVq64WMnYCfkklNYlYZuESiVgj4Ddar
w/WVrZtUtvrt8Jhgv3bU29aS5oV/Lc/6IfNi1xkC1zXmpNrVHhLqErH5PkcNEMJ6ZlGGRk9IaTE7
Xd/zFC/3iH6t0sAB/Or77rlX3W7T7343hEE64KdurTIT9ErwNET5RF4DhTSd8VXicmK55+zRFFzL
HykpEOWHJiwBqNGASoogpGdQIdpvlhmPDn0DHLwpqxrIwV9JNakx1TGgIdBAyJvydssgHQLH/qnS
DEgrUGkpSXOOP+E1s3C15CeW+OQFVDALwRaeCgJluwc5no9uO7AmvajefiKIP0TqDpW16hD1UgVY
HtrcVtm4pHfcn/lrEMZVu3jJbHBeg+1uT3x2TPjvbpB1jYHPIjNFoiHDDNfmbsQftG/83DDUm4sH
/LY58aDUqJm4R+PFXF6B8Cju/aIRVWiaLqnKSUhP6eeYqbwR8+jXpRWbLEKrauMbA2kSixf/bCAB
V46JlmZqaWCH3yo2vl8PK6IlpD/PnwAXvIZwuqnfXnjIQzYD62Gm81nfN7IFtnGyEF1qZobzwGUb
l8BKEmUenleXJnDHQ+oEA1suIhK4ln8rOkOhf4KZ6aIG1zj4zI3SKxAs/Qk5bc6uwuvZYfDMoL0/
+LlEbdu27EyiIBoiAawXMVpApOSzmAKJf6s8ntXbH3YQp9V+01hYT8jQQa+1NkbVnTWFUj3rLNmu
vwqV9oRp0fr1wwyXIMJW12m+oFs9i1iWBFlKyy+1ExeNvihsi4soCjljhfuGneH0pDDG/Uyc+JkP
NcXTbUMvoEL210o5qYeGHVPqmOxlMkJFrjzL8d/zc/FC90IPoidjcbKOvNL1cOadFXqahUPQ5ERq
QJbH/k8YazsUitd/0bZtbAAoHSeGoKz/Ew6an4grdtD4LfhIOW+7sVQrnIUNb65T799No5A4TAN3
U8KQokeSliUrxVFqC3t3vhI1Y54+J8y4tSre5i2WRaPi0EISruTZGnEDvIF5U+uoodjl8+Zp9vld
UtQaoyi6w7zvlBanmMAn6ELENU+fF1sscZrqM0qTaqTxzgxcB+eu67C9xoUL3yAPVC6E220q2hLn
qFGoTbZsedJOwLWoHGyGsiSWLlPmRUxdL4nEh/F80rIi3bcatbytkzcLFawu7BwL72CBasOfklXt
f4JQF9DSjqnnXWJ78BIiHBOlr4XR7dJd3Yh0WCt4vix7IvbRahJvv7TCWnT4GlU0CQn5xhoKXykH
QT+ArGoSak5AMplIV37AescZJNzN7BKX/o71oCKZOnjWzDU82LwydW95HE3IgZjao4HbJZP4rzfO
95RBL17oNdd36ZlzbD9yhRxmS5OnMk1XJKsUe1x2NBO+u2nw03BMRkZi2Iffi46wLu0MVVBWpRiN
D/4iv73tbptZlshSB63TXudzM7o1Gce3Z+aH4ce23p1QBjyN5G6QLTcsGm5UFX0bgqeIpU5YJfgH
s1n1RGf4gIdWJLcamfEaIL+Fk2c1fK/jZc2oIdh7Vdrexk2c6d/Yfj/DGNUcjNA2+UmMGok/Ws5H
C4gYtiIMfXJCXIKvhvSwkxlk2su8jIbXsNgWjC/xYpB+gxe77PqBoW+/xHoDsgq9ZMwinImphcCc
AsmUjEN99kCtU6ux/DRXNzIbBlFcAp+XKEg2YoL/IK/uqyB8HsLs1Tg0Zz9zdXQfsRpSuM9RVSPr
KK/08ZYfL3viBJm0YJotT37EN9KLdNSPvJlTaAyuJu7fXhHdJr5JKDygm6DYRwTc/q/JaOz84OW0
k65bEtYFTxO5HT1HhdneyvjMGs+gjq66KVe921Uh2w3//2Njfq1y17Di7ZlXiSH7x4faGaBTBaOh
Mg1Cz6007X5iKyZv9PFbqx5CPZ8FrIk91G0xHI3+Wm5wQc0dLAWBGT7NzFu8viTZYN/a7BKxf1OA
Ospo0n6o+HR4y7OlxHCI09jGVX8txVB+1ioXOhkW3Mr+N07dKeKbD89ycbBmfqjm4vpr6HJuuh1p
LAEm0EHP95nx2xBajha4uoTBc6GYaK+J6VgCFGD8lnbIAQj6cJC5R1DxwuhxXl939HwKwToR96Wa
uD3Bq//djYusztBGSYLTR2mg185C43c0BsKB4lkuw4BQVIOvEuXa2K0LdmqfL3znK1rFbP6/4XXK
6c4CBg5uINtXhKdiI7LySUToKjXz6Y/FOVvFzebttqxhNxyvg0NfR0W2ennNX5iRvmx2rXOMppbm
6a/d1hTdCnV0J5HJSP1xMe/5m5zFCHpOjCoEkymnWmctBzRmRvuCTRZ2umOTD0bnShqomWiAJgw8
Zo8efgXesFLGn8EkFU9x8sFmO4tb4NQ4yT22HLyR/GhZks7x05/yFDzUGAoaRKNcpnRsyflbdrjp
6P0tcl7Iuv9YVpFteDPZ2Vm3pqbvNKBJBUd/I+q7///ZxU4avpzYBD4Y4aHttq2slOa1MJzW2OM0
DAXxnFD9W6rUfHojXYS+T+xz4nGg91SsLzbzhRlVUdIJ+e5pw9CiBw23xdOYuGTYWfPRBq1OH0fN
rHKLShp/48WmgOihnZh4gS4jJxtl8w4SP1/sGnxg4kp8aoVAgY6YOGwJezb6HQ/aM0jiE9rrdeYA
WjhxuBl4XxCyqorPQK3DLYZmr+3XYAeE/kgmfedx2kGzLJjWcZzuZ11PaNOQdD5C7eLK5OidvcoJ
/+4c8u14llXEBOC9KqXAPibD+k36th5N7dm74M7LFDUqd+W/rhJIVIfkjZqq0sufugMU83Gjcdmc
tig8H2x2/TNZj2i3PyskyPiRNQJVFZtlkWhj0D3ODkO3xMSRhSisVxJFeYRABpp57+W3BP8SiGL0
BbmzAz3pYtdAlrL8w0pgTqV4fCW6yxDV8kRA5JHVX/Hl51xIwljoXMfQcnKkUzNDXXdLd9jFJwpi
sYPKJib9BIAMX8t2h4uqFZTmjMCqpBy3Ro6CTaBWAypkFKkFDKo+QnxWTEmfdLvSAbCLHvC1+E4v
KS6rUBeEAhcgY2Sh56rg5GqNx/R3DE2sEqM4Hj4fSHuGrO7TdN+igsXc6Mqh4t9E94QI1bSB6x10
VDJ/2Fgn2URc97x+GbBZEd/Ran2ZdTklor7PC0SzmXeVBCYMMW/GoNJ4/PBf7F1suzi8aVVcBJeL
jxm6g3W4r9pi/dvCvkqNn9DjtgD1HAAPcx73h4wQ3GVIrCBeFDhSeaddMZw2KypBM2IiGVmMFUhw
nGMXVMT+Pj5YHaCNiZpOlJ1x3+XKf9j9ws/9eGZ16t/E8Fld+jAUIYmCb7uDNNdfwprxa7w6R4Wk
ePgy81ScmPHFGgBik7s84Hus5YwTI+7Cwz9DaEuSCL37QhVkrXp1IZWr4w8zCYlQhoBEBi3hHrbh
wC8U3PzjYWaInBos2336r2qd3XtRHi4B/riJBvWJfXMcefGC1gcTER7E0jMpXFJdDs3qCDMm+7kf
4ssPK99Du/k/UA3xjCegJn8RzCThwKYInN1F65jlwPH66v1C6dgiEQ8lSp+G0aNxYin8thjyp7SV
qCQm0DWuQ4E6jVtq0vb3BO2YKNhd/KyKzPOY1ykBM59Le5z5IwLnXdRJ//1Ikr7O+1Rspc10C910
b97YTu4AFCaL+6hzWXVLYZuLfSgg5CTQO/13DXEMQ5fZFCWTY8E111PvUJYYooA2tv5/lmWo/iQh
ZPLaQHFn3drw2FOsX2Tl2vKlCOuarpQeSl9hMdPdVqcHiEG71IBqo5RpniBA7tGHK2TlSSYEWMbm
lCUr91A24V7gXOu+z2nCOo4ugKSYO8gKEa+TmsVeQVMiVcP9dQZBYMh74KrvXRAU2oEjMeQQ7Jmx
1UFAEwHIulKL0h8hEW05lX1Ax3pWV04bWybsXhoVCt4y1CStG7pD2YLBN7W8y6TNV2Hpb0drPCxD
UEFpUS49O1BAwZFN6Vpzm9Bd6Ldhb0OTbWA8AVdDwU1ysWFCwUI6+gJ3WSSnr2HMrhf6NmtU1DQH
Ja6geQdPB/MsE4DOxmrDbCY0Ccqn2lGZYyipsGHNrHplYtUT/6c0TqYwwa1+LgQbWTV1lydiWYQ2
StI+UjcAyN2dgA41pfVPuddfrNvSJoVykKOiyGnLAfjak85qLXtWpXDWTeE5c3yDpjr/43E5GD7c
pWomzBZKv1uwLjhPeSEDWluSWhrI8jj0XooiWcymoxAqSkIefjESD7485YHVzeSgcgmqu0yJi4vH
j+CkJYc7xBICh1z+YMLzlymJaxezlgoLr9tCgmHVCzqyOmx+2bYM3rtEatTd01DFzBAJyHGimAg7
B+yeXKmb6mt9y/DJbLbzfXK3va+j9qnv0NnCyzmfaUpyDEJgeoCUoJjeLZl3kYy1OInqgrjNPRWS
CrGfiuU4Fl1EFAoTRYr9RV2nyqqCm392Gqjz/6fiCkJbPcBH+fGNwb9Zz6EYfG71RuHYt1m1I6Od
J92YR3BuZfcYE9KDbqiOVQnLqB9vvvWPzWl746YU3lx2WR0zw5FnBN6S8tsNY2vp4yI/uYmoVTy1
txNzQ7eIBX4ESzUtlETwrxKv0alUAQxcIEr1w4VGya6oI+fTrU2QMNDZXvMyU8DSVcr3MwfbWJ9P
q+JRQRUELQ1SsmcZ5m/pQNYcugTjcCvpfUSuhRXgKqSRqys5ay+pW2J28olfOylI5ylxiYn9tNT7
MMqbC7hFLVw6ql0568RghWHMhaJHnmi63+n2/IvwiMJigEBIdeRiW9081A89hKiVkrzejiyIoeUk
F7KN3jND72GksaReoSt40Nhz/cUwkzl4I7ZPsyuLqTgsRMg//KP6NSYUwMP1uqJHn5C1GkS/kzx7
xI13B3lIZwfEns9VpqDiyvjEYvAA3ojJy0G0HqrfSlCxAHBaHCfb96wSR+DbrafheeNMzdCHWyg0
YORp36n3DQ0uwYujRmVLcqEyaqwEGZXmYNP89mdbrlcZjBID18wnMdBZ/lgzqDFbzgR39dCEh3nv
wbs40igU6wE/RiUWGqImfwbXng5YZGnNtquEO8DJtal0sYJXd5/67TY2daKUFlTkuZyelVeFjRlQ
kpEfUIZ+7T037ds3hLuouO5gJPSWGMK2EH6LwdEMBlOXKvDxlLnfV08D2V+ySPuJ4YySR0IRBL64
cqjVpvv+naeIJ2e1XPGoohLFFNPkYDNq6kVU9Jzee0I8sLTkmagpWXeB5hngwt/VMfC4tQeRtKLe
H+SAXidG+CJ9rKtkIRUd02kk7hXmtK0Eu5XKlfhDI1WnjARHFZ5DHF9ZJbhzhREtJrzu/SO1F2Qi
rFsqL5gcmqM9vJHv/fZxBIdcmV6WdIg4snjG/LLWDsZbxt9KRwV7NxdpPT89pPp0Y7J4A2WEWbku
D7lU6RlzO9xwTKfN37oXlgQ3RgPBRzP3TYdO4F0LFtq8VcDrhBQIcyVv20cF2qcBTp/GNFsWeoBm
XEgIiXxx5BstkzyCt3VaKwSCrVFn6QKXDHlqF47xK0Ge7XZW2XJWyobY/4JNoMjzY97WjQiVW1bG
c4/5ii3Pdf6x0mUp51TsDlOfIKvtNCqjS/twJdvkhyKSM4AOWK2wFYdpNPAv3QxZFf4UtTX619jX
GjIkgV4oDyrU6Ub7UDYLS5A16Tc6oou4zo2hF41WGVW6G6bV7zudkcG+kfa5JNRTOSihR4jHhnF3
lVNoYfnCIf82Yo2lBR52XQxI2bDtG1Bo7bj/GuoLaes0vWaIwUQocyKH+FL39UQURAZCX/SBz6O3
1f7Ls/WCJAWvLWCRGQNdkdcCNxki5UYTDgYCZQaebCIeCzP9/0HlozV4RdAn+s06PLFpcR7yM0aJ
K/K2TPcFL2C/+ac+aa1kAHzFLPlXxw9dz9WDaKqO/9P5WNehbv4G4RaxVKhDLIfeEz278xnRa8SH
pTXsrnu1LwuGSZPnULPw5HpYC19vu2jQw0sBVt1zYWlumXihAvTyRO/SPdNZxGJVDUNAfql/1m7N
XxgDHTgNaPkzgcyY+dPh4dgNE6sGjLB+8Rgt+F6i6N1CMNgQbATGC5ECDrSXNT/H/WJV/6zP3ulQ
Iz0iTdqFmQb4UVAyUHJ4ousqJ6p7LdCieECQvsG+TKvizdFu+ycwSFGrnOmIzr4EHMx1z87lqnn8
qPszNWW35/b1X9mzYKxMQJ9et1EZdJ5hWCoOqfg3f9//ffvxXOuJxirYSYjIfEFEY5h4P7GIFvrH
9qHhQ5dDb/oAvopoYfM27I+AcUvG8NcX02AyLwkLt004Qe/WTvo1LHrWjRTeVQGxtrbAPOP8s75T
sZ0AsZ2D872hDwfbH2i0XOMZi2Gr9B5bLzYjDvHvDBEo3k5lBszIRP6BFoRcbKV3AJLvXcagqQ5z
399t2pey+zvBRAknDKg0S2h+VH1DsGIUzIO2bWzO0zSr30Uul0FvwRltXYBgR932M7fJHBtzjr3g
Hx3oE1WlXCs70j5owrlS1EeAo34G8FGh1b6F4GFoLdUm5gkGWLGtUpROpMiXly+lgGhLcDkJhmGh
wTDAUVSmifb9wZeIV76mXyZsaYJgwZ9hnDBT72zGO1NDWI+YrhHn+m88G09occfNfbDyJAGMONwr
f7CqKWJG2aH7dt7j04cCaF5E3XMrwVtp/qUjSb0A1/UPmR0Mc/lFveXoxOWS2cZPdKWh5D8k414Z
WYouUwOx9hmA3bAtL3P2+lal3aWC+2cVGLvhliP/GPHsXufjvhuP/+4k9BX3G8VMw+/UC45GEofH
SPIhnh/HiBdEV4VoPn5rJ8XtFAESWMCmKcEF8bXM0qwqHijlXYFjtrgQvKCFpPHn9X+yIbtKum8j
Jp+Ys/ChkUmYFg07HzFRUbuTf2EK8R5nJk/EGw+D/C4m/fFyAmQoBHZr34iqjT0hAJy4B69AePpG
A+koh/2e+FxUuHSfFH9rgOUCdgS0bmyGEtHemZKc62CqdRM9EPfzMT9c2q+LSMlff/QwXM9mP9Ri
7MOiGNt6706VjIaoC2+e284Enw1nQVgf8UVi/2DPh+ux2xO5o1gPmKTVNWY/gLSpH34+6kkqt5Y1
zjYuHDYHLGE+b11bXHdXFkHkkGfudvHkkXp5G93gMHfix5muck0n7/6a6doQUlO5xsbZyVFVGiJy
HU0daWJCxbg6q0u1JaTO9/ll9FSvzCoqt+0MNu6a205d1wCYTehV0IOO2ZgF1QyPBf+rITFjDD6s
/M9v/QsNVKdYvHSBLelW1o9eZaDj423wwWHJuaagn2uH/KUG0/v3gOewyN0z+c0UF06bK9ns+xTI
l7pkerRJU8tJrc2U3mbs8KwEJOSIS3XcHXVvre1GFJTsZuQdPGMRQuQTFKxgUlFEpZ7vrYQNCaCG
3czE8ROMN0rY8hxpqKdot1B4U0Fkp2gaI6GqHviEJSKRh581T8ZSPlvKOYCJcLutapAsv0/3WPMy
rE1nrczRMH5tVl1JTfIxRYvDzLlrV7mIKMqdEFK4vpmJSr8ilEKuB7JDv3zfsp5gLojyjHkcT1NE
QnoOkxq4093sITlBhmTuSMQsSGRH9riIQ2n+mczBjZK2c9ptrqmgSqDfBRDdbgAaDe+mPZU1WSwD
SkMQ5wc9smpDKM5MoXk18ueBhkVjdRolumDLJ3cnaVDTwIzOxBibXAlgb1QD1Y17YY280nmJiP/u
VG2fxhO5zwVN1ylPrDq2sy6hqdFww/oSq4NGgdcez3ir1pZqHX1ccO5h5FQnv6Kf8o2hl6SpMNkC
QY/e1V58kX02vvhL/T9EcCCb0cfaGVH7UpMFN9YRdsAbAJab+W1nvuJUYud2OuJuFNTcn1RsnNtL
k+kiQ+EMYbK4VH6TkoGM2mOC4dU0aglzfOzTE9pz4qmxw2KnTTojFFSo/O5FLNnR2rDB+ytJqnfk
Qm2lKglvdZ5IKlDJyh6TOaZkhgxyxYeOosRzOw8gEh94UZGxx1WX+qYNiiSG69KA002OAD/KTwaf
5BlDQU6EdW3WqG7Z6NFuMhuIJcgTmul9nw59lPicCEwSDmY14s1PGTO/CblqhGvK6ttke4Z5LcQE
N6r8c4E318BT/mrDXSF4XiWGiEzOh6glZWMq7S24U6kBZLn2zeiziXV6nTcwPGBl5hhCoVmDUgpO
8UVvpcksrcRqe27IxM4/qY68sgRMi0X5hk56KneqzsZT0FNwRKR0GQq+sVhlKTWRl/6VqawaupmK
d5GlD1GeMZQ3+5lZtgHR0HcsPZTnuKrv9g4Nhoak4+sN+repgdbhlxQJ61qM+i7xQ0OH/N0Y/Tpf
rMkMZMGmWAzyFlPzGI/9h8rxlHKChObhbovO/D8cLqWtcy7vENmuHacz3Bhue4k1qeKbWw0VjSLn
LUF6VbXWo4F5yhs5y2EeBii4y2+Hxs/MPeV1Qv+XEjTl31pw0RzdBGw1aV7dEzEve62os+kqjh5D
Kgl1+RjIpLvfDpymE08yCvBZhkB15mUmD6CG2x4A4xdkyKdjhOddwkpy4iO8Y5IwC2yvR8aAH1Gh
EKx5ywwPRq8XUpgL75Qz/L2xLWoO7C++Xl0MZkbfAayp5NLTb5o3h4d1kbhAFbtevR/ExVPlKdy+
q8JtmMxkadYJjPBB7vKLFTqb/jBZ0fzqErE1LpWBYmivsiUjIw7lvxcamfeVUbRG9aZKeO5rJBEs
MBY8vdJoTdbUw+fsxrd2540i8J5XGQK9AoTcEBI+UfUhTh8RIZVz4PPhT3rMJ2C9X3jksMX6hZGD
RFotEyOkygRvH8j/s2yjUdSxO02wj0tETFYPPklsmaj3ds3zDMdbXNwbXtpt7n81BMJR6+iprrVB
WTfzFQ/yQCd/E5cwXomRV38EEcSeAItMIIulmab5TgK6FObw6KyK5YTRdh080AY5rOyaTwgxcOBE
1Bpj/dNe3RLpcEqU7hfIJmgeR5ovTxWQiikpVOaHljvqmLQFeUNf5tbpr+J79PCzHga5gPiDJPr+
1Zz61yUDXA5E314bTUqOTvEtUseRzoD7/waste/ddJhI2rQ/1e4xX8jBfh1+LQcg9Pseosu2b58T
kwCwo1YcOVbVyMOsZoTco9yX7srgthhzh4FPKv6bD7J5kFjucayzqm22oRd/eOoZDcTcbeIrYDP0
dioAf8vRUOVN2dTpmirVTkpP/Cxgw5Sybw7G2ciL04o1NGksI4F5GIR+YlawWuM5y75AFZpVoMhP
OCswAnhGOz0BWbk/GYOBsUvwu1I1snYJeRem9/p7vfgWtn6e9D+3i1ta54FaKBDXK5wrTwylXttq
PG4xYHN0iRPij/y68zDGv7FHTEh5tx2EGlxEXWGQLE2nsvnmVCe/Nc3AgTHuW4vJAiAJrAZLLmkx
17H6RR5gR6SQOpaTFEXSSP/fbVXvlU+V23zDidPpY/w1cvPoX1RIzEOUGlJ79IMQuOX1JNs7ZJW1
kjuDFwj9MbmWnkkS0s8C4W6MpDBd3osFou670dGYHP8iFrxlznwPilhsiQaakdaMt/z5hUEzRI8q
shu+P15AxuZaTdr15GBHf0/cAE5BSQsji4o6C44cK2s3FGZq2GTXGvqesfC3Nuaw/gimMut7TBg5
uMcrp5Tl0tNrvQJwm7ghQbd3WqkQapSW2UbkkbTxUlxdH/bVKt1m1buP+X4N30tKQ4ZgszmxpsSN
l6mlQOb3rQNUYl3hwA/2NJNOJR6YmF7a8UIG/60rZglXOdrYnJbxlWaG+cJ10aNf5nCGGIzv8hOI
hTCFQb3TH8foxaR/dFIuzwB8AwDq4YulMec4yjAsqxjDEoYluwldqhuTyTERYb1olTKhBC4iQM7g
+DxkiZHu/3jCyAOthXaxLPrQlWsM0lpxVLIPkA4+pOxmZUPPPNc/hmpEvSukf48bOTUQhf0AQZ31
+5SQZpWAH+Ks97Sc1qv88qrXCOEWKz4cS3gCGVhWksAIfzmuTW7AUXeThv5/qc7jWi/bVixjxWeb
zsv4BxnT6tGADrFFrHKUsD/1tKrISUAq60vhn77OthnJqIdRqU2waA3WPXdjLfhLr6cisVuijvEK
4THsD7IDvRs5azzZKGoYgNnP4UwACAzz/HzVvODimrh428UYLjbA3QeyFraG5cwW/TpVgZIG+vPC
MWLHz4lplgykip7i2EeFUCikBDT+Rh4I7gIVoyELOmQRuMgYdxW+EorxyKB+fKzvbtgur5o7b61s
fi59ejWwcIA5d4eFpqAMaTEYIG9ju+hngXqrqLn/oJ6yJI/pX/hZMmNd4h0MAYvsTrK21fwLz1AF
tP1t3Bm/wraStNIT2+WSqN7MO8K+h5IuBVCozWC3LhDzVrL0YcFUlrVKsViNgY/wOMhp/TOAMsQf
ZTUWuyQ5EdnsSd3wTayRwRw9yvyRxl3Ddhd21Mgr8zCvGziCzvK8RvYuZaHQ4HOnhCFwbCUq+DRU
2iELVMZZzL5YtqvGuNCe6EQlg0ljEkVvI5kUqqJ583atSUe1+O8OArL3QmAK6RvDPlM4UP2j4gu6
VQUlfke3fbaNPOzUyMwT09iWXmW/Zo+DcN2sUvfTwN4C8URHVbBDmn74j/DjvJ4FiCbKOLsm1LbL
F5gHPQ+6nsNbYBv5tHUZ9JiibzJiVuD8wHyBPFLV/f+EiEFOBfVdL7Ndc2o1Pz7IP1RrSUg2JKME
0+11d7I9yoaB1inhgfmbNB6g/wXzxpCGKkQKwQRf0BxdEeUKWfofMaOaLWXx+e/Ct0Bp+s82khIw
bFVvfS6vxVmXoen9pzHW1HCHEgEW+8TNmSu36bsKTR9WsyYzmdtQX7PKXf+ncceU3+AqU6for41/
XT2uxOmpbw5gpdOF6MM4gcV2ftnr/4zheyYT3YDeJ2rqh48c19S4gsItuAiegkLSVSJOYHsD5Q40
tGumdKuP2G34StAGSzgI0uAXGIL4QIAcJbiG6OMC4QTa5rAikX/lFAQ5ix+Y8kOT16Fsk7WCoXOu
D/t29Jzj9FkwtCpY249EvAkGTqDfWKcMCmsb3pJKDkaGUn+W3VN66qxR9wXb8l4Lc49mmH6lENLW
viNB1ShcVetT2/nUyTszGfM3CrSY0fITlhWcwwmaCiBQy9VYDDhEaXYbCsQYnCveyXAlAMt8cenT
tUE+srDRhVSDM2WWyVyL6dkSOH/sQcamlEWnahxnXqKoCcEOgQu9l0AplwIDN6aCga75EAZC6KEM
6Kl/9nPdCDFrsCfPWJIhqluNkBPY7yguFVzjUyUXRPx2vLSxFfaND8pujICWZ1Ek2n8NoJlWBpgO
vNlAX4Cq06cFKtiPjNP3AoOXgMENVqiTZ8ILNztC+Lsejm4O1ZrovTO1NgVVVkY8PDPoyQIJNNHb
0VsyGFMle7eiUFr2y/9ZstuwSoVyBriHJ0XSL5p8FqxP+nyJcSBj5jSJlM8lGOW8zQj6yhSg3lGE
yDne+zQs8EpgndhDp8ET5GbBEW5GYkeWeRs5yhQ0PW0vifIkwQIR4C0ZOUlTECX/AKX/3My6/6iy
S41YxJUNT9IABY66Wbte8mrdhQ6QzTmulzJMzwsi+0Sh01qbzECfBlw2VXOhRoM/sPT97dddF9B4
gr26dMVT6pabf1U2ydxD6dcKzwDV6ZJJcFgvy4OIwIggPNaYZBvFHjBoNH3v1ravAehaMh3ydgXi
e0uA8JzuB4xLS3ySQ0GWJFHJMHFvf2j5fCTUeyzqZFwEwLiE5Q3DJ+oADMrj99gOTx2pacB6eqw/
VXQ9uKx20MAexix99GGImS5MR9WOMCbWx8PXXakzGF3B04s4KRmyL6fQlZ4ls0GzsRGJYVwuCe1W
V//qo2nSTHA8UZfA+nlDbbhkgVeIpQqArG73Vq/pMRGNmzV6/hOGHzN4V/1ccKkFom6mik1E56JL
p0Oqme5Go7fc0ELYLwVWPcJ/eq0k+RaIj5EWmicG3FJXtpbZjLxTcIvTQfk4JgPxaIQKqoTu5T2B
KBa/y2PLoQMUgY0OIsJBIHMOwnyfrAd8vUIqrGfBS0HDNCM+rhNVWG+UYdZq7T8ze7Fz8y1tqzEk
4DQBZ5htWmhmP39TvsrHb6Rpdb/2sMFthBo4jE+xJbzBSlPrc1ZWT23Pp6mc8VufwKXB2UbLG9Yx
yHVVyJC/Wyw98hDGtUqwbUZZvCS8uyQjCoLHPGEDIMjinUEVMyU77qbqVDYOS3JN6d7vymECMfrB
JnCycoQIJRW3vJha99xRyEF2BJVPq317ruDnz1sDoPqrurm7CzN2ea0btY2GQYOub0L/RMPB/xh2
iNgLGB0qiG+4eVwTL8HsDZSwtq9v/MBgeXTfF9anB/0ptSRg15lAaDGKdt+vgzKjjmLD4yH8dqjd
g3m7ZSeKDjxBcjTYTSM7L3RBkhjHADtEiL0C8oV7AdxCdaZzlKOg/jn0SyNy8otr63I65lHLjH0O
xgWyHZy4YuXD2O7zEbmrWT9PuvVYbfRfJJXc37ehAlyBWAfMuhU57i/XT0KatUfj011SuyjD+qYs
mpKdKD7Xebd7WeajWMxrgOBUbO0oITCKUSoEddEgSkKir0EfuQC1BdmdGFdDq/5Y4gwY3fa/y5mL
4Qo9KZkS/XYYxS+r4KzjfcuDGNU6f7mvIm6mJB8aGiP5lLPhWj7Bvh+WuKkoPObt72GoggdpDZ+S
b8W+7aEvBJ22XmXgsPtJHei5VEOAVdmOi63dl0+3NEnsxqcWmBpyL16ZWdGliJZklik2slTlDGO+
/Q7Eb6MRJSAz2hDNwiXEePW6thyBHAeeXqrzkL2HDAVrmFXmO5gs+9BBQDX0P6NnUxqj7uVIKPY7
G226dkaAWQvk3PjSlRRYfiWEpfmcagGRzFyv9Xj/a7C6XiIHRGgfS07mWcRnF5gk2KjJypNJd5Da
U0v574HhrvBEkhkGUmppYkefHcWieJRpYDasu78tUf+09zyXdPxbQvcBKmL2MrLrW6x3WbsN29qP
to7pX8uwfFGa8XOo/PSK1Z/Dtlsx9mY9O2uq8QHvxbIAbquDdO+m5dzB3+bw+TQ3NBaEMtq+sbku
Qb4Tc6U63JZ6N1Vieo2gLoZ+NJE62Z3g9znPyMMtuE9S2oQhS23uRRpDcAA+wa2AmAgnjSjmDiKA
MBE/z1YQZm4ylPrRI/4vsMl/vrhGmo8lXVPvJoRtuz2t7pWA6recPxBSqVfJoMw2HcZq1jnOnqiE
h02VDAnQ09TKP57P/vmM7sPpMPQQA96HXcXK0TM9s/JLVGrZGyqbw2RH47SPixEz/a4eOiZYPl0h
6oqVMwMHN7aNpAgr3slvQZIKRwBdtfMVfnzbr6K9LPspOceGCQqcyMYL44l8z8xB9eYzWCE+8QKL
827NymSXoVa7YXjmOG1Y4gi1YUVt4hUajoNWtGkaoMC9UMoyJeqZmhLBTwcwhH2bFgKwKNmlY1JN
lFL62OufEdgQiJJYxq5ijPofSKm748FNaBcGWpjmZHBCE56EZ/7dkbKJ+/J4s6y1WBm3EiEH6h4D
LCfWAOGRjvOoENtYDezL/FXjiW3EgwNHQ+WVEbMMg/PGkPROZjC9Rwxugmm63vE1zGS+2SQwj45I
AQ75GL1BDY6xSBG3E2ibZJL0bd8rTfPMqQibi7n/xd2t/KjekTWDgoFQ4RdfRkRmac2bH3VWDLRP
q5fgWUwvZLvBp7GaJYAqUh/6ZzliQuoWkJJaTY2pONnlEat71F5cBPM3Tn99Hk0YZjpkpIDgIDuR
SjC3gn1ArRP4farYN3sz097Jyz03kVWqwz4OXcLamU4smZsOLVj7x30PTNvSNfKZ/kXwY7xr1wNP
2Yj0Gh60m5rhIjkERHR+4/AeKV8O28rov34qdWAjmLakFcYnH6rCJ3yZREh2qyN3YgG8Ls2LDUy+
e9A/EFLVOpzHQmHw1p85JL4je/zUh45yauN9NwEHisOrOiLlTF3a6IBnlFRAKcOCTlb18bJQe09R
dRXGckWHNIoA6vRvkLgCpy8RxOvMOLniBrDbZSxjh66SGO0Ncc/WHGaZq4rL9Gm6DnzTpiNsJLnY
WqFw3wOJvW+4kFszqqxOfhBnUkLcjKhNhNbomj/ZalQ5KpfrpN5ne2s25HYitTNw3wqXvl0jlwBa
aYLVFr06/SuCHK2Kn1+f2M78aQO+P1sEMx3PjkP7m1YXhAKkgVZBdwBvVwTl2+QxdQDdPjCPMsDB
lkYAdLJtXY61CNkrmjI3enKNuYOzBybvDC60EKEtJ47Trs7ilg/4gSZRVrv8oHf3IbW8PdKGIS7d
Uln2QU88EQ3iwkxGRxzctA8ZLWG7Y2DzigPVGMGXLJgzrc8+AzM9+GBRpCKWLccS10nYovzwA4j2
56llR+OU3XwZKoZTG1f9j8jCII4UyOk4gJDUpsGWPam5wEuG7eWVpHUgi87x7zoX6FkNTtE3uLmG
cHJmHjKIv3Rdb6txtVKrv7JUh4lc2bQSAoJJZZZxMKET6Co12/5fAW/nL80KPiE7Ahyky3I626qx
LxDyvW9fHEPwWAIIcWsJx2GqU8XDuD6+eK5V6l/cj1SsGu5awb77Hf8XyS1W5KkPpqDTSjSkfLij
hzqFfqCmi5qgWX22Nbc+MMH4G09au5QR8aRqUx6y43PVz4JvLDHXshV9NcxQuqau6DOExSfnyIt+
eG8uKo4XTqJOLEg1UqyJCrFx6Sx8IPHwUQEd+sycP9pgtdgYpdbqTSO95c2p7yc6CjM3II6NjIaD
ZNo8Zf9JSC8O17Qm07PByj7wWHZ7eTRyHMALmFgGtr3uCDYZkvvFvy31U3n+FQ4PHUwd3nkQ3sGC
204lTHH6XZFtMLvWJrHF412NrilUcP5mYzAPDnjzcaO0kNHb5sMqlIPIyCD7f2ACUlL+SJy6mdBY
DBgOg9vYQMQsblH82HZrOzj5IaD4cvcGT8xctwHJ3epqzYNOI4izzSvBOlyXHMh8v+vrT/d2QAUv
9lFmhb7fJD8/2jRuktHjSyp8oSKMYyIYb2o0fy2LIqMQwuWViMnUKIrJIUka1G4haMZqjjVwApQd
SGvdXDzm+RF7G0W5NIs8JcF+IPH4CBvh4cNRSxIXohXNbi5718Km/GycplQ+IlY7HoVKr4sTNoEo
+rjNOijw4Iy/vE43T/IGTpwesmixhBHy/Hdrfr+SD76xlcuzC+jUcDaBOi11I3waqXfrR4jth4XM
OidUBdKC+amDZs1Th4EnqFhhzN4MauzsR0dWhRMJNQHpf/zcDFtiT2TaoebuqO4yPhEgVpPcAa9T
UR5rsixdngbAxzq4bZzgJCr4vINU25cJLbhEcaWuazXZnjTwjVjGDuBv3XX9ihGegmAc9hyFgU3w
3mya8F0BAKvnN/llc+uRLmOcetpbob3Z7nbN++/+WaXzt01OrCIvvR66s8Yjh7OtgNDFgPlyjWmi
lNBBKyICc4e+5z6scadN4fmMk1EqdPQ0aDtyl9s1bZixU1bk1O1Fi2GqzxNnMUESODI+Cc0fSAOH
gV2g3QgltmMy6/RBIMcEZcq7JurTuSR5I1Gks9DNeAU+44/rl8kWgcDFu+giUm0wGYbGaPn6YmDE
LjZ/ASKODoXKy1i9pj0Nw/hvMwvMvH48QztKndjUziEu4hG64faWvYMJrgKrpBDhdx2A9jDf3SfW
Hy7p8CGmwo0lEAVV5x7LYSH1tEEJkp1OLsOaI7XVaHwjzifMWGCXeBbE47RcQ+CSORwNd9200jAT
5Z9R5iOUvPrJeD8wopiqpGnNw+5Url97PKrdQmjDV0RuTy2VjCj2jCrg8fwLTnKLX53D81iCshzW
Rp+Uf/d2xq2qF2jufqg8MFK647xwWWrctYgV58s8N2oVZRRhqvFVUl28dDdokf89usRrWbUCVMlK
0XwDgoBo9OtE5AJ6t/t69xvOZZPvb0LFZzWcDA6ALTYEhPbEbJYUNYG3mixABepHFo1Y/nkrhDIr
oaQLi7eLgfTSitdwEEmID4AvViLcEqC7LP0bDncbqqYqI2x6XxFFYpaXbH3lzO2Ggl68Ki7Ia86w
KqbyVA2oaG3WFzDpt1vOzsQkOuTTVBMP5XjpAUguD1EIlBTEDWCOtSyeatKbC5JjGG2FFCf2MIJO
3f8lHEX2IB9JLEoqJW9ajhL77UkFEZVC80fZu0yRdJQjAOt05Auh6q+SKYbYndYL4XiU7D0t7A2+
f5yc3XtYQksEathQi9MFOaWKT42WwakafIdHwBO7plHFGCfeWuUOUbTL3h3IGULTcmTpNhuGNBU6
dJbRfnPHe4Vl1MoJeEiEjAZCvKSAmzDnujBlrH9YrWzPvs1hu5VHsgzrRu17HVUkHeA6V0T1erfH
PNBFBA1d9a1m+lqrCPV9QRbN6iKwk4dv/4o+Vzz1JVxnBgOr9BVy41QqJeP6EO+qdKMstqWohaHX
5zePB+uHomHaesM22Zz+9uUlrHZCtembq5cnL5d2QqvfVPcZj70ZiQV/y+fezrltxz0KCBkVwUJK
Y025EPhOKuceKKHYeGpcXvuVrYSacpm9cUjG+RgpjHmI1FqcvdvUR6UmoisDLduqbWHNIVcyDhtm
c1licFDSHs6bxLjrFVb3poXvf5/b60YD+tlcVoKuOjrARM7zJDkgPupURu7w9xTdSmSSOrLOGSOj
FQafnxTK1usZVC0YPx4vdPVHIUJJame88sG0jbOi6rnUlQRISEyw4HRmskN65VJX1GzrLfRjF8R0
9RzIeCv2DbKDptmWmFJeTmsRKhJ1esm0J7zpIvPU6WiOaN/gYm5xis/34WJ6Sdzl1hOuR8svXpJz
yW707MpzPyRKj58PFse4XeGNhlkf2wPXiyPQ9yRbg4v2rqQ8e3VxSH0pnGxcqyN0fXqbODKv1oeG
Qic4pm+LR6feYu/76kOAthL4Rh9LkB/qaH6zmp9HP2uvXYmbUsoNDwas6OLbxXVB3PgbXSOfKU6J
i7vLredTTjUzRgKlc7Vvx7M7AWjtkqVJZj2OuyzHAJV6axbooDp+OqbMxiyfD3ieDSqQiyf8ob9U
yshIFaK6nROXggDU88MFmn6MsSP1/Gd4Od132jMXFcSCPabnTaQNVKlGdAPC4jXX9QAh2zZW77ZN
/31kGUNabDOWDGUP+8wfE4oti3mT4Yv93lio451xV9XsGFrbrDN7F9/uNfYWElqU/oIxPKnrVX1r
RiGNMnqLFPnCjEoJX0ysMcmuCVQLZxFGDmd9cGgWnYfrMiK80R74P0kaxSeJPNZKScasUOa9Fln7
wMG3PlbK68wqkyjBhqxZRhjgRl1iuDoNz6R/K1swA4MLv2GlDAGXpsq4alWYFuRzrb0oUQSlG/u5
Rf1HNaVJoFeXbRBToisL1+msmfjF7OUn8zPOAW3iYiyAXG2+u0lW3eNYtTgr85WTKIHmmXxl21ce
T4PUEcj8xduIAuBunBq9kllJDG8HPZKYunBDjC8GfEqPMgQdWnoiJCLdZuhaQ0Q3nQHXZWokYXU1
b3Qa47RRejo6JXNFvdJ3QMCbEvHcx3vt/J84UjQJ52zRsUK3iwT6alJVz9U8hmIAXK05nSNNUJIv
jifKHEB7wck56cNfK+Voaw8Xfgay0ShGkFNVEq3GTH77/WwVp+ehzxK0i/eKrubQefKGEKDtCzCb
S0YW7GTbV6szoCnJa9E0wUscFrQHhHrqLImhAark47X6i7YxM1Qmaq8uOw4YB196fCAKRX5/i2Y4
iwtX8LncU7Xys0wWq9GP+ma6v45TmmWRQpy70rHFW6rn6EK7Gwv3T07s41qU1Uxuk7Q8KlnCIzNv
mmxBiwo/IcXKtVEIeU4Q99JtBSMfXAbN5/cZnPhy3LHWz8/+DUKEcfs9c06huisnbVa2VAgTx8U2
JJ2vwLXhtFr0kJpMqLAk6SRDmGBSNpcTVaujIiqpbB5kpJjaQDx5l8YiOVFlh7p1xQr998Ei8myv
VbPjFfrp8lmc/fTrSj/n08YdRzl6VImev7VNHQ7hwC/6kJSrQJcHqgm5tw1X02VIjxlcuJCcGDVa
mD5vJ3gCw34o1cyD9GydDsOZtms5E2K8u2WvzCPUv2CA0UsITwbBZpcRB7nDAzn700AHBl7LlnMY
3HgQmmERWv5yLwuqGZupbqiFwTWFnC+c8l4PAzsQm0neh8jhpqOgMqTlHDtqqmCwxPd5BL1FGMoD
f10RcDUscWyojX/m2dglNxbClGZ7FX5OAfvcNcb9LfgKT1B+AMhLE3Vqp+BryHKW4uHDZ8Wpqyns
kpMHbrAgfSe0H/rl5WeZV2dODMZQMBYwGYFvRDcr/YUh2vnABiKpB2oq0txNePSdpJyuMiLewCJs
DBUsJxq5UUuIZpU7JNap1owwMc1vBeI/dc9gasIPCezdbr+IP+FFR6fBhoAHe6FkHSEmY7MowBO6
MQFXCfYGWUnX/dDnBlu+KeVm0S4UJRQtWJZ26P0Qj4IpKZjAvlYK9Fv/YVThDjFu0MGfbvmXwKUP
/u1tacp87KwQ2qT1mXIBjdO8RUTfDz/nd84EveoGz2grG0QpFVidFuMPd3MJFfVxcEAVtVshOHF6
hTX00URA7K1AH3up2A6sVUjpum6rI76DKX7RhMGyBy99XuCEx0e4MBjECuBk/thMparNbiMl2DkU
ivWgSCtKYSdjoxpTHAQotxuXAjPLWT/8Vjrpg3ojOu1KZl2EBooMfrqHrZRgqA13FRf0K887Y5wT
1+6vNJSUmz5sdSKhGq+rIoyRAU88XRByUUhlgx44xDc4gvEOAYhMIi/Xb7rTm+bIq55FHSfIRYSZ
OyJtthiduxxJja46XtglVqz127300q010bkxoVvRxyfqV5mxHbqKaRK+MU8BHSuXwtVg3MHlUPu8
2ORULxs79bf7FnQhglY5W8Lbuc1b0Y+JKLmgpDJ1lFFZr7WbWhLWasjz0SRFdwdeUB6rCqclfXU/
4QH5TGQbwKK44/tI15fNC+M/Hcgwhf6PZo/EbWGGolkuXRvy0zsOqaDDocadTRYUKxOBPaJvD5p9
wwtG1ez5PgbXEqUkdwjza337AWFLNTXoJZaMw3ePacEDs5fTOqzTLPerP/miB2T1Vrd5QqXmTzmp
mg3YEqjpA4z8h+8AqD2iOi4+Jkh4EPbqllwYjSerDGmlFyMGMLblDLER2LQv/3GKM0wkzk+7sqnX
rOGRMkfgCk5SGTP8kUEfjL1itRhmhExbRRYYbXKNI9sPHmePtybvecc/e3JOlE+5cJdctkLJMMWb
osNLp5ObKSaDeKhwg1LwbBP0x1CBccbcMZMWw/TlEI0abI8X+rcnNTkzsEnq5vztppSYobdw07f+
Ydd3khA/emwtjVI1ySqybO3+lZ/LieTMAxvaCTDxLt1py5HwpuUvPqJNWm0qm3ZQsi8iHDNw2h5K
2DlUrFevk8d6jOGo7Y5UKV+efPtMNz80bwoxPAzoSSG4jvU9YzUT7UqX+IQdo0nM6xqR2yxhL2AU
PHVR77pTQ8HAv3X0jXdPIILdakMKFzubuuN/jR+fCHkHk5srANRpIUpnZlV7klgv5hHAiTshbzBW
nyyO8Uapumr135Xn4Chqj+IgdN4dAabakWsBLvp6NrltAo3OT/hiHru32OYWB4G1prD3FpVF0Bq+
vL5blM0iX6VA6gahHRiMhDgFUS2v0pscvU8Xi8RQ8f0yFwvnFYe2MrIVAaVoHZRHMDtexuBCIgh6
foXR40WNTc9T3h2xSZlihGMf67oFwL19nHnarTqqW12MDfD2tQYxzut2g+RNrovcJUFwmvaOxQLR
jB7UyjZOGt8tYr6JV+tg6CbcX47WvdSzw5OD4+wgRGHcekE2Y9eEddK7iCo1ZFoL34xuv5Z+hEbI
2+6fVUAGt7w4hlk7yclwi8268I9+VzqI2JDUf3IQMcRJ9NBTQHyct9+UKolR5HD140+0FBIo8E5g
h3zgM5iwgHzmraUT9VUsNEhHqpJ1aSzJ0eu/kUnUZ+/fDRAsq8UfM2JyzQdwsGj4K3fj84E8vFcW
/ZOB3dPI2GpyQOZEHDKKNZt1bVqHEnQeoQvBXvGxzxUjL0aE1m+PR3GTJZP/T74C6mcvVx3H8LXy
q9ob2PcEXNdJM7n6dwte7nIYIDu5rQGWSbh/x4xOfyyzJkW16GfT/aAu9DQw+6EyABooRlWrgwKk
PoGenB2a55fkmARvaWIvrwI6syHx/TCFBh8kUMKLLyNFWWRjAnmQi2jYvsupxPRnu2Z3XP1Nirss
PRZk0IZoHsamOiNXpV/4YQ4LblBokdWY4WQYz9qHHvscrZ1aXeI8ZItYqQ5LzbPWneGkZMAPeS+u
sABa7Jm3gSOC5M2RgVvvoA/6UFNKiJRXaMTCmwYE0EgpBlnG1AO38J19Ih9Nx+NC9EY4JZ3iJn4e
hXK1OQz2Irrf1KF2Hviz7CYjSY/KJFtQxxkH3SPmq7MAafVe1vdiWby4YmDOISTTKypl346vRAy4
yywBprZaUs5M2R+jSMJM5xVX+wehJcUOIsuKkcNzXZmuGNLwohGcgYWmH4AMnA6gj9HBthcxC9QT
PBgPjcLeiisaBS4GMd6YfaGJqgE7qOHfgnqwxgYHIkTQAHPfNux7QPl6ULsY9AKiU8hEUdvqlju/
q08zgjpIER6SZ6mblYm5OHkGq2+WPFKP4TWHGdLHTLSEnCn764wFIalTNNqCBduyuDEblRbOncka
HnoLtFM60d4YDpI9L/N1EVSmJa++IGyMkg6P3HjnXCwJkHqD0RU970lp8Q57PHNkZkPWxwXSEB/G
9m5EkqFQ4E/wYvSPId+/tRDBr0oBFMlW1K/Mc8spFe7JOpI9I1ECRdieOG3xoY7Y5Cp64jCnaTHU
3b71H2pifaCtdxcaj3T/C45ydSU8XHnC2s5XEJtlwcorwiivdZ0GOZqhLr0fi4zsZgN/J7BtUWeZ
o2kl0DvHpJiMmM6KVPoipR561hbIL1k2t/Tf7tVl7AcOULAMl8353LbnroMFO6QAvlVJOnWIhA09
Kq5Ay0gKky5CrmBolp3AmFoj4pcyCFYSmCtHfaYXjPlmN2AerPnFvb4XJf95EnWJ6vkrnvJ3xNqZ
M5l2U6nY5hcCljC6UEZmT4rj5EW22v2Qkk4FNyqf477XwL3DUlJB6k/v2zBwMAmRV0l9D6vnzAc2
1p/LVCBgYL3rJrz2qyjZV9sTkW42dvMkpl3TRmWWCTdYMNswfg8fxUcHZZ3ulF63YzrqzJBsJ+Tt
XKv+59rqxUldpVdaFbBenonKtn7ghD3YTdGu4eIpukjM1yjwlWidN8zhtIbMqSmAthK6tRIkQbps
VJk+/rnRsgk8ZVPbebsymu5/Y/LtqVOvK52lNDY7cFT4ObT76n4EAzfY7FPSbUzKJ1fiawqAmDN5
TNltfKv7tn8VbTlU97+VxIAFiTFXUyVqlTjaIDy8RQ/MJdGzpLJCKPXwTcWtRFM74WEHlLXtpPaD
l9hxYkgzkVd3sBf3IUpRNdkdeo4mXPV+JRtRncfwStF+UPwo0zQQcVWkkeFfQ7xWCTOj1Nze/MeP
80t52KvhXxb2cEcIXvyC5EA6TaG6iOmxuEYw4yTRxGZF8Ri8/OHFvVi2IG75z7uNnQU6ZZKNvUT7
OXIjSlUga1ONftIFtwVpqSoVgrbrkwr77r11rxvxkYBMO+3q71mR5bVvA3btLi3O/zFLUmenLPl8
E5vq3N2sMe+Y8dacWzbcdgn6rk16oBsjRY4gyrOmwtxAWHNLW2N3qFc2nSg56ux3W8J3iJ8oZST4
cCP+xBc7+gaCmUPwsHR+azaMBJ28l6EeluYyJRRlpi/njvEWKj/rYVk9YzmiR9iyqRuhTpKhJr+u
pE5/SbcnIMzTiIdUV+RMgXx0IcI+WnywrMNvvJgs79QEAt8O80ObKsWE4Gs24YXS81XsX14dwdmA
ofSm8hTMqdhYiGWR+3NbR3j16U6EdQ8DWhZPd2zeh0HBRaH/BA6R5e/l7tpEOEVonJCFbXZuFTZN
19mDBfqDie3+JbbFhMpv0R2qMkxFS4Q1+4QZjfINoc8j8ElGT2KYffVH9hgv2eWFFx6+VEW+22/u
0Gb+plWCf5sUm6RexgbP/hvLeuGXYNVRzrB9e3juuraU7RUWehsKpaXc9dpg6Q2aMd0xb09a0Wj+
xuWCXWICC1vtzaHFLZsjr/LyRvuTLVQbkQzwLsvMl4yyyrw9HslF7CfL3cybuRfmRqZYFkC58m9E
PYyFgg3P2YDsMcs/RRfO9bhK/UjU/iusiaZzErS39h/MVRoe28L1IVRcI26udlwxgJtKkSoWE9W2
Oj0sbOCquSihvjBPYf1nxXo6+E7ngEAZABJ5+3QXktTqd5qZLSCJesbYXC8SWEdbp6KMCYt9VueZ
+/KEAs9f8afjcH5C0+XpxBLvxcZW3RQwHRy/5kBYedD+yeSuH3UweeeCTeD5VYMIXjcwuQqNHKBy
+x/XScp8f9nxcYuEJT6Udup1E1zW+6Z1zc5O67qJpwwdC+O3dKeA6fpBHcjhfFBk+eLo4DPXDGwA
tgcyER7RTPrGhmpBptSTno7WTBirskku4CzT2wr1dJXUdCIpN0ol+Rt6c4+tFoypIUSYxefRXXfc
TGKhhpDXrVKhOYQ6BGV5SAITlWBego9xk7mUk/0mW2BorKMEOXoOPOOrWTNA0rqF2t/YaYhJwQX/
+t18t69Dfh4aGAxnEET5XNoAiv1bh5GDxDkJav6lF+2YSOrHFiy3odPsaMbgVGfBbSuu/k8FtS1X
yJ3xm3OzNd1Fm5pvuPcHd+YmuAhy6KJavK97h7RP1926x1RX+OVfQ8sVDPLE9MX/GNA74pwdD5sF
BAe6XtrNEY1OyGFqunjtt6/ULUxtjJLvyNIztKtbrjD6wIi21GQ/4gSVkIGNRobZS9VZT+Rbr/Us
d1oj5cJGomXODWgKNKePdtz76z0r6cxhesUovgLeeXB0aceOItFUGJJs1cA0ZKbphfnwHEHGs38J
j8BHLbGVnWirP+iC36bXaruMWsyWW7iXXzG33b7BhgcGGRlLD5AbulILjGgcpfKQOBIGzBnrTfog
/GOou/5I3hwcs1L6e1VvzdY3jya2VwG9/SldpT1IYXRjF/m25MIaKzaCQwm6V49UslzjsLKWQcVz
xG91DQL3+c5t1ekvh+Qu/o18YPrJTzUrvq0sbzzHCgQyFSG9MgMbTq8SkZf9dziq00JElM70zVhF
srRNtos/Wy5D6JXXrWttmkwoD31pGdy93VIxmvf/o6Fnwv5CVesqSKteh9ve3pGGvXJEHUpCFam/
6sltmnky1jYPi3OmLTeb8A1Hmtq1nDXbh7TP08LsnaxaHrAKXES0/RwvyaENofzC4zQ7vrzgGQ28
4cCLcGw/cLPFLgi2+edkzSoLf6CLEM+QEIlRsyBFG5yFY6iMDy3PBJqV41QttLEBK0UGvxNRr0O1
SIV2H/uJW9MTr7jvkPl1urvVINpRt2AM4Nj4Do+TVNFbiUhXhJYQVOyuP166tA0ptQNdmOEbNZ6i
slPDCR74FxB3iIOTZH9lvmhKg4kni9EnT4lbXiaQNmJUzEpkCjGJOsPFV8xU0p7eLOTuAo+BMEMM
//esR5/OQVI0juX7rPSDnJmQQm3xoKmiQo4uYrYW3o1p5D0FOo4vayC1jmh9jy3LdDECVSQvivqk
uMrbYHSjaLDCtzpIhANHjidjOyriE1KGw2kmjGX6WqzT42dMAaUsmvDrk23lN+JpFy96TNnWilhK
h1wQn4N+OJKGfTBKYlsviMiW+sKr1hj/MP+/TA8kPjSQ6igkB+KaMVwBnBylcFhTjMU+Ka7BtZ/W
GZdDHHmp+O9TY6UZv9No3mvSe6swqHo94WUkE/ul3hZStD5lzi30OWbjCtnh5croTaPay8XoSNoI
O27cxciVQ5b7gUkHR6NvcuRusniLIM/0uzZbmWA9fjxb/K0jMo3zKeWl1p7sswk392cUIiC7un2u
RpB9ElS3d7KBKcsBZY9rWYGX5n38JAzFoAQY2ZFb2mXNYfvVVD7jMq7Enf4mz3ZxM0ZsbF2cMv5q
XGtdjy8cu/p6jJr9S9HXHAcVYBvOgweYTBkEtP1INQ9ome04vZGrosJ18DJ39QVIBtZ7UsXqMro5
CggnZPcklrSsR2MkFIN/nfHEPqLst66H6ZMmqOsWfBoENJ1RtrmklT7P+OcwsOeV8gluzM+p8eAH
1jjuwk1ZvhJUztQpffOPPRdwYl8Yrgoisxkg6eEsiHvlRmlX1nCsaeD57KTCY3p5sQ6AddxnxeOr
ByD2C2udaxTz/XonfF6dh8bqvv9Vgnx8fk3XD1AVIPuYeyl1hyGS6o2cG92nKLUsDGC/CZLjqexl
wzFK8SfUsLE8s3rzvUeBqT4rTmPVH1a/Cg7xYz68Rl9MUrSHmOk457i6mtb7ce9bN0bQFjTfz2m3
+sse7RIGpixBXjV9kstX4StwNXsKps+KRzTBTZCx8yVN5q7cet+TLs+PFLFu4plZLCa3fkPYMqgY
88jCmgQHLFM7q6/nqVGcHTAFZxVA/aSL8xDXf30SBebbjQGg9PJPjkuTGhV4N54OKUzrfMj0VZhQ
+vN518jrYt1IN8k5AUcICTJnXPF2jejXdKJ4inOi4trVAU1ro3Sqgk7dHLvmMrzqQ0gvap8xalqS
0pM+e7hjk/qkvOdwYBaI0PhU29yUNmwlQytBK2ljj5tf7J0JERh2gVLV2sNgQ3aQ9PPalrtxR3LP
Uch++VIdw5puaJFnv4PZ7Sk67u9qR2oiQJC5quKMeSnXMavYWJ6rgA5OutTfsqectBEq077xCdaq
25nOnUI6KKCeKSnoPIpFVrfQbnVQM5hCOEzCJm1Q/C5zz/GG7p6ADkVzoNinwKjTqwIbkENPSltP
iNkED29CH6xcZ6Y4oLPJt7ECVYpg3TCBe8EbPYMuDUHUvMNmGjkQithyd4ypF9UsOg7VMXjwFLYU
dJbatBSu379e5VaETTEiT3Fvevl9UT0hX6pzwu+kH4GTEqGmSIEjI6ghXI5LetB6KqkL18HCHcuq
7MXxSLcDFiy6aP6+BLJEfrAUvZFg1hCMJjpS5yzNZer/dVYWY4NjuEtk8iOFEEGUoRfJnxLpCmmk
ANNmLZAwLfoylnoyE5xUicAxAMw6abpn9j4qr+lObwghj/Y9ezzm3E18BqXLsRKrt3J1KLLZNBTA
6nnJBapnxKOxGpWvWPLfHVxk98eMiivETEYhgudIyhEbG2Vt3OURKnpckKKCImVqq4bSYfxsLcqR
dTwnEeQ+n+7xnZs8JgZni408rmA8ItkWOuAGAAD+tMEGwBWU9eLcZQaUbCkvFJjBWJ+mkIOMSnUO
OUPOVhMcaxUAJCwSc2Gy8NEkbCG19smUm1A7xkOqrfUFOvV7F5a7/9Q/3TwLl/HVXyErPcFGM9fv
emiTZZlK9XguMmtc8mrM8/q1ugkEpMLbIF4rRD6CCZk6Ihs0WhTE+r8dZoY0xLiRgyO44+71N539
BOcd0Khc2qh9ESFWkpsezGLdHmTiPCPF6p2IUXTlfO0OM27WyjI6W3APrJWNsuq/VG+RcFCwhP2J
dMmzTKRYYlEjlpl73w8fvJ+37oJCoHFzlzaEnQD3p0Wr8oHNJOSnf170HUaCpUiLtPm7wTa+/LLP
K3tPtlFk7RQwZK3o0uqNzhZhEQ0xboXLDZ0K4vnhMyZqk4dclbk0GWg5wkzwSnMborP81557TwHH
d2riK0PJJA1fUXlMOD6j5p9eHYBtoIphamabb+jdRHV3kOkLOCFkHQINJ9zcMOGFWkjcSWoyQU2M
k5UUw6KovP8BDKrrAAOhex5loikWeb85gRJwi6B4AVbE9WO7kMhYtvFoK8kjino2aWyOLZyfjjat
TW6x8g9xeHvdjLimH9cizgOmAF3wE3GmyKftIxbETbwH1YtWrINiEgySuhRi/NI3NubuJiPA/tpE
m9z08xiEZZ5bp6YxjI8jLbv7WGDZmTwBVFqcKSLBqRZ98uewV6J6R9oYnF9vjk0WhVTT9i9k5U/0
K3hmjyszkOQcSWhrs8vkEQQ6AWiaNa2xyLWIGO2Ia9MG+8E7pXHp9aF9K8voJd9srJdrJ+CEryhh
wtnk8VnsLka/6RQ6nwAaaZzEgjX9yhUK3kiaLUYdmBKhTC1tFGqnwD6nPEnkM73T5exj35A59wYi
r+erQKQI6tzN+dNWsCQUaKxzYJXSvg8oasxcKpK1eaJTK8UtjGQdOPZNRax80iRTFB1BQ/mSMJa4
BJtR0Hy+i08C9DzxPov4qIazu4n1a1FiA5on+vPlP0zegTCuEWI61eKVUavOmqbbz5yznbQoxw4C
pwMrW7oGp0w5PTUFXH6u+MmXRoG2lJjkvRsssaKSSxFHX9fbf5Pje7GYz17V6jLobLbp9Rrvtlls
CCvC8pBsAO5GWd5lOgwClR1r5UugBr3CPECItYUew+DEaCE33CWtHBb9utOvc6rJ7Q4mNEZ5ztS8
Q/C/30YLjLP93uPf4Ggv/+IA7Vuz+o/5Dyx4Di40UfBJudUh8lMushxMl7OukbLAccPfj82GAvdX
9141YBIP459YtDm/3TmWXtwsTZWAXoPowVIg04sSN11KoG0rQ6l80bhyCHGL4G0efoyUDIxOW5H6
eP7oiaKVZqFqubqoZan0i0bBVvEZV3bTQpe9mQiRGFxT9DCd0IMdMpJW8lLN33WvIZW9y36dWiw8
F7JMBjLPBesCL1NrFcrYF16/YWdEgZKjKwyuQJy6NJEZpfTU3JQtvi7irF6mgk3V/KOefy0Mpctm
q4ksDwGGjr2aqEsGYF6A4Rv9HB16r9Yz64pVRaqzUQAnq/1ReH6v6YWWMgrmTBIdw8uIFEvumCz5
AqZtYpbt6EGjQU4YcRfDmyBDe0fVmjBkruLA32wIO8WYjRDAHOgUY5CdE0eFUvgXMkCcpBBnQJqP
ml+EWe4Zg/vqY0ssP1XufxCRKWFKbc6AcY5SoNE9uBNRTQzkxoR60sJ3kXobahvqx0hrtXj7N+x6
nWnVyRIDthdUeWyINgRmLvTdLJumyFU4s0ivGtp+SAnuqpWA5le9vyijCTO0nohJY6V5YifAEClp
wrqVNsNjTO4o0vKZVgpJkKT5anVmvjCX/yFO9AvWha2w+2B224gLghLAv1hoz5rprJWCYqyeqSYp
AQ4/OPhCPAN6TYbl4Kivu/JCmlBgtyT9uWLGvszl+xHii+DzQ16x6fMPGs18oZCZZQjuRjESFFAF
kxiwZ64ItcSwIfFuodxm/PUKgYpcg43AIRrsPg34DSOqxTv31Xu+k/PLAqQ4pq4hi6Az97GANq+z
O96hLC+HMNZszvN0ETN2jjVEMynLGmnQJaf/cApyxasb6xTjFje5mQtOrhfvG9xeqfEznUQu8rOc
Y/ql5gor2vPFIPaYzL/av6X2kTKkj5U+QkJdnQa71pME0V6r3OM2P91F53XZgEQRC4f/dGCi7dCS
1XVqYQMk9chHHIBOeYWr5X1kJjk5vQEfZig4s/WW2yuEzgHkSRMp/xVkI75DOKm+FWrTM0KuS7gE
DSHhMM+0bXRd+Q8uh11wB2TCmmRwnVNYooIRlxmKgerTTEqag2l0lFhYKA7o2itPBCKpa8TRxi7r
LYVng/Ux9DEZ0ZisWHqIWpqY8d7yXGCcDAr0IDmUa3aRyPizATfLp3z7LatpwobhslcNJ/MMf21D
6IRY0IQA/UzVrl4vhitEDK9ZyYMRIHdn69KTyZ8QVr7YubLQvyg/Giq4S+4bpgKyusW0UNFgUV0O
Vo0V2Rgukcy4wWn146XZXAzAuhinnY/fR6H9CedcQ3q2DkrU2kcT4r7/d2EOHE5VtrkUcqLsYLNE
IUSk7pMwMEhV/n3WMQ/u5GtzN4BMeSD2hvlxmRMPc6IaK+1y46fak+H/knydPOVjyZB5wbip159I
abRUZfD8JKKDT4OLeY2XcPTUEE2l96m8bY38TxXlVpR5VLLcYjifu7bGqGmkDCZRqc1r2zhvFSwX
X6bPuqBCEd0hywDQupMbJlv+kRVueNZeAI4el0rwBxPTaQoQgdUh4kAeap0waTsKyMh59ivY3Zti
CC3pb75u7u/l3pZdEPjr+vPmerwraupgkuJpZju40iCdgDD6bz9foGjAJ8nhpGZHM1NyLrBjP/EP
GSDDsvWT1v5soq62RUXaw79fUtx6YyMwFlNM/DdTI4adw9F9iH+B7bc26mpxNApKoXTQSspzv7AG
gIWN8oNteM72OYph63SV/7yNKiFK4fjmqc+Dt9o594HrlKLI4PZJvZm9nl8liIzi96atMvjK2r2D
0ne4E2qpxqBXy+WRKYFbcmtzJsNRqXQs2toA1rsGWi6MAyAxdoQuxOiujAyX9qE/ocwTTHnUeiBJ
OQ0K1DDMy1B2figJoV/aiLPwgD1JWKbJEfMisEzfcnMyP0ynPXeXJy00m+hWAAiZ7VnURj+2sER3
A3Wdz8h2WWwjLCt2KRO65QUrEbnvBhb1xXUqYZlykzFUPpWaGxL/5zs+IeFIMCoMCgicfOCNZuYf
nQaAe5A9x4dt9d0qPN3c2RqiLjXrF60IYDP37asLaJgIGVxl82fv3/Vq+juieBPwkz4iMHRT8y0C
L/yqak3ibLGlw/sJLXdRqMTwKNPks65vF2oD4UEgvsgEyXCz2lzPP4Xq0MBEoQ5gl2qVRlvCgyeQ
R5nGtohVE4L+LEMnGC1DB/5f7cWKhg0d0VCLNGwtazejJPV04LDZxKLTgXnMujrpuqNMwafB/OeE
3rFSHP5EOZdG9da5BtGl2HwGZORe35vMfDF7KuNpEDWp+8wNWBnvjTVewFzKuRWcZpBk7LaapRw/
mXhXsax41SoAO6ZE+jxyNM5OFG5vwNdJcHFEXLN1BohahA7ImlJXNaBzCO6ca06Rl7eKRhixcIqp
1SW9d//yKCNlkqDLT1cRTqCOi5ontSjlZlqjlx8vAb5EGLPDsroAKaWL8MQx3y6cFPhIqP9Nipru
5Ea3N3PA6HElZ4THvNyDHFT1WHUjC7Kp56wdbejJDKQUs0BEyfsQHQSidp7hijKqGs9o3wd7VQ/A
CD9wX32L7zxr96yffUlOVeqMpznAN1s/MIdLT3GlSYdEdSelfo/x5Bt/RyvoGoGQRx2ZI0z/4QRu
qAL+rIw05GpqHVdggzPi6pzj3/oBBJ9u6/D0RwNc+cRI8mmQlllK87MRcTmJqlBkISvsgATuiHOz
BN+A4fvTVRAxoCkjCpVSkYnw2vPh7aRyUp30MwKiNKgvy33jEsgklNhvjdwsmLTKImfVKCrJaNG0
t0+fpjuMjHM0otnuhhDbE0GWjKLVCcCM/f2RQF4GLfBk0ovCDpB25Ttl+YQ2/PcktoIFDw15q57O
L8kATgTqwiveblGMhkW7QrBfQLyEdWaSkoSNi4OUMtgV0AuC8/UKeKeGJeNdojSgcStDfEKp8mEU
CV3UhmdV3usEofrNHUZdsMfkgtHD4lV3AKT7bopG88vQZlUelH9g7Hh4xfgFq08EHdouw4GHQa43
fHpM4BZ5dGSlXt+BptrM3I3gQsXCVsz4vBa15lyJBUoC5O+qVcpT386eaTcIDnlxBbAAvCsohURV
Z1gP5Pypm1nlXbsQOwZhUloDt2n9xlljo0MLD0X7whfSqEcbJcFLVzJTDhC57lh4W+xbqjxnPhvR
yhQcepu8asapImSzhphTbPAqJD+lGkjMuSewSm8c7QXlMV/TovPkj4y0xmrkPvbI/+FUPb8dxNcR
al6SJcBwjU3JWUfj+kUVGTC6FZh0aP4m/lQdOIYA/1uk5U7X4CCshB0n0DzvRosyQO2SR7Eplga/
r8OMZamooyTGku+wRuyWzeHFUiJ002HeRINSYwyhSRVnTcz3c24OW+a7whUujVg76bJkdxVzuNR0
N7s8kl865TUU6Ew/ieu6RfFF1fZVLJhIYOy+vhcXu4cSS6fPaAlEqJW4X3AMAZB7sOF8uhcdZ/NB
IHARK83x+zjxsOWUUa3gtVQKqAS6L2VmvGBMdBaptpMej7Q6szlktnz8QhUGUf1AnXRVBCQf9YTa
ok9bOKu63jpJgUN1Jr5QLrAz62kLNXHjca66RIrWJ7ClOQrhGuzMVitnXpGvq7pehfiXfSvCDSvs
68ixk44iWBrG7YXFAIy478/w5hVJSGQrDIu3bqHUofbUOhMrQRGb5IuHMZnUGtL9oLyQYwzaE4+7
I5BEEvR48iI4zDv9yis5nCN3PvPcMegrUGOlbxujzaSYKY3MbpL9xzisV8TRmW0jnxDkZeQk0n4u
+xw6CxW2d3hv7mlUvUFDt5tLVlu5W6veSJDgAQiHZaQ+3rgpf01oRwlzF1En36sCbMKyRg+9J03o
aHl1MAB6qKmHegjBzc0osTgGMBELIjf2m+BCXQim3RpV0RUM73HnvA2AP+Ff0qhR/mOxRH/WeCKz
N31WaElXSLItgdJ3WJT7AMZxIoYa830zzWALj/tbyUmWoQAAjyVIDHhqTK74Xe1/AZMAYXFUPfuR
hrg1GLIDW6VwgljEGKbJAw6ZzfgR7wx8iDKCYYw1do4O4YZziSfnX5KtpYu/eTbsDmYTzJCcacEt
zEPosQ6baWkOvuxzPBJE0NVDTQJVW1NBHBiHqjP+O0D0hp1iqicUSnJZfuEOBa10+LZ2Ri+XF5Cl
3PP+mzssRjzaTyt9XSR/BJI4nXDztQ8vPX0rXMRO89u/l15tPp9aE6WqHnKX2i8nluMoQJ1ROw2d
FODICr03KGtzUzSXTfVdZkZefj74hdmAAV1jxabpxCmxXzSSrneII+orUMAX8MvJaZEcFy2RdteT
d3ZEw55f7EFYHEynEAaN33F0HpigN+k0sH6IVvXVnSLQF6XAOKlPnahsvLXcthnkJA/auqrNJHZC
0JWBSKyWKdUo9e7wPBTBGEwswh1Q3gVXMAwQzZpC4CvUpYCyWsSGteB/5riMbnPopy7ALFijLTvy
fmPdqZ6Ey3XGDmegXyoE1jEMByUHVGwwCH7z8HZVTlnFCuxOrSsfTCLMvlEp34JPAy7zlIbeq8Py
A+3DuIIqHcciVaBUrvRb6LpVPn43aFf78QtbgveGE1IwFaMnk+p5Q7sn0Rb4eresDOS4WwbgqvJH
N45Gt8sBtsD4COP29rcrILdeuoFejUqYlDOZYzZhCulMffaANpxLebxLRsXNcEBuDvEEDNTyszxp
FdcAyrmKnj/oqtaogi6tvKbVD3itGH7K710IRXUjTgoDfyQTOo2LOERYNQffyuz1Kq4on+Uj7HhV
PyfPRia5EGTqUmQONMBqxxwNiLzmmTpsKSvxtwsLTvDvGaAOGRqyeD5XkPxHaM1YjDaHv5MI6wR/
9K0jZdRVuQKDaaIwUy1zkDehbEJag97Y8C4qnV7NYleotdo/d1bQGdcKWy/xltnXE1J21wCGyN4M
L5sZ4xS/HIwJLoB8JWPqCagQwdiiFMU2B+7GfLemYNwdybhoxMfmKHhVsbv+6K6zNA7nMrLjTSvU
a/aW+a7hkeZckyRNup881Bjn+kU0bq7cpgGUVdlskPsoTikSDtZTgWvM3cDWA5FFFYtzn2HcK8Ay
eoEZVRYuJ62u99350SgbTtPWgjusHVaSMd6wA1g8Qy3CmJz7qmJ+riGoLsHYwBe4NOEBhAgbnlL3
sJysDITGfnX7n3OXiuSzfxCW5m90GIXalBcJ39rvOWvDlkbJyWMzRs+JW4kPehaSe60TXGF2yIoy
4DSmUWh9UdwPCu4pDdGQ/HZylGsHRamXlrrtpzW5+VJR22au7Oh9IPKD4b+7dmGR6H5JW6A8YISa
5o6Sc6tF+meEqg9YgjiTtT8UAjOlgtMKVNwrggFnqloR6SWnTp0tY8A77MxZW6TzlKL2i8hG6hf5
fDPA8ptlYt/hoZ5cEjnZVJQCZJ4HLP48F043S4GGWhls1Bp7z9w5dtgmOFLK0LDwKH9kKMLpOEgN
g3nLoHwmd+rIdEmcz5cTAh5UlyvzHJWZpR2nWfzMfQ18/dwk8XXNM9euXFoearpu07oNhqdleFvo
kR9Mozbb+6LdzM5QyQKHaKSekT3u4u7LRykSeb9PHEK9g3H8iMb3g8mvjeYBRO/kyF8I6Tg93NYp
Nr2benHQG+9M0wXyZIIcWJQ5JYKbOxbhMf/56S89LrsqPi1KQ1iEN7nQzb5M5u2Hyu7vgbXYBmao
GyzuBQEo1GqGcB6Zfk4HPkdsh+3UdEA28Jd+UVHjkwfEwd6pZumguGv5C0TssHzViTixcVYA25kZ
pYCSleWlSViLDjfNPY+7MsSEZfBbysxpr2GkSELnBznp86xH1XXTczOMb7JHQmVxKKVnHv2x9GkQ
AlNdwt9I5VwLPmuUuHiB5FW0+nDG9oFMh4y+fNcy7+dWSkPG/6jgbMpMeT+vNv5QRxTyy5R/7Prw
58tiYyAC8qo40uM0ZddYEH0f++jR1DahVtrfSigs+eNLJqSfnKPHJwFoE4jjD0HECaiT/b3TAQm/
cf3LAd5jp656SEQJY5FsQBHNT0pBIg0Dx3zYXU8QMFmbSFShmNojN+pmBCnt1dyox3IjWXbn0rfE
Nj7cI9rde6jORL6sb1qEJhQocbM4ZFCkT10NAotydJZWFOGHIzvjQT+a/UNLT4Zk95o/i4NqeDyM
xf0YaTNE+bYsI4pc4H7HsQBB4s19VAQXZTTlrgEF//kOXflPn6lpo/415UBXYPKeVMUsKTuSHC/E
k6SHw4EF3/UFDTmTdi+XcHLWjj+tfLFHnV995C7USYumtLQIo5l8+z5SUoUIwATR5GIkYgEZ2b4J
zhFSE75eBGSwocbxKPSEz/HBZjB5LmArLnkJtkbval9PsYm229Ovh/eevDFEhMP70VWvPh8w73M1
/fI/Cxod+NqKPIWgiyQSp3GnaQVdVeVt2CWZtlvKmlR/Uh2uFcQw3pa2HXIkCaFBg7NaGH7wEUAG
X+Os294pwXKXeHWF8M5dwR9amxhw/e/feZr7I5OWXSdNvscQA1Y9ywB8VsiS/YMwNTKc2MgZesZW
kDRuMpF/s1Pip17IL5mE3Q4e+2MYX7OvXtxv5EQ6djkAWunWDU569EquTMm4bIf+in2qMwyEeyG2
fjE1e6NEyiAqKVAVwBqkrgJ3L1Y3JhTKwURjnRm8Pd5/ztnKFAjYrtWLn32KKcLeNqSu6T+Sb4dd
b8LJeeRUyRAIMJ+uV2847FzabsXsKZP5BiGrGiPQO9O9hfqvhTbu7QeP2qsB7X4ZvfcNGLZAxuWU
ajZqvLWJw2QEt3A+CnufgRvKv6+hY1eBvGb0QS8jxws6jtwyS5fYAG2pTEAynPZKtlEOKIudUYHS
mcMPl6RwXO7MsdIiKHl0tWuTWfPYzhz6UoHgEO7mWwGWwkQpxszGWAlxSv90y9PUyZOrdbiaK83Y
rIykAnJJiDZrZtBzC3o2oTtcdUyiuTBDJXGplhnWn3gfQqRfzzgJyD1AQWK7FKLOAexYwldp2J2I
XU6WDjuibHPZYlRi/LsDHh8QxYT5SFrlb8iWi3OsLsp2KcJ+GDOtsbu7tpyVTGB9DKMDsgdbqLI5
QCzTUxZC59ehJaZFoqPZkX1IzlfBMN5AhmGb0UP0wzJb6g09EKLp2SkCG4db+JH86Ch8Et89vWkr
JR/ZJOe4iAq5DOmKuJvfv0vZ5ObSG2WE//k1ZA2qSjQAd657bI7aiNMBZqLmqNn3m9DFllhAYwRw
6Ij0CnYhvHsHaWkCjRcaTO2RDFNPD9B++W1iJgGVL6IVzaSHeXEZnH9Rq+UBsUKQMmas5l1phqVv
twFZnRmQHutEj99hfVHyBj/fha8Y2gqNn9kwG4xnFtq+toLmGv1QqDuamPLBbHDvakAfpceaxFcD
i2D32D82kc7VXGmDmBxP3q8El4AM2e5+R1Lkh2C5rbCmve7z+Jv0VVWq8jXlcLgs6R0KCwim7bMh
mwPR9vM1QMgwUVG3oERy5idK1UTebNGa+JxV3bA6asbfnsr3eWNKSo87vePkCbt4st+BlfpFY0Vo
bCO0kcfOP5XmHHEA1ikYuhfsmEIqVYj0GfuXJ1XEaN+DHQMKnYexQf5GcvnV3aVAZw6WTBmXfveI
ikME4KH8NHxtLQIyTc6RVdCySqZzRUvnwc55mMruF83Aq1wW87yKpVHYDlH5sJjxzgc3r14GsPaR
XJ6/LBaQI6G5li8ETqC8xqqG2C094aV4cwSe/77fkLTtR6zzK97MaGCT53WuqL2vp1DfRmrZ6nkM
tvNPCBkFFwS/hTzKkj8V/qtmcmJDoERZYiFrYnuMpDH+CcPG6vMWobxYCAiC1oZrsTTVgH2XiuG9
TdF+Oazvv0mJt6V2XGBYhej0KchY+tJFc1mXgU3l0ixqq4i6T4I0eL48Dl/cpuAOXpQbumZKmMIw
DFnRKWs6yiHTOhHtlC3pS/HEj35yy3eA3W6BwJ70ilLxTQKGU1BbFh4K1Xg6YP5x7SUEAiNXr0hG
zbXHawq/+OJGq6aLCINLEYmTjZfLQuSi1RzAN/axQIzk+5mjwJNdbE/j4pmeiE9dFmJmm+akErcN
azSlpSfvp9uBimO51NmG1hnynkig7n4kIVXVK/MKvhwiHE36VnZYnh3bYLcRBj7BTsEUhQcdLlpK
sF1CQ2k3Dlv+pNKJMflA5BuVHtd7ZOGg6oxyr2iOMy7ls5472gUUEi0ZaNnNZa6+MUcFBkN+U+xg
fEWbGw+Fxa5LlaXbKB6SBPRuadcEgsgQt78QPnWA9OdZH2hi6xpZG/Xe4/OLeOVyBKXahbXitF1l
kNrzbz+Luz6k/DG/z1u4fV7Ftr1u8Y+r7Rv4cfZK9NNk6HigkFXVHDHYbAf4MobWGC4YipLmPAjr
UiRMJg9NLbQgSJTCemQ5n46sCDPg6SDXqBWkwhLufrKAWnHyB3+JGXjjNGhBWeJf/PveA9HurHmY
wwO4g9yltZrcgQlh5Qd1m3O5IvuEMDxK+DKAWJjRA47CIwfw8Oe5A1skY7vcZ0TQHAsZKN+30ZJb
b0kvY/i2yf22ZJGIrXIyTgtArSa+ubv7z6Ai+UnfqhHdtY+3NRZzMbZQOtjSSctW055OIWPCZdqy
8dIEho3chOhshweHbInd1BtiXV3YH1cOo1uUFaJOfvIseg87xSVAOe4ZEKHZeQxwN6YvXJNMxFzu
b6eGkIXepqI3aTeZQ1WtJ6+jnpHS3glQsMPXv202K6qG2zAGKTgCi0zwW/v/IzNJns+flG0oZRti
zTeheCAfxG0fFVenvOK//wsRB9O+XPMm/ig3p/6nPpWMCTO+FlaoOfQCLLmF6vFiyE+ZVd5lnoUY
p0v/S4bDdppO6X9V+WFQ40Ak8ZhJVZW0CNLY/DtvJYWIUtgINvXf0PsAxj1EUzYCvlki9qDHzIDZ
Y/FDUHNgYBrHAMkdPPb7f67e/X59p/RL9y+8U50HZyT+HZSctDu/QcCgq4rnlH8rEsuxNBOdr0j1
ujuiGnre68nUAWxYiO/3386Y6o+vjvKYIkHlf6Dro6M5hArXmK3sWzf9dp69uBvZ2bHZ3Y1D6Gqa
F/WWJiyJPuGAJCHVTQy9F1OcghFcuBJ5M8HzmWXS/Z6RM1RgRSFZrudUEIGSwYrw45ouo/Wx3vcT
wzwZaw+jxKDoIkepVyhgSZuE4nKZJE3GhYr5hP5rtjv5Cr9plWFP0sv3oqD6BwzD6NPOa86CDh7v
72a3f8GAjEa2TSMGDMyRSCaFqh36zdjmfD6HcIvOUIOoJ6ZegJXow2mjSVHk0XuPf+9YhY8WFP7w
sKEtb0eM5ocIy7Av4WrONmeDIad4OSsfeM+4Bx7mua02hwGnn5sO4HqZlQa3domPD0iu9xnJfhjZ
c69Nab/a39XpeXN5VMunbb/ReDONtUbt9W0BOTKKTJE7rH3ccFhqvvUQPmmt1gw+dWh7ixf2IXX1
pKG+G5Vw7zDEW9mehmSiq/vllymwAC8tpdhm9kPA1+6ORzLuwk2GgkKDgG/W10x7gTT7zPFqjs3x
bVr9BxlmFjUYv5GwxHr7/Hld1LP/C5GX14gdRhb5a50k8SQv7i1lKvAcjiGxGEEJOurhy5l9XsN6
r6k6tWQadOrmGxrruVwXbno9K3pobKbgTSknmL3v1rMtkfxb34atVn7vP8mvaUZ+LIQitCTW+HzR
bVavGc8xHSYAoFfLu1aThYdSWgkegObYOn/PvLLpl78Bgh4EZJ6fYzXIKBB3npFbiqngE08fmwj8
+202x/3RqDzIDAtTu3pLoCcPP/YHaDVxzPSXVn5POuoTE7EHW8FZiuQskvxwOBDNKMVdRBEWhuoj
79Dkb0/jH3u7j3fx+rOTkjQwaXg1Nw+KBx9NLD5knu1k77K9rcTrGQeb5h5RyRJcr1G2aifCzbiI
Gl50HIXMU1eAp+Onl4WbWiDNcyTIwhiSRs1f85eM1Rr9axo7hO2BgKcMd2WIZNXgKz2dXewU0LXM
K57pIAypXxz7+Xjh5ou0rQ3OAqJgxr1F6qHecEqWWYVIV2zEzMYyTDPBPLJSapF7WICJ/q5W15V8
yQiq5j7O59lmZn6SEhGdZnIgam3sIcNeAU9I0vve3Mt3ubop93xWf32JFli4jdX6gxL6iRilB5AP
isUq32XsxBHDpUDx8BsC7EyxYB8/xucTnPwJrVuXrDdeRzhUl3WTmJXRC+kH8yAirchUgbH8Oc4p
l0f2aMbpbKjhpBtT3jhjcaPuy2RKheQnjO97510MOUrUts2V5IIf3bTdm9wvn5ueiYGlaGEubc2y
J0wrPxEJ7f8LAr3D9MDy1GPPMMg3tttIuB1yB3h/b2Hb9BVTwsS720pYxxUxEHZfJnmAeRQzvw6Q
dJHVBJKIROGJMc1i6KcgrlSGC+V+nniQ9maHPciRlCMWdIAgKjt5H4P2S15j2IfhuxtCJyGO1DIt
LgazawcMQOUwywN9xgScr+LcoS9tFDkP0q4jRZ5Joj4BoIv+qCExdgPYE7xH3d1mR4vVSojrN3vt
RXdunO/EaZMtuNyFbfFRVs/FmL1n9K973qlHz+CWJxctlZG8lYjl4dFgWc5tVlUJyDe8PsjRHRfU
OBLWKiOEghoicSJT7GOjy3GDF2o7VuiplbtiS7Yz13JJ0m/v989ovBT0vSjaHS0+YpT+XciLKVMp
gwJ8rD1D8haQouPcAITci1gUh2CTwytOxNtclM1D+RHeR6eEaceOGPg8u1sGjMYxmgxBVsK7X4Pp
3HSU2qApOlRgkYqIEr2P4EwFW/d6ggK7V15cEYX/8QE/Hrfy6Nl+Shzf+t87IA10T9nI1TQVodZA
rIXNfyoqv+56nypU28hcvvlawKoMscMjkkoZX1BoNfNNRhGiI16CQv/gBHcRngysrjogfwn88BY4
fSyzOR84FME/WLX50jxGsoSjm98A8Yj2vNi75h3+7F23tyDw9h3lY1sCKEJK4lwrEFeNBFzbGJ4p
txvzKPCFAWPNBYkmxhYxpT0GdZVIXokFzm4M8Q9K4KM1ZVTeFzKDNd/uLaEuT4Aj4j0wFDjs+gCV
EFE5ZbLv0u31esYc5wpSdouDsf1Gj999JDsk+rNafTb1gAKoTkVCU/RlR4KA34+857BxQr4O4RKF
9c6Pz0bdlHVJoRKi2vSFnaZzkdiDC7mYy5W36r7f2KHJuJ9j85KjcubyCtt5FsPaHF+FH5rttq7+
VacgP+ceZ1V+SV6qDaPxOX3b0NyGjDC6894F9C3Lf+Y69I/h/Kk/RbDYY6w++jIS1xW4ex9l5TNP
sCBjl2MB6nj5qv6VNxdrB3kbjJqNEGdWflLYONS0i/T6EdT3XIdsGiFchAROYfAQ5V2Y84aOFAL/
B0633UtJ9+4j0pHeqOrO2CPsXokxmMBCC896rH1DeAsh7P16uZYzDlhIbJPtd+r3W/gLGR/PAdOv
EC7bXgBCo6LsDrQuzOfsLm4PaZC/xppfLH6DGndTBU7JgbBXX69pYtDAuctrm2KXT1ohdeV0EsAn
InvV+6mMGC7tynhoh/5QV2SqGsGd/5D3O2iQI+RQdr972rFY+V9uqWf3acNiDxAUFdaY7EYD0NHv
2D/gzL8SrNyA66LosnXC2kwKMZBe6NRyCbU3nTBv/kprB0uQOAUM960OVqNZP8Glvqa3gveCnN3Y
+2zmCHt67sy/gZ9BndxX/zG9NYojylkil6xld6p2rhv2uR3eUtyNiMu0p0O0FTOq57ZoBO478ZJZ
7Dqw7hbGL+TTJsf5r1ZzYzX0w73g0oaeFzFSrN1rOeA1JZIcoQMP6nb9OvM6SDltBmwSnmCm3Mh3
KlqszdTTNO5Mh6nBxxn5lRqQO9AbbQaa5LXMvUHzhrbhXv2jew50z2GCCec4I/hdvkKKBwmnxBeH
8EinDhLmaTZQ1LQk23GG8kkgU+141rsX9golwlXEp1WGYACX6t4GGe3E/l7kkuzteAMA70yKhFvH
dw237wL8g8veP9dpnQov7ylD+tUInN0g7KV4ByThv9EEvnqezc5QPhfMzyrpY+6J5a5CzhbKaPWD
mGvb58How/UErJbGmgaYD44rceeuuH1ir2N2RoTks1Npq+BDVsRaLo1NxTQfS2+K8hFT33pbUz+y
d5FF8B48o6v+KHFvA2g2rtka/kx56OWffNn0SY4x98l8f8EUgVgnyNW9Q/fTzUGaods7mxbTrLVS
oxnEMZVceKoB30BPnc8Qu214QEG45RpsgqL+3XC1a6pUvSzParJvBfPKAVTLA5y0bYUUqg8V2NYo
GNHi5ujSAgPAx3+DxAkydJe6J4DsqRZtJluE5x7+0cRoRHgXG0xrt7xuNnVyjFJGDnwEavQnZK64
yZHg994DxJOYR4BbY3jQjwmIv1DoCJXMfwnvv0aL4DRncUyEc+Zjol179wsCPWWipCXEKAyUcued
73yNq2CjCUJ1ULRMlNltWS14Ddci91ehUYlop5zZpcL+dyNSkjTRXV4x2CgvxqrzyXPUET2qvxZ9
2Y3erD0+nsrRtK9F4auVBBQsIeLl3xVEmHxzZlAMSHDCjOE1GDlUR6BGNw5aI/9M63kEneUAIFsa
WG9O1YxTUH3sB+PdASn5UT+u0IHStdDybKkAm3DF9vPU0GEybam8HAnfFpcRC3/6E+pHiWa8UI1Z
8PZVR1ovh/pI97D3Jpy7cbRJlpZg+vAe9b6zuS7cliKuPgmBDrfjDOIBPUm9AAi6qwGL6NEjPNXH
KWbDG7zVo4fN4bILKFcbHdL5wLiC25/NZwg139utlzj9K5tY6R/Mmbj39PHMaKEE4EopF00PoCRF
pg6izi0JpLGsj5x5DEjZoRf/KtDfKvodPuJonHQTsuRtp7KMJw8MXZWBnwpaMIu3+1Bu4lstZdFl
BrJjGk0tNE63bd+doVYTpf/1kXuemJMJ2p6fB74iEPx0F0P+FZQ+ex5kevMyBfDPtnIU75OJG9JO
YtgXdwEVsBmXP15LJoBTwVg6nujRP6ZDznHJigQH9Y2UDDU6imHLvYL511liF9qo3TEk18jwJlZT
Qdazr4s00sxIgtwMnAL2YOQyrTTIgmclQXgHoM1jTaNCxb254mwuOzqY8lHVKdmkEye7Vt31jObC
Y9wMYr1Y8GF8D5eRxAEKZwAxl9wDVGTt+BBhOYt22laIqJWLtICT8dAt+5RY5JiLZh8hWNjxEady
ogZ4d35COtXIco3qGc1u0IsakvH4yVK2xGTUoJo4mgcTmcoMfbPsmXdUZcHsrodNAs6ccK987x9I
pyjtbn1Q8OHUPrLk2/IMFRA6mUwo/Q1ykiJOPAcHnALqUh65ZR5CK6vQiCKmpRgjfMW/CTjxZPgn
D6cDunR863jor+9PEa1ueEGFKmVWh6od5GYoFEV2J6NbsZ+Yq2mJU7BV3aSbVs6U62/IR6pJ/jQE
ANdBhfcyU1GiwjU0Xh7Oypt7naB3GD46DFxUJ62cJrhs+SYUAuopXMdVfgat2RMs8XN8g2A4h6L0
cQ86Br5e2L2cZGXGn2tEOdgy/FKXr08NUlppERmzh3PT6wT59mVS5GBiQErFiuxKaWXSgypds3Ly
WJ05DS8d5cYlPnbfCaiPLu2GciC3JQFQMpIPPbXgt3tRS1XCSdMFFT/Az/5/cmj222MWRCI6MM8x
koomLgJsOmK1eXfcRAlY7Zq8Trvb1rF6orl/GcXU0FZdEgFyk3B1ZzfySIh0SUrFT46cgWlMOnTu
Q0o1WpPtdpUaYiWnp8E1pvHWIQwWXPiKMpouDrNj6zqhRPB4pGbCNiDFIqWD7dzRyrVsBRXGmcI4
9mjT/vLiMcHeCEJYewXZY19LOQDXx1H7oxtPBPUvBJtLExmlIzj2rCJM3P2IEiGVMJzWNEiRi8sM
neKfk0geiX/8eOapoxKNogpTAwr2TwdUSEAgpDt7ogzUEg9/46lyN93B5qgikzhumE4d5hk20StL
S8cNVyikSOHccvjl4Kz1RQP6/ngVLTMefv8qTyrACqkapBY3V570C6ranDlsIp2pGH7dVKb55qvG
exSnjL5ctkBFmvhjtEkn2YU5u+rAxhdTnStT+yDyj8QafLKS1G19VBwJf2+4TThCOLBb5F/qtGFr
sJ6RmH6Ne+0EkJaH3ssAZVnjchfNhN9VnCxvJCeG3qB7CEo/6JDQRcdsNspaThXTzxajuRnFt2ut
miESI+fCwKT1j7J5qcpvM46PRUyv9Y1Mb3oOKOQqJwJe93d3rVUefz54TdtnMjKBnP+WvotZfP/b
Kjq+6D4ES/7yIByYhFd6IoEFHHnP63X6xsxnucdQhieWldOle9jHRHlecVDm8/G5gzEsZ2eN14XQ
tNNoD6XSA3c4VWxETOY02amxgLzqYk+WjZDjm+cqid/JO5cZUl3UXwAHdYYOE33K/vjHm7S6eJdX
3NdhlnXiXcCuxsJO7pME23iEqixEvLlh/QjUM9cEJvNt1MlJE9FJqAlRMpJIyxsl4Oea30EfMiLQ
h5nxLFdca16suwQGbDMMxavOQDTE27LmM1cIlcyMCvVgnuVzxrV0bdDVsHDN3Tkx6PV63CRJ5IW4
Yw8pi8y6zJFh/D9pBo6OHScaHmhQXLSkV0sVD/qRqyemf3jR9kVxfy2fU9FznTzbiLjjsVFTWJya
PdHLm4vr+okVU7c1bFXKUo75prVrep+I+kgYDXqEVCl5Uz0qYw+JBKpNIm6LKJkuDB6y2GoAZt/Q
B0I4DntRT6dDr0FFssduxPjhG2JV5D+YUL064xmsSTC8Tj+kVeaObHx0ihrGPJFx0NDeljblLQuI
VqTr8vLWMlUOUd1gVlFU+Fc2nkhTCnFmmOgW/6FnY8UGbiVOWhwlhhZ+xBKggNSbx4gQt7siGEd1
ZzycCkarOv8vAT2VKZtcHz2UxLemcY/2G/hqdQ9alM1mdNUfnDYWwXtRQIqPOxkx2+Ak0XgiidqR
jcCdMy2SpuI92GUzOZi2xRaEN0y9mEcZSXuN174yDY2MQxSmKelw3j8/LqJVvX6acQtjoKQBBXzr
2ursEUZskuzRp6RhSAag9nVprJAnLlmrSucSaa0hOLFDKMvUkQfmo0R5IFQ6+4w4oQvEMxZ1I2rk
5NL5Nfl2oJpPLm81IE2NETJNhbZNs32TAEvHFA9+R47wxAFX3Z21NdL5A6cPi8RYPrfpw8fPluhQ
GH6G43VMivie9ua8rZY0yVQyNNJlsvTRpjhKzFtJkSCo5qoJao3lnnsrzncbcyHXIcHAR70s3K17
z/18+Obi6ViGIAp6f/7ufJw6lh/gXmXua84uk15povM49vzrPQ35zMjzurPhauTIq1Rlu6dO/tp4
rlXBLQvWgm6pSSY/Q9xB8XvYr9rXDlbGzLaHCuOw59PDpitnlbztXVFSVfjeDVmJEq5VAYHaMAfN
5EfKoXJY5Qo2VHHCR9yf+jKuooGfO57jAY+9FN/hiemJJKjUiD+bnRUI20YOnS8Mbnrn1E8XpXLF
GnQt8mwV7q3k2r5R0iuXSEl+yw/o+aWaNgv2QbMQL6yffD9+WurrAV4RS64E8vi8IMvCAvzQHSal
p+E6ePtx5DQYcaiHjjlSxz28smQBnbSbEQ+89FAWdaQ0VMALuY+0n9dxuT0dBQ61fY87mHLbeNPS
wqq5vJE6I2jAnRfSAVg6UdzXdGsHOCDZI/G4tph9zNm11rwd87KLF1JZE3wwJSv6SQi3vimw+LBM
ad0TBRuAkFHVA2gks8cfLbCRrMhojoj6xO4MnlX6IrPcF/hvjkY1Colz36H5VYCgH4egL1JatLk9
Ieo3SqKnHB2TDdkXwaIoNY5QKPVuLoEmIuOVEF/1CkmhIYW/XnDlGLy7JDwlpnRB9eXun6niuWzL
NMVp3gVcUKKfgfKIi4AukPdFaz3qp+eIQSfVXXA1OQLfdpzSTXKqHpdHmDRm6youLvcTNO8jVUe9
ZKrJEXW/z0GrTU/iGfdKAyJ2v6rcbsjk9cSzkDXwufI5TgsRAZIo+rTFNyRM53aqMFDq1dBtj9++
I2VcWXygGReOnvVlb2SKptlwXw+A4GCKodTWNGWNNK1ouOTblRPGx1ZkX0pLSIKbwmtnaBmfid2D
eS0hRdimIZHSgqRUWn0LOtRMyS2uXp7qAC/XvU/jOa8NKDN+OLpBHEbY9cm5JFNAR+Qpw9QR++hP
DOls+L0/Yz9gguah/zoQhIY8XSAUdl3cqQezsG4LRKC2R4q29q+OgcdROftCE97PUIHsz+pWsQ6S
nD1aLzilXWsHOHbRTQp/sSgT6z4nZcRvwDw2ER9+EVIbUnUoKOCubymrzN2Xgk27B/XscWwcVyuI
xmH1LEm6OVqNXWdKt9X5gXDughf7E71HVZ5lZo41JWMGhlxNR86n18lGY1IFCh9DkIChVgPu7hdy
cXUEfdJokrvdHTuzV38t98k83Ll2h+5e7gHsWgXsdZ6dUI6Mx/bSqYxjGLgHEZpTaWGbUzdmfWUU
9sROM8VrZ4zbEwQ/Q/aEt93W2xunS/x8LkvdQLFECrDfdJ29RjxohhpgYVlQh9wMJnw2g+ZfTtpF
Vu+YGKwbgTbMa3rVz3oTMZasXRI18NuRX341nFU+1eKzwUdtv0gnXVfuqWG31n52afJuOKW5J6ua
6dyqX2IKKgF+PRMNwXvLrYXWhauEmunWCb0bOiV/2gQEuYcUvblaIQpeFeIGmtFKleNc49ge1O1h
FvBaAC128ZcFz4iH9ok7ZYQnZYlI6/XsxSJxCOXu7lSXE5qRTG7FFxzn5MIvwxnOF6U71xZQxi+h
ycpqPzJ725Wz6j74KTQvJ3KVFRTVf8iOIg00nReYgCTvSL8lcgtJiYFLYSusMXnvpTdlz68zw+h8
druSnPQYti6M9+v7LKp9H13O1u+DYyKwRHlp9flDh/gm/8AtUUQ4KZOE7QdRGisNhbir+0JJ5qjj
6Q4x9PfToP1o5MewldJYdlWt4AdoTeU+4vPTDVGNQrXinN4gCp8fkEJrvXQb9/SnBOxfeHmEQf6c
TL32komgn30nLMxF4tmDwgReAbhtaJiQfsZLg2LFAmM/rvL2UgXzPkxrxR5FJG5rMOzuQ/6qu9ka
OTyxUQhRkfBgb7B3d0WliJTXjFEIHgbTB/IrI4yiSxucgmH+XgJR3dux/Yy6/RXY5R5ouUxXPgZI
tZHWCnedI6pzsfotihEUdC1J25pyDyACPB7QhIgp0NhGOGGrwBI5ghYlgioZf8IlRE0LVIgiuqMW
lnwC/ksYRFNTtq6XHoa0gUrzAtBvtgJwaNfXcfgU3lzBR37EaahHJRNRGb0tnS7IyDomsYekRtwz
i5yh8EOl4HKypKPJUCAGoYByVFT+l8m2UE5QSj3vBu+xS4pTuJiQTkQV8S9HI4eTBXgoLtgQCj5m
EJaNJCOVw00fDbxwlE1+y1pqgql5Q9/HgqwEG+mGSibz85LyYMINeuTJR6u9fZgU2EqxzgYL3rT5
fpIizPLaVUsfHkUForg7xoWkrrAwOGcmnEKbkfRJZkfs8r2SoxDVg0/byoToLaiTkl5dH3LVeYaH
OorInPQC175yHqbfKRYvoiV8RiEuy7Mb7lxZ242+MHrr6LLx8iS1L0zkHkcKBJ2NugX+P/9lrkT9
VWxGnk3xUk2q/RBFp3VT7a/SYahxJOSmosPFKQZjIbzyfiNtkSMW4e2AW2K0qlUWb/fgl+mKfpAC
AhT+XL8n3xiP2pp5bab7DSrG503s6aRyTQ0POozzL3SNGqUiiPk6Kc9/+BjIFcjfjmWhFlo1u8Rz
Xj7jmcTkoiEaPiOHzCTaYuDdwsOWmppQYtIYFoh2ClHv+hHS88vRzBkjAsdppmoeqhsU92RCITat
yQL4rMFW2p6Z3F38SAn8CrVUvitxcQwSmd9fRHShEVEB4dLevO09SEBq5DdYXs5ehlfUCBEnyRS8
6bm3xOj03dQ4dQ2J2U0+c+esKZh7a/4UzWH8Q8VZCDZXaJzg7XhzYNghkAh3R5SmmO7X/1xxeqES
7vMz1RS13QQtHkw3hGJB22S8tWG3/zTVyGJKlSJ0HeuG+O1NbFRsCE8Yupij73nvgO/eqRiIdbIN
fbdLehZWniNAIQ8s6LL4qhRCu5VQ8pDViXCoC7AZukquTEoP0HDqCN7hX1LT2AZwJXETH6M7H0QW
mrpRcKB4CoXXvq2vqgR7Ys81e9+wzcT4lKGNyK1/oKcs648EReM+fPt076DHR/81KEa7JPSG3Pqf
Cvag++kDKsXK8jH4VDwN6Yn/cJtEKCyPpHOFbZepL0MxpBuUKgsL9htHAwTNKZOzJ60a8G87sNI7
X0mU4Utaca713OmjE+iiKIq9arWO6IoM+MXJdh52SqVA7B1wH6TElrc9HV3KoTvwEEvTPgF/grqj
sFcrMZ4zDn2ys5uP75Ml9R1VVuM3EnhzUFC5LadIZPyZZg3q6iMlSURREm7Bo+DJgAcnnbPAzPcz
NcaEV2k5M8laeuQG15UElMJUGtaE838fUfEwRckOR9mU4f/Trxwnl+zfb5gI2BoMBnm1M/wDQxgD
hbi74+4/ykByDnDdl5sVXcO347OlijUj0NAxq/2mXOZqtimt1sTj8E49fl+9fLYiA3RiJZh/vAtw
kuhRAWd2upThwWbo3+k4admxxD6kiU9D7DIXKm/VzcQ1Ph/5Cq69Sx59zeyC50Lj4KanAfPj/0i8
h17VtwsyhxvoLUQNNm8j9hB2pxGJFt3YuT+BgmST4bWoV8QAmIGNzpqZBQNrb8iK0+o1YYV8cof+
lNmOELkAlW/J11yChliuoQwYzkdi/nhH2SJlU9uImdMl0ABWMzx0LZ7GGA9ucBQpUn9RcF8ZhvcZ
V9Y38iQEOH2I/a2xjgxGq1Q8Wk6Dxv+GfY4cdcLalX6Uvi7n6SoMSajKg8j+i0l13dTzpijq+tzu
cgrWjK2otN15rO2+S0SMftJjiPBweUh+tBQAd56s6VnM/IqVeNg+ZVmgvOpn0o/HqGnTgPN9FiFi
SuPmpVpecgkjbHrkXiWvciWlaB0V4E5bOYOqNE83FPB9rMYGrlFHeh2d/8YnSpt7BtPoL6i076L0
OiKS/3RmfEUwj2uncpyLgyA3H6aeJMVZ9KdoTl1NF6JWw71J5+dqQlG/Rh3j8UciZ1StdfCkAwI/
V5MtZE+AjfhdGerOEM/hLaKRvh7u+Ka7NFcglYZxwQI6jdYlM3XqoBNdEXOyR4e/qw6PJNfxppMv
VzfWdVo2LZdRCm794PtjGhscX4Tjn8x6a6KT3haRJA1lVx6SqtRBIDWO01+8iE2kREOa/y/ZR82t
dV7ywlY14oHcjSBHZLleSTDXEsVWTNfvMLdk7XgBr/Q6fAb9mcl22rBTTmy6KxH+kUUJTjuxMgUQ
LcUNfh2jm7+SrqakP+5ZXMTzrCLdEh2ejGxEbn8/qmkdIlL7IibCf5/AGX0UimJwNk2fe2EPhA1x
jzyYJD1xloUJ9Ae6sfUT0v9IHv4AVLJl5dI/YbVz0JjSvhCk2CPvO947+rLGQKOTKDT6ClMqwdOF
d4+fBFnenONyyV97/YlI/JclWrc4S8bCZmOlsmaL1zHwnImooinFVnEifMhLlAwbev+KzTZuf7CB
+gnUWrkpliGkNh6VVR/1oUTF0nVEQUhpbUJOEc44T+Io+eX9XsCqW1ewYONlh6Hnj+upz6yw18gV
xYGavxkl+NhLNIpN7KQ7wkeXmxQZiWUiqBKj34h5tu448niKTOy8Nf2Yn/nbml0Koq169Hsoa790
Gg2V193Q3C1O+6upZSK589CGhgzaCb8j0GYCjNNeXzvD0dsQuvXuot3H2YfP516pHdR41izuRG9q
fYPotNy/JjU1t75UBp7qm4PZT199zv8TiD2Mn+xmlTGlqWVOuptJu+ooy9Ctu3HpwufTcn7YUlp+
hstRSXCBm1mLzvdJFO/SKCKpJnuvOOpbcgqYDGW2LJuz3h+CLuc0fbHD3nrklVBaqmleT1RNvjnl
IHGIjn+DE7ghbm+T1FJK6eqsgmxAookEZnB5xgN/+8vnKc+8YHi9APg9z/EfPvIv42nmXcnQHfDr
ySbgPIDxp711M4qlgI2UlIBOKQOt/hATyldfTxxpwiDHs9jvK7mAiQgVwEDFC8WTGLmqPaA541lr
NtIT0zWVN9zE5FlAsd/wV9VnpE0MwnY0WDoaR7H+yhSjQSC5w+ELTg4M8WqZxiJ18ypK3gmsTksu
zxjnFfVCjckRL/WQakPw7xlReuDW/UwB2ATiFXmJiJODzOFVzKA3fK3nEwWeoryDFu9DX6wJxkhw
hwECx8C3ptlnIA6Hl77P5tUCuLOfF2irqF+hNUbfPThHvac7dXM94dlad+cHE+FUgM1YW1/Q/kDX
0asFfuI0M5ffhUsmxsj0J1Xm/3gsZZGKNfK4mYbySZ8GFxcDyTGWONa4JqWCbHr7+eIe71zFwGaK
GdyPZemXyyVi5UbJOxZCbgY8uejc6ezK1CRpYoQ9FYF/kBYS5MQt5rt/H5I39OhxOYKK3k/DESNz
VfuIage8dLLX7mf9r7lxQhNkssYEIPIRIk+11mpOzQJte65oBCTj8rsmybSOqbxS2x9vTGzLTn0p
+pZ8qbPmTqZdh8srA7UdjEDpuUic4f8di09ubN5HvNQTbnTc28Qy1R96EWRtHWKm0WD8+dOgwGtk
9EoluzFixhhCh+IHWhsH7PnUt4gGGjWamWCnwXT23sMQV1xxY8KbjfYLRLFfOL5HtmdWlptv0kCf
x33ZiUBxlWELFxh3HjDPWpzW1k/Iec2dPuPDTLygjJMMGEYgD8CSxujx2Bu9BexwBlWM8w8GMXwd
1mmLdaW8cpbE6MpWZuQ2BXRGQMftaJ4ypil6wT2pId7aXYWaALLSwS71vP0EfhO20OJ8cn6zldYP
SCK9UBrpFPiiPQvnbGDKKzTt+tFSv37YJ1+34RKQq4NMNudzfRtELKRCEJ0ato5+N+C4qUvdcYIw
iKORtNtCcZV8S+ENUDKhuAtdkjqXC/myppScmlrhwUrKU21IQdM2C/gUIjMaOXUwSFCqdVscINzI
3XaRt2Kb6QLbHIfQjrirsTuCvo8fARy7YG+XrNUL74NUUhRv435ytj1XoFAFRoE3YaLmHR+QAfiW
cBM1nNDG05n3V1uDcK8JbX37Gloi97WoBaxR290cF+b+UI4Z2DCYZZlZADqrZreUEkU5EZOOSU3X
imlojYtkCK99J0yhwJfowV4C7SBnR+YyFPLE6ryt46EUM/Ho+kVsjcKTf/T5pOcRMI80oeI+CqhD
YaRtfr4j5WaCHbfyBS+Ki5ZyKXAatNYKVEQZVDB8YKXEu8t6IU37PHn+83bp9X5fE7tH/VMK0g+5
+VKIQclOQ83AngBusHBe502vUAZiKwfna9rXF/kDYfxjTPI8Z4veFtSMrGZvtTXl4F82gtcFcMgc
YBXa8atW+vTO0yL95lxNNQdGCUsi+BhCmUyFyMS1CcSih+jhzzlkSuL3rBCsyiWKy+o5I33DfkX0
jMrPdymeJDQ6CSWqgAFJAsW8AchTWa5YZGLEizcuVRsuq+W8ApMu5qIksSklKW/8Zal4n/AMEYCk
LsdBqEENNqjEeuXY1RH6/zQoviAjYbFAFi81lIeP2igm2pmQljWNKNmKth+mbCt4KdBVXrc4FOxl
oDVHHOou8Pdvbi0OjFq4lxaGqoybzC7s/pJ4/FQaqSzsFaMmP7oLKWZg1D8XymdL++Y/AoD++z5y
+pO8Wyiwd0LKT50/ZU7CkFLSHviaN436/bi/2DWkYi1GBRrqqOkr+SCCqLerfY1qsPe3GnzwnPje
19XkSB43lI8MEK0OWuQXvWIZ+Nnkwdhro7ChitCyD4irVNt60JcCELozj5eNqHbfCPto3OdV8LxI
ugao7y4wnxqJGfUSBHioDSNfBCbidzWGweVtSDsvT2z4N9O/0AuaKSabd8CtieWqdEMDON3kXOhd
mOtvwik1kdLwvXodgjK42kJG5BbKTWkwzGVjprISAqZoT7SKZdWO2SwRo2UN9R9x8LMpj67w1ip7
VDI05IVj4XvigoOmJVXFWHTrLSYLrgXvF6saLIBWF63Z2+tlXQI2smT9lGtJxaYDDdrjha3EoYTy
1k4fnR6k8WQE2/VydHBk6HCyAvo6Q1CfqN9C3KX9CrUZUmsfUhXrqPq8EN71OzEH1nGq0AB5lLfZ
n2VLxDGphobJYWmAXV3nwLcdKXsTp+qHRMWT8TT+fVHALIoe3cC4hs2hLqwuf4ottTGaTaYdXVNC
rS80gCYrHVqj1RQjordqwaag5AqkE8sxBGoXcPUy2BB9lVVvXfePt7jhvZe8eLaAs5udK9Vj355Z
ym7pnkPm6V4ihUPiOvZnXvrNLhclobZOJXDha2hmeqZ0GsJjS2fjmEtK+pkQC35XwOZ2Yf1yi4ec
wTGCcLmwbSg9YFYvnMVfT5d8afxnE0PP+pk0gCmkmci7lP5oLl4VvJVBFLb0K/KgXRzXJx9LuilZ
bmmR+TpGnR6lbuS1UO2oIFgR0sLEFU3J6rN5FUN2QHNgYsJo74fQcaVtYKPIIm1x12h83nyltsbl
1VD4/TF3uDEvsy63/BooK5NW328uI/u+U88vWMwZhN1ihX8LPQ9QZ/6bBVetNWZqD7bPSUeTSW2Q
g3KZmg4m9FuS8J8oEk6sO20dMKvEAEJt6+he6MG06gis45nPhXuXUSCM82BMaBEdbhDqv16opRjl
ao1703KTsayqcJxc928SCkdSfHNjFG0xSP4vHFDjiuVMTQTx+eHEkztEea2ntJP5OZ5QTATqZDsC
YOmbN1kyQGxT0pWIhY4jEj9dfyCvgdbww8MNyijV0kXokjBUTbE2jCI2yTf9oPJ7qjIsbO9pwh92
A0BpXeFNQrHCaxt96rxIXRqMUj9dusIGC5y4ugYiXhGnzBuHEoPwQgRDke+tCazH1nU+8pAREPPv
ydrq+k484RdHsDyp3KbKo+bFr2cJd3d/A3CONED9XRBrlRGpgHcM21fKTqAYJ9+3MNWWw0/cLFM/
AR5peIrrVZc9P7M9yTi8V1FFxw2/KW8GaYobz3u4n6pu5aSWG8mPBaDnVhmsBahZw6aSfQ1dmfzl
tfZ0wcskQQ1tAEqPCJjlHm5NTKyRv/iHnFM2ZrFaqVId0c/ILJFVrZNE9g0+Ka/5+551V6Uz04PI
rm0CDg+3hTk1mmg/ZJqp2VzCxc2EtbiRq0V7wYOZWwXm9wLEAVdNdBU+TcZzeRx/qooLU4wJzpDi
8SwsyXkZ+038ONvMrsG4qJoXy7ac9cf041Cg+bifIPrYa0TCPTkwW/CiykJP5UdoxHA/rDGHtd5M
+g0rBgZhAphLbkVUUHYbgUi/DqHQT0VbYb5TV7dK4X6SwbdEuB4qlpkF4cCpd9Q/hNQ07iXL4u1L
ZRmhr8hTAmMqL9n5ubNuD1jLRf+YRJa3eqIfDcJ1q3A8+1mPSVpLdjSWBjV4BAs93xXgIZFgCXVS
dq8lCJOLLLGZDbUzz6JiiMA5cBMkvKLbMscKLpbBN8LujR93pn4yIk9k9ecPV139u1Z0IXYPbK7+
7SFl//M54REZLg1PmVoXjUe7oKZ6iUp+1AFibuKwf70cT+zBhcWJ5xV6JxojE4668HLKVaxTqAYZ
bl3DK+vAMTCxYMzKSVrvPcz8vFt1d5xZ5k4C+NLhIXMekyb+RvPxVyh/tFAn2K0BarKqt5kdhoPC
PF7foe9sERgVJMQlDj/8iwNA2lNTvEvpH+4nom3qO2VikUG2l49QgGxyL9C9u3JLc7ZA5aSuDGr1
KbT3/Q9NJd8v9FjX/dWWT02zRofCYjbP8JKFhf2k4Xix1HPVYl2bJ9R4KX5cU22SV0dAuXH5Ay2F
M+Kef4BpgxjYUibT+GnJp0RkhH0gRI6DahktW7O40V/+R8C/Ev1AQIeDUFBTy1JL+JH9YmlSE7ds
YWi3EPr8kTvGbQ7tLGXKPe1lXBekVGi0MA3iCXI3iUpS+tOlMX2fXSWOD8MrLluXMjNS0y2CdFNd
WG80lPvktJDLjwIk7VC/Kw1OI6zL0T12PHixImMJVko4CU9Kv1n9Zh9WtAtvb/BKNlWC9eXxShts
xrwDepqwaEpDJGNcaR2cudj1Vj8r2lM3CxLPc+pekOzIKtdys20mVS7PjPV+G8eACBRrQnwWwccp
sPeJCDZSNeyJOTayWKrPkY+YIqQSKg3SyoQ72XNwsW4oefZLZ30HkeuGE9NviHyHiSW6WiJSYIcn
PEPYruglRVvNAIs3RvODCMCs/zyJnpOdz2UT9vPAeiHmXrWP44oFOkykr9wLGTHHanU0dfYjDVrr
2tT+pHgBaFeIbd85VEXXLalvqrfBZDxH5+McAkcxXzAtXtBigLkrfsF3ReSjfhMXfz1XMGX/ihmc
q0zf08kZp3PucG6D+guPoBjUkAvHljIwSCm72kCgiTCRbuzoKJyMDvgLRWNviLJaMGBQ30UtIiTT
KmKqbEeEN1VMzrP3Q3fXc2Tyn6btZ8NGMn91o6fIlD7agkSpd+046n3g5fVIMLQ53Hkx4sr+obdk
q3oIqeJxKuu874Oarde/QVXBnuQVsoWpZ+7I4+gF8KwM+sbYjoH6V19wi3MrsrOomBWMF0lt+LyR
LWpE8UQQ9sowMOYcOT+dWXnUveow6qfhjFcwEhWQKY127+iKm5tn7wA93BeFr6YLzy5ZDiLor4zj
oZj/pZ4FzavhjqDxcnEwMccLYKwFG66VN2mqc3T0jm78/eh1iJc5fyrb0N3DLXpLY/B7ZYI/aMLM
i7iDODVIMggg1gJwUsizoUo68VhojcMo6ZOKwphR6I3qcsh5xqKDHu9GzUE1j8UUxL9ja8K4Wsi8
CgE6yWAmzxIevSaO0fe7GNm7cydve+JROVtVr0rlkKrSUauSDHSCSVQQVQMuE15GbLK43UqUxgaH
4/ed4FP4N7Zocy1Ri3L+w2cy+9y1PKevhqsk1aUC24t3pWmrcariWhJFSWbp5OPUinQvV1yo4FX5
y4CBVgKmnBuhM2ozdq4g+0y+ENI3LYhQwFf4ZVlDb5QraTF2iua3+G7PDvxKtI81EaeBBxGCsmzl
fwOE85O99DLpOHBAa8SjCQQj2tIGz/YFtC/SfV4g757xrFYTJ98ALwZGRSV4kb2HOTY3rdyuajfj
9Vm5vFg1EN7oa4BKTz7sgqteSblU8K5tOnj8ubk9fxkQcnsSmnsJmKa5GPf3rU8PGtk8pK4irCkw
6Cns4K1E8nP+bnaU1FOcIdsHEUvP8nARm66cMRCWPW+mnsq0fPoPeQZjyJWYFu1prsVvH+92DJ3r
oBxs9uShwG/f+dSCBMopxuPpaV4vRY39AlbXQGecKyTVC872R/gTijXRZ2gW2GlXgIUo/R+15iN+
4QcYaJDkMsC0FKQjL96UhBn1Qphld6eIsQWXlQ1WqCVm73oEtmC9v25ys68eM4F0RyVF3P7pJumN
Q4t2DX6ADqitpaHPFF8oOxpuJ0lZ7MUdzgdLcivjxcb+VZQ5CvIM7W7bsicWrfwBTPY0SRbwbgLC
qoG2tGnb1VKATYQ9wPe6Q+Ai7n5WN/Rl3aJkHHDvck49XewlCZXAS0QvirGnvjUyElfhvRWuMdQO
6PlKspQLgW5NC5Y9r9pSDZ19gZ27NSOcwix5KILK/JQ44Of9Ln8YZR5IifEOPdLKP/BFVRrCLsoa
dR8APgWoTXwpp6rC7H9Ez98PfEAsqWwOxyt72rWrZp8p8T4F3qre2XDR3Yf74h0OuI/RTRhqppBK
IbRl5FQTefrDTKJqN5yLAcewM9k+8rSlDhkh2P6MKZTDSTTq/Ft956a8MiaDPDCZ5hzXMKSU8eXG
P31/mAmQ4m09GwXsiIVymMaIwmKahQ7jofHSAFCvHuN/KiEYRPZrOe7rPeGZqrrW69cQ3asmQ67n
HbNZAcyrFMVzOMuIInGhwxzFQkHVQWPkSzVvvSZQS/0veYogekOqTRVQweOOSHD5ojVkDo6rznJr
muIMwRdsLqyq6Tbnk/uqYv42r305isl4QGVAzsmKi7nMQ6xWyjz7s+X66S40asE5BZcnQg8K5q9x
qFzaDmeh0aBIoH6fLV35rdGQf5SWTp9vvsUnHVUKYQPNaMq8fv2hCjtMP2wrorugU90jhJ1EVWgC
rWTo5KerteATfVXvS/l8FDXJd7/mpaK91n4YjYcvsUgRpzY9zdxCD0HglxGMP+Dech99pGnVHa0A
cKaS4XIvxsAnCM+nQqodJEDs3/chRHbQRMWFJtQEo+l/TA/eNGBfu6/5EgkBxrx1o4M+TLByfSHm
sMDKzKZHKBVyC54T5Fpknu318fQOXilkN2xvBvpNGS8bvLqvmVKZ49sxhgmF4k90jhz6WLKJj/+q
VCAJHNCGe2IR5OlAH5LWPpmc7vXQ5y500cI7aKvZNn9WNWkfL2OXq5UuX2EwhNY7EvMZpYp0Ak/Q
ZZ8ZtUKnCgodGIAjU5MDMbi7nky2zoClmE/co7wArQ7ca0mpywY4UEVi6qEhk4yJtm3u8Dsxwr1o
fSrMEFl47IpTbhbY10IkwGqTwmnxpyrpXjHwKviLQfzjCuZvyiYfPz8e0noruoBcwQXm0VvbAezB
rpAWFZz5UIWi49VKVXASuJ4ti5qNJsF9eLry1AoSVFCXhjA7JjP48X3Tv8uf3Vq/mOIofZEjA1xD
xghb7m6i0dH9rDk4mJQ6j+bmhAS0M7zlD1i88V8Sq0CO1L682pvY6QCoadzQTRAHK1KoIFGUt5li
tUyIgYWWsSUJPo5dkrbjINACrQXMrbhpDmAwi869J5gzZ7Ik2G/FHHJzW2+qNVjCQe2iPgEGPwvQ
hoXgqafbizI5BqVTy5YiqIO3tP8AMbd2VSot/aZCJL/QceVB3nS3TeYnnBQdq0XNgfEa4iOrxlCz
hGqr/cjglvq9fNYFMapdFwTiMlR8pwrF4ENliM5Jf1qcHhHpNqSrjJhR7VUmKAqXW29W5k1VPRn8
11bBGRL0qLX3s+eO7xHDV4jH0jWarV5R/y2mE4FEnFDhSkFn5KOGmEqJEkrbpaRrWeYGRv/st7Ve
udKZ+gVCLDWL+vGecnuA6qTUs4Hnwh3uLkpdfcvK4vs+CXAvumVIF4Q2OWwMttKfm4AN4kUS8VwA
L4wC6L51haGhXtZn5/soIsF8AUPkRLI8JcHBxbmLhMIs6/ZsLxyxejrlfv65Bh5W0ncA1fJ6KgQV
+4NP7Ph/NcH2qu3nDD1LFeUrAzUlnKRB4XYNsuQErVlUEXsNkAoKsOsTYzyj1IZswg1dvb7WpvBz
d5Ykuihl81kqfUhPOxkpRyiP9DSUarLFlxv0tZIaXxPsbpgzaYcOLQq/IGKGTEY6lXXFbVEwtpQX
fMmqb3yqy0/2QvQZNHLUr139gvxriZaHdQnAfrxFyI2ttgEfCdQlI9QU8ZyBI1lnYYEwzgyfHpHG
BN3Z5cgsiqvW7KOkdBuG6rYNmpukbfv2Rvs1C7J6rsht4kpQPYu6o0CTwtelpS2pj8yTLWlf4+l4
fytF0/fb4XD3Tl/fND9qvsbe+pJqIDvpZ47tHLb44Tf30qZ7JLeyGCyUxkZwzsduCoAJDv7Udbez
Vqh8lv6PD4SgDki6Pup96BCLM6zRv+R+/72SxMy1iRveWYwf1f5TkNVZR2IPAj16y4i1Amgl0UDV
0RenngBtjrHSw8XSwd/vpqWFGBAD0bIwMZg0covGZxwhkfBcN8q7/t8dXAx0pNpoquo5ObJGXCdJ
F/f1nI1u4VnIN52ISciJTkjJbjiMSa3OtcGnaNTESgwX3l8ITHCubhfr9yLc91J9HO6SXCB+6qCI
YxIDT+a1h9I4ZkMVHTmpqlI96WxufX+xqEVcIwujIYM88UnuwvBvOZpOygHDxSTwSR4a5OSQ5CAy
bwsMdNi45qVk9muodJOvxN+7YoKgmRobiV1GgS5uHOdH8IjWyWolFX/GdhqO2rm6jH15nGuKmdJV
SsRsBAkU66ljreGCpeOBb7jMxoH6WPwUjN4+0G5ipTKMKdtH6OT4OT/63sgVNte4XLvv4nC//sLJ
m/suKbrO39AYFk3PUUgPeVnwWj51UoavrLEKxmbw8VFWRqDyq6gUwvYUWKDOCVlRCgB2zzgFcZsn
YhFDPde+CZ6yex5RH/FZ6hZiNJN6cPdONmjpzPIcho9Q+pOuj6QkSsHocvuuAnosymcRsrYqym0M
AalWWz2ScYCpD8MxaRZa+9dgrP5bmv1ZbCvZ0gsQE28DHsEDsD519jGy5kzsrIOwg+Yx7Xz1hMRu
4ZGO5+G2CmlR03ib7kRUASMLPcVF2Htzt261MAzGvxl7mpE3dHLCvRl12S8GhKWWKziV963gBDE/
gBQuUY/biCfBokVB9Ud/8gxLz333c2BoFSkwpR5eAB+pzhKF1ZXHf/fvsMmONz/BNt+J7XYA9LHA
onEpavp3rWuOFgf10nbSJ6DTSEz+n6mPOS+FQbZfJJx7RnewrIY79B6ENeT6baMgJGVJ1Wmac49w
26YZ/F68WN/rWNzZ4I728FbFuwIIC1DMVkMcPyv5osrwN2GtT9zIu2O3gJgzINlvaw7wmBo3v+cj
9t5hRAc8EpKSauLAS7XMUh3O2NU1XXjKMZseHrGg9Xmd2RRm3ID8y3gFimnjuG3qGDr9eEOJu/ja
nsMzQBBBBR8QVBOm3py2xGuKMm+yB7g+/1bSdYO4gPDx0QCNQXmK715Sd2SCUdMaLqLTn5kA0sCS
nINbEZdc6rdMdsAj8u/sMwXOkiUKEJKovb5F8lpW5OtZ3MI//SDMeALFwkxGey6x+Z1lF1I0sNMr
l/mQ+bnPMv+1nZyAgVDXjbJO9gffzFZtEhc7sltqMHnxMayiJq8g9tygQaxh+ffdUSPUc7GtpaFJ
2pm7/jJpmolAJMacsgj4O60HPMhrE9ceLfikEr7udRodCdk7Snhl/mjjpEN+910+bimdgKX7FxYS
8h5BpRT+L4XHBH971+qTsCJOmQMfGv24knCVF0xKNAI/7IqjpCdant6oYYlfrZoPxfTKw2HDh5x1
SOMBwVVWvqLis91hpZYwEkuPEz6Pia4id1z9+ISdBT4f1TY8g66zNfeaA2XLrhSOO0s5DPTHyl+m
nCIMFyJlDVxMiGFip+fEa+WxMEFlAjf+V/EYsNlEsO+IYHDUzXX7SjfKf9MXux7zBSfWuVFvppPA
K/BLLZ58sUj4/cjlj82rZJPZ4qxzcOQKby1i6T7fJMqhZXWTffo+FWpFQo2YBEple/4dZabPkN7D
iYH1sWA4yO8yRwTNm7flwGW9YPLMPdk5t++hq3EIKd4kQgyKbORzbHqjwn4E5o4Z0kUTyXB0s8FU
JwFTAFn31u6jY9Eh+s1mIUlWaBpvSebkTHhZ9x1xoUUrkNzXm8/bxiqn4I8EuPtCkY+EwbqDnu4V
FA/CLv/SVvpFa6+rSMu8jM9pFeQXw2jUNhbbMNYoIu1ohUAmkj3lBLUeyYr2BzIaE83pOIJayssI
S+TF+G88LvyKIBs9AyJohQiIux0twW33gMLq/5pbyVtBRoQw1WxOQDRva1gfpU/VN7j8XEpXwAPT
BKMbxItF+7Vpft8FlsioanZ9VRl0ZYJBQhL4u6xAFmkCSr+RE4RvOgpDLAaj85C0bOkQiQRydxh2
XrUOaG9GeS7FhdufafnDT9hJxcbFrgt6WIwHXFcfsgPOO6TpIR4eF9dNJJLDS/d2UEgAjwwk9cSQ
yAYwRQ7zZiAsz3hZcvBF0s8oWpfBDkhCMYAsjFqI9W2/3rAKSJE6AYbI5ik9fy7VVpC5IDpNMttp
bw1m+9Iyr+ijmf+aJXx4tHvE7LPYzlPe+VAJD4q1HJYX/kQag1vqwt+wrG3L5kbo6ABebKL2pMM+
ceRBSn+58Gw/DVp6fCvTeL/9bj+jDvxI1wWt6zqaZHl3/sAvwIfWOEXrnCV3kdynRcIdFEbd36K0
OhtrZRd5iw47MsFAQO6HYoNhSehRJA6Zk42CIGWv1gxw4xfHgBi81XchmImV0CprzLfu49JNaofC
SRlzLrHRz8s5apdops8HL1FyYd19/a1l/p2fFdOrxk6gbjqyQz6TSu+z7TE4C3AC3xdVgWjJuQAT
ZZls/ePqLt2hZFrx3Z+DEkBis6PH53gWBiz3qX/P6crKPADI4qiRsBuPX7D7wXdPebRpjlIxj27r
I2XYXJVXPaZLo5307C1Q1nbs2k/7pXZwC/TLn3zoxm658nwoL+gKYhBYYfE0APQwfo0XVdWheooV
5gqT5KKZzvEyOdNFpBGh1RWBJIQs24K8pyA+CmnjD7fkTwpA0YCVBbrmBOYMK4QoLej6bXp102ap
AMtVj1soWPlcMNX2U4+iIFw0LsANgwrDLO/5+hTRwAW1kOwG+qLgFLJsYpu5yFh9LUx40lt6I/+t
TfoTEigckdslqXVSBIZA2aA4JaltnnsOcEoux4t+L9lcvGESWLiRkwGWkYqLE8s/l3iWTho72lHN
Gxnq7EvxhyvRC74I55UAjexmMhnj8p3KY1DYH73vfl39v7vTQBJSDLZC2+1Xo/TYeBFtwEkOYmZr
U906os6Z0KHCfLFpkEara92CBiKetl/g2qM18MAqVpc7PySXsQJu3rkkpGVfuH/u/oMG8OOFtt9s
jpKRzXDEvT3gBLjDbkLcyhDl9Zfz1wuCvX0e4jjITnvLTtzg3TOHJ10cUc4J0fwIJlm36wov2U0W
j/zK8Ln1R09Mmq1/xOoUy37EER5XR6t0CDecbJbUV0fXILcpB5dheLr5ZdtUcncSrtRTqUH4N0rs
I6vHBmDIePlHL9sZqdzeARo34Jced7QlsGqFx58hnHfX+GSXUX0f0t0PAHgW/f2ycTOz/fKD8nhq
LLBdcTOxv1fo0nnbRKQVl4NuBhmNuGAJzOB5jDysrQGFZlxM+dc5JIIdlvv9VsWjMz4VC4W0nL0T
yxf6z05pSC7vLH/AlOcB5kDjjQpW+ZrE6hkq1GhaMzN1lqAig9VZ/E3iCK5NrJId5AtvpUpuDyri
WCfOtLaROJwPoWZyxBprp6TewUiL0tm3SNB2FDPJHRL36fupKvVZlTijZ51Pz/MAqtFyJMBgqJOT
BXj+4W62ICyW+Fi7OLUtSPjUgqZ9ibpeG4kQObIBQfhp9sYpIOdZpybhGCwV0zrebRrXNIM3nd2s
lgmUtZRimRHP6yxPjHsD104IJk3aHpJuLXf6u856u0wY4KT0D152KhKdgmhg6CVX0jONdIL9iGuI
Iu+s1aVlCTCsV5TvGdT46XP8i23Y8VULA4DDjRVhxUJKfnP6O+bDyAMnzmzVi8XRfNCPNAxGSkvA
m6LPsBzESCWUsKnsa+eMkrh/IGzcd9O8brP7Ayb4VecfG0QUHJMFgiz5Q9/AhDhm5xgLrawiilWh
acWFVxzGYqoBIxwSJzqqqyAocczEI2vsV/txxZlZ1wniA0LtFAgWNT/k/0BwLINU6sswuwFpuFYD
uFeMlPySE1dIKBWZ71K0EyBSjDElrz4y7E+DGfDOp6tpgCsLb8OyUHduNffBEmlNxsrSxX9aMBmF
oYpHs9itBjlcjU1K5IROmx+Gj6jGSpkqqcAOTTlSVmvZTuXL3683E22SoDRJ1Wo5VmV8ez3Ss1GF
svYq2aMYusTzzB4cdxBQlnBz+vA0AXHdpJZkWdkMHv/ghx7jFHcPAMIYREEJnF/e0K+hwtisIW9a
QjDZT4HAfzYJXv5tOBJq6eLGRHTBmPbC6WWIgyqLoPisZh6/oV+2bbxr5JnyNru6YKdzc/adVGHT
PVJRBuMSlGb9ZSYAvS2XcunFmZ7ySv2PloWlP/yCAa2YGj3wbjbFSGlUUjZ1jixvgKnuJWh3npVj
QzFjcGOBg7mfBqjH3voC1RayQGyHOhis/xfhiSsNHWEUF0vHP7zdbGR4+6zokDOq2t69KYB9MqqY
9BOXkSIHdLc6XZ6AxM+C3z0IUlOOCu/G3OnL9KVm6oZzyb0DCuVtBzLgjA8xE77HImPjFk9QMhJx
c46MCxXj4YU5BSvsvdJJN2Rjv9iQMeRxBrKceZewUZGPvmMk21JDbnL+Nsv0L1CASspJs6mOrRyL
PUTdEI8IJFTOYLlgqKkwJmDtLAYYX8zVoxq325eGyMAO1DHoaAtIqxdstAhv9bOBARVi+1SP3c7F
1sfjx9q1xqnX5AyU2b18WHeNUmxf+Mr1sfr21ThbzK+/AKyFjtNn79SPbtG72U+5xWx2049jhmPc
CgWiuyT8OkBRBH14a6QY5Wk68CP0r0E42u5XACIAU47wBY9eD3P6fQsQJ3kQotwEPCAkoQvk/ZaA
1vlhsYPIy/7QiGRERDvJ84NxT/wTQIpdbI9xycvuH7GumVxbFG6AmyRnxlEOSPnHyXFBI14MiDj4
So3Y5q/cBpwL6//QNsmAH09T4QTvdRJVjt7pIjStEX/YPkDpalrzLavoXMlsaO0AFKeuqCw00gVh
R2NJvL9UST4ZBU6K29HMWkAIUcGALGTgFg4Cb/Yqglq7lZHfgmQDWJbHzMJ6VPB3utoqNYJacDEu
KMnh5T5ToAl2FP8UjohEOstKG3ikv5wkYKDIY75JHNVWL49BFwTBCKWpxdMGWSJl+ODpj19sSGSi
IKc6KF1IM8jd6wQa8gtLQ2yIt/tXLbhnxqV4+kmTP+6JiHHtPyI7N+pFhlE+lzbT0O49CgGFqyip
EDMrwtmxqb6wQRdf4d4xVfdYeZ25QPYjKe5NrOBhYRkFyDOObU+iezkZauxZI+cjfXJpapAM5CDj
1P0MxlfeW7Kvjzu/DFRGcGuMMx4utoimsNrvJsp4/Ta4wbCmwZnIKtgBS/id+Qg0tZaA66IsKa7Z
JWq9NsITqTtpN0N2+UhYMlMu3ateUo8u+BZH0ErTwBxaLezWC5N0h53bvDlJkfSs8771QRseAN40
QJP34+RWI60iWBtfklZWQ2x+Qf3ULytZ36P6tROSleZCzw9pn4twTd9THo8Y5+EKqFfBkpgypYR1
CQL5oM22emvS2lq4wlFOXxf9xxojTJ+zYE2nvLcubOYDYL+1rvF0Un8jbANw9gHaOaL0CFDtfgCf
C+ZG+kS62xqKjA6X25r5U+l1urE2EFDuX/migt9k6Cyug+WLt//P1Mx/OgjwopHSmvC7Pbl8pGFl
HM6MLZ7d/QSQQdAfrXhBkH97MisOn/ur7NWj6Pyps/++73tNS7nX4tiUe2+F/fTA6kf0bWFpoyph
L2Q1F+CX2LetVh2bZSszsWTZWT4GGAIMZNTI4MwUa7YfF/5H445auOUecLVt+1dWmR6gYZ9XO9+0
Ej1VJ53CUxfUhIa+XT5WfnXPZI+eZDHvc+CYEmRh0VR+bSJKwtZ8OSwZnOW2A5nqDh6JRN//CukS
9+0TVM+T0TJnvsiKYzEnk025qbQ6mRTIpTesp2a2RuMce/KYbFRI1aUVhEXNX6jkRWwdwzC2FEgk
nhQX6lVJ5fXtx3dldy6yFbA8YpY8FU4kMKOgbKnnKPVZ1JXiTuZPoRuiCEq/jvzNd3TPvXUnAVh+
785StleMtIZDKQreVWae9MiTJ/i0pExFQfnzoDtClYAz/AW+LAHA5nsGnZ5EQDQivLkVKijZ8asS
Wal05Ogt4yA6EoSnXbInmPVvKZG/jAaa5go/pLVzvdilR0AQKyGjN7xe33VRYiKDJZo46hQe21rS
oitqF/IlI1RcICPVYlw1/4fJOWXklr1605OZJWaP5deZBKaVqwUjEuIP2/9JQA4+k8T2oXmaN+oa
pRxtjSfZUVl5V9uHg6qFtZ4OqAgHw+YNTFYwl9B1BHZI55qtAy3FF36XjOqMmrQdJZCtRWk8+c1K
DDyBGZHT/9bfUmuIDDPLcB8NQSKqLvCDBDXevAHLHVpjEMNnN2uBpLLPmKsBlthLFvlvO+u4oUdH
lgp74GveWbTWbuiAM3tZwKt+Hp0A9nTxZ4+/Yu3UVsUqeo1mt2i1XPIBzdsxIuJ43bI7DM0eL3yY
5gHbc+VPmbCX+IX/gJ3bgJNCOa/FMVH2YjSNI5CDah2v39LOlQLq9kENkiUxs0Uf6oUd5Ly9GRZ5
G+ybS27R47phG/zZGkNgWQRMpOyvFXSxvzW5yn00EG8+T2gCsN4gcZB8O3BpUsELsFdv/V8cshDk
gAByFGCf+Y1B3gGgP+iJBmYxFC5QdcKVa2/8NuhiA+dVCKFU7ymAOPWrRHzJimpRfd6jgj+1SBZg
TFQG7IwmCJ1zkT5PTYmUmAKz8JABmz36fsxjS8d5gcWRvqTq4nzBzZL773MoWur3zqx89/Mi+aTX
YVva/2eQvZGzmMJbmxvQZEteuVEEHZ15cfdoHFdTedAIxVW1oQ14EJMCIqIoAii8RoWTc4pigQIc
9RUcVgIhoOz4elFErsCJ+rW2PL3vDTEs6rsKOXU+tD3qs254gQV15SVZ//d53PTQKOrePZmndSCS
4Y99auN7qA8DGb6qaG4Ekxk3AZsTPz3zJH9SjxnOr+YEg09GA9R0tsm+pJ4O/x5ZY/VyU8rKTtYb
TuGpqipzhdC01QYwKyUowDzssj6OZkL2XoVeVDbW1Ls+pWT+hn/Xes6qnNgx9LgyXeeaVUtjBsT/
otQvxKLJCmq31Afq72BaCllRubFsuxfcHaa5P9qchNrrMsvV/b/bEZeM3dE9pHXZsgP+vHPdDObq
bsgFcuFA0veZNi5uj4aMMQX2cHhnp6vfqcvLeJKL8aoVfLFe4bzZtC6fTuL1tSjMMguVcUYU+cX/
YqWyz9L6Uj6dmItcjRWOIZsvIc2qASx6ZTEDA4Ar7vb/bUXd5/8CxpfpnopQ7kqiDWOuOiqOI7yq
qBBg3MivsehA6m/W0Ik7wY0adhNZyeik6rRFlqfZaCnO48vkwzsYzckZOe4ae/hz1nh16n+LqbHP
YToBkqMBv2l5VxfHbuEMFxWmc7US3hYbO8ToQYfq7/ib3lx75xIUIp8HiJRoatxyUWub4pwH5yvt
ChI43vnXxGdyKXEFMJC7Qdz3YOPDq2acyTrnR8euxlhthcB86f7/60LOdzlQjZ5rxwWkSTXHw3fe
rSta/I3C6woLL1cHBMR7oSNM+N8TrxdH+LOBV7xJTzGa/m6XtWgNEqfUjcgW33r0EbuI+UuIichw
ybuYIDcapadIrSKmgPquvx48IalOXr2IIZvSX4EZowz9LNY0DyhC9pvQx5fmbnhAhjrl9cJu1+4p
osuda4KXz5DcW48b8q/kojAPYZtolnUSt+wM7k/QFF6oyZ91B7xaLaRyfvRtkihYAWb6pIz1PS21
q91ZmYGLHdWZJ8moxYoKP0YGNFd68Gb7sFYQMNqPjhoTLXZx+sj8TeACyySU09V7JSVB1TDpFwE8
Ug9NZVk823TFcqo9rJKChr/qH4zRjLMMPr61Dn6pLQCZMan6bAX4xj0lnYAJEt0DQrSEHBMp4EUA
ADu2nBXME4mo3zIDTT/1wbHgatE6ifCCGW4kTMcwr5U84FPbcbw/vIHSyMfkqAfB/rqov6Vigt5x
Zx3Z1CNaS+sK4uU/8l5IR0y0KMtzVzGIVDl/9pk7UdBc+15DxfYA1VFzczJJ74V8O7Kqze6NyOTg
q9UYq6n9mjk03KGGphGHOm4C9/DWJnU+M154UbNcKlpPSGGpyu6jcqC31+tMJinSaabKYQOCRNWN
iVAMy80wazFb1Kka5WYlH9h6tIZuLiCCICiUKLCLfrP0IQqGQeZTNz9zuM+SKBIbl+kCLGoqcwt7
WcLVR35xkPS14CW5bcdkS7wWZmh8zr41UMT2seC9BjkNhd6EuqAcNK+DV5AlJlUV0SX98nE4LYep
QAUnNOFys1qJ7I3R9SWxgw6JgWwAYl6ADwYVsgN67PL2bOIWa6oXWKoAXk+Qb4tsUq2Nq4X+twh9
jhSiISLgZCQ1ZwLw8nHAHaawTsMMFA5TYt3K3WF3kShC630B95B3J6txq00CY5K4sEHX7NEj5b0u
VymsI8XsJIa6TqWsWU38/Zapkt4t1nIxokkWF+BP1bDk4kreBUHzFhEom5bbo0KZ++Z7LMy+egfX
W4bMaTzfTCLxyHgVj5h8vzhZjaoAxqG45eFMYJi8hx84LhWvuIqOaZZoKiedKnnZaG1ZXDGk4DRf
ONjqtqKHaOH/JrLVIkA1OaN78Bc5Q0umkJGRaPkXBGMbPiX1ru2rsN5KwmIc0ewyS5u58wRM/TAm
9VbCvHZyo55R5khxRKnACTKNIqvDpFNs0k+XgrFGOglWFV7X53bFuXgvSHHuc+MLWf1/cLLjDELj
l/tJEJW6CCJAhJYX4Rf8IR4RKKQlWP0HMFtJARrBoiImJApQcu6EQr45hj+l5O2oMuhE30KW3B1Y
ycJVeZU35Vub1C8rQWGwh+staVAawyTFfgNqa26PAEPN4NkAgCg/l6VYCZ/nbGuWNXVzaaUDOo9z
E8XDMI9dNzXx05rBGjaY7/5cGyBOmPeNveuR7Jdaq3/Q11O+c1drK0Org6tZSyN1V8eIxP+KNaeU
k+IvlAnFaNepaAA0WGBQdTq/H6NXuWaNd0e67rheLKgvhwbWzOsA20P8JE04phpwVEtGmD6FoHlG
pJR0KdkilO+OsJY3NbFbk+FXP2qIqw7a8meyowfbRNbJitJwV/hJ9jUglyk22axx+nwhHVAW0KlZ
eKzPOEkwDCutP/u/CfNQcKkOHjiQvQ0PM+brSAnBZllVUFkqRe+ZNVFlxJ1IDsPADIsSCpX9/ZpQ
c6K5Vuho4tmbyy5j5jSUXCw4SbRZCQS7kOa8a1xCjNTfxiGpoMCrtlNgWH1KyWNE5LFFGJsGNpeW
z7isZ4n+3P5EP5KXkYEBDbzYfPeVp8Ftt7tnm4rhSHg2VeEJtwsd52pwvuU7Joy3Zdom60/lbxZ0
YW3dM+J+EryNZVIeX+9h749xj3U7VXty6imFooYt9DOBUEKyeVIOd+Ik2rYrLS0uiFUTjeUSISEz
b/uWvSp+ayDJncDfYKtu6+znd1Wr3HekZnDME+IGzxV79b+d+vCALIpJQD0Zk25OnpIl3UtKotcz
30fIGg5KVZKUmWb2CivN/4UbcVrwBmZCvIx6eZscbvSRnm1AzFLwV5iQ4hR0Z447hZevwTTZvpX5
yrHKtayGk1diXqUL6fiR+k3WL/QKVUGicbUAK0HwSS8j4VxH09yImqOkhcmzRWTm492BYBBvjQoQ
5+Y2S7Oh8/hRa3WbIg0G7TSjb7+DP/yUcmZ60aGhZzJr4fiLnu2gx9KgsYoOH8NZ/FSAQYlDkUkp
bnGIyh1nPmTWglCgHR2KXG1Yh6ytoKSbgT/JuOxfJFn5zpn+MElTr+TvsuneeL+g7S2XNXp73oXl
gYMr27brziELlJuLzV/kSw7oL34r6TH0nKV4z5j+PAi1CfItpru7ZF7yOXk+HqyvhwXL5sx83ZBK
INwMZYosCWYEPf+FTbM0NM34Lm2J+/BkUxnc+KbosamaZQlRrTKBGGp30Pnq2h2Doy38ipgj8qc0
gMu+ZB9GK4gdNeMvU/FAliFl4Ma1sZBE8xPe0GlzdWA9WUxREC8/1liRBvsh2jG2lcXmMDvG6d0c
XGS4W5TYvZ6FSj+7PVDIJpVNN5XbKGTgxKI2/N1cOP918CnPpo5bQXgrtjd7F+9VeMIBpI0Wri/0
SLKo1TOMpvIIRAH40uUV1pFMdAnURjPCzp7ncZPRtIaw+hm6Bdnhik/kxQleDv0y3Lg4aG6AlarG
9VZd35+2iM+bES0DyIpeOnBfXRM4wrzo7i/65zrZ+TpD7XHl5O5WG0QhE6cEmSHcZYpR7eh6K+Ph
4R1vq1XT9yzE8s0Xp3sTKDZLMtGgUIyTbyutlav8+1zN0tb5LF8J2qix4VC3gcLTyWhHv1wEKjde
LcbJqM1+as4nHJ/6ym7EkMpLt0DzxpHY9huixV9sy8HC+0q/AF5cqNhfSvlaHWk/DlRvKqaqU6YT
wOiA/uJPPWnK0xCKf7FIQ1qmKzpywAlzCr9/zlI4bA1gCk0ZiQs1Gbrl5ZoNhKFqDpTKDg3c/NGr
ATpQxYikQ46U70MBcewlAzfReo4pb255lNvuWswM1Lt4B5Qoja3Muv7FhYg/KpDoXnbScdVDlrWt
+pke9kYjIgyZ82UkULI1WdO5wUaKbS0pyZF/qn6fXYuHzcQT6IlbPN7Tyew3D5obMEUEnxl5rZqA
MrDW/20dgolMOZnEPRYEwfE4cKkWIkIgc8doxzw34Rw5zEtblpxLf/yQcJEVCKQoj1VdpHiFVt6G
i6mdMLeexBmXBVML750lUmfPMj13w0zcnaWiS5G3Xco0IF3zPhc3hEtd5exk2mZ/gHTJ1URHHmNL
qfQh7Ypq4YJ6KbWWTX/M+p3CSefRC4n/c7dl4EMA1gzkHu2OwxZyIS0mzResG1s8PUrsHIoPDrZE
61NeCajJOFndXHFHAnvk7jKS/BJgTXB/vr8GCCEOUBSf+ASDQmTd63W3hUcAc7ft4TTwVcB+0CVj
pVgxlWk2glNJ410c8aXZyAiZE/enV6zqIy64XRX7gFry47cqNYuISEJNXtLLZMy01jRgl2zwBqKk
6xisviqob+N0o1KAtfooc3BYm8xfhI/qeZb09mfZYjq+v9LAh/fwlnGDXOF6JegWG7VSbw7ZHzvg
5wNzr8kDNsx9qa+Rj9PinzG2n/7G0q8DsRDZbYExQC5Unrf5yf7gjcv2+Pqra1UcfAwyCEFTmxkV
jiL9QyK5/OxM2QQAsAOwUihLlI4LMNtQI86Y5GQZ160SfJqcLzvPfAeinvVhhnhyc/sBP2UqTAz9
TEuNXnv6Xl9y9OYG/932x7CctiPlTgCegW6WGO1gcuSOeyRQkoQ8C6cmZYpiNpO55fh1R7dh7hER
GCKVZohC8dYUEM9BEHq4uJ/VNf7KNRMKeeVXAi38usNG6O94voNkBRnZsDSoG/zw67cooRY9zpAd
YbeuBxnYHBxQ0wtWcIjoIwiNK8z85fNWCzZN5fRZuDuNVTjBRAtvqBsGCGZBYXoveW1LgOcTxN6o
CcUbJqNqdthLt7JsF2ZxsNKhBPRDWJYWW/9MpVJ5OSNo0RH/n4SMk9ooea0S65X7LIV7WeiZEZ4D
XXvQA3bnPFLGBzY56akLnHR/ix26CWL/WEnXKUI6XX0Ctmrar/P38iHM7NhPaxJdIk+Q37utgDbj
tVlCq3xKRUeAWyZEm6KlaWG06H7yCnfgGpGO20c+PkSaeXrwvT0zXCCgBRQl5DFYoKBp+/ub6OMk
9s99vMMUge2Y0RDss73Dh21K/WIXvCrGfKR6oFU8HZXPF+ubqlL7ApDcxFkoexwwzwdcmw24yVWm
trxsAv2xS2c4b5IsmJUc+ysSgeVssM7NmkYM4PsHJct4v0f+QQbpB2MHj6qM2TDh5tm9+6poaEEx
h2MZgDlxbRiVUpdlLPUOZYZxh0W5iWyrWvNeVX9K8osZL+kyi8ZaUGZeN4091kfiivnV2JeSWSGB
YU2zFs5DvJi6+NeesZF5Xv/1+dbDQzc0syU7FNXSq3kN80HK79wBBo1KiPxZcZDEqFRxOiDUSw/b
pmr8ZjiggJZR37OZAxPLUpk+glzpNM52E2eu8T+P3R4THmtNKh24AIjxDgjtRrmBHCXWNyRxzKku
GGh+YSDZvgJ5Pi2w8lLd07HBW3Ik2Za5LfAeb2+kwdfz/ilHxqwQJNAFewuDj9pLD3kpHa0M84VN
lgQm+bUDPkR8Bzl1uEnT8pB39WlXz6sjINnGiPZOq+DEQzxawPfysGq2OLzWAKYbo9DDAREbjV43
ThIlzQtrmcYUd7N5lrcJdVkSjhDb9SFflrhrGnSCq8pdfYZWTQIl8B8mTZX1RoOTiwENk2C19foC
HDWn2P7N70qChNXXmU4AF/fFppxVNfNjlyH13G42P1Nu5mifl+/ecev4HOF0aV+5xo7MYHOW98Qn
j02d2I5LwqR/14VAxzEaFh/qxP+lreel9NbgMhMkqUpPndos0X5ZF/bm5xL0RuW+E/29qCisBiYI
2Sd8YhPnbdfGXUoI5lW+J+G/qspm1490Mf+qNz32tbMCxkTbLK5TDslz3L6IBbyTryIQSE9wh/gJ
14HPGctiK18AVqzsmGqv07uy6WmJo+p7fzNJZzdUceh06/TF6ngGv2QGR9t0MB281A4039aomA4r
Gy7a65XF8jgq0xHSB0oViLSzhAnqYerU8X+yqKAODFvypvtfOYV2FyB36H/JzoM4kY0nZETYtqKw
dG0XibJxN+5gUXePzfQsqKmt7FtmhkW2pSoKZcGCsaynqSlSp2LHzZeL///6pAmOWSUjlKhxf0Lj
VGORXNEiNPWZwLCOGSkYS+dwoap2IL/XCMgTcfKu/9yXK5i6f9jsLIgIpTWfLkUsDL+2veFEWzRk
gZUwCPjiwawSWJbpl3hricBUqn09y+8GdBLCRAZOk1zAL00ZhjAi0bWBnOJP8f4VuSJ6fHYRB/g+
zxkYVu27IlWxjNQRFC6kQB+JmI3UDkUw8TFSR14dDIssPKL9GH6Q5ZJxR/YuJ2S+JQ9b76aqIby6
Wl5D90r7DcWsH3n+xLDVvID7t1Dh5FrSKVw6nY9mNO1FGKVsqdrXPEVIEhf4o8azsyESKzpXQa8D
IyVTidg+A9OlX0eRVj+BukHSPuy8FWEEf1Bb1hwrRn05nnhYlSit7UrEtpzk4rAw+jypcQCjXnHs
9NgS+B2ua78EGrwG2gG6j+5p0e6UuB+zApriPMLK5keQviKlYkzWkfEDf65rmATNt6v3KdiRGcJL
3l7y88cKqtS0N+nEtcr/Op817u4vWk82Uv5iZTXTc11eyOEUe2A4CFudAcOh739YWzHqa5JcPgkA
Qg+IDv1DmTH1oRJUPjmFozKIj4wMrdoj55vSy0++foeXM0vpGF+msfZrh5VspghX9eULj9qljCsb
VVtvFGhoustDJODZ5nO85CxFXriY8WoCvkqqP5DOEpVdLbE6E0UGOZEq0XpYN1/SFIwb/9cmSnMI
qUoUBSmtbuQC2xyPw6W5dFu7iCqoNYDMh9VSpqeFL4Hj5XNIQLg1V2RHNPh9I1aeaK4+/KlDkwpY
VrAoeVkfrGaUamifCjiX11Kl3Ul8WNEluMpeVo+//joa+Fkx/QiEEY9cmtC5GGIDs4cdIWglZ+VD
tsJ6+eKgR11ayptEhQvzrF52BAvsO9KcsVaKiZ4pAlvfWYh1ydt2+dIf4aHku4dpfcTYU9ny7sX9
7d1zLDvO/2eYWwacnSxa/9+Tz3UWKMcQ2F+UrAvtT9TLa0RcXLLU+gQuQNOKU7EbMXYk1ZOSVYBG
VCnoKlUbMRpUiar5Lid4vAk5MeAs1aucRqAAPSrQovcaT/AmnszjjFo32dhHdtqiVFnrjETyV2Z6
ofI3b7n/BuiEpcz2htFosdsGQV/M2CUK1Cp5PRkSwgckAqsI3D0IRQRjEKmLow2mxjeCv/3hDWS7
TvzUYbTillmn7fIVBh4XYMta37BXG9n+BP2fQkPaVg9Pm1XGu8dbxa/faUg8KBaQqV4Y7IHkgLaE
aFIu0bB9YNPHwG9XDVlFqd3JEkPAsckk8QtAtOFG0PXfF8xFKrX/QJs6kr6sl4hfPdNre9GTilpG
ZOKq+79yvq/kUNmiynnDZVj+oLcqSrThyYZ3HyqJSyqlmZSS9NvX58sInQdEZBxaqA/TFkUN4kjo
q/LXIhSiuRryriJbpIb0Vadlkh7Bb1o919MyiLcZ0897ENZA0i4SxfLSz3+/GaymBnY7oZQcMe8W
c+tFATuV8jQsEODBgw7UAkfMh44206ROtcWGggJdzIl56uCtLn0+vqpuaOAyb1K1B3M3A8njjWxi
Pmtnxol9O0khsav/hyvtS4j62vf6CQkazQbUHO3ki1Ceqd8EAqD38BhE4SnwXCRKh/sdnErgjE/v
XHMhPrVCIDjWe7avnVSm9v/sUxXyzlmfyDpqqZap8AWdyvcGMECge4Re7C30RJDT5oSIhL5uT62z
w5dlgTWm7ams0Iu5H7HTnwDUt8VB79voitYELv8YaTWlxN+a4x0YSrYU+jfKt3txvVLVxoMHdb4m
wblq2H/v4D3Fxr6FrdC90NblRMTnYgTk1OSeXMuDfQFzPR2t+W2+bSbCvZyNkcr0LcbydhtEd/zx
Cpwc91q24YT27odqsSxCj+xNMYM4aqeOC1ZzhlT9itFnx5dLt5Mwnaz+jwXl0MC9urqYrjHHo4hi
WiTcaVYgru30htkGpermR4edegcs1XmBqGf1SvMikwu5bJgoA4GcJWHRD362VRceiN49Mhu66l9Y
deV4zc3mUkgc9RGiSUCjRLUCJw8oXs3OZlh0qCdQetiZP6Y5vEWWVHqvPG1w42myA0DKFfmJ29aX
cNquXKHVcvDVi8B/jK4hrQnOaIFem3lux20GZbSNIQ0ODMgy57DBfXsgct0To/qA7o76nUZbw05E
GH2ghcJjicocqNaCHVnjN7kMOGjfppOnM56ro657EicKGchivkuJJ4TwQaQFDTGeWtGvmqNPEjtr
qrGzpxEt9F+PkSwmIH33uxHnItt+HRmcIUODn2pM6hdwVfOetOfNLpz1aB0RwGpqttbKfrxIiCk/
3TGooDrzyDGnnHDjyAxCkSzKBHc3o7DSZTkhwJdrMe2epSeFRmfGVIcVoTQFQIi4goy7L7K9hB/E
b6IGMCGOQw4UkXpUFeD3Trl5xnx86YS6hwYZXIvMAzcVjQ1e5AdIZFJ1IIbGRgwjt4OqlZkLteQZ
c0MsZGUJGmPXWVHgdT9vUkXG4VU0cbCCh3pSYEPThnuPqvvwwvakm3YyGIRQqQFfkQeM0zJGeaIW
N4fWaTN5x0j7wEbWruqWjl6eoyiPyr94YkYolINRV7JVEFcvC7/NtzMsSFpUuUlo1PoQIe7MoZvr
bxKJozRH/AgbrM0/LXnSUc+jEu8grF520i3PJ6/JLS3D8mBQ+FHoorK6ySeBGTWnVpQwN0ZQ8tEC
qVbrDapTJ6nsdED2FuhfEG70R+A78hANdT6rO/Yz+eovRHig4EDTFLEIH1CFMrANQg7P9R/5O9Fs
c1UJhMXNav/Rcl9/ELSh7/apx6+a2SbKHIQ1hEqe6TviAMduS4T53JaUT6dFXU0lBt8VT7mrkpQ2
h2sfzdoJ1LhBpUp+g+S3oNb5ydcTBo+S/bPZLnHVgu2T4TsPZIl3caUokBeKBP9GcvCkyHfM6bPR
e5Lk+I2RwYc/wkgj1EOtM7Z/cRx5TPbjsh5HmPCMazuAljzukI3UbAkumG+TIoKV6RlbPc4GTzgy
NlpRbauo5Lx8d8F3LPMZSq51dc5GJgixgVtRrKWZUrYv5Ul5c9/98tUEBvmoQ8PTI95yircDVCyV
ae+A07B4tZUZJ6uUmQEPidPx/bLgjEe5WU+Iey6My1csBUlS4nhFSci0IJI45MYPqxhIkRqQCTxh
j65Ym0wkZqgemznd9VcRfEfExv59/ruAB5l6HkM9eb/9PVNqrKGzFMAPKnAwhJedlbqT7K9q4rPp
srCgKbTxxFEnNehvqQzXkPWb6vpBCDcxc5FxWiy4LmLv1Kszyvo2zRT1h1PdR8fhpzCCedQreZKo
7L8UAjJVn3+XcbsohkkJlSrLpacFQ7q995Q5qX1cCOw4Sl7XbEixO6KZ7fUjhhWYbKvKmU7dKPr2
Hp4AoV2i5pQdpDfq2gNi8/iA8WcgUB+NnWrSOyX4qzDLecA74zVCO1IeEPV16VTeqQpVCjBDXbYy
HTeVT32wMjphjRWb1/gKFJ7Vv+GSb4HlFrsAJoOSCq/Fa7xrOumb3q0zk4/7tuhDdD191CGKY2E5
U75X343ppehnyD8EKoWt5MKHNAsV03kfbSnVWYeNDxhsoUJ8MCe2kGVNS3HqmdfKNU0Up2AcZem0
qFVc58ieaWG+U1XVtQspUp0McY8vB2OMOMrvb89Ag+XL0HTMHptRM+7xGI6lxGo0DDkSiz0+utjq
v3JtbEr8agkOewcrssOqStOiCgkbqbN8ltMpLnfJH9TQACJ37amS8PlkUEGQ1QO2VkxsB3PuEAgL
V2UGR/sH28qR+e2CCBkaXTrdzZ2YKKKb9LsZ1o4t2B4fAqkTleIzj71jDUvtx82JdJZjh6hk92Ho
yfXE4XvwWkUzCVZ9bnS0rlYW0yQD6ZYxApRaVm74of+Vtt12AZthWYzO35+UF4m4Kh17Ev2InvWX
pxl7FsDe5ASbY6roedJGl7TBVRk6CCA/Ra518aQWSb5/wVgNTaZevIZBzWGT/W1dzMiYsF23t591
7zXwIOn8cssLa38FoXfD08qchK/gNQpH7DUXuaWQzIOrnam1q8opObCDweuSaJuEdy2FDISa1+eB
ba2VDFI3hsDVxrwXEntH3GM/4yRvvJziLuSWMccn4LyT30T5Fvqn7HkIv9zdMN9J88xWml/Bozc1
kJhAx4oTqkYCCqADNLEtt75nJ4JabDD7P6lCv62MCX8h/1Cj5RVQudLN0VvziyGHkT06c8BP+/Ln
DsjzjMHGczibIhKEDNn79Qjf6iuy3OwRxt+PNh0y98LR8Tmza4Bc45OQ7LZOtp5zNQAwDswYwNkv
ZEq24AOi13cIZGJ7AnO/LlCJ/4JUTLXKXGQuQDr0/AMSJOFSX3JhkUCzNIuVSZzPYpX3KAm3RRye
EZhaql1b/oFoMCD2JkrhyFzmM5mOvYA3uA2Rq4Wh+hvh2Y/mdCojiaCS3aG85XmHCILxDOexZrpF
eZbTUzgf4BlI2RTwHNVMQ7AkhrZh9ukadWrTaBJRAS4mu9yEuNvOqGaDkzMxPdOFUaTxLx6oS87y
7mip1ky5cidMMdrYkpswOX3FeDlrbf/nDPss1MkpiI5DGsTnTp92/JSm68t1efv3zEY4/6FVPQG4
FgAA/fMIga6eKTj5EhbwBYTchyh+LniBuAmdy9LWL6xBtFRnt+ZcUfdDkvmMj2zpVKG84giIPNmZ
eQRypPKHXsxADiaVyBOVezp8ruB58ncSGh1WJerOfsJO06rr6mEK5BZicRWIRbnpu/E4K9/KK8wE
JKEmd1nqSK4yRghL0jnwrZVaGYDXENrhoolA/ZxkqyvEiFafQbSIhPMA70KE+N+XELa0Q+0BfjJa
2p28xEIEsi+obXOO+C4W6QsX5c3Ghutp+gWTgw5kv833Xf5y6+hQ/XhlEPKsO/5vFEV+fywfeevu
T+6yZSf0Ipi0Cwvyq1g+JXhdRwPICWb8pC6RuzOf1JKKnWpZPZElQb2BEnI7DH8kHMsQH17VwVEo
Qy3g0H/x5bljaKHJOK8vAkZzXt2nKRCr4kPmb9/oxipH+TaE22IgYEWIjDaxR8oCX74qaYlKMFjn
cmu0pPCUh7LQsMRLTbd0DeDAnHFvmIGUH7ibIYd1FnTnC4z3lrNrV5ZEQAZeTfxukOrg/fD4LVs7
p23cTv3SFuaYj3QV8+ijOP6vovR2aY32S3dTwXD2WDIktnwgBiKGfEnNV844awuQdn8F7GqX9Inp
h1YTc5yW3Y2Fj2rykcaLI3sVieJIIqS41rfX0U2ACxPGP67pIKygRzCi/QJ+EGx0ajbvUa7GYsH4
lkH4jmOqAQkjVp+0T/ifz+2Ib/ekDF78ZyDnAQRYOf1Ic2A7yKntabdohrXiwML/hahqShK5esaJ
a6Gqu3jBGM9eJtjvtk3+cVOq/9oHabL8wpvUCsqVY6tdAyqjFeLnLCUs5TWNt+GiNqgnZ8NNizM8
76omUzwwtt3cdOYmSTXZUc8yfQV9vdAftu2bFPwSDCruUCjMuDox+n6NrukOg16ZXzZ23n8BJ23+
atVPJ1lA2iTTiZJhhu5eREgCNydxtMJSIbJIUWbmkqMQQiwDKXLzXuwjtc09tvMpLFY3SsN9XDb/
rXXeZkJ5GiX3koioBKFp1Vt1MPTqU8j1jVO08xhTdLeGcPtdXiv9TclES0qi00+kxwHxELpckPSS
lnlcdQusmcw1gLS5lMPAGt2AZzijQ5fJYF67sODmk6XDYbIW0Fii+4w4uT76Xyb9bnevb7x64sJ3
v91QmzuTMm1FxiBXg4cb69FLd5V/BoDlZYmbWXWqV3A3x1AlgPfHPv/mIFP0cL9+Z1A/hI3qbFWj
zyyct5JZpvnQFPbiUzDP0W7wWARPVHiUpoI9aiJAmyF698KAXsF7KJ4nLTPwVdZpNWWg0dsgbyOm
6X7NRQ6GsPKUXiybEiuauPZEPTZ0Vx4AFKNLOre5dL4WXA5y3vyNKR8rl8NRELDUuSUHPA/toH2Q
ZQ5tlUVtToe/UdPHabTl6IzFmilio8f7Oyl/1hB5b9y4LyM7xzTnvjdQCjZHZBSgQniZfEjWdLPl
t25SB6h/r4GiC+QysA4CW43AvGNaEHP2e7vVVGkSkkqDd/VSzpfK10ZobZhyCAK632UEM5nn8MtB
re138zauzaFvAC7umW8RJa4XlZSVfQM1f++uzrjC3W8l78/gA98QZJ522+yUGFqAjU6aRRsUuif6
O4/qOR2Z3PIyM/S49E1naU7oevHXTrbmh0HwdwLWsgj41ZZWbUXCAr7AbexlX7MWuRGXHG/Bll2s
Wy1PH1L7HjI4I8f8ly5b54WZu4iz4+I0cMa4F9Yxd+0x+xPhJiCRTtKGcE3+9J2MKCAcp86zQdtu
/1h/8Rlpk+X7tXzgOl9EvG8o7MO9PzSX8WKa2LQ5dwQVn1Z5oCJ2w1T17Z72ioCAAGbjeLfhk5hr
B4aQKFMEnZn+qiJBvHvtItbqTqZf9E8zk8lRLGo35F7+uSrOO7BYXSKj2Xm/K3E17B7Wz7uaRJ5N
HPIHsAuJ5a1JF+O6vzLMPhMEQQK0ty/ZWpJZpk08KxUHCxi/peNpgjM/0ePxASmBJnLG6IoEU19w
kLb22eOBsdDBHIf6dk0etX5kvuj/Als1mgjQtpO0bt+TtAZ0G2XDZQYhsSOk1Ct4NnIzECyb/WDe
MTDIB5pDIcjsIXiMlLEBfGsWEFl0CnlJEVSO0GeZU+t0X2RHbhuDFQdpoq+3xVSq64tcj/fyBUHu
kYUlktNX35R9490+t3XHDAGzuAokI/opj5R2ZiEDsqH3Qt3/T23pWt+FUERWpIrr8XRKs5N6z7ZT
4oTCM/V1RfjEUaqmWmV4N6NC4Ucd79xGuUKV6qIcmzpanhAy2Z8l0hQ3n9KKVMbvnZ5AMXtgd4iu
7J49Gik1/xpH5IyK7epSHX2oZCiN23FyCll4xyVJaSmS666b5CLk7++VSNmXVg6QG8DX4Icx6YX5
BW6Nez3JrU47DakNqRm1Pbk9eJDbXFdQeKPeWpX7PKmF/fo6IKO8PhZDw8wc75jPlq59Xt0NIuQ6
thpxhNTmoa1bAzb5V8LF9ASizMKB0aV2QDbeb3m0Fh/IHnQJQRYguzTTYdyGPt2UYdesuWVGeUTb
9+g5JfOShklPdgWzV7t7L2xbI8azKrLyYTWa99UNpxCjZOPFuegzPqJ3274slQhPQXTpTESuw+SF
5su/VtSmQlgU4mPymUzsnBIEmSmOU6DWmRjayS4APhSzt25i0zgi1XTHLm6f2AQdOLOg4c4jd9R+
UcMIyk5BueN8ySTTZnQKqWa+ETPfn8pqBaOddiSeyuUOnL+GXnisbc0fAHOTO3/Bh351dnoTTSCk
Jdzsw8AsQMrU/e6RXKF9zpPKZYqqbA2sJ8aikVEV63YlwW3fluNsNaokXLXu5XbsdOVyx6tJxWJk
sYJHESYBYO7ZDcO/bO1+euQY6rb/PhprHhYMzlxLVQxE0oMfsoKGfZsavPjYc9lzbSVygVN+/0Fp
uxZxyaRkMUfLZclIO4nRWkwyYdbhXcwXGuSeloKogtOaRY/3IloE0tKrQpv/IGDfAqIubWLSQeDQ
xmi7G6bssdKpiLhvUV7xNhoSETYQvqNAuJyPP9/IH62v8b4EtORSZ253gWY8neXONPK8vASaihiV
NNn5wLoqcR7cmaytNMsIPUpPscLifN4/azcs0jTA2W3nVD6yfZ6dvBG11Z8mGIn1dmvLernYTKVq
dDzXm/L0r5hk4wfjY48jX20KhxUBd3N3Kqmmw5ybSJhGBHcZ1rHgmcQXcbKG6iV2XW4jQD0twHsY
8mNZRtgTvTdGkHk3mHpqXIvxIh/V0qBEm/PaJtNDHZ9+R/X78HA2n3TCTBfXiruf6NciWnw60vNw
ZMulDMyENo127WmNbyVhIyF6b09JCryWJQ5txMzaQEqPy3QKv5vUmfLOmW/CT6aVRQMAE2FygJY1
t0Sw+1/OxYlYs5umsfYaE+RlVZ+BRgCvkAgJ14rllA+ZyUYfIX2KTv2dd1hCfrag+s5hsSZQa1E/
GFnKdpNZ6Yxo5uyUuuvglruKzv7Jrrrhda0kCTiOKEAVe8WCwZtZnhEtP4Y804PZUQuHmtHl+lAK
EFgJiQAstsk4Eten3Y+iun3mEDNVTmsfgs4UBX0j9tgxWbLGlYfZ76ZV/kw01IjFynRq3h3TbSqr
bpmQL/i12owFqbZ7Dab7CwzDUhtb55AfRirJU+u1PFG1KDVAlKLaD0tNeERhldiUJkvMHmnAOeqr
4LC5fxjaDFT1ieZ+OF9IQxChKUeeuNfVqATNL+Xp5tKi+sevay1NZPhcqd5BR+yZi0i24UshIyje
43vkAflbwYp7LG22KtqJYD/FVUnpZ3XhAx2tPtduF5WPitlMYtkyMCOsHEyD0BeNwPHgZM27L0LW
SyH52LmO4oprR9Rx6ArpJmd0U5EBTyiSIr0WRN9IbmgjS727Cx/gIe3CjJVgRPXtqIz2GxHrSV/x
wDBt+7fMyF4fqFE047IsCLeiQfg2krk+F2cb7DDuW81mXwJWGo1eZr3sSCz0xu/Loifmicd1Yc0O
VMRR57Ec6zuBWbYL3TC/By8SBDGf2c3BsOWotApmGqUHM+d7AM875WtRrYgCEJbwe91U4WmfrwQn
mQwwygqkI0eP50jB4gjyEWxdT/kpdgxqa/UKbKvppEoYzO7Rd0C8jeNh6F77FwZBRq4DLj7j30QP
ZqoQHadnCoY/Wvj4mJP7RTHAZKKhsze2nMXd33sdfR2iDfk83cTMbnCwP1iK4RvPMBb03RIweZoZ
HpKfrdqaI3L/nZPWARz4ulXdyDGeyQhosbTArPcNDHzBHxRALU5EFMupcj3XgjxJAYlqg/IniLBh
Rhqglukcgq/doEpNu+8JCJMnFMvjmwfL9jQrA5EQqJXI3sehMCXBnB6HM+VAkxhIGkSGNCvsIrId
pXih4iovseHVVdNvcnQ8z568FydjYrhc/x7bstIXNnpxDiQ6cq74wK7quhGJh+zs0bOCZSlj8HW/
NmpigomIDf8+NJFkeFs7tib3QlcPUSFCjgOWbtvXHmst5rQut5GII7EtmF/Df3G780+GVi8cocG0
AAWYL4QvEBGf8aIxvH7Iyy7EYLSAxo7IxCKBK4mh3nnz8xfd+jMTnxCdXL7ltTb6I6nuO9vmBLde
sVD0Gn9tXcX5SvQ9zDXG9FD+pykff6Zar1UhXqdeHqjVH6BG+j1TcKfpGEzxPwOwRa2dgcYPlSYO
UQ4YyIGJecl8BdEfE5t19eIhYAs0Suuxa3VaRMtaGgdZky9fv69W6AxE4Cac4JPkFutkhP2LNz9H
0XmMORQ+LZKjQwbUBRDKOuJwEqUgOF9n/mJVlCEPYQa0NiVEYlKQmn1r+aaAKmaMZoCH+VAKQryo
cy7PlNmdzz5sQVNufiK9IAfL2zrtMuhShzB08zQzldovN1w6ZeGhSStHHzCvwYjBy9Ll3wIaCIcF
4Wk37aBKfZpmZOeCaKMkg0pvfx6oybOa3UCrty5nfGsAH4k3zthD/Baqpbk+uMBdb/cTXkVSAloQ
2FPPaBhEQ6UwiLy3kQItYqfWHk8LX7k+6oz0ipRDHzr4cFb7o8fn5NbEePpHAwbLazf6NgjlDxUn
a8yjwsRshAMJxZYh6m8wq+4PKtQroH2vuQXNqwPfzNlFeeqii6dNxMthTXX9Pm6qXkQ9p9pJf2D0
WurZ133gKivRVzdmolqUXvkGmYlviIsNebFFh/5MwC/Dxbmz6vo8nX8RN+qCj4uW/5yHi7jjq77l
KQa0dMdqdKIEu4Y3Wf4VySmPhn29d4gwNX16pTVC3UQAq6RZ+nUEovL/bRXc9NPyyzlcQNR5K5OD
EZufhMxBjtNiMxjhj66bHQKaxAJ/BMGp5bF2iWL0F0ED6TB9XktAzda27ziERpYLh9i1YRRo9LSt
taz7gcOzKNta5esUrGaGwC0mAL72waEQZK3tt8LSF4DBm3AhRbE3dfFbpBTA1JjdlY0qmVkncppT
4pfMkBLB3RBV1cpFgzetgg9YquNPyA2xhECq+W/vIMChAyFev+6P9S+IJFnftkGwtsuQeauGs0zw
p0NTkAcK/ihqYtBQJFWTNMg43ZdQCj+Cbr9aFqoosvHbXygztps9YFEXGvLAfbhrCEg8ZjBGVc7A
cukO92D6+8JudtjMGgeRaOS1MGK1Pt3Jd29M4wBtLZPD1CgH0aha7wtXJ1vtd8qCq503zPAp4asM
vXkWhjegu5um8vIxciI4sSONHR7txF0HpfizjhY9MUsaNJSB5Y5DcCuWAcdtxE3Vv9wxrX7jGgr4
qndMeSCAqEWGFsaFBZ/m4Y2/BQMuWA75Tn1yd96ng0UcCfn6jIWqESe8pSHWZpOoSM5WLIvZm87u
RO961Sw2Wl+gojz2u7Nh8Er+zvuiQy4Lqn3d8lKkzotKrLL2eUK+2ggS7VRAA1Dcwfky0UI27L7r
v7C5vl/SL3d+rNam5Kp+2zfD7taUGFyegVMtRyj1dXZsRn0YMPYXxQrlZ742jx4eRfkAF59ef5Ue
VnIhz6K9S3LcXJsCmO5OIpIqjcXU3MB/oL4hhDFv3BCiQRV1I7h/wkRETFWLvduI2x6xU5h55KFd
syz6tCpaQixj15pHrQXVjBJqTyquvc/8OvRG7uI4ajZHLDzdMeCo8AMpUAjWjOQVG3WwKm6dU3As
422biUSU+j5nIvKMWEK888944DaRKYkpLgpJYdP73w0GrEGem4Z9yMq84svFo49L+XYTdiRqjr1Q
9X1f5oiFtRLILY4hk3oarHVv2hfBAcAinxMP68VcFQh7hKQaQ/zckjssamLOr2IPiZXa0X8ipsTf
rP9TIOlANUnDz27411wpdLBsSGpZH9SZD6p2pSJbV9iNh4x05vHaJvm1S4O4JuuSBroPZlGdr4Qi
tpVY/DqNMNhvV7dTEBBVcnikQhSqGmxWg+5VEeOWnlY5JUE6dmtbVxYMve//tzV58dFLlwTuSrU/
32tj98XB7GtKNI4YhHKHnJ7d6ntp8xLQqO7JL/Fr3c1ZsUSqWhctZj0AvmAQKvga0z692ggBdPgT
hduVZqNQPm0VwxErw7Ktld03opTWHJWtqYvNwDHBK+BPwYUcAvG+MOMsEMRD+wC/FBDxFvZlkz/9
kacNlAwyeobn7hmRKLUjJ2oz62dkys5dG4/xLnshX/T5riz0RU5AQPRNXaZTSPq1yhyhExIxlCaQ
lnsIIbL+ZG7objrZkBn+bL7YpMEvkvCYPkVmaWptosb+DdY/cu+9NJwwLGacvBPdCFIE/5j7o7kf
S/vb9ejtArTejHxlq1zTmMTBwf1NT4XwmjosygYQiG7dXNl+4IyXqqGa2yBgijsanLZgkN/3SyxX
cS9m5rJiXmEApsOAs+QHUf9PWMaj/h90id1UKd20ASBCvzx9xUksW2gneu10iESAzuzpxnqW+0OT
POq2Sd+c637EKO7id4fwf61i8PC1oEaER0EoPHMP+FqtBZc0Isa1bXUvstgUnJrYvEBm37O7m652
OSO1LmVJen1RGxZvyqTE6kK1kwf16F+p+dmXtf7/BWQSchOY5epKrmakINkgZzoxd0sanghQVwTN
NbovhALQShUzqMuRA9atxzJVmAcHoWEupxp/SWzF9qEZORAsWyEuBllJyxmolRq8FMHpqHvaNjmT
jzuV8/cu4NC4EjTtlcRM9a1MidxG3D3Czlm0gYogLswvtwjs0g3GVMRdAq7mU1B/0p1iZO/QBs/n
73pIkYs0yZpdXRDR74z5GaZCvogrsYk8ZgTcRLFHWxoZiXR+/FejE3UTNgj+AJR977SZz2zAXQN1
ngRSkg5haQKtTqutKbwYD3bqoI3AoyZwmxcEtbrhbMIv+6CKLJu6O3Nl568vNl6EamBB6/cqVJJI
/G7yM9HduNh2x4Wy5HXE0eHoOV+wNtiRvo/d+C89Wb1o3MFhebvajzrKZKOFeEIjscqadxpeWDrI
qnqL9mmqbErR+qADYsSZKdrVWwstWl0eABI+ChgqhgK6/IaHykzRIngoSeYtCSI++kKM1WPe6vlY
wkftBaH7DHIapJMRHHRrmpQZXNycusWR/iA0kaVbpTneXvwj97J2fe6ZgxeyoNwVTtJs5dehdP3T
W34jDzLRYV0b8hHdJnjpMpv15ywhnc2naQf0IDLugfff6ZMYUThRZQUOxGaoLiHYPksSSTInNQXE
p73F9laZWOLibrJacYA/Y1NRFo0RSp/55wIimHHPRvcZLYOiipbxCAwYPb8ocRueklWkELp3FE6u
oN4oN9zTI4yhjuv6ZE50/NdcxkOeKZlkRWvVxPSavIf0fRf4+S9R8KAYTIIBDSiU7qjqa0/91cue
6X1PFSKq08tYXubhBvzgxUiALdm5CxFf8uSzIRkth89MDM5GpA36FwOxW2i+cCcD1Cc0qzqV8u3d
JHeZNKaRmpna4OTM4X7euKK6I0gl6CODpYlfjxoaM7B39wahz70PsmaUIWHnxl7wZuiwoIOi64tH
JTOWENZVhUMGVDnRmsYwHFEjJ1ClX65bfz0d6eex+SNK7nL8GL5AODP44GqqJRqGoGocr825CT8I
/ESmrzOOivH4zN+3Lc5+J2eIH6GS0OKSJV2b3+O3n3WH38ub+hW335rwuBMgyJ0OQmcgAKgK52jb
0jh903L7sZTgOplMoaDawEb5CKR3UYJCfNFsJojGnZ1U94e6lPmEAYYkvdeRapVrG2zgA2WbjrYw
tvt2+mOEZkEtetlP/Twn+kBt+qdD0LWYEiMgzi1BCaqX3kH9U3xyY6VjgD5qCV/MXvjSK6YlOS0K
u1kWvvZsNF8c7pW20vCTqmfU7usNqxftQW6SFZltZC3Wirh+m7VQ7RCf0exXOt2xvjS56aeOoj3o
+08cMAlFDYhsPIFhUGUy6DAkt/gZLGoYCGoNooKvN9xKC9HjV/B5mIdAdaHOmR6ZJ6asE77AfId9
8V7A8Vd1E86nxAArKZBkw+3KMFG4M9deet4WZDxicE8W71rM1ASJ9Ms2A2QLvxZAFHY9yLg7N+mJ
iuX0jC1OvqY7+atGovaQo46IZ3WtyGdXVCt1JlQW2hRFDXNkO6wsogwzndMa2QPZG70fS509DYed
h20DIwErPeG8lcEfrJXRY1fyut75ByYnfzefahOpkb2EUlUPmR27ZtJcmBTYsXK3B8inVVbYWfDJ
hN/1432NcRA6Eb5vBS7kMT2Sb3cNR9qsuClB+e5svkXKDtvTdvdk1ZAJCm6W20CycQ6feHf4RBF8
0uN6+p6lQ33wp+QOIuZkf8Tensc2c5vX/hp3CMLykpQ5LIvVmd4MoS7NjQeueI3i3QUGSa0UFKYT
VaAnqrme8gqypmTu80ABRNSy9MXMzryL6uSRE1nm41ozpxGAgffUy6E52eisZcLNxS2C+Di2lVd7
0N/HL4DycIShCF7vtlt0KmB2XNaNgNdH2YXlDvReK1V1eRPiCtHt806POmRkj9YjOFi0T8USkopA
OAdgeuFwhsO/zxpcAmuwRe9Cx5PYHOVwTjE2wtGT91ugu+jy+QSsHXDS4LfjlMtZcaOjsRAyMTaL
Sc/EpzgL6m4CTCw+eFU50fekXI2WLLXT2Exg0Jrym71YmpQirXo/GONn+WS3laHpYeAkAzyQTe+s
dJ/FL3uMFybSJmOyBAu+m+c7sEAM21vtkJBjJt3+Ph3RBmEB/k3WAXVc/S3xe1YnUupDwop/J/6B
Cru2UmetkQxP9RQGN9EZns8DqT3Q1eUktLdhuNnuzwlzj51fc1L/WjQwF11baPa/fs6GTJ0Cqh9D
b0jIqsYpDBmbtonmh7gWuLy89A2NRzxvxQLtBjp+oKrx477rE4r9yXWgKBPY1JOtjkST/8nLgXgw
LeB4hnelUr0tj1IODlqdS3x7jD1IXrehIwi4mcUKp91fQnnxeNr8PxRXM/0+McAURtdJ7EPetWIl
7k6KpAQLP0geUqa6Pg34PQgssM91zd6YD1hTZcfr6zGzp3wJJIqTgdvmpdF8NFCCDjLb9DanCYSF
8lIIzQuJcUSkkbp7FKxwo1VBaJ+AZucqY3dSomQ9ez9DYH959B6T43k6YypXl4gKQcQ4I04SeJ0g
VbIf+s3INU3q/gRC8t1Cexh5jEofbiLGnEaKHVGhXrUWIMvcD3HT5K0VB4FTqqJuThAfUqEhZxRp
xau1elqI9dUt+X4Bpw3+0NVQQexTZz6MEa7zYijMpKH89wrzAqD2YBJYm1ihz+BiUvihHvkk9pl9
vt2yS+PEKy/pXEA6x0HOwVVZ5BfMDgYFeChyFmXxTjdPW3RKy9UymZ+kIpSjdYp75uvRDJ8IHRoW
gmL1JX98Hr0nh4DiVer5UM5wNOupEFTlCc0tV9d9w/JWBo/s2Zx7GeiV+h3M2XvxEDdVu21ADkcx
gf/tMC1IK9jjGiWfZPhqiZGAIUOVzJrdCfTuhYNmxMR7SpF90gBww514CRg0vVk3zcwR+cX7a8h3
1g5vNmtTj7QI3fT4WPD+ZHm7iBmb8CX1vuAX2XgSn+MEOi3noSzApIVgms3MiNCVtB1SOKBSJ/4D
NXhRzEBwUMXbgNqV0n1h3FHOXprdYBnm/5UR6oQawBSB1aT9lCmxf/ioUu5ChXtL/k/gBk/kNLHx
ECoFNoiwh/XExudA8QPRPAvYRG4Fjjd7e7sGmCEwFS2+VDpwMhtIC7bxNBN4eHnXxG7wLt2/e4+D
OzuQLMX/tVJkHOizFaG7qceQuZklH4AN2iVAOPbbXxmwjPfqL0rXFAEER7qUQxRyYfAJENmznXwU
CrWSFIFm40nqjkfz7eWaKU7HrwPO8jqlGxY/kuZVb9EiH6ivqGz4u1jgnWyE2EQMMhPRiq5ulm9u
PBGt1do9zp7xSRZszqm4ntpZ883yj0xwHUUKfD7HZD/EZLSC2/DBM1v6QDDM/xuQ1YZ8mRgSqukL
MR9kzCkBfowFg+15fyPGOaFPPvS2MddsO1KnkT8yV8ObWRtNrGbYxeFB68cvAswDX5hxKidruBa5
c/1bT/esqWdUD7gkTKR5ubOMCyt2/TAmMOrBDZtqt9uS7ydsHbHz26rgIaUnW543PcfuNuR9Sbg6
0GYXVwlQfqwKB4zqwWpqd208gcyMosr4j36S025D9NJiFZsRqNo07GZd40XeIWI9LTyo/y1rMcnF
5Tq1VX0lHeb4nReu4i0wcAOjNg4tnRqihCsc2d7QhU5xzH+Y1ttWlobcyMtWAZAMn1B2gKR+LcQv
OBGtIJvn4ljgtPSz6XyU+hBssAaOIbT9W69C8qnWmdBJNlZWeOSNvoLclTkLXZ+7NresUK1x31sz
0GxaWugdACiV5DUMGVnHw9Jn+jEGf9vs2laKiWO9MlJBir4NINHX5ejdawM6aFazAQddfMXM4Hgb
ksx6sIFp5dWNujhSLx13wu7sukhz7+E51fLj0QgOTY7yFydBPcryikHDFYLHd19LEk+huSIumZEK
eMghrFb01M3qAw8ndBRos6RTZl+y9mR481A5pQd8TbQfatzP/Kl4D37e9twmZ0SnRJJsDTNwPiqq
W8xuTLyTXp/ELbLWHpVYMOKjd3nCajvI2YBO32LNPpWGVPbvJXJ+2TtXK8b/fw+a5dM9NqtCq7mU
VqS5ogia0plK3BTv+BHpgMjgd2gNyQIW6OsBrmSC92vp+2rE+MSJZ5//34mHeiASHJ67wZVsoQWu
Ud2lgjFaGFoq0ICSyEdfSyNHI79SisRmkfng8ozy182N+4i4OlI2HcA0+oEktlU/o4PtH/3z2q5X
NO1bs1wvZE85q9muP7O0baoeHYJNB7z6olvpDAd6wo2L+nkhIT6P7VWrB1A8/RyhB9JTXQXPj07J
t8C1ScTbx6cgxVI+eR1ohS45y5gT24mmy9XwG674Gk5lHyGwLvWiYLdDkcqrLZRauGpGUdyUO7pg
sCjJPG5/BTk2QHvt1JOd9pSaiBSwzBLKsdd5phSZHhptfDDwTjofX3PZlfi3V3+3M4yRX7vxGZN+
gNXujm+MORgzK4HH00tTtPtcILkhr/Fr+VG0wQJ+A4gbzB8nOBcOhlmulyJFadfLNf3gsvIe8c1w
Xpp3s6KNZtJsJ4KsjZs3bAnHpgrFhbsmbDMvSPZ95eYngpBeTTrwM5DWjeZfWbl7WnPW//UhdnKe
j2Dsx5g8Ojnz2hpv1mzWQETIWtIkT8l2FDrNwB091i0JpyPAkK3d/R3xTr/t1lrALhmz8ql4l++0
bNDhLDgMF1Wm14SCWcTRTxxiNJjk8VbzwOOYWrjfuitFMrfKncokOp2wX237pF3r4lbqydkbwePn
YAANXNTZ86Wd+2oDULXEBILRZpjxtf/8Fgh3Jr23wSfFbSRX53zGERnR1B6ohunSDZAQykz9T3YO
qgI08pWZI9rCsh2y6xqnkkfCFWfZGNCn4ZZm8xQ7flR5Q0D/kBuac6J0ACjhXZaxpxqhIP20qfqJ
qA9/AGSy6QeB5h9jjhTY7cV5BovRdIiF8yxnBdWMbVeHFxaCBkcCFRommZBXG5nCjdx5T0zBqnhq
ZIJ9hPD2kh6ZwYc3wRALz4jivWOrkIGMVULgnKpYQPefdAyrSdlbygta2nbGvVekyjaBF8ccn5nf
Hj1jVigPkbjiHzd2mmPKBL/7r65u9Ls1+xEdCyHsPwnUaGTq4m9dpeL5vt9LHb2qSQfRhmLYYAAZ
VyJZC70E2Nv9NHEvnlU6l5/bZwALIp1JZ5CWVk+BzFPw7fjT9isz8niTECaeefXnlqQ1fxBhfFLE
HnDtNxjrbmFSh0uG7mdVTzUrCCaecIKbPF/tpfN9QI9s70Za7YEB7NfdpOcc6GrcrXVBotwCm6OQ
et3eGWgLsJJwXJK5wfDKaDNjotjhQMwaJhPr/XRECN+2KID+o0ojF0XbsT7X65F9oTuUPpNNKE5D
q2PKdW2frjuM4i086tZ47274wzUjqWXzz8xO85LD6YUcAtqYQ0NX2JLPG1ALpG3kSnCY1t7sk6Yj
70Syhd+1K2+jSLtP21mskN+jD5ZYyJrqkwIzrVDdGtu6wGNgoyol7MLlN8CuBytWaom7VqLZZ3qU
HPcv7YGbShKOZQL+a9yX6mf/OTcfNjChPdsnO+rvyP4FCcp2pQJydu+Pnb6gsgdHhh1NNcP2yatt
FGiryUI/0GrFp2jqJGV9lFmjwibAcBUAqOeknqt8lJ6sjaomFFK3HM4KFpdwmEEPr3BoCcLcvULY
noBNYMKkjEim59nkBaRGgMT5HXc/NI7Ael3zZhrWDIbkL5OUJS/bo2Facpp9wigdx4yRHA1KUwMJ
7Ip48/ouNXeyvGqeR3gGdrE1GlyeSx9nAHIeQN0OmlvcfJCEsnglU23OcNrfRJ0sYQ6OS60zWGMP
dcQGEbxHbn4f0XhcHK6k5oNJYCIYv9y2xgS5EK8DvHUAWufV343OajWk9PHDOSgwN9grHPPapkvP
/gW0oSpdBX1qp2gLW78Ey/A34W0goExoD7IwPGteq1RWoeHjkFLRxzDNZqdsW8pdFocmI3OVx+Lt
fFdhivjRHfGsIq8l8QQWHb3/ZeI7Z1zM65r0jAcQZIK2GSe2jhTJhrBE1lHzNOwHuFJYbRy7T7Ss
vLUu10T7opQ7UTQU1m+0g7h2C/cJoYm3NejGT7Zs3LlNlz4g8DzQEwFdKRihWxhjOXyBHnsYiP5x
5/fID73JhOBqepO2eB7+EWOY9FWIeZqOgawCXx69FrtCkMWitGaNWL1isMBFraTF7RDI5THEWD/2
1iaGRcU2Uu8aLPD7XEThJCoTsL3wHafJPdY3kw1R5r0I7boQjFZ4cI8VjRDNo9hK5H2SUdQN+two
P0G06NC5BJvSzA7M5skTSi1MLUSq7neFjKEkJkLzaeYFixmJa1T+ByUKHGHUegKZJRE1lFkq5KWj
ot5zj40bHUtc58MP871q8I5j9OevDvx7m3zJkEb7hDbmb/CUyRjyRuDKn9bsB1nLPCLza/Na3lPE
1cmtn27EP/MDiirMAeJMDHO4W8GXBobfN/d71l2jG1cCjrFfbjmYW/HBGtl/hW+IqEI0bajDN5Za
YMLipMt32cOYe0tMJl+g87mf2iHOyWGmevN0MaibCck8VTVxejZpe3+0VRhHXiz73NOl2nn47TQx
NLcSmoWOd01s5HuXBvZVNLxpjkYNGogi/4UdQAgX7UQK/8672AF9lhrmOWU+5R5qjk3jv7vf3qBM
wn/Juhciquq7kCKRxzLrIz4bze8/HFphwaY9HTWU+5QYLui6HWYUKwFPt4FJSNruXLqkY8ihdY4m
VaK6DbOBLuJ+n6adyPZbH6s/gRlWFDLSN/K+IK3X04MJfV9PwUpSjDFSSFdCI00gbRYckhKH1SmY
ZGhHFU2PQaHYc24HAQtEY7dlI6fSNE0I9Zk/HKZ9h7T65mz9xRLxRCTLu43z2JPrrTuVGqk0B+bx
57iFXG2dgw+KUBLjQmR2NXlzSZDwe/my4xKc2LDx+l7wfy9hR1wxAJ6AJKiPC0F0x+O5mSPsyS9b
NrOilogr/r/7X6gAaPJBsm100qBbjXVAWm5FJmqf8VAG47DRJj8tiIGHREFT0YyJSs2PxUf5zT79
OMCuQXyTcP6RtykIjbHTY3Qf2clx8qXX31fDxCWS1iqPuyZnfWMFaVJgbAtzI7DYx6/xpOFKq/2i
FhfBZUaKvPouOxWHUmXFwNTm8gW5kPZZMd7HfvEtdTSRnFK3eWooGCWQSjCzqTVqEULhGakUEoCc
fJKKz/WkqajmSCwdwnTefZIIm0XvJXPSzlX+OELyASQ0eWj7iAq70SA4PfmBztIxCicNnPW3gpEt
EzVlNuH87No++HdIaCJ3JYz4G3TplbMyp7iGlfG82DIPzo2LW0Bxd1c5fNLsA0Kv4t8TRaf0rEOJ
E/rYOQrKLhEaqKisNJo1SOFnsESgQYt4INJWv55KCkArLK5WT8nH0uTL04H6EGLDH0Uk6/CFa/6n
9iTErk/qb2IVrqbYZqzA32yscXLFZdUeQL7ew44UutAQKbmTUiwwbSmmLgbHfTrjrn7+EZ/cKG0U
9sKnUKjT6PmR30PSFsm3ooNANy4+ht5Of6r6EoxjhYLrF6Z/vFBzZ8oHcE94vv5zSDdJFtkh/leT
1lRvaPTZh5Own1Mb9UOvVu8PkCybACeVpRrK1FaV5zwn33qCmUn/xJhAAkuAaj48KOejubVHRCRl
yCZO5HokQxoTJQajpsvQNqaK4E9KWHTie0cJ1+Mgr/ricf/y9LDx/HvhHMuhYBiwbmhjTIJBgx2B
rfPg4h3jZCm98UyZGTZQTAbGkoyh36qpEwFPZSJCdFdG2HkVai+iG8R9i1LU+YfBzfJjgEc+VzoL
XwvrjUg1jSrkfvcwqE2UzuGY4f/SsUn0k8GYuKxgRlvHrpRiHYuuzMeWX+iIzJucwAmS9pwA+x2d
EhAPZswtYdYXQBLEQYd3SiwN0GD4xJwy1ePC0645050nSi4uj5FulLGUqwYuCdaGj4UrWSr5m31/
DguNFhdn0N3FiDEQpzvUdhpJYVywlc+1vm5yZp9QM5byrihRUiMFKjqu+prwyGe+kMjSqHfrX8uA
6RsSxEc5T/kyN00TUaBS6eFZnQ/D7uoLQtCd4SvgrMD1p+I6Y7B1jZMqkQDHQyCJ4BqsDbkAma7I
f0Aw86lbVDVdGhYDKT+LVzjOHKepDCrSkxoyhR2J0VA4baJHvSfygB/F3g2QdhVZppLh3ngFeDLI
dkPUJH/31Pj0QYbvqtcx8pZGJlqwww3BQX7+3KWPV9pGYn0JRmlknkvoCn6Zegy00iRvc7TnnEqs
YlnpYTb5N90o8oZRuAK1YKcQZS4NRGqtzc2YyRNs6LarlXn0D/3V4dUfy5fBEDBmGTipIe5WzDhI
Obo+FdDWN1IxRJs3PDLC/y0/pNErKipNpv828/6BKK3QofrJRLqgF5nJugH6E3Kz1EecVfy+sh+/
XQGzlEK0B240onWZ72eRsZvky0p8AwDv+P6r88zClOR99ic6tAIBOjgs4wI789/waUdOfysScKgV
3Q26r/UtnWNK1V0bkCcuLuY4uO7FZRpXWx/pb8L6nXE4QtczMg4H62J5v4riui2D/KH62584lFO5
CE7GcGTvBBdUn16Q+mcZHjWLKzxBFHM9RfiuqDzKZACgMv1Yqo6NduypjRwdjMTte1/l0Lnh3KC0
Ivr1ut588uemk7Ym9EpViBN1ZvcOjYmRjXMH2uUceNN/lZMCI2nwTsFnRaVznUgG4ETCfevgCD2S
dCu7glHit9HHvqtOMPKej4uFaJQorI1uiZ1gjezTEGgYYoZjBOhUPiJRbuHsm6zs8fypD1x3rlvr
DZh55d2HqONz7lok7xXeXYCbZjxfgPBE81bqdPVQO/A5V8rEo9V4K6kPYJpSu+x29fVi9YweCXgR
QwbXq0UDZ8rp4+Qn2ymsxfc4YnjNAcdYS9bbnQtQZci8kTrni35WnM1uGQmRt7ZWue21TPw/BEGr
CLo/2EfW4GjHdhd/LcEZ8jYywfemU0e8io3m0xSCeJ68od8C+aC9kFW5cPz782kM2M04vUMyRHo9
HHJcQscDRwVjKsEFlUFUYp7L6QD29nKgwtm2tXkEv67AdLT6/Yth3xKnbnHTobH7aOfjzvx1/fpa
leaffZBtXpUgNw/O7UzQm38k0G7NoEeuELGTYWU/BfHtG7ABCt0bfAX32Mq5Ab/wU1de0qK6RSel
Ry7IotMEAdq75Jps6XfX70WtDOB4oH4DlYxPAM12Lv/BInE5r8wVQTxsHc+QJrSVJdh90ZU4jC1W
2Uqfc3LayPnw/jvnfx5sQCfcK2G2BTfcvwShaZWODwPvV2tNFLQ2WFuQKTWKDFunGKlVB0xJJhgc
pohWWKQXpYbI5SByf+NEUmGnixrIDaOiiRSLF8QQenyplS+x4dDpDtLAbDJqkB4LM1+MCMJqPjAu
0rjQ0ZtaYrrd68SeoeeAsUgTs5v6cQzTJA6KH8b4RyKXAl/nbalm9DIMi8hPo0Tc4cJQpKrLfBme
VSTz5ojlIqes3PAQ7AxpnZDdKxwTicMvaQf10Xy6jYaKKKP57wS3x4soViQGwJilcdn8wzJs/ujU
jVESc7COe1KGoQSa7cfE9qsxJxeo4OEaDoHl3AHHBsbUOrwHAKD7v0RudIMAT2polQMvcaJ5fgJ3
wPQqGwZpvSxnne5arEuqN+b0QezWz886292jrmd+Uw9ceuoQ0ov9sN/eEc6FEDDLpBD3gqrTbzUV
/IjWWANCvjAyDLjBp3oJuINa43FYtPfOgjjxU7cwAdyPd7TnWk4fcHPJTdNoawDhexUrFXHceV8O
lNrQMosirUnB6MHLY/NSqaoOA3ihXi0oHotjEstlq9j0MbSJgGrCnVCa/0HRKpAHXvybA9AiPGAh
VklMpY195p6UXJP1LU+4fhbUPY/5DZMdkTjSioj2Yb9ydSe08A4UQx/FvAhSlvPSPuvxsERMwrJR
ZmA6uVyOP5UZthPgigb1Eu1RDqIYHoXcWOqi0jc1fkwCnx/NP235vgIw1fqHcgAbkHI0nuEe3zrC
8S7rXhpu9fjc6lVxgxnI07n4KQcnfTVKiJ8FXotEMKWtn2dm147j0li0oVtyEBNuPXm1EVG8nUwP
L5dj1WdAtvbLl2z9/5IjAJnCWn0O0nUqj72wWYFTmYxO6MoplwGcRDOemKIBMNL7zP9ox8yR+H98
CG2BE8ERy2nZj4EtG3sGeIOr6Tq9XSpINSWJp1o03PK9Jghk3zaulAY1r988Iz9ittdubE3yqtLW
eCv9RqyDhJ5pEquEzgoFYdTEKZERAtw/omwdgF7ntY6gYnhHtmycuHI176Vh94olFU3Z8J5p2Erg
XUqmLpg4ix/F2eGXZnQBztYOLtkmCHt4BKlydHBgWE94UIqHc/FTAFUajd4Q8QuwHK4nNZ+w74qy
J5vpb74i5Ks1FMV5jOssB1x2+NIjCaFE0L6g/VSgDBDBEUWa/Hv2x5oa6DGcuyK7oAwNwV6d/FPb
8QgdSjPX+q7dOhGXePiaYvajIsJzjp/ZqBDapbFGZph1PKJN27J6Td63ZX4jUWNepSmbo25V7F00
rOpMdVYZJ5GQdB/NhjDGc21aPhbYLouBZM90v2Z+dw3Id6nOITGrk9k1gpau33uEiH+CdvbnStPk
VUT85fIPamHOh+OHtaTUXRh7W1SCGcZ3Aaq1CnX4/CpcZSOj6lTYlTJfZvBV3erx77kGc3EDAqhQ
ulItBtG3eebrAIP3OPm+X/bcsck8EZjrzMTtMbzYZkz5bZB6BcGmwyJ1ieS6//XFuXoixALIjwqn
aDoAGtDuJEWq1Hzt8PCpNYzhAX2ujCiUXsIq2v28omjM8Pj+/P+U+ju+eC2kmvkk+Ii44XLtvXZi
vF4kAa3xumB4qV9mPnO0d/dPizjMeMNwqzEqzhK7BTT4o7NRgTfevdM4FMEwVmO2TJXdEAyCKkbK
zhRyEe5z6a7LNutvH0nt22r9AYz8ujyEZPgZLDULlpdXYDgleNvj4LmW+fFH0cvNb4nyl+wyvjk5
GTZil/Wje1WxFynQJVqO9isCEIWPdu9GitQ8gTH8fDXxjSxKdWtQ9/Dd60wpzpvz556uFeNqw7+3
8Xx9thGW3LzNUgiceVeZH33lFWqFftB8Ql2IInM2vDzq7f4C+Zzx9vceIG6vCrxzdENky+9KH8HS
Amy9gh2cev3cj/0SKw8EJXhqrzMJqG/kRxCr/FEfvD1kgyOOs0JYMWm9gKkaihkWoVkHs9KzCnZ+
v7iZ38IaaFC/c7XzGK1eOKkiapDgkMD0QYtyIZwHhEnrNtRVkb8DtQFw+1ZJDjsoVDb7g/cvmIzm
+nGRfyZP7qdBWJ1SR0bsWXHYKc1xeoPfWo5oum57B4W6zBdDWp+O928HPa0yfOwqTLA03rL8TfB2
Wzs1cHB9+YLuZ0051Eg10nDlACLLd8ZHYjDHfTufAYRc0uIf43BkjuDw4rqbEqk3bofX9xQ3tmjd
+S750VgIFwaXZ0w/ZJ+ExEhb19vhVB0gU1cBB0SDTXKXxULcE6tptpLQ3DpdIbsZstDrCTWS+fiy
bu++Wu0knsLbRoMox0F4kfvPmnCt/zKK5RJEZho5VtIdx3Ec6Kbq9+8mMHa/XUPuoF3VpJJ2oPWV
8es4gc6GVsNDuG7jrANZU1AqD27gxouSvdvVp66utccLXQxLpXWmyxhxlWDXiWWIJCJmPRUccEiX
vbcR8gUidGB/oA0yLSnkUT4FZrcOT5RiBnTFkQJ+HDfrs6UHVdT+aZKuiejqz6s8DipLw2N/DA9U
IzRHsGcoCL72A/p7CUT+qQEU/NKUy5vOcxCmEPN6XNv1ZAaX6IOBLMCvDYJUbu5xZ/9gif+8O7vl
TzxvOwD7gnsjDkQI5mQ0Az01lQLcKqnH6+B5ste6jpRd6TDCUyjAPSbyY1PBt5GMofxdGvuTrojS
VwWf7of6oupRbbKz0RTLfQ2X0vWEAGLnBYLUZ9AgwXzQ+SsgM/G5fueiSzoRIeQj46IJVxZ4pQK3
t7BtIQgUhOiCYDUJTv05h9eVTv1LzP0RfVwTWaDdInOZ/fvP/t9MDTzS8NMkxMY6DAQgSPwDJpwR
I1i7V19TD3sc+xV/8vYYRsOTlQ625VNqYxuaH6sYZb093tV1y3oAIZYKODhQe+jmW/vEeSFsCEOO
6KDXgycty5+NOrWHlfuC13Kwf4DH2yqDuSBPvBkSJNQxtmZqrdgigE8dQvxuzC6BnV+hdd6K+Uir
t/dLjFfGrpq7HKraHYQBWcov3n0op0njOIV7z8bdfpoiIFSV5aBzyhjLuqKo2aDImH45sW1gB+ey
F9s+JnbEdWQ4bGMIz2EALt70xhOxFJGeweXoDeR7AKaCyGl3/Zw1SLTsGrEvkQGU1zfB7FAgF0re
fDAU6bJfCEgeBnATQEmF6XffoaaxmtJcggworcqsDkC0dusGf2RW9W4vEhcGLt4nIOxZVf7Z6zx7
5Qo8siwCBhoQ/tZkHjAGmuqnPm6auHlh4YWRo/IwVJPUVrT+nZjMleKotHql9Idb6FmutNUYvZ5x
pgXtfP107vVoTWhs3VRql7WseSPd5N8RxDSJRUCUZkZx2xbelMnKtueO3UedJTVFeSmKwjqDeGYQ
RVRPW8oU0HMav+Ym1uk3DiLz382xSyo7BWF1Du603/6lrP4xXER/GxnJRDsbONO+L731n40yDYor
6uloGabPErbAEtHTcK2ajDRYXOFT6e/oI+tHvI9kmjQfvUDfnb/SYSmxcL6ZDrqf6DL1qug8Fm0T
oCvfpM8ofIKScweFtgUGsxL6PG19J0UvwnPpwHdd4D3EOrCtaeQTLlHRoZATYrlZJtS9ESdM5x9+
nHlScOx3mpeHxZkFFykwq79RNwk4A27Vm7BxzaoMjbFXiEuGT7NejJ5gsLNnR5D42Y/bBUv4LBlP
qwsosLB7QDRNSIxsWvQDWvhzHrTydyjA4FJ8pjb9oOVK4ZhppCMFG1l5OL07BpoVYhAIGbioM9Wr
lwVQ7w/zGNGzju7J/IXzSh5BUamdHzgROlkWJFXANXiDEPmSSHFR77Y/0yUnf1mucikNNQXgzTjf
wmFmds+T8V8NFLBgj4k6bv15fCRpdj6/dqtcLZZfP1RUX7e8Z2B0aQDthpSmNzHBBgqt3c5Q8gE9
w8MsAlKzUt/BgzyN0pZWssgLASBXUrGlfJkoVq3m3Rp407cf4Cnd8Nx+NY3WD3+fdYOFXj8QZ/fA
0TT0jayUvNco+zi1FX8dR0WuFG+GofauFdj3jyn802fzy97HqdJSJxG8BmBlRqwGEu606euLlSs8
Zej1/LF9CjsFLMw5jzPK8IBnrs76oG++VUJYLaNilfsyKieU7kwModmHUZxS/F15ODMnpJaRMaa6
M9tSN5Um3tbi60k5rhyOINU0xQY9moNe74SMTBRL+vv3b+COdDwHzAbd2eLoA7vXoM94LAS+unw0
/Ip3YQH/eNIRfynSoox9Dgd9iuIU9v+Tul/EgV+4DBZe0ijQmLchyrsVezi0qrekLCERQdQvmGKR
6khGG+jkyWjbGc8xV07EZgHc31qJbOixt4B78K6ZQQy82vjVEfL7hPink0BVKjwwghOWf0WoNQp4
Dqmc26TK7s+LCY+277qtZyxZc72uY1pXN5iXGNRZQ3G1YO0yD+fWhnPvW6BHoEqh7pwIdqesCMSa
SNvoF7WZat8F9ZhHHnKg8TtQ3NcFYZ563CLoOXjdJ390g4kKWQLcZN2xTxZkBCGegs/hxALXSOHa
ApvjWJT8wjn2Sq53SMeleZOyxzNoIGPqCVcCaDmTx9n7Z1d8el29jqlj7Odp4GjrbNbGi3+7nA6u
CeJKNPpo8sQZbNQ32DMKSWk7jeV2MicpiMjIdKajhBeAC1TBVIPdNhlCxl9H96eiynmOCGeJnwYA
uqrLc6luxwrXUVUSklBD7CdKKfbgPjhXWH/sFR1L7szRHp/pQmrsXQIIfdMJOMfWs8xGAID7Auq/
s11fnC+hSZaav096XKbRm4oyGcj67cL8sR1BNwaww/egRVLjX1F7bYfeThIj/MAX2lOZ0oqC6A+c
N0Y7n8UuF7Tjxu3cRQACbcqWQ1FPcGaBtLN+0kB9U5ltJl5UzPVMeKe8FFREzmxpMEBoYGUuIEEB
UEppNbHRtzdZvqTDzIUkhVpfwhh04GE+UnRlMlORXEvYmZ0wiY1QidnXJbdPGimLMjpG2n9ye0i/
tgacfyQ1fHGJjfQaM1j3tobAELvFnMMqEekqYQWBUhmpCgGNrfax97agVmpQrUCRN6lqTIPo9/5G
ONULIScqZ4iZxFczwDN8xHFOkEZao0wuBTLa67lx0gYOt7q0bnlDt3dJIMQ4JPtHbivM4+YNfyRS
rJAbsRmhmOgI/WjGvf9jIbSmS8CwpHF2/GLwbfquTiCJuqz1TYefR8eKRHazVId5sjCT0+WrHjIF
i6cMySoaIgRwjf/9VX0kmXAZO6Dy/IoamWdWEAAUtbqlTp2TQ5DMLKlEG84HPAg3zygvlDV5GInG
OIRE/sb8QObkWSR0X8zJ+0bQZI70EbYkKNNillKnqKKpWeWDrJSFMS5yPJ7dH9Z4eoAid6cBINVO
NiuuFkMBijUyQdR+q/O/kAruqfEd81HxYf0fqlPbc9R+ZGLIp7uO0bJbwjc/SH+BobBWaknirEG2
Wrvd7fiOF0QXGF+dP/g20TNDIcIZdhKKVL1lP+/qwjgwGNK48g9sMfrug0K97Hifnk1FliwJys+w
COUTtLbUBdNZDQCvOKeJGICaWJcwlOZ++3t+Qqs1GFjlRFqMC0BMloFgy2L50QA8Tzaw2OpGz20s
WsuzZ8iZGhExWxQR/Z/V44rmVuGTunkFIdFeGY6ezKctTDsN80jLAcaNQ2kiO6d5NeDuKjx3uN1q
QuFZekZjLF3C/Naovi4oi4gDkYvhiVLZ9bIpXidYULuxII0IGLFAt8cykz1jrmD9DIwEjUxO0CAT
F2Nq7GHcAnGkhbvMqRdd25PcoIMwFBfOvXtpXaupX07RgQY8yupHNsMBTGhxFMy02D+WV6CzyDGL
9u1uGFQQDWDX0rvuMqvAyUww4I6alBtDpwcjsAjwFIuxSwALiXwJRo9rw/ZnwqPBbmY3HE032Ser
5ErMmbc4Tw4GCK0yiTqT/GJCWZkZikxtahTLmC+8SGDieaqwQAHZLVZiVuapkFJX+6RWAp7sy0/C
3zZJWd9HOGVJ5lm9vsffiHIc8XOqsIfU1N1rgntt8UG6npTkW9HYGseCsuSo6O6vZbDLbqb9KLbr
vz5USy4Fb1D4ahBjoLf26maYLU5k3RQfzFa+ZwnyUAMFgfy8KFSyQv4uk1kHn6jpEh6eS0OhDccg
Hn9iIRfZHRFWpSOsbt6r0dBvL76GfM0rKT0wVeIIRpi2EUSgejEw6dCyjblF2De+BxzYPgy86wni
HGXjOpKe5O0jua0gqFPTWxUfgSUZH3aue2I6HE9Zvs7EKft2uCzlu3Av+ORudW17HMTZn8sFwgtE
uEGSUxSko+hTT3x3EehbHtk3F4N+P3zqcV80Y/0YWKkk0MMKRGzS7TkX9BQx9hNVCB0Lsq1UQFrD
WA5nA5BYNPFFlTzAs+RK4BABG+lrF+8YcTC1KayKRzdKCCL7g3JLte0PkEkdqdAhuc3TJbKMrZdr
4mVJk6gqhjDWw7SqWRqs2DP2zNjgrHfJlQfFPEYyUnUlZ1YEDeZzq4HZVEQZJpyblfAXn2N+rAd7
HUVEmhdvL9imh+fjrwh8FnqiaMSD5964nCT1cY/C9O7c7XNpWSnsL2n3XGk7jqHJchtOKr491A5g
fpxqLY0/ORvjbw+zO5mJQt6ghwNz9utEm6t0oIHlZNFE6gdKhbJLtYbKT/bJ8nzwF/5DnOUkDDIK
YrujJUFI3oClTR0zorTVCtYziVaVOlMIzdyJMHlDnhO7sO/R82iwliG40mCKjIXnjZH++FH49DBi
TiwI268aR7POrXMAsd8YdKdS5SsDAGrcj6XfLPqL5TOJVg9FSxgktMFAO2T983vJLc7zQOdrNVRH
+o9LVZCImkmhJTN51W5P1801whn9zxvg+d1zVkzckdxr8NT+pCp302VABl6AAxB2ZU8GfjZgBgsr
6yYV2y5Y5yAgfM8xZVKsS+JBoR2ss7Nm+4kh8JsSvPY9px/KmWeHH5etDvEQxhWwmZwgI2tUePwF
7HFQRFleESzavBlTBte+U0k2ZYCZnKCKNjktoTTsESu7TxZmGgNAK/8JDMfxmcHkcVqblcd2rw5b
8QRjnbXusTrXxS7Z1X9RI8U5dEahxJawFlFTWfg1OEKvsbQM7ZxB4535zBMpUUe9b9NupQ12kPJJ
KkJ1nw4sDK+LZ1E2qOmDCHYdayDwyf9EfnRDv8AfWPYXZrKoplCLYsB9k+2yg0lqWb64+Jb60Nt3
hdT0iuhmvmogOLFi4Zfiv9gGRuN1bl53mjA5aItT5rSp/xNgzLq+g0v5qSUANfGIWZExPtGAcMQ1
U4J83mEY1PjuOueLZzVRVAzfj6vkBHUmUz4LaCyp24hoQCSdohzW88t0RYw6MOVBo4ly16eJTFzs
eKM5plOAgxZ2nOhGypLGwyeZSRmCKGvfHzeC6b6OVMeW1rMxxAmgE+4VsEAqT8SBWdpZATMOxJw3
kHODRYSw0hsQZY1ZQTougp3j2Ywgn7xAiD+5+e/T3CRvl/8tXyPp1fvVFYygREw3n/sGBSKq8U+f
GRds4QR0vCrWMJw6O+zJSkpdT2dw6FHq/5G2QfjUOo1LG9vWDeTG+F7B2n8Kp9Bu435w44Xjt9mC
WWNYpJk+C1s25YRWfyIhZ5RWml4HCqdp+0j83earYaq4qp5g79jcsXdU+fiJ2NAr6MzIi5+bcO+2
4/9hIrO8xDWGv7pUGqhV5IppTixUJPV5gHocPa5+vskPMZpgNYZmPDf0tjrYc16p67BQ4y+vkXt3
hlSQVhiGIdzg3Cu+gIIwSqaYjxlIZQeoGwiKLAKJp8QcrJxMi2AruLlHEUAlz8t5lOTuvEvltDao
FfuBDJTc/qLLuvHwu5GiEwkSiONOyIBpJjDGQJ31JWuL8o/xiL0+cfQf4Q15HoOF7ogpn2wtCSeN
LgtrXhFDENFCsbPVGxwiXpMxH4dZSfmJz8VbmG2XIChCx/3jucEP9qEOsKsWaKdoL7Lc/GJdX+bZ
hHCSLX0pkkxqUqF4Uaf4QAbNsNg+byrFPaKfUVYWkBGAuW3zzGZr0UHTIFf9k4aXcXrqr1seEmG5
hhLPOv0w4vX6NIMoIvHZcZXKIoUZYL0TsSWWuL25lDNuPbfxXbj0i6z9aI7tC0CQPPyxgNx8tVq2
FBFd+zfNh5H9w5QYWLzk57RHFyEw8wKXcWrLB/e//SqcMwcJr53ZwjTRZHOUQXwQ0O2uMZlXDmx3
x9qb0aUDkxY2nmPOTxnr6VVc3PeWBIczifhaU6f3tGA0Mfe7eXGhh+0frTVJEhJHSZCCssGeLYK1
uureX1FeJIh+1jpCG1pCY1zSVYP70kKWgXTcLH0LWxqS14f8/Qyau9l9NVnf2MESazvJFjTT2d0z
ZoaqZ7UoXWuY+aS0tAxxmuQU7TdiPAaVeSYyF6OM4HgFlBe1QYfnplgfPBDUeIUPz1DwGVEx3SFM
4e8yh39Pr9HxE25vUEUzXcVCQMpxK4OlNbvqPRNIyPlti4w6hvPlCOSx36f7sWrNz9v+UrQLjdgB
1Xgd10uibtF9uIwQfAnSG4LxCA6JvIxT0StYqcv6gvjjc+0iS06i4SMOsdPq9gsZyg7+2Zj9oOTI
5aCM9UT2RsbJe9Fo8askZxq5PMTHoagdvaRFZ3dQPETaBZXCK7y9ixhLg+r6O3cvR4Qo3Z+SZsw9
oRAyWr1MBHFKWvSzbOkRq/9hYXqkQj0z0BGLxaspDtU7LprVkuqGp6lHBhHYIW/NefkFPyVzoAS2
3n+hx3IaJEtZuNzn6EjslH20jQMIGH3moML+5f4WjPNbLhKfznAZYs7k0QDG65CIrDslbL3Rxca5
9zDX8Qj0dy+5+a3YmTfDoGOPz0SnNqXU6puJ4kZTJJmXLq7mvHw8cFPm5qWMTMKmn6E5s6ZZkX2u
SleVlZr4t9zGP9kq3fctW+BzGZZP2cx9pX5WSxWrBOHPRDrwCRO9qMf9dooJzu2G4qNg4KI+Hhzq
Byje6OlNsRfo65bcm+8DU3rDkmnkzPi2IukZls2stvupQ3DrIgn5qKs0YUdU6OnUWTpYqHMAXYOb
5RVfJ3+CVqym8Ib/5+liizV4P8i7N4j+9f+EFEx30WmHE2oU8jYeRAb/iDYxnTcd7Li9VEIl95tQ
2QdCnf7OAn/C6FjhnyfriIDEhVdnvcEKYoLZZOYuHBcgdfF0iNx/CH8THKtkzwQn005TLZhWWUJT
r9+FEaD3CZGegsjlsIH57GIeNZmkZyC4SnuvldjEqxNLew9jSkFo4SHyK01ZS27mhjNtIHewiKtM
MqpCzAI1V/ygIeCugoxu9T6DFbVFKfQP3J8Epv1c0LPwSMlzru+YULEGs4vzcotbX0Ioh4aWlWoW
UQy5bbwWctnvCwJWTV5AIIs2+HAZqGutzIJlcVSsmDs5RLp9MKnENNPmeFYHfxGGtLyZfQ//iuOu
9spd2I+UgpSXfahW4ge21P10FJL6iXSXo/9xAahwuRE4wCDSMq7+749e37bMwhKTVD/SnClbeE3f
vM4UGps3el4xuvvg+x6Rhra1cnB+QaPGgFlr1dcdSZyzyImbEm2qXrkByisyQxnbTsMupTQUZc/a
FyoevVVgHztopAigwj/w2nfm2EZBnEUfXejmyuo5gDrSibusipqavF7t1cPpBMdQQcWzxj+SaLEo
eMBCew7CnwagiOguS1NWrgo1WD0/eoS3qPIr0FNvb1+O4jnmNCTNK/viNy0c/pCpq+WK05ioEzQH
+ooI8px6BfqWHli6VaDRVJqINcTqJVrWBuWIxCh1tCK2uQBLy5g406ZDD0c3dAljxWZOzI4Nrdsg
jnuPRaVvWVoOAinyWWFSJwILP1pzDhCkx7z2lUIzgEuwnJkrCS+23+wRWeG1C4jlv9PpJcM2Wbyy
rhJbL0UgVJ+oq21P40OYEfru3WjR4TucqpqCWhEj2uGO5FexeuDL8CzFTsSrkiAHwcW1oZ/tqx6g
Bfvm99UWuSm8IWh9D9xlDdtFTI226BJCIFz39cHAOI6ll1m1oG1mgSJ+zvHGhGkRAj7m4+qMKd2q
SJ3Hw35QB7wG1HwlTF+/eczK06sHjfBdT9iAuImDgwG+DVBsJw4wIpXOlzkT8jtVAF8dnbTwKlg0
2T8EqE8zKn3bnhZClHOq0ZtnA04cq0wGc3B7X9R+LuHGdjIrk5r8yO2CxdmuAetJJGdaFNHlJTcH
+gHw8avhFfpEMya1pkJ07yAFAR3PetDXHl/RBXjawOgQ8PKYT490UtK0eF2JCGDiPnGQ2dAkenC+
+uTaPFCwh/NpNXLpevniW8HaYN6JXIsysdCq2WAOZ9oTAC2z+NppG33Xai/2+yJ1PRUXYb5iJ4jr
U0K/SHk3gHdCpVmsyyLcoge4ZXHoLgGtjnAsaQ50Ft+Sb2sAUpeBXsrQD9Bze/L89yXQMpHuc/qx
e+MSVs7Tv2lB9o6+g+9XyTvEDW5RgV+Xw5cn0A3Znvxu4aNRUAF+mC7+fysboi66znLh8KlmQ4tR
U/rdNhWuJXiJ7qWFHuF+6HoGaUffrCoZIdWDpn2OOVnVTIibjkaUs1CXttYl/yFq8KpU9Oz/BYiR
Nf8sdquBTV8N+o4arYHDkpqKf2NvmmmwM57RBCf7xwMkP+bi2Iew4iKcGBILeyz/sdUAGzLKhhGI
avSBusHLH6Z0ahPBl5FoCgLcO4FDvelMikycq9Qqme3m2dX1zd8aVYschOD7ObFpzpEz3gxzHTvn
rJo2sKtadUybrHIFCiC2qIn64SxncstsiAsG4Yt8wxVa0TPJtlUnaYdXn3EChbxEbK1ZCWH38tvR
qT9xr5T2H0BS3dl6LgsmHEYO9VU4wuPrBQeIcAuFYTRPING+zk2nl7NTAAjMogLWxk16p9vBG2IH
vgs941/w8wcO8UeMGiKUiUOo7hz9J6Ot7SBLeuaPf+SZoNaM0zBAlwwNpusQBTqALu1pGTVKcxl6
WMAaoiXkvoDKoXXsOSKLwGPWm9S3YVrGcZ605PUYT9g7ZyQOwDjs9gWCDSnfYyN5utrqHESAXKXO
GT9J6hNMsO4HzSzf25HZjk5Jo5EOsd988mlLXX2RdYxuH8y26uVStQ/rPeyqSxFkhjuXdadV7acm
GYujl/vypWbD6EwrpgdhcjXmPX63MYWE/2YuZPNFV+mLlXMRs0l4nH1hhLbjmIaw/Pd6sqeDWtYO
rBFo8ZHOqTrh9+UALKXo3WqUCNtfLji4ktJ3J8jumwpHvJVjWHaFvJ0ZImEi/WqqJWm/anguaL67
tSiUDBtpXWQyyn5fQpkfBnmt5PkDX56B9TGIZbFMt+4UqfZINC9IR4GfvSJJi+XA11MEaefFIZeG
O9QsDisup01ZaXG64QDe1y2dzYtZSADq2o09/8RXsw50G/BlYMDGte1o6BhlqBkBCu6THQB/g98A
KA2ejf4X7ymNEG+3ypkNEzFy4jXfw/Ke83BONU+X8mtlu2yKxY+N2AUzT8uf82nUrbJEUjpyxkol
plbyo0+C+XlB/JuRiMJN47s9kRKpTQujj8eh5bWqn1uls6fC7pJlaG3qkYqtSEGtMcgepBAzO0tN
xBW1PqYZmA+gvWv4Hue50fmG2PnFfj7dtWPl4IVDC+lX3hVAR29XiY2f8I6pCyL7W9PalMU499Nd
T425SsAv5VlCLBVULsegpZom4MFyCDrVH3tamcE3wEaX2JAItnhMsTbMClyGk+TRn0SBBJReST45
6lmAXKkxCi4Ttm6vIBbQgPEWxYyJvuxOGTM/AgqDaXN3J2ao1oRBozhQ0naSXRNni2HOACuIxq34
bIpad9oIytphOlg5ns4dukMoXT2mc+NxuR/OIOqSjf75v+tRCuUdJ2/4ebKDdNnDsMXiUoX+XLZe
RBw4EbTjirELDl+0BXNZT032ass5VXwDJaXos1TbCQ9M/fKUr41OL0C1jdgIoEzZoVY20VeWIuBd
xsaWIk8sTrkdeIN2LEQnnd4sBbCVVTzCYZxK0fMJv9uWroULoQXQ7uKJW8+THpa5hpu07Hphczw5
UHqT+DdAVsY5f7+QZO+KxsGEI05ZnTsOl4kHDnubJmwNmqmNUNlngiEtRv52xdBGdiY0fYxmMp2x
at5ksMpDPP1qUDDl6UK4HyiTatgc+hJkrWkol2sMKOrPBcwpNPDqq37L1LQBhtmLbMDGj2yd0XiL
iQKSLwTYrFcfXZ1euRkKoLVyFtaY0BDiBCDaLumZPJEa/xiLAnEBZYHAMmthfcchVBEGiz988qhb
Q8lazL/GHiQkYtXwPoM7ZDv4DkBfOemeNCrK5yGIC4dyEtCEPPJnI4VqpRxi4liV12beD0u7DdXZ
wTjs/RFcjYRyivL5Yu+/6T5Lq7xYHCF8OAK0IlXVtKEfHDIScvx30X2rVeozq3FcSOontCHOWCSz
zz7JQeDdh4EFSAOSiR0rHCAKtHPXahoJrMIJokIn001ddMGnzVuw6kNPOERSETUQ98oROnJUhfOY
S1P2QkNOajBTj5DUwGyqTphcl58Bc56rwp1XjXuye4cPwOkP91oP3oLIdryzak3Jcmk4omEyNrjT
JJi6Lb+29EOai4fgPNRxt5QcnczCmlwjKGI1NXLBYRU0w6S7Js2Czzg+QyjmrV8a9gdgifadTCC4
Nsi01a/pa3sdEXzzrNHj9SpkolDA8iRn2bqI3/oYTVoKA2Y/+Xd2NhtIRmHUxxuXkLsa5NLW7qF9
DJxvmhYZ+Sz/ZXNkLX6T1E9wa8NyvClWDsgTVeJhIvUqr2PBTp8rLtRDLPsMkS9g2WPZJI5BztP+
9PMC1nczIJvJU+CaVXM1L9sdbkxdJbQdvj2IO+m9Yq1+MsANt6aWVwuU8TE6hwa9Wznr/FDwnKaU
M3x9nTj+3KoIWLa59dHV8JXOeJJvhHmwjbelMCW1bWQJYCWoUbCak9QUKfcvT/krzoVVZF6MFqsv
HGGurx+4CTC9Tmtuz8uDFqlu5o4acYzLiePWK4Kn6N+BULOyw1xgu5CjvD5g/mr/2hXE7IVUo5FG
aTKqZB8bYSDYasfWIh2IE1QMtIQ0uEcTdRFqBMfPIJZ6S6USl0VofLjYAgxaclRvhbQ1ZdrU9BR7
kTNnvqXTpvXWyYCEwa1hhEx8wUnc8emvxnMzlf+RhzCI79XJ7VNsGaFsjRSxbC5ugLbOmT9HiTmM
s5eFBOnkijmd1TNCtfSbaGcaDoMUHm1dRF+hOC3c4o8DvgK04/dYLE+2hn7acJArkEodO7BlC2Ie
JP0KgxbZ5CSQTlRLFc0VH05BNfFi2t5FrH3u2Gu/FAAjZv5G048eoRxs7kuycEGYDV4BOY7rXwnr
VVYagPsBGyNOSxiLpxWovfO+GGIrUoqP/bPdU7P0x1EasRNRVWYI86kjP8C2pnWW+qOXB/308qA6
18smy308HEgHLxJqECwTreB0DeC3FQt9SVUy9/3fpXTqhuYICJ31KxKx9dhuOe6guP2Z0mfRwqPR
vYzI4xaZh1mKNffXg/JwgfSn+BTkWO2bJjxRaQ6l7jjcj7tC8rPb8Yo5sSlH2+Jr1kTV5xORA2o/
ieSKqCGi64HZ4jIpj5LDAfTLGR/9y+8Hw/n7e05MuZKE3LleP8aSa4ca9W1jlooK6N8qyuqdyWQf
0zA1EXaYm0+00ND/5ZZl1Qb+jYcAxIlZpRfSCMkdyktGq/OZdr2V5zPHvx0LKvUonJwSPF82qJQt
6mVWOSsgsQ5IwmAJsa/cm85N9m1UnB4RozyUk63nR5ssaFNF24sWZkBXJG3jcGMsNuiZoroLUL9O
M4MhnN8HyFNH+ZLXWoVPuEAYiKRninod+cpP8sJuCCylu4QvlPUZXiAr1McjO2rhLV2kWrnc7QoO
BgiUAs4oJ9BbyBfvjew/nyE4KLksoCSFrF3yZuPEb4CYeHwP5ayeD+4mvn37uc7ny5wiTlrkxH5q
cL9kgqqRMP1MYOt+dIMQuA2VACK/6T2B7W0AqpxBy8sw9Insgz+Bk9gISq2ud1GQ2xgsHX+6YpYU
B6bHmpr33XqPp4ZMNIch/HAnlki9RzSU9AkiDERQe6xy3DM4QmBe6Bt0RXVF1wKkSGA+9/+94eTN
LJow4lc+epZIB2QhAUf0Vsd10PCv0fHvVcMR6qUGjQbNWyurlu7ncqSEQ4gO3333M+6WaiBo1zaz
DpVuZfhO61MtmlDuY9tZaiFU2GzetjKeJ4rSup1RmZ8QaRkPKOeiUoEXON2m+jkPGRlFXhrjBoiz
OsypsSZS6yDhljOAWRFTPBfjzYJzVrrD2obzTl1f+OczDBS7I6IhwwOlAR67rTZC33Lp3EEIrt2F
cX4IOYDnLU35Q/rZV4ZTAPzBW6+GFHXYC1eN+jSE30kaB97VUvw17loNastHBuZcLxjwKxY0mNPy
9AHADtLRY99+at/RtZIVVqArIDTUDqXfgGdMI9/QHS2LQPcJs272Y23HY0Hl1xWPCLvBn120cPdJ
TEj0Ii1HNcy4dc/qtF3NMVK9JlVs0cH9hh7TiS5nJGwFH/TSunAArZgOKiIE3CsnLjVMpGNuw00O
w8flJQVctb/rBwAPNwGj3rGuxsUpIKXUVnBXLkO7MSTLH+qHh9s1N0oS4gJGIaxJuHnuD+d+n1yy
Ef8qQMCOyQCrHzWZXpU2y+u553q5PhHIXjCsBqg0AcD2dLiXwUbnc0Xgg1DXN3x4kB3VdEvZcUnO
/Icv22rBJVbkreEsgdPqTJb0zID8QkbXryMTf9W4Rs1uTYTlZKnFLiPojy2rGCHAtAsAXxU5l6VJ
K0nl2ZvQCigpiiQ2OI6c2zMBAj2QiVkuWygLs+Hw7sffQ0B0nKCfzyfADCxbzV3wrfa8DjO69u7W
BzON2ZLML29gWthFJHobIoar4+UMjcKBVUFIj1e1/M29yy8ddWqjZz2k0PrbxjQpfuCfYPuba602
DdET83dPswkOuQ1jCVQAnZIbfdnuNLYPjYeWC03NmVnJ/TbGE0OFcr+PYxJGiTrj1ge9yHuKwQVa
6viPWt6oDMk4gzPeNFkTioC2C2cFgqu6sSUD9qi3x6fa3qldSAHahO/QSmDk/vLEmriLC226SmS7
4ZQHiInPB5xM7mWdkQxLtT+h5gtWTrPfIc+uxC1gvinjoYkzkJNGIC5j6+GMGLZmDPuxdj3dQfnW
gNwRN8mlhZU7EvvTMVCQ00V3QjtgGm99YWxnijywfRP2Hl2tIuXb8YhCRaNVDr4J7q1UeCaxG82u
qAhZ7++OrWgOAXhmEPhw4eigtzCsqj3OVZI5Cg0Fut/UFogh9GupWbciscOcM+vvE/U9yNoqtWQT
w5LMbXBXTQhfb9IqEW/+kf5TfkaCsbjWvkds/M1+Z8sf5HuefbDTPuSWzVNoIgroCQF5Gl7VEQe+
EbTwHu8VgZstG1h1WNaVGd+USSXLrt+U+YmY6WwG3BMza57/aBglxeoHS/JRGwjsKQgSwBwCM/ga
Uu6IdVhhDIT2Fvzby+sk8AE4Jmt5g9OG+R8dFJtVXKhJF9F2Bxw9f56dQAN1TolINapbbsTWDF2I
7VBWGGo5EbbsnWcGv6J9NeBQKzShvP3dM+xzHgtp086eiCW3o0F3kLRVq0ilOv8KP1Mcb6/9Q/kS
3J8pZSRXTyHZ0OSqTfUD+sWbGCnoCb/kVae+F4JB1vc0O460JDpOYiCA+zayz5RsZnn28H3rIsve
DE5Z6DQ7P15QHnbohRP7UGJwMnhm64iLpoE0J9xQ2g/dTCW/9yRG/6+uThvtSPlSeQNp97FcdURI
pt1b0QntrV0fXYJdQDMj9aeBJ23Pu9guWg8d0rahmS8QGJ0A7O+BylhIl2VU9LSDiNd/J6Vu1Dw/
vmpLaOP94Rj0pPpeJpvkbILdXjGMp31nYiHrm6gMtvkNS2HvhEi2dnM7XayH+jlDQ0sjAV9bWh0I
Ai7X7u1zhdXoVFuLYtOsYu8/JjSU4I5v4RhSgUpcY37kDlPKZfn+Re8sV5685bH6SRD85p+e+Djw
JJOpkZ3Hy3xz6IQV+X7lO4DOHVxNP0ikv4DhgCFogN4S+2WKh8o0XQLqGf1qW30gdd+9Kg1bQy/b
unvJs1jBGx1WElb5gRikJ3j17StLfG/EiqUUSpfemfRowoeCDDjOpYb8OCRGGIXz4dbzyCXAuKSG
gaeKjCZ/WBPq74umgED9c5ddt+H1Or7L7+IeVgqD/J9RYPLKZ6BguDaF1qrhIjoqw31K00j38HbE
7WWdlJBxSk25l6rkrMkyw/PRJ0vrwgSkJBN0Ad+MP6ArxSbh+i5TugYma0dwFmED0WA26faqg6F0
+2ZuX0LKibvweOIfw35rO6XCrrAxDKPf0iXtLp8a46gq+USZze14ZQkIlwj3O5jYJToO2BNdGNKw
JsmJQtVYorDxxKs6CAngWVuv7CZ/dZlGZ8MBP3bti6/gcHronFkrAfWB1j6+ajmIU27QNDNCevKg
t1czBwDV6xXZfNBNaBVGOv7Wo/NonlrP+KgUXKZhP7l7bXx+lPmENOGwHK5Y0tKiy6RNWAqH6sSD
rHz/gSlB+uNGmf16GqcKY0B1O3X/qdNlGtkET01mVBlLbMHdWe0TuC4U1ogDSAQ9CfFp947+G6aR
XrhuOf+BQXxdwtQYo0fNrwyrompqHcmfd3c76HmW6ysYdJZDeZL4Li9wCyudQckza9VT8jgB5CAK
gJNdwHK6B+cBNxWs2RO4+uZ6l9Mv0AGjqSmysIeJvhVWwB34OSvuwy4H3CKvNFtuYPmzSrjMQ17i
+frB+wEC3v5njdA5S3VWeG+XtwZDnHdki+prHqGCAylsOhmMGmG9pFt3RdgyOUXk0yulIo5xx6sV
wS96nZPnOt7Qdblwt0Tz5nCsxm/PGOHaoYcDyPu3aPnlDJzTT9If1wtLDHISYZtjDysjbLZ9lPQB
6Ok/jGwEutEZvuve0+vfUSIFTfqQ17puP+jfwKbGtJnFJXLGqx1zKdx5V+lJjB5/amymtk1LKVF0
IA5prWJROekLhuBRcx502GtqfEGZYALD7WrRgFMX/2wzUBLlVTDH0gq91ST0h+CiRrbtSnez0hVb
nP/vbaf9PwvHucTP8FsEZOd0pbigQmPg4/+1ubygbvIfCdhcN/Uz4g3xFyMgDWj/jaVRlots7SU2
m4KnttXQWrXm6PwkbHyz3WxCg66FR1u3xpvjEypKz8Yw3YexDAehYmOoWStknQGi4kcvtFY1GAAF
j4gmEnB3uep/XlwYcSbVMXhYopjtwPGKNvpZG7lD2YR0TzMmVI/ePdCctBswonRYHt7QSs/YERXn
QgKJew6wlyM/Y1VlT9VEwK/uN4aK+8ex6PBz3/1a01DOwXdBrfxro92HrVGWWf2Hm/REwUSrJZT8
ikbox1AP6TB19+XAeOXsv1zeNQ3RMnxrVwnqVk8Fms8KaKpcLPQJdZv3tS1vvW/2q3+SgAPDFQLq
lfiPdVp9PBq080k9V7BS+yq1/eeTtZqC5afJQbp+7jw5L004oy2AC08R9BHJaiaSztGu8URzCJW+
9a5fUdPlIQmRlPuB25ZI6dHgLyzg91eVqfTy7X1SHK+CvR7l9TULMUGYhQDbq4lRsYxjck0Bz8M2
ZOjqOtFqOjlefxKxWsJBJnyrOzFF//4FvdLICxkZNZq9qaI9i96k5og0eM9yv9MmsFB+lyfxaa2q
sDfJ86oCjFy/FRDe+pxzCwuZklUWCZ0T3wiB0M60MgNeyKWhxbY2BPntpnazx6o18+dMAIWu5ERh
YKlnTvNBNn06Waa44VisHecb6j6mOy1oE9hWbrPJZ7ZkEBsFdPdz09YaU0AJ4XS0sLZDRiGL6eFC
W6/mxz9jJM+yxJSemV53rL0U9ZYu21BNe8/i7+vND9kDY8RjGpaAaRRB/oWpBaxzhwvyJTSSIXBE
RXNROEvgH5H/mrjOe9VdHT58Hty+ZX98OMXAy8x4//zhBZYyv/UKhB//TlEgIxcbevuT+1jsGp1A
IKqIxA7Gx2n9/kK32Q8RZ1kT/yZnoBNHArZ2i5WQu2LCz6qrszf2TFbcimeYoqvHfFAge3UIEWO0
t1w433mh55sS33/xZbb43Jf7EjqivNcUvq+OGLSS0kaDjFZaC5kAR9M08oq2z4SRPVgVgiHyS/c4
gG37MGyIDr2/aAuetWBHI/QJQL+sdVmigorDIWf4N4HgkQsfWI0NNqp4BgCGLjzvJ2S5dT39O6Kc
vHJRkLdvJMp/ieFE2dK2VEomGFH66wOp2RTSXZ2ulYVhPYxvDgiyraXj5BRYE1XeknWRt5Hd+ZvE
okxqJRZQU70vXsKdNgwVOko9XcnItfPneqo5kYuobVIddMSdhvuZJD9L3EkjNZDKzSWXSdUS7CvD
KIEGlgQH7j7dtBgXuC99u+DF/AfJMISNri9YgIplimFgvjE0nk9VieB9/xZ2TT+YhEhNUN02xrNr
DoxPBEwccx2EWsunldDmC+ty14pI5+VV04NUhOLgDgLmI0t5YwyggMAGocoEZ99uyE0QOW2nBOgQ
6Ad0HgPcHsng7uWYyttLkdse1aev7m2MYuq/AGRcM/4JFzzT+bYHafB4ZPf3zWwjY4BSNpSFQvPE
ASq1aMFzoYobWfpDgKMU5S2QrO2BBPEozhrND4c6dh/9eUtQfWEkLYxhZm4dBW812FYy1OKHQv0a
iMIQpi1EglCriEyxX3MChTKc0X54AmYCdhAuHDwUj6/58c5J4gEal9nEzzRuLo2b1LcgNjHX5ej7
1IfBkCdMZoG5BZDqHh/72MdRVIYAdbcjyt4OWCeCpXVetuCOjTTUcOylgu1Clx+A01gsjwlmy/Ii
mtDkWMef6ntDT7WOHoCJtNfVmcjuOFckdSyRVIQCWEU3bnXPzhFmQZKhffn1Zitrgi4448Rvni8B
Dni0Vj7fNa3qLj+A/nF/t8JEgQ27fC6eeGNrVOuPF1Dko4hjYJD2vv2tm8aafmGr9knydwnzFxZQ
HEyhHcmMKP/+qKYalwLY6hR0Gi/JcJ2nocqTiawaMaFCeWMl7IOHv6cjG1x5GHjCB7461J/pNApx
ubh2r9dj2trGd4x4Cd/CY13/+u8RKcDaSfD4SHqtnS3dfcDXc88O66qxOxYMdd2DdDhTvsynAMUo
3zFvooYzSjYe8utPWFsgs5U2Kh2ZNIaf1RiUnVjgICiHU6SIxl0rNV2u5I5dtpgabsyHS8NMC9sB
wB7P+s5RUCearbFT1qhACS1/+2YqZ/uUxzNcsfIhvDCiCVEmtydBSIVfoNq5URZ5SVVbRH+2hflk
BToEnQqtN7lfgkKFI4PBeWOG1eh8mI2uHuIi97qytN0q87MwfBrwf2QAlq3ZE7O61GKIacFwV3E0
uoRpFKy65MuiK3qaKI2f7h7tMO0XMtCpzaCVOP++FvI9JSelueG0xZNLaA9cxGYuxpzapPy9Rtz/
8wE1I4SyXvZi6ffiXCNGInNS6BBSte86jDReFSLsyCcNiGVnj077pjZpj28sOuCNBHi/gZh4f9O4
AlwJkKkYCTIq8FE90H6M7NsxPATkMatpUCXYUBnIAo0erCZYuH7ds+3A6bVkt6jodndAh4YZsE0W
ew8FWhNDRq5T1N7nLjQ2M82wkVmn09n0uExKw595umjT0uEIZ5QJfJiJMdFnNl82KeScoqiWCZTb
zwetObm21sc4FIuZJ5h6tgw366wxPqW0dMOn++dm2kAWAgwQs36UzmnHZt2FtJIbto1r+YU2NkeU
c0YZTmO3NqiUyYp0Y3FMBejMvGzXz4j1xxfJObhQVu9YF6F7mjd/BqAiTIaNdDf277jcFOgbhf8Q
eRNxQv7iZ/SWeUgbtrEe230ISTwuC0OjISMCg7UJJkaXofhRCE4yveZPM0VVy7wZ9uOHV8madfVE
OKO+yYxA3lnsGL7HRzqopJPOVqmhbytoX3hVoaWXc/RQuGC1Oko1Sb+0VlkFaZ9i2lFejQKyife3
jxKvsFTJ7oClIxDMkuuWON/ubBrP9GNWADqxWyVrSIY22w3HFTn9bQjqm+yvd6dD4V9xPk+8tK1L
qf0eevBudLF5PFxP3S11bhFKGsCXCgUcJbgfGKcGjXaKHfm3aGuJ2XU6KShqW2vV4AXLOfvyZWvw
6Hk3aEo2tcnRRwKiIjoFGI+oZFgfteJq0DcLmSvTO/OG9oakxXv+G2O6g7zKfcD1fu0TMFET+VEk
ebwWC5i4QV0kP6O4vTsvJ2Osd53H+MshJ6Lu7xbNL2ZH1XLsOwORdpr6VKWgtuRIjkIWRGcO2UaB
XtntL6EqZjBcVgS1OiZO0ZvcsWa4Tge4T58/5boH7YiF85jBm7Z1K+XCaV/RDhsPnWQJOXcnMejY
AZ83l46DTBdK2buEiLZ9tCjFB7s4v1hf7aE3tFfssDUqkmh+qq7+VWstv4b+XVVvTLsKzVk1Au6Z
mc0fYHLDDKNVuGV2bOhG+NlDJba6pSTCbECl3C3F0cpiUpiaK0D0tVLzKHry/oxDqK//i1VPijUa
E4kMlqjSF39YeorX4OPuraUzdxb8xpYGkjVr5jYEoGfcBKc1gyKnjyg9yah0YApeJLJaeEiQWe08
Ko0XzxfOEuwa9OX46FBWTmb0H8HW9HJa461X/HLbBGZ+u+Gd1ZJLNbckExD86a124Te+NYQlA28T
ZwKYBVMqyX2rEXKakd82Fn/5qHnMoNy0CewX76/cZiFHbprQzswVu5xiDYx0TEVH79kfzk9NhuwD
SlERMsl+cN8czhoyK7yJk/0DQX/zP2O5dvOni0bVInFPXc9o5ZAh3VCCgMp/19naDv3Pkk5uJ7LO
7nlp5nL73hCbmsyBBwC/BB198XkBN6DvFaqD8mPKmyhf8kCBBITgiZB9FFUogcPlIGXwTKddCnQ+
TJK6XV8l9SivCu6MaTAUZYVvHFWwZjCtVX9wel8XSS9fuwAULFppMdwRqBEjG11kJdSIBBSMMIbP
fegSDIERWZ8Ej23udxNSUSgISfgFuQ+cSU6t+S7pN8LzQTKoDxpErEuuippZO8Mqi5utOobNkDgY
0QOXyMsYVj0fYxd6rIZUw8/PN0Gr69DgsWtoVtFANAwsVXTvXNkcEOJeSCW4ejdpz/gNR+27mhwV
3JUxIBFFGc3CCQIAcyrfiy60JPfFaj0u+mR0FuxeG9Z0EzfUb2+vnCd8LMicG57T35Mjxrc4ximx
6kgn6iynHlbG7jDq2Nbua/xSZyDP6vxzYMgApXNTKAEkhot9ZO1lcNRYiRThG54lmlHLFCXXXoSK
b7NyWJHdAFiXQI4z8zRsr15E9sfuuJqTvoWkfNxrTbPBfZSSEU75AGVyTPdoUQxIm27AktgAA6xf
1RrTUACN8ZIaimIUbGLjeGw+YaMIBjaPyRjr514luQQdjjbJbX2qQ7lk/4tq8ZpbOEUXu3WDVJ1v
pBWPfl6wjgzehaMu5Bqu01mDNbz08vkMpREHbZcbbLUG3D24aBMQzH0RSvlCUNDj0Nf1Oq1HvJmZ
DwnYGSIWk1Frd/k7tOAjoTS6eIr6Qg2XqsFacO1+Ni/Ks6D8MwCYP9a3dRnGx+bZlYP2Y/8UA4UU
qusDShMXk7ZJsa+JFUOpJBdcYcffJbtPevZxoUqkfcFxyZwFEvR3u29mJYq6Gt3kF6YrYdyr+i1t
DolRYgiYz8RUjKHxT8nCtz3d0gH+Qs8ckauyPa42/sztP7Z0tpzVcRaLMYRdJ9LdDiruE8+kEvz4
kmGhh5uwsCPyV5YdTXBVlaIirRV/xh0KpWtMdQL4dFqLQyJAfg73HMo9oTrG3+Y3MTv86yXziBQu
DcWNx4i7AWZ98ryG3nhlrqW3AZzmb873RUf5+BcuElazDFnfqf0aGEozGEWpLFJ+zp49/WBzWD7u
f235C4uBGBvvI35H+s3DPI/8k+sEXDJaE2HGszH+L8JQO8X+Uf0AdyAj0hihSxwv21vBaQ+2SGKA
NqymP7B6kf+apeWFqbfbiCjbnTbZ85VxwktsU9D5h+Q5t+w7uV3BHNDvpcBP4F5QSjRap9fXCPtl
6+WgG74DH8all44wyIWR/2hWSxreL1+5BiLESQ4d6bHzBT4IOXW74vU1nAYVEBafriA6mYVLi+oN
SK4DZyHBf0BY+LBxtAvtcA8ZkgV3nZsnOxoUdVpSSUnlm019pmC34XhaC6ZuTvTqvOIjRFJYKWll
tbvZaWMx3aqQKK5iMVO/FQaWVktShHjml3MQq/oOHBTBW0/xXNpGcjU4wDiDswi0Mr76NZ4EgOY+
MTRrkuMF5UDAdRKN7STc4v4WYstF/XI38HUE68T2jy9Wpx2dACqsYLyZrce6B/T3UbwKtVfMd3rO
hfCngY9J67tBUZX+zF0ZKVGg7uvzHObcsOnzXE/nTK0zwA9vED1xs/Hc7Fa4tWgFU5DEbya6IOSx
yzes0oaSr028eg0C2web3myym0iQGg0FUMJ/eAId3D9A3zz7VUTViQ9XkC/kXRNzSnJ7oPVQFWUb
6dt1g3BSgwBnaeDS40lc8gcbS3FeyoZSfKqz3+Oyk9hP+RNzZYrrcgWNOBqhWM9dsDGGm8ihFSJ7
6lgs47YqMNhGMunbJL1FDcLzd12TYpaalIPVFraERP8PX8DmMnTBE6gRZ2FpQL0jFpm6XAW/ZV5Y
nOcLXXYcbR1mSALWNYYg/TGtYOwX/a0M3Pgou0M1+9RVmFkYqLNVWv2OaDM+6t0ceV3p/qqRG0ko
da2vXFmIf/7BdNIxgsHjhvN7LIr7lltrLSu5X4jHb0+5el9gljEtXOtI82ekIh3RIFd12p6eHWzE
THRaJmNf2pCeDoN6jkLudOiU30CvjGdTDDJTT1r4anVF4PEnwoUcIFxCaPbdqvl3Bjdz/pqrVGBp
9oOsKOb/JMjBex5zKjWfniEateFUY+zRHXBeXovsAXzIU1Y98HF8NIlk7wG+GAkrwG0Rwf6Kf6Mw
US7z78MFZqfwEMxsscH2McxOFKxiy2T97w5RKet3ztGM0KmK+6vckwhuZBhM4AxAvJrmBGNZZD3f
a43KtidlO/dDBuFD9EfnKm0G4hc4+VPi8+H8nwfS/p/vScE6kUVvpz4cPhbXOMc2oYfiKix6X7P9
PZoYswGUSkyARl2iSQU4PV+rmpFbkXM8nyTuyluCej4v6c6ilCsIpEjAxsazov4iwRgJsHpvVNta
TMTdiULuyVnmsQNI+YA1QE+6S/TQOsjfZFk946zGaOeHi0ypxsl33HFfnE6Lfrr+DqBwVd4mVLcz
afK2WkhyYVtFUkNJqb2a+K+nJ/5rzUc8DRh2luSKkfY+5i48EtUbzEufbLdGpPdfPRZ/bWoA2OkR
y2binpO9z8GUDW58AOXemCgFLwNvd/hvziUOQE3JMHzJ6x2qcpFNioeuZQs54WlpZ2LP7Y5EgiGR
MWweqSe4d+NFpL8nw+MjozM3cNceVgyLTZTXVdfmoPAjU3tXf/+Nl+6X1jfq8ysSSNTycu3RodDZ
j714G6+6vti04/zM6YV2j8x9clOzkFVoYP6wgaR09ZPi6e4AqNXq3xjtG+/HsBktkmFJFi9C4sEY
iZid+n/KdsUpjbAChTKEU8P3Pl697d/gn7rmPH9H68qFGgvdoYMWqxu7FHy6dYitfQYEFwGnzvXU
FGnuSrl6+JROcLpsCCSRhSqqN3e1wpAX/klQLBUncnDp/n8WFLv4vBdP1vwK44+ROdN4AtDaCSYy
iISfn93+JcXqghw5rvFH2JTaoVgXPbe4ZdLG75pY0xIOwm9TZ9dHGYqsZqxF4NfdIwU61BLWu2zF
9omaz4ohRgNb8wZ4+hbSaJLsrXJ5s7D8o9mMH0/XMiRwry4/2LR7PW5FtxyRydqn/1A1iGwqFgNF
XZ7tLJOcE4lk+nxjjaOwxB3Cyrd4QflSC5CgeuWLWsiTJIwzOk5pOeX75v/SwKnEYviJpOy8F7eY
zwvpoWOU5KvK92tOl+hnlInAAPFfwNpAQxB1zuR2ZhET9IQZiGtzhGewImIPT0n/zmqc+hxASEJb
ALgTELu6SmhGGOauBDy/mhWndgk6i9AuHJ6J4yzfzVyKQp04deAXlIBMGSW9qvYZyE1Rg+H54Ina
aDSJYXopKYipNbOstfS14vk2m4FLGl/49HegP2qk3sKlPj/OUsLWzgRd+txYBX9P4hKkD8Lt58Wc
VN9nhwuP9Bl6axPXr2nFsRT7fMn+7jiqDEKFWBC3fpO1H6hgk4v4QxzhTNzTRAsJxqtEC/q5s/zx
QBSEiDAD0CJX1Ab3zXOz2qgRWk+Mn9s59VbG9GTfrj/4cep0d4bJW/QDoy1Fz5GjiYf32scotn8B
8H0UZfrbQ8rJwJ7JJ4hVXPvIzcid6NXOUWunTw2aH/BQbTxp3hUcP/eNNO+AHSya7AmzdyM0nL8N
kSagxHG0vyoysvRhZhfsaIfZ9bNDKbpKrRVPt3XLdY52nVO3VboPxH8qDAW6bNgOwoUCw0iZKLnI
Wlo7o84enO5sRwUylysH5guC25ekGB5dAmj3BY+TrdIQuy6F8EWHVfoPhHc7izHNw2pQLGmM3VNk
kHziXeYxDXkc9iTIazEPHra6Xsy7pgfjZl4OmyRI2f5YgXXBA6YF7XgvaZO82YfFbqFBHp1T20Rc
eF+bXQkZd60ih81OVGyyjoA7b4KL0WeirAhnrnK4/vlxqrS3E05ftnMe1Yyl/goBa/xp3uPDQtow
9JVWX1TdLc4zDmc7Emv38vZThDHLaqlC1l8zOYI7Bo77d4fGCvxo7kbWvvI4A1WXz6POa+JjNfp2
XdmQmUaIYKMcfgssaX8IdttnUGawBqhOl/je7E9Yd/YYOchmYQtVp+wIHIA0UU1BIC44nClPI4wt
Th6VZhS2icDTZSYnSK5JpVs+2vuwbUHBTCaNZq5OH3oNiPPJnXbvTWS3ogN+bcN1vGCfA1hhGwsL
JgLHZJzzvmxoAzkiD0rc3VQZUjg9DjQQ9O2En37yisJFS4bIvnZzjwgy4r9gZg+XlhCAlyWbDjuy
ydTc6HsKbmcQlYPN/BQYSnC9Q3COJzMhqpW4Rb4eq0LHTKcUJ3YcSi4HXSMg2aF6zMGpHAqjMJWm
igtoYNZTsqOBkn/zGKG7rQwi83fJEJC/roCLrkuBsiC0IL3i8KXOxnKtVvSopach0ZqpanzBj+N6
ApCEWnh1qUHph6SRwM4pE6p+HDxqn7CX4d4DwR2eU+vd+5RmiXlFnLV6oR3hGxr1MADNuRZscCNe
4IaMVLKQf0RSUh6HQfXU4TWPFW3oaJAvjkxGvKPmVBBPM+10fh8AZpnnKN/aZdBkWjG2TbyQh6LK
n6TcZ7I0/QMewfSC+xO0qoCYxsTnjLU5H412uYsKeUaUdSnN/EO2/LB9hGAWBvwXavJSaVMyTkS/
3BG/a/ntETF/saKENh3671bc7P28+569HFvIiJT06WqJ9cLI/GpfHUOksdi+RZhQYX5gfqoNuf0q
BqOzWuJanLHXLuiAJSrCbhF+aD3OXvozFkJR8amRNo6SeA6l0SoUfhdkKJ+HsdK2OXa3QWN+i1NN
0b3uf+XkQnhX7yxCx3mHLU5ZK3HXUi4qKAiS7iiaagCq6ic8Yd4IfjmjJzkFfOWSzmf+JGoluyKW
+4tMv7Mq1Cw0xjNQ7iBfUSkxEOXtqbPHj45x38GgDj0MPDb5Mqzg7Za9mEpBz3Lvrc3fw2QiPT/F
ujZwLplN/XHD+wBK7ZA/ZBFEZqsOwRZOUD5EeDO/E+vaRI48m4kLEHahGKtoNdDj3bbOHALThanr
I1w89o0478YZMuO8VaW0fTzw4haQYlu5IXLJXciEUoTKlii/6EUG2g480zCIDkHejYEv4vT73iIM
pMuTMkVtCIp/v528H70K/DjCVpoTeDoHLUE6KD8dYCbOs9pnEQfPKmWdxrZQTqG00Q2TXqXa63zF
M7pKZ8r6eZ76pxJ0gpUoA/MBc0JzVhLf0uCnIiUEABbw/MNs93cL3SVMOGc695yOAKoWo8OsCgB2
/Jk+GyisV1FG/O6nqLYZ6YcBqzwqAJO0Hw/yV6luySngkjr8KaKPYSN3WEOVk+cP2OBjBlZ2Fajs
wz2vj2cl0A1XvBSHkvH8O4Jf28yhWaGyH6+r/6THYGeuzsiYJIYJtmc3w2/kaBLXD/0iA2jPjNdY
pNvr9LqKPX7331TJTu8KPeNLDke2oVG9l7DqWJWA0DNAgelBAzUUqTLOzYDEYVmGqJKJ1bCncpV9
3o/Fsu4jsLGuD4LbuZJ8bqliQQ/LrC9Dtfy0MMA1pwO/xuHRWVCDekw1SmjlAVIgfQEKKD6x+GlN
oE/bu4sn/tyRhjzSpngENZ51+dsj8x4Pw2WqoU2P9+3ll2heAIG4r+aqVMN0OupulBalrEtsiEp/
PYx/k5sQqp27L7PCcDI4SEeC3AWTj4zwAbd4U3PHylrD4mxIBVWZ5dZWocjD9aiXIKpAHcSFCPK9
J25XSM1HCuGeA56YImuymMambU3R3gMCUZnTl2jH0gx9mR9G245hEoeFrCwO3YRTP9dM56pMJ28H
I6lcesA0+GlEm12aVYBpjU5sXLWAM+QGqM63TeRKlaeFmskChtSoiagLmduAnEJtgMOWxcHLBwVi
U4GHzcffh143TzkUlWZ8zK4CxzeeOlAMXzgrQ9MyYQVZrlKtBVddNUlZzCyENR/cDitsUkRQuo7B
HV59cKAmbbM2cddwdPHTFZalHCj2D0bbm/xdrF3+YOfMHGcBb7Ob7OFblnyLvsZDOqY+TKKBsZ2y
fsrOugSaWjZmM2GZcRiSbagK6omE/+eUPInomNsDZ867ButnFmncpxBhS7kGZtF6QHW5kFDA7IiB
CGbC2qo2TksuK5MNHW+VQasfsmrk3YMx6VkU5gKvkY6gPY9Vv7gBRtcjTRqRrJ8KU+LkbNUN5USY
t1NJIuov9A3+PHDpZKr7GkvT7bnWf83OIxDI91lTe4OkXtPppTlzbfCLOBIPLl7l5wWv/dJ7NRC+
mGtgoqCt4JYWU0lEsLnn7SM5nx9aJa8wh4YNz5c5DnIiD6Ys8UKPP5rTFisbUdnc3DKVuToBrJG5
THzb6mLjsZoZjr7kSo10n3oWh85lEzkttGF8Ngm9j0JXymOEoJQFfSJrKFZ5BxKG1Q0DcfljdAGu
j9T3t5FoIivkHzdNcAgJWda/C0+clQYLBpxC7Jza9H9svWwLt48/f47A4tNztxClxO7P1rA+SNox
CPDamRpIdTxjlmpkHGbOfSfxBO3oRKDv8YcPVrmOynMFihGrly9hjAQCvetH1WnFHTF3HR5o+jhA
S0pkYgj5ZAP7sj8wivl8AUzB/cFHh54ce24D6NJGVxfPUmP4pMypathQApIsMdcVnjMTXsP0K0da
cLidZ/ehTFIwSgtrwNuYCD6NrwvOn+/L2saRacRgSV79UeNpcfDiJRswWSjU42NMcNHkIa91QChr
ryrKdE9gETENWMy4d4WhhPBeb8re5kda77YsOt1/t7YYM8srOuloBTzmmr2bXHx3yX8bMlZTQv15
WGHglkDNM0OJc6IQMwEBv4+n7Jz53HeE19TK84rv88J8NKECLQ6QE63PxB+HNX68xTxAqNZ6SsId
CrJPXxq4czrO5FYBb7s3AiPc+dyToelVS5rLdVzWAFe6jpopcVC5nJyKCFX2/1wtL/DG29gPcJ1i
p0BaK4nvH9aW1ycnpj4NHQWo0Nj1ECWx1aVTcBNLBpQJUcXoC92WlPSOB8pQVW1bmI+gakoo2H6c
Paj+9Em46UvuypgORwxqx5N0HrKdb1gDhVDg//bL6ys1qvgTdUNvPj7U6QZ/y3dVXesQ79UvX9Hm
XAZcyf1R2c48RpQFf3xEItqDx5nwUwijBpFp2MYlTKol/QZHYQhEgBQd9v2WszhaKABO0IgqvDOL
vhHK6mLCcV/Rbwk1v811W14iPAlB/1oC/LqQq0NwVE4EUQwtn9F7bcsyZ3ecga8l1wXqfIiMAheL
BuELhkZ9CnJg5lzOAxN1uzxAzIdZw7hr+EQM9mqaAx/r/O9negfW4zKAJzeqEsFE1Dg1RGN0Lz/9
YUbFYxjRUq9LfkkftHjQR4bWx9On6c7A+u+drc7dRMxZAeI54H/IfZNyeDByHgrCGhK7zhMIdhtQ
RFYgtHSxGeLR+AWl4EbMlPKBX0Eu8zu854VsvABdwMQYX3oYdnD30UnaW//J6hrda6A9L4Js2XB+
G3hyQsqs+7pelwcVGlHGX/tVebEAYhUskeCXPMRvJDgRRGbqf28V1jsuFw4rnHjKry7pFWjDZ7/u
nN08HfigufyWXw1iJbPmGjhkGfnmC0gRR0aiPWsP3ZZPHQRk78FrKpBGKdZG8/YmnfYHpt07VJkM
UoI58Sjns6fU4VCvXsCqmOYmnyoX4RuCHg08XWNHXqqL7PCkFxu8kWTYi6WkRH6gOW20UnMch6tW
+JIu8jsAzZx3PIPc92Vnvg5ifAkj9vqKuhQNWd1Sw/Nh/IMdJjOioC7MwvtG3G13pcKTzTsTPQ7T
cTHPN8scqI8Y1TQInJ6woVXyc/Setryl/PQWmFT4CvIlyHTmC2I8FUJQw7GV9sxzP1bTtR4bR8fR
tV6LQHc9thVBCnQ3GLLk7O3u8dQH3FI/ZbynSr0PFjMVdwlLSjIfaRlknlAk6MKx0Ats0rQODrCi
aCc/dzH5HQ0O/wUOsb/i2/r2AaHDU5CsfLE3hs0q4UxZZah11qQYznIQqSiGoT0DzJSx7jIh0JeG
jg227VTJV2rL9X+ZVgP/SbYPy2fyRm95tL6LugPXhw8ToWOwSWBdv0oc7XcuU6U4xrVdXUVuYvW0
1jzgHiOPwj35MvJgWBLCfQbOE4tKzSxiEExT74u0v98U5jxfW+PUwHH/Kn/iU2JptFSAHViMnZ77
+GPpEh8icPGNFojppfKeVR5XE36/5G7dLZQAXRh+EUHagkuyi1kU5nJFE8HpDuXPbstVy77U01eh
72l4XDQ9OiM+eXLCEW/Qy3qIM3kJ8d9VsgOVWQPMU4Zg408e6bLU9EKl+7EPPCqZZWWpYoZ5I9E3
CDKCIf4uryz/0bGHk/uiA+DJawpGPf6pxn9U+pto+JdtMQAdWbpL5vydNB2Nzkm8R/ZatTqTE6/6
91pK1H5CkneaIbAaC5q20VFazg3VR+wQ/6RBfW26qUqOrTfHHz/uhY9eMY7DK8po2kwGJN6yfAid
9v3QkAqtZK5X8zHhQU/twdCUjIFw1x7frSKaV+f849N0XPLMSezhDO9sklBicd/b/totON2oQsqA
EuFYOWEVlNOopkVJCFTnvY07jfVJhTDiGsVn9zniNpR9d/2RHr2Y6qqafrVSOHOVXUh+fEDJobPh
bjd9zA9iQTNKvHAvUFNR4O9yxnKcU+8uhabh5eMQ5aPs8pEsflMDKCsJzFmvIWdPsexZrHT3+qZ4
QFoInXOvobnv465i8giVY3tlra5B8m3i6a66eO+6rTY72zk2HqHaJpozpjVAi3EByNMQxarlh/R1
irKeTSdvk8t7JkT/+OyHfoH99fwhMM759vKuMGlgkOrwK7VHuTGAMsPjoTnyYcqRY7nsjg5cKlrs
JrCPhIej4SnOkz5VMbwig6DhEJO1Y8wc5ExD6vJvLO5rKCC18WdGSxUYGKIflqnOccYFn/MoT+fH
o5w7pYq4z8vq1kZDVSCntkyQe4RHuq2kNauN5LZe1EFvo5lxW4vkIaY7JmndWhhjyLVmAdII6tet
K5z0pz/TpjZHrHRfY5rCJYPyW0w/h0k3EM3FmW85Oad0yHtbeoHVT+uyiAeqCAev7oJHCsS8lNLy
9g+N3GxK9HJy/1++7FsGYaxp9Tn1BR+lQkQ3izEEZrewWcLS1luuj1eEOhyXYFRrViE48gXUOPe8
dfJkyVR+58Rswg1Gc1YoEM2GwMENx/vtwZjYJWeGTKFcGjdqgTgZMoYxxJ6h13kpe14nS3ToTT73
7FJQCtha1s2bMVB0L/Hit/zDeoUD6y72pBRrw/ATM8ONWCaeLxLG2xDzxGe5mvV2DiyqGtWwmPpb
12cEdVTLD+PBVWxT4WjJrytR9rK4IFpEmt+s7xI9NMmdlakKzq9A+pxFI3YCnZCuF5ZZOX+XffT/
3QatkB6vsf/WcRrran0wabE7ylnQFeHuTYJwNuXuLEA3FO6vYMfhO7T4fU+SZviAiLLKdV/fF93X
oxge91pzW6UE/LWc7RsnR0g66iCujJ2AmjEme/QitIOkRPoOsZo9ZzRZkUTAq7iUhyMpKdbmKsWk
br3z/afhROgDLFp+XWWZNHgUCgYmiKT49rKjS2m1xlC/TWjqt4KrZ22k4RXIi3uso9rBBy3WsevY
yHobsDTki+4eX7EAyZPMBPCZblfC/gzaaFG+xPStirU9Gie5Pjonvke+5G5GUMsoG4Hq5I6JCC22
dkR9SzEH2w8u3VX1hWYEee3xotjHKuTRktybl/eL1Go5PaukPqlE9pNHYQ9sVh8Jrfu9Z9/HhEGX
uixLWdhQvL51dC7y4KSvFPpY6dzX5vuvEYMIJRXXanJNyV7iJqcshJX+yCWk46v6/FWJoruD2Yj0
W60bmyj5OhhmzgDat8qe9qjYSOTDvPoJCHzGLUgNt77+P2JwbqE8jPNZGg9CKy3do4JhOwNAwpop
WNq+llHEDshySm5irYnXKn8D7d5fUA6Bj0BsILbnDuFN49715RnuU1SQyuh1w4JVz+aJ6FhxCA6W
WlL3FiFa2ZFuV9Iu+j4nUyYVBICHpQGevqmuSuth0xprdGcF1Vo1pGzIiQFPc0a5FVSEBchEs1Bp
Er6iTWDAqMXWXXOscrmF0mvWgbsHdjLZRjWv/FD6VuVbtzHWpAFoj1vAI8DwsjARMyhicCOka0HA
i1bZMn/3r9Vf2SrkrMuoXjO+QcRd3sXdLXa4YppQGrRKmhOscgVjUiUdsNStMTAS79kP76WEq9SG
xlscnleFN/hvcqtBoJdCUFpAje6/8ME0nuHQXYIH4Wmt6vMvSYSJJpvfM1qStRFD723soMIUKqDE
E1nI7YjbNJUAc3Wlb8nVoqMZan7yml3SbXaVmHcOqr9b1yiDI9Pd57CbO+LBWzJa9L62wwqksL2N
N9P0gnY0XXp9FNGw7siS/hvv1jJY1VCv0T0+VzMLlD/bXnbco3E01nI9oaAuIjiu1HWx5xUyX5ol
YmAETEfekBhyk4mIecoTXgSaSuPE5wDd8Z8EG5H+fYCniddGp2QkMPwJfm4JEvzwuPycVWs6su89
hyBxFOSReQy9roVBh+coe1boWUv2WIJu69Xfebup/lz77HjSDLWv1X5Jy9cDaBKJD5HXiOmlVCvY
oxGcyJROO4qxMOy+oS7Q7QX/CT0BC5dwJ5San/Gw0NHprJWyiB/4a8GnSJJQ/yGK8ZBxif2nvPKY
JNrjK4aPx465RuhZk/5WaxOnZ/nwkLGApSWzQtUKYFAB3WIE1trIrDSufsB+pQgWGIcdBvsKBWK0
dgeODk5miQwu5c+9aS1oyweN74TIwlBrxch5y87JocK/e+4ZdvcLarXqyAL8IcxV0iJLpL51GJwI
rBIa48FZPWu3BOpUarE77TY11Rf9OlpYXPnmCKn//zQULeRs6FAk9CLy2agsC3PJIbn7HG1YswNl
jolF2eeGs+kHTTlsax+518hjzY7RXQt+0IHs0qEiRKFVWy1PX4wkdF6cOMDCOApXqy0ZfUotC8va
1eTG60fpnmqWxwVI8EsY0SLUbUgawc0IVl72uLax0WpfyhWt30FuloCxLzM4sLYViTsGEfDNTYha
+Gu0BTv4gnE3RSjMtYdsSkSWn2935OO5twuLOmSrzkv1mLWcSo6gms28MSie+NU2o+yFRpnwD7GB
N1CqYIAh/6aTPXY3g/8gW3E/wqh3Kf3EGUiaZu1jz71ljZWtrS2D7Y2jvtu4HW3uxpRb+SsXQ5c9
Z3axT5ji1DU9BeN50VVOd4Gh++ge3ZlUfp9wOm0R8yzx4B/Xh7tFIuepvTu784xT9ojteX8Dc1oK
fsfF0UucwuZRfT9DZPO1bWAA3GwSj9bQoJPaCYMqTyxbN7+g7ArNyCjbPaHxxzYja7J2cYF3EYAf
iTfAEOZsAZSfYZpF4XO/ZwZVeNPOD+EfpVMjK0/yYXqbw6z3bQyzeY7HUPB6+92uIC0pBGYdETfM
991IAvvZHxMY5q2pp3tSPDmxXxZYFBQocsFSgu9MyRyXA/VxUtByOU28gtQ8kIvduZVs11VqcMrp
4u4WYjCm06bhrmxPmoySGkdTgcHgcGOn5IqP8A5Mfo5VJFotCFa4NOIOi3U0gO5qPfLK1IlCdxct
9+Xi693kINfXAEkUQ3KhzCKa88QXMxMsAyLvWawpHvUY+zP/adWGkBOdTdnmkTCpt5vewGzCDlzt
yysc8nH7CRjIwisgLH7fix7rh/UEhkdSLlBZ14+Qu6NFpntf9tfZm4lFqUpE+ROybje7b23qiaGV
nHOsCgP9B94M+ngn16lDAZPUZGMrZokZ0iWceImiEj2zWl8y9bRzVeu8Rg4YVmvOOpybV0QYS2oM
nPZvM4YdQC5v1DQusNy1Liba9mH/3LVAKn2ztxC++f6ZpdHznXIZZK6K3jNB032JOTIRlyEE6Hxl
ysA/gd3lrutZaG2yLVIOR6DjAyB8mp8fPMsNg+B9ckS222GjayJsGYza6hRVbKPd0OEBx0UhyYZO
vRyKRW3tisecSj2CZ/PaTk1QPP226ADFUwiLntG0u/m4hXb0mXDWJ/TMg9ot3CXhX5jMTZLVu5jD
gUfU01DCFXBe65Lc3bFiozzs8ZMC8Pn1D6DnEv/HJ2+ou4jqP4MH3cYvi7Fb5RgQw99+XdxgIIvS
E/YC7/GYvzm90ZG/qji0kPMfEr3dq5IkIW7jyXnGIabX8WDsP0e/BxG5GH7RhGKm7MhpdGV3NBPG
OfzpU57FxA2bdihnPRo1w3f8OnQ0ff4o3Gj/fOWPWL6RjH8Do7dhP6nn4n7hcqIYq2j8j0ZoPLNi
GA6tT0p4POIqdtp5nqdp0DGhJows/jr90p7tslbM0lqzdaNAGihqTPl7bscoiuBmxZDbsiWj42Vh
kjcR7vKjw1TyfDMNikrf0Or+SnqNexYg252gRhvjHsIRa9/Kqhe1oYWLiChbb7b81I7E0GAiHlaB
Aw0M6RRjeuDZOr+1D9SALJwcG2QJZVZWyfqHrllNHyAYLrAxU2vQYG3AMqifvTDFx419Wk1o6arH
utOrwmLC6mM/OvyvkPnBdvEJI2K6SQLL0TdPinIgoOnpnlydN4N3479G6/mJMgrQT0Ew1Q2+15KO
fIIkaaMFlrsf6vzEOYDcVOQ6uSz+YbnH6Wn5xoAjKkk6iihBIsLWoTD7kWo6AV/LAodQNTwlD+aM
fUJh6zME0KxP6Sx5DlyC0OZqZ8oT0dwyY7guea446yh5zuAMWRt0vu/W6G/wHczxW6telZKJXva0
njwLydZJ/m8sSel5iBL9s6in55UqV+5UjGpfPiRJ3tzQhYmrwNXJ0LfBwzbwys9rHFaEvIiVitgn
yqhyoh83bu8WgRyYlEdfPJ9IRw2l1jp5UoSiFQq9WuctEJbvOektZLAoKY+kbTlA3XsmRSVNCtep
oRmsDe24WVFD8TxFROoNb3iCJ7pXw626Rpj11HXKvw3eniPDHITn2fWc4S06y2Ha4+3vj7P/1fHc
bKunPMCEWCuDSyljaq3VnyCUFMg2JjAmh+jS2tdlSg9F+W8aSrLOCPVg6x66nTtP9bljurwqymQF
EqWuhKkhIUEzlGg6kMBuLb/tKKa70WBNG/phYbnDCOp7LTDkYtFdQhzpIAhrNrhBS4nnF8FxkR+c
ohSJe8OMjCOSJxL3h1Sd+t3iCqN7NoviFYgqjiqt8jy8WSGA3BAghwJicyLy1S+/aDL5HJV8PLU7
6NhRopcuyE5UCjXQW54zN2sJ6Eqe1BhQ4h5rg/pDZYkybQf3pVBb63HV4JKyp5RiLAADkwV2YPGw
UUWfFZS2TXBfhS5oEHSlrWDcEvqtLXsp4kgbX7OAL71tYNiCXvy2YQdbDkcFnyvsKxRyM/WWKddp
eT/5kjl7vELaNBfzC22JYC/n5Quhci2/Qa4+XgwMicR1ywSamjpdFp8DrTmb08ifPcawirQc83vb
BaV5bKMvmUgRHlRDpDbDi3m149gTxSqRUL3uq17p+YDTg/PTr2iBXWybE0Xd4Wrn7EwPfKTRTd0e
GhBgGbfTzMAVpluYmSK3gen34sPYu14ucu93x8HV3DmElagqSIvv+jIVvDF0wvU4SZ9pQEZsMdH1
KWljk+6Oz/6Va7NZQvz+OdZ5yWSO5dRgL9Y+uE7OSYvtFRttswwtbTBwMZcZl9nHmqmFVeNiOT5C
XdfL1pbaRkqbAreoqdnlgMky9KXlctym+p+HIqOts/WpLA3vF2LSvZ9H48XPwc/qoo3VSauW8Leb
nqlMX3nyRiL4ZBeVzWPhzmv/Sjw4iZJG79xKXoz0OOobPlot3xctgmpiNIu0VnsYfnQOkQiYdf3M
opM5h27xadhrDJNQ9qyhbpkhHxE+MTpwUdP0i++QfJLzXMUUs7H9Yl1rY68VcsrygOqiUQI8s545
eSw7G/tfGfKRXqlRsne/5P5XYSh93WKP0QDMKxbA7t8gjNgx8wP/HFuRwBFA+vZQIWlbq7U6NfG5
OZjtGqSi9LgE2tbLXRZZouMwIoL32YRoJvyf2mXd9MDPdNHD4pN/1m4G1icaxbrWH3qwboEA8NgT
t9ZpQOZLL/lCyHZuosZIQeJnXEv+1k63dvXLiDddsa1gJX5tVRgH/qJ+W7MT+YbXhpnl1HpdIyYO
+r43Faq8euyW+TNRxliehTDnN4724MqQA4SmlVmBl6m5L1ZHx4dz4t7FgyekWaeGUeqCSc2flbka
4pi1+4WOU6/lzqyb02sC59k7IsPG1W1cdPrZOCHYKVF1KMYSWjDRwTDh7mZXdp8WTal5P68TMTR6
nPl8NaXhnVHh7qu64zQJbNs2NgvK/znmBkOCPR/XbGwPLZZzbpoQlsoD/aS6wPFdwQOI/VumEiAX
LHz27N0a8JR9eTzrUrw9QLhFG36IK8NV6PmV9kDP+Zxkoy6yN4hHB8pk8bQvdLaVxLr26mnqoKJb
ev5yp0VT9/LsNJGu57V5l+mgkh+PbpD510OoVS2bs4tvoxapovQABzMthigX8hGOmnqJnHwY3Rri
C9qQGRAFbFKr4GPBIr7+43C9u3IitpbKbba0ViEE6x+/J2tu61hY9DR/3nwdqJcYgf6Kz0L/yf5y
pkBV7U1Uyam1KW0lZ8vU6E/wLM7qpd8DWOXldemOPo98eKxOkWqsYrXxWqZecMpAbwumwkwVCIYt
Hps9KjVUBQqujr969/FE9XflOvEoxszw0aQGgtuqqJALcAxZcp4kZnTqO00Iu+rndmlUb5lUxyys
TO0BMnsmLQzomDWw2l8vKA8bYDcqbP2csH1fgozr6aBlLh/KRVjj5+WmG6Vl1NHejTkJSF+NalC9
9EBn3sw1oTJftyuU5PueDxSN7us56OmV+aRqY6GDKibtuChHwetTTh8it3sr5JciBaSbt2s4n8Pl
7P/inKa2WblATT/Lt0xnHiMbZqtPBaPqA5Td7Y7FG1bxAwxqbE3jDHCtct55KD0Zust231ISayzy
Kra2Ttm0Lkk7Fe6B6hKU6gNldMQrPTB36OeNHGsaaDGc7YdGupSLepLW5V/tDWG66B6vaUAt0HLf
TydS4TvxZOjrktE4WQdJHB5rSQvRH6SgY++8qukvef76/TZmCM6umzMGzX4ixjmnHidTyBCmiCsW
U2hTsJKjURnej3NjMEXgfAIZg4mzPkU6y7bwLMMBlOO48yawu8vldeBunqwgeAQ+wPRDIRjnlHyc
WA3BFBLwaVGdzvwhJcghyxvtWgVs7XghO0D6NbqzT4tw5e1qq64SPkfNg2OqJB3C2wEb9hEdaKYV
1CEp2t9mh66AliT7VMfDkIZHs/NyGHxuvVP7qlATIOFRetskOxdW54mDZvzBP8w04W2t9whcpNNn
zsYxnDl+stuEirAowRg47XyUAFqdKURbT6lHISX4H1j6KXV8+KfgPK50WnvstKa0B43Uu7srQ+c4
iekojkp/e7gmOBfkClUTv8NfTMf9JfSsSXDMhylOR0NFJar8acYYw8htg9Gx5YL6cTAN+8nljq3Z
d8IYSI3vmrptXMomn8X0fNA7woHPe0AfhqO24HC3UAkNunrkmqlYXmfCgG/Bv3nIs6o/JkQQoTSn
vOE+jmvwS9eBtEEKMtkbfio7QCokPAbSKAc3O/nNQhAIJFgM3caaI+M7m/FFLoJBTECh5ofdDzDa
Ldcb1mVejBJXQvVuv3FpYiaXox7dzy1PR263FuWRXSdpDf0Oh6KZehrj+KFQGfKjfYzdm3+GFU8Z
02p3IcNGM3A/1nTTwMWAPVJQvyBxhfqnJQEAfN1LllDUTWwSAf0gfJ5eb4FQaCQaAIjtiHy48bu2
AAqQqzcGfUV+6CWxJNnR7fMEpsYcnY4Ej78jKuZK27s4f7DvxcIuzMVapo40XcsjlggbzX3SJtbP
h6gsAgbiQfmOSYTayP82NQuxhIzbdHG63XLDka/q39EGRtOxmZFbXb6VD8f7dvme/uYW9CWDwc0x
IMMg4Bwutpqu8KaIun0/HROV0b7Aj0B5E3EstqHRWJa6Zu4X/Y/mCee0G1EBjGuJxfA6jn6WBNXe
PT4wixzQcjLigd91a2x4wII+KWfjRBQquobf1XI7KnGq7GVVDz7gL1JMgTZlbUwVCX5b4xz8hq1F
BxYZ6hERusgm9T4IITZiaKu9tIu7hlHtR8D/4NAp3J22yNoewmTE8HFzpkjO/dtMm2XdfWMywSbt
EVL3Lh7DD2sUJVLOQhdrh2pcyeQGWFbbdbTPX4o6n+V96vkvYs1lZtAnOmwp6Xn3YlNfF+B/wOGi
W0Hcui0tCFu27NTCLCZfPm2ucDGl8rfU4tCGaTdgeM2rjpK6G9VOOPFCMTNjx/BklTY2rmlSUuQk
Wlsjv1ethWmViheJW8kRrSFAUSFxGNPihKL2MmbvsfyZorTLe6bn6aGK+l2beaW3zk+ejZS/G3mI
mH9Cx8GrlebiszPF5BR1nyjdGAOkIvMVhZpO8HClHrRuNNdLBn7ijWmGCcsLytw4z/rYjCpvTsoD
nUSnfAUH3QivQlKV/Z3GSpeorjsgfxyB2cswXswNBOO6HBDOR8Yai6J0ObH5D7LgyGzrw1tTdDRy
T8iyqHuV4mPhvOzKcTuhIiUMtgFZkzynfd1fizwFWb5qIaRLD5ptRp1FoKn0HxA8w1BC/uqHcWuq
SjUHfcXBM8JJF2Rc4ec2ABBt61pwpYepYmWPkEU/AzGJng65nf/vMk9+b0b69srGWYOQSfWQaPFd
J3eDr6nZXLuGUkmS1enH8Qk8QJZ142zKCnuZLUq9dMwvevHfFBEOYayIe+yQN0nj70Pi9IQk8IkL
xvEfs1tFaPvq4Cuzm5XL0lbnnVr5EocI9f0jLGNwmllx9ZbbPBPqXjXxiUuNRD8U4SH1BRClx4pA
Lq31XZRHXisuGdQqwGWu1wKVvMTzEqtljZfTPPusJKJy/8G6pIcVtUuxZ9X7meJcENiX/wLgVQYi
NNSgKXLvgG8a8xS968yozgvDidfGwHQE4QySVd1k2HUhOuT/ER/GLu8z4SynYPgVNWjJhYIr7dxp
EbyWd5PF25ZlrBU09ZKGM/6PG7PDei2U0mFO6m6r4sdwrdsrqTZtdNr43YTEsZTVrF4dCufGwG4a
cLz7nS/mwz4PJyTJtNvO58xH2BL852VJrg/yDooi3AAEymEpUwW5HFsyeIqwkyDqylUuAqaBzF9w
+NbPlqdKyndGKMEy9dNmKYtcJ1ICObWIHfblC6YCEs/+THaDQtauL+fHL95EnPh1XSXXosKFOfo8
TvMRePoE07i6cpUEOD/sl45cUpDiZMf3y4CI4glZ+QGaAhOhoNsHhnjoSRI302mIGSTLoNZpkVwl
upN5pOsjR1eDLXGSUfJhGpnOylDDS6JkDlH0kgA1OMLSq14c2yWVGRq7NRVxWi//f1CqNlhKBLzv
78V7g9B5v2Nt0fyKQn2xwosLQ8Ez2hotncMY87n59sqSEQDL7mTi+IlZH3hbx9+c6bHcxmODsag+
xvkyW+W16SMgaftnqhLNeQKy9gURRN/efR8yvowoT/7Y8NUxnJiEOutIRS/nnlF9PCvyLWGB7Ti1
rWuriu+s1H9/s0FXhM0jGtHF7/mric6s9sI5JU+Nox6UndSlTmE3n09IlXTdxV9Ngf2J4MKeql0O
WDl4Jw3p7rlu1wVM6MPniH5K0pTRIB9FFyLK4GIVHqyCN/RqtVzwPTQ4zb7FxlfkF7JZ8vsDzgxH
EAceF8bcVI56LJRLX3DfYN43Dacd2mirqij+FMvPGhXNYrZ87i18XUjNgB0auVNrmOlmng9iEKZC
0BA/bI8X83UndgfofLp0pF2/YSfkiavyfHhytwiz79toxB4L648tOHbh/Z7yh4YMAAOrYO83uBKE
337k5CJi4yHNP6rVBPrzF8agI4bw62oDp6O5ALkOy3kh65djzlh2jqOySiimuyFrVyLtj5cA3/aS
09pi8xkobunxWmllYGxRQsXy29UcQ6Harn7QJIgus8QlTkyikcCAH9Uz6YGAwDRQdtrDT7LfmYhL
G6yce5Rrz+HHwWQuCqvN+TLNDLGn4KRyhD2h/dkPyPr5XQU+eEPfuSzIqqXlpcvdzyPSJD3Gk7MD
1/ARpFIUWoRn5svAnkhH66nse7b2LUmB4pC2F3kBZUw2eVbneRRxE06ecA8VmFPIWUnYHx61iYZp
fVHSPpVzClTPjNGlifOhR+QxxoLjNp/Lu2XbVd8j8QCo7acWQewDYXYGhpyyM2Q6aq//Wq+gsJ3t
xBrBcv2Y1KVfDDujUo2MKNOCVIqkS9+XpJWhj8MWwU+HOLK2o/1Vv4G+NOXY/aehPcVw4gYkwu88
MwDgwqOu8SEYblgbMyRczpa8g7StzFMTo1mkHS9shxUA7eW9RWxamgHw/2Zra8b+gGtii5Zi74YW
XAUO8MtewDEGosmDVOGsh2Dd8ymLMNQuKZ8ZGRlkOFtHm5ccJ1VAqXLmDJRey1mo+9BmX3/Bet+m
tmD9UWbGUESrBGmU19oesRjeEuhrqgMaZvadde+8DgykKo0ukNTJDpA2QhfPBR8YEyikYlGm/UUE
emwzm8G+Wc2sEMpS8U9GjGlATZvpXDO0Hv/u8gUXtSMFRNrCvUq3bzfcCCWnhTr74cE+GqtVEtWH
RA8X6oajyO8rEgL/zGN1lT5A+0HChKDNgsDonorGFDpJ0wGAvQe7qbAF5Mm8qmWUPCwbLsH+AKqs
AuP2u6ibf0YmfQ8f3vdZhc3tVY0K//uH4xGfXGU/U7KI8ESCFFmK0rz7vglKk3YJ3ZoNb7tCC35V
/4qrkr+uWuLhIcW++w1gVDiLharyCnN1aauLPoTSX250VHVGBAfmwdjYML2TyAYSmFMXttdZC0AR
Hl6EtRfmIuX45iGxWBQ/ua9Gf8hTH+kOmQVhlnqqXMzQPpKCxFEUXyE1eSvknV0mK4Tj8hwxidac
0Cl5FQ4CZf6eukpmprCDmGNLRB8E5DDdCCuGMlmr4Ci/SSO+NPoBy72ovhtHT6kJuXShUb0hrITD
uY7ms+NQFhRegi9+FFjMAib+T5EGcYgVyq0zdJmlNUjVO39yzJnUQhXgWuv5OG4VVo7MxUcQx5s9
moq8/k3hIaWZ+cIF3J6Nf9ifje5RcTvmXSEf1fvk8pV+V3dQx//GfmAlB0y5jItf3UsDwO/3sxWL
e9hl3GrXaHfFRYm4k2wQ1P5lq1wj+KIMeAQQblhF5LTL+a2P9c9nAMYfQVzGyRw7GtXMek9MEZO9
RglFg2Y0DWdhOy0Q8ADodia82kDIyV6nT5UdoOFx6Jwk2JeNDzQT3JxKreYC4AvM1qRii7vEm8QJ
WxJLKmi8FpBSfOmvxfEC6ASTHFXQgpUj/pEtNM+z8eJkhOzUxFCRmR/nB1TlKHWzHCaxhIez378Y
69A1Lr7SLxAnI+1xWxDhv4Uyfn3LCFLQBOEggLHLSNHwWT6oZ0XSC1TIrQy1c30W1nYFyt57ed03
3fuory7umrxU3LQ2NIqLSbHQBOFg5DSpAbSLO1Z/x38Je48u6eWKt/MA9t5pc/C85dPqR3DAlf4B
d5jAriX8GjR31D3epcLd7rJ+niU85QjEz1q+wCO5+x3Tgab/YSpSYKT5RJux5c2YK5W9s/Zi+Fwp
R1aXXPCkwN9yTcQDYbrbjwSe3+sMwnXeXJ2Y3o8Za/tHf574d0HaMmjQMd959g2JVQHK9qNJUUME
JEnFZUIQ8cMFjOy2PPQjVAA23eWq6eTkutkTa0HMqJIXgIsMY+R3YYcmBzJ460h2FxHyXsuvfE4y
CXLEBBc7E+iQBAqFeO7Ly0n8Ro6Z4plYJmQYhxFQN2l9etYK1dpKfWIaGs7WQ0HldgyA7gPZGunn
zQHLXB+vCNvJo31c4lKDtNk//Qv69YTwGz9z1RBIfU7i2j/nIprOdnAEyn00wfM+V2VZ70dYz7e+
8pKlXG7GWY+LGIDNHpuQJVaSiMS6anjdK8nmssgBcszww7nVC2hOFnJhuZkpGlFsr2Jsw5BOnhTP
k7zP+RfIg6bFWC9y9iOfOD0dBstZgdEi+tF3Tn0Y0PKQXIKsXOVrINuSkpoimUajmRVjFDdOsX6P
Usb37U8q119axtpvyp0o6k3VuY80J5CY1HwxCDL7RSg7Oub1/p6MlFM+caP5urWMc1bEliAIatne
n3yE4CZG8OTNWEcG8wo892JESoA3II0TrSw4loargF8u7YfMTrcqNWSqUcw4W573SuGLjmu8sEPh
W3Lj7gsUuZfaDa4nN2opoq+Oj5s1U+NCDDRP4At9crDoL8jp4Edpt3909+CDgZmUeIVyUEXVq2Cy
Ha70l99iN1Kc1Fii4oquG/dxG0DPRsPx+92PAzKBTokGCdsUwjMBUPKoCaBixFMbD95RCzBJqf++
/avm+Lt8s9rUvGF0fdjS0uejsxJsHyEHSvElFYVLFzK+dfZqUaf5iayolYHC4RYvxZ5RQkwt+v5u
46xLNuACdRrQ4FARu8N76uxj10bluURMqPrXK0uDach8Qvhisv8yXdXK/XdNtfI2Z/2DR1xYzfKg
7oEAD4+5504lW+OumnkoAAJ0Zm+IiUdizlcQJuYP+48OUddUPoKpmUb45QV6ysaqP2cDhJTM6qVF
CmSfoPbtudxfiOX4tZFQcI4ZGF6Bo2UOWEqLx2Pz9yzKt1gLBUnxemJb3wvsrbdYjmb7W1Gc/3/K
WdtbEYYYxLpb5UI/kE9yi3D8TMyb4Y+hzgXs45hjBHQVd1aTBLBultyJAYubjDAqOtLYUxGDHIPI
qiUfnTafUY/Knu496/CXyZ+oJhNrAnVI1mr2LpOXq3ACXWVSL/a2xHvZUNqBaof6BZZ4A8cQa2+7
kHilmM3fEUamDRrB+wqTx0D1IS+988JKVFiN0qxc6nczVw1BMHRHsOxG1HfzdexkV1KbFEBoevZ4
kA2fh5hM2NDpGDFHXYsLi6V254+bNeaX8xPDXDEf3tkX00FoqXZBFAZBrmxuJygtq0fb51W1qmHU
P/t0y9l1o0HC5RUwZ0i/AGWfPFzAtgGntJB3ciDkZmriYnIOonzCX8yUUzFWfZLpp1aVsbM+Rkvk
BiHkAZKHET0fhtKP7mW8SMXD+83TXYAHhpGc4Mo0ELad/79W/NAKdgHw4KP0fkiubw3Ijetl4CpX
SCFYa7Ly03OmISNvT6Ud+uLpKQyUv8yavJzZ/eLYTQ1jc4Nm+i8MXoEeu6Z71nEYG/jAlZQy0XUL
W/wm0yzoK8RWTXM0NBCJsfUjviDIGJ1YMCOECyjYalaqBUJyA9bsgXFacIv8MNSV1NhQyYTAJRCL
hCIrL7XiWjgqjhXatApVutnxygzKUqvaoqWBU+hpE3Ki00TOAqzI/0p+0ZLFEqqj0z8U4ocXMkOi
WUXXztPgH9MXGuLWbXSMEt25a1T30UqODL1Ga9u2ScuIu+GA7uYZaXNuTLufZJMQ1dsBbT+Uo7kr
x0pBDhWvw9nYmVoJ/t6dkXOOXz0VahzAo1FI9MjEa/FVXoJ7/txqEAs7X4Ebwt8+nCXR0v30HBWa
I0k2Rh+9CinitH7FqNfuOEP5VhA8uaDLeUm4uXbrIER1BUOcVsiB2n9LWUZriGrePT6vJqANh7VW
BYYpvGNxzQ0Z3z6Vhoa3/IISTeAKG0YkjNa1ZUhcxixa4MuWB1CewhKiiPbkO2vCRn5uFXxFxeCh
IKMuV/SCjcot6QymgT2OhUrSY+NU+pcTnWgko5M3x4JuVTbh7vN3QCdN+aIZns7tOrza7jR/cI48
UW9UAh3ACbSks76L2rycrEZ/g9iwJDarAsABvaAc/1cgr0lN4VP90zmegwdsGuf4nqQrtlc1yJG9
ELoR/WprK66+KZETfof5s7/Fxy7a+RhwLIGMx/Sm1EM1ddT9YTVVZUPfV7cH0CNym6HDMm5F6/bF
URqw81iiedSRlB4TzBLTe6YbJS7Pn21mScXpn/C204R0sgSitg+2K/3EjQTEjbWZ+C8JYQwq7xEL
BbkeqFQl8RmfMYvZVo70coGJ9mSDLuEkWEavbgeVDXeZX3lggEyY/W7RhheiSpw0u3XXUVRN1fBW
j1ULJ61PYyG33OaltVK11u8OWtLNRVCCxY6ue5/1PakCqVqzz0qedklb4NvJIy4h7LXqxDE2xrsm
58OAIqrjy+Tayir+fNXH/q8E8AZf2f1HoNkP0TqKMkHt9KFG6QcFp7vbrbPZHbaz6aJRRDzfrxzZ
D/3bOa62/CCUlUPQq5kAS3Z427brWSHB/PIdOZILctiydsx0cmwxCppEarx7uIw01tPi0OwfKT4y
6lYiASx0j+n5GrMR0mXGsK595LQulat5xjYi8Sg1h6lRs9Bp6tLnLZZwiTd8mTaV1JHHfY/801tf
uw6UWfnoDuk7CpprFd/vL4cXv/Bq/Fo3EuPQUZSiiCFa7lhy6HXjs3AMAR7Axp44AeBMVWQzoIcj
24rgpU/k+wPRt0YtCWVjEFm1E4K6OZgGBDOzvE72A9TkZ27M7++10cXMVBKDnWvnDHuQCWhjDbQV
YBPP8R0EwkShUtQUhuIR3kMlDBrFpNYS5q/aYBKZZ9FQS2Dpl40R5yQfVJXX5k3YCv/dR57qGCni
eUjjZGHvfbp9rF3QPDfttTD2ZsULIyD7oM4sdUc3guus5smTz5iVg91D0QaIz438PvmIIPkpg2VK
0XD4v7hm+u3SbF/8ntAhNcZpEEw81Zzq0J9csOKnCmbmb2iZ/wAWfyjHXb3ZQsgbnYk8F+2Zpl21
y1bwpbc7sg3ENHM5wRPupK4XxQaFaQl2gyBfS7qS7B3qnK/cFsrsuZUIPJ1TzpChANO/hqxbQ6lI
TXq1ZOc7TBEgli731KWGgnj/+/rlg3zsduFEFOkWN0Ome4izUPOupZGFIT2dgdDqb9CsRcxyW0jG
lhT8zADdGhYj22JNK9Ywri8+gPZScbb0EANDXx4qCWKE4V64u7HRNAOLBvUolNqB+ye5ZkUZN04e
i0hqPQhdL41OuGepvgXMaJSLEuG77UM4ExemIiSvJvs5w5WTn8oVuuYJBmnf1hvpFAg41MkCfj9J
AB0GfBJUU0c1cUcyqwafOcQgYd9ixmmsIDXlHEfz8+tR5hjAFM4fM+znP9xJn8BXJ0aTL3YZ5CXH
Wt3J8JZRuxnGmKAZDonqy4tmqTkxwCrxZpQmUJf1I7eTHJH7/gz3LWSW/SsFxDxyCcpWrU8XEAnr
mpYussXEkrhArdi0DmuipH6voMO9L5Jl7cmx9yk89manYvACpt9fuItBI44A80l0q+6mo25iQ+lU
9cfTa3NJ1qru+TZD70SOVu6Pw74Nm/V95FhFOjaRmZT4YvoCc5tFSVQKqfLIjXb+67XNOqBHRugt
qhbxUXne1ja1OVn8x+2Lz3xLl6mpkkNs7ZAoLjSX4YGZi62XH2nwMA+l9txGiHbZFqt9rM34rnkM
r8Uf587k5T8Fp50HtBjLDD/797cjqChhpCWbxEst9vXFVgOG1+7QNdJZ9THMIrL0Rtp+wHLaX7m6
qnDDTlqvkyiT+35TId0U9eKLVRoyk3KyLqg/FzBoAmnpb/SqEaG3CqpHzwHdqPsx9cUnrdiJz2ME
iXB3fRS/xejDSDdyYsj2Y8bfEOOA4Ww3DpXTR0AXDmsqEQgdOyE12KMa3fzOpPedqlsP03nOE4B1
LRQ9mCgKtC1IE7f/An83BtR9a4q0QC87hvtMnQF8bi/BcLw07btbCc19RIR44K1+K5CR6tOsPKKw
VEMh8InArcORukfBK35x5y/vJzoWlUr2dPxo3s81LPfb2LlDy0CYIqCPrapjExH5YdilTEe9kBEh
pbC8yfyPcdQphmglBZehxfy7X4p0qceBjgIOhMZv+NVeF4cRpaVrqGtnNgtHvE9ywdS4nwXz98O9
iU335av2QAgdBzNwApykzYD1oa3fg3bMvtRddfIUCoC5mOzO20GJvMLuIgU/1XzdndCh7pvoUbX+
0eGK9YQP+KkO0xRoZURHdMsr4DkYp6JeFDgKAWQQQdxIvlVqIm32Wj2yMH75Fl0CCBh8NpuBJsAK
AqWMyM4P1yj5cjz+ltxEg2XFl5xBb6Dar9p2Re7XvwXVr4TFlJSklUv2op/6wh2DeOldw88wfT0K
OnreQDXezhUIHgRAmEjnBgsDTucbAtDpMEiJWGNnQlSpB1PaWJN2WpNzvy4OeVLhN6SrtdWz38Fv
qHBHNMFSVLB6x3YVwpgbu0cjUcb8ObqPjiHr6ZnbKo1ET1acNutbDWJA9mZlqNr18sQJeKfW7SXc
MTxeLpKHp+fCDu0Rki03p1gKhwlX1HzdhHTqA6jmbR4Plx8TfXaEvZrzfXgv3h0HE+GEkKpfwP1R
8N8Le/9LPY5cgkg86zZLsiVktuygW5rVe7G8obe02GNESmtrHjJI1HB0jwtwwdWP3vYQp2iDxjhN
MP9sEYfNn8z+SBDy7gNDGN6eKHH7LcptQpdxXmJTwjvAAuvKnAZb5VgGEunTmxIZNBd/btb0Tbka
tuRp8ThI74Xb7lp9YfRU2wdyVsTK1CvE+goEQPg38LPsBor3XbejbHtr7BdZF8sZV0vGnet2VFiY
rs/uKGxc+w7J3pbIK2pfpjjP9rqgEzZJHKdkXOMIpXB8l0UnVooFYPrWbCkmRf44gMeGX8IOqlmk
GvcJK9Jm5Ud97/gKQU+qe+6ykIrlluDE7ti/aSuLmqLDjZAxm4zRM3jgghTgRKoZPi3uco+QSorR
iKPdTtwcVlNr4I4AMYbkYnvN9pVZH1eEDl5WFmsz8pFTtuktH7zmJCLPyCfQFhRzj4huQPkUYkNL
G5KaJAXUMH+f0me8iTppNgvnr6wkdIlrRWKJbUMStZdvyOaZNkqc8NXZ0JaYI/CtEmO2H6ecwIc5
WVU2iw3evPBzZllArJ1r8xkQ2eiEGEucKYbzxEtY299zXtQhUaBsljM2j3sxh2b99za/O9ED+TrA
LxLoryHB4rKd+l6IHWaFDyjtVHdn7uU7izQbnuZmAyjf4tPnBvul8a9hJpy79rbqGIt1uXQBg6CA
ch9t58C0bBZCCjeD01nPHqBx+u3FVSZrnBbNj2dn5r1glG4zr6i8ikg88DwNWTVScSyksT6ZS4cw
4rEjuccyZE02bcdr2ByXuto6qksv4wSIonqljGjiJaJ24T23Gvb9kWlxjyWEjcSzcbf7ZQtgKwGR
K/JsnJqFmbRCx15h5dMUfSnl+A0n/iqFvHyH9NfPu+Zcn6Au61ceRgRpYh81vqGJivL0ciGjemJr
YR6tJy35WPSneSLZ13spl71pWqLFY7Qm5UoBshZxfz1an0G31y2ReLNoi2wT/gR3PTaBrg8zONIF
aOXLDH7rSwcw2mQbSd01aMLpZjgDxaFdTJhFdcfrPnA662T2cJ6vNFk10vyzZnV2H9UUv9UQputH
qk7+S1LfTr9eLt9I6WWXNf938r2yE3aFcA4QMuvaYFJbrnRY2EmZ9Xh7GzUOyC+98fDDE3151f9k
ynG2gxBCXWkUfPlYlsM5owwbBKLhgYCGpP5VXqmz6RE1QlZq2eSnPEvGphHFdI4Wgd6DwXPwvS8k
5mK2FbRKNMq9OCbHudMSY4o9mzAuvXZq9v98dpSEqBCJiV+9NAi//v6ypbJ9xUvERHRqTfHiqVz3
rnFeLyy908qK9nCGZO8qTL51pd13JafltxmloKipdSKucYZ0SjkS7Re0tkGSbqf0NSGLy2m4Yb5r
oFuljctmPOiqjzWOG+7dmoYNuEUTW+VqpYbXfxBl9hQoF9xllnNqYvnzxQEJKh/eWZo91kCLyiuj
t7vCMoG6KUsrnUayGAR+LgD9TSqj/bGXehixz9LBr0kEQIK24Ar1+ihdOv+Tall/xZJPRFzqUiGP
HtqEW+ePQKldfNylK0tH1xVf6b5AUTfDDGh+uO5dwCjgrKiew/1m18nzDP0JksPuve0NrU5oOK1l
Rqw0/+LBqSexI+BBT/0Pbfh0kERbUMMpXRasYlgUcDgrUcdKKlmMDUYC8CzF8pfFDSydiRd5KAYw
6PGuzpRUK8s+Vo+qIavun2oO9bFudWMRvnxPyZ/MpRCRVlcEKHvS630C8NEkT+cYg2PN/AsZ8R8T
QGNhjShQGNbCJE1trPoMUjla52cFNZ2A0GV9mzNqVEvDxwCQIe/TuQzbt5agq7hvsH7byVn2g7n/
tyHe2xFfdGEq7wzP8rMVKKdZ9amtruJEXuThxF1W8XJPKVfVACg5zOEpAZBA/B5Psqr48Od83kDy
6o6aXWVZfurSBA0lCvyFfHtEH3PfzC+xqtEFRbdFBhUuwGd3uVITMojT57XgA57V7fVRl82j7VnQ
iIYlUUHZhtzRpN5rBMLL0h1IB4f7WXAihZ91XJ9PtJN1W7Bwx5AhxxZpbtb1774U1O/PHowFc6JF
0MX+N3K8hTCpAl2vXtWtPnVvDmgwXIkjfn+rHjWzv9DRKViXhCWsprpMIROXVcUiK8jLmHoQaR5u
yVRduAfG2NNVBL1zpevUTwLjJ6ZF0Z2SEceoqD0s69zxL3753FVTzdhXcwU8diyHx2sa/lFD5PVT
4pVm6LkRxdrPn2octatL0eT+CjIjTdlbFITysFHLekAMKyEtundJqalHweNBJcIYxL1L7VPZdNPF
3CGEtFibW98PPvsBXzrMIJjEieD8259fS1nxAMkiPbHwPSQAVVgRe9CT6amsS4TrWIxW8NpgcAi7
rmpOXzmcRIQ8a6OlHT1lh7KmoErcpmL/4d6wZlsg6iT5bF/Bhu4+IovAQ1la5qiUUpNi+LR9YzyW
di41qkNUsEd4SWogAxWb0dtnEISFQDKI1fqyMAIwfCzbmwtGQh3bg7OEqoafE7WIPomiB5MfFKB5
eTO9KUrbtkcX+BpmkiSoE6r4tJ6DWFdRQRld4viT4nOgy6s5jSYSn1Z2q0n5wjnoqoONrcsbE3go
ZiXxI1HHWSpQ/le2jgTx4QAVRv4wJ6hZ1FQWAPP7MLkCm4vk4w18kCF0cslJ6okstWRIwaQ2a8Au
OwWfwppDQ+ktr5MHwIpKdSj58Ez2ut3T6HMPhu6rdCfdn1oDH5LLa2XgWyUUyS3UTll7p6ZtdeG+
WVY+oQszdntrQBeq+l417tXCjNqvEJkzMGRCR3jXyWx+/ny6JtoNiPX8oz8+7Hx0bma9FF8BaPO1
jqUNIItXvwHuYR5OvziY39Ex4xAP8bCFf64EpcW7WJlYcVu1jztwOBLgMHCoKUflRN/C3rY2/NaY
GHec2iWkg8w74f76I9cjraFwIqw1yryc1IS13oZ+EdtWScv0xyLwyBauXIWv/L2lUdFmAQjYtEce
L1n/Ikq/EFazMa5Wtkngpx+/EfRsAr03hmysAUGRBcAvECwyZHbXOlEERw1jT7uSC+iBWLnv24+h
ZFJcv5cLFskEzXDMTxjVXavZxg2mMWL8+Ebm3+9DKFDYs/0flnwhFSovL8uufMxZidamxKlwVC9G
MvOhVLnbhRY6a8A4ejhAz/141Stpto8Fsz3xQuNWRikgCHNbM7gz5T/GUO1d1hoOwK982TjHNvA4
zZKo+LF1m8C4bg1kdbNNMOkZeUl6YZn3zWZuSGnsDP/h3PA0N57H9RBeARfA1brhUlP5X5DvJSvH
1khDHIkl10STH6CSUnsyKgvnvab/VXvQG9mgRFCJqSlvmK9SJ236H3u7Phk/eQh77Kymhjej4lnU
FJjPDaE6lItRdG6HDptwjuUg/AkfZ/rayjmvCjKZoOIOmczA9Z9lV9SopXUsUXuWwz0phJ3BPjWO
h4j76PmL/rMpxqrCpBsYb71JhUSydNpVT6Zg4/zPYVNqwNmtS+t1P6EcUkiAYPoR8aofg8CEJ7Fq
j9/L0UW6Sw2mQEVKx0gqHa6DU/Bhj+ucBmR/lnltialA/s5/3GM0k6sG/tHahUJRJ7dCJyMlM/Wj
kpP9ZzLz53z5jPC6ODs7XQIC4o0Iq2TgLFVn2ry8UTs8tcLutFhzugoOUaJcppVq0druguNC6q6z
mMl4WaqlsThgqngzc58RiTHY+Je8IHXK6QE881cos/uxbPr+gHdpI5KFyzZYhDUBIjg8O/wiqBQw
smnQEKCL/I5JuMhELhM+FjFmRwDTVounJvhYV4PiKHSl5TcfV9M409kqzrdWIx5CPoBNjAK5o3ur
ZldopA36tiQXf9AUeTcv9VEbNp3+GWejCcqujaUkE/3sl0poJs5hBSPHswvRoXSjzo9vz7dW3DIm
FtpYY7Hwz9KY3GUeVGMa7FHSsrZ1JTjlJ9bYzFr453+IbZn1gysoSU4xxCtnSGmyMbOsuSosmmyH
g+5w2KLBygysM4vFtHceBH9eNuKAId9XQHfq3wvdObAJzL8EYsbTcGcwBT74o4tbznXAOUiXWWSM
TJ7EjgshF7uM5icNkSCsVgJOEbN6v1j465ZiCb3kKJSbQDIw6kDf/dDbMFW5X5SlS65b1hy7Ry1p
6SaGoqB5da3DcycXmdDcMBw++uPxRHuiinaCD2bYBDqLay/hUJ4HMeoPOheRJs4/G7TubAdOe9El
JvReT6qWv8DGz08GGqpiBBfPnxo+F33T8sqzDf4bIwyBhEmeWcXXeyvV7/rzj/3+EyWcmNxp6l3U
gpqK/EicZanNtrfBN9NLA6m1Kge9t58ZT2gPAJje7uOFEl7tLCpkRE+NH1G2D2i8YHXNea8F3Bak
4posXE+Ae67ML6L58RZrVUeqjkr2v+sK/me0FJx2Dhtw9yZIPmObx8m9RLVv8FsdEz49i4vk9aeW
H082GfqejJp7tX0SN5aJ9XILThtmsYTTQ/OxKrgCBsUTs7Aov5m2wEfKnG301ReugHOlvQ+Kdyhm
EbJjZwo1i33qg9BRoZnYH27KMKTyDnSmhvr4NAJ+CqEl40PojOeK6VVRHCSXbT1wyqfthCntT63S
ptYQqO0ps+pPjCVkguJW0nb4DOS+vNj/3WmvoU2G82JaUT+8UqRGskicYrxPmm/xxDGaBrHX6POX
kkNfMOEsFElg5xwZNhWfAGiEmyM4xkcbvrodPxoF8ylYY4gPPmkM9A+VnkZiOViOja/5v8WSha/i
uOg2p3xxah0zaRJGcpSzGHZCnbYHKiRBTYxbFMKjZ5x0bRd9bBh1HeSFz82dY59XLafPDlqp50P+
fepmOpIUtToPxcKN5rHv9KDZ5f+DXjflibo6zZOEJt/ipgF0P+yyMowYgguPOfCAirwcM+w18ZT6
fYxgvGljkxhDXU1V72wN9n+AcWJPPGHECH3wzun/VdQJnuT7Z+KqDsfmeEjfr4TZuLgRLWyk1XaZ
gc+YukfzaJqOzFQckbao4p4FeTBkltBR7xbsmufzqc9C8PW2zaupX8MYMMU7WXhYYzLQVR+y54Kz
b6pOZd9KWtHt/2MkfdM45ZQGpgYdWMYfVhdei/jYx0PX8VH8sIcDH6nCy+lqT2y+Eeb4l2i9DR3I
dX0tZ5nMcmJ/zSzl+xktmUGHAVU5PLTFvkQdakDm/2z5uHafal5yuukHyXD21sAx5QWtVcsDnX+u
n/rh5MuZPHLb1iC4a+Ze44ecaFvcM07lHLUGTBJO6+LzRlkA/xGMTyfVHRiIMsj5B6nOnRVRUCQW
iuzDXk5tCUvMkgWMgnRcX9/XwrucpyLZvrj8svVz4mIhfS1jeHrgG26zI0dk8FVVku7AFIvbR/3m
TuYQmOHytQjXJsH0g870g9gyWLHBgPd4QIomaAL8/vw841Zk7lOZ5Fgiu7vwzYz5mK3kFljYtjNx
VbE1qsgTW8BE4+74zRC5hilCoShDVsoLTnbuPgdu47i4AN69GhNJXa8DQHHo/V9wfDrFnD3f97Pp
Sw8W5Golqjgy28fr3UkAS23mlF5gHU2nZoAOWQACAfZu3lc4YpM97jzkx1elTiTaUMzAqMiEarOy
heS1uuHWI9usTQavSo0KiBzWiTdNiVI78dUjB6c5+K0Gcbuvyv8EXEqq2fWwEO76BlepggXlivr5
4R6lcwzdLqm+6qe/xM0YBnHNN+QxI6NYtz+7xOnD63wF/PFh2aknH5XwPrCVqrbwHORldioBXjEs
5I/jNCd7AXKmhTTiwxhRWR+/PWxEX5EP2Af4SquQ0Gkm1ohLhqQRltprmT1nssynCMtQlFFDReFJ
LpwhjImu27nJ7fJjQ39n40mLY8x7as5V4Zp1wLN9yXuYCpPVtIP/Cqig5PKZtUk4R60S7G5YMy6b
Kva7z0FJsnaYAoF8ZLDHce4JN8U4pueoQvj/Qus+hvu/ALhEjKgPLcL827jG4gRsGIJWDbnRAoE+
xTMCo7DRL0w5xmtMSdwt4pRjOjvSpj/3+AnsvhjMcEONzH4smVIEJacUsVTqerS1Qa7/e/3E6HNq
A2LpdrIjn87JWoXahu+KGyMwrQJ78xZtF3Psh06S3xh1VitztVPw/PFK8G/e4Lzk9AKJwkvvrduL
pGiwOln7bN45rWdaeZtWXp41gfXvVisqYGWf2H5t2cDwlep+v7WbpuA4/dxejl6y5ZEmvWNSWSKb
XgyufOqecIIWWOrwzTHuHDhkS0O7LhSYuOwiILLa4EbENLI/kwNaqRaHNCmKjZwSeWFFGj9BMSaQ
bpJmEDxEs+i+DRCWToTN50XMM/KQuRfEiEd6JA/r1GX/osa2S7xBqgwyMeIUxuHY7ImbShB1MnFQ
iKzPShQ+TT6EaKsyXy+2jfQ/74v8u5W8Zpv2ZFDpgpwereESXo1yHb3JRMYeDn22qzyJBvUypoBE
DGdE0OdVLBTML6Ji2qaCPVxjaEKdgrtCgYX/zGhIZvr0BVt/eLTUDKGPobkeUF4tOWmRrcUXY/hT
T8spFzqaAqmtBzfZPDv5MooO0OZ0Y53fP9baaCwtVnf6J+mYttdFyxw9SUqS/fdHX7yWk9Uqryqw
wlNKkkiQmCDEyBjL91laE0FRiOl7iotbZoawPWbW7paewZmksV294CqE2f0DZ8tzm/5L281Y34d6
k/dFBag8B7ZhDGstaDKw79ga2xxGI5kpfHdIBjbmCTx3xygaco3NRdWouaWxfW9+bdExWFioX8F3
IOPQNZH7V1vUCzV5LlVUo8+B6Rt9tYJQ/f810bZny43QtxNVWUDJcx4OoDQo6Bzrj82KD9BPSsmy
WZd2kWoCoG1XwpWqSDe7eTo+6nez7uTDh3g50IpV9LVNEaoBMCCBkoVVyatgVLm/YL5GoTjdy7Gd
Ar3trrMlPYmOyg8aqlugNGEeP1jWa3MFvOweKolTlJg5w/RZ3ukNENf+GFVmV8kkFq3S2IhGyNNT
JQTwvlTqALejVUsBnx3Mgbcp4lQJHKxF05TXrYkmjdHu89jLg5eqiZrA1NKeBOkGYrbXpEtzaG0p
Kp7iJrRp3F3V6B5DxhJcl4jIKCYL32viS1i2ZEJZxRt+tn4rnaezgt3I7GsJuDRKHXv81Qs+wKoP
emR8c3ZKr1omnfr86t+ULsKBc08f48XPh4d0yvdJgzJ5cBk+LiK1KG6LjfwWa8s7OJcO8TH0ScV7
HIZHwhelP+5JzI7mIk3c+zPVKWIk0IAVREeIjfAJtWcR8sNAcs4/MPTZSGpiHoFksDi88mUlEDZw
E0hae76g6OEe3IDqfEaAi5b0WOB7VJknq2DG0c+mmpCHwpPSMFxK8oVo2zXKnx/8/12IV2TOH3EL
hTCOJKCVwr2AoX4E1y/sqnKf1fe8i0Gk0/nFX0uOyvI/OLIU+jKaw61nMJyUefkKL7N+Wat8Ctlr
7SxM7Ca77XscfRa/oCX1J5P2NUFCDuLTv6UIZSH0GDOJIRY9eeBAH2e+nXk72LKqd7fGQfWVKTpn
+IVcLulZjkI4XBQWJKqZYsL2+AlAbFaEAgbaPjuakwin5W9ajHLe508KyjtOn/M8/uFsh+rU5Pur
tYNELxvvyfOKrl2pxXEHDkm8TAYvR/PqXgkYmwCn94RJGvN1ee19Y+ssveCcSAJTg54DJszBQ0iY
pYx+mjIut57aNccRGVmwzaYUy25FUJdoePV5aEEu5UaPEvGtqz0Cy5hNfub0Nuj/m4x5SK7wdDZJ
d45I2nDLfgaF7OUTqMfsn4vZrmZFH78ChAY5Frnf1bSnNi2l5azVInaahhQ48f3z+8+yIlIqZd1c
DdfQY1nntvj0d2EB3PXzvu8gyq+/yT2ngBjvk48lfgYYABuHPff3IgOUyUxOiRYOo0kwz6n6nHaL
bjxZF28jE7vZHSg/7NkQhJa7wvGFywQIDkql/iTKhCppZXhQ6yAuI159c/RIB+Yy0f28cpAkZr9/
VWNkQ6dxjJ3w9p/3V/gv0JimXT4xbmX9miPUFq1USOvxLuxh8kT7U5NYRJPoV3VOnQ/vN8SDXMhq
2yd0fpXt0BMdLsbVGdMstqOBqXaU7G0Lah/fke/yFc2kZ+q41tIpeD7XwCzPrvhBOXKGqnLxQrdD
PRbTfmPeM1yWGAJnuT0GxuDuHHL9KCgFeIi+7P2Mi84zEyExVmSxqoVZdja7Vb5cD4/5FVIgDMr+
99K19L3z4xnDEPiOCeiiJl51ltc/yrl/KCOeAGdMtqiYYHo9ewFaK4o+5o+GIwxPh2RnwHMSyZZC
PWgaXJWosoXqMIQ7wgTp1NLg+SqjaFp06jx/YfRL3saWeYTyahm16s/+CijdXuVnrXVLtaLTk1OP
l3oplcBMsqvrCxzgJwbbKKYVRjvG8W7mqnj/xWeDqqJm5JIEUnhdu7q9hCFSZtXZvWe3KV5IQqaO
fzIKXQxfcGweuRbNNj2bwiGAp6BjEplE7B3c64XOIuJG3j+EqK/bNK854Y//JeUtN9B2tOn7cFs1
tMPvZ3TsSY/D4BGRCTJH7MG9d+6dnkRg19R+Hup6WT/LcdjTnizdLKD9w/GmYs+k52hW+s4iD1d6
/eYP95CiKrjCR7jmrGIKklwfRXaOOo+Q8jt4oRyJiZx5DiMMbIeECMvzy+GCkaLG1TaN8ieNmQz4
080McVilIAarQJjIyGsSrz0vSKlxkhlJSlzE5qcR4ur01mwxdYj5706938cfEcXZC590YK129MnX
VcGas23dYjbCHLftiKjrRqzy907/TfBMEIBn7jwiFVnoxQta92KTfoIZLBac6+2nSiyl+Mon6+RG
rbSfxhZTxL5u82Fs1txveLsEV9yeNHgTbm9Nl1jgd2CHPEbc7S6hi1F6oMVxg1qUAI8WaUomCvhF
3b8VpDcoYoPO5BXytlJINfkfGW1XTnYRs0bVcjmU8XmepJ/hX7xX2BQbJ9ehGUFWXwu1WSJmyVXf
FeGzcS+dcsnkRzhP0aDaQkc35Rd91tVj+1PF3VZArrsKs4BNB4UV2/Q5sDrq/k76/AV6ArtKtxvZ
aGy8yaa6VqDDeqvSEvnBFI31Efg/V8av09P1bS0fUYhDdKVE9FySfOo4oyJW7N+4T7BD3dJmp1ZK
/tWG11hpe0WYnLAaTi45U3hkyaspjdstiez3o207VSOp5DKrHxntntRkfC+EHc7aMchA85L4dG7L
Z6vKjjvssFTZlYFZ4HOtzshX+GVpqrzk+PXxuoEU/GYLV2H9c+ZzgB2lAvwjaqsfyY/307tsrMOs
HynEIf6FH4SIlDMVASvMu97Ku4arQYd2yTHcEsD2kyWPbOBPYK6aR076VrGASwfMQJDzJTcQYgyb
Rsf7g51snFoLU/6Afv5g4U6QWRssyJl0fT5ifIfPd2y8Wds+DAQAxKzWiGmpmse9zSwp7YuE1d0z
qp132v6JFT/07TcpJtZbZSsckxKH+KT0mX+dEpqmSRvNw/oY3L65V1gxhupYX4T89E4N8P6QeEDu
902FHoIVhkgInYkOaNAIF85DsFBkS2/e1Zat7GEfb/AWl8wxleJBmdR0X0wP7ksUstugSJDDnwd0
r3ujT99c94FyaLbEUz9/EcQWcs1wPZXBv+G+Is8jwJBDhcVKMbrwW12UwI+KVe0r1kOm8I1hunTf
hFPi65qJu0wEeb9qC73GatolBuDEDxazcw4aI0T2vMY8WFe0FLhj/6LTleKGGaQjrMAq6op7bFuC
0LxYImVAnLuK4DmgOb84Cn44Vah9mpza4tDr9CFIL+WqdhWWMy+io0HziLT7Ymr5hwzjOGjWTOe/
XphAWXzPzghYA1m9Gydvo4VyvF+5OVZZk1zMUAj1C2LnVRTdTgs388dUgPLj8NMFMIrAD7PemlkZ
2Uk0pGME4JzMg2sgbnvZ5gNI4ucld2v1HPXn54TylYUl7jDKqjQUxdrFU077+j60hom5nBMybGAU
EZmKLcxxCcyc2sWcGvpibgrDpvzgjzIKiT5vExAPsAOT8nfBhFeiMFAaHM7jdXRdS0hB5GxyVAeX
Na+BhjZJkbLwFlG9BmiITusnVVN1FB/gBNzEw0BBPhhTW+lUSNarY9fAMIkKI82R/CdEcyBtyZnw
Q0+zUukk4UTfRaTtcT/H1PwR+Uip/q9zjiGITelsVE4cyAdEZmNpPkl0knrm6wT5Q+kwCxjFuZGr
GJa9ZD6wEDYkU/4TzpMZxgw61xaIbPdQk/HAHspYQGit70wYqYXlmzITZlKgcIm040dOU3JPhHQG
6lG0CpyfEUx60CWreeCrNIGTPnzWz52FIW0zEYWIdJ5sUwFpd/YR8yyW5OgXqkIgH4lQn2265jYA
rfHifpc1QeCd5jPq1D2tK0xcZIxE2l0cEC4VFm8E9jbY2Fkr7Rcey/hakkLvgijWCUe5ht6MXH1n
oYbPhvvHbphDnxrKaT18tIvv8VGBz9+6U4hHt4XR7qk5zENBN9ryb6nYK99JYVRBHhB0NR5M1+FS
DBmeDcmufnSawqeVmtGsAXSzu+IZ5UbXldpOVq0i2ds3lRAhAKB8m8R3inGKJYqo3bf79g0wGHQz
lkedeCws8KUSnu+Y/i40BLtNGUeZ/y1GKeXdzGNoPrU0JSNNIme3xKJdYY47YE+EdWucM02kEBJI
8KOh6x8UZHYzEFd97HQ3w+K0fZHIjFZQCXo32F+KqNwMjA6r90bnoTFf+h8BLpzvBNyL+fCNs+6m
u0YWTZbOq5FeG1F71T1Wvd+XZTKLWydmP1avIgSfrwW6nT6w3rO/cG7giOIcHh4u6WVBJj6dxqdo
a5z4WO0MOQx/viJtWTxpJYm3vn8dNcHGjwpqM6YlFm2UbPrRrdnPyoTjwnmikufbUyHv2wclh1Pl
4noZmaP+PNFpQ3RyyNsjB0Twfu+1Kw8I1npIfvkInWpKdBlNoH8o4q2yOnmHgWeMnRtb0DWXeDFe
CjZgnIwjsWWuYMducHRXekmp+GqgwmZSK1xgeOv0z+YHe7GMqaRbFRru4njQA9OPVtv/Rav8lPa+
xA+WZ6da75ARZdu/HjK8goRaHtuIclqd/y3IZ7QznCYM7P+cHzQr1H4lzEoVK0A9BbYBIBXZF5qT
ZW0A7+odIBi2TjI/UA+YtFHKiX1b9BuliFtsVfofg1AaGynttwj2xBYwrEm92n0FivVGFZ2L6Z5A
G7pB9nZ7hWPLXlOVtvO33NVd96iFlbV29HCLJ5Tw7KCN+LouwkXzDRvdhH0D1KVHre1Bs4N1DIlW
2Ov88koTqWitFQVe1wah9FA2oPbobUOfAUophSJmQBCcwol+4eQL5nuGHbyqT8l/gr0kzZXLDONk
/MV+rR3fItwY1vYnEz6zWlrCRCqL0TPH2vd3LGRDDkpXaz/OVj2YUcLRA73QsQtrA8SDk4hf6x9k
NLcsfOCWfGWlVXxgBdmAl0O1c2G9xQO3zHgob7sODy6BHAHovy25fuCTXpdXsQzXNhOnfCLX+nxL
KAuz9rHHqeoe/3wPIt7tdavEf2rbxWXqrA6xB4x5c5RiIKzJyDVv7oTbvdhxxJ8mrC/k/9uJFpuY
4iA0RHiuAiPCJlh2Zprnxt7mCKiWy9pSw1lyR1/bpmJ8rGHw45zidTmfm8BwpaNsdaz7gm25iuUJ
Jt13lUAx+M18NuFt6UHLDABz3vxSDhJsAEgj1XWfydj5Cr/DsZaxUeNnBvIBcgEW9esyWkQWK4Rk
BAklSDWpHH/3/7o3cIwZfCJGuWvXDSeB5Kxvxhy/w7LZri1EKPDk3rdnC2ium8DzUBd47kLsqAjj
cpcLcHAs/ODX3fMvqxV586ZGWeTuEcCCDBaLdw6kiC+mOGZzzZWiU/B0K6W5PS/TQ++CCZZ4uFYG
yRW0zZTvaZb3zi8ToHjVo2ig9Vg0cmDyMcPuAZZiwpeYtedgJXfqsDPgSz5EHjhWxi+x8lw5rWXp
i3OgYk5l46PCcDoa/t1L/M+r6VVzInx+JPDFyt9tcRDbhtCDH4Lm49hn9RXi7ztrsYTPstjUwHXY
M3qJ+ODazO1qQHqtm5qkeQvEy1BaQtOLmod3D3OG7XdNBZp0LA8AcDa/JHml+rjLsxYiLkicQ6ts
bTEJ+lV/OeBwOo6xKidyK30x1RZtomDew6rwpxrOtNjPHItQtYQzQSyu3fRDOpPkwtAqc9uD1D9D
iBdsxW1YvXaxzmcrit1RkvANCcW3qygX7ye2cslY2o0PL8Mf6MZtOcQ/CbvY3O8lbOTsjSyjtlji
GAWIDR28QadiQmdojowbucDVeLcUtnUje57GXZ1dTAf19WX4FVdfcCaXZhmMQWEcgEAIHoRAGZRW
rYpbWe/rhNb75kRf0N8vpZGHNADEW4q98FJu7/ryFig9ZKtQuJV+SFlUx+7CtcaVPwmGUQNmfxd6
XfdVxYLzxCXXUSK0nKu4URSI29pXLuEXdRl3uEozpcrgmoFElS7LI0IFuL0FkUCUMxWp6KH6P28R
36h9NMaaOq3VftzGlkpj/W+UmZShl5GZKQchPa3+DVbtOxbC/PQ6tlGowKDSKptkDIIVWXFaG0Qi
ew4tZb+34aG/8bpNDcP2flj0rguilM9Qy2wsddlG87KGmjjwPkK+kF0v1rxKYthSaQCeW3O47/34
j5juwuBKY1uQYYGME0Tpwj1nAUzreKTHWQR7onNYAFkUxV/ru2vPoawdp5Q6zsjX3UU2felPUnPQ
iovg3ExmM2UFy/a1+b7u9vNxOu//CTWfbJfoDWQxbUgXJU6iOryz3SR4FkmDhT/7p/ISEQAdV/3n
jWYcs2XoKqdwCefzI848hYHfilZy4DRBtzUitWdVPqzg9r+jZAgvjRZ3/+pWaTVh6gZaPghf9WLt
9bKxfdKRQ8t9lQjNj8Bd3hHNPvDDos6oL8/J/d4qc9EVm0JXDhH8FAvDPXx02SANqFDqTIRO5y5C
Mwg8ku+2KZeqwjpJqIDiJfERqL/z4u/srF6SJ+f8AXhiFG8dvUXEyoWUR95M79XjJ9CV99lvK6RK
Z3hi36c7dNjWPt042N/hcAnLFNEzJy+kZQzV5TJxJCxupEQizpcck/cRtNI94R4/Pdp01ud+g8om
lf8mtRdmBR8ytG4lv5086nXZdk31zRikRcHdEKeUYBpSwRfGFw2kWBKBmIg+JrZigh4ldOQGnaui
MJBrzJBo3KkWqkz7yRewEg9zCvEOmvczQSaV5aVGM1g3coyA4XvyJ+Wty0d2Vmt4n/ZN0A3fTMSA
Uog0ES5ColzHfYK/bWquDp+LCqUJIwKuUfhHfcUZ7z46rJx4cAUE1drCm9E72VhfCHHWEpugZE+S
Ya6uOmTo4xuX5HCyuwxOQWaUTqun57XI9RE6iMInPd+lBsayN+CpEMvlJI47i1WcYDpYa/qxuwIu
kV3oURprxXKG/E646lyuRSpWsurejOjn58HXHGno02bRRtVU7DM//bd8XXDrf3tUIMOgsLDGz9XE
W38GCeIKAMdqq5i1ttkyabJVu0uIJSfnix02RlotBKVK6dtWcpnVOi+woqJNt4f7RfxD7Qe1ueum
65bR3p8XpvIOLJfMnsNl399LGdOjgnuteh96LuKUMKiOX1770Hcs2JTbgP/agF/q0Fi4SJsfGv41
YrNMVxCfO53VzCXpqu/vHbk6/FdglPvs0+2PZZOfauLu5TR8Zgr8Q7/kaT+fTMu/p9UiY89cSsWI
Kqz/sDXvVTlnOJ5glN13+UAD3bpzsZQETmnBipM9msGA3v/cIbwTU4MjOyCLBPvdDE7Sva37I9KI
u7k0d9rc+R8nG5ZLVOyuQhQXdeyh8g6ddUK0mQS4c27XCtbKZIcxm8cY53mezleKkPxN/ytXmd+5
5pJk6k1lNUEpUh9n24D8e8mSpDdzApXUyQ+M6szC+hbQ/P/q+yrP04cjzqHcKhdRDevEYURZ/J3i
NcM/xIgVEj52Lcmz0ohjShtgbTl3mgXQdzpzFa3YGr0xa7/XfHp8iGZIJlewfxUSfe2F9rowBVhB
28gnWfLIZV3hJp/KmEiqh9KfQOf5Q3E+fxpOXNHzMuUoqhW6azINE/V+l4vLURnZ1EX5q0d+SJcc
FOAI64rQUJwSkVnqWDau6lJ98849RBnZuryUuOBwmMkoWeT2l8OuFjilLFsotrcJdiSGAxgF6sGh
IunFyGsCjLtexpvYKVeyI5kAPM/R1/uMaANz7c/HtzIYOdXKHqS4Rdb/mAV+65g8YyQvsQwSZBKf
zkC9jr7cg+y82R228Vr9XD5aMx5NfJ3gSwNhgoCJEOagjMYXBZPP5jKmh6VtfpfhXYtGKe1Fi6OF
5htTnyuGAEPwbF3YFa/uHBX9N+15EnTlA7qt1DQpxlitilyvKdiOaWXQuxkWNUem5eTLRMkpHdKb
HmBSJbE37dLnchTLRAD94Uld2vPzriC2d+tJ7gDNO2n58/D3F+SDM3jsDwdo0iypogs0jhNVpcaw
G5Uq6KnWc2My0N1dkbwe98TwNZ3i1PGH8dzQaVZDZsvp6LhT0MqmzUK105fAPDV8jn0r+2oDT5t2
PHaHE1GnFxYCGyIjEA47XJaPulJ571fL1BBLE4wRrJdiDz0x3BGnJKaegxWNe6n33aN5LM2I4c6n
nvnlQIewG0u5hqZDcOGFNcYx/9yS+JV50KPoJ95i9xNwtmCOWjOffkSFv7PKCN/1t/NrMDxhna7w
AAwqxUVIDWAQfGOfZjzpGBISjk6wEIHBF3GAjMNK1g07/jmvn7FGLHAhAiBB/70iPZTyG986RIbm
WD1/laX0Lo+fos1/xQOaUe58XZPYHEO17S4yJH+ZP1/9fJH56+Yj38n4j1XWK1felIgw2+OYchtp
gssUk10+ImfON4ZOGoF1AVX6ofyXHS4+pEWoP5fwQ38p9h4lxosbw1jkmb1Mx0MSHptY+OKxnhXG
fKabc3rJRBCJJw92fo6CsMq4z8I5/djEs4wTFXxgC7aIpKJRgEU+bBkFQOR7Gs9sLNj1TRYRaNKx
xKOorvko9vpOd0IUswok0tsKVNwskVf0C2XcoDpaC4eDUaPV1SlSH4VGSj7u5EYmDNabDJk8WHCL
nxJRJoCaTsYxYbdb3ssZ7EK99OP9LNiwC9FcE0+96e7B8aXOKomNL91oAu51iOykpnNF6yBseAVV
NAlX+IFZ8UFGfCp5ZrXsJZLnSQxxt1r2XnimTbRzRFWUKStxw5u2X/0IuhYcinKNcQEqz29vl1ss
QUbggpNiYjQ/ZkOkI/YL68bIfKs0OFOBQBfyhH9dzElmrNR36KCwdikaAZHboKTrfNFz8DX31r/k
PRy5B0xy/QClp3pIvSLXy3UkfNwnutQ88Z7XI5/UnQlWGAys0Tvz72b9h7xzWDGqu+S7uH28mvvF
pzeZM+rrvCopi4T5Ip2Fv38aQY103/fHbXAmanjlCBS5GV5lcHVryKfoydd0i/atyXAFeJ8PaNLL
Mu5BN3WUJTfCdFY9jtjzXTwO9HDzsDkTAr97ZVWb+l/HApIieJ5Do/y5GhYiR9M3Kz4icHmChwJp
XlpExQtVX1JurWGV77Pap601X9Lrngpxx2jEerJsRPFoQe4Pg5t20IWrvrJ1Lygawop8p8N/lAdW
eFQeLg5Rd2qx1D/5cZAn84H1Ie4OuQNpTMXnRS/o3SouB5JpeTRsEyXccUw50rjGk0R46oEUYea9
IkV9/u3FqvMgrS6JM38vBUt0JaDChwQRwRmNJSk+9vGVh4JZ79AQdjAqMcJHtvhjb8fdrTaES8Ks
OPvpZ1U5uLQNF6IhVEdoKgD9C9oyROc+phH/83PyPuLinwhdh1b0u464xHqS+5gPNeFDEi8czwnC
eztCRcqH0VSjb2GH8eg4KDyrzzGkLfj4Vivr53vy2mer1WUlS3CLMEORgmiUYUCBlH65BrSbLMmy
19CRxF0y2m7dwz7o/JGIbDkfzKL6pfiChrZ6VAwrivF6XPX5A+1AJsqzBUpABFPzAckd5XaZPWD6
lX8KTwyZCD1IHNf4AG2WqfEnlusfBRALGElBnJ3Ts+QJ96m/LvjPhZblu69fYiT79WuJVcOQ2BmO
TbIJ7N3QwUgiHIEGWRUJADfduljWM4qB2vy7ol8xw6SbJ15vIRKxqTsnDhntzLymtdzymDwRR8mz
rodA7IIwwg9pDM3xXWJ8omgPaJ4jBXAO3wy+Vugu70MIcuHvKv2hN05m1KPMVAuzkW6P8EcNC+q3
u8T5/7c3ry73qK6hXR2RHC4BTdDF9zHLxDUssATlYb/VHao/hDhu5zGKh8lF7Ay1DjCqpAwLUYlL
CpVabs9Dn6fCr38bk2Qacrwq+xuA40oLnJ+pMPk2+4drD3UqBwN3wMOpu2mGFYPJG+wCPz+aGGra
pJRbLz6yzQ2f2DhtL+f0e7IAcfS/VXfol0r22jo6PE9CcfQLmWMMJPnKxaeC2ZHD/YzFeAkthkKq
q3ZuvbmsS5C11IjXM0ktuTlbd24asedtunReeOrPYeDVVu8OFM3LVt0UvrdqXRI5rhsPG9crhDEJ
AQl2/LEbw8MiXWhZCq0zOFhlhOAOx9bFQhy9Om9NO+4ixVaugVo0e525qNqXFesRCDCx4SVPtdy9
7R0+0GqGD/xgRR2RGzshElGNK1Lk8MehpvbZXaDm4/WaPS+1mBh+OXbW0HZaNRv+H6cLtk01hLxz
oH3L/Oey300shbQG11KACTtGyoiLLcNVIdWeDNOMpxz+nIYgI1lU7Rdt8nqqHSdInpOspIiAH969
FccP9qi8CR5mXV4d0eLcdr2pCgNgqcaB6Qogl2spJLW011V5oY37d6J/ntjhrRvzAdoRrVXP4n1N
ej8qCmU0nN5QiEC8HOEj3AgCnBQxsIWajsptN0PPbe5TZKrHtDkWLUGBz3k+4cKL/91AAuXlOd/U
L8xe3Y+NOzu/t+8Vet0SIrwithZy/lRTM9BDj7ecbwflU376te89JsilRS7mK1ITtm64KGtxmzSX
vL8KMEuOyhYBmm6J03GraLj+xpRDQRM6aHbF59Ze9RE6vldxKtF+MKd3Sf6pR0qQRnNDuupTnj6F
ShQdz+/eFSqgjmMbsl2s1vImCxBfZH5K0t1RXOvJJsWbsQZV6qPxHc8mT30Uk1Hah03Cwvvyj3sT
Ic8hhzsU456F/K6L2qVScK4ytg2/kSCbHSIQMBk+Bgw9OPEW45Ij1e4RL2oLRikSsZBLdkc1Zb+K
AJoVQpZaCPDFFy4XKl6Ku6MYv0/569WYsUmaLOMDaAE+KkM7/3HnxOzSkCLU0Q9nSrdbdmaN4rGl
3N74s+B6R8TK8767O++QuAMPSJRvDIT3tFShLEOXT5lf/kE6wB3AbiN16Vp1mKGQodVZsZz1derQ
YWHVA50MjDLrOVRdzMkcmemF7A2jC/vHqQJnRl35q+z6P6aVB2frFi3eIANHe+PJ+If2G176nCgc
pIhOcd/3WyVhybVpPsNRVyRELFnn8PDDCso0rxvrxPoL1eoSYur2Pl9QfOJ0KH615003S6nb2MPL
X/M8teUhbdTuRMEuqJ3pQVAI3r5s5paWbBCT2TqsZnieFkDCiVxjzVJe1oua04KJUfocn440cL4j
ZpfZecy1luf+jVt2nKlWQv1z6Vuj5VoizP7xfiCOUsQhGCOc6m3kyduIteMw9OFzHUHLxmDoMNSW
durcFtH5CfjkVd4rVssQhpQ0VB9R4gLtVsYscxvg5+UZSRD95TW+M5Lyg2xdPQuKq/7rhEViz40p
4WP5XoJkfqvStAkp10B+a7yy9BFz6Rqad05EkLV8NwTGIqT9QvjDCUcPL2diwDUAMLaGzVR1bs3j
4j7WZl+tRUoWnPaca+zUj0GBegBhwrThznDNDfrax/bks4pZWbK+8HhHTdsqlbibsrKiP3T+uCFG
HNaiDC30qgsTcnvgMaXTVzlqlJQ2e+xpX669eHD78q5Q2vvgw1/zJNw/Sxi1oakg+HW1kp6Q3r0R
exCkpqlynNUBccuyzyF6wmrvQtF6D2KgH8bimCDwM279Wg588vMshSjzs2+nXVqsJHTSEd7RngaR
/MYVt70At/KlZ6j6ZhKpYQ18uVhLVk8+Kl1PtD6NNP8R2yXnVKlpDldIIkfq8K+yYik+xUeMAoiZ
PMNTK55fyFYlFdkM1HI6gqHPthz1jjXS6rnh+hucP7rKfjPM2MqsVxvKQjsuIwcM5GYp22dWQTt2
cAE7qnHtJsMC1Zb6uDRj7FpCvvIb5yb1YNF/047ZrwswfTUZTLRA9VaSlkr2zcVE1ZIrjdzPPt2g
M4x984QEoNdWGqGBxyKFdoKMQ/Efj58JZbVkC/oTtFyfAO6o//j6kGmT+AjnWO0ymVgIs6Cv2RYR
SgB32eIiey5ny686Cjhu2Z+9nW+ztuY1cunEGR6sB4OylYrBp4LvyeT5op9jeBuqwDkUK//O7E5d
hJVpUDLa3s4M/o7zIL5vKsShb+bxG36Dblrg8YH3VYuj271fQnCQ4EwBvlPvaxJIL5ca2ssNrB/H
k4XKyXxzvISTTVTLntSG+Eiy7pIoWSohDP1QPuRC2VqnO8QiG9LCDCIMZjooa9o3o1Mkfju6FfGJ
38hwBkricUonJwb/gXIGyALKIzMfsZ1LhKH5+X5LiZhFZzlzhTGqdJ2vdWTRVSAxqUfMLIwmMTp7
HT+QrWFR5HHNWRfBkYV6DjuXhe/aBX+LrZ1sZvnOZvGsT5eiOqJjRLrrvqZdEEY3DiARJSXZFabU
lCwRyvp8qeifEt2XO08v1yAYNMgfUD5YiRtlqT1+GGU5VYWeonnr6hL9N4hthjvf9hgkFA8JAiOi
aXCDvnkQMB6XeMZUH/+T0XubmUaUoOng9wjf4IZ+4MwjJLULPAtZR2zKssUGD6gL/wXloHSePEKQ
u9P7Wsea7w9gJKH11D5xgJCuww+8XV+Ev7q/3z9OBgWucz7hUuRso54ige+pJaSM0xXOFqHCWdkt
grxuFigu1ePKOUEXHn+vAF51r003MR2KR3m1fhT5jh8JgAtx6q9GQOci5w/okO4Jjzxk45UoKe8w
VSAFS098gQ+wVxuDnT0iR0VvHhWqyFP5BnJJAAGkZ7G6r/+g52zKWHdI5tcfrCPRXQ3QJ0KD5m6B
WAvFEm2mGu2ZDJK9V0QvHwZ7YFN43TOEjTafoL0/pg30hCNBqOVPB7uGM5pDeAOZV4SmOnjyuH9B
yvhRWQQWboBlVr7g093RJRf3wilAWhbkkgkW9aBi0aE59rW+A7YALhFkkT9h89uH6rcxwaXib5YI
w49RqNeww+R/NPsagKUitLcuHMMrAuUo8OdedWxlNYwV1XAjox34VR9VY6EWIlMDf77ga89lTPM6
OpGJXEYvef6EC4y9iQUcHdJF/mxMAgnPLPMLh03IRxq4u4xzrC8orl+05uzN6LrOdBBndaKndTxt
E6WgNSrV+XTQHxw217K4ODf8KPugU0uwCAa7DAg/FsH2vmtwuhZhGKUoC+Ekh6zszFG5meqcs8re
hY3NKS+zJOWkGOu2lf8gEsec1S+G1t1DX2jVEUFs3s9sUMLEoW6Lqlnlgq4Rjb+MT9Zhrb+5TxyT
64Io4BP5ARJFXu2txu9Klpo/7PZdf8oLwjePJLRVbcVnsF1Z7f0qRKQfrjovnt5TlN2lF43vyPtx
DEhVnDzxu36N2rYPhWw0a63iRGB7PHKUgt2/d3euyTGgT7XdFrtW4YOJ6Mm6XQSaW1BJopiC51BK
0dVKtpYyOHCKsQzpbY1bxM9+jxL55a9StY1UAjfoikjYH0rEEXrF8MfAFh1JcU21kNMrmmSaRV/Z
xGu5e8Sfme/948GAqQWgWpYEhy52uC/3CH9vfOjXBvroPPHl6XHcvALbTRO3qBDFnInkAseYTIVI
KS2YMJ3WnEEOnScFJpILFEk9PrSSC3S35w9bCwSMTAWmyqofXrkxgdUX3BvJV114OqCwLTA7NIGN
yEvJ59Ig7UFfMHCiXGWP8CBj/p9I04NF/miRjiejQUOTjgF4pE2KZmvUvuo6sexzSBFYlCC8CIf8
2IFmsCKejUlh6KUWjp3mbKcFjEgKtgKlDXVUgnvzHpChKyH3nBJYboNs4zJCZttHf2ZcVQBT4CCt
Q3yhni0yAjmflqyQekcqoJs4LoRr/6YQNDx8QNTmneaS/8FUqgbaJ4rPAFOPz2xQijTaXvKm/r/4
ua23NNE0UiULQBSm5v+SdkgTQbVctpdhTglphWlo6gjFXyij37s52HBdFgw2l4H9gr599JjrlEPQ
xBQUOMjl5Y2YVoSoRFsZkRng8YZWLlq8fKRia9qk5pQgcD7EQAP32LAJb+9UzynqBeOkAD7fkxqQ
64EcAQgDUh5er4N4b9aLWUBiGJngUn/Ipa3mciybFmc8DgzmgXgfh3tOTlSyD6rmA0m+iIxUSFf/
TUFa+rPtRKbXQ9JFIMShyJgNPt0WYRx4u6Se/8Q/LFfZm9xVxqTl19q0qcWcKUbvVf++HLjIfgvM
pXBAfxW5NdiLBaO0911OofoZCcsn67PvkOxyDyQzqB8k+mGvkLOQ5tb1F1qWIUJ5GMkhE9hCZ08T
zfrjmoHN0si1AqU5HtB44+PmytHlRCxH4BQVyFcMRjD1DCDogCq/vh2frt76vbCW68mw6IkGkmo8
tuDbq+AiPTEZPw4Tb4PH9+Oe1tppqQUSam7/xq3ZLExO7SrGW2poXQ0bAgPJM08n/RIYb2dKFDa8
0m4+3GccyCnk5JYj1bgX41+9GaP+5A1DfCjDzMultSQQ6f26A1jbD4lZHm34T8GxnaJ0XQpIR1nb
sTr3tNAGF4i3UqWtzdLsH7XgLXqhxTgq4PgkS63e3oK9AC52w3i3SABXVuSchYwCmk1M8kJ/Fu3v
TVVr/bqbrCdwVYcI3HNefMajbdzQnjpCJOodG77wE6kMb6HzO9u/lF607ILCrnSdYzkT28ynSjqY
FZmdmeH6LaXvMgWBrYnVMjDQoiDPwFEgG5Cw3AAXHuTKYEeZfw7bOyHzkD6pfMkzjz6JMbXNLyKU
YqdU2OPDHrAo1f8TpV/8xs8k5KaYkh/ucxIXQ660tP8nJtZYj9dYcDoieFLo6G3xbq5KxblGl24i
be+fzbAFiRP4wUOXkKnikPpQWxW7WNAtWASf0x7/7QFQJQJoJYpAChL+QlNSZm3xbLnpBZL5aiOf
kSHwMmJ4cKwpMvNRhCYKxpmuaz6z8vtFUAWaqQP44fyXG6TgRGe18FCN1qB3K3YpUpuxyxP/tqSe
520Xmf/xGTwItAyqQouZ9TNJ0de1iu8/4w3a7dWkd7sY9vPaG7AHYgxtte1aHObMWeUSuK+fWeej
AiNmmHKB1bkFdLAFP2G3K7V7iZqnPgpgsMaNa2u6oMhiBiDoxiPLPNpu0pFYhDhqPXha3OdHLjXv
bSaPlwPCRPy6Knr1BoTohHoMvwRJ8cnuGBeuTXMNyM5q+UoB63IMDmke/VTrxaMdqzvqHDHITnyW
yGGknqKCoO7BCWgUbwXllLLMxAIrktkUyEztMLh7zwv39n9v8DYn6EoLPzaf1Hk9gVDHr2NLLfDB
/S90jnh6KywUz9m/JsiHVY5rNb0NOZaAfsz6+UdAmNmInhKw9IDLuwq/+Rtj6Fjt+YF/hWvQrxzL
tcQ7MpyZSzKHyRfS0lyy4MS+UPFS9LGF89O6nIIU5HGCBtarKEsEAbJKir/bnwLzv70KncS+iEve
LZGpMel3h9KEXQeCtlePwJlM4SA8m/0bHIYCIgFnZOtpsKg5j0MczXgfqjwHfZuwtq3olNDR05N7
Hv636o32BZ+AciO52F71NZYatL6kMBpJKIFlJxqxPOESD37cgUt3PhCaVIbgGLN7g+7et/WnaqV0
UubVmLZSLX12/zn7uBU2Is7mKJRy7Y1z4m24qmTOWaTe0L8o051S48bawPIeBjnIBGXSgdw8FAU+
q0ZfmjgRfN+9SYpVsSsI6cn7MX6w6NdVmrG5dm4XBGHuCdS6+3R70IUAE2nQUPibnvh5/z9qP/Ms
Y08iCU9gFkf/RUdi007ESrqSbl7l4aiZA/fSm7StlYiKaNTWhpfl+Bcj5gcMUw8GkhT/kBHXJcAP
pb4D6AcNgZ1pPPAq9cfvk0s9WXJfCjygodnsTCV/EPma2AJdA3DKkxr1Ghdzvl7kYdTFORNENvrF
eCUsHJZYoeZfHYBtPJ1K3p9aMxHewBs8uzdARBlBAz8KymSpp4txLL2wuiL+U0kKF6cxlfNKOhix
J9ZL88HS3fJ6/NsrtY9/Sbv0ybNJMXZEe9kmEoQMRFDiTmF44MyDq05YaLy0y0JEn7GSicQ2aBmf
4pOETv7b0+Wrw4FO9MaulFk5vvKcGcB3tGhzARw+jp9FuZNfW/yiJC+SjzAkRj8uDCPfpI/cCIr5
jpeXPh7jvUrm6GwMMHXMVs154hAqFbVRZTAKMD7QpMcWJiVmpLOMPTB5kiwLCSxOwl0WrHgpebMM
zEn0QT6YMV+cxpvXZ4sacycgdDm+LMIIwIuakhxaEElxsDu4BylRe0g+hhtCE82OFGXAW6k9ZDpS
hfaGweDiLh9lrMokGmcJBDQ/neIt7nP7PS0sbfgIXt8GLS7bfmUaQO8iS4FKkgmSQghn6i054CK3
68A3ljd5x76CUdcI6PdwJnqAJ1nlCShHGRR7AoVji6JLp31iudYhDCo5kx3qKwAjIlC2gAfzrPQK
vYIw5YV9Bx7j3vI6XBqCxtQ22uIcj/1lZNhHe/rThjCaej2m/Bn18w6HLzAmfX36TNSSUueFu7CC
V8ZYj9IhYRb/U/A/px6esYyKRn9bhKDU7v1PnCPHrx0PI4lgAkKRQjt2mtO4gAUdv+jtofIkDcRF
twsl47cZcrwtpUGOMNvtZFPfODBDl7DFGSyxMIYcFiCxqvNm7JJlT/T0sQ7NUUwb9td2bMt5U5B6
orIn67P8CPwtDqz24sIfrD3NStKam28f1/sOElZ5WTUSExg+poa/iHBZ/RGLyB7e9L8FCy/0HtJn
ucrVq0teZsK2axL/FNGo54o2iQETbN0QtAlGONou50bm1lWUUzE4td69SVlqX109C8qVbnRiaSlC
PKo+wdsNDZCK3Yl/F9ueUXDDZ/NcQsTgBEVX+XZPOeJp7TvJWKECRdm53f+CmvIqAm5TpHaGFNMn
huWoV4NLs1UUpMCYC9ZVRRo7woBdtuCkWw318XRSlc1m5FB0mT0jMaM3N3VWaPOO9zdcC233ULKd
froOjKCbbZ/DZE9oi/QJJGDxk0DGEDtsW4L3qg3GXeWuJVKG5kw+4CRD0+QTeNLT8WiSOA10l8Aj
MFe37e8K2ZsaOkCkBSdcl49Z+tVaN2cUg0ep7M1XtmrfF2KUllTsDXGN3EOJc+FddSgQ0IUCXQrJ
T9PIUqnmiLJFOKmgiJ61/UMEWTWqSJfbVFhjVgj6V4IlB6cSENiNpp5S5AIcyLf1ip/OHsiMQGFc
PqZ9cCsjLcZ2zWa9EmNcQISCoOpsI2u5CVqCl+ouoDjJfsINY1q1B6FcQeXcTTvn3qNDoshhsVrB
2M5WcXxG+SyMAXKqfR6KAkTXCtUvMm8bUDUmEf7AuXr7Q7hfRNdOslYmbAj6Al7bjsxlY1ChiWvC
M0Omn/uFCS4/HpNb/rMxj6FRv7xaP0fQIoFZZxLFAE0eemWCrO6qsOmun+BQ/Z8rxKJ2ax85f6NI
eNon+5Qp34Bj98WKPgP7aRQxBQp0YG9dDFBriVsfZeBCsQchwmVw7kFfdGztOUJyQXwqKXLPhsba
FAiFrTHpiGG8kTkBiMd0tyhpGPpeaiOA6ERzO5RrvBXq1tfTIJubbVdKGKijRgpcCFXXanyiU+TK
bon0JkXUY39MkJLzbwM6xtxlow/InXcTYmWaQMjTFFuu+Q43i39+LWq6UMy9I7nBiF3rBwXpPKjD
x226NjMQ9giEydwKQ/z1YL6UUvFYhguLo4fZjdLvEbfvWhL5uK2goRmASYULPxFcehcLuNC0ujs/
CqBsoRp5zaE5xaencPg32nEJnXYtxvOIRvilQNTaH3GlnYtD95lSfxp/AF5/w9pzfYE7OyaEaXXv
Q28N/+N/BwHRexj7tIE+4JV1pcwUcdL+rhifeamMKsMJXfDQk3v6+6PTT4BvQ3FbzEaxJQlRF8AQ
Qmqa/2KH0h0F0GNJye6p6dFZVa2tMHbsMSRTDbyinedVzAhjvYKTaIVXtHANbZK+QC7EMYEzaM4d
7Acxam5J3Iq41Y+xWigaTYCikGwoFihVy+L2/FPRILsZuLUkSPtTt1S8cpmZXvZn9aZsN8vMjrHI
xXWHaNJdFlX0Bto8nCE/I2eYpJTCVRGEJUFdetd0/mdtW7YTbomYLdMXXGRuR4nauKF9GtHnXWyO
9ooLgnmZ+IfgnqQwM92UuLyVT764YckAt3DjZSmi0Ug7o3ikdwMrl51EWEhKFcgj47Yu0CtUzWAU
88HABX/RC/HE/LMzECcORodqENHHeHQg/SGp5RD1KsYRghPjgUeTtxUeH2e0WarGaz3qEtrTNjF3
KXDUegys3pnA5pojnR9F8E+k/P5tHqhcoYZgoryXxUtZJw79Gl6RJKSpByZVYeNYhhEK1Kq55Qhj
mVNFtlyMi8mCI8s0o2k8QC1/yHSB3NUEqZx7VN3JUYYxpf+YWyjrVgi/o6J1jrfotEPTnkAR9FE8
8Vn7Xj7W+ikAVCneGvMd9jDyCECaO+fGFgB3Ar8RKmuW2CKu/MKYnh90UfC+zeGclJNYpItcXlor
MYXlySDo8uU3/lxabIMdW/Y0klAiOWGIREhtfAxjtpEubY5UDwraBi606k3zUF9tRAhq+PQpeLlV
7Iu8f5WpKmfjlORkmwxGGNPq5SWhzlOlLcaUiMN0WHCqmQXh0XbN25A2DlQ13pC51o4xkAyk+c8p
4wgFVFLHrhI7c7TbgtqzjmV2nctQ8041VY2JfDrZP2XkHq80fm+Ry4cIcF2zp+fBeuNH7m6OabGb
+jBOzKuxleNUum3n0Vs1kl8aNiZtr+VA7W6u41YxqrjDNq1TQAm7zMIbuoRieB72S+mdw0FxIzHQ
8clo2AtKeJRbSy/+KNU6yfTvdxCVIP+h8Zt/CGxVcxbUEW7NodfVX+2osZHvbqzTCnPlBS3k+bul
VbG8INhoSWxA2EHGHLVMWofYsYZ/M/0FAv+mPgn7KGQE8mml1PVOdUOg/dJQZFZJwemSZDi1157I
P2YaAWUXXUq/opUyajf70GntxhLw16xbfgy1CWRqyQL3rUgYA0Al08e28jpLbmhTZhLmPvEassOz
Sl0b7c/IASKdPfXDSXRaQcFc67FUX1StVkBIK1zTOt+YmbcpQmWh+1RaQMv/3HEH3kqL0IEMQH4E
owW6tQ3vZTIY6CV56aGD2ySuGfiM7D4hO2ChocGyiTuMmwxKQFOIXvNYPH5tfmJzYgimS5ZyUf0E
KGVGzTYJCApj9bsGBgj4ish1QtpCoqxjjZa9CnH9nFFTKn5aA4DWoYGw/sPEbNV5ZP+PAx/d0KRI
Ed1N9XQJyX8nLQZFHswyiRNafn4gLjPGYOQzgkTE/0rgLWYfdHSjTJC3MKJ9bSp1fH/j984QVjfU
la+ITghPPhlUNBs2z/tw1dVIbff1+MI48Gw7NowJl/fwVM+IDkw8smqtg1mrqeNoHAtVb4yDa984
GmkKF8mOmSycMpc0ye364ld3DPSaqM3+0FW5IfFbh+kwwQeZHBjw+Mgkqv6st+R03HRthjnsihaU
ssdhGwFtglEwBmWAiRogjxYTAXr8VezfmaSBGknCdXPfuc0qV5TCZDDSxkD15SNmGNP5v5w2jG+c
X4I8TXJioiCNlE2uAv8lQjeUJNNsGEJZEUAATJgTyDmhNAzfIqhrVwoi/Kj2kf5IWvD7RJCWFuZd
JkxeS63yVS0VuiDX7/P+BNtix4KUdgiBnFgkurLl4240YqCUNSwQ/qNGeBBMhhMZlPRZkNlLFiL5
NSoMrY2RZvm/pbCAQJ9Xn4tn0YHnEoKDb4+3VqHQE784ZAn2nrbhWsdXesgVOF2MYDHawZLRGRLX
meNUB2tqUJrxNmb8IJERKE7z+RqtQNVIsAhNm8JF+7jz4ii1u2gZGI8NvSWJCgU+U3RGxuhYPxRB
4aVJPk0R/oVYO5IA0yPD46X8vzloU6nhWxHunT6JN2SS9VRLVjVJsO3EOzBKCdDp30Gx94HcWtdr
qdYe42r6G9o9FZ2Od2ED7btp9vEYFyoMD9qIvATALl1w6vCFGNiDRGdDLXoQE8rvuJHqhfihxxPC
wEzsEP/6j5nk/VvpweE3r6tGWeJ1HgR1+AbOjal15YisP5SbjpMsOd1SVZr43+8pOYZo4GLG21b6
qnWpshJzEt3arUfar5vz9lFn3DB8ArSY/2tDHSeaBi4z8/fatNW/n1IjkEgIZWm8CsHvwOVin1q0
KjkndW7k54g4fYARY74XygBf+AYmfzQVQeNoBKiP9z100gSa0wR1+KmNm1Ir0wKT/xFdZhZI3Nbm
SnyNKyKOkABhVPczqdeIJPDtymqhM132t8U0hcPTttRs8VZt7DK8Jg214Wo1kveWjQzxg6zejbXt
tnEWe0fF5VJeVO9xHBEkWIOHK/mNvQQr+wa9b4lFH8TvyliZBDPTXAJdUIFwaFabfFGiYQVQ9b5C
s2G1L0oSVICfFQBjgbrxNDd7UoYajiwWKnOCCTifUYyh4Z0ccf4UODNnZULdk+30fkJd2j2t+oNR
V/Znw/xls6KYWe2OveKACPgkC7KoNWNts+wqgXNdZCWmbHnigz+CWHosNk/3T68VJ5n6RlD/JBhY
xis5qc4yk3gtZiWCSaefTV3hb4Um62Qwl4tGp2ksQWAuo4fSrMBhGD+s5L9DC2H9IRQeGnZ3ViqN
b0W4xFUGb2yBAlXboMqtXr2szMFKEaNvcLC07sRPyLcTJlKUh0B0WC8r7pEJ3+NgK7WuRF5iBLqc
TB4XTUqtKx3IskcOgOv7xF2FUY8HDeBBi3p4SH6hJmr5Jg66XW9x3WhdbaZqn4yRmgrswRxvYKK5
VQTLb4KzUa3/zk5jG2EqY08qivbNMU9XD9DCuOkiFR2lt1NLiBn9gZSnmcnL1EHwiRKRdQHYsQJR
jOpvOfusa5KLOWQF4fXY8+Ik36OHc4U9nRr+KFE+ffWzOf5pxM4QZ3MVZk0xePN48c7blSJnRbMu
MmCniB02PYhd1ZFGBzz4m8Jcze0riB2sqGQzNo3qU25U4+tCohDPe7/wSuljRExtrkaHeasa9m4n
QdRFH0xH2bQjnfnTxMQ2GrdRdhPpDc0XIyK5mg2T/KgZzXIbvHhI2/7jbnbqsqUK//Fh4okUMzzE
/r6WNNgmb3kh26q3yeYjeUe9LesYsAKTViYG6XKusZ0cCXbAYBXN1xomFltsLXd+VIeHj9NnxNKA
a+Y9NWaF16zop7szZTSwR00GYp+2+jOfcWNcluQA7RX728Tl5DGrIm+Rhj1ff95m60VwbVpr/j0h
XcU9EoVLGMlz5+8PM5KYyrGcdAtEIFyJT3mpfLj8x2M0eGOeXGye0vUv1lm/1GsVOAT/W4t16dJY
4dAa1c1kkrBYJtaytoYPKAwIYzFiqEAwYPWKfDgXHCR9X20HGSDMUx9tFrCCWpDOpF9vvJL65HEf
GNv7uLs834WxtHboZGj8qOoT4pvJkSnI5/MN06Q9u/+BEQ2TvxpbIeRKogQgCBgDpi3x4OX0zIRZ
WSpKwvRtADbyKnxhb/2IGnYlMuKXg5cnjJF8Fskh6AHMTvW2u/7bZOtqCy92EsTFOiEvoKUXTJdf
YrELNTRVm4leePNBlzmQhOaV4Sz8a+nPBDwDT7w9AtMnS/SwU08OJ16Fph8EKBZowIXX9hunB58x
IaDOTsRYmPkRoqvxETWxhw0XVbh6sK11HI1MAI6Jn6A5awwpAASL/Z8f74jLVjjLH7X2i4GA0TBg
efr8Nljux54MQFU94eDB5ksD3ifX5JELQbiyebHDwEpD37gGOpl7ymuly+SV+ndfwTnk+5CxM/8E
/ad4m8nWN+g5J9ZSovb6XlbEGP96nyQzH9+kIYVf2HMVwwoG65rE6m4K1QzKoe8B6BAKW4/pB5Km
Lzq7dpxuIOXSv41bcRs+8YdvtStZURWWNDfWxbVg9Tblc52BziDqLP/ZBJ1rNM+tTUoKtK0SmxXM
LxsYqMwCFCJYjcPNB3KMC0lrmzuYAwXIZdV6ArJHeu0j9IhfZNc6dmo5lFAmyLKMjiHWC+kAmM5Z
Ntz2wqDErgNHvSp1TgF6+LUpps12/TPEW3VbB2TCMCygIsZFKwWBFDTZp471tLWxkBmoJlzipjlS
f1mFeCT2nYkPpVnvkAeI87l2NuCwOs0FAtDfK3BHyVspC2Q4L4wUD6ELgBp6x/puANDvK4AzXeFJ
0nWX+1sX0Cw/DBoQWSTIXh6OUWE+GNyVsmI0N2ur0ThollNJEImadBVxz628gMa0NDm52PsAkEUe
nz1E8WG2nuI447RHhQvMIjVSTE5OilOGtEdOXwtr4ZRutMBx7tHIFEAJzw1zmiZC1NbcfIqcq97X
Fr8MQS+M3poQbi/CZSxvw+yOhPgp7vvshtyyyDxaJA1YCtu+OvFDxHZn/e8pvDJh8/R7x0exMYko
h2KZMxhUfs2KDCXBPSqhtFFM7+8bB9RDtQTiV1cnw1+D3yndpM/zZpxkbKRcZJ4Gtma2Wgpq3ce2
UBPbiI/UF2UOYd3ftRZsXJo97wNAU3pLxmm9r4ZZi2mVgeB/vd5z5Yum6Oaa6biMGkQaHQTb5LnE
T9WAFyVq8uS+BK6tB1zxZ95lFFZqzOLVA9oPUpwVpY0cjK6rW6EpXiNlgimlO4LRL1m3Qj6DeNy0
DOBdvO8xOdxtgPpsoJRN5zqAxcZpqFdD+dZvcc/VhpcwvaGSrOub8KcPhbhC8SvK/Rs1C1PoZJ9p
NpB8TgOwFN0ygYmRNVd9X75/d3OavrE9hnhuJIAzgezsxfdVFTi8qlRAMIhpcpPqe1HeYTTWxFJV
voAEZuB6+x3UlR23Wx56AU1w2s7XxlCNxGTDqXRER+roZnpGktDdCGkFMsxsbujHgkWEpKJyXNDc
nJJ5cfj22WSZlh3M0xHGnXZY6EgeLFOctR50bz/uK8MhPxzBnkBlWmfoXODYY+GAF+KPshC5SVqT
WIT80A+9Ash7C2pvIEt9C8bKenE0klLuEvKGHgxC3WK0cKuBvi1L1q7Oy5wenj/syOxeQXH2tH4T
+L+CFBXyQr8qCog5GnauewqkDyZBjif2faGswP9wx1nZVcKOHdFwpjyuBEz/1vGkvD1Z5ZTBVDhJ
hyxT7iBC+XCpFjlPo6pggw8UlpNzl75l2irca113moyi6lvfjgO742yu+te7m9kQDezLY+XTY7rI
TzLuNS6rzn5U6jEKJpVPqLYSESdloo6SP29RN1PTh5jvFu9O5Mh2cCTgTG6W19R0mgvbasG180fJ
YPiOANk2sot8wHTXJQ67N2EGl37aP5Rcofvdy2HezJYFvneLoereDZBhVT2phwfIa2D95vXdYhGi
5Yw7t2CuaemWdV71HVNBxRgbs1P4lS/hjSt3BLJdijmqj+7LG0GPtkU1UhDYmV8ZHWO6TYgM8Ik3
0DlxvW/OiMDoGk7fHuyTfTbpt5M8LV7BKGVmX6qepj/27MJHvAeyMLGWv5clAWSLCSdpuI7dH/hd
OAS9bFkikthwa+krbqoGPk8lbMc/C2X4kzAUVjBFWYh5hO4j/kGGCiEzvsaNLm43ucFRks/tK387
tsQYymT2DZaFtc5jM3YvGvMGHPHuhTG0hYQxR1lejmJEzKia2wZQm5oq0/a/CHn+WWuJj+eIAJlv
7GDWjzGBDXzbiLSDVsQSaGzSB0jwMfcbmAlcS4V2FwlAjlM9EI4b7Jg1cWq2ZAYJtwlN1YcLCFkU
HyvFY6/l+Iu+Oiv086oErWUIvg97ijNevej8d/Sx4WKsHViqRhO4lF7/jtmWNvtpTN4OC0C8B5HE
rS7eVBpT5pYgMF8xBDelqV/2lWT+/8GuanheqJls/I8SYk8IhFu24PxkVeNu3GTtaVq7yVwly+ya
jZGr2OC9+ofsFPklf2l1L7PQ+D0UvYZlGlGYN8PK3SXV3h4tDZzpeyExYgCDdGt+Iab96TtzfdKC
sDm6qo+8HafmlxG6o1S+TRDnzd/j1JRgyYAUuqtt15hv/aeyLC4sqI92f9OVZZBuhXlc5TmHtZF3
qsZi68LGtdZ0pdhaq84+O1r5WDEB6yHDsF9xvcrRiy/HL1EVX5hyvUi3Ibj8Jdb46zho7nwSrlcr
8DBCnlxy9aY+YmavdyguwpGAgsSVWmOC1OnDdvo5hFn8agzY+4RAOy/Q0TQc23GOxVlYRrR50W9K
DzoCnSUpa7JlJmqnPYlCidjL/IXD4tGcKgpud6+l3jpm8CI7kuu2uxThPXBG5OonFsgOK2XLSrBW
Quosc6hoIoAH2ubvpc3ueLK/ODLfN6o6jw5Vpu4EiBfM2WBbU70KsqLjCvj1r898vN2m5NQO37pt
djYsi7Q6PAv4563WfUIGiJN6K5Elq2W1cSAAgNVUADzUTgHFhu6+1Er0zE5z0nPnQY4+G/ToHI5p
lbL2nrEuTkb5xIdUlvg3hMTJhUvv2WsGc4aU+WrlkIGZ7mSD3gtNHSFykjNbesm0wjneE2MVqEH0
9bolXUYghGGYZrms6zZ1k7A9fvDgs9cdxakap+LI23nctSlMS0Resa5JH0yUeGny4C5Qq/yAlSni
I5yXeovIPnqenk7WbWXH0k5tDjKsh7nf2ncaNZhR+84Lx68m1Q7qL3X+6fRJ/jeoUbIMpsSu3y9Q
w8ocmlloyfaLO0BKgnN418OcsAGRj73U10YMyRXLGP8X9XQbMCG21GFwEy40tVmy6WrhmCXwRGXm
rPjyi+R5IrDbs3mSAd9VXvCgqRvFDiNYEdfMZY9Pmo85Q+W36hUMXWoz65eagIyUQCeQaFtyMZOW
B+3Mk1e16acIaA5kuwx9rTlum9TATd5VzisNE9UsxnOevrO/xcxxMPOA2BZlWUIeZAeimfxD0kiq
2QNTcOm/hWdKVa7q7GvFaH15QZYF+wOdWIaUq2+wOWAmS28chTdlhlUlG/tqSIIVuu+DZBfUyZtl
5gfYkmjnZiElIEwzWYxLYm1RZGNDaNTqjVFcQFnbGFf4TEx/SZtptbq1puYvUPai9g6DeMQEkIsZ
6X+05jtZcpjOBIvfTD/9cho2Z61OMBDK6gAL3VpShSu8F1xbudG0cir9trpownbqY4+rFigaCkX6
fc4NBy3QmpC52HyMoQ58fRqDQU7ACwxTKKBG3MHWunAee9kS9ojmHA4sCSBsz5Gal9F8IsCzRIjN
61evCIJZDYnwmc7a3kFg3olv0u09js+y/LsqBaCvrOv78JCxlrCqtH6bPOwd+cMuzUXM5JEl9lzw
nvagqxc4CVykvOfNIl2kB0TtHd3JoJ/VvY0G+F9oJ2SQx7215HzBSrbXfML2CPWr1o6Ox+IjvW/9
nE6CfPhaM3DuqXcw7hAJ/s327bx+/wd9H7XOB+t+mmhTz1r0AZ09tHoqTpwDkpTdb9nMg2/RgM7c
gmLd/nJzmb2v2lKQqA1Ifnn+ccMdUy5wsrmhgopFFhxUcBQ7Dw8GXCBHVHDnE7oBcaDI4Rxz15Qp
hV+XRHE7fUz2d7FfAxRyU1/OwobxMSzd9dDfynTEijGMLzNQkmCUwF5nOw+7VHI9hTj3gCWtV/Om
BguH+mNvZvQyabDbEclgkzNZfazrIcPM5BIBcH0ZGu0/ezKJsg76NGmOMb1u928l7zIY9LnBgDiD
Dz14K0371dnnYVa8g5QGN8krwW0MVVd+OL3XaOSQPB1js+NyIhs0Tqlgvv5uNh+9Jyn7cJx2JP0Q
qi3IH9E+QlkqogorgQVHqLadYGLhoiPcvx8JEz2VT0V8KkkL0APnBDzLd0GrOkSxA8EDo+ghaHpb
4bFRbZPzG6n8+QmsiiI+ZPSkbGaP69VmtPuXZiltQwZTknqkSAfz8hqXn7WjBubBMmwZWv3e1hot
DqEMmYMGx6Rik2Y2cvz020pJqvLJYEN3fTchlC4P54N6CAzdOITM40/AFSs2qV9LffA3A5BN4FHO
iM4tq3N6hLaTJ/EsaSK8mT7E/TpM5nIT3o0nu7oEQn6G9MNpmI1Pghr8+4mhkKOR8qf20zRiO4Mu
nl1w0iGPwVrMJjj7qHqDigzna5mNQxHSMHqKDOhWr/II3hf2IqMxImdEOpWkWIA3U5iyR+NDvUJf
OODIlKBjDKtYkT+yoA2C/Nr4SuHGJfgv93y8IXvbpCpW0bbxHmsJeZRT+SqMz3zaJMbyR6Ca7x30
HknDIvn0F/VElD8BViphWeCBQbOX3/pvg1izYItsCW7QgH4z2A7aUo5+fnNIFWvpiGpDftlk0ApA
lv7Eh99xuQr6sS0kKxPWFlSadw09dDtojzMdbRgIa7tvZ9zTJ8ErzW7JuH1iUOp22k76LAff5Uxc
x7ikW6/cdrE1iymds2yGo5dr4cB0IC/nDudTT7tI8fEIc2m2f/2C3/fqF7qIY6MwbHzVnpoamA5O
h3QWtXlZg4KOI17sVilg6Rxd6sX+Ea6RdVFM/d/vDhGiz0iI7cyEOaull30ejzH5Si2XvRbPGL0O
wQc18ysgUEmVQRYlyXFWttekfQGkfzK/CQpYsk4QRXph5eLKENKSc2UQPvThAeR1nSLzxHPd54rT
AgGdf5T3FIYPUwUDrAtg0F/hhe2E76OvDVMUP80cEdW9aP54mTn7v2dYU2fHIXVzA0m6jqDVKQG4
b7D1gz4XD9AbzF1UbzodREMu4Ax3a/HWXxio4k601evICcbOdcRMsJYfGJbzRkncvdlqaKndzpcM
pmOQaH59WrGuddsAMpkEaHpQEZ/hlwERN0e4qSixHfntfj2Cl5V6TZFLLoHGfiXo+SyXJFK9Bm8j
o5qBz//DOqegspFty7T/7RrvcSzTebplv7lMpraTfgjB0PlHIXMHTakReKGdjH0rSbS5yEQunasg
6BhjGXBzb4HQCEY96JneRfOWmjnFKdLRtvCB7AB8iJLXaQ+HmBXyYD3rF20lW/oJ+wfnjS3qs4YT
x6RsZ5GYFR6uwcuXVZbFkmNZpIqj18My5zoo2lCMmHlzraAvGKAVdw9evbSmknOV59naOFFoxMxr
IAUXTYjgcUvYB0EpGHKtf7KNAiPajLj9etj8hasNkEyP2brpUj5+AJzrzZjlPbqW3k/VfU41j0fq
uCMO5bQ4u47fih7+YfKUb/uxVa9A6zGnHO+D4//5FfGgYw3VW5Imnxn7m96L3bkaSHLsRCTHn0OB
X5uO/o2MBspthZEx4s3Ydj510wWjKrT0+0PgRmGdoFzriMnKpJRHUeLlp0xsE7uKcKg/wzqNxI2H
OlcP1Yt4A+cxMC8zB4M4eJfLgn5uOx8OIPe5eU8watfMk+c/rRUN0aCNY1FB1L92e8lz+Oa+mlTH
RCmNIKQp4RkeRU64d7NIjYCXobcXYvUGqT4izEtUMh0QivmikvbsacCQz3qsKn5JmuzURIdobM5Y
ZMxHzEWNGAR2S2Fkm03PookFlWszKfI7thnx9QOqfpH95loveWKCgZY9TlgQ5lvg2ca4Fp9rGDwo
JgTYJNaC0GCX7V/1eXIuRaqT+0yRZ4WzhQIUmvf0afoEN0CHhKClI1LfdxJXIXIwk8kMAmFvikSZ
w5vZXSEBVH5aPTSKRg6UpY1mjsUvIfji4v6VuwMUvLKmGULZO6/sbk3sm7QCnJWqPeeAk4VDQKF9
1Foc2NO5fN7Yg58RvAZu50+ljaAAyL5diDmHyJtCH6y0MrjEPSFayT9JyinMsL+Y3EhFFeZSY88V
UV4OQ17grFGYj4ODGbCxxXfa2U0ZADj7pGi2y5tLd1iLm2QvcvGECQHmWuwwzPTsKZmJuqEXxihK
5Z+GaqcXCbywcKRWO/AyT9ALTOsfpY2Fqi8EB0oW38VXp+Z6Jj81yVT6hLao+vCI7DZem6nY8K1l
MuxIPeJ6z5MgcpGFMIT57ZNj57R077UkIk0rqjE96KcXNaeIuO/RvgM4htr9Cz9Z9eyb2VT7jNot
eOY9f4m3HwhADnGz7ZmZopZZU2n1g0UkCboAvGnFgmS8Vn5F45lVQjNHp3oSY+/YvnBAoeKC315T
XPxM95SmWh5Pdz525unjjIv8aLAd1iVYhcxDHaEcqQcgy8mg8ohHfZ2SNTzv7sHrZlu5Czdh4WcW
Vxfa6JI626wUZ/mTP/V0dvxNL6qj41KwPM97TOgIzCCExYkh3If0BT90XZmw/UMyhCgpDSC318C8
hdVShC9m/30eZ2eMdYpnSKdpUspT5LS7Sgl+WMYC6R5ytOmSYtlowxsLVEFjoN+E0Met1qpjZYgL
RqmcjuTA6gk7+SLcn9TRhB6UXEQibKTvhfqUALVDI75Go8cYtczTP7cq2y75hUrrKN6FkIvmDWBv
1EZQkBIeRfDfX91KAnXPdL9cAW4XHlXEktgx5EUYCeWrRh+A44BQYmnIaYa90/Kmvlxg5WDYbojd
Qo/efL8PUl+X7Ts0yKE2s3QasVssIqdCbVnXTK3A+Afk1QTBv72HrmX2tay8446astoZVbkM4QtS
tSgfo1n2JLPHW7OeNDwipUFARBStvcO5BMKf9YRP+dLzqWD/F+/KX0Ie4Kz8Tf0F5hEp1vPeRioq
C8li2CxDVf6PABh3hKny2z2u7yBIKoRFY/gX8+OcyiTPMmQzFcSyNr+RswxbmKSalg8sw+AFLoK6
VirEC1sPbqXN7qNkWqPwVxikgnrzri+by4sD+kHmP74TWXZKxRHz7WCDe+9XQbWfpNWc3i/l4rX6
qwuJZ6XpHTgq0PyeFtZqA3ypG+nTqNMS8fKH+d3Bdud/I1wZokMI8zswwfS4cjkVhdtqXaJNGvOr
Tl6IcrqIhHi502PNeL2Xo8JFMwdHOYFHP6QmwzmWnGM0jmfZYoKE5N5vpDuNdZ2mtDinGMIXcKJg
x19qEFYYk9qktqQlWgQ4wcvjPI/lKVFa0MeLfJgu75qZ2YDWM5RqWLJ0MPjeWalduTKX0//jpImb
4kvwWjaux/1SEkKDYflRA/DdRtykMBejECo5YfoSOXq+2Gy1TzrCuN374ee/rnf7JOtnG+iL2MEL
bFvsVu+ViFNuRLtTfI+gStNU2vzVTgXBQ5uldmWdr0Rg+NkgUdbWMWOHE3dwXKLTOlcQ5j2oFwJJ
D4l6dbTc/BC3hIfT+WzmhTzrPmUqjgrUiSMt8AgpRcC/IeNHq/YIwAUh6KlyvY5ML1uJg8KkzxAK
id/vGAq1jMoCiFZFyluYoNNIWSrIX+wonABHOAHlKj469zziYB/hdqb3wq5SPPRG6iFUkS2I4NSG
K/w387SgprwXRgGTCrqpQoE44KsLyRTrU7l0KeGz6L60/j7Rq8aTQ6KTcYx2EdFE4Q4H2cvDycWp
bEcEEKjIsXIW0md+8V+6gK2FL9QY0PuzlyDsiMvr//PGMF9FbdEAcCKpAjhpORjZaGqdaXyr4iv1
dirkOQ2GPxXee3hCdnQh1gwCPjdYsixyTgDbTGTrbE0YSIpxliZRY2jGz5W7k2UnetJ06Onqv9d+
PbW6X9bSbLlV9nPkbxnKVeHRLDV4DuzJUdLpycZisZAQtm2XCyuZPBm8L0DBlqZHpDQ1m+g0Zr6r
JJFPug7z0jyE1rs8OaRqeB8z2RmiZetn0RKISIgykVcFP91S4WeHP0ziHOf8mGBe4DbrGSqllyj5
pizUjLUHGWBxyW7pG12/fI6sTkAAwKavKyPruu1NEEasaY00nh30stCQqP9YfWMNEkcXEOYBacfv
fnhlaezVFetAWj7OyPUypfqoYhaZJgJgjq4JrzxV15wlMbHgF3xB0/7nemA5QLyH3sAmO+3S2zKX
rlZa44u/tmCJv1PGtNIO1KzuY5g5tbmA0C7aGEup3j/YUg8GRVmIBhHDXcKZebNjV0zCZ3DyfTZA
9MvtYC5Znod5qFAC2YZdenjxZGhaqiBhfJRgOBm7qGxVFbnHVKkm8tD2riVnqqHtU4IEho42oeE5
L7tXVu0lboKgvMaggk8Z7GPbtfCag5CYhxIMQ69BlQpw3jLVnWb42VokdaB/rNQTZWIBp2FkiuQv
dtNb1/RoxvWqS38+bjddE2FZ5FRg0ZmXCSzQqHibwJOTiYluZK2xkETXe3a67dGIm3Q49w2Tclqs
JDVnM5BQMNq+aQr40Sz2YP5o4lHvx639zjp9kj6D9eTqvD8Ut2IVY8HshehEU6ukqMqixMK7X0oO
tzpglu+Z0yf1JZqMJaEoD2UGw+IIkne8jQufhEtSahJu6W4W4rS46iS2ei4DNKVqggdlHAawPBUp
Z+m2RLrDBwlyJM32dC9md0leeFGqHn+ZjqGy9dpE9DW+Z5athG1MJYx0gH/NdcZFFCPveEByfR0d
pIMj/kvGvQwJUZB4Xqq+il/+HTXA2hIoZSzjIDe1l/fTu7Uxd4lJWSbaveMbQ92CVFsJ6+dNfJ5B
xqYoYzGGV4vr8/+kuG9RF9S2gFikl+OLdoz07NGiNga2EKe6/f6c1KK4dgXw4sfwa/lOj2OrAbi1
PNcRRgG5qxVFQOmlTkEqwS/ix37MEvJY++9yT+CRo9FBO1+pZ9271yG3f10dgm8+2bpuk6mHjZao
ov05iqqL+HlRYBzGXmOhrA9+TNKplxsqfkQzqRMgESHkFPWUzHBXdtOc3oAueT9uFkgxQwIIoVZq
yu7hSQmiQzx/gAv7ppmeXKAtHdGpNf6HyHQp+mOtCa2vmRuv8EruKdkxjrx4lrqaT/HUYYu54RTb
TimYfdvxIPC9WddD0hOAjnTuy/WUVpicqvUKXzovHYHMew88whEv3OOjfoJ19TjQsNQOfVOHl2c5
KMEkWe4fg1gMbzBviBJcoRKk5LgXLyvDZbwYz8Rnce6XJsP2/QreVelwpF+9/579v2/HV/S6GAXV
gsnrWJEFb1T+DKESp4gOGj2jDVkBxVrgoNL5ZKFv+eY/RdSUtJrfPvcKBE41djFG74BRRM535K5E
CtThusbYY/Y3Bf3SVaVfNTHIROjVUYeF+/0RpupU5szLTZkUzbmzIFlO7s9P5BeAGi9wsh7L0v3f
idcfZenhQJNN7kcdqyQ70XsXxAF0rtE8zmbke90q6/qlwUqOwrbi1DerPSNzka63eFwRa1NVbV5D
O8ohResmkU1x6faVxxYaJcejtkAGtCEWww0qL1Jx2Z8bw9aB2dZ/D/Hr53kiEU8y/ns99ZdNi0qK
S+/NYZWoNd0lodODNG5WZLrfRHeOcCq36UxrnObX/WhdC6LhHZyvANFtljY7UQkCswA+R+MlpS6R
5PCpN3yoYA8sBQtJdujFF1FU2ZfHvYQKpwpCq3C/Bh2xdoY1cK3O3HR+WFjL8t7o3joIamJBEzfG
cHHFXisVsgowpYDUkVbTElAJfimSYDRrELo6rB7m1NmM8vlH3VdoeKRLBq5CIkiJ54/ToguyFo4E
Z18QFg+7skGBlAH0+/o7eIoALPLte7oDoVJkEHpFGeI8O4HnwdUzb4RTEPaKtBpffAcpn3Xcu9KN
C/fC2j/Pg05irXRzva8adu2po3/4qpOFXBHL3p8FiK4bL9Qvo3Zvor9qRCWAVTwLeWA7rYje67MO
QGKkvmCROmtDa7aDNUmOiKnbv5XWrVOzOnKRtsklnL+gA8kasvjbg7Ky+PmVoClkw9vTBv1kTW+3
WvUa3hFJ6GnWxS9RXp9WiJuQfG5xqjlue7xzfxSf8/m+/aFR19bjwGUCSklbgq8CIsi6LKY1zPYl
Uq5dtx/swtZGWC/hDDo+zSn2RAMmpEugdFZfOQz+mqU/0m7/26+bd/GOshC01xHIRkzu88yb0mqH
/EiQMELNQhibZi5rZ3A0wp5lmk9je/ARICX1P9RP5zmS+isKE5mKwS82KbZsSCYyzNUcltDK/QRG
OnZqHpMTRCcriOpiYjvnMxZnjgPheAnZALvGz4lmeUgm44uHCzijTmX2VoDd/kfgVTKjxSBe8Yad
rF4rwJVXkPed/4PTy29BR1GrIDWxmKLh1MdoOgcRVXIeWFSs1wtsPA3OWMqaQwdDoAyhHaP9g8kp
u5JQbMkTymUf5V9+dRFcuqFcOjJRR7V6r/C5AEHhfp8RyGsMoIMD3Ud4wewxn+ZDb/0VZNQ6aI4N
0kVqJDe7AsHCJ/DyhOLQV+3RoOFu6k5tsT3pbyzrwNxrkVjWn67U+R3jhhwCO1pfvP64EHGftP9s
A8AyWI4RRPJwpufUwNjgv6UJ1SvrXVcgWm1AOQ7CadyGSIRXUzDBzLmxyMlidXu+/dghzUy24mkW
DkZDq2+lCOsnK1NC0c6obDzSBY4FKrIIokZaJdSg6S9LVhqtvW2n8Zj4fOF4ES3Njrya6SSLqIYG
64XSFMp671J2/zZMJxfvorb3f2w6KYUtysyiXtKLsyeT58+6+QI/Fdg0o2rOfHt7ODRtxE8sV05V
LI4qD5Y1GB30S4qgwoyaYQVMIEBrs4XwQvrmeEPNLgJ327EMKPicdWz07CHjEZvQk/QIPpcT/QjU
yGMZXjhPqebMRIfc2C0VwY34Ai6dZhphXBvqK246sl4+rbKRA8QRpaZw7LAQ+U/+hK2ha0SdCrh8
ro3s10wo5HeL62gvFQ0gJIEDQ5i4hJ9kAolKcvQ/zZz2goRLEf/LZguBhe96rHn6dayi/PG2dba6
9jX8gwNiDmOjUpTixTURPnw4FFFFd3jJpjS37A7yZkY88QQsH/54OM9m367oCX9pspiU4U45rGWR
/Q6AURSOBD/367V59RqVs1iFLNx5gTLpEMtWRwp235qYbxGzp8OBb0i9yUpAE7vDxATATYscTpjw
f1PJ1JcYg5l04Bt6JL6Au2GC5/nPlys5iVdMfL82PFZTIxtvI+9uiE3Ae77mosqo22tCPjSeqLaT
2SLKFox3A9Wd98rKE3X0WUHZ1H5BFy8BBbSHKW/0Rxk1esN+WfVUyKEgMFSGqPx+4nBRCQcQsfa4
132MNoVpHd2F3q4rj4XT2eL7rp307wai6wrfR4GkodZrKnACRQ21v+WqyklyC2EJBZ7AsXKbPk78
+m0zIRObpiigZ+P85NbDyPhlYu4igXrO513UnjgDK2e8kGJgbZHstts1q/9iZXtkpnDB2wotuK6M
oreYlrqK8HlWF74KTwV9xksskt1Gc9S2rUi2Q2SQq81Vm66Lpfl7Z76lHXjRgLWdWpf9o530nJU8
p3pEEZJwz5THKfVfl3U49LgiY6qML7gQcicFymyxHx21SX3n3fUWcwW5j1glayT//yiyM3mWrjNF
8Z/9tkzTJPR4QIPWJ8pFRwTL7Jw3yTGez35TMYN/wCNSOvfNWupOFKJs60CLmJ4Gkie6TdCPdOZL
upl1D8R/k8BtFYS9B7NHPq/wjnSKttKNGK3lqy5iIa9aMVPHga8URH2OaVRRknb3lwI4oEYP2ta7
fsS0jSxDH7mvCriNVIs5qmKpfSwjdf8FOyI7OWVSvL/1FXaVuitf1kBHzP1tTBVYOmgNWllfy4Ky
Oo5rHuS9NiuicUawtjLgawRnlSMegLsM/iL+/puwXYbKzq5Wn7+njoT7WQGAgJKoFkx/JoVn1ueA
VYHJbV1+4RhAjb/b/QWZjrKBmzBdljmQxGw1kO3JYlxaLjcvApcIjHnsFeBgv3Jx6/3uvgg4kGa1
RTnS0ANxXOiYa/VqXU4lIqQmnn2PMVQK1/2U+SeUZ81gY9VkBRVd789AgezVQb4k+q3yMjhemPhW
tTzbb8XsoNsVOqWM97xqs6GuIwjqMyQo2lNi2cg9XpETQMTIIpq5YMiB5DEQrzT0SxBKx3ztwdzz
7IiCYeGEkcLd5TE3eF7IlX4soIYIHu8+ZTfN3nCn7pnzoYwmWN84be7BNNFVyLLT9O+U807iRMpI
aN1zTGn8by4FV8wBC2V5GVLTJMfP+ihQZKrc5cgo8DLMEpVisatl606UtqaNW7aF44Ubb9EDf+9b
gbQfLtUSuWBYAXU6Dxz2MciT4vKM7SBlMBHC6j0gI5G+4jlKNtOAQlrqUdj4NUsdMMAYn5kF+uDH
t3cJheSc399SifK9pSccf4G0RwWW73ovG/tA0dRRzzJo2fysInPJ3XOippGfT5lSYb6EsjOm+A1s
1UysjfYGqXezq6zY6jLE+ZFpvrm7WWGD76b3a8g2POr1VzTgngjWlHeW/SccVY/cJKKHGj3eKufV
ceQ6PelQziydC97OJvmD034B7SiEJdRMr0Jea7+weTC0EYJ8JmIOVfGMsPUa5HKK/jzYHIWy5BrW
cq2opfW9KYSZinRfNnThs8H4+EF9ym0Vhw70N2ILGuiUrQ0b6DEDF5uUReZPfY6VDj18eXMCh6Ja
vBlmGwWB4rfiZ6DNSLOW+gbX0Q2AB3vGAnW+KztD61uN0q39HypNmqHUyoLL7hpHOGJzYXeJuQRQ
aW8wEGE8LIMBDgq3ZuGkCxff0m/NCAxcjfhQHHHBbpC2BVxY1QatYTmCCGSev6saXure2mNtHIko
xA5Os0CwIT9o59u1a0ucV20kGsQEbZHJrEZcvPqPNLK2nIw4/4i9jVajV0QXK+Syd+AxG+wj9NS4
EdrLZv2STJSAm4DWUznuGhTXHQJLgpiZmx/z3qcNbY1q9JkCBGR7n8G+GQ78gLSdFW2zWd6oGrca
MRZdJnGXchXe9x/hG0pEzctmSp4MhNsFfMn+99uiZmtXm2JJciwiZahiEu3TuTLlki0Ddwme224Q
AxW4XaEoyfdE21ZvJEfqH6ovH1v8yEKFS2rRIIQ/xsuHulnYBuSUbjMy8TsuF14CmYTDWbUhlr+o
ZMUzz5hJSAeHRn5YAc2HU8iSrOX6snpBnr8EH31m//hfKtoNc9/RdfAtmlEb7WG/eMeQi+Z4TfSP
QagW2YGHT6bVMDtXMyv+Uk4yGuHYqTyTn1T//pt6P2NoiIw+0eBiUF6NtjUFrD7u15uTfAfNmdv6
FZKhkIJ1fVBdryWmz78SfWJhvmG2BDWNLJjl3paD4Mq4Y3mJnmvA618eaWxuBW9NUqlWfVv0ADZj
KPfPVp265ACAFmU8t7kFgrQb5bNVUbsOtsHVOWBODBtMuEpI4XOf20R6l+sMsmSnGtF7XsAjvU/g
wdJXpi0Pzq2ATY51jlVDESWoYPgfDmCiRi9k9Jnf2iY/4xzJYlO/LGVPHXIo1W428/8M0pAZy3kp
co9eQe7zpEL6ekaCqFBKNZovH9hEyRnhwtPjnW84G2MIbgxpUV99Jz0BEG9MZBXgEwYAYY8FBgED
widq2jR7k1LEOyqbXeBIjxktXFvyMO3l/1KY6nWNRHRPERx9cKHR0TIYMfXTRU0MFcOggleko8od
hWu1szB/eGaA0QtzFaSD6JH1p/ZMonjrn6P4TpY28vIZEHue0mIYFjxB6ghgRMBpd4AHQDNjML5U
aAYeCJfCRkZH44AqDZlnE7XQoMQIfpEPHfEDBzQOEO/BweB+lW5AqhRQ0qToknVbh1h4PN4+BcI1
KQoJnGeUtdww9mheWnX5CSBClrB0I2PWn+rXbEe2+Rgyvwmu8cwVmUMWmtvsOGwUxM/ERiMMUeAx
KPTzc6D9nCAXnKH+/zvV9d8wJYj4vfKVh7cfvDBcfKoUbiZNJ25sgcWue3vceKIGj9tMJ2idjXDe
9oLHQb7JgpbSacBppCu+ebjwO6A5FI2IrVtU6EOmHUokZL5/PoerMk3uyP8OYeoZquPjpZvpFKXg
u4+w3OI/oyxTgLsCD0SADWjRfeMONhmePGyBpho/HJHXpxVUsI4AG87F1mJ1y47DrSq6Jwf3f+Xo
AuNEglXf7ji0meLArtGlTK/4xzP9W++xclFwACzY0zoFIx1xqja16vEE5FhnC3NzF6NPuIomN7pt
kMF4v0IinkHgZ77jIVNGVR+zDFyLI9vEb7lHB4X2Dc7lIZu2JYlyVPUiXszlOX9/v9pT85haqM4m
pFtrnRuYKPUoZ1wm/UsaVdyt1sRLlchMBi9QrtdWaNDW/bcNoHsMn0pbtbIQUHRtQc3o1IhaDDvS
aEeJ+wP5+Z/9Bnn/CTSCxc00OHOw3+ZuOh+3dKDMCqmBI+vJK20vaftW6gsQa3NKxWTSFf9GJ3/h
uADzQUEVa2ML+loL+656t00jwwYK2AsPmwi4J2nt0O+vILCYh2QzhStXBE1SZMj4oD9Cx/Dthc+J
quiT31U0LpxYo9Z2UOGeSqNpFsjtrJR0uHInyspStcSwkmJEHgMBYHuB6bTW+hRMNKvwGRsdL3oG
uLfy/QnRGtyNQkpfalLXKv/NLRGbHj2koiTZu9LqSuI2mhWWcLmRVcnT2JBSMi4hz2MyeVf3aoJo
Iq1Mc6sY/okm36xBkG3FqV6h70RNcFUBWGO+RQhXQxsGnGz4up8NI6yc4orZBF63SBbcDpGMEJK0
u/TB0ngOt3IdyXdnGSTpAUsqYkEgkDRmiYVtzevS6cdmf7zCU35t8WBs7XiX88OSn6PL9to8m0JC
dl2h7NpbBhsqYwlzSs+OXDB6Jbw9jmV9jXjBQwCuTzQXrFX0uWcgK9CYQ/wLSgRxdf+cuapJtcjf
bYu9Z3mGyQmWplFTj9mZ2BTIMApF7lJo6YT/8drqOPFdpVjoQHrAMZMoBqxx2ASOas1I6nQ8AefW
Rp5PNnsXEXbIWXw73wiIk2k6qVvbWj/TCVbwGJcNGDkhuG/8ePOFcT3f0SbXPpbJ6+NHNZaRuSUJ
VLVuJ/CsBi5/aaxTDqAt0UcO3PJzF8oUJmccREDNG9lbQaf3UntM8dL1T1+W4RMeQRErzuwwAnGL
00DqF902i3tobKsJsOoccKvi2Wo4VLDksNosLnmhlzKS0RfZ7u6a3XU3udp6CvnOmdc6xpu9XP8H
MHM07/FOA/YkBUGCH+kqwgl/Kkqhqd3y8kIjZbycGUk0pIVVA8rK6ZsA1n1ivgJd7EqEG/svyYnB
Dl3Cab+5v+/bUTd0QdSGiFlxmrITmMvBrJjFa86oDaKXTX2xyIYuWjzK/Zu90b/o+SKIuPE7vy3i
MF2GMjt3HBK3nQL9YVSmVTTQ4MgR37mOb1hPe3UnmeOfG15AWl+vYqfPru+twvdOmuEeYhQiKWRj
2AbkNF9eqUIJLXKb0y123acwJ6n403fsGlxRIrAsJPjVGxcvCqOGdYfzpekoOV8NUp/bctmmSYl6
mfjjpQtX8fyZwz9ewiaOFibIaAQDKTnx1i1o1hqg00ACAHZoCLVlCCDPbigVTUrXvouZwJeCP0Hq
QJghN5w8mxnE6AXrRCWHL2er3jpErINRNTSsE5/gzgXG9/1uJNDhIY95fEiR8HNl556PEBPI5AaH
RWggFudTtQ7etcmuwtrFvaQ4X3OG+cRTC/cJSqHsva8ynwld9n31+jKAlM6klsl1LWiGbeKFrxWL
9+BaFPRbe6sVKuBmLRWbRcn8Li5GzGFDQ1rMzrzvy9Zn00zBo04A+JC/pNmwA7CFqSMPgJdjJY+u
QHkTbTmMTdhjkLCoEKsndgI8jAysXMKOrAB8Qv9b33AeLrFj/C8rbjCu35rMRnyHPrOop3uusk6f
ICepHIdFg3Us3rzzLIW4lIVFDwcio+Wd1qcqzXCAuvUDselZbHCc/zR7xd2amy0n1pHGB+t0PvBM
yCKH0P/DT7Rx3nYG0gLOaq14La/t9asM9bkH0TsyIYyDDpyDfBHpsEC7x0K/uAY2ywDcDntJi/Hg
aTF8QjI2E2khwzgC8kqU0UaR4roHvT/WTiNC+DESCoRugc2BLZO7Jcg0QbglgrjEPUDUyX+LkLH5
abPRZmyiTBcCepL1zxgXziIkCxAfoa7cxxMqmFOpCn/wSqtCA1Cj8bglIsE/PQwSVVz2JtTWd6wG
cCxn4MkrGUAha9RdB0dtdZyzM6BO5Ig7FgVVbVujZUu7o/91noJdnwJ6aa1qQzqvwRjIr8ztnlq+
vCjetijMvIucAebzE7XIT9cEf6GZ7Cc1TIOq1erUJNmXqFZWOdwP4ts4wlQzRWwNRQKqQqXnBn+V
6+O65Z90HoS73HXjUNDeQmxWVdvzGVt1eqv4rd08VHtr/hRqVMekWwNUF9qet0AqevFLuKUx7eoa
lPzBagmT+Z+WdpMQcQLXmCbC/umu8fBMbzFh142FpmWQ5VHLKalFBJBg0y5fRdsCuNUtYK2LYG6O
Zy8yQ5d/SMTllRoB/VA4dLvvkDtXL+dqL7vf7b5UFcN2yQJ97CVvSDp7yjxyIznGWy8uYAOB8wSn
kdqEUwa3OruUvWBb1Tza3daufOW7zeIsQjus0cKrEy4pvHLg2pPrKUlR3SRKSKWepYWpT6u1jUcU
Z3jjtbC/xjMg4n9Y6fGzdbifjVZ97wceo0I845WSFr20a1EwSUP0H1RUCi+XDewf7EtjXGIAtf4W
G+4zB+nIaihy1melGCjlfdi//dXivYa6/7+Honc3SLAr4hRRJ3EHFE7mYVNXecOgA2GspPzBg64g
D+9Qw7YCK0mf+W+7fKFMWUaYjMFmr4sRgLDK7p1Xo7vX93/cAP47MTUQH8EUe00Zp82oVge8y13c
t/FqHm4T5isXQ+4GB1YxJO4+4EDGQdp7d0H1gOoHRsDh4sgkBXWdPAGsW7dv2fLkWp+zC5vS5uDE
14BiVFVPDpHz1UDT4CqBhSR5djEISOWX3fFsB32RyP589wz27vDakAbrVFxJoA6Bim3ycIKzJdFd
vVT5jqRLCX9vFn2FwRPSoiqBCdHM2RXKSPkm+XopBbazGQh82GfDXZkfoehkUabLG94SabpZ6Czp
Hbz/9lLjd2CPV2Gylt9AltPcGNxzk9uqzgBA6V43k0vkjjpby+urPxI7UtIFV8m4Bp0CvZRiPL5R
11sayKWIXAtzniQaHdk08r8Daf7fEtaeAA1/7ckH6Z+UL1ZbUf+D9yE9KW+uyCeBsRLNaIJkayAD
UnJrokae6xwJrHz+HooXLbZEHigts6b1Tgo350FjHt04QQgB4ejLauBvrgstiInGRC6tOHnI9R/f
HQz52zS2Fwd8wBwDI5g27z0GrmK+eo/dyMOfXtdq37c0lbJTvmEVer74PLWMD3kd3d/wD91RS4as
T1FUVN+lo7oYaMS9YzvqTYiwGb8xdCrxodrtSl5XX+fLHt5TERtsyNXPavCyH2dW03hbJK5lG6PN
RnXLM5nm2byVf6zmi0xR5s9t1pDXUDSVuEqQynOOiUm5jVkVU7X0SccorFJ7q1IudfjTp/TYX5yE
NhZO+OhLRNYjPB3PdhuUHAR3IScu2/e83ldDiaLlCzXfZ1WE/OpZfm3JrhW2QmI7aaSyuDOoDo42
yvzyRUykabcTvCfCbSr8/Qa/vOJappF+R3MtOtXBO9v0oyKH9bjapzmY31srl3Aw75r2NCph+NcW
GIGvx7Ljq6tDhPvFACJsV0FXLH60pqIph3d5Im97UZfA3/ekJ3xhwhVKKjSAN8nlTf0VxONTtyGG
z/neH+2YEoVK1hgc11UxtwCHPO3Wcd8ZM21hXbmp5WNd0rAZh5q3g1FD8U6Ib9aJi60/KssOSuC4
8/vNNZV0Rvj1eq/5N837lDzXtsmpuhxewMvHnLBYC6SCl1vHOe9Ep4SWxCTFXhfHAYjuZUynvIOS
9nkNJ8TZi8zGyWyM6rtNI1oyDAm1SYTzmw8Iix7vvsIzD/yoSOQFolUnsWWACHU3EX+npN4vJC4g
Fy6Ce5vgGMT9S8m2FV/HNVCoBsTOqUcrAxlA3eTJEGaK8TpzR0yilvpD7whDsDOIAPrxAmh76LHZ
qeNCr6mcoNhYt+/iSmN6DeOrwP8udRqee8n/eqeyLWyev7Blg8j3GZYyFtFgQUTe8bNBIeAoH3jz
zOUByRVJ8/jF2HNRf1H8muSVCFQ5UFybeweuNUS8HcIFTaaAJeflT6xmaBiwVbpO799aKYlG1PLy
ivTFq6Zc+43xPTYYi6uSjyEYI4xxYa/RDY6Bp8Sr23k7ZKwHhlkqlnzlDzDi7DwBzhQquLJjV+5Q
SFFeo+suJewLLcdRZGp8Gss7BToYtmW4Q49gzmJQtdYxcnznMQgJ/A9RPBuwr9b2P5Q/YYBDC1I+
w/QioR0jlSxrCAttqZDZXojoobJ3sIIzMEVPn7O2rWP9OHMS1DGDVEs3sK5vz7E3Va8SjGDFBf8a
JL8RfiQV87jqzvpWyWQKGsxW3GjUHxn+bmJFMY9hbkPg6YMqeJOWv6dHLuVswKN5FtqQ7/7XrKf7
NRAsjNYZ6vx6YAyEcetyDur56y5XcDGjYGH0gM7q4G+gdgeL0uYqms3nINzwrD5NhTvfFM/yI8M4
Kk/C6PGOrHjMROifpFj8ytYezzZ+9H1Dh30DPRlRI8XMCLJuZi2+RAi89MJ0MF1Rfyc9ISIILvC7
hwyAxiczZLeyNDmgZZqIk4cjwpyrX8kXnCHvDiKoKDtNdDa3tCD+oDQtqf5bJrQJ3lLlzuGBwh0O
v7WzRu5/Pw74b6ZE5lUxcYmomJ6hNLj2GBbmouXl3bypWuDlyvQuBGLoTRdlGHEwXAMaWvNBqk6Z
tklwWyfV0jxbdcpyG3E/aWCD11cKomHcq8Uu8k0oRvZ1bp38KLjuYnSh7jS6TCo1stXmIc1msDjF
BSM2LLTtOG3oq6sfxEBTVzGU+R9X4PI1IviijkjWxle/AqhbLWQtYlWXxIoXz0HUWkxiY4H5Sa2B
lpHxj+NE8PLZ0nUsqJqzUMyKCPqqaN8guGbGSvOBJh0tP+pvZ6oN6Hj1daisA4xRaILbe/7CmTy6
g/JfhF2QKR8dD19frwG62IKYKs10K+yAqBXEealS9PtyAz2p0s7s98MWfWjVmvuFxL6MIpsc8lQK
5Pl41aqDWNEez2+esGFEwEew5wsFok3M1Lwr4WpMvfWCsLtCArQd4kK3RAUEA8laQmGbpgsDjPaS
zfMXDhOL9hEckY7WVRH58gtM8n5d0l+qTouM06WAHH2/+nh3lDitqTRN44OVASb1tLi4osrx3TY3
TZUJsJteUDyd8SqF0JRcXcNOb8lTs1j8CmwMYu+aq7LvftmNyDh0Ceaq6AyaWAmaHx9TXifp90YE
jrAtfX7rAPtQzcps2TCZtG6WEJPLII0de7MiISqyEZzSn5XENXa1oJmY2T11+urakxvLfShO7r2Z
HUWxEInHgfU1pXqEt+Z5llSafJ0ol0LE0tEmhD9EDFZq4RLS0fOpo2dNsvG2ayMU88mN1wy9EoAb
swRYXYfKLpRE9UUCBGidtM1OkUEGHnh2YHe4IbgFdwu4jriqUnOz1f3dsgynsD/z1gbmRyQ90eMQ
W9KYYE8Y8Wcomnv4vOAQWndiwsJUrXHUS4MT1veMYwixcHfVRpg1cLDElRN7qo74kwl6R2sJ7DPu
zvoXeDVatTOHRbWbXex1PyjjcPcY2UzACxYHq5C8XoPxA8kMZW8jFon/URPC5P0tfJhqmRnIF4hI
ybn46Ap6ORCMz5KpgN8ZGdBJxGAT8FXRD7QudGMw1Cxwf/3jsg3dmzTc5zBDjgFL8AtZC+X5ILBp
QC5gr20vzb5+n1W+bJTrnldMfIZx0pI2rrICirtCyIjIcs6pOW6LukDL0OuFdzJ4qAg2P4jhG+2c
HDbmrLPOlMzYOhp4KI7C9ESGxaeME24l48YSPnxDwRWcwVplWHi+vwZT4/eNRS7XY5B6fDuCXULV
A78lJOUVI69SZAbWyjKVPhuwSq6ZNbXrt+iRjY+kna2gjcU8nDVX4wZQbOAyinZSKd2BXJACc8/6
Sk1PrwwPCaGWJCAZZ27VXMbu8pXSbp4oVK0mWGnMEpPL10vkd3oBdodfL1LaBhxTiQczpEg9yo/s
re7tj3Tz+z1fhFwf1uuZ/Omjlgl4taPIFvP2/dTSfFeTrCDUNrU6hfIb7UEgs+ltvUvvWtqKsiR9
aKJvvCNNDt2VNJVOHF+8KE7dhXDBD6lJD7yIEtYJ+1ZC2o7g93hVjB886LmWgQDbjrcotcPzFowt
Hdk4jC+oPLqHNCB1Ay4nZv3nrPv3EURqBD6CN3kqHSPRBlHMuGfuC6pXylP/lFe0pCkf0HJckWlV
jQSqqLKwvGMRzBPwtC1vSaxdEKIPj15jRmWzEjU5W6/cDJa1XRQnJMPESCLFyHRMMGLAXSrK9N/n
K+vZ0Wnp6JuqkOcTjgHDmscLM+5OW8LNl7eI1M5ikm2S4D3ggF1gJ480LJ+uLGLhTKPQTers1vji
OJdb0ME6BV9RH0QoFHf18C0N+vkhvWJDKfnWfSnzVjPVALSQDoN9P60zUggrrw52GMu8JE89164/
I/1YjPN8uAGPo6UtOXgnZJBGA4YY7/bRKACTrjuV8f1Kky/H2HDEQZczB/5wla7iQyNWldx2x39F
EzxF7IvYjVySCCurjhtZ0J5BBW/ecjfDrUQ3JZiJOB30NiSlgHk0neBpKntJG3ZK1Klu91RM0TfN
lMCo7P/hxlbQBfPfrhwUqj3iSYOEZNWRRoAdg/zQZ/WTBiXRG2GxV33Xl0yAmAwqDtSltC8wm2AX
jACrGkyr+l6giwrOaxTTIULfMKnMvSbOfpGYFyal4cxqQ3u3IaYWSnNEIUJvDBFOSxm9Kbo3LdNG
vOmD3oVapX/N9aYJhTjNyqBNJfQOwyqdyLHRp9KhsR9X1vR6vEZH+dRZth6CWMXibh64oR+W9XYq
Ze+ZPLsx3zHCD09FlJ2PfXQf7vGhTe/2EYqNm7IoONlLO38oc8LWM2IErxgHcdcXwmzTWsHcgrJI
DySnPcXxcTFdM6lF0/V4SZlu25W4VuIo0aA/kncyLYh3GHJgjDVaQwG1bQPgT9V56reZ1nf7uoMc
4NDfBg0eKPUsYxgpqrV4e9JKnNIWoTsxSGYaSH5NoQ4JWm5SUb9QRXAljKXlT8XjEPlXAOAG36U6
tdT42zASMQ6SfPCRfCMrBW7STV/uZ/zGg42JUEWg+THVX1Y2vXVQzKMHWahJRnC84B1+TnHaz7Uc
O+HUm5DE2NgwIyZoxfc9rxsaIJhuUjzwOGkV2Nd60kjabGpMcJQ4tLbAegiCD7wXqmRMcnzyjh09
6qg3bf3RFD+WeUTEq+DghGhO6B/csSXbF0J/XH3SK3XoeFIAkS05cNJUL1iZdIVg19mDhDoWfIpp
RAor0wVax2nwNZ6Y9/PMXQvuiRZaNnagv11o01O0ve3syXKybYg6pJ7sY8EUDroqEOhdTO3h77jb
jz5xqTx+/Xl351CMEHeXMmFdcSQmZyvC4NT3fBox3TTnzrZWt3olwqqZTNQ3usq9pBNWkrUfbg0A
bUFdnFMIwHobtQqp7MBX3ff+4S2MBRud/4fgwwv5Jqx8PVDIfk3gR/lricj5JGtAR3K1a+cyEdUv
Xe7l6+RK1W/9u34HNVRZYa65BbyuFp/rk4/b/3pyd/KFhzV2eQx27HyotziwQ2qiBPwij07ovvTf
pv9DkmyDRHPeCVVi2I4OzAR19Nl5dnxyYkCIN6WrjmJ0gd2NFNUQGCXceyuhGr50varJC+mYpfqB
12+sQkQqg/Do1qPV5o6btxrEeeV6SAU/E0qDTKDWaJ150PE0CG1qgj4XGOzLAlm7miA8GM8KhX81
E6Oy3Fw5RMLIiC+l1Ux2Dv9tzLcgOLQ5t72Ukdzj9kc/iquzTKx5qOECIli0FtHDcBBql5Pi4gke
6xJ5A6Fltfab/95PP0Ae96ZXuTikAKsg4JDsxMcBg8hhTJySrSbcDF2ykvpwpz8Cm7xCJ8KDewVF
Qqe6z6WgC6A0w+EWMGQVREjo7s7VtseYwoLUMd3AfYYAbCA61ofbK8YsxnBm7cmuhaiilpEayFm/
evZl0XSecswcyxLvhXHdFA1mKKpocYIvTCZXiKl9Ro+jyHupK3gMaNczeP1nXopu5WNLhcK9+Gu6
RvG/8lHSkeB6DQhUBAIhCRqiGzvZDYMHzQ03l4NGvSzGMf70s9vJ6/uumu8Y7auTPZ3vN1hgmPRN
PbxoqHKr+3LWYqBUl908eA1gmK0I7q5q0NQhcYgyLow4P89/ynmlV/qASI5DRg7S955YlXNzMMPy
Y4dyPvfQ/Uokth5WpOGQ8vgde+/xix/uIRmXd7gIgyzllZJLjgY07x0vpG9TvdgfzVLd5ClM4sHz
PAtguLF64mXncOlcs1Wq1HI+aM/1yetDbsY3Vf/Y3pVmJpbUBX8CMY1rXjrNIDu6HjNBu9c9M/O0
NlotK1DQiUtnyNM7E91Lo0EpPaVazBJ7nHSC2Eqf7S61bbFeZqsBRTzsIJkVeUqoDz6UUrNmNSQB
GfdfwUGAG3UcTrwQG+LYF0qL704RPzs2H4KhIyja3rI56OWZN+veTRUZPzKF37graZBuWMjuGMrN
ZVLXic278x7aKr68KLB2jHZWONdgyscvGaRq7/lBE3Yp1rC5qyVTh6rDOmn+UYqktA9lFUQ30Mzg
9rSqzwZuTW140F07fCcugmvM8JduZYTOO5y0co85fFwkkxOKLTp6uCpvgdFUyJEXQ+HEKM+1c6W/
sFgrM8HxIXFP8A8J3T0WqL4wr++wmVQ40EqlbPYeATl44ceuzOKkK5moBrIZu6pS/WlBqdit7j1K
GlpWx30YR6m9SPNS44KOjlAIDh0YW55wb6pSxM4sHi+vkZ8HJ3sXwnOAHwYspGkRzlU1O8hWjFgn
zBckKC2HrQvCiS5sMGL69c56fs0ycxL3tCXjNg+gIAXTo2k3S2vPKIPAdwqOU2wv9Y3W5VyR8vhR
YG9oIZv5YBFjIgM0zdHsy1GCjmscBNqnl9dfnqVnt8BLtHrdTIV6H/BfnucVy6p3qP/VWnM0+nUn
yz33ZbWtdaVwQEv8ssLpA01jNIDSuQml0+Kd+12HshMjkMUeERQjOLi56RQaCDD2ok4P+9LK3sxU
7g9bA0kZR4dH+4inPReV6YOqEB+yUAqHyejHiuplKL/6b+Z4w5stQf1QsrzwqbSlYevxmxc82XH7
tcMYwUQEcL/ZktvwMGkRBL0tSiL0LosOvUPbFr8dGWZZd8cklnqQpOpfebH8TwjkEaSyH/FDfd4g
6mq1uisPdFjkaWWq2bVrwm9iCscVGLmY9vyz1N6Jgoruy7jDD8itqzdopnHQKUkcVMzSe8V837yI
VmiMakUgw6QLPtUmpDPuoVik3zn7oEUaZdCPbp78yvuhN1isnyM1G1wH6e+qa5ks0bAonFGmqphF
dk3o0CXJSKSyFgwb6iVTyUcfk26A3DzLkMLP194qlw3xmlwU6zFRaznMBdY1htWg7oOB816jmnNZ
WYbwWzRguE6uVRkRgbNcA8k8hVOpKnSvwhfHUWETrTfl+zkk4FqzwHt+vEUvM23AXKgUbOA7KlHP
uwTPtqoj0EuZ1MgQkxejBq4ECj4xdWHNzwl7DSU4mKk46ivBYPoH9J3HMqqROtHv8p0WWBK1+fNb
YQmEtseObp0Jqj3bQVc7eq2x6TS9/F1iyhV58G12cdx3a0/K4ZhzrjHbLJn4CsfrFGJ+V0VEJBmm
kH8qLjN6Ld/JJxVF0PYQf/rzVl7vaUev2y1MbSTO2Z3yRd/WP/vo6dOoX+Y12HhRORFT3JHIeBsK
aTn3JpEMPlU/7OvJm6PuShbfkUAmdVLBsvG6PEWsjoZjypSAjERRWG2bNLo9NSBv8Mgsq3+meGgs
G2PdNSmPr+Gun0x3e8mus8TkwN+odjUFjHbpaoPA1cGWw1uP8nu3t69T6dq9kMK+LqO3/zjEoUz4
UJsUGtK9E3iz6pTMlKhKVQenUnWvT9zMzlHXzfoueqV5pofuQS8JnIrSN+DttgGPtczFFd04l5G0
sWI9hVxs4xsCvO2iq5OO2w+f5x3atOESPA/zSL9PAGKAbujMJbdoF8iEqSby5HB555FQ53V5yEEP
ICeBc3Mbds0I+SMb1AFKZ6qp3AKf275WXw9J6EOppG0y7DObSzyV1wwtPajYBu4x/CMue07v4RoV
ipM2X6h8e3Ai23o/qjrxrjj+ZnfRxLW66GtuRXMyElUZlLYUc06vwvEgyPT9rFoUyYVBKBoyeeV9
nBieTPEOduaOfeoANDRTUP1Nu4fRjOpaiK97VFO+jR6CZuXd1sGm/43lEYsdENa24/cl8pYhPAIj
+xM3XxR4VukzLv/pNU/CFxJntKHlOoiLL6ZYYcoZMieldXfvbHOehSbiInSYOiVRcdV05F6BQ4Zf
lkKtwg2U5/ZXOPHDmmwmEmU8flQuaw/h0dh9RAZIzZ3YAGVMB4in4Ll3tDdV6CGMJaupYrD7eWDp
SHiYQQwonDHDKSUCPSYIiZ8qtMRPV8h+lTjEr4JKvGm/HSMSKsw8JGnt8UbgQAzjGOtd5lgi25T4
vuLSUw0hKnOeeQk4Mh6s5+QHCJpt6wnrTfKdjzPOOfTW4AE0bTydA+rjTT9StUJKZaHNCJ6dOueJ
blCNqXpa6bCI0zA7DpukBqv7cUaeea5p5y9+qniqa3RwFzfgKpSZbxmGJcO0Cz+peVJ8eekg/i1L
rTOFv2LS0nC9iDuPSSDUuL+mrIdJB4y1zdtyxWcFatNXOYb5uXfqp7hSOMmvkpZKGXtfx63EMIQs
bQY1CiqYJsObaMdqB50dQoOjLWKxUI3cajM9R+bsLJ0ACBgHI8X9VkO9bso7BYFG0xbxzcH2jLOk
cAKRD30dzCH1XC/VlV8FlT0sCW9V9LeJvqJXgva4oNvZ4fFkAuQWdvnqKshd823CvaOMyRaRBjyJ
fYIG4MY/PNnC5i1ZQHL+/lpovuzPhPNEUW+nfxDkGHni8cXMk6watTQqX0xc6s1LKeyA1iyjDc6m
KeuJljKxRy0CirSaw0xhHeijVxQV70X/6ZjW6b4Jori+zCXeddyiM/3gQfpvFnfEVfGECbjg56uC
Iz8FhstKtYaUOZfqShmucNJ8sPrsnygDRf6lbNwIkBlLfvIHd6R/2wHKiIsp0YhzA+wk/24Xu5fI
pPpQ9AEVUYnSISjE/FzNoL+Ea/DdNHU/qHfr8leDtOwK3B6ZmMwlxLVea6I9LLALoC7woODyWDlR
CXh3oeHsJIxt70icFPmQ0zWNn7VaoHuD6jF959gk/CQChWSmXUK970as19KZJEaPB0NZZAzIB33E
xJAHgLQKJAVobS8F2Jsut8tyqXU76+cFkyuwNq7rMQsh6tUbN2xdc2Ukx7aD6iVncmZwM2Wwd2Hu
wdf08NqZw3QNg795/YJyo1zspzMxvRtUA/dt7i3ZIXR5+bPtzOkxMqpHISvt340sa+CZqnffjy0C
XtgHV+7UUWLLG/E9ph6esXoA5s9y5soGd1i9M+XevONDhjjkp/VB9AUsUH9Z9woo3WWO8XhcM4Q5
mLvfIazvIOcKwDNpuvWOtjE8zUtsrI6VRDMlWY22IVxf/iixJjhgYwp0O2evOQOMZmy5pj10Byri
ECYSles2CDbIDyB5Ed1W3MCof9YxIKsCLySnPZwHYfCTPk5TK0l5MoJfS4u8mj6JAeM0xm2XAryi
DZ6QWQ6jeFeUxMK/VBbRej6pw1ZzeUFG6+c/x6m00kT5y/0cAH5BhsvNfYQqMM6GtwyIe4J1+ApI
qEdkwGseCK0UiKHhNU3Uuq9/3gBoHJDZ7nv/b0zX0KZRys/PokqExwQjXN+0Z82m1AK/G9UP4Bf3
K5DC3y7vwBnrhdSsmADRV4f3t2vco9c2A1RyeiHnzypyXJcoGyjq4GdZ9TjgTSdN9YjPiw38xbsh
1WzDDWaciIUUT1zb92yQe43d5nnPVRwUZOo1JnSA4NkaN/McBCsf+pMvKQ5yQrlbSJTeyviGBV7/
RdelSRHTQlRHyJsQM2jlk1dXD+iogBt/xZWi0f0nN0/XnULWXLEjyjPU1ovFq1/386fctBvHgx+6
NeCNEGotawSVmaS7NnyFXNN/nRi+9U09CFEyqPOUrZyn6TMArwQ/5cM/QR73LXtGS79jiJRf/dX6
T+Ta8EFqV0FpLNJ6FxvtGuVS8ltxF31HA8/HA2NUZiUCH223PzZgiwcYEIF24OI3py6TyHEJE7Ue
vXWDIYnrLPNE8O1gCQDKVLwySJHJM0zRcbcVaehBpo+8pKh2etbI5RVfbWbDp/KTYxlgJnCuJ4tr
1K+lZtEawVWuWPdlDHOvmZ09DkBZ8Ocgu+TXnzCBDg9EAlG8eDK/69o7KSgAjwIusoQ6BHaGE+Av
NxU0GMJLyAM8XqJBAVhbaclMmiRIBBTLDh5+O6sIJiDNJGJ/pJfqQCRhvr9hPj73MKf2vkfTboRo
SPR5udV/Oid6n3b7ps99Wu6lWyq3utWHbAE+QFR3R3+C5exGKzrGUq0wrBQlirK4oGcpy/ZeYVEI
6oQkvWzxO8IfLioluqA46D2MlA+voP1UTYKXRp7W6Pa6hF7rf23prnJu+x39kYefVucd3C6+cznm
SCjWg27YaSI/YU4n+JBq2dYkVWzw6G7SPUD9xQnEDYC9LNQo8jn8/cLDU50jQICPFyM3t3u5dQCV
jewT9ccYzwtaQSqIqW+l7tXO1COuHz6/E4Z869ULrNTiQED6CcE/Xyx9r8hYc3A4ZRimfED4yFJQ
3G2kk7eROi2PyOld6DzdUIUDN1g+xLgWYkZeCoavAfTkcB4nQUv/VqKm40JpcV2rxxnA46lTEzFx
oWHavyjaGA1efeOafzbep6WQjf9w7lCNGZ0NegDj4B0K87L82+RUAgxlK0ROjCStnRsB4dCajw7m
rbOJAjrN1x3dwucyueTFEcdR6zqBFlb3v6weusT4J3VIh21pb4WKYJWoNWNRE5Jc+E9ca5LlOXAS
ZtamiR42lj9u0oAECZn02h9hsROrOq2duncfnltXg1AzmSsHfRIijtziETh9TShh3O4rNID4YDUW
fNX3yCX/ntVbEzk66C2fh5oA5+xDf7UKsgbndoohspf309S8+91fHrkGhODzPa5Knu4UZVHOvbeV
D+LhAfBak2L/Y28KzzYBJPtZprd2N6fqAblg8fuXBVENbvOMcSxw31mzGrpBzYwA3v9cc8yQosas
fYj6NfMjQJNZlPbuP5XfvndxXXUH2qX3N8TqaponS1BjcsPQ8I/t7yxSGd6jYP/u6EYsrLK8xQ3+
W1YWJ4i4YHNnwtAnfaV7O6Xr9sV/PtKFQTA4FzGGVeFCIKa3KkETrimGgI8y7TtkTaher2Wg3rMM
/0aW4fzLCifXzK1SM3mbj+P9xEXV7XYyckt/bAzO76F4nj3P5O9mLhyXVlWH0Ch+WR6KBKjiCs1U
0ihkOCSiCzDB6kRdvCkG2PnwZ62cOnMfLYlRz7rx6nwndx0pd+zh2KO4VrwRgEfnHeJ5hdZlKTfw
ahMHTaoINFrKB23TOiULHTH4UQrpil63IUIIAPDtdSFNWqd/J1kKJHx04/w5COh2X0SXgBbRcHMT
di0e8nI80hgJS0GjABixhYPwDJd6hxElKvugbrk7TpBnhRDx9Hm4D4F6b/5+WgPG0mnUp26KCXrJ
3Kq4BeZBpfdJFlVFiqGbVCSAyoPaibiVcCPDKBb6pCif7AW1570ApHDBUmRGX0lg2kRy71o0azjl
qHfu1We7heA9osjKKgjk7mR/8WOOXNfJoW9WOyvkz1oG7sQIiA0ZoaDKctzevt0kJUzo1yQ9q59A
blFMo+gWcAr9Px+j29raPM3NmwJZZ1uLAQIQE2xfsVmKSDTNojbaG4JFlWo4Oo2OxjIMb6cZ2T2v
BT92b0ghDPWyy/qQ04+lp5V69XzvbkM67DjM6Juz1Dd08XpflqRor42KKMPp5NaVjh45xon0laIG
iLtai8SXzdmGFQb/OFNzFNXykhYw5mJJRyHR7Fo6UATvQsE86JVVBkg7Zc6sw3RRarDnH4gKJVNr
frBu/UEBeJ5zVNcb9js/IdDaVhrYDuoeUEniy/UlEScaYtDdjHu5geXELBF3MuRtctMaigCfbdvE
F1uXc7I5e5Qbldot7fS8V9MFT/f3LbUd6uLHcZI5rOz6gg6wRQ/DCgOvop+ZBdOatipqHNMbdheI
4uykA3vk+PQcj171ogG2pSdK+6N6Qpbp/SoiSuIPgQLdLKMn97c0MZhOQkk4RCxLxC5vcm2EPY0P
wFZdzS/50+9BjxfcCnl7bQsi5j3my/3W1Yx0Oszxw2pvS/ZMxDjt0erOBG6MOc+we4XzbxnR7p2E
AKNNucXd8DuZiTicx9dOl+zVIgUa/znNGx952D+Bn2GMfGdjwFCDi1FAA6eU4ZMey8jBYTd7GJVD
k1QkuVk/tn5V08seLw30xIzfl+QfSiMbcwFUg0X5LlGVRv5dwVsUae0wDSSPaZ+ABRBr47e7/Ioy
WW6Tnxv8S8zScyrSNN58wvH0Pof0QXqRDQd9iIju6cjo3pvkeirretafNUQi5Ux7koFNSvpUrS04
sWzNBriWWypZwl/LJs9ZnRqRUWJkKcEvVBlC9X8VGyyX2Sv7pjbLB3CqBPUXB7azobszzFrLR/O9
grswfc4Ej1DeEbsgBt+WO6UA14ylSxhGISWvT0+Hi+DFgjtxiojZL8SekvK1KT/nABrPVlP/PTCl
1LBTFCsDc//rRZmETz+i9w9Nw+nj9QtqXpRHOct/Eae62G1aebgI/mX0Nla/i8iJ/+TsYJjpCtHK
OALxtSVTKBOhIwe1EGirw+3ZdZ/sba20Bx+mKsdB8YWtr40nk/KNJ1vmj34Sti9cXA5oTrx9WbVB
pZ5ukCVmQDq0UR4oxVVOT1Of9iCJQ5j2AS8A/0zxH7Rk1gip1jk+f2HlrfAcRLKw6RNnoFxSiS3E
PPACPWUuLV+w3U6ZHZ0f08POEjgiJlaJjw3UIsqWNreyE1JepvTER3xdhr2+0AN1rPGzgabW7PSe
4ZSvi0QbPocPFgin91rfWHp1+g75aefinrKycUa45UfPQdZ0aC79oANgIZGYT3X2UOS8HMmZA992
Hzmr0Th77sDN3a1PteEWuzZPqX38bMDy8ka6bR3uW00XMNw9cgCkgpDly0Zz/VpYLLRGRhhwWx4o
lWHtm5xmBFtvMCiEwTAXohnrIDrVkhRTM0s4UrYypwwCrIP7T1bADq2BbOLxMlA7wtuGfA8b8All
9RGVH5VV8bbux55UWvYtCoY2BTfxBJSuu2zmI2UG08IgLS2NI3YijiQ1jfSFKjRV/KYqDiWbtDqO
kAFhB/KUrO92dlTDS7zFtipR6etzBuVSdZHu8mQz7pWU3TakhSDwhDW87V2gOPZhCDfLOi1LMeAh
YWjbApKK4LJBD9d0jrioiPxtgnER2RmFkgJ1EExD4ZvCrBDzLZTWRVm9R1Aqn1tfN9qUcR1MI3R6
z0gV/9+1wtR+pERvTzB3Ntmft6OglPtCzUxmyOVYxbwLpd2RzA/V+LgIZDQaMf0hqX4SvKJsNXNT
MoorYQZMwunNQqQetOviyp7JjG7EJW/fisPeePTcpoUYix5h1VDG3hujDxCCf9GvhGjksgAp46nO
53pWrkYrqWv8ysYWwPvc2G5aQIWv9uAaLRpJkosUGuMcZQDrbJb7GsSNEjocLJqvT3MYsh/jwCyd
RnQyRX0IQkuQLic9T1MRgiOrYWPU7qAj86c1m5OGlSiGVc3egpnu3sKrbKJQhVi3pR5PbkSvL+86
yUR4r23pnzSx4urfryAtzskPpI532vSqNEhcv36x8f1YHS3y0XxU82SO2ekO0QyXwxpr68vCgpgk
yyGyKIeYfYeS6W97iQfKgu4bC4mFhywXJoNjD/AQZn8O45cwpL0EqfSCxpHzbMDBwgJpwN89DgJL
X4l2uUwrZhECqzZTe5gaVBJA1Rrk8LkhND8U8b0cbzp8H7trGfDeOd3NQ8nPG6IgtdWnRDBk2aTO
TZHxtIcb6nH2GA5Jokz83vEnbDqqUQE7wRGoPHXTuX/kNsyS6PU3K/tnK+XHb7lRffmyOrgIYP7C
QJVnICDBenvrFvpUWsRfDLv2Lrt0UuQ+318G2vzxgbqpA4kJyNVC5riTKjxDf7uFKpOPzBUYYj77
1zEWSftAZ/aqe0OK6FIxsXgErOlA7zo5czvxCminY1QgW+MHO+KTTZfAI/5i2aSPJOB1E0hDx6Ml
7+mkqvxDvGwQUzt6YiXJkxWPh/bz0geDyCGDZ1t0oLauEWyTpmrkFFvdO/JSoEIIAS5wO9UQzO5x
rwrxo9psesA5kLFbo4P1wEIIL+qTlO1b9/zarT+HwixpG+w8c2FTWzMN5KBf9xtlHINYXotUccPs
tSgUu6wBhAtyxtaASZEbUc6iCc4ANTY9FLK66CyOMkXECqC5AvActrbtqwW3Hr03j7ZDxlxc76/j
MgQNFjBLhT4he8y9lJTvaEw5hE0z93aozycF1wlE070Wm3DbLVFDMfJPdPHf+pkWggC8a5fekrxN
9EmX+FOCP/CLTx4HpawdTuYGRmBZYUQyMEZrab5uyDfjXs3s6XYU1Figy104HqdI+noxUM//+jnl
esaCLFp9XYG5Ses3lnWwP1kTD+wkz3EeTDtiBxgH0HeNPvQhV8jqNSzQn6z3Vk4oTm8YGtB/oQ0k
0KyG6NcJkGUgwFp88rPlxXPdvopraMsezG2LYCMDstkPRwhw7mayAKYAHYcqzwIBGBYTU9sLcDg9
IDlP8IhCvcKOWvlI860NBILbC+iQIEV5hFBGQeAkJ+uPS7xcWZoJhSHlu3qAhQnxF1DCF3UadYIC
TmXY3ESZp4J9dOqfJIjadw7ysA6dVPdcCgL/3cqPJbqjDqzdlqtkJeD/jg+Zhge6ajN4WSohluua
hMDjGUkTi9muLNYoPdUHsvGiZgH1aelrMVbo2hDVhoXW85UT+geLYvyGLdc42RGfXKp0sRQxRsYe
nln7JVH31cewjURN+28oURwdX06KkJFiOo7BlQMaUQ3P3MkdqYI0JZ6A4Je5FCdS95T2vOLo5aC9
jevYUbmsnqymjn27zL1kxSHeCm9UZ8HpZJWZxtLdFVPmOK8wO9i0Cg2kFAy1kkhLSJEVJ+5bSxfp
KooyDGbZeV2JjorHbFHCntKojjaqwVHQC+dsHEJaL+8s5Euy+Yh65TK/6k1vi0tjVOqPeWJCbFdC
oGDFpORo9gfR3DsHm41C8EF446bJsydgSCec0xmq/Akl3Rm9maqqJyIJQEgEhiX6Oy3+vWVSFJIl
HC/R8ONnDxKnQJTtMc4qrNzJz1qP8TdZzpncnHRk0yAjkjC8kugEc1vH0PE+OPPdDmVe79mcke5B
hnPF9md3lkoZZRf4oJOJmQTl1N67cTKUlLAwdjYij+rjk18jIfT6QWSJuhHHuylml6b5G18FQL9B
U8rO0+sGqeSJsfA+iIqdyzKb5Fm8gvbftnUMaES99qZ0NO9nRzkFtjz0KdbN+ClACit1ADciTkhH
LXUsKo60Ybo/OtU0rr0UHfBqLBv4GGbhrruaH3KUszcnf5Dxf2wGUxEF0N/KKm86TAXGv30BBYIn
wkFsLfFj5NqUlBadnkLSNIRlxs31w0aqy3sjjyUmbAT50K8lPqwEuvyVTW/a0PfWHuvMaSKWvpHz
0/SwpWMbYQCz+ioIBlyyLnn8X0+GF6g4jVk541YTEg1ZoZZz6asxGmcl/H9J2IyZdKmyhQKb3xph
upUTe8MYiCmrP9Y6MF29SD/la3+dGmSK+gLIdLrascuVEGPDRKSDZ3/Gr9uviBog+G8W/Q/UEmjx
O9/eFvfOYVp5SMLT4fgFx0w5OJL3VlelIwwbtiFzqO7ZSZbIdoqatVY4OjgyA35YlmY6jIZBVb2M
6dMAjypJGtRU08DaoUff4yn9KFhA8je3HjDcufA9NFo23mUsZhxrAsb15VA1H3MyPeVCNhUInowp
PM80G3EA8Uzgb7gPZC/edCjMG/uNLxpyOJm2M3F2A402/8yJ4+imSaLA3053yDGcNrq6xEL0EsHe
903WUYrvvmu7D3iyy0dOvRNqeiTtNzb8yLNNpuhCd6HBkYfH+wub7XW+ZSsLWOWN5YgKrZTbQjfn
xcwpI+pr3P9I6WrvyPmRG5vjIBQ1P1qVYg4EIydBcwMnM3XLOPddMdpUu/G3rltSiouUPmiSr/F6
8sTUdN2IjHgLNcjP1aA9dwEX0YcvSqKLAozTFZ6rSzyBQ4X3ntNxnS9KYp3HUxlnHf1n/67x7Ea6
xSP7F0R8yXsWGFxlzfV/mKIKqF2ZkraML1K+HW++INFsCZ/xxiJ0MlRIbePopEFHB0tkczcudxoX
7XBX0YvTGxBveLM2RVJ6pbZ5ZWhBX9jrGWswmlv2IqTZdEV7qKgNvbWYLz7QQkk1UgjIw/i/5Lh1
UTyPuk1zL12ZZHd7gnKTUjdNcCXv3jxYMWrFmE/CIwDKUrpL+Euhg/uEW4RD3UCc/0QmybieEcUA
pqvBeGZ2l271bnD90d/+O3EjH2rWZ1P9E7qZbBGwQnonwCS27KjtvmTDqJoyZyvNxjdWeUB0Pv3z
Qu6PqPPeDGUnOGvqHLo9FFa+WF+vc21HGzLGkKWwL6LuruOlKTmPeJ4DoWteU3fSJQY93X7E933i
ZqPqrgBp+AuxcJFAZRfUptV3Y6v/4GVsYkbZY1rZoonCblWnU9/fGXWs9z9CNBFnY9DxCQLtVn9z
BPVBEvtKffnLBITrEMvYBnKAb170uelnqUdes5kWrB9w4MQynIMm3IWy6jbyeLu9Gf56Kgguwmxe
kUSHXPbJeAcFFQLNYA0nspGg3TPxAjse++lLhsU8pjOzUoNBONndVg6PowRTiNyxCi65R4MeRqRz
MLRC2fe8BlUVePTqSfNHH3K5CSYgBN6cQ7Qw3qNBwZMvItOIErptWCpm1oFTn082PsEc1MT66Xs9
b02xLSpNjWdgcB/cmy5L5g/fD0RvRfVwUi/zNe1zSNcUNu+dL85HARC59DjVoplhD7iSLyC7IwYC
wdAuU+GzX8RW8EUAcszJfs7W8L0/5jnV0vJ4DSBs34xeMOYKk+9afYymcuvlIdmnUdoMYe+XltO6
8L+06BfeAGHaqUbEZSVThPi4bSawkqP7KhMfsUVp6B3whtNuOF40NusoY6geXB1dEyY+QRPGv0HS
H1Rq6RQWMy5pWiwYTmX60RF7sR45cp8+VaBv80y336NFlZBTu9S8WFk3Jh2XkJA5/ENtgl2mC77d
O1i9p3WoBS5pXFt6M3bMKdtbGp+10F/K1cHIyw2q+QeddUBtpvGhcKv0M7HkFbfeEDlNlvyMQxHz
cG63sIV/g3CICPK8t9Fh2HErbEvSL/Lb1D+YFWCkTKme4JZlOuc9K7OT9Elep0NbjeYaniM8CXic
rGLCrzZXvB5ryITuwq2WNDWMvvkFBHvBseJBfn0dnsoEUaon8R6j7KyaJPvyyYfZN01SyrvTupAE
JFzg5T54OObatAA8ocavBrNwk6Af944wP/pAPD6HyQopvr9iliQkKEJgG6szSR4IUDsDpmDIgoPx
Ln6hxM5dgiaWDZTscCu6E/sMhDSXynQT71gSNZah3xO2W8cQJbG4NSdKY62yvyQW1pYn0F5t37CZ
+aoDjYN8jtiq3Z69+7SbHXWczGf9spt8zHCHgkEOqR8FoJA4PIa8hC1munH7KZhDMKC8cvB/nm1s
zAp0w4+KVBoNqY+CgJtKfOMJBflkyKdEXiqLBVavRSrE200wdEkRZPxIGhDBui0B5Pqb7+Bihshl
T+LmJbB7NYY85GqpVzxAEMJ/WM9FL3YuKRrcNaE+/wqJ66696UZugOW4+zoSKMpr1WGSN3xhV/Wb
iX1b2IfGJLyvy2Kdt1ZuAY9gSVzZqutEg1Lf1coKC1HWdTivS16HWBB2VMbhQDzfx9ChBTevXmOV
AUkRJ4vK9/9EWsm7Ey1fN9+MhIA5fCCKZT82QHZ11paXaaZ51M8m8sJX2jNjHesmpeaPnoi3Jo+7
i93eaNvvVBNUQpl4aiF9AX0sK/hQQ4dKbpmhlD4oGHlAQ8hSE7Wm38L1W7BC2MAfEur1k28GMVaM
njCWD0kmPMl2okhClcjWe+IDD7J/9oC3TEdECdy0Kjgzf14lhV+hHijYzZfVifuLaenHVMq0jqjR
7FL22b1YNSvPAGBlusZx/rooP7u7Mo1S332S+sxl74b+d7DehvcMlr3xgmWIrZQfeg1H1oFJfPK6
985TC8HyIRlovQLv6+o0XwZUlMAgo7N4t76hoZ2oDJf4W3QStjDl2pi2d1ViYWlCb836GLp94zUW
VWKNSGricL8ayLbSXGwAQL3yT6A39brJatboOgi8JQ4LR3mqHWxkb8xT7sYRGVdDyxDaW2lVDWE8
GvUOkjzSgOLaZHIZ5zHm7FTK0h0TtrOqw2Vc4/JIl1CsVyJUeBZu7z4Hlm1mYdzcg3IjGFsZsZLf
vwoTjwYJdRJIjc42oXE1vDUMJrGk2fvdNw4HDd8LHX6zq/hvEcE5o0ibTGe2G6PqUSPlMAPDkw2+
uSeK1hcL9a3fcbpCN4lWEUaMc+385Q1BEbm7opuh3tkktFpuWohhWzc9+5nUnLP9ju7ztgYoYb9x
T6tZh0OmqbgCRHTlpJQhDIxEjoO+++YGnHBSiz6WMr+oGnTqDQr8UMuTf0b5Yl67S8aDNKhThETx
l+Iu4m0qB9zcBaBW3DFqTzk1E5RVo27gZdltcD+GeJ1TV3buibJNoYpgI2/+o8662xvi2ct9tlf2
a0pYyyEofuJWIb7Brayf8uKrJsuY7yaijoxugX+e7iNjt67GkVtQ2VGeWbNW5zgKmXhCUt+U6OoT
FrxrvBgkfVag6G/m1I9IyAOYIyRckZcLEq1WgZ2py9djlQflYeoG42+KZ8ugXQDGfblaQzjlPz88
dPRU3F7nKuXBu5rd4fp/+FWD4pBCF/blkRJD+EgVs9Meqg/vL0Xs7X94PVxvamyY2ex0svXq+uCu
BZZcJ3WIv2IKIPTo+NxlQcgFOPKdNIcAfUajBox6PaoC3aUlBmRlndeM7cb9fIVZrBOvjmpRqbe6
/G8xTH6tPa8f40VSYWImYvfy2NfdQ5UkdCD3fLEfWTrMWhMNKh7ZANkvBfg2bGInUkLbXiq9Xvtn
ItAGRckY4g7ii+UtINz0qbcMD+TU/CAT2HTnsZhmUvxO6JffIFPFKsRuPy1viwwPnV26BCScgg0X
HYpwA2wlUTixD60oiNeoJbThIrOrq0TtOU/8MZww7dCLmXpQEeFRFHlLqVJRynelJ5CxNf7CgdfV
OIPGaarQtrzzKLUs4D58rvtGiW9+cB67ZJ4sbj6hrQsmvR7FBKz/vyUfoGqry/dGe9e1iL/4fUq0
/Duc1n5PwNlQjfTKy7O83TW0xtZIx95PSR7FXeN3mK39nu5DqT4FGs9YTdCFjculdG9kpWqgFIyy
AOoAsDq1AXK6U5Cq+j3/yd4PaXt+9+odx4RlBpGAvHow0pIFNzxseEUJ/AyPTnnGBksyEo755zzG
lV5ZeDK60qizMy+7qLBHvBRi/YpIWWqSYZs+s9NEme6qhz0VIHZnfcrqs1TWcbjL0XTBxGT8h7zY
z98IKR7q9Ay8XoD7pA73dz2UZz7K8vsxS9+CX0o84zbM+/FffJvNJF0nfUL0HMnwbS/UTv5M/tht
7E9osKQOXV3I5tk9PRTuLcGNNFPL1S/h/0MB+kg3CtYzeL2YrNr3/hDJc06yckjMRkY0a/lX/oO5
mpgjyVOdLKHKyCIiGasOB5xctpa1vcrSJyiSbq4I1Yc+CyZS11DqpWDNf/XtIUIb5LhGjI8NcXF6
9V7WoHSOq3FqDQ6YRL5eIitIsXlOACPExlgELrpEtsK34b9ygwuP4K5gjF199KCnPuF2fvUl0L/S
KYSMMOge1VlATO4aPkGsI2GoVcg5dyuurf0YMdiYA+LF3pdDvpVFVKNCF4ltQQ9Bp5FaCc/2lKu+
gWkH32iN8HRd2U13uNwVvPU9K0DS0yEliWD7OjV2b4mA3AMoe3+ci5g/XE4PFPus7livLlRwJgy/
U9mxkdlQV8fXg+2lIiS8E/o9Z0j4D+d6Y1NqqNYn/f0ZYVGrCvNzalp4axp6QKv4u2qUHVi6pUfO
u5GGiojtLhHsKsHj0MvofbNerlzq3rQGvgy0ZjUnrAPkLkkHH3KK/el3N7UoliPF5NgqN5pQ3hJe
wt3Wg71spr9RYh7DY/MiEytn1jijFwh/sJtFNjZCkQYNHaI1tYr2pCkfmZgUoG3rqklqvcAmod53
kkfp2shRcZdelVAtZVEKBBjI57y1R//YC8H8yFCqTATOe7C3EZrhnEj29UfPEjq8fXCiNlJCtAF8
0on2GHxkr9VCNnPqNIzKGvAf0RA5JohDLRByzwDcW58z4znp9RRgGXKAKC4S903P03LNDAkRPdHa
Tri0gM22iyDueLCGZdXk0leB6jEQ1LvFs3HbNXBgHjFD2LsGH9MQfi1Vcw5z2Y5/xxPISpLYu+Ms
curKJPXPOT5i8HiJgXn5HTvKPYKIrxn4dnCRY0gtv8Z/40IJ2tbnqitgPK1MujgoElGv4suzTR9v
Mlf23yLXxOrVf1oeJdN4g0tef+x5luPKniQJUz/cYnkhFVfOjB1DgramT9gm9gvq7YtvVE+N3tr7
B5jYc8dkSJfPuVlh3lXU7PThvT4UGm6RSQdDf5I2PlpRRJ1vEYTfujQQ53nbltvM4zDNdR/FBXIS
qr0jfHAIPxpfX0cZVQ7xe8iIqhA8Q/rcyt4wAbB3Lhw9WY6dkHSXFK/mZtg9xZK2CiB/WegWySu6
FK14FYDydOniPCpcqt2H0l/KgGtQD09XZ/OGdzafZvBGaoG+6XNeR47Y4QQ67v4YbZ2JbWX/70Vw
jkul56Ee+EIWK4icclkHF36FSRiXJM4M287RxpZmINOE/Ay0dFyA8QKgH4FMkSipus/xvsdITg0W
QSDlUL2x20tmvimCvW1b7BjZF4dtEOQSLRSi2Y2cyVPO19IRc52eb4+5layNI1/hvjQcvibkZYLG
zKjMP7RemTVpW+5y45AyQKOFBmmBN0rzZcaQBaFGOn53J75KSxynYsqYdTEiZ8Ejvf3szzPW/WWx
RARO3gNkjRzBZpTFkF6wpR/+dC9gm9WtoJoF+pF/EzyQtJH446HD7H91tDtkEWQIdjwx22HdOuK8
QElUAVa+nqj4SUkKf2BS6L4iM0Z0O5fAUecd6hunezGJK1C3qsp5eIfIX0YjZE1Vq8Ee1DcGE5lk
16bhivygwjrmOjm3n+wwqb+tI5ztleALLmXgwrqq27e9bz+ZobH5sJ0PO8ikNs3KV2KdEQef8pVF
6/tcJfYchXg8vXREzlFtgv1GnYRSmohsdMl5Idh0Oj0yNSShG//aHDOo07RRKj7zVYrIyN813vWH
T92NqAjXNb2x0G4YB7lq50uPDLXTnHCGEXTZULc6nhubIau8hnyY1xHeonbzkzCoOq5CENIUfVuu
VgEtGW7A3JoSBwkHArtZsD0d4kqioc5jKCj4yalhqigRhmdmr2l1uQwRsKlVo+CH38VnTikQGeH4
sFN8tx7wJ91qhFA9xSx6Lmu/jVreNcrn0S89tW574mSVTeLxIhskbnoyua2wmQ9lBf3LuDhpHvfq
XO0iaJCttfB0xw8uif4Fkyyv3FD7QnwkNTWnx+hAiTAUiwZBygcbhxLFchDya+UKa2JvSIzW9tIz
fzgC0FgTyGmZR6bbkWzcM8VVm/bin7oeUVZtF8z6/1txXUDFIhGG+ixGI/oKdQdhRV0p6/cHpB3y
XLtzbn33bakl816Rh6nO42av+L4P25rAXxvjGQd2Un2ErpM+zlG2kAhOnW+oGc/rnD/G89ssI5Dl
E/ukP7YOE3dBUGDiaCEPQpxh1G4auCPkT4T7OuOP2q4kvFXhd2WGmZSnaasJx7UgsWkkp+H2PzG8
Syt9ugDhL0yPY6QWQR9RwdMcusk/fAl/3kE5EWNb/VBxDihos5OmbgKHKoHTqX5igIDz+x5e6d+z
T+E1+74paxrqIdjJoevF9wz+9i1evg7BL8pLc8EEsGOGO7L+v9guKupPE0U3DFgbERt7q3aUEuI8
Ty1TaDD2MHG4JgnJGsBcTv3gFn0gNoMjJg+qcRPIMacN7kRnyrdjM+Z5hLDB8zAF+ezYx8RP378s
KkJDkB7E6aZtcla04Q/I9qudweaepHBWytgVWqqeFCw1wR9S1kOJ+f9+GIhQ+OfF3nTBvjWhOg+F
H+ZEfpYgRF9d7VxQm2kOHCiP68ABXJLgTKyAZcK3uYP0jWGz3UznP9F1DPLumRdof2704mfZmweb
D7CPakOP0CMAsVXybbHIQ5BKgVbjTpq+HPy6QE9oN5XMmUDFqoltoPcCBbylkZZoSRzQjqtSaIEp
kIRYqO5kW/R5mfcoBHXcCgEsYPBnTGLtjxhIDmcZHFbILyOQk1jEhp0rCji1y0BOsOrjVf4gGNSK
fqF8E4oyjZZOsnlmswsD+TZA/n9XjVrBsVLTmclNxYgEfCioP3CRCP27Qv9DwddguTXU55fhLaEG
8AvNnbdDRrm3t0SrV2ipyTjXkv8tjL9TObF+RhMhYo/PvCqf1SkMpsoOKrY9r5eV9h/Lr28/13NU
70fUfT8xohv3L1Z5p1QXfq79ZFegmmSbU4BbJHRmH/UjXmVlKVSYQ4HWNYx09yYp2r82mjZAEtad
vgwfSPJsPoUDL9gQF1wdR3UZg2faOgZZ2vxytwVplfKr0Hr0ylR9vu81lA/icC5qbAq/zY6jojSW
Ifw4NhDNROwmc8T5Md3bAWaYmnox19oNuY77ISE7Y75Q6BZHQLeJYjIOzV7DBWQV7WUKJvSefMrP
Cm2LGreSQMkuDoqltwHEzqw9zexm9douibsJw83yv7vduw0aR5HhJv4lux3fSBunOceG5PY4NFuo
7MJAVK2tblWrE4gpU5lO0d8UJP0/3csk7JxotSc60uekTbseoEM/BpKUjTTv20IlXiXi6pO185mf
2gkZQfhDawmRVcqxoodV0dLpo81dJilHtlZJP0TmyU3/Z1qKN8jSYgy0CSPrLtVMInE3AwW8AzKR
9N++ZO9IpmA+4Crm1UhYrQp3Cf3/dwdsqKMyK3DvuYadw75P7gIpxCjHDn2gEwDfOYQslGD4FbBh
wC4quOYF5CPcm+qnNw2fnI/+hIh0EEKiSbMrJFHRGN76NxaxEi1/wI+Wf8ubb9PzTbM/5XVGBCuU
R3MfrGi2Fmov/CkdbPAtXjuGvheWVPIWvlZec9CRr04RazYemvrzm+v+2dxgmP7e/nzBih9CkUfB
1WDEnf1Iq7n63p29VbrbUsiTjD0+QbAXC3twAXL8KHp4fZm0trCsZV88jbG2Q95X5xB0ZNXLlQ11
UTzoC0X+9e90K6h6RUJ5pfJ9vot2bbRue7okSsn/UzG9z+ZW+uJJC/z/5Obci7KSOsBrC3WMOqvQ
XaJqDPjgQ7WCmPlxGUgHVoaJ+mRyEk4sQOsLzdjcQZIi+KO8IcGP/llUGmmgA+//hpZXVN7u4sv+
k1LdJVWkKaHZzPPs1Qc/ETSbZAWZa+08BkcbOSOO23/464GzB7HTeO8wJ4sNuIx8i4ZIAVzWU2od
X7h+kWIX4qRNonB8vLL3ooSj3mDgmDlqL9+IKGLwzcq8Lx89Wr6fJ/hHctDCnzQakkPUh5Dte22c
zK4Bribq5cAHek03MlU7OpSW4rsqXSnVhYDpDl/yGdDn0KzpniuQkUd1znAgBBjt+cCk3gsyr7Oj
jfQ3FlVgX3NzQInbSoCyhM4bhze7Fheu7rBD4M3RphzoZthGEP5n1M+LIOfpQ1gQGvMDSb3w1Ty/
zNFlhAJFzZBUyMPAyr67ffh0S4qNKQst1OIFAGGlzIJV9DjRMxAdKQWHDMB+++xtLK1kBrXdzpqT
Ay23OG/8o6Fhhhj2GJTGlKAvo1goc1b1BqUJAUxi5CjXPZcyuhXUR1ZptFVslMJJPx7wLvB2205B
o3NklbtsfgPiyikYvuvAblOR4S2Riumypz8Jbtp9grFnuBUYi34lzs84Uq9aC+DE+js7DDEu93FT
s4goPEyy5tWznowc0MYntbf2ABxwMDOEVQTBvOfDX3ReHa6rVGO5nP/rg0F2JiBafRxMvsUm/B/F
hbHW0lfSzhdA4NrvrYd0erQ5S0aqtShVHLZhh86t3WZgrFqag2McDNFfG0HJbkZjH7WjK4ntSVck
3/2o3EcLZf6IRpEeFRNxUjALa/1yHC6veJkO9s1Of7AiBqbd/dquPYUo1G2AUbAnI/H2A6EXPvKA
if2Ig1hBIKUoG4g5VG0K8bIWwpQ4ObwXg03z1Dk6fwdqQeqAbytWpP2qK4NSCMbNYCU+sHiLqhiW
ctgtGWthvhAKvlbENsoG9THQEVUuPD8EAKZOzrNkdqUy7DcfkJkpmJ8R6KHgdV4QLWLz6s18Kn97
7H9qBJzePn7gcXSYbYA1Ni9zN77f1VtylcLY6mlZ02II/iR4dnd2OAFMLvT79hISY7SnA+FmtBQa
YqNmRi9Xm8wKbwo1ncxyu1oHrHESYYUyKKs75svMliBGpUZgJruHndLokJdFX8pZH22Fij0AXmXH
qQOR4vRmQ6zxqkA5wXT6Byr/73vHeJ5LHbmjbK3AL4hXeGJtA0XgtdYO8pjAHB9/dFdW3lePYnQa
lXvpMzyTH5VEtlHIwur+8aFrnJYarZMdSArJpyZYu3pW9Acgba3FglBVG25X/ELHa7bXqMi4cuhV
uj8QeY3s13FzF/iWOJuHr+S9HtPcwo2DbGDB3pwPwibvyP0pET8lRNKXANNM/V2ANAEvdmtQb3Gg
9SsGzYjhj41V4FVWiUwrw54ugR8KSWSs2pwmPtXGvJqe26vFYxNhhGJd6W2Bd2/PMJaEaJFMVzND
N+DLzERbviTKy0R3zcWE0RB/lOIeYhfVMsGbfFbG+6Ay9v47n1AGGSF8kWJYSCZawfTRG/vgG8n0
sBd3glJZrw7lEvJq/tlxCInHWHu9qOzbKefmHgaTSGuqarBdU3rsOQceru9RlTcdVxpAUIXU22CA
Kdtu98mw6ycFDEjEzuvXxyPYi0E+QPMr5PjfNvnBi6KJKOeTPF6oeE2h1AokNjaHZfx1/yXxT3eQ
/MaQ1+gi4M5d+Bb5vIoa8BFNycUxHfi4J0S9WDa3RDJOfxvhRoG88w5PLEYaZVIDrzQIUDFiLpCh
mHZwJw6OcWDxKT5TpaxM4KALeKtANku07AHbl6XKG/nWcDj9MLbfCgRykYHmBcoaIGbYtsUBedE1
0zfJeNfYnblzSGabmFysKqXqIpVX5i8At0hFJQbEg4RckYxTdZIhVOsvXwF+pEzx8N6vDBV1WCJ7
KJSP2tBiQm11h1EAYxdwsYnBomzvkhm03VCYtzrxNUCmiD6YvLo4nn4NP/8T9Qmvjj0XfnFBhcty
8BTUTcUegnA/9heslg0AEK7BP7lieTc6UitMjE0P4eb1nOCsLyqUJ+zbVxElJTycRgRk0lxYhrZ6
qDD9RYDS+vbORQ+V89hA0dj0U2jnYn1tWVNBjs4ArQwndSK7wKBVof4qWQKo6haz/0ZK3FwFxG5s
CQn++019wjytUEzSVrDqH0t1P8vJaT5Yww0VLLXmlt5jEtC6AZCvv+3BGoLcBJwowSVYvx1oG9UQ
RoCxVDj9WBKS6nbOgVdEulc7xd0y6gIoQK1E5kAA8yIiB8fNH1J/68MjHlddNW96wXOCYOYsp+oE
CFOWMb5BZspvk+LYiN+GuKD4T40EHAENpMNi0dF5fjOycCFTkfUXLs8axZnGnHdA3EbxVnRZIxW0
C2SgQ20lWFgsrhbaiHkdlqTlIM+D82pKr4ujS6ancH2vaKVziAc1Wnks4aSwKBimbewgQTl6a78I
M0b852/2dl6FbsCOaA/wvUmWKEs0g+tA/Vt7Q0HOGBslMwXRCGxAgrAbeuyXSMJDALA66E0M0aZv
ZAHZptBDi93t+fFXfIxEg74CxBhQ84pvxa99YK8ahcbUOmGKE8qI7L43TUnHDCex0Fx3ZOqS/T0/
ItW2+eBQyd8hlvvF9Fjc4F8iv4crTezB5rFAsEKjAtSrjf0zSdUiolT1rCdbRlTTgTYa1/0oeIAg
2M0tNsycupQr/8mYo70pJPoHee9tbRRexalEGozr6lnP74R20tskGSiRSzKzjGNgHzvynGHlh7of
7bh5TxxCu5Bn7PLBGtidkCyo15jFVNUnpdz8x8Nlfw7to9/8AUwm4r1e91XpUulYQOgF/5JolxdW
mPnGPyV4DazzzujacvAAFMSpxm6FaM0D1DIMP3Y9Kgia7yL/WGzag5GpJwcHBBT1JwtxzzGpFhfN
AYWkSkkItAkAJfJV/wDtVuhzZFdg3JLw3jn8lLWVf8aUu1+FZWV+BDxArDw9I7XK2vlRTpeDDpoa
Js7RKd/McWPprRwOYYuQj4tKAT7hhnAa6sdvJjcSBiTzqj5ao6OyUsz6dHVvk/Hdc9VZlAd6HbXn
xsxb6N8GXZvvvKz3AOSsWMeXL+WhAPns/9fS5QY4mfL5Fa0vlHlFpUF6QKD8DQSmfqCeMKj32cdJ
p/MPaoRtL0TdLiR/bjZ4MixmgHJpB6EauY9xTQmHt2GH1fB/EahjSTSkt6XuxXY80tukT9zk7iZ2
BHxlYi2PHpQW4F7RA+XElx9Gd2f0t9jist98I3nizvA27ePLmZzl+MycOuh3Fg36JoZWAh/csYIx
8dwIslxDVXFQB6E+SgjrqGWPIAkABV39je3LSqY8NAbw5tI17cdbqujn/gxjyU5QyBE0Fo26Xk2h
MxpVEwh8WV5eiXV9/6cCztvhlVq1Ame7WZBc8KyV2e8qsWmhOp/I9PGn1uyJ7T+NyqxICEdWfRo5
bk/gWdiYwjBMAZFD4+AUtxIpURLm8A2qrOOB6VUxOIMSTvwBpayemPpQdZSgKJ81Rj68qZ9A1bi7
AVjcyGG4/s7zeSg1Z02qKv0gbv9K45y3XJWsvzrMdkfBrFAkux4Y4GNj3wP6+nt7VgrgbdPXxRRT
JRMJKvFw1q2kO6vkyH7xeow6TAoJOX5raO7yYNfc74A7cc6mLKnOqh/l6U1MhffbfyoD7j9/FEgo
LVhKfuPOhiDZat/FQthXXGPAuHNLFu+G09HO2ZnmUfeKUecaU/Cr8X0afjoJfhox0Lo8aGjz4ge+
f4bfx5N9+HyFyYlbBKWq7MvL56tOb1oBcme1uLLeijVW4Ai807+7eIrZ++Gyqq8SD8hmg7j8k1h8
w8exNR82M/8tApePVpBKPdigECZa8m08l5O6ypye2q298OqmVj0npRMPCkd1fJnncjxMFVX2j9br
VCIXOP3Iy2DyFEZ/SKQrxceBHbhEI7AsjEMHaMl6FUS0VnNtbAIpXgEMb+NnaeQw3T7brb+xrwrz
zZUoQd/5UIeVFeWkLc9CPsV2bnzfIrwIM916ymyu3x2yZWxHqjjRw26cHGdxi4z3yDCacWvAoseG
XSSrdIDt6thZ2MqWg/FmrCPPSAXmG6uYsJT/bCoMmWDwjnxkmg10ApAjRDxRXLd6Uz/B9tFm/DpJ
kUXbOJiZ80J6p3D5lIt8KAzOK4CQ6n83FNO0yNzCtYLs6l547ygJipGVrpB68v1WpW3Y3LMMqHYq
SeW88NKeyvgHUVFeHslmZlsxeZ1Bpds068Xqfoz1wypQWXJEoiMhygYXu++fmjsFLVhHZJ7Dsh/q
tJsBSL0SXnhDa/zsP+xRH2afhMm2qR6NzXM/3e+aTedU12LUDkn08Nq0Q5tNBFDTBr2qptAJYGtp
4JReY3a2xm/XUWRffLXw22r2ff47I6tQU07Vb5V8lQVlh8b7I/HCqyVxayNNHfaBvRZIcNVPAN9x
P9kfWKq42e4vXPPYWBN0A2vYHH8z21eCb71uZ3GcZFN+/Ew4oIbFHi3ut2rH/SN5i4Lf9StYpwQk
8NXfGy7UY2NBpPJhLE30PrVdZSUc1+aiP/FqzE+rXbIo5HtF5oezHa2eoTZogBl0cm6FIghYmYq6
zyBWhs+O/+2mr0k7eT3gUq/74eQCmPoSeps1enrNnUdmhqZCWK48RYQNzw06s4OIi6MWoSQTXXN0
fLeCdnzTH2dmapDzq6fPNcLHfsUw+6gD7ZtY1fVXA+fQm3v8npAaviAqYHY8Sb7NoOg6xl30zCe8
3OWCQ0pfaatyXrTavFub8zeB0WbeHoxpt0aPT6/e0bpIBFFAGA51SUXVuaU4wm+keg0EcuWmJcln
t0RYYh+T0q+mLGdp9vnLRzjETMwbw+zyM3lBavTcbvB4tZoL1tEu6Q6jcGx6NI6r/Fq/wuxvYq8w
gKWGClzxIxqMHXHPa9ALycIutZj34AjkUP935EqLM9T3/+IqDEG+eJk4piPBuKpxsrbghvfqr1VS
nWCeRTvewZrQRDtm5z60ubwecjqr+O00/Dfm7PO/5DNlJVUZylm0WG4oeHorQi/qqq8t0WYPZjh0
DTJlAHt/QLVyVw9IS574xUu7EKGdrz2bIY6YUwV+os9WwhQxJ7Pqx+UEy63q4+c7/09L0wRWLpPt
GdWzsBlDMzjMk73g9QX5wKb1ct3qu5RlhXSIXOOj+DLrjUb/xKwP1nCH/ynKB37XYSbRFR1zHk9+
l0s4PeNjyb5cALzNFuOmXGumUVofXvpTjeGdIoSs2XcgMbXmAqQPDvbL4AW4/iCtdcHkhmJqtJw5
7gWBf4raIPV56/wdF6HsjaT9UkxkAoJEiulw5iaZFZQVd57I0y8LYg8uoN45Zwg/dib+qg744Qev
uTwC2fDqZGlOerK+NJF8KuHJAxGmjxew4VhZl7Czy4xqays7PZgR5TgDHFf+Zz0onIixDUfW2ILq
HDM4eOTLDpb7xopqxjbDZQr1a2evPY/eqxsR4BChd/vBVJBjTPkycx2VWrTBf9A9MJZxLEq9f4uD
x2URwpmo/qSGQaOF8SxEJb7myJ1MChictb1jxUaR5EAGxJYJI2RXCcVnvnjGfuqWNnEve5Sf4H2r
Q+PK6olQDAjwSIQukyf/Z6bHA9w/6371M8xI9NdqBwt5nxOP6z2WXZYqgquvretFw4gcL9bNqmDQ
uvvljyRFSBrn90xLBXjNmtIaMeLNsZ11CehyTZh3P+pzK3NPZdyETTC4gmtg0/TPftM72+RAnNIF
gtqnv3wG2ORWVLkwy7Z1ePEFAP51pnRMTyAWemB0fd1a0GTidzN9OXRZhQZ3n23zb2VWKN+VLM/m
B2M7X1mnVbeCBOMdE61upbYXOtxdRvv7abCf8R/o/4npPYZUDhe1P9aoAydErPTVzKJ1k5tdTHZ8
TIvwcJx5BbSjVnmkuNRGAVFy60oos3mBtkCwoP/A2Nmk1Y2R9ZbdK6Jab7hQJsX+IQTUezilWOiu
Uf4p9S1TE8NXptIPyDCTGkUvTIWMR1cLRBGS0esvpAyiiUisz6ttmAkDrG62cdTyok97O6LFJWWx
LwH8U2hMoHIukVS0/+cqBq3Oi6WxjpOTL0LoPSvd0+xDW932YEkSQJLZRIf6qBEl3bJ6BppH4I+/
5o03i16WMJ6+Hty1e+EV9mDmNPTLBe1a1rWTtFtLO25rJKaLxebxBf7OVnTuMfp2xD66lvvUbcLD
3FyaKNoYV6f6RdMaqw6gChEbaxec2UlQNZTmWEIRZi925oQVkcLVZSL6J5edqp4+cjmqswyPxAjL
iGTNvJAo1FInC6AFw7YDHk8mAOY+HBFANdsIvKOD+QWOXRYsTzb/KTOWPvaQLHMt0CPjhfxhOYEp
LWm5Sakq2V2fnTu2ssKeHq1mAnkdmcYg8fbomNgeQNFmhFw+YnclCRLVxorjch7T8IHiFO/kb517
+Ior+qvH6XmQsu9p/B0ABVwWYr0bPe2a5Nk4+nZLWlpiYqqjbv+uZiLOJDCYSw5Vy6MIAAWEAju3
ifMm5PTSU3NHnY1TTB1E9UMmmndaxmsSpc55LfnHqdfYflpelIk4HnTzRW1KdE4LSOsA2hgyGF8y
Uylhno7JObyibtEEY8kOO/CQywYResF0R0Ceg2nbt0uKHNVAFk8vtyGZc2+MQjyahzw+s0iP+TDE
2jou/QpgYo/2IRGq4VMAKUBrSUQqYbTP2EzWdUtB3Qxz3Zo7PG8AKSkwLLOCLd5Khkg+GN2EXx1I
RAlBtDtA5lF5CgHzn5aGt2Uri6Oz5gJf2YM/XGGYOrMNzGoZ+Z+NT5YBHz1xLPOi5SyadYFrhZmc
tQTjjR16nHaFd2rbqorcxhSNZQYqzN+K3ozLUbCJ8Mr6ezKi2XpJnf4wjm3MVIqxFjQlSQdCT4je
3SHoU8K0ls1Ih+09CiewN+tpcSZ6WqPJDSWHx8xQo47D3puXJ30PvWFI+Qns1PswAjMebdV8v1t+
ibsDWfiekTpkIDdRoHJbg1VGzwsS2xiH7QrShtX47f8c6ZSKzio0UOsjnnoO59qCplvDk5UY0n2i
iwdf4CQewOc5Ex8k+2hmHRoK2WYwY2ca9Za4Z8jiS4yhl8K/RbaAoDHggkXgdliCkfwGqocO37uG
tda/c6VlpTBEzO2XhVEAJrzwvZ/FHU7gWYTKfOL+F9JSKYrKW1KzN/Ql+CQ77MeZ7HfNhaTFxHQU
Mc9uryPPWR7v+xsLm1A2oBeKLZY3Wc8kAbJMe6Zdc+XpTWljVLQTQhuVMgVYCqMdI79fs5509x/9
q5n6HCSH8cuYLY6WUMjDFhPeZanFt85GjuG7W0gXjEo4gUHhWPMGTTHhkOJTRmNaK3gwRv9tW9+n
274jQi+TFnmbi0zFq/jrONPeEs+qa+WeCBF6CBa9iQ69BoYczx+kV21B+QuAr8yMxHCiE8S7hL01
eqCkM1h/mNhL3TCYUvnmzTC6Gth1dMYU+5yCL38EwHHwGwaf4GkhdXi+qZE2ehDsPyZhGwxnFrWq
QiigSolqN3a6W/mU1tkOMm7Bcw4307MyCZVt5UgLwRjVSgbMKx+ZlOhjpIGoRyppg19x9e+u8RhG
r2b6rMhtWiTITBYkctaAZbc6CvGVbd4/lr9OEesjc/bWGxj9vEIaRidcUiCPa4YgiFVRsJ6XR7yY
Ey1M1RRFTZlo+96YLDjNl5sHAjJQi3bi1guwyRKOc7ZUiPTJpb4FUttUeVY3Ee/lCzOr+iz4Ec0p
O3MZmkBk6ZTp6iaBZqyc3qkYn7b1gsEiy5UEoNVeYIGlYRThVXf2zgF3Of69oh26zKrige6f+92P
O7kTzSKdA86pNgTv2LZqwLbinBcDAjJrVWAVKWgzojopXc0L3m77GZavVC3pVmqXZliHc5KjyeJv
PFesgK04HPs2cV7+X/EMKOLqQHUUKhoz4Gb8+SJVMzFAdQA+2SDTN7JbRX1uKGGpuimc2w4xgEs/
liMOzwkVjBOIs966ny1ytDtChh6C31/6v7RVEY0ogjTHZRYl/tqnSaRiRymzQ+3zEZ2avZERgXyq
fwF1zpMEBPeQhBordmIwL+0dp2wBl9dCB9fP6ttdwNBQOLCFPJRyKT4FZb1XiHpXEgmThB/0lIN2
LK2zXiFcb7BnpgCZkK/7BUoc98qS8QV13RSuX+hpx/PTm0E8vMVqVNN1MldOCfhRIk/bp796MggA
wVtNdkO0hmLDGuMK03uhpJf/Oe8kCv4hGCfauvAboWpCCpnTe20LIgdlzzDD5j6J/to46aJ9Hdqj
95IK5C0XLOPOpVTAmolI4aOltR2JFJRvTf0KTtR6XqeJ/aIY3DryEg2aRPhce/yOyh6vhzgRVkpS
3p1+t1yIwKz7r624Hle3YalHI6lw+MXMpqU6Ro1PNsPe1RuNgscTBEa7JoXfhvFBVagQfUPPrZJ4
YZlzRHvmmJAHH4WoeQtxdnsB4aJ7F8ogMnsXnXkYfzV9e2OQcrfp8l9KwoFTrd0k4bp4jzz4prQl
skPyvtxj7VQuJj9FfgPfwE6PHjGXSUJIWeWebNLvCHSo46h5MqqqIuimV2G1MvPf2Zi7HBmK5ILn
JIU1zp+wmJ9YmPMj9EyzqmfkVtncp7SshbKCdae3lFnCOtBTxgYYhmlGKdz1K1hoikfAjnxL/E1g
G8BMN5TQzLJOVBEoQgyLZep2Ud4gWUCn/A2exR4ju27jgfI+GNvsRokNrOK/ExBEf/dVJgRop0vY
qXo8i+CIQTLvEtNcGBhrijsmNYavI2zSdW6uofuPLelFXEwGAHhOPiFmrsAEtgpKsw7CuhCF0M8N
zhsqsdE1Y5UNfKy0OANxb1+n77Kc0hObHsjc/8HQF2rRoraXoOz+eIraa1MP2VRJqKJhG72Whnik
3vDNbaReFojGv2VfooyeEtrtkajxgZboIZQD4nrQL+bsO1W3wxBBGBxJfIA2hQyfl/JMJZuimoHF
u0rdOFGaJybV7uONTVGuNH6K8etJ09t5yrgIwqgJ25xvI9G5nbP5izlFp3Wg8SUlh+1p2nV5Ri2/
d+q4DO/SnxehKuiLyxJOkMsqTlEpMi+hRQVPe43/dZAOMyXnDZH/tXcIST3FnJBfBXZOQEhgPwBD
NQDgxUIBegL0Nm0yTjcxnOiQH1Bg+WBzfuvVm0u1uMo0eSV4Pf1hqOU7G0hsnS5HrQdovAXw+K6F
llTdMYEePV7gtwKOjyxFID0MIalztljMXCTUBxG9T1ObB0MM8CInsbauJ5vUoQiQ78mN1NUogS70
hvmpvHqyN13NXGxxLBhGc7bVUE/qnroyn0Fb8bu0fMIvvbCtVwmpyZt9HcoAAPo4LFt0sOEDxe27
xczJ2frqx8lvBNWMe1As53kvl/SuN6S4laGJqkuLcbTjniw7LzcFflBWpkhUekRRkzrUDSOtri3R
nOqAnGIKbIe+Szbv7ccPeNGFBu9v3N13Ofmv8drxdjvQBv4Aq0MKw0Myt2ehWP/KGWsMa+kTcaqG
njE5ZLboFKZqD0/FtfPJa9q1RCz2UXXL8EP0xYx6/nE525ZN/BSOlgMgOW2j7KIHpvkChfPh3xv+
wTL7MfCFS1X8Ipkx/n9Ty+4lcYrz0onLukKpW1REvNrPoga38JxS0mDnkuaHuyD+qo09PleRHE3c
RKZFvx5EdLZKP2g1U1ya7dm9prCIFIb+FQHQpwNF0dYMY2UxXDNdTxe2qvkKvbJiHP0YTn+4lxvz
gprcaJ9vNaQtCkTmj9en/WUtMwIZTB8UUI3rVQZ/WbrweSC8PX3oNGBO5AtVvc7y68h8TtOIA9mS
uG0FjO1eqOv0+286nWAL1iLz6q8deIH3ULBl5L/X+PcBRbQd8izWeUp2w0EdcoVxYieM4cqx9BHE
9/vDOLF3JZUoW5zGpcOfke3AT9EhvSZ2jhxesk2ceTOgXEEGJgsDwpydK4XPBWppgHUkTrOl2ehP
WUYhfyLfRHOIw79g7soyhGgFX7xLmFchuu8zcHuhjzEbQynQcy7p3h3wej4egT9/LvibUtLt2+MT
RpCLWOTLqTyvXnd3LKPASIYI4cjGJRgx7Jwp3RIELxMb93iITNU5XtcALenRwRWaq982EGdVCS+P
pS/qYp7AnIiP7WsL3SBZtH5nGILVi4ASGGT7nV+l8DXOjceWISbW6ULZbW87Wdg+CJpGIFAcuhtf
Ck0Uo0IcHEo2S8eiLUgZEf6iMxV67dR7czzMoLXB+hF21NlEaaj0TD0RkX5lMgr7QB4VqyZUC2rq
nsCDgD57okZj9VZFzpB9uQmki7ezToFuIwJ4KEQkvI0xBOYDfbSezAGWVoVISYSGW0sILDyFyuxW
dsj8uQANsUssaA3mDpMdZE4VGFMpM9ltrjLgqkeqnPhY6SgaWDdwm48bkOfGB1ap4uIdeyCTkdp8
1cclBL/Rz9Q86UUEzl+APhwzrSR9CCjWW9w7xQAjigBmVs8JBxohz+F8hVeEoDvnjtJznFzHDQhD
H3aYUXeBhtanaUSh6IQbWmicdvbtV0yUrphE2mbgeRIRs9w1mirm7s+xLj5w5zMjIEGdiwskRDoP
285y/GY1L9btRitRVNJf6nYSyRk5AbMog5W4cxk26cr6GhhuUGEFRVYmMHw1LWKCwDpQlGOyCta1
hoblLngrmTw4tQrmRAQ4VMlIeulB9jdCK0cX3mEZOF4cyD0FXV2JeQnGGVFESdRHC9HJ9mHxL7b3
KG5lpmYiplFHubYv8MPVXgIyYGPUKm9RbLcZYuGR3OA0fDd9WZ7xS2wkvXQWs4W9uYhkNPaYhoCd
jqwmRlidqR/R+8oWvRRdBBd1SgdhMyGEQnBf0ixi3vlqAMcLDTl+v5IBrz85p/IAzTOFVVmCJ0fE
jvhS+wkbWl5AKbHFlD9R0WsFPvTbG4gex0NJNXQHVYMJ99ayUeZhnnlseYy0ja0Ild2SiJAlkOxH
cM3VtKXRX9bONcQhnutoVBXeZlDg7/2UjOJv192RI0Zm4Ibh7kV6tmvw5IBkjn9+CP8NdQl2UEMj
F7LQgeU4uTRTAZWAv5weIBKPkGVPB5E5917Q+w0B+4Poksbx290CXEmc5K0s6iLaTC1P0MerAgNl
zOYvfAzdvBLiO7rqv/3ox+Y7FcT2GuTfRsWvdkaJ2WduVpO3j7MUxLyD1aZ9XDhtf6lFuA4kBBKn
ficOEoyO7sQr+nFFaWQ8wMEKBMlanpHlqE59dsnk8KBpCTALqQ3lg9RZ7QV2TkBF0jT2vCfu1h0p
eukbrotwRVCIKm8RAdqEFYHMDQAMfQuvjclmUIcGSWcimHapKKtVVgTptsAknsxGLNvjK2BIumkj
zJfsO1EW0msWujyjizFieqpJ1hTFDSxmAaJS8PNR7H9Hi2eNfnM1qY+s8P0xAHWDqrrAVDnXJ/NH
bAN/VQdjjyL/Mco1GrO9Dd8pKNOd3Jmqnv99TZy0CaBg7H672DCYar4iavDIQp7o/HDf1bkf3ysj
8ESx/RMB4UeGt5d+b3EvNPvVqxnFPd0BJ5p6c5Cg04eflGXlgIW7Q/gGxm2TV/bgypyDcWc2nvNH
qBJXarrPbcNv8a1Yx8+4nyUOqal6wQlKGCv8o6pRiin4M9cQar/UHRy4moFqeK/ZJq0jvyCvq/uv
22OVMwz/vD8OaMcz5aOZKhvLqkhixcrcq90IMAi1SgkW4c5GDpDWuHEavYWUZhCZSx47kBCVLPvl
g0OPUxFuUx3DJ4MFYo9CW7b54KvO5G5ygyiZi2gwl+sD8sVtt0bjM579wc1dZlYJiw1jRPVzw20g
iOBPmi2x9UlFFgRyklxATZZGrgj2mPOmxevkZpMjD1ug5gtGVnB8udpAAIDUsqaZN6S3tOP03R/b
aQ3WPn1UlOl54Tb9GQgmSKKUrkfmQGRzEaT1DmtRsgNsIeuijI4+WSFV1bINaNyPGWH0g1ooaRSr
9AQ3SFHeBPrxtLMnyhv5qI0Jp7HEl9FtCTzsdZlk7d+AiB7nVU2+Xv7yCxJpXadxR7NRMfRu5PHO
qz2pADKcEUh1E/yTaDE52O3CGl2COOiHRyHyx9YQy6bUIlVKiXYDVpg5EFMymyO6XWZQBzd5PgcH
1s2v0QUM5+dILJdD4Atil4m+GgpZm+WhBPmdek2wKVaKl12UprcgAGjiIbtMrcuTzjr1FMU8o3Ng
qMAiROCyLCgKT+9GtPR11EXzpsr4Q52bULo74bqUQIomdr6l17ggidxEcVxnoNyF5n/oH1X1iwYv
I5eSOejwuslF4qBuiJi5L6CuxfjmUx0yDh/In+0j4hqRomCA3ktpLVDok4BrrW3V3zCIgd+W/6np
a+V4vLacm/AowLoeaU2sSXUtjhnNDETDZCyReqBTf2gyHm9PMDEJ0Tx2cME0xfQQVofiARc9PU3M
TrxYo13k1d7GTvcVIChveoZiNae5egZVX8COsF9Q7hu7Dw92S1SGkq4C6TvOyiQkhSvXWZfdiJH2
4pxzpT8Rqhg+YXe+fFhMMhi0lpWCbDVJHX10xcRuFY4G1QCWg7cuKQKz2xnOn2zK1qM9C/FrE5AV
b3WDdXssBaNowv+8yyq7AHvxmoKIPdUUlhOrufsAUyq7cviJZyA1Hn+uf2EsSIvhnuB2TrWmTQB/
rj7+r7vs9CAvoVz9FIOkriDRWefPl4BeZnMneIxlK+milD7MCqqvXPJepEgAecK1BUEI7bnWv7tu
WWsWIQ8GoCwxBXKcc3cRpPAJ5rYARcsTVasnHJlZWVSxpulHjIJNM0IbtoXkH7fSUTMwMoMFId/4
WUAp6E8wa+EBIODgAOzgWXu4w+CuvcUFv9Sj1ElC+jVa5IVhUCH35h89FC8C0S2hidpPvgqh0XbF
J+RE32FUZM89prUWELup7I3NUH4kNfACn68SbXXBUM5Hr0+TZS/i/v2hzxqZHSFdbVhDz2CvHB1f
G95Ez3xgXFo6Hzg1HzpXSExTgUaUSlEKSVePmO1dYMA//wwLzFItQRBGXrdYYd+dUPBCBi2m3YYy
d61Ov5Qu17rO5kTKHRNUcsI9sVqjzOoTGdspzdJo2IW9ZPpgWka0JWgpoK0QQovN5JGcTi1fHHnA
J1IBlbXpB+9yAFrFCUwZ7MOSDKc59447WPYsizp29Ks1hi1AKUybhXdkArFqcwP2QUOPAhvFuRom
VgE4bPbz31sIreQuAxkT8D3enf7l4CsB09u2z5bdwY2etE7yjUu0TFwXbcFxLapSFLwF2NebKIaO
sXsu1IcP7YJSZIeJepVGdHA4JS7VN1RvZYSaVmuInszRQqvLEANtuPqp+Fj6AIYAHJR7MHVwoZ3+
6/STFMThsKSCrdcsEJpw2IZPPMjX9LRKXYkD2Cs2qx0P3DIjfx7ltrxXBay//xBLLTy6SbWEeyUk
lOc1PR9bVSrsz3MHihNRpigQgqiy6X5vSgPpHdguNhBfpY6xwFjKCNDgRDV7Dp9W6n5TWm0mIzrs
E0ROgy92pWVyKE9+ligWSB/X57KDiHMZ0nOJZPZVTH73pqQXnImd1Wvwx0DQtvOO6oBLEP4uKLx8
WqLhMC/ultKermgxSpkAJkMcbZaAPLcksOq7YQmwnkdVcF6PqteOX7nk+SyXzrmZDzvT5MZkFzwH
S4KQhuQe69SMrOzdB8O+T2imttTgqCiULlH8FKg+b+7vSMB98HXjuG2CyuK/zzj2hd4ePhYUVqlY
spNZPzQjle1DfQukmmt+4jCm9tTVcllZdbk/cI+Y4yxt24rSOAeZUwZsarvL9cxrlhi2IT+G6jeW
MbnTV2BmjN4QkhkKY4ptI1bmlc6+3Pf+1kwcF2zyXtCe24cnT1N0FYiNBHPqaujmDe6Fwl7xhCdz
EO2RNxgxMGWUJNShD3cW7k5dKAYKf80KtwYS/hUKsWFOOa5HuMr6HGcHYN4Hc0LhRi94tS04ooP4
nMm2VFEsAf357zAxfTKnVvK1RSYgKTIe+ds5LxvxhYwa5h1MWod2hbujlOwzXOb+nkYqBErfl0NR
plH/JHBnw5eV/NV+TiFUsWHVqpk3jmfukxcjb3vZgZLmQ7a+S5Z5423dxiuia/Cmld0TFDDVVAW2
d7y0xQvcx5HrhdNVVpq2W9XqWfbabofdA26mxKZTx76NQxmTJbW83mMGAFP+Jcy6vZCPyjdcbKkr
HdJnpkvK8R/KPIYOfAGQn0ONoM8tN//NbD6zG2WXfW/0Nt3gOZD2C2thCb7m1jRbEeLNPcZL3F0T
Phxww5v9F/Ps15LXAJ3Lix9fWTCY2dmPZ0ZGxjyZ2AhAAEZhvX/BW5qkKULu51501NfB77Ozjawr
55D3w4GdeymdjLizF+0warMohOBCa+hG8/9P8FxkDIuVtvmmev4MwEdlV0hGQ9kAPAMLCRHJQjc5
+Strn6UhAW9zVXltd2o89ZCVJ5h5Tx/Aqyoz5l0znjr/PL7MjRt4E/ZOqGqEA6JE6A/l4q5qE79o
91MDcyrl99aAxf50AZNXCkKbDgEj9FFG+jzvLY4dwFsCWEmix7lDrIJxtYoyOkp5k2f4uBDS9FGk
ltKYP+nLzBQ24Obt+prhxaiBbzfoW2qvNbtUEtEFD8FKyFnjAwVjdoslpwp8RdA80GUMaW8vTWGb
dnHnhP6uT6oZ4ffAbYAzDYL6m9pqvOqeNyt2GaoLwrB7X9JMa6UpbEM03+dP4X19naworTW2qqBQ
kP9Nr47j109ZOq3YpXftowHoQWK/1yTJngG5XYIIqsy47So+O3yZVVQMT+sHwRpRbGRgxj1A6Ptx
OfPyWE3IK87ZcRFASzL5azBVZLVZTDKI1TJjpAqDPv7KWPvMFAUD0tWjDY0ITYqjZ/3CHLCHCN3w
fp2NIXSxMufC0pkY/CznTgdr+ckZpozrkjp46aWycQ0GYQpyUY5NWqK6BoLefdLctB1ieBzXFmgP
hm6/wAPwEGKMENS5yP2zziTmkPjAKxsvXONMUPSzle+fEKhCSAmtNUG6znmMJ/0/c1mAl+gzTy3a
eArk6ORVfctqdt6OLRlIqAe/7YAMVcyOGBLui/rNW/63yo/XYY5rD1R3HKLqyVGcBndPYvbjg5LZ
dHlEzh9WDovLRqhzXR3f8fUy9oeywUykinv1gBS5uTz3llTpAsN8zSPjilHYjH8k7gFM89WrEHvS
RHTny6FuXoMt+BvhwsjEo8zQDjpD1YWniffhnnPn/c2/z9L2nhhLmaXw+6i35tMq7ea1pMZc/B4J
Mii8bqMbl3fxdPienWav5d0hLVmJkTQc3piyvr/dVbzmZHLhdosVN5y6LB9yJgE29SCARlFx4WYm
7yGQyKwkJV5DIzulqF9yS1c2Kz4GgMWsWHJd49ZyfxSETJJkIZTvR1xhzTtn/wPGmCmxNARy7cCf
mchCXm2xkEf/kNNeXFGCnvOVg4Jkb8YEnvR6QWEJUNZp7/6Y5QJKKWXMsKRvF9zdRAyDh8H2KWC7
N91wy71zvFI2sjxa1C7qsw5jHOzcRJwgypo49mZlWzJOOhDuVm+OB8WafuNL4XgOCJbvQgOKhA67
2woTYvNxiqJgH9+xS7WGKKzCdNpybjbfEp/f69iJs+k5/Kn3clxY/ID+jKsw5tUdUt5MU4xfSrUO
g8cyrhtaS9qFvxwIl1i3b82PVW2aGEYQiI28VeF0a0LYWeIKrJcZ6I72AX/q6prPAWayWAlOr+qA
mMgmVJUEe6MopcQJbhSCLwOLInTPHNq5GuHUAw3GIgjjfUYp7hNBW9RicZw9dsXFBrQlmxzDr/tD
q8SmbrBdFE+hJ+DiacrcykZG6fnLU401HG1/LyCJGUskZjbMAPMp5CnRHvoHVUXxPW4PzT3c3TdG
1cqz3TZ5k/EOjhYpplNOZi4q/150M/7X66YgBsfZbzcH2LnREzNkBd4bdVfCiP9UMGmzSDyGUjhh
ZNpgl3BMqJTu21fJciTzBuCfecl5YZehsiFucAHwv81aRGsAdO6+KUz/QpozcsAXuDnlGuibHGEG
NYSml3nmAoGYRppdLitoiVJyZ3uLJB0DV8FG27RMYHBdTlvb0MpFkULW9HxR/h2KPKUKujAApz2w
qTZbdNWm0H2mLL74yBiCCBJJ8DXEOMi+UGyOQNo7QBljLsu+oDVfNz72oQ7jLwjc2kbRZxOKoUra
3XVJt+W1LfK5nXpnJZRtqLt17nJRx7jP3paPdxvc6wYqiaZjzdXnb2peW6TXi5F1Yl7JwtFHehaG
c3s6X08aSeIkD1lRL2nBBz7optliEFc66ymspNM6ZRztmRuYZIn53636IcA3VoCKaq90IaL7KczK
W7SFtN6cj2KMd0zXhGGp2czNLhuZjmf3nubRx7Dtsl1oHpNgXVl3DgJl1+IsrANHWp0Yn7gCWr9K
TTPG0m0d0uwgliW0Z9o4X8a8xgYEoBe4xsw9f6klXAHcpxE8Ck7sdW9ACc0taxT5gxSlqjXkGL+4
cYxr54hpLn99t/PC2RE7ezbNVUXZhjLweOI0ykpiPVaxkvHSvSDfUfouVhvmKwfOqWl/tlpZN3Le
kOlydubxws8YrE1Gj9OjteQ/e3YZHOSpvlMpw3TW1cy/8YURLYN/WQduWIP7lTmjn9+nvxXuNXTD
PqF91mfPKmgXuBhrr2Ypqdda64KyPdYZNGtHTNdn623jJn1PuZ35Jbhx1EveT1eNI3X5Jb1vBEcd
K0yu0b/VOP/9e8cF6ixDfm2ZBjgKv3SqoyhkiVFKH8JZQx+x8wB5Wv0HihaolIk01gSryeIxk4Y9
LCsmx/79e0bvLZqR6Nxs1d5zQIS14adwzNKnGuwyaOobDRQ8S1IQBWgVDmNRd7bN+A9z3MkY5qsc
VLWR80G/+f9DD2WNXQYKrfZ6bmm++VX/AZu2uD0JZ7hoPT8yNYZWH6cmLh4GLmK7wiCqz5NQhiXN
a2X/KXt84Vk50xbABhB6AdHliQ1MFrb4WK3oiCPXskxw3dNbYQdgyywahEZXToDl/1j8A9DPF6cm
DcCvhGB80k7MPecMQ6xS+jJ/hRd6Ioplfxq+8hbXPg/2eJdlwj9cgx0fSL1JbbL6a4mRVokgDJ+i
TX4DiOi3tAitv+J2rkBeOX2zJZqdWpw/nzBth8KhPDMebwgB1ZEGjOS2XBGSF/o2OaVSA6+E21/u
zXn+SQjfEE+ezSXCWBZTMzATpLb9SfcsgyRVeJ9pWz7yuf9EhvNskLNMTSUEkDFaI+VdkjcHgm+U
m7i4GgExFBBG/Yn/b2JxKuBvGTAFcCyZf+n//GfrKYpT2FEMKAo4UhZ90mABy3O46YNdMV8PiiQ7
0yE92WlwqnoLYpV2tckOe1MuTzh5HJms2pQj4/WIV+WPoAC1iQNCKfcvSFrWpeoE14MPKL6+kTAp
nIHwwLgFFSXxPTy7yDeax+tsGe9DwjqEAAcsnNpq83nvsEfEJfXad/kduoHHi+Zy5C7Z2m0bCwkY
X7S0d1yPW5IE9ZKVAEMJ1a6brPjUomVVT78MV2XHQ8jncQnV7gKyTtW0eJtXQG36D8o9ANZdPX6L
Clku/O25D6gO4c23qDQXZuyTq8bSLoreL/Puw7MB3eL1+tD3tkCbE5QnLnxXKZXfpm6DHLjzIor5
GsfixUzKuesAkHXHSaO4ekzugvi75ZdWhYqVHBmAklZvJhxPjddyJSgLJ+exIyawHeKyWvDJBEVK
sU1r5YhOyJ1BtxbbmwCNzetnLPczgw/uRcsgu9b6C372x26FKG6Hsz9Q7ugboAatrh6nAISi1Qov
kjCVaoiVFnjWxuEYEhCVO4bez8/LiNv8tQJMFVN5zpClcvUpIT87VCvIXh7GGgLySJiKxe4nqJq0
Y8D9IafIBtfPLHCLRuwK2+3EUlQD3+EBqGorzeIf7HvZkfOuHWvHs6AqZalrSwNhSNzr9lYeFFCy
Yw8OyTQHP27PMj1ZxiyomQODeZorD2DklVGMfdfjztCYm1jRwteyw4DkwdpYa7+A5mphzWfr4UGl
81y1QrjrAHjzBswj+YJi0TFoBYX1v0GyjmGRt+L51k9qq+i00gZmux6pHAuRTyd5BryNZIYiEYOV
c+7jn/lpyQcD0MJrMi4vTKlJCteBCylXSa7duag887NLxEuJv2T8CRKgjWtwFHmCra8pVutDoe8l
WChH/hOyn9cR5IUsHjfPjH5FVKGFvDlghKdXSEO6CvjdrFGNDjkZ/qhDENtvHNUgkGQnvLAqZNcf
HYjxXaBpAlkjhJ4HCQuH/Y4K0MH9Nperlsx9SmBwKWy7bAcZTNksJ0wAnLB/qup5NT/6OvLTak+0
+j3aG3ImCK/ylmYG9YJ+8mAnNefweuiv1bJ3obAQNTtYsNmjOJ/bHkM0giPKRNEItStKSmsHNBSF
5O9xc6V7FdFFh0VcYiE3Krm4ejflqvS3WV96MsCzizvsfzL0Ds0npbg8kt8Kbs5QvO6Xjyjs/xrj
xFap6rRg9M48Xh29J370Xhr2RcRrXkg9O/7xf/eCHrDmCpTPcKAekPkpFiByXPQMAV/QUpn9e1lB
BzO+8ZcOJ8g2gY4M6IO8oCNolqoFVW97cJW40Cl6pnx0HvfQku3WvJ/9doFqSuv0t4xYH4XTo90R
dl+N3OyBSySiz455l/TvC06ju6OoSwnNsuKj3VWE1oo7oVc03BSRIhonPMlMEP/xtSIB8RPgTmMg
ICvGCcWBesH8xvELozWf24smARpR1erT+kyU5OB8vn6HwdGrZYPWRG0GOW5FDZIgBJvtJQ3+0HhR
GLQtw4NjeMKqvsvr6XXKCfdHX7Eo6xG7iFhj1xs5mC7vYUiOXv6tTWyK4B7z2MFiwjHznoJhC9EH
ErwBf5n7nQlM60YpFJ1JhFS1iIlU8QlGW2q/iSTGJaUKvzfwrRON0957lPcK3n2cka2eDGd9WljQ
kBf0u/OgTpEoEkI9DFu9QIO8FsdbZl+qizKbmF0ZFyXNxYE63RRTVChGQPOA3XkfY7Kh51EZuRwC
0s40CJkl4i4BXLVWCFe30HuCRJSyl/awbJExHWv/Z6dv9prEZfETaNakaWtTW1pvRZXAED+shy/g
JtXuBDv4OhQSbEMZhfPnRuKm7Cp8tgRS1GpCvqgPeROHUjQQ9wmstg6+tGNHqD5baXGw5kihQfPV
rgjbGsoA4Qsqz6Qk1flwD0rH14OKCXbJHPAdOusuxmlRsUJE9WYEziYo7EXFPpGyD553kTUpjw3w
yDEQnmOw158H0MyFacQBWtvtpnOdXLBz/JcKaU2UHoD+yY27WcEvuN61TFfeKfI24LZv0KwCH3YB
JJPALucnURlY/XcKf5pfCFJQo2iqeNnhW76zY8p/oEwVrabj35YtAmcfmPgRNNXsBNW7GPAeKaPY
ooK0OfMDiqkfA6uLouxtKYmKDYwOawxxU0QORdtk81heZYHRZQrj/EGoNdrDypApOIsxXix0p+wT
42/Q8TJUL+fKYovyFhJMYa5T6o3BNKi93ZuaZCVLNdDCjbsJDH/ylvaCmmw1q/oMpEnoC9EwzZ0r
7hJuduBtx+YK6I0bGZSfjHKO7FG5X/sGCiBBuSuftJs4dJ7uY+lrKaSL2FEjetnTtHSuLCM9mNyW
NnHEFmfnhPEjEeigPDqhw4Bpdl1XWlGScfhH7/r96j54xcU84zF2/6EXVt7iS5eLgC7Jkd9ibdy6
Cip96aURALYG2zsTbSpPjMM1ej3uI4ZVoEioPR54ETDZ31/D43QkW9dSumlekhrTx1yJnWbjZKBM
eiVbef5pMJnMn4nOvBLHUDpQbQtPdyG3I3w6undo6Fc+IrVjpYJEuJl4BturXakSjNA2IJ2KFOq8
uMdjnQC0/3p7vHUHmPqriOP3zwXc0OuYtWiu/tCdv/xqR9YZUzu3RGmvFuefzlYEvujqYqWaaiG6
IrtPKRhP63SjcjcnYEs5pV2dFldKQ1q4E0Z5EBLROFE2GEIiZyJ3aLes3B9mdn8VHNxh1Yc+usnA
ZfZyCHFDIP0h841MsYtACXFBxBIEqghaKCv2SnbdaZM4ujWKSIv8EqV2gAP8NYQbxLSns2LxN+qR
t51+Sa7y+hQeUWEjfMd0pr9PvhYdvK9AzJXI/IArsrVyDRnBK11XYsZkhgeVMSCQn2R0nPsO2shr
zSNfpaZNLJeE4ISn79RHa2TBjeayKeA1AqyhZ46SbxGm2P0zwD03qShYPWPScWVWa4uazgSX6ZKL
IDEDlG+8DjC/Hl7jB9Cv/a3j04o7rH8KHCSa3EKcbPglciiIWJnerEzomwCMYFvLADLchzlfohA6
GPKFq+Tw1WS6mmIux4HEjsQc/egI0Ea3KrywrnvHfjztVsMo9UIocdCt76ZGmtMNpW6z7458kgUA
P+gI+KQMf88WV3Whqs19wuLdJF9VzmWAB1wVj7eFmyhA6uNtRrOTUfMmigp6uPWAeqy2h54ovjmv
IN4LHWIzSf5Q2wxBah5KfiBeEHvs9NJ7xkHeAybgAhnp3Qabw3TqXi160rFIGjL5QdwZpiynuiSz
NoJygJqjYtfkzpUmI7c3WZ1xxF9TBslfNgeDzoQEWAVYbL8eNleTtY2wui2VijqAmn0vYBGQ97JS
2GX9Un4i3nZgETHGKTAztprlk2Q42bBg3/bfljJ6KZVVb0SxuROYP8xMejlQYwOM5sP7naLy8Obr
6FYGgLJg5U8Lc9zs3MfxjpmiaU+/UuFsd2qD3AWHZzjngezWz52To0R137BfM1GTlxb8Iuhu4rDo
jH/U5D3On0VAnURHgfddio8iFDtWq0BihJrbZKYENCrAjE0z5HFH/cEU7cje/kJ87Ch3SH4Mku3l
8EkTh22/nemxCTlBGBUuOFghH0tvwPttTkxXJqIo3mzFHWxTedEETHbuc7bKe2Bz9Iql/JN6rq+P
y3rzk3e6WVq0ADSCeRly9BUUNTfwN2HFHfv/+cYKmuUWejpWrHJwS9xrNyfjoMBMN3Y23yjvCYqE
YxXDsDh6AqQm7ylgvEezguDdly4OfNdEx0LzIp+Dm2O4pchcMXKfXMlEMQPm88nBca3ahSRU4c+v
h2DnMuXa5kJZfQN6zgdZf2lbzOHIFBgaq5kxmhG7+w4zDqqbPUGOnkwsyvjer2gY3YobWAyjSZPc
D2IEkC/OvZcCm173C1Ltx0Ng7VZvtFJO6yxaRxkePHZo+nTc17i8IQ5IN9qu1T/vwbvsCDHAkmTj
GQUMfD7oFpDvKchyTHM6tsMKWT/b8DzofRwLarCMZIakHwxrQaQplb0OJGOZ99RVrIwapkb5YB7y
YxgctqAUBZghpA5APXf/iooXeY/k5gZKmtQ5RuH8/qf8wBZF4TLLxFXoszz1jAkVSp4wkuwHJxAo
VGrGxDpfOUL4kluFYsIQWJ35y7Rau+3VlKQVtX9r4rM4GNxxO7DeYxw/dfbWU84oVxYrlfd9+O+Y
otYOtVz4TYm6YX35qQNH4a59ljOmBMtASBYBEzm97c8nUGLpCqGE3cn9naGNUnsMSsNiKGRzxSYr
2KV2oovYNF0h47oZ7VbUB6NEyfia9IXh2mJw8JQhsNIT5PyBc9fqCBuLCS7ZtodTKBjgsAP+N45s
6t4gJ76pn802EUJfl2OIIYpPEVmuM/Amv8d/vj+gnLbtb0uhodUm7yQLuTU1lwP2mKvfuDNNPt9M
1no6/BPQ1/zksGn4ybX6tegbb0Mln3Dz3NvdtK2ZqtR5Gh5J9lzN/hcwft/bykyUsN1M72H3Ah3Q
LRZIdVQf6FkKUO3C8IsKzFM+dma46q9mUstns9bVL41X5bD9S64GrrPraG0u0xcl5TfFIsfZUDJr
zT6JvKFOEzxPVURCpqe0G1RNcVQbeIWvG5V1ZdAiKNVz7kGAxOSjCwdn+9Nj2vaYXhCvKbKPk7wC
E29+ga6LFWvrmRpY02+fx69boPebjE7RlaLxjcC63OuYZk1Jnn1F7Us2dCCOc4qCf3C/e0n9T7zI
XvO/DTDdK10eiIqWZstqp6Ttu9BAErYzIlKNyE43AugwQqWSTfsVFYvG4NI6hH7Sa5FS2mIPo8GR
QpvxQwt4Z2mwWt1FE7YrOTW4K5W2Fva9Pg8p1uY/m+BILrLKmqh3NIxfFLnn5CW9chjQA9/eTRcI
KlhszN5a6MZNW3XbHHoDK1+VBICpGPZymLKXIFvXNLYczkoSgPbBKK+5mwgao7I9fABCzfdBIlDZ
b9jsa2Bk/IH1Z8v2qA4Th+2IgmJeelFbss7nJeIj+kLxG/Z2v2cm5KzY+WpD1xdrWhi4dnHLaQiB
DfH1AN8pAXSE805TPNiY/cIQjv1DLqcJq4DGTLkjK6EiIPesYVk10ARBd7nb89E3QEJeBwdEMKeW
OzUqjNoTOmqK6Ydny820d2tS917K0kgIRIwSJmPdnByw9bnvIyjjXCu43w5lXnxv8DktkYOg1sks
lEwA6jMz/dntYF62RrprPdrk2Cd6ifhDEOv3hOO9l1nVz4GwNxNqXgkZcwa+O0d+lNjyLQkyxlLC
rY4mUMcJT0tzVpQ9ELhnnXuS9h0qMu+8b59kAZxwqNFWsOmnu25f5zQQAEYGSjSgAH58GV/JfRbl
D/JcFBosQth6BTE56Mar3fG6c4lFsgN5PJtCWvFwqAFcufGfphznkHkggGCLs4HR2LvW7vwovu/N
+3y11yBpzhaWalDkHj+recR+1257jfMqgIp/mEjH8q1VmFt4e4ezVHxEpskYSR2xcn/obqBnALt5
bEcNGdas7Zx6pDpVdUIRyolrIbObJguV/jwLSJKTTjWylK/4FqbwYNm50tY31jaeOYgU2VotaFF/
p+z/9cg3hb8QIJPXUjjBbD9ziknBJXMXI/jsgXiy/joJdrzAxrwQvgMSnu4/QtzuWq6jV1pPrW70
f0pzEldv8XPa3s0CqApqjjqlhjx6Tngu8Mhsy9vosYKnxpj3sP+QX7E1V/jDAdwPA3lqIYsypSVD
J5xGx6SH7kbEtNPiAque1XpUvCLzMBBOYJM7QDvxTWUdUdXVbJi/XqoRYEaK+X2TxV+Ko2j4BXuu
bUEQDOZ6MaDACi+BMuj3+lIj9+ZmaM5I+VS/dABYjiz/W40x5OXtvvMd6R6OLyKSQHo8BzrEkTdA
LPMGlUoyJLPwYILLcvsM+UURcc11/i6F920ql3EFyuoZvQBYPpX5XsvA7l4ADQnX0i6RRHFkWRqY
+EyTypbehXBuyjNy1jq4fWA3CVhx57bdJY+cAYputDEmPQ7iHu/KT+aolG3eCyHu0EiyAZpuLmXb
JU4NRu4QClynAn0IQATsSprGjVK/tuEZcTLwgRY78l97huFo0mApFZqIFSuPbaZeId/c8vajZn0J
bn+x7LMVXRDalkYw1On6GgvkXj+DA5ymY5pfsigArS2b1TIGVG9F+1zSHmMspflSNyjEBdBy2QQL
xcju4T2fcKjJN6y6/B9E6uOP8TZT35ykAjbp9L9xK2yKvC5WBFKqPQyYvRYnVxcdMsMUUFS8zBFX
cMDmhGb2NUrKZlNM/wssS58BMqg0n69pyGkY+p+Fr6WYpZi1WsrFqsT1ttax7kbGZS+D9v7zd8YH
4ZH9DCUY7Tn3G6i5HpmaiLB1egMIuWtdmgwUzaTtJ4gGaNyMA/vA5zDPV8EN/01IUNhxEx0jV1EN
Z9uDuJ96/kj12XTxpnlMguZ9Ei/OAjJGHaLjAyS6JSb0PuCymxAf2gOFp3G4wMHA+hOyh5u+SclH
ULhhBuAGRdmhMYsIi6+ydOj7jQdClB8ui5A468Vofr0AaEtfhHqCyz3WdfdfabUWY8IHlSZKZPa6
iGm2U2guBRXM8bl+OangMioHmr/yHpqSypn+PaxtDUk49jbU9/WGMHTouEHQjl8qLsiIWIaKzpmL
nifAIDkrQNeYL6bX1ZTJPnnRQshxL9SHsh6th5wptO3+kIujC4U+B9SeNFHnDIfr1NcIzfIODzmC
PBrV8VY8ELRt62qdk7XWWsE2qHOoq1J2cJA02jHLw1gF3P/WhYvbtvQPAA7WWG9900Nzw1wu3h3v
a+dlsJKSz5Kzp9Hh6qcGimmAIgPNA5JaQn0KZHV8vz9vA/q8dYbzGQ9Wlo3/Cvkf2EOF84IlyWnd
QpxM6MsBfjkpaBv7VfTaYndWmjBrXb5UWi6ARMVQvxdRg4FLTWSzbHTp7iuhzPOylekR8LuTVP3e
9tVMgc16rmB5R/0hChuHu0clUPg3gKwrgSqP7viVG9a4QoDHjjn/2U70bh0TDmj7ziUmJ3WJ/Rby
AnZUsqk/SD5xAL37CaxJsVznvqWtJopvueLOcAoa5LF4ydjUkMV8f9+Pe017nTC2D3ZtjEHtjm0G
5imscKrmuS1bb5Z6grasyvRoJD641V3YQ+HjJa/eM3rwv8abUKqHRBxBTtx+eCYmqJQtN79vP8Ow
bwwlHbRCxZaCxZEYGFdLzAE42J/UMdzq5iIS7dDGAeTDGzZXVgd3CsyflTFZqzn3FvQrBNOjJMEb
jCPyRWhbHltWJQAGsGPjSQl+IayY66qPDiHhnwJ4yqo9eiylNqdZmcv+Oz6k0g0mc1Zyt4ZrD6OM
bMRdMLz9eKPwlf8yCtH9q2dGNSFg/uaaxJvgiRsiPba0vSzYFBLiXRXZFAwRUz+2yl69zGvchOL5
Sf3cXbnJwLO7pngqNMToUu9Xw5m6ryVvhHUSBWmSey0HyGAP0Pjr46eaW6zY+7YpH0h5/u77GmU7
zTAtOq/LcKPc7QW43KfB1g9cA/VH0mRxoDkUu45C7z4ZDdgyR5tSINv/1WhhlajtdWgAtJ+9rb/F
rxAMyio4AvQmbWEeGOwiqE0S3H5wC26yerfDWgVWztY4oqVSigEL15SieRsEB+y6Jg10bfz/Ho8d
KC2ghSMS1I2XFBjuyv+mi/F31WFh2dvQ+1T4WxaHDekSxEVDb39ADjrNnqKKsUE3HalZbC+I38S6
hbw0SI+a3x4ZS1xB94exVVBMZbZ7pKh324wyuQ1AqFAmLk8A0DKxR90He7aDlzi9lrSSYdAVNRS0
BUJI1m0yCu2AwTXlsWFnQ9aGPpQwrHdolyUA+O12U1niZdQ8XZcSyWn0wysXsdL575XpbOLdTUzz
Vvu19A7BU6Pv+k636k8OGr+dlpahjg9EWCJAp30Sg6WjD9zCuE7gbPH7uIjzyAmrpXXAW3kBzPVl
3WCp/bdjg2m/9JvDx4KIBzOwd7mr9PDu+UgGp3ir5aZB47R+eWmkSKl7XKNuhGMrM2otSA8Bg1P9
NAV/X4J4TZN/8qmsMq2pVHrzuNnvm64q7Jko4DeLNpSTX3A6J2B+leWcOLfH66kFSByEoNDpRHsu
UFVV8X3dC9Y6T9pzJnFLkdEx3gAyElytwg6O//N+IWpO6L7zPnW56gDjfyN5Nhe+oCKUu9z/v/fh
LpLy/yKrJof42pDCpGWBfT2ZoFIpSoFaVFqCkw4y5hJJsRVPsiRl58E64RrDiSlNp30XPrbLhMlo
0QHvI9yODY7C30n9h+tzob87qyl9ycyDy+jcnWdIMODyf8IgxLkrFH8H5r5N86Hm+y7fyF9OPzZR
AR5bbTJJNsxoVQxsez2/mQv0Z6W7dwK04QWeVMiQQAjiv9TrvGJP45/y2+LoIPBRur38KPjHOtIE
VAXVWPFFdrAF8P2jZUsg6e0vDhHHX8ALh5rDDaTLqgozpxNKReR++1VEF5kVGU5HKGEyhWa7vHek
LdmG55kaWOv2GU0CjxagQuT/b83MgYc8t/rxblQfhfL3ruZmdSeH1mLTi6ascBsplYuFo2xfEagX
/bt+g6TcBoTp4TvbCzxqHoznccmu000lvBz4UA0vr61Clfocn6/rOnU2ztTMgqqYYLpcLxVOWA6X
EADRuJUyNnoGaBPB5fxi758yzVwzll3uqspHf56XJv70qjVqrH4i7zDWu5hFEWAX3hYBWC/Ndb0Z
t9ibUkgxj9xR6kYSpdNUmhKCbescgXxEJAeRBsCPg9TKFj6CCyH1ng/jWgJ5oC55eZdZH0l7t/zl
j6slO2ik5Uk6yiawdy7JiWgTdQ0MFf3mQRt1KewBO+6XidjFYXVrBGRID62g4za8HuAGrmdChDgP
P284P7gI+u6QLW8hmsq4lbrfkkxSXb77LdrxWn86STeA65jb4qopzddmIjplbg6LxqDiskz3hhvS
mUo9Q0k+OwobTr+OtOkGZSfbF4+8ZlP5s2ieFJZWNSXNnA0kZEV1DP9Bg4iHFaVHT8oazAYBodm7
t0UcNSr0fXwDhpBgUxPca6FRYhOIHUSdnf4PwV4Q6kJ3Rgt7N7e4yRLJhgaEVFi5wEIJj6sYiUx3
HxHluKhmd5PAOnMMTaQniR/2BulR0FJCMlG6FwVCLoB4tDt9hqX3m+MkDKIzpMPkp4i7cx1FMeL6
dZ1VjNVAY6RF1cYzZLrgXG4Icu8YmTXinx2BGgUDbxXJJ+xXwNfylAI6obZWwkRokp8EVHl5PgGu
hEUNDbAE+Jxot8rtkPPHSqGnSeaghEFgAHFmpOQvY7+Ogz37tFM0C/rwAwTG2DUwmbiUMvpPtbbg
ynk11gz5wV7qg3N1xsYlkL9EO8t7dNOQpAUhrbxOwORDXMk/WmqzXCCIfpyQVcrVHhlpYevFp+5A
6NVS1OeB6olAvXFffBJIras0w5bc0q7zU2nSw0AqP2dt+xajhRclXaWrHhmpropzM4DP6oOtv8xj
f98ZCunOvKbiIqGqmNOy8wENv+yi2JRjacix7GgjUpgbUSC9jiH1WpNf2RX91oY68I2C49rY0/zA
XnKSrWhAAqPT43K4FZzVGxt5XOYQ2ic5La/EBK8Rz/Q+qWLQL7tHkGfm6qcSy+hVpE5LMAxYk+nc
whXPTscctPgDN6HBo4/gmQiOatdMOqEc6UoPqdMStErhvxPrTPRThogrpRYVtvI+85x6M7aNLQhO
cu97OKEApPwzAftc8zL9pqfHTDqG9NJ8ueh2lY4TrIPwHB/QiNkRYQ7cmn0VeUgN7u47PPDDrZe6
9c7yrdWeUJjixD4amHdDhXNeKuMMBfuDvFgxAkmRdQMjLoJI1ZbVoAu0AfaVo7rli8QbuBUv/gRi
ApP7H2cVVtVjOYEHPqO/kMBN99Jp3iyi+l082ZYKhqzLIsAySysKEyTqNwWu3MBSiO6CDUJdPYWm
WO1jRy/Zsuqqm3Oit4Jh3300Av3itTy4t5u4uwSm/gYLlYlI87Z0hIcfSJQrdKNj8MyKgJuWuq47
JW8vJcxfsCewfxr3TU4rbZg03vclwf5Z1YZG6rlL/egJqYgSmIKZbmmC32zYA85PWepw5o5bNPII
WR+tjOsUMR2SsxkH7vqNIG4eN9bpbKnzRtWV07lX5m61rqkLBijjgDeG8Tz2fScm6UBdxlPtrGoD
te42Vynmn5j7uLDjGowjOZrCcwLmxxNCsGRRPZpeguv3eU5HpQuIogWLi/z3RWuIav9KKs76+wIP
9r4qxXpFyj9pDkEp8X9wBiGVzowJZONS4qv/QfnfEJz9NXc7ciyw3pMaPJCDB8audGxY5kVyxHoY
BvkbPDVNizbTf5Y+WMPpqrs11G4/dc1wMJrlCCzgWNodAD9Gv1JUc/DGpkTfPd1LTo3SsdH9Coyh
0pGJg8xxnwscYTzNK2Sw59qZAQf9e8GIBmPB2Allb1RX+rGv/sfhWo82/zrsKZM9vrRHnX6VrOvF
DXC62SxOtM3Ve+t/dFulpZu6tKpr4/bPXSaL8NJzicCuh10LNMIj82GL3AjTkdsLgdB2tIRCv90I
gZOyIqoDHvZSMCH+ELhqDfWK+7OFe+XQygKGlm6GA9ntO3HnRQEQMa1saixM44XWBHlRdtGJcw3F
AtJnKJ923l6Y60fkY1RE5KRE37IuZpfX527y78QZjHe4WryRYNqzA7AKGbiKk+kNclKmJAmejrKs
0Dg88pIpEwD6TVEFWUts0TFRXVgpmVymmGYDzYZTyXZ9gwOCcFQkkNzk4xCstp2RKJMXQEiLPICl
mIAa319iZk+nuns+oie6//FvlWapfQXjIAMN3503cKN0O7HOBrzJFnHkfSnXbjQyPhVNGq1KgqLG
w5CPD/x7hopy2pfxUsXZza7awsurbAcWg0KzxiqICqq28K/EVrWm2j7oJGi5BXWGhrlQ9LNtiHlN
U+mwyNH0bqwnsxxn+bl6bdUVK8UAUI6xnjMNS+XQrGX7Z4MObRcOa5l3SqvHD7XVISKMQfX8W4An
YvZveLJVzxQcYQP1MrucTD6CrPNCY2VqvDeHKY5UpMpd3w3+ic+/7r3VwBcy1/EDagGlJE8JShov
LBnyzOBBmR5MSg2cEEwvaTRc1VL8Rpceuw2XULu7jEVP14WyCRie5GtK3VpY6/QW4oS7/ahNYQMJ
HCLDGHSn1Zb4EQirEssjlNd/Jzi6WNAGakFSrd06iIokVcyJuuJK0U4wjVHgfmdqTi5IZ5Y8Raj1
tIpsGb7J57qqPlZUaK1oQFKtAkehjFnXvFGsTo45RUDZu3XRilMXyLEPwjHvQ6QzXjdhPIFyujVV
D6zkekcbuKHOhJVS/hlV4QW9LvFwpnPACb4T/fg3DCW7D8HF7EuKk7HTpYoXCkVmjHFNJkO5ORPY
i7c4RwhDdbLq0pAoV3pzubbUBjEnjE6Ki4s21bMl73ZOrbL/XhRnnuVvJxKwju/19AJSn7loeV36
ybgIevIECJ8O5UdCVs5jzzoVdVkHv4VqXVNeyw6iu9K+pH7Sq/y8S/uIdYK31gRQN6xi6fZ6uXVC
bI/+Edv25R+XShD5wPunbaU1yrItdSKe2fcarqtdmthPZejVp/TNr/VOsL3SbxsWF4p/r+EoUP6o
eiquMQYGVgqHXoKnrR9KKYZjdDbpa+6edEvmrU2hJZD+TATkBBvo2qmTr9Oq+0xFYj1rAjNxJYZH
MOUUtYGPoOgl6xHJCR2U5mkwkSw8woVOeHJ+1vu7UHwv2zjlCThpl6EpNkOEJ1UuI5kndhvp7ftn
cG4h6Qz7H6ApTV4zHOaKtOFljTcUJYJWrDQ35hforMxLyhh/YfPzJfpD0zL2TVvhRBNMFr5BmGNa
B8wcvqVA2fl/2uYothdwZnT6EvrGTgpze27XmT7ezsCM1qJQYWq3KSxTBDrHhZPNrPYIWHeCJ16w
tVgLjsjI6+0xXj1W9rzZCbt4WRNNFdnBfSrX9Bled1+DH2oueEyoTfMjhlh5d7Cx7BNDoFB5g0Kw
9eMPLm7RgGfHkVvqAETl3hUwtqfdwoNegXbIjzt4P3qPM1XWHQZe8C4IRsCScrJZEu2zQ3EaNvaN
hs7eHNliQ9HcCk0pR/zD1bEJ2UBTnO8Gs9qgf7AUlZIGAP8jv7sKYS2XZvzEF8bOYBsM0VhhWcZr
u4/0PdAcwLSxbWzhRl83fuUzlOsCmoMF1nY+e0f0SMZNAoQ5n+KRgLXu2uZF0oniMIaqFX0YwaDl
vZkUHAycDMhnF/BK85ST440mVRVZEOYig7NatffJd0+1KifFK67NkWu7cxGTTSdL+mSlW9kIV1se
t9zMY2ZxlK5Jd2SgLj28943f2jzUQyfIoBfbiCVLJJENwxErwK3lrICqCt0GD61+0H+p7b/KlT7b
7M9yXurk9OPqy8IEaKvecq0rtvgu5C1KMS3vWv0IQxxKSvCp/tfe/cDrJ4F6L8MzJkzo3ez74q1a
pW9z3pEufYICKKbcYD1GpZJQ477A5gZWmVsFHtHFAoSkUNBoUhjj2OsE0SY2Wl9AOsZq833IQtVE
gqc6K6ePw2RrK7Lkj08/45cq0WSVwd2wOo2W3WKPC8SJ4hczFjsFBANuKoqEvHGQnd3TNw2vr7kK
XYT8E5EhyhPvGRsr3Tu6Im+2gDXFPf/5FsZBJJNtql8r2xNF2Zy/BTYkmH+ysJoT/Rb0S3xQfT/+
IZhFW7LbuM0RPaiTfY0BKBKr1xQpAh35pWRAaGF26VeqT01k/GJ3iLRbJce/y4GgPXZc7SwcfpvQ
aFqPMheGCaWR+BqIFN9QoPichGxRv8sX1V5y80P+3yjIutlYk9vVpk4XyhzjFNf0L5CxgULIErik
9FGPY/MgyUb3HqpqTKBPL7aIq38HS+libmQsXSrDDo7HZz+AwInFf2XnOLUJqgFwniPQHhLZikpO
2oWbnzFl4z60eg9G4Kp3HS10focWr6jdTSxE2hOl8ISmxo0cfbqREIqcWTj5qMv1YY8RzSlMUboG
MxOlc6XcyEt2XqKon8nvSHf4UkZwe/tvifQdOXwj/KqTaA0Zu9Pddf1NtNznJB0tB+5k9o5k/TLz
/IZEreNq0gK8pfJFvx9e8SeB8BpG3rWIuE/IXn5ZuTpAtl9PDrZpz8KZ1xC0d6UGGhkCNEl5k3HU
0H0OqYlkyi1LzSkweOY7/04sKZPuW6UfQq7mzcEIfQlyHBrs1FDkkKSf0u9n272wvTMhjJub3CXs
OkLlYEfuA9dyyMnf26jEi3e8fLUyQFXoRJAePjnFXk6Fli1ua28+w3+csZIAoYZH0MkbTWT3v/XZ
7xaRBDX16RXp3ZOhZTD41u/IdHbSFJMKXEpUG0CiW4ngEHpb4OtcA1txl8OGcOYRSgeyh0hjsl0s
2y73/JoJkl4eME8HrWPSc8uC8zl/EeaNn5Dk6x0JkofmScjjB2DU26wnun5Ivx7xdr1sh7a7LOBu
6uTBClwKi1hq4FXwFAU7FWMYP16tKw1hBzhy5UJorZUwwdw8rz9ugTvRRM4sg0MYShtcLiEx8r9w
ziV4dG6eMAGZSu8a/rHmjtWgICEliLOJrs5fcbTyxDHFPPN5i1s5vVNUj9YtgnFCHEmwMQzczXgT
AVkMnUZEcXwR1OHdh7BA2PxEaEtcwXRQWJ43ogz+tUEGQd2XD9UJ7Ca3piGpdOA4VH9t3Ifj0Ooc
ru7IltXttbRPFmqKvM5codPHQmpE4pqNJgYqB6EApo5V8nNygTI5WBOJtNyHOJAyVPsrHlg4Sulm
OylHKL4B9YE0+FLU1f8sNrfZS8CBM1XPrxPCv7/SIRGBFPAnsVleuU0g/hFzapHbaaR930EnKSd8
XOZIeC9ckkNEih1iJxsBv3RRlfXzUUeyogcvycY8XnXB7au/d8XpWrHS4biQYiude9oeurRx8RK4
pJ4e8CSPRFIBz255td5Cpc8cw3U2mJjxpp3AnTXEst832Ht0KCdZldkXHAiwA/DQdb+3gbF5J/UT
HZE9XNAaFox4/Hl2gg8pnC6mE6CWhjWD0Iz73sMlSxw8g2Br8xFU3sbwrVgkRFTiGzxwmgTBIgNv
u01sQ9hab6F2IHZSpGLxFkCvFPMGAkXmemOUX8+XXl6PfSsvEhgdq4HeJBWT72+Np3kuDt3lqgrA
CU1c7529J3UN+/6/WvOr71xGa0REGbQaHJBPPUZqvHd+XbqmpB1avVO23JFTY7btvvs+oY9FpuN/
qgli4GwQ96Yw+6PalFegquO3IFSIGl7DB6KGZHsNnWppkCTILPMr+D75O9qje6sAYX0A2S10xosF
lBN6YRqIDMDJKMh3VO5+Z0b/pT2jzEWKfLOvVjgIS5VNKuz7xISCcSF6O5/HZmJz7O1y4t9u4mMP
do1a+EpjDdjQ6houDY97omGf1CqASzS8VAdWXUcg/na43y7IijpCg9KMtH5adaF5rd8lT1+blmjK
DVaaQAa8ELifG6w/Pwsxj9NqIXCD5O8coYZLvV4X7wdopLUHu7uNqK7HA2aaUCAhUSatUYgjrzp7
MyC1sRCJE+OAe1mEREif0Is9Nf5Ky96gw1rYtg0s2spkFfKo8tfTszctYWT5N2p4Fd3J1x9lYIcE
rzVhc60kJBQ5kwoIKOBDkIXqJJ6UDrKcStedPYD5szlzH9e3Gi+3ilO1AdlAZyvCoWFREdgR2CFB
iMPEBNxSXIqeSuuypINFLIcB95gVvOz1oZD3CwtWtEprrWA+1/LaG+BFnNPdjR/qBxFMXCvPtisX
QMAryajFFMlxdcHcufXyvYieK2BmDTELxdPFot7WA6KtmqTobunlFcjJBtt6gUMEca0nKGAjVqcN
Mue4j/bBiAhv/MorwnJGDm1Se/FXBJoF7Cf9+sZAO5Lo0ARQ7jV2tLThW/IZ8YsTYj2/vC5XvNjm
Eb4kbo5bcpDNC48K0Ecrybk0Zsueq4B39lz/CIxXg9tX+0tgWv+Hf9YfFXFdZG1dnqvnpE7/zllQ
7NjWcLEpwKf4ShIWR/SEkVrbjrsUTaEe8qzyeDNOMbSzqZW6A1fKWWijw1vL9gxW9+KnCd8Xj/p0
sfHA782/bHSKQ5Ks4/KJ9f7t8z3V+KD8g7AfRmOQos7HK2X0FHT4F3luRzD/v0zbJSslUn04f3wX
OxRLsoui3hm6e4CdiKbxnblKCkofU7D6pw/cwMVUUpipo6w+49Cx9OEy0WrP+5TokEiZhXcqj5S6
ufifP6BZj6bs+z1Ata8q4BmJi1+LsyFUF1iKpNgvmPOjeRcR1rl775D6dyVrKBNT5+84xDRBkvB8
K54Wg678SVRKtVzNd90IFUYhPdSB+QBmqyNvULPZ1VvJ1yBeAgIMZGnPfLVc8xlfKURbq9mnPMUB
Wizc8W7rSYFGHVLqBI4eqkuQeysE/TJ6aM5Aca3KYBZKC8ZQcWkzDjVowl9U9iRMaep8PVHu6YPc
mk9Dc78XBwpD9r30b+mhewW/8Reer/ewYKnWaoNNy/hSdH51UynMDd3KXfgY0dTcWgU1oss0xL6Q
zlSfRn14BrnYlBbg63JkR1OF332c6WNbpSsdiePCs0O4UqZPjq9nh7rAMZfI2woFNRVS7ZrwG9cY
FNx9gecbp8TznpNcJa25190uFs9zTAC7KL9oQ6/ZVIA3Xm9k9SlW26BHoYAOaXrSIhXY/4SFeVop
/0EqWJntD7FuQOhI2HmUMHydneQD3n1KJa7pBmIDDL8v+K91tbhaOQWpxDBn2yl7hM/RjVCqFUl+
7IvW490UTuNaSqbnha9ifD9Nsaj5PlCqKcdsU220ncod9q/7A42/v3RtHc4ThQKvWl3KRbv2P1KH
VoddVs2d+NYlV4O0gjJ0DywbuCcqTL4lb+U6sIG/Bbx3c0UKu1/TCZqKHWvVFzAFvHRpzkWUqQUS
37kXWAGKs7cQRyv76ME+cJ217S6MsV/ku8Pfq67lO+8ialwmiSl9RHKpUJ7TFALNED5E5HV1oJlt
xyJYb5L7NfMIZF17LYrMg0b1Et5aO4uBOcHFomswawJfdJ3qJzMCvkoNhGNoFEMplKOmcdnZGxUH
O43jLNRjqtFT9eZ2SE9gE4Pxap1+7mLyROMMQ5wtf0kKxAAbozgPiIWJBBCwqyUCjn//Ym5sXV/t
pgHXJM+Qb2AmQuzUQB7gYeQY2OUED44WzDuitFlkS3s+A0OPaxLE+meRoo5bCWs2kSbELR9qqU92
N1c+ZmJLOlzbiE4bMzPqtHxzJpb3bDteAcjwT1KnWiNPHK7r7MYBwZGYeGXlqDh9pAlaCvVZA1sl
gr2P0FN4bIxoXZ65iMj/lX+wufOwSEg/TEHBzP858/v6RA5oFtg+45Fep6WFSivAZFs+kNKzSRW1
EsbkK4c/4HgsJ0rLKax5CYf4scxp2sSno6Ph5DUb0CZ6sBcnfGTWlyEhPUzxFs3dfTJwoyjqKoxe
fdCvXAWOztsu2U0tc80dkFMuUAlHPpoYjwRTUKHseRkwp1L5m3jSKYeg/8TEGaPND7CnUCqJZPmG
suhLcCthpxkgtNIr4b2bjJeUGlgME29/w6vgW8WMdNtNrF+cwWWXZPkgBN3ost+WmJF7iyyy8bwW
ebv+M7MCrctCQTnKvp6sFdNzPEZrF2rsihjTCbi+aRyMl/BbWRbVY6Ii9Cjvx4C7ZL2dNeOYd7a7
3HCzx8d06n9QYbCC4iKocuX8klYvZmH2UxCYwC+6P2sWG42Z9OlqT05fjHZ3J/COaNuUqABJQBE2
/ahPQ10OiKT18IGJy6AD6TcKBcaGHh88GwJ37W6KMp7O8gpjWlMFaYoRhzjgqqgW4xS9+0BHl1Ei
KskUlgon6fWC/zIpI45hnF6t7IzXJ7NfRlLgCa8lSjFwOY6UiVJ3MH/80ZG29a/FHkcpJMHtmv8F
GCkT8DHwgR/WNKc0xuaQtgHoskP9PCkR65fUIXminCFbYtLLBe2pTsGP28ND/bRreo7Lwg9IufUD
XW/FW57WCl/RPg0W7AKeEqrsSzH5DTOQZTGFYqo7UWtPBCjOU+KzZN3NnXWlczk3QWsX7ptrwi8m
ngtMguETgPxWeHabWl2FkY/JbPAr3VaPnT9EnSBkMmPYgf+Y0JO71UBjoyM6k1Q1pcREF3Tawq33
GyDnfqnaQcopeiyPVUMZDRegzwkc7fD/Fbrp+JjWA+rOcDinV0RVp8pA5ET5ZUW3kUYnoBlv6T+j
/eOC1ebBRkcQpJmV+2FONKuOE2bYQYy88S7R4c7G25S7lDTVjS3K16QKegimEvz5pxllvJhgKcY6
a7Myc9+8Y+Vq2/R7mD5aWAGMHeDEBvv8CunvQAN5OO+y3M12eljJYJWKaxf/29GTtgDh9MVU7APD
UZNiOq689K4IRzGjFoUYYe/xXV98wNEZbzIRoSRGcFwB85/Y/u/CaeXgJ76boFhCJD/J65jzKxcG
Jtadbswl9LnJ33r83y6IyfeVlvIOY1ZKZe/QHwBMgZ8EF7gJBoGD5Q1VfCmxfhHVJkaNC1sMZU/j
Jw/h2XoYllT5Gcmml7BZFGHM7LsPILQ5u47EhcwHX5uA4V0BPtvtMmUK0L1k2GDlStIE1ODQ8vAY
7JvzEz4mb9OpiKO3jrKcdQjat3WwPPGAQgfXt2OMnhO8OUfxym1YvWFfHcHsT0Y7rVml8mijbr0X
v9Q63cdu9ecVMbnu/9cPr8Ql6FJjctzTCq/80ozdvcWUqJfKfcBYve5WZGSPWRsCTyvqaksQugSh
T8zoESlxVMbRYmljowRmYSa+7HlNvkYuYQind9TBf0OJTGpltbhyyQQgjcUOmvXzRJ+RVVfRL/dS
WtqY/V2zXCx6BAmZc4Sz5hW2GJgqWsNIizzgZy8VEYp5NguNa5H0QEpi0WVtf4gta3MelY7w925B
CBgqqz3KCcZltUsFxsehWjvcxWkzz90dtPUehvCGVOwe3FSl/fRjqLLgXz+w5NtRbgNhBjgOy5YI
kLI7lvkT6818/SHo6G2bwBRRpehhmj2SCu6wDyNrh7zM9ASXLio6ctsXRdRt+rYtb0/ocIqk0Vh0
XZW0+zuo+quriQ3gl//yS8jLRxb2HQvlKdeSrPphGavBx2WD5SC87ezh/bvUnn12JYVICcrqRqHK
gVSek4FAYGhSOjZ1bTURRm9aOBpFaW9aa42HTVI0o7fbcovfDGDtg3QntwmxhRKbc79glVtOME76
1Xk426P17eTIHXXJnZ1nTM43vj6rPC63p3AhGwOsRjfw4l0/7PlyPON79JtnW+uCrgH3aIoB+a2T
Jy1wp8w/soocsIRceBr0r9s3sTSSbDYIuZGEWjcLCUBMOG7NGKTFha03PosTa6RsXT8RQ203sTvl
1RrvRFGKL/JTu2T+dk2njghcwHoiSvbTwj7dFSaxjTeuWNjC9yOQvH1FYxCLqCo3a/LcFxjdzFg4
EsrR8CHBzCElmZGlz+GI+rxAca1bR1n6Bp1BA2dPgq8eQujpHzebWoUIrwZ6eizbOmDEEgQ3MsLp
dDNNw+sI+q9q1NAK+DpPcONXUJ9c5L1ZzxkHjVJBcQmrFuOTIfNPXnZp2qfRERidsII7sY61hGjy
QWKx61FFqyWtW3cbfii3FaNnAcTU4IT6W7UWnZTb9cGfVldQBooWibhCqbz0dst9fzcfSX9+Saej
yhzXcPchLU/GlD1BD2Sd0q5/ygscnGdlvGt4QyQ19+zc3MMx5KVwRxhA8TVUgAx3JTmr+c+s0maG
zokxBO4EMSBQ407REegDmBwjyHqRxAb5o7/yBIqFjKJEk8mjVfucA6wmfNoRrxLBUkKeEdokkirA
zuX+idXiAwakBVG88DjAOKFDxLa68akYVuwDOrFII1hZb9ShNQcplxgA4nL9luLLIl29zZFPd5B9
L7xk86iVRQ8IRAZxe+zLaThqi/erarU0jb2BnHUjLY42r2GUdmUTFnYRfTabVUg9BfaEg/bSC8bH
i6qSNCqjuInWts9K0InZ6354MhbAuWOBUyGFhP3ftyxr/fy2SYUWiKKvSM3gKnhlgFHANroELZD6
Ihr3MrFgy3cysKsThsyECtIFej5BIwMhNg/5L3TEVmjfqXTiGn4sKFVkZ13MX9i7oIPYxrq/tpT+
hll1pIcbJdTt9hrn5zpLAuAFvD/53hC3cNfmYRrzkW7hbE4R5P+/9CoE2ZeNWLFG10sEDYgGFir+
qXYceyGbRk+EMPzmrb3lPMEIc5ueDgTrcO8coZv9kOdTz/MdfdCQ8WhBMvPfSgN1Vrm+siQCYSEy
8F76IsJH/c1hxBqjuXrw7rb5duo4OtYvS9FctIwQmnPMDF17el/ulZ8IUsmXAgp75c6toV9DJ0Ke
W0qyEoJ77dm2pJsGH6+PAvgKuhjomgDsw5mpEdCMUUL+VFYiZyq7wRNuWmDqDn+2ON6V7Gy0Wex1
6jF1AO8Dd+pFBDSkrlYuOO+Qwlm7Vo0c6e4LYMoWeap7DEfLWswbMp3waruqXIRFzMYhRyo2oZgK
PTAZAopPehKVGd49rkROLnF1N0XtJHBNs4xHu1wLQTTu6/da7eZsRSk+3TgrmlqkTaV/Y3sXXRRB
DsaEMY6M34uQ2XzA61TKUI7/s2L1vBDBjA6PcUBFyPWD3QgBPn6GoUOcd3OTvbArwo8C4/7G52dp
4wuN8Gs4/HbeM69NJyGdsEOhANbSnEwwOLjrXSew3XnniWqRdOFatnvFGgWr15JXPXRvK+KoEDj0
z7LuNQ7VGAa+j3XKX9ZkAIRtNP/Z4rsKF1bl8hl5NUWftxL6VfBKtj461P487ejf3ilIieNe+JJu
qUn+9ytOexlnCPiH86hqYLyk4O/OA16NTLnh+01XHYlf6MrFI4PIQXBUHzjauSoxAuRRU41V9CeZ
xkdk83Kp9P+aJAYcGyt2ygO1jO4P8DfMg9knRmwr1vK24J3rKFS6cLVTYCVbbHfgboRhjdzyW747
FEW3Ki3/WmbVv1bBNYuX8P6ZazrKMKSSApAZThHsLVw/6QjIdrbxjCU3s0Rm+oj2I8K5vml4WBd7
2ioFAQGAvmSBCCubkExZ70MpX8sU75LXLbKm01MGBt4yCOCz6Kw5zsSKnEdHjgYhrLvHdoY8e5la
F2JOrYdfBy+LHN4TNA58lmHMzZ6xOO9DpZRwyQ0VaCUxDTjPBj9/zeb2G/hwcAcxLYUmaQ7jaSuh
R7RpmBzhTO5PHGAZEcnBh02NWnftot2nLJ+UX+5534gEroMyNnWrDOBxUmJCaKTur8pTCSweEXgT
nbHc2DTrGzvL6zuAyziRJXO1WIEn5J1RHqdLS7V6s1An582E960CwMLj/4NKOtq16uqF7aT5A8XJ
1EzmYCG5kidpFQNh5PJ3KqrFwyqTH9LW+nCXWFZpK1Jnjk0O7C99L6uD5K2qMDF76E1CzD1pDVRb
j3qKDmuQEwzMIjIcNxHannHvTkxDoSUNAig1c4Y3HshiRk6eEDmVela4j9rDdiczKkeYgU9sFkRX
7sWZmNJuJUISFxGyRwep9FaWwqDgXaIbeOWkQwhRYmis9rQfPLbLoJA8QjiOVJ+HYl8Ck8M4G1FW
ncoG5vSN+SXNYKLAFIB8nGVSa5oJwnT/2N5/6+OcPghdvOL1UlMy0YiXtxSQAGMvfwn4s0Yinrnk
mH7527bEUf/FtbZ2PTXqkNHIAotoqytzLqU9M0HWMbqecMZzaTJIjR+6elCQ8DnTOYgdLYZ6TP/2
x0YvgqNaYxtg4EsxW5eJxJw1kutcv4pGY+fkLX01gD4vyb8Vrfhuu0zY0K/4tWhPkPBXeErCYtvp
pXnj7q9EDwUk56NlUFXJQm3W3oU7LgYbTTgeQjgRpUSgL7RHVKTp0T3T7Iizsz//MZBEXB10D8N0
e3nguamUXnahLmc9Jc3Jrd1y+vy+hJ9HOVG25EcLT3SrxkE+EjtE6pbJJMM+moWDP1LLKhAC5q8z
05eAyqeXs52sitK1+j6vuyuwSPpJ/A8OGAtzNuzlcdEufAs40ySUKoOCIZlVst4OT3RbSMgh6Cl/
oREGHyhthqKNyZLbjs9i64KzAiNIqK7VWWC291a0TNj8/+hxvSpU1XTuQwudyGhvaIKZkhAmHrvR
2Tl/DiiHHOtg7w5Oeo3CR74SLC7oIr9UxZincbmSx6BtAeTldHOMJW2jM91j59WPAhdZ2GHdFf2H
IzDIpqTUL+fJW3TylRleJfCdS7f8YdWYLj7F4hZdolXMZsXcN4tv1fYV10VHpNsO/POPV02x0H1U
owiSbGkFmBqF0ozhBZVGe2wzm1668SYgLHwLocmKZfrf7d/hVU5u15gpKSQBoH+DBt6PV+aYmv1C
z6Zk76XxQq9SAZ6m25ppQA1+l1nuDHiFhpePjmwNGps11uhfcT4uxVraTCchplO3Gwj/y5zC/k4D
DV10YDB47rf5Jtd4hbXGr6/IpciOkiEkO11u0tUvB/gs5iqLiv+w9Yxr3eNwernbSSPWJ+YnLUyQ
otYG5SlQ2TXpVFoGPEFCHDiGXHC7g1pr4vyURqXYGn3FGU3V9KoN+F1zUoGLnTdg6DApykQgxZuZ
WDW4JzqCApcV/F774FIryRc+xdDgpVS6GMpZRgcfA7E4tXFubhcaWDLVm1PNTTHtZ/woi1zvkj9S
+HML8Uk24FcWRWCV2GKCjsIVva+V1IIzUaZ3s/5Ow+YwdP2mhYJXqItsYeJunITOzmvutqkvQQCa
bKJO+Td7YT696OxizMMTSM0snX+BeY80L28OJX+NxyjInG/rMs+siH4ZieiQ9tPnTnESU3KS7SBX
ZDxMYuYUyILwNINJcHRNN2nHG0s3v0ZJSu4Xu0R+KBg6wSjU9P7mqe1b4YaiFi6rYSFvayAilql/
cVVPDzdWDpscwC57rv/SVkLmvJUK9df9V8sfq6cWtKiP0y3tAvs5G16+4buQhMmrzG0gtKJVCtwr
otrZSSNgnkNJXKjdNYNVeLqSRKToMM32RJ2c0hvwqTn5IF7Eg5DVXZqSYdg+FtHXKXAYzcbUFwyb
YWZR3lUXztlu/+bPFBOoGIjF5sVvvv7ywrHf5E9q1/+fzDvXgF2IZ8a6Z1K8k5pMeAxpgU8RO86w
9lOfzodpV4soV7Erx9kczVdwppWLvHgi0VkHU19G5E38G7oLRzw8BeYGJ++SsQFG3TLbyVN3zmpS
DmjgAJ35GAX/+M5uE8qd0aAoATylAL60ulPp0q1w1rSl6MdJ1/2uYbF8aacpOst90dVRzXoukATN
yJpR8a8jq7PGnBHF+VjIleHmBs5fvEfC7Xg9ncK+58iSR0M33ee+dvSO7NA3RLB2PrOTraXgmpm+
uvJoj3SEFubeIEfT4LsZLjcK/dKzrBLGoY5YeNDKPBZhy6HgY4ZfdZvyCzwr59yIpUlM5ksaffiy
ds41Zg0fnjqriObTtsK9h8tiIpbsfLiE8ojwIehEbnx6o+WChOJ6Lq3S5IoS+wcUfkpDJeh6oMg9
shNq+OQG4fPgow1J7jG/nE/G/fqqrM8qemeMlG2Ed2IlFqhK4Iu33PvZ5XQmnXaHat1bQiXdPbcF
Q09yIcR4jJNiokC2lo+pQ5+Lfj/Miz9/kk0KDYzBiWHopnaUuNxLANBO2szYh7IGUCuPkOXAZZg9
Tme0xTl5tHnLknTag0AT8eANhbmnXIE9cLl334CCf8Mh2ft2IEg+xta10MNXTVMHbCgrPFUKNmly
pFwClJtESH+zm8e7lvIadJYzlUqc6q7d/ZjuR9nqcurAKs9bCHNMneAH76qDY6f4wY7DuxnlATzt
BGzALfZKyN4aGhKTdSJ41+fYceGRW9wLwOKaLY7cMNcZWr1gsvtjXel5LLvmiXOyNKQoY6YHDfXj
SLsGmotALJwX+tBvRaK8mdxhIgIIAxKsqYspywFFjaR67KX1NUSRKkbODu/e38+w+H1Pca3oYz3t
51iIdilqxVtaAAInjIs9miAurmKokdIsrsMOsw0vUd2dZOcWT72NM9w5QA74dC5KysbZT+lH9P9h
9UwC8Y8iCkfAw3ezZLtqCcLT4Y24vPywh2vpBQ4BZkHmBAwFvtKiBGmiq0C5JIiPoNZKShJqZGjc
URxJa61pTby5tmmqYaiDAB9tWtFjr+0nC8T0Zj9DnijA+6O1l9/EE8ykPDuGXT9K+sL2HpwxlV4x
Al7vE+h+jz+9zPW5urD198RqBVvs4yxloTDb0gbxGnmmS2TNaC5EESUDe6ABfsnhwPCGBql5KkYH
mbvdKaf/GElUm0kJXmnaxT0LjFDCu1tRW1axNyQ0CP6sr8IZPlCf0KRjPzcRY2eYLOXo2ENNDgio
24kBWSKneqyTel+mTYQGAbwd3B/An8p1XqS3Vu7SP5fO5PFpFGRxSp6+SlLIEBjZZECbdQwBg15b
m2xttO8A9vt/Y9aDpS5Qhm/JydWX6+yPYjWtkGT/2o1L0Sc3XP36kVD+JsMvIW5oe4Kv3ieJDuPZ
haHXbjBaB6JgfobHZGMcWsLvsfQVW36VR0FunCuiHDzJDXRa+mHppv2JdlqlFM2cES+f9xAT/Pha
sazp9Ke5HrWa2bkyMbjKr9gGDJ6kZG/CavddXLWJinR2yWoY5vx5yFWb1cu+LRtNYtmPsFlJEeri
ab8jDN7Tw4A62lpfP0+9PtqE1a0lm2Q3D+cX0F4vfE7PBFuKWvLU1TlJj9OPqInoLsVdMDCe/d/C
FX4M9TbGOBdfXSz1Oov9aB2dU1sA5XbP4xIdbDnmowUlvRj+r9YE7xNGWEU1rR2uRlIsh33JYW6O
eex8ahamN9FXPngb17/sE7RKn4DBsXWIys3fYjmpNuCNx6iew6paJPgEpWoQNXk0iTU2qkYywN8s
qVH3ViDGc8ReERh9aOpftD1P5QLEVIZBaWzPlXb8Ex+Bsd2jx2/MLgI+89/SD08WQLJx33CqkqoU
43KA8yR3s4VJXGTZ46LFZATjdPeyCB4J8JrZtJL5bGqwYCl7ZHQdi5N74Wl6M4JHJt9amDtxpJW4
ziYm2kCJ/BRi7a/aBbXSjul9DZUFJTtNTrOBT28p9w3VoYo4bCnQlwdErvQvLrqAfpAIDVivYZwU
+ss1tDlEXQTWDoMr3OE23V0IawF2CaIeMlJmAYsYO/yFGjl4jV26zcFxsCk5Lu3TALHJ/0kgrs3K
Vt+9dqcrSkoF0iUfRZ+d3yyp8xdE6ZLFDjzu/1qgAD8ROQ0cniAaty1SQ2DV4DHU/7vXuOZOkY1M
l0u1rXEpKvpRZPQbV2NnrLV/9KHcFWAfQCMnBOP8dJhqz2SmwtlnCa/dx8jjRVK5yPjBy1GZFZ4d
vLHCKERWD4TMkWzFPB8EzCm1ldd8mZHJOvG6k3MO8PX54T6gWks+j47wljw/RzELCmGP+sPWIExP
o1P8YLSaInI5vJdbl/8cCJh4kEDEKTaJvP78c2hOgwETkVUmdWyxvia/yUHLbfHOra/nZv3R4kIs
YbNRQueALzBKodFw7kx78BdctP38Ac2OB/7eMLl8lznM6xgMN/FPMZRVZdWi5jIZk95KXOOnmjmf
rN6Aq+EljE3hMZQ3IKXgmXcogxM72NqsvzMpoV9hfIqMHnwoNvIxDvLhaHeBCQ3jiwCCk7I+rTTS
RdWplqggz9Wn6e0TwE7Xfx2UmSCG16KzlYvF5Y/ery378GyLS0PM8lmONFoAB2lBf+S7B5SMeQIa
Zm8PCmmjpFi+sLjN2N9NYdIroiA17idW/s8KWdQAHOmbDFZ8XP8msMqkJWnt6GtLNZLOy6gj04OG
FxNEGfMavCfkkxFpzCCO9QmnIWh6iYlCU0UOXaIT7GwIj3UkL9SGFeIS+3q8UlwnLtArxSwxzkdB
0SptEYOHoTUwjn3sWPmE27sjNvsxo7B/JLmTIK7uCr6ak+SN9TFApq4sty39zg8l7Q4/pgxUQmyl
gO7MiR5apCumxEXGlB8ivTLYnQkHYzPmDxbNc8qG5wZpL/UoAYJR3zWIpFKPvLNuXpV/JozkTlIo
bv2SWdUoWU9/WB7BlhYmJI050mzhYFCqVCzUPsJ1rZ9ufJ6yvxuNpNeHVXT8ItHP7j1cl6kIeU8e
Ktl7sE7Oi7I+uNGJiVDZ8PHchhs37O+ZjlAitajkNiBbxKGtl4YCajnt4pUG6ZH5s/XXvt4UokoP
/HWqBoOkn8Lktys5y+eDtQJdQPEb+C+KiW2r1S7nGcl4R8rzotadsCRyOvdXwQysnEqMFTAFPrgu
+8NzMqAbH4VAwL9cwHPicDKe2Gv6W/8No/oHbzHeUz0k6bBoNPbkbfSiJGt1FIRrUwKQWB+QyVJv
LO1cc84jy76rzaAbRaR1bClogAEy+sa4axF+Jea81nRL6q6fCcEftfJfbPothousfgrSMNgboiWp
C9KorSOOEhn9I0aaASmr1V3vmwJhV6YXLpjDOyN/yPaeD0MouPCB8m7uCtFtoSHy3dokSLjndAnN
sY37qeWVja7hRCHBhCxZWKrOHocIFFXwN5ZSz24POfvmju+Ure3aL4YW2b6Pu2aA+FxYFMDxgmmk
P1gVbprSKbkfFmOymEC/VSAb4ECJbg2CDiXSvk2VAVi17fVRvL4HBtWe+un4vFmy4YHI5VU1+agL
bQ5VnJGSD/3x57oey9wqu6EJhUe79ycKzl0yJdlmLxTAs6/jkrQLzmp6BHsqgesGdbU1nEVCyMoY
Cgf003Suq04uI2uLYUvzULaBI3+XX6eR/h/Mrp/U+TtExEnHJUqi4HP5RKfuK0FvkueDPMKSvpyw
S1AIawzzgYe1XSZEQpkl01hXVeHO2vqKwpvxe3g3wgqGuqlqzz3h638L8tlLnTpph2jdTmytQVzU
Pnk6p1QXMu/fZCRDzNgeygQIdMAl3+EDoEgm63dHttzSlt1ihVA2rAL833VB5PhWnNbnRzian5L5
JaXLMPQ/Gbd/BK7qzj9cD5OUQt15CSVQixyEmyt0r/at8LhJ23jHEvNUNH7li9p3tPJ2SzvggGNV
aq1+/t12Med9SgdxIS10ECFNUkJ0Q5/TG/fBe21JIvhQfqhsdyUIMadjN2G1AfXqs0Z0jfWmlM7y
devbU9WS7F8nleb4ZgMlcIFwacLgRvw70xJcu6YRc9THNMVdp3y8rKxl9ilPFWAHPlwZ1+KdWFvI
mIp7OJtFOsNNqCIbHNrV8a00rAWU7NolZ7v+vd44JgWfLv6+qLmCdHlgQ7kkwxEIHu7uYJOlPB1k
MoMotUvSDNy8GImZJOhcy4lc+EiBQChScBppRnwW/OaYtUdABaWb0XnvEL+LlxzmlNphQgDtJ4HS
UBfa10s+gHAYgSV3h8vX9+rnKAWAIzjLezCkJVDLQC9a67u0gTyLonIN7DqLQAd+i76Cti3xbq7P
y41Ez0QGwsCNASvzh8oDmc11e/6TL3+qXKmzUyIF5hQId1ZDtQlO+LhmQeKIu/ySakNm8VEjoP9x
Wvu7JmXi3ebvxm8ngzsQk+gv9iPmuiMJNwIADbudww9P2BbjEVH0a1PwpCL4ZZIUvOWkxjDyxDCn
7/RXqm/BxmCFtJCibXGDc7Rp21KiV+nKKbNFYFqXaethyuRiud4lNNRlCsxscLa/dK1RzkVCiL4L
DtW8JJCMibaNFrxC92E6xQ+fligeZHXk2V/I+yD61z9810dguzH1OjEOLbfmpaldXlLGZ6nsBAqq
/OD7Ai+sqpWTeFkqO4/Cktjx9O9ArAv1HyJLFNBXXK++oHYU4Oxzw60NQFPnHS1x9eplVbUispWg
FA+bqesh5dByxQKmOcYRPpmPistD1GY5bcSBSep5mbkE9Cp0N4jUkq8YbE0H2hFdcNJtmC4u5xzV
AGWc3eEd0BbQrFq01yHbwMYcTaZAK5AWWT4+jHh+vd+FiGe32PERpWod32L1e6ZWwYS4SqAHz3OB
7QkCWCdWcDUjk0ECBaa3b5gmVnf3/lXtUbNigO0ki/ZHeXX3g6AMWB/QC+hfeGGBBKcVJkARCu/U
ZBRrVLK8A960z3kohlvjlCoxUX5GoTDhXQ/sF7gsFD88sStX1Q0IcezPiRESmoMhbtAVG14pgdnX
v39WqRRSPmDzPaq+alYcC9AolP2ezmbxfv+8vgi4O7dmLgfZGeNnvNM/XbZC6OsqJ2zCVIhohEON
ygPKT2XOysujxKlY6IqmNNJpu5OHYCL95PktienJeNVnCx9LmJJPZpQw2ycaCSg4yDYeLZ+1IyYc
48EHaKx9m+cyFXtU8gvKn8HTzR/ylgqxuXqEjvICLjTvChcrNosuhzUXj4fpxNwkQFe7TqVA4ElN
QIMc1bhzE2JkLfqBt0BXZSL63IWDjamWapj5Zjh75BU1gsozbFAeNcC5/aIFf1nuiqQ/z7VO9pYz
BZ4gU+RFkb1GMfUkToRrGF2bCcuMXYKHNynQRazGKpJ+f4OL5WFz78wYFjidxmfv6BIPylQJARVF
MzUKTVHGSXmJx9GdrRsHuO5PNFWDYyS5+3e/NJnRQN0M/QxQJeEXV3EcuuDt0i1EeJR0scl1mdLj
t+QgbPzKisoeRz7aKe3DD8V2Bwi9uldzF9A+iMKx5kevtp0n+YpH/Ao0eDQNu/l1HQBeGirPSWsM
FDIizxgCDzmRPRZyxI0+nfTohxA22BftXvid1WoCTjPAJhKwEiKBeU69HqdzEKjF6J8JtWI44y0m
gcZ8kpng4auHRpCcdyo/din2dWSKTj5bYrKaqOWTut0hHF1CQ7p+03TXsHTvrY/y34fh/MOmPTzj
uUXrRLb0dwcXK4cf+81V+i71php8370o/0booz5kc41NCb192AD42i7UcX5d8aoNgIhUg2zoFO6B
/639GG6n3L6ilf6HGp0Hfc+a4H3/vXhp4oBgxsxsijynBtC8IbdE2nP7cA3tqBRdZyWDQdmHbNsx
Dl+r1ERLvcyBj5Ouq3dxUUrboRMVWnrM00j1HW9L7LOz+le5jr0vmV0fQTEq4E0iDpzaAcvV32rX
2FvRdmge4lzXFSTGbM2wXuoj0y6QNkKuUx2jjv+2gNr2ywcGPJNNWz7Q00Z6AwHNi5hDAii7agff
L8vqSqcPD5w9H5ejTtOxlPUA9OO8hwoAWs8BoGZVLMbn37SatIS1NGP1/W15ZXtr36wDfPk+DUTO
SZdob5nzd20PWeU+mfUOrmrVrWRF+XG9nS16nbmU5+lFtGhVrXVbrDIle1P7GFf5s/jZB5cD2413
s69aGmMtFzqlzcsJJc2JC2LgX29S1mF3jgxYfB35PwiUuxLW8bgjXB42ufnS0NA8VLh3iGLhEvqz
r2aQZ2cxqgiwRKUTovI1o+VUfrp/P1qSbFkuTdCn9Sn4ZYChxdNxV5p/feqfQJMjF0gtMue/v1lQ
A03C30FNg1GNLIviup/ZQ09jPqRg2q85LjCE/ork6Er4sXPlE407rVR1x+M5iHL7Hdd2wvMANpbN
rm3AWT2MQ6Fu3FQ5nTpXJs1jdlAddo5U1Ebgoo8G9sRufM9qQekS5a4+H+lYH0OGujsMG0nsNODK
gUXTP5F+FkCW0b9pa48OpocCU6iruHgsGyCz+xY8kiAEXJXd4doa5Rbx0sbDhmnYxgeXQekpBLV9
WMsSBhbZGmwgmSE8LLiXlcvc+8ZS256Of7nZbylJT2f/Z+10H8gxDmE8kD2SBjVWMZm2BZEN4iH9
JDl8j94pfoqgKXnFc0JQtGOg6w9pw7syiN8h8YCbj7Fj8m2bYpjQmpvKc2YGQQPijcQ9dZKYxZsE
Q/yzXylgSoO2bSn4r0SfYFx2iM4HiiajUjO0Kd/Z1yo0Rwh+JPv/7cbCpTGUi43We6F+9wVVizhB
+4ZMdtcg5a6NEFBMCq+e6RUEe18mNsTaxdV/15w9RkDhv+GtsaAfRFUxNt8YZ/rtdGLwdStasovr
vZjCKC/BPWln3Fey9qeQryIxTyZ1zgSRNd9Fcf7KpG/vdIq9W00N7jODnSsvmWgK85F0B2eLt5Zd
ea2zbYZelM0f29eZQhMndE1JYYqDaoXY2QqYGElqkUnBhcijo2+2Xgw0hnl/cu1pyq2/ErIn2MQV
Ss0POiMWUgrYedkbODk8U8GiAZCoQ+3VGrgDwzYKHF72Jc7FmiwpeEViXjbIAK5aOFe6zMYpcarF
9gCRnFL+ViMMOaW3T5chDlWgi5qbXrxs424dA7YDlrrDInsYd9Y+g3eM4BYTVxWx4jCplNyKZ8bq
AckeGbFRj8EhWdsaDe+KC8wc8SPSIIy6Y5oj5Uh3Bz9sEiXYfS59HrnTLlicQ5U+O8WIjFFjYnWu
WUDKw1QxfkzBRmIQm4UGEzbEp31zkMnouNyIG4JtkkUWTim8Dw5iRiUk19uLJuw3agdIyZJdvoKB
vU21/Q152j5cWymsOvGmbQ4S4oyMQJsdG5m8Ev+iy9ZDTRb65X3fBjORpN0eg1qOo8KE6hOvJ18s
joQu52NVe3w2FT+CIHEoRDMPvlSgVTqkxfK5M2M1kEwAQ+X/kgNXs2rdbeGGTl1FkJoF2H+JsDbI
6UltEPKSFOLDhk3goHCypM2hxr9ex4/83andIDrlmnIz8PndgEwdktASmGw8FOHUv0EbhfPbqJ3s
C3xiiDIieurmUX/NhCVxCWA+WAnA4h2+WlbNvOPJtgmFQ5iBDakvMm5qV+wNpN3gMao8ibvxNsjD
9YYaJpjz8UEWzw1Qwc3HbghEf2pooEqY+00MlOUPaoszZoOGj2hn731cou1APDWhMKROqmt/Doi5
UndYJKi4afw67VzmhBX+N0LOSOwZR26yK6OZsAeR5Z3dRw1Knria8M9LUsKofxYFqgKR6eFVfdq1
XMNWOjdOmGSe4Dp4zvgwRBBa+oAW3VABRd3mSWl4CjgXg8ubF0iO0b3cqXEXcM0ExvvgUhZUl2SM
OjKBs5azZRMmg/xCRhqWWeg99IM6sy7vLQsGhbNQ8h3alhwcmYVcDfFNevek3+ArSvtQhOBIewvD
j5aFPIScEmFcRhyxK6qphzYbHmsbcMUUk38OA9oizWUrCbgaCAPjiJYcErr/1ohubudC1RQxRiV8
LchNLU4a0kFPTYosoVe6ais3mW/lbGlgrB9zstyEiojit3SlH8aVj3IRYaz1EcF+AbMYyCiySMrg
ITmxsuEdn3IjqPXdKWjA0T9XGfzU21C+MU98224pF2Xfejd7omXRt2CHKVTxLDie4vx8fqKdgP1F
6jDn+oXYP3FoSXtU0sLtJeNrlsAtWQPiEZ3o5vD3TAmY/lGvfTpBWWidQ/IlFOuAgDCqJLJi5gRv
qHbCQfnspPg8gWNSvGGsFTbXlP4Jy5o0LUfKQmWvPfqYEw7O9Pr5BmfS14kQaR+QOMUFw5wrB7Qr
ySdvSixljwuDKZkgLBkDpItyInc3/JJJExfmRV5ZZYj9MD8cXUUlZOHQ7Gu9jBDhhhfPbjk1Uc88
p23p4o4FbuSn2gFZ6rrVRZs8MN32lOpzC24kx+cMTo0rYSnqpzq7wBdOpa2n8xhqE18pcONCCdsV
GfuJN1GblK5YYGbtYUtDFqXhbyOqINmAiKp4LtMeuQETwfOWY+latmEotSPHf4xYbBQLFoYGBSv1
PmukYVHPH1AYI1uXCwDfFhW37K74kmigleCW40h4gh+Kb+LCpr+zWxXkNhQ85iSsKn0xye3MiSAG
lTiH/UOySuF1uvBFofOzi4aIHM1B5sK8SLTD4fWs0yC2PQ2pkqk8eWjoVCwB0x/BHZyKlcxKHKWM
vQ7RihKKbCbExS87JM3Lda/drxBGIMoHz3Q8e+1J2o7+mAH6Kr1GD30JusnwXvz+klZab4YeTjmL
5+Dhuimlkpnns5cxHyx4doIzTT0kQUmfqpG0JA4ok+XOmjLOjpWaftjVuO6kagO7sHQHZGzsTI7H
UTdruxSgz03MTxTqjHrXdCooqLGdcnQ4irK8XsTO2AS0o+eA126GXrNHUz1n7OtZApfb+aSFyx8c
xaUnfDoc5FvOgAG8yvksgd7W8y7VYd52KjDzSaAood7q96EtxGpv0gzlB2WDYYMYRe0ETa6AUAPm
WPpC8DOM6xwOtA4EWO9JZaJ59urTUKfolQN9coTsKQtFtmLV5Yq1F9VJTLBgCtnzG7YW5c22zV9U
eB56hW8TZQ/AVXppxUBmMoTLNTgEnBucwaDJ9RGbMnZrQNwL4oKElGkhscC2VLgPUlyekQlkD5iv
/hYlHtwTo6u8dARMgh42cjBst1iuX85ZRwe2a8QVqyKidkkbMlrrkUVUr+Rnscq+tD0YT8GgXbXA
tTr1KrLV44hH31k0kTmf43i5pNpTVO6OnNsH6jRYIgDrA2hlnbkCYF/ma60V6XF88o6tX9ENz4Yp
/XfWosqNIwMl6Vtl6Mfpu+l672LOvJgIpH9YhhFy6aBHKLIfI6eTKjjqXmme9oDNUXZ23oNNbBli
1DMKXRjEsGwT/FiI9gssWb06dJ6lrAktuVgLqmWw2nqVFXMbqOn+0XGw5FhdkiKht7l4bHOHX85g
w18CNJ/l76ks9s5XAs/vYHQ5VFAe9+Sm4NDm2hGzBY0yuscXBG1GVt+NmMXaTHRJ6il/OO2XxrxX
brpUMcH/+fgDy3XztCvHK/EKPVGH7aGNHGjdYEr7aVWznviVP0SiT8MvEIYYq/m+vwfl3XvRfSZV
0ddb+lDRO40qM7XGR92kDk+XqbKrf1KvkcijcFvpgnZnK68owJZ03Lae6L9Ey/kK5kynhh7EtgiU
GDSWRE1DAvO+PR5PzP7UZcqDw0o8aJuFp6aAd64i5coqgzpbxdVxVazO3PwLKK1T0rzFyKOmEt/a
taKz+WDxzWaz7AQMWAluvCTLeezL0mBYmu3W4vgogb3QWiWzBmopR4NZb5EwhV1I2QHCYsOPqmxC
qeowZ4I8MYG+EVCEphCyvDIN+LarrwVsDyuOyfxDCFbvUnXPKMxRYq9hEaXntBA2SVTxYDwkMN+7
bEsluGsiL2ihZCq6Nx+45VoiAkeF1n1nhfj6gkm8fz851lVMP+1sIi7RvOoukyjHTf0KqNTczIb/
bZ6N1xoOEFRAVH/UmxwLDTlxtqKXkxQp8+qdV1cQwPMEhTaNhCkuLdYGDoLndOVCj7Qe04p9CRB+
6LaEowXRcN7NXCwhDdxtQEmOkaZZ/oniNh1oW6UuhmFAUnXCuOZyPjF7a7ab4DLkmZzry5P+N6gA
I6BTyxjJl+M8hv0bGodyOe65leMXZV3ytQM0L648c1sWYOL3quaW08/KaB28sUKSJdWy/8eYa6TN
yHa6CFIn+VNNjndw2PQMpi5EWy7/0rt2+eFWDaZQ9U24GwyHUMGT2g1VECtutFfQ0w1dXdRGckGv
7E2zKaGsOuyALuNGlRWTe3fkiH7nxJRaLQv779ctT+1PZYM6hkNHMOxNhEmCV79VVhqJiY7BVZ+P
lnKL23qeEXwxK15y8+Ur4jcVn8FuE7R70KwRbq3fcOKnhFQsItBJXHbBRJ+i336Dfc5PE5lipoBo
DY5BUC7WYPSgJcE/Dn6s6DG/qoNYNmKw1sY468vnJFblltJSQLH7ruAFeJKtV9ok4P0aZLFY6E/S
qnyoajLLtUMgCqV/yLMDwOXy5mMxR63Ac0JuDaEwX11vJE9dd6lwBlTd3lFG5Ipg/tr96nO/BAKr
nL7dSUrRQw2/A6YUmUgFP6X4V4N1+8aKiU0pmYRI2A58Pns/uPdv2/2WNDEWj4nRfM1CDuB5HFbz
Z5a/88jkTSbyfQoxWOxF2nuiq6cBvIyBO+4ufNH5nEIZSYyk0zwq8FOo5DiUL4334MebjjIb0pf3
++X8Ixf1ZTrLtynTTHk5ds+wAWvTubuQOF0c3wy0Jo3LgZJmXJ/kgD437CXZtw1dczGLebkF1FJC
l2GejBcRN0dGygX9vWjwkZQ5//PjJOoFWb7Qn35yWtVFE+6bmNMD0p6++SOYyZuT5gQIcWG9weqI
SiKZtnHlBF9V0xuv8/oUJUrkQU07zRe4xFMxtFpxVOnkWJFvEkwRghLmBuyZSZqJKcyqND9b2hcJ
I43oQVihmlOZYFQsWQ51vm2VcaCvRFjOT4hwrkP/MKxCwV6IqCGe+OlcJpIM17hcpHKmW44saQAd
tYwa5iLUtsDQuRYpZ5+rj1xcJOOqnMWcNsnvznlzGLLlmQUzbZwSA458Yil6BP+yUvncqXW6z7FZ
OQQQn+zq4tNo+JsXwfJpFKeCJBNCLhwps3FPZ3D7N5Q6eynJufWRZZXeDEcNW/sYcshKGdAhQVuN
hvaHiemOxE50Iue6sBUMrZokD/Ae8ZNTbvZCXYGC5ai98KUDkhIk44ZKWKONlRaMvf+YyEnsnrZY
7msZq+ApG7yhjHdUy5TCqv4+tcplZcEFKZSgWtwPXsa6rwyLxEpg5XCLgxaB+Sm/yxt/Qv3BTaam
WSm5jvMVLNhaDC1sAfKfjnyStr7HnNldBf0PqWghJjbcKTik6jtqOPOEnQZFHinDxyzd0v1hI7RR
COV2lCmFbfqwBhXW3V53Vccx5pvldxwpUMkyAvrSHrj4+5SaSZLxXH+QB1RtECSvWwvfKapaz+ff
lf49PGvDo+Huu2XNgkiKG0JaHB5KR7VgEjI7uP50mUkHNqOSGqFjLkBYqvdN4AWN8lVWYeA0jW5I
OgajFd1VCPYrHyrxlsjrFvK/8Gk4t1bZBB41hUahswAaDXWW6o2+hLoJ4VjldJ6sUzyJFz3BS97u
eiUWzRFRvICe9eODRH1ULVeGEtDpk8DLKb4MCVhS9RReVfPSRJh1Ok4DMqKXuWSB0w+COJuceMk+
K3yv/sXCxxF62xZD6e79lBBypdphjcFbJ4SA5zi7wnZCcRaLmIxOyiijgs+BLQUbgSFwRbO6mYeM
0Oe/jx21+3YaIUTBT/b3Kw1PVnUVjl55xZzi/sk3S1FZ5Kiib+9jQvz9krOE3isxP7xhfEkseVVT
0RupcOS9sUm/pkFCsQAM2970rxsi2g4++y6spHvgWhUamXHtiQT91z+kMZJ3SyVXWgYimqeL5jQS
bVYs2UURSOZE9M188vdoizvviOYfvDDRbXpgiuxrJN5z6kBetyWOgs6yJBRAHZMc9SRkQZSMGa6x
WAB+Ohy/fB1aCYQBmKcVYr86BQx1AvYG5fjlEcWt0gkkpchGg2uoiXgFF+e0dgh+3ZsGyRIpYIdk
15IjDGp43ca+U53FHUflvK1J3JIeg0YD2Fgs/U1yo++EPXMUIwGAs0HOyAuV1jUEADjpGykIuT+8
7PlpN5/JNQEnB1ylaQ8dGjXvXpm6dSkGEDuQC9CZXPRsWqp1W/yL/H4V5193kqrxf6wEKjjfEs7R
32BiA4t4F+maK3spANU29iJqRpVH4XB2aPqXb28XzQoezHhxvVs/q/vuo3HudQw7pQJBB5axqimv
zu97B6ilzbQ0yiGQX6aoG227hJ1/xQc8w1nFz7/eRWbbNzyETSgoLvxHQ6IuqqdeMq4G713qn5sY
w9h8jY4u7lnEMYwNUdG7acXgFN7+e7pQh6mKYsukUtwxVEsL3aFIU2vAH/NF5CtK9uOW1l0TseWa
oL7wJv2b/ZLyNixdXBTBmxHsT6vbpa/zR9WAmomGeXu2CbUzImoGT8u5XFyK9tRaDhZBlqob7d/V
fWkJ9bHqxAJbpxNAlTag4BH+PhGLerlxKECu/o8YfikInqiAnM+9UGX+Nk5Xu/yMrMvwd+kfmpq/
B+zPUIFJNcswcd/5fBsd/TL/nOxIyTGEDsPqvaFz3iWxA4SsvI7/I+aNlZL98MGIkDuF6dFgazIh
j5Y7xnhzPRoeti/svDCwSTYQtWE3sk7YbjE0n8juTeqR+fhM1lgetRbwaAHnXQIAosORMhwgZfgv
xQswracg+Tnjw1WksZVqPKPKTaTO2CqWZ6NR4ttRbx70Rob2Yr8NoeNS/GB4Rymi1CoByfEbFYtS
7Ginj4e6I/h80R8h+yPBwCvGkEddsutWIISITMCtStmQLy+TgZU8nCwvMVxh9OMFo5bQSItDAYB3
8vVNIQMpMFGNzN29KOPQ95dpeMBhrDHe6zsPoXIz909jwWtlqW2vnw9u4PFZ4zyXcT7RoWq8BmE9
21U2M077eEe8hLlaAC+iZoyODEOnWy4KMr0zYIcTwqXldfDIQlEqhPlwTXkpt1tdj7mEVb6VYp4o
xcSacBq+N74GIPyMviBYpcW9jE4eWafWslNa2iMon3YwJ2QRmvzfgQCsI1bwN/raKChSLCY8aKi7
TUVp0oFgBh2UikuK6v0BeuCCWNSJunKj3EKz+RIGZNnZX6kD4o/UGq5DVBCxKQ/1F+XleOePzKKb
FC20NCoK7hMW5sF8GWGomkU6GstS6DykFiLW8/H19t3tHeXSMJ6TlsCkpSP6DkkptPjm2bve+KjT
stQEi0ikNUFpz+8kolGf8lHO2MdfgiovISXwsSNuQr77OY/CcUgMsDdE/zHXap51CSGKqyJvUtMl
GC4k/zbxNUSASiFKELp2MVVR2z2lONPx2Gz4NUbG4+Y9Ai34AHfxonQ7Qm9cI6Oj7hlhcNRx7soq
AJh1xPeGaIF0q06WZt2JooKywibTtYE4u4Dd96lVTRpKtoWdU/myv89TJWuEKrTxA1Cg4stnbRpX
IgyyTcPNuqmHTWFAjkY50RmLUt93SrZHCS7iD9FUQRr8ErBgK6nk79B8XeYSiqr8kj4wdWFmAA06
0GlD3oEswlHXA4flExbS4Q+T61mB7ZMD4Nqaii+CM48VLuAD1btQCHKAsLYieIIaZ6uVp2pLOAak
X11DMVgrkT7BWA88nH4gq8kg7UNxk3QEEiDTksPR0nuNxhOGxmnI3ipEhQcsEoGUQN7O++fkTcve
yEyMRRo+MGjfynUTEGieg3kzcsdXS5J/M2FMmutQ1+QgcEqLAF2TuKO8xg62YxW4lxb3S6ZGSO9O
T5v2+JK3BZHF+auebACA7HmhF9CtgsB9B1I+S38+Ua2EsiYcXlaSC5d0bWpHMypvJiQiAkBROXMX
4v2OMxnTnAPyamMkx++m1+q9dpQBA0+sLlWRt8C9OpvSdvx3HWQGKrLxswwvJk120GMb2nsPlYsT
FwZU/K10bXAPY/t9pFbgW5smooieMN9eF0r4Fsm2kcy/HffkFkq2GUKWlUkWTKkKcIkOykwSHZFY
8XpCpMs3Onqdjpgd7Slhsr8jsz+G75aBx4zZ33qf43TRyigVKGSUnOv90g7d58ye3FqZFNfn9vaw
EhXqqCg041vScxoAfxmCqdzIZ1euMFBbDq2YzYmUuy4hiDn/rXTTGm5mMTIyMjgJcdWDs9TXLRUE
rHeOhPbuQuGoXoWQs+DYHyj5Y4DxJtBV3+0m/TDKveA2lesdp0ucpLLEhHFdkce6ZC/Pl1Wd3D4F
OwZ9FYM7/085+IhUp7SeToEQKstvPJH5DeU/YgE2skooYY0PhFBG7Xva9VWwTzTVVb6xqfyuZZJT
CQ6GG1O0KjNytY6Zcn/gURg5TzpM3NzwQtArjgl4UXGD7uwZMKE066IIJuKBQWUQePfjQsAmlBMq
xvpnb18aD6Zd5sewGeVynAZ7SyDh2RJmtSVLJx8RXeDLkX9WVFT8/z/7dAQ9cRwCqMZKTcH8YuA+
fYkJHFNUVCoapB/2G1NBO0dF90mHmz1V2xz4o42KRs3OmsuLiPt9pIiVDjSZ/u0ZZ07x/9wdxY17
R0LTBGlGkfbZA4C63QlnS/yp9ksMCe1PC2XV24hmzMRUqU17JIqE7M1pxPm8Ae6OKT4QncRH5xbu
LhtjGXzLfcae4wUmfPzMLGZblZtq2Zwe1a31iusmo+kuli0SlN6C4zVT9aJYZZRQqETehC8GI7gf
xqdVLQWg5+VdSKQrtIrxQKcsWy+Xi/J63YIgtTwUZPOZBpyJfU+WqHbT8UkYRAAUsqmQ05YRLMfK
/fvTBDbXYHFxCIWqnvRhJJZmzsB0NyPT8gNhQIV7Ay+xatw3aEKoFr675V4/jBV/f4e0BQiTd1uu
ZBcp8I/R0AzVuOwNv4G5/btZ6YBjfM8GoI6hY6/7uAbA0xp4XYtnu5Nb0xy/T8Hk+8/+EQJ2wMrS
aWTz4qSr+jlzBcrvxTUON0vgt8Bm+Z3/w3nHxvrLyYcqmEY3q4sUtPhmVXKgS2AdLBThB8W7FlDN
0x6q06wBWjXapIoJsBXje9rLdyRXcG3B8G+OuyjSCJceJEByMJMadxpbE6m6THfl21YO71CUdRU0
ZlRLbzx2xKcIs85ok22nfWEr2ZVhWAts4OfiYboP1mUq1ixxn39Z9feYpzbzO0RxFP6Fow74MPnh
kZis5KEWcLlOHyZgCK9+twXXEaTy2LEArRiFom+V4xUOfjvlfrYfrD6uF2fgR7aO+qQfkfvBsCbF
h0m1wC8mtcTryNXqtm2MTB6OVmRqChH7c1X7tQTHznOO723cgvkoKuQvufne5vxTFDCHwwdOFFRQ
FZYmpGPan6GYn0IqAZkx8q5BbGB09BjUaB0293LS1eoWQ4OoPk+JzU1Fj1Rtb/SwK84EVfdvxDda
swWIZzfVPCb32WwWOxwD4Z0l0Qph6vo8l9KqyCuDqr9YhF9GMBFB9jDGP/bqJbySrvb6D0lW4MIE
6TUHaBUpiJ3WGyqV1dZj80ibSpngjC46tT1c+HOkuFohMdBPEjJuU6sVxeR7rD/QDJcL+FvRDmtk
LlvDH8ydWPSGYlI8WI64noLlDnBCKvxUh6wG55cOHlPH8pwbYo1xjDmyzwPIgMG4fHlBEl+F3V8g
mHTqL96OOB+SONurJZOU3I5C/GBmh1Ark1AMjqrnj/D5hq2ms+YMlY0KKhoXy+MnZvmb9A3Uk6hf
Gqf7r21QAxt5JSFLoDcgrDec58rFSA9dGzugpYpjpIKaF3uy7V3MVrb5JUiZgxhlfqMzeRGxrvP5
Ao5bUruhtkyvkt/IwDLjDwEBIE1bZdHynpKFcsXytHDwblGDuIttqVBwJxpxkkZZP47NjuL4BRmp
CK9UYgujrbFtIFT1uTtjip2MbtvDNyL5KeYu6iR5j+2lCoGe4c3qIENd7GYt0o3cc8M0pQu2alTf
BQXgGf6nxomqCwGAUoxTqeDI5ARbIA6DEYmPIF+caT4P8qUmDXBs+UBsxW4S6/OhnDKuX9Sj2jUi
ZEs6IHSzo1/7ATLjWAHerQnaf0cKzqpCvdnmJ2Ti+d+yTClEs8aSTpXpRZLffS7DIMlXb1erihvY
GUksKSJVnscKg1Yy74lWMGcez0xshxpxM1dtErzweGMv8YxEfpHsJ+ipxIy7kGOiuJk6Wi9D3AUM
L/0suQ5i3gbpe8XM9pM6l22OBEcbaYH87eHHz2t5lUPYeUa6lSovvRa3ol7m0Fe+5k9oPWoo+ggm
mWlqnXuDfT8LiNSTtsZFFVPdXbhAzdTzU22CimFuDZQDetnrzHZcGo3tSGhHAGlyDrpteGURGx3U
D59u4+FuQUOKucpZh8hzojb/uxf/9EgcNGGr615lIY5joeZANsInN3iub7Kav68ojYs0wfco7feS
69D4xmNjk3Dk6RFk+H99N9atXZzCJuXrPcFi2bOLSKJlJDTt5OEN49o0rB6cHMiUaCiFFgXRu0cc
7o/mUoO4guYq/lO2LqylYH3P/CpJfRqx1/C49GM0t5aHXGq2m82OqrYNADJM/8BifVkrFZ+TPCzk
yOWYC0RPqheIn2CdR6unrxxTbx2Hs8ycjZR27GnSmBGG8FHq8+NR6uTVCKsZFVdOotO/ZybdItiO
uBKWnEWXWvVxy/hYjOsd3R5tVyaK10uzcl2dMrJfuVB6mVD2PqwoNcqD7vf4yAod9GYD6g31DHxw
u1WF/NuVQb1wTlx384eoyybUdGtyxISEAGff+jsvUnZblF5cmz8nBgfsX+jh8wwS0aINwMaSvk/Y
Src3ODRJ6ZBYb4adQ5KADHH0FzmkHu7sfpeZYEtuktC5LS896zl2Y0fErBybMkg5qxM0JcVI6miR
YTLiOq0SQ+fxRNk+NzhAOwXd0ZjZ9PtUTmQGldrjN13RzuHnPz3b3lTn4QJXmYIyR7cNYAda6HrX
jZrKCj9nTj/iprw9Q74USgtmYBtXKjWooG0Z96JiYTHblKRAw1UQqfI2tiXV4fzP4ZPOqjL/F0f1
ryfZyatzQCopv8XXlpUv8Ax+uuTtJJP5WPJpCJ1LkGVrNFdo0BIO0w+eHY0VG3uLLDQvzlf+PW9q
zTcO0BRR0MzuT7xqKZdqfe4sRKxmf534nmd743bh92HIyDscOCccvhvy6s/22NUmpA9Oi+frcEZf
RXKKGC7JHAzfHTF0xrP/S78LwUIOWJcqrwtNi58auI2Dw8Rx0qH8gKp+KVuNqNmuGCZAKJvxX0JY
0f9OfIRNsepm+w5z7P72iIaEiOL1lMrUONpWSpW2im87AcI/nKlbbY1cZooVsqTCXAbF0K4ZlCgZ
5p6fo2Q7cckDGPYwQIe7xYvRDT3qx/9ptRUt2/MxgYJzKX9vWXw0/gAsVMDUVLQbzK/RfhgDrGgC
8Ly0lB+epILhYdlv+K42XZY1lsOrnWfl/yHSh/eCDL/9igkNjI2MI7EYnWUx1FJ3TAV5g9jC7Lfz
2IMZ4YTcnlwMFaHs3nZq7twX8KnkQBCdR1lfZmuTvS0beVCZjLrfeweacEusAy7ubuBO+w4L0YIB
drfxVwvvBd6//LdIvpBEDUeDJAC7HUi6A4vK0Sc+2KLH1fFH0ogf/slzhyeyvyRSTaXVkfxQpBHJ
bgoGFyO6ifj1zA7gmS7K4n+PN584SA4M14FpP+n7V/8XhPbYHz+LeNjYwSyxTZkNdtfwwRpprcpO
Ynhg1Lsh9DxXRI4B5W+4NtFlXgcXQw2tU6+BVuEMUBkXqLrZr1UHmPa24Ksl8hVRcwXj2bIUPQQM
i8eiWuTSO5kv+rVqgomHohoh69vRBU63gZZzEkzECHWlICV3tBKTsg7x+56dB1XookDyt/xYxZuK
il5V69XUOiasHEteVOQ9GO/PLP7PoH4I/VJ0PsWb1OmyeGiYgaSKK8us8/98UVHRbKGlJDSK9rqS
YvMNlwVAzcJnFDksr4/c/dYpCcBtqXnWq34+CXmv4SQ8LlP8+J3RtRXM6AFl1i0GjE4vg/2sMvL6
/YiwslDTMc4sPf3yOHzKeNtesNIfAntDbLQQ3zWbY9/Ahi1KnavSeFWYhJtCcyVlQRL+7+Sz/lNS
jREwLQ28J0myeqj/ePNnalPgQI21gzOasZSB3Qo3AcFn3nDLGeMf7+YGPyVCBOu8p6t/OMTAWByu
3M10a8WvoKEVdWohuKEWaoKUActpfbLPt4Bzy4JMetlJTdg9iP9MHwcx1uF1kvCo59/oetXKsBrC
SEp28e79fAV9wy70rflM3/mGOofn8RxPbBV2DmGUrH9acmaxAMnUs4a/69Op3TxwQ8RCNzgHl2Oc
7OdUsfmjOcj2OrttbTDMRGzQtaNm16SF8Tx++ZR0SzvLEy9pQLl2V1b71vNJy1AHRo9R/+sWsQJe
UD8oImJ907V7WjoiCDOFxpi1qPlCv1x074GyXB3jliv/7Z/Qs3MMrPWjxO8xKKBssN6eW4zIrPrN
DCIDvp7bpgeeQnl085poVsI2v3YPxh+YXD3DiplninU1wGDMSKxYVrglPOuZaBdcPyRDZ3NE9AhJ
EOPu0F7aXyUQRPjptHEkmOS0gMyjY/cNSK8+juSnOs8F06JjO7SXqHawMMCzgVj6xYfqjW+S+TvY
Li+AVKe6+emYNR5OKhFo9uFPT9l0pA5WO9gUUlH62MRlpOPzSKRtMXtArI/vnGKZLp1v6U9pvBnJ
i+6D2Wk+rinZrvBlVrTsrHjsiroxdEgKRdHSHZUuCjJc4dYeUhncZdu10Opoo7eUeeAirklc3DZp
7ZGT1jD1LPhabsYc+OY7IP6USSSiiuccLFGe/PmaD4Laz+9Zo5zm1uMUVkQWI543WYoTOuGYSMYc
GPv9r5WqoWZvB8YbKpXLv1h/NmvT8k2j/Wn5AakuSC6gmwBD48QVyjlSjYs2XaUU84uGrnCxWv5N
9TduIsNAuMFttSy/gIg/A3iaTcU9USzF7UJuTiQaKnEE+btmXc+hcyHSoOl98UFUGb94kiLtZ0Kj
bg7EEvbykt5yl+YPeQ/kp1KxLiSnZy4zEBU93Ns7AkifmTSxZFSMrkIJBftGkFl9bHRNpb1GcphC
7xP7HIj9GDBzgSC+pliNdLdZF9taj/pcrQ1e/6eDIIaTJYKfLEdX1cJtGNr6QiHPL64zj6hJvSCs
f/ojVm0OeXcHCFOfqoot58+zoLYCJjAzfpL4p7pvIYA/OvASzg+lJp0Ju/BDFuoCCVv8ac/R8ibL
Nh2Guqzx6reSZAJ8iAv0e9k83BI8zRN/2JDhf9mTgWNMyZAEC87Qk1zzacbRvoClhPAVpfv9f9Yo
SJtqsyLeLVoPYndohqRyCWfNCwgO38per3kujpEXsiLxQs96KscRuxO3J+7780uWKCxtxqnqSncf
YsK2yTWslqJ3XMYcGD0/M8vDSDsmHictMuP+JeqvMuTbMWRfIiomY3a4e4qlC4EI3lHN1AEq4aqI
78vPkRuW02GJZYRmbFj1CUDGg9UiTQS5do70Iyns9vzYBLf7F/VuWInu46KW0sZVX1cJbPdV68Ug
w0MlEdyqOA0eHPaKGYDuPRhsCM0FjeE4AUCEiP1UQaTxKcsTwyIRtBGfSGWs0pZ5naM8sakHKmjJ
ChlB9BKtmBRbqBil0neI0b3vBzipkL2WpE6E4ByOjPpOH9qtfTytA4ogjiCzMAc2xW65zcGvc16N
PDt3CLrruZDNb2Hs7H5SJqNGrCjJzh+hn4P2pX80QvBd7HfI+ti6Q0Q+7Dhb8NOVWImOa5prjzHz
nSn76pvxW87/VAlQ44c6rLorNqFI7b5TAWLFdZb4XtX9v7ffY/3oSUoCkEkZXCc/ER2C50dvmDNM
yzNh4YGgq6Pqqg+LuB7VsyvX6hvziZhBt8OQRk5K2TE5u3cRZc31/PnUE42UV4WYFB/QS7RoJnXS
S3n6rASXWzf+n+1mZhqsLiLDgsTJPO06T1sTovpUatJNdv1BpoD2ukRyI6o6mzgqo9+q8pvbyTlg
s7ngX65uxWNPiva+DzYr/Aboc6Y6jCdCZt2a/HDjuZ0UO9FWk14POFe8J917EtQXlTl2+w7IoIB0
PgHIaTGNAjFkF3f0Q0lW2I1I5UFMuI5KdD7prQssMipe+b0rSHj1gmbEMmhmW6VNWMpU6Jry8bSI
XPp1nNTXTWt68FkYTmPuHDApamu4M8GzWLh5HGy9JtkCBnPwcp/xg5kG90lswTuAELG09vz0K4l1
IRpw5Aoq9c2gyxUt8l9OS0CbMQu7CyG3MvdKsL4dFtLz0oeK7gzSP0MMGVaab32UZK5i+mKUEFSg
bcWdHZSz3xF+tRTMC388v0r6L118W4yavT9VGw/rIXkiVV5UC7s5lFVVGt0+IaKvVRZwxPneiqdv
crlGFvBPCN3i1MCspjYbLc4PTpiWy6on15ECiJe0y1Rb2WPnXfwK/ZOxhGAJp9Vdl4fvKTOPT1xe
2MstdITGTGy5Er4nwYAQMG4kanQU+UQAHmPZHqhcCCil0f1rQV9NgY2XrncsitlMt6u5SDibxUnh
YIPlwkqhhGrocC27tLBu+x8A3R1N9I7MBoBBJA/3OncF1UzxkR/jSa6UVcA0gPHgiRwQFEG9wv6S
fxMikMwsR1775g1naENHOEV+D6iBjuq10lKzNeEWItgmeaLC8AQWIm94f5ZpBbU4+JT2IrFDsB3n
0gAa3hkDfNG374DigScYcdcwauxcjiWaXTRElHv4aLCH8882M1Pt21e1J7uZDEUyy1n3EvGTn5uy
RbSLYYDQTAundKuSK6qmmNP1GdcR5jqcBUzYcZ+65RJpOOSBBTU6UBYsdVCIOQii4WwWZ1fJW4RB
EXJ/D0t8Hfm43eR+2dW3DqC3S2MEO4duIYJ6dJrsCObY+3kjSQ1yuPnRhO/u/lPNJPbDRzKpPZ3p
TrtRlWAPQxh9NFxLLFH1Dh2VBN4i22OY3xNOJpeRE4vFdGdvW4xxazAVZfis5kaE75NilvJVVTVt
1JKGCRJmtP2mc6AYYL+ly8kuHxm2vwNToZ39SZfpbLSuxUszXER0QazJrULYhp1GH94h/aB7JXw1
ZYg3+347QDvn3VSTY5c28/yNS1ArAgKb/8itNd505owFHaHcfG7jq64Mn/I3QAsLjy/eDGumJG6o
1FNwTRu4KE+4BWa8NhCHJgHxQwA72EfxEb/eFpenTDdIN3Wi6pX8Kltlkta1YhM72NlAQIWGdLG9
F6zACWPa2QdC4Xg0gUHCHEKcduF4yT2p5wRwidYPeCdjJjYfylVr26PfZm+lA83NPBCBhe3wHK7F
lMEPOREAKBz1ia73cXl+7X5QiBh2xQQ6S0Vj7Wb4OoM74VYzVVePwXM6EAM7PGN/OSKD02+d5Rad
u495EY70B+97BZtVsQIMtWjUkqK1A2mtz0IsAErTXZSA72UKBXtszhFcjv8NoUqLjFwTuN5XulBd
R4S+ohIgl0cdCMJnRz7aLRRYw434KN/uZCgpRl5peVg729NXvC8ssZJrVEbdcm/56dhYqte4zFaJ
g95Wsyzmm6Y9RwG3/vklddGsIiHJ6AfeccCfbxnQqKzbWzVHXeoP+L0H8pukxlDttGJQpBST/Hpt
dO0Uw5Y0DoZGr/u41SE4XsXN2CEraHT0+xt7HafKYtgKlSjwYQ9zA3DyLWUcnBahb7yNUNO/6M2g
ibfFuU7QqDjSzgLEMWXizj81WNaYS9087VCrUn0iLG2UsZSel2vOIa9py83l6gDTvQf6bIPvdaNh
SuhjqKZmNkrxTM2vDwHcZ+Nr+xqHIZhLNLRuXuTKBELd2XsSD+ReNC83iH7rKrnWThKU+vx8MPPk
/wC442KDIQtik1Q7WKw6LCF0irnNrkhEiHCL47HRqoq052OvK0Ml/DDpBSbFBJEzKjIOdxNDL3HH
Tq+ZzlFhpoIcQm7jEhQlYE4kAZYWTA3pbNa9jZNC2lskfVo1jab5dstdCxMMjysB2PU/AAgQSNoY
7F5liD6cXvhzJ6zbtYitJrT0kqZ9n8mk5OLHCtL6YSF9MIwOwofs09tMWEq2yeLikODpseXBpoc7
REuauiUmqZhiTFrvF0fgr7myOSvFZ1YhF2WBHZIuonMw1Sv6wa+QPmPOH25yRQRGEBH7gHrPR1oF
+nyddOegWMMPtP+YDniLk9KtYSPSfKNWzmIIBGr/OzAxke5Aa/r87ShLEynhXYPCnftUx31gjXBc
Bhgpjs/5kNvQJlu/TcfTnPC/3JzqIOgulnJn5KSZxzoIIbM8tKZyByLV7wjglePInpTX8zsPpfIr
vSK+TGyFF/SjvlBfvhAS5UhSdUx/2eSaC++TI0cxrmDdaxTjfsNQnkaOj1EWacGgo1VLcHHPGsA2
91COPO6BcwN7MRo53IkeDxL2OYzNSAkEDrXsJSw4o/MNRrdTq64uiswDcQjPdpZd2jrIu3pEhjfl
m9f1BPV+vGP3kinZ1M/nyXNLBF3B4e5uOFQQY3r+7/fgCg2x4qPROctmq2Bg6RllEzFM5OirDDYV
jmBX3S38smAGP02KO5kaEU4C0P7Q6pH1UWHKpJHfLTj+6dLW2X1QDJTqBKAftslmlrz7FoePHq7z
+S02AFOjFDnyfZuI09CvprpsunsZ1h7OKH5F+PzUos6ttEDUNQbvOifwYe8OOwqH1Rw0kzSYCDrJ
6FO1RB48nSrVVbIjoB5eSdzX9Y2AQalUcgtwKAZc04bzunD0Jt/a6aHGuNUfNH92q5Solq+ilBUB
TGwFQ87c8sBEmVizxPn17DbGzLbj24ZVkadfym0OR2dczjGWOO8BSIceMdjiFI81O/LAEwNZkhB6
moVus/x94BcOfX/mtHvgWQiilSyjpi4cuB+s/fr4vM1GHp4Ztw6+BSVOA1LSthZxf7vn9XgUJ2Mu
rofwnmTMR/46g1n35Ogneldcr0NbocCBQNb6JKct2rrkv3THmWzQtyCuDcdwxbU4GIQyenM3Vq29
0Cc2PjRP6iAbQUkZt+DwWxfuyg2wfNXwZ9mfvqeEyHlpkaGeiERnr79c6oEyXUZ1LGaMtSPwgMOW
FkCRD3xJxybQsiNGI76WJLU40ExCQ2eC4s3j+hwM4RmHkMR/i4zSuv/uzAHZEBjHmh2mdb9apJYb
lSHvxKYpoDW3NbtSBguC9NSd4OyKnPKdyDchG4LMkKkVhfS7ZPOkaWUlfAttYGq2U1c/iuKiPuoQ
ksqSxZJLsDaCN9s6gWnHloaNRvVKqho3P167mRGJOLvSRHILmDsii0x5xSMAjuDX6nC9O+4LE/+u
V00i72KVFLWQCMpdQJIPyuG9UtUmF4Nvr88LXW9B9BqihbCMdSTH+yDrozX+QB96H5KuuxZKPDI8
u/k+8p24RxPvtHVkeLgVkQR/pDlvuaS/iYOcNQYPN0FJMjDcMiKQGuBnYA4gt7W8duScHXuJqOWU
YVxGV+k1a1Q9/frXsIGjinoymb2UvkbXX6jXaUCpYM36t7epAQGUwBeLtG9sEWrgFerPMcTJeeS7
72M78Ki0DO9FEXO/MKBuug0aHnsgj03olUEdGiXk/al2P3Ha8JTPxaT4qQKj+punRgD+AiqGzgBZ
bqEeIXOaBR4CZpuEQ2bgXKnjlFddRKya/aDc8CnJ1aFFdtJ7t4FiJlKFIJGUubnNmPG3l23iMt8H
A6iH38Pfwj2JNcx7OaNXyWEI5aUkG2TEHI/e3y0bGKL45avgZBHEzE8/DMaSFUQ3d61vcjbPWgLx
XgjLdnRjN/W5ZG08ynYdBtaarmKp9gWkgK1hH2HsIkg4ctgSXy0EWdrPm1UwSCjQB3W+5mUSbAnt
OjQ2jkxRzZLIr1Sh1XdxsmFBA/enTzfX6Z/RbuXPWIENois+jB1SkRkkUJ7aIj9/cy23WOWWsq7/
cukWI7565JE7yQGuAZZJTrpTT2xTvj5U+8h3U2JEf2lMvCBExXO8KIT1fUuo7TGTXuDEzNdWBooQ
/mrG8xKWinpB6qlkRnRC1qkhwy6DAm4wMEYI0Fc1CjPQlw6lyTC2yRdChquVdVbexPHWm3Fd1NUg
RslS1i9j+tUcoQMdJsrLKNJjTq9Fzk9cM2/xbvOBBCpKqee9R2SlNdqUyt613yZfTrQjCbQZRa+7
+3MTol5kjpLs0tbh+GPE0WmwMKpBSw14WXUcNwehtGfAiiVgclxCG8ga+ffZ68OepYZYW/sun9g5
zXGZU82GqXUxuWmL83ELWodBMdq/NhK5Tk1mTJPjDYdb5rNKQNkr52vqMiM3qdPoPyokdTBI33ue
I6A9h3nzVNnWfOi0Tj4gP1E2Rq/L0U9OQzKdU/yl4S6dJSw31zmpsCxtj0RYoj89HM5dhiFPfSlc
EgKHy0PuTnrW91kGH+okj0lvjxKbUfQIdLth91FO1jeeLARKX7NKtzx5dAijkz702RkXdESRdotE
qHOpNG3hfMOAoXmesTBH+BjoeD6yrbSOsiEmEPfzplw61iQmJXguk9RSFaAveeig0AOJSR5Rciy+
iKuOETHueYhkKFBAlVANWuklxbKbJZkAl8DOWGpC9QJLTUgdSiOdYwP1pzcx2inquqmAvJdR5FY0
UkEY+0o9TNmxPNlzvFwTtqnLdu8mMPe6mbeeQDiMPRDVavwgE7t0XaoopAbChiCw8dtj5eClfYig
MY0ik9xVpqrrUgKu6TuV6h3OFp/BrOwnc/h51rS7v6+wFSf6uVELjT50dTY8Cw6JnLg3sziqU29F
Tsq///i1bDB9bDYkq+Zp31M+3QvSUQx0/cs7Y5RwYtMywW/gYhFTvT0El3ZizX7YJ3NmfzGJrLKb
akMHbh5sqBLc5D6uHNvbGI7mzBJJy5HGRD0zCrbbHeb6fi6cTDijLa6yI07K4Nszm8Oq+w3CGqyf
B3FWab65hf8CTqKT4YmFoxmBKh+JwJI+Hz4URRrqMNadUbb2T8oKC3Kz+Zz82gJJ67TAKHlJ/Fmy
CLedKYgUNjz4p/nYCImyYETfn/ximz3vW+mk0ifowawHji9MX5h4nBqBNWsTee/YQvPEV7aCJn9B
WS2shRzSf5Flf6XG3ppEJnRGfCrxn3rkItwf20BoOitgh4jFDnUdRuu/eeruNWjFlFzKppX7I05W
wlvW5o3TiSGTdlEmzrQQ630YIu40sfPRkYHTGRt8cIg0rveGnkhOGQBO4XpJaO/pbMQqxMNUxegu
nauPdDhppNyz4zyB+W0M/2//HnoFyqEluiTvoDQdkWwJRIzpCxEmp7lsMcVIfVsaHmnyqbRPiHym
OCsflOPGQwT803o04/w5sii0qGKkWesdOqbieuuzlcACKOyTrQ/0gBSIAPwhffjQdSSWuqGyaMcB
w9+hCfunHw2QWZiIaeSbI7Hhyc/VgRSL9t52sFvoX0DF4GGHi0DoYTx7OFz/trI7SW4UVfvTOcP+
5eXRqg2YFrRB29HXd8M4yGfDdPqydMz51UqMYBDjmsOyZechGbMRGnQjqGBD//DDOHh34PuMRTwr
5LRA2MAyCqNmrqwjPtVLQTeQiloIn1k5MA3cpspVwdIwbsQ5EcFp0DS2tO3UX0cAcT3ICjqn9Xhv
2u2Qnwu6odOXh7qRgqhjTBKkjcEtFk5yn3uttT6pRttj4W53QyB5Oo/j1af20VztDiO828Kk8NPS
8R1mR5nJSPSEQJyqrWI1UnAsRL0MNET+Es2hGDsYgRXbnPYF4W6Q4JqjvCiWRyeejswTBSVsbKA7
49ekPyG2/JSD0upXysG/4dPKI+8EU5VkRsuMyuWTZTMqoocCz+yaYyjK//SdDfJmKeGNBACfh715
LCyQg3P8joN2u51LgJCu81cKSt0PuVXwLoGl7mHjt3MsRZCq1qSf01I2G4Npara5gWq526t/EO4T
XT3CO2LT9D3NdPI2V2ntHF5qsIWGIVmsHHJJRgyHeEaZ/JNEYEgYHF1elLKqoMeOnJlCXYkrY1Gd
iXjwkepJPvnAC4I4p/bJ/A4mF2KW4KnmvBh2PLAFEyJMBRkBrkp8n4dAWOPRSEbmYofb6DhXz9Hp
ETBAzpsNRCXBGRD+Bug/EUzIhxLNM0acJsZHlXv6JysZ3mY8na1hYHEajmoqWP/SPN0n1rvnLcP1
I2VH3He/fCL3T+jbknk1MAW4nh4UOLyGzh9yHTKxBspBnJGWPrsbF1p2NdxgDzBJ4PhIZz+SKrKV
CBl0ugwweIodieKPH0xMxrUSeEVkpyln83yMUu/fSsnr7D76dB2ldyNfxHLk9mONUDmF1fhdAB4N
LHDd7kBPlm3k1bdIjIUZ2dN43Rw71Qj8EfTjLa7vpRYoE2NV9RsF8pAZE+vW52gQZ8/CLn2QEMAy
w+6TRhBVdBHlUqqwvMpQosHEZUs/mM8hEK9WA4fJKxvB4CHO0VmZrUcejcwpupMQD2p93umc3af2
bVy4WZIQSY3eAcra4/HeH1yjphtIC/S0J0us6KMOnL0uGTJwrHBleYJZuyeATAovlA6YIMI/huB/
5/Q0xj4e8Zw1dErGVH2nNj05JyKbUjwh4xGesSUVP4pvxNbGeiZ/LrPE+sl31cmkG9n31poPXWNa
+vQl89G3a5mmPje6A3lPBw4qMqWN4rB7clOEoNikpn2HXj6KekbP5K3d/myEIgaCa3biOCjUYJAo
8+z4gCET9UYrzFKGkfoevySkXv2Yup6SjYlBqBEhDoZRJ4Q68hUzeRI7TrMW4zTtaHgSf5u6YZPM
GgCNusKL6A4GtjuzsyqdeXjVbF9UgZI4H68Qrg06hY9PEPJkH30kWNoNzdOP5e+oxMm8pm24hm5i
dgc3NPAp2zNbwE3Pmdyq5KwcAsla3J52J+OyUdqQGPb1NY4pYh+pTxNouHtpFWMgTrRYPjgl3AnB
DWjvCfz1sG2zkXSwGWr+jBISW/f83CLFEsDqir1SR65u9VCoiRtnbJmWPH3tvPIEc9HrFaGLprxg
xHpcUgq7ZwRto8wetlPGOHwiVuBZ/f6y5/k69Wya4wLLQ2K7xyA4guVgyNTRSXQPSOJ4c1WWdUMS
ouyMgEhCNwOX6mI3tvUSixehsTNWJSC0/PHxFplmBKCoGs9FH4yn4FdUpp9m4L5lidHddLNJiD/E
BNiaGsiGv1+fdNFKgjtuDqz+URhwOKGzlVC3lR35gmNrxoDI2L3axwsWlFjVi2GYH/Gn5WpNxbbz
rjvhO+2zkGmRsG1uTrwOx6j6lvnYxHqzNcVbXTfux4DVEQIKLkQ3S543O74VhhJd43EsKR22Pb8o
/yp+YCyiBcFDImvLiHRz7sBRtva90j1Ea1b4kWiEw3ugIu9A5mjXCjixa7LnEuZQhRRwKqhB/UA2
zf1fnHejh4lzNfybgC2B6yunq+XnSbVAodOFt/wruftsEghO7j111AdJVClMVVZz6/3t/nDkpF0/
/SB1c2f+TBQyp0qksttsx5VJO0vUrxg5vzKpIJzgksdzubBfCC1a+eSJaGnfbbK3JKnHYD9O7sYh
/v5a//gZeVPJ4xy+jr6RZRUVJnnLAf6/DGgFUnnTPUOqlf800CwAR6OEwHSYZsKXUNYquvEA1pn7
C/VbX4r8StuJaQ0npgbRHJC0i8FAlMOxs/uylqBuoqKBB2OA4D2NsuHhD3jxU8B9Zvd7CQd/+UF3
iSB30yrM3EsRn+EzikHwv7iCmxaHgktShS3HqJxxSuM8OkFiid6vgzz64jTEzLCFnu/Tz1zbxsCK
ErSiCdLWqSPw/dIZrxmIjSjLqyEnQnNCcd2nM/Y0Vm5U0vxsXbY+j45+NUvz3ja+3ADn0bSRAclw
huKkdjd8zVDyPhHIx3lMSVHqi16bOEDPhgriRSa77SfwCecxcKrA1nSx3KBIsvAzSxltlK3TbTE9
G8rVUFR20KtaLPzhUNVe0bXHtxJmkCfxgUaTXNJBnYKHUva2lYhwsFdpEDJzjyu3Dsf0Tdz6RQg+
shEyQ7E+n3jssBY4Ml+SGQs+qS7colvjPgdg63Xa79XGjW33a5AqinSuNvdfbo9eEwasp9PpSyJu
SjXM+rnF1vb56TmWamDanZt52qud6QIiLUGBAY055kko9Aiv6C2Vn1NkYcJBbGN6qCaB9Y5u9aZI
4/ADXv5QQfmfZcYwFaB7nmJOiM2PfHLEbFTNDhcvnabMBLyMA/p3pVaTDJ/NtsOk1dBkwJJW5EsD
7Qf9u+0P6mrUZfeNtZ1i1m8F2gjUAT0eaNIDAucj/LO79gjWi/k/0mKHNN9x+Psux3TUAvMF7kT/
Qbz1hbJDiYEEk6vIn3oMePhzHgTkvFok3qUsxo52EAyOQF6Jq5F5WYMXS/f7i1ik3J5ulLFgoE1t
n0DFwE48S4lfZu0pkdLpb0/qnIMqcxNxlTsJqPxLlZmltAQZBiWwqXdiNsOVzn8K7bYVYaqAm861
vHKaSX4l7GQCaVrp8bEjeKlxhMFS1C5QVdK/VmBn7Xbbbu1nPPkseERXE34yo3OrYlEEsJj3AokW
NBguYoQS5RE/kkV2O2sfWCSSW+t2UPKb+JVkllGzrph7Tr1xn0z+2/lQk4ECeWYDvBNBSlOO4+oq
Y9E2J0BZeMbSp0u0W2aVebSThQ8dE0BI+vFChtngoXbBUxtD7XfMCV4+e5SwpCrdwmkYNlRyntzP
kmWFMWaw1upaTtOnzo71TLKJUFyO1PZIy8xquClxqf0oB2lNxPiud7VivPn36uKlzws1ePJBrFgS
UxzE0dfSud2ddkANFJGLqFlvvTz+tHJD3vy8aoFIvV9sDQDiiKPI7UI5msOpix/7NwzGbyMBD+Zi
VOBoSz1+lC2kK5fuKh1CLlWdEqvSY+c3igRwYHpcB1ycK8ZOWsFZwqiVb4fFRVYGvxEZlGO94dZm
K+xrwggauQDgYzqJbcBqVFi9F4R2epuSxcEe9euyOG6e8IuUirKCw+UdAQdXHFQemDqeXJJKsSEG
T45wQuSS2PXRKc8RSfS9Wvccm28YNglKKNPuP6SiRyYHxsSn1S7HppFLDRqPmRTvEI6uOt/EpFWP
1WbbcguQWKhmi+INssMzi5rMWVD7m2kx2emlIj4ryv8+DfkDuUvMI4c7M0a9WZuZXB+NhSphoyzn
eN7i2VHxSOL4uEOv3DmT8OsWSoiOm01SirItpC5zTLdfiLiWfMerhHUGG5fOT1CIjleGcxBNkvog
HC6v0wywVhvd9vBtkejCqF/JSrGiT4KlrY4+4V8YLTdhkd4gWeyFNDU+DZAZJCg7ZWDU/Pp8oTPE
M2F9sHJsQKCmh3Z8QItK+DzEdGgaS3ejjMqHMoBL7xqZtttlpH66Fy9yxc1m2T5ziIKsTl0/mCZE
65+EWGm2Ol9oP3tgEHbPDYnzM4YCP/38qTP1iUOi+AQCMx7D+Dq8pTTaRwCxPmV6cQc5g3qq+7AU
HD7mn0J1B4j5UrjtNYCiau/Ozr9oKTMWonTPv/HxzLIlNVPwKts+Lf6PtD/r/m6qYxH5bLKWDN/z
viJH9WI1o05NaUGL9nf29xD8iUEk+XBoJkGKhBLSdZRQhS7t7+XXMZisVxPIGFVZt23/OQFZnjIs
jLKHdjBZL3ioyQk7Y319pLeL1HtFKRghr+CF9P7R5l/qdROvSKEUwXQPMbABCVTIaNKiR7mOVUBY
SdBDLnIr5AHyZTGaobTdGEQbfzPJGAArKnSuTeVhFcmZ96eafNJE5jrcR52CShrb5uetiHCP/M5s
cUgMwaIGZl2TYwykJh98rjmyc2X2N2qFZmdotznZ17HFy2/YOVkj6ZsHoR+CNewCfgQMZvYaSQXW
Bd5nuyE2qLIqIzJwYTYRf20PPKjX+A0jQgMdKum7NLXqZ6S0hbsypu0Jdu3oduRFcOm3rxlfDYzW
97dF0wMFFNKKCioNyRhtRieMQTKHQj5GXJZinS9wXdwYV3rIzMluF5gtrYchxUlBQjEHzxYf6Jlh
zk1N5izfsogLttXs4amALzpT/Oeffvy+qI9Klfp8yl5rTnQO+nUZ6Qbp8Z60CipjDg8dC00R7Z8m
IG0YE+JrYVnc6PEcse630t3toj1TSP07OWRLdqVUSBG37VrKVIhSctFUgJXoBin+ir1QzBnbIPAX
l9Jsu9gOvSCygrC58g97eoT4eB1OkITT9beuuWZtqbepBcdHBPgVNSWuU0Qoua19hEGPJ5pFuLZZ
vvkAlS1eClBWzXXv/PbHogWbzT+VJzVsBf7ZZkc4VTHBFzjXHQ9n7W2OtqevbnDbHaiGRl1EK7uT
kuMeHvYt9MUCgPqE98ppnsjH7L/vbVCkNCfm2kzF501bZQOjs4mol43eJGfmprigXIdecifFAci0
BQwXetwVnNZ0O9AksDOv1qz8C5/HIhpPBnAJrtwLGYsY87DA3PRMjYy8aGyyFdI+DnNqtztQf/SB
qd4aDlf9MjS2VxIBiIaY4aXxbWcjpKy09b2yK5bhOEQUHc2orhQbNXO2JCtqOq9pdV91CxyfFE1g
kHLCAEC/6Fnkl8aLpTOtxA+9nmXlBZJ1iuspCW81LQeWi3zdHEH6JKtIrwUq4ecRrmt86qCY9uSt
7e+EVBt9N+XIehGdT0eunqxB/BUCVMiJalScwkfB89wittWtrjVBMQm3ovrxjByF3K0qqBRdWaqC
DZi0fGrahS6YukYNvj2XtP/fyLHEcPpHPqTBziWT/VKbdejlusQ9RIVI+6GffTl+MC128zRDhnf4
LWcPgsKgjQmX1wp6dLvNFwAIhu1WnEHIHnrHBrbn+VTQvsPtkE0iAG3lAhPA8T4exS7b3yr0El/a
dafCPqf+71h5wr1a5xLRPgIY08dYNClNA7X4legvgC3DT6dRDaV0JNM3KX6SMMWcPlKo+/+31RU5
Kwpx/xkaVXdBClpNUZcQgOtFW3XQ04hXtr/z5h+/1Xv7mpy2rP/JyMBXBfBSljFX49Pb7iYWg0A/
eJLQ/FnZ8VJObp0z5+vzTg6kZSJyjMVaXmlWoYv1GswEDbm8WIigqSOGPDscLL/h99smqItXEhsV
q4z99uGydkChDlE1Tc3nE1EEqhHRJC2XEZ9MzkeT/1veaQVCdCd/tvL+lKU3sRuyIBtd/31HxTry
3qscC5ixYaNvmi0Kap15Moou2LqljAzC9MxFU2jtBujr7ab75O0586KKvQXZ4ftPBVfhWlraUPRb
ChtwgVjNLZNuUjML2R3lO/XvsoMacbTSnaCFbHHXapqCdaH5RVnJQOiEiYvWs/PrtuEbe0wSWNSB
NupPcS8JPqN1Pgj746ywigdxb9ZCoX0i63P/1cXoY6sh40sRGxY6eB8CtYedLQ7dNsgKOPrqElsY
6KZ8oNdqigpHr9eSKhnABE9hdLPA3l2hsnUH9oOQ57j+daSYjQLOAWKgW4hGWcWNpzKhClenVNFt
JG61FqD069eIoowV+tnz3dQxlFMyJchgfhlBHw5HdbQIwxIQs0Y6rFFgWctmiYENgAOVL85XygaA
6cLnTmmwHlCnxvW5y4P9kkuF217DI3gFu8NvjXgEuUAFiHVdt6VntXuVtDxx1tXON1ksMRTZreoP
t6D+pqUgpul3CTmgmRGs34l5FqvB3HFprRzpeKKP/hL8XUTS77kFrMNSDGS7gqGVPYrRsmXtM5K3
TFs/lGSEYomH06M74SZW+5D7l6V5yA0VOa5wZwa0/iw+fjNPDE07x8gkxL1cCfFdufxAu8YBOet9
LFRc0wwXAtK/TC9fXjw7tj3fr5kl+sQnHXoGecjlbwM5UBkfw+akTF0Unj/47FozuVP0QtVn4ZRA
0ZguxeoGbGXoJPvGk7p+ecagws2TgcT8sp1OpB/4FJ0MHvWkHMQQiUonvdJ3OpKIl5u6HdPbjQ0w
gwJGfezwNvWagA4ZQoH+inGXeG6KyoyihfkJgkSo5RKfwVgoeRAJckp7WjGxLrSdY5ZVD4UawHcs
NfQIv5YRS/twdLDJhbw5qjXjA+cqJDEN7bunSuiCokBRgtHhlUA0Z4ddeleGJExYpvJUZMc2Zggi
UAyc7MI/1t3iRW2iiI2qGNUSte7KZjyBZrmAnjnRZJoQXgMa3hKomSHIQDvhToWV6ILLEgnqL99n
TghO7pMtHgNrFEUFAUhHXu7L/2kANVbxhv95nA2nYxRGjfv5XO6IqhDh2DK+AeAw3gFL94uc9IAE
OnvaUDr0kVdDfkASO7kDzh5FTP8Qmf0O83+sb/iLwHOzer7GCpi4Sf16zqQORkyMIhcm8/EKaj4N
4t/HOBzjndQ2NLs/V+CzFNulTwvVuQ5Vp8qtQgqVxmU+R8BCs7AzQfA/6YXCixrX/Obnog7hU1Uc
Z3w0ubqMjd0T0I3yx+ybA/zHOLbBx2GzDxkJr3b73+JYhKYNQ83up5Z2PAEfFa7tCH76LxCkvaFs
EwssWC3FchLp8icz2j1AuiHtqu3LH0jlAaiiSxinr1tQhODAT50yR2RCxgAl6bH5bZJLb1VAMQ1G
YWnYNLXSHTGkRni1xmmyUnvCOhG054VEfBzTgbkL/PxhG09ArwFMU1TFH6TvUr633Vm3KoHMpBQu
mwJRczmHRhTfB7N/QBCio7LlkMqC1ykbMzLN2sZ+13NQvOggdvHyeW/B9H1Jnl/zTGp8NvYLTL+M
07qspeG0tot95Rv3a2ZWZAvGR5nx21bKjLDX8Lytr8Kat2jxjVubdMR6PggSj10XBLKAuQgZfHyh
IkWhRp2zMx1uD7UMyAvkuBDa2dpv5fj1XVeWiVwOP1EQAHdQzSMvNM3mnSyxfnMqsccuhfzPj5Wy
jbphSILYzX5aybPST0h1cSoxeqGAHgM72QtD8t3LsfHM6EutUk0RXlObA7KssbxUo8QaxN5+FALw
2IhwsL4A/gkUhJb0s+G9A5p+8wht7yzZdblChexF+9oVSceMjmDPOTm4SR20+NqxcEepftiqSORj
NLZF8x1SIFK2i/37d628XmsJPaZOlWyI98yRPVD+NKBR4Ki9gcY7eLj8FAIYZRYvYsXV4cprZkKV
w3bh6qOzR0N8ugzPhknUhBpO6plYvDiJjJXf97khwn4JawQvHhyiFazKcPYeaFJGGLl+p8Tm/VsF
KmWQvDF/X1GH2W8LMBocj2PSjIf9f4E0DBVf7cewq6RXGU75C1/BaKQR6dtXtJqTdrJrXV+ZvciR
ArsAPAhKVo8EBLcRa2bkJFczIu7hRdyopPHpaTPjolNROoaxda3UYSQHmm0F1xCz/rINk4vyw2qR
oA7PZ+t8chdSVcNIkhzMy1umNvYMtviI6hj+pgQPUjQs5kpAXVTufmEnlhXv3URiICE10WrS0gkO
Zuk4fjI35BSw6tYTNJqcvve/hG1poDf6fp2svlf6QUZmHhSqidxMfCjGd3T2dMplAwpkN9GG1CiT
+rAWOvdjEXWUIj01BweFj05Wohg1GmG10VyXlGpbPu8Xesd3vzY6wm9fos/+wo96y45OgATty9mH
n1uGbC+2w8p6jQlobb/waTXzrduGUK3BH4t3yTp1fEX98AIS/fCAWzBEzYDkiEIbMewIperq9Rsy
Eou1rEu5yEMYOxWurCRmH/Vfj8Rglbr7onEGPMKKX5qKLEPr5et/DrqDuM8MhVWj82j9x8uwJu5r
6f0/b55GtGY9XT/fgV3wn9fYw7GzJnvkIg3EdNLX0i7MN/FDPAiCtL28N1uD7hUlyf8pCGZUIi+A
4H6INlwx0AfQ4Nl3HwceL/8M5QkJBlcSXBSrhqxInc5SmwHVqzmcmzH9hBDht8+YcsVN37ZXfVLL
zirpajOLHALoEAKKPr+dttRUGO7kCosPf7kqzHypntReqZCQd3sp2iDVGdzv/p16+gx8drReqJ4d
0BH8u4nmF6GCG48Yp7RDXUKRarQxK3u3g4HufU6MjDMucXFxd1YX83+1qAeA762CleVgfnWgBTCI
EfKnycaZlV7SuFQyJFC3RXjocDtPOdPc2anWDl+wpM3Y+pbAFQutKDHSFDk3Qe3by7ZfYiQDmrmW
i0ft8oypyCkN3D8GrOZRauyzYCKV3IzUSO6Tbqb07hKAM8U/4e4UOOtNJjUFHQkejchBxKnCKNzT
RcNG+qkZD7lDjiaO7PWE+mje2+q2wgDGfyVHbnVYbKkHn3AYLKkpBQXF0M5H1DlYklmvUDn8mIGh
gMSKsSRzVw+GGQ2TQHpcuarjGuLcPAysxT5EUfKzCXl8RktTB9tWjEObuxO5jOeYS23dEH3YyF3J
u9jbtoVa3u51d5i95h9ZW/yjx/U34nj6h7AodR63GTQxMVd5ljDpsDSEMe8odCw4e4hx7zhMJhwX
8pGBsLtDJSmOBFYZ/2o61kiDRnTmm0wqDDto5RGH02UZlZcSPy54IVk+qH/kZWrj54QczvQb1Dc9
WfLrSpjt1XW4oHMN3iDu1tW7Yq2ABJ17Cq0BOJM50E88TOzqJEMXIkxTkfdPl6Vbx58bxC7zJo+U
CRbqo6lAjUN25UwJ4E9XVfmSyaqlzo7f2dMI5IWr2vmaFPxadBLUa2O6YMrTeLfpBYW/qJiSYmp3
n0o7gWbpqufYr7aHcCrQ0ef34QOPj2h8XQOZYjVbivmPl23aw3ADg3UbXVpysoy9SYWDfoyEV3Sk
tIUVOMNqwgcx/m3lS/sg8sob0OAD4sedmTB9/NwDbbnPULcVBYHKn+oMDHUCvR3MPVZ5wuGQZodK
s9+vWgMccEIC70YiCCQI9xqS1JmWz2itSAB9ql/XSRnHIDw6x0Eywgp8ewH7haV2VFISOnL53fKP
0jvluOsBfRcdaCmvpZgxRvWhHC2GzJCek18IWVQoQakwzIDrulwfZJluaC963toamod8kU3LgLDO
ICQObc1JgFqxhg9qDIUdJvYlQJ6mdxL/+6QFdcGOrPqdvFDH7kXW3fThABCnPxHJndmiE+zBn67G
hhdbi48Asn4UkBWlwV6BOKIi1paoOGig6HMcLIPgvmCV0Bd+Ke2+Nnm9IMu/kLEO78xm/YvJ+Xk1
o3bg1GR2mC4BjNKlH1yAM0bArMYpWVJENqkSWAbZjztxUkLi3keLSp3GgqUhRIGN1oEutKSdt/3j
qc1T0OBXaeQq2ZK4JwLcjWgQHkAd3fmdYur75X96Fac26XLClhMi4/iTU4iv7pdEi+Z77n/P+29G
aYC3vT55kwEf4GWDma/nl/vxsj+osz3aFh9b39u+1jX3n+/LozNRXeqQqnLNThO045BLZSJm7ui5
O1zvuzu5p7LgC93RyLhv8Lk+mS/YxuxcCyMLUtKoQJEkQR2VsPoB5n6eUd5Ft8vpWZ13XYadrwqq
3i0QeFe5qIa75QBlAI0KzAOtltYpnxuj7h5kRWLOL1LGhC1or6YMVuXuB4t85vpqM2rAbid7mEyC
UO6y1/fO9BTKKDUtaNqqj97KuzX5Fi+//Z4W36J8s8H6m1tWbqk2QNg2yvwzCCfvEU40dt4JxopY
+Ey/PdtiasWqMB+s8Vxh71s2NhUZhh8KwFACeZMhV5Gx5emWDIvIoX0pVn+rHuruzoOhGl9mi6SM
oxG4ecvHoIHc/5uRpHD4zJi2U9mEjOWq9LRk9n4CrfSkkOjOuacopJNIo5ONYvfn26XWuY9Hp60l
ZLYkEbAE8CxMR0EzkCtqLv0NXhS7X2td6Q1RX131sBJzmuOlissiOG+OBGvD95Lwt6AjyTISzqt2
fMT1Sa13gPFySWwlNNr4nuQjrl+CXRhHcf6UQGH43K0WzHro+NGbYbdF6QU8NwiSHP+l0sbn4zJR
az/ESxgVSSqfU9QQDfDDI/N6vbr6Marf5UlUzJtQe3x0D9DNJvqljfNL1Llpbjkb+uUXQAYg44yn
kYu74wvblCGUWSYe4mk6hhRTl5C/NOBKQtY2i1GmaEUY26961WgNL/e1NMp8fUB3wba7uImeZuZ3
LRhfh9aeSPXNKa4mWllSyQPnq4LH0eiuSClSFq1AFNDQfjAwKFPWhUkpIWeT+YA376lKLqOL/b9x
cenXIGU3dglbKHM9zVzxQ6Qm8jqdySnnu62mOnIDQt5ytI69s44Ma8KdjqsBs+gs2rOLWDCF2wVJ
q4jkcXne73CfTOLFEFDPCjx1ic63RVAMDJk9TgWb7cDt5OhU9XAVSnH0lVTU59NgdKlfg4DUb9pZ
YcUu/GJJawuoU6DhOpOd6wm122AD/I8WzWBnsOoct/8pm5T2SLDJJKdT454D7/OnbWT0iyiqV2kC
prKMEUOsfOf/0ghk5siEyxdzSmP7/3v1GjzsZPBn+Zz7ONvn9fHVzBQaH7WF2iKsaxuhmE8DGKlV
zxPjJlVTfWl+5tBfMZ25lqtDmCU4xOvRAN6AnLaI85bfkJD2E8DFCCE+Ev8VG7PK0g6C3QvK9v+X
d3dPUxhWCGCpsfyddsVJDPnFPT+DgQaMAXX2zIzTSTohHOflJzs//LOHfQqOWENfIk1Gb0qCfipi
m6N3KdMA1cAfz3SWGrFiq1wRNldiRbV/K5PHfZhcClIo8c6iBXr7TmiJMFnwIAkD6492xwJE05ur
7JIS9snPuhfN/Zfflc00CfwIBG7GCshnr6Dwevo8Hu3FRoAiZdbGb+1OMce1B/cWo7Yt/LiJP876
WhFKRoX0qerBi/NVzCdt1+XbOOE2BJKX2NwiW6rXVapXSV/pmhvOoXMUNf6y4CpLck7VPQuaPvHN
QXixwFVGxanUEIM7L6vMjtsmNj4xHUshWn5nVUdx5WNYh/JajUEPUSLrds/+cTxkonIQ4IVXhFHw
HcxVxM9K1lk269MrJowGuoYIkqhk9Zcnr7I6qDOvATr+wHee9ZeP4kzpvA+TbSIn+tDfLzCdhJeW
Mw1wdDbMkOp1zqN35cyEkrq7pU2H0jQTj3WHv/XhLxQN3gVixJ0Dh3yJ1MjvgLSx31dlRWxB+Q4v
2ogaQHy/5V/Xx2k/SdAI6DKFgiwJYea8sLId2kKsUPckHolOB/8QERugWSt4yvFTPfAxg0tFtxKp
vF9rqnhn70f5yd7H2QbLV7XF0tufEnpNJ0c8RkuvgaUfOX3L914hHwsNAB02bac5RnMpk4pxsiwV
DX8/vMVtoSYVoifXdlTzTMmTW8OEf6eu5ivxSQZCUEbd311hFdYCL+wyOMEHS3+df3EbkZ8IhHjm
t8glwHhWlGHYrXM4VasrrMw1FKHOYD+ejLGyLl+4U+PymWwy4mBXUitNFxXxr9m++5X9MJy9W9k6
99IslRnRGJcCUlI5yMAd/qtYWcTukZQlU//4tafz9TX8zjTWrVunZoC1vb6omgDCJ7EuS2dTbXX6
W9hPrum+5ykRcmJEoCtg4pGXb0jMgWPpeo+xCrYr+UYXI7Le6hcWz2qcTOnyqSSt1342mZ7oyEpH
pPRg1DwRLms58EB1zJRtyPo/jO7GucMc/l+SRh3ljD9VajKTsWXOy057aB91OkTg/q2tL3IKS4s8
F8JRzktby7tDfTHuT6SXcFbjJcFPfgc/yNXRxvsSuyQxrJFjwysy/U30MUFxsKytrz17UhYU39Lg
WqncJGpX6vt2botxSick06gLYQ621Ngnvi3aMiQq1nESE3UyIrrJjQCkXM77xD2i0capPJZi72Ps
ZwI0j0j8Oqae8en34VicRN54D25ozM11IpAB14giRpsg/mP49jCcf5YgdO7IVmQPgYzEtV/pKf5Q
Laubpm4ksWex0JLnMdoeQu3gW0LHj/8FbYZWoAJ5SUUY/rEmtfuTDZfEowLTmBz6Xe9MxXXqwzXE
3m+aDVIoawNYRIXgAVyglY+q2GPLUscBuo+GNX1EYzuMR21Zx5rWvaoVXNYsf96kcmTqvHx/5J3A
Lj5j5oVvHw/KI2Ul28zOtPrC4pgOOH4pt7QN7QpZgV50mCmBM62gYYaY9ABZ/t5rtAWxn5/o7qOm
w3bHOZNJZi0VwZBtMqajXgIed2v48CdDmXRY0K02Q3G1TtbR4QBEGRJn41hT2/kQESiNoieEZM08
9JYyinExGE43g5F6RLtkUHak1wn7wJY7cJpe24hT33looiuw+n/WKvO9C2t7/23DpeW+wIJVvl4o
4HvH7QU2qeTe5uiua22rocz1BKQgtrlY5/aAU6wbCaLrsIXvRJRELMDm2OjyafxAqareuzdE+7/0
IsgVk5DfZS/xvfWDnVLBRPWV1G6jZXQvHiX/kOfZrtqiHQCtSS96Vek/xn2MqXIfsNHov+dt8bzR
6GYuircfU9hEjoPjTE0nE6elO97ieQ26cHwvL5T2T5exB1RDip6FohltMu1/Yhn/lbySDU9I7NQD
6MrI1ct9VamZoZ7EH2irT1tt9lKS7ZI88tjXrolDdTbkOg8ikI+qSHCaQa4xFS0MXsuqHodzm6PY
0uYmhVfpkHdwU1QJ7RyKNC7WPvyYvPP4RjLILa1QHe5QGubVy9wH5nfx4E3zodOsKU7dDXUoVUk/
WQHmUl0wXnlCrPz1ADgbQ8MpIYx500rRbJOjpyWbVvPlevubTEAi59skWIEHsaYg7kfMPBgb9Pxm
jirGke/pWH1NoNR5Tid3o5vAZelqA8VPuckrsCAlYa48BtOpaUJwEr0vShzGOknpEpElK3g+ue40
jgvLc9pka5syivF5Lk8b2LvER5rCwpd8JI2+LPzslGjJcJ7QdI9VeQz5eq6TtCPJ3ir8q2L3pgtw
IrDtGOgIn/2+6KkLmxT0LCiLyHR0Q0ryn6Xaj/VkeRMQF36tY/3IR/KlYmDhQ6FKfp38zgtanIy7
gTg7v8S+hS1muAW9jl+EYcBbmuItILUcMQZsBrejHsru/bywMs2U1PAVj4C+h9qH/1W7d8vl+GqS
PZcyM2lpXfllwTo6tWQiQvUhqpPHxmo5hUOoRCkQhWma8zBmM9DldJYCZKeJgPd46hMIC/FxHUvs
idZX42j76OhvMnFcW77yHSf73gE3zDm/L+pUqQ+DLMK5dgTLck00nYNKArh8xTGuDjtPwpdqn5za
7XBMQKLZTVVmNAxFGnkCZEiki04rEv1Sc4wvkeTQ7Reu17OVAgVDzSp+FEEyI4K4YBQ4OxXexnWd
bzF+FRSr1em4pr+nMGLepatWq6hhfTDWsa34Xoo5PTOzyfRLH61ghoBzYcz0iq6PiVW/UnOmGIuA
2YAKG1uff9ynmyJjvuoCaHbYe90JcoO2Kr5UxIpbNMcreCnvzFI11ijZe5r5ctpDTY6X+g9Iudk5
eKMCw/I0r7hIA3jQDSJG5StqPYpSesHEf/6hMpnICJxnRsfdonSkrJgIzMhnh1zJwHwtb9wtQvNy
FGt7Jk9ihB8I9JOZ7ruhFYBcz/sDRjlJv99ZSMRafnlBIXFRK5qN49ObW8ehpjn6jeTU6PWYl7TS
MjNzErNX1cwvEeF69W3axB6p9OmxZn16YEGaOTyQ7kNaL93/C4NJRBBFacHUYGau+Aqba6wmwWHw
vsh1RWfYf7bV8RMWTc5bADTnqiOXzoRNOUOybBYtXv3BHng/hYX+NGrYe4UTn5+OEZP+jLMhyZhx
CCp5/VMm+Mbe8/zalsP8e8RzasaWjMQvATDZbfEd768xWB7YkEF4L22uYhMR1+fs6NFsoDiJygJo
Kxd10q/jijO3gYEg6c+2IIzz/HWTvcftR/uG8Y3hD+/ha7f5Df1d2GUjFA3q2rIDrMjzcZALaXK9
lNRDEAMOu1vrygDPDHRA14bnMQTkWvA8ZiSir3e773yvmdbPYqMTM0xjbijMw1/MsuFI2ZnFESaU
QjcTzZ1kmkoKqh7GrxJl1GlvI4JQNuMD+eJgjsETo6BU2D8WLHo8xXuTrXYSlwk0vKvtoj0pihZH
Q6oxXF9Sqaoh96jtRTDENDdm40DgYBl4LD/xpn37V/35PgOeVHSC6P0CWK/1P64xB+eJoarVqp/Q
2Ty0Q+L8aRcCPfStUhaCOUBFm7ELdx9+p2gHDWtuajKdMGeF41vn2tNuKRdlb4Bk/iWONp84oOGk
SHjAivLbvLJ6u2l9m4zWsR2fhudgK7/lvDhj3t77heCCa2rnxDBoKVB2Uyh+0YiQxWaK+W4gXa9w
Iotkvx4U6f5gXawhoh4e92iCMqGRXgC11XGX0c9q5BavJMOXpnI2bDvkCgr1bxQQPeJWqmUDsapH
7feh/KKPQxcEMCTuLTlTS1wlJBOqz94IIYyZOSyBj89RwakfyLnOtCg3xrmN4GFRqrbj+4Id9aqm
qE5BmQy0ec2JR5MrbrR3TQC49x7vy3Lb+i0Uq0Ys88awtioPFPjEAYMDMj7LUSxjLYTvZhVN5A8S
Ojo5m+6QpvPh6JGOVAdYTogcsTrVdyNgeT9GhFhEUymL+HnaP/WSUyk4nrc2+RnRAM1ehJdpvMaQ
m0rP3Qv2XAOIfJxDgGm4oASV2ELQM51Yvn00jiqI1noBxKLnahBMbcN8d7Jrvvs+w8gsJFilIVxl
F53muTcKRN3FDeCQfIg8fVxrl9ZKiZtMklcsrkYG0hyNaIiVRyflCnFa7vkTJETFwvnOGz3gkUV9
AbKpJcXy37NE9k8g31pW9AuoNv7f//PEM39bVlV+zU9W+eAQtoTKTXtB2dYFolkq+N1mhtm+sxTE
lndk5gU3lt4CCFzCtSm9RMtGwTAoRW8W+ZkOZUJTKinrTDGkVRHa8cPyPP+QIWeQjFnyIN624Cft
10SS5sDmbLOEWyvUA3kjJ4Cs9tdo0TCk321/SdfIZb2UKYN67WHWlR0zTsOS6KWHnMB7Unj2fG9U
zxn43Bf9Gf2B7Piwzy69Lf27seHG48kBNQJWixn906KQTojXYDwcKiBrP48KV+lmtrOSIVYkTtK9
MK7jIL48aIvGIqeh+IqqLzcU1y4HaqzODPLIKBBz9ij6JaNUCfPNPgJquYcUNvnhmXubvS44LUuR
mXaynOfhZSqccx+uQ17CFxuNnpuID5KDD1DI2L6l4FUVZpHYl/5t1BnYPrJRcrs/ybbAQrIirYSa
2NfDc7GMZEXUhHkVXMTCwlVPqUtoROqLB6ahuwZ+L9gFdd4p5lR1arDzbfrJwcpDgAXNOTjmDixd
Uao2Rr5gyjhTs0a87qlgMoUlr1d6/C/znpBZweRv3xYvqHlvPzincVt7EMFGcjjDUT3o+ObRCkeJ
AG05o0mgd+hCkYsjpPzBaSSOhu8kb2hNXIZRtJjwY+DtlTCH/K5ytMIR7MPWCuMUIdXvxRLfeLzp
nyDG4W7+maunsV99rzTKFEvAe7fkHvJxltC133DeJHf1pDGaNqLUZDIrI/ibj3QTiwA/s6/zT4lf
hlF8iR0JmzHBGZwRHVPQAMsEpPQkcVw6zMAzwXvrhM8iM57PhDdGSNzgr1DsPoJZCuro8pJueAfD
Y7hwTEfE27tM6muVeNUUEpYEyded+N/S3bsUxSof2wydT3NiM2xBIVpmL7ATYsLt01G8CZCgZ8OZ
LbA24NBGqem9copP79WoGN4jqqLUaE+16YItuHqsfoUi7yaG0rT8KnugWT7ApUy4djb7tIeiuQj+
nUOnGQV5SHDmon6kCDININX8Doiue7J72134cocn+JLezVOmauOTDtZinFgqK1wMQAB3abWb5u+3
kUEn5eLgTKZVVRQWFLE7AEbSpMRs3jsotQ+qGUneeljqSMr9Cjl6ETf9YCgToE/aDtVb6fmjR+U/
KalemzeUeVuKds2MvB53Q1uAmXxjQGyXegZjj3KoFLCmeKAAGvqxCZwDATygXDQl1I3puHP+rnLj
8eZCSRn1gsLXwzt1CB9zg1rlqeibkggvZz2HxQofSxXAAAvzMQld34WX4ji+EFQZllv13NhtuNvh
MqqOhlj5uwy679Zd0jUblFKB2OfhiQE9CqsTeyswk4rrj9rghFqtKP8iZEw1EH0HPZmyn+pWNog8
/cS/ZfR47imteGQWUHz8Hn7go0wj0GO+oTMwtOZFZeunQw9KrBQxCcUB5rm9yKK4CkmORkDPJCVZ
HdZSptOG8E9+207UEKRJWcGF8lkz+2Lu5kklskxuW2WAY1nsnELJdHOwZV1vAIfVL+fOm5A0OsqS
A/yKN3160CTjuVAIyUlRVA7NPKiciZslaIViUn+eaWZAZF5zyuhIkVJWxsvUv6c0QVKoh3BEAxW+
AYahDv0l05MJ8Ld23+4jYlfJmv/Gvnuj80g9NMBQnET8RA12JBJegOG2gskcbGyBMYZVWX3/0RWu
Ums53GvSEuVmQcj7zS37XA2g3TGfPbX+4NWBXqPKh9+v+ozmIqkKvxPpoKz04xyjGckjohXhtbdw
nYIPUGrxLuxY4pPAoh+/fCUO/8uAtwVxkbW2owkKerdExAyGPxODhJBxYkDqzkh9Khbz1CMICY6/
moGdaTQkJKjI37zP1uwhthY5nF8soUlqrz0hTACWIWL+sf53ZT7ItlEY1JIWAjyPkxrBhwrPgex1
I8K7XFwWz6N6Z8+eM/iBLTUcn3YqbkmGlkhrHj7D9qnGHqvfRRT8pShW/5oLogBEwCFppfQo+KCg
WSpu8jzggl3fo0JQFnQJQn1SAEn8/jXimueGNXrHZF6doShfZyyePLdvaU79GKvx1XmSpMWCDYGi
XAUpNcUXUyAz/nwh6HLKVHU3FPerkl5J0pbXgqyhO0vcenfWKlWzrtFVJqaFM78aNquLy05lANwg
3AVtx0XPXo1p5iYfW24OdBZ9aN+jZXEf86JmCERGs0TlVxenVqwqpHrNFRRQjpFomiUpppVv2pVL
w2LhAZCUg8c4tGfoCxrQG/g1HxC4iRxczeYw3zcWFRfmmjhtYDU3jKnU8xPawW8782jqqVDaDvL6
2au4X7tW1IuIeyyOELUJxYexGWNtlK2jjPPMEKSjWUZMxyEBOQh/goJ64MVfPVDqnN6GEyodpooH
d30lyxAf0oTROwkUahqiXO8YReWViL9whHFJGr4KUsJgiOimS69n8SE8ggWU9ypSjGEvopcVlRqq
78JZ0RoWoXPHmILGCWZo0wy5ackOFLRhSHC0U7Efo0lzHHcPSVWPs1i3Wnx0vrxGQ1z3ooqEOEaW
+ZqXFK+3+GWiLLW1HmY2TRZpAbYcaM/hSE5W9VGp7TN2DQZpn6IruTO20lXOaCh46Kr/zdIZ3cNi
YIENrWG9seHECnetB0B4HmL297uLxk+BLLMRn53++Ipb8V3dFN0E2ezFYPG/dRtlj34lpYZqbXF+
l96jYzc0ZTrulubJDyoGbzxid82ILxo17P7fghEm8J3AFey5B2ZemsunOlXqvEJ8WYo7ixxJzIrp
wttcNLEUSsPTEfcmy2Y1kCPEn8P7vASFIYwu97i31Lxs4Ed7AOmrbNqfc8Q47KLCK7cJUTvDP06e
/si84Ac2ZYKIDf4cwccCZeoebLUkLQvhXco7VB/VIjxzyeEoBASapaT95spxIhNl55bN1vs7gd0X
FqtSqe6vuCQnlBRO3TyE1zZNoqtQYbmiyWcNz8yrh4mUuxoOCFXFjmA5YZABBTzTqdAoufFCKHgM
ZkdK7914QtmRW7GJLrJedMplWQxP2tRQl13TaEOhd1Qfb/vSLiF7bsXPpLzydwavFkIFc6QbZjIO
A9lfmDC/6cbI6bnkuRLuJ5XG4HmTimjxdTChneEw6roohsgpN7Gb9je8ggyoTvV3Un6weHE5/mzq
dh3Ni+DAggaUEaR+D7UrxfZzcw4e0tln5RBnXzHUia5wpHrZmmcI9Fok07eEeexQmAbfSKsjbmTX
aqAiEp5jMZMN5exdnt4TaV4iUofd6r1TZ3eKEoNcEzwl5fLNVHwPFfggsYe4VnvfBZgTlEXzX7F0
vDPMnIweZaMUCmb2SQiwIy58zxszimKFczNmVfj2srPOaqiyrUd+d8fmnBR80taylCy80Q44Ajz/
CtultxC4ybe7Qm/7xnSNKCknVof5FZdRjpdjoGN9YmRtEjQOEmGPhmjonPcwa0aGYOzNsc0zhUbF
P8NkCiKUFSSYWLRPugqjpwUTUnPY6hGnyHEo8Igl6JMx7Ng4AZWK5Gy0hVWt9yqPE1WMUP276THi
lNLkiCZzWb3QOQsA4iaiGYCY/aI7/8ZdkzOOYh9FI9zKFnvA9BS0yYNUq17QuHcIFRU/Tc2rrlF9
vZMaDNik2brq1SY4YKhRU3y7/k8qhnl9A6dflUjzTRZ23MxRqa95GhXy0miFV9sRC+QVatU923iY
VJdl1kXSyVSaMX1Z1ZgHc2AMoif+NfSMOrK8VsyWj9WLtycdPfWpGOhHT5cp7fX6/xZyNmxEpoca
9OzlQut6tpytEhk+wbGowYY5ZednAosf0t/qvXcwwb5h/lUV9VkDnbRs2vK+dSr0GfPXrQJuOQSj
pZlg2IUod3DRRpJmMpaNAshF/N+gm/wHl56LuA6WvyY9dD4Qu9Zds/TxJ0HnrmUA/wDfhP6BWo9C
ZkMcCTHVzY/kDauxhtgabdIUj7BGq7Mbk2uL1PQSbruAq+dYnMXG6Ij20jqw9cSfhOqIctEkAYav
1ckWj+ICERSVdXW6YNAvlv7E4gv2AEBvkgxGiVtQi66ZBPmov1+Zyc4NU5lAQu+NwzoslRa92vCR
UIkN7QsZUEjUmPC1LjWBiD/2DB4VkqYoJIsl4hkN4OcYpSsBdCWsMmwp73EfCUrIznNtbgBB5z3W
aOvt+B2FQr8xIbdFIqrq0mkOx0bw9tPxM6HmKPRaKyTF9gT1vYr0kY6da7faTc0hs4FFWqH/5Vdx
q8PFzigJYot0rKZ0At2iRMSo0PslIixYMdUTURhvlKHx+tJf1SkXK8d3eNRVAcejkvhRthFf4lFR
vTFkWwNbTzHelYCKs0TN3CANWOksRTU+PXaGfrVo2J4Tv4saX/bs70cplIAyS21eWgCv8FUB/bje
JA/lWgfo8ZUWSNNuikzEJ4Xql7W3V88ERuu8wGobW51DEd3EhNCyfI3b5nbCUpQteQdK/f+EFI+9
9fMT+2Gkl6L+nuy6GwSx48YxhEBR7LHA6EzHsMHYA3O6rh2phAgDjwvemrUhQm3lHhXNJe8pzDmo
eZKTkIZ7P3DhdmYBJOxSZzzaSIltMR/8Fqi6zfCtZUaRF2F99E9OjGObg9TqKFYmskV6dbH82/Xj
Q1jrPYc+uyUqPLBlNrienSeN5WEvY/4p25JA9D2DoKXASqADfrOzKCgKV+W3tDlHeUMgIff0ZfDS
7KrNPwTUYHg65KU1t4znrGE+MuO/j3hYkkaDfp+ciZ6N3tt2PfD19KERB8shfHS3n6gCpKZwTO+t
XhYr8M0MCZp+PnWl+ODADQQ+yrhw5ZFCEBXOWKKAX0qXprNiHl/ypjuNC/kS8ue2CFBEHUuLZY1a
c68RuXYrx5T2DnnYI3I7OQgIIvR1XNYpcAs3+r7G6w0wekkhTuh6+sVH7Fow3yubyrRBo5yTm+5X
YEG90IsFH9ktO3roal9EGR+dJNT3/K6GHBv1tsvYqEPPzzhj8/6PYm43TJblXfQ/lO3PV3w86nsL
CjImKBddeU5X0Ht8LLvoe7TO2fr57QVgmjk4TZo9FYTgbpj8glxfvPlC+j+KZdguYCdo3bhOypOi
wVgQc2+BabRkQWx55VA7IAX6YZEwhyKdVOMboRN610IpBz5GRiIK7L10z7eVaCOPDhh4Y3DNk6SG
owLQ5x+4opFjLIuMk5H1sVfkfm1rMN39ey9YweFIrqym8AVKMjeiHjU5lta82DmZDdehYj3SyzH1
PSgHDZGlVnMpir0aYJHE4GzZ/IN3RzIyA8URI/ctqWitp6VQ6QpL/0iaOTQy8xZS3Yz4StvoXuYc
KgxnHXDJoX+2HQxuPPMUXKeqaUQwLmyA405X/mKVcUD3nmcCh31xPK4ztMJrIFCyDip+D25rsEnn
3CBvn8hODP1qsY2W11HnY3i2Kh67dVhhOd6VgM+zaa3F0rW+10GF6askfmFkZo+7nFqe3qc/WVfd
1b7qpIfI11meqbxcD0IMAGc5e2mmY/oRhy9u/Ej3iJgfp99aQOh8RKr7jG6VjbdEuNPx+SvMXVF8
bKZej3ZVjEl9kElhNwdJYH2VqocHVouidzVouuYhl5mj1/S/gEgBGRvnQSaL1H0CvKXqAY3ppkpQ
G4nDRlU5oWstRvtTkUMaOX0JKfuCyH88j6sLbBzU/Cy/rh2y31TWKIRRHdOEHdntj7wvudv6vtA+
ej6zBa9cCttGsdgaeGwoiPfdaVeWV6z0bYWwdMdxbPYVqO4KUj8BKR+TKdMCq6TuRI62Bm6r0mzz
lkjWpPYva9+vL8ZJ3jn7TeBtiHZrDULF3CzO1JBuxuouyzA2OBh/hCURndB1yrIndDWptt3pGJZP
R7195QWjHndT551El2Pzne4vyhzm5IGJyl+d3GTQFnk/aS9iJFXhxEuWbwKX425NDrHy+Bo7/mSG
MTXwGV0Hr67lI5WCN9qlmqyZGCA+w0XdPZumzrxhwSABW1OQSIQd9S5SXKZj1x80vko7MpEzMLmJ
ris1/L4aC/RJvYHW08qGYM+j15zOAQykhlxVhH5elVFxSUqGicjeFGgl7hPxIzUM8yinxwWawR6t
+ZIJ0rUTkOGCwUM0udPKpgVcE7KxeK0JJda6/746QE1759syB6bMdG43phS8QCzftyyY0/Ss4Qtc
IhS/La1dfSaXe0Z0kor6sAlGaLRMGpq13o+8qxB8K0lE3clnGyuymJhIbYW/oh4FtBVy6vz87gKs
5f3QjQYiC5l6HP7LzEjEFAa5Duf8aC0VFHkW7q+ybhFU7ZVnxn7tZrP8B+i4snbBKTqBhibZDZrC
J8Mc7e5u7whjLL4c60Xvi5SyEU34qGf/Izj8B9xGltUbcO6gK2a+oofglkxHcBHAVNvj4PpZ/0K+
KxeUhnleCvkqMRMf37iSzRHq4EkGTppjD9hndyryfpmQ1rst5i/06OD40R84EGwSl4I11ug4ONdj
H9BoUcYl6vaMkgMvQ6KSRTR2Ud9xeZJoKLx2NppoFLsGEEYf9QwAvz6ljRGocguMeVsSJ9Q7dpr3
wYz9/RCzSXuOWsWULGkk9XKfGR+rbbBd39n6XcLjykdJg5trl0J534YNd+dTXpTyN2ZLLGSPKz2V
2Gp+J1ye87AFUEBI/wLoCuDr5KD8O/J5aeMfsFT6lX6pEQ/iStayXAps8kbEeCSmn04C7xL4mI9g
vQwH3PmiLvlmEfSjKeEERusP6TEb9jm7BnVJUOO/Dw4JyZTsp95p2pD223rWppDo7YNHZ4E7ClyV
FbFB4aMMdYvi/Wp8wzCyBGhH2cWqwuCauul8tuwFdUKBatJNJifIZY8XrlRx800S/cq3qXHu57Zj
7KAZXHl6Uyka7yFdIROEDtGdKHd9nJIPHbi0ZWuvrFaKbOv94rHL2fBTojm4ItfWOfqn2km6Z1a3
S3cQ11sCNNS1LTg+eX79jBwjTQ4HtnzJZgp3UcCgin5r6mw75Ig3lTEKek7XDdzT7BEv/RM5aqOS
F0UL4wH3R4leWM47UqP9XxApzItFqTjz7S4sDX/zssozNX1kheqnJI+T20bxq0shoZQqL3nNFsJm
5kAluAbe49AGBL3JALzK5Ae6BoIGjm2Re22m+DO0P9G+VtfMxDUyHNh1gEWp+Fn8+ikKk/zcAC25
Mb1PsCWO56PcbN2Gd/A+U8ZfAD1oqxko77a0VME9Ie3j6eeBEJYQpwPQ6YBWji7hB2XSwMGbJgNn
lNA0yvG29qKkms/f16leMvd9OCSGxM1HZ8ObmOLfJ/Hosgq1QevBqGZ5nMfk1zbY2Mjby6p/sZfO
ywfLUCdOMaVCydNqjQFTwBTyRuAMfcyUrmfaPksgiq8OuzZ39kylkSuhZzvf+ROU6rSz6wvnVjii
YfVBk13CwJpz5ORWW427AHpVjl4IldEkiLjc6WWGk2FygWXYLRfl9M8+IfCc2scD4YlIZIl9lLse
b7fXzTXtbc6chI/QD+WQDsbbJVhg+/3UdiBNeyp5kwfatPCPRjePPzlAaQPquVb3qV9aH47zXNHO
COOZnu+JLQwpFGkWDzbG6dig+7eBMromQfhxe9rNah0tAaoP5i/MxARF3F4fPKyrl5LZuzngrkcE
bS8OxwEpCLTvrkgQZLpgakkRNgzBiLdehfrujb65s+xbdg4yz4qYu7ht4s3yab0WUaPEOLT7lbjg
rOpPrIoYTGXvwvK1BD4fXKhz4TEAPjtwZ7qVAwYkDcEvSQOXz1ICDTt+wzF4pqi+OT70iqm8Cl/+
s+qyToVSYsrqPGbL46PW2+gNo36pUFVnrNtuXyqEU93+phw2+2g0shwxUZAu0o67fy+CqEVB5X9m
MHgtzr/cdv7V+xsGrvFPxj6b6sNUAUgQcsBTF0jYC7225hbHLDCN20vHXq9dUharmg8r8XugmkS0
deIeubTpsTf0dj1yzwXyB8UjHbvaBCNAIRvkb0C19eZdk/yg9dj3kOvAoFaOWNJui1Vknyk+t0ve
NwAny5S+MuV4toWrKnGtuau5u6OQ5LUki9zRCGlhxnuSeksqfdoCyWk1T89paj88nHuDxa0SrzcT
FtMC1xnnRgTHYkPEZN/m7RbUfM5gvGQ2Vrd2GiH5dnBx/CLc9cT/y873NFTzo5z/DnR18PHOiu1Y
8etyKmPRZiD2gWo26b/c1U90e9y38bqaYhiTf6C5E6VsPk92jO8Ehadk4Z7dS6EX0q8JcT5ZNXli
Gn9v9SIhGLJhZZWfU6sAxdBJWJTv3q9L4L/8AnhAdZJsum44iCPAkGPsCJMAE3t1ZpKQ1Zg2gb2t
zTqW3j9Mv6tOV0SmfTboWE9DQq5K99XJTK4cgQzu6C1CKdZbF/DgfTLz82TdK3RJj+37G0WMCyjz
WBmEYqVAGv2XifAYh2VDrruVhFoGqUYOm+Sa+BvdEHQlJDAyXKCGa2fIB+b4xZWpdB0zaQs+50xK
FdGlQkDGLAccRaJ6Xv6v878LrOReiNOy7L4JYOvRiZXJEbKK91lUSXRFNq6QHvVRgJo1CBywlveh
xnTDApuHdddLHrUs35RLvQjKQ+ihwS7Mj5MnCyzFd8m3jnfMahmqVkAzSpqhbhpioQPf7JYqdt9+
dKP9lRncSJvfW1z8MHY6U8HRrSY9zx8nWnmrDj10doJZ8PUmtGkKGuZvdU1RnP626ISXazvEuhCa
xafnxYfESDFEEneLgx9KBcIpCSS5Nd0HeqH4SUgiO8XBBDl/hD899kKHbcBwbRZCy/gZhQaZjwP1
AN4dBTKmI5hk7ROZ45LdZSH6JZn9/BZkjQHLkNZowmfCdFRHYk3dE34M2OEvQbL1LW06jycq3Jmj
aYkyI38cXvXKDAqno6T4rGRNEw+nMoqhtlODWZZmcCmzryCiswm/T6C5thfjm7iZS5EQaur+SF19
OHLLZ5qLsPN/FpAsKBY7F1jnimMjJ+nIqXM2PBpQp34e7M3Y/v4L2KYek2SVzYqcMfM4uBKN3Yl+
Wao12Au7Fzx4qtZPcuqLRjilZPl4WvKxSALRYaF5PnH3TArLSgU6pnbXBnlL1UpHOvKCsOtUJ9US
PoPkftyQFIbbTa/wZj/GPc8NkT8gbywNTkGMVxe4tmaIBHl5W8LT9IlAjtnwEUL3J5e8YoTrVWu5
7/fAtGtLFFdP4OB/vZDe8PqDPYC8NFhyGuVTWjhrBznbNCKICi5DxeMhP5kgmtrQOmKv7z9L85a6
D8uX0huj+4Gj9qffrE9K9ZWAETUVLlHAwXYhi++D6E/1kMNKuW2tR+pzmMQwozmBiN2yGQuY8p/R
RhnCKtCrzslkOdS8egeP/rpM9AF0hcmcSUMBc5VXbqlsbjtXp1EOMqcinCu8Kl8xEMKebmNx189J
0yvCVP2gEO2bSYzIZcILKEHwz4kAtnBf92d9sNGzugFpBYrmNmyaT4l110wZWFBvvHedIPsyDjtl
+3WLQiU+INtDZZ38tSojxCp2dg3yBQyehFFoWqTuyWQV8+sYdWOQvLJBxbKMb7mCOA3xm8+2uz50
+tA0T6reIRtxHaXf+9hZFr0FY+hmX45wUXxGlV+bmjIVtc1gvu4XtqAsvHKPvBcn9KRnjHK5ICyK
oi+57mV2l5zRfWPzvFvBE9sQV281p/FcUx9n8MfhjYIRBFmW3hgdyoO/6laQobvOLHta02vkRZ5h
mOxgykuMdzMl7OTITf1vOxg9eky2pQwY76AW58Vjxi2gsc4rXLR9NQakecsbV6vejxdHmoYZdwOQ
vPHKob2ZHIMPZ5xCsMYg6qYviqQyCGkyBqw1tFbsXr753coTJtNhHZsPaM9GAP5zHy2GOIdCYpeM
w93PGbwuEWJMhTSXYsplO4sR0Jm0HWK3OcP34gasLL0pfuwCgf37bEek5rdgDQPWTw56i1Cgd/+/
uH95fjGUSmVb9Qiqa+nT5aycRM01/LhpHMCjX53Q7jETf20TPGNq6DmmzeRFIh/EoYweiqfMHbN4
XkKzCdHz+Ytass1xQrp/WOa4Gr9qyidQ65hBDeznfqt5F+Y1uoI+xaVKEz2PR7+mMuaeikJxICEC
kiX9DHCqzf7LwS+rj8fCONlgih3klkT21KRioI6J4g2bzFhLfVntriRF1KgukZqVzo6esS9cezRU
ytoDWL22m4Vc3HEHA5oBAPq8bIbnCZ8KZIyox1T3GGCqHJ0jMac5GU4gwVzOKEXhLm2L+i2nBvbP
UwytsqaVabD6scyPn6YW+2MT50u7H3tYOTDKY0sxJmX/a19f4lfBsjSQdw95Xm0hKe4vGzcc0MQV
cE8LwCy4b+8LP6hPxdV1bzjXRpfdPVW6CgvSX0CutWx1Qh0YQPK/FLB/FOuS3kU6opNzYNCxMh1q
hPDeCM7ReR3Li6OtzrUxb1D29LgpC5TrlIuqqgSyjZtrzU3LQH3vOCh2VYDuEUoG+SfflFo1r/43
cDiHe53aU6OHSVjKuxP/dzRQmb3ZxyxfC7vK6kgMBLabe5s+ZW7rMA3L+wMoqMD11dz6808ml4xv
2CjOSzwU2bn7xhGVPIYBZBSXiUo59mo8+PVJQvCSR1dcJrLtqX01O94FsDgvSnOS0muBQ4lVRAN8
binvY9DKZYXMFThvSVWjxHa9qM32fTzGhk3sKMwPjLVl00tpsU5czEJm1HwrwKrjZBYwjOQFNPZ+
W7yjmfwdy9VeaMxC+G+yhtJ2w898uH0vEamCvmT2DKXAr84L9e3iUDBfEk62qF/45XLTQxTIXkJv
utYwNNJcfjjF04OOONvl2xz7Sf/hSJGWnl+n0l+o/VZOUvVLbp2ZAgCXmcMIcmFmJOtwplY6/5fD
DrXXRoKSQINimwmdMntabr7E3WbN/X0NAZcMftr+c75GLBK7OAM5AtPfdOl+yGvJimHC1N2PcodE
PaDmxcku0jqJ6kH/Wtt1ba09vORhcD2Fah3IgfWH1bmcFotrPVzk+yu3w9hteg1UwPOuJ//FVu29
2v3NdtDxYCEtaknKSMd4eGKkBkVF78o7eg+nwQwsJaav5FWnowZ24Pnwdao8lUo2S653NBXYGkgc
lmq8INA1VlaTg1C1RnEvk2i209o5uA1W5E11L7S+tg1rHX3T338HTNr4upcbGsU6IfMfSsbQeZMJ
uBGgsi/5WMqehrgl7s+8GByG9dz/SfKgvezSqvP6FmVQ6En1gGQUASrsylkRy3AlHNN6O1/thNei
6dpgyCwy3FzTBSuL2LWswI/D+2vO2j1KcBDNg5rG6hDpSPkx78Q/MfDSGW1TY5J7cjXdJbX96rTa
8vg76mcJD7d4a7lU/Iu/mUXMaFcD+LcpZ8Db3eQKNp6z4jIPLMj02sSsQA8w8UyRWBJvgm/vg3Ys
4OM6Tp8FUZFf1FOiibel1NtdJIbY2dmdP0y5+QKVGTKIsMFXw8WuJWAjUotXXtOntsAS1qz3XQfR
X7eUGX63Sz/c8o3Y72yC7ar2MQos6KwHYoee4FRz3pTFbgo/fdYkrPVsvhmRqsfN5uTS+F6qy+Q3
+YkViZdlp0B+FU+NOJA18MYtvQyi1hP4LbJUJFgaPMbx4BawM8IKZ2FsimzhFc6l+ReBpVQJKjOl
Jr1jGJmWvMYO6LMdlYn9fbjZ52/4aedLouGK0ziCJ1s7fql51vzrpMr3v2t6Cw7tzDIPDHGznn6a
X/iSeJMi0pJP7YZkVoTBKUi3ney3RSn6Br7x0/fKoedvGbRHmf0WgB9c8yaFLhJtSBM//WRfAYKk
jsl8aVjqZw8524j8HK9AxZBptsX4HohSqVzPZwMh6OnG1M1xmXTbbxOCCIvEZLF4HJn2NL6hLMF4
awSC+uw1DH0fUj177BowQup91cL5E2UKYMWbSe0D8oi7el8HHXPKldTmw4H6w+K+4yLhSwlfmY9j
hkBJsZ0/J1Qj7hCSX3U/3dKqzQlxE00sdPZX24/VRzeE0bvYw6jW+DS6ojMv0JwUed/IqBFzN0lO
OhQeAEvwHRX7ASWil+rxidHC1DgYd6gFkfe9YqQnGiLa2pr+dB6WPFCN5KmpvcIRO1jA8OMTdsQ0
rTmTiLxpeq6Ct0jvrt//lHtN45+MsadwssBfOvUJg2PRmv1wMKr5BEnR7UD98LbQx+o6+XWP07Cg
F2WomYKfszGi8EcUhr2nUKO6kJI8EbvsaYy9w+u/6MWKwerblAnfOWfEQX/+cbUI98C+icA8yFuR
mUZkWiVyGAEsgxFpNytFe1Kt+EaLHR9QbkSZ2COCrH/1ZxfDlDQbqqvV/DvUCm60yP+g7p/FQGF9
zI1JexZF6nKTj5sRHX8/IMnedl2fKcrMVyCnThiuXuBeGUnLmibZ8NWeXHNQGHh2wjXTvuhd7z+Q
GulTQOQLQ+sxu5Xe1YIXO+gYQTDRvt3NzqTMgF1zYQpSSB2cXLGp0uH/UaP5vihqTvK56lvynqgz
8Tqf/d+gbiRUO0RLCErk/TY8ZmFPVxmVSZIIhaBQbBrNt5Sr2orfyj3xZWzGNg1oI6/+v72J2eUB
addbJyIkqZEJWaZyaudl/XGtK/FfuNsyhlYZ+C9kjLPJKurt1hkE1cqGBDAJFb837/z42KNiLh+Z
VG2UZ9Xng1PERv4cKIedUOy43cjzjLKFmd0otAerH/2e3kadFLMtnNtk3Z/hv2GIwlIHUv8vT7KA
ctAjH61JSn3wMzmqbCnBpWw8ySP5LCjOSkd2dLZ8Rl7216LsDPAOMbn0kbXNUZmn4xo4s88kmuPT
r3c5mDCzwIfpfDMpEm5DgLhNB0lJs3BOdwzjESy/wB3Etfu76kE2RRSTOKf6t5H3sJKGzth296fU
F4lVEX/zo21ZbdfFJkve2NcW2mXV5ZL/ut5DJldyewxJLOAtoBXXNX7cnCc75SuJ2+Bvt0z73GD1
9tIa+48wHPmlOoIdOemwM8esKyQOgnanzXGXuM5NRjKpvaaa/E2+98PwlomRGjSlHGVjYIV80l0x
nSD+CfWJqpEWLtkAO+k73/Dyr4CMfP+i3Tj1MxFopyXHefzXv1X1CIwtmxVgLE6Be2U0J4DckC5y
MM15lk4usjktY68Dodm6HEc9PQRHnFpzv6M2rRvmoB4TRVq410YIDdbw3BeTKX4c6W8LQkZRsYsO
+nyoPPE8idVBotC3tBHfk7YGaFfT3EGp+xtZM+wiCfYKqsUuU3LJcfARt1PREM4KSIl5KoBSuudj
wVXhJKaKSE60+2gyB2xRo/9bv4oAtwG6PBpwU3jwlnZKndl50vsWqBa04Xr0/H5q9Rm9wbmFkQMU
lZiaPtauevE2CmW7D5l2knetB/nqjK/K11Nyrxx++WNyVTsecqNJSVkBVVzY0LUNbbPbM9qc6Ghd
mPjPhCzxyTAlq2iHkYl93qKgpFLCp+9UsIVVTpvWBvKJbrKhBAzTOvcvGjSog5tAsfBexKZkRW/m
gsDRQRWVXP43QtXDCSNOZGuCopD0Ix2d85oHONrMNiviCOert5vWdGKYlC4cRC+5sPRIBEY5h70i
0SWaKsglxqTnURhPkzBN3UHgndY4bvIr5UWfOGIKRHRJymg6Yur3HoQNxVGKESB1ViaFI0QiQosR
FMyvgMZf973EWs9qtFdsVs3TmmLFOmjfoUxUUdxsU/y/qDRTcSsz1sQsvjxK1HO0GnYe98Ox8OKX
kdGhfOFGHTKEoh1ibRuPQQNMnBMQ4NIc1V7Ao4+5zHQDKywOzDk9adzvXdQrusGsI9oNnUJcU18k
bqaU944AvHRjFt4YoDhsvbTbDUajokQi7tRpYv4Pi4IDUGI04pGvEXti2W3OM+NQesqkh0R8PtiL
zJ8q1BeIjxC4UjlFUJBhfucj/FbtehLsVE7wgilKjfHEB+mDlIuvwdsCIc646vM7zGT8Swn+hAS8
QFoFTVnseQRy3+CQ0RXjlGZJsidLkHDYKBQvbIy9S7OcVRo5HjG5AeMBOKC4P1PBC1YcLKFUA6kC
wIK1p1ud8fHGrM74yuxvTUtpObIsmHSXU92bT5obCDAjvqAAxAvVhv8xt26WuB4RNIWnlZFW3BJl
2i05J/EmO4umw91tYw/6a5pzuldwkpQcGBlaFsW4dnVvz8BgHo9Yz1eFjJqd0q78l4ryVDG0BDJr
ko4ISTepphh5l88TbqFCmgF5dxaL3gqS2E558u76+L0pyDzpVPyi+AKAil7VDNk6U457IBtc5dX6
EAQT64TL5bJ6VkAG2MuMbKBbfBmO1yVG+FAFh/zhcumxb0joMMe9C7cHEIUGUQWps2mZcm5P7Toj
MkWNIk8M4cPXMVj66KNZ+erEscZE6DWyssJ8BQnS8cpdSxjjKIfAJRd7ccqhBc5Gl1v+Wx3Db3JY
l17rdH6n4I+Yf7N35m2e28NuBj4in9JEYGxDVWLJATUDikbY5o1BTSNck81G07Mf2tbCth8XnasM
PVcJ1W7Yl7eJGGE+qx2mVvRok6CreCWWMsrbCZirtkEyfvL6A6YYm8ab+N0Rgudb/eKe9/P3wAqG
4CS/z3VBddYsvd0ZDsxxh8rODqWZX3FwW5vLZgmllrhvktdVymL9O5javulWDrAXdk3ucWfJnyAu
MOg01aj936dv4iMRUiRoGpXmk6SQNja1LZowTQQ4cPB+bZUEWeBG0b+4r7KpHwM7W2gnujN8zL7S
ESFrXjhDnuUrDo4q1GDe9DDSoS6euH0KkiFX4cjAf21afC1REE38UglQiRkSUZ7iSJ9FVAd2LGK5
+8VZ+HtK+I+iolAuM8Vp/aQxUE6hPITtmji2mBUCFGymKcPG3Sn1JzqJZPbrDHrASdcGIOmYW+Vt
Pp+0eJr+RurFHZP+lDF+MbH/HAEsnr56DukcZCjD9eimUNCr9//soppDFoYqdh+Xzh+O35TzzWr3
1ch7Y3ncc7u/C0XQCvXqrijvYy72lU9SXPmR9v1XGr1hgxyes7uSLazwT8L2wPAyqLn6EDrEjbgC
45yGWdhyEoM12j13rXZYsbQdtm4Dcd9KES6EKieNx1gl+0nhn5vkFZEgHFtB7odA9WpUHgj0k4B4
9RS36UemEZ/59VD3JDLtv76p9jECu19YlL1IVa26usqfH/HdZbOS5GONAy8NPUImZ6AsE5hZrQZo
lEUN3c+L6qcQftx2FH88Ork3cNH/GcKfUslVn2RGzd4G3mnb5OCj6hshGSPKtoRQMhKG68QLHZ8A
02WlubnTmngtNdOnxp7f6RENSsJRA4sMIrpc10X74VJh/EMhjcIWIBB/tNaDtRtgIy5836OpQzIL
A0jdOirrS1AWmfcvlyR+urUsZzLhXsPbaJFMSQWLZlz5SEiRhDt4XtSRBL/9KFH2CM6NglLxEEWW
+krcj7eGCl8hmTojhilp96CDy80h1PZ0eY9TTuRwV4gZwyuwvtY1ygNOowieXt1No0vRIi09xLKt
/8LxxSeUve6VvomdPnIrMJgWvuarjWsFzZiHpzn+PwjVMMZAmzd8X0I7kWtes0/JowjNSPYrKtAv
sv6nuRlAKzTwoDBE8bJlKLrZBA2tVMhMB7Oy7/JEo4skdkVl6+Axn9079ZL6HgK23zEHNYHWLwzf
7AwvyBUyFnEc4FJobfbfsbJRK3yTCzkyGjVem/piv5nUs/RY+5IRXSJgkR6lHKt6POCh2gdq9+zs
+YnM7+Qf+RGNUUgWJP9exeHHMQRRGlpqtngeJRzSa15Zo9uiMKnLJA+KT/v8apzeXd+wGq2dlTyZ
j4BawMTaCCn4Z0KXNPFQALJVYHznAUbiaIdsBpAAAtL9hD0m/gKUJlSir2SRGNh8SQ4CBbX8sDxR
EwPm3Wat5J1/N+SGaHAI0ss9pPKXJP8Qaufm36igrV6QO6lQXqn78geg0evK30v6dDSwnlULZIhv
sFurZehqjIO4JgStex3e2veH/FtrRnGCyfUbgT98pHkMmA4Oce2gUz4FJcPLbCVabAvi7xodUTcx
ZQg7FudJAEPhOlyzy7FTMJng1Foyvw1Z2XARW8iWcvOhQ40mxhwvieIFLG5SgWucGtH3uSfZV2pB
/wVlnTqbT4PiB5ZzopyucQdb75gxLBOFt/zImb3xNFfXbfNiwb5385siT01EurjassZyvHBarjGY
qS9tbUXm3xRREMaD8E17Nnp5hR3Jtel9a+9Z2ouuLIusLjpXWa+oqNPLxzCg9qLMbK6V1wtj10Ph
OfPPNZg/SZHUBWJJAkMBMG9cBBmtyVW6OKyvC2ukboS3yjgN60/5hqGS+4OC1WUhFSkvz0sVQnPp
5JQSMFNTLwmmtXTbyKKzulHLiDb2AQPb7W0rmxPFOaYjDvdJ8mtRzy4GaFNyE2eeioB6AIAg/q02
ld2U1dZ4SGID3XNaEyZubEJzogomPFysSflGFG3DoQ/KVGIrUwmG6cauzndbJeDsSca5pRlaPfx/
oagh03A5D6CyXDdQ+GuIbd5tFngdpD89FUn/luzfWVJoKCTprO33eRhoBQUPBo+P2cvdsQ2oBfHv
r+55lwIwqu6k2K9BuXLZSRJBAoAP2Po6rmpA4tG2ttuLdLFdzeUhUOVDAgqp37SRGZCA3zZHnlHe
+XgPBwScLGFsci5ZdXJTkvgKE4NaIEP/MUt/8EaT0JwjpSdr8esejQ4+/mUhh5KNSq2QjcLESDGx
daKhl45NiGIHJlDjE3fZ6bYjFisbIxXSzBEf7/v+93SY4xSGprMo2zb5IStzn+Ku0yHsklDbe0h/
1ItfEI9GM6bmVxX7ILwJ41jqA7wNhEBPENl844+uO0t2g2CBW/wwv8g7uHQIWW3c053E6R7B9OZn
+o7tT6hJXGaJ+txQflMUgMlkcBcZQKZV/kHpg/5wCmSkL2i3dSgfXoK/PwEhUnOeHYGZSi/VORI4
se6JajEplEYp4QoCJUsNAWK3WmJXFPHLhs6Fmc4r9a/mTHB7Up490X+ZjrGZjie4y0pjDbvDajHT
0VHI2fxLh6mOuT5kXZHA+gElUHCVcolTv872vMQhWhE2hOHk1n5F2pYnBAcCr0OMl3JnFoV0FEJ1
htJJos/5sbjejY759PTLYI1AVSjGXPIu3G/SOS4ytEawazFaYOpH17CvaHrItN2bJsHkRNv+GgCD
4lc/dIjJ6vN4kGxj3n40ImeQUlfKFn/d9ieyResJNSBdrAevn5/DFgAqNkjzDdIAzhCWvB9qIOix
EvvWrfvB+HD/l4IvhpTvVtoIsTNzzecayErM3+znDcg+vzhBXnBAZSirf12A+nicML9fmd/kFB9c
HUpUfs7rB+ZompF7URdKhVGacQUdkvM9HwBECbV/TIoeDe5cEgT8a8mh1VBaw/5GL/gksJt+DWQZ
Irs/j3btIOgIbx8lArgAV2PJy/jNZ9S2P/7D8lzx9zatJb6qZawtwIlVfWX5PLUjhX9XDtk9OWsO
2ot72+csoq022aUH5O9TV9sgh+GyD1i3XHQPN1cBvzSSmLAU7GqvsYTYpLhWbVu+GQMCFDEcPWiy
vPhVclVKPcTvmjE41zum6AizWLIVBri2UugjH6f+wX05YMsv6nEUhIk77GbO8PbIlp/DIwnmeVlR
eglnk8e7lqKcvtYaLQCdSeulo9riAJ5FeMDQdFLBN+c4It1oanBN2mkPhiQEbqzrGBhdy80u3piW
ZaK4/pdthm8Wa27FT2qkq3v6QNor9A1/drKvV1LZMg5DxRD0Nz8Vv1nKrqlcl728ZqWOamv0LD7h
uXyYvtkF/AhpzbEzAnQiir8XaoR72lvcQYmD08l+u/CBtdHt9nDLdO4kK6fddanIMf6og2Qd627/
Tbm2M93Ppv2J9LjaWNMAuFhq3U0fhymvVAiXP8W1l7kWaWBjhljbZLF91jrycMYV7RPcBpQ3Cy0f
EXIHf+tIHoaArwS0XaeuKQ5GDYueFDPmH3X6Wr7UDQcnqjZ1Zd6wlBBSCxPEE6d9vgfOYn4Imm90
61RmusiLX70xGiSRMUmrwdBEgEIcRhlBN4dcuA3oChQITBKZWr9AkUQVGZNDNrIPo1AXwmpgrLtk
A4LQty08tPqt4Cx6NHuc0GbsQcC9fB1bTxY96SF/mSkyRyfZCKvgQOdKmX0BnI+zG778eCbDot7u
CvVd8mdZ+BvBQwLkCZM6BOlu9hXEWua2k+wB9sAzA4TgG+YempXB0bsJAJ8NrhFb25opO0RHfPvp
h3xGD14BxOwPY3amrHWrsr3fGjjcfsKJOEiSiU2eXHHTbwvCo4LzOrOdoK0IbIVVTZj4mrmk9heI
zrWa99+HrSr1GTEzAZVwnzRzXgTme47bpC3RIkZCivg9wbu7c9Rpd1uFH23LphcSZeNSuso4TMEj
zH/bg3Fq63CJq4DAMsf4qpOiPFxfj75xlYS1wwxa81SdlBEuNf35Rb/7VecgwjY9Z53e+jtyOe9m
4MW4DqQVYX+gFTLVBh6ppZ+uXprBLGCf8Y2cHiKLX6OtAN/dMqUQschhovuaRJM5BxLrcRpf4cgx
W1Mp+EUwDM733jLPGWp9v4d9NcL+2vEOXCzHRM+VlqFzVEXwu2eKexlzCDblW3VCwu5FRT51/Mz6
oPQMdS9AnzbT8WPNDz3qWq2307FEKPd6uC0VxOlJoQ14/A7/jaONfCKogRXcKZB594eVIlUlr818
wvym+TEUb1/2DyZsjZE0wU+Q3AsRUlV/CG2j4XzvP7h+Ew5e/WIMPgERP2bYx+/Rl0yGdCQEuUvD
Mie3cjMEC23T3omt1wNcInOEnF2dOsrKHV+j9Bv5Mgz7TQVpipAnLbiElGroEdr0yAMmMOXVEsCM
U3N4k4V6YhJEsk7eaimxXQh79x1MRmqUhbL9MFqyb3SLO94KCL5a1wojll2I/BEozFFV5SjrlI4R
uBvMFfC9yLM63sPCNNZRx9rMNJy9g5rNkqjZwvEAFvZyWOiyOiyvjYv5O63vjI3olFek9fv4LP6S
82+sQa7J8Vjxj2fwww686BjXXf30w94sgw/HAcas4cFKm8uMNq8Sg1lzi/+0PZXebVQaJc4RBVMp
/pCeVfSnLGKDpSkH+/vjCyLNzvcjRWqGILPdjPUIXC+efa4TahrYPpYmn8tU/Dw/LO10y0eqJauV
1Jxy4ofipwtYGrVkD70wWXppEzQf2UCdd0lhTghTnPzIP6eSH/Zzc+WVp9azeJ+2do6XgHVPsyoA
Ota28686i5iU0NcgnkubuJtvroED4QTDYpySHGI6+n9axB6nEiV3IzUI6BdM3/hhalpGp4qU6CcP
a18ywW1RURgGyVfeYofBIyE8Tj1cQOlknB7I+IxdLpjKLPTCHhAG2L2wf1rolLOUAIzpfC4RrLot
v1s6JRhRZKren46gP3cbKC9BIEvUYeMEgNilSs6fCF5L5hBOi+cV2wXy9oYfcs/Tt9Zt98NS02uR
JIefNsXa6Iig0bVHGy4RX3la2lTn5/LDUy7ML40ai+TYN0oHPH0UiUzZa6gwrV6jPvZEc97SmmLa
K9BdyWHF1IqVrypp8lKyV/wU8UyFkWwI0ARN6W+0w+YQq04iaUj7zqEtmJWvkXZY3iyys87C0vUx
nwEAJdnCI+OzXVWGJ3ujP9D3UEwLU1wpiKqsgsxxNPgiw/9PNzNLno/8LMpDt4qONm1xokNJze9U
R8oP3tTCR8KEr7JnceBC/vxyZTmoAdvslpR9Pt925sk37QFauWthcSt9tLqcQ/N8HD0Wq0tWvTa3
BY6AAUekcNX18wkNhHRHcmNk2NaM0+XAO580L+Wg5r4eqndc+qySByb5VbRaD1QS7hxAIwwx1AMU
C2313nnzL3xc8HlDDXbMpqEazYoBxB5ffAfGlYdEuXiTXfwy+DyIXXlbpDgbRaXTbWwLbOL+hIT+
3G74ADafF7lqTKrT05mlK5t4iPUbqTbvbrJph0Uwx7uqfnmsXae2enbdq4+A+ehM67gDhPlI1HjT
LRfsoM49sKTEtPmpLxcgyZLVhkXSI+H/eh4BZn8uv9Im2ztXVai1DBpzQDBYahfp3eJWHqDdFJbU
TgWehJqiFpBPmthEHkgiSEGKEjBCQtbjHF9/xyfKB/JnePlD8XOFjA5ig4yOJaPSuU0KvZcno3G9
oD4z014TV+SBRZVKfUe2w/aSCsCALu5QXzAsX+XDjSqcOfogi8WFVKuowdF+PC3YFAk2Og2jYeKv
JfTHhg7EbuXRxnfx7kZz0VWMPLf/nuygLHfSNL3ooNKviCPPNNj3BbLZMY6vADec9qI318FB7ljq
CSnsRbe0QwzhK0I1e7UMZSE17wiO+DAcS0rFErtfyVdLUqqPWJWqAK0DZguc77cBE6hKOmg9CENL
8tg6QPLVNxcOyTMcWLyLB8+828nEAwMo71DxIviPUJ/aHDBJEpi6MJi2Lq/w3LAws9xChARMDTE4
DiSj5kbDtr8JA5jKF+QKMkGc5GKFd+IUvTM/HsiQmiB1Tkzf9nhQeF9Ya3QT42wgWzweVWG3XCQQ
EvAZykPa9DEGjnr/itiKUFjsElIw5a2mB5OnGM3xphguM/Pv31PEWeiTZnrzAVAHnB7ZL+rb4xBi
KSQtc7h6FDTqq5lEWSTmeS3ZZdKuxjqQnIGGykSsmlVOEa0CVTtWCPZ6qUNKn9CQwzEApavw2f6g
MgL/Nc/ScDsCrM7BluwyIiXQZfYvldmk5MbzaRlz3JP5seKcYczLj2B8Oz7JEJ94jD+8W7tOjvNM
INBnvHPsUZ7pVv9LqCY91G7mpdmg4YGrQt1+n07T90kb2CVtym/g7upze8O/6YCrB/rPjKkzodDq
Ielq2QwCoREWNK5WmaciFC5GwyEaw8nPY9emT/jWXIoX3Xfd142A27LDsxpkVUGdoXUwd1cjXmpE
p+hZkctzCbW77LQV9ITv33Z/Z8zNUYAai1G1CXQ6z2Rwmb/Y36/rv1l7PDO8u16dWKmBvXD2rHAx
j6O1LuFnXpWoWZbTIIqyqCGAdcH7OPAbHA1YKxTQ1FPHLCkKSSr2+luO6VARVl4Og2GWG9Pt9RE+
2QAgfSYKzV0OlrISzGGdG9AiOzfdm5oScsD0MNkXqVateUCpzb29hIdlwZ8Sgx5ld3C+ZA0RbWlt
IrV0meaZPl3N11eSAOTjVLNJJGZONTCpFLPIxf/tUkxIcMR0HdQZq6peeqN8ykJav2NKu4FZJOIC
ok2+u35oHCyVTxVa3i7tGNDVmaryppbZfc9Rxprps2jAuUfpzRH/FBdbw1vLHBdgDKu9TTO/Ttxi
ppAeaniPNSAybF5nxlZoX+Y6iwO1OiEapDxCiBQjAWfW2Fw54/HYskJyniLChoipIWYe2RWzD6lV
6Q7VhPO35SP+AWKbwlH2bWBE6+scO3OCFQ2FkyUpdkm3dQ53InlPrIXHKmTFy1H7I0h8aLEYe/33
QRhkoX2paKWNX8k1YLYE1NmUfp+i9Giqh1xAxqGM6LD8KoZMdwUzQK+XPzRp+bM8B91R9xB/qpS6
QGkxtY+qw0nC0RXBlSk5Nnl7mMb+nwudkm/iSRtdnMI7NrVWVnsRVUE8AgsQPmAvYs4dR5eerJ7G
8+FLv4reT+ejWKofaj6DO0bCFDNScc4ddhFNlfOmx2JNadUgqZU8Z0vygPvPpNspIpxvmnwEQvCe
ioBYcQ14Snrm6IUBjN9ZavXU5L0/roBZksa+UaryFbUnH1XMhGQrOL2ej3jr5DtqltI4RZgglDOv
9mqrsB3A6heMuerULkvuLVJaXq7+GuFFi96t+uNblwXaWJb/4iOZNn5zCZ7vlEiyOltKQGN7x59N
PreoDXYScr0VJIh9Ix1M3Riv94Ru7h51tj44YJkDiJD6PFvKXcTalGyUCwTXTqQzWwjv7zunBdGv
Onl0yPp79/cp1mszS4lrqVLHZfwIPQinrMcEhtXDhqXzhZqWXAhC5TnH0bTRGNfozUt9at8QxnBU
sLDnDLALWjMiDKaLKWkA8rsGTPzh7X5TE2iG/2KodNdxWni0NRqr4ztNZnvLIVEQEIg0d6hMefPh
lyrsTt7xeFEXEXSAnVtO3L5Y2+fqiGoJQ/J8URRuegTtSgJjHHZIdetBYniULFPYxNDQT9wUtsLw
lFPjgWG2psgCPKDBZXL3A+ooMCuFDqX2C6/RHiiv5hC/J1j6utFA5eIjTrUfyN+aaOhNJAG87UCw
m9u4n6X7hPM2NB8lGcSMRnjfusNAzSppFlhkcAZb+MD1zI+MTyLceswMEnf30/OZFFLTSeEoQFOw
GH8gsJr73Vnp0tYMMzx3svXUwIgopp9L/kYnnYpHvNCXMrgRnSUUlP4AQDdXPTXWrrNAVNb73C7S
NvwKs2dEjHfsFcQ+0DrvaY02htLuHJXJZwYT9wfMSTT6cVp4vi1aSwRC/Fj7y/ecz9PMvFS+lhsx
7SKTyeviPaf923f0mmBAcSujcZLEjqbjCMSbl7aCDv4fCSmARCHfR4e2L0ewELgepb34gePONr91
mQJP7nN+3cIS/OXljXGXZfZjVb0usb0AsLYPPEkWfe2hpyCgh467ERTh48yExcA/OzcoCSPheNmc
vnH5soVEXOtKQEqid8fCdN7WgxUMwHvnnGrXmRTWDr5MMWY/fvp1VFhiENpLHBDEsw+E6Y+mVk8n
icuxJeXElqFLpQaGQGGFD/O14NR9v7iH83J+yuTNswGDJRLZgPGJ3IWeSJfRPNa/g019ULqRx8GI
d8HzBw9OLIReSCwXnQfyzRSTH3ENgQzUtauh1RBgggBwAU0I2PCLKwygnEGxyKuk4U4PfY3tTghj
3rbsi8zY9Jo2IuAi2xfbVAQR3NZHcggjml6+HrUd6/zrDZUvd7AWVIc81Agh8KZJzDUtDur1E/Zz
E6Eca8NVAJ06KGDdB0ke+/S3aTl8HTeW13h81b1+er1b4ewNvArZ+rkCnn2pRZtwgc2Q/UuatMei
pzZwom2FQzJZFh3RunY8qM7tb4mnJfyJA375X1rhjykzUALob9zIbRyoXHtnQtCSlqlxqP27NCai
7ahrNIX8kYwjSUG/HBqRRperItNayQqkZPk2QlY8EJPMO9amFe/wFvZHArWj5EvCtYb+bkWOKzas
MO5ba4AhcNtTSdIoN9+cC2fqiDztyWXvhCAHXacJJjwDL/ITS9UnXcVzrkx6B8W5MijLy8+2mxZV
Wh3pqBc1Azvmcm2O50iBQq3e35ddpSCcA5B/kKj9f9uPsBAXP1/szANCCmuJ7WsJxMqwY9ol+sUg
EAT+cfCmCFUYsh1Yr3iuSmueHW0sexws+EaTXSDWfZ1TOEVnUy2oIAX7CFLv5YcXsH6KDV5k4eQk
waM85Vxs7C40jpM8YhjjlFE0sBvJE/gNrTsc4wAqrfUIbpwonwSE+SuEYOKEjnDxtlJ8wDPRnqu1
AfBP91LwpA5c1A1ldg4A+st1zBX1VVcwgGBVpuBm6PVTLeQG4DRn07RHiExXO7hy7ejLnQEkW4Mh
mos+c40uVeDyST3PuiA/4pIP4REooEJCh8+9z0t3MaZv01jCiI8uihCuxH1kMhIuSIMogtNxkwvZ
Pch/nQANLVY8KnkbLE3QupG/c0nozzKEfxuEIxGoqru9mMms1KNazdBSqTLNNeR/S3D4afFqHgbN
kzJqLO8h/aFMjF+OHS4d/NwhehQqQApy+0Hj3Zp4JhvqpCUQjdsbN2JsZ9Tm5v3jxHtLUnqERkcj
yRzK8sZf5PKLvDzIRY+aRsbDPVFJTaJxK3sdUPewLZiM1Z9Rg5E4LcShDe3mhgY8v6k6Z9/HTXJI
Gc/QfGRsq78nSDEIaUgFBdodSeoXm7cT3jOhClCAJDg6m/RML6YMskGP1LlJD7rsH2wsJJSsnTiy
BScPvvqXVeNI0GvGftPs8N2diil8fuQxqOT5oMX0TMgbwPyNAmdsjIrRMNXyZoYaY+vpqdmceAnS
GNJB9ZEBo2oTliIfmNsRTQqmkQDRGlCrKlGrnyvtw+Fj2lrWRhE1qgaptpOhjRAcFrrLG8uEvsUi
GD5aE2C5hrS0lMg96nt3PKDk4cfZkzb0UPluAmD+eBCjZA3SgenWWfdUrN2koTqCFy18T8UVTZnf
Do+PPiZVt8zceLI4wL9OAcLAApg9avwZCFGM3H7s7D/OD8VcrtlhOGh1/pd+i91EHXSrdM46rl9P
qeSYY+3fde9ujeWZOSgHOOsi6smEAOevYyABbq9CuTHdAaCrHrUFXcRkg0J0O/qYV2Th5T3p6wy0
NaQVhWrpVpG9Br564v3LgtDITx2FgRCz1oX4IwqskkJlp6mZQUfhPOiZSgh0B9kikBra5ujLSdS+
1yklZaCfVsXLvwzdV7J+XEG3fi8Wz0sPq0eGDRzT+NfzwurpJe2fOZVSwDmTuu9ih2hWyosDKLPi
gqjKBwnnZiXOj6YCAaJFhGzrL3m8laaObMzB9ftv/jJ7DddJ3uxeshSAtTmJlCKok2Cm9gqJA4Vw
shCmWAwqiTsYIZtclPfkiqp4gSZjY2BuZ8jsSuIN5sC4OCcClRqmyK3Hqbp+a/+oOudLkL/FEWgS
9aKoTjZXxi+BCh5dmwecwjpLozx27NuxZwulxNVrAwjmrCILn+ls36GSbqqRJkYUvVG1nZ0F7hFW
X8qVSBcFRNPgb9SXndJJN4aMSpovJriMyVw32fA84y5yTBu36ptegqZnTuU0NZJi74htX6R6GfCz
YZ/c68dhMnBQbEIyBDX5dXLB7QO7EalamYCT4b59uv91BuDUytz3uh/dJU2WQ+DVqaSCuDEdsyh5
+C7iBjlRNfuhAp+amfpy+qNtiRIBTnWDY4cDC37fqBojq+carE4FSJJ/cW9ykduAYNNWLHoipJPX
P3ZAO+9gMBvQn43wopLTXOvTdHYDRMV+BFqFB/6sWcsCgFeeLJtXc5oYCT50UNHwLJallDY5m4dc
Ts1/Tp3aC/D1jpWE+csN8HuEaXJwOSmDKflo61h3mbVbKl4Xv4DvYEz6xf8Lx6mrUwBpu4iWkGt+
OMmer1dMJpRFtROYO3CBUhZjEeWFVankdbcCTSoecRBeONDtrVsi4LnXQtDlAa23kWqIf6E0uMBS
uoimP+mvMy9HBwX0JbR9EviY3XFwPpN4/MaN07LibqzBBx1pMHKzHyDwuQwg1EXdbvh/CSBm8XUM
IHUqBDkFV6Q4BJiOCcbAbov6lB2D00e4K0pj+EFF646nigr7IW4ebSSDzCF2twdVbsWeQKJ6tv2s
mSKGRHB5uL/4GHhPEszxtg4rVpIm9KFF9GE50JUxmES9RkpdqAuQExASbHE9JV+p6rqmpwRykrSC
BJB4HdoWFJBKGVvMrZFmGudm+NdWzDaTMltx5UhBBIYacsI7KnaMybILUUW6hfXc8bFsozyDaQKn
QkQEWyTivoHkrOrT1GKq8xu5NgKMRy8dqeA6pZ7XVLhC4VsaG/bTcKjYTRVogcbg+2ip+7oyA41f
4KfTUlWTBoSNNCp8gvMp6dUtQ6Ucxz8HdZ0XPGANpYq1CDep6zOfibRYoSjmvgSnwBGLwrDqPD+D
5Mc1/d2qVqGuqdm/6BXoRmf5Boa7zAELkQqQDmWBu+vbisKIHGdshOipYRGMBHSKy5OOjHIOUdLF
Tbd5XsgP+ugV8DORyABKrrtlV1nCLm4K/jR/01qwtdptbEixnPS7/G30wu6jsPIaYxTy6LFd48u9
uKNJQdPf9isfYkaekiVvCpFv6qn25EZImBbhBQP4aMzjLzqMW/RYg3rS7JCtP+Tp8gEYxAyKcp8s
41//1ERD2Q5CTbJpBROXkSLJz166fRuTv1yvpWjNr+uJlL0/3Oe5Ov98qViCqwdh0ZaIVgyb+tQs
/k6toCF4XwXrxstoutixpBT4F9kzx6aUNFChg3we7B8yX6q3MpSXjnmdNOAAhyf4bs2KSfT9sLlE
/IJgcWJnt5SmzN0bwUDbIVeOkG4YPOIsifa8+mcN8qGdFMmKqOZmQkYhkRhhEgkniBiZS8V2zyug
9MzpeT7bkI/TlHu/GKF5xzR/yF4qGrx71Iow2Vrl89bCM8DDs463CM6rYKdRj6S/Sw8d30gObBs3
qONygdGpE8i0YwUcH5XBOaupAsniulUgwCNCXeBrPLrszuKpYhWvHwMyvraQWEe4/QDhici0juoN
e7ElQSMB4iKb/oR2wrmJdMOwQ+k6U60FgOU0IKhXCbYOdFwKQQJp4yKtwM6jaoWIUPnzrNb9ecyt
43RkxK3WYmKDcWaUZie98eX1AgVDcPsXCfc+uSKKrodz3mOZ6eF+buoMtUCihlvDEHZ98xOZxxxo
JCV65irMqlrZoIuca2mAYt6vkG6AN5D+mt8U5Noosf1AQHwuAJYaAtBRK270q5iWMH/JGWlQ+w/U
BXGblGI/1CjNx2MY746OPKgLZwHMgb8QTlM9bUyS/HUVcREziJzbWgNjCk5qVA+WNfxLhqmA9nGn
BXlWyWtLvoKOk2DPS0+jjwGkSXBbktWB4TFsYNCTrm+c7e9Cpx6WexiIppGgwtQez1tJ9Q1l5yno
6geKa9duJZHccUEpHLNiU5a8BOIZC8PraLWiKTWk4zdns4H0dGNg7ye+ciIKHkGHTFZS5i9joHK/
uomX60RkUpSZ+qQKLa7HGVSfGh+XmSwYisvHJ5aUEIBSAVzgpPdkcgaQHegEb3IC/gLmEe8uwgTI
VdikD3Caaki42BjHhP1CCe4ya7+mMggdbBx2nQkwNlzH99RDTIk2imLvwgGdF0xyp1WAUrun+VMm
y6CxE0Pik7HKt467fFaovE9G+2R9re5mkiQNVlkF3GvPNiWXoNZ97WQAbhk/Et2fS6wbkZSXvpe8
t34LP2/AKrXeDQ8GmZiKFbs4YErX9//FKKDY2zZmMU94Ts0OdHARBHAU9PBi2XK504II2EZ5BMfT
ZV+5Nh8voQygPWV9vKE1ZBoYfNg6PFRXEa0DhOy4vfB6Vu9CVk8btzm2nNR58M0Cs04QqZWsyc8g
BMIuw/QWn4ao0jrJREk8bBN1ZRqbncsXLxZ4jyZW1G9N8wxPPY87FbgYk0ImCqkSNy3nl5OiW/lh
yBiSKQe8FiHvE4GJKTWeulSD8e2A0Hi/l86PCPDtAs9+67PiJSKoAgN70F1/OUorI9xcJxsCHRfC
w7bnczc0/8p65FH5r6rdUBKREtOQ4Yv65jS1EnZ14YFf2ecIVTybmbOgYmorDtoggA0lNxEG4WhZ
ktv75zSSskAgEquwb/8L+tfY7TaAwFYvQu/dfdEKZsSm+4UYql1297rywdUghokXNL7hue2NR1bw
wVQDvTzAWb6B1mAiOs2FDnXgnEVY/m4gW0VwvRjRTxMZc+BUY10NTqm9SsxFIR9Q5EAHnW6SJvdc
NHW0YN9TGPySUZVmG1FQxs5wBnbV+5PYnr6XNiCXpuErjvzW3j+9NeWygRbsj+/+q2B08dlCC34X
DzC418KsxGu7nxrwdO5BQyJOahK8pfQq5HYSEeSLLckqsIi+gGbniENCUy7EYmtfNr3iRGNuECFq
9Sgm1o1w2JnFQ8rmfNuIzcevuwvm1ZlIZxUEJO7m0EjVtBkvUW8/2X4ft7DLUEWy1JnxX9Equ9l2
PxLf2/ewZLMCgdsUTRwR8ci5HH9EdQ/bYqkt++7Rfw38161ufh9zgqts61ykw181SXRJj4/IijJz
lCW7FYUXgjVDBFpUxvUL7+V5P/VAlwMTaZaeMqpYYa3UG54zWC+pmGchi+d/DeqsaUOkb7UPUOOz
g7BXWT5K0+XB516657gSHH8PVI9VvGT02/LsS0M7ZC2oBJumwIGUiMoToET2CsYvx8cdSzlf7IOH
LqQhT641irFdAInn8K2taH98ERloqh6gIOajpLk3iKuJjqSVBwTRhppoXDs0/Wgh9W1yjOJNND/X
LDnjAFubu/30Ok2+dBMDLvvo5cXXFY9dSAbC0dMA9xj+66XnWN/Ygqmj/1WAtF9u1AtNIUIxxLbp
NFH9Zp9v2Ti/PfvysBrYRH+/u/oPQ/IfuXOgNqMMxP8WX+u1ly5eCN5omw8BkGNQpljpWoAk1I5m
ME2ahPT0Qg1OiNNSuAFUTB1KCuOaPDb3oY1Vd2Cfm7Ot5pOOC/u6Tdzk0vjyG/URdNtA0FS8kgRo
8L5PJXlWAlGoCQKUm4eLQRlJAs+HAhet7wIouRlWHf2xhUwcUVB1gOMR9PNzAguZkgR/bTjmz8mE
xkAa1KeQqtskaJh2q5o4Wxs5rBKymyCPb8HewVkGgJiwhysUi7qrN2V5B3tkH/xLHopMwDxd1ddj
IX2q/+A6Of/oIUVmctqH2yhgaosLrYMCd1JhLEItmvXHOxddMG0ieyhOMsjWCHt7D2JmzaRloZm4
wXk2nzsq9jZQDclBHfNHYi9WM4xpVjd3MzZvcMDeEEqeYaZBzFgZC52ONOrMc0Z3O+ELhzax0aZE
4nh3ncA/i9IKglABgTGkp/hBHCUVG2oiEH4aqfiCXunJOwz+734bXicaJtFlPvqFBMHiAV9c5Xq1
46gLFsKUxI9NDtgrKIzmnYz2j/kR8ayp0lRaDLVKdziWNuZ/S8NT6ZvlmbDacbGmSTvAseXkqbzI
bZkttpUM9kWhxm7AM3OTgPWBH5A2HuakaNrMHcUw+gbKk82cGTEVP58DaD0PDO4IiKD8PW2NopRI
SJIHxprCD9V4qT7nayrWe/wx/TzSUoWMqVp8Fh8xWGpjO8Wcbiw5stkIGwLU4uDyAZCLYVlkdgF7
8Ae+Ag8jF2Ly5cSXA/9A46CY9qNE6W8iC1dkl7Z9uzYw8x5oxd2q9lpJVzjgjTLJ6d93yweugmBJ
q7JFDFEREoCGgIK4oBrH3RF0iDwVabJEI0F3XLW7SmOyUD86cfibySE9qT6yC0Dt62t67aWBad2U
j8wTuUmMC47h1eE3F1P844j0sBYhT1Ij+abnphjQuoD9JKjKBn4d1DCHejDp7h7jFfu+35jCRefP
RbxXPov2YtRudKOiBCV+eR6KwmIfwY3wtOrXPB7AklY8t23e8hiynZL/+OoytUL0Yve3qZzqqYqO
tSxM/3fUa35L1BfNS61DhTXk9PKTdjCcn9FAF+zWrhHcB7x6JBvYDksFe37fWX9/U7VcbJZmlVKu
3qQb1v1YsyQdQ8zzP0PPAQTLHFw4zWjgC84yiiAmA7FW7pI83Hyveukdit8CABiMP4l+JNYU6n3N
T3V1vvuhZ+iHTh4VM+bE+qzqNdeLTSzeY2a2fwtM2Y3E4thW9Xbjz1jIcPDetKUS7lXP/55gj5DK
QFFY2NMw3xvUDcpqvObtlOZB78XqRRD0N7jmMCsd39qIMvz2iAK6+KxSoDRtoi+iALGVUjquWe4a
dDEi5o5czP0Wh31OO3NNcLGyZ84Fy3PE2aIfR6ZLxfAgYjaFH+30o+OWYRiviu5MgR8lc+SETvWm
3jyMvfLQU8fYrZ7QYv4WDxiX5do99A9EldnuJqou85bTKb+BxmhPF1mvtMWT+2rHDFq0s0z5iByZ
qCYheUhTyF9xcAfwnR9ADESXiWmfColV79DHF8QiRvHyMQN/LBZVhv7bcEKkIM8Lq3Bu7lNPVhDR
2/bfAa2Ebrs2xX4diZ1zMP+G5gtNjU/Neaxb9mwKAkqjT5Cvk1mbOtX6IXUuvQ1egUIvb2vo8t6v
m2tdJBC62ZXq2h0YdHuBqxIbESM8jos4hOZO/RbaeyPP0btvTTdeqUi4afNW6otqy2Hg0Z3iBy+n
FoFwD6s/apcwNQ3Pd9Sx3vvnghHG9ovUNoU69Xa4agyjnxxkUXQAKdXWL3eOhmguyI1xgaE2yl/t
y5Xh3m8ga6tF+9Zomp/efZCbeFs3pG0tTsUBQHc96DT7gCr/WrzTHE8XKTFmBwuQuovGa2J404vB
BJdFWprJr+80owmkxMPaIrzJSvCvJWgKTnIE9mbNCI+YadXsAjMswykoBFE3j4Eop9hqgVEcOZR7
uhKvXJfzlysrm0FSJagApqzJPjZwiS4wJjmQvnot9h8Kl9XRZAqc/HEi2s4h0AV3Y/JqxLw7WQTb
oVOte5JCkiJ4Zo8e5vhntjoH5o7RdOh0y4HD8J9bQxC2GhT6MVYv6pkPXwS4IPHptJAEJqY+rwN2
s/vdJ8E2RQn1F3hhXp20iWir8gmIYiwQxNcK70WFGJpn1Tp0JZbKArP1LXXxCzXkUyLeHRT/ELUA
ZpJECwYciRLiTwDRS/MJrqaGApu8rLuWA7XOqGgA0F9mtIixOwEce/L/vv9C2t66jYR5mp1n+JVS
ME2vDPrhqQ6TtZv0DK5giGdT4lXtR5EEFl5D2ojiZCTIwK8SFnnpyvhrNsmiNtGXcYtpgnOW1H31
Q8sSNsPt/hq19C4nq26+vQTgv0uTHMulw3GSYCWjVCgKAMz29P9Dz7jGrPtgmJ2aLNNqE6Izsh4v
cvZY1nsiKX5pxycDeGPIQC5lxqbAvDR4v5Ubd62FFJMP3i4brh/2eHZQOKwZ+U8yV2b1L8JRl/3B
gsH+Ij1JHJyLl/NuYDPNFIThvIhK88NtUbkXLFlm/JL8VDvAYnvlEi4CCN/D1OMkhn5YYoGK+rcW
m5kKyczkSGSp/pvhZFnQGa3yL2OCpMfnvf/DjYBtMeWSurYU09rg4GhScq/MrJjaWjUixMWli+on
ALcz4zibGqjf2Wb4J45SK71IDl2B0+v4JyAXgErA7Yu8oGpcdu4tDfnf5K6pGIJv41nu1XOyDmWz
TYbU0jf+M7Yc6duT4X9NJuuxrMHXSPJVJ70TS/zxzd2h8rOLWMPw82hwbfoWBrnZpwKDH8G6kShK
oRuTGSe879Gp+BhDTqLreIultjF27KgkWo09MohjjZtEIFL9SMV4bDZ0Q9ruGOAttwQqxLV6ilQM
n2uBthtKG39bssSafTMCYt+Hq59K0HwtZBTMNItmKrpsQ8DjHBVRrGh1gWLES668JyF1XsIcOXX/
h4QTCb8zsn5Qy4JDIdr9YBoOz524c+DLxiAjNkddaOYVmOp5MYv6IBadrW+w4j7CXo0IH/DO7g6J
dEiEgECIotdjPjur0BoyN+vy5MtUEgJ3SWzEI4dWarsBf8aMktZoY4IvaNxzGrqGJlg3DnHmPBOD
5tAdBc7Z1O6nNuBvx1EaRh8IE5vvQqOUXzOI/ANt5pXH2mIm1Ludxc8Wkv5MacZW95vGakBPHvc5
Awhiyot0KyJgyrwPNOME/juK2Be+OTvQ2cWx2SQ/6xe6Uer/7tkrnJOFS81QPixtNsW7ZVZyiYc0
cP+wF0yECHa4ImdrQBrPCD33EhBK+mvr7kmi+9AxozaEfJHQj/I1XVjoCtH0YYXAfqKlpzBOgjjW
bBHA1lezcRM9/c9hUbROmMWLt8xUNeWoEz330uX3a8hCHCIaiLiroKbBFshkUP2FMapnBl93LlDf
fVslnlSOUR1DsMbuMlhEekKkVM2B7IC6erVEN5NKwXiSnaIFxyLmOuMlgvLe3NvizXMNqWcIV3rQ
b3d2c07nWv5xLtFDvJxck5aLIdqqpSz+GNAyNLnvfkwKl+gMW6IKEsxusFEZnv+SZGlFzF9ysFgm
Ln33apkxhMRnFg/V0n3V1xX9xOSgF1TUWj6gvlQrWEfAUDlhahBcfCTwytNUaaDddBASiuKulWyZ
hZNURiBh8b9OVgyJrF4gmrPRC2HqiJSb8ODGYTyCuJLKaMatk+TrkVPdmUCpkUrr3bxY3LXTAY5S
bwkuoepmy6mBnwwECbv2eCkFdht9lCI09etXDZzqYO79SXhq7EOHi9LGHcUGUfekmus5huxQZUdD
RBIj1mSCwzLYMdXKIrgt3Pw7VQ/FmLPLfWNFg01rWesNKaXOYF8C9l76jZgunwgyWW7reDwRPzo3
dZaap+gdLaITMwQwKxPHGFbKWmJ3Q14aiu/bueAVFYfRbyi1ZOV2L44YznUBunpZmv5Eug3GzlCD
1Bqj+PoZJHKlCYvIhK+fgRBNY53MS4ZRdLJLgDBI61ukz6Wy4U6nZ8YtXcrteoHmZWULXl+fF4XT
iAXfSpTjS5cvbZmIJoq4DrbcAD50ZnStVtjQJaGQpUp6UJmpF5GA3y9bFLv272IeMOMJ+yNnix/f
fSxUqscKftBPRPFSqaG4/cwqXFkdt0nXFy5eEYJflpr9QObOYADcbH7kHQF9oujpFspBcMTVO/Cy
tWwYduRyJDuMpX71UtQCdMLN3pWrtFVE+sVdX4mNsthSaRKQUVj6VIrsMHWuwhktnpSZhDzjm6UH
KxrjeKkptkkStQS+W4qYIsRhGKc/pX5BeDAc+OvHSpIjHWMelZT8yP5s9djQN2UzFYCvEDxVaGuc
FAPMNu8Ev8Twb4K8KOKXdglYjAq/WEc50k8Ta6c9z54Q21Aj22IZ11QdflKTYTZ+PLIZNtmmgkll
Nvua41h8NG208yTTDJghvl/tBfBLBvosKGsVXWag2xx5oMeaZEXQ+RrR0a2dmftS62kSOWfvDUly
oQYunB++C2XBwPNAevku9l49q+3oSRHCyQwzWxhEC8pzOX4lw03OCOr5LBWkVMkxcqAfPE3bjllT
SabVeO31f2f6SlBgS6ZmT5Ly0kG1CJbl3mwIghL8QaKiDwJFfwV+17W2kBvOfOxRrTSV+QDZG/3k
U/piCGyGvTLElhjWssxok9ppo7CxUBHjvMRL9peFWA88yebLpQBON2K2JvS9Kunlh/FbIkNUzdc/
+znrk8Zq2+nR2/fW1sJBsNCGzdUS49XuPlu9mcNGcG+G2ZZ5rNAZsabfZ1WwlEDqotIFXDvy5K8+
8SPVPta5Blq4W2owbENvfwD0sPqwpOSFC91GlYdESRHPDwVQVhmK9TEFMu+5oMNjS3ZcJm1oO2I+
6g+e/FMjAdDDqS7KdsLCqT895J+PjlZFib3GJfMGuW2TBCDjLQ6qi9diNtA1FS6rzCYZyzToRRJ4
dzKyIwKAd5oKceRpWn/LdHD3jo1p5eBxTkdi0SWOOK5gHE7kkL3kAFNOagM14t7st6BDix71nKxX
3q2ouHv0Qw8Vi1fSCb48gbdVJDDdTL2Btxqmdq3pxBtnsN55N5/UiELZXh35z106B8o41L7SfuFU
/yzRVw82uVuR7YG47ORmzCY12hRIZ7kSIPkZmT42zJZx4wSH5FIIXgF8qSyPaMz8bNNgwcUIIbDv
zKXYQwoRKs+WAvogb73MrmGqnCfHfR3p1H0NouVyx/qD41TzeR45uvLnrHEoYpD6aYyYfjwLYMiE
pgPLKoVbKA/Nxy38gVaBq4DTYZYiitah3eJrBe/zaK0gRXwlL+LsYltPG4v4UJxWM5AXacWt336b
BhKur0yno0J8yesgkxyUhjb88oMSysftXLOGdW/BwRYyONyGaYaLrjzscinBV20WDXCKIVJHuCb3
IwnFvYfGkUMcIgP6mUmJbFD8nrUuINY7gAs2Q4hbGzMRwE/9X6WFuHRrraXsIcry/sNpctkn3ClR
FJvvrMV9661ifP14J1kDl46pwhMP1NQxsH0NpYn4qR1KTjlYhQp+LZiufxOHSnJ1P9/T5yADaMAw
lUkZiutbCHD3iDTfhUo2nRrh2z9eu9h9fqUZuEcipm/4CDe2hxqOd0mHH/O1fGCMxfbaxA0RF2aD
teCMN/IimvhPIg/B4RFoN7njijWEL7szPPagvqte/0yZ/W7dCpW1q44BXYQq11DH+D013Ll9NWko
TxXVznLbk+xGysINZ1qPFOL8TJm1XwekdQGASVHeTzNhIlenKKudRliz2PttS9WeLwANRfqgr1zg
sLYoQaCL6kPapYyzJA8j7pRu5JyPor1cgt+rqrk/eLeVSEJFSrH8dn71ZPt2CeAle/T0K29PAAC4
vzLEmJwQwxjBOiLQZgZZTQxjTWyNho1u+CwdL+THJRywvNqB4xtKtz4FMdgHP9IKcFvvJuIFLEdi
LGXh7iEyTPm83vpINv40N9G7hH4ozCFdVFIVLNtfD7PBJk4laMyAnwI/h53mjIxFFFmT0i96OFXi
nL07AQphABNOn1JXPPBQNlWd+h4FKSX6MHz7nmIElRlOAujN4Ee1wdmEC1GuqyzeHaMsX+6JueRy
gczgQGQgC9/LvvkZ16dqBrt15NfaQr0J5x1hoOGbXl1mhUIRVVmxgqXgUhUthgs+G6vKDT7uwx3G
Ky01uM6XfaDFJ/J8xRbk/Rj/Kqi6S0GskgUbXSggtaZYBIBttSjcszWrISqTfwoHMUUze+CHrSzc
WbkLtWstas+cHVcfDSu08k0dsGSZDUNUgxUBW1MNrbTEYbQ4RcGvs/gDJRKexaLIm4vuqWM16xpC
DK4Zol8UvvOU72gqq4kML0srIaqiIeU7Qb8H3GRJLNyIs+8aOshlofoFaZcuSBTS1/JvXZEBdO15
Nc2FHPydUz5L5kmLv4DfiEzDuhXYYSkezWxjJWQu7byZkj70BZnH2nTXnIaaXYIUhvjdpdg8u0sO
XSSX6dHRRdJ6vTAygDq7UlHoSCSChaXuKz2UoqpsW1gqW531K48RP4kZYzS/hhaRek8V3pzLw/OY
sN/r95jm160tT5wU3CbzcfOelyyVRDXSAFSJRuf3hvFdZnvaJNGn71zzP5tWTAdcD0SLrbwRFtNw
ySl/F4GLbRWrbvlY+DfdS3tPTGhBgiuB+ICZ7mVKjAJjC3VuE+vLcl2D8hEhH8gUL2RMYsDRQVEK
g2NOCf1JF1SZ9ng+Tb5aej+DhKdZYj+qTono8uy/LgOdP6sACDvhB0+0Ip8F6TiQ2VHfkEPJNHOb
akbinaZjnxevpT+8+xyliWfqswpXHsQA/KsfTlEDiDPTjNfreqgY8OobN/NtzaEn2/zd0btwjaNo
nLDDzDSV/02JFMVZK8vhOw5apVYX/UUHMWtoULx1dhu8znh9hYc1OxxKnk3SWyxDf5yAePHlwtDH
w/05z1Rj/J20TWypfZDZsXNdZIDJNPKNPgNIZwjuLjkEjTobUk50SlT3OhirulD3ZYS3EBba/AKL
y0SkOnEvfyv5SSS5I4F5/7dn9ixK08pF+suOr0kuYIoGmJgkkYggGdcZjH1xrtF08NavzxRhNyQf
JbXNYIjB6tXoOx9LWd16QtOP2CmMWSWVfjHC8bLuiBpspEJtU50pp0J8swX5HhFj392k8XFRcuJ0
zQdHYRJd3Q+kPDoEEfxFY7POYKwy5qO0ktrs9fJhSySCrsxnJy4PKpjS6KYoGDh3D8wo2be4OAmv
OGBuPTk+DtUTzBdk7eCWHT8SYMCZvrv9QUjpoVAS7a7Deh2bHwxfaAkrFuRgUX4mXMs+8EIgXHQ8
Raz1JEHH8oxF450GfemqDVGUFi6s6n5nO9R0qh4Yk4PtKzyaav1uFCl79fIHuywE/5dIyPxTQiLD
Ic835EBn7xxM8SBIs8uZINzP3OM7dtlhILcaHfB/fN8djjcZUZWz3CgN4PAU/8itV9GMtmPQ6K8z
D2rwvMuJbMmyW0fMTRbknjWZgXUOZTN1A1PNdFokRikaZ6+avA8cdLBGXBlI0Gql6XkRlYYzUMar
Oj7rMktJFVlZks9qhLDZx2utn5rufE+CAMnoZ7rfQ1y7iclpp5mZQ+QXsdvXIdoNFZo1O4ojGstO
sKGKb9H7u8kXaUy17PA/qFnOSwxsAHQ+sd+e8h7H+X8QlM8vGrj7729QGXHv7ziKkBmo2p/JSAHd
6eHlZ8/NJ+6us+dkzI7CLcbqOYoGoP9I/IEiKyalE2i5GHKOpwSy4stKoHWqyH44DcE40y4OARfV
sveLgePtcyE2i6SJ5W9rb87jyD8B5KLmTQ1clDfdpr8TyYINIKa1+Ju4mwcjUI74Rfbncw6nf/IN
Zyv4Auj1OMtmApa2MFIHQFRMqG7Vi7JWdHT++Wczx7I6wcoIhXsPwjSHcm9tXbty6ozG+BwSuSMk
eRbJfA1v7ukIoU30UQcnnxDkCsCHmZTrupULM/OKn7eAGQ2GndQsA3yODtflo5WCfFpVn6CCngj0
Lflf0c1RFyDSlADfAdFtoz7WdktDoSx3oTEEcnRgqXXeEz2lSm3/BHS1dn1cVTKRXSx0NWRXcXy4
EME87WAxSiq+EyLxnFT2cAYWAgnJ/6mwfPvrEqtnEYS2cHY47UN1YtHWV1y4HF0wmqVBnD42PyU+
hxvXCQ85lVy6cZ0FamsDURuFWQ4WK0rSTmAEdz9eauMdlOVpOTSQJ5UIcX6CDp5wP4mshAQ67ScF
rTl3lFW8ny6uFQ/KhuohOfYU6Sytjet6Scn9tTZ1ZXmvi1gANv4fHdG2KfCNWKoyoLIRwqqUPqYC
PpzVinCgQ0+x9a1CDXUrjUmpxXXBxo69+49lg7dhW53BCJuDHuB/aMn6eOlEvufwiKDVPkQDcOqm
BlGYdaMNytqSe06qriUzqqV/GGx4LE49qCMtlwQ87EUE+DgrYiYLc3NwqEeoZAYmGYhAQttqjhTo
lY4TQXCZG2IhUJ70IYnKgGiF3krIRLT5eO51YzMfAA9Og/Drvg9GovMDyvhAS1h3OYcP2/ZNBRub
2/8exK55DNiRcee6vTQlAeV6BNHmjpcV0Hnk/VQoBErlinvGomCpVrZhD18zk0521E08R3KTKXN5
9IBOMu9H4RZGmhaKL0Tl6QRWQeXEoy0wqurdgsVzmgT6riWs+iaY3bXolaP8KM9EwrS2RrLMqWnp
15Wj16eLHwL7PDbXjiwEnSWNKsBKIP4ktpKqTUy5isqnnuLR22x251yl9DpBI2cArBThQAYmew6d
CZk3aKis3QIp3REIv9/6gUYRjH/YyCdlq8TVhYtkQLHU8S7UtkKQ+pDbIQX9G5OfJygZRR+NCkdm
7dD3ZR5M73PePMU6PWnMjjSjZL898PRS19QJB0D4B5oKhHtN7AJvzeCuFiSuHO/ZgVTyricEGGUa
wazugnVp98ypmbtodQDjXmOsPDfC/Ve6qLfXoMAiQLrtY224IVEvNMv2Jf6HM0SHfq+uOjM2clFf
zypKgVGTdb9SY597P7/OkyY27TUDrw7caqgf1xLYOEWmGqV0aemz1vUgF6ya1I0NprbHBjXNhaE7
LFWFCJoIjxYn1gm0yY/esraW2gF3KNBVPqkOzQlgyvxK2yOIVDMVUBrJWkqxLjxKHQVX6mIe5CsH
NznyHUaAeEyMFVkZd3BVTaChum5A59TWv0NUavvRf083kEuBIf4fjHxuRbCJJ6f5zHZtAcc7UUe5
LLlCrik5Lp8jIby3dzrmf301rLAxYsJE1eBv1tIc5hqntPxViWCHbcq6gWYLRPrX99NKslvtUtav
fPKQPEFshiqZXAO5zeKPnHt99I5a1eO3e3HJf4uUdO0WO2KpiGuPEnycAJPPwbfwelrpFBZLC9o1
X5s+6ASXwG+RuZBL8hqafQwto+cC8k6FhopttF9L7zlahaIMoZ8FLgmy42M2sM0U/a8bvUjzXsfX
RlHX9+2uR/gyBgKlcsrEZ/fbyWvYQKVifAzSmbl0zYRwczR6xORbLnxvXw7YdfTYigXuPoeRSnF/
fUkwg0WYkt/K+GenzAeDnsnrfoOf06EQaK5Gv+t+CY0eIYA0gHCSDCP2CMzFo8T/9rpSawvqDYSi
QR9+p/xgALQv9y4CmaSBD/49fOW7iFI0a1iXR7zCrVNcLoFSemcSFk8QDI3NwfUSDIbPrMaJNdtx
iYQBfafS03ZxA405yyWcDUw6PFNz6D5slqvmVfej8pt2zJ85W2h9GFUvV5Xue8lAbnbeCp/6VsHV
eqjbnJ/cOndrX4SMruwowe3QYVYwwvzkrT1NVXVgJN+E7HnS67TIDBhpNwYS4PB6yFicuWifgTGO
pRVI8A0R0WVSSi3usdHjWDcUQFMSPaKzpHmM3ErSP9ultp81uhxBMUnBhbS9WFRiQaQE69uTXSt/
py6mFZt/3QcTWUNWWC17zGEvjQDRfToVVUI7xP0berm/JAADm3N7UnG68T3SUoFFE/c86ps/gILO
ykMGFZcXqiZi21XIvowVdVYufCvBRlS/zft+l4WpzVX6m7GrROXxSv4rLFFbOklcG4fb93RkpH2J
7gOGK7N+wlcSSrkt/hzZ1pt4F94r+L2Wo4bt4/5xqnHH7G+psxpqWYZOWo7J+/YQCF9Tv5FU4PRO
YbPWPO2AO+ZrMwdztaR0bjxtjS8ZtYrdpzML90q+VVkM85N1SW7aL9AfkOcbXJ1O8tXQMlj9tE43
+4Xf/j6HngIzYQZGeyGdBPWt66ML5VWcJOU1Sow/nq02vzEa114jEZfJB+HV0MgdXbS2qt21dO5t
dKn+x5CM2lkUKnq6vKUj/goOAknVJa9ZTsS6678UIeu5SiZxCYpcobO+eV5hegWsZGvwKpOWKnV/
d/di+upBX2QKQxulmAJvfM3kpYmrg5Ubzw3xfFOR3C6ux2K16lxSEsxBW5PUgJBNIP6AgrJekGgg
9raPMK8KWnQ7KqwWdUgYm9gP4oecW586Q7HpBOgwH6kAKyTlRSgxVdlHg0zqYQx92PlBJnV1ABom
f7vhzcqDya4LHL/sw3Z2iNmiIL/l6EjUGJFnrFXpMCjivOohXn5ORd0Xoq0osfDOvtI/aoGIyChd
OjHJOQqeW9bugCFOGlvq5nRQt5Q8ui2DrMipWmYaLBbLiE3fyjIanVjdoUoFukTudrF3DKf8v2L1
8DY6yP6BzcRtgw7plv2EJ4cSpIipHWZIHbf7fOvTeg4c29DC+OFHWdm2gBIOPBHPQ4r4sUIVe5qR
o1rjN9GeCAL8KM6LHwf15W2SmVlsBrReoJraqBka3GP16Kbk7WuiXy0IDTGrDhAT51ekvPypQD8X
uDjzQXfy5WA3zIKHcZC2ByMkN2uwp+i/pgHjrqHD9F8gq/uJpHMx7nJs8TVmkOVMdkQlsL+4vYQL
joJ0Wo+r6FRelcGBbnEuE9XUNoY2SZKALVLHyJ51cko1dxbX98wboXpRC11rsRxv81c+xbR3cjY5
ZOPmFVYVx+N+SgT6+wIb3QuBU9pIe9iSkOCGLI2tv+GLVYSjyNMCGRyQ5VwMxuxpT7yt+rERbZYe
uPb0Z7rlRi/TtTD9T0o6SEprY3df98oVnUzrs6k5QbL1QUc31BvYFiq/9d0HFDdOIdQ4FT4eV8j9
yu+ClKPF2BkDKO5E6usROwxNCU6B3mMs6O//BPy6lBo/+dsIoJHTJYq3kqWyCSNABsAGo48ndn+G
Zedn/x3bm7rzhWzPYZP/b3sKWyIZKR511NrXXGhSvi+nIqIOPBYXeBt3g/IWnR8Lw1+tsLTKiiYz
kd4ib25MXy8OX6kiIOVOm2LXAY5XhljVrA39VFToSIrKWRbCziQJTROi128cnYCoAym5IbWewXkT
P5PKdqM61oH67d2h3eqiPzWx208ScTY8fElZJjH1CehYFw+Q+QFNirL+0K26SONdQG8A3i3ElLzB
jb2lyvCOl7Cp8tkBj6D2jfHoU3x5AvbGhIBI80/FY3xb9tYFZ/iSGkhYy8aarIo0TGQsvlPaO10W
CUvN88dpQbK7Y3FpOAvK7G95R4UzCKJfABZMU3+369Qqz27cgFnwsRnW/54+t6FI8Yw6fLsvlK+k
TSl928vlRQmsSLs4PV3JKr+9/KDbbAKefRrYijWmE/N00YKYmXgyHStGJu4ikn5gxc4vsKQKY8qe
At4590fo8IBGcmUIsBGkkpSD1AyAJdzv+PrBTdPAsnRc6bj4VF/ASGHvNhHDvWYzbmRP5S4pBc5k
2aNMEWT1YfJ99nSsInYokxRDYywtcnUIxASIsCNE0YbkUcCSoUCJI8pc6YSXWux0Y5uUbwpgBsgs
HpG9RO4xkDdcsZVsLD6JptpdtRlmBsfFg99407p2xn5K0pRbtiwEihrrkKBuNqHJPND1+u1lAmNh
tlrWUdaHTQIC2yhh4OCNdNERYBVYom8s/s/ZNroA8O82p3lBYgb2kQpN1ntEerBXJ/Q2+p5B6hCa
AzXhSUkLfc9sWmbdCHVGGnHR/cjSC8Q9c5D9IJdqQ7yITKt95hzH4w6IOTUgp+nt2JU8buUEpnOm
16AxHcZR9XURFtpzUtHhfEVmo7m3jGHO5ezfja3jH0Dc5lQqo3EYUL1n2OvD15LzSueIUCI+oWk5
2LAp2hv4ebprpcPz7235ufDiz5F4ygtx80L8A404y99tbgh+Q0XCalUigJeS02wWplkxRRysgpt4
/Ne8AJHHIIDJsdckthij5G2MdEi3B9OIkAbBEL8aGK5m7qJ+0CxIAaMC7kBqhu+AyUgUjBB3C3oT
wwAAY+c6KflUiDV8I9shUrgatThL2Qjj5pzObaH+PyE46THMgH9JmdnkPrl2mGYa3QaU/W6HyC+4
TagcuTMfN094eMzQbWjFLk5dy5XnZmMRPstsg+cDLcG4uIxEgG5T9DQyI7hVowHu8NHK1YihCSBt
MWzidm8fRFAHDXuHdi7P5WRZwRbCqs3Dy06k3Kk6QXBQt+EWLimWR8PxCmoRLW+SjEXqjfTkzpqq
StOUzJBc7YDy13yT4U7JXe9zS1WnjKMholV3JtY14lHcsvgPTZ+CgmSijb0Gy+aAPyCZc5NoHIUG
OmWwkc0GloEISFJVNEJXomoig3sZz/cnRQ982WhEkP47YwD4qcH3QVUaszMh2vBgGPO8JsrVJ4kr
UzfmD6XIvR1tPf4rRWtTFkkN2XEpLwnKkLF3ov1gQvkFMB4HKHptQleyVuKqmeICXhjPU+tIbbbJ
u021jCpyeq536z0t25xnVBgMgtVI4y33WG+EcxO3GNH1vx2jZEJzha2GUCd4P/ADXtCUVR70/08O
tH4TT30xZ4raWqPlXtGgaZELv3N3SaevKttJcuPSN/rwGHWKxmDr5KC0NE0+I8FGak2aIla4vWpb
4aZB41m71izFqmuNY453EhGXIEMuJ6ABc2yI7UOwZPp4u6Rs3UQH9rdlFHrSGzfy2uURL1HGSvCo
UtuGH+XHWIcTy5BSx9R9xC+foLAjtHWxsLO00yoJxd18CRgMHusG1PfDi1vM26XgPYSBT30AADAB
ulJ9A2mScQxrxBKSIZKJLlRUnZ/12nppxoJHTa1CsgmIR/DvAzVGodCy6aosixIbWpDO8aKpZmcf
DCB0NnuEBDOwZSXcrz0/0cb+0mSx/6qNxgiQ7jmdZYdIIK8ndYtOXM4CccNm8MTHClyU0fUp72rX
zkoLANUk7NDNKG7/RlFQIBNHquEB8ZjyFu0XHqXFG5YIud7djdVntGcEuFoeRj1joLqJnRCwlGNh
7wWHypk6wylwpAhir0MR8wGZKqHjpZSER5owD6/54iKuom89RB2EJeCJNc+wv+/hq6IOKGH+vjIu
gwQceogDc7+u3vvTvdM9JVJIDF2Man9+ij5htTYd8JzaBIVKOEMgR7N8OH7eIixXPsLYm4k/b1wd
uPFfjQVAb416adGtTQiVgFuxDx46Hhp32KIESPn6lq+ew40xnpoVvrMCIREGhgnMqnD1fi61i1yM
wkObSG2gpYA52ASMfw9/NvjZYKQzpFNn3Zy0gDzyJ5sXFeu6zYLFLvaeayAX6/WNFYXVdRfdfxvx
mPw3FbEsjYXn8AE84ZJzhX8nQfgWAU2LHgfgt0kdX+1K464fnrDVZMYkbRMHjWPvr2h+kOdwI23h
pxRFTWc7bsjFHZUvA6fpYLOB5f26xsquJzJxLuXRXoyQ95LjzaAUdH8EDNMoBZ8D5Xsp1UechOoj
L4bAVoSkoEqLbpdk7VA4t1sUXmxLctsOKg+xM252X+wFr2EgVzZLFb8Cen8ly2b605jCJh7TZLP+
flqRPGHOqIiz9CmL/4pmEgyZxyEXQjdBCfF7JeW7CvTgXRk4moLvguRKpL0JMXQ4pA/pcPMAX6Zh
Rz3DJABEPNbgj3o2Fugf13fSUTZSJU4GA9GwYbyMNztNwftSq3ZIaftXcHe6uu7OKP9uAoxhqFPN
smFnBPSxsuN0LF9ss8BS4tvcM6axgfqUR4KU/WpeObfiVAAVruAXNNMi2x+/sWfbn3j8sjUvcLgN
czEuZxWrpvVVeXPDynBcb7nZvVJlK0opYtfvwl8us9FRO+jq3J8ObRJnSnRSJ0CfSTtHJwCel69c
uCj4ikYj7zdbja6m4uf0rwjZqLe+nQaKjd4gAkzgoDLPDxXYwL4TzOz7q7eX1HEzcfoF0b6MnRH3
mMS3Ki4hmvmBPBO2bBMklUj5NKMwLIZFVFjLrCU9KXhplE/OSwkf4BoXakdfeZl5V6BCjPHq0Yaw
exisFuniGY2aR+DfpGgYC1dOg+DOuUgt3hypKKLF1IV9JaH8XQ1uD+4ZNGO/ButrlwAGZ/qJM23A
lxNdn/biUuLPP5Df8aKZRdUaB6FTDNor/WSxwyUFKNiiYqtO+FlDSWzzKq+qVkXY8/TJRHQVQwal
OTdysdXQS9pA+JxxEvLUxYYkiSWTmk3gRli6ur6wagEgb93/DUEfi3GlMwldsLVbB5KSyfj7vJBP
PouXvomNnM8FOVLK0EzTfpThsKUhu+oOx7pV78teeDDWH1xrKCRqnMwJ5wKGcgUE4CaQqO12mP88
AMsuQVa6o+ju0R6bTiqfgELvDr+p3TvkkjFAeI8x/vvwr7/D5BsLj7zQnKJ5SYMB7EVKB4ogMZjK
VFUpIDqgOH+/coplrf2rqLkAFsGNxQuPDCkN+SEbuwjyxdWM2ce14D6K1fjx0zlJvrZ3H6NplkXe
YeCWgn4XqY/9ygxLyS7l0oosAur9HdZbBbdkMV7X19fng/nWWbYqHra8fI54JvUBd/p+eeXkrywh
Mwbv9PipzCJZo5EM1PaFRNI4mZhYpbR6YZ/X/bo/4x0d8hBkw3AckIzQQtUl754kH8IzssmPQJjw
Ox5gHokT46PTuUNX7egjHc3ZW5UVylFUGuKSW2OndwG/u/RIT74KRzFyQUsuRJXJsyro2b4MX2IH
jrGwFzOBDX0/NYhD2rynH6lWuW5GJhcSPoYP62gdFPot8YXlONOOKmJHJp9fYUq8MlVqFQE014aY
qQIccOz8lfo6q8ND6/FKBU/gvbUOCqRTrgovYFQa+ZSj86sY4fO4hu3/ckyPP57fEWaUkx0bXBVX
IDcIBAeat3+U/JJrHn9tC2k++NeDQ1zRNeoqpvlfUf1EbnaDjKgeoqsn3kaxM7R9P3rkFKxZ5EKk
tFwdZ0+NXTvbtLytFv5VLVeyYRcBy3Vdv9kFN5AZCY1zuQ66RM6iWXEKMuxTxCxQb3BbUsNQXrOw
rQZkNxlwaakmdRi8i/wt1nGEexVhIkc2Oo/DiHzD0s68ptQ0pIBJWVADZUNey+e6Eg9CHC8Y93+j
wnoKkKWpvWew8mDmG7jSxlCbJ2KKJuFtTO1i9TtMHUQFpQO6y90dE6JxC5mfJt2pKGWR8AZlh3TI
Wl419OC/dfc3LUNiIEFeqjLbEj9ELFeHcMu78NVBxyv3Dazcp0cyIsPe4OJVQvNafspMvLinAzr9
akug7taR/hQGxPNqwqVotGZKyJNDq3Tks7Yl04ONiwBaCdSTBREgQCw5n3qyHsAC7KdLZ2hELFc5
Z6+JA3b7ZmkwPz6SzyPdHg8pVC6YF0FwryPBBP8rx2SRF7QinKu/6f6IuT11qhk87ttXd2sAwSk8
K3vsTc7YCNo9/Mv/LQd8G/6v2imx0fBy6Ji2XTLr7qnE0Oi283GOuYunuEc6AUUcbTrbGfiDXZYP
Ay7GIhQ202y2RMMh2FeQkV65Y/f8ZUzLoEwgE3ph2gN20pGpWowM2PSzEMoklkVnrU6/tAtr5VzT
8KfGlKbOFP37OfIFMocOi0MZ6ULNSvaaYvSMTyav3+nxQBhXzDspenfb4o4LIQBjPmUhiIApWf0c
4if46LIay8n9OKivMetrWLk+W8DDygqras6rYiyRwmVrM3bP760LgqYBfJrcBPQJ2C6/bRIa8oiz
5TzJ6umbrHSeRVMeKDvawkWhDcGOkquseyyGjxpf0DPF7Ydbr1x+7e5TL/iRaSQiIKHJHiHq6h47
NZR+Q2gthIj+mDLwuaoZB9Ck82I5yA8otgeq9mLk7H2iHKjXqwAq6GTAxurYGCFfdBEGNERIBoV2
G8jH1I9mWXb4WZoYPiVzLlMbgrShykd7LNx7m8f/p56EuzRFYYLp9QC28+HKfdrOo8zn6mEXyywj
VQWZUHRkpvOitirNu25fdjpHV932m6HZdJyW48AfqGKZR8eJV2/lJsxlSyKw6cYUJT1QxtvDs4yn
wGf/cNQMVbXT85R1qzL/1Tg+Lc9c6rJ7yfGvzgs2y6Lb/1GcOFYqnoFjcJG5zFZnfbpM+4myGrEi
2MQtWjrspEPVbHLD/4DNvxauw3GVuOEbaWLwQhwBrvSNWxVDdFDlNhkFqvxpiGgk38Vr4IkuqEGH
EUULHvSKTUgq15UdU+D18otMSLSAnh5t+Crs+nGzSQa1b98Gua7Rx4v091GHwa4nc0hq9nmDmbF3
QZnczWYqzptwfAklqJu+BOUE63hkLdqAVCIS/rB3FMO06v6lzEJQCUihKTS2tRTYswdgo3PjmJeE
nq3yWyonlXClQw4Rmtk3UxQImf1lMApzm28a4knB7BDMTid7cOPQOET4mIXMm0YDqgV6GganEsIM
hjaLwcGBN5WunGR62gBYsA+mz/N/XsoTYx/9N+ONgohORVlJCwIjzF1mUBICX6mdDJFgbKyKm4SQ
SI2lh8ckXVLbFiUn9C6/EVDjuvfCVg69cw97Nbx43nSKkewSD7kB+5iTehJFuthgP6UW+q6Op9+c
B1CiKhMVSQ3nCA/jpDW9DJVJ/ZaQJLhIgN2V/13HPyGT/yc3dhPM/9LfZKf1iEmS1fmBNRyvueH1
iwm2SdqPqvODg1VxeXFAqsTOcmXBSKi9DwJDSmoJ9P9xCi2gxu5NokNaE663g4pXseQBRr+qbwSj
V+LWtT3HxxRmIuP/vtI/8mpa/Z/OyzauFwYjVhwDaPO2tuFs/r4PCU0KsABGuLQrfoIkOKQLwaH9
quxubr7+8s6JyUkklJVJ9pk5NpQerrPy3Am+W9b9JHL3pCd+qyrKVgjN1wIMBBqD/M2FkyibdUP2
wxEevFT92eX4mV72hvihHKcXvWo7GHM55g6iYKAW8E1oQK/6HHbpYptR8r0bfSLacRxerMD8VWUg
EKju+hvjB4AFphvVbcr3lHup49ksLnSBjSSjlog+Ypl0vbmjOA9ej/QVp0YPFCTXE5k1JGmJnYr0
ySYbNtG098n5Y+kyRk+gxd6dyTpaLLD1UZjQ+eoAN5Rrn/VXsWqduqeqTvc++SKeuYdTzffTJZjF
SWpmiu9bt0zLRxvZfrJ9Sd8gXb4M/e+NqePGwSU58sV1OxHVsCowy7Q7FwIMPhNLcUrHnaBzUhFA
nC8RpXMgDMkOzo1InKrX+mdbcBcP3jpSoEtcQrwZrXkfWlt9yvMW5EpYeWBDJuvcXH4D0ldmZDYN
TBDVZ4qC4xvS4c+yrdjodHnVGDGzHx2CCJD2vpIMcTHAf2whCI6aSTPGRB/dmrUtlpHSEt7X/Z2f
7uVzN/RPiZcEiPOGXyfaVtxWR72x6Z557/3x5GsG6MppHa2/DXVR82vcH96MsnKZ1g81PoWA09xk
f3mWlnaY5js0icoLtQoJBt/ASGxJTYcu2WsEj/uUSffu2Vi0VUl/t8E0CnShWY6VH6W7zd0pz648
p3HnLHJbIMmeg8o93Btsolt5Mp8vyAj/TZ8UqMsCEJOokafuW8WPKBB0Vm+U1S7QH8birz/lG8Rn
kuCNzskwl4DnWa6pRFIwITxpsG4UpVJiqh8c9F4aDqZY+hbQNUdUrFqpcCT5FFiEjndMB4o9k/PV
8KYNsL+AspBjac1t94fBrOfr7t4b/ThV+RAjOqPPZto1m21r5w7zEHixz0hzv0XAsJ4iW7cIqw/x
edGGG0OJ9J7+nktBd4biwOzxCnYkTJP5dqVfmyqPxPtJRWdPshEsEmqsiCve2tujBX4N5o4EH4sE
ZDpLn4UNXGekfS24S3YuPNMBwb/c8/efuMiykBfLLb43IzbsUC9jqtVLAbhhKzeYdWsrxqEvbJX8
hpG7fxKGPowBdccXpDqA3F4Td5mWq/hruqBaEiaEZQm76Dcm6MvVnowDq37q8hOiaD+aoV9CEUtY
r1xJWH86kcQWce1pdKKhaxfWqqPbIY+Gk2Ri/eqNGnDUK3pzIyt1PjTHnzM+QU1VUSabXI6rtP4i
oRsY5g94om/1NOFpNnU872eqKQWkSfYhvZY8AeNQmriyEZcJisRYmMwdqgzyghtHVFEwOcTwhgI8
F5/LWDu7IZym011kpR0qVRABv23J6yB7ti2gMzStrhz1JkuO9ub+1JbTtXs/uoRgJliI9ZyWZig+
A58qQ4flg7/dmbW8TqF/nCy/VfBvP0zr19Zbv9QogsihJnqwlQqJeNKZxpgrUlMBjNjwfWQCBNRv
bWgMnf676gfYXGTM6XgFP1Jv39hB9uboalNCfFE+pMPqddqxvWlyHIEMDHKvMzs0Se4gMjOJUlMm
bWyPjPGyu5dTbujuwLj+2pVuELWt1uXNvaQqvEyC7qSR/bfwLv4NWe1ZJ9UBl8cv+fW3EZ9l9yCB
7xr1v0C+Ty0j1Am6vORysVCzwPVlbxkQirTvVLFjFuoYQ9gn/j7h7U1d3z0nnvFzZpg6MFZkuILn
bI/q0i+0n2mE8q1ickUs0M3VN+8RkXLN2dPURmlG06K/9S4sI9AurCsPLMpPI2795MkL3gXwCeNn
A28+63MYNq5dQsqAs2mylsLaDO/Wv24DO7fVUosHTe8MtnNWdWMZEJ6VXxxtduLMkApwiZAaz45h
ij/6s3ATuuV5AxPPEUOzzv4iAadNSWJk2Gyca2yq80A5hI8ZuX+uMhHEEG4m19Tu7bhqcZY9rlYI
T9a8nvYkbb/6guOuFt2HX8p9r+Lvh0AKIUUkUtsR6P1a9RkIhYsca4j+8Qu0XI3A2cxwViXxmu8U
bXSGeAEcmkf5uVyGkO5zST7vwfkkzqbnSYjOm7N0f/gTv+1XsIMNU1DDd7RKvOJqt90lD2ms7sXc
+rkGAsu2ocevMsdz2cXQaLrqUWSpbBMLJnGaL2If6vqRNhtxeRWACC59fsDsJMvzXCg5nhlNFLjM
H6/3ZGnTIVxCVJF39CjOmZs3SEhvzVKsR2/cct3ba0AEaUtR2IOn8TLF0LSgtIQyaCzEcXTY9gcX
/vwSCHDigizx3WUNyHAnvI4qY7pDXMMxWTWExK3RHqoceQwQOyAygivFk2KZ48JFY9vxjH/qr8++
HPUp5PA6lI5Cd0mkXc3+gAhkThMsJDcU9dmUt0gYjZZjkxTFoCZ8t/uZL+Hy5nwlOXrHmQFG6Et6
6K7AWv41GKsuzEAu35lxMNL3kQCa7mJNogHAiC3iNKl5mFroIxMSjXbOL4oXGpRax3Jdx7qMVfnc
x1ulrCNz/rqjpfO84OvlEzeFOKSaqzuceacF4pfFKBdUhyc1k5j3/0jF6lpr0wSy6Al/xA9F2ZTz
qaa4xuPKTZct66kw7iVPwgJwpkUEsjAfdBeFG2EzwU8kUKi/KpF7IdpOcVH5qvKDJxa8hbNBV1Yo
nmrgrcyVebfpfFWJubfKslEeCHUa+pQbhach+uyVlItP16j869Siy2pdzx9LcA7MxiSFHOkWJs0l
J0dsgCNLg20kznmSDeuqe0Nm5oipm4CsgAjqGclLdG27d0vd7awzDSj93PpVKYut+ApbX9ms24MG
DI+9WG5RJgc32gUXoP5Y874eE3Dhc5Ru1QRH79+Ubm+qxMYyeg9ex//Ge2yvK0Np0Cjn0dKeMBJ9
Iozwp28a+jjLygi9dEyDXohMWdDU9uUbya9iY7Uew2J8wCM/0RjM0zVj1yZsXwDnbQe420/9+9w6
+096NXOS8WFkgIk7DTRqUIUlB5mF1xXvdTSfcS7C96ENUY8HUBH0T7Dr/8VVBQTpBfHJ7j54sAbl
bYBJCpHCMoSfGlVNymaBsOdiVSMTgC/2k1uBsjWwRNaMF5I7RXSXOnFUKlYoC/J7ItASRLzHInjK
frfzgwXD3hjTU4Zddaxh+Ka2Wd/eQbqCKz5Y1k5Kcc9AXnrmHCaN1JiT4qE5wLLS8JTFAhbVhS2Z
+V7yLcMuxpHhTvByxgbg3n3xpNQg6Bc4Q8cIz4I3u4P19RE4Ol3N9RoTO1TlOUww6ZBmT52jB0KO
JUeXiMjYVg4DpK3SXD3cdQVagF4T4C2RFm51kFO4zjdP++6hiUKlUfo+dLRhUdj6EB5r6Pf+afOc
xVHwFkSyuXNg+ooTqcuRhdmYaUavPp6sjppwRBWD2CbWnAY64uNVmst5SoZgiYl1k+zOaDbNbVIK
bjz49MEZ2K50m/RzYZQ3wSxFECm8+DgN/JEyk/M0Nnl0+C1Jfigb0bZxZPOlMFQNHMLEkFBlQ2EM
FbqrceF4Klz86vH54n2QuhZzjFiWqeZ10nXIbk0tcuLcdYZIDmQaQFBXd/+oBnVPScHbNYkuJCAu
m8+AqRoUwKNWAlS6ozoT5x/kvgbFhN3bjyFFnwBMjdSu5qct0wWkO98wgKkc9DUTcoPLg3HxT7mr
4SPio493RCta3g7d5oWUWu34PVGMW8nlYoZWfvuMEOe/O2hhKBaWfTNnWuitJYe7kFJCgkFsev/A
rZR0v6I8cX6/N6aASYKrBNO7hiMofApcnqLFuqQ47sUKCi3EnRUCg4n3FTYzImfpx5QbimyxXXWM
T39YWFE4kTuTsNxxGpzIYk2MqObwRVRuL6Mf4xMvlyGxIKsjZgdEmWdmu5bV6cYP//LnND4SF2Js
GeXtnpODb6BvmucPOTNZo41P8C+iZt3r1w8YT+XOnDutc8YD17F22qB7LrVWgkDlJUfsX3k0JzOv
oUGgZIPq8YF+ladkAfNvP1rOlu9Jgpbd04TCN+En/27jLafilO96FiR0PRIdKdecMASB4Ud6baUZ
i7SQyD+7whW9TxkjcsffDrlRHGxr950LI3jdH7i5HuCCVp4cotscWVQsrOnnvTZLb5LqrrRpmpGh
K4NIbCVGPUGdPdf2m9cyndCEV8u+NYptzaQxv17T1wAE7PUp2/SgiKHptWXmNBnOQHawRn4fKrh2
Rp1xOqYwXPNPLDUxE0GKfkN3O/M53OwWzlShzjqVyOd5MnvmrnMTh8S/X9a/tx76OpiIcId/k5I2
NF50QPtqjTOnfQHDYmz7SLp0TruCMkPMZQfFFgjkDgCoDd9WUNilGSQportMpkXsyOWXFqK1Uqtr
IgjP9Up09ifxABDnKJ1jTMsWOUStCpPHF46r+LGX9L0UQctI3m3Vy0SR8LJ/r8qcAptUcJiODiA7
STqy+xB6p1mYHhzC3TP5ESz5xFYFIA+kOz4DitTwOhx2N8FOMFiBD4jflUKEyrjdqsF38pxylMEj
DTbCv3MDPNGdx4+lJBQbt0m8FDYaAUG01LpY4jFQEN216JhrwuRhaFeq3lA4ATQfHhv9BwXDnwRN
trErNESZRj/Mz2nVoD6u80K+2Yh4qeBsnL7zeMrfeRlH6Wb+tMkCxOwBjin3CdPLNAY4yiOVRaJg
0e2v3QRxc4iaSYkUfLdXETBUqkou4Jgx1HZf4ALQRVyDjb/h6Qitlqno8L1q+gCDFz9vguvcSiBm
cTvUbGA/0yk+SSQl27dxYvEapwTr2huLBBWQZLKd/ccU5xxaddOGCSFmxTqliGvdGn/f2wlgkqGa
ia1slOv+9rJuoR4arUScFKly0hlR8q7I4FwC9er6VLh1tPJrUp/7I57/W9KGpiLD5ttIW1fc0ugJ
ayHzgoD1EC6y5ZwIvMentH6JtoeNWs2BUU2MKnNemgCO9S+F7tuds6RNks4bC8wZ2mKC5PzPAHB2
19Jq87+gqPJwsVvV/ATYsrWZ8jskqU16ddd7GBvk77xAkobPZ9cg9GPvWnOI0LF7sY0idLJXN9Vn
6mTS4Z/7qaNrvMIevoin/u7QBoDDOeUOeGaTMh/ySJm8vt1T6t0Ukk0ulRxZMnDKVA46NeZ3jEax
w39i9mNnA+e3IJlgXqu0IkkwZST6DAKACSXhti2uv+l3Ke3P5mCm2ni1W4pFz/wXAroMQCj6lDyj
riqAXF0gBHXbpYFvalEJcnruclaLRsUYMXtKkwVoazm/gbGTC94mY/cXeDa6G7KiinYL403hwhEH
0FZB8YjthXqp1opPXYhw56ySwLCq6W/iq+effv5tvLKuNPp5lrYEeLiS1JyoAg8ml7X3iigkBVWN
bPXmFlueF3l++GYW73s63QD++SjgOUt36kt15O7FJVXP5PhgNDzU7ugMvp8EBs9KBruOZTdpTnSp
XysYrIWmDxsyZ4w0XxMSgI8XOAzqkLzVKdMkZ/G4f8xHJ1Ef4PmFnBEf3KV846vD9R+JwhPBqegg
gPPaCjYjX/zKtDPYR8wkniFaciy9Kzk5XpUozPjI+psXwEymMv8q3Goid/i3MA/L9LX69lUQADD1
BUAmxKq7FtrOVCvqqVKTJeuZRkI4JkMFqB7NzBj/ADoQn4TpfSbmGzR/hoDPZqCBzTN0dMtlv8sf
A173sbhgVUcre/6wErOtS/yOMAdR+oDdUeBvo3aOZBLZpBe1u8HxBFmck97HGwCi9F+Xc3Qq/CIX
Penqoxan3ti/Bv/cGZ3R0A0W8BW7mlO29Hgj6qQYvjAswGbwwteHjfl1/Me5GXik9ZH0rhj6wmpb
qAWqqcISyqxUwS6VPgC41RL9d310Z/2/58GfHt0xVNvIouokwyjb7RJqbfl83dPbZdMo0/o04tUF
w/c+C/KZzqPwGU8pIjxxUG000EhAKz7zRXFb2X0ecCbQJD2oQN06IAqZsPjUsywDGDq8Dmn11Kg7
joke7j6cjwLSenR9WT/INNYMBy3yO1cQbRRxVrTcUYYrad3LHYCMj3bh4C/N4H7lnGaFvig6WC1N
1rFw1bn4+8M5F6F5hT8s6DdTp04LQmtZJTEXvnQx5A8+oKryI5UwMnQNSl3Hyws1A3e9vuHw/rrw
vihGHePkMOWX333DH84mHg9o8+xSVwUmv0uL76ao+vtmH2YhqrBed89qXjUsfAOQ1VoSVk7+fje0
mbVmPwXqgkaSfFW3Nc864BTgVy3HwUUcvrCL1kgwGt5nXGS/EP8jhM88Z5Ce3QljrEzaUNsRI2jh
8QD5sbQRgK52ano/qGFoJ56lCKBSFi/e6Vgl4sIlMfe+q0d0cLxXfcKqfQnG9+/ZfAgZr5p6kt7f
W3r5EBzNXnnlEIBSx6AmZ+TZSrzmizjUe5fpuL9xnJU56t+TezFastd/vPMMDECXy+59HCkk4M7w
YqaPmPjJgHrFo6Qef6Nxo/raBhqJhsd8UGq1SR1smOXdBgd/xeddTu1zoUH/yWeUaU6I7aLcXw9p
/4F9t+hg2BATHneje2+vzFY9C5rfm5+mrnX/NVmSCvcfKZdYSuSqvShyUN98YIxxSeF3d2X8CV88
3ix8Wgo+L1qHhghPfxZ49khmb/hvztdhfFlZETAF1jY1Jb07EhWwij7UYQVmp9nmYqH45dFd3Ryo
gshNvfe5f/ZIseeNFP61qLPZsHU3aMdXGMV1534eOyHGc+ADlMgtKQ7eP7PcOXUlnL7xxoVLdWm8
gxdtYKPg/dZD2bieF4TMlbNwhv3dE506WTkbQ945UZ81YDMlAXshTeZY1YMXwn26n+d/X5Telwlr
R2fUmBYtNV5mFrytSXVjTz9VA8b13O+Z1cBrPZsZTfGlSH18lR+3jqZRGDncFqc3ID7a7vTfWCLP
u73rBndsWWFuGhggl4ZQhlStQjUczuMaRC+1YEXHsP8cVkqO8zSWKG4nfqf/ZyyRC98K8Ndpkz0Z
KgnxqH2wTO9zniXd1FS65BhgbXsk7C8bP/QNmZwPPLkznc245cIjggcuWyNNpC5/2belipJpTtpt
PnLxo2D/tNbOmLmhQDrBh3meaK6n0us8OhXu776NDwkz4AeouFmsMn3/5cd0A7xZNvb3ylF8p2sy
qFQm9FYCv0baV06w479pjzMzTMT/ECjRtFX/BUK2y8V7pKEhGP4HVoKzA/9XUqA/ja9I4ZNcZnPk
JCkgKSMuHEaR2C3QXFpIx7VvbHdSErCCkZxGT1266uvIlV+sVYUpemo8SXS1f3kur9b/19RJCVdu
nNApQ3nUFCuUT7SVYdehHK6JJ1Rimr9gpbNkCY+g30nJBzUnnb6G2cIdyB7LP/rCcY6rLg7yN2Re
LPh3ej/N5ytkp+rPBKXCT36bOcoojlEYuKZKIuvHRhOK7Ixihlks1cX2yfgYb+gNbd1FsVte0i2p
olQOulkjv1KAMm1p/9ujcWyT8NNMQf2A59R70qCVhw95AzpXHkliIVsmzzjwpqmqhRioD51IdIa4
HitINTaWirZlve2bZpSFFJaDWaAISXQFH3AO+Gy+YZ27GhK6wdiDOYv+hr+v0PDk02kHSwPVgGb7
fNt0MAvcqxv9teLihTly63MJpufbJEud7Fg2ZBAdfLyjvITEvFE9K1ad03sluvfHOygfTMkM+8lr
utCXW8Mdb0vdneVMQ61y42QgRbnMOUpnIIrYJANWZs2lEXPyFKYu1nR42yzPqwwII8WeqNhKEljp
joJ5B4u7G1H1iWgeDcnCq/g4sjFQKybOGtCqLiYn/6mhgXYYi10kJXoqn4+ekrn0i0frUCUPCg6F
aid3bRn3Pzd5/ztF5VuNj0pFkTbSsYCXwof1rNTKapyjPOga202I31ZUtqfjDCJAJdxuV9blUZfg
Qpz1Z3s6EOQDYq/7AN4fCiy0o6YcHROpqi8je6hW77GDjkpKzKvsiQ6IgEpMEw1kxLHqtAEYvFwg
25xKxiaS6v6HJqeTBU7KglCWeZ7NMMDNe1RplJ1XrvFJk6G0kZB4eNOYCrZQL0htQ+XEx/61Z24h
F8FlS1l2ba1vLuCR1QFHXw5ifZAviM13O4yNP7BjMxY3yNV20CWRhJCf4kS5ZKv0GTSr/c4/yysj
8F2DSqJL+MV0LL6RrHnu1KQDk31Un8w6i/et9TFdndMot6Cdf+HJBcU257qoazZS1avC1UTOhz8T
6pZmygd1a9ye7Bx/jeg4gTO6fo0UW2HEJ9EnLZ9UHP/k5maubAPfaLi9LndygZaoqkndE39v1FEZ
ChAVC4fZJsmFLvf21f39ZaxsYfdHQxk5qc9Bs6hF76RLGU2jyEYBYgDkPUtmpqrSPeXWldcIhaN6
SKxgMt3hCMMSSXApdmLH85d2i871LWKXoBqFw1f8bQkRXWyd4K8WUCtzjl41OHDLrR3Ll79nj3J9
ymakEGCyPuly4PseBzNqAeOuNZo7KLBKb6QYNKrZj1usu8UQtrRXyC1TgwhYWTzJEAbnwf3cr5N5
8Vwi3EhCO6Oe+jWrhPqruSE5zKJZRwTj6xQgi3RZwHW1TYnjQbE/eG9j/se7kdXNX3v954Et/605
cLur9su+sbcp67N9L9FTrLj3HjWna9igZXajBKyHsoTG1fQ5NZO18b0N4ql/ZtM1b9ft99rX3hsw
CyZpiRs/fwlkyL/OsJ6dwfxsI0KxJt1xYDQ8D6oy9EK+qY27rcpSOvAwW6zW4BYBgSFDrx5mzXeD
jcKXSdrvt0lP6zkxphwlmCtLwcEg3RYkqLSmDD4Ccyf96RARhi6NfpObxxI+NoJTCKKgCoQj0kqG
vjBnRcWKqiZ3Rb95lqnQKJ29uP/pKN72Ugj3krHsnymqquClf0SRsVspO39+8R+YGcwu5KAoco1Z
gKn64+MTYdX+GtvcnsKjZLCDEkP6PUZKUJftB/NuD/0r0P75ygauUpoEAHEhkVFr1UHmUNytin2L
TEMmWGnyQYD5oLWZgg4JiueR3BsJQhhvduVzLzVplpDaF0xb8BpGJ8RtvLOi9sIVQbcxRzgzz2i4
jcLiGZfCcuBAYTGzTMXBnMLOUHbH9CjO8XYrAIoBW4VUgmT83+Mx4nFgQH9dhfib14TE55B3apvD
4Bh3aPx6N9kBon2I+ymBaeHcZz2xrcJAMtfTqCWxLolvRGqG8rAt9eRR5Fb7nU8xKnIl/I2RCfli
9iH9Xxi7laxewIZm4H8JZxM79q8xH4yI7nm3v2z4CW/gEJtd5CkRx2xou/FbpHDa+fqJe1kH5umu
A7KaisQHGHEz2bjLV/2LTgcaWSTE/NbidvZRMl5BkTALsiPYjqnHTVl7qfkZ1v17DUoZIpHD0P21
PItM3Tf3ARqORcum5EdP9iP6rrCNHCnFGuhNR1usCVde5cEmBO5D9dAyBCBY1HBLKrB2jXTwtZMm
86yGtxD9qjrNpW9W2TCRJTc6ZBpr/WUfCdKeINHUxD7AJ4RWO/Ii29im30Hb4HUsiaxi63ER1gss
4c9kLWNCXWf6sUA6nwOHH7G08XBzbrfrDVfwXr4T3eXKc6RUSqlPj1FlfX9jDYejCRDCN2lLMAkA
yj1GP5SqmjX0bQ77svh9B8Cl2fBxQgUwPSqwpXWzSy/pkPhlFNvG8OmWQz6lgizIEwZvU7i63r75
ojZDmeC93c5ulYXfn7eSK3fSWgnHOP8DVcO9kuTcpr8jSQSTmASooeaRWFOnEPHSl1mLV8OerBBl
A6td8WAvGrd2KlIBOv8w60FI8H6PzuzkM5rNOQ6CLeRd99yM6IZscZBXRae8ZWFw/eKZlwo4OLS+
UQAAWLMRxZt4K/n7p84gJldEiCSRzShR6BUhKEiL8M6N1zBzDz9E7IX0lsybYhg1n9HIptBq9ZCS
CJ7Av6gGyL6TTvelDHTzRi5T7GroKOSp8F72tH0cO7d9TtyTpOJIoMETMXHqFsYV/kAdBmHZ4G2y
9MsZ7GEkCtwsu29fZaphz9MkGk9YN85p+fkw2u9hFUGwDf0q6/9J7hfVS/9cUedxh5NH6a1w5Pi2
AOJkKMjVZ0Db8RAAhK5TMTlCyEgHwBmbxkHDVsrDO3xGEv7eDTlPmOuAaJFIBLD9ueD50JwpN94q
odcCjLVkBLUIDvISZjRBrx70CXN+f6JYti2Azj/iIhVx4sbgiVTgxMf3GkR2B1xfXGUsj/GrxIbP
KQaWc7nxVilw+4U5yHHWSf3lzadbpUXVnyTzxSxYNRYUoUgQd6q9G2Hb9FYT0MOnxFaZ4YgFg60y
zdChGYkIAWq85X+Dj5xaDjtoftCJKLkgwhBTr9UiYT7rcY5QjL8U4UCZ7vZjhMqKTMLREwhiNpx0
noSYhPvSZeTI0jxrSEYaRIhvDhAQbVHtiquuwRzeY2XFdpPTZBIgE6v6xN3OYLCXNfEK/5j2W+vX
m9/GPUb9UGPZjTVl+TlnMagWbcNozWJetpZ5lI3dPeL2gsvwhvG3EJf7JQZ2+1DFp6JFWz6BEPTG
RAHzlrmBfj1Zru4Epn5R+80J3k5ANAaw9uPfDOIItX5p+5BAzDGhmi+OKBY4pDq6ZKvoolSLUQBY
HUjjqn1DvTq5wWxYiuUV1AfUiKBeZalzNHihDXrcCR9utLQ+EPyCSBLmWnqDZ1WdqI42K1t36i9o
89YoOtkZ61I9OS5wu666vhahDQF2Un59u6hmQdF2hcV3xdccD9QiEdsMS1vHGcI64xmDtUqXvo9g
QOxkUBWAtOgZdyHzmWxZwUliQauTlPNWecq/apHw9qiZo2veA7RZ5WkXIumumr7BpTKnjkTrv/yE
G+M3bGMw8XMwFOHTQXrRdJ+QctkRSfCQLLRv1Z2tG9FBGMP/qBWjZk/K/Ad15f5T3NG3aq7FJYau
3yPPUXz7BcO+dzcv5Ph15H2ayegozVQzvFjhYeeoBVOzxp0TaXIHZeD0xYZjdu+5YkqKP0SGMLTL
xe+K7b//AJlfNRlew6dZOXLfQMeMuJ14ZQeE4wP2fgQUhvZQHGKV1EQ31YIlcfB+xS0v/Jqt0DTl
gL69vmquU4v6i2SnRsx0mpH8giqWLwmASDU/GmLC38TXcLhgTLyzHUN262IULfr+9AM4mnwMM9u8
xF8vJWBstskcMNY/ctB06l56daKJe40fBzUgZcsudEE9Kxs5tKx00HHiyJlM/w6vwoXSxEHVSzeX
opWk3+TGK6uJliAPWmIUs+ajjmtd6/sQVyjHfomvCwJZWfX8nna3oiHTyQxtZrr3+IiszPSfInYV
kIXkGnXyM40OmW5CbA2+wnC0QD/k0hNJkbwywKuAYS9Q+zUtPi9bJFi5PR2qsi/b3xii9/vbmwwO
hlDn7VrxJfy0xUm7RJKghk0KT1tAU7/syH//bhtaVa9UKEY/AmBcVR1ijZyrLhiMNIhyRXJgZ0jn
n1NjjnGkmeBYDDr38pHlV2p/38tNXZOcA3hHKP3D4n09b7PqEs0pYSjVgzOWINh2SHfSAPIfQudo
xakjeRXIuv+h1K6to4gogjaA30g5bPS5Ty+ojKMYVJ0OKXHVWWqDNql1AvFLzOsTgJ3fx+avO6B9
eDbm69a+hBOT50zXIIF8d3v2f9QHXAHscLp8Hq+fjYVu9v2y0pn/A6tzPo045LpfMeJBPFYG33Eg
U/uoqp6YysHUX8wbRnf9HyN6pRKmWGkw4l8JpgRbOEm5Xo9TtsZoD748XYsrE7TnHNOUdm6U0eAB
kgE/eUdKpHfpnCMx5U2dmiW1CyEO2EfsIn4CbieTHvC7wZH140RKfUAziHBOj2eNdyHOnc7OG8li
T5SEh1pMfw1O4cWhmAvcCXFV5PwR2VJdFfXn0/Wnge+LrB9/D3pZoDFjUdSpKq6ezaXRCQ+EtKqz
bkeNqGxW+EqFNen/GnZiA51iWVPPvi+eqX6NLi8AhWYATAx/Q7Lho4UC4uz/ySfNw17G/12fgRcy
cnchW1DiCCREC2gmBP3dRtaep9FLo+zqmiCfFxRXnfYb6NF3U3aW1TxsAiZGcMJCF4KDStJ6x4qC
P1LE4NnlP06jOyotnRa+Sx5+cqP6y2a9TyPrfE+7CVyPm/TyuQoMiUkz4um3032l+ZNmT9HWS55x
Yv5JQF+hvl/pMZd/GIZ88y90z8E6b2bFjjhUTeDEMLKcYvr00Rk1TaRbcsR6ikaPOXg2xHTiSIuI
CS+GcjGFYXAY+A/Mf2MG6wBspg1hZLZAHZ2PcZADM2GU13TylUPTc7Lmrm8e34Ozs4t7XP8H4K6J
1OctY4wbZfW6rKLAA1COBlu5ttdYwMANXpP4VqFiRpkcfsSHwRsk/dg4T931ualW70dXis6fzhwU
huT8x1lPxoP9oSfc7csRRJ7xFHYnSEWfh0JIEeTpJ9WOrnuEnEXuLpm8ka4rqajbShE1U1oUti9b
iKsdzUk/ldIBrxhYj5qmGDhhfsFpUngqneGkVZlEXGlQvz0hLZkwy+9Te1wlL3YebHHXS+0oX4TP
wHsCJSG9lF5zBzSfzirBkhG6zN/011Sf/E/xgaAeopNg/Bj6rDCEGWfQ8pZblKFPUBT8V4M10jpo
8/Xzv26F7mmU71J6n8MyfQM5XCTuzxlWE+atct1nGT+xwK2Do31bt8k1UvHMC+pHqmZKqHWLdpWY
4xBDzHKPGzikdQYXInaPgtEdQh0h/6DYhJW1Fy3B/D+RXl2ZpQfh5tn9UA1jHygPeQUSnBcaD23g
2gkVskwlpl18/rn0MbIe2KM3IjxI9Yj2NsizeiLyvVlpIUA9V4KXwwZkeBjuVQBcg7wSs4v+aCAL
yyYt9E4fkGSVrCEJuXrHQ+91a8jILjVHJET86l4ue0cQI3MfgV5BivEvWD0V4tDrKWZ4KdDzKMhK
5qrr1OtKlGp/m0xJLA9hkBW4fpG0KSppRueX5Ax5gMnTrcoM4UHVfncp/tV9AQOh8FQ7kBihxC4y
7WGX4jZOHxJjeiMboLkb0RlDZbfqAQ6T4OmSfHV2y2smdievyijKSHrD1M3AI8XVfmc7aTP/MuQ7
8LtFcp3W3pYUjets7BJKE3aMVimsJ9hXHK2uK9FJ5o1pMKJihBafo9+A784fHzXs3E7g1k355mhu
iTE59Mlvltq+P5Q09+X+IsP88XWPoYwUCSpT9U7QDSELt6Ms9aARn4Cst6Km447B5NgSIO1hVLOr
KyyNm0Z4Uc0TK2GZCbypO6II+p/ufp/ePlzom2yRivU8raCxlnrdeMZ6B1TUfDBlweEB7a9xFna/
IsjrgGD7XM+GWRQKkxiBfWC0U+TlmbL1owHkMW8Qtq2zGENpLfeyZLqnOJm8iLEL4riP28E1tWUR
YnPyYu6vAKQTQTL89xoiiqQR7TBeOknb9lvbEDp77bJr4lXlm1kAFF8Z2lolrl6R2g1Xkc3uPY/l
RAk82sWQ1Dteu1XlCGXYtbkPJ5/5xT+MQ9JNMmyXn/yxJDAbB3rPi17zsaEHru+FIv0wp2D5OWo+
Z5EsJMbaNh/41noQngrG/Cp95JmMXR/PQWK90JkGQzOTVbYJ4YJ459aXOdPfv3q9BiIAEc1KwA10
zF4HGp9Dp6FrTQ2N84C8T5EwPwUZv9kxGI+hfGySHFQztiXRi3y9ILJtoYRz4eIEGdOkSV31tq+m
ODDpNmSV6XJa2/nVg6jhsqhP6zZVKYFaK++CP8Lil+oJcepMj8KvmV4TdO3XDQCfVLvBLa4ERkVC
qYjisKhZOp4etqoaCU98W5z6ow0qlz/rhgpGyl1Pfew6WS/bywRZfOBs6rf+i2zEwlO78Gb1Gnv3
0VEpkO8F54WXsHV8wgkgpYBZ8hz99Lyc8MYGp6NPKWa074tO21r0pFXadf7fSVtvB11Q3Ssj2DiN
i/eozsERXk3e9QPy8B+F6LAPwuR3QGX05S+ENlANwrTWGsuS9CfGdXmgLbogb2K0A4mEPsMZdy7s
DT7/vLtfpMh4u7P3ChFCrIx1dihIQuUaWpaWlra4QWS+ZEQYxWRrndyJsG97I6lomluD1ht3Vzu/
j1fNWRGvLvcCkmRT+OcYObnUeJOkKVb4bU2QUfvsXFurC/212WCRGSF37ghqYGFR4IyiixlIgiXQ
FXezM1SpDN2gL1+kRN9xbNX5kqjA3fcA5kVb5JthOS79ZN4FLascBY+rNHS47AFq9fXPx/OoTjBN
ymiB0M1akXqBzsGNtKA8j0k+PXAE9ATJqiwmsilNrRAxVnr6p5I+tuQNfFg7j5lubEr/BXI21O0x
RwmQKqwih5QC+K3jwHAQbo1mvaanl6icuYQRGzG1tFiilkhQh87IsJ6rXYSIwWgObeduEKN7n7aA
tuPEXQBEGsY3CEEkqjgGuj3zQ6thsjm50RkJXio6lWHCOPVzXJDX8olFx7mGpUJsic7OxUKOtOqy
IQQj58RDu04hJKhhERbKSZkSzlYKIJseBzSe1oY6wDHpTVhL2dNfu0rBZreFb2O+1fM/84y6ZrhG
65p47gMmg9Qr4ke0njmFZlv9cssjHZHfKKtloiptULdC4U5ENgK6ih4iPQj5ulFvWdCsLkmYzMsB
xhV+lEgqMY6sSi7fULJM/bKdpbupKB4cmEZvAITHmtu8uyYOI0UWuswqWjDIew+WYBMaDrgBSCbz
Cx1OA8HOz8QZChkFwzjFzXG8p6L/+Y+ymxVL/FCLpD0HdbRCV+Ybk3OlfAdFc4r7tU4C6YJFhtN5
v9OXuGLEuwqaU+ACC4yk/bv2J0zwj5M886BB2iA9Z7OGVgzC7UjBp3WRGbJlk9A/bnvUY6B/Z+nE
b+y+y0uOVa9xcDxAt6N0TEWmeqfQrzPF0GT/OBKzvF5BY6efAisriOQ2DrRFSR4VUtutKsedwndA
kjVdht9mReKAClGqZlCOdsDD6c5dy3Y9mENsi9aUgJDReIm9nTbKY7QVAu6EylBGTAXxNespGMYd
iJJnjABYF2/5Hvc9G6zunZhei7H8ygpdsTtMsSVihHVT2VNzGnw9tWVdG7EZqo4Z06TIekDivtuG
Su6z+6t1nm83yb++0pzBFnx3yaXox/LzD5ZyVYywsz/FP318WvME61ay80ZjvbNsqbK1puc587zo
WmZ7/n2vWOnkpf0YYq6ZcDRyl6gdjaMq7YMcWSsGn9/j8EP0P+gHKV1TiENF6RcbfVBsJpLD0qDR
03W4dpmFv6QyZMyuHxSFkDk02dS3wLkR2Ll9vo42aVqtfWaPmu2KlH2Fpj0tLEngMQLE92C5S751
KtIFRj+S+b+YCynEFYQFoysEsTLcGJiYNClTXCtlHEBDuSfKoMgYdzEBmLZLobmQBzCyoqRpCyPI
5rR4IIA+TArE9qGGTfK0VsZjMt1TdGmbzBPZ9Gd82BL80dz+etVe9Hx0R6UNZtVZpqVfauu+b1Yx
WYU8q6IouLtyNhN11a39JB+RqUFGdNW6ORr9zN5PSbrmX744jotyxsHjugpGhl8s2wbqa8IhlPTW
aEISB4NF9mBwLgdUnnY658amKENU2YvXVaJZ2BCOXvsq0BoGcgkw0fskOV562D4s1LMPAXkaijvY
T4vk2cNtKHtTUBhlxBWqKkCEcyw/Z7oVn8YK7rCdwEsORFWSzXt0yHSp0Hxu9JDHcslc++g8SFGw
JN6CIZQ62/Shyw+hU0FVPBrY9aHk9Lj4Niqyqi2g1GK8D7PMR0Pfbmb3X+8efouuQmfFq3+kIHyn
HalseQNN6PvffxHtflN8P7sQYq+6p5X8at7NGbglya4haDbQ8gNBJ2Nsxlbcd5vPvg8Q3EKa1lc0
2TVFD0LqoeRfBer97kawQao/eq6jMRTBbyPD1/KCzRmGlt4pQihamTHPgR/6UZLUvVEYFf/+0yEL
OStminGYgXGf//x8XeTiTb+EXh2eR8V+KECizmTfJOCqVlFL3LGr5sM/6G4jlqx8Hz0CR/HIzXq1
JBChMvIXVTVhOjZFzVc5MKEuSmOUfhQgakZAIOmbInMnTVc5MHywTMzEqmFUihNd6SRTTRsFo3uT
Wi1MdoYAsy7IZx+qaf0CK+JC5qtngL9zfuUYmwaMAtzlCBa+ibbbsZQgkOy9Z5mNhrnOScJlXyv9
46Y7C4GYJ4aNJ0oQHT7sLBknu6NsFLRMi898P9Bai6YEAcyha+8fNrR2C1J9bis7JwdvZ7D9Whi0
82DGpTgf6C6OgJFJkemndhxySE0YABvaiF1sbMVSKAmArAFqOyWuKUxUVHZNc7HnYjnw9Xhuj4Yn
pp79xO5foD5pjh2dabCTKrQ9+Wq8uxXthPUxEUJ8pdjb8BqeA1wvH9qGwtaJ9DPlTWBKHMBlc8YK
MzsuGV7lcueBsy3mmSvfUrQewW3t105H4hsRcbcsX/wXiA+ODLp8uEDjwRowZJTtDbHs/E81lRrl
bzcs/sstagZU/DgDB7eSoiONU9x/o0vGzcrcOburV9ppo7IVsiCX4NPNBrOY0gMTmUJ0xLPUIwTA
RqXSoyJbPfHSne/D0qo4t2AQ/NiHP+Cc1829tSu7Iy/pAfuQ8fVYV10h5DNcMY1gyO1noXPtMIFq
DAmrKrMJuc1l98BVxR9mL3fSAaeS3f16UmWcGew22dcaBurTcCupD72Tyy184ZRC+MVIgxuqB/Gh
nksMi+qnESgvim33q+oK6GUGilYQoZkUs8Pmqvzcn5kgpZaq8OGrggfUqez8o9XGoa2T+7u10r9E
TJpiULM43KOPVZmA7C5Czp+f8C8wag7ooEm0OBCKUJdUwM5b/Zh6VUpEW9mgMhA3MVf5JIdJqbKY
hXVTkDcHRL5dciLuKphuKm2CurbQKUXhE8N0wtQ4RLziQSRGgQFbpfL0MDMZk2SkG+0WHdDBDtsO
dbQUJacRDf/tzAnlD+t6nQMPea8doHN8Jc+M0mqd4vwa+6kjOos92nvB+48qHPSKb2GiPIvI/d2V
IUa2R1TfGRQE8S/qANzcxAZp2uJjv+zv9duM6ZnYqk25nl3XqtGZViKFlRfDXf8LmPX0s202Tmso
OzEDae+jW9KOmB/5xdr8VFfA65bKV9ymOuLJGI0nzcs2empT613n/FJEG2vQN03gsZB01vyEQYdS
00I0Xyx8eLvd+uiQP+iTxzGhDgFGtslCXBOXgxvqJrfiG9X3YdjAGm7rVH8uXTRaeIrSdJD1Dnz6
cg/BY3xXdcZp3jKRtMfxXIf6vwVW+6dRGCd1d2M7NWEWkWbzosUvRBqld5PgJQtY+xi7tl4yKYEq
jR9D2DAw6P551e1vwE1KUCanqLLUcvB7cCwob9cKD80Zkvoie3MZKBO8vMXlay2HyMhqFNJupOui
aiQxwty/wmDbeGXiid5LzouiTO5EVbiGtxSe7zVM5qh8GWrLZZB/furANkTxmtLKCsSRU4M+C8sJ
pfAsvEDwsp85xp+TotOjhi5TEe0DOuK3hpk72vQm2WN/bdwJGpQMc2qWKr8lBdTYcRSAhtzgfTru
ByeZUyAVLf1bNeub8VZPFFMDTX6Dub7ufI+ElpI5rHALX03ndIm5pLJ8KZmS37pmJdj+mjK11YCF
/pSkacamhvkCwluJUHvwjR05aeAJZndPSagV1Lr8u7FbQr8i90kZdMqIN8OstjJSTtTSJfZpkjjF
CZG96zOBbglyLY4MSmVY4n9WcudZDuXJi3jvzIHiOWPCvTA7sz8CxgXmJW13P0zmDc/LsGKrMnUD
uCDOk35RIVVge5qvNWGhOgbROY6XbQ5MAFLC5Lllms3whY7UaYG0/BIyxF9FU3pt8l/oR/WgLxZE
l/1CHwFVL/z1IAGAoIaZNbK2HqbRygohnO3RZoSgYkTQzV/SLLwn2FXelrJ3jLr/l8+KO1ogbsWm
m8V3lasBHTcxJ8QYEKG5kW8niy4tu3SRIXPHya/hrJPCev9uVMxeWCZzVri8X4BUHqjrdBojdgao
EA30TxR0eFIJ8kTK+xPPJ2Kv8xRLxLMjfi25rUPNLG+gY38fyg/bqV70Rt5e02efLKPrQteUg8Gy
NqegP/6m8ikeeH6f3mYbfvRIRzM5L1NZPpbOBja2CNbEwdNFBN6dfVJjL/JUPtxd4Tk90KTmcuKt
hoOiEFyCGYZp2naPJTi6WsSyv58g0aeOtWhqrAnr2K4cs+Pag6WcV1lakA30kx24YbwH5SHlZbuE
aI8kjmCjEJLO5WLvqEl7vkixJT1Ts2u5K5nJ8ETuU2x4EQi4fcN+4yHUqM3mSRH+omiKpZNkcRM4
rWJXJnFM0fgFOLdzidLU/Wb23BKiu5DtXXiHMzi0Wp9pdbnsYqUX0DggSNoTdlzTp3+x51XfidBQ
i2LMmo02XPsanwTQB/9TDKdrHxKkvpca6jsSsLhOFMSkd/PE4FCTOhH7KrE7nHQqi8ZHxQKJPVR/
93tR/nuh5I1GlB2N4D9/3GBKJ1YeQnNyCAI2R9EZhyn4Ri6ZPlb1alKMPkd3/x5edUFQw6h64+yK
U7s1XOABWjBDcN+peJN6DQRDtdMAeaIrWGBf61q2iSePIBgTpMYXI8AQ5JsqqAj8LarR8Urv9D1F
iB5LdbCmv3s01vl4NN2o2FQO6kExEOgtLAJsSBSBzGKlBSmjX1FDHiXPdGBO3QLj7bTo+hXYbR+P
7JP6FWGud7ss/q19COxv2ulaUQS3qLW6fh2TA/XtgGUgmxJuQ82973sKRqnfDu6+HWBLkVBuUnbX
FbL4nWVblmBR1q7PIK7OM8gzNmNjB19LyJUju6+PWCrXe7uvAboLLYLvdcr3EYHTcsDMBO3Q3Fb2
oES42uNYWza4RQBuF9ACzukLz/PZ3E6USWB5OerQhGXy39ex5Aoe1aoe3cm0BHIWZEv5SmT8CmRA
+D0MoczyMTgtpmBKUBMK4iBHRaCOWlLY+chhaRnUz+diAm6TKTHB9ovtKXdW+qZGsFCwW44Q38Kq
yLoalCovSk3l0MihZVPW8Wz0XD74c1arQCF2CgXSqW/sZdO7XnFQkrpY1C1kuOp7ayo9k3vmAIxn
hEmaGqkvR/zaero6DjYkoSJK9ODI9PrGtCWNlCoUnj0zmAPE2WLeTFwv7Fguz60b7l0gG/sZz7dp
ehWbmMGU4boioBXQToQZd9hbI2St64dU+MTQOYciFLrd3bAgerqIdHEAWpXub4JWFwhcQY9RfVR0
6fQ5fGCML239AS5s1QGb/ifSqJ9N3N+23MdPqp1HXlD0ftOi3MUjmTl9BWpJp8Y6/H9+Nvty+kqF
TpPe4Ca/bViZEddebtTTMOYqgFKTuybWhTfqJW99x/7igBGl0wrzohaBjkhc3zqPdAeKyojGWiUg
lD9y4ynAMxw6QNs4SGEiFz+N9ayr4vLgoSFW/tQTfmEJsbgr60zYTPOIE/Jb243uwm5FYwrlUFRU
mfkg6o7fIBhJYaBWlgMH71tDiVMLMQT7ZhRCytuHpH0mbEkkf4CIqJ+LObErlNuwYi9kDqXliQXp
91okzBZfc0T0QLQTmm60tL86klTqoTVLbPrP49dDPb2ze5c13Yhjqa4X9g91XnGNLoW+FxlqBoPu
Xn1rX0S7nuXkKJ/79hk4hu5fQmkwzhmlrmdI0eJ1+59XcoZGGH32658i/UNHg2W60N5fBHcwnlZ7
K+5CU3nfY2cwrWUNMI2G49Rn6dw5S6KQhqu7Te6DVdNjX7a980GqJ3xHpmMIEdNGq/olLMxar5w0
zACvYh0MbBcFjo4oZWhmtc8ErLjXcH9UCx8+DOuuB/Nzk9iLv5V/yRXw2TTfdG5iqAEep8rFbIST
CL2cxx5Ctpd64unjB7+v5XyymiYd3KA/XoLspZBrAuYpJ+dsKpOgKrcZnNpiccJuXVnZ3SWTUWI9
iGJojbLXpLnNxAu/XwUpt0gO586xKeRLFaL5C7aD6KrUCpVQ1AkDaW89e2TXm/lQAd4xH1l6cTRR
fBKHe5jZrp42ELPam4IFIb9nILZLtnIiBxe7YxpXJakcKhTDjDGK1JfJl2iWHPqtUmB84Ivu0Lo6
fqT4spvJaXQmnllg6vKqGSKRhbe0p4sw/HIPCiOWIl28hVwM7npB9tNAHBZtR48v02F5wgvFaLKt
8xU/5l6/3LFaYkzQHOuaB6FYzW7yLdB+6VtEb3Ebnh44ik02UZ5LCjXqPjSScy/1MCW98B5tsdWy
MXdN4YrZ/xrNI18nrl46ZoOKOIxS6XVRGiAg/R4enXZoqeuWHods10xSQyTxfxxH9sR23KORFEw1
wQ6PixrcYT21MSEzrHMOy1yMcExnXbPWOzzXPrgJbgyoI+VHC74iAvWUtPMVPTsPBo9a90RMCK6n
UfZNGCfoQbfh49EAiSgH7i6psk3iJlMhjsM+CVKA0xkGaLhaEzf0ZAXVTM4oPqC8FudKb4BQMONE
xd1pPx/CDwFwp9uXZ6EUlvX7bkdN4TsYNh+2F5ETeaZdUtjB+bT8Qe2vedl/3yKOG/S0lqoZIujV
InZMkuJJ+AIzg14ikvZwxaa3MS3wpibFJOtlOosdST3PDDhLmJvGsjbH3HTesX8aGfdSnw7c9alT
835u7cRA7dn+BGKFpmdms3kKOkXuP9vMtue9RlzVemL3LuEsrEQfWPYmiAIm8SG3V59Y9fG6v1ad
0sXBD++mWMQ00/xZiCQaels1+Uv+845MFoA3lq/oHaqpgfsD2XsxEEWLfMx1A6S7MpkZ9BQ5D1K2
aLWxldJr6yFuBz2scD+/zCtCHnXy8ScPCRi1pFQy9RDOCXlo6dUr0wCofGn4CwJRsJ7PwWmB57xB
BjQjhLcvhz8FmMbqhC70cWsMzdh1JdEWAhZeiTDBKq1rCcrh9KimbU4zhVRfnDvxR1D87VcHyGp7
nG9hoy6SYhZT3OBTRtGotxZ8/1ZSETsd3SYW0kuqEaXNkgISwVHpdtEbbZJoaKEck4fXGGLB/gA+
1A713Xaq8TFd79vT+jK7MWZsKge06g0VMRsFBW4r2+r+yTw8zhGNZUNTCb9XfLPVmH64H7Ce91UP
Jd8iurb6cBFtuKf1xPpUgD0qHARFuq8T1ZJwJzBWDVbqKo9dL2Ng/X7CgTqiUDdYHbo9fN8YvxbY
L7RACw+Dv8PQBBGfKdatbyXDF1NlrJx2gQVRWxcQieH9++/T4hhNyC4psnTkUDjgEO9kQJQR1+nG
UqKsHxvusP2nsfWwR8nXCQOMQGpolQHiX1xXqyG5neQMN42Qnv7tMUpLeTSadxqZBQgDDrQPS+L9
EaN3zD4uEM+ZZ7WBB/zNd6ERS/rAqAiSLAF58C+4P+XggteLBuRHoGNmFiRp3GEaJzF/37JApXvq
9QmCRe7wPh0QFq0waGV/8zHyU+VNO5COo95qu8I926gQIMv4UzJg87CBSu/AfKVGcMeX0WjSZalC
n/7rEf8DF+qSBauEqhBWHfqysYdTt52TP47RUP4xYu1M5ChdJazg2O2f91JX8vc+1FA7FDq5tGm2
FJNw3tEB1G3to4GOMePR5sFlI/r9rZzluEIKpZ1r4cy15ntYEFMfVGw6CQ8JtdDOQwNNuZv/K1NA
BIBCLQHfuuoF3A6UELee35SUf6f87rkzCcg1Av5Sm7yZhWe+i0054Jf9gDxZzAWlMAISHJs3sKcr
sZdSPA6tccrNp+1Z5vTL65V28RY3Ve2ODeY3TXnBxDbSuRMmo62qrX6YBXDj3Qxhvf02gU1Juocf
7sogoZrAXCr/PX0oAjYflm1DZBa9rTn9xZ4CLa9nwLnie5Wkrx20FQ/Vr3mQPIbEaEJoU70v+QSD
Z46e5RdAHK6LWsyHJ8UfXixTvz7zhNL4BlSRK1xHYc/J05irwCw5IfsektHys0434zPnYRRm4Z8N
5p9eFO5gqGWRzwwNFRw2HKKWT61swzwi+GWDMjar5JmG2TYRylTRJPJIh9QMO5apFvoRr1bf/X+Y
qM353OumxTlVv+x2a+EZgG6JqTbVz7kaIZsRqtAVHO0BkkTWZ/su5RiwiM08SuXOvs6+Es1IXt41
Bi5lRMqWN4XgA1hkdPWzNmiddC6SdXJ1GpOQT0nolw66zo3ki+GpDcAuLQhXvT6wKi0jmYaKvG0f
xruhQSlVkYTx3EWZubjVoWjanlFrWQluhvxkefBn4GLKKsE4fw/zb9c+JeWM5s3f4Wi6tnsYLBWI
PAJCVVERREmM00MB25JyIHq6zaClyxuXgg96kNEVG/+ZpMC+OezVFFEQO7cIQV3scn6jDYUKGhXm
83Ez+kJKBQhBSWZkjNrvfmBwmwNUFzIQA3my2uqtLwl0uza3mshS1Vi1EyYH/A477COC4hIZPEs1
09wmZ5lkHRkpDgYzplYpB4U8vUABuB9+dhmsbqA/xRxNKCDesKnODrPARNWmKDgaGf1oO+yOMr/8
l979FTqYHOhY/2CH4sqorg7spAnWWqquFZ7W9Wa26DKKpP/pPAm2xeyZ+QBdxhsx4itdhEe3Zqos
L0kEzgR6HCoksGJZYnekoiJlPXGKhzcLcGXBNP7CtEO/gUOZw6UDhH9RZ0usraWnuLjHOc7sCG8W
03GJTnlTmxAhqAfUJNaNpqTteFKYNAprfgpzwJYYGa4FpJBg3KriBe9YCxpf3WxPqOE8Lss7HQbO
MoSdmoD6UY+soBOiRW1K8qsIW4jTOKRr8yOOLY9BAsHJevNnbkQ/ux/554KO1QVvFsEfpblWySEs
p5dJS4VNnM4sJLG2wGXp4ujYX+3xR7m3+X9jaiO0C3jOyzWD98amD3+H4e7rwHE9Tu55ZzoBx5IW
rHWL6g2h3vc2Nkj400LkXJ7CzWEzZcXC7KSHeNaUHXfMUklTwreQZYZgmOddBq6qt5kLyQh4czA0
u/bxK8tIp4nRImKNdBgkdJGZ2EYIbyn+aLvT8ZAfy3XeJBzUMx77YNUxx6m1eCVhpz9iZfK3Oeta
fMegt9h2Mmg+pSHiHiuzlhf1OUivXLd4wm9v286+9+qrdLvNxe5r5dghpxYEuZIEQ6L4H44j30+I
F00R/QF9dzrOZJX8Us33gu6xKAcezeZkHxrGxmDQQfl4EfkL0kZDAYKxhAbQeZyJ5e7ExHizg+T9
PliQ+BfvjPQDu7Ff8xIvFUYpZhN8VAlInqapzc44xtJDvKtExIM2g445SwbD3Uiy/B40lsBUlKWQ
pjfNlQDmFp7tylVxSkrFhwrCIbOltsHbCjQqA/9uHZ5TCWOmBig2OUZpQ3+ACK9qJlvPOzamjG/I
QtZFFsJf2mLbkTGa6i0//mugYmk+1xcOQvh+N7SbUEabncKa0DcANMWPj1PadqeaQxUXXX1Cai8K
OPLdrCp0MYCZbmrQNfIoJeoAxqgsPX+ghsV8VmbYfY+QbrCQr+mrkBZEQyQdLGU+IPfEj/tU0kjc
cUd9wPOOOSD7BeWeWFDAPw9lFFIjmFkFLE7ghvn+7OPl7qvzm6akUDeQUWJJyq/sNHtZu50bBLeO
+P786KXohNIyzjPcCBBe6yTKuslFatYzXJvLDP5Qv3IIGiY30a70xJU/MvEhX7R2DpvyaNBTrxzt
aRewTmT1hVrEygMNKEH5f9x1Ve6IMROx0yGo/Zc5094FRmYBsqLF/UdNBEw2gWsuHC+wsERGD6JW
KSxxvYhVVvG0rbhUIj9jm9UIKloKC3MB0tAXm0j4hxcO2KIPEcBmF3Oaerpi/AZXmwad7DBqp1gz
VqbZS0a9OFFGs3nP/OOvxXDXNFaDyYswQ6FgUmoqSXjsF2/1z/G6krRRCa4nWLQfWd4xP5jXjTA1
dip5xhZL7gPMuC2s7KSR/QtKcL/Yj8t+oF+nRbFTC/Ah+G6A0wz6omqeqG8JiiWrhNKG832LxrxR
05xfrdgI68qkm9w8OBruVXmwszdy9ll/LQFr+7XiTDbdwUZhK/LSup2NKsZ8T83bXQSm+FtRERPB
qBSqUAcy/Y4VSf26m7Fr0QlTPvS38i1AYbWa1uCpETdg19grla3QmKu2F2vYrYqYvEMRk+H3x9gv
7U08qoVW5IYzWoiq+vSQOOuMH3jIqTjfYiTRs4GApBUCWav92OEoIYOW+Z8YomtDkDznvtXjlb+2
YwvMsPLRCdlvU9yq5a+yG8NWXvC3sklFlalyOxR2swwmloQWbnSYlzVwrON+K7rwM7zljgq6ZljI
9r90l4TxBkaoGbx9hzrradXOofLPsOZdgJL1Xx9SFLa/OV+X3Q6FKZD0PvyncYHlz9Sx0pPoZDpn
9xAMAb1KTxZzDIGF2QpSP7mlfQNhKvHdKRa8c9VW1i2LXdmEdBnGG7d7R4lsqge4sFjXAqC3wTfq
O5/CD+95GWEI9JsI4ru97NhtC/+m93V++NIoJeldljNZWQn4tS789bOvnmK8pZMsz/YsaszWyvdk
Cqtin/8D1MnitTHvrjgsnjQRtAq0zUyYjdAwu1ev6B73OqrvoZOnp18PVmXj6sFfiUMvAN/DogG7
E54c7SaTrvZ5RXGQpOz02RDoEW3M8yGvUTpQwBTj/OizkRqBJuTfrIs9tklxSGySCHEjoUAnfPkx
XnISyBOTmlkVHSwgI6k6HE4E9IZgdJ46wS5uEDU/a/RedEO7sbsjXs67+0pJT99TUBNww/+Fvbpe
ZGtQDJNax1O3xP/lc05XQuFHK708R7q78QcRwZeJdap5QrOwzS+PHmhbPQJoeHiz36wjZNWcvCJ+
+wuWubD3HiPxhiBiFobLoNyPj4yNKJ61EYSWsyrfoF2OvqToDYWbjwDcuSSbzqUZUK0VgCv790Yu
a9JYv8Y4Zg7Vqp8u6g+NS0n4r9R1RxhWh1gnAA9G8xVDif/7lkywzu4xFGJxjixeIX7XoJGk6ujt
WVpG7p8vwLkiCkv9sTL53iTGN4KRNsUnKLfV3sQ0aCQJE9jcG1ty1ccuhe5ciHzRzXxhI9m/4CH2
cKl7X4CLjhxfVGYrgK3j9EVPsJG+kfL3c9Ile6f/wTksXR90OrJeQL/jba4E6C/0mPmdMMfgIYZW
FAWJ8JZLpn895L8bA1MneVMm6kg9r71DzooQokHOeMGQUPYlJh4iSCw5gEOgFj6XTtnrQ2QFMhj+
CDXMRujykMjILBsXrG//LKRTH4/+sNHm0PrxE4ZmDfpfUD2POkt5J2rvmvi/CDCV/VyW6eKCZE4+
inyxuwT8aHTD+f3ac6CL35HoUVtFykIBO4gh67OTgSXhSdH2wt+6SK1oJ1dK0MZzyLfm4z9vJmG0
OSXAH6n2dXh0QPTMtj/Ygc1SnsURN3rA3SHrygDvWSAWBGebkTnduCal3df4wwxQHXD59uXq+HPE
LtB4zxyzDEE4dDYIm88gDU5sQqYE0Pkd5/jA2nIO9BXxGSJjhKHe4vy9xG9fCIjnGOMoTmr2XSNu
L/CX+FDvdwlAzOz2NlaDbgVGMEGqp25PMu5g71k+1AvYgvV0PLLLy8oGShjfuUyGRCUPNwI1H/id
j2gcgYxWMNWCgHNNEUTU83og5yqYyUcQOkPldrdGfPnAsxjUc0098/KYMnmc+iiQJU467YaM/7CI
Xfz4/o/FBwTEmaB2xTTtgKxfywHTL8XzVzKT6cTw+gm41+vr8aLO2HQqYl2TDbY69A4/04Q/If50
gQDmCZmo/xirWn3AVw7TEa26qAnMSP6KmIu6cRp4DXH76dLGJg27Qd4IL/YEjHBKPGAvTeM3eS1Q
ba3u7340EjPfZKhl0dbKNTmEXfZp66JycxQlR34p1juHEu0rX7M3H12dIUCkHas3DzK0eEjea66e
Djk/clT/p0mH1dOj+O9i1pbVOjsjDPn7a5m8JW99YcFyBPVE/UqFQp1dNG17GVZsh638r29QEFj7
Y1kuU5XEMrIe4TQYkFGshw2s1SCe0Id36e7xv2rD3Nt5gSOZihRemPp3Ocqfam0krGnDMfRf8hSK
7Np/6OJ2RrcSS1r8rxK3gE/EUsd89MEIpNuoxhYxtyGoLdUO0lvbAx1VLl1pVee8TTrgnURCzK+u
tw2oe/6fBpm3fcppLQvVV940s0bAICzRpsVfps86QIE9u9Etx1aMqhNpDAGJ+NG2Iyo7t2ij2jsJ
GmQWhOY+rhjqxgBozCCWFNmTSDtLLIp5RDVyeUDXOs/C3g9L5DNROwuiaOgBU5hwFa1/fjBY1823
Fthj+uEFauPrEpYJyYYQMvA9c0sVs8SunsSmVFeBWb2B4Lsgb0ZYn8KFddri49Dpghcw6Cx8gJff
HZzG7Z8WDe/fjeB7RKZ1Smgww9BHiOlvksUA1nd6C/tjG3Youz8QJ33gBufQIDSUTFjXOUXBN3/+
/fPYVEv0373uVsdEJOwu/sCRXMJ3o55oEnak3h+9788st+opKJfb+73Lxi6PsigD/FAcVsBeAs+2
ys0bGxluMP+MyRZeri49/9o05ai0cjmmY6iQKbvHYVUWMBzMdR+3322jVJ92JeMs4Oa5AK9mlrRp
ir2gOzIM1hadisk/72mI8VvqjFC4Dlnrj1o6g/G5bw+GSRU8JQmYMWHC81CzwuLtBB5jB3RyFqfU
nxojr+fPLcgqx5YQPCHOSE3AMHr9EqcwYtme2TEEAOofFr7rI6gnzLcu5cflGSV/V14iUEnru586
76a+D7s3YOnPKfwab6jTNPs1uCLnXKTfEGtTTBHp5vMEf+5JnC9961fvf1DqsMDh3y6YI6K+pj1r
mI0JOwh0QE85obTYKLL607ahbtwUOoKzJPzSV/8aK12Jhz0oHEPJPeBW37bSCu6nCBFVeMDmlwcc
v5vKvXPlCmKxC9Vc3idDkDYUS00sR4pgnWH8vJdq1TXMSbDQpjmxIrDVHQiVQ9MWkVTVedCCx02D
Fm+MFgBMpij418OOO8ONGOCSFK90uEYgXWp46jYxYdfDHIwB3+9sR3Xnyer/gbriHheW0g3dfp1n
b3/y7E64NsobjxMUr4e+OQ4fR2PX/n14MS5o/Q0IZujD7PXrA2Z+a2M1hyWHhN9MNDs9YsLACLaJ
nRWInyvCndnwry4Q8Pr3NYH83Ou4Q5mpjg13A70NrVxQMWzn7AYmohBcnnKu2xzFHFedHkax5c7P
eZxFFAAXAREwUJVUBDYvPtU1Kj4p1777xU2ZqLALntQgvL/wZKmJQnv0vozWMpGf6MLcZ6CkDQxE
+KgD+VAjoyuP8ssEc6Oi2oyWEXOYyYEc9gSrQe6gTOApwmfT8bKMbgEDiCjX2oZXX9lqd8sj+68k
v/ENX8jc3ftHF7FhFDB4NUUczCVPE6gpp3gW82hOhI9/zC/ES9RJimYsZeOEhSAWJdWJmbC5KQ8X
ZdtgWrtFpQGvg0vrx+MjZV2UBa/5qruED3cqLsmphgTr30CFR9cWKfUlgCxnmP/xdW7SX2ipDlru
5xvb2aHLrXWA1/SwLdfVrn1mWxmClMnW9pHs3JdW1NK/+yz13cBpw/Q3aRZ+tRHP3/1gg22KKa/R
r3mfmwhdptrUI28nXxyvjvLOUvY6ACGCXp36Zu1Rf+JGjauQ+LcEUsXWsJ/EiN75QMrDcgNLLSvE
J6aIiqerP5KN+KJwh9cgs77J/YgSvgngXPny4ehg6clIHF7/3+JGyN2rluQ8cNUxxgKwB9eitOrh
USIErbswQh4+I0S1GlJ/VN35TOB1CKBp0tA/p2RE6l4x3m3J6aJ9SlNDv3N+oCB3cr2VZInM+Ctf
/pG1AoZ8tsb2yJnoDt6y8Z415X8hL/ebL5BrlbP1L22ST0Yuxk+EcvlinM/6MZv+Agm35bvC858P
G8ENwIXdQXinKRYb3yxZSOy41FYUq8jjAyxgywizBExUH57PvbT8nPa/7yDPMOIzciRl8iTv8T4V
a/LSP9DPMb8l3hZUAAJ2xAMYqXKIKimRCJW6ftVUr7poL096ghLaT+eGCt7Kp69q8FHCyrnxtZ0/
Qepix7e66bRGinbjkEzEeAPNp0Khd4bH7l4LKQg6Ynl5D1g2dQ3NuPAYr5sUo6A203V93KXDWjpX
KFGhr3hT0h89tV3f1zRlR1XSEb6GO83LkGrBnbIj6BvkfbORbZ6PQJ18Mnfp5MrFyYoKouiAOUcR
rCicKhnGekUaWf3vVl7fdy9+AxPAQw2yq4ZGuxkSswTCuTgy7TvZETq9AiqVNhkRVScHr3lTrZ0z
TIgQKp6k4Qh8cUFJTZDlDHUV2dbE+aciKcOWb4CWQyV3Nc24Xf8oCe2gtM3TqjFcp4Bauyipb/9e
yjdzKocVuopEUUHFbZupMlGN49FUhrN5FHqI8NkoA/O2+NMuwqNVebHZhr3vZ7Pd3MwdiVi35xRA
FOUNrQ1Lx0kNmrNmrobNXRHQxVehB/GFBn33v6XZIdW7QDvb+6mihOb4f1h26ABjtFEC7igU27qG
CxqL+4+QNgmkx9D5ImQ+8BopRPXXk47bQfllYiKSo1eBFqxGDrbCxruI5PtFo8zunF7O7hVw6uNh
8Av+1gxa/x/2ea0ozuoo9G+EHAz4EBVvOHnY2WS+zpZRLLIdZhCcbv3rIY7EgEL04XwEGCxEL2ZB
5JYASuYGM/tS9i+KBcp2qDbzXUU4TvVI3NTWtFTi3Ct4u0qJgIQ924JsgqStavO/NnWHf0VFK1fd
HGiucIcWalms0lmfEhJ+R4Nr83pOzxIFiobdBgydDneGcqYPzQgZpa+VB0ljfNCZia6L9U4+q5v7
9SF39ZcnO/gMMPh0hfiZyFbsZdWunsjeWtIh+e3gGg+SQYs1XCM4EPgYJBtqJkc5MdjQHt1TX0GJ
4uqj4fbT7bSSYLmZZiCQqoEoGuejhnVCMVZxqhEg5GHtUISYZa3V6rqFLWQF4NZacoiEAlK/HDPy
XEg6S4OxaAJEZVrNDFrgSs/GNx74U9x0tYy8lD2zuOqQrA0qEyyr9Kjhed29o3mSqVU19+L39MEr
WCCd/Qp2y9Ug0WvmHlb1mz+4gN3wlzYfuJO96/+WNE0+415jPHp7N7U1+OgJEMgDoBtTT5U6oha3
45gVq4KMKIDkzNv3kgWESt1MMQbJ+kCG73yyjdhbp0FNbfenAY5rIUPr3sv7J0hF3lGSU3O81eY5
FiL4/snC8knoZGTatvmkxiGU5xynbwE/VPDcDLl1trBfE4EbvUi1exHnKsIl8UJaRm7JrujLJ2uL
aw/DVpDCvEkLtMovF4IS4S4SKRRL8vQJcIc4ewi4M1piIZco8Yo2t8x1+VedUBwvBp83uK9lUchb
GWu0Djkt+N0KemcOX9nVKqut9gxienjihqdSMRkpM9CFWFdjfE2lBLmycOuYPPMCTpulrKKYrzyz
/wMp4gjFAm0BxJTHipO62AzVtw7Yxdnh6g9QfZb9IyVY3B3yiKvCmmiN3gFeNExdVHb2BTAhuVV8
TWcgfuLXkEdqCtv+g+xi3oEQDxT2kBj9TrH9n6wcRotFEfvAQdGh1bDZwwjHyfpIy6uDdrqMtnA7
c/RGWNN7psWaj30BFD4Eg4uXDUwmaDxyfmacEFlZF1dlGjLAzAqiWSegnX0ImauOFGnp5YMbQjXA
Ix5Jr+itSvEs7QTRaiseHAZGXD0UscbtnXQVF7YfzdH8kJWFs2Rhb+3HJP6MQ0zcxRnViFsTR0bT
xLrNKg+o4upGfQGBQ/xOGMpU2PDDtozZExo0zu1z6IM/+KGUvFP8a9PSTPVm6pErxLNrrftptDlP
0fA6vYUEMD4a9CI5BZslARD6nEVBYwxekLmp00NQ0BxYSokxe4Y/kr9oxlDzUE6xrhSRCekqnTrf
xNSCbM0rSzULaRTkynEX+PvbsE1HiTeb+k+W94tSVaxbcW/hLlfTBS7Kk2gzxUmtukFHQgl4QeGU
aNsDOefJq/D+si4/ibiHif3Z9rMSSOIZrkKGibE+KYSCQvZopnjkLQE4+5rizylLaP4pds5Si6vg
YzLE+naYo6COCoxkzwEZ8xtVXdIffD4f4sn5ZYXzxhtO4pRfD3c/t/JCqBXzBRnOm9qBciBKdTyA
jrMkWVlArSV5mLSYH7iwSwqtY2dSyV1BrI2kdYDTeTIms3FaMyVs8Jcq2SNOdIeNNzx7+P5eS9GZ
4SeM5gWAKmtmH9wY0uZXQQgd93cszo1TJzFgRdBZWLcr06KC0h7sb/4K8Zb7noIZqMRS+qGQHB+6
hwGbWAX12spYDL+6PC+SyB0IfJEf+g93DmEUmcZI39Dd6lMqbLUsX2Zx8Y4fNXazdtR7l6n9NJbX
v1Aa27Kb1VXmsJ/MML864abgkfIKE36bKkf5n0JeCzlUCDY1xdbWZitdUX8q0PILgt6WnrewybDp
//E0kEfPiuaCq7M6AxJNN/l03UN6Wt/pGl+3bjm7nhGBjgUyf6+aNyIhF4kGR7X2zfXxG/XoRNcl
zfZ34iFOTct1mcLeYEN9ola9IBnuFGqr0xbf3pJYAXKvAKN6vUhfETIO8WzOseC32j7xI66qP9Vt
WccCxTuaB1G/u78RD8Z39HDGS791a6ATw0el2DwiJkFX9tP2Y0ocUWLtsqbcFecB1grQlBBAAZ/a
yjl/VatWCwXmqDqiq+nDwRfoH9fQsIZy0st5Wa8koxp7dDFONfH1AuO6MFY58Gtu191FWJ0WwTo7
v3xaA7gLArpuEJC39vwWMZKmZc37HnkmOclCzBAQHeDktX0GmsMxseL8hadjKAocUq6Cfy4uXbjN
DiSYmQCpE+aYtF7xZ0BJRJOiaUMed4N6CiPioh8A5BcSbjldeXyMq4Q2uVG/qEXgrIQ6wWyopgB3
ihOi3l5J7wJ6HvXNJByvCyq2kLu3BX2D1bxpuIgFODAkgjIL+Yp2Xs74gnCjORBOtgUPq0QU4SoT
+M0byN5FourdkNON/utm+x2bJD1q0/nR1y2Y2S3PYOk/wZXLGXbPx5I7M7MVecoEktfn0qrg1+/k
IZcpfWeLfOHfx2aH54GUSHpQR22Wf1fI8M085jh3iiOmhEgeqbxSiHrIN7L/FM9rucrdL0ZfdAIC
4NA/SYgM8VSaC92PttsaZTVhTXGWnEJ7kKUgpkdTDlf3oLMXH/8f7ncvGMcZlbqyZgpHA5WZtxdX
Bcofl5D3JDHRfiVAiKgAhbwzPMpRtOV0vVGaCW8eKV8f0iku4mMHid6jvpNMXaZ/KbSvSTrs4a4B
kynrrjh7Le8gl7f/HseD+eRlmuwUeTyfBSW+K0JcnI3meDA23mWAungVe7dN1qLTCBXltbcZT7km
RRoz2n6rkdjpftuhoQs/frEhZbCcPUh3g2xv7DJJrPfKnZv/HGDUIEE/4C8JRYVAMvNWVc6+wVLv
0ZXQ0cyGdXsrMY+MoJo6Qd6OKsmca/0AOgQpHeAxODYk0SnRAHlUugwevFHvLgi4UTDg0U4P3op2
QzyPgtpDivED+yMBTpepVdyegLdFYD0iYsnxkiq/FDxldku0BznX/rRjo7dcqrkkx3trnjhbEwpy
aPtPgDDK+DhSXqWx3Do1BFmVew+nYkAiwwnpwNmRXqM3MUgu7bpYAzjbxJT+LREYvb5vBIYJAXmX
L8v7FPuOvNn9X3k0dewmr+wz8uVDwlt7ggmBYpYqW+Lx6mOnXJcSojTQieBSjMTe0kvObMvr7cqL
ZyiEUmPv1JnRzhvZwXJos2iWsrVWXnyWmuKVUTnniH9COV4ZWARR94ElaBXfpzgQcSswaC6Xc2FC
k8jNjFDg4B6ZDGJPPlRyiddJQU9Q9PPCqhBDf3ewwfYq6dM7xllD+hyPZYz/pAGLt8sYP/8byGbb
5pRZlNZvlc2YNi/U7I/cqghEtQCiut97OpMY9/6cUK6+QyzwqkS5UoVAhSz3msDanj1VAaihZbVR
HRJRG6ItvqPDjMOivSOHcvqr6A2eUFQ45EZYHFy4jx9ydqPjuKbf+FYQsGz4JJU8CLeAE0wtahre
oVPH5rE8yjl1WvIeYUgjnDgpRuC/NJgDgXVAHFPfMHdQIU1hoEoHIrADW7cvmU7i7kWskGvydqVi
SO5YoyGQCJBzsdjtdn9QNgVGE+RzQBbIF5xASAFq+vVPVt5+QxmTi6sXA/AwBFLXJXE+fqjysWeL
io7f1inhYOOr+lvvzyqRjd93Wkj0s+3MmZ2aU8H4Ta3Gts0RRhOQrxWMnvio/yJY2bWMLzfCiwDZ
vh78sZg0Pl0qMV/iR4PMDGnE4P8VrWguB0jqbSxv7UA3nv1dFFgdx5U+YNb96ohrMkX7xZvvHS9E
z8f3KbJXUx1zMY6RZrC/z+6El8NVGPu4WQdPy57ddGGyzZGdTk401JFeRkJ8iY7V913TxN6i3guJ
eOX/ZMUiNorzq49naAMIOccmGXRvGC4udjHkbSmJtdVFSIw/lmlmYIa7UVJhE1h0IRmA3Dys+GJu
XR+jdL3mHJDwPBgBo0TfJrFNBjyvYnNmIchzQZ0rfiBqd0NRe1Brv366huBYvmaTJizLdoYVbbde
iY3ANxY+fA27LyArwNzogKRh5U0rwrlTHmm/mdpwVxnAjLwh5BzK1arBY32GHxCYYNZGilKc3B8J
4hZxI69IbN4NLXh0MmRFvNrkeUmx0hzNRM1vWHtE4DrHTco8+lo7qHlGK2vVJ/VImmz+vBr/gRZ4
EjIZCYL+AFCr2aRQDnVIwrnukOgsUPrhoQ/tu0KuAuqsOLNuh/shOqG0xCMXe5tlGF95xq1PncP8
llgrHRtdBRxNhz1pxk73aVI/aodY2PTTDiAafZa7l1V9TLpCi4sEAEKDc12zFElUALW0JPpzL1DE
KDqKeSmLch4KKk5Ts54x58KmYEuruyoe593CRRc9YjcC7X8Fer1THIYj5iLKb2awSZbyh59a5saq
bLsFPIUf8LqrmnyWP04Tf1N6Neqh6QswXFY9wQ+W2XxrV1G+oe4lzIa3rBLEl2DX7q58uIE8R26P
jcDG22NKNXtURBYihBnnGMScOuiB2MOiR4NvQkLg2tLRjRHqHZu7+38DPDp0ZD9XHOFnV0jSZ+Mx
hb7xv4VpKZFMeh1RI113iSdT0GGvZsZV0s1u02CvhxqIHNqfYDWlzpY+yVI/IJBi8enyh1LXMuuS
IZxR1nI8YaiWvkVRbA69mTMIhr5RzcYd3dSVWj8Lz1ouK3+KvG5sUZ3piBx9iNAWCdHInTpX6nfZ
05l/j46U4ELocezwTSJD9ioH2+TtgustggaaT2UC4envNxUqR4rLDClailY5xyZGtVPa5LAWW7tS
02cSLdZDtJJwGmu1+iOJGcm6IsfaqAqG8eEO0omojeYEw44uaX69h654/XNVa9tolZdI5RPmXb/M
V/NgtinvJkRBPwDk/KO/tXnucgfqmGRKnRDLa6z/4nYFcMp/1+fR7GKAfjXwK517Zw3pbkhCRIOF
jZLLMfWyRj53Z28CqzZ2WCzfIEsEYAfJVNQa/No/2sR0oOZEL5gxqS5k2G/+Mvdb76w5nju8vJ9t
u9bk3KPlgPbN5Rp+/RgFXy7nkyfp+4IjGf84MDvbZcK4o912SnJEYAVWAzpQ0MlVUiMmkiKlQ3Nb
mkxdPyCoEjmNeDkngav85QgAjmlconutFHdwemfoyhWo5GRjgf1pZc4bXlEa5v7aUTVY2jgM9CR3
rtURDkeWWOMOs9HpwT0HzKMn5IYeuGSSRJEiTvGtz+ddyE7FMRp3fB7/PWSCMKOFihOgrOeEpQS9
iCaX6g+/VCCPGN7TdyZ0HFE4aNtr8+0P0h4jA7Q4qZRwOskhOtnTLASlzgb4C+xsUUeWyCmXKdVp
xHvKFtV3rrxmLixxDhRFwhlpkSWBXhl+a8j/cReE1Rd2ZwA14mWMG/ikTXqkTa/1spZB6GXJ2ahl
wIOjf+l7zc5eLg91AWuNqYdXMNuk7LNKsmaSGJUIsJbdqGIFGf2ml8KmyA7SU2HPxXiI+OB0KqyT
mPy4KmL6hFiIWuWdrCktAkir1WyEJEQue6lwLp597zwJzMJQ7c1K33FL98bgFlBPr2rAabVpgmRu
iHafTWG2YKtrIKzv2nxIl7NCdIZj4Y+25ljqGmL06pr/YhuKeampT+IGHoczSZcm+yNTe0tXvPvR
6v1ghW8HLwSt4fpgCklUtFZDeITnytG0LiaQOYnJ/qpF+BIbFXIx9BcvTFK7CpA8A38wvIGqRFT7
bqS1EyynlEEvJwNIw57+ic25MRHv/oJt0yoWjWQluH6mQ3KFnF0cUIO23UX7eJbJS+MtLN4Tv+1S
hzTm6xYpzyM7D049u3FoJnXAYoWFvTRBJxL6gyKkBojE/1Xq4J0mt3DcPzrkmwL88Rakq2kictnV
yLYS0be0Fy8Kj8pySRDSJMcJsd/srrt8tIAhEUpzY4lfdwin4Qv8kxK5VEVM1GdghpxImUb0SWGQ
wupdCqO2QuSxihvDfc1teGn9irKJ0ktxBFlwYBfOlxtJCN8TvRjvvQ+gBFVguvUYw6OZwM9y43tG
haAWUI4nGD+0bewe1z4BpJbLVmQomW6MX8StJCeUYVB7a/27f8+VsaYtPAJfFFcJMya9IdqeK0UC
JdjK34jI2iqiVEpIStq5Tfh4Zg8Q49lRSjCNAZMwxpvEC9m7zt1c5aHLvFtY5edz04q/5PonXmH8
EZcpYYoxgMS8jFRbP8wzK2SbR/1th8TkaeUtsxwZMihcw0fROSyZMIPJ+7mvZle4caE09XOvJJ2D
z81dYw2FDX6KD5ROcs2sII8tRL23K8M42BPaBH9HbKira8e3zpxCQVjzYX6AkIfc1bz8iYitJXB+
Md/U3dm8wafysw/ZogEPYz5IE26o4cj9sAZ1l+iU6bjWl/ADmwAdB4cgn1vT1oWSnISsbVoLKTBQ
QOr+l7n/ubVWVFItg2sXLlHdoL546VLaRffNSiOFRk8JG3Ecb9tMDY9UBiVG9bvW/Eo5Xq7rrzl5
LT5vq+aaKoLNlkxoxFSo5UMgk3LHAGANMH2pOuLyzJEapb3ZiHgzqPStNDqIJiDh85qv+mSF1DMd
sxtLqDc6ETUeUXPWfExF2obKfCai0zVDZegnAkRbd5oDI+PRn1pCzEfJScRs1SAiHmAtlZBidOED
6kbB8RJxaWldm12WjAN50ppQ2At+nwlHXJ24V0Xlxytnj3oO8LUY4B6vWRZLjegupvOcp21KufQq
YyDIH/2DkR5/mq2zwxsLwcL3Klf960wGXeCrizx2hTh2WK6ZC9ETkhHAS8mf1TxLqb+vljD0VOHG
HNtopR7F001glJg8BOOSOIdLJbLC/MNAICoJc7IpBzDN8vQN1Vl9Ah7nKlVCrMlfRf5aN329pXEb
Xw1nNLqYzPOTtI/0g4o97hw4nmcVevePhwyGokSjpvkSgsgCVANm9OEG3zH3ylLPmix1yWeePKyn
hTYH+gn3ECcQFHfn6h/POHLqlvGaUf6iWoXzELHauSyY5XAUSyuCAHgZbXSE7qHUoCGVH0GHPd+4
GTJM8ILEAHZUQ1LpJuc3d3lRmYbTI8FjqJYIVYzgXu57gYqRkDCxhyhBMUAc1N29Wp+06MA6ARqz
Mu/04EutaEbXAWTrSvSkRCyPEFfyA/e3SH4SDrPZeCDTE/cnlP3oY04sYjEdUhUPWEEJ8iaybSJO
grmrAdCkPpYmXD5RO59kTk9UpoLi82Sbnz7GH5adTrO8BhS+KboyShcZZ00fdPMBRye0M8TmjUsz
xnt9VCVihebwD8Ah+B7fq5uSH8gQOzG3a5p3Xh5SegBe5Yl8Fy0gICCZ+l+NnE1+t9yKs+9jV0Wv
XL1rUB4Ai/CLgnkSeObsATOSswLFjYsn70oBU5znoSil+sFOP1l5GRk3b1e0uePQTc9kOckQzoqg
nlfeRHiHXaX7Czp2mz2QWhvi0jUh5KWkhvlBNnwWjHSTaFx2IZ00uxdy6OOsb44llQIzobnui0fj
FC5eFYkbv+n3PI4tLRr3/wfK/4psGK/tXpLQTske5bIbkeDKM6N0dUXz6OnbC+0JmGTN2Iyf1byT
ZCBG7a4cBQxwCLbjrAcs6G6bVvHSk4etwJ9tfA2T8Rx6wvyQ1UmJcDd0YNVTqmqvuooZbifqNJUH
e/Gd5Uc7rlt2G+6I5CyRG6JO66WEfq0zdfYcdoYSmY+p9PlYo+KTsoyB0/IBYu6yqQvX5db5NzEo
YthlVqUlfnrov4mEXjvgdJ8ZmmgihGJfKtk27jxce/V+f0811k1SrM28n2y23GwC2L7BCzt71MvP
D0xZw48TxpO12yZePz0/vr4pAsfQsqsg/4tpU0XOhOufWAXmjkyrorTBN5UFMwSpsytNKUipG9DZ
01quuqtiVZQvu765KRtEbiEXHWA2AL05ZpWRMjsD6Ho2EPsfeFKP5ViIhz4LaH+a+WpRrSPxNSd5
EAandQb+XmgcAGhBfXbMfMCeWcIU+b1UihGDntN0VyMEHrRwvnZhE6YEVfgqRspHZGYutfkqrEop
Dk1IhKeZ59t0fIZnrIm7I1ApTOnEwS3HCJMMvMd/WlkprQ2CZNhfOieA8ilbgvzDDT7gswGjsfn2
xZGtDt/laWoGYnTHqbTQjZvLkkTNqS+1lxvCY2rBplc6wRQqB+4WGYDaWZmLIn6OgtirP7TpvsHv
kD2nUWq7RHsoxJPHa3LCsQC6xsERlQFuv1ui3jRRfEn98J5zn4rZnX1ybzs3sWW59UrR5lcuDRuf
EdS3xRlP+XO3CeeUX+vyPRch+QpYsbaIVvNN4zfOliBcX057ZKnBHjAoiC66iC/eiE5eTXjJuz4c
OKrCgHxYUUxAi+TAKhzoqcIvhfK+dVOUMP9w12DrtOnXMXvNflqJz2YqkYIq/8WoyetA7MgsCWII
tG6ssvG/Qd5qwfEd8WUHnCkzWz+JhiJxD8AO5bGOrV489fcQPcVnlZSDpXYDyI5vmfpoEN4k5NdM
34mCcE6vSWR2YdzsqdU/0rpY81U1RuiwXAjGq0gOR8nTmbK78EE8YcriPbdt0SZSxeVG8Q+3L/K/
UAFFM1gY+3tdC76JS8fUNoaviQdwoX2bbXfTP/YclOEj1Y9p+xWkTGYdSNxsVP8p3QaqbVSeIsKm
1apfarKrPQj/53ZoDLdhvPpUQuQZq1qgbCQFcDFlDLT6VioXM+iL+U4lHiMSfQOqv6c5ZGd2s0Vr
WQ7pDXTf8DkeLllx4dpdLUjmhGPDlK3V6UGDXo8hTKQVYYwLeHTU2NcDAL3qL/3GzHzHWPS1gz0p
LemTj/2FW7yx9j0ViOQmuLlOwj64Mw2EOQKlU76m5PcjSPK5YkMFf5jtmDkqt0dgVeu+5TP3orX2
1vPFApLA1qxsT059ebGsSyUaT85BuqQLszu4uS2TkUZbflqQ4afWINdoK8FfNNyiXlCXeFwpbk90
HZ12e73kPAF0PL2BU4B9SwWWjJScicQslkWAIDXD7Ad//P8tB6xm0+iQGR2vw20c9D0UbsxH38Jn
bOMZHEULu4WaD8JgUDz9NOkANbfWjK13QSU/LFsLuOtw/ml/cjXN6Cd8ikHkay0HVKn3B4E9xxJf
rCkAIF2nP0PsoUJYhqMytvUe1uge/hogPN+bTZl88Pa2PrIk+7kQ9Ev2/JiAbFGs6oPZWnqzvfOC
sH6g/PLNtyDOmkpUplUkaa4iDzZ+KHZMl52XLvGcsS2BrY+G3G3/Gl323r1aqoqwuRFQi4gYa+Wf
LgIqoOsAJyjmRw1kWI7bEMaIirme1+gQQqIivWIuO5EbJjD1bwG3ro7gvKzKqNLBj5I70gLWfjUU
yD/+JYhJk9AIirkeGa7XbzBvAwyoic5zKy0M3eiIvlWUO125zOOeNE1zYhbY1LRe1heaEwzIoQHK
AJ5Ki7vXAtNAO5UFeVp89mLpZw02noDBNTGsnNlgIEDwNhH2T4MTE47VPxA/e/omu+FrFWvlVaoA
OwhpNR3PA8weH6gvLQ1Tc22a3g7T28w4ikCdjhhehhMSsYvpAgsMAFWeNIMbDMV8PhPxoOt+c50e
3XOEDIADTZoH7iS17wjQiTleLQBjZ42si9R+/3+kiUMJSpt5U9kt6Wb6/u4S9h1FkXN0a2bScuAK
bVKQ87aif91Dx8mRywM8H6oqH7R9QY8rzZektvXoITz7+LAGCPDMuBoA9SoR4Wt2rdWJT8f0CTP9
enPTEUUuzFthEQma3AStvUveJVJYJGw71+Vcrwz0bBcEWmb8hNmCMdTWBuIJn+pk/a0ABc7TaqKA
uHljm9WXyzCkzw9xaYTR9rD31DvsU4A1vP/iTwcWMZwvOWs2wgKGpk9esOZXnGYBY0utRsnNAdVD
RODIgwZGJkG1qw3aUf63uf17pwG0K05iJkSZP9CtPnPS4xDMAypnuRM3z4SZ4Jz7W2p9XQsVcCOJ
KhESB9D++EJt3aZU8OWZ++px01RaHmu8PZoBRGOo7BdZ5xLkZyHQCUkxDK0873lxS/m1JBHNZ9C2
ZwkJqUKhRT8LyJDoAyXw/XL3ziDFm4wxX9qb21Iv7uaRvieNQed6G5MkWjOrStYQqJqwOz7zlGcc
3nItVoYDLWbn8Veh6B6DZYfvE0Lb0k7ljdafga0OR6BDHBvi0kOgDMXITwfisWCrYiOjgTBdl36P
xSGykf0ehIBajc+M8eCI5z2vj5G1LV6skfwRrzz2b/TwBk1EOE1WnMWK65AZK9bQAo/kCacOn3CR
jBiHJOsfNwn82qN4b5SFPcn7hYiWMms/R4CfKz4VgRZyBEuDgcDehg1LS0r2VMQR3WYlf7Alb1OR
i3LC2G04uMl6UmEGSqNJiYKSSD/wqY17w37sQaCDVJD3FSL+fxWjMXpAaTscj33l89I1nCYw1+7R
I7oxPUlhnLw3N2ESa2sL58dY+1H1g13GXfMBmRgYcfM3+Q3gkYeacf7Ywr7oZPDAEp1lBeybpGL1
/SVvuKN99ZlIAlYFwahsBD/9LqvKs+9GGzFhcx7Wf2xhFXnOyk4jZdPdoax0+ckZfxb2WKnhGJkR
lobhTV3jFW93Qb+loqVYxVs5RdbDAF8+hxfdD/IugrOH+NOop63g1aUCTOddmWxTQ+nVIsZW2XtF
5PE8V0XiLfjEFRB7QzXBSSNPJgTEKRu1xnrtBFafHgw2itMZ98tVRwqxkOR9MD2vODOvfV8pOwrZ
nx9VOGOXvZiaJvYEqqMuN5Qb9jK+M7kkf233DDJfIG91cS+DOgYlt5LLpzTPBHeBnwen5lvbEowo
2qeQ28B2NDrviAEJbPonvsvG6YdE1X+y9Bw3fYcGnNXyWA7xjZuY0i4uhQqmv914fzFtpP9EhILS
Q7z3DjM/1KhCVnrl2jxZM50Lb03sZoW9v25M9QhQAATRVeLCLnxwAOZShjYkRksUPzYk6NDOLW5J
cBlaz4mgQDkJHGOe9rwjt7sIajaoCXNdd5RgVG5HXxHL3ZRgkeGj+IRwqQ1Izk4WFQ/3wjjQLHvd
lP4Py1yK32NjPNAUwO7sSRBVuTXj09q1dflYsId1Bf4MhYTzmXfan67BjQQ7STBn1QdH3vMog/Oe
yVf1ZrAxFL/qv5WEInF6bHKHUXQOSCkiJNOCAyKP/nCxrBG3TjmZJiKbFH0aMokGEJXP3Klh+/bZ
bPiqiQO5KFkLoyhTGtBAvYBdawX2oKY6Vho3f6IsyAs9thf7M4nGySwczlH0MThtzbiNLLZhVtjs
fOvZVnrVnfH5m2vAEjXOn9TybEgeosLnut6PlIfq/OGyFYncX6V5gj35WY7n18DBSM7Czpy3dEhN
2p6WozXk9aC6S5+W5wda+ka989rY3DEMsfbUQz+VD6LPHN1EGsjqjyrguusks07iMIBVD1hL+0rp
Pd1+IWfwGxBnDQFd1Gae1ambfyBWq+Hg8kiCMyUOGshBK9xE2utVV4WXRKToDKx5m8nFp2yhm/eI
gu0mfDe6FkCRMG6Qjph31WnN+P6kFg99Jtu81cO162CEixaUUCaP8128gMnIq0osTNsWf8k7TRz2
/XbSGHzGcO1TpB3DmpHqnsuNNh/ysZrCS5YENv2CRWWveJtWcq8Hxfxyzq++Svm+h/Z0tTGVXlzc
OsR28QgNQmsbSHiG3gjk3nWO0bR3dp5GjyEu4k0bFiQPb36vpZ7hz50/2kZUhSg1wglWzCB+UVNe
ACi4A3wfUKSc++Cx3VbxQqDUqKCmB6o/tUV1iJU7kRiFJt9L1qC0xynThP3gM8ZGK7+cbtZCmGx1
cKkKcyl3MePkOS+9JtunlLg2U/h22CQZOXnv9icrUvTiGykTi8zhCF79vVdEvrQx9yq1Fjco505c
okGYkBWtr9s73Dn635ypGsw819sEGaOZLA6huz8SfdgFMBCjncqiONzdmY2SE6e2TrGWF3Gyjdh3
PDSsxespAqKR9Q5vWHAq58ABF4Hcs5e8rbx0d+MVkYBkVfdN6Xgn7uJyksghAWeo+UL7QBR4FonN
VnkWrjCPWlEE1yk3vLoevJmc64+tNQGIHSo8vKQ/rPL6crwpyP5WgyHEyW5fi0Lfm7FybuFSpxmd
YOlUz1hJZ2Pqx5uP0LzoTaElqld+wiEDdix6WDwpVzURJxVbQShjhXfnSXUfMxlf+HQf3Hww0twx
DaxfHx2o2vshJd/6tN4twYP4X0kp7bLzy5SSG7gCvjyvi1YGE8YDcwSenqsfWrwX4QdvcRZQPeS9
hZj1QHsHqBH873pygzBLEUFYcIQTfiEre28SfxgO+bXG4CfcZJVd2uBy6rX1GIojCs/OGHniavSU
gARYTnXsmRVrjjA4Aeff2xdM696izDbnZIXCgq9Mi25A6M/azRSsH1lzFVga6HCec5e28oTRrpX3
bppxiTPsGW0KOnhU+IalUCP8gV5lg6JW6Rr+D0r7NHT/3WzSRw01d78pDqIBzX5vtGS29D0msqlG
Xzvfr3xNgFinsH1wJ7AxsvnR+hvFREztRNxZ11OGFJD6TE3nUtoU/6oX+Jspcc+CSxI7UmowJSVQ
NZr6xZKOWvy4ozwM4vgRT22OBCWwwUhPysfhXzDAVZk+bAi74IlifJcfpRloKSQWMVkSjMLZq55T
xwYUTpZvZkzg0qrUMjE8mz7d+U4WoIWx4KVNl1x1cMdhA5J4aUHhWgsJbM/0k/Qh0kmMAaqeI2I3
uzwNgq+zHRc+8Na64X7CGRIAIlPO7KskCO4j/UjNRS/sZP6xZMuLCl8IVfx46WQG4l+c8jFiZphl
OJqv/6RsMVouqsUnNb14PWhTSGm9k3WXj+kX+pZq9dB83FDU9MHxma9bfcvw51ScMU0rN+FNXkDc
q1cow1KWEjMzongtCsGumYApG4gNkqe5Or0cSMOh+cGy2dko12foKUra66tiEjI+XSxf96+xFXtO
zFYMXNfF8lQisOwUGE2Puj3buSL+ZfXwZSI9+7szIYfFiBSj8E1qk+NEtbRSMxcPQoehoWzEEOdb
LjhZ8tuzdvxx21cBfiBS2qfH8cRZmDW1EZefM2Y0ziSkzRZgRbKXci/aUBWaNYQUSgwoIzIPLoO+
XKi3KUKVYryes+rYdZSK87XBhn05eV6DKKDbRfhqMkHTxG7SxI45LMOl5hLvDNc8XSAo5aC19Ymd
8j7zj93KltmX7Hgm8yKJScuu0WDVA98jUpJtQnJZa+Er3Udw0Xri3GoPz3v4Khu8kX1tFfodEwt6
yowNSLxnougC3HjE+Xswo3gj8dxt6CGs41B/xAFlDj4rFoL2sz4FYuLJ6JBXNtKE+FJXXFGca89u
jGK8slANYytWgAUEN4DEzVz1b2ex2Ow7kz77DeMz7aTxXJA2y/WxizPoj6la/TmB2BPtAs6glWIQ
LcjZM1MeCOdMjMCjtb/A9r4JCJWbuXiNLtP50NqhFaLaVb9aDzuPrNOSoDtpEQO126Sl8F7nqbvZ
+5wfiDN/WS/16yAyhTEoYD3C7FjBHrD1POtizKEWBeKHbtvpqNBbUcWMCFQiUPGOMJk9+ZbBvdTM
07RUse539j6/xYw+9NVnYuiFlYp5V0C6KkercbpbZTskmcC5TDxhs1GyL/sc6TSlMXs7FDkFxmne
2hSgA1yLgRzTOMLj8VsiVvgB1OR5eT+c9EOP7dy7kWdS1x4gDiQo1fV/q7OMRrpEyf4ehV87aYgz
r78obZWMK36L2e/fqBPBSwRJNEyid9LGKnDsdRVyOfEm9Oakm/pX1BClCWraA3bjtejTVgdMyBNB
OMcKeWzU+pHKYPifmCuhsDR1VavqK55Ale+HTS7V64XMrT+6PBQZTolgxdqI63Smb6Cg3LDT46JH
KekijChcY0aGkKWrmNpZd8HNmG343lIgPPL9hbPJen0nCdh+tsVTTK2yEsi5SELNKMvSI6tZbGNi
nIm+Q/IHXZRO+q2SZQaSGSpzFbRn8PnDs94xp92f23rHpnM5aH4NitYMmKTMlFBbgacOjMrtjHvO
eyz7m14i65KC+XBxJjrDly308nwDFLSfhqvQO3vigNgElnUQd4MlFjYXev0H8xAlsJM9JCjoQlM5
CJbcw1LZsSH9xJlchH4K1pi7jkZKDghl/h5z9Q21ybpzl08Rs/o6KhueeAOgDY6RB9aqr9XnW+ij
OuhVZks//Wo04KdI9xBf/rBw0cpO3OHAyiWAmRq5KNMDMivrhS6kiL3aMxdXMMw3MTNyu6PaZbxh
3GsgpFPQE7BhQcvRaDpYPL8AVPTfCLw5kDCSy5TCIYXHmnFu9UOKL7W92yzaMTaq/D8HltWgJPnn
WUl2Dj+UddoQ5HAuT764dFfmQByMaW30J1aHaZfKWez26LRyOi3e2arRw1VfSUyzd+FrSu5aeAJh
VVgpIRp/UB8uhCAwcufoJTIrnY9Whdi593j+WuPIxcIV+qN91MymCQHKDr/5/MeUg26y2DGXGW46
1IXuddmRy5CsmSMv0Ob5/hVal8fSpJjC+GgN6X0YM9PttkwtjI0NZNoNV0xF5vSpiBcxpkS9n2QV
xqNR71U15/DdGhAzyl2bHrKHRlU93xqJDvTSV7AbSwaWiCF5BjDnLHMU3HD6Cp1biNHLXRbYvvqi
eBd0mpQf/uNkb7AutNPnv4TKL4u1GkpgWTP2vjp7wWQJske6TJeoLjlE2qWCtSuMgj7pFxS1ls7X
PzYX8meuNbb6+g5I/xSoF3CB3VgHoRpEvND2WD6wyBwN1ET+HZXihQDXMikc6UbZeKrxTv24bQeH
XCBwx24Ka5yK2jjY0R5iNGVyp/RPNjcogmKFKD+WPg2756OxbCynJmfpnYO72JTq45+eyTTZn0in
r20J4tSMKSaOsVeAqJSpG0NPP46eFG7wwPjTrZVGPyyLHjd4098lEwai8t8+H2YymQc1kUbrKYQd
q8QiJppDssJ39Dq989h2cFzyCDbEbK9nax+aq425/5Cc8wRYGRpYkzgPDLLsNeRbw5KkpMNER4Tk
NzEnwrt5bYO8YMMjo8XXm8YEZVQijF5eEZopHCPBBNTIyf0Y5CZ4OGcXn+BiPzzbKcXu6+qzOYCf
Djq+mXSNxngE77b8YU4L3v4vg86nQLWKzi5wyIjVeZR6xtVFvYQNB1Ux5AbL0fwdkpMdjHiNiy2p
dxm58Tn2U3ZGhufO3gz3hwNvxfk5NjLmTMrzgqAV2tIahUZupsF0FgaVljyQ5vjk0jtg9MSwuNpr
SZg2lcv9E+SYyddVK3q3UmG99dkFOeoirRR7wQN019ISWoabHR0JRDdDjAMFwVNQ56wGE8LF+av3
teZH/GX88WFkpB5qWtnt9bSg5L6kKqNU3dFtBjUMQ/w9+k8uRD7gLd7eLp2wkSnQKFfv1R5ElDeI
0jm9NU4fwI9gOKVLJDVBmxpJIcxYfknKJCJd+8aBJK7Jm5o7z34BjTCnUUFVN/9zGRMYZyQdSJHH
+y3QvjFY1Bsy9KvCAjaB+KQM8MsJLlgDZw0H2jDOcunHo2/FCIJSqRP3h5Z7FJwDAAauSfOFouHX
adyzTiEhPyRuBRXor8oKngLp6599rpO82Kf1j8S2vf16QaJHh/M2mb3RgO7qkdIJbGF73rE4YQ60
5yXGiz7uq/BKPEhxaiLRaanILcn1QfvLzizEq+AvXfRXFWDf0yLSSltN/k3fxxAclscfnWlq25OI
fZYCniZQDTfyBoKmjIPW8Us1c6awPOjwkzzMdDTFoxP/7D90EcX5A4tgx+G+CSkoI4Ff6pj6izUz
+2rL1LisjVYA/5RkphoVkj49I+8hBgSBRl3FHoHf7cwYEeTocx8dzamzHhdXpqfv6Kax+4MqmiGQ
VTzT+nv7Q2YZ/3cJ5YiIW4QOVtl7HXhiz3FR//4XNp1t9tQ3taBHYu69w+5Yl6E9x1kTSmopTJ9Q
d8aQmRGF9mk42/9iieQLwrq9pKH19CKcAHbuiiUhcthqeEVMoj72HooHC4GsW+tUkyyk5B3PPAW0
ALMqzPBWaEYGcZpB0NdnrYT+4+bi5Ei1VKDYXpMSGdgmUT7PVcH9MSa545zjaKKzsnuvYYm3Zp3D
NMuaco/303KZOiU4hFszio3My6H8WraazJUtNvlcgpVeNTlWAcZ7D9AVZEAS5sM5dBdIA6RvZ40g
Yi+p2Ss1OeoRtQUXlURxltjySRJ4xD2AxIaoE8eh5meEZcXO/pL4yVd6F2mDtSkILsmZS/tUwwFz
4tkReEY6eMDswxsJsyTMdi7TGsrLh26PJUWigHOnR9ZdRoiDD2A4FuQw22UFQeorMEcAYGBKSJNL
yWaKicNwcORRt9Vt60+2BICxLXTjTAQMKDa7PXvpBwd7y06CgITK1pEZx0YOwuN+PLovkwAv725P
GIzyj5/n2BBkH1h/WW0uAVCcWKK5k3dPc60GGEHA+/vXoZrDqi0swV+2P31GEy4JZ6MXfPmz6F8n
rsWq6czM3jCDZoDoYYjRpWjYmXev47YGF/8quNju2bpnLjX9jRO5Jq2h8iVv+vmyeeHyn3TJ5xS8
eha6aBLk94LvNHunxpR98rOIm4+aoE6pY8B7PNvy9k5Zi5XnMGt9smMcSIfU9Hr83320D5QrYoOv
rhp5vNwPBf8Tly/iXj2kwxabLkWljRsDmpyU4ip5aTb3thUTaPUp5pZa7ekgKmHIDnbfFnQdr4YF
s1qEq71fH58s5VNkY9O+Idy9bAZvawrwE9vNgog4bIBiH10tXthMiLqXJZISGUbJolBiNW5uDSm2
qs2e0utOn6yvLG9GESTNHUDEmBLTFU0Npg+qt9td1AU0MPsAAVRpoFkyNFYtwHDYO5PG6Sh1uiug
kAjQf4hB1Bh9Qtd0sr512AI5soZWTmp6BYl7RAA5eB7mp7cYWxjSQFRuPVk1jLcBsyWUrUI2GvDF
+5hKXBDwrzat6nVVp2SMUZeWGz4P+tf54WmcMTiwEe1vQhp/DQDzmiMsxdQSX5zwqXQf5pkRZE2J
C7/vi5+MCj5hHthKeFaTG3iPMoTaPr28/GhHNQ0GVaBZpd4FCmAPQFrQ/GMGFsaCxSZ3MXDHcvRu
NNniOz7/kKS2GZ1FXNcOdori1FBDi0wXTNuKauuC7POrO6HfI5fLzpaywACimlBxItR9bLkMdNQA
0FOOl9qyXAD4rNuaUHAuYmUmArNuKhAEvfrFppTFOAmZRc3E7UqklhsrCn+fFJYrYjv7H69gfBDY
3aM6NgKV92E/0tTtbkcE9c+S8Yold+LiarjaXpQBJTrnycLFMmc0W8VIEbzL7NTDW0LhXaql/Ul7
M9kuY3Gn4JtC8MPpmaFplioVywZut6pw4jUQbI9aRxTK5LLQHVixikxKakQdQCfCLEPvAH5zDoGs
biOzGndfl8rmiC0TbCVzKmXKhtZExAxH31bGMMHvAOaRKIIhX0tzJjDrmCzinIWDDFikc83euBhb
QmByX8SpKGNDe+dda+tTparIQKCBMd6C6TKzRK90tTxgwdS6EE8vg9r/M1h0TEUtZPP+TOxgpzax
x3+18xSjVJWV7Kr1sd3crpC2elhiQ33SnKgcDoqshtvqr5opdSXGZ5ko60K/zyxStHeaPibeLIg4
nSNse1IOWVASTjRL01eUUYkC2uz1ZmVZgsq+xpy22zGQvtITMrig6ARj2abuBcHGA8Jv4Le1K6wV
diNevx81FmLdbPw+rIZYL69JJ/+XOM1XlgT1PrEn9atIrmCkRCL7ugxs2jPJko+FtyyI3WbkPn2c
BDvXZeH3olasXKW12UOuUwRxjKqHiPOUEorR4ymO7Ee5+v/iASakGCMIeaXh3fnSBhUbUYwc8A3S
DfJolCHJj0MwnR2ANOSQc0Cc8zXekvBppkfmrnL0nxoGiJ70m7p8aqrRQniFqWgtb19FQSMnIneu
5SRII+lmytKsMdsfV6viFnO91LLP+014C6V8EtMYIxj3braRanRH5qGyEhhihJDy43sWhqL0SPNP
efXr42ZlLWD78y8ty4xNMpauXsa3rpMos4406p9CyZ6VGHbnGSh8WiQGkQKuHAy8Sy04eBM73fvS
PHhY1gMxcnn6ujYXhkvS+BOeHV/Je0/b2JtA5pLdm+IRkjT1NCO3aGMR1ChnksGqITWz/FA6u/hz
5m7dMDtu/xt3GgoyDkZrQS9LlQbem0M5BZ6WKcL1iavZqPF9WmY5blPaYu8obZnFLUOAINHDF6lI
2q0DnVVn9TWsMyjV47of736r5d/wsRUFppa9tiQJKxi1JB9kte56xVUgqNkZV069/z9CIZyTSLKj
+EfOXwPwWEScAyLTpfxAdUaR1zIOGOI2UXqNVVZ+gmzGplOsh7QrvAcDYluj2CrysVeJv2bs/yrh
I+05e14TYELD47PMe1A642WOf4OTl9NFHbKYUhxaMsGZrrn76ZQhWEW3ONCTrVG2pIByMr9pEEq4
efOaVWRL82o5sy2NfMwIq6LsHKOeF3NSp0U8tDr6x1Lh62EpU6LptSfbK4XOADxlQHWifMOzit+q
RdirxSU0VIalF5wCGXxOaSSUs4Kb/23xSQMa2QHwCi8F0FoH4JtbP5T0J+FP/q9/3knUiQfIwn4t
LJ6LrbbRmRqKjGEq8DgkT0Zyq7HhqXVy+hAxbHtU0N68zKaJnZf4oCX38oXL2nRq/KJXNvgAKrQe
wZYyFXjTdeAhdI+AtQKCa1pvhsttkGkcMaidUWForb3h6VfUy3dH/Zz7LkFA79w6A37r7xSOGxDa
jgmEmKAqZ7WGJt8r/DOBzVCU1Pi4amqmjQwOAeAwC5Vu9Ukg5ZjsowQzIzsanCt+nIVVDbCAg3No
RQEGg44hYNpPHQt3+wbMvOOxxqDqoxUNEK6z7fkML4m9TM4E1hVl2nDHDB3Vncx5SPGN1ow4G0xj
SW4q8FMZautbMTECw+va32YFBc8Nis+vQkQeagwdu+b0XUF5zjKykiTnj1Lpt5RH9Km2Z7ebrvlP
zsdrm33HiOqGtMmHONc/JSx/UKmQ72vKLoqbjwXyXzYTymgUGXC7sXrxr0GvaJAFSaKS6EAxRCtc
j5klvBK6G49PZzqC0AVPkgzgV2bl5/s9BKrrc4sugCqbv9wHkSt47S77OpS2YhLRPSuEHTOvbILs
VI+2tSAUiXJtCuy0DgHP7wEn/vlTvMPiyjZDw/JyDsU6cl4b8B/Z/9DBPXDmXC/HdAu/mFZwR/52
lZ+EVTd4Gf4jsZxHXGRnMWXEql9H1781+YQ+ekN7NcDq2rpWZgpMO+24h1tLqfGsZyCkH2mG4XbR
awhwK+LbhzmJIjWh2Lhrnyf4fCKeAFfIro7N2IWWPg0Z4JqIN04B0ZfnLipOEx0P/QoPSrnxzAcH
8XBkAyCvv7LgF9bf+A/4Ld6ZpAF8gYEKYkSNnvvFrWSnHwnN7UVkekmbGKdcf6T4HR357QN91xt3
r+JTnRR26y4sMQ2yzmHtlWmfmMKzGRf7CZH5qdOZ/ri8ygzJ4jbBA1Aov9UmXSkflpyZAO4OwLyv
y1P7T63o82qb6AMQSwOEUNe+HLFzC1s/e3Ir9xL/cw0O5fgLAUclCn1KMCU6xCyR0VQEOqJJQuov
QQAOznZ7Bwn/NWmWkRN4E0uW4NGhlKgulHlOIKGOYVO+yJzzXhOZ4AAKToaOVaRxtCcZrY31GrVl
cQ3Z1j0fAz6mYz/eI3CW0O8mzj0MJxOXyhY88wdUq0G5Emd2G26wf2RlNvM0cC9HhV/iyxTqrGcI
0smri6OEbyxGuxxKLfUKWID+cLmlFibUMou4qG003AOY0FUS3lMUD79OuAPMdhmK8jalCxjSbDyw
FzIexiwtnuI34rp6A78MlegHbzEB7JulubJQwYDqzdVQflkqU4zbY+Nsvb3q8X0cNytNc6IX3pBc
7n9gjmaJXq5rxMzlV/NtTmvDKxIYJ8giB8gwnzK1SXPf+GOfZt9PugNiF7nBhAbcA/3uxipCKSeM
ZUnYnPzJVWM/IWOebpiAO0BSqtU+e8VUnVdW2TUaaHWhW5Ab9vs9xmNq2aF0fMhvblaLTLz881+X
dPRauF6ZW8StJdFfhfMYNv73jgAExiuNxK3xkLoUXtRXVG7TG//953e+i+uAroV8U/v6YNfJhfF5
zllqN32V0Ix6Ma7OHjUCeQH+7RhY7Yz8f/p897knBDprJSAUmVL1yXD/hsqJC7TrGkvIhGNsXxiK
4YgDW1+wOgwRVOR2nPG/tVgVG/x9mrPvBJNcuxWBZOijrBhJlnTZiG7Pp0c0G9XGrOYZ08xOlpSS
F5EhU+50XNghXVLdoTV2drYlO7GxQEz8QHPj2PHs7hU8Jwk8Wjiv/lxBjZKpt93A3J+dSUlIU0vE
Vdw10IO9GfqhGcTKBqyevV0x3AmiC4ojZ2ofTBQ4Dx/f+XkSbdspbsQ3SxzDfLGJqafKYBykw/lb
7R6yGJqgHl9ii0t6YMgYyGaW0pL6H7w0newfao3wX2ceWoze9XAPNPsPvqL1tPNNr3/2j2dAyBvo
JMIUhobo/lJwK4Ymh+tgbAJ+i3W4V0Q2GeynfNpqrcBWBiD3hPiIqi435WBdc7HyC1kPBICi0yAn
5SisLpuWQheZV/spT5Xiazh+poTevsNxc1a/+Xv/eAeUFwKujkEN35pIeIhotbt0cYFmVa3wd8or
RxYndRmHgVuT1Ht1ercfWvo+f61QHcmpA+U4aLHk4K6vcU6haGyMyHjDEu9+5ZGlHFuz8QDFBpwU
RjYts8PH7K0hapqY2c88Npr6hx7vl69Y5ivxbR15fpWA+8psjjLZuG7u/bNWx1pTjYg9EQL6qRAh
fottaDXxlI0KSPUgCGJHEH5fJ/rn9WKFpqvHkCy85ypAzIzldH3KbI8mFa7pD1haEd3+CtI57phf
Y9oNheBH8pK07CF5dm9NNlb55avz2Voq7xKgNIxWVp1/xo1y9Zliu4lKAvFRhK78qeYE19aqwi0F
rRPCICB4l5n1tQcjZoJGHupAW/h+fHsB4QhdpzkTPCsy9SseshNa4o14di/TfkV3rrz9TiW+rJkV
Gz9g+B7J3pw+G303Ch8ccCGF20AphDgoaR9NFi3KPwWtav2ARN6JG8J3yMfX6Wron0N7QxvWX06V
3dBGBKh68ofB3AaV//1BeZ2sAj+q1rauhs4vHnLUDgYAS5Iuap0o2/76I4M0LcI0hMD1dNiPRnOS
+ep7Sv3GfMVElDIJQDCyOldHWftOaI+1dM5WwoHaT2uKkVG3cWerrBQNjZPg+TXLGqUwDFyzhsv0
M+dr5ulExAQMgRqkT4g+A1qWmbgmfAxZt8WrwRYR4UhCR+Sknh5MEbQMAZCiO4IoWWLrAqGfRztO
1Uq6/kUlUvrVn/V4Z3hsA5hLs8PmLXU724Lidzc00e+4UAjM18FjbI8w4eHDW7+Dr0+183WOBbzE
h+ZbcLAqhK0UW8dcwfYJqiVRVO1kZntaMn3KONqc1n5WjS/dnve/p67Nk+75/lL6v7h+5I4wztPo
ga+vD/I8VG+TdT8vgNoMZLSpK4T+gynWBLi1iJUdqB39rsYOUGZHFagZuGE0zO+eQTcNRZV2CHsS
Po2V9HsWjVZAD/mImd+l1tNr/ocGZhWSWklXn+XG8Wrnu/2ujXPn99CnNfZidUp88vWvZM86a/0+
yL+Z/cqepodStfCLaoQ+Y2uvmIlJjVg6lNCT6Qe/N+c+zwDrXIS6gZ+ynbj5yeeQmEyUW0GYfcVw
r0kFFoc4aFHsLcdtrttpA+fvSyhiQLVHX33mXyTivVXWmMF18Me9/5JpxS8KYnwOM4WBHLZkNvKX
UNyhTMGIKECrbuTDZNqI0wl4yo+r6byRw/JVj5BQfKw/xzXCGxjc3rKXYlxNw2qqV7hIZEmkyPQ0
YHz4wWIDfPMAEi4kMGMlpIPL+NVkWJqD3OxmP4ZY7nnCkHcAQ00egut0hw3TK0R5HpJVga3sQkm0
V1dn+QflD9q++4wrmZhcHUPrpy8ApzTOh5EeSdS3DYFTWaQour4xc0484tGlKCsMFV0mpwzuJDiV
TOx5tvTnnnIhCEGl1iV6NrYAmh0nD/QT8BWNPu8j86BZjTcjjmpJ0LB+BLt0XsJgvuH1qsDmSKlF
0GwfEENTZ9mEUsYHzanPHe9qT+27dAfOoMqCsmGtqhLmqsNGRv0aT5Vb+0ikuqoE+y9Zkb+CojR7
i1y+HOsQBxq+T0pnPpVn1KLLjhwPWv00xNl56iRs5B4J9Sj2A5Lfj3dil9rNbvhEV5dCe0A6u2A+
ycD2qcMQ45pepwdbOSHpWoqbR9AKc7FFExNs55IB8qrEVuMewqcL6FnTcnvDJAJYu9dhimUOMIQU
rg6pBRzvEyVMJnWNYimkhsas/fMAFKSj82Nkk18XDAbh0LRsiDNdsBlccJSmhQxi1q6gHZs1plII
QB4rD+OHNcgpoCeDSlpzvobJgRcWukmdGKTxluE9b4CWnyTM48NMXaK3cvuWu+q9ZC2RX/15QzUz
wMP5/vP31z6ETJvSzp7npukm3fbplsCrmEYMkr9ycWMmUIkGqQ0eMyBxB2zrqHCz1/1qYxf0nJe9
AnHE41FsBZ/HtugAajY/PezYE6PkMEc74Xiwhtjc9eASuHuleQ2ybw5FrJpVcs5UGWAE4BC88EWW
oFPgq2yhwOOJ5afnCr/SfbwjWxvIN2de2Dl9CbxF0Yem0YwjJpaZOVGaEkpN3Fcu+qZjH9tlY90D
RcgrPCgjQ/7fPEATOQDyXls3VXuKCtNyx1lmxLS49Ib5gT+P2ApZ6DG+Pvubt4wCjYZiuYQz/EuD
iYjJBKj/ncBpySy1iZKLeMXGxQPz8XrEsuFCmvoSJc+cR7nrtrZX+EsPr61DNa0y10UxfwDQ5ahq
WiNSnPnL562A1CIpaTjQW/D/EAZ4O9rtKFUmjR9SqK7v11M/+iANrG1o2F6cS6LR8wZMFK6gkCmb
S3Pzfga5a3Sf08H2+SSaOzjJxyf1jtHaS7haT+Owmr6pMqDj4YeCB9oMELMKlyIWpZY3GQmPo49I
tDoBlqDo2zuhZ6+lEWgmsPSlISQs/0NQtoRKf84+yiwApPmS5GNtddLzu6NIngMzuc6nG0XauJMP
b3Ml4VNbdamhvVDoA3DcROuZ1uoQwXBxMgP1jZrIogvla3v8IRcy92ZnH7RAk9qiOYjwC58ffE8l
KCaM4D0qg9TFEadpQnd41tBaOP/Zgz+E60D/e0mxSpKlaY+5UA+2LGRysim5nRWjpGrhvFISL00P
KNGnrQJRXqxZsrohLDrPv+i/qm9q698QW69B0+siPJbCgfNsCqf3xfbz197I8Q8841kdtcenrilz
MfN4AdcpEGsvhF099i+nfOYRzNuRYUP+yQtxyLWUp9pjm9PwouykxUnb5IeyFcoiUYeJhKQQwLWO
+VyDzO5sbmW9ZQCp1DjpKKPHRgkHefVBoszWvxJVWSNRnYj/1yxapF863ed+yk507vu8uriH+yJo
vXF0XFc+dHAzhwzTV7f/H2Ipb0D8qEZuxnvp+Ht47UdtOXjYLHW//9Tdogrfly6jOPsRS3IPqo08
j2tn4a7AuyUJMq9t8sIl/J/LGCBmh2rjrd6O6N9oXZ2xorHXdJKvL6/4r72Va7rzzzTO7lrzAagj
UlztzPL+tK/J635QQjXbxSdyDObV0Q6WmsdBQlsvvLfsWy4Y+JNij9fjRYv1RpFZ2upDq/SqATR8
mffylSpTjwRlKiZNVuvCrzE416xKkXVR44/Aafs+KQkwmjtrx49xZW0pNOXikwnuhbBfDpfrPe8K
2qUSc9gu3bHti0WTGkNYHhBITPe36soTXtM8Gh/nn6ACvjJrLOcwRm7R61Gh5qE0+gfOEihx8B7C
lRToup5gN4wp1EbTZI2YWwc0zInk2P7z4ppIZ4Lri/l0t/PQ8l9Sea2TerYxKQQMMgcxZu4b1Z/z
Doxd+q415T3UlYcRXD/ucn9jXKRXvtY1/U2Kjk7YISxwqsDCFn3/9NZktUI2fREnlMlyKjprMfOf
b3y5xSP7YSx8J8JwTXqHjlwjBKN8QuKJcfB0AkGwOZFdWucxoo5sNTYXGmGx7zxUjJBDwyIUbWBj
5V0NJxOmoIELOq3bkcLz0LwNlCn0lBdYUohk18Gj/2FFGi6zzUNBKpMvOn+kiFgqIBzYeMSM/J0P
flE/WI/67PUeSyF8DMXKS9X8cfYezYc241RqemX/hWd1jXgk7hPJ2dd/iY3nBbCsr5ygQesYr+gm
V2wzPZ3HIPjoCpqtxoa2+1nV8w+IHJKPDSeLtScU7XNC+ei6/fkszqUZ6m4fNlMRWI/IN7rB4NWd
gHUTsBr+cXr7N6uc1vbu7sVaP2F9VMiaz4nQvQ4uwLvbRVdDilJACYwewY+fRIYsE34lXiNFCMel
1iLjeq4V8Q33g3JitoIbp897qC5L72vP9+4JXRf9WH43ptAUNvFxxMCbwLYMxNyhjtU//WmWPvjx
h8VpFAjrBAjaszAzgWdN8SmGWglemGFtLpi+P1ouw/Rj1x7UHMrHn71evwQDPylk8WjSF4wIW+J6
pTu/LDBfvihMtdvQgEtGHNrru+pVBKusY/s4D3RVqCHHM65KU1owcz8ycvlHbE/l51fFNqsVL80l
4jeknFF68NlxUJlDG6Bosb05OKSNQB+RWSbuNC7WR4aa7qpNLbRWSbHWxuNuf8bWQ9tluYRCHo5/
YkXV7IMCzNygh9tRGqKyUcVy/6dzjQDZJsT22ODTH2ZsFJAV4UeRcQ/ItWEVjB/4fioKd6ktH636
JaCNT1DgfiX6bftIHFLXNTdaXvujB8jfza33aAbdx/Rq7M3eXVEnZ3mDzE5F/QdqGid2zSjx43BX
TXBYQU+8Di007SREIZwQciXs44ryq0Wv7BdzjuAYuYrAEtZHyN2RRdaExf5ej2oLfGBni6sbJ4h8
HVKzeUU0C2ufa79YVKCFvRO9UrR/3xPAJu/a6hsWlLpN8ZQ9XwJwbEomWhzbfevQjuR9JFhLBJBO
5Z7IZhJ7UOvAZ50ZZg/8qKpUi+/8txJve7B7KGObMQkyfGAhiM36tGNbJOiLmOwe2HJC0uSrq7jA
VMnY3MhQepRDsGclTyzdZyw8d0tZRyetVIWtwxEdXWNouLaAaVDSFnQsgSLyIo2y4FC402YK720X
bqIc7BQYkcoH8ih9BjPxbsJ28F9O0uZ2jRo7TzVgli27Y303ZtRXDMPWfmDK6/O8IJgJ1J2n1spO
kIybeWG80TGhktoRi2aeSopbqTXa4u9e2LO56sJrjuZEoROXj0R4AALk827EBIrVtrdqK7d/LUOy
q4YfLexVx2z+bdbaQI3fqokxB1WKAALIymVEyb063P73nkSMhZ0X1/Jj9gShYYDu0IC12CVhgXcb
itfUvqmrVIUw0bsDgMmjHGbQe0VJvumgyUY8yXNL5lLSXYFiU0oYb/JFdB/ZQiRG3GclQmOTYjhg
JQka+Ikp4GLhCRR5HqZBAXAQaDlIs2q3GBj7769N8IVpWqzkk5a/WKSbSaBgILZ19oMNUdo4KeED
BRw0m9QghzrG6UCcm9YWXCoiO5hCppGHEKoGdGCdyCBbxN+nl5ZD8onmEryseFgwCNbZN7kPloBd
5t0J2Js0vUolfxEEAiWzoaNwOPQFvMtbyFJtvS46rk11w4k//z3nBbg0hKIBywennztG157dWEmq
v6QAath6AuJnfWXQDZL+SFWDX9kCFZiX+/HyC3ECpla2ovcKifUbbHxAaejuP5vtCwRmRuFmdqLk
HiqUSQA4HzdLRv1Fh1xd01Q3+MqN9TlObB4NxUBCXP2DaQ9Q5l1JfzbnSACgS7ojkmMdZV/ZiRTB
5tX9eSUdVV5XHjI8W37l94fog1hnX3zSVyPihOwN35TGlAM6woJ88Jg8nziRKv03iLIECRW1s2MG
nPzvF3B9sJ2HPCu+lNUNiLSTiM/P8+ENSP/R357X9lohhC9yHqAGL0zXRap6ZmdJggq12LAYc0IO
PuajER2mgES/c8UrsO++JEOHAv2L/Ge0e16m/rPezvfhPwcoNjAT1fCQy+e7etq+x0XONN8DgQbz
LryzntXMPN4nV4/IFkqvY6SRt7wjd/NYc2+ggRt+IUYjjpBpcv2Nb4YbRlIAiBefv/Y2R8LUJtJk
JZTuPDjtSAzW1mX9d6sI5ZygGyO1kbTz9K5BOnvlmwKLKsupzZ3JDoIXaGL2deeIvpTNoMZ+2v6H
SCmTylgaENqa93wxZ95d4826cbjfXY9mNLtCKW7uaNMzs+anB/YDRaVmEWAVwiSwdJaxMELp2kB+
msrn+8mpGnM4XFX3G83BZCpzhkw1Vqxbty5Eh4z8aOuM5NfASkIsiNujvENK7oRM3jHpHci4kuok
NXAZPahDoubTBDCiZVE2akgjWvdkAXe057M5/7QJLWNsyNmBms/ssTA3AOiYx4DyMyqGe+fIDGLL
duD6n9f46lN3GFjmLQuyRDKR4C/cheGZcKnqfPPqqd5xCRDmEiMkEjdvrZiPoqGLp+HeKppJX6eK
YiihVCV+ZMveTxBLPq1jfSawYk4fwLvY2jdtvdjldwmTpNK99UssZZhDMU5Mc2NhalZVN842JIB7
JFwnBwrd1t5eK/Sw8LM18r2s/XXsVh22RCe7Nu8E7KLmoUdu3IauopNwGvRvht3gssK4jOxLn30b
iVw47f3PiobpNH36gswXQTP4yM+lu60GkePwznJcEpwUS3BomYWZw0yT8+3/r+sdVmeA7i/NL/qD
s32HGvVAPbfQGPUxVIy5DnvGqm2ABmLf3pR7J2OVf4dnL77ngt4Rx/Ot+mq+1wcns+3QLESHtmCX
Wo3EPNRNotsMlBJ/brJMyLFfyJPxuXD/YV80H47LxndSsw/WpBHZ3JIbxvcNBU7CM5a4h0KvZADX
5J/vUGCYF4EgbnLsP6i608xA98GalDRBk5HeE2vh59keQx4khrLlJqwvv5gbRkOhBYf1f3MAtcaK
6/vRfrnNa3iz5cDH/gFszEUaGsf+R3/7vRr48+AQXy0zfO9nEps7RpMB2oKeOHoPP1COVq5Bchjf
2nErxjMZXojTW5CMylRyczzam/GPYwpW5L7H2zLacMZ5yD7LnRovUDJ0yZugDIdj/xdep/Z1+OVo
ZaGyFI9+u45xeTXrPK87WqmZP+c5T04I5rF+Eey9B4CbtQjYYx1WJw89ZGhr4XbmE8vdJF30jOHC
rcdnhizpQgmpIidC55MCPlghyvaYa6M7s/LpE0sc8xO3UQP/TJ3MyY4dZuZwGMw8K2gVeoRUDbw5
PyOfRnXhxXUmJt1ym5U7+GbErE7roskbiVDEiBna0BrxIzjCBQ7eCFfECaOS2WBCoYbZYotRDyev
qe9H0Y9j5Qqr1GvAGrIkD5G7eRwTat9XS2LnW8LQ/LhzVqCTcyUJ9bxNdHfB/Wwj8x2wbxofiMwj
wnYPWHEdN/6fMm76YebshtUJ0AcrpJbct/jdpAtCtBHm/LK+KucG5/oZsYB1MXBzeTiYkcnSLFjf
McyDA8YPwoA9EYYrurIpscbbbi2LEQaaxzMJtRft2shRMrdqQ8Hfxr6U4w4c8KnLLlyHm3jV64TI
/m0OSI37dQ3ZSWQQHesym1LzaPPfXI5QPAY8ZSUQZyaTPnKz/f83kjDxmnnz40XQVSpkRu7c4eBE
UIF5InV1geeR2J6q4TRueBqDO+SjnAmnPbVsqFZHulv/1AlSqxG1/APbqgKGQiN4LQJ+uLeSefVv
HWUsKmIgY9kbEbvrG95HAzqNa1tRZu7Ieybzzc20wChBB+r9Mq6MUCZBzA59HRFJHhPGZe/UpiQo
jmZhekDL6OeRMjp34P7NcI8mN2i8dF0rtws99KKdMo72s+I/9LzDTRBbwXL+lpvGonPVCTAEhgPj
foZvbHA7RTHrBXoOTdYrvuGBqMeONS8cv8nRkC/9Ysoi9z+nnWf+xuhZOftXKnVqoopiNLvR2PiT
Fm65gk5u6uNtCSmjxIO7J4hj56HcJULeA3Yi45giywKxbZnETM/aYqyb6/EA0V0+6F6LidNJyyRb
1NkRffPlbMpOW5PANZcVqgY3qsb0Y1F6Yi+Cn/oJKGPM4p39VSf8jkzyx8QcJGzMaA3lsqeQ3lUb
JMu5dIKKjjXx3IIXId2WkVqXWLDR+hmL5Ism/rFapaHC0m7C7h1CvwC5qTKtdzbwBwW3/YK6eq8f
xuXlGcJGwk+RTJDW/ttTdwScLCnMqYwAsyTixkeFHmKO+GB8UfIfan5/UF2aKtrDl6miAe2FPXjc
LrJsrCedzL9bMQcpTtS1jC4D8rtQ6+AxSR+IQdT/QFkJPnfoGCDlYgOHI4Xrp02o5Sx/t49ERcJ1
bw3bh1KKOAxqiEPP55I7Ytq3NnXHd/z8G2OP3IeK4r85WR4WULb2WtTHkPUOf9ZpwrSVN2FC/Jbh
aW9QkFuSbcgyuLQ7raNuJujgnH1KibhCMjQ7sq4D4Yj1AOvBDHOAlMblLMClafG8r3xve68rL+LC
S9enkOg2xuEI+OKzKevqe0uKyQ5MpWGoVrA0DtiDNiPPPWD/hH8/hmJ3C4TI3H7YFPj/eHN6ZvxU
c79lh2u9FZy0pbLilCfOk4VZIMD25Z8LMmsrUvxloKruPDoZVRXaj7USSAf60m3LF+ium5kImzAP
tKNDCM1kVKqz5M3XtOJL8iqWBFxzKifQzzC5qnrTAizJn+uJ+skWeYD3SVUQXTp4N7E63eWknty9
ftBrIkauZkjeECtcp4iFizgVRaFo0x6BH8hlTNdQXBEABREJNtQvkiKKHEwBBjMf0yZkMRgqy8ob
VilabNtUen3VPiEELtp3SJeQ6pwi9h3RiMAgMHCoFlvKiX+GX6kbd7RYc5xnGHJ1CN7/4oxkB6aN
OGydQR4WPY4ikcnreBLmGJ70n04uGItv7/bmqq27X61sOCiapcL/9FopISWglwbek/LFxGUtn65K
9g7E+HubrJKwkErScyau8446vwJ2Jwyg7BabgfE7dVJ/K17AvxWnwFTNW9txQF9t1KGDSO4uOR89
QMyGbuVBU/TgEBYA9MkSLauS7T7DeBq3lWGKSDz03ILIZqqjp935KnYJf40eschuee+PCVXUXKdC
3A4aLgQv5qU45wcRVAs9mO5PrtnlIdgkCFdyJeZxSjjBTjPjsY7E/m1MYV1l61oh/iC5HbVbLSSx
0CN6Sp9kne4KNb1NjOTRMd4y4Q7QMfc+C1RHAMHF6jxwvA9OoR+X3zJws+7c7m2emhCTB8715ozB
rAQmYSmwKhAoZOAOXOep85npxYhovBtreYa1vNtW+UvT1zJr+8daSiyBRMhoUgfz2zxu6sUX89o7
nS7aJRM6yhMNISXZLce624/gtxmPuSzBsm0AfFgHv+MXcWGRLggYn+4tXTovrtqeMBQFZjtFmCzn
PdNyZQSnvI787nIk0bIIpXcJ5hqT8FSYMjpnCJiHWhGmyVC4496wn4UAmZBZsgw7eEn6cxwBtGab
AteiKJeV8t+EBaZjnCramnTolD64+IssiS7a7p8qHo/pfDzFRGR4wfiIHOgXiE42HJhHujqRDfCm
g31vy0J/4faRG+Uktxq4B0su0MmNDFBmvYEk7a7Y5/H8ZeRx0AwVrk4fzIVTFOMg2wvp8XQi5l5N
fWjpOBttEbIpgY5OHWMA2WFECbDAhNFGX+4D29ogRCJu/bXeBOHh9+1MPUYnmvHlOvCVKs0yFUKz
Zwaq/ErSwKkXV6YVHvqC1M5hGzSRsXhJfvk76sEIiOpVCIL1zvkNLyvjEjX/bojChyg+cWQOFY4t
IPzH9wh6GmoJoxyjwK28qew8XtntEvGP4dbnoKJcZC0+ZQeBO3+uCGrCuHv7Oi8pypZBizKQ4AnS
3oL51DdOtYRUB4yH839nMN4bVwoUJO9GAP0l+3wPsJvYhoGsHrWOyYQsD1clfZgwf+LUXu77yXfa
MMUtey/RUwk5C7FIG2hOFaLcuhaCwKfy6BnujBfP9sBu1/6Ng1J/wuMJHiL82k35TdYAKIoI6ZBh
Sz7Cg8Q/3M+mVoW1a/TTXjy4QzGyx1TIH2nT3Nffgio1pns7gcQKlZNEq82aXIyWrAPieZluJNaO
lXqb3MBk/xO17BDKZeVh+Q7P+yNg5QN/axMlCmuqoEdAfc8QWDDlhUZC09Bm6pT/M9JE03FjbwgC
+TEIRVT/BMrSfDibC04t7mpW4n7EWLC0vDakxQtzDLNzN2aXDdO309WmOnEY7kbNbbd0WJGvkGhT
6Qerzd6yieEQx0V0NvyfaC+j4fcTFyEN/j45zH2Ur9v/vYlOyqBzOxysCtm7cl5Nc4Ga44vGFRSR
y1GzubqqNIhbg+MoH/6YmBW1crc6TNGZQ6J3hmjpJNJOGo/s5sHpPYv5RD0OUv/6Raz+E6xdvgM9
1aNL1yz2rhPS1/gcKfBtebDfyJLWOxfxhbOtcXz/PSBhXmlpZBSpsjxnUfHm8x6Hkhm22rTPmF3s
vMflrjdKxIPhEiYDXNaFdLrUZY03tS1bZdfTZcV3180Nc7+/M/iVxJG9h+PKQNJxom+CFVhVG3kp
b8oKossYLqmlbhy5y6ym0dxtaY8GfUvpr6Snb45C1ura09ORonso40x10TRxsx8QdnS/YpPhTKP/
ULohtddDyis0oGj69tdA68gCYelih103RQLCyfM6SPUoaDnj0+5kdit0Xqw77HfLkbjLMW/Lirlw
VJvaZqxAyd73YcPeBCbbot0f9Nd5jxpX5WLCfzE8tx01JFemRI5m3+E+3aubRCKLHyAEKIAZKeRH
hyKu8yp6QAqH4ltqAY7B7PuZHXJpDzVngmq9ZeOf3Jf+Y6cjwenigQG+StK7mnSuRPI8yD251dAj
euf7Dadgef1UvisGyJnDYsxGPnBQ43zQ9ZKvSED3r3iIdpIflVImRtE/KJ3VtIcvqeOsMviW3Sh0
KbDs/ZU4vEGGhuSUBO64L1t+GD1LzayQ3Lfh6VesaDA+ecC09gZw2/ZWGuLZeegE/puFUgKiQQu+
ZNe4kTBzocBjuRFFmJGLFMH8AhV2Nf+9flVioOUWevIqYnMVbCf58pJejAnzYC5fWyNN9qgAIgDC
+HPIeHuhxbTb5gHn9LPV0cG0ehWzOJL1NcuqvtZp/CLnAVHNUv+8+inwN6DGF2dFPRA42Z5QKZEq
e6iV7F0g6b/w7wMivn4oG1eG2lUNSaYMza8ZG3JKaGoIrmpZ3xQAH+PxylgU1X7n9d/MzG4pS/UO
uyPeAlIZjJc+YBB4/EQ12cPp2dTAph+0IXjJrcbf5ci84kqUfyELgHD0Y4tnQNFt2cMWXx84+v1D
gnhK3I5zYIcygibuTN0WpoQBmq0VZlDpiO35kuG9iTS1wE1hw+WfU9Zka9o+35ebYLIlKufGgJ0Z
B+WvnnmKYLxG07bpQ6X4DOzgNZwDvx+Pp9dMznkxiYyLw6Jjiau0FdpKi8/yf/L+piWfXl++1gE9
6+ckbXlz4TYe08dCdYCsnmOoeGbAepYy0XJEDdUfaHPozKeS0HgAt0/NqWl3JZfYV4XQYZBIkYzP
zbyqCxhy8iHQpOh2WJTti0HDrHzKqEqutTyFp441tcAFI17/HXwMN/DeNRW/oLF/tZv1DHpYGIUV
dnFmxCeSqTgjYoWYUmsnw5wxBoTYCA3Thsiet8onEJgCirVAuZ0nIv88IDyGosMHHQOeaCa5y+Um
fPuh6hf7YZJwePzUHMOwZhMNk5KaUB+hyx+BeVJW3BdbPK4QZsw+6hKLEd7jOltLKInWFDrW0neM
7Iy8/LOd2FCzCmqOWMpsHYRmz/0Gh1hx6nQPfdS5xESxXKSsMgWQViamYWgxkNokbrGZCtngz6ZE
j3iPx7MmwhlK2PO9VRBbUDq9Kmyvfsr+IWT6eDxw7UsjquiVhGm2AM40v8ffwHwxoOmczE6W2zTo
W54iegBIj2CxI8w1q1is0AjPC7NebyT3Bo2PtJSbtdAzKOVPjsmXOr7yKREXksWz8ur9oJDoEX+z
bCTJ9mXwQxQEsjuytVt+JFMTMwyLfLaERsqeG9E8k8uJcOZhiZPM681QEb1kBSWCDHO+pnTQ3AAG
lJL/AUxOnHjXWOva+L6SIH5Ahkh3TknIFBBKpV4MXsQ7pHW5/qGwqRJ+OswBU2PZpTMoh/mz/tfC
AALUEvVJBEhhfxqFbNa5+2LLedq9dicpOT6zhqmC8ZDf3ptcY7f8InCpKx+ScjRVcni13OWI9b8D
8HmXc0wQAM4bBmh2/ykhWR3oArPpiK2PFCVvSsRpZ7byyCE7rUehKGjgU/XNkXibXGmw+faOeOIt
NYtFhas5hGlGoV6uVqg8j8Gat2YXe5sY8Lvo7wYrZreDqAhLgzF0lMQRaI6+TBgfKjfzT+JXRBNP
eEtVtzySx90P8LTV0m3TfRUeFGXHoN0O9BmnFBvYBOMq00uCFt7cSFTny27Uuhv89esz288+nKAB
PwI+K3097NiPnF25HmdWsFFA00uA0Se55+Il/+HzRLM94mZfRRwpRuQA1UMrGsmdC0wPxdcW7qu1
INmte4tKlSzQgCneo6usyclFEotZpMdhysGrBw3xxnv4UhJy/1GaQuBBb+dBOHi6BXSLJMB79pC/
jDjj9/Ct87h8lanlfHUsMdzMn/GV4eLzaLWV700GvNzs/yXxVePVQ+cKfadRKCcmSPBrRDf9HP2B
NCYzzqH+SWT0ZZfur4aJA9jMSjzBp8EiPD+Xpj/tjyboeP+1rcv2bBEkmsZQ+ZP5znwQPhfF7Dtg
XC7HsswQImqDpuonlSC28rFnoC5L33h7HYjErmt82cmL9LSxnNIsR4/hZYiPeX4oyQpUdmTbXYVP
v4Tzi5sg2dsq7GbM7ZzH+zKXDvEAipTbREGzc7ak4Ciir81c32Me/fs0n4nUSAqJKZiq5S6S7dH6
HXYF1lZOAbvvr+Xv/vpGSKAeS5EYKzwnmh0QecFLSKCDgRw5TGcoReoCsOrtJDCAGFx2/HZ2RAjI
UeH8lkchqnexD5FWArog7r5U6/aas0V6I/qWyf7TNaxyvRmWW1PaQrdk1BE8KR/uCzJ2bkCr6BnK
pHgGF5KzSqhkTN756Cdoa6LX6ehjnryjb/2sRUxfVZM3qU0lB5Ti3nhyG9z/fYy6o5nKd2TjwkRT
+u8nSRQmrIbYai0fc3BT7Dnn27w4B5LROy3Ca9wDsow8LvFwXilcB99vW2w0GVCCqhxlSSzrW/bc
ThkDN+Rl8un7IIcp/JfRwhOULFbOZIXWLNHQ+eAQHCHOetbkpcjGktw0rK77wJeXT/hmQfpbsHaf
+4hoNurmEMxG6HR+/W2zdnv/ip1Gj2+e5jrP8TZ1hIYyscHZi1RqLgrm/yVIU97qs4u7sXZ/COvy
m4r7n7fM4qIrnHkJBscHirjHT+AaZOFFNJEuM5HeNsSQ0if/M8+SgDG7NYppAAFvNgReIGJH54w+
ef3oqw2sXzmaMwNG8ExocE4K7QQnM9iHNc5fzlwpIL3VNkh2o1WsVaTuRdX+/U+8hM13Z3kmVeVI
vpC54bv/Gl75hVuxV9xDOS9TozpbbW/9uKtt6nj6I12W8I4/xwLjbBOr5V9RD28YwsYjNrQElYNg
+b5OawrKVUi2y2VXyQ3zNffKmh5lu+BWgPfl9V69BtOWdEFZ6c1svkMf4wAzXILqeqVceO0ebU6u
ZCGDYBccR0DyL7Mv4y0Tszf+Hn6Rw/biWo57IIOl96qNiVwL/Q6ZI8HAyFNK3wrjZnQLos1KY7b1
ZxxK6dUjGO6+7FZ5arK5TuyCpF1IdkZ6ffrIJgDuooaXOSqIvHzdKwgP49Q9Ho6866qFnckvYD+P
ISt8In1VpeeI6ZCJKm6pyMkzzEJj9uwxOW1pc3edBIdiWKf7Xai+iobyFdR0xaMeHeqWN2qLd5n9
E8Z0YFuQYe0r/sZy9iHXZefN9bWAGHv5xkQ1KP61zM+KBBb3nvMVg+G+euMR54CREhkFeL9z3ZIz
sKWtZSgVRWBS9RUwaeM5+AXBhNzmf2ATmry1FtVz7C1haPqS/XkrRbSb2sLhtcncpeS3nKbAQzxd
PwJqWQn724as+Q7tQlACOEPtWDSdBZv67Y4btqpszaN3KPRS73X6OAQEZVfGB3+PGqEJga6Jn0Gw
klhjcNGwi3gFBBQHPxhQYwYqeQlsWGThkQn3wgq2MNQC3FEWrb7PSZ1fVIjIrL4ssME+B4OtEXL/
SBopPcKMR3eqMNMJ5yJzNOpCZNxfdYcAg3Kg5Xlb6hLdCy+SleTMt27+Qp4GDFaVYUNQujCvR5BJ
UI2fk+/2qlKh8E3JxkVPWLmg8IXyU5FUrFBSZSxpuc0xe1no00jLpjizgICdj3WndHWptZetXRYb
VrULndLT/jbJoqI0VnIL6HvOxQGu8O5DczIgVYYtfIxfToaszxTCQPCKjA76HJ+ujs+jOH5BNs+N
hlui6y9aSGIGRRAHcHMdGnbjReaoof3jLObGxrwfIPEWlhONrIqTtdCP70NQQs+LbyIts4FOmWgj
RxdaLwa5Fu6ZdULcUYLi7DrLwdysXrQkilVsrn82rN8mTGx+B/opSlFDE65UVYJm1sSoxVsSMIFM
V0+ZRvLjfbad1PspqcYoyEyBZBIk/Ol6qFgPKftYWQUP24ENv/PfP6epWg2qfP2z6+PFGzRzrj9r
B80v8bkkU2B3NIfQLvYSzuRyJecIfculUdBszBATKhd+mc5yX5xFbtq/29XWRrA4dpKH46u7Hc+h
/OAPLdYgrMVTB3fLhIjrpQUn7ZhC/60Ei7bGoFnaDXi/Sl+7E56zJ8MN9mfPNAlv0oPfJvZlTpPN
tKXf7yFB7JmT1DB0QJOvH7IEBoreCGoFI9H6318LmGMb6WBP2v6CctPLjeiXanu4vUUpiEeyZROT
60AUsdTleNZRUwG7ql+1AWV/44H4V8WtRXTOPO+tg1qldu+NSDoPEfUnjEuuPv3YgY+AdqaWAoJ4
VYmOuPJduoF7x3inW1HGdMHNq2lXV3YbRhhIcLDHPgH2TJPxkfiyY+E8zeU4jSAdUBeklucvpbQf
qIzAXKij7fegI+dKZ0Ja1WQ1ToRGTQ2fP1NQAdKbV3y482j9a5+JJ+AL4Ru6nMo/srhfpVhB5Tn1
1tqstVg9MyJOF0J9P+3B88w2xBIPpEpfMmNh8OTW9yHAxsHK9UBBl8OdTep+DU2sAO5Q/MWmZUoJ
F637T+wf9EEmgv1d6F6wK5JrZGi6R60EipT0toiA9OwzUPsSB0ojvKuZgrDn4tzrpbZnyWH+n0YR
r7zJBdWKzwmA1PK+oo209kqMbNuBuiHeY6KV7KUq2IWseXey/WkwRj+wmfJ2g9cMjdgwtDs1p0i6
bcrwisZM6tGKBmKanzBTJwpsQ9nydAGdwVK9q2a0TQUOPljGCPslL/88zOZFaxA5hwBFftghQNxe
UTYTzxJdfxwkd7Pd9o/+8FMeL0bK0eQ82BuFqjfvI9gBN9BtXQgaVS0+JzJLuGGFP3hh72/FVP3v
UXh66oxMjFHr8+y/Az1Bn9XkUADp9+XFSf/FxMuZQ4iPlGLv9EDg8EDWaNvaqqxhDdfoVjUWCCaT
xoZi9yHIggss2SmLQm7vEGFlxA6oeMRkY/bPEctM0XYUa7kQiuNn/SgthM6wheQxZoo4xttG8k+3
f3yNbAok4z3ilgGU+S7ZZzxyaMFkMpkjN2heZcI8wVpNsMXQfsPSsceTlC7KW5nI1s0l8pkD9uKj
kaVE5KiaEOZDOXIVp9zubUWSd2nPiaSZKRNQnpKFs7e8wV1f2LnghJhDW/DnvpoU3B3ARdUZ8OIS
neZ0Ccm9GCrMMXPNqE+a6YLkuzKsxhW1tZetc9jz2lCTmrp2NnJX1/vX6ahBQpUWhR2enGfaFbnV
0ySsIjpWBGuFCeSGZNENnHuRCAjZQj+nG+9yyWc+gzpFAw3OlhJ/TyeMC880Jpb3IVwiymqSgIm3
jTPsh3intCrLTAmxiOGUscA3bOdpla26wboPF5jvIpMd1CgB80MNgeQHASEfTiE9VpXUjqVLZZ8I
5cvHjt5EBtKw8TCs/dUMudjOGbcf9xp2RUCIUzmZ1RRWhKZJZV8IlsTgkHuQaPO8J7RGqV9Ysm4O
N7MVDtNc41XiZFN279ld2V+7ZOsnTUGn2N95Q9DsAonk9hxLv8abszNC0X9D6KBf8YXeYQWdX/0y
wLGsBeqdiiNN3GNSJGSPqWG+JWOPCbPdoXtWUvW07YAxXmDoOKoBP4fcqHKMxc0Eg/daVXlFJck8
TcIgSCR6G1WyXaipt7gaD9o86KveVtqZSxtoK3wFI65mPV7HAiF5wl/k5BAliP3XDIqkzWI7FRjH
XnXdyepGMzbKIx9V+d1tdAD+nZzXFG8KsCelRxdkMb9jfMY72K9OVZqUDGJCagYv2xF5VWeWjweZ
NNHHSo0K/QS6A5tMLMsnxbntD1KCS6jZ4mRpVREc7qdkuy4dnFh2m2KEdzPjOHeSF64YAne+qJR+
JwO9TAsYsFzjewpIOI44oOoOl8DlKlaCsLFzmrzvAKa1nCA0ORgOwA1+HXMPa8oHQgJiUuCtr0IM
lNl4APfWlcA1sggyQ7Bq6ceKWoa1w25xMVKlUV/XY9cz4XTu5llidmAiu5YdQu5uxiKQI34olxcX
Wk0Vx2QVI0mIZsEsWSG6brQkjssKpHln4RnuysYElPXA69uJHchp48uwRZ/yapuQiWbFB4S1Gqsd
gbQOyBfpwzcvfvSrF/WgOitHVSjauAxoW6wGK3HI/+JOC9nn3MIHBQLzOXBdgz7z1+0WYPVzOEBJ
ismvbcI6a+8GoB9lRMfJ0iShCPfFOcQf2poOZGMicDc0kuCWkI4RP36LrGtOUQehHgoprjPWw5k2
VIhGfXoSweTGIgQ9QYl08JzgFX4rDnjscEFBpc7PCBX/mWS+ODoP5jlEaDWxmYRjgnK4UMERHxb5
Av5l0SnFWlSGSK+d5zhd8QZnuiudeCU8K6vnWBSQk8RKJjEgu+AB+s/B5W5TIZk5V8jUihOf2Foi
9R0kNIGUiHpDEMS2eOzmOZWfazfXXqbV3lUwClNx0bdylP6JeDg77vMvfmIWMd034QiqpCPNe8d4
GqYqeL2kteIhZG+7xVnjU1/7P8AvFfvei1nbe95CGbxRhj4cd1yy318kQK/Yj01dbTaKjjVtfGdx
91xHr6Qc3dDW7t3i4rvajXwcO59XpofRSg/1XPca6EXJ0TYbxDI7UILgUHY1McNMnXm+f7RtM7Mo
ooW8LAzxwZCLVpqmwRPXxzRep/5aMUN1OAP8xaCJ+3OuC5gsRbbXKLKlXTT+bYCGypGgYGUm13AQ
WZh7I9f/Tna14b462eqcyZoWHl/z+BidugFKsNC660O8ajzQzRyFrQqTdsO8q6Ep5m/PdrcGDEKE
HpgDyCEWocixkU2Rtuc7UGcalbp+YH15K2W+rKXOcMTbjNqoJhJwtnGIHWciB3T0qnDZUJ6OYHiZ
uMeyjPJsydpb6oCZS5SEEC9SbNNC3X8EB4cBfVLwYWLLlo3GTDhqNaGoVYtqZQaQM2rFqnODmIf/
SNedrdQhnIm5OF/oukR0pNr8zxnHQLnQwIYrF5t69y4HFYuR7UHw4buwNAolCHsa71iQ8Xqv5Q2C
kNJ5qDldCl/kgDsEpn1z3Jp+uq9+XvwHxkgF5inHxzMWcjdthIlGF2hPStWaypXYU2MX62kZpDky
+bQxJbK/x+BVW+8FhIbv8xFooy6pP7LWvFI5yeFiQXQMBs3jKeJm2ta8e3sgh8DyobChgsXHTZ8K
eY5JAtG+M3LfRLFvGfW+X2/nALmjHX2vNxb/DRKI+zO4SObZUIRIHFNJxSRRHtjodo9tfeEP4TDt
1Mlom2k72PROMQGvBeYVDuBZiPxK3PsGLLk94NzVTqxWZYbZ4Tm/n8A8L+fJn6lTQ8OHx63HGwNd
4sTkcIxpP3bCZQYrCU3m1mAFRLd311oZTuQ1ma2sAL4cKUDHSRrUUEn9Wv8aFrwl4w1QBNvXWTFl
o91QiERbtVbMcOMo2HME4S2bpd9rnuXovkDPjZYMuZNDYgH+FLjKU0kgViVZGXuMFFMtV9tbUw1+
e844Pm+6Jq+OE8yAmbx4guCUAjwMBx/WojFx0QvmYa96BEVo1LzteNojGPLxK/TdP/iVg+hvAI4F
64rfyvY1BkvjN1T8agCZrrqfcwA99OpSG5YbFfb2wX3yL9FBMcBVVPVzG1joJpizKA/piuBYVjpO
LhO86aZYgK/hi5oShKEMqqz0CozLYhTiWhYGHA6smqZ2YzszzVbwb8LeYnRUZalqlJDQJxAq79K7
3SqQUc5EDJN2vJabVulKcFXYvymDaoFNW/LqKSRZCShJgMmGMwWmgp87zkoT5S5FtOB0gbmuoFyI
PXxZqul/2SzopB2lsMvQuu8hy1RWlTHSFmz4IhBWqZO6bDcqy9wb8KR4Plh0qmgyLHOcDkZx4OKY
8Vr4FzoDYACRsazif4YcBzasUPwjCBUKKKIGTjNm8gWr+EJNA6cqUNImr1iPtvokZtqDSzL+Vg4O
w4aDauO6jF9DOCx6tea6aTZxHnfNpR1S4qZjMqWrndx3qL3tbuPsdJr2pcZS1PVfP4I8mXszxp/z
gS4Y+dUQfqO4pmdAeDKE2lpgNEwhEx4KBKLATbyJIcrMUyxNk9mtDRyj8NfaizO3QOcQzL85ojRi
j77rtFk2iSMo9Qt6H4IPzN/X7qX8JrQkp2vH+JMQSEjijU2m3ksF7vNrQiaDZu+95+R1h2aLV1Zv
BFWOO11mqIRinWgxoSVjZF/ghnhWdFfPjjCGVDJeRBer+7OQSDZlKDR4ayjhZedqXUE7DS2B9as4
G4JudQ2QINYBzKnC6pDCFu+oLpVIN6ePJQxHvtVdHMQkMERr5FCCH7t5sb8jhsxD/jLuEQNnbSKm
HfVFzzPkQvXFVeQqYz0LHL3ijbJIRAljEw7/EJYBMasysZChGh9P9LJ9KaxrOYd3zkGQ3fYe0W9k
5W+JsjCzPvRmvgiMIoWisDwqDv+mLqUxW4hqoMSaUsmQcVs9ANYs6KCnkdDx6auvBVkvlEtgCyT9
u0AhgW0y07RdBSMQyPsCwAwhc8dwJYSmZOLJjxS1ync1CLp1rXUFv2CYFwkMKR+9S7+a8xx5wjim
WJjvLqbjTt77OTrFyKdh5Qxv8aV3popLGXf8SpvhayqLDkGH4MjSus8L8w6ErLFs1n9j+tJvCoos
Jnig2MQ4mSaM+cnO+bOtFq2IlzjDeRTychOGgDy+lF6i/24pJxFVV8HXnaMeBoNXhXk6bGpq9jfT
4ulyXYgMjVOzB3l96aSc9DciSxIQ2HBiblKnjKnjr9Ly9PpmaqShPVnkV3HFurDQEcc5FgnuSIrj
zpZbhs0zbYDVUUhBdf8aUak6Xj3y7oC2g9yYJyH+FcCKtW637uolSKLyqS0VuYxS1louL3rXjXzM
6k2pYiCri+qe4xiJ7OgloV2S/+fGawxpykLCZyn3nQH5daoXYkma9biOWx6B9DL+szupFTRXQoNb
/I72mmHgFlqX2XAvr1xJtmto7sQizt4FQxh6t54AgtwDh8ApmPPHdQOrYqBhllw+ryhbaDDPA0GA
rCKeAqiVG4FSdmL+ceBd5AMWcN4b3jmmutOxyixUKw4sc9WZJY5yAohEHPifFIAzYNU9o7YRkf8e
gcyc3JXu+BW3psTIalAeDMRSLbXOFOLsuvN9FmZ6up4P3cn8MQCiY0r/wSt7vzoX8yTtSqUGq14Y
9OPnGTF27f7mIs5zlk7ze9j5O9FufI21f7KASUN24HdptLrqGrGIO3Q0EE/qLTLHkbu26p30aBKK
DFd0Nr9NomYFkyR/yMGGFfqdoPEtkAWW2T0VyiQ8nDPrdYQVPYWwFUNZCA4N/1rpCRz9UWqmDBMV
KMTpq2Sekwr5XwFlErAxZkX14IKqCgl055Nl1qQZmJXnjgpt+gI8PGaRD3N2EC2tTHVipEoMdWTa
+UN0jKW8EHKkJLbAFY0Okftp2ZyPzXLMbYcJ3dUVUX3dO8pwEA6aZgF+6jNxTLhjqjWg7eRBLgF6
7/TGtmO0zCS6k8h87JUStA3fYuTwgdjIzUDufaceP0fK4nCWeQjz0fMeiAlLy4qk4aJB05qxtVfC
Yvq0ggE3Wl5M70W0V40/NJ9ixClMblbg4Jc4luYid+fweqLNMOX6RAGxKpROstbwfe+9nFVaix/m
pp065nAe77188YvAY9CXMhiOTEMLcPQTbIT7m7JdkKXnJR4BItoGjY8yF9UTFPDVcwoimPuEJ1e4
6SSlJeeoE8VQGuvffnzQ9AsLm2iLO6CowEJkEYEY/z3xvh5FRQfMBGuje2+lHBqJaV0QVPeWEoYG
/dpB+ABeIiMsO4Xm99V1Ntzbh/pXq/RUFsbkqRwO+xaZ5/9Qcvgg3KBY/DMXLKB8UlCpiXXVpgSI
dk9kkk2m/7F9OAcEga2iT9jvtyBiKNTZMDuYekttgOgbT/urL6AafIiIgE3VABR3s86LyT87om2v
oWJzLiycybFi+0Usv/xi/XKX6mvC91WBfKGOHWjhvf59nDmGv1Vz57atp0fGFTJRXY7/FmcOIvwV
ef5zAj7WIKRpaatNGkbp4RYt8gQX00+5dfII0AxdRKqcHL/LyDfHS4l8DweH2b5HG2a33MIQ6Kf0
C2KXkICbZFsqdvE/BJOmts3jju02Y7RIAddRC/ZLaFKuo921fAVZ0T4vL3Qnhmg8ZSuXn0vJ9Gy1
03IcFYUlde4XANkcittVDk61FWx7jzG/uM3A9yVLABH8sBXKcymOmOxAeF4JDzBxkQ4FVIuoKuad
zJG4iu6mJsgOrNqa/xcR+ik/YeVMpRSMkqgjrVI7o0gjslgDoogSs1D7ydG6c20RXpYuAZDoskOD
knWL/HJ8WlGToM6EPK0nhxFGmjacwqcsuGrLVhY+/b9YLTtYXJwLLta78E/eTH+XV8AT9B7BMM34
dqb0BAf608jLfnaOJb6uG/PMEv4g07MjeJHM8Wlv4159JWX3CSiS1mMjFJo53pGe3iF2sTQ986Fx
rM+n1d2Hcj24wkpEQD4f3VoTRnqodfdTY0gl+Ju30R7908YD576uMSTbNZMWbwHyridbXScEATMf
Ga8Q1IbnzX6gJMBE9wtpSYGBXylSqBwQj8f7mGpJPHeOS8mFVYDJI+2XO1dhoB9dH0IWIoSf0M78
ghGVEb21znFaqfsz6eKS1wxn+ODFpb/r70jA7OvZL3PLupVeIEaH0Oc1vkIPyoYNcLSzWOnL83CJ
5Vgtn/pVZZpIAxZSV4JaDb0HaG+2KSsTuSh1+N8ebZgISEVQGckdwCLqXXdjVz+MgNetaJREc9Cn
dtm5l3nSCgHQUAA6J/uCimt7P2xALCpd4j1dDFx4km533sKOps27/qnpWXTWZ1Fp+ToFv2TkLwiJ
6bsrmX4+CFSHbkCfKGbS1hwpeY1KdU3zNdAll/EQoe9hx6bjbp1+Uqf9eSvoMKFaEfmM+J8Q/Wkw
TBky/iQTRxbMCmWluuYhFxH09phzHEE689kq2L2D2IleEMIkujRaEgyYkXSEWl6jASOXjMKREuUX
PHrBwoGpTkODD8pQCrxcR0IkruUSD+UmoAiIadLQCOnOi+P4s6a42sOEM0Um43UvsIxJE+sA7qTw
7gzKoJX8AS4lx5GVUhYTIqf3TZ8vPH+1f8hMFhVKyNv3cCcNza5X+6yTO69EEDOvFMi/gbWwZIPP
owI5EnZbbn07DW8bmunxUqGc3a6vWRuAEx0TtILvtbqHNL+GqIYKrdM3K3y07BwBS286qd9QnwSo
N1K6/Pld2QKNhPIfUFdW3PZiIz/qra9f62Zw6DlANBfl+OVnk6mPmzUI6qcdUNzkps7VB3AVqgb2
in5JXMOqcQ+jBlLr7HW8xPy86z1hcgdKxy9f3voVTtlMXFW2VjHTPYvSUaLJeEuaJno9X7vVrQpb
nZd4FQjW8JaXb0tVDxFf27vEU2b0L3ZTwAvQ1dFgJUoG7yinz97xtMxZ/mxjHFYZBa0OMaIkc3xP
IZiQJCof/TMj8oZZDqmYLijVKza5dL1yKI4M/uO9iwt+41GC4J/9ZVXajheO69bSAc/ytM2V+5Lt
QyPyDxghFpTKy3da+Uvn1dMO99iPetqyh59pZLvuXDBzjpa5jQmdcBHXVk3XP3m8NoKn6aRmzZGs
4T5T0fqog0hU7xUI4CEOXBMWY1RsnQCLv3zV/yvGQrPqBaksZZFku70YNc0UVyZJV1+KofJp4QOy
nUM1UOuaUm6kxL/bxqSVwtUxTPhHD4hqflg1IDa1SWw24Bj2UDkzQAdsQLh22pyj605ag8HEibpZ
Ld+tUd41CXQvqloQpAKrGEMRaPksbc8HgXTD4kmo8sT6JcNTmrnFtfpzLgP0wOU0azVw1jtLuUDH
YXHa03bdN1NA0yk4NWaukIH9oOZkcbWnkYEqUN06rIpphGMpa8pTzhe20I80AJ8eUye2bZULVt4n
NKqzSOZf0y1ZUeEnhQ1nmca8zgJ/gQH4AILi38F9WKLW5vwfMVJPS4xRZBaQyWlTTVOAR16WTYgZ
sO9476GRpuk5m+DmbOFoSgmayfjW0Hu41Meiiz9c2B15PE8r6tKE8CmhAfwr76G8BCV1wS5xtPwz
M0RPVvz7KBom4pRmr5+f6ax5ML7O9VMe1wS4MAiVnIJqlicQ2FLvMQKBrxBmRbzWFDoHPInNzKu4
G729QneeD+Y4PNVBcYTn5wVPc2KLsZxxpvZIFgrL9zXZWiwivluLMiQGvzkNnog+AQ2y4wOSCwcv
CEXhqyZByXqbkm6rEfmrwikkQzWmRPCvLhiG9FYAUJCjZ6ZH3dPEac1uhZz8OH32T85ZuoVCFCAR
Yb1mpRVB0poc+ebqdZRjKab16voKY/LR1HXG5ilVH5jUDc5WH647TIcyPkudlJTeXmfjc+T1gvAD
ypGZoW/cgQlCcTe+JcjcImhSY7VmOAZpUZsmC34Z48Bn1iK3BUaT8/BK/DXK4Zx9QwH2pcOrQZ3+
o0yhvz3gkRLUrM58GGFarRoIPuvyVrEFbfd4TNQoh85PvBTnX8Mpcj0u/tXL5nuLoT4y5Kks/Mk8
4XlubND2zug4nsqPjutLqL/uUgWyCvvToKd/fIGMzZKlIeUMUNOY7rhqtrKwCJHpO92+gGwyoitx
ZKuVRdUmfQlLd8Pb6NzKjynmfZXXnO0P44iR8gdMIBDCyWOpx6cmKgDgadCM6iDO32XM5oyc8W0C
6datrcj2kqu0Pmqb+Ob7HgU0IgQvdgPOIIq9wCPcey/lvhb2bC/v7LOtl88m+3r8w+Ae+AchdYI7
CvO+PJ9zplJFOu9pbowCAeL1KgL49LFXyzhaGD3Qeux9X4H42rIMspvNKrg0iBDE3PVIzQ0ClwaS
hcxdWUHecMU9pp+D4oaaxC7jfEGcycZnQhKWRQIqvMZFxbpVapBNtVC0aVAQjMIGSAsTFFSu3PFR
PHqTeNTGN8ZjRKr6jFuh6zBiO2VTCe6PRNU6fJqZTbjM+je70fHD9fGrWemACUpT4Bfl98U2S6oq
QtVz+wb3iPCpvMp2U8MCRDCyJA+A3o3qW49ciE5MLaSCV9SlXqUp37Pbx4trqsBfWInbf3fRTORd
5gEQGdgXlZfGJiLxGLcdW+nZc20Ie/4fyPFk+hRD/4I4ZFWVz4pffYbrWMKak2GfIkm1Hfi/ByEe
REqd0/UV0ySqrUTbHE2iOgbVY5FLJf9ttU+03nqXF5+VMcgGiighY5O9jdJ7FR5QM8ZlsxMh9RPK
Qibx2gEfQzRIWfjojbMVje9jgdPUy6lU1VAiVrjE4jtipC5TbkD0zczNRivnLa8FYTfou0Je298s
Ll4rCA+k0m1a3w1+juQT/dYxLxNmqn1Y1rbT9hK2GwQAkybHY6tDhRVR+sL6no82EPNHMtuFdFDb
UKK6+ZEDKDb4IGJZjJL3jeWfJae8O9KLeZp/1HF9aILAEYqopnO0JAOFfj1eXpQemQKOEKu4IQmB
5VRl9IIGNJnGITi1GlLasPLksjPAzdGkdqTc3ol75uZ9b9IK1CYRXTnMUTLxZEaznUflJBxC5Kb3
0Zh3yjvP1dVahIzdHZJz5mgGxxT5bDJ/AFPFdVA0BpWmCFkhRbCGGZtAXBaMm5bIPLPGoS40z2be
W46lvRHwjWoAl+FdOXufmCxKSgWUo+amNkCfit1ow9uxo88SSsHOcRUWvrJkP0aA3jXkbbIOxE8b
AEczku59AfPaTysz/cLVxM1ivG+vqX3l8G+lZaL+BDlp2Wzh4ZO+vvo7y7iVGeS3ZOtWFbUhnEpA
nE4nF+TR6vYXb/plE36h8diCu7JSP5vE9NYc3bz9St0J2gAb6MctvPbWysHRMyxypP1KwzRhBSw3
IoP4QOjgGgUKWX27Wd+3p3DwlGoYNsnADFNlgjGU2O2bt1LVS3y8qGZvmhlQILqibVuKTIcMNNFj
StpnkjqgSzPUTO/Hxfqz8OjSRb5zoXaRA1IfB/GIcQ5lNUbXNPWJTwMXoBNI/MSTjY+nGXpqVWoy
aCviYJp6UGAt9JIdVUjviy5bxUfkd76F7tsb6kARKzCtLOZPMUiMKErOgfCi3Yh30rwL+YjwXnC1
u3MvC49MoLIcioS/LII+qCLDPK3PDQa6P3HzacMfrOyrLerFVSdRb9GYc6cUAsd+i6+HpmZTZfWU
DIj3TQTojyqXvMHrqZe74Df4lwGLsOQCJVSQFjl9nuI6F/qjpOynjvE3L/vXMVgGBgKJ7qtaLWH+
jUs/b+oeNO/cHyX+NpCgKjapjq69d+w4zPJcBgbd7fOmGYSIOCpe6Q7bhyPrFoMzC3VwNGu/EK10
jcl2JwOGbX9L3OiGPH3LPKdu8RLmCe3Fes63yI8uVpgro0fUM4Od6nudsaC/foABIXD61A9KHM16
O35nIR2I0pGhkxF2NB1yrShSQtofsD/oq6HaZdt2/tulbm9HXt41RSyI3Bt5Xl4KJEM23ixE9bdH
K51nM2rmRbzJfgXPdbyi3FFGk9M1yGMj9Nyz8Nbrhbnxn1TqlhPo5ua9JtqCSchLPkolSAwNAFUY
1b1DPuA20ChKmX8al5gpg62oyeB1qyTmaIgYGrB75is12s+8CYi/sBifWjDDx/Lnsbu/FkcY+lfk
W0eIyMlSjlEOoJ/zdYa0xQeipl7l3xRrHj/5hB2AFf07roMb5TpfSzGwBYWYYRZmU8DMKxYE8DAq
/Bf1a3iIlLAiCwSnZCvozrV1J1wwoxrxeeO/ioAhuFI/6/pmjijlKyiLLwGpkrTd9frp60h3gULW
7gitSqsMjTrTaFea0z9/06UPxENizpcLEH4kPY32FKRCITz1+huGQ4uKFOSwoluKBANaWEABGY17
fhSt6W3b6guk1zDTAfwlu4GwSsw3rsPK8V9+5M4VEMNTjp/7HWkDw2DtQ6POQElhshYrOf5Jjp2w
/pkKeuEL1ZNsnYC46KCQHqSF9GkRrKwTFg4sq84MauJiHNbTDeYqgLrKD64JZkGidGGtIQPyYZqX
UtxVnTey9yMrKBOqnthmWpMvpPEW+wjwy+rmo/fR6ZvZjDF9+aklp9aGIQE7th/crxPyJ61eAIKP
Qku3zJsxceUzdSSWv1iOgYzE7Hd9q9/YqrBRutXngZOfwap6Ax1f/PHi2qGJpozZMr4Mrg72dZor
9m7GSbvkOuPrZr9wJyRl6uzDVbI0yaeljr8Kw3tnX/kcsglSTN/5Z4iGClXgy915eVpj52MlquIQ
C5B95ZHMR07I0l2m1IBNUkApHXsW/rPnSSSv6P7nQJG/AdCVpUZdINQ7GF5hbZ38KRPTZ5juIIGN
xlBQHvVYkdgpCyVe7zm03kSi+aWZgG6AZuuzbnuVuvm8ne7T3CgiRj85ZLO9c1s0pxWXgOSSmhuR
gppGakL1gSBNBkuWbr1pGO+ewXpX/GNj0u0QzPT0pBRaYhgWIq/NtoPSsidWe+IUU92EFufYfiMk
ZuGxMVLZKARHyucG+4u5Cq/ruVhvljyFz94LiNxK49VNT7ocdCKtB4GMgNCTuDx4NRvpWIuMmJsG
lsHna1xTKcEpPQTMgvDJelP4VJ+QO9uGUlwkq8Z7nb7mgdXFqkl/+rPAAcU5PxIQYStsqfQUPZ62
SQjYnguO2OVpak1SJXfjvUNJixOSQCzZwgcs4uxETRW9ErkI0kWqDurH2l9/bcJavNJ92LUB9R5L
yPsc031KFCGMByV7jpgRajU2MutCjX/UoRFv32Hfw1WGNG3IrEM6xudJRpoAlqhYvLnrjJY5IgLk
36RAkVGuflaFDH4Ao+KJwDC7J/8Pza2+EiX+02YxaZwrx334U/KyJXuFFt8SD0YIQp7alnn/g/7R
cRDO3dB4mDp8iDnHQ1nQGg29jSrPUwLu9sDdyEjYMs69C3xN4ZMwxTg7e1JqC9YomMHIiSriDfif
kzXNSJiT7z3YkqO2CSDaayubHIVza9vV9Vq4kiHGbSpgW+Po/KS3HySsnC7MAkKu/Xite+saJb4t
3Vqq1zazZ/OEusCQCJzr1Ys6CZp1CcoMJeDNnIbpACNN/gW1Aydv2dB5SKvjxpFg5W9MvGb9q+7P
wwSuyWTc+xOhNHetfaptCFyyoHEJbCUWIXgmEFpSGpOR5FaojWrmmyGVJfzKk2K2n9EDurTxEOMl
zdIyvq49put/D/lYPAFl1dA4/rE4jij5mv8ef18iIYzPUBgjme8hfKlDfKS0KnK7GBxSsEnrYFjf
EZwjoTZhRtx/XQXrMC9lN8PFM+WYxGi/rflaoxKKcCdy89CTO1Xp9v0cIfSSO/3zjyikCqOpom2B
wkxtNBnIiUw0vitObfaDrlko27RjjRHJhr/o7bGgMzwB1SLoSS8DtR+wvuWUZcwqKLpSv4NulhEU
8/VrksZv1BI6kmRf8uuvdweFhrYVaafGUo7yUsG+Y3sNhhAZSe6f89rz8Q6DvSf83jn+6O3Z/AI3
94Iqui5os/s0L6RkNu5jMNKLcebaHVolWSch0mBR4JAI2H13RrWTatNmq8v4z2gOGBFPqrayX03r
f/JOMelKGC95aQOf4LSCoLZY4SspJmo09PbihgWZXVMxfT2609S494udtqcnURI7iFeB2QjdbG+0
Fh1DFQQ7bqN+g16b/iI5AcGCadb4nrvgMPo1eyySMZsVQoIysyJc8IWQPJscnDIKHn4MunIqFuHZ
tvxcyFvzJ7XytAtPEVdz1gLJ/V7oDCBRgaWGbfJ6mK2uaTUGJCCuTS/1DdmYR/GErDCkyvseenUH
b1rM7dpUJB5+3txqQVbkprNKaPM0jqUeF4+F/aEpaztNpPjv5aFGTTGNdMkspHrQI6Rt5FtFJkrd
FnRsdZQxyeduTjIvEfJoOtlRm522hozH+tOzlm2wGAGmVTA0+BPgv0kSxc22qXhWRcC1ko9QrmjA
oijrsmx3MfMuPxzwbS1TniNFkelMKOcrI42gESlSh7E+DxVyWChGwYNcxBXzRjx87iapGB20XcH9
RedjInRVz8nADfGO8sVYUSeBZHFJIP6DDzkOnrBxQ77fAE5t14n7qvwmhYyOmSS5UpHJugvUAQ/L
s0D/pPRw88qvIxK/DuL5W9PEEUFssiu1/9wGvhIO6AnM5u5EgAhD5kY0UhZ+4iauC6tUj/pV99vY
t2Ox1CCTcYmKWxFeaVxNUpmboj2nk0d+eM6q5jPB/PpGs/8Kq4r3q0YFKvog8Rz+7097Ai4kLBWh
Df9qe114EnqEOYKY6j6Mryjez0qSXjoaxfFqromrpD4pMGTotfLbhcJ7/CXsd9+P58qBK7jvTnl5
TWQjYVE3ygCCiugc7qVlLu0DiHTgxXg/dQ5hGfshgG50zIVYrgnfP5ZC5FmVREIf8NFRJHFTPaCz
7hABTW5cq3NiyMklFWUT5yXAP5n57WQsMt7Wc0IneY/2r2H8PDRyboVXBpKTAJI8lFv9/KDwuxI6
ei09OQLjZ8Tyls5/TCk+uc5Mp5xL6TzrWqvBqDJtsyWoFGg6NJfa+BqZ8WBKo4Eom+Iy77dbrCXW
+4Hh2YR2lh2ye0dYO1tBC3sTzkAiHett4m10icA5OJ/gAIfJLmSLzifz2G2mecRrrvn8njGhTG62
U1Vt61CF7lvWMtyFU0TNFVzt7MEIs/mK8D9ULDQQsdUzzz2zNiuI3ob+4aCtKCuEiX6S1ObUX8W6
ce72YctuB8xp5PuqFpI972a88lnPdbLq/jAuj/nOrBYNdan45fwXhNPJh6IITMUq+UH0yfKxHteV
F4F8Jhks5Xm29ASbw6coe5HrMsAr4P7YGbaP801ghYEFMBMo9T38VoNuYqwUTvKqUAUIibtAxihC
rq/Eyt8xg/AChdMgao1AnI367n/LU0xYGYFH2IKMAdFlRBMF/TkdC+lm83YKAypVQo0r1/3B/xSH
WQB+tPPCTYqdOGISHf2Mt3BIetkyCffvVt61xdXw1fa7QXYlhMS7F07Lz3hmU4ysHTZuYA7bQi6N
MwQuK2LLBa+2c/hrmjpN6B7Udv4PzLR8FCrBo3u5hBnt1bjQ2xydnaomhsBxLxigWGAq9JYEBTjl
ODnDkASS/em1bE3cHt870KSHBwNCyp+Sj1UeS9bFnDE0nfKOrmGHPuyjbf6RYqUSbxvcaX1e8FKB
3anThPZYFAPE30i1wpD5xLVawp0NAiDhcxQguKAaVqcsjrnoxbga1fKMknY7WY1q6taDOLj7tAzl
iGM5RXXPoCT7Cl8rqqXx11Cx9o+nAySr/d31OQnX4x3cjDP7yQ1gtmwX5kyE27sx3z1CkO9cUeKd
cCXpRA4/90WCsRdwY8gnhNYn+Tw3BL2IcBZhbZBXLdVHHsfdnW2Mdsn08mR1iQlLR0s0d/dBeIb9
nmhD0Zuboa3V/gh7HYQMtsRNtcO/u56eF1qOr3ri3+0MIz0xJZuYM8/uXZU+tAlvkevZ6qONg14R
K66XdPXIQnQqjTjRzw57PmkFTAp1w767B8KBJYiki12TbfpHoF6PC9NiBRC7P/kNr4u+fi47NgrZ
GuTgW7DL9uh9ryB/pNsSjks5XuWpweMXw750DXgt+MzuElXXLnWvA/SpB1lw13lzJAIWYdY3VMk/
yyEbeDdwSoo2XtcqpMvMp4CbJNkP33QpZJj6dYpviAZT/ILx46/FwMevhsRgwzW2UGYn+TrQ7Qbk
0MZb+AX2sG4bWIhbMpPYGWWxqN9jmm46vqN0lIwthlfQgrKJJgyQrZGAkDdXBrR9mfdEhRr8l+Hb
7bV7zF7KGr4ctqyw88C8sKjynB147lz59BsedCF+UtYv7EY5G7Dxkeh1GUxDct11Xr5PqvUlABa6
0J0AeWxglKeebuZiphlHKjzDdAuDyPGse1OOfKm2k9rRIt1eXDI8TG5uNjDu2NSYEdhLz6oK/6/R
tmDiWno2gDuX2wGvi0XPMPr4FTT+XyfRNponN9A46ZpajHwXGnbEoiLDhyD0Cm4AFcPObtdo+gAd
2bk+Ynu6J1ry1XjB7L3l8KDcXXnWCFxInKNz0oRZ+nYpaOS3nMgX1JlD5x43kGLuqkIxY3Z7bL5b
7ovODqZs9Gc4zppvdhlJx5QEi3v+jLwRD7DkoCeCP8Dj2mr/Fm7TZJl0piY5uAk6PJI4srt8DFMR
b/wQIvOatiX940O/5g/fRPRUk2GCCT/wL69KcVzTKA7rF6i50nd2RIyGNlFW/mEStoHnQKpXJ51m
5hPvOBJK5TNtGZGQULljnHDP/5K61oOONeJWhWFRJE5HfF9osSgDMUx/ATtmJB7uzvE4paQKGEQN
ONkvAakPcDm1sx1+PDT9HBGEFDyWLT+bA3PUBRVQcGA2R8yiMWbyfti29qR5326ZYknoEHM8BfYu
Bn80Ym8tM/Yx1xVzXhs+qM4iwhnAn5hplujBA1ENTIfHG0puNpGHL8JQVxs19Od5gxdpjZphLjx7
KtoVGo6ITtC11VstYC2VSSebWo3YTvD2jLJrPpglrboMMbm6iAwMV3r+WNy1ssVuB8zvafQtaLpX
grl0hgvAIP4xXi+bX7sa2O3Ogi0RNAcngsrWyfcOxhRcoyV930DrV5iTSVU0Izw8ZWn7ev5V5EYg
2BKdVY44LIGeGOmOSEOfB6oHImxb0aSIqtmjCC7K9YtJNBO6uS0kPfrSJuSGcnVpBsUslj4sZYnm
MXT4AxFa3mxCW9jyF/sLk6Zfj0gzQimTzQIoVCs6HfA5jzI0YqYveS/be848+6Lyx/v7s8LRERse
gclJVPbFQly2e2eDBNqASQTj/yYoUcXNCpL9vKIoiVtU00Wq7umPs2us04WmHKNm4UgP0Ak7ldA1
nj7scOVNZ4vemLsQSPGS/36jUgf3DBg1N6K5Xzblo0I0+I9b7hp9LDudw9qegNjsEE0JBL+t4PRI
WLmEVn4hhvxTr3WtAE1yzABYZlb4vXf1Gr6N1s/+1ZglFxotrzRy8FhtbYpa0H872wfn6yQsNGh1
GCZVKSx2mSTIqe8k8AJlpIe6qjySYInFYVX1t5w9W86HYW+L8PnGxk3VK5DP1gkk8odu3NCeohsL
P5YQTEaW44IjIY671QTXUH5FcQsk3zzSEIIrl0T8h3SVmgvi8i2fkXyq1a4vnZvh71XiXzj3KqHI
i8+c0nEi2VFKVsPuntzOsqJBGBcnESAbjSXuy1Fa4dW+GsXDiB95wYv6RBFB52aaoYxVpWfUrS2k
w/Sryk101HqqEkBet4jKOa5qPenVmzsu9cY6JpjuL2gfJ1C6sTadjVFIsC5Ufno/9a0dK8F4Vw/c
wwbwtzD3n7CfQJgfFYlW3ARPCsfa1N5khMqcrjNgd8nDC1StZAOmeTjd9vpwSS+7pJ/Pii0mIUeT
ezhmSeZ0jg0flvdVTIXaohzhUbdlwSEMEhcMoIuyRtBUdgVrO0t0t8E+5z1J1bjZ2h+0HzZxmhAN
wpk4lBCKxsGOFX+8dxOwiRcMjNupOq8Fc9WZhUI1cHQJUR3Jrljw+R7sJHCNlc8vRq1d6C/rpjWj
nZql2mdAW6YKdSrkmbT4tqhw+LpD7UlDYcjz/PD25DVm9moZFD+/GCSO07WHe8H+6Xz9LCjbmS7I
syKVsjzgAcwJoG9ZGxYLCU2OKxXJvnE5bBUYv7Yo60n9ZujUUGi5hjv4EbH4wzmfdihFcwqj8eqE
0Vbi3LGPns1guepJP3Bc9qhn0vEH98/J1IwfJACyrHa81Qc/clMrB6I18dKlRTNLJDgTcBHyO0xo
0cK2eHagnmHKnn1t270QQ2v7iJzJBfw87Em/pqSQWm9Tcugud5yasTF6TLxSFwmsjPuK+yQ/KL+e
E4HG65F4O6vR+gpoHHuSOU5A156ca4gLmJDJuGediuvobzFYRDK9E2OXkX1M8dD0o5IysJC6Qtf0
6ks9htDaMNbDftJ2MD7jgeEczmXc1UV/hFGN3hPrDH8/hqDQoAijEtH3KrJYMPpFvJN3cGq8lxHe
fYOsbJthFeHPzDc7QvN+i3Z3bHgN9vEKDS3ntL35+DuIPnQkpmWXs8b529jWl/tauEBCigZrA8WT
zCnb7m1zQr7Gi4GEntZYbhyJfrsopHXckNZu6qoE3/8Wzq4uT3rZeGu552bLGo1TX4c0WVAhW/nH
C/qllQjymgFeYvBE75YDMbMLfk3pDX4ioE2BKMHkLCRDYeXujKkL7eRGvpNSwqPik7m8utE9ws/N
L19PVLCMT7uWFkguwoAY5VlzzM39PHMzviUaiIc7gy1gEAySPYEALbjUq++bTBz2CQpFK8gSL4re
P9ld01AkBfqlxVb1G1ebspDSX/fCbAerV4ReBddWSH0qXFFGBdIPP5yIQDPIbq88pMWERrtdlOvh
VkmT0UtDuT8nee+dTg/d6LpBO4R8R1VFoSA+wjCr0lXzPuMNYdMumjzgBMKOyvj+xUI24JiKDRdn
T3d+sVyp3pLfvrrRwxa1Q+euXtmSte2dHKSev8FjXdsivwa/s/4MwRHDYlYvl1XwsG5AqpnxbzAw
5eEKzzjUhigeZ/KEeEnMhSkO4sHDBRNAhsLhN4ETLnvEJXc7OT6XUI1O3iSN7DNGXANSpdkO/l4B
aeWlvfbQUBxGdhp+8qG5urhIswwSziz7p23Gi6l1QAeybaPeepGHJuephIysibA3q1R8EFC7gmSy
+Bx5y3YAj+xoNL96dviwM25EsXyC56P9b7R9cOoNydcMKsdwE/bOEjKx1IGk3kBTTQsALbyBcF43
XrQFgw319ysD+IYL1MEi80zyK6JDc9PWlvzIXJhI4OgH7wWm2akGI/jEQuINyb1mXFO+E2K/HO/0
0PFCvbnruLHk5M3nXqoGR6bFaSqYDVwtTVaCHVJ4awh7Hftf0L2cPQdaXF3DXIRvsstpbEPN6an/
rNeH7dwnGkwWOjhsx1mLs3fV+hyceSvueNoKjVAKp22pa9NgxyOQiewOrGDfw+rT5pIG2ygIdumF
9YvxTjOMpTJf45jPI4MCGNrilsXvXtXhETy6Zw/ouQKPS9o4+QPD5bzIdRizrgxZCPYBoDDcVRjm
7iIoWLtWxBuskknWtbmx+omRDQyhOa0bv8wt6uMS/rLxH7TXDVYtE6JnuzregDAozamcUiifyT63
IHkMU0RBWPgKgJ7fPLB3GNGmO0yECn0B5mWIxL1qZR0j3+0YwjJ1VQZzJj0wQ7l4sn/XXiLC6ek3
BCtQAzlrOMuTPMRTqBju7Wr4RH8bKzFW/P4gXRqt7zXcyWyIW9luURGr0TH1IcI6CrVMeAOIlfHN
4couQ4QwPdCXfM9smBdRQ06Fkzhj5q0bP7IQ51NIaCs9iVWDSgzGsHqByROgKSaDcb5c/c+VLlzi
cazhEBKBd0gjERdlQirIsL4zYrArCZ4X5VOUxf3LfgO0LksDwY/kwsjDChjnbZk/53VssCW3TAcO
bqnm659+NdTRulmMcJ5wqU2R9GVji0nWy0h/dXMoO2vSDxkawdHP7tidcLW6axboRgMz5F9xbpVs
Iu07eqCA0F9Nq8A0jVg0T/FfhtDqkGld3CUSHrCcfxBBEYhbzneb0oOHkq33J0CRKoIAvBX0cLVs
aFTguX0v0ZAwwO3xTbqmmYYPdqtoXNm5ocF9dlZQMl3vwUudWxBswAvd9qmdLdHT8x4H4OPpeHwY
KhjD2ivdOBqFxVmNnCjBPS3roRuTCnaqYiSTM6zeOk0B5vboIghFqB9OIgmRRZlKbW4KaKmAMbBL
w2dl5JCvCI8dZfRxJRN6NORgvAv3DG+4c5XEazUwFnZkrA6CJ5M8Z+tc2QPssYBaZo0GuOVyrlTI
o3s1d+NKEx5h9GVsk9AFFEZyEx93ORbpsgZTfT4WmXjh32x2/HVPZlSZ4CQHf8JBQTDM+k+rkhIq
95FQZwe0gfexxtgYOCoWXOpRGhG3Xyr/ekotxVKHV5FuIO9fJQQTFVXBm+ThJIxycBn3EB4l62nt
uKj2SBhUR172ltqZZhfzcYuVbhI4aJfyf8amLI8OFgHJ0noHmyPBfou73DgEJj8qVfS1R5GDY935
4RQH/kTVvnwytwVBYCXAl8OAO7NHoUbszV8yGl+s5ZJuYw5WK6A2N4TI/OetZSewp5eltgR5ih06
MM+SvtBLWKYa8j38N/wn2j/lr+9Qq31F7wWjWaP2yRULYEyqchiCCyixNlHx+3li1jLlMHKgXsjg
ZpjqLMAe4B5G6Y6zqem8lN4fQ84iiHPZMMLWyaVmkWxeTvkarkX3W108CEJRGw7Sbt6cUuTtP0oH
9FOY2gipr0fnbMGGOPbWElt2K7obi6PmWlihVXnwXZbBAxzdVhpZ0wzeN8csKI56FMQ/9TMpwxxx
dFdpXLReESlHs1BbioqTAM+a6P4C85L2ZNNHxpLZ7nGZ/1XkmHEuZnfCIIEvTus088xlsvWAsI5n
WsE4rcltfCqI62Soo0JuPTdfUvW/ij8BS1N5ozeNsDy77hLrSoWApVx1YDQ8dF3msX5hXmvlIEZq
LyrBEccsSzVrDjNoNv+vWkM5MnAR0zMW6gdfFMbjXPIWzB/BsIGmaX6IXM+07Y6VBFRxlvCf0Unu
z4okVZCXS2ccDkllR6hMyb1V7NmNk91Z+4rnUIaT/Uu9va1fOEuFzLEfQOL/4g91pXLTHojuQ0L3
Yh1ERqUH8W/sD3MMh8v2OdwSTwLXseUlxQ3ZO/QL37ZJRQ+PCp6a/YJjB155CxAyJsLvARGBnjxr
NWb2PThw7/uFsl4CC3GBgm06rH712jjTSOiWbyQNJYfoCHlFJEnHVIZiSwwjBcnZSwDuqMAMfXGG
UWPIQXadjO7IWneqNOA6aqxPfxAHzxFSsmd05r7YyGN/+hgu12xAZ1THn1nfWP9UQa1LtLgcGlMo
3inaDaUdTd8KbnNsuOIK20lsrSVu0qgf5TKOSkdFdgQCkO3hyeic29R4TrkFJ26bHglgEzHvhbD7
6sLGA5qBhODFyJOIG6FxViaJfxkzVHqdrZdFQf3SMu4ZsFvT+hDkJePERfFB21lkbOmCOA3Fi5ii
vW6XSu5TMVYc+CmbZrvHGQMbSeO928lTyExVIzV4/Rf+mstKX1opgPpntgyKvb1oe3L73jscq5zi
2PE398lc5XiVIGnW5nYpISfc/O0pS/AVwo9/NkbCDwie1Wd1yLjOJGyv8WKLu+lcb3coULyZHEH3
kV9oYvDny1geoKP26xqn6i+Tybv7Cq5fkwGd8U0fBOeJMs58NEINL/b+pHsIxfeD+Z6vC3qAn/t3
sTSM+bJCNRqlyDe3N3lf5zkuMiAIqspmvNAxSmvsZ6yz4ZdO4Q1nIJG7v9avT0Xryx2nWotLvzvt
v2TgmJYYWDVZutO6ry+ayxBayElFjczeGv672JZgEivrgxxh2I2VhBssoTsaiPt6mUOHW7Bx55jS
FlHhpavAbKgReDwR6AeEhU3DBSAjxBeFOTGAwGslac6SmIcc6mvURQmP7ai0cT1f6WJQ3NzvMI/K
nHd2EXLdCccqjc+j6+mvshduWBbwJhuINj+fQiA/RfoXMqO5/xGYMuAOLtCWaSTJNYFsRiV/NV2c
5TcY5Qj/e8gjMLVpfU6J91NUhuERRMialgy0yTvS2fthQN2La39E+XEerK1ZWAX/5vy3ey3y9QSs
LHnmKrGfQgyQvrCTzzpAaC8I7aTa9UOX8rjngsysNrGov5HXYg/cZpdwJfg6uLBFKrAhq1DCDoes
qL3ZI0TJhYQmRm9v4gBgUHAUYVC8uNc7j5Uf92EubZq78P6AzKa90bhj3goKNZVQOsZOl7mXa97d
aNj6c9R3KEzLX99/A+pibx5/B2hvDWXhkyph6LrnvOZWDrYbyu2U63hUYYwUFYEwTd3x6EXCNDmx
Rop4J6RXrT1V/DDjBbSJMTPm12vvgcvnYSWbV5eH30V+8vphQRuE7qUr2zD8moUBTttYJqw07L8b
qA75wikZHJDa5fw5UK1GAkqyYt1oP1CG48BrcqpE56bdxWIK32ii3k8zUM9l+cHRZm3YGDbV7spH
AX0Ub77PQhCN0yDVYGH9kjv4EAYHc0S6ObH7c0Co2jvbksszk38Qyd3E96ryqsuUyMDHcsRsj7Wd
byuB7xk7UDzTxtHuozO+TAsZxUMjhMzcQLQY2Q+JyOdHKcLWpsmqM5lpKyWrm+0ZrvKVHgbEOvhZ
EF10CzvxTdeSOSjtcKIIcnARCAW26ET8/ZHec9icB7+mfZGNmhOJbF1/E2qcxJbZgL/c/ZLCHUpz
xs8aqipJ24gFgL/G6pDctbjByAb0fnpQ+IpYQueEUuVrzzxe++R637Yz7bvqefn8oT0R3dBdv4D5
vFUZHZv5VEN9txfgM6O3+/Hvy14oB/zUklgZ9i5UxQKPy5Cw3lfNLp0lfnJLhAkqMkAUdtwELEQ6
CZ2nGRleycVJnK8v+FYM2yjmVS6R7qJu7jtAv74qEMvJZ4/DSwWKYVH2RYGoxwtHZoz8jDIhKYFq
CFtJqDu97oo6fHBFjwBu4+bH5IYAWDBiPtBrRD9APpKH59HoLChv+jEYiuAKjjM/rINB5ItSHTkt
YxYh68nsjsPvms0GsiMTRFh9n/06Qteu8OQD9/oQmcuCEZa24IJob4CGp41LSqZVGLEKG/3gT2sa
a9X38G1I0LsOSUPnqH8qv4/ay3BYDsTRNjh5pUK52lTx7v8FMT/rTxUCpdFH6cjjzCGstFBXzIoo
EQ4SKwayTpYwy5DbnKSldYDVRWz+jlPaVKeAEL8DX8cvxlDC7R92RQtgYvzUa7GhwSV2EnQXFoCY
JP/TLHhBTEPAvS6WCX1TuFZ0/eihEuRYSJQ3PpGHEG3ZSNoc7igs7S1W96fFqgJGB0kTuDomEENm
+eMqGsbp9sn0UF/Ii8A7kg8J3FDY0MPd3ckjQn2iJJ+SOKdfYZPCpP0lG2C8b+JWixWXzZWNZIVI
gPE8e66C0cIvy2Zg8DzoMMtZzExZj9l2Vkr5KdRvkcl2rPzWaGsLrbWCXmTVR2fjG9CnDHIHQKnE
/HpKaAzHsSsDpzM/0udvQMiFoBdxMpnYp6gTWdVUWzE3jOoDOQ2MajLml2fZ2rZzC5vSwSiw+K44
pZrdmOAht9zcs6+EAB8hfeZPfM97p3zJRP5TbPprtt72Mnx4FkETUmlk5UZbo/tZWzN1+N2AkmSF
CneUP1YjmFgzj76GeixupeQcUi5W8a0i2KOrACydhsu4cMtFi0ZBHKpCGmhJ7TJ4gUAStOesOm9M
GwTmq9CezrsKViNuhEFYryOpsrvNvBwQ8vyg4x2ZI/Gg2DwL8EpJGjBBO6zJPkuTxaFwdoOODGeY
d7vBZVaz1VqftMyeEoPqz+mb/arDiIRhbFZA7mycgWCoPBIwkFeKtzHvgyrRMBePFzbVwl8hsVH/
gRYB1EFj5MFNM3OKurBY2qhg6aGHjj0TSq8IqidL7VvasDaY/oLeDAliBCiwy2e83GyXWy4vT3Kc
i2AmPqw/zqYj9fLXERlooJFEOimwJqnpxfDC8KPd0/X59TNnQ2i7ZEzgt9Uj6LZXGcWsXIhL6Y6L
OvC6t4+4du50VlGQtL+fSaTsFt0nKg31jnjufJQ9E8hoAD9iwT4WhGCUdP4U6FD62ZqByJmTdLlD
1CCQMXxg+6+/KhRMXolupoYxhUqWWh5HKUdXt9VdTAOlEmoONIaGb37vRBpY6vcVr7ysna1hIpBo
5WBDkGTzUq8g92TxjBIeI7stjB8awUi4hCZsfWKAbSc65Vk6JryTLDL2WKVkP/87JKT4iPqA0pOF
BR4MyCKiS1mJ9FH7Miii+7jk1jQOZbrSI5rhsqEahdfIzGQ3Ph/EL2fLznTtm3+R0LDdX35nIGs6
qEReL3vDgzxA2m7oAPVdZdmf2DZdofRP1h500FaivyM148WfIlOIk9zQk/1wkiQ7Vj9pOqtEfhbz
RbNg39gncHZM3FI4z+CyYIBIUHUDkzz4f1fsTRHBZhvqCZt4r3VOUe+P+WDrXBKZDGi8w94q5Jbx
lohIi2yVCmBohgwosJ0NXRSTQ8RentuOzca7dvlnMLil/PUJpEdk/7SEBwx4IyEt5bxxq+kVNRAe
utH8a08+SlM5D/gDFWoDC9pZy8X1VAu85uBPt+yC/oAzAmWwIwHQ2DxI1oyejoy0WxkGcN4BjFiU
KYN37hkvlgGxb4ClxT+CsdKS0P3I4SrE39duWBJALYYmkEgbkBvseURQTffbcWzr5PM2+H0Y4R5n
673gVJZ/SvXjA85YAAwgd0/TIP+rhY6V2rw9aVwqhkXr2O2SHcoykzUCx6nComXiTKUGMAtTxKIC
gys7+guqhGTmOwsOB35v4P7y2RJJua7axvQgiIlhlEmvpLjAzh5WI0SMN5hDizSE9ckecTeq9nro
amJrQwGKUbi/NiDzpYSr2yawEEZj8bxLvOWQcWKJs0iV5gWkxUP30qweGtVjtzJlNotP95NdxbVO
QM6OeINO/yRbdOcO3xhgLW8hh+TVBOb0W+4C8reBpMZ9tFWbpT9mr03aHckwyduhTf9UD+cCPFnu
xfwNMnebnA3AK+hEsiQD82dhjCUzNFiZeuHTaM9HzsyMjSCtIDxIdxbp9MeSfVRwOOH1qmfoGKyb
QnrfzGAE8qiPOmIN7s8GlEmrSvwu6ZVDeSL4NxeY10iZJm/x1kgkLm838BMlirXnoQfdA2Nzk3aZ
6RIFPgbu2aSthsR/egB2A4kBGz4fn862z1SlmVefztvRlmIqWalMjROf9tdYroAS6ox01eW0nSog
IRkasdRqzLBc2tSzlTwrQvwugNYKwWUu1N9OId/cN9DZZAdivbAy6dTpjHXSi5vT75vKG3WmkwEQ
VR/Sy1z4uemJwwpnvKDcKiqr7xQ7hDGzjjFjv+pvTGBNM6ixKiflmoqvDm7uJiCQrnlXdT/+7wgw
T55M7+y8TxWQFTB9DetNIDXMIwoXPFM4JjruQENaf1jeixA/R/b9nfoo8LsOM+7+KNKv/P1kra7D
xTpBkYjOYkBosLqzggXzhgqsZQoBzamtk+oV1A1ZvXFwayqjUZYPuRE9guoLTd8KWrLhns/vQjfo
P7Gm3t0jBH28vCwzfASm9nfjqeKQ08P9zi7RseYbz9X87aDRPBBkSAOvxxgGV6aHuLoW/QbEqPAs
kB+cePePky5UEQWlEvym8GCbzAiXt2epra0oIW3h2ISrwXhtTMgBl/vfgy0cqPeWsBfXybUbdXO7
tzo1AsL9+Jkfr4Luqz/0iyXejYEo+TecSSFIU0o7aJnoV30XjaT0jFz7lYjoD7UUlR/TFKCTnbKn
GsN+re6GryPypu/Wjv8UFCTFfGrE4l3tOUBHn3uXDzsFEg0xD1fllV3mbbAsgtObsipbb2UmpA5f
D1NbIgV+qZ4jTdoWuCuYppTD7yffLdwQxHjf0MAYolIwVIxmYc0T/U/VP6pY9hlwFOUNE8YM/pRj
Lrw3LZqcTpzngoAmK+9Oadb/AjB6xk2gFMNVcvmpwHiAml7T9J7sgwoNqMTvaqLkyw803RBdTEdo
rtNmaBOTHN4Io1CRTYnQSQKAYOqMqldUJGJlfUCdQydHsEbCIgenvGpbq72ubPhdlA9CB3csus1F
6iT07tVkKE1Rw4+oX3sU36kPIvrNUSBVfpOmJfXTVtRpPYSXdauGFlm4TJ/ZN9tTb0fIJhPAzp8W
ZqJutk0UFUbLM2WEVE9ZIyMlQ+IvHVez1nJ9XFrtoXKX/uXHy3m9Zs1zLoZStS+hZlHeUW0xX1n3
c2fws8VADBRGv/7iKUvhdNgvBGXLYxinYSXsf7pCxSqYjF+zB2mTCZiG6mFBRHCxbA5bPYxFJ55I
Rg5gRZeisnIqCQqvRdhwoWKuqrMgTPrlTvOrCtYNyAdt5D561lrESk7xd/5WQYIHWSFCgXcfknUT
15a4QymDyG2c0AA4odJ0FQ/Z13M9tZRbys7ePfgpgwq5GEF23EkiEKvYV8vREHkhMkXkq/Q7v1nh
RH87k5b4jV2FkIcO0DGvrma1bX5EO9Cq/QpyOmb3/EHyGSblmhK6hFNU0L/0MJRlbVZzpG9rVZhq
TAGAYq521H5SEiY1/miGK+Um+TH9eMPJGMAygEMD6vPCjUTbbpoEvo35+84tWoPju/So8o730FZP
jryjMGCBLQRg16qNm7EHELshNO2S3f19qb2UCdpWuWgGcsuj4CN31RTml5nM6cdWUKIpmC0Qo0Fp
wUIewxagFfUnU3dpt3Zq/VXUYNQ0biAuexQCF+F9R+qC2Bo6JzbPoouxDHBZFHui6wa6SrZlM+YK
TEikwmByQIIRRKRo0D3swiJSXYSm6ZrKCpfJCQ74ccWdo5/4GcUyFeYE8WC3sEd6DqAIu5DYz6et
8tFqH42Vvjo1zBHVX31pa343EOjg0q6sfpVfqQ/DSAcpbJkLVIdoEhLXcdf+hrsV2Ew5yIwFME9F
57b+INvVL1G7vxXGy9TaR6r8lGE1vznVPsFA01eHeYxmtMs6XXcAItwC9S2fB2Vq/2cjCw3pTkub
kCPsGRjFs2goYTxJThfpbYCH/6homyeN8VXN5ocmfllOqxP1g0nH8ziHF9EH9cd/c+vs+Prie2IE
smoEt23DpQ7JkZAri5Vqr/g8WmyRJoK0t8g6pQRyGLe5ntcQ2C+J5CCyIuLex6HFb9hBVaX899td
Yv2rDoOaSgIaEruO1HaUVPTkQxRa/z1nV60lQPQzbBgG209QJtLHRhBcQXSYHDcReoeiBolDJqvg
JZXKvwhZ0GvsdFJ7bsimP2fyXd0fP4VxlRT582Pwm36wx8zDhlEaJmPCzhX47cnoXWDfjYeSmgha
io2Wf2qmU4VFEeFh1fCMZkkMZxw30vKBrVyDAW+c6Xt4Eal3uZVqUgLfdHlNSjRtoGnXA2pXY8OP
qC0irFaSCA6imqv/A5Xj3cbrxARgE8Bm+uAiZEKTsrhpXUpDnZk7sHQQX9Bng3D6SkmibNmlHwKB
GsK8A7nbRXdFY8upYMusKsF/FUzH4hzhBXneSSgBQlmPBbORcroqy972jv8sgQC1ZtiMzFvuOvqR
xZjBJgDMMYJ2TGOhpMszH0N1EXa4mGeEZRXSPJ/8qwYIrQfhq70YRNtSYmKshk9Ptgxir0Ah7kUS
b0qI6E3KN5bXrHRRPH+pLjfUbe7hCoAUMLEXTOkrrE2Sj4apjoKW2lj1y6yrEr/a5tVhD7lGVPqQ
ZtZrVL1qO48v7mg08jDaNwS8LhFwM5n0gDv+tBcwmLLZ5yHvCfN9CyXPpRSeAGd2g+TlNMDt0Dsx
CRfhbBqkznHl338yMUm99/tEbPZMch9OpYjcXjnScpfXL7LdUWchth0jiq64VxLsYC9ZnDF4nrb5
ZZUe95dnr5IR32d3J+3JkyuW449C85vO7CaODhXSiR1sLlYgOavKROh2T6QCNWyNy7a8q2IFNFqV
MHyHM3G7BrLzOuJUZ6zydxVCK/oLcz3HxYFrFDNtC/UYi8XXWpdFzZqSayvOliIg8N+vgjNvYc2p
blyyz1LK+F4OtuEwwkReBhuCaxmvxjE9807qZGs9OcHjbVrVTevrkqMAkJKr6YmlQjIE3oV3hAWU
1wa3LLo0XNIkYGU3rJ2KGo0qeKFWvj8HjNGBWNCdoxHZfrA6QCRjl0IJbMPC+2d+7iDym7975NKa
IX6MJjF57rdD25d6B2gVtFk5liy9pivo9STc6VKlGkyJNkjR+5CdeuYbZK/Yxsn6nycvpr72A/tR
o8zZejESVXngOgF5ZaVYtv10CUMOdKeEMlSRuqOL+b5iVeVhoM2sU7F12YZDAt1Vw2hxFbb07Wi4
9AeBlTaC4YYS0713oyjD00xBXWY3FftVHais0cVAz4MSKo7lSUi7XUPytBnm9MOOORySd+wk57E+
LZS2dnMEibA4g54hS2AlyV8hE9SppOkteYaFtOJhz06LGYbLp4o6a6x8j6YG5Zu023IRP3E7l6NO
veOGOXFWIJ+8iRFtn4YyysJb1QN0JCeYJcfkNGsD/PbXMZ5PzGE5Kb+xz1ELnRpiFsaEsvQKe3Ty
RWGxH6JH+lOAhyafcnknue9C+8FvfeGHMtJP8xP+E4HWhxYQfoV4BS5FKMIu9jXRyi6msHR3wR8i
FuQfcx2oh6kcGp/j7C2CVE/mir6VdHp0p613FqgtRLmqZ8MWFi6wK8yQCG9COtUzzERxmyDFKWi3
Fv2m2NtuFSEJDclQLI/MnzydKepdkRdpLZ3U/3pnzv0B5YESpA//HSZJ70h1Fpu9GogIr0Qra6Yy
bLFfY1q66+gTV3hqz+V7KoeAyQ/2jqQqmsCmsDpErt5BKQRX3nQrHgE0Ug6sKjz6cKqqzuFbEYjX
kvBeSx42rY3TUONQZMqVW5LUi3mojjZKBJXOGuAd6/W7Bggqk/sFRCVp1rkgmetpLrVZd7ybgM4z
IANnXtoIOfl3YF+tmy+Du3nkn4P8LmEtqOvp5X9lU8CWrTuDZNE69RZpXCzIDNbC/WS/9JJNpktt
rFZ3Ay08mAyx4tCLnb2Aehh+LcOgjBKg8r/WSo/yAwfKAmOsWOgWfNy+21w0IVCWxLCv4UI+wWAz
IuMajNXgxhPYVdiqZIuObsc8EVRoPSEwRmlE2KRYLHMJJwtQBR4hR9Rv0egU4HQ4/5pnZf8ChsMo
TsbgJdi4MojjOOFpfxRYPJVQkKiyYFy4vlACSHHRIzDMOpFwzct/ISqZxJOfb0rLEigz88QR7Bb6
HKSxqSdLUR0i8430NNY7xL+bF0Qk53T6wgZ97bbMZRkj+3hX5G7Eiq+JjntEMbjjwg5jNzf+LzrK
jfYpj2PJptw+YSbJKOEgqinRjYa6/NK3W8jh9Grsyv2wTUFtCYJ6E9rcrJNvIEWOln0EKtEqJYuR
ii5QVYBTr6A9C6d5OundxebNCGUMPdw3VqIN5cgHhiY+fsf+3RteTQG7Qt0RML4tVSY1Iu8vkKDt
/4BCzhOnYLQ1w6NblfxV9wDv/U31zdt7uizWRcTMIMPZXr5XTjHK1DC33+PFF70pT4pCwuo9K1MG
w64hEPsw2mX5xBAlAPdhkhHocpibsLEliqhk69prnAef+qQzihvQA0Wd85MMTfVK7c9nsXccU15B
2C0cEDfMoqmjEZY95QUzph8rYO5YIDlw2Ejp/oAH1R7jj9scWTaAB9Dn6Uop5y5gipEm5pllPFNn
95Aw+jCa9++7rimv5YqPlNI3+ZRjT36Afs9RxGDPNpdI4ROMhUyoOl83XlPVLpSv420eCBD2fwZT
nhs0v4iDTXLvDgiNTOiyK8XC+Ng5YxqNy4ds1GTjdlLAhBxsJ4kkLC1ezNaZpC2zrhb5YNuGOudx
I0LgTENz8EDF/dB+co+VuWBz0qJ68nLzdq8cgvycRLVW9pZqNUmGxL1puCUCNB3iS1TEX9gI8h4t
V7mKWRNoQW52KWQ2hJy7rJ6AmlR8/aU8GttNqKFs5qNjmhC/8l4ufbtXXLr0Z1OcxgZIIWEP+/G1
1MROqjaSPOZfzhRfaHXJ/r1pMsNaKcyayw+H7edRK8IcUHxqagkV11hNmL0h8H79vO0MQhFERnol
aNrsU6QnGnAwPPvd5Yn+frqvG6IFGGqSVFFdCVzKGquvvaLJck9TW6ZfEc2FZMDvbu0KEeY3TUpN
ofqPyEz3uaPvhlE19m8bR37j5SkTRz+3h/eWhwGVw8oTGwCvUArfKoIyNzDpyeqkAiZZK0oV1UrA
2+/05CTMmBb2NlShqvtHMZdmSlKTE0iSqMe17dUhFId52pBU8/Fr9hu+xLZ9Cn6B5pSAQOlKRp56
6G4JTnNQSiC4CRC20+5vXRJeHN87XHohWazQpxK7UuNOgWUoTkY34fLTju8WfBkbjT1z81R1eO22
jFTlz9G7/MgwStOWaqqfQYgR8NKTUDiKnVuxJ5dbs81MCymGwIQwdfTtYu5wqysGKVq19qn6pghS
zlIhXoE0EbzP7VgiBbXyFZR2jdnLUzi5AiwyFNIqW9udIiB7ds6U6fLSisYM+gTukLGtgxd66rGk
p1m9k90TyFyKgIFHkLDM/dCUPysETRiL5R2u48Xc5JYKJfhBCM//ceU/LQSF+YaXx3zFWOvkkNxq
B0nmQvMqlf2qcEz8cp2LCXaHHKTrh7Kk2o4F9tJIZUGkLWNQfqn9zRtbqKiSPw6gYopTctPI8IX7
qDkjv7gxLq/xlcql/RUMTlk6Sb/v8P3xXZxAYtEtHGNh1nYm5vrcPElcR73K54qhmDITZvRlyJ5w
KcUyPLzisExBF8beqGiDondTlHAtorsxOInB3d65Jb5ozoeEuFYb3J73WITFNhWqJq9bB4ofSLW1
WTaZHntEVdBfbc2nOIfvGvRf+fFgZPqRa5CsZmm2MJECP0ZI/Wfzh82AdDxDTVi48Q/R5fSffG1G
ehSs2Pei1RxaFo3H2yFRL5Cp3EnWb1uA0VsJmLiESJfXi2gtVQbY8Up8BpZgGEkxsfw3hT7s0DAA
l3g9lVu4RxbuKRj5Hmm7OqDz2z9Tk8W4+erF4WSy4N4PjWPDnoh8uQ45BQyIh03IkH5CuAeE7rPI
ZhNJyP+H2WLj+SW7mk6Xq3HBU2hoQ7pqoIO2Vv5bYkXs0Odijq6fD8bPxAobcRkKg3uoyAll0hxv
G+q/PZS9pzN07fu9pujteAq9Eegzo9gKmbDscXh8pcv2tBDpdYnLKphDfhsejeXhWhkvm15EsDoX
n1bBYm2Kr66XodnbyozuawptOD47uiqb8oHq7xSjkSMhzZwbEbrOhWS3sHVqqQq8L0D+dl65TtVg
E73zckKlW5+JKFC1kQO11PWAyT74tsdklI4zVvlssYOs4J9aZZboHR5/KejvT95wvkDuqeqrxw61
6KQZH5VYlKhU53WY9OvbVNp9O1Fxyp1JF0ut51UkOS+QdW+UxIa9E43ggr/m4uenK3/Ho4tmkv7j
kSkGfIGbnbKd6+/MnjRgZz59as7ThftzBOmOi0c0ekKpWu2iqEy3iLez1P+01zVXni90FznWeu2p
6K9UgnupkYMaTi9bAvAQ58Z4d/wU2xfPzBzo2Ov4ZUeIbLNn9ek8YvQgiafC6XhAJGYrPDPT0Gu6
UWYsKcAypGyC2PV06lO1/M8y7IPKbqJUoOLrbjx1A845//g3ZUWgkOpjFxjyMwHuOt5XGl0vH0RZ
H8jWBDwj/yQaTlkwZ9DV4YUfiqKazmNCOU1xZEFm+/Fp0nWejRjP+4SGlN5iv1TnfXdrCyhxnxfb
qtAgTU8lCyPuNmHjmGVvJVtVAeP9+FTC5Mu7VRiVxSfIEopdoz9KklEKmRKjA/EeJWz4/U+ZCPVk
/TsdzNKXaBGd+PtkqbCi1YbcuGXmXkZg7EQZTFzZAJiQAKhQNVn9FsFr9siOQY5xSIOgXR6C1X0V
GuSrIysUEGlRj9hQJ8MYHPy6vO17BcF+nLIxTDet/SH5fcr9qB95jmg0+rP8ympRHGIknoGS58Jp
n+kgjZrdhGMD82c64mCaZRMIAgEqg1JQlbMKt47DQFWYq4iLF8iwIw97ZOFazNfJebMcHnmPDJj+
GZiwbD5r/KND2SuY9nZC3iIXvyrVNTuUDGlOTTJgC4fmBZlqXATopoxZR8hYWnHGvA6pPwe86Ou5
sg2yJOhmXDSyqX2zQfrfHVMjsbjGYmUjbznjasdkw0cbwH6vRYl8cifKmmGJ8qaJlINWCqlsxBLj
t0jdms41PRn3vEm+SYxk344KQvBCu8JsrtqJDyz5+wjD9Aa9TARvipqIV8D5/XX90LwtTUVK4t3e
etONWbgN7jLq+aenHvOsKqFjV8PrA9InUx8mwyepABgU9XPVs4Q2iBP5Lj4AB9g7+ffWmE0Gd1R/
2psQVItVM6yXDCBFKYDx4OvGrKHd0mC0GOgXmBnWoO9E9wXCYrLzKbuZk7d8pSO7U5Hz/s8h/16M
1vaKS6rA8MLePJmhtHO05ndDC9PHOh4luLconqAlgDlAnL8UxpG9KCN/NTDMfrfXZm75LByTXCZh
asac41Nx3jiGgHfiGT7bv/jN0yDf3WHYyg2KxB+o1ivqRUOxCn9jQd4ZztgDI+fH/MbuKaBdSrxk
o3tCzCealfhZE/gbq8cEIt7J60+MGxNS+64HKIHiEl8uc/kzAvFIQTJ4ktdD1s6t+hqntkfQkWCr
YpFGsvTba2SDqkOaGcpbeVLHEKiGbf93XjrU5m6Y57IArpsiwQbED4msCZOWmNQiKnA0WJrMX2ow
Pdwx1r+e9y/ALMwd0yhspbzK6EEktemJ/mvEhyo9iRlUabbV6tXBF314jfdtET36fB6PBxfv5HdO
KafSTR4lqieVskmwsQENfnEeyRjPqcWgoAC+I7El05r7hx34aDZwB3GU7zu2sPWicfMYjAhqD7Zr
Ha2fdMAEXo4zUO0sl9NVJacSRW6b6tCE1wgDKddwLTXa34ePl8iKdqGD3p+RGTNCAs2mMCKmQq+m
Xop0gbu91LdkIASs/CIG8IqwyPcT0UYSFK1WtX/ipJYTX0tUyToBCAlkrnO1BpF59VEC5rQZd506
BzCf2sRmyjckHkc/hzKmw4MXVo5IT0Awi4BYeS2BzxwHGJu/UlIATIIeQalGVMDF9Y2zlnWaPD1y
DQ+cmiIleIa8j31drfzWtGYT5bQvVc1ApCWF4qCNNrPKreO978NTBSQdECMQ6MhdcX+eQpa+iIr5
/Wi8a18OxYkSwY9uowN3SueXayd7wbZPJuUrscFz4P69Df3PuloBVc/W4w1hHACaa5jsg/kfnqZs
zCDbRx4NLH1Cv8Cc9ZhU5rqbWXiIAIguX8szn0XU5pOtiAABOZe4H6DVedUbponkcsntARk5cEm7
rrRU0lsojAPmda8hUek0BseUudA8iiLHI3HomGBmPUJZr3EXSzi3931a0RVDbLh7AuJSl5S7e1Pp
/wlPXealwTi5XWLY3aPwQU1UPT21hlfl85l27F+Zv7mcINi7Rqv2x0QDoblhzBuy7g6MwE/TKL/V
c9SHc/9yDGjCYPgk86Wl82d18IdagTIkZXSsFNM0nqn12mRy6vHriJ74KI1p9brP2fyLy1tp+Ps0
HWsJwwCoDCk6UqVYkjtCzlnIs484xlIcKVvnnJO6/g5Mor3Ms+w9AZssghEosRBAwB9FOy00bwJp
8twxzPAwTLg+wsgPgzHIv8onlVsdON+iwYBYxPx0Q6ORtB2CLc36GP8IfLXGra9Y7vsRtQLx9p4e
g1rMLyhPUeufz5Xw5nkh++6V8WcJvE0ksf+QTD5y5nnqT0zpQuAQKvxbcsZxN1qnfroECejeFj+w
b4buRT5EOVPY1ZlUwTTvx2Vq22qHbKDA8PT2uuopKiy879LMbW5o9tClWXCTLzCcTgy7sc6sACrF
ZF2tbQWBjiCSOk97oMtXgrBL1Pf2yDce17x07hg6Eu0MLV3C4VDnrbm8bibIwxFjbu9DxAryJ5Mh
7QjSgILoud1wmTplikjHAvJep6tXHJDZomurPattNi/fckSYElqnvcLpjskPx3mn6ksYEFzrLqNZ
0pG9dy9krmld97tFD4GFY56cLqSqO45KI8k0Pk291rACretjpEKtpAHTuYDpvn29GhwM1G5sVkY1
900LHKzxfiTYpNdUUl0mxpOxpUh2YP8m02wNsE3+OsQPRYAO0XBbiaJGXC/VDY7HIC42Py9NcvBr
YbJTiGp3OfQPWog+up/nBeSD6j9mDygbol1ZmwHqkFTjvmYI6ZEmseUuHtojR7YCiBxImORfOGtR
GdWZM2+tQKe83tDP/PiE/6wolMsW1OIO9q/2DSOvcZwsrFZZNAfDBbqoByTbekB1LyS5BgYPcF4+
2S7z6/S+m9G4O0yQGZAE6cQWrn+Gyjb6eVNWXPJmiR8uTl/HBBNxBiTU5OmCxqgO1KBlOLRIke1m
ve4gYHxBlLJ92J6a/4mc8IR4WXBwRw6L2GW0C11AC8hf0DUg0bPsCgb+aa+0kw7wQz78pso8yS44
X1pF/+535JHFFk5cL6oWnHYwSa9fjKmvK3kCl3gd++Ti/qVXycPKmgM8YGWgEFJQ2ezGsJt6LFDj
nki4LJqBfWkA9OJYGxrpqcIr77OSqmdr19mH6wd39gtaS+po8Mre1qiKH2x74o6LTUJsiyHjzJvM
Z0gw1jAB/u892UmK39+eA0V17qu6qh2a5Y3ODPWgdQvCi4QbuLSKy0i54L4uI/3XqG49oVwPI3sg
fxFxS07jV3sBwDN8gUUgVkSv8b0pNo8EsTE7pJR2kbCxHJgAtga9laEgzE711W5s8RF6FEN/5hbI
rRygc6A3O/ZaWD4bCJt5Fbm6ddc4CuAmzJ8HKBqcVS49HAhoLuIqtURZCQEJQVEEWM4mBSqm6h5U
ShjP11QEu9gfB69cGozR9NAi3hPF90dBr14OQLDMk1Loy0VwC31gGgcMye0hgKznX3SzUghfwHwn
VMriRLjvvXDVfu6XpSbLBbNP4bfjjijCozwViqG2LdavTEeOin0OORJlUYdphDrwEFFa0dWQbm3z
UMgcXuxzcpF7RQ1XjURgWoQMBcW53AOcepB2wn0RX0suvAbr2ziTd4nKcSGEC8YIQV/iMqklG/wP
Sj+Gk8y0ovTYyQqCr1aMGsXdJaXTz/ZJYVXFWSbsFhoGG8o3UsQhnmxUlKNpJcJ9mxis+dPWFRVL
VKt41xyuVOkMbD1LJsZpcQscZ2Xw2grn6867/zDRZJyM6skS7HIw+YlsbZO8zUvTC2g36ouPZBkQ
JqW7EFm8UcoJlSW30HwW/eFgGeriDjLSWXtjPo08ourBDSMG0afmpEP1H/I65NOmAY6l5goZiIxx
Klx6iG3tBAxhsl/YPiYSFoItMVGV3O953RPYnEOKTHNDBj+tH3b+R7Zpp3AkPUdq3oWR+8yAXqSm
wwFb05/u9JB1BeBCYrwBCRc8sahkgwJXo2S8mrz1B8lCNqrNoFwtYGsPZbUmN3fPA5hICtdboRDB
XpESHLCi+aGFGiim4VBkhueYbIcRrRUj8YTmo3Fj+AiSjE86nQ+wH8Jf6iss42yqQXDX8Whs3FmK
ceUG5ddjXC/k5Vv3WilAM0nZmhLk9AqTKsgq5TdlVKkA9SrPQsbkhqxjsbhPP10FD6oTZluAzaPU
H8gb8/9I6i7cZykUDYb1BIJA5blHMK20+MLUEJyLzwf8NRkMl4nLcZqvqWmZ6i1XrwjXVJ9kBj+J
LzN8gEpMawx7pHnr+cyjBD2/bhQo4BDDXc4nbIfA0FRb1h/O6FQ46ilOA84iCX7jZdmVfQml6OzE
VSHcediJjuOc7d8ptaw5ceKVMrIsjQazzQ8nKvaOZ0BZEb0xOUEqgGh5bfwI5gINdxKRJrnbwFwX
SCoQRggZJH5We8VAdszB5JvwwhTS3RrLjifPGcG6KZcHc0J/HhvnfVZyZXFm8/xboctV8aO+bWoT
L2O3qXQNz1lJyLbvY18bidAdOZPAUGlDnAJOhDn5jalwX59WtbQzeYidqbnevLmpQHhM8TGB+tmV
AFuAuaVdTNqIHcw3rB4CaXcZskLeP4aLpaMwXAODF2IVuiphRjI/4fhSS6MrjyzmKBA4XHUK6Rka
LN0XVctV+fQoiLtXTALiG5kO815hibdX39+0LziRBfGf7ZMIRd9cMu/hwKdultx4fs1vpj+NmKPJ
zU+3UlndRfxPynSJ2C5HojK97PydMaD3d3NCYu2qfmfG/0580Ufm8DxfZoTQDz+40i74Y4tMHr2C
Zhf4WqOCEQwQuerpGs+/xvupHafadSc1TX9EP7XuoFrTkuwGoY7YhCs6hCJlxD3cLxopLF7l7zcR
ZOnd2RJfnKuuQptoO7q80nPYNWCNH94ZjCKFRBNw5Plo0FNNumb1utJnVGD45VJI4dkuHZmjoDsE
dtOCizEvYDU/5Y3tSKOG03MJ5JlrNDzM4tlG3gQfU4sIhXR9YvPXuN2mW3jY0HsHOQy8mCRHXYVa
rC9XxDd8LacHJnThUFefszWcF9slLTx6zBVgXA7fpq/tq9/B+g6LWHHUWocU4HuIwuLGW9990sIy
vb06sTMjPM3juZbP+lhzDf1WiNqBLZYgEmZR3qE6hFLW/BNUV484c813dLeIOMKJs+toH+WChqJa
8GHtUSiHSgYGY7vdn+V8ah4fDTl3mzedArm8FR+OvDiOatVCSmqz8jG5RWHk+IyR6ZGsyuQ0ZWwT
iwaO9mtoqk/1DAuerInTHP4qHOM195ujM6aCkJt43/M4Io3SsCWoI871dxRzXcc8lRoKJlBP5pZX
Y9EW/E8aIM6O816wawK5KsE0ETmTQeptQ4m1eTLagjizMhYkRFzI9LkAsQrfyd2OKYQQDMV7UAYF
ypMK5q/EEbWMsjezglOY62FC/v7mIFmpsPaP0pLwFG1eYvZtqK9Qs5F8RXlxBdb1BD3aI7ixY8th
DJVksbXERJgUWZcIdscGip8twr1mkWFMQlvdXlUkRFnXX0EviyV263BlF7HGCw/MKjdJA5t4iZuM
LWSU0yPjwKF9KhdCoq322F97EdC2Isoefr1poE+cHiTsD4bLzs4tNIQKdHviymW6UtpZ71yBtMDY
4B9k17c+JJezIuyH55/q8ZpmxBauzzlFOpNm9zOHM+M6xUTBXDfnwpIFcRt2OI5S6ShBWhjDPs3q
PFEU6VSzQdmOVuzrLaUTaoWqAB3y5x0JT7UGUY8oUYXW+Tve/kO6OhbvfxtA/8YtOkZwNqzvN/Og
fckQR9NA5lLJW8SCAVodH4uSQZchAVpGvILaSyn5rj+j5+DKzgp+HjW3VP98c5yBJzT3cQFoAxIy
WRpIK5l+aDBgRy4jz4TAS6+PBJsFZhF45fSkODABGHOKRtT5NwptfxjS6CCr6/nQ5A9hAhq/ERoz
Abzx4CaXqeo9jkS9rpGl7qS4FcbcJuipKvLKm4f9LPBhu1gFyz97Z4S2jG6Gxs1yYXwcR54kQZxo
kZHT98nqmBFuYbj070QGC0cI81MMLBQQcNB8BkyEYHUnpQEfJLZp06OCMw4Vf9rw00ckvFTBLqLy
HwnNINo4hztYKVqduDNgSa/6IEoQMqhaZoJ0fNltWkV4BEF0tn5PmS0T8fmszlRbbQkauXAbZOWa
Ut/gYDiWU5hptpw+RjiBnmgXrbe3t2nONArq6jFBMh/8jlT+lyR64iCwfrMZX+vQKW70sfJER32M
WF2Yj3791WFN9ojKLLTxwnCRSUp1vpd6KYRI0SVC0L8ZttevSeWHRs+FHO3/ZHS12UUnULCTUdsN
ah0sWfj0tSz6Nsvkyw1CvH4Zmz2MaKAqmru0eH9rycX89M4D9Jk2Y43CB33UcgZGY47EtLkRijuu
dS6RTFlh/02ESMTetgGph+/sdJvpM6ZaYr7VQq9nZS8o2bp36BZLhvsyauT74lwY1Z6+5SC6BULw
Buezx9bbHj37V+ZPQ8MbURRO8gYTQKHHzxpPtRWmhTv4UAXIdOjIqOAs/xyxgFxUrwsDmS8Egsmy
PMEhLgLwWVIDuEJ/gOMfCQHPAvy589M8DQ50HJ+4KIYYv5RaY9UN83/NYzZ96j0PEbs9oSl8ZZqo
9KwhtZ7kLcc+EN7YiFa4+npjbPPtmfOtiEHyQzLkeFZtNAdj8O8Zsw6fG0NZrPM0tzSTC8qNtuBY
TSPFH6wybahHCxebS3d3T9hXLcvdxt8emhK6GAfU1LwL9utVnNzIjQrAlDLJIYngoH3Q1IZSRTqm
qcBd5Um/yhPnIwtKBrqKXhXs2Q23fbvV6SZmiHiCeKO1h6b/4FTjUdEOSz5UrSdLcvrnqV+mIWcn
nxZdcIG0ShC4JYExzmd6F7/ddm/+SkNZOxLWIc1UW+/lEK4GMTxYHXc8KN00cBK8iGmMxzRo7Mg4
/etwWJ1ODoeEr4p0WMSfkL9Ep24s5rIg0nsSNkO6jCZ+AIqYQmAaFhFDUrb6eQTJB/1gSv1myBMt
pdgtkweKdBTTXiGlhaxA/TvAJ8mS9RgbxfLvfpLFBIo9J0dPzB2uWBKK9nsjzEoNjXiSBb3QL0sE
wc/aUpnB8fm9y+65BOhzWOvwH2Rs4vzyKZOrfCrfE/KwH0gbAGFuuW+axa3Rzfpqacif3qPjzSz0
+sjyQaNvFDEFss1P0mkEXOVGPMZDVKFI9jARVa+QuqGUWaYDcTmr6BrPIpzkkUHa5D0lVVbf0TzM
Tt9vKQk3cSP1eXeyuG+FPcAQP5nw037Hr9rR+wrsVIfW8av7d7Q6pk4EpPG6Bjbx0uB9+DeQfQB8
9nMfOmj/JqFKiKTWz4YwdD3gqHjWouhEpW+Ej7i6hyPLTUgYLBKD61/lTDJJoGbvmFNMPg9SGZLr
UxMSLiiPnNkQUQOHcWon1e5nsJ4h5cSO+vH/lljnO0XS8qflwTOZ9g4bOYA7eU295rpab8ihdXtt
y8nZqj3qPt2SWO4Lct5r0y/xnw3poSkKAbHqB4CcMmZHjYtKgvzX5QJ1rfRILObikQ2t3omdfv/r
DIxksO4H5z+m4Be+ccF1U1lpFGlqy9xu6OwePKhY+y//DvuutROVUwhig4MuCo+w5QdOtjQ6WrEa
D19Yo9v+81cCV+KVmi4VEWomxII+UD2Wa+EYKK9IKazrynY5A3sBzxoS09qjq01ft3LwnLfBbGlb
h/qchajkoPqB7Lkd/NwJTauc4ASjxYdiGtpMppOUb0SGbx/eSUD+1On0+eyOYDqnTATSHxAUq9Li
SoWK8FKkIq4z8A2CVR1OohStjQhMOSHEHAS484llddNBV5LkYF9mSlJPs16hyXt+0WX71Q3y4XCy
ue+DGk7SQd8bapRpPKCZqXPJFsTsd8iRt00hp0qGRTqjQPWDILsbwrt566X/0XlaviJqXJPFwVG6
GnXrSiYLD1vgyXWuTA+aNECMInA5vLqTvAzf9PKmu0j9Y/2SvCcWuJrJFCQgdDptZBs+d6R+l4LX
cmzOH8M1Om3vdER2H47d5a6SseGQKh64+x09ijeIRirXpEZjSHFRKFNnQvQnQGbdh80unUPetfT6
7ouovkTcSHkNLvz8IOLwTa99aJf8uuXLehi14phLebKGOwy63hLyYypMtlHMOFpP30cUhm7GRqLS
wKc7JOli514ZFN3S3VVj+m1MOPolrL2mPC3mHNGdEZF9FSafE9CNQm1/PMpYiYXEcjd6hc4Xfb2V
2GQdouS5kiTxvhlWL0f/NUU62zMDjHEKTXoQkkYUlBMvFom0e+RDwukxTutBh4wc5JO+f1Wjzzzx
2H2cMphy8nokADVMtPRBUO9MuO0aGG54eeX/UpqqY9tu3UP5ETp3swdUZIx8HVaIbyR6Tg81z32V
AS0tOQRY4iV+edZNgHBem7XmVb8GCAyOY1pQcDaObKX/qF1sqrs+Jrg4TihlvR9dB/OIoRM07XOs
TZwqdLfo+zmCPkT97i3ApKWW+EV/zYw4ZjyMja34mu4xEStJyx9Ok3hJOnBnyrIpd0BJFtD3eSWk
hGghHv41EM655vkQeplBCIcB0b4iYXE3dj+MGloAkU1Qqd1gYJC2cPAvh7AJYeSZIVRXSnxxV73b
yTRoxex9e8MWoH6l0K0SkpUorYybdsp5n60NaOAiX61RzZmDo010N3vBSIncw8jFJzIuxmkxIRFz
taWY0A2GNPu4EbYjCTrbnWLZwmgbg81xMTgzZF6jKHg5rTSZKfA/aZLXqWsahbg/Ys1GFPELx9cS
d1BhOFVgsoSzfLO+48K9pCfwKucqrbM9pJp8fBRbDTiT8LI62JjFwLefZQPP0vqpkLIUUn9uC2O5
ZRNSD1dP76cdngW4TIfzIaPDW1lmg0Os+YhDFCRBzPfkGkZ0jLxqitCwv/yCqa84QPbtudAiI0Ii
XECYV4HgCG52/QstgyPN4vN2yVUCoGTD9HgqO3iwYAXlg0UqOVptsS9FVvLWfg4XroqFlmt9hH83
gTzbtNbN2V4tOkuFZFysW5xTWzAPq4uoo90O6FFSU48G7G3HzF0CmEhhQ9TxO5fAULs4dnOYb0sr
UwdSAcF6iXja5JyyloSuc+3153+NKt6mrlCBFrTmel8IGhrC1Ij5hcbJ5e9Crt8NBcWc2/+j+ix4
IxM+vrCzLfneuVpdALbsa15mCII6wO1NAPlMsaCLg4O0MGEaczVEfU1be9hnEZrUt5pZdHYxIYPt
1EJFcydd4pDtRAdqbhB7jN4eNPuExXc2V69mYDhCeHovW7IrTtd2RuEZ9/ln3MY1cOr3U/ef91X4
gZfZrjLWX1QECiqtFDskjyRkuDLGNqeYwnmdK6qTlhjdD3cL20zPtnVVEtJgM4X8dQhInEIfyXv+
ked3i0PoS2TvFIZ5DoVtpo+PMF329/DqxpL3/40wvPiw5bXVbyeqk+IsvnSbu2udLrKkvrYeJibm
ks6aBCzqDIFmsEos4pxY+Ax8MNVKr+ll8+NUdeoIAaWPHdl08aM8RaGibfygVdr8RMCdA/U+U0Y4
csvlEJY5JDWwJygSn2oBdXYNWioNfYLhlU4gaQnpJYaYquD5NtYJQHKyx+WBoQ04BVRnUmTInDNt
sPClALZLfXvvHmuWkSdXL4DYl3tToGzM+HCl5ouuc1uF9sshSL2BKgBqUfaFFqVvdwMy2MonA9AT
iRnS+j3d0mgBnH94J6p7VBVIwJAxEtXZR41sdX9UUPu0IYeAtypnART2NyoYaVvttLp3Y6KI6Kfy
rgx78KvGPrVN0G2R/1BmeM5xsL40afdsnPcHEql0Nf58gcI6OlfRG+F9fUr1kVDdssceZC/zHOao
yBlyXal7XUPXePVEhrNXcL2TtOfAvgdpWGI/oYP/RpxJGdJ/zkB5l+FTtIDTiuTYmCMb2ee6YIQ6
YBe+qs1acaTxNKwfp4tHCfrQLy8pkVw+BC90K9EcSFnApnH+TlNjD24bALUkbrL1muuOy4ind76z
3e3rK9ULwqcB3/g1ZNDBE473QLWbt3OkVbW8YHTxRIT0xft042VLJ6cWJ4FAqKFAtdO+t4VYQE5J
zqvQjkotur67PwnZTA62m5s2+W7ZpThrj5WF5ef3iml5C2O7+s5LkNOypQWDC9ZlgsSq/6PJtnO9
6eOZtwtYSQWYm7ItdUNzkIsLFzGk3O4tGOAV/+jqwMU2nKrQZA4a1fG5Gtf61HDnBO7sg0K31VMO
3VxkUNpndoswJxYDnYP6lU3zItq13UnYgI0NYkOujQ8x887JuEAUEv5Cqq09WlRJM8yBd6yf8qGM
e2W6Kkx+KQ02E+FklDTcjLfRMrWUPHJ94QuBlFlLC0RD9SOr7X+qHS+/fEs6+phgYI557m4XanV4
z/UDSUjn7DqMChL+R7J/6ao89xtmrCnFX0m69xUarfzyQ2mu/02iSHO/C0UK98vvO5eMDpI1lhDO
k5wxj6Mouumwh6RAEA3QlTnm0vM/djEbYo4G3uD30EKhtP/Yu2lXZTui13/wNb2/n5d1NqJ0BCMA
/u6qKW3oHyMpCoF7UjavJ7z8E5WP5kXjP4P7ZiAZ7KG/RBV+ES1OTiIr1iIdo+JNv/aUACZXB6uh
3b88C5K2yown65ULYKgF6ru9TYBJXCQHIrwnsErqf32Pjj5FSu4Gsp5NWqj9y1hSxGfqyyT+ht0H
JD0nPrYZRmi8STDFB1NUys1NglszkQ1X4mNZsDhNGW4SPtgAqoEcnhvQm+ldiY2Jui/bNcROojhC
Zcy5wivhMEU7H2ByEIJEMsnS2igHybjmqa6Ev2BkkyobC5U4WF8yqijhdn1B9wlZ7/kLfFYWVANp
edW6RMfetMrXXQPe0KA7c+Tw91ZqMjXPUCUDbrvm8mSSSjDichzcwqthUr9JPbyl86YIe0ZgwBAn
5uvWaMAA57YKLWqVxLKvoHICjPAoYMINoqTVygisJXxQSkBgFe87QhgCIs5VCUQZjALnkrykpWSG
vMTAtSylK/aqlmczFLrfFrBxrAMoIT2dIwG1igk/ShkdvYwIa3MSTqcnDS8cymUVtyhRJkYclTGQ
QsbHkhMxB8dZ80Fo0SucxhRUmIZ5UOO7cVfMOmQLyeE21oFNU4zMWsQ8N0sfe8dXX9kzPEoofaVA
0Au5cnBOnV1a6SLBxZ5saH+6/rSFINhvTncbl49ix7XQL/DKQjRht1vZHF4+ForjOWcVDbHyl9Ps
3XG4Ov6mmRzm8i6+I8Ljf98+RrAJ9hjGtiE+vOqWIiDKgdeI9cTF6GptGiwl9/2A/KZuOVPwWurk
u07BMSjVMsdQV7YNykPixkVypnJZEW5cTIyXs+f62eFr2Dw5zSdSSjtWtLNpexDV3v1DePiERBcM
Evo8jv/LW/4mLW1GJL3U1MzjOhJ7IecKe/pyhtnQgFHvcvez1jCucq5WwGtQ5A9gc75+0znVitlP
AM94Bbeq1fxDTecFwKOLAtE9XCI7Q60rp0EejfE/QL/gPxZ9VB/lIoVF6POtv8w/ELeKuhSzYyiu
JB+4OcqO77yBu7B7ftOGQ2c7feWy3eDeXVZq9AQYOzGHYVQf41DCyBI3cwmFgc+YYUqqTZOqyZcV
WETjbooI1aTp+3aGwmOcJx4qN/ZFd2nsVHzQzhfr3pdVS8BrucgTNoJEU8jBM7c5gWw4UPQ0GGjW
BwWqu0lPRuWK08PEfSHuhDxN6oauC2zHTqm+YmwIlKgtIKWEYSnns9lhNsykbnKdvq1KD1J8Pgyw
jaCoDnBlawxhY8DBP3l/ZAVptsRbefcKp6dAH3i2yI1F6FeFhkNWweml6DP45Sd+U22W5GoyNnpg
hQSDaFe82gWn3bPCZNMADod8gXpvWNTmq7l21S3iQXiyP82Nb4m+Y8TwOqZWc4iV68oRgXzhEAIM
QwMqb9ayQts2hj/YwbcwkAVp7E+S04YWF+DcqmYbIho7TvG7NXbYxnkUiy0mMaaDm3wdI3AEMyEw
puDPycdJwKEVYIzq6DhC0x1GozmEUoH77tRDIcgESc6bGAgcbsxDuEVsM2yptc5aKpSi4BDMbtFK
hEkki+R3MZxzwXYouiqVZx9wAYAcHK/P8VLxUIL0xC9lTtk74kkSVOMaN7fTX4p+fqht0Za8+iMg
hw65hvULL1eT94whpxvdwyoX5noVKfNcJlYcwjpI6l8qkZnAT/jZGGxGDxU8EfslscSiIN82yOmv
7Khdhc7EXOtJG7zMEh8+2QEYflDnWWb9XP2lc2nfNcugA34XNhPELMSNQbK9u5rjwqLApMYr4MVI
L3lauDCdKhfVjxJpjmeHWTGlpX4aYZS9Jn41ewoK2TAqs46gyM3r9er6Y0xSyJu/DFq29ekoV8iw
wgIrOAUD/ak6FoQvePuDaqqcVGGXM3js0lUGmvsTrQHESMVLYTy9Vjx7Lo0b69Ph+KaZVgBrb7fO
LGBpXtuAmVjShWrl1oYXnYJ5xrIwHJc9aXWLawdLhFyTxS0tLSgTj9Lj/lBaPmod8fSn9BF7WX5U
HH8CYnIihmhW6XvPybOyPogGu8qhBeZFo6J6fxxieQMg06P7CF+ZM4FjYVWVCL6XFnyUpR0RCU8j
Mw1Zfinz6igiwXymODCBVds6oH4gnnL/7pc7gwl0oVAMaMxUk95Aq6iLxII5v3w2rjuk7Z+Ib1/r
92UmNOgeu9goiSiEbioC1lpFEWTDP+DGIiQhS5EjGvrn6y2Bbd6NzfYJw1+/dVzJXm7VSdHbNZI6
h7eo6aMyDxQnfoOKW4YAb/Du3jNyd8TAHFKdJqs7zf6KlWLy+txSicdnWjwl0rWmJd2ZDAah26/U
6XEHiJz+WYK1iZlys1e/GHs3cwLljNZJfozdjEEAXHUcVw8FLuMsxFPTVf/aZK41LfUqafFwP5gO
+no0SU91Ijf9qNtAjkyGLELHKZvppK7H2gc4sGHK7FLPrAE+/2IhwRJrvaRVxkL0TmOcZ3UNu91o
VBfISR4ii7Agm7s4mFMBYlAFH5mc+QF0PbibpG4XkvCz/t4sZ7EhBRG3psQObhCGRtLfInvs9Y7Z
uR5NsAQHa+on6QJoAqrGdr6WYfPekQpzc0pdBqGHe9/QEdzP0M+fqkoCp8TCH92D8DRKSiAcvHKf
RcjOaSdUPP4ZGvPIwhrVT5N3DMR7i7B51qtbHGDu9YKFXzFNOSNsNGh+k9UrMG4saG+5y2OZnFcM
Pxp8+FVm3MCem8YJrFuAb280cmCLKOEN0VzfWjdc1CeUvpGNfD4WIEbnchYbFsYO8ZkVQ2zH8OP6
jyZZdQfgFsQipeNl9TVYi4e7x//K4CMCC0GOrO0bcIkYt1YVI+36MfQD2JgveaO7G/OZNj+vTeQM
1wI2Q/EIFKdKLO3tufcvZdBTLmNbWNm4Wah0gsmZ9bLe/D3nrX44aQMAuexAaJBiaGzd4dmkmn29
Ux7Nj7lZONIO2xWZxtMdvekYsz+0xrxEIedYoUwt50wyFE4lVRH2RAu35D9cliZkOMtN9zFfENro
Ym/j3ohsseF1cWFDkInLvpcmioeRa+H8bx+1lwVs2EpIPIxf7XSPh9K7Oz4ovdUux7RkheX8qKAR
+2DQkFNShxBOCbBFXlOnxg1VG7QunPUwqLSD+t3tAxCNWhNBJc0Ij/kW34XfbPewWvfmcAftZkkw
2V69l9q2br+auEE9uNpAuOQpoY8cprL7NdprCHF42QJHOQeUvO2LGjJKuZWT9c28ANZmxJwS++F8
hP5HvNk+bsPn9e6tvpTufCob843nQeWHdUSENyIyqdbHuopjsB6hJIm0hjhxFhuGrCrI/UC6xbyf
JbVlJkbDbSoHiiGEc6ftg2Ok/vNkSXEw5LXa3nWKjHTepDWef8+TXUy32ZFyGXfBZG6dBodbIc30
ZwLxb3xZ/9dB4tMScS6RW7yi3ban4IETfBS/RH2eVOPm7+1orMCWk21HVNiUjsYyT7FzMvO2wgE7
oEF5/Uy9byceT49/9LGNVSH/Wen9oRA/1njpuwQngOPLbA2DCq9Ald+FMQDtmz/pPrk0aSRHaUOg
vsQwXnY+D5JvqFgbqpbA9fZK15DqCC1T5t3BgOGXCPiaN5H2NLORd1UsbC3x6ePRr+p3UOuxwizp
T+5TAPa6R4fI0V4PtLgzd8BRGEp9fkizWKdZnd2TkwRs7LzPebc1SlXjBGhab+Q8quEkSDgE8V1v
xmmHEaUiDrw+6GNuPGRqSkFtRQkQEh3aFeJipFS9Xyp43yb9/arHc/dLlT5wiNMpo1OBYq+zzJ0a
z675nJ7tfF4x8Z2sn2IZpp+WaWIR47R1T4sHSgTDGzNWknlHVDfZ+ZnjYYUZg0zpj9nf3rmPERbx
HxR2KS5+sZqDCKnMccsAPpPo1MXuzdMt+TeUl5awEhHBllHubWMCjoGEvff5ePmwssW3kPpjOafm
I5szeb0eUE62NehYQHFxLKtOFWbjOrYAKyjJGbzVLLGlz9EmeW5h2WlvqLMixd8sY5+dEJjmco9l
Le9Kfs8K1Gvx7nSnqXhL8bSj/llg3WRGCHUAM014SzmVATDt6vcepdR3GR3jJVpWJg/q5XbDNmgs
UNWOc130aM3hwRLmxte/bU32nPNlPqT8k3LpK6sWjmrToJ5EC9NsfUZfirnIWaAOPRCb4WZz1ydC
fZQcsc2wpOKqzY8RXWceTmg0yLN52Omiv+oJkJyCiYl3fx60CM3UeFKSHCOE2ZCCI8uhHwSJCpo4
Ok+Fmfe7fOA7s30LGcblRbQNRmpMvFci+89Zj2mwoE09zxxo6p+1DunzjwSVoS7l/cfDp6roJX0o
V3RltmCwZp9Ar71hfResb8/ZbjzxgRzfD6EJBaa7PGNTDg8OuFlmgG0hmZo/uKtPRippfHwi7k4z
AfVp1hiz4ykPanQhI9qFREmp2QsPhk0RQQJ2CXaaZSCwmu/vr1MQ3qGK+ajxqNW/HDDsItq7l0JF
jMgcTf6phRsLLr4+cHr6oukXvmkNxpTrzAZghxTvRKAPUgHtEhe1tMjmj7moaE8ZJYpS7hr8ZzRY
WVtvenyhgTrbm/bgCtS0wT+i8PlTIKmPW+z/zog7tYAkTA0d/8xAScgSCjt67jgNXwXK6Ifga8Ia
O9JfgbOl0VE00fOQjCAgSsx0j+lN9Noq4PKqU+uX5opQ6P3ISDFIWi5N7aRlPoAPK513keZHQsqk
FHMhRYnaRoHTGNHBs1VVMECroLdEbe7lIxfmZ1yGiE7MtUKw0mW3XtsLK7yzALtaOVK3qwipjnvZ
s59kFkLvaz7CN89NMArLK02wGhRoVVN+zPUxwbokLoue5GykUxo/jopeSglh9X9DID3K/rWFh/35
IwQWaLuif+T/lsyr6JONiAOX1bLR58IDMwBS+0jIxJvEjiAOBkRbbaJOZaPRbPhAONuh2SHUneSH
k7laLuKqnkK9zz5R6ecmByyubGWfPOBbdmqFD1cyWDVCFVTuxBSVnLWhgH/uaZYX0kzv9rTUrdn1
tGFOkJR+A6v5e7zNdpD7cIgBwk9aJIk83jQaX8m1Wp3dOjB5fvghLcG8Aq7qK/jBl1kedwGP7Urs
p8tc/7zrLSnuX1+6lfxVU+9a/KlJtCwtJTVs7APQRKamG5ExiNCj694q1nJ8i53nQZMcI/OvPm56
QuXejuVJ4E9jrq19oZwThDR3yQKd6xMrd0apfN9/5BvRgE/pz6RMwpzIIQgqQVMr9gAlg+I133JX
7sOSDrVYOubHl5a9JZsV/HDHPP9vKStbfU5IRvrm9oXolchB1iUJpA/7Lb39o1BQ0qWYKOn81SXB
Q9sjfPj7wT3MLnHLyYPPsPJYNlPoBjcvDlU8V48agwtstN6e8Ojz/DyxqcUBjs2zPrhYzD5Aw/T8
dNS4Yo9rrfA4nVzGVPAGe7pv1ncXb/nWskTPS54N5H0/+a113+WJyJV42NfB06acjyay9ts3xhJO
jZsCzgjFGiwTxMKCXBuUpz7iF4TI8cHvjHRGzl1yfj7lEYiTUOQxgYsvWP0pbiXwlYfPHOzyFmD9
c+qTlPkESFkC7y4icgSElxsMwJeTRtJIYTPLE0BH1sW0O19x2SjlbR9eTqInRCxtEIYKMicTSJFa
IiAvzGY3V9RpvuXRcCjIZRku3pLiEj/P0pkHvKTHLK36PobdlrrndQx6yccNne6hVSFfFK492/lj
YgDPLc9/zv5aIbgZu7Aadka+e2Wrc9JkBOIdBNIJ+KERnqviTXIgujoRTnkgTzTtOXD8Q1zS32kM
R/hdMTo3bjzvKAe52Cm9+SOdTZ+0kFYsCzzhTuGqW02TKUkYgrp2BdlIfe5tt4P7wdkGSEFc543k
il8yI0VV0uxl66jj/vIYgG445fq2J/v3NDm4aRwGv8ALGoT5XNIGW0PLHGyxjG0W2FfNCOuggNWx
kaB9hfL4NAc+tJjUV1BU73p88B1mSsAci5w2B8fQGofw/BoEtXbupsEXD8acyl1Fqs5niLT1zKal
8ni8nWd3EiuATIyB+w/+UOVzqcXgC+2H3JA+dLeCyCxCu//dx+kWUfEWty5HEAyxgjw23Ock2wR/
+UDWoklk1f11qTH7si5Lt5kiGwwKH52fCSe0PTYJglQXlqh5FX05EFf/Gr0q3M3tfOWbUSOGDIE9
4VP6djvYEopxNYTdJH80vvrJyN8LX3uPDXlx2dLv+TJKMig6JwXXrq9XyGoxfTDpDji1kt3ElNhQ
0iVQjvX5RyHUBRtrPIsZrNfVBgOYNt3sojuwQN3CxDcuCpwCj+zgDXLa/0nTQpRiYFRqdCxMfJ4a
8XDmpGGQQqGJb1TgCa12mHHOodkE+w0SiZmcygxgOQjTr2EcbpPNQqK0wrUdQLG7tvoI9yIAbv3P
GRZnVZWeO/VK95w5FbLgEiwyxQoZ1a1utsmPn7qi74Lq8M8xX7NOW/8L8hBU3ebqoxnYvvvI3myg
8PyJdbEzyXO+BaqBQCfXGUUroPnzV85rpCEgfUF+X8sy9/pYcX7dvgr0tyPGZYEOBbyCrt/O/As4
l4AMjGJjXSbsSKHaC/TbIZAun7SuxvK0atx5IAoxHBY6s9M+9ZaDi5cVC/8Y6DMjsmwaVUcoQN+0
b37TJ5+Dy3D/QTLtkNLYLW6zhYnSKAtE1o4RrwzRbRDMRXJYbOOyU2zsD11kClTXkh3LC+NJ9/h7
kLutC9ZAg3no6SIuGLYyIVvCFVvyEJ2wdvBIsdNhc6MWJzQlbyRiSdPjCjlM31/xZ7QqH+fUO+Z3
+mgVGgIUS+b00/Ik1jhmBcdM8TKtcPZNa7fAvq0M/TcOheOcXpXVMool9byoh3QHHJu0NT2WTbq/
OFJ0iAQLIWX+HZ+grTRHEhuduVjUMSdt5rN67OpP3YU8O6Vo4gsPgkxFZjKMI/yPWY6lx0+87Ier
UwnGICLUlKTstfcO7yYa54a0W/3eTD0ErnaLxDDYOWTlAnn6r/487VBEfi2mEjUh1czdA7wcytZs
hNqws4QMKHrzKeZU/yXQmW4TEjrR/DYO+R5MpkOlzR62Y6DCaEGVDjKrlka0xrN49jUkvuut+wZr
34lnY6fu1FC4RGSHaxDwMZmsa05G4VpKWn/eG5Y3d+thQd1XzgZ6kzMTEWvLkTrl9cxAP+kjO3MR
kl3Ua43ISVpS7ii91ceVjJVwvBZwI18EPgPwFmbQkfrjJikYyyFsxfSXUqqIQ0xEODGyX+Jsuhh1
5T2xndfSsyjxHZe/oSZCyPv4dcz83PKASyaN4v/Ag7is1NrQDBfWkAj4gNeKfyhf7gsO2jiB2AvL
VZeBY7amhuWpONtszrtI4BHVwGbgrHd4+0ky5F2d8bTtHUAR1VCoUvB/9Zu71+czZv9yBP/yib3Q
5QK10lWimCP9e/RsZnQ08WNpy79sj3uXbC1lXpyjlcNBxwLYirF/b/V2jBo6p2vEdl4CxUtbFcrV
D918Q6Qy8Pi8J7GWZZC35UKuV1ysFkZnOE9LSWxMIMdJcsWIYVuB6LKfgwwWPRfWUN0xjCfeJx5z
F8aDHPwvi58oux0KL4KL8ZgmkJ1SCBp4l18bUq7JtXk46iXFeSyMro0ZEc2Mpoly+3haipt3ywLK
T7+ppboDIqBblj6agKOmrAq6pZlE0AOdSVwKs0RRSf7wUPo1yffaibtUPD9W1Dr7ooPmcjLFajOK
ycuVxM41JycRupAzs5V+ShJi86m8pBkhn+iwa1uGIzWUbg3xii48tfaewxupxkKyNpDKG0mXKGlw
RQPNWQx+XCroU0IQbGt2c0p16c5OoXTh7Basb3Wf3w+AVhDrTXOuWzatUOy8niju8s03D//b140C
uWWMnade1cV2NNjfXsYzbUzicF66wsr8RI23c95A9MGcExfhTYYexXi8AqlZ2U53sY9oV98CUgRQ
zAoqzN/iVnCNmLNYVvtGn+xgFwPp+RKkNhBy4zx8L6kA424aqphJje6AYX3NGqqjV7Tukc7BdD6Q
h3Inn57MvB4OOQwHDHQUMy+KPp8rKtzGDHilTPnMl85zLNQsKfxJlf2Yaml/xdfMlU90ouIz4s9t
KMXpjczYYazCivxTIEqr5rbz2oU3SxalQI0slz6aRsWknOorEgC1mgDlXXukIPKyP12GSCL2rRvV
6SrkW7OfRhO1t+P6dAf+lMz/WVzPsgOpT6QFqcIqLnxI22XNZc/u5zr3/++TB6ZesHsTW81Xc6BU
+PsXdrVwGRq1WCSuPhF6TBzthDZWzI71TH3GOIRjByur9LQQe4b7xwMrQYs3f57ULhtaXjC+OsUB
YVs0+W2+xink6w0AVeUpfIr0bIYGypZpfO82CV+GIzuV7j2fpwCLqBZPQdXaFuMug3F+Y1L/M5eq
SCdMJt1b1yWVDAt8NDFEUrIbe/dlSbfNPr7AQ2zdtilW9ZbDaVFjXS+smkoQms2otNcLm1wLmDQ1
FcRO5YbyC7W63YwOG6XSeh8V1tdZWHRNLrD15DdFA+Z8KYepm5+3HmZOqOLqPS8dfj33KKUyUO+m
wbFLyRRRTJWVS+3JxuZ12lucTemhEO3JFp3+c4SaMoQsER37TREgrMZc9ogUS/Alse/lTZlBmLs4
T1aDnAMKveDE9+S1AnlD8X+TFK7G7d2WFrSqG3WiXwTOuLGtoziSxviSq7UbnI0+l4jqNA1t49O8
qWhg4d4CNgiVGKst9JbrDcsEC0vE82XHaaPhkRta+AogJ34Mqjz2+zubTeij/lOM3EYCfy5B+4HW
5z6ezbJlEC9Vvpuj1Vx7D7pb1tc0ch5GaJfdO8ZNlHGZb42hctEVGgYPY6vF+vAfMsskCVUlYQKW
HIc5GSLbL4qs5MTEnMhUz9AYh3XXiw5wipN5c6JBnj3u9yh3QMXisR9OWMqyfeY4gdhXarWY7i5A
srwBw6K9sPBqK157uC3iY1lV09OAYbcKmiefbKZxMBJdicEVhzj/61fUzooSEMRy7PSWQUIQtJdf
xRN1zOSx8S5Q958T+eq1V22RvhKoWY/CnZ1XQcNEw/FwMOyb7p+2BOiAhgF/JEvONYM2+LSLEi6l
RJLLwUrNuwxOZi9NVy52s6hQj9zfBrez5pZoio/h1/dCdbmBhNB2LPODXz9GxC9PfwPO6GeJFiD/
TYqagZBQnb49GLdoFC0Cdvb1B1qQ67vRt4+lUg/WoR5p/vWi5YqFUEERGr8lpeZ9hpu4RP6UHky3
3Xi1A4ZCQQizMKDPwEjR6zl/eWNNNudW6Y2Ow/T0LeJi95NjIhKg4HwwpdIFy4HnDomeE0KXNPdZ
yxQZ0K3iPBZueVE4yVjmt8uRnX9eVg15irOLwRnT0FZo9Z6GTpLL9ILJv9iIjXzfdGxyiDDNBTbq
T9MLkA/YaTVaK9EWCWpyULBPiNBW7Bg4Y9es0Xxgj+tDlsrIL3foHjTV5tQHnV4vJvO7/csSDehA
OJOnzkWw7Yyg+yd8uEcTgaDWaKzQdSOAIOMjdKBNuN1OXmVLdirQI43l6hG1C7bT5e7N0oBE5aKz
+WKxDz7lO1iEZXFtK9JWWezrk7RGqtZST88A8u/OTR9LFc4Q0tE8Jq6YWQJHIQyD/zfXl5Kp1XkH
sesmtNcX8LwdUHStNpzj1/Xae8zBkGEJjp0Ao3pq2+T+te8ksGmiqe8m7A9mudjPuxVUFNBAjbCG
X3GrWsAjEvGuty75D1U3yStc3/jqKtif3P4OqQ/ExMd7M4R/WS0AMhQlCH1oALVEpkHolkSHJYXb
npvQbDENEaB7CCYtHzRY/os9KDZHWXwwO0Js7+oU4DgTMikh7kuFAq7XJi9MhYbdpOxb/5ZXUvFP
ecC5TXnqDZxHyhIERnDwtH0Aql//gxvVhz/tcfihEG9mr9nf+VawP0HEYhS4nuX1zRKEBphTBZBF
pSm8mxADj84lQV3IxcjljShmO0NMdzpQBcF2ys9oMK/gUT80AP8ptXh9ADwuOw0R1RbsI5L9SKFR
sJVdjcCiLzCemQCvY4BgZOkQQAKneXGcSm0rqabtPFl1v1bqBrFKv/Ex/0whZHV1v/iWJuNdm9dF
6QULjIpmadFFUW1mKhfbTOvwGdJ2D5K3Sp6q7HPTYgY5XE7nrlv1OR1wN2cpiOm3uirU8fDoBuBY
XeJcPYimui3Pio+lAjl2ill1oENbSyaa+oGBXx4DD3+kqp4aJw4NrecbWWcjGrE1J4EDv4Eij0Cy
Ohu9bhCpeVZS+6kHa397h97p1WgtM/W65qt0waOtSy31Gme23OC9VeombmDc2rqDbMRk6N7rb3K1
n0LmPBBSTRQe5anG9qAfH6a0GVBbiDqVl8RoRobFpZahX160kgPOtgAyVA1PHFUL4rumwVdiJG+X
ODK6/7/RE5+vvmZ51/GtJQdnl5AQ5DwCHpP9+N28JSkgeb7+rvzSnNo/mChA2xbgQfeGwLwgNKhD
GAbu/0frp2yv7wiy2dzc6YqS4124KgAEGalF6o8EiUKdSzNMfJoSV3A1EvOh+jbqZQEtcKaN4K6p
3oPkyX6F0GQvRssKxBXzjdIzjz8joLbSmmkElS6WrMdM51eLdNCU1C8giLVv/Ia8kJEderBhqjdM
nNCdDd42RFq3sudzb6xN89Oz6zKdnS+bSUArNPAmyu5DCa2V/fGot8LnIlJPwcqFVpz/ZmBMNhr1
RMCgkHvHUjGsymUIpsxVB1Gi952RxdySMlCXnzwhs/SbmXWu4QCvgyBPhs55+OR32cQ7mIihVoDY
rxtpSLIvPz9I7vZKCBJsfxX41PS7oMurfOYyF0djV9oIs5gJbLDTgvZ8tGdQBEU9zSwIbAFaqOxB
BBTCLL+xTbfpH5QDwOiZRIZr0PYQPGmklcQLv15LTPh0ET91/GFur0P5G19uJ7t0i/UklMwSRbNR
+8H1IlO0Bw6SuJbukf87RUm1Weokf6nvVIBfX7OQRap9aqTgMs5bdERkfDwCRLGTI02ksgGpXwU3
g6CLHg4xAS7b0CvLQjN1/YaM+5UzCS/kZTkDPDYT5dR6NP9YUxb5nT6lpFHSjjnBRyOlsC7FPY7l
O8mYuWTb5+2W4LYmgrSv76dVgL/evBuSXwXcz1PPGVAXKXlGyVAslxcuq2DmvwFp4vLeziTlL9EP
nxe/fj5lysZxBC+ESY5I52iwdK6VeKuBHQ/y9kmMg9jVVd9BR2QiWVXCd3PsIvQO2Q/LBmpJBcVD
xx1jUfblqB74mUwTxk8/HQwIWGDhhLtRRz7jECHW/jmHRK5B1T32HKdqv/ALchgxHt5RGPDTfcoJ
abtuB8E19+XuQ4fQpy+S8YVcKgQ3rncFE7qM4bu2ICvy3teOWkY8Yf2Bikec0iy7EfIs7rLxRISM
HAHYRN0f2dystKI7pIJO3Q/pOYVRKZo4W8U7v4Krme2g24O7rvynMb+HLvDLXYFoWPWFNjhai0a7
rxhewdZxK6MRgs8wrsO9ctfm3FNf5vIXZ6IMj+liclIM96r1grSahO8ie6fJ41Jw69OcOel+wJSv
4lL+OPGC4D2cXdMevtd3GFQHv0oq97/v7YdiyTmH6sbLsz1Pts4kX2yzCNLe1XPD92zA+7gPn5zk
4sis+aNb87/eHrNRV93gVwRA6H8kqPtqvurFZZf35tp3RTyIAqgI7dqWv+R7AhbBijAbPD2T4WaR
DqXFkRUIrflmxDwMt9w4xzvK9Pt3JQOGcJgM5h2wdsYuoJW3xc+3LRMvULwg3itFVEggr8cSkAvu
RP3w1/9ORCyH1bH+BBGVnxfLGLR+owBzHTUSAN7Wm38VYD0EZ4mJyNHC2tVHoj6KbnplSJuanZ3J
YXz1e/nr7iyvYEbUVHVh3vvLgD5LfCcLit3Lv34ylHuFcRNqX4uilw16tNyzzdCEzBAPZCPz7KVU
J2XWFUo1jt2o9Gd3mTSgs1OFU36ht959uIil6IMx1xJfDDcjRFac0alsy3fypR+iQeGdkOP0O8Vx
YQpuBFXaxqQQ3g4/7bQaGKqgbZ4fZBCJFv2LQVOGQ+1Z9FU2NiLLB8JmNVhuZRK3cNKXHYI2Akcm
WmNm5njrqIG41he82doVl6lpIfpArYknF9KlZ3IhTXMriHTiHtLOe3YK0+sKEIRaF9R9yI7Dclox
EiO1dQky7zC6fZrINZtNnRWgQE9AjNaknKja1UhQ92IhaZoEntvWJlbkIqZzT6poAN1PpYlIe2aL
luvYPKOo5Xqgck2f/SKeOPzZ88hp4v420wOJccD65MMX6pY65HlwjS+5yyHt/VrFBBScQFZC3tbW
+umO2y7SGHLID9LZHxX03bzcqoqdJ0HHQkxf1iJE8WiQHjApRlBmDznZYwyj5nKQUKw2gGV+r6Rk
5xFU2MaUoyqseznfw6sSf2KuQoUDLY3qahWstC5dw7r7HYglsX9drG99/LkRS2Ir3LGGt4WdfPy3
MN6PRpwMh2acGA/jdC4hxfzY0pjvUZdYaxWthpqUXg3qdEyQ4TfsYOgyntLCE1wyfe6UW0UwXDsE
cESBJTYXJo8goZPWMhUwrxLI5KR/fYsoV4sa+jiGLttzhv6zdV+FjfTGNIcJULRUmlcFtXDw3q08
m/cFlpfxz3GtiJSimyirGpoqZPDx5bHtGaRJtpTYEk8qfa76psKDRYuOT+V359P6oqYbZJ7xXDTH
nxDq9nfv+IryxeGvTyUiEkN+byx80ImPzoLFXOH2K3jdHATWChgP+j+Co4XNNZSb6CihtXneKXc7
FTu6uEhdeJWVN33nMdf4qJXimIiBOjevIs7jBbGKLEKUoH6ZMuZ4biNAo/PBfjLgyxCKziJd4a01
2v0+LC2qCaSitcU6COMY2BFBrcSNJAgS06/M/woivtG00L+9VyDW59fc4kWSUu2HaQFRW6K1apyI
vdgymQQiRLgoGXH1huQXi1pBu/TIRDpn7OgT8sbRuwAIkGRvALA1jKky7c5HLai1dZP1nTiOFvAl
kOY0svqyR1hfOw46r4MwCLbMySCMnGnuAWNNWxLx0f2ZE5DeYBfiikbKj7vfT8c1qjCXtrKmgrym
1LEYh9rVyJi8IYcIQHv5r7EEeQCbjqhg3ZznjFU4gkM9jaqpFjXoKLgxnRhgCnH+wo1lpYCe28MT
K8T/appalQWb0K0h7FNqHG8Jj5SGVkaGeRALuKcJlQRPdxLfSm+1DE6ncidaPwdy9EslSB17MHjy
esZPSjr8+bD94DgPHIrvINVRapBXBq3zwESA3iuIrs+ZFuwiea4mpvY6gDc4XcOdwIrScDsxwcBv
d7wcRw5QCI0f418Rw21NVseKcfbaY21MJbuBJ8tlwkhV6a7QnwhtzrismW3KI2r53rm1TPZftWyP
XBg5+wpKBBXoBCf2cXlZkUxH9COOSJSxWIqe3G4DiJt8cFLNXTtUdBCLUgSNJHwhG2jMNyXnQhfz
QvgZbTJUp+QkGHWdWl+Kl94wGsL0+hE7MHuOjrtljOCy2uqzYOBK4LVbfWUiXbZYjCCpd0F3JlJh
jJADfTCPyMocPkcKI45eeIl9TZKEhs3pLucIhvbhXrpdnf/ioiydHeQVO7qUZ+RMKSm/IEkeHIW/
bSJehFTl8UhfEXO9hHWh0LMk0I9VYBo2aJwQ5bFaRt0+dLQ066cjlCAfZJo311poY70Xau2VN7Lq
TqrAg977dJ6wMzP9ETUePB6bOY6N77ptIMMOGa8M5tQPri46Qk3wwZQzNuTAHyVR6s1Yg+YrEhnc
L0By/LK80kS03GC88guBmfqSe7OE0Daw7MybbBNm1HB/DkuZ8RzPQfULGPAR1ZtLuNtiB0q/frxS
+MLjBDfoHM56lbM3nS5niDJRDUMuBw28WufQ0Xd3tnI73BN6aptRservOMMB+imvz765yYt95Rh4
DXevB6S+CWRxD037UlD4xTC7qtJ7zbx4FrohMfTR3argMvaoQhwXD/k7J9Y3F+5oe49Ab9iZEah7
CLddWvmZZHqgQqrymIDqybQw82+Jtbbqcs3iJYDjNAudVmunZ5nff6OHbs0Rdo0RfCEaP6ejdf+u
98jFWB7FPrh+NvUEbZbUQbBroXmc2LFgd+HPxZxhO/ORkP60x8+Xggu9SKH1UDMb93l4PWr70LKP
U0s/2+xCPRmfWKy9R6GCKtp1vEJU3+fc8iJnCspFpHlIbS37JNRKt7GGguNWVpL7s6rzS4cYcDf4
ZNvji9nKSRVGUeIXLvDLtQk2a+ZRsnoZAjoJU3IRuPw2EorPLe5LKTcFctlvJGBqGOcqWLWm0yHt
sulcRjwFuTQPYzLPfOl5th/3z6skxXWoBknRDrdyasPutsVNxmURNeGFnlT+rn3LQHoqlGKPfkA6
8KiLJkPX+4quqJicA8dB0Wd1Jz+X+c0/Kl9cublsijSnbUlZdEriWQI3ODIVzPdeemcqMl3nDgn4
o4It8QkjurQKr9kvMhIscFWW4KqI7MXAYkQCzNtWGZI+shHVYZSoDI7mFY3lPr4knikKRIR3BUiH
cq4+5SObwfHhf+eOurC84RlmosLhPM732G44RmS5HCiLAVbErEYZVbqDFJZIyF7lHxt2oEQKfbUn
s/x+OCGtwNGZeuVlTwVidDSZXYwH+zQslxsMFpyYpv5EPzhjzdheG1fB1aoY+Vv5NZwfjEW9ZdmO
UIOvHvuYtVrxjbzzMjoMg3XEKjpE8slmYwwm4aDdHM1SK2N4/l3hwFZQE3mcSiWeBkM7LH/aixDN
XeExZ0G0jRea0ZXpY/8THmZnrWlPaO3VCk8BDYixf5CwXu9nzXEdX9GdAuJUmpyhmCEaBJH+fxpt
e2NQNsKb26V/mWsgO0SSLowj2soO8VIp3Md0sTlDllCByzuAcaRRcKF92ajWGIWAvutkHdanRCtc
UA2YjLjDp011pk10hdSHg06hW4RxG6JPV6/b8X+aNvhWlwCAFgSAQezFl+WkKkO6N3AbmleRZRf/
Mj1oH/YahpJf9HO7GbgPPBO9Jeox7iLhXF65KuK5m6gnNdYzd/uvfhERDHmCaQerGCanHPmrjpn5
pmc4uUVlyZ+ES3s/jVmvafsIt7+6b4PZPL6W8E3oiC7eXS8NShGw2pSKYN3C6RGljq7LUO0K4jED
vouJPzdo731m2EmhQX/x3ksZ5CwoljhthOE88GYswVYc87BsrOMvshsMEorYmnSVov2kC41yGNE/
TYXTWqFbIuprkZph2VJhy8lfMAOclyfcP4bVXeD+Wz2E2IldauOXBYxy/sgXw+lvHty0ypNZIGIb
GYaUcM6zfvyc9jVXfCGPwzzzkZxZ9bbuxEfUKV+titTWhbu5tsPMqRehAgfGxfqefz9tHUQw6f8T
YFKhFt386KjLsJ9bHSp8BTCQE8Rzv8BUvUY/Np8CmkF0meFwsjJ/s31r3H2UCLaTA0NtXC9CFUie
wKEj+W32SApusxYG6t+tSSx/gtfIutOJjWE9Z8BwTHdXDf0Rm8g+QnOD4Kqax+6sc/6EJHdZx8Wf
qroIufIRb+IyQHcCwK4lTVrIubn29jkum35LWcJYjvWrcUpLBNGEOZItHNGwpaMJRW32ZAVo3k/E
lNycn6hTj7paNp9qhDhn+/+14caf0pwNlWhYm8TJy0viyl6YEWWjFZfeP6b4CXo0jyyHLsHWgym4
akTPZ4OAkOnkrjpOCzFRPEZBAfCovEru0jry0TvTYnjtcEyBw+uXWkcB6nEoZ3Gmz2IDuOgHR15K
ha2cwNlSYdj1Ej83Hx2C/KHKGOJF6o5CjL9jbPcUsytJwu/Fz1AKzM5CYfW8/R+Thz6JwWhvsLUC
LdMY/WMHxWjbelOmeK/rq/ZETHMZN5kXtBauCoE2jbAgFbOBMTH3brlVn73A0Y1AG+3zC+k3QTTN
gNUJ7qJuWWpwQDiqHxlRnkMZxFaM7NhFxzqGpY4HAAaCTl6Apn47x997VfQQkt8B1A+vFQR+35Lu
FEAmOEo0WOIHU+8H7A6gNxuN/1TD7lq20ueW6Y7xuc/7mhiLg4FdArEYkvyCRfeCY/G0GIt0kVl9
4H5xF2YdvQ4w6IsePEQhpYqqzZPUqpJ/e6pL7ztIBDcBwTepgJ8mBS86pYhJfptZuKCWra5QJMpM
AdIWxjEGSzvOu6qOUPbfoMglpRF9yDb956QZHLY/Kp3arLBXuPMPwpnkRija5lZJEEd0GLhX35gT
FsTZx7GFiy4FKXqFyI0RtLQPJj5I2dkmsyMNwC/hqmz89b/IDjwE4P0DFGP0NtBFnopW5aRc6HcD
+O5Pk2ako7W20WJAYyKjOQA8WPKFYHADaDgie9giWCZU7VcGxoRtvmVrNdDpUvkKH3XGhzB6LT6N
iKqSS/G4u8BB+Y9+UbGQ4u11QH67Rwqx5Y1IQe3JAnrA72bnLuFPioT/zqszPkCiRelZQFYZizGM
iX5ji+qAR//0TFAxJnVEhWELm7arvOaAXBoNOT8a/kxzn5eLapz1nqe2Beim+bITHeajeNF9r4Pa
BSmi6sqZeQIPTzEll91MXsVKTINCggBe8Y7LWMGXloO3hRtCviMeMI+Jn2aCK/go76mYtz6/YN6/
L0x5OHRN3kBfMq+qzyGzUh49dBllkwG4xATuU51C19AyL3PDGpdPmBW3cJA7HxSEG77ggZwLIbT8
BHCAkG3PcNQutHnM7tovkLVD9Bes2oXZdeHTwIjamYZ/YmcYudfJ7pCH0MZ19LTQnHrq5+BA5SJn
YSr4zjlh+wkqB3lUp0DF3s8agHmdyitHWzGLxpiL5l90mH8iLi3TptzCp+wk7VHLr/2hAOJpjqel
tXvw/ANDvJehhea0XajDXXaaOEIhXobYwBZqRJVnyZI6cyn8vGzXnn54Y2nSxiy+4qEy1SvQL/ni
j6Ir0OOjybJlDOzgOg+9rrR0BfMY7MgrJIFkEERT5JsxNwKv8BjXHJ2xd7f+UZUeU13OFBY1EB5i
BCOA6RFmUUZRvfGZlfq/R3yQiO3WaIVT4Kn8UIIffGCuUPcO1fnYalTcCFExhBmMMUtydbpNLxSf
elurKoJ0L8d6xkc6Lna5sKJBBt8SiSJ7usqlB02VaVVDrtLuG96Rw1yjJJHJ5xzTwJ89xzKugIOx
b1B4qrM0NJ/Nb7HTUUjxIzalROtXxG/NxAyTq32kAN644tWmaE5pXGqO/efqhsx0sMG/1WwkNwi+
QxPofSSO/VASrQ6Sw+k/UEGgJSzfjWmwj2xt/bows+FzZJBTQ4noR/hsHtqTSMFj/kNX/y/xfbxB
25xfFIVP6NKANdceSN15RfZhBGaw4cBB4+ulxZRWNIqwOGoEAw1ZyYgdm3mb0E6hYg2b0MJOAunr
E3AcHC5gI+sfnAz9oMIVbHd1QG/y88fI72xPEs8g+hzOl6Xq5ryp3B2GLgDlek1UGFE4ZbthuZco
KXjDChTuS/8QFSdb8f6VBI3uzTeXHd67CiU8f8xL1fJTfKE9PkzNCWSOMMaSv7rPPwOLBbGIAAn3
JwaZD+8RIStC2s7a+0KZLuQdSUG3DsQk8Le5SFqBOIvG4QHNsHcpzkO6MqVamiGZpsh5O0+ik9bp
5TkvOpn1gMcMWGBQ5R+07BzEc5ezU6OP7vGiI3FN/DnFcqeWywD41K8vZ8rfRQDHGEJ4q/xShTDh
OikKUuaIpEOLRyOvssB9/KJqGBP1vOqDFlXBuUL+E6hN10nOHcj+vAhHvrYfWHUbSkuVP8KOy7xF
kjaIYc2a0e9c+RJyb1uF/9d1JPu7dOnH2JVA76U6hLRppNc7GPxUHuris52c5/wLJdbsxcRD+esf
IPlbQPD3x0j76zPg4oqobMRFsyU/K8f2z5qYm26URv8171t3xEU94aCcA9ULGZEwz8w9oKP06e9U
SbSKFb2tS1BeJ8frsU8IZcCIv7VZVisqDtoGd7wxlzvQbCJO25veh1A+L+DkIEsRPvKk+/EnLilr
pX4tVMRT4zJXXi5WBgcUgARgzXtjybC38KCrdscNFE/30f9KxJvS6nnj5EXIErwgHNmOZjmQIPna
ZkfRwnRLMzehCMrcxVYDN5zSF7x3Cgb/44vP4f41gDUtPqhJFDhU17tMnoHxTJmugrW1H3WeiU4g
RAT7dlumLt9KLeDH/6Aeai5J+ESHhU7S9+pL1ACygO7lOTiwXvSyhWkCF6hClOY53uQWkyAOrMjW
oQFDbB7qrB0dApswLkVnqRY/p2bARqyGYQqW2JZf9gao6MUOVcXzGqwPSjs321ej39ZOHhGFULg9
Bv6TSE/D7J+gavBzJV9bn4jkM1ieVrK2CLVZ4QAexDzK7fdic74b3jqX0vfW5EEKcSlCBSnimCxs
ToDhbHmBBvUfwhkIRwGST7x3Rz9Ru0C8CTWzqZUBXS/GuXVfNhhz2FWIkDbfcBTHMrj7Qzvxz27R
eA0p45N2Y6NtKbZYUUparTyVXxiMCl3kkO5AkujxClEGIM2L9N12mOWNN79uIqkryE7bjiibXfb9
7JaqMGuX7FTmnfvWhStBUadWVXN5OLUpknWoQZDP5m5kztS+UrhRSZvG0It9kVt6MP02LG+mVIJ3
NnBwK488y0gwFbPyW4aaBMe0wN7NFcteEwVjAU0PpHCP1kvPHp43TcfQmFZD8AVqvs4Q6TALC2FR
TIoucT3ac4I0HJ4kveEGagfkHqMbN7TVRvprkcsMABe6D9Nsyfbqobw0vfhd1qLFRBmXdSjy3rCz
Fi9HO5cX4ESRMpKWvFoj78mnpPA7W79+9zqGtJqtdQcB+XHk5o1n31eKPmcjp4ZOSM4NUkqFoTWm
dFk3dCp2bHSUNMBRCzVHT5DNp/Pi3bzHNobBkBkBlXvS6EaarSjBGBlBaA2X6PqOV9HsfIxAULn3
9PTv9AQxURbGg4OKujD13sMzZcDsnrgjfgPQPdqTN90+hwsyvR4jAozMh3v+GBbkRZbQ+NWh4Zwt
OjRk+F/QRAEdAEuN2WpM5400QitDlKqjF5VgdybiDZAqpsse5/YGmOrSoku9dPYqD33cl6kbPQD1
eR5X8RpAkYG7uGyzW4RBfX1ZYJhplNwhq4SxClUsoTaTiqKCqhxs2VIEsW4NlayNswaNoXeJxi0J
gosETaYnbRRau+J9laKcEcRUST0oejqjOdlnHGbCpKAU69gYMR1x/0m4b/DqiNqG1XQWPNjGDU43
8ea2/XnVgap4Ghp+SQAyxei0uIfPLzQW8LFJ395K/T9QD+LwbMZIJ2F3sNkizR9Hd0kINmXGLKWW
tcPxpu359h0ksCf7zIvD9SMyxO80f5FrnXvFmZxwli+omo1drluqYiaXUxTf4wfxZRpCGeg7vvz3
KPqEdLuM8Y+ORgDh4dOvEH4lGlz7AoDUO3E7+0bmdwrP9+7S293meLN6pMHOw8WmBFcjPtcXr2Vb
Ri8Vz2U4gxsW7b1zWSPoBwc/K2aCMSwb+EboHuCL9ViV/Ozhii0np3fBMMR3SjKKxlfng54c8zn1
wjPa1Gml/BiqWtmImZsIAzsQnIpmj/W1Ww32vy2y17xTUuFA9KPWXYplv7LibjeUHeWkE7UUh63y
Fqflg7Hc66HNb6fRzyCIBzdTsIijEDOKt1NxsFytGENyk70kS93rF/mST+5HWj+xAusC/Y0uYTLV
6Fp9WJPKOmvr5RGWhePedPMBGS480QY1uKlcumF3AWl1ALyttXvLYM6SI8Dod5SdiDdY2vdGtnaN
RvgpWJE0zundS0mcoh30QWslXV4qP+kKNnDmPSjJcj7G/QxhyLI4rrV4jHcL6MXbp9xEimHh/4GN
tJksAU81/1Y3BmXO6E3tyaLldAs+qo2/cQ156phVsHQWlc7watUlLvytM/AfoxxhAk+NepkfaGUb
PORJFTgOQ8tV/tYcB8S5E2OBh8N3D+HGNI7HgAHPbWQiqlszlSZKfFXeFxVmzNnDLo+iPBFWIRaw
1H0O2QHvcmfkoGrEyWuAedrcY3PkkG+kYcNFGewc2UKtqj9CQ9PA377LVALqt+DGzq91tuyS320u
utNt0thl4/0IK7mxq0vSBZN/852u/hIbM5kVC9CDN1tJFzmVFATW3CRvyz+z3iZyamqvqJGpvWWc
ntfduxtvwCAts+dFmP0dBJPqIMkWiiFwP5jJRHELXVYT1AJjJNCZM/s3I/S75tYySLAiEfiH6Rh7
upHoHDIaG4LnmjVnU9ATsDpQE4QCqUH2LXHfLDqbqyflW7Ac/TAsd2ojhOBt4ys/O5xYmQ4hE8Ch
QzZ3fj5XQwkcqJrQeUYIZEKv5gOuPdnvPpHn0/l3GRqC5qlkW1RkK4tZO7hONCJ3/IgFi2EijRPr
21Vkt5Ah9EfeGFRQPEMslb4nQFplSVMbekBpQMHXH3Uwjbaz9yS0+T3TyEgd3pcJJgipj094c4YC
5HgyBTNirQX4ptD3KJVgA3/+t0eIOyLpNYvE0/PYy6WYW/2uSu28qeNlgbM15wQYXLhhEZSYmXWw
/oU+42w0By+DeuykdH0VNc71Zo68y2PzrNp5FRadpxaeVGmiKjqb+Fxz6kRZvQViDIqKgA5rFxUw
WWlbRxqvpcj3zLdIMiMuVVjzuJCDie5TbW/W/Aph16nrzKJ8ccBWXtgCfosB8Io83xj2uoD+DQBt
HxOpizNbgCXA8BUzRO3B7T0QA9L7lQB2Lka+CEtWJ+Se9VgKPsEebMrQGETkSiMIPuWj5AtqlAkX
s8s3FF0fWxEIhGgN3rRjO6fK1rniz3xkPq8mj6AHdY4l407s9cF3eNAvVhMdZN33oy5MGhFli8D3
pfyQqA8B1Jl0NsnbhtOPsz3+zbPUWKKoVH3oBGL+wSCNno/z9q1wAsfg/mucerC9ArRIQo3fHAzx
Qlg9JhRmkjaQrEHTG5gdED4o6W2w3tXyAk+RhXhFnBCBvqln8nWfzJScgipey+kfdVJjHdtGmo46
ojRzVpJ6eTfhnpXVDBoEmuCR3b4YKfXPCdnTFhHwyAfsHIUKVHBiTKQlAaC2z4oAtDtqsVsc8aQR
lcS2vCXlnGsDgkXZp6PBE3mfyYwBr9H2hcoCNfAf26K/vRhRJqPGljba2q7D6jSbG5K0hIwnwx/c
QOOSWVSOoWCjPlzR1zH2hsvnzQ1xpMb6cLggjP2OK/nDBJSHM4boNhbf+aJMwwe5dny5fwsc43El
8/E7V5le61VLruz9hmW2ofsxYbs181t4CDk/g1GdLXwHRkTTMBKZvUVtHBeYNlp+bV4fpXH7Wumi
1YG93SqME09ynMdvcdGznH0K+D8eglxH9RY4Ea0xBK1LlWgEk/kqkPhxVTcxgozSEmJQZhPEM8FB
X1qbiBsygURL6vBfiWpUfbf2SnsAbeFdhpxE677CplLNEZLOAPvykGiCOZA/jz05Y99Wu/OENhci
4NwqAUQyMW/iaGrAmGe+x/mO4OaUKUqfgHfB4NjZ1XdtNFVGhAC7sw4+IIyp/Afa3HKLbmQypUuC
F/79PI2ZESnmnW1Sk/ccJKBb6zvRpqm3LQUEyXub/ONK9JisS+a5R5R5r1R0DYyK+BP132VDgOvL
RUSNejeYe2BrZMtNzBx1fBaXIogWk8HE5TwViLDKgFjSXzja5gfHeKCqbeeFC5B18mCLV2wlah+j
PmFQy8EHa0jX141rYRu3hc8wr56nXXOWBMaBk0dNdsjlVHwuuB5EFzJ6CRNCoAdtr1mn5jGZ/HQQ
stpwmdulJ7uyy5YVJ/4ehCJNJLEnUZTBsNeGHR5FGb8f3/O9HC3fvZFrNVNUYJxFLUVOV0Wt9p6t
VUtfpI3BepxoZztSJqmsJX2KuxS5NEogTiNiXfk7PxY3QgRkI34pKysfj6M27KJovr2IQ71P2x1j
V70EM0brOkDHDe0rO2Iy6C9iXhQuu9kNN22kiUWaqlc8i0Up4Ap5EGJl/FBOPzIg4o72THXF6p1u
YNy8hcject0hIGc/gchJLEZr5HKVCuXw5572jxC6Ft36Glb6J/Gqg6YphDTP7Z4TxGeTmLGaK26u
KUGtZVfYOjzv8Ht5P7lU1ulVUz6xgK+6aGs4SX78UF+nFY38n/Crt05BOlf1KNYw9X8V/o8OEzuz
4FF7ofvfDC/tHWkV3HVugl3VOvcM1qOzc6A/7Ec75JHKbfmjMNCtWunKv1ZlitsBYBPyW2IkaiHA
dmZfk6A0PwCkVtsYcpRFjMUvMBwflcMQEe0CXu3pd0OoNftLvXQ8WRJXexy4RAXmE4CZJTemRuRp
L766uf9+VxHq8KpG5qAXOpMzm1TbggEAWXBiJecQ1It6kwjU5WG4TLg7OH+jgB7qvw7OHhOefjlP
W9LPsYm8xLT8C+b0RhiSXDeimyoPwUcyHLWbdhejuKXp/7G1oYEobZA2VUmfs/VAvesxcDxferU+
994ivuPHqmWdYrJmawl1ga4VXOre12O+dQPAAEe3nfmaSJ7E5dn9U5wXcucoyjcBuWWLkvd2JqXv
MxXFgRqediFFVV9R6GboUmmw9y8DMtkh+HiiMMRJxVmfCELInv5jSXm5HmJUCLL4wDKn0nA2mQd6
Z5h188t23b6tHUvPTDk4SXYIqbQwGIjxqE9IDnYGW1wTNET2h85Eur2oV0Gvx8PZy5+fGM0dv54Y
unJ5peFYUAYiGrrK9se7Hd5/fKH05Nc1+tQzZnPLfSmEsJdtRZoLAK//GpuFNChyOH1iK4RXN4sM
z73w+wX2fqYQryiz82DhvWw8qIrl+glLYc8fiU6eeFY8bKWi8jRb0eTEOqHQxeiVCbI16MeGD0xc
R2+ZOzNcj5rw4JxYXax00/jotOnExsVDlcOkonXhGMEbR5ZoRo42Xxmn7riJQZHAX5SRRCgR2lkt
gfNCboU3IHQ8+OXyr5sTuWdABkXAWwW2KTs5syw5prKC9vI6G9afiUNzP18cbOC+PFrUKYwvJplE
5OXdC+O0W5eYvZJQU+5fwNbKcA4FR28GgXFvS3EvjtecUvne4oRrqm/JxCl6bnbcW2EGmEMnrsqk
fojzE9kzY4VFf58+8ONmDA+In8DoqPPSK433uikiv0UDgolu678YI7fXXAuZleUB5oPmOx55VxUK
bvg9ZpPhyqupTqTdKc1+c0ePIZTMvzfmGwX5Nn6bQE+xG8zjiL6OSEOuk3uFKT3sh5O9gk16zJJ0
i5DbvW2Z6j8blqYwq0oJ+NPPSNgpYp6KAy8H9j63i71gYt8Qo4mmjUjaq5/gPEeGWUImIr/8jHdx
BZYsU8JJYWZ3J/3EbW9jTvB5TJ8nSNx5wtj7DyHfe60sh3bH8B8OU1Jm2G1AvusPJLO4pUxLlaBB
SCHaGaGN12XzgNBHN5k22i/J8m5wdW4HAdP+oWFKkhiir6H8kImk7TNEiKqfJ9PRoNQvSr6FiBcT
m10HLD/6ZnVv/W29C2nGm723eFaZOwztwZHcPP8rZlpvF1Va5M51I9JI2hKLa2uM4qAYJHtix6Ff
ZzwueiESVztS6qcOZbrSN7jvwWmxchsNhCwIjwnU3zuqNpa6D4F3KpGLW0vi1jzLzNi5cOIz+DTm
KF2EQguNKcbSpmHQajMeWkCY41SM/KThODjkaHLusazVITMOJAIv7b+9AGXJlS9dZ9YHIHKluFGF
vU6peKKEvph7sBhIylm2oZ+KYjDhpksGFRCkPM2PL0xDi8mdzD+jU+uELCTaCI5UUnNHaSpvOVcF
uTvKoXWNx2WzK3o46PL9OmJhjiAVhK4/vs0p27HL1iOyJeQ1wFMfEIGPt36TlsUx7rOK17s5JnDx
e7x6jKUPBMAOBMCOzeWevqVV7Bc3NfaZMbYPPapY3M2aPRLvRw3IQOQL+NIO8hKTCSyAeFcWwbHl
jR8ajmIRxLd+aus7J2j8SeiqCmV6hdsNBzCP1zsxglTeqfKUMYANwH/J8oQCl+4zXJO81X7/U0fb
FDWjm3/Pk+WpoihIhpEoTKhIm7zgoMIexGUKSrokKzrB/5iwToq0n2G4sVZZtxRymeax8wuiD08b
RJkdL3uJ00bBiTtrTmIrms6YRzjO2v52ndH/0dW4zx+lAL5l2sF7nYzYLyuTUNuG1Cy7XU2fRsBE
21bAPM+9E+LaARCiuv/HOvmDZX9tL0QBFa/KTpAmC549lunDdFp9VbfmHxWEOc/8+FhvZrT8lZa1
qUiwt3sUPsO03UjlnvzjTlQ6X9OP0u3rx/rR1BZG8TfmOLH0s2tqMOYlKkaoDa4GPIhJhsTjf3nj
+6av1jB8pTRKHlU+alw9Opn2Gkm6ZTuJ//KNjh1yJceHxMa4dTj/2syFFxvwZpJd+tshDp3AXhM4
nYUAIecybO+QbDgsErtMXVihUCZ0DnbjzfMa7LivzMMwuaqssnSPkTJLrZqxFxNTcTphWIcqCPKs
Y36l8SBOugTvpryDmfidMgD23/FykLuMRcjTcXf1z5rMx5tpWsn9LVgaWBRejeutaO0BpYcR+Enp
Uoog5AswOuNK2vUXBfpfZzUan5m4cJ/y3HI8xFz3KhBqiy8rXYHkrDfwDexVW/Ti6tHU+FGwh+xe
qoX4CvjwlIj+Ao7cFtyQaBL+sq4WO8n+AGq25ere5ekk7y/oDGUP53fgojxyCv70l85to8DvTify
ettYrdZha0uTNNkE5baHCusz7PvPZM0an5E+vjjv9UJkaOzTf0Av+4kSXkwwsWm8+PcXnTaPbk1C
qgJfB6G65dK+XhTC/jvVtKGpcjIhyx2uVkjfM4FvAdxbqknEcTZAqn5naCCjPovinKJTi9ecD9yS
Tj8nM3anjwBkgB6Z5l6x3myUOSaqBvFEA2LMblBbzIFskwFMBhYSzGvS68L+Ar0ippod8QGtpNRB
2XN5fGtwrwKSmnKG60jT0ZjjTXSnYUkcMjQMGBr5qA7cuPejP9qWbYJdIGipia9V1+dh54FzsU9K
5GcL0UDrD2Gis9VoFFCIk9e8Cl95zrZlzCImWadW3pL81glgi2BUeYHLh8Ap7BLPkY+b0hnws8QY
V36OGShpRVKXwe/azJ4VGwgcCStGVXyiw4zZ7ElvFYmmEKNexZMwLHQC6O1YGH6Ld0O2vEaK046B
DI607n9nmUiSyDnix9aBXWXGAaykvyxx8GHhAhkeFCVMMqwgdLafCnbs92Z7mPjg1AVIO4p2glx6
J2dTQcJMs4/e2iK7iaPV3YyHFEyohGh/Wh/VyhdKWm6DR8Pcgbt96GVUVWMpOisvGRihHkUd4sZz
Y9tW7i6FIiY57IvRNnhd1P8wg054cIJE60/uz1WAkncH1XBFY4B40TmsAbiaF1Xnu8rolI6m5Ahq
x8Y+576l43Q4b54OTt/Wil+Rqskuf5rPFKiIXKJcWa6Or4EJPigSzAOk9EXjl1c1WTmZLOkGClM4
HSoPcrqc4ta1itL0dpnwTjEqgKxPwZLOGeTbEzsSb53QLWp8UbYEVMKHnJ/rM3v8KvsrYRUdvsCO
Jslhnn9eyee1JHc2K3eaRfDv+a0tt607L22X8V1xPlV1LrbgkaGJ8xsWEIo68XcBbibd/lNahwH2
F8pM/Y99ZVgz4qTEI1NafHtEOliwE66gtCsL2U8p9UTXiQrQY3zs1Z3HwiCDN2KzoR1S3uBbAJXf
ps6kegQBLuy7mLClAPsorBItwyPACW6dvWnV+SJo1Ql66PcJKEvCytgaSZhcInXAAhnEnVGK92Ua
8+E2ilyJROl2rGTzNmyJKDXob6xa00cqZFnZzTpljL8v5Lot3Xeigw4QCd3pnvRAd2q6g+VGyvNg
v1v4/0P2DciBWoKfoZPxZL1FmzmRiRfGsXJth2hLI8Zyea8D1nQB9RlDOA6tWBrzuflhgug/LOsA
jhC21dVCNAzHg5K1EKLVkn9vhCbju/DP4UVx4MY7hG64uurvBeH0dpndgOqMuhWyg6hRT/WGN0t0
02k3m0VeQksZM45OKbiwpDW8/zNadr28YaW6021Ba+0X8xc/rJb1/ZsBlTGOxDRgCb1WAswXHK8V
KuRdWIHOTdMFUe5DN4vODTrRTbeyGDyh57jebPCR6uis7U/ORPu9UAtJxnGE7yZBegH3GmGyTabL
Ai5qz5sAZsrzM47685Yo7IocbGzTA4GeuUQN4rxhrnJFcVKL2H3uD+EVASq+5QfJt+DCjDnYuK5V
yH87S/OPsC07DyLNEP5yIRD+68KQeZuLvRMUQl+Yt18HZaj8fz3jvNW1MCT8OxXByJ/HHX/SQ+hK
/FcD5hHPYfuJyQzSN/YSkgZdpBZZ9PftBpevBjGB6H8TGIy9k4P+WRRbgBNYMtOCej73awszgpDl
8Q/EnZufNE74vomXeRdHOmK7MMI5qtt97jAdwjezPtJ22GnqGgdS09esLUHqLHhVlBJBpYkFhLJD
mFB8do9oA+ikIZ7p8ME7jvXQP7YmMBo8VOp1EyOv+y3UVx7eFDc/JSeZHuiEP6E+V01/SH17hc+L
jRnH0vckk3+Iw/Y6GqHO4/rO2iAgtNbeHyrba/htVNkUs0o8hNQFgG/QIWKaHL+SjPXo3I09XUMI
cF2/gpIz3kZ2RGgMX5oSaoX28ivOXUPiiP/hQflEqfrStyXfXwLw5lsK6Zs1Fv/+NEVGlQk3HxI6
MgolU9x0lnJg2mOgBU2S7QmuOyT6gtHfOPh43qkQrfr7JhiYplXcutWPeDwezMmIo2sjf+o1w0eM
PaJo79iJZ+VP9OhSUeMcgDCwNqCUJTh0Ed8v8g7Fe3ENEdlntCkqQ4kof4Uruqzcl+7NrZh4livW
+zKxGb88Ko6l6lnhATYLlE3KS1ydufa7OnaOJQBAeSnYyxPpUzGkPjex0byKRDNvRNSdm91q9iGt
S3XTvjZKtFFU/bMCVyTG0SZdCyPxHOBfCgeCmLfFevn1j28AUAPKdnhQjU0qfawguTirgJfVicyA
bCW+NB6qyHhHycxKYajkztSn7r396Qr4E9QNDxQcVhcYpzqf5PpIBh/gtcZjS8LRofDWT1TdmR3P
xFfK6SRg2ADMqcn9rvWofsoq1LA2ZH6egArUh4yAoICsDDfLxJen1drWG3TVd6Vs7JAr7GhOUDwT
bMgt07ksg83KK9SJQrke4X6/WXKbgZazodCNRfvRLY5x3XLRff7z0EmKhq8zJZecZ94hEi4ozFFq
eo7OWM1wkN4NdC+kSuQEFpxwG3iEGGCHAp6dRg6TeBGkrCP+8ONtinZI9t3o7bnXMib11JaV2+Yr
pIxhAJSWCFU+OdCR9otGY3rGkSfD63ueWnf74zfANPoWVX+OUSQv7clvUQDAFPfQUkl+DWOL7EIM
gr4gb5F7QVH7wdUSJ1gR9R0i3NEM2aoRs/dfGOy0tDOhL1BcUBpIfsod0d42+W178B6RvEnoWUat
ba63I0Ku+toN7gvmCtDoAouBRDHM+A/dZpYzE7ZppikxzvUwQGffT0o6om7pgUY4H4SyPbbzgn+S
VQ+QbzPaPtLYuE65LRevlnLdt0oCUbgGK/9Ap6wUuYIlF5qpbJil5J3AAyO5RZ30RphY8VbOBTdD
fuOb6bOBohjwn11hKvoPhHG1TxRDvHmekH7W29ZUyxRpvJSWrFCiPULb+sRDRBqB83sG8Hsrh2DL
NOnkow69B0+hImCUwqSNirLmGrOhS9nHc+Fnrk8rZ+vg3RQh65aUtMThFzaWg/fwhRPfi02EfyP3
AaxScW2cE8odNnoqXSLYzfPAMNlNt06wA518oZofI8cU12SKQvchJZGNhDdrMaVPN7thAXZ8sVjp
ON/1ZviuifnHBUvN0GTj7AxiPk7tl0v8Y+D4zWnFG3HgPgxmdM3X+qGzkcvp0pJNFgLQOL7mWfhA
KNuXSKAiwEAR0/8R3GSX35e0ejc4+wokV1QT2B19B2U9bTnr9Zyb4/0UZxKEz8CSapk1PhPI1tmd
233cOB0RNIM6hzVobzTrxBn6dVr+UeoWY04l0G6Us5WuXq4ahyI6QKMmx4KrJOkQDZCDX3dfsdJD
lUPg5ZXa2z0BSbaMoYjj7w+06AE/cPBTInYAwwv1haNxTwIpS6SIUbaQdtnphq/3nCJC5Pwrg48R
UI1KqKgJuM3GM+6a+ukdUU5xE12j8mOlfUcW5182x89dHA48lZhVQMPLtlElgTBR/6kkQpYq/WTy
HahHVSKq4naPYAK7NUF0iqm1oo4ntLwkzf+jCJE/DxtWjpASmcuVNtU0ljlp2QdBzoRBg3Wmsw0h
jj8Cj6WAZE41Ny3YJ8NDjF9maoiIlPOkJgw0LzYn7vb3RT2/ALYwAHGXuI0u2aX4tAzvjvJLuAdz
QLUG/a7JBZNMi6bGYo1fstGaKVvVc99gavlz0jVSxOYUBqZfDsfH9iEoTVM09IljJQifL6chjVO8
IG/aFxs+Xl0De5flEKsR2o5KCejIlLfX+74Cu5SrLB+qpdWjkK6mvQpN2cq/OzninBKtGfYbbQCf
/LUDyJn4ui8O1YBgUlaNcqAni+gFCdJ/qJIS+slWxm2xJh16LJVZeHhBGmAdVFZ+zBDISi3OTePo
5wnOuc1B2e1NGA/FNDx/PEULh09XgsF8I9PFSX8YGrm16zSTNYzJmKB7lbH0RbTuPLRQCJVh4K3U
WD+P8bdvb88cmhy/DZlSK0O3VkNR3tMQkBEX1varuA3DGfZyTSHyMb0oX8lAobiHKjfBFbnop4pl
dy5/NJu9ZeHPzoWriWzThSpxl0wyOm1cqJzfb+mhoOXMDByZi9B5J1u5gNquIXWCNW8OZUEqWbof
PmoUYHLTfAsjPyfs5SOKcErm2bFhQg3K9b6LIPUm4pDK1UaKj0YBha1BwvlbFuq4WR6znKuT68sI
bVLZNnPO8kqj+vqAZhLwDuy3W1V6cQjAbJeRh7LUo81GmPA36ajYUU701tKNf/JvMsCYWlnVsguP
lxIWYfsYRBfFR1pXYzK0nhfZrIcleSN/lhmwsxffBdlHgBhlh6kPGmy2+Fe0vypUTTsOHz+eCrwn
lz7gTXHE8QqqxsMaz9j0xMYPuNQf9zTI8dM1slLMknC6XBTHsZ+Z0NaI224epwmvBhEJcMClykSt
PHTgnowcErG+qjJ2YGy6qv9en+okFBlr/858D9ZnYxOHPVc7cUUvvdOtRNRaNBhdpOSszhBO6oZR
3EjvCdTReyguBbFU0NEjp9FqnnYZB18Un93FV7cnQjnaMwFJlOWmQfLGTLyjjGXBGZoUcYaL+3pB
nO4O26YGR/Kl7cUiwHweGnL1uHJShcuU4MLi9S1WFHKMTTqPlvDb0Ke9LKJjmC/sBDYSVUAAIRkv
qdhbIz3lw38mbm0SOB+XbREn4XmuaZ4ZNicVRzZmKpFES3S4dpEUqHHE52AHQM9xaheP5/HYYyU1
Kuf6olhvT9qmOfsQmHFrJQyss81/d1QRknw/KZoXq+687HIIvLx09LaJtuBmrZfihmv38fjAJ2Kb
HzbQCH3OKAXDZrCzgsGzyAgasUEqf+ndN2iEHEqKuUdmnjY/+uq4Aas6fCRNUknaZOmQ+QEPRD6+
KAKp/PwKcoZIr9uOPjRoMAFtLXzv+NjZNFDO3uk7yGhsGU4VpKwPIoiBcyPHrauE93laoMB63bY9
umsMPUEAB3vG0MJXqbNdFV3v1oKLUFBkje6azcKU5yJ8sqNCUbo+Pkpn/4uGZZVkEGwFjK3BOVJj
4LHEC72d0cY6/T0/aeoot2V2LujuI1hHl0Ku0+r4uKySHTk7xPV0QaBrQnfU8b9rz9iWQjps/5ZF
8aZ/JSI/aXF7BhRMB57ln5SX7vlIZQKQDJ0Dm5pp5XpD+wHCEsYnwRqesc6EHcz8F9CqmHRPLhyu
xA6wS8SelVU/87Pin220qzHcXknNPmWMSuTmdgKX546lFAC0pFvkahzfQceliRP7fKCwXyrAnTHE
nlN0RQPiCLBI26Vh3usF7AdQtV6OSvf61xjYObE8oUspJUvmrMkl8vYVhkKUVNnTDS6zHRBs6xW2
7Y62tS77rT2s6A9t0D8J70JwgB5CRMYbeefX3P9/qY9jaAji0Xle+gk4aJYYTfE1eJupWM/ytYs7
gDZJFVsnwpQg7epZQP/t9WjGbRnSj0A+MFzbucfuK/heJiV8+DWNhAOvOvOsZxmf2AZqs1OW+YAV
mLrsPJa+noaEzwO8WV0VGs7FqOp0liaGeiwZ9GyUWO1VcL7JIwUAvN5DXAIQoLbMc/lnWeyTWvyh
Lbpp6c7Yx44qFEtobPFdQSmUpWo0wEqcseiEpc1Mhwr/UFiQTUESqa1+EyuiY5SPRqN9Czw56asb
e9gqPB/DBqTG8/A5agmLRs8UqzXZiXvGo7l1bN3q+fGkur2ZBP6FBEGnaGCc2dTrEWalZyQJT3zR
ds/OhxujQZhnztSA8lBD6sU4FVLMUoponOjv3ikGd6XD7OXbJyujU0d+uWXRozQmfC5NE0tLag9Z
qFu6UOln4ABJEnRT2MuGAwM4UlyAsE5MMUkHCqxOj3ZLoy/PAgAX1bB5ithXQZpgWxu2Vbn/1R05
bs7Pk73R1vnvrhadTi/tzbtRKah5Xmg/mB/bK/7IArqc5PPLSht+1bL41lfE+JdjeuVAWLIMQuT2
+sL4QGr1RNZjnIXfrrUlSJtJevKpfV/bC93+YHNogmAjoJ14rgRXuExUqluWKE6+9+0URmXZY5r6
atJCslhIWpVSywzksT/eSW2xqzKHKC87NrWPDgJDgL+5XQXmfTwp+19aNlYURt+jsb22I5S+hdgy
wdhtQyVkuX/kbZ3Fk9Y6s5C70ywQTJBreTxbZbfNRw33sUSwcknWqGja348qubVC1RI7L0L2znX9
ON+IzB/zUhV3FtcbM00fROgWtBVioayuSh2CESnvgi4SVoM/Sk14eEmM8++GqAJnqmV5jXLxAJQN
FWS6ctLRE6VraHcwfp3GnPmzdNuiynoaA9bX/Xn1cD/scfJOZuOXPjDZtZDIaMqgiQN/PB6TqECZ
aQ63qmSD0sKDvbxc9g9NqP8dftArbUDbyBrvVs4uT4xjUBks/a2eyOg9Gy7CxQAqxnJI1K1qeEQn
cIQf6ebqyhPKlYD9r76adrIwheW6TwB9xO6ywge7sC+qOtcQx6AlIucWf2tHNne9VQbTelUa7jHU
e2++kqg5WnMADqbqEa92TNZxSshTSOBqfOcUukiyc7BzcshTJhm8smz5Y6FVQ2OSXO588GA1C5oX
DjQ7aYVOZMcmpDyxzTaPqt7H+rf3HtYmR15tgJGFV+RGttfEBuhDDNIPzCtBaUByd6TnRGzKeP5K
IafaPimOeM5Be1eR3zQTkxh4NIt85k3I9TM6GuaXSKevo2zJetG/SS4BRs+mVLAZXezccne2MDwG
5RRw/IAXaNMUbq4kQrx1HYz9cMAsKH+hTxVl2H8aIFgwK8G1BUVtcdR8WrEBNxHjpR4vM/IZ/g38
Fu+tI09b8+ULu4aGesej+veUgAk0SdkDzhWFQOKGyfWl7vkIJIRpg+tMhaSTQDmhhesnFNVei5Lw
0AFYQuSsMRfxePfd71IXTXNm17VyZynSWX24CfyflnQGsrHiJhGUDNDrF/bDGl6QJ+vyXsxJpkOr
RRBM5fZj9Kl2pWeegyUsaqSeAf+VD/tT+LO7GlbB4ZMKXPxPhS6ZXhlfVs00YZJfQdIFFvADT0Gm
ow/JtWtEQyAMHoJ9bpcGivGYIbKXacpl470GInnrNTh91va1rbdDX/nXypHy/x+8Hal9ddW3FXdW
dG0Ga0IKj4jEsXUq10z1Bvg7kn0iJRxbIgr5Mrt11ofVXy23mMD+rOtAyhUBwaZ1/UBeBgVK61BZ
94qd4SpZtsXAPFQRu/srxoRk5c8jvqR93m/shlPZ62kl0fEPoOykXmmcrQqjxMvHc/uB9OpiU19i
g0wSaMKdW3zV/it69d9NA899ub2sCjeR05gMWVNxrL4zfV/NwS+JVYZ56mO3DTryrKrnzRCE9Ylb
mo+oupkHxlRzY/sKlmnZ1ab20Vb0L8/V7BO/oenslfHPFemhn8qExdpYLhji9kt9qV/gXlsCIgUJ
NRy9RnkL5puIgBRSIDzN63aDcAvKk+1yt4JoVtIzyczFnZl7XSyBJXpbeHgJLEDnQ0vjV3cQSTk2
c09HViP9AtGQJgbiJZBx1GV+4x2iq0YIb3vK7Duh8w3rREx6bXZRHvk2CVS+MhWv3vpoaa7+AhRl
TeuJ7Bmf7IhmERuzHoDFUFGcq/fYjPei2ccKJ9PMpw+rBedqdSikNMofoQpKKyOyjHmOTs+1tU1K
Ewh6t9+ZORFNX24X+90y4fPiHMODI6QQiVZttSyiez2oZSarHtH9KTn0hpt/mDWk3DRDyxxQgEda
jhYDdNoCP82YQIFr7iE2W6WATrP2DKHEE1ynppulXhyl+j+ZWWA6ALGIkQbnNlPKOmmVBpmgIPNQ
6l5ny/O10m75Y1wR1wekHBk/Hic5SZIc/p+BxSBqG2BySO3TGS1Gpeu3xI7z2J9zT4fiTC2ZPtGt
LwdfHY+cNGhA8zh2KYuNsWdOEn/NM7Pf5/KS2vSepLggeedDYF2xNu9kvksnMxVtd8dIAVh7/JyP
rKxIgtZQZmnF2HA3Dixj2AIjdqzQ1dWI3GVR1EOjmpSj9H2PSx0Gft4JwZW815X7x4JHDF59bwpB
bukf2ho04PNQygKsdsZ8CWjo2pm6t4b/1M5iJjBIT5u+7qP3OLVtf11BLnXc1DhMJUaXZztiSxBA
WISjykTKBIWXwSSGwWUOECYfbpy14YhEoNCbm2dVAOnwtxUgP0axaf/RPO0OwwnpsMPmea9s4/Kx
cItOEEqR5gkp+bKTgoX3xIgEa3FJVHCBbVW5rpzlOLJG5D+NuOVYj79+xXI5lxOiOZ5yVfHoHU0c
Hkr60ry38gLrvKcOy+nBoAGwOZdx6e2nGKdISv+B3m3jk1fsIjzMXqB0leNqEGFy14gBhh0JtPCi
5s8kWmh5YhoiQdjx7jvzWeLUqykZFAHYjYn0vzzD9wCfAU4Uo6QnHVO6216qSHekWfQp1QYE+RI4
ApwEYa+KaLM4GBX/r0Vtqku4BNm6F3czH/MCD2BvSheKjamwLLKkLAXfhideyyHYda9H32a5dvuK
IT9AV/L2BNQ6MqgVYFXvtt1D4GrA4KgC4FpQhPwLJV9vMwfaKVIDGvYMYrJsX8uSdNzFUQIo63Yc
g9RlDrKGZmzpMVWjseT0CsuE2xPZ87SWqXGOI9c1VWVNeURUgoNX/OvAWVzQNeRbvZdYXhYbHUh7
+QsxphsMjx4K+XqkFFEgJkkwY4GZzL/OzBBrNMOaBp/IE8LhaBpsDIUcUhP2pSfBCIV7ZB4OrWft
TF37x33t9Z3O4XmkfsNno4F7BUZhDdbUWxzCT8RzFO03jmT24tQpFwcXi8M4sLa8gDi3gbEnttel
oMsPNqYtNI6g13uQqWRcMhKOU+ilW09/T3mceDiSwYEXLkIHOE9MigExVkw7eC5tLVFLI+sjEGhO
hbirevwzwJfxUOqRylq55Nfn4dWEeZrUodYccV6bmxJVsyzSPyvtTMRMgR1TilXDA0z8fKDu2pyz
WDrAjtDmzaO4ilmWuSxglTV67nLtMiP0ArJc7YDFH04Fga28WAD2BJsR78Bo8UvkzOJo2vMZPUR9
xlfeS6EenKgF2Ry37WrTvd4p1UV/5rTdXq/xgiFyt5aiGtdH9Lyi9+r7kSzbiqrX/Dyi7xaqRjue
bAeHdjkX56tE50ILx95wH/WbCFIwghkaMg9wQwfUlmS9UM2WinOj2uJH2XebKkON925GsZveGl6R
jbLSLjxISO3gV2Hf6IPVKj4OekyTd38SWrhMAOYEop7p42KLurSzph6u0gRz8kt1q08LUxGaxyC1
I2Li/slmZrgYDZHiOYG9r1geeTD4VzgxXJ5PddY81fF3fv8M6HselNHs30l5mIwNWASuHsVi13NB
Ww9ycgq/ORWbOUdTIdlg0aQ5ZBV00ULxioDZPd1St2Z06IvRGmE7ExYW7DNt1YCuE23kagYhcd/u
Cs7FdJ9FnVuYe0TtkzwQPVJ7gwY4uVRGZ6MKAKARfrm+/3UuSl6dnM/S11HZf5iKdFX+hDdqqpW9
5HstjAsR7Q0b//i2j2ux9/vEYUspY9pmHL2OdoVoCYejU+Cflx/IoPWLJXN668e8m7sDzts4Shlf
NlXZ1O84IJcF/9YKHeQbpqkygOR+ZefKXcIckTEyN5W+q2ODQxydoWkUkltzRJD+3h1PWuePUfLJ
o4ztaHV5yeiyFiXF1ENgTGviujxtTGnvyck5vfqSOMEfEH9YfZb5MH1f1yWKAoj+35W2XYZ+luHy
twOyGXPqfUAMBr9nO2uTbQwRA1cHfmZ1wWr09318ro5vh+DhckhvFUkB8YWJXAGPnN3bBMWu4ZeM
QMneu78NtCKlNZAPPbIMSrIe95JYzZhTXSw0iCM3WMMtLCnD1dbYcmbaOz2t/cWtIA20GsXfktU6
KZ76wADpQYh0NXobfUqde38H8ncmtUH5PABbuMFcxSbBfki+iCYBoHB7HyBhcypUwghcqMXDisDy
rcbOH0wCnqeN9xI5Fi3I0auBCe1FIrUw17SjT9EL0DAY8IbVyTos9HitF8mXE9s4FYEXxP4ILo6s
phjiZgVK9ykmXqiwtcy2Mv5I3TKpSblHixcsY7j+j6d2noO8KdGsYwkl2TI4WUo05FrwrOV1SyPA
lWFu7jielQymDbkjLw1lBuuABquNEKi4HNevrPItD8x39ei6mlcUttIQBu6OigOyLwZoVl6bUhb6
iX4LRaElTL9nh+9tYTpymjUs7KDS8ft0MSvYND9yzMv8A6P22DeC8cCACI2iFcAjp14+kYWi6qWa
tLww6BmVRMDHMq9PSTD42HLScLxt1h46VGhoj0ZlYW00YfK1Q+3Iflw0rIskamI5pSPfGkLs3huH
I3MorLEsktG6T/KtK2FWTuZ7aHBQxX6umwKVqByFByolq5cyHlV7HWoxQcVf0R9MWcmbvxA7DVgr
QLuX8qRuwp+7+grBD2Pw12qaGXljnNblSNUOW3dWBpsVfmoXp9GBo4TCshJWDLDpelTtNdtwmT8U
Hd6Yzqiq4/iJ7OxhSSvd2t+etHLK7KdxPJ8dLZ3RpvwnhqYPTitlx9PxCLgsEsEMeW+0d0iwBdB5
5CBLova0ZBm91Y2RRVldOk6XnVSCEeMTt03ln8y9yLLfCFKJ+3NTkWqU/2uoX4gBoNjQF5um0fI5
gA6VSGO5f3zWBIkHTVDQdjqp08BzrjGQjSZJdstUk/LKwQpDkR8oiT0UFF2nA4C9UASZQrBfSe6O
AYZ6tnjGVzk923wovI9FMBf1kmM20BDGugyDXOmVRqv17zY6CYHKU4x70wi6Qk1qH/gnD/NWjaiT
hEiDKIF7lLb8Fji6R2p1hAPq+CBwTJL65BQZxwrL+0I8RkQ932nbX3PeRzTlPcU8Z4Jwq8HuOoha
0xlBL80WXzDr5IZ4oG2+mVHf7E+7z6GrHG4uPf+fAYPl0ftNpePviffSINRnBamLrl86w+wxePit
elwyk0UDAaUTbbFp0ChY7twWxcIREhI/6kNO8NwDS8wKPBtgyqMQbRFwIOdsDJbAARvihliGGVuR
wi2RcPbLj4a2twVJpDawtfNynUeBtS4DnT43f2bbFAtsvw8Ea5CATBItZpdX7J3fZtdXsmRFduIE
6IN1FALwd5bKXKGkkBAHpAmHXOcCzcROA7sQqbf5bogO9ovOabsvjvhkF1GOPwnb70mlSF51VCVz
zYqZKfHCPfoSB2ipdycL8T+YY438kDnUN+me38KxssJa6KzxKuYcOV1GmRXR8Odz1a41Qqo/UtE0
uta+EiM5S3Xi0mKdHKjgoplGlXcdxLyrWgMuaKLQyjx9eKgDqZND6UTk2PAnMh/wc1Dx78H+phQv
3V44FDEY6a+OlZ1OTyd2jKJKdp9l34KDAdUs+xuiBLGTJnB8lKvT6FYbPHGrGpTd6aMtpEriY888
3CFhNZT59QnDJmjkNrw0HfbnQ6OnTJGFf/ockrOrz7zfV7RtezyktOiWNIymlxu3NakYmfljeSfU
AXUyHQsLbuddAhBsCbzF7Vre1yKiJmQ/1DKs1rvoA9jcAfw2uhhh972URgoIH9kw9LN+9iGfaddC
zQP3KHfCRBcJ6jOA+h+Dzrw0FZg/LVlYbAgyCHUArt88wF4X2P7n+SjSPKn3Y/vYtUODKmoFK41f
9YI0ofr60a74Zoko8GLY3ggbLopT7RCbEDiCHeow8mdPnJGqIDdsbgnPK6Y8l+QLxBs4xyASepi+
QfhQzPYPYINJ4gzTX+YDpP2B1RyhXX/hXxpS5w68/O+Cp//KyHMV/CSwQCec9wNwaB52ScWdbybV
1ivwPlHXO8UP9Ag6qpm36AyfdFrRJr2uZGASettk0OkPMy4RwmaCpxZJAjOZpuBiGPs13HzcM2Mk
6WJJEarcLJ67yxzosak9EQ4TvebKXyFKj16paoDDTdyndLOabsYRX4/NgT4lise9nS9ImBgch02t
qRN9ibaGrACFfA6QbhaZwQngxrUxISJU0ZdXIaENI2XFMxNZWnPBZIJluCcVpE423ZXjnhVhQcWj
fg1kMsRqWDD0KsQwfQvM23uq6dyfBvnmhL2E+Z8zyrYwRAR1qEGmEDluV3WIQDcfUj43VJiDC+Wy
fq3p7FeCDIhPibX69JT+3xN8v9VugKxQJH487NrijKPWRt2JHl2mko574CpXc+x+s3xfCJYpLlTm
geCSPbL+Ew+TEFhrM9HWmrXSIwate5qhyceRXwhkXsmvcQyre6+gYXWLdDUY0z5hJ+h5pEcSrXRl
zGKZcoehJrffAsJyZ0TQUeNxQEMcmeHzACtV3pYvCu805hnrecNIt65kHvEyZ6zA2GFhbF5AX6M3
4l9ZRRTqXxmkKvrHX/boeCs8iMXp/6L6GfGdCcVFQx4Wd7EQB1JMJ8ihTVeWTkcg5D5mydHHPDWn
hhjU5oE2w5GOt/0zwJ/f1MN+GMTapR7ks2I1fa2nuBSWE4c/qNnPaJ+FDz7jxQiuiT2PtvM6MgCK
e0Kx7Pdb/Of5wEQy+aRq0PZxQjlCHY9SgfGcZaLzIqNT0uqRDlOpfg78k8+79rN8P40NKCgKuqMK
k0xkHV6HspMiBIIeK9hnTz9yhalZBqHo4fMDnvl0yH1MGfbeynyrn6oua/O8U4URke3FiVwtplaP
jDEB8OgAH/Wt4T3kNJU0MSy1hwec0JhTR8yAeg/PoAPEuBzdM15WHO1Op2oYQ5gi/31ONFpDilue
FcltlsWEn1TV29YQH9WcBrvXt4fCI9p+xx/reeRiIIFo7U12eO84UtPd5k8G5daCrCS2/v8CxqOn
2rjEzeRTosWsw+kENPmZtS9P+4w4fEiNx5/sqXcUal2RKbuh8wwexQ0wyru2krHAmP5NwwchNN++
9fVhlbEuIR2RMVesWPhFsa3VsL5QQEwo6ltH+HlDMyCbKEfPGYkpJuODnbF2X7KhMBlyIGvl3K+p
SMiqsqEdtU3TVhod+DsiwcNGH74dhLkaG/Ip58uMQFFYPC+qiv+TN3OOQekFW5+Rfccrm6fevCSc
MrTo53X/FpTWoiMusiYM8WDyXAhn2OvA8AlMzx1EsmWOO5FwdqDHaFYkJ8ZFI/yWxwCAtYPtgvjh
S8DbI5fXA7tQpaZcMfiLmn3kbtD3dDv1IW2hFrGkvUnLSC+xSY6yoIUSYj0UBPoJvhREt4TGRNhc
XgAh9De+N6OK1kaIufgAA2bdnoMkxcGgngbdiWiAyM65izBI0NNsnmvvmKnORrzoOaWo7g1VhMSI
aqCZXNP0sEWkQfFU563435kiAImoufZQ3G2PYD7BfOeYQAH8gsw96CkGQZaiHyit/yfn1Q2ZMl9t
QG900EVJsG5B+x3sv+f9wwBD+Y6Js1Z4nvwE6qIV7cDhBiq4NRC2wsL77Oh0q6HAWnWWW6ErbG5Q
jN7zEbfOidAP48hVdH8Zx2XAUVTD2UEFo/yWigZnkkdAAfB5dm8ZwzgWN4uoFK5GaHyHm1iDk/wW
YDQ2MNXnLWwH7vFsU7aLa2zorCouZiZp45CB9+bY38tmwtJUy3McVQiPhDBs5zNv7bjoE9n8fubz
h5si3J49C9JQk9WcgLtHuDCvRmDMwEpTS4jklHiaE6DSveBc297OrC5/WrQe7IGYk4uGFEhgQ8nN
TaYg/usO5xF9pttO+PUyPQPVjz+3ewy8kmidpuvwd5CjZm7h1tfognS9ETT+fFNe1q7q8pfX3jf7
MAabehMCrgDRREDL8knLGWrbJPW1th7sSimInZeHQ5hWTjRe0ZHu6o96tEFJIVDyiu6DC0HDwmQj
yURve8eeeF/aLJ2kkrA7m2Yv20Biz/k42lRNxMEat7Fambb2GrNr0aL34lQPFV4WSUrvf0nh/oR5
8sDfN57SHW/lE5cFgGUZFl3SIAOBv4BWiciJJg5bo1CAkqhzQpwajlmkTaBkLoQgNRo3WdgghSWy
WUibprHc6OcMFmGkTUcTkb/WF2SplgSHcqeu4nS0VB03BYLNAzcHlq+AqIlOJV27xzp/9KGZhjOC
Lblgi3+SbbMYjlgNYWt5vbomC6UkZIddqj/KMkWnvBOGrJzbxSIfSx4WO85jhdSFW94lQLKvrpFG
T44fOzLDJ2RyQkOV0R1kUpWf4/qRIgIlVP2BuSwOxw2LwbE6SK6dK/v5Rnk4XCMTtHA3TeJ2h4+Y
HjP5ICBKIW5s7OktJIK5njmiIZUhMdqLp4D9Qa72tDaomVJcsrFDOUAXIWG1jewrIaEYN5GIx9ab
tzf2mlE0pm9JjRCaI8NijJR4emj8oaiBX8PuWOfsIAEJn34gtJ7F92r2NeY3yORU6t/KrssESLyN
+XAAPnAF6L8jZnlahrVdRcQn32moFVBaDM6W6VkkdxY+Zani9FcRLUlH8S+VOSMoa9dT4NLDl6EH
ASHOToi04lZQFKpCwc9nVU/BY5b0tOXwVu/d0/abPiHQ98X4e5Lw+wMMG1KHAsmzVuBCs9ATKEqF
SOdQcwKoanhChI7xoe1vSKpH7j8it+ykV/NMPteJ1thu9h88R26zXWy00y4dFNGxAv2IsGBRqhjw
BhK0M08MbhqhIoW1nmsaX+Tls8j4YwSi50Fiv6+CRSX7vmojCW7HO+IMmiXKnMeNIi3UkQikz/Uh
nlLOEMSpl6wXoXKfabAysAClemc76RUEgrgjYpvwphox+h6yLiewein4MiTPNmTkgOuH88vttffg
+aFuVmW/NGjb1nkpuiREEU6m8hC5dDKf+Uh1GdXfO1GaxzRWfeznVBo/Qvo4gCfSJk8Zl/InIToy
ctf9N1Q6eEDHAUOAyMeUkYUZQBisXSpByzl2RyxqzYDwJD/yRczSDzTYl5XvRW9A4eWVdwvJTdia
QmlfteeDFuC3EKHTOug2P8xbRI4qhFP8sb92bWN5V/oL8/LEZnAclNlUaeJ5jZYmvSWQsJtC83Vp
x06VC5/3x63rsqLK/HEsnsjsVIYykHkKeCNIFd6UlKZoEMCfaRVXwvIq9kByO2u5K16Q60uRiyuj
2qk1ZP+zmo1vga/HShc5lQEUSdKvYdj3Z1R7yvChs2aRyAauoeODdOl8Kkvh+eKaLXm3WeaAeIER
VmrEQn4x/AEmrASG8/T4kRb2m9ggB8wJ8ml8bAV/XaliDQy0AfiMUzc7n0i2h6RVhavwMBixIIXe
Wr10nSQXC3Fh7pnU7ZpgLOcCV3SlLoVFfTbMqx0DEx+q+dZSjqz7OocTWb1BMiS3L6HnDHGRbwtn
Idai0E4r2gn5jQyRRi0wcBNtPYJS7Bas5lQ9S5rbzM4cYxIJkJ64zo3vbLS60YWGQbhHftDDmyeQ
jyf0t8MZXN/M2eGIXRWnHitPFUXh8ECx7kx8rdyp8z/eT2MG9SearfN6hQ1HDP3C8Ssi0ToT0f5g
NPicvSaC562rfV/VgKhc2AGUTrn17dYzGGxQqdgNjMPRSe3p8qf88gqYwzXREhgWMq5lBmks54aZ
q0dZL2/J8YGxNq0Drxj5nYz+0Ud//5RZqn0OaNQIJenX/B5EWYB4dW0AnZo1wXWMzogBkRN4x7c9
/JEC2mQumSUl6bRavhl8UrnvyA8F7ht0dtUhwcZRrrJ/lzpvNK3CMBAt6PHrWTwzl1c1Usa0NF9R
0ycf9mHVIWJCAfjHmCpceLWFBSLJIYx8EWnILIRGsqM34HVrVvoGraSXEAN6oBbtvpz6Ps6cHM6H
vmlsFf+nfkJtQaFy9AGouWwMtYzvvFtSw86ZnEogy3MedfePza9PNqa+bGoOtguxrLHKtmbsGn0W
b3Tu4ydTJaDb+Ty+TJ4IN6c8IsnCKWAQ7DYecEzs/Pm5zttJjCwAfpWi1355Oxjg7gptDLPu7EBu
cAtE1GnnTK+Zhso5zYXGLZGNd7Xm+3E2hKHPmYZnjhUlBoyP8+7OqyET/cQfJQQfM8UZLrbXLgHO
KM5D64oZ6Q1eu1B7Ab2W3qoMcXRAuurYsNAYj4tqQAg99FVzol8Wb7KcLn8GKhdJVZ7RshFVT6Ah
2u2PJsrSt8uPgVoIviwqdDKXyXoTD+lSC1jIQVVJqMWbBHO6ZlkY94mPTw7TPSwEwjKaQuC042j1
fgSO0qJzwSjwWnwtDq386qlgXjPp+nOkOlNVxAUoAvG4RSV1B6OMXHK9MH/H5GHjoMh218XOBe/Z
2ibxfO69hYk50v+gN5npu2mFXzUet/ZFvNcPN8wChxqmSgFo1C5Gl8srXu4AII4cpV9QUd+dHwKb
zYEJxTtaii3hFoQz8bc2/pduZbe0qVuRgXfRtDSjw3r0/jsVdOBLt1UIrlaLunVcWPkLQeSL9Oqp
+RKPjfE3dfhLqkLTfUwgm8jCOXCCeQqSpYgE/b8NkSgpD8J0bCzPkGABdPSIe2DPp0YIYTMd0FlK
gHeWNpK+Jk1inoPbRM7mGULINnpS8ID8MGrCb/aBGbEawKcBydb6QQn7Nb2GNZmqAxhQAVVXSxL7
1/R8PSCGh6Hc8/7sUaao6al01VTuM5VuQofO64d+Df4JkwVUfi/1bCDYF8CL5vNHZLiI0UmNNAPT
EBLY/X7baoxu+StIV08M8zjOqFIyo7eUehmrQC5layQ4zn9KcAEimkyGz9nZFnzEpp5FCeN3vmAf
ZXKE79NTrLawYg11FrTzH+3MAg8ITYlyV2Xv0q1j9T8oJAW9j0PY9vXidVUUoie/4zOPuTyP/ySe
a2ogXW4YLrHlIT0TgXiqQXJZeqAFXwlElFUxuasSA6ANsuEHs/lPjlWHmFgP0dRslMZGHD6YXdOj
TCaYDW38mO9AAjmuADVBv00bXQC6hrt2UIYXKw8l4lq4ijpt7wd3/HQTb5Sgam12swJr0uzLot84
NrF628Rzgb2CIWhWaFukLCkvpnIBogT09oxOxD3UDAY++8Y6brbsTirCpdn+L95FLmhC6nQSDYe0
Ai6MHXbufeflsbRu/rhqj+8fqn9yf7rqjjT+beqlYvbqXsHsc2CErjEpmuTPxnwkeCzRUE7oWT7L
9Z5W6AvZPpkx7TXlT3XxY2DoctPVc2apNxPMvY66qwx0RvL1Y58VYdTw+i7+UFUk9hRChp+jjzop
rWZlNFnYi7jLy+Cs1YJUZXL4MCQFgfRlKG5tM+izJMAV2IdhH1qsM5qp247tpOoVSigOoeEAG4uu
yIG5zsU/e9x+BesvP1KzoKaLgkgUwgCKlNqOa0Wa4RgFCa7hnD7q8CkSsOd/bKvG+7uK2ypEsUeq
cdtKhfFSx7h0YGnBPUQbg2JdZ28YVU4CY6CqRwN3naWWeFDvKSk1TrU1iKyxhdHMHCv0yDplNYkX
Dw8F7UvG8bu4Y14O9o1yz5qknDPS1UaO+E43YOZNsN4WIAod10gRpByPxqRGJJg25CIc0HROTvs4
XxZgbC5sKquICigRLwDZz728aqaNIXSuv5nOlRsXp1tZJpVuRb67fgB8SvxwmYwhXxVssHXcyyvr
mpWc+fjlxpdjSKO9/f5LjWH8myloT1+iAPvd+/yIxQl2dWzeXyN6NYSG4fwcQruKc81LX8cJ3Vpu
oJLZdqkMFXPglcbNFKm+KF28ZwfhJrmubqA/mJLc3fg/rsqy/VYz8sn2ELbLGXSkzcnePsqVnF29
CWGPI3RcOUwDOGkpIlEE7aOYdYAJAnAMPoBTqnaCuPHb0w9ubhNzdaI9rFtGobfV9bwPXc8K/c68
mthc8MtPhf49ABsQzXQIoe8xGdzm6b1MUhrpJmzTI9l8X6MCjU5X1Z9yUSUwfJFCtpJ2ck79eOGy
9HjKERswu35jkmwJhao9VWvUSs7jMKvPwRSNzTSFSzlaVa02k6Pbf2Hk39NeI3bGcsiWkbSFsGfn
xSer8ecMujE6LM3yfk2Lc+3D5hKhQ3FPH8oi5TPPXAk8JrbjifFfioLlsy9YXdvDZ7LvmQMb93lq
PyUyXPTzRHj7zZvQcK6nbAvNNYA05SE+YzupFGU0EBWeFmlE/LjUGsQk/vW/b+2n0F3tMg31T/9n
cXjruG4CnBaeFltcIcSF4LKPw+xoi7qJcpbQHtt79HgpuwLxt0laXCdy+TxBg/Boad/qTD5fK23V
bTvJFdt0BL9TNXlvjv00P/DD4SQEUbCSsws44h3Xr0D0mnHARspyUcarZHAC0P5679iGp/oTJAhH
16AwVh7iXTu+tHjZO31m2vshodC5IOPQmyGttlBWTJQjGCnjCgHie9z+qvB5pVSFzmgyD2dpEZSz
HjZCYuKFLoDQELUjpUpMEEtpRVM79GeDuLLA/4QDWmd8H3en0KSc5CLgNkQvO9XmYA78lR2JXfHY
vkbDbMziXGoQF4p6oT08K4v6NUa0taBofAinF1nWZA9CFu5XomJsUmDy9Lehd94t8pyRopBp/Nfy
ZXVX0L4/f7l6G6wdna7Pc23xXLGJa+3DzB800CSrWVXk9vcTyCGf9Ty6nb80YjaPxipjezRp2b9L
zoBKKzuSlLETCOQynYMKjVH/Jvwr4z6986RXz91PyQBNrDczcH4i96Kl7/iuhf+SRAqbMPZe5VAL
yPY/cbCwb2B00ovm+lCS5Nl2G2R1+M3VNCst2QuHlpZ/LjiYQivfty4jrnUg9y3w7vx3srGLqMOa
5w5sJwzfQ+V3GTZ353HRSy+/f71KAv/TXXOESseNLg+OPR3hlAkl+t/vJE/pdrGKHIGU9x1R/fYv
YSyfRfjQobI/B+mMxSqQRmFoXe7sX3ZUMQElR+03Gc6kVdpS9J6l6/Jc1ZUSPWrHVOt8epbvz/VE
h09K0M5nGvWAOAP1XbWltdf5Vk1DqKksp528LIVSDnJR0k5WEESw5yLgCsOM3KrXgRKjJPRQ3s1F
2joqE/85dD0iWS1sFX/82cxJR2kmfIn8Y1Dg1h8bxmpUVt1MdXfNZHF/Wou1wyuKf1NSy/Wb1Im6
rwRSb3l44l7igeuw6wc3V2stOS+GOM7vP03LWpalmARGzsIrl5PuCBTfsOGtGUqXE9MYcdVmnSxX
rhmQ6/QEbP5+zev068OQ5IBfVGilmQLZzjR3b0DtVLJy7NXJ8ldYvBMyql5OZ5EneyNJ18KZBZy8
Xw1Pzv0xyuJGMPUcwR6iFVr8VdSw8tjP4ZboOo2aTSoqGxU9LKIkzVyqRWVvIu+JEVf6IIaU6rVX
iAqGj5+oUYbYC5uEtY+7xFKy1tgNmL8qgLgxcxhj+Ksr0zvzeYOtdy9n3TbwLzJMf9fGzWYM7qf0
PWgBL1H4g3S4s5o/s9JTXiejtmIU5U8xgtY84+Md1pgLL0SrY9b6+fGaUNpoFlljU1NzOEe6Hj2Z
/rYt3TwwbBNJOmyHSByDXkPJeACT32SllkatkVY4RZvt4+uX+EQLV2IJ0YRZy6nQTEEneK3nmq89
GEZGVctXL3R79Ytnl3hgM9MeJuj6DUUninjzGpR55SF8hSGOZd5F/cAHdkwFxLnkwYoCFlZ7pCUg
klK3GFZJB38hKRbtmcjVr0K5Sb/gZj7ykYO1pnsOLfX/g+pnbiJaKpWFBQ1BXNCLJOmh5+3f2Z4J
Nr3/R1DPjWEQzChtwa+jfEnc92RLMprmHjM/PhWqLfEM/Jylrv2PdUyzktYNEcrsb/6xqMr6z0R7
gUY+Y2owoFMxraEgyJO41Bf6jbqp7LxSQm+ycw1D9sL4Y6k8FXN68euY2SWz+eI36M606/KgqgnO
lE/KIyQf8gS9ItrrH7UkGydwvUASasL5VoEoSjuDSl4/kkG9K1vtfSWyb223Ux+HHLDg27aOTaUe
ERiHGcl5wbDUqwM1gQRN8FTmX7aQqqixVAMgARnLijoqR9SLvFRvBMON3ufAYhFOBK5PewpsOcE8
qw70NicUob9SrDzzwqEUaPbYpt+T+PmW4l+8uXOrcUnd301dxPKwo489fkWJdc028BJgAVtZSua1
+X/twfYM4NGWYWHGDeKaPobEwABNhLbSvgPbGW9bkKQJT54AowLIuJSQN04gyosjgCva5DR7pDpS
fLksJiUty3+R5+f07QSSpAyL1SUJSWByubbY6XU0Mvm5o6BPwl1rnka0YdPw+aA0XEKa3NDMVvnj
1knCPbGn9oXXR+MnVOR25A4A1LpdQbAuRqHnaqp0YNOPAgrYg1DC+Fx4ulBoRcuhLa0QRupRGoCX
Tnt0w20u3R6sZ/LoYlI4ijKdRRHr++/yrZAElWPCodYuJpHOy34B5G840Xx9dEnkKDmxZyp+5bfN
fK76d9234ndMRt9nGf7Jbyz7e0QO5wZtDUmTbee1b63A0tdSo2FSwibAb3EdMRv9GwiQcEQpLr8c
vW68KCUfAueXPEtOhMmV98X7L4UmaWHv4B8mMPwPDNVEDTS8XQg0k80jx0/iFzF4EhMVfqAGUWt2
CoVkcneGunLTphk9LNZ9EAquE2HSKUM97tVUs8Vi6UoezcJytFbTXiX4gPCmEY3MsNHp68NdqPsb
lPqYimIRXhRKVpL1eodQWr7FdIeqVlTE38GqU2yAYGomOOK2AjLwVoRHwHCxA3jMN0RJaZ6aVNQF
SvlfPeQ7PGESerRjOSXAuNat6CVH7oCbv70wbn67rfWAMBENAYfukahy7TkCkrBctg72RLmJtZ2G
XC27KVf234ZmCLwQeUBzc5REhOEA6X1YP+54XpXouqMJItiAlThm4IHLgiHyJ+AE2uOdhVtx1ivZ
ybaf6k2QS1iwfBnmus/s0h15r6RupYQDlgZMsBCchgvAlvQYRd5gMXVb012i/89046FKbx+76AGw
C3BJakTX//tN3pMUk6hEdyj358AvSx2VM/s/ix9kVyjxs7iQHPfKHiX/YnicuiU52RAwYdlJq/pU
SaN6fmzp4dP00oNrA/m6BrElUyK0FlBTHXA7wf1mUpFXiLApkH4mHb7Oz3I+LtvIpppnOyXh23J2
IFLQutMltQ0hh3/2VR1L6o+0ySfMEhqx63WY6DhMtbr5GfaUiSFya22KrcXkLX3j4CTwjZa+fkx0
KRiGjJmLbZJz4QOtv+Ovo4Or8K9/YPoCSUQmP7RM2FTU5Zdd4bBGIQNiZXUFOepecyGTi5PzeLs2
vDxTlJCgyOuhnHUZaOGcZ+SaxifFiJaMnH8r+C5nj1VLZjWN7ZgAuHA1f+q2+esDP86/glNG6zLx
4h8SdAityRy04tcBkE5w3R+9JXcGKeJN8n0FMm2P716FOmjCvmCubk1DZD3evQTiqjRc2Bj6ozKe
NzymaSq2IMAzlNZhQX/avl+6lPbrKzfk4T3YdaL/zitXDyRJGBUT4GiDgWzX4kJpnxP6WiNtDrrj
uDmjcwGZxbA/FGj5I1GQ3QYcxz0qkgVHhI9zFKLFsjyIeKvIhgk8cjosBFAZRLJMpGQVjLXPuoC2
SHKn5nCTdwqa3ckaOwoUUKKL89Fg3ON9pBr57GHRSIkOwwR7kztVuNN1NoR5L9Iuie+z4PbFTzRg
x/Gi62ez7jtS/L3Bvw07RNKj7O0exCeEbjYKf8+22WhPnusdhxIZdxfDhUum67VNCN4Sf7M+W9y+
XsebDjPkc7oY6N3dOSSCr18lT3uPRer3Tws4/2RuoJzpHnV9+aFuOE1kZ1VTq+1g71OGFugY87nW
2w1CTMwBxWgP3M4nzqnHZeFm02FAvMAw3rW6pznFhCZRj+adeqT6mBjIc3YA17qgq3acJSZLguzT
W4xUj5vHiDoO0r+Cjoh/zwdyNiLgv/dBj13e0Dl310T+groaIQRIesePzROXvTM5MzIHvaKXaUbk
xtXtsuJ25jGJLjyElikP742l5mL8Y8004BoQ59BiKd8MTA4XYLniVpq5dni74HVqB5ZbfCuv61mD
6t0y/EZeUiwRk1aePqAQvb2SS5aoJu65f9Lo9419fAHiMc90xhWTyd5uX8iNzMEfX/8WZGZFVfgs
hMHTc7S9u9cTVqohExFVbbmb6sSW6XZkfaaXIVcKCK73uqB1AkuRrmE8qR6jSuUzYUIHb8PNQZ54
zEWj7itdJfa12mVBD9DjTtYSiLXlONoEihQTQcVOy/jLbXW20bBQjONUJf3iK01pFmYN3UUWSH0a
Bc4d/+ckI6S5yCAZnKIxSX08Q1kje0JDKNc9zPEk2pvx5iNJ/FHkDQRgcDkxyyvj7wKfMsh9kDNo
y7WPbyLiczqJrgsGTTO18x2pWINrOWZA0I8b8stM3hJ6qOuobexCpUGWfXhW7r7U+nzNMlCv0d2K
wNsIYHUMy5GU9dQA5ePViP7V+g9DMjU7nFZ7/WRNKuAexzm9JzrFbvCJ8rR+UyEELauNReNFF/Lh
ClG7L7ivGJlb16ALkols+59CA+akzlNrpAK1PfWRwGjbEseh0a1pSov9gjGpps8W6J4+2qJ78wfG
p77/J0SoA+7CE/IHKM6duUeuiv6nR6IJvh+op5f05OPOjEU2wzhyzS8HZT5vpeI/tnIhFtOe8yeQ
pk8zaaZYbpo0WW23GzEiTOn01k1Ulp6DxCM1RHA5kNBSzmbpH0YjIlzCSJNOzH/wqtzv/iIuwt4/
gvSKzAJca0QTwX4U4LxFpeDF6/t1FJfJTsjjViYmKQ+RuzTGYAdhLKmHgPLoqVKyc7I/Adp6t8wy
6IpgqtC+cepeuvJWSgYDnADK4ZmkbmX0w2NJuBu7g1pDpebbV3+sDdUpvQ496vQNqDgi/Md+RJ4d
vjAk6FZ0w7DNBL/IDhyzpGQEFFVaWSMQKQf2tg/HBU1y299A5Uewa3tTRZ7EzzxElVrhbvMc9ktj
ROETl6wm3hj3tf6UZYzAOTLoneS7AvIKl5zi8BPDUiUCV4Y5RwYA83aK0/LH1l4o3inSxxa+Rtg0
uNEI91grAlDIKPYBgj2mDUT7pqU5bQYAkyp4azGPi/gHP+6LydyIEVDSTI/S88XWoSp2Qso5omhl
oxcNjFl2LIHiXnyIJPOMv5PQ8XubzwebJ9TFdmH9Eee1h8UVlyi68sze2SMV5zXMKrPaYzuK3302
p20OO4d/b4PPaUqVjckhZu9AGF4oYuzOsiWZdGS8rT9JmSGjGwDUGF4C+52euJBztKvWKU2a3jM2
dxWJafL+Bj02DipWI2zqYpmkcfcQ1aeYzF8MSl1Znh0oKZTgxiIXydHDR+grs341HHIDZaGEzZz0
XnPZJ8KTLs1GLOfAlrUIJ59mmhG0FHpQ5751iqw32rhtvMwNhHXb8bYu0Z2ZckeddMH6sHAdOl+M
mZ9/DMmgDQxJzPhm+GuJM5KV1/v/rnpj6g0X5L08kyVGrdd0qmn3+v4TevtME8/BUghNab6WF35p
gDJIhPkSYoayEbMJmjMT7XqxoO6GBjn0WqalEyWmDO13OKazU5FyPwH7yQzozCxBfq0pNZH6isJS
ckq96b3jRMCNvbQaOndTA44Vis4Kq/0JaCnjrCo8vBddXHAPTuYhOlhGGGig4HfL7z18I7ZHF0BA
49lymm+wdMCxFQcjkYyBuEXa6tU8F4PfkiiBr6hhlpy9AYy+KGFde5rSMfN3kLTBnFgqt+f6BQaM
m5Q7S0VOYRblBVBVJCCpvTOucl+EpuH1sNME4PxOnNZT/6agOyKI7B8aofrQGtNlszXS4vC72Tv0
X5+5WEZiA0Z1RsMcNvcPtE2aKXLn7LN+nzfStgapUDRTU/M79fJhDB4qOSOPgHRfnL1QElHa3B7k
vkkyPlaClJHWZNXY8XsAzGU/3rsJlzd3g+ybP8bqjxj6TZF6x4+3xfOjGxSMIowxBBLOvBwANHkC
OF37yz/pIsCe8ta322Rv/PAQUcp9R09i8xRWUu3fvk1H8YVBii4IeilubVupo9Ti6BFxj34Vgn6n
PKvIYejpwQHSF54ztqAmT7DodPwrpytPqOr2VCCXszlyhXyIwi/IpXsZFzQVN8i5mxO1FijcLEXu
0kvqdFfmkb2qwTZw7YZl1Z7GB8gfovLptyiDolyr/Il8Q76Hp1jlEx0NZ1T0c3MrtShRmjlaRZTL
5NNkyZabzNBb+7htBMeYb7e/u/qUeI0vk36QdbkuaA6C3krIwVwfOXDy+y6U/CIg7hQ8OWbRdWmu
x2XvgAim+cKS+nEMwPXnZnK95FaBZBVEKjhWNc597MK7njJCzia3dk6BL+hApHo/GOBS7QoZI0iY
zVL/wR+/NMRzZa5Gs5mlDeyYFyYcar3NjmBv/o4eNAOLO9u2idP47vdCJ1kRPda7Dlah5vtVIoi9
hQEFQztFZEufJXHIzK77RKFmyCKiWeMq0fa/EvQqD0chYZNEJ0jIdiosJ60NUEqAWzMcmO2+QN24
32xxF/OE68aRFtC+E/HAoZ+E1wRtsysNA6rOfBNCh6X+sGw2YpS4P9h1EEMyz1jvWig+N0S77kNy
9OvXZvFwAsC2d0flRF9MPmKxNvuARQS8scPIygD3RHNz9JDt+TwqdSO5R7iSq6zRX/i40ozl23sC
8omj+aDLUlzk6+prWWMUb1lXDyeJ3MrdyjcaQmKuE9gTB4KfiqMOyiJaGO2TzJoJ4nGFvnoyYd+2
wsDWik2lMvlYZbFyzxR+IYonOqll7rLjo/AMqKwdfQEi/6uElFq3mHfGl+KHvmOXglRb9ewywarj
zpP8cu6cPhc5n59Ad7XDBTvz0HyuBv4rq6TC5hvy4WG6UpAiRb0ynxpO3MGAUCva2ElMGkHCU+kn
FRfHAIAKQXQiKRPakg2M6KpW1PJlPgHSK712upK+jn4oKvHyBnAgL6WPtQWUe533RtsLrXDViq0U
nX5ubjm52t0cUyD72NS/FJyIkUqLu1Zapz01oysDf0cxhiE+e7mp8UN68N0cEqAP37TMSpj96bk9
wJ1Ld9nzd9qtQLHito0fqJT8BLPPyGcPV1spQ1p6+uHpgEk/Ofx7a5d5FAWMPfqk8iE2Hb81yk9c
TlE6cb9QlVTa0Y9SqBZHwGDx7AenG5kkBmcLNAKL4Nrziia1YewmwsH4ihM2TglENhU2xvPqCpOk
+n7ctKKuFeu6u/wxhKPgIgNa4efLV3fUPUpTHuGb/tGsiKgBcjUHMuimVOh7tLTswDdUfPRS9g3v
RyWZ2IicGKFecLe6wm1C9gzG9jH6AQ+TSVon8rrv9d1zZT8w6w26Vdypi5khatbUjWuR56c8YO7S
uxa4WypXtPvqByH6KsFdATve4sBHNm/RGN5YKYbtu9Bw1NiWepgCJnPMT4K5qE4WNA8d1lp+50y0
DiVqa5rZsG0k/1kA3Tk1kOtsSZqYmVQg8iQ9Yh+mw8BrGwmegAwyGOhlP6dIjxyQ/b4SmTS5H0FI
a4dfjU2a+KnijDO2N/wwf75ltFidZlnHJqKUn9fx+gKiASSxQGAUtJymb/Xqoar4AjcUDFrb4xxY
lqNgRLId0SwVKHmZOhpmqfoU47x7kxvQwD40XdkHXFs9uaq87YhhJzq8ldiRb/OIR3I2htihHGpP
vGu1qYXMhoxxF0VVt1T0p83NErLL9PUHuCaPuRJgEJ7gItrPYsvlvPl3o8CeCbbNdykAP7M3lRst
/DAAq5ykKvTvR1RePE14QsJQs/Q2FkIcm+cWj2FNxnOS3zFAlomxEu9Jo7GnPglkYV73BshTkvga
Vx1BHyEPQ09HS1ffWOB/+yqJIqvaRlbl4JtaSCSmOGxkxswsiiQ9/KFCmNZG5eYd1Mtm41csYxCt
SMcoUGiZtoUxTrzP8ErxNkledn0v6FZUI9S1tCUps+7elt5Lt/J8+MGU1qPAz4RxeYec+M7BRoSG
hQmYTGPSAPq5UWiE10OxuCQfG7jGpTpD6wbxZlA0YGWn91tQJKsYufGQphpSKPRpz8Q4wMkn2eGa
VU/farLWeEdS7tmr6QaTqdRU9Pf3yVFgPUHtWo1JOkxEkBX7QqAFQ/X7YpGYrcF9I/DXITQuThwA
Yl0LGwFrMWgIYaadjg0XFPPJk/rFrCLSLPNYcEaucbtH/+7KK/v3nBpbUFTM2V2Q7nym0NuTb9AH
SREMjlzse+XZO8X7po9PyRYmoMT/2CzZLYgB/uSyvVqtxi5rnR5jtx8/l5KpTV2Aiq60xNA+2iQg
Hy3w9Q+2qTuyameMCOtW5g4rosMhhVHvnI7un1ZcUaXmKAabDa9O/wSI1vJ3ATpMDh5Y3gufUfxL
c4IK0Qri18P/I+KCqHZV1UiV7MDxEFPjBISUwneA/AgZ9kql9jq7q9bYQYdkD78CtaudkbvK89pR
Pxzf0ciOHCBAiiWZHD5iILpo/Z9Rc4cF3Y3cIg3fsK0PQxhZVf5qC/TL6cdb4drYiRYdFDYe42b3
CBzsNgKcpMjD9SMg5lnPAE7lZ6nlH81GJ38hbXwZUrywy6i3CIIme/YtqLPXGM4OVop5xPjETC9E
xqEgOIbVdahKay/C6qnjRZStkKniwM5pYCMnqVlzlBNTlJeyoBOFdIPJayEU4AEJQuvL3QUEZuFm
kGkM7cs/mujDl0l3ipR+6ru8PlqwrgM6Xx93F88v1qdYwU9VLt3Y7bOfabf/4ZKTMeE1j0gkcByC
QrKPH0gRkKAPcBgVOVcFECCDLRliUu3X+USvHMqjUYFjHPx9xm93LPN5qEndrks19RMll7pmVDkP
IyCPtrUk4bHhrX7DSCbhNUeJMT77Wrq6G6YlQ6EcwOmYPrwQZiwGJseNndKx/IufacjashK/5CHr
TqwwQDjpIIApZ1oH5y4qTlDYJ8sJjX+OCG56+eHdw4FkjJON+kITV+eW4fYau1loOG8hUN4zcIWp
hgfWqJhbI81R4DKejpz8tzWCm+loxT0tyb2T2JhIayWm4ip+gyRXguC6714YF3nEOQQxZzsOQJHA
VeR1j1wCgBEuRzH6kzzYfjDM4Y4TA0o2URHLX5v56OWz/GyVmhrIDkI0DgBRkIEg/OWINHZT6boa
klK0RCsspb3GP9Vxxs9fr0PiluLZO07v5l8abSVNScS97vRHKxeQ8wtxdSs7sNy9EoF5E3bDF/IJ
oCrb9JLCsy2qAhCF4oxEqPR357u/0i1Tcc3Y3hnRmToPbSwgRZCRiD7/MoooVn1D222BT6dChieC
xeJzdSK87Hhra1A33fIQ1XRGhhum52soN/MbI/FvrG1p+xozTTYGdKCoM4unfR+P9NNlc/mTZZOB
zrrGg4+6OVxhmZcnIt6otHOxevi9zUEqf5E0BnHhf6WZ9EQniyn8oFfroMoJKud4cPSboVsVezUq
g85AbRBbMooKQ1YKCofTIqjQUpTNeIpe9ZoEsmvLplsadoDug1gp/8bocMaLu99Y5eNr7Q6c8tWg
2iIVWxQJmp7aOdC+xAm5FNJWzXyvxNHX2PGCFplgFear9EwgbwcdFrIzToXL7/Hm1V5UlRJ/MMzM
3J2JAEol054q61RahmpKG9CNOH93ibTbpKxknnwgF4av2UAR1k0wWbOZmyu+L5FgzZiTjKgOMRaw
8HgBnpXs+tsabq91MK9fBXM0oM0qvmjBCH0auaq+BA8FpiThJPO1EGHT9J+skIvKxdHrdG6SBgDO
1GLsY1wE3VV1MepNJIjNBKOdazZI+yk1ZhMgq5nVEmCCzNwvnixW6y0Cql08ZRaVizzVlUvwVmkR
UkKL8OVaRctC/+FC6L2KtyFjMYOQStTH+8GppyaDmtBuAujYVswjkqa8m0d0aIPGsxTzNNUPDPoJ
RZGbWuog17H/aPIUny+W4gkK7aRzFJFXL4MuwmYojrpku41OGGfCU1CrTyD6a3GQxJd17+3Mji0/
cumAGzvvLHwAu/+E8zjqN9Iw8xgxpZCRqe44LfsHjE3SF1zdC6BLDtZuGnMPVloArFmQFU9qgCna
uScM/ZkCaOcN5TQQQXsP2ihFkhK4OWQfj1SgH79o3LXh9NHQsp4uhsA295e3gsp7ZP8+lvw5lGDb
sRjCpwMaMhIw4EMMLuIumMx7rL3r9BXAArBNyCrwa0rHcnfe+xy6GJMsXh1QYEWSQywyxQ7hYEvJ
eN85SuWBKV9p2lDvQjkxdhPI7mgmMfTYjAoSb1f0QNODM7CE6aS67whXo/tb7m9v+RCYwpxECkzF
ZPLWs+v1NijGfa/QCDGUPxpvBVLZeTklK+T0v7PCoKOUVP02luWHiyG22H+LzpOhfjDV16IXZr4l
9HzTiA2pRp5m8kn5yAm+xiM1kQ6P41JJR0T12w8FYr0ET/Vjo58SOBd/Yic3vpsKQvNGKKjVr6sU
zFoD2iEI2i9x4/jzg33gHd8jDqe4xWRJbmUMBEd0Mi0CIi2v/4OPlHkslqieNKr5mr4GQ3oAtP6N
KiV2iElYueZLOHAwkv4K90GjcbmwSD4gQDu2e/HAPZSWlKaugktwp8hZX8Df/ohC8gmhQwtvaCfp
KtLZNX4JSzvpEPTOa/riSCNTIR4wbCDe+t8YM0qaeIHioWrsZoU20LFen+ZLH4DmL+0JW6e5Qcxs
lOBk7klmlqhNeeL2x28lw34lKMzGwu82Wi0/WnBY+qIqGWQYsag+X/IeJ3W0SIDiOjcXLVPmGMEg
eqn36TeOdLWzf8hkhbad0dezOHHA3KkvKuUHJ79k3o40wtnAsapW019AA0xgAtAGcybwDK28XwcU
C7CYJ7a6bupNrvNh8na8fh4Ya7p8e34MFYx5OHiLDnoV+N09Jz4ZK0sYWNkrWp14fdPQjWVLYWEX
z2xdIHs7zLpkNNZ9pGWA91Gjqq/vemf4fEZ4ShPugwN266oQ7HGzdjaVwWXiMdvxI4l2toWk3Ubq
dYADqWchWnZyeW/5mTcQWR7Qo9jpe69KMnh4Nfq1jwgFvG2q9ttRNGGdghoUz9rD8r7/YknsgVWI
9fbLgEQydF/QhA+iNRv5g4lq53T3ZxODTl8HPd6LQ/gZeAgkzXn9QBGHRCI0UpFktNJMNQjZT53a
a1rT5btJR7ddejhNGJTpyboqhrHudH5br3nBB8HGovU3v2y0paNCLnFJSRRwTNa+KrJ08AMvTt9J
IGuABC19vFzKxG8xi+Sg7DdCUjdCpuRsZh70Ibaz5OaSaZ4HYCDTcgUq3K9ifOe5mOsfgh9tHU8H
YHgXqvqe9B1La4aXm/ubFpigKkqUYy15u5zqOy1APlBHELGSb+BT8derLHeWn7bpEDhL0GuurVTh
XcQjI5Cdfu5mpUimAQaH6IKsGt0GnMX79dI3XuZ6NUrMuudNkH4h6txvv+4DgPasf5LLPNHQbJfa
ujTB6zdMya0eUg9SldQOGQuQYU5IQyokjroxSH+CTLKNJJWZTMDVR0jksG/4xhJQLv6fHh0mSLdM
GcFf6aGF0rZb6mbd7fWBfufXouxEokDKRkGnIpvqr1zSiRCrlc+IM/1WG1v3uSpMCq9phlPf4HOz
Z/1EtpcLSG0lsqHT73LMNC9eB/4+buasUCigyv16KY23goKxWYqyzkNp1Tx3l3xEzyWuOnOUwZea
PDx+KAallTo3z6ldD7jjecllGCL1TMzYpkPQILoQ/biIRJrrYjV03Sk3hGXG/wTznaxLnoB4pUwu
TprGiK/+vasTw48S84Vr2sqvDc8vg+AuCP8SW8PG3XK7yL3T97ANtakAr0CHITuLWE5m8emBfbHF
1XewlAz9jXdhzg082l8IZpD4VQxAEnJeA6hoLZMEIFj9aRaSzmhR+PGCixabaTNbBdR/iGoP3JKV
MBUfoeHnSzYjqroTKhI/xugdY6c1Z7/hqc3wSC2T8W6FctHMTi1eaKYujCUHhswuIR17CP1uWySX
eM1yr9VwGbLlzkA2oG1GU+ZDNY7N0GHFRGgPnpdKalkUmM8GV2PRAhRcYCIF5QvjObt/uKaW79vA
DtDct029xqflUKrIieLeGzG+bmM14foEEuHRGQYct9CftExfZK/JZqxHWrqwPw5Ya8d5mz/+TG9T
6sd2nYBPd+UskQ+pTOrAVeduvkbGq1U/y46QjIFCx/AL6+GshqlqmY36CzwpcQCdZ5jIJ6H1PVuE
Qin8a5ltqOhR7Lc7ZdMB1VkkEaFV4uZ2QniZxY+XWEm8f1LG+e20E71GXlwVufn5RVoZmDLuXLQS
vnruZqLTl/xK8lLr2fX9lwGfH9Q7f+OBGuLKTVW6pABoSckMfEGMmf217HpiRCh5osoKyiT1c0El
uQ2Yb2LSIiOa2OaQWBOdI48dlFAlTIfvt4HcKoJrVPVg57AEJWLp+EdWSaegxVanNpAf/EqTlhr9
rq2wyN14P+aYXFxlIoV5eOS7ukAuz3OA1oTVhmjswxyCCEkw14FcJZ/+UHnIT1qJ91kcbYGUMF4l
9xPxB4RuVs9fked0kWiSIZBXFiYuAgJ+zYVEAfo505UhxqRBrfqZ9a6T3wZlGdGp/+mecVEAL7pf
R1YKCmCXdHewstkPLerlP0GJbMLP58TdM+P70ABLC/n/2GJTFJ1S5oepfKmK5T4DInetZNyMxPtl
Sni9ojPCoXkcEpT34UocR2fqcxiUX/wOU5HH1e3ryFYUKftnROVSG9FofaU3E1i0+GWsKXrq43fu
ZnwLC8gSy9qY7Xrxv3hC/tM5HrFIjXn/vzmCiZqFa5vR+HqE6gnhxPgR4h3prN+rOPpi/kYvwENB
JockdhBWosBa3apZBw6LJuyU96wC/VvLyQNowfjHlwQY+GPlxjGcNE4GMVk40L2JKAqZs6fq/FPq
et57pt7gUs+jILSxzRboN7zguDx0q+0hkGjzbwHD6aEJZhqn8nqkcsKM55DM52Z/4eRiPO9ZEp2e
DX/3pDMCNl4AIm2tEFO/XariqsVeJW51fEHtF5GJ9JH5PYlrF7WXu1bkXxSWQR3d1Vb4mwyssIzW
yQSqBevImCptb/ZWHYgoEbyMRJhWv3IM/pK23vscB8X/ZtsKZV9V3i8yiJjAhi4PLNQ+ivLZp2Pp
NAajwKzJrY2gMCqsNcHRD7nGWOnV4u+Ot1voT/j0Odz3aUIiUhEd3r0a8U9RS6A6mmPzs5skCmiN
6NUPaRP+/c3YLfvitkgkewY8sZt96zImLBX7EW38DCL7KoB7OoYhk7vI3wiyDU8tyQGlbhubj1fV
Kb3i5Vi5+Jbmq4H0CGd8cB7AuLevsuErX5AgB88qehgyCrNS3D1HFh37Dh8V5L3Kxc+hdEv1YRz1
PO5leAd9+iKddZUBXGlD+Nht+XxVUvyIlDq1tUo74s6GfsrV/SoH9oOvd/ZVCEmh8TqfpzGjxpnn
umrv7rdblhxUjz/8aae5JJtAkJCZREVzaUtFbIXwENL7tZMK7zAItoZSBEfTxDhqCoa08RmxDcK9
DYM2djWjVVHuNdwb1ZxPmcWlvx2vJAZmkz5vKxwKfqxsOs0FfBQfaTWFPNFnwM4EwDIOwRZublsL
0G4Iv27v83orLSVQncs2EBPZGm38+ZPljjFuHUa910WcFmlK0cWcSUDNA2fI3IVcAcWJ0lHPQ1pI
Dpo0Aokx39zwiC8UtFY0cppuMZAkGN7n2fdO8HBnFc7YgMOohvmxNDnz6dL3OPZ0BrxHMN/qPD9o
Kzti7AWckiM3cF4s2/d6ntVmGzk1j631zcN49Yyod6iky+wtFdRMgbiKy7hQgYUu09JjKf4cNy7H
UZ7ab0Zq3mJpOoc0m2dz8xFDEtB13aKlg/9ZJT9N7JjNp67VWKFdwK7qFJR5XerGvKRROdwfwEAv
zqy3xl9Epsvj7d67g6C4HNr9IAHTpha1ezChFIlFIl0r9lWCfYxfEF0hN1bljSHgakqcvKYj19KI
TJPawnG0PQ9tMp+k1Ku9iHbx7WSUaYKFjSc3+rMmrPX6EbNrzUbbFnzOzsgEtHozmx8U72nYG9i9
f7uPTkQ3Tb3a6uLDbhcKLX5N8PYCTD1vtW2+lp0obMqVTNxScapeG1VNhoCM6Mbz8KXrBiuGMSi4
1ih5GXu3xafY8VZ7FdgQBFaf5zdUI78T7QbzFmiDUrANNRkKPtSLB+F/tuvzt6npFeCX89BFc4V+
KNDay5wCMw59qcy1Itt1J9ELU2Z3ReLXiQiGu36q9RVnx542pjmqU9EtQOYGohkjvUnzlL03ugk8
bOFEIKa08/ebipYTMeK6EhelAvyldovBcUUNmU7xsLa+1zZ/sL/8LmB/wwPm/WJUPN+F2v2fAECA
B6pFMaKNptCF9MzRxSPGdT3x3uNQe1jStzPG5jaZIuqQLTijhXJaAKwhZVOehFusWLAspX2Memnz
pYqidAt4Aimx0uOP2oxh/D89nYTCr5L4BFqCZvaIs87bVeDk+ZULJgGIR+b0cBZiJJJiMftMcPza
N5gHr6ogfTaC4wMuDJ+os5K8saJ4ccg1JNsMYJjeHHkU/SsDpT5cJO/f750TZfNvG3C8X4cc77VE
Ve6VWWKRwoOB8tUyO7gXqtjb7Opp8XKlb1AfIilOzu9KCd/Na0QcOZQck6rPoxT+tc9mRnpTL83c
29V6o+KAOxpWanW/ukP8SggyKtnbxd29bIzi3LpEP+in5FFYoz7jZ1XvI6Pzn/aqU0LWppki9YUc
385uHa0VAQg20AJkhFkLGMHVXgUhFURMSLF8NWJdzlFgpfrR4JN7v7eBSq3Fd9VBOYtGxLtEdOwk
kfOX1ZumUCfmZbgt9FY2Qk9Z7EC4QT1y55FaaWp3zLqZMkqjAFoa9so3uY0eA+QZrKFltSQYiC3K
0RLScjBNmDmm/9RxKhWB9P1vIkq0q0oZeGgiUSgDgkcm3wJN31fh7rQxD4WEY7IG+uovaUNI3b00
7/KgHkGkz9e/fjQqiXUBZD5OI5S/wehIMokaTgBimGyWFhnkNKraLC4Ur3hNoo+gLy68+ZypZAIL
6Dmu+hSt0EqAk363UKvTWS2MHtu0vOSTI+4fjatFVkllfaLsDmwtsX7ERaRlEPLgVJKle69v9S5k
Xmp1XNOeqZJoXMiUPxUTpgGZPz5t5YFHdftaIRj4g0OzO8dAKW20BsZQvAvhIUebeusBJYN1A117
6Rg4VDLirL2U8V6T0q/GNjZAfxsHPavx9KSePtZLVLGOYlquNEcK4r479voGfYVUSltPwDb6cPz3
UTHFjIAUn6dup1doG4dvKS+bwtZbPeHfYlF4KG8oVE4KB13PbNc9XMY9smi19LEKjaJLOVt+zg9T
TIrL88W0kPKQHzeic/put5vddu7X/xKZa8EkLbeJ+lFbf0YSVtgyTmup3o2LsxcGji4AOkmutkMz
g7ka5t8UmLh5LNgsAqHuCcA7dJ+u9Kyv4WFa+KyEC8fsN/xhGk2xADqZCdQs9iRwrvXk55SekOPI
1oMWraTglJa6UgMYg6L6t/ucVbCujwLtw0/FDI6d1Sy/staOZQTWrEdQKDRLgDjd5Gwsk48j/QHL
F23uz8vRYH+nck574XIMGd3w5xdYH5F4GKwQ059+wF7/onR5mxkg6TADyc8eo42gCmyLqwtzU2Gm
9CJV+Imvf6a2dwN7t+guFgt2RaN6J83kL1rPHp0ldBv76ZhMOJvtJVM2sgDWekZo04GoT57rg21L
qe3Owe1eTAUsZcepBGUe1IN5t7rNhk3e5Un4ojp6YMkUhF9W0VhDoYiqgoRVOaK2PKin6o/d5ppm
XGHlc4uJG0SXjza31HJTG4HwJO0QEckeaGnkNw0W3s0nKlhLLUs4EQcjuPRVTJv7W5LyPyhimPSA
+FMoo16lmr80+fRiVxgTHbqG2UNNHJmLSRHnnoizLHEob+Yb2QZO9gcvBskzWZhCU08NAWZDbfph
VMsWc3GJPZTKQWfIKC8ojGHBbKuo+0DuzFljCzzC92srJ7CCvkRpgCmWugSS6VqVEHNjdVfyQcON
I7Ezq9sB8ecMt48HjGxeWR4O2r/NkncghUG6pmlRGXSx2lTJq8w8txMahv0YrXg15r4bP1vmGsW2
GucI5xx6u2AJR+o0rNN4c2Lc6AtlIBZW4q5sk94NBk9Br/Wl4JAQjIop1XIBogLH760E+H/QgVWI
Bpkz0Ec448ysaQVWnoDzdZfMQbiYmLyIIxPaQ8LX+OSRVV1PIeO/0BF+PGzBwUO075U7KZJrNtFc
FvJLpQYr3P1nvTJT4VDrhBu11yVsCdR1uAn4TTKOzZPEY/GmSRtcd2nhnFiHBp669Owg2VSb2dz6
X4/N6aIsXwwNGyxL8xT3GmuatkW0d8tPqoBSw+MtWihD5Nyuyqtbk/Pgh98DpvPp4Xqc+umQiHo6
DgWIv5Vqe7jY3FUDsImQhECByz6qVtnw2NzvBdCt4iZxQbzINMXB2v4Qtf90jharNvvQLNbaPY0n
NqW34548ldIF8zisgTf0p2BAzEhja0iJLJAb7PU/jvCYyHofAFCmAUmMY68apNnxmgLBO6MYZ1KJ
01MUu5e2b6BoEJZc9TddT+1WhjN1prbOAReYgjGFjKwGpPbvWVio3rfWm+K5rYJSuORnnuboIMeU
2NoAJh/9sh5RIY7AbNBmGfAVw8Wxo56NrRkXppBE3IimMMKack+BLHZKvym9DP2N1NSn5d/vKt3S
YiUOFaXxMoVPqhY4FGO1txNqEJBbwRsYwoEVZ9UiqfrYDtvw2G1waI8lFqJTDZ6hi1/3J+JXfxf5
IGybE1ToCNIaCX22Dn2CTgpToVEXJGUK4Kl+6WM3EPEAeLaPE1uoz38I/eseHSWJhLjShiDAFfiq
2iKwKk4VacTSeFpB7my8f9ieXxCpQWrwg2eRJKTF3UoSxqohQ39hyKZRGYvODQJy6fz/zAqrS5S7
3XkhtJD4VFvOCv3WqvpNKc7FyeiQPQnicv+FJhxc6XbQWF3UA2llljhsAwXE+r7YApeclc4kTNUP
VptHeOFji62wLtWWISKFEywjFmQK7aT4Kgzij9nnl19+vulQPyITRBqXoMiuF+xoCn5yHKPmU6nJ
M8In2PgDlfBEHrOp+yfLdH+2JjMy16G8nvjERBLLK2xSm75gdGdhS/ZTVN0xrkxKN0X/a+6Bm6RQ
wFYJ5BxcyHKI3OXD0hOkcHeLtM0/so8cGbpyzK+gAIJFiQ6E9fJdwzmFjEwYYGV3o2R5Tpw1tZbH
fuw68Ku6qf9HsmCCF50227wj1FSi0eWpX5biCKwmUM0vPjjvdwCvgT9qu6CfzaN73/Uid/kYUh+X
tQabOHSyWtUUbH00LKBQTZZdPvu+E6+OubgQPktAjBkdzMMjCWqjSEW1JkdzEuD+1E4eVY6gaqPL
aGtIYlzFNtd+RMyS9jpa5QphEK16VfWHlx3PwsYSIbpxPunxw918b0RWFa6z67foktwbgZEFxo+I
HvKPOkw/zDAzBosFLsB8HRR8W5yIT2aBZjIepUVZQOX+AuiQMpeiMxslFN1JFOfgTDSne8+gpHjT
EVMX6svxjKKac13OCDId/H5dsJBtRXDffRRZ7YDhw5brKDAYWud9WgzUwchQJ83HiRCMmhzSl7fO
+DmRBCYuqlbqtP5Hd6PjWve+V64TM38hdnqVVhHrRUIbooL2D+E8Uzg4eTR8U25bjTiUI1Y5IDTH
wOLKBGLn1togEhE5MgD6YQKaDmgTFDH2Rzd6Uo122rF1E3Uc00IJbGBvuwJ/sXSjpZ3B4JDpuDDT
Qkl2bqWAJs4IZbCKa0Q0Qu604q4oJcT9HY1UQ4uvECqyHqyOPb92u8A2bTgA5GpfFqNqiT1xBnrj
iivOUiptLh7QTPi5pVb5MZPIE5O/bRIDBlxZh7Lw70pveEerWUP2+IcSAgB92yZYNNDwS0vrCsy4
mZpSjpJ2c26Wwi2Tw4rTM+MGmexjeh78hENxsUv8jiiFAQQzTf5F/s9l10Umm8pMIEPu9d7poTw6
ywGDA0JNLi976U+sVM5slgf/DFby9bHeT8HXe9ZYjlKyiliwjKoYVUcnqLNl1d/yD7u9L8Bm3VfR
3hRU4Zm7/NScy4B44BYSVV0MJ/V0pS2lYQhLQihgs0hkHdrg7fSybnLVa4rROSrYIf5TU9CJkDfl
vByio7lJFptlnOQQ/ieDCK89tmwzGscbOpLw+E7BtGo+x1g7LEEpyO3zTdCO1GjielMnt508X5Y0
56oAS9PMAEoz3dPCIyZ8pbnyIwz8YA4M0ioYx1DJM3wLvk31x9e7TuBxfAls8yHMFzJ7c+XV06tO
Guter4VdWIaJ+pmuwiDWzcIJ0JxSbM5vI12w+bqV0nEy+BWFksz89b5+eZeSId+3v3jk3YARwXlQ
nRV7KZ82M52svjLq/ZtFI13oITg2H9M8PBydF9/2x89YTiFqGPTwWsuuSrGRXg6omvvSAhFdHqU0
p9uTaYQ9yq04lkSuKLEJuczcQICpkSBGAT8baoz0/2RB4NxGvUzl/w7yZkgMo+TX5Yn9PaHT31Zq
G34j2yz6jpVsu0xJ1jcb2p9do+Jad9i2lnw6W4fCsBAAipiGUPVRS7J948T8blsFeRehY1npitsD
alVrrwKD16f7CvpbtQce8Me1yhBSpdR+Muw9rO+0+9CJGOZFpADcsRzyVjkR03W4N5N4ymNfVN5v
aPqGZWx6U0IwYpp09pnifgvYyinMWBo24Mq7ag4oE9tHkbPoEAChdpaoLvi5S1DuyTQUKDtwMqdg
/U4IbgbdU5EkRpWRieV9pNXEwONZVJFuns5lc9X+4E0myTc+rotSHtdKuS3QrviS3s7ETFLLvBFZ
uNAhF2ss47weiM3EPRbp+km6fJO5RmCn+2OwQAxOJ7x7s2wQ2VDjpmZHO6Na3kRcR2hcCERypSel
2jkqhrmdLjv0tEuuSwWUl7CHhIUGUbKWuRorRbEPqZlaxafJOHjxEWjPZdSdWsn81SV+XXRA/ERz
31tIDfVUw5Lv1YunapEqbnxNQMSX5ubykpJgrLwxdW9e8t1adUTsKGDBTFWHI3grJq+rAwt7c63t
/KyWgFSYifFuWL3lmiBZZFpa8ZcWipabd/SR2IsXZVgq7IU2jZ1b2b70bpKKVcy5LIqlAm1Bt5TZ
TjlnyNvMAkkECyVAYfmTjT5lHA516K/oE/RXiwJDDxAkE5FEjwKpQq3cI6tYTDKoWz4DrGK0Dqru
hAHILqyRPfe9A0KTQpkHCLuZ0mHUoRlap3DVD9kEqFmooqX7WTxIvcw10XwQM3LFgcS09Y8i1KUO
sKGVkt+/rBRwrcF4X4jlcA/fIkP1B2lpAjcJaSdJwDJS6VC8v02lYv11WpANAzJNJXePba/ljcLZ
KxVmpAqkB+7tAzOuQytdxH0X2zAK7x1+z/U0mOxokGw0AiHQaeWr5+nzXgZmv+Hy7Dk7oInTIomu
rzYRbaEDVYoeWjzeYzUoyH5MpZ6yZJJOeFrEDoIR9IU26gOSFibqho676EuklqxVe6unTUMl98Ec
vriixVVeuHOe85pz1SIMMue+C7IERiCz8LZW8ja4UsLAtFFK99hTy3QZ6gfWIb2F+z8rp/9ldeHD
b9iblFV/ceHL6fX+hpJ3yId3sgNa2yVVfuBTTRVDldaoJ4Zn/2EJCtl76/emMVYXNhZ1QQ3RFp3D
RhSenzs6PEiKPtKzi/TaZ7cK89GVR/OvEOyJchF9bW37kPfhAkffchIAmp0FrixT55+8pu1/CJUN
ukSR6kA+rzvC4sDugVk/U1iOKXFfS5wGdZ680qTLgjr74OCQFNsj6G2bT30d2S6a8ELuNTy/OG+W
ItuGwOIV4Jf/EnJ9aatx5cfW14nRre/0WoHAxrRf0XAUth5rYn+KhIO/SbEZsqrm5BLY5K+sg9u6
pWgQtl6WlmFu9sUHQmDU9lx2xdqQUY10qgBtXmHeNsM0P2iRXzpk+SZ/4yaOQwURhH/Vhrw+kOEc
dpkrmy/50dIjmcgDEGxXl7jwXd9wOWvAFTZyKNtQVKkvz4ALXlHU0UzIB7cdrka+v3BrO/yDyDnV
b2CWKjv8/z+gFyyiwCKQCFzLYP8YKMAr25loOldNEmisMFv1AIAPE1gy5/QGmJq9qOE+YhekLn/q
+AfKOJBiJy/fP6at1b/4HjOEUAnVonSO1fMZRWCydEo+Onq5ANYsS54Wb8ps3BAqiO/GnDaSaxCb
UMh6R0Bdk8XlWGnES56TO/lcaX8x0+/AsWLOmNCIn9ZMzJSfmVV4M/ga3x3Mf+JftZf4oHI7SfI7
ilSGdZXJWPtGUheaP4Vj3VNdLQEcXLxj5J+0PYnigtV2KkzSxo40KjqgUnoV/O1muAwm6PwTrySY
U89xrS9SloI5Lwf6KayBVb6xG8AfXN8sqMdqi1tojoHLf1bw5SMoGXt6A7hzDokvu+YELs6DWKW7
00QuijkBrVvM4BCzsPq9eayyAKmegpHHfeNsvCj3KcerouOa5FUUbwhcLKzQQMuLnVs2CRM1Qz7R
+qXvsLOZdawltijcHfdx9VyAlECd88WPlGEXDGcQ9I5FTbbn6bEhbsyV6wvjLQzRfSXUkmE5Hf1b
PfWAJRRXKBoWg/VqbIQijOqFCXH1hdAS+Jkn0NMGAuY3vVH1C67CfwdA0CUElttIcY5zWkha2tMi
NCPuLR+DIIUngZJcfRFX/y1iwjyqhmyZXrWm0YcUL7w+YYHrhpYn8lZ2tW77+M33vWzuzAsGIlQf
zT0bJ2E0/ErbzcvxhxGwodTS4H/x16Ts0TdN+2ae9kduJ0qYb2FT50s6Xr+V4T7gzdYY3SszS+JU
LhRugOTeiRVVCAkIf4d20+CfuP9Cgqiyc83t2zxPa+Rpf76DxHbBPpPTuE94hFx+dJ9JaNakKxIG
WF6V8NwHqAdeuIEIq+XRvl2wFxRRRKxF/9LRyhw9GRgTKB67Ogwl9HibHR3+u89thSwuNuVD/gul
AAUcoKtCR5jlN1eUI5Pn5W8zDrC4EHhyIn4zL5LeynChJz/bDO+kIQSGNglJvs4K8+iGYvnQK5ZN
DYxd34F8FQ6YQscm3zpC1WnJUvW6hVRdawUdqAOLNugqpoMzdfQn4B1zUsukPxFoGALynjfOGDLW
8bFFsYaakv6eyTlyxm/nigtseCKVyirYmBZtKcifciCLrw6sz2a+P1tVZhw0UI4IFSkdqh0FfTGo
cryE9eCpFuubZsrqcb2sOuclwJetA+gxT6KG2jYVD9VPCSujS+lxjckHfTOy9owI851FcvcCdJAU
nIL7UISwR5j8rBGakuu3r70SdDXk9g/f+ymIb4npOTZAB4Xc2vRAWmoQ4iC2RLxerCgO84FPgVCO
S9h2MOUJyhL2z+5t2vopvQzyNedBU3sPzjyQCiJDbNHKZ6cCdIBAeDT8q5to+ImOJn4lEaQrwkBV
E41K4k4c43qZX1nrk8zOlFne3c+nKQnHfqh34H04oeAgrM5RoFnhC4KpfLlRmeSYcvisgf4QLtSx
iL1SAmsYGX2GrDzBdYAlEwp1o6zxeqO1HUV7LaRJ8SXII1JT3ndl0iFyJPiBkOAwzX0OB/TCw0oI
mOOmMITHYkUubywtHDcgMcQ/lxnbEJEs1+WnDHsTzYxUkPDqdwyWLtnmmIZb5DyzQ0WB+5sUns8O
GSa34NzpXcvyrVt9+Eqhccr9K0ksQRosX3h+4fgYZsjZMDoBX3hAmJmbx4Xp8lWqMGmDOffOthTq
Mjtj8MRtvGN95Q0kUKfhP7lgujuKnjkZmo87eXKgLKIHEvaKnq30JG8mzhY00kERFWBPfIu74Pwb
4pTDGqTSARuQhoavdadVf0HS8/mhxrE6eHez5NJTx+id6e3P7lwRNPQaYTUcRLal7ZfrH4Uenlfu
PjplmWizaU1O2We6vKdYAq8g4BuKdnK/8T+HhHSyPrgj6x/pwr6n8piU0wTz59LrW3yREo1Lh9P9
s4sGTG3cpHm4FEMhrxwFUgJaYG0WozDPcJjOaT5onIFvxhv/6CfFH0u502qVG1H2sNclWU4ZeDna
RNA4+iYvgTULxn2JPXPyj46uU2GIu895uAEGSir3bWE58v+yWITX58/1FjjUDMTXf9qK575JBDi7
Qqwykja2mHVOllKKX5z1VIzkgawu/cyh/pxz0b3rFMxoUc5Y1xhviRkJDGWUMgpgLl5aCanOD/Q6
OlXio+3GG8td49UwY4ZVbQKB+MMKST6jqoq5flcfehhGLxbpCBWfXd/gSYdLdAZuYHKr+/oo/qGl
KNX3J1/Oud8iAXH0znzlp1yP9XCmvHQND2W7pJInr4Vj4lot02ocRzpYT7vJKT4/EGWVYgmJXGCw
wx2hR27bpmBdj2gO0jq0DzpdXJjfG7nd3yIZyza9YRHNO2Wj+0zI+ZsedMB5DZijSRKHW9qFO+/g
PX8ba3RROGqM3f+lYw8gOhNHZicWSqh+slBtgwfECPwK1UmxkgOGUd72LcrXyiAueT1c5jz2ucXq
2byAPLdNLGwhqyzrnDuZs16xbJS4UAS5kK9Jcu6ykBSvDh4WpE1c8V3LrNxiM/8qap7Bnlcr3ZiB
xMJfDBRG813FXWULj+POf+ndEUIgJ0rzamLmcuxieT1j1a3lvx44rnYoQ/oPHewta8ofKPkqd/al
oNDDo/NjPAyaHp9XBdvFjaQalWuojVzNIp6dV765bNDauCURG4wC1yfOFhkMFMOk0kL+EAFX4Hho
olIvOzyTkE7MkoMTmnf225XSwaZu6O0JuAKoe8UGAunM7KeFoDBLZVwmJkOsuG46YSREa1KjHhG7
TTLN3KFatEVgUo/jqijfR0frQOE9q9aDG+E8FCkq/CPomZMsQcGD5BrzI+sT+lIrIgRt4ql2DKD3
lQP/KJLa6JnczINcn3hju0q7Z06l6dG8b36FH7gIJ7FneljCEIrN4ql4PpKPoEroN7Zh8U2YJebN
FJA7WHi/6aP/wDosPFvj7tfndZylux/ZT2VymFnQgtO57BZejxK8WTuVK7Old8zS/V34Tuc32XA4
WbHswrENX3qgmOKSfwRu5cJ4UMKKVBo9LLxbmbgymDppCkj2DnrIuttbGCgiezC5wvLVF8ZlyE6+
b8AzVdrKXlq4JRBlxtjVoRB/3Q3vvd+4HJ4da1y4XGHJPoDJd+MJ5K1OMcvvXXWdlXcy2PuMUcTa
MoCVeReApoakWuPg6fkXqj1r26yCvCARTB1h+761oziP4LNH723dg6HGoJT2JR4e0srJRpFMzooF
IFAtjo5qAF6iKG0rXh/J/m8uJWs21OvsNR8ScDab4hBoecsGM/q9xjWQjTUBzTUwqPolTGAuuUKZ
vDFEjhWXjr3Sn1VuEnjbYa0ooJZBFmbolk0tH/Ok4HaNUcDEKyjBWZiV/DFIzh/xs11xKp3rcTKb
OUCUL7Le7x705oYdVoS1lJKOrWp6yWx91ehnTnzBWhRtmcRGZQbeNOKelZyv4+iDsoqKLfQfemLp
n1YHyvtIUl1l1DjA+vM0UZhrYs74Dp8qDOufYByEoDwh7BnsKUpKwzpn//hcJvH7/NvrwgOUm94b
sy2z3VI8k/3Kcmh+c3mGkjfOJ3KTjS5JQF7L/Q8QM/FxwOdj9lWARpOLNwJM4oKYwbVdtCTD3fDK
NFaoURQnInMYmbK4rDP2kAYKGZpXIIANNCZRGjJGZQQ4CIKr5qLP1C64aGYb+Z+NEcUnmK7VlIcZ
wQs2igcF8YFvuIUdU+zUDquBrJMfJuoS6M1VPusaHXjt20fF95kV7Y8Bi5Qxw/6QbzWYUIpMEHuN
3rt6j+vNpgNFWaLwOoNLqSOfPOZahSGMKlX1nhpM93VYHgIWPDpuLquSYwCSyOUCfwJ3YyTq6rw4
eQOna06WhgOsc7sNNRgxs7xrR6ikq2IAGLCUbCP3ieROoYrA4cd4ZQ5cvRdYsQ3VbBRTRu+qKeZj
fO8dLogHiq0I69IaerNZxIeCHGAnAQc5VIITXBbL+SH+exaunG7Ad/Q/I0gNCV2JPglwhML2KSFO
rWYu7xw1Rl4gaxj0wMxjHmTQhUg4sH6bg1ZPUdbPakpIacJPEZNK4YKsrMpOtLh80IXBn6ozbXL5
OPIoZAGc/AY9NYz4LVoXU9BnVxkZzHKqBktGN9YWdolrctNexh/x68x/tZKuPfTJ46SQIY9FsrgT
zsX/l80axt3gR2tlGbYCILr8zgLfg3+EQjP6KDPTojjmK4bClp1wpp3T3Wo+jEGErCMSKPMRU/DV
JyrBun+BGk5qNKu5Mhj96h90PAAsVxscIN/h6SpfTl52e2jFLcRhY/ILr4zWWxm35BiwAtV7gZEO
ryc7alTgJutWLqIojLo5ovQE3tUV5cacxEFKUig5UdB2Jka4p5TiQZHM90v1M715cAiyyL8n3zAy
inWPJcRDeFq4sHrVPVpj9bkCQyhMIuIa7azexFBCfzZDwtQkItemMOVIthYWVkpI5ZpGHY2hQTSU
Gi7YEchxAKwlR25fA0kO4ikEntRyJQPSOakUno9j0XfTfqwUBBPzcT6eVwVxFpmrSVHGv3RDQJi0
C4aleERVX72UrVba9OW3S90pIE74NBJJqnk+pmGhbNN0lTS/laoQ5TKxFG1YTjHIdqt24Vd6ATcK
m6BkoDfO9fdB2WQK1yRGmZDDYQT1nmrxt4DumxbNUFLOllD8DhVO7FMhkSiZMgVVti4z48OKHl+y
YT/wW4N0WFpKI+qJx9zmk6mMEtZJ4G3/UhJ73bLA13LJj658/Vt5Q7xDw0Ox+8BfvRACQXkrDwXf
qF8ULf0YW32lZgby+5B/ybexIF93PA7tE6m+hLW+gVS96pK64IjD9LI2DbKiINd+oQq9XDoBG5Na
bz5NytrVQjiOaIIEXA+DAF104gd0EmLukNZkxNuh/QOLz5EeLbWKB686FjDJQDIEtrD/Y56lJ/NU
LzHiLS/GqEH6eHW+U5pIDxv1WJwCfPNsj6gj3CP7uTs/iV+V3UykKJpPt25Vy56SUSphxCGFyDao
VMYZtEjfsIcZQA3/A1yBrjRSYf4i2tisz/xBZOcZHoHIMaRHuQQ9NrnE02A17JtWoxQrXhHzyg0f
z/lLxCEUxmEgtR4Ft3fOl6Sgz7Gj6PmHO7EidmeTXIiiCHnPZz1+J+ywK7s6kQxj9ah2G9B5DNmn
LxNrG2jb2eM4OVq8ew0DjnHMTX2gsk/4+YxNThzQDbUiACV60vckKnX7+JiLh8FPHh3dBquhZ5Lc
+0oQ22FrFVEK8wHQt4eRPrmseSsVwkAxxZwW68IZVjJmJ5MfLnw0w3pEx9nLiOZnqKvopF1KEHUf
Kc2b+2/zOX6GQyxwhBAYZmwCnggpH2jAxAgZXFJ1IT+58VkKf46hgdXzOIAt5Frl/iHaeuOTnn+o
MItey/9y+3aPp3ZQDTpozwB3kkLV/Uo6Mk5ugo7FUZlB3E2BlQxM4NF5Eup4tXSvCkDSxO/9NaO7
45+YtsRP4w11yEAloiI2jP6GaSoz/hyNiUA8Ed4hoqyJ4WgAspBVTiKx3JcTdjj15p5CQxwywVIk
GuRSaDRPgtweFnd/gI4djoV5kntFtTLaQN+dSVoGaCi8Tn5JTgFKvrmpQIhRbExU/HSUBcXLnqcq
W/FMlGC795u1hr6wab4kZe/9bA2m7yxoS32MVINVbFyJEUzx9SyVjo+QFOpJaQg8w+EgvQ21c6V3
GNv/HDGAH9qI+IDeHK2lZjqXa9Osk/0Dx2KNZpSZH2/iyakuxk5mTVdJAyX2WivQAZ6qjSxP0dJu
4tMnKymOIBd/3aAMviB++q1IXhwzy4c9dB50HK9uMJLpP9WVqN2QSjO2p3yxIC26e22A+hXnHjco
+MdzJHC3/1srfVBwQBIZVU89ZVhU9KMhGI0/4R/ole1HoQYTGt1xd8PNFlRQpUaMgvt06gwPXtdd
iVRGeC4j7IbKWu6nX1GSrS57ZXw7SAvSZ6+CKebhOqVQkJQKNjetutgQXSf1K1GjXjLK41OnY/q9
8n4iNWlfFY04ZjKSzmkHma3BRhEyDwr8Ykdu+rk2Xfe5OPzLm23p+I8HdwDxLkhIQbQZO/LqoHf2
X2KzfZ718LiEi4mq8tFvMctO3+dBpDOj/cHLrSTymo3PopS69hybfkZskBXO2ZVPqKfzmWW4IFUP
Adc3VWLNFLZKwqxokTM41Pk1JhMNwgTkzxsrVusPDxlUGKS2Tf7zwP+/YQ+SQRJplwVBFrqxMHOL
zJqfh2IpRwjGk6P++y5ItyuOepWbhLOkc7m4ruh834HLVLb0gNarciti9y4UGBEt5/mHRjSK4nnE
yjpFp1p7RTjOtJ38b8HVbnOnRW7fodVsbAMtFrc14U68rWQ2F2JgajKbN6/IuprvNQhXkOAWGJDz
zDsHBynMfMnbtaAjWAutteJC/vUQAHGZBJ8utbdeRhaVIPidMYa6orWY6QvlqF+4RpoByWoJVTbr
eyyE3dMndzZQ/Sx11B0mDFxiUC3SYkkT+xb0rlLQNAuBn9tlTeJAhPHl4+jGEvF9UeoL+PUHHn+f
LXHjy5bTR2IccKcqZ/nn1H9YyUYh8FzsejQTSz6/DRpsbpNBr5vG1zDfdwcfKyj31GoRwUJiJZfQ
MkEGQVD1oQdOyC9ih/OrsBzNjrAvus3dekiWcAPbNjuyhKf+a8Ugdq7RQVRaLIJrLugADZSbUE3Z
0IV00Bg7bwSpBusk3ZBhM0vVK4uTnaMzYH5UPbpcVPmY7jSRXK+Qk2BgGUtAUGQDzN6xDUPXTEG6
CMuFOIbJDguDhg2ljxPdDRoR45GDE70qbJn9GcDx5cbSWVtFLsP+hWn9PjK8U3LZ2t//V5oxZlBN
eZFxnYgmeyw3jIi0KbQFLH+dV9aPylwFbMh8BA0wDuC8OVgG0NGixkiPwBT8SJEDU1V2/RTsQCaE
5uvTiojI5TByIbkYTcfNKpLDCW7IpeqT67AxhVSf4kVhZ1+zMJKSMW95P9zpvWBabic3MPbYxHh1
NuVe/daGRR0h/sRCVgmMjA5q9dVlKXiUdxM8URopU0//mRyeVjqnIYDoIIa/rGlMGC7QVWlCNFkM
BjPTjnhD49fEtETcMSHTYW8Rpj9fnZ9TaydyYU34D4DoJVXUWiNcw7RTneUgF4xxPofM4Tg0BLpm
73+/hozcKuhIYygxT4ujptyR61RHNU4o68G1mc5CZCjcqJiQjbhLcG8lUymp82oO9uvjdg03PFt2
x3AXCJVrZyvLY6WuoU8zR8iQIsjfOqtZJUvawP09kSiYqsf9y2Q8n93uq2BLQ6t7QgyQdDOxRs9T
rOo1tDguCNTBXuuMz0BLOpztigWigdBXwrwg2UvNUbBKbcJ9dkM3r8QNPGoKz6gU3BH45K/M5r5+
XeKtK7Ot7k4ztjWLmr/UZT8JFPbnRrA9drpn4t3JDGgSi4+yXCwOanIVtX+8oOP6HwJw/m42g7yQ
X1a3sIdrq248WGCL4z+46WaiGw/yT+t3aX2g+9ssuSz7/BtshaIH8Dfiyk7BLsz7bUN5LsnuuRde
/+Tzn/oIMe7K9tcuRO2w4rfl9xsJL3Z20+Ul7VC2x64K/1yXqaNXFGQ2KWVM/m+7sOw5lBWOk37C
OT/Apf13cXSwPlWTww6pNBCRYM5DMF5LG4QACghHiLwdFgAuBLPQGXWKk1/J8PZLARxRUdy+Pmzn
HRtcIjtPqt7XkD8CaKl9iwJB6ikmLDS4+SAJn0me9b23qEpMVAG99xRWpOnowsx3NCFtBmZT55mI
aliIYyY6fdASZRataIy58sIDCy+hK0uatRMKPfSIbmFJ71s7iEOjCayzOexuN2hDMX3Y0NBc2BqQ
KcR7J4AkWefFP00isybgF1dgXS/47xDgfCOU6UkGgTt/lzWrpxjHNVkxSbkmpIRLKDZIwxERKcxx
YoxHb3gVQZbCyKktCwFWFQ8i4yqD436WbnpKEsDyFxPJ4mPGYFJrcF42mDyWbPrCr/B7W7hPecXz
FlU5bXk4BYeBSk9N5pNWus3oSvnAWWU9fCNA18ijk/4BNwkb2L1J3XDnFMoBx8UIPhaScHHQWZgs
Jnj7FRy48wyPoeUQGBTfz4Fbp/HEMWv19OaDj1Y7EJ3TQUYXDhdNwZPIGJkVaGuGKIg4l7IWu4Oe
TIHfdXX06kpL1VuNO9hUrcPzG2NkXiepzBgEzN2O0+I07V75P2pvMM9NTNnIbSZvLSpwbnvYIbCX
qZRi9BtlFFBxOs+e6A3riqB0LcB6E2s9HooGasaoUiuqV8sDT7PuV4n2qKI587to7qmMz6RhLSfo
wAlaSDvV97uQvPNw+4DlH3bD+CDpTuggBTLEKMi6+xBuipxD0ZqqsyQUPCNyCFhS6ueaOmJD8rxr
/xAXtXV8t1lfcSqhbDYSeN3hboIRyVDVcuNCaLSjkz+TLqVlxcpLqI3TQ8VtAq33oJsRC/DJxpj7
qXSMQu80c11TiXzlmec5N/Z60IKJeXpq5uIWg9+kSy6XwFFOsdUWdGAz1oy8cFn8yY/O6ETHDOLh
tg4DMOcWZ/zLqQzBBeM3daWwUFCo4XJ9hVD9suyg/LhlmHy7cWeznk2rLoTLU5qAjAdL2yLbdUYJ
ojh2P2IE/FvuZIIRKzAbLP8D/BBTnZbbzK4aJAvpaJImmUcx63LWs55B5wi2mTs/kaj69KPHaiov
dEeOgY7bqs7Ij8Mdjs1wFB5grNSE/TaG/sMFVwPIlqSedpqbUGhjOuWum6sPqevEFgOBbREdMEfg
mGbQbfKa3jcDgxxNpOFO6aectZAtfG7sOxvVBrc8UuiW7jbqLyiB2RjAySiJ4SpM0hi9fCXJxiYQ
0OY8Yi9i82Ee7eNr/h+zCbP3rhlqeaQPDEpGa70m+ATNWCK0T2H11TiUJsMjcR+nZa/ZM/zBe6PF
yXIFWxwaqG+Gkz2NMLQ4eFUzqAMYrMi0f0mZvr4+efPpOB8T7+p8PztmB8Dlz7S3JZz+u5jtUNJi
kAJeJVcoeZBD6Fn6DeEWqK78OsYWfHOUys+oVx/DNMuX3OKJkygLKSCTwnQg+lXTaIZaO5MzpLJJ
NsnOgseAlwJKYSsk6cN00oKK8EluBA+01Bgl5+YqED8ZCP1coOwkW50GjXrmwwJxaENEhZtqunhZ
CCaICyNpnbKn3rwBmE4EbAUfkOCff+n+mjkcXmkLMwWpE+s4mcGy6KfPummpxGAKfU5r/D5oXa2u
qXWnCx0pTfU3HFHTxPBxk1vSNSowA7jTRHmpWoMAhAQXt5V9GDcaYBSlFmbr9maQ2qkhkAJ5Hydo
6wS5jVRZl5zbHAeqvhztqxRJRd9mA/ZDMFasHt8RKkUdw76SI52CFWphYLeJ1jpeTPIqOFrnyuLU
iR0Igi0OwncyxFWBkbsMAkhOamTXdC0S3CX7BPjusy8PPBnIqYzuUEOJwASFltJ/EHIBOBiC82Ne
Dw2/a69+r5PSz9Yj873w8SYQrxsnA2HCyBTk0T+AX1oaZvITlW0pXV5/9d3HyqfeIapVc27imVr2
xwiBUyFw9THF6cvb55kn1nZIS82cYCHIZAyJkId7XuzD3BcgjNvZjdgbK/0ZgADhMNtrl9h8Fj6+
PCZ4hsgNOh551xyzM3/O0x2CcBi36gjSJPF1ktM6S1E07UxIHDsUwuwiXM8So2HJI591sz3a33YI
VGmmNYD9rL7NBNUkN08l+JUtAshSLDh0mRkDAU8Pcn3722tz7oFobSFQhWCts6KdlTSxuQEv+nLb
k504SNgHvr1ZbgaEFsIHshpgJ7v0JZ8v6ooXPPusztmpRMnGl2irCle2soQC+ccCltA+/QGekvk3
53B0Dojxut3I4oqrIDIqVJwpPRw/eDxjNd4zuj/X91PAuJf8lfh/WpESVVjZOs0bCXzeRPlLBUYK
OqSouV1fN9si94RMkL1hR49zqry8BbixZzDzVNyZRwpXkC0lrGk5ix8XwCDNGTObcNNfw0ylBhBC
FcI3Km0oICIzhu95Y97oJoWRmgGZuqjs/abN6PZ7YsN1+tP++YL1J0bXVEo0V/m1dM5QqflQw6WW
5pwU7R8IcdK7voOC5jYR1oxPRGSovF5sCUh4sDz4gkv0O4rNSqW6K65C6Uw6UkXymB/3+voGtSxD
CO+niqfr+K+i5/9QjCcQVVU/4MZNbNSx6yugxt8vj4L8t+epd0ocAY3xVZ4MtDsgMYDkc5lxwLb6
pJS51p2OzoWOnNVXIO8K9XCHQUvv5NF+1DgrZUzjCl8tv4X/baBpexW+obZaUfn8aHzGnijPjnLi
iv6MSN2cznIY3pbuOAZnZ8EEr5qfP/31ZEVNmnrDjakZz9EreYal+BJY/f2ykFn3Zo1oHHyqthHO
TzSijTSSMvBEc0I3MaSA997kK2kS7Q5tXedzkwWzpxVR+KTxpaBFdJEXB6erm0v9rcewm9X0jiBD
jYjUdq1FB3q6t7o0rWCfhv9BeqZ8gVVXy5uk6+YS0X8zGDNbL8XXsvz/IJixyEDUUvrnyszxL26V
yUsOntkKBUrpesVIHiTfGDO2OkyPJ++B3kg5Ki5tCEgBnq3X8zUd4/ZQtGO5yGzBKkQ8pLnhOeJz
5rdeBhzDkQEXK4evn4F8T4PcdCgp2ApAbcx3QoEs6QHp49PHqCzcyQJkJ6tf1XMqn+412/bxSCVS
a5cyq9eCnkiss/AB+aaK/4FzAexXBYpL22eV/gM26zLt0DJpeK6vYlzzmXBy7P3MFCreSqEEXDuX
gHvyUew3M9T6zDydycnc+J1csm+JUkOJZ981AAi2EqOgL+D6qRO9mb9Y45mG4QhV4tDowrSuiEWD
8fQslfEj2QntKw61gPDalgWtD9Desx5hiYXpqYFFqXWJoZd+o0I6O5NVf7kiOUfeDtaIvHiIGqEF
/uZVeUfs5FNMCBBR9aZva5jlH8CcjO31wjTvxRoG7oM32ZaVjp7ZLYRKSuSHCEKThX8y1v6JWOZP
mxjgjUP6QUsOeCdXuONmAJtye/RY+mfk8Vrmp7awOstbQqjn88mGipoS/eH2Obh7RuCusOY74YZg
evJknBB5wqtdi0wgVHY7PNbkfGR1DgorRqaJl1IZnWd4eewffQjkEX2H2q4aDXauWmcPonKHjTlj
f96RtiXKU2pDjNa7lqYKGhZ6zmJn4EfdwSrJJWMoLkE0hQHm0a7Pc6Pk4N3o0JgDT+4+eulEI7iS
Tq8bNpSQxy6sH5f64/tbsH0SjJ928KfNtmwJyVt8mpaPCKhs4YpEfCGkq8Oyu3nCaCxkcMDpFmSB
8VB14MUk4T+kHg8vADhhZct9lW8I5Up8AQTBX/jltBdCEBs80U57b/u1+j7dEZXJ++qjzDzyxTpt
LzjIG8lOyEqnC6nkMBusF+rVyHMtN09mODcsEy5F7DNp9fr/kiEMMh5i8PqVwFkfcIj3VMd7cDTK
jpFlOVPKPSJuuGHx1WVClTPOOgs1EicCZ8QkgBW1lOD3Ex7ZxEFXITP9mMLiNaafGeQUuGF/rXMM
yfNPsC5tgbtIwJaFtk9qpPJOX9bd6CI70lsRtdotlS4bjdYla9r/uFVupEabxOHTEfWr7xP0f9n9
fhy3Jf1doPM8rFfpzx369BJd2E4q9Gjiw6zTw+UiZewdXGsD+SP54qx9muttuvPkNITrtGDVBfXk
kwVj3KfGlI8jiIUVrXGwg4Z9EjD9f2j5d3IKmKiAf/KkUv8d5PTGhake643kKqUzTppjBc0yH4SF
M1fXCH892o8pH0lMgXZZcgPRTSY2NkBhMAI8APqWs8HybrpS6bekzdw3yd1i4mgFPb/3W4x6DoSB
yhAwWJ1IbIInA/Lmvx4N/1oKPtUwIRFE7bU/SQfxCLJPjFxhaFpGm4+u4kmvqdqldFKtMRcVNQ69
Llr/Qjn4XjsBquViEqzyuY09V8o2T66M2GP859eenljtxPhdW5vEUULMAg04OnljoXfisxib58Ul
ORD1tzhWKbszDZ9BlbnpZSdla8DhZd8f3yqrM8NI6Jl+yds2LUgk4vFXBlMyIIvOvsJ3TWB4aCM4
1LX1Jqmsg0Xw4dTH8xxQC/p7e2SQS3sv4Kd+GxxuMRzk7JZ9FBoAkGnBirweexq2gQMhNrvDZfg5
/cvDfe0lP9frKSRcXvBusTsq2tIb41zeGVkbFU/JyGOB0dkfRRaOwfZc4ruAWADAdY04JZoRzxI/
Rwl52Uz+m0cAWXnkiSMCftJdd1vPpUexLa9HiGM3t0TUveiSRnHShL/s+U8Nbzw/1hz7Ga1PVJgV
D2NIvUtCDHVVPc+II4P4o3DfM6jmLjMN/FqydZfKc9hsChVW5+/uw5O9nbH20RDjwh6z4XBq/opV
P6Fj60eCdjAM2wwJFTGE5FJ2hYqXaGSoIrGzW7zqy+jhyUxD3D4E8Rbtc/n5GwU6zZchZL+eS/l3
iljMyArjn6jiMZjra9br0lUI5eqyjVw4MDkik1oBdU8Q5THbk+x/2PqeuvH6KLFQBQeZbCkKOZC9
b3ey+mk7arSypEQigYNXod3APso3Gr398sYsI71LvblodrTJkEvjNMjp22D5yuDl7QjTBdf6yyQp
jxH6soNmvDydNsarBZnk0jAyOWA04vsWijnPZvc6UaP0BTFjnQWlrYCTkUk/ANi61KekV6YGtmxq
GaGaVsCwW5ERR0++y3K3gt45q4HR80BoCoif29td/Cx0WD4E4jL58PS/KnOCUI9W85JHHIta+Goz
/QOUVkSekLB2bVALO7CglxnTUPMzye1wTkk0OjXdjSF2+Qwk7sEUw8LYU06ytbHYPjs1Z2r3zZy8
J6Bc67SQCSQv/K56BkzMN7fFElsIi35Sw4sCGUWxs6brnoMOLZXbiEc/KasZ3tSHswtQLsKcoU2U
v6danjiJG8rlSNsWbrgdU/DDkKHwLem68yNYp/uTsjGQgb64giLgoLYfzCgIL3fmZYdjK1xajtvk
k8dMexyfOodLNLpSrTEbgz3lU96KX+eag0jo4i2w5/PfNMaGBNYHN8OnRu+TNxMZe0lKo9cap6iX
C6oIhrvP8mKE3RjQ7+CJCZHRG+9wQmiOV7LIRQsfoycYh8vGTDRq/XAVQAgPvE/K3e5NfjdzdO9D
wbMgsUzd1IclVuMmA1Ke+LaVCjgFAClCQq25huAhnKrJC9+/BFEQt5DTgCIirKwq2SRFOxQJAhFC
hLCGfPs/eD1x3RxYbOBvAXunPuyD9ZRMbjeBdlN0XrwGSc23HagsNy49WXyLlcDnYgtZdH2INY4o
4g3glV/Xju4SbBKqwhXV2PsQdi6lW95uKCu1qJb2qlUNpnE+KXH9GRLJpsdGHMOQhSBy+TUkfK9K
7NSZ0KIfgEkwTIslvxlwaOV5UInBYGFiLCgLO7byiUJKH1GhNU0h7oWrYWwxJM2iGUxhtZ3Q1jL5
VHHvMtJz5PboKcDGsg0N7632JL/amHDoOcvGqg463YPElevfHdWQttnMpclgyBoiFE9bdFfKfWd6
EPIABEBZDK59Kcn2pbLQGyMlCQglEf+RQbxhgLPINWdoXUh8n/FHm662z+atPjBpTa+DPCAP2k2Y
O2/lADC180/HzSXeS2Mbub0tZd9Ckc/QJoQ0tog6Z2p/LVZXCVYyMvx6LelWnsAKxNNfyIM56Zbm
IcBSs0aKBfccdXq42R5Lcd1EWcfyNXphSgMEOzZs50jKRDSmXAVFwtIzN4oi2ZZoBKaZxB1fvdx7
06w5+QAIJOdGEX9787mPWu1nANkEUnLqVTBejDfoNdOTxG4w9hB8P4H7sshsf7wZ9pkHgjfVNRnd
PeryQd7fMykSqhmvBykuM9pDC1h/7cuQ2L99AlguhUPVYhwBIG/GP72/TenO+n1CxG+SMRKKrfBI
bs8t+jDDOkeHJW4dhK5Jfz0ygq1hk3nr13gOQYfvP9C9znY6xScXlbQiWJIEj1nDDPIDKHqjDWhc
zXOQ5h1RXtA9hKFGEiNUWaY9VtGGwc2LZ8bogC16zPHXQcllUcQL3SAZugkABbDqmrNkC3p+Xpox
aPeRV/7yftmjT+u4BtTqMBrXLBa+9XAn+QaYt0uTA3XTX4F7A7MipwJ5CFtRufh8a/KlRamb6rRk
pW5jJGDCajimaARQi4rXZOMEuiKTGdQwkBhAp40ZPMovDu+xNP3eXRvOoJR62unmwQ0uT30nNcVJ
qVKai1ogrQ3B1PAjh9hFSGphbQqujLVdn8yLyiC2pqjR9H6FyCDL22ZC80d7rwnxsuOxZ9I1zjL6
NLJT7sYukKKYE5xgO7+/vFgAhMhnk5fMju38pXwPoMUr3hQvaofpksJy2memtn3XZS2HorHJdKHf
IRytEUlMUOH4m+ilU9uI8rC9y9zbdX9omeU76Mya5NJa2Cqh4sqcqUWJioxq5bTu7rt32RFSL+g4
gjxTQo/t7Kd04Ok8nAtmJMsZrC8LEz+z7+Ggs9J50Ve9V5Vt0OhbgAP4M8dxyV43pPAB0HRUzKbt
TWfJfsWJniVvi6wbY538fHr8P5cbRDSwvK9M8slTyamjkfuoYPDGClSUAMBpTP3phJJmDJwxoZFI
ams+J+9ha/qJYWTkf7COVanwaxI76GVaF+cnfqHsCB+Dxpt2pHhmnhF7I20AuxCT35BMUimIdXVn
gHStYd4PWoJJMLuYVLI063LU5qNxb2JQimrss0xfkWQABnjL0YCIYmgsN6Wxa/GdK8swmp9tK7/9
xK1t5nlcKaXeadBL2Po8EGC512t56MGxDyKv1cNwp5Vhzty6+HpMT0A7Y6zEJAi/AjqKR80e9/JT
JxGa2U2hCWOgLYOZsSmnKpE2yZBHDiUcCr2qEoJdcQwKiHcRFYYlzFmcy5NLC9U8zCaA+FClxG5a
b3BaqmtqizEMt1cI/J0MJMngsJjItdq4LkDM2MK+JXO+v9ewYwqIKHNVvu8GPMcfTZOYve6BD7n/
Ayzwy15rskXV+UuaGLsY+AvAJXUobmm3yy+yM2qLjnRSvhdZYRgOKIDwaDN9wIyP1Xxo7nnIkP4q
qSVo5RieumKqsaVMBm2GdeBoAsMOvlIRdA1oSaWqJqJVfAle3c/nNlXB36nOtuUj6FbovhKXOUHE
ffdrBaNn8AGq8mDKKdjJmlWo5cc5viT5RyNZ/C4IpoBbsrj7KwNtcooYst6SYlh58ONF3MONt3ht
Wm7dWUEz+q0mDJ6Ox6VLPo1miRjuBXxXaOFFqLNGEnGY1I/dd2kL7oUtR6x2nlF0b/jYkXKn93Ty
EhVSdeC4a81aSl8Cmvltvx9mG1ZBe0MZA7qsjz+Qe9XHrNhKhwAC62RnnRQtmrWMtAyueaNkcdG6
feef9sKIdkjIbo3bX7qSeemFivlZ6PJHTwCromE3TxwpM4FNunNSyBE1GYw5NCkDkJ12qVBn0Ufb
JjxXmhV+bRm5ICc2LuTVqoi25wK17sOeQOUPVVbBebomC9Ll4XHp4DQgGoYoXTvrhz5qAA3MnkLe
ueUWurDNEWh/Ho7K+aC+yvgdCrz9/wx8d/9lOHuIF9910RMxo3nDAVLYR79QSmwpnDl4fCDe4E2+
o2ond2ado1WQ1J8Ub6Z8aHose5H3vYeQY8OWl6wFvoN4gAdRLNZb02T8r18F85XSOpoch6BEbXNL
dKgnS2TzjqaTMCZ61bvVwyXb8dNd5gx60FvstBUOabHRldkK6RfI4pOc7qTDf9zhhatFXZum8UPo
gWBChefK3B5OKjiY9QNK9M41sG3l8lIEHdJEItl27rlEUGV8yjTad6r+qn9GKfnKzvUG2NyxQ2PR
o55m753IVV9IjdGSnGYqNhdeyEv+uZ8FG2ETvu7cHrfCwpAvA4ciDPHxLC3AJrY+edjBC0nXEB4S
HcCDym0iehWV4eG1f8g06wgDmdX5C78QV4V1iszQyljbvW6/zEYgLBz1C9P2uTMWvWvpg9H8jmWi
JY0dPYvQnKL+moLi1lLoLVfGz5IcfB4AnSIzuGaZeEjZgsKbNbaMAGU5Qqk+V7v9A7rrbbSZScXd
p0daooYL7iDhY4YJ+aHnR5ZNOQ1sYUs/LIb4vD3hoQUbsPcsqBMlm/u0DzEpRtO7v+C0kJEezEqG
7wYsxfDleiDMYW40C2J550xix8VlfYEtUU4y1HuUajtWM31jQK1UriKscuylYTIgPu5DkMCBI7P3
ZUfzzGz85ffICtEMi97aht8HkZToMMl3jd5q2INy8/rpyFKPClM3Q5QMkWI4bvSxlhKcoUREipTo
wG3IIF+/IJCDZ7uSksNcTcuiJuDVYck8/Mr8XAoasd16ulm9Y7N6V8urSv3ihrwWVgKuWDxK0Xdv
DHHjCVzT6AJiDBoaeRQcuSxO9exKa3imC+hx8u92dYQa7tRcfdl+iYi6pidDbIsP5DpxhMudH0Mn
l4uPOcWqy53E4PFO4dBcKD67wjD0GZB3js/gOa//j603jMa8iEyBZBc0vGUHd04++3D3Ss1nZzyp
0oqXV8G0XWu2d8NgSKAztiHNOzEt4NLVXQ56QBPkRmY7PnXzK2rPtsC6FIb7j6s2T8VeUgXYtUxQ
OY4ZAuwa4fL/pRjSqdqgfbcgVqFNqKbgcbXT9nK+aUB/CJsPhJWSi+cPEcWs93WngmI5Igw7OS5T
/GdtBYGZ712gLhcFOYxS+R/B+xp5fsNxsJG34JtYuIv992jARM6a6Equ+jYyHVQ4PuGReCq7Jc2B
2ixIwy+GjStVR1bBopaOJPsEqtxk60gLnQddnjMdyRgGDX5mDm/8YRqhJRNV+8IC5qNnrDEk4dtQ
vNkzYXwrEIfvx5/SQ4m8nNuDzc9vjbMbZFomQJuXL/IDHvXc+pcQ6fuktKXhdx3Kuc90gA24mt1O
ivrahHXgkFASgYv9LE+jdpozCrnxDksfwLZ2D53H+F4DhFhphsnN4WmIZ8KoKP/k2rAFIJworHXk
dsnf31fmkeP7AoFUHFa3dfv5a7BZrGxX+RHaoaFm5QxLwLzIBw6YI2sQWl+Xss0ABn4dQUhqBFhE
+OvUHEldjbANyb001CxghizW8lMp2zqGqbZxw8rDo4WeitgmpD3JLOxpXyaYmMe26Wg2665AxOej
LU7xhB30i3mCOf/Va3JEuuXfmq88WQoWk0A8szb0f00hhOZHmy6MeenYlyEp6q6M9pOSkhf+0qMu
kOl4ACo6615t8QnBXT3W8rXLNOFJ4kl+AKCVQeemoYOUhw8la/ZAw6dg2/HXbDVC5vsVaMPUH0rb
0bGWHDF6K04FTyDfiOuD9w2JGRjdvH+O2dTPmrE4X5ZxUsSCj/F45LUBBM+VfDGKMgm6EXrN2oK6
vE7iWGU+GLJsAoAkMclfPprRVw+1YZzKZykS+QMQnUgzPaCZrVyCalAJDoARUhC+qzul/GuldY/0
QBnEE2IlCG8RP9Bik5vhS0EdfS+kHEfplIXC1ZAwN2Xmf+J5zyyJhwF9Vd8fnNqry3g52H+fwv+9
rty6TwRfmeMz9f76nxG6cAZdhRJFTYiud8DPUiN4aTXyNuU4kqo2m+HxLd/rgKVPunnliic8VA3n
/XNkib38XoTJuOr2sO8jVfhg4twOAWfuAeTfyKap2HcQt/nb4reyrOvulUmFZqdNgO+Ook+ZLe+M
ykoSkMEZk0cizYHtq9ixdxzZEgRUirTIn9ffvWCwAQGqOO1Soxs3OvC2rxhSAsU08WreDqbst3kY
DQ/WBGGKWKv+9cIHvdK5rf551Ha2ecvwF3h31ZqeNpNxMfHSi5lSuOSnrQ9TlHzTguOJbNRO46py
AJyZXT2hxrkguCDZZdj8fZaFcRqZ6Ljz86Z1EUBntbc/Und0sAHzl/dNLAuMRK4biO2tygh2+bnx
oj63GzlZ2A4sthTRl8vn5jYAOn2kgYvc7qhCriDEaZfh/Vr6cp4PqUqoOzPZPD7GONbFLDsg7ZE3
Iphfg3mDPJEemWInpwjtJPnvlfW+Aw+hOodrtwNno1oEAmQHQTsMTYEqEZvCafp79B2mpijEyim7
0EIQRnwL7SrVNDTIe5vt8QCYy5L1ayIma0Z06xORAl0Mer741FmWl/4FGYkffh+AzUK1TtYAD/cx
6MqQmbSE7vIvE1e7+0cShx8C5p5r+B6JDY0RyraMK++DJ7UM8BE/aj6JSorfuz1fajalu/fW4Lg0
Q0cLx1b4QQ8rjYecB41f5ERf+gkOJ4wg99tVKDEjAoa+ic5NW9bPobjB7uSSlC0Oy5dBanmtl8C4
cAgAdZ7G7jwqucbA3pABy1f9iOZ4vXVwkxYn305DsyMUcKb9GEtWikmZ8I4e+EjWlPawhjawfBmu
f2ydEYFyUDRIqq8GTy5wuBkcvPUkWEgEa982VQR4/bGs7h0o/thkuz9u5+zDd0rJp5Tk2QY4YSAI
yzBiOosjrK8Rcdku+p/XO8VHA/sIBg0qr1ll9QmKBfa6rZ40nDhiMRLByar5rqr7EqU6ZwzdtwNv
/vwTKr89lcrS2drBrNfGTE0RlaJwans3sXbUPEZiZjEIz+lQF3lxfVFv5DBTKP+aigJ4IN+Y0REi
KkA6N4Y0DdPTpEVcWjKSCdnP2qobHs+GkSUxuDvVK5qhfFSsw35i1lrrmlr+G1tisFiWhEsjUbNR
Rhtxh5MAz7BhCJ46JYCKreftoJCFIJGQS/C/161YgNFPwE7fiWO2lmSPxPbIO2tksa5AaK9EQnSN
TnIeV2+H3+KULBIf+2ROEDcamI7x4IqCQWmlHDj5GLIN2oiOjWaNUq41jerEzaicQ+vRAUe2P5M2
wySFyHKxaU8DI5YMJQC5vpeKi51EwtozPB3UsSiU6mhTz0poDPh39X1kD/QQovUlU5jTyxccy7ud
aupxMuytpnhOvGNnxjaLXHkgd8vcvk5ZJCGzWmojeZCIG7KXgIzvQGIO3208n453R5cXQrStngCr
Cot/Z0mAu8qGl3zKYHhDyxwEBXY1mciu9JByGrumjvgdF3zRjH6j8ejwMlJ13JQdY5IwoqTzflqU
11aURaF15NoDd7CIgej9ayL0B/q1Y8YUxbfU+GTdkLX4D8cSDQ0Fg94XznhYyPDJJFGU60BHAhyT
yOBfcRXPnEnmnZvXIUa9Kl5y21zs2u82+flk/SddVOCLLoP4AY95OXgj/tIIDKPVjgffxTaUIRZk
ckzryTP645L7xNVjymnD4iGNvtpDDh00XYVngZojDJOf2sHtkUrOKbxsRAB1Sd/zLTKY/xXOF+PV
BPV+PMN0zOLuec8OJyALz73yDaKjVDtZ9yRWTQJK6A6Bj0yxXxoMYO8Wro6nwGd/5uR64CXMkrk1
18aCSmAse78wyUeeYRiCF4q8surC0VkkH/296ghRev0BYqjpJXW1d4A0IuOortzPFAN8fsOYfajq
mbfA8978qbg13lCetNyjap1LjZb/8OLXnwtzEFifLcCLW+GX43wcn5+fqUJm4LswINgx47J2XtFu
S6rUIWbQVE3ygK6dvYPR2b8bZTo9YqaVBSS+Vs0GpQb4kITCTyF38mVuQ78f3AuJcr6X32jPjz4m
Kl7MsE7bUyjXOjwIBGnQc7r4ncQP0nim+n5yFVQrjJqveHYyb5j/c4gIVgF6OIQjrmdPw0p6gOiP
ZnaQ4mR4su4MksvWFr8Yz/NohQ2d3NGmqRJtHFuIxEkPy7+CNzN6NXUfBLmlBQn/5Ua0Lyib6Cz2
dFD3tWYCei2NFisMz1H0ieagxierGfxbScvtdwKZVIFxKI0rHVcafb8c+sukA6eguIkhgBnLfbOS
k6kA6tw7/dAqtNTZWi3sW01Xc19oDeUB5GK77fiJh+8Y1bi1hs2GtGr9DS58QUEMFj87DGDv9tQO
fTCDbWrhCSGU9OrT1KRYU/cV09UOVZMtpKmBOFtfVcRQNnGEppE3f8WkT0fD1xjhhYZwu0/RUPoL
sRhJdGD/LOiazBwegt6HOllGfqTiR7/ZGYjkgDHC7HZgengBdfvcJakvDq1v/lhzju46+6u3ZSmZ
2OWfxCQ4S1UsLeEuITORq2oNHJXF2cn02mio356y0UV+vGrZmcaVzM1gPSW7Ca83sPH5dVtY/1XS
G6cmEtDVxMK6eKJgQna4CceJBzkz+0C7rTO6dE4sMM1SLkhUw5MtFH9C8Uq1QNNBpk2iJcgDugiw
eM+OFUSTcRmwjQ/UvZoZ428Eww5yQKywaOAZXvBSpAVxnJw1JZROj2SF8yGkYTAZrFXvW5rXacgi
etNUZ58l+PJ8TyUB4b0VFBGlrr+OMd1WFSki+fujKvhF/yVIbc+CpqZYpsu7eGRknL4m3VVl+c+m
vO/I+eTdG5gRLNWbm/yLzClc2vPME4GOEMdmCdfCArS/Dnh9QddLTxwRxICmGV6tJfRQXfuTlG9W
q1BPJemazl2rWzcchfB8uHm34ihqYA8Uj/Mn4C/RLvzjd7SxynEzWWcWQm8d4LrpsAIs7irIzoBs
1tKFNLVbely34H2tQGToybNj9c41kLAcL8jpzwZd6kVbbLxiZqb0OeMs9JkVQmY7ul+oTl9bNrnM
05UukpRHwWVuRRr0rg449RD1NMJEEmOumtKawIQxlQydhb2uKlXrjuAjIUVk6OKLNmvmt33IPab1
z/WjVBBcR7MNe3tmndA5uw+/VTr4BZG7mhOAU1dteluxlVCKowu83IpGMQ9SvtKyQll56aFWowE+
RnZcbxYTs1Lh0l51HZHy4/lQmzcjMKkASoAEKrE5l7hMrqLEGbGpJkjCE42aRBi2BmWBg+ITaC3x
fx0hZcDYHa61FFOpftpdZis0Z/0LEE38w/TST+MdF01IwMzilftqBT1iVuaoaZ+4J9VTahBfLx7h
/PbCcsFRClhruYGjOs13DW/ql2vtCVJcl9MdULtsOkm5h8d3D3SNpA8bDIYVwbLRWdN3wvMImPQK
3rVLUCntDYeigHa2M12QIaEzTOKGXfis/tefRiEEyJX4OIo2/aTQSxUqL2AQRkG9SNezgltOH7Ea
8Aw0QgRHYvY6B+s+QsDoTVxjJzrvQxyUaJInWO7mWAZ8CCPnGbcnO7qqGXV1UJjqG/PRDcuEAw88
x7epfipyEMubhPEz/yNVWuyRPsIyKlei1/TjerIl+8b9AQtywoKPioSZ2W2yFN1kzzLJB4r92bz0
UplTScu+NJKcjkpOwvwMCWQ5i0tug5I5vIkTpPZDg8jGzqg4w0rnIWmrzMuDQKI2hu9YFjehkE2R
BwSPD96fWSmUAdiVY6wbER8sYgJSg3x9SI8mBlGeIMzAetJkOkV3tHcseDW/ospy2OkCHhMcOWQD
2XkTA39nsSkTNqGkDMVKcjn9lw3575M5+DoSLC37X8zqhB3BeMcP2QSOIdjRqynvDaSRYyK7F4Mc
4SNzI49jvBTUAtYo/oBwGzdsIitxOQj0oVLfofspdnLG63zBEdPzEQ28OaaLZZ2T+kJqmlU+J/nf
xuzYf/g/qLJWgB/XWKXZE5/Q8U9I3QKpEKQPVGNEwOYiA4HoxpLzCJGu0lJJZEkxiPPqgl0IIbQb
QohGyIbpfFW+BJVAh79n++nQ83YFq1UwqPVXF9lwx6GHQs2UVgDMXvZEWlglP12YiJ8JNV2tGYuP
L/SulVKX8FJY1Bhi9a3r3GX9O45ssC2W9HH2PXJMNWUb1q520tsAk4JI/0miW8i+6Cw+LwICZA3j
LqXcP8AQtJUF+n+WR4fpqj124agaNZsCaD4BEvf455IqM1CIjvCNmih/HeY0io6b1GbbZLC8s6cF
0Niq+YyvMwbYRKMsZQKyPjP50mmIsqhjQpR9kRDJjmmxOlnqOAExEY12h0RF8qqIjFmPcGIBXE1A
fDTop4bu45cJg9f6csOcR4Y36k165ZJcFd7NtIlPl2a7KtkBr/rLg38H0SuI1tRtHtV1kgPJEXbH
dtEZdU+/wVXBrwOPxvSYhnEc+gnJ2JBtj3xI4QeBKCKIvFr0Nh9PR6c4grpatPsBtj2sPoK+NksG
0r9pkwUormGHgPAHzFVSeYx2g1SlmHBRdgO+5pzT6yL3WBc4c+JGFT4TOXi6Yd3pTTOmEtVjRiuz
1zWI9ZU0vHM7fAh25xJKmYNRNR7oqrknkQezT1VLSF1TQDyLGDO9tBhjWNoQvxvRiSfJOaRX51QW
gGX6zu8eGBeprqnZRh0d78LUwkYkOh3yf4azmtVoDh6ujLqQfH+G9YfYhNV8yssr6jfzAR1dOAkm
TaX1wpSqZb0pQwZ89XajIlVRJ9iWumN2IkpNEEoGlYNagkb35rqhTCMjQYiwZu6Xr9LVNT7TLwj2
9sjYFimhr7LvL6x1ME1yRgc6HmhoVncDQjcFwoIW+ZgBx+6R0SyV+7/jJLfmt7/ozTwgzZBUVZPy
N6qITT2saDlDiAWjrEvbw1Ck5s7G/wibmMtUOe8EYeV+bNYwM685CEsnK7GyOo544Li4NPtaEyfB
6s42zYwpmxOziruxtxiuYGU+6IVSUUlOPPG9a06TMkz0RqyfPuJRu7kZkGcIiJqPNjl+PfKIbYx1
neIeXziqjfKA1fPw84gStSIaZqRzXamokEziNTm7BKzdSnaCPmZZAQoYHdMS0ed7wyUq1CGIvivR
jhXnDNezDQdh5u4BHtjJvBneyj30xLJ9TZbf7Cm/K9XP8aOOu0mBWaUqspruyHU3s55OSXi+9DLG
U/MAEKlz4mRsKY8gVDqco8xmze34XRRAaN5wFxKLboLvkNs6L1lkYjHcglzD/Wn0lqk8UDCoGluP
DHYO1Dm0Bsiy7EZF9mpnlz4SKDo0q29leyS1dBqwHH89+ZGEfwwn9lt4ATfIB2XSzOHIaPN8DF4O
kjieriNRB6iBFr1uXlD0tmOzc7SuTQlllB1tvkvbOmCrXUMoNqTUuxYmAd5Fy8OS1gLdtz9IgJGM
98iFRE8MyPxHkv0LCPBd1+qlAZSZaf5k6muv+mftyLwwXwbSaucEVZmdAmtnsBNINgS26LQb98e4
hQrcmWnaL2CaVCVjOcD0KqAv3YAyW5IYZFPizxLxCOQfnnXWNVX6psDqirbi7tKVpe5wpdeCRnE5
CIls66VIBwwgewNQLwY79k90ARKcZyYHz3MdaHHvzrD8p+HaQ3rrSl+QS03J6aXH6LQaTI+eZVdQ
09bomLD40Wbt9Lp5uWKCkJv9iQ94uUfBIAKwL9sGfPHWlnaIHedfolHc70hqwL/adIPt0FY4BMaV
CbzY7WDJJfODgSF8lLSm0auGHBsmKs3WKHq+M4alD5uEqgOmX+zQuI3ugQwo0v7o+kxRFzJXdTsZ
iHiiPWx27k21Atlg8RbpEdpsr04rGyLry2Lbc5T1BYR8hGAj7QZk7JFcEO5gBNzCKkcoiBuZzkbB
APu69dPoA3tDLdk+NAZ/LOuE4dTa8FKml3X+C46eqh0T0mwvtu69FLKI0pUFkFlQusQ9qhUkTvM5
f1mtCKZSJxTFlHuEmTvqLZ4906rS6gskoCx+7ElGFqfgrc0rwJKkJKyMUgJu4WC48ceSLJYN1Ng9
8FRIcIN3C0xDMBA0ezM2vAoLBbsQW7Jh/HjU6eW+PJUVYtsx9F+lmWbcvs8BL3tjrjxY0gCyMbpZ
Tiu4fjfESRj5jhiDySjNpnxjye0jzr0koxybLpaTqssZKB8NSHsyEKsYsO998nDbjgRSrhHmjvdk
2UuWGB7H3+TYLqkvYAScg0IvN3VMsLgyGrO11tlUQL6lrUhN/pYLxLwRfybO1lhFE/86I1/5Ecxu
mFFTNCR1v5kXAfzDePIxxkagjZiBU4x47p5fXE+CPwQ494yzfDbUmZ7r10pu9+djumvWvNsH3lB3
TZPRkNuS3oUEV5SYDogC5CduKm6ImuG1nWn6oJJhjFom0cuH/JMHpTMQ+66hb3S6i8F5b4EmIxme
CZf8/h8j3mFf0Fg8OrIOCUTnuGvaDVlF6rgmLnLxRvHyTW6//FizdhmI7yW7P5ahiQt1Tv2zkaZZ
pi2iWp0vAVtd5AQ/0ycnu+/SlO4p/8dnVeFqTY9KVu4w0tNrZENlj5Qd/mIm9IuhGzHWCLdBQxXb
EgTdw/f+XHGaSj4gUdyqMPFHz9VI359mWhyVxRL75p3zeWKhoSv3N8Ye5jjPYJG0gt3PCZr5gxNR
Q2vy2GiT1f89EriGoT+lraZlAl/XM7IivbkMgo/dvG5WcxHE9nSql3/g/eNnPFTp/uFw4M2JqBbm
Pkrw9/3upaXbBCdftylXf5GF5cDwExBqFQrw3Fp5F3SM40SoIYN1zlCw2jreXdkTOvu86n0IE/R0
JRjnTY3OiJQVI8pLUZ0pABiZreTnFM4Du9BLaVfr9HY6OBFcGUg7b0TlSt74YaNBkbZnjLP2pQJf
HAEmjwJuC7d3vvdViGno1BTswEE/Nv29KdEdbYPv481mNWCLP9OIXFmwwBQSIvyfwkv07DGlCmEJ
+5UpU+HVTSlITUoS10F6FQBR1BeNOkvwgkSkTBxtw3W5frr+XNIwV3Gty3Ykkac6lAKpRjFcd8Ii
tNgVRqmLnJ47aNRke1l/K8HwHElGi7GjHUFr1HVIAWqSjKTHwk+Ks38aDz2J8Ay4UCF75cOetrFZ
4m4D92RvPmSxGRjPgOM3zG1V0dS0nkcLRmT6u4KjuC5wIlLdgxVmqIJoqsWplSCTeiGqMZqiYVJ3
680xjwJjR3dvmgWqqNDdq0WkUAHhh2+P+NVWCEyDqfDvpe47ewkyVprVuMVrKeKbRF5LFeDppjYx
cxJGFWiLMa7OkD18ouL6uUKB/hbr43GDP0umQZo0ZYAzC5Fj9+1QNWrV4Enmh9aT4h/CwIjcj58s
1+hGzY5jTqOWZjF5Ks6hNRvZGFYMDXcwYeEWqretkwMkcn3H3Lbi+xFe/Z9wkJMHsDYW665zFlZC
Mdzm5JG9vXkSAP+iCNRxvBWdGIyRGyiVvTy6FX67AJZOYuwFb60cfXtzhcx6sNUTRruG90z/wWBH
UnVBSbX7A1btqnVgUG6mWKyokcdyJgwB1lAd2eVCMsDdh9YUDbWWkE1rkcBUsDRy/5TA7Lmu9UlI
bi5T/3KycS1zBirMb5V6pDXNFo5p8SX55HAfXa6ubBBxLju0KVsi80v0n5DmxthkEOeiYRFA/TrD
X6fLnrO3ELHZD4qqB8MY7q3K4MpvIwUbxUh0CgwUnDVS6GF2Jtc/fWIlhRdDDe+Jewz6+wpxpkvK
/tz1ExaH+Ms6ZsrFPlvcXOC95cyKlmiLkB/VLzFTXOIvcnq4bWNmG3Rm3u4Vq2bxXmzlgGxuAnoz
X+3+Ag0PAulhFmrJKAN7ow7MiR1aLeP/bsmD7oFP/Iai392mjruMJcZ/wWdt3jzAERVW5+q0mqBD
RqwaFOo0lpiBfee8hHp1gnltcl3+AaTK+6+gb0M21PbychCMR69LcU5PqmNPKxdPS+wW8RvnjKk8
+eRRdTBd9kxgkS6/hGM/5xiuc2qC56IaZflBBeX0dLL8mp9KjgE9QmVphJyr5dROFr0p7Y6N3SME
fNF8ywP2g6kiQ3cxYnto5hO2eBW1jq6uTKrD44myApxaYyxFalcAPNU4j6mnAIs34UYcPNWJH7cP
Sw6Blvzl2tELds/VDC+gl9wB42YOoKDkzO6qzeufC3qQqeuj/cUuIeYJ0ClkWKkboSjm4KHtxPtN
ywCrRMn7NbalibMsBZLz6siiR0x9Te7fIqo+WE0DKml6pnLX+iZtqx+PaK8coAKyxJ7lKK6S6uAG
xm85Jqk83UBDVYYpYL8fgePc3L74+4z/57ullMMm2XiTSbZwBfW4KYtVR/jxqUeUMV1HfUrN+IIf
a6g+B082vCXrjz3ZIQcVhY2G4IJQHi6ppvU2svOS0a6UjLf7D4wPRvbjLRym8uFExF+Fc18pXAPR
lS8jcppKNZD3GcC5GX7jOKpUkeFyRn4AqAycy/GGi3IiJV12dLADNXiRkAomrxRBCrYr52GaJKMZ
X2a5LPzDf+wHaLRTFvJLEPR5zFqYvpHNAwizOo2pVmyBHl25J3/FPwbr4fQa1VANMU1GYPDzDkdS
tcG3ogfyOPvmBm9HXyfpTPkqQPvhAby8tf5MrmFFQ8J90/nHw0Tf8acfEKp3MZPwOQbz/reevGnU
FuhtJ6rdYGHGgBC804tvzPesFoSRdEgo3RKZSzmyXL4wWAiHmhAa/3AByACdV15g+s3Ob6XV12G3
QWkHZHtxpxNP1KGhkeUS6G+8mqCDMMBc9JZgMiBjtlxipBrKrphFlzmLgGpbOSKA/FLHFBFunhdG
UrIYKE2nWciTVCacbysvlHcPxBVEjZ1ssn00yCbgm+B2nJmdxBdmFtzOGusOL6UEuA5enHJCgK3f
V9pMvB9uwaioxmHR1I5E1sRgmdTz1ewQ/5b/ixtwIC1ZrRDGiN9IwxVYrGcLoDjX713zU4xzib4N
oLM6XyfQuxkAKLzD5KBn2TPYaLS7nZiCpZ6/suVQixGxeFuM4PXNGAd8NyeDOQrRDNrarRbpdMTp
zzLXnE0rrEjTn+yJlmedehNOd/ODpHcYIhcs49RX6HntTuOiqz43lqnaoefeagTXyRQHg2gXDJEN
j4yE7aTnhqG4+OjL/lXjTVvxgQKnW8MXnDohgFuIFg0lJh9bh0t2ycXtShTDMnZ+X/RYs1R7Lrqf
A0sJiWnLySPEvwTX1CgM0jK1suVGEZK2lACrPrWDvFnelPKcL8UISarTElfxEU0o4KCGwUvXZcGQ
xI7XF7wl0D+IttRjXTLiG7uJekWj6azo9qqFQUTjyEewwzrFQ4C5RIzhMYBUjvE7UolUbVW6smyh
jskz4HXOJzQGoJn2bXtJ0i7DLynlZV7dn/KNHsI2O1S0xaxYNnPaETJ7VLIr4K0QXwSc5GbBi6KH
G5wTY/7pG92kb1+xDLvnPq8qkwhgHooC8caeTjebLyYQEscTRqibPsTq5ZZDEQaPkx6WdNQ0qlBE
4u0QR9FKjakpYcNCirsvPYul28oy+vvweiwS4SmbRai34xFiD/WG0A==

`protect end_protected


`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
llIaOLbuybqQ1JQ3WV9KZwiIlSa46gwOnWdIZzWkqoorsM/I5ukV/lYcWsxKTCrKWtBBWu+YZRCL
yoTwafDix8UULWynT2mmrIbsPP16j5zpiw7unt5Cw/BBgY177sZW+Oi6f1Vs/mxe0/BLLXNG4CpI
qD5vtR1L6Pi+W5koxe714cRITcAOP6AxPz8RkMlcZvTO4Lz9rblIt+7ZT25hqRh4xBYxVbVeO094
5qgh5gTZSKRb/LqyqOy7WHVfnrkiDOqpNCTlh5fiHoeaw9XT2IdKiTryIAtLmJObVdPsSl5JBkLw
soCSd3u/VAba3mtfG1tnZQ9a6tLM6okGx8RMcA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="by3h6I7oY1J0GOpdkEkCp/E40J0Hho2eVANO/jF+Mp4="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
oIB5K5ZeXNm2oQVgyernNeWnSnSozji84V3aLUiNp2zw9Ovl8rMnENh77L7GHNo33n20KlTEnX2w
HN1PK+Oky+C9W/oEguhon3EB2MZrNdBe++ySQPqUoJqQBElQaqPosz50+gIuMNaC5EWWuprkc014
RRnC34tVhC4ruk6bhEJvCCjWf76VKNi6C6ntfIeFyuwX5hNXzrJd8TZgv0nAlz5qODub7KrJGtOq
b0kOCVBjqfU0+dxm8hM+5fEZ+LteEUChN6hPv059ve5/CdngcPIp/Uywl9gegXHqSd/mLdjOqTQ3
dmcf+VujnnlOGmjdm8OnISwRF6ok1ChHdVN8Sg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="8eSOFS4laNP9Xno+fleY4/s6yuC95xqBTMx/iiCnCw4="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
SSo9tPXK3V0icXo2Bnb7SgvwojmKoRsuFC1J7WIxf0gEPCQnYUrUNKGSkIJBskTuZpIHETs7R3oq
Z+OaAU00wWAI3CJQ8yVRz4pfD+gCvHeZehEFBemqZLrMbZopOSzyiYqQxfBUBtYzecgiVHHYrm55
Xe2kwHXsiiR6/lNNCY7+HjOqk2NDFVsNZdbC4MQS1JTtCWbpy3yq5YFPu/aJ/ghXPgRAfOB5QX6B
PQqBW+GrddUM3aiH7IKk6+SJE+dBN6tvtBDLjjAQM/s4otH3sl3XPqMj/akQZPcsus2cgZCWIouN
IiIlbZVgT6pKTlNxOUl0TskjebUpGthPiWfqvw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control xilinx_schematic_visibility="false"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="51tWS+Slbyx/5Bvn6FT6RxFVPynIpuysQnsAqq6/rfg="
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
k71leBXT4W1IHofX7hTC4KM4X2aanurYSF/A0phMyiS0jdwPbSDMWXsFW0CUo9z18PJi89E+0qIn
6OSPom+q5PXbW8xamuzL4gxLxDrTjTAJvVHLTi0lF/qfA2mcxqCp6s+2btzh+PMFUqFDswH8nPMB
0HBgAe23yBtm6VAvxzmvmHuUA0Mrjqc7KYe1eEfL5E2QQ/HJvBoQxjmBCZYQZQ8HbF9smPuMJjvV
mRgRCAc+vD3AH5wCGUzfgYSAS6PkKbUOgQ/8b1udz4qmYnnIN7EksQT+Vnr0pXsZSPzH6XjskPUS
lScLosZ5U5frADlN/MlPmR9XGdIUf1ITI0hWUQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control xilinx_schematic_visibility="false"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="7HBhv82hSwhZaSFndYKNrSTV5DJvE00I8+lFbdCOHx4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 288144)
`protect data_block
2E6OZjTEOWfBmWCcdvgsnNt8mLo+QGMs7+d7ngTkDgd8aRLVAyZw6EQk0P1J1+XS2Fdv9ismq3Yy
cRvSrp5kr6f6aB+qe7MGi/agZA16+VIN3J//oUTCGjFcUaFPxe4fiH7PvOp/pAHtFpz4m3IV3qzi
owEmBtF1OW2U8Q0878oLdj8uaFmNDQn/osLIVN8uBE1yHo7S09fbfJrxJISTDe1cMHRlGXoNs465
N89zSElt9XlPEYEowpEU+MocFSWTGFX9px9tRLtWJLufryLQgSj7MbhC97wUYeFCoaSmBeOFnAcq
cSrrlhRR9xRDnAf1cnhwWsHUtxhhbItrP652e1wyRkuRWnuRwH5n4K6CsrxsKBGsSnDV3sc8IW7x
UskjcLCPOq54gJT9Dp3OR89Ia3ff7DLzuJ9ER5b/iHIW+n/ASRXyWHP9BEdpJnuTLGCU3GMAkeh0
YyVTQy/WkZIYaWB+kfUVZCH4KckHAbaCn8GI9wb1Vpm2BwHW67Njg28KKKkOSSaq8oloOc1CQgPp
QOey9S7JRmFq/HrDKqBm+GdHeIyrPeEgZH8pNl/1e/6UyYvEmSwncucHEUk/rTcTNPApd7Pyh3G9
jHlpcvHrS6EBTKskLiys3Y7cu5U/cFwbw/o/VFeXzXavYZvBp6Oej2e0tRtLIaQxpcSzoN3U99uH
a88iXljg9+Pfq36Rx9dj0QRQMaunTFFOU+KToF6jMN+tmpdIoGTnDaL0baUR51FSG9TV5LFqylPH
yhGI+medJjWtDyFtYioZHMsQl13yPNBiLfBP/LhhO/C1E09/u9h6P+aWXbUrJwQ9xdnCvbT5uu0o
KOgMFwMMrC3VJWawbJbwLXXde/4ij49EcqMtNE/Wf2qNIFl0Gq5di6TsMf/u+fdOSX2usKbquSpN
BzDFz7CG4ozfymyzlszhcY1jVsyOXh8hxpxog2kVwbc7QPjAyOTcTCs/+JynKHBQLXhrJT3xjfxB
ryw7gd8PuIPdYJmn/lEsvs9KNDDLsCNLY10FpM2DWTajkiygS4p+yW6zGLWA1MncJsifxUG1nYo/
GQP/oB37/1/eEzqHi7aVZ15CagbqmOvfRCEHONPdNqh1P8JWSKz1gVSYykEIHZP1c34sV540Q/k9
ahZRZYjMype86tfThQgJy61EiDcSlfclZ1P7g2oO2zcyYGRFIGlF8GRWOCHw0nNg7YOE8Tc8vCGI
TnaKFHWXaRldrlFKpxgct9A78IrPP/dNoyp3do6sYynoRUEGrQ4ysHiXNIPf212IhFNK10PNuaK4
t5x4A7o8HiM5480KKePkUVcUEzQf08m9qSqHleoJ34mF2qe1np8/XL7XYyC5vHq1qQTYRt7Xiz//
Kln0VQiriqznWwnILyUGmFt7omqSdyGDa7gh6h+e3SmZT69nQq/rrNMqLR0FUhF6kSwOYz61BwBo
Doa43uLmu5EwP2Pq2Aq74csQfc5/mszbGcKqj0Opbnk1Dv0CJ+WP6BVmNbM0xINvZ0f+WoeBUUdK
X2PmIbvNawQqvvk6jE6F+ep9ShkCfDglOPIkfER0x/enKCfTqG9FY31Q6mHwTvHzUJ+v4bxQqCgL
ZCHAPALHSFvW/bGLgjGSJl9nRhRG11nXW/Z8vqqGCbkyzbcAKKk9rc6ATTtzEsbCmvuLJ7HCRP3T
RwH7PG6frOShgd3u6AZeVMNdJHQ+ZkfzcoYV1lhavxJt3GuAI8KYih7sxzUhfXjR87e93sMeRxvu
b5SegA8tA72bMria/6vIsn6KDFWcdyLw0ObHI5Qx4NT4EEZ/XvYU0OprCoQ1ZuSV1OEYCZsqs59k
KI3bHf/Aw0/j8w/ufTZ3KFJJF4hgTcSAMu20Lfp4uEShvBaW/0THCBXEP4vBzQf6iN6c0KmIsA1T
kfpLprhrhc8NZo2/loecNbLSix1dzAMeqFll2XohMaOBTOf7sOUJyou6+/7/jZsYGDlIx305gorf
ZJn3vO2vWIYZjWfbKo+fSID1d9LfTrR2nFLmJ6omOiT/DyuzqaDjSrrFEu9WyWBCL2je4paqgpWX
MEbxTkuuvvTBzTuG7QoOZFdTKe4JKYWbGHZ1N+xVYd5KprPNtEeUQUG1uWitc826AgoWdLkl14NU
+zvZ7fw6wuJfw0oNncenb/o+GV6u2C1UZfSQUZWC/SsK2e5uCNdL+vPo2bzghwBFXOzVGBZP9PMq
bVXz55s3aonY/kWUNN3F5QOCZ/ZtOTRnsnmAsFkE6mP6xidlUdZRQvQfsM07Gzs4G7A1VhGLzr8q
OIIr7/3u3Viow19Lqn8xIb7flRgq+zDtR3amUldVSViMtndwnaJuLXJIPin8hwHu7l8vwVNhIhMp
PJf2DzTbgr4xEFTonQ6yxMeOI8dHxM4LXnJWPJr8vh3UP/BSz1FC9UyCpMzeYyXzdXTdLhPCOac0
DHhZ8f2Dl8/s/eI30Jd+9i8xMLWmD+l1d1aeWn5ruyoHZIDUccPms04y6cieho3GnRIfJsoNsNGY
BDY1OCBxKLLjjfmHpoQ8RbRFIvC39VNbEoYuW3Q6mX2SP2NKIl+dykC4N81CTKGkfywUnQJp0Ej6
uIEbICfRMhx1KBLF1cXMX9OSQJIsZmWlRUuVODPzpQnBmvkJ6ikPI27TFmzlcAbM/Q25eb0yC5I+
Re8UsPlRIrs5TyptoRlZRo2hkXzPzPIyf1iKUGhzQqfFTgsCAF/Imi+4h8bbyUi8QpucN6V9witO
X2HgVIsDEoZ91YubLnygTYACSAL4p4XFacIP+FJKqAu9CwmJb4D0uUswdQ2JwRs8YCmq/J5khRnh
/NEGZkhyV4SStcJsVZ6vr9xQ2c7SXgRBuI+dpfGAe+Ua5D1hig1ZRlxZ53pAn/TnOn9yJSsaDYMO
ti5JW+12LKGR6g6d3pGYp88gmd3EWUauGwkW7tS5OgtxGjaj69RV6WU0AYYn9lsp0+CPTzknjIlI
dG4wJlcqUvp4ZJiiPgYxTpw1dGjKdzjLR4xVIjwGwCb9EhJe5/u67UV4YVJbBgPAI+VlqcKqz6Aq
EXR3ahGD5sJz5HAhQSTyZu/Ijd86LfcHw8wqrPUECNG6f0Bfg+aOgvNMbssLOHVgPdaxUj8VGjaJ
TgQiuFc8K87g3bqkFELMaZmVyo0+PiPUY8SwIK+j5zvViLTS1U5lLDWo1KhHTGbriAHMfjIBYbYG
S94nBo28JMtw6UZl/6o/pNkbahCH+VYOZtirSeAmkkebffKJ98YVEvxYnIu3FfSh3x4pOLnCvm2P
qPOC8Mh7xR5Udo3uIA0dVDXuMICu+LL7UrOxgQZC/mEjPlLTy7eI7t9mQBZlLxpM0CltaTlwaIWZ
3mHktNUjQ0zbxuURUPr0SJ7bF5yr+Aja78y9nuMNh2kp0y53XBWs/Tki7sRoDcPcRPyNjLNO7Rf2
YVoP/L7wz85+Fx3qF++UN1tv2tubyEYZFkhrbZhRZA+xfJxVknSGm+PqnsN6jJrm5ty2xc0KbcNI
Fiw//N1Va9j7VWL+9PaltVOdPPKUU5hwW7xxvoJDbmGTrSJiquf++yd3g2UDsa1T6z13l+ZhKQcW
sntHBEEmff5t25S3pApWcPGdwG1OA0ibXbz706x2H0DSWQ6eDnrz2S6DATONgPZ9GMJ+FbFNaBED
D7hqi+5I3Ve+ma1UdhnlEs+fPuyof6JOFcDYaZIhtpb2/6YDByC2eW78IjBt1xVGVVmzH2fVjz37
E8aWGTju0vHMDuc+6dMzyy2bEme6kDHTgACP1yPlb5HE/gcRz06I2wX4Xz2sPHKlMX5p3MMBvVbF
xo812YwZtcentBbTGM41Rbz06SS1ZPKQ0CYJWuToi5FAW8a2jyuQvuyV9k9WbHjwL21HN5dYdPBz
a8rA6dEeHL6TmbuPTPnLtwlb4Cojn6hYOD4i7ZMVA2ING8TvcdWx/Da/3TuwerZdxxD3mq4yGAcq
ue0im3Lv9MO47UpGTvD/yt+1dZfUj/cAQ7FKdOWsaGrC7ABohAgsVBN7U1xUvfnwP3owWOmM01Ea
ha/Ko9F0JN+061Nln3ZPed3Ky7T5Jx8mlA3vVfh6WjybiICwspYbhDepEEKmePjeYWGb2sMJ52An
tNYWGWY+i+KQUiJO3WfE4ZgBk27V2FISM5I17dGwUFqr2+EOgApFISlnROCagXZYHJL/ZzlFQwjN
3t6vmvqUFOLPIEe0NdRjDjSM553Fhwh6TdZmEUDvmitqKcCwId8ahaaD3F3KwDLBUop4eQSH86DD
+Pe9UCQnqXS1cLlQMw9EQeQ1blkkvNCl6pUGpznHDva7DeCpU27M+oPk2GXOIidgoCvUPOhMx5X1
Qu/eqSMPAxEwNfQowPukCAbXEaUOL6rr/WUd+qAu8qeh9XzDgrDegyRwMYzBGsXNkcUae3QH2BBW
ohOhBVGcZsLXHbXyifGQKWXv3bSQu57XKMz8Kaa/+P6CR5yPwbe6p2FHhTdXkuDdxrsw3qDBMk7w
uONqD3IBHZaABuZyvQgCSxijt24jsx6x2IFd7dHKOSIpI0s4Moyowulad29LZG34BWHtGMGkKird
BEvtfiZTClxLwZ6rsaNYY1G7zLtViSrATrKq/KSasYnsxppvGJInRxjMEZ8V4+d1e5ByLMBg4p4M
skAShhvNS9vj88adJa5dB7Ci0p5QuaP17WHlslTtsifB63ZnAAt+Utag6ERnJFGuz4umjCe7hRCA
Tmz0KsFw/KPNlQUFuWWPhY+pZi38u/voV8IEDk0KS9na8HdM64eZSMvp2GUmrRM8KL1bdk7KSzkV
k2+PtJLDnir8xqn6y//Yw0DG9rbeMDfXjKRP0g3mKiZ7jhL5paZ3OUZ6zGt6bDxeFTtbTBCbUcrc
lObNQBEvlkW6lPlzQCUNK4ERO3zV7zf5qmMzBiDZvch0zM5pWmtHVaqqWJGPbD0CIpD9DtZC+oIS
J6DuL6qAWLVEu8K+y45M3ahBPIZt9N19PRuC+JSU4FQBpGXn5vnZwrArmIjfdPJo3QO3MRMOPS9M
md+Q+aeMuKvchgJGiwUMbi/CzpET/NrYZwr+zXAI3LLyWF4YD6A+hEGplr6BMpiSt/T59VyrvwUp
PMMsvFdbdZSNLz0bOgQRhra1aiiK3xsHH7VLqETZmQHVMko2zeC3At9qnItexccxwkc0cOd98Bmo
HozhX44W1yySaMnd20IGhdwYOPM8gEwddBLPicyivPDbu6tZ/HT+YL/ZyIu0MhtiLgBeFJlZ2n2N
SqhvZ2nZAvaeIlqHoFeRFynZndba2JC9ymgQXnsJeuqoCAtlTyz2D7D2ybKUtpYWGsc7MC5IxcKm
KpMu7iFYimQLdu3PzIiJvaI3A2Dl8NrMrooK4tUkA6hqlvZfT5maiK+sdWGd14fODQ7zVsnIaEH9
ayoIXPPi+cOmybv//MkRf/mXOhpBynKKonGj+0Likx+8cXMqCFrK0woxNFOiWt1xusai+YHq1J6a
++WDlc8BsUhrH9usG+sUuEYHOlt58GNdLeuQG4AEeqekUKByxFw18LLFSyGKjDbIeABh/j/X1ACM
US0P6WXVYSHaD3YOq2PzivDXcZIlp5wUHKR+DvxKh/fLdH4HxIAWiFrzsgLgKixRfv7ZWUIqXKwO
VuFaw612900BJFQaHHCeqfAHgFnuxAKF8xIfXxS3oI9LAPjx69aa0SfbKs/XmKZ7BQVfJXKIrKXp
y9AwqAs4IUkXjOORVuk2D6XXaxSZyhwGRJJAMj4CAMTKHOgP+804YA1dncUDEBmykJcEQ3UnkgyL
/iJdVP+foxQvtcay3qLb16GqP/rTxtQtyx4lojIPyp6tLhFYS3/LkATHhnBx/XVnrQEOuH38G6nR
WyJpaaefEsAYQkVUHXSMFo05ZH2NUSZ3qv//cYvGsnTNij3wdDu71ZO1MkhlYDIyfO0rUReCtoM2
RdWTQnBwFUA/mF1jYaTz17O1BwH0djkAucnHDXwaL+SRn6rVFvNp89jj3evyR9jdb87t9oUuAWDw
/8OzlHpYu0f0vQmTIkbqx3y8agRZGFFNPwqnI+Q4h/XaJG4pPZ3i6B4MihHpnh8shlk57O7wq831
QQbw3jY9OizOWUqvF14V0eFN6ZOYrDRpKqOpbe9z4BgtvPt7IoOM54c5NdU3hKl2LD8YJO8PGunv
Bz+PeS7LhEDHI7y64nW120/PsCOqbPYyC4vUWug1Os/qHbWI9Hj7pysfViV2GlHj036bTBiEw859
ITpNDu7yJIPqXIMmJz1GS59TYbPiz2tyXY/BrjBsQ6VU69P2exRwGCBzulcF0tARCFj3PxVy54UD
udL0FCtEx3UqeG4j3CkQzpxUIqSPaGqARdLLik1WGu6X59Qkj1PY19XovZYdMHxQJFEIM4lSX7Ey
0xgsIFFC4KI8FOzPC8VmM1aO+z6uwkmlXAZ4pyOIz0yU9eJZc23DordmL5TzFkn7WxcppeE5Gf5t
anqUKe+mosvOivI2sdjeUUUjkfs0LKiYeGVMd6CmBukla1X/1jeJCdmMMg+vvbuPdLD42gdArO4M
2F83pmtD23b0KIS0kRnNB4LawoFME/XZPdIGaUNpJdkZIiHcNrOzNV0dYNyO5Qc4MP3E+h6VahiG
l5BKUCMkqkwLP5NWghrYPQtKusehtOTSZSAzaqeB590S2XjTdMDdh/f+Wekdv9jmbJqqZHy02uzu
Owot6VeDlTCR6BTNgNpiQbLGnEe82WlIDFBJjK0RAOt+V98Z42mPpV2iJ8h6HOhZmOJmUoiN+aig
Yb1A2b5MT9BwVt34Ta3p+mJGLQlVx8MxHqvCcvx4jNfoeyIWRZCfod+XnFBQCswwpUAQQmRSjTBs
76AiRp7ZqcEoJ9e7I3A+Lag7RxRfGLAaL69MUkmLUmULKDLaG8hnqLobBb98Z021fM0ESqefmgyf
LR3g2LnlUknXi4cwSEcDOzTIaZCDf3ES08rzgFFildzu/WnW/4iyeegAKS9f+oI0S5p08lf0wr85
EJrbe7odRAIaTA8mvUAHkaE50c8ypPgw/HqFg5B4ESm89Yu/Rk8hpZVNIA7r0YUQr8hY5jPEDg3z
Aew4pwIjUHXYYEIyDtj3OKtsja0x3xsg48/y+K8jAAsh2XAXFBNj6veGrnNNt2WK+Af/loxZFegz
ZH9Aqwu7VioWsTEg0MutGHat2sdkrqyEVi7keJISdbGzsqqAl89is7E2BGJ5KgXjX+AIhqUO0ryV
AqdkfxmCarhP11V7GagmSnw+yzehj1pAzTmTfPpxLo8lhpmG9msN1r0jk+EpoALyyKA8X8dtgfVj
WiGkGkGD7a27S7LibLY9wtykbySk3eD6zcMYjXXKj6eMRyzvkzo7cFbKwevRCw71t+PS+Z17E7AT
oxxSEqmY70fC0pt5uepuXbms8J0ktMwzP5lLNJDBl7o0sigRp10NS8TpeikTLyn/UxBwEPAB0GcW
Xefv4uydh7DnzAnTpNEphICb/kzYp8a3fzNoY5aN1aj/tU1oMof6eb2hBBb0xbrGC8ZKnHGjuX5A
as/M2WovQlJUVTcJbieZaGlw2Z4OGOPDnFOe9Lq/cNxtoJL/XJZDviQIEpZSAV94TOV+jp3r4goE
3EOimvA9ee/KuCSb4NUsEXGmd4vuxbm7cN40ODmFvhdeedUYNq9FGcYJ/fqxjloW/M0l54xH4QX9
79oovWxSkRHnbBWp707DccAF6QnpiRXC+drvAVNXyY9mBkD2q1JysN+tjDd/rhR/eNGes3X31Y29
e0CIvZztKxv3abPcnsSXTu73y6Yy9DA71rffRF2KTh9rPk6guP6RpKW7TRJ6SiqGsXuE+v+8384v
nEWj4SGc0OvaYDJkjNPwFLLleQPqQXin0h4lfokyOLgnI9kjKVylaoT2j3L+9f2OLDdm/qLPRVcJ
MRtku19A7K77MkqXrPIpA/g/rpv7Vt9gq4KJLNjJKg+vzwfJ1E7v3W1qw7ojRtaJEPaeJRvpj4uk
09rYlbHFAzsGPWAx9SwuaonFO3+5D+KeFikzmHKxsjp5z0Lcm8ZIFTYlRviZlLnI1xHnF/D6Zxzk
nfGzc9vnbrF2PunM7T25xGsGSqa6DjOm/oPSfBO+4cCnmfrPjg1TComnzg+NLNsYEPRZ2VDH0/cB
54avzrHvmWhMIaUIZGSxZHTMPGm+MDatzzeQej/ofanxD4Dc5Ai8MNAaiIUoMZKxJeQwZDg6vxkU
U+znC5PKHpqH1IehtXiFrNAt/vCvxBxPThExqOba11bNpV5qbzayFvYrtonqCl5MktZP5x1Wq9pR
MEOcyCm3CrFtbqklz1OxlBkJJxK0tnt3ALFwwIGVOWE9zb2zqH3HpvQNmWqUPdpgx1MptLBsFNke
EpNZVFNX4bEWfvHFfefGFZdXvaatwwQvZjkwwqJL0UsAuYecfXai+SiwXY9NqDg4ZgAy71t9TZvQ
g0uG2tq8QZyN1/nBx4SeowDxninebh+1kruG7MIW7WZAK4etGztCnM2smgh8ig0vxi8s8q4MMTJa
1gcx7EHDVrXp2yPHDM21WsxSqwf93kgLco6d8ruTPl6VUk1w3zDG1q4T4V7TwO20mnd551lOKZQl
HCCqwtujdoRxnnB4FzgBAneO6wJwVbTEvI1L1EUeUQCGaRjEnTs8XBjA+0am1snRu2ky+Kh/KJEA
zpWaehe/bkIayqMqAulQNw3RQtlXQ/DlL4YoV8iCqYGqfK6fzWGBVsX/H6xy4tZRGssZq9pBm338
o/JXbg4FvX2k+jqUXBe6boaURPfnB83XWpggbuqPQFbY8ocaZUyUjrE0zmVLtUbxqtIt8IIKUFe6
DAlXW+A10IPrdHpSr79P8v7sLwGn47Fwxudi096RJ6lOGVBYz7xFmNwD23ou7lmvQWQU9qJu85WV
38G23TrdN8HYSfeXX4dIHGdia6qK6SurWcCCtYLkoFbdECyxHyB5VyCmx4epPIDJem4WFMi30eRP
DHofKCm+I+IP+kQJ9gwk1iZM8Wz6p5LiB4hrOltKyxDIjhdwaO1glgVhiMfYtodaTNwL1MRj5Y8W
wZmcCBTEgZL60H33Kbws5HxMuLWr4jjU8J8zVxYtg/B2IR4bqPMWx7bHjTbUJyNMLWXSwtmXO2Fq
ddI0MwEorsIXBu8WsEUgmZMN67bzNenIj0MpG/ux04QRRG2kTxr4t4wf+U9A3XSvP4bHLeE3PZkP
dVXEGAiFzrSNKICUtRZjWfOF3G7lmbM5nDVoYxIbLkJqMEzdIY58oN9fG9Flrb3LywPiIFswChmw
NU9xuPWEN9OQ4+cA07kp5xtEgwq+SBXOD2rYcfsVoKNo6khroKePp3LYnWsI/H9nKauEyLRkXgsW
HgmGUnGawuO4qDXmxzPfwEknI7iypIyKDE6qVTx1D5hc3x2w9wK7gHa5kQLQ4eqxcvw1HwcZL4kl
5LlPs8TTkoDV4fXdyrlxfKbLFTf74dFJrz9G8mixiLEUSyia247b7efR8W3hwTCzxV25/IdOgArZ
oeFS74UbAYX3AW82LZP2wtv3tVixwt95c4EmOn7vnrMJDO+SNz61USKh71G+LYLQHB9Gj4TqebdT
O2AgMsGrFuKpWLQ20J2N2JTVUEr6xPJajQIyMQLhYfYe+XLns6mLALKX1ZNXYL4Hp+/kzSXGkAXI
Sm04bLbYc3ejKU81oWDqrO6olq1np55KNYciCC6n239KBhk8kg9jIlNvyV1GLK9H5m4fbmR130/B
CFRLUUr8CuE89FcukuM2oOKPfjAlDnPH/5Dj1zlRLfJ8VjvVO5HV8a0p5hfou3sdntZ1H8O9Ablq
QyjpnhSXnnDJt+xf/Uw53wn9pAHk+rO9JtMaZhU0Zv2rDFll9HpsGw9GeRPcFdP/vAMPnpizRZh+
zzJqNIy03oXdQRKwGhQZ3kLLKKy3/WYAays2U1XK82Szcu3/Supvmg8TpOJJXuj1ZAUMgcp0Cusz
DKF+ytDdyHKZDth25yjrGJKGBbgs0gW0A5lQbW5iq7X86pU1yzpsUuZ0Hqb47rQLVCq+b1zEt/Z1
aMtO+vVCK0eXPnldTtN9g7CDOxpvKrKCgnRdb/SQKBJbqau91V0IE+/ZBKuwBbcIhw4eG36O6jHu
XGrgF9mzhCay7d5lTfsLyBeVHiLTo9ZGVa0ldF85tzFJILu9vcMWrG9jXhQhRhNufyJOQ73+6FZ8
jhPkIzdfcre6Xj/MISUk85iiFsyTrenZVvHXZh3bp9tKxL+BIPgOtqrXA4iDMEGjP8iOrmZle/nd
y+pIBn/vVHuxTe3Or9XM7yxxUmmo94jI8zEN5CoDDMWe5ZGMNfWTg6eXqwtzcI6sU9Q685W9lgbh
GefrnWuX4F4/yMdxJ35y80y1yR7qO/vPbb25BpqhtB5912mXTq1Ga6qwCiVDrk80F5yYO1F4OkI+
e6ESi4uzDHvw6m8oWqR7FMgeb92vFjbiVG6+ZJFxMSFN6RV4IhQK8qiwyq/TmzvSVAYXLKQvbDQ2
q0yhlhoiDXUbII5OB5RRCqqXtzNB9YlaA8U+AQ+V0W/93QXXv/l0k8a9/Fa3HDgTeM4ZMsBw8Eho
G6BNUjzrg/UL2z4vrkEr2bFAizueqwDwbW00QkwHiSsOaxKItJk0SYhXbvDbe7hxLsE7JnMRH7J7
QHOV0+a+r3yzKeKBnRyUCxqznxcw+J3FYKPkCWn91TQRZWhbp9ZH3anNpPNHGh+wIIHekeIjJ5Ku
R+wZbRNEhiaVfLHY/KwNvTU8iRBbS5CJwwtTipvftUHSPlK5jgO5wNSP3zWdwCAf0hJL6fusn5tO
PaphBex/8V/vWDngM5QC9yMCkZHI3dsuJ9ziDdC9nZrlg3CJuOgxZfpyRSj/KDXlCOKjyh2YEJAj
IE9IX26euMHiqnmBJ5pAi1SEaorTc1IYjmctNGMd3dB3K6SOLxWnYRYnwYRfnxXdWJiSxzV+w0s6
Ki13vi35Uur+2aHz7TLmLO0+KgzSZ467yd69Js9uzp5g2OZwY9SWrJBTsjsJY8BaXWn8z4OPT1nF
Z8LAyiYhejIjIUqApg/b6inu2pi1CbGPhoKAnxJ+vLw/ByINVBWNbGIDmyk4yRZF2gPRdLuC/4eY
gdip+RXR3RcM2ro+yShaRpo4BsLfYCD3S+0volnqDBQSD8D3tZb6Dr2xei7oRZMGVT8CUKHeL4Rc
m0preRkaCkpdd29jyQjOF2akqFF7UkVxiCjST+Vv7pBK2iDSXjN/yJU3PBVYYD5mCiEsV0gnP0Qn
d3d4oDI42x34LZqpwHFoMCOMjKn+rLeAUOuLwvkPFer3RFxdXWE2gRRRARjiM2cn0pPQ2sL6wE9T
BHriNcR8Nm9lCi9l5ElKPfen7ZW3L97r5ZnUAcNjyKn8jQk1azAQuzcaB3kbd7h/4Mm893GPyCRA
8YX5ADg5JCP4nNFH5/kF75PGZtBuKytOGQMSbmp9wAiskgDIq4g9Rk68IzdaLMpNQEr0f0Rm/bDs
g9bpNTOJOjBoNSfisbZS0yVOLq83HtsFHU4FJBL79eRH0Cv1tOl9v4ClqKU4ksyYO7QgPrzb9mFS
k9lPGTZyt1VJsxgcg2VCfIijuL/zU65ZGUinlAsjHXC/vjDC3aYV4Qsd95IUTQGsFMOD/LCdfcQM
FFfqFc2Dcr0uDeLa7lrmc3xY2nervnvixOebqRgjDmoN6ZCqqBrP5+956NBHyLasWd4EGQwXl302
b+Plvu72ToDQk5r8RLiNTOYyQmZuiujT3ixhzd3WRm8iBlfvWLPgeRqv5eGj/PH5ETIEI1s8Aiea
WnWkvzpQjD+wr/He4t+lL8bdRLaVVV8E+LhCnI0WtSutKXgk9W1WJF9RxKwDXocMuBFBNu2Pzz+t
0vnwzXhezzB8/9fe42zUjNt36DgtBI4ds/tiNHHV+f96Am5/Hz1hQLbh063BGEZ+Zvqqf9RmlxhY
0sqjeuDtXo35G9MLqf/+dGSy2fxmu9DVGem4pCf0huLqrMq0FpaYi0+DyDG2yg3hO/sQlkP2UyVI
q00Tq1Vygi6GanrFUJpNJdU0l890jo3K6vkTAFgXyvxK2gO76iawXeIb+RmDaOkAKm1MZfdt2W7J
iZhy5VXo+zXHMXyis7T5O1tlPacHHScVCQJvgUpZAaB0P6zL+2Rdnu4A8S8ht3asONwN7JMbc05w
KNeTO2ORg3f7YY9HU+2MsjFCOtohkQhIR08D26i7+rDFAm0A4J4x+5D4BRvip6hogoKGaoycFsqa
hcKdtDdxaMow22xUM4WtNWNjsP4/pSfHKiBZ3C/y9U9lqyv4ByalyoluPvVjJEqj3EquwncWUN9a
zKBD9ErOPdbbcPkSO56fZIKVFhTR4jvnGkIKH1rrYEU1Yruif5VvJPu2kxaxoDzJd/HhWYTkXWRL
ALTGoG+QUsVlCgarnbXw8siq41kj4Pxm6dkh1dAtbrtkKkq29bI4s09uRTX5fSsRRezxpZ3BY1Ms
A7jAMkSNmUaIG5mxVhlIMKuMHx20MMPhmM3J0H9fYW49oIblAJZMtu83Y2QSd/3skYNYxdk6USG0
KHZ1NNyUCKHusS11GjSdp3wYvL8ezk1Ax+5fgC2r6CqLEF37RPmzvNT0dCzemGXi14vCEEN0YOhY
y3sFUGVabIOLXrieKa3T/nlEtyfmGJ06KbxRrair9n/XsYMsP/c2lQH+7MECA2Ij99S/KHsdNHj/
lKmdcVfJbVdX+Gnq+D9N0rhdmTv4O5dmnp+Yi1mKYX9WniEbSIfHseSsM8LJVu+nD78q8lgZNkbd
NvBpvHkkVjGsVbNFhvJ+0JAPgBEt3XXkvIZ7d3Ogzb1E3D1OoiuiMKMjpLwKhjMA06OJo95YzVw3
U6v2bi13QEewI5bHdm8kwmoBHd2G3zIX7+dQlYzTDFjLMzzWsGvs4UHNGbc1xyR1GKXohL6G+uNr
mQd5NvLOtQL6TIzGw7Xc17UbEs2mEKsj2aOoA8vgGAgkLao78KZZn+9SCBWDcnzCAIQf8FU8kqzM
MQF6fmaPUGwn7jGWbFHBT3d5R+4OJ+dtTpzPy5Dn9aOl5UEvqBXqLhbVW+f8mlalSOwtsgbxy69R
Eu/8yGOZnX4AbDFs8hNu80wX9EWOspJVL5pyokJsu4WLe1Vh08cZY1PVGa0jARLfe6/0jgshLi/o
PgL7zuASGiYwr5qqeX2abOzryAkzXXRiXz+n5nMroUlECOvk8BCmXrFBUyLnA6T5451jlD3S5y5L
CoQiuqb/IlkkL+JjsF4Uqr9k+cL/zN529uW8VOi7O626Q94G7UQqkfPDpWfDf9BP9i1FpdszMrD0
lJkZi+l5+wLjpzuq+8sjT1CMCx9DWxsf+9twsoFRVMiBwKTsmhyIiIR61DW0oSr+Rrq7h4W3uTJd
cnetZ7ePFkZhFKexf/Y2hTlRs7vEH7s2b78WdTruLdCwwCObOvY90mVlLHbRBiUygN1v2WXg7Ln6
EQythEn4XZBLEBVV+k0ALAcTI59n7u6p0D+sYMCuAJpzWKwY/Hqsc1K6yQ9Mvb6dp0ItKB+Z1OG8
6NIr4ma7E1GYYuGgyjAIHVMp+8RG7HU8yTXf+HghdZ0czw7ERUjH5/6iOrAO3fHVvCR26ADQAVcZ
qWI9Uh4X98bpDHFcDz7HMfx7uKRDpDBCwAmHcdgHnYDm+qAQGKPtj3LGYaM2qT58jJcJFM7RqwsQ
bC3bBi4M7jYVR2mUnlHCHhUR+1i1JJNsr9+GIvQxAoJIn305FUEfpvfut8dqNe+AzNWu9TupAR0F
B/Ivt5wtjzGxnYU8jawG+8WIUh7cR49XKkyNFPKHY8zCWcouacriDKJw/8FxXYEdLaIc776Jh0PI
6Ztbq/pZqEeCU0/xznLuX5oeOnX28HRQvWxgpE4SZBUpDg63LVMmnbWpKHRC2sYEegNAQbJ/E8Aj
HXmR3U0TBaimi4pQ838LHYMK67lNPu4IGcvj1qlDm6y+o+Jy/fxIXNPq+sAfT84C7tRQWOUuVzBo
6YW+IJUKgEQZnjK4JO+4rfNZ5sq9hUAv8E/Ubf4egUZQZt2W1Urdc6Z7joKdlruzgdUdPu0CbBL8
gpvHMyMu829E2pCA0SHVak3di382SKvvsOIo138I0jGjQQYzKLeDol+F9pobfsQIBAiQjzAVunHO
aURiZbVhqmFHMU9p3NVdnHbjhyv60OFUb/TBGdweV07KyctHWTDVP8pe/6gWPyeE51Zc1qLUaFy2
bRqCyEe/VpY0ACuDlZOmoq/Cer5g4GO2Zj77Fryb6MR1Y6jCtizF/OeFmDoS2FABtd4JYgN600k5
83+lWLDB4K3NEBdxMWJgtKxk0UG9y73GkIeoUG43oMBJXw5lYxhpCgMetIrqKjKVqIEVhXDnYQX/
1wULusx1/VRbMcpVR6KSX3NNZRD6/okSstfbkW15RebvEzvsESnUcEdT8sqBzD6HBYWvy18/PVJz
M2SWnoBItl3AUYgt2yvL1On+gX90o+e+sxdgpqw/QFQS8QmUNmr3xcqnW+wFRU4lmMXsIMlDUyjz
C0cKdubfIejNeoMLPqgRrahc1NnpiW24aDyxc7U4zDskWlVGCdetNF/i+IbneVtBcbAvmWtta91z
JPeEAKyycz2Lr+vILpPvRZqNuKa3D8ksYTVEaWYl6PgrT8BpGVAif+hDha7HP8PCbFHrn30NVb4s
QeF96d/rcMtItxB45h+jtCnMllK+MQlpfp0R07B7jTNcwDKCxVBFKRszWM6MhvP8WxFfy267sjVi
wCw010vWehcAM1rDmzfWCCZ8Y7HoWuFd7LaoUpCWwb3xC+mXfrvAGyg4ilVf+Z4KwtaDWnrRK4EO
WyIr0xM+R5P04XV9fRo/wQ+JWkRjwZW/bcxfBQjG1sZKzBRysfzu+0/VM7rWtzAJ1eIXX2NHBGUD
AadxJcYloZSJrl8kfFS1F2ahv8PoR9jKUpTQCN/cCoarYzVGTrg4RaTEoxos+MdT/bttErhrJock
QHu07hfcHEFUcapRxazdfs0ckIul/H5GhgxHYqyi+RCqeNq3e/pMQEulZhmvnvbUndD17K9nsRLF
dgLjIfjKswtr4bIykRdX2dqaIkFiMyYhcsU++WRL8itNob4idOf8q6UkNXB6Kq06tGFTb00jhGSW
9Ig5LDm0yEW+wxUYUokMRhdiZgT0g9TXAABVJr+65gj8y4IoS6PQpZuHQaUA5WlAwYD5rz05LDQp
XtpDYiZBE6W2IxfTRJ4TrVje0Sw6sTfi/mMQ44ZfbdwYGd1k5G5C92EfVD0v86nQi+lmcvSuiAUT
d50WgKJPXYdF8vSwTSHbrZdgGRxtNDMOmK7fb4rkVY0u2mx57zaYhpZGzlrMXN8Rp4uFarfTSyqG
o2USC780MAYRStpHfnISs51T3rX1/jDh1H29VnYjdwXn9VWolVQaUaX7Ld0qjnT1S7LLJ1rUlSl9
qt1g36jbZBPwL546wb9As5DqT56XFPPqXv53KqM9Raejilh6LfLfQwVP3u3rFJzi3Y+6FaCQIW8F
57hQkoeoRJ/d1JQMbPUz0zFhXiZe3cfxVEmdc6opuburSOOPsSw95TRcxYhpS7Z4vYXRXFwKGzC5
26YGV7Ela7Jgp72L6QZj2gVGHHeyenKcHpZLScRd9jCNpnXyucguWda67/RX0c4/QvNxiTo6bSpg
NHlh8uhkTxSMZQgtX2KCUNrh9qdPjEzXgjydWkpklCLQOhX2XK5UQEnFU0POZsI0bHYk9F4OJaCp
kMthtxV1BOCmEWfRHhuRkb2hZs8yC61VxO7mk6gL/gagzMKO+/+zp/ZWCAWLImzuHXo8M1UZpJdD
0npmZFrZmoSu2GeHdPB/3crj1aG+9sC+qw1076mFBrfvXvlpP1zCsUcZtt5SGk+Z/Jblw+9mpC3T
lNzSIbUGiY48g46YXqOUkXHVtYKsZY3SMT22eeWLPaqsQh4fIMQju7lAwg5C+nSvlakPtFl5dwO5
0xQ517J3k9Zv+Y1ogwzZQT2mqvTjKM44sNxs/DKFiphn/8tCksY0JSm80eExxv5fwO/XPgeVbrlM
vleJP5oZeg34vcKYrnsMZ//TWbkqq35CUOSjEk49cflWrG9Oqp1Fw/lm3hTv9i8l1fYreLelO21T
ItKzxVZ4hDrDNGFnjJWP5SUbi5atT3soWWrUm2Bx0q5XT+VuUNSoHEgRHYs9OGEsNxoMHmk4Wxot
cTEdqEGSctqMdtCjMjK0kMJZulb4cVpFUMntJRoWEfetKHtczg5kVn1f6G7n7SPvcodNVgzSZeDm
bW00VgQc4G4JvnJJ0yPsdP2+xAkWl/HE826s0qZZh3v0vcYDw5rIyc7ghzm895+r8Wyf0Q34k2N9
O95z4Vnbx+P8vI2e/cPEnMG5d9sCkDXTH58VMXUNYm6oZkHD/CsC+cn1RiE/2uXr+CY1lNkhJbA3
0BWulGGPR3r0UwdiahNBJyMU/Y7kuUeM1iVKK5yn5GtOEAkJ3+pEK18TPVSzQcgSXjfmD3rbr/nN
MuzIOVUyEjbl4Q37Ge4dUzTs7ro7VjWWDwFZVa/Zo+gEh0Wl/xhzWgdgmJbGd4KsYwJeP89qJIQg
eR5DCm8a158mpnbjY1+xrbrF50rAszuYANlBXN4hiaUFRH07HkVq4b1ETOsONVhF0q6PutAqO0MM
d3eNI0wD0jzsXOEz0lINE5E8hvBnaFZ3bmNsTRndqC0LKVg0ql93l2j3cVndgVDvDXk3EyLwWQwE
Sdg+g4vpRZ0R9qJ9uq+NfU0QIARmkVpJykTGzYz2ousq5//f7OoUgLU3ej+l9ELEEyQqkIDTR3rW
Ab05uMqWdpkLnGdQ0cEoV+EecY+c3o1XKcEW+DDSHa28eqdwgmd/L2wuLM7irLLuak1foMPZdC1A
akfBIIepu2PwJkT1OtAyZcbq4+h+QblWGUllEqmaVtGkBl1WHhCcV0mktIEmztZJSU3/WNboq0mi
4xcPvDGVXrY9bhPFtOm2OUFyla91Dyn+8pMBRZJyqmUkN/snzZ/hX7JSjkUo/ZWqzuyEhxpAD7Ve
ufiSwy1jJ05c/BtUT7Y29mihC3CBuWDGCPWNZikDL3Lq2aLZfoNMXrYvSzb5g5IzeywMtd0CdJbT
U1sBaZ2MSwr6HVBVb0pK2hvfyncCn5x2aC7dwY/GiRhLLaWKPxn6yr8NQ0U6XYW2iRJaWRlszwyc
sguYOQnFNH2pQNThunc+4FKULfB71+RzEb8DLS6gCGs21ZyqURpY8f+wbGRmNn3F/sA92CduwaRS
1bYiBW6jfBw3XWFueOzuAv9rWxMkrrI6UINjKXwHOSIxz6hqof1lb12RnN5IqhgNPjMcmnwyK3rN
qIi7M22lPpYq+kOM71E3eoTwqrbLm4pdXxsVGPzN2gp9aQRBLSl0evWxIQJV7dVk7GqMn+BcAbW2
sihqBg4wf0Zcv1P9zaM6z2NnbVw4E+2npoBPtTk6gfmMPkfwzrWTO5gC2wBxWBAxI4J3zjhWILqR
/EcoNK3BrmPfbfDLFJsA6AeL7kgTDZpuN050u2wnA1hIEmbBQ4TlUuYgEwMO3JgKRfqvkyYi6vjZ
/0ZgAfJnwMQF6Bo7kMvOTwzCiHhezZuKelDQRLbPlyxM9XQKcMqAMpeB1mRyVAsmGIG8kH2mNgBi
1m6hU2aUha2tHrw9SV/JeXBLRJWyXudaK3oQOgm7jJren04W8K57TkiBUuwgDRiTlbkNYnm3vVNW
Y47zArODeUpBgJsVASGLdP8MPH8agrQqo/648dKYUah+E15QsNwaWez7Hi6fmDAus+ZiMVtcPN2B
I69SYJmMyu+zhQ28TRtqIAcJoho3gjQrx+sjTcjj54ATgSCx/yeO8qed+xDuIxX/0N7tTwqYZVad
JfRuvUnn2FPbrFYsrv1+/u1NT0ONpFedkGXWQ7c0RcXh6vMMUxaG+5ps1kXjXXliKqLV9lYlCA9P
+rURMh9UzzHp3/pEao4sWgO9STffy4umExJWttJXLDeT+ZkdPIgqI2e/4brpvfAs8+GWs9pMm5gE
dHPrAl9IgYXjSUFwftLww6ajWRvJVpLDFadRGfsSNEAqMrYOb6KkbKPzHqejgu+jx20mpmqp+33Q
I3VBxj2nmjxI7GYAZlfztpJEZLj2G4T5JcM7uWDVDlCK+THV7v3/weR3Bs+aoJsaP8GBAuL0+4Ci
y76JTEPe2TAIthtEl52Eo51Sd4IsXQIygMhyQdf3A3pMadOna904qLHxPhmSF67vcDfnnJ8EJpIb
WFjrNGBXb7RN/bBUGcFUcfUXCxpMZLJCClIo/kAaDOI9xK8H1tR0ql5ri4y5iG05Dxnntal8cbEB
qSu6Ac6NZtLB/nTh/T+Bgt06vWGC7jC97iA5hJIFJsYuhIGbeN8aRRkWJoicaCkVloSqpG/HOjHe
OHLdr+GJ3QLz5LZQ3OMzqMPU0q4W4ntl2c7fHxWm3s8sbHyPSHUE2EyfcpxxoAiCbPH7RC8v3XEs
fFf4K60r2VsQ4kWB+HlxGOuC5hUbQodtsfGdND91jOC9Hlf1xJFDBYMhfOaWCFbapehwWQMYzJS+
eB17YbQU1GR5AcKIX9w7RuxEWPYzseKg4et3TTTJJUfwSoZkYYLCM4kDT6pmL7DhC8A1HF6gJ8A+
p9/PKRPT4B3m3bBjSthDbyXI88/yt0nY/IuOBYChjJxEJNbr4J+EZCxc4ME9XXHDtyvfQaCRMVJ0
d6c4e+IbjM/pW83ilP6MG2DIh9R1jIfbsfrJQCOqOkYFNA/PLjxxEOpyUFgwDJc9pPoqjkT+SACf
PlrjL7mgjoZld46YbiAxIxol+PKGx41FhMn7JgxSt3NsbodlfMeHDuqrTXrfm9K9tW4yW4UyaHaO
1VzKJv+eNkeIxXDg3FBG/q9LURWbAC0e3dJGbD6zhxk1xzX4KrYxzeE6INxkmAccXgRUXt9LdLxy
Mz7HcpEItcOQeg5FKTND/LygbYWoXriup/WovaRF2xKdmsQ2LCQLhn2J6ZYCobBzOxIZb1wFc/eu
JEspy4B69TYde24NGXqze+y7o7TO0eEjkL4osmphvZQnOQXqF7iguyur3chQzsom9DKwauiH72eP
FaWwIuYZGMGw5s5c0PeZV+gXcknly6e+kk38QQJLERwrHBZRFqKqLPBvdCXBIFPAxBASmRDGxJTP
aIPuVJIJMcO4zt11wni3z8fFOOlEg7USaZ1bAzapWjq3/5UM0X48h0aquGJp1m7pHOusKCI8fF+1
0PVMfmywrp85YvEjKZwU4ijTXymnlepQLM4UuUN9dl6F2rs32+O72vPJLNvV9ZeXVIJrHlYZ1fhS
rVqFFK7qwdlLkrNe4Fs/QXipKQzWOcJPwqDQER+xuSyOqVfG6MIQNsY4dqkq0FTa9WLd6Pqr/8gj
9Or+ig/yIQKR3QAPTtEilqjFubcS7b5BJRDgFvusOSo7+PGjTDI+nXPirW1ajl8zjpkggeEUcrbZ
Eqg1wU51ii3iLdKy7WgXBviI6r9qwZB6O/9HxnVuxCKbDRCWZLwUPuXewQXWTa6DWQcTE1c1d3Fk
CPtNYNs3d7ega8OynlT6XvJ1Y/waeW/COqQj0F//HDojWFmOHIkwhmHYgQqJrFSpVvBCLhcBg77d
33ddQ8OQWgpaH6Ud37Umw2TtLoZGP6nhN0BC91FtV1t6rxtBuYjFhCDTMMMPLOM4mhOKgSkNpUNS
DR4C5VHwTaInl6vildsci2vhyz2efpo2gsCyIRrc97J7i3DL5fD7r+LK5mtRyELwvM+gAGPjnlCg
pp6Zhef0op3ScXE8hsl5Kcmsp1A6rAz4krmU/znPLnZ0hgAtFuk+dGcwQQENP05yPmSzWacUkOla
J7R/EZD16ADObFu3is0BInXxAM4OePdEX8ZnH8hB+595wTHKtsFG/eVF8Phumyctj8Pq13xGXhyV
NUBZ3+2pj16YxfOYaMUMoYWrmLdoxnGb3bLnST5txJz+b351Y/IvS05PG6WYoXX0jC50ELt6HPCZ
x5sSmShzKJEtrQqoSQwyfV1ZRkYlBjSNSHUQE2J5T25R+4RfgxPJEsfhTgf0YA6k+ta2em9IOkwY
W2Gq7OptDgFyCGK7Aa1eI72OKkxp4j/zsRpyKxmkuAroqNRqlIFmUlw2QN7F08gN4dyxRzYGQUK2
dvCuPwBwRJm2YHUkzdfhQL8owGHlv+E/m7F0wtYitI3/ZWTShePTjZPPxyxuyFqnNLctohqhO/6u
XTPCwDIcUM31byDZfnRA/EQNBb6BWwjZN/acuzKwz+5DFZI1Vrvv4FKjZcDXGhX5nj5K6QxP/JaI
bNlt3JZJEG+fHVhClVVi0x9Tx5krNZbx+/gtDDXDT5Y3sPRJAJCmCM7S5tu4uKHTNRtZkbjLz7M5
t0+7Pb4lg7plrQQ1mvW8fhJRK4pO4qn6XcG4L7Fm/LaA4d3EXNwcgG2J7eHyUdytv/TxEQHCT8ln
qKAOaoiuncpfR0MN9n7Gq9sBl2dP4EkU7ieF0XZmeBCaJs0ZjtQ0Z8hQHVM6yHbNaJ3iWxixyXWx
/nuuXJzyzKjXEvHRvyhGKFqdCC4cZk4Pw84IQLCHPPmBvz/cHadoKLhkPava1Ikcfn9JDKAqjl6h
tNTL71Kk9oBQMFAMfXR1k8irmGWXTsLbBfu8UQ18Xj6oXxoGwHhH+nI4JeSVBLdTu26hMa8IHCZP
XjGWydpitNd5DPQKx07kGnOGj/BC3g4+USnNjoAP2AGI67ZGWn1sxCJYWSvkZ+/9B+k4o/q6g1ou
NQYtIhPMjGLsY3icR6/ShZZir0vKxvKwcD1RN4m6CEaLRJuk6F72MuUagr1FM4IQwgH5zD8M/etq
lgeA7D1EWwWI3oJQ7njFf7Y6JzNwEw+52+cwSjJ2vZ9zkEHf0lzutOPJlOFC4Y22vIwtrfx2Hf6L
9U7/KZIyWhn1FmCAjS6faETP9syB2YZSxiuK4ECWKYwKGAzf0cTTTuM3H6bU8dsGlk8DMoCXdqoE
XpJoiTrMw6+LzYe7id4hSr46fb2bKHXyi5ZZn1tGQ7DADBwYQoIPSpVezuuXpDvhqj1R6Qmgbwmk
XWhansUotgy9swqhuj+7lYl/dYeHgafYvwxh5ZD7g5Ms8TTB+DrzSxNj8OPSCLaTg5O7nvqz2HzY
vr8guJBW6QZ7MP+RzcxMhmDdOBdGuQ4peMAl9xMEliqOituLNPEnoh6WSUw768ammsNJ5weqGV7n
AuXMoyWzm9xTBMMAheS7IAUuz+Z0XEktkhhPX08CsioU4L7tmJu2lzErhcp6tOLEJ0rXKLS+OoZ1
il2txyb5yHAczd7dDXSbGNuRKIo/Sr5VD5dBbBGbh/UCSJ4LbMe1CL0NkNe56gf6PkF1UNjOHfna
3waQt/G89jIof5DNDlxN/+ChOl15/mk8B05GeM0EiDAs99GZ40A0Ez6VGVtNHPjHwpshfLBz7G5h
aVEs7G8G100+fwGt9HLYHUWC8nnP3rbEiXm9GjRjfUIXlJst9PSMOx0Xekf06PH2z5BugxuuhkDR
EPXVPUVLvkorbqJzKvPkqwKBmONx5bBG+fCDLFXVXXC8YKI1xYKW8z6wzOVF/DQhhPBXCydl1w2c
OLnBcut82nib+9ISl1Xl2k25kebR4m7vOyiMt9pX6+ks0CKYtyHz5OhSzFKNeRzcEAfLgfLME19H
Vh9HT65e/OkbyNkPznM3LHZz/Xx84R4xWhRu9/iA6hrX1OZ3CFGujEL8sn9GZQAFSML4itKmfa/0
AiK3Q00/SRnQ6dUs8HO8pqEqy3JutKsAIl4uu4m2La6B2CpI5t8gIEiA8D/U6UHb5O1IILp0qnrH
mO0k2eLmrgBAgHpFhCao9pBqZzAH+IRTpj7Lqxo1dKbeysel3lzLlTol3bbJWulOqMCC8pWHnG+L
xG2O5bmwvJHls7wkaxWZlCUiK2dIezr1/aExWPKNkfh0mT2O2wOJHAb+YprrMY3p0D8hlyeIRnfs
cfjxq/zB6ZXT/odjZ5qfQVTxF8m8RTA+Sy7jXH7Phy8MCYbwOcbo01QFUyknJ6Pn8fIvAMQQ+VrH
fmENMUZapCBXwbFc2Tkb06ApJE47rst4FcFqWc/XBBwJCIu0ZAVnmxJhKn3nZyZk72FGzll3yMj6
uh4mw+MOtJf/kVBFFYNFSftmeJDAuRJGYzcmdWgAKJA7TD4VdPizAOPUlQ97lr7vMTZiveqUwi+g
Xxk37aK0mTaKL6VfUFAFfvxwDXeMWZX51fIZWVewsvTR8fVe2UVEmdig+35XPD1FX0mNWyBwlALN
Pl1Dk2pCsI8wlLzlM2YEPxgiZmFkXwVsxCkKxX7NUYzjHYy5v0HRBw2GAnE5aTMks3zAAgzYY2qc
xzc7+FTVg6AAwNk8/LbdU76M0/Nfb2M1HJrC3ElfnP5PqcodS2dGk51WpH9imVxQ2hlU10iSJRDj
oXge/SrJjEs1MvjmR0YGAFb+y1RZc7P4Kr8IjVj9la0yKxdpgjs+nlnNtcO4dgp+afBU7IT27JDH
0WxNGAWVwgZiRMbBpyNCo343BrIqF/KXTAwE5TmcOZx6AdXns4DkpIxZQKJuMU2qKBGi6c5j1Yic
h9bx/T7uwYMTzd6Rvj6HDofHEUDhmcD2McEcJb/9J1ihKnOpu3SQE5DiYCL7gIdgP1Y6aMUGbiQE
sfjWyGmmp4vMacDbqFpnGTwHNxe3Amovl/yr+8N01azq13MbWPuZj0k7g1mSCPCYe4EEr4ispzlF
7VrlAmFneZ5STGXGPF/P48sQoMM1uGbRrkuqzvai4EHqtP0uWRDs+wiKUmtdA1kZwLsh798Z7C2Q
E/v7tQkbXpVcz/Q99L5bYl35H2DgZLf/kcz4nTmVFb3SWev3aPscRL9HRWcumRfzrb0fo4LTN3BG
m7Mn0FyV/kMiwSo7kdmI6FZzC4n+Grc+f6fd+79U5bXRyxmjCgT/hqEDmUGKD0oAY3daJqybmqAG
S/VAl/NbuEocBX5BjHKgMyxrlbAO89xZxBnXyRSLOMOqKLgzUM4apeNiO07X20LJiMI67Xg+EE/c
AvOT905iJLrU1j8TqescECA89S716gN+Jans+Av2kKEKnOaKPXaSWPDVwR0bVl7svgCXLGo1jfPM
nwWiJfDau0MREb6ZRuZ1Ot3l4eZ0ZxbQgIpX46VxaT2GItUgBgQJ1p0INmYgzi+50S8c72iBgbna
AKT861ZzyYDk1iy7rSt0I2Ok+AN+oYETbcK5bOwTodERGW1kIpMpf3FKOYLdLMNAXhH5PItQ+RSg
9mlTG614o0FzNH1ApUIhqtV2Qv2HCdca7ZlEzM3AOvzTodKwOzlGCrQW7mLVHI9twmnjIBhJHwKH
wDYfhiK+SMpiiCCC7RebzmpDHsIdhTRGFciUdSwssb9bFtJUh5pGuovm5gjPsgvxs3MVCO5oSiVl
RREhxpjDiVUd9mLS2QKRtoNx5U/O0rC/ISMkuTCOJC6qgSIzFI71mMH4kNn93NbHB2HEE569IY7H
4EsHyiRoD0lHU/EHt+K59DSySayGgmkiIpiRsiIfiFYZdlIfH8WgCzxI1ElCnOMdZzT9WGrbJxsG
cZp6dS5UOTnqUu/OkOvp6ig8bZvFvx/1ovslAqoMLvZFrZ3LIfhKmKo6CEt+PvU+q90b2aWwpY1g
xpjMZ5Vg7tPAWWjBxUJpcX/+m6rcMNWdlGtKnmmH3owDTB3lzgNstWtjsL1VhZO1qivhl2XG3tDk
8H0lbEt6y+Dw1npaZ6Zb/ZV1zSsjM4FTc9rLFB9GOyQnqgrKAYi9fW3m4qmArCdEYcqJlJxT32dT
xjd8QqRUQMsbK/h8omaJt9wnYEeOZj3Rw6BTozP3ncgdvkgwKtc8Sg3TQSppJFu6ea2R0pnbAOHl
zgbAPcQKUhOW5DRThe/5XKXj+L/Rjvjv+1nMPB1prqQMziYHO0RMEPy5gdDNm8Zs7sgQD5vTyLRt
eGjUOcv3SiYvIadbZyPJRfz5Up7fFezcB0xmPePezflPrnnuWlaJ5yWilN1KIHVtv/qHosrH10NE
2A0YWk4skArCccDYjVNow1aNfww6hY6cWa0dzCCF8TDo9lwwblpQFIwbTq1b8ejZ5jmDcDsoL4Pe
4Kzq5eq3wlJXYmm58FqaFV+z4Xpzl2xe7wln6Tpi4KxkU5p2parE/DfG9r3UipW7jiNKztvE+Ww5
XC7Y5s3W2NChJOxpWHTQJpJFAO4AQWHzpaInj7bJ7GNoqcL8K0DMWNXPzjGXtrQmJAWEASmIm4vx
yxeQVM0iywfPREIHehtiZdbafCR37Q7P9+zqBFDe4CoWzJ8yUss6ULV/860GtAEuHw6RtKH1fZCN
EWEU6nayrXDdEUMU5CbAI3hZN00jAaieJYe7rtZGcUk1BCvhAGgZ6MurnbpLPtiNfdk54QdYYmBj
ga27CNbuO7YI6GIyu1C+XcFT3QaUMmPlnKkCt7av+bi5X9JtJ7J/teejM2ukbrgIcK/1munW5i5Y
xitAEnQQHC/ARsNkdtxIvdR9tU7XdCaMfW6bzqep+7xFHPLsRmPP9xwa1KDIDTOhf4mpHo3ObDly
Ew/0UIFgD9fHfLzp3JZlJF0ICsmecXjKbnf1lQU3/rbzFheGSSvYo7BICdtMIfy0YrfVNxIy1kZC
qFLCk247gAlFfVSWCmDwntwrW5FRUi0cTaHZYfT5Kanq0EX11iDbbvyre3iTwTdUslG5k212UWYH
bzNgBQQQj9hD/c9K85WHi3lNVY4rU/YuUltjGNAhKHJMSzQLtWbbUdyRfKhHlShp9nT5IyRLsMcL
Hcm/tJTf2fyWxXzQv5xol1bDHZI6XGpz4z8hdGUveeExzHWg6zEJRRkpbR6zoHM4qGitDfihF6WD
D6L0PiijC+jiLJC3eazTy1yQmgnpxizF2tXb7NoDun0rUjCwJl9mkaTH0V/uISlk0gAHGsro1FGL
daGDC52X8nKuV+1YGsoNL/qmGa3Z9QeA0AizpEMHlR4rmdO+LxskiQpIL3mKP2lFzcHobNE9a7o6
OCHaX19jEdiSfhgBaTNOFvjrmnJLFQT0uCwLm0xvFB5dY6aG2+iGsDCL2+E/Eqjj86RqorZxhECJ
udnPXLGNfapoA/6BzLbb5nhFEgQa4yNRM++Ca4X0olNy8y0ppG9yN3TnEfJlrdAlgFibA9oy+WHi
oAjuix5rjhqjYqAbhUfzpyc/Lz6q12Y/htUluYpO1loto0lNgdbwp6u5T1laQ+DjU/YnLKV6yK7l
dMlm2KzUFfpVtGp061iux1OmdTKIUQc3C+DzQDB50B7vsUZ07D4zbYgNudN+6DwaCi+c7pQPaoo5
s5CLFbQPAL9ijun4g/t39u8IldsY0qgv+fRg9WTYmgAM0UWnR+vLpDxkp5qmn9LnzY1+0BDA0DP5
X4z7m3nR5/ighM7viP1sDSe5TKPMSdBnsC3OrwKbZrU8ZDQVQrpBPLPzA7ocTDZ3Wr2/NRQ2SLQa
WkgKju6A446pCz4w4WQdqGrEoUFBlXrrMcMt7mTSZtaDyLqldqgDjA4SbvfZJKePuzFeKaSal1j9
VLcCF+lTRlAk7ygmj05prRJfgV3Sr3KLGh6UE3SASYd8ZHAG4oWHKLyfrAClZs5UHdkKw0R8H4B6
pYe+jcx4nfJmv6SQu/m/47nTMCDSgY5uaQ0ufSx+N3CWECe2ufbf466hgyRL/2G4iVi5A/xc9dZ6
PuUxfGjZYpGj390s7WxU0Q+5byHMrDE9z5y72xfBt8QuHw5DwWIgXzmAOJpQIppeYZY6FiCW27O1
Gv/uTvWz0jK7K/BrR8FMGEQvtclsN4FTm2DnLRru8b22Xjlj9nml4g2LplPg2Zy6UvNMpSNQwgzJ
4OnbCfoIlNT9v44JHE3LpCGtVlh7SzTYrjRmWhwbxv5gjXwpc6KRiSs4kF7aM0eHdMoS/T9CObkv
yq+lh6sihX/WaacMyG2BcV/BkkgpGiza3BxTlvu80TaBLLNlrNAgApPvtV+Fodp+2CpRSo7S1N8p
YhgGKe9fjU4WvXTihzaztMhdc47ldyiSmOtty8VNnZzh5CnWfunXpq+hUJr+eH6blyczdgB0BqH/
j93gV6QFn1+NRVC7ndw3KGR18gqY25aMkJyHwoYCjhZB2DGWyyy6kJyOdn0sKfQoy0vpTR7rfQ1O
vgi4PEObsfn/CVPu07Omk4VeLj3qj6HstKDQ4Oc4tqwFnur5Q7MTFEmZWJ8CNLxWFcQazcdhhmvR
yrLbtvfpMq3tn/PDIgXEaK5ACezMBPNXvP8HzqavZKFKOIINaTH5C9kb+YHL9fXxl9aU9pUXHn6K
yd5VvUFRJ3LbvFtg4Cge5F/g4edM2l2+ajR+nRpPn13mbHLowOG2Rkk0S4RQxtgSPHy2CS2SKzhh
Lk3ywU6i13A82CcDzJTE8HieH2ewaLZySpFTIbF4+pK8xgi62RjrBu/vMoJ2Putaoferk9ddf5jU
gq7IaCT9s7PZyUS8r08hYa6NVmce9rPTsP8sRk+FE1SRysftvYOj4ie0E70bKV7aBg3qhSGqi9kw
zDv9FUn+m40GXrQZPrVGDx4z4UD7H0xuS8ztqq3QRcgp5/Dt2qjMV1rZ3w2ZK8SaXfS26Sddnc7k
zRKVgQYySvi+HekJW/mNpwVSIeubfD4Rb5hAsNLD/phZAoB3/wr6CK54l6B4g/PY+4y3C78XA8sW
7veo+6x0WyPUSrlSagmEHJPC6VLO69djyb+hvwx1o+7w95LdpBbtOnhiS3OnAX617W7Jp9xtlSLk
ti4TL/8g/BcOkHUNg44A61L3NkkkaZpy4Si1t57MAgacfZQXJgBW9Rli5lg/bwnu87XJiPWchcRq
jtFN6PJLM5YBnN70cdzIyNHA/updJdfd3LsYluc0SN2Z5ugEkqzblKyStBP/5q+4RJGKNjIknxsW
9Hbv3kQcHnZ+oh0JYXdb3/bYxgWX1/fhOHzaZzn51ZHOCJAM/EWoDuZHfg9VZa/tcFRNnoslSOow
ESOY5F4xeFh44Qk6J7xyq2+0nxwsxjCNDaGk8O4TBcdT615IK/AE7Bhwm/+HtlXS4beE8Vxvps68
p/g7jBoIezqBwCLkYO7Hmz9d/60LC9LgsYUv1Kx2xC/qTEHCZuPhWfsILKZGRUTIkMnfoCwdpd68
CBNS8mpCNkRbaftnGVQK0yGWTNkoTk8xTfLMAwJnHSI6uUlk/Iwqx6YFpHO9uIafgXVbL2bm0Nd5
EKEb/wASBFrwhqwxWOcrWWvqISXGu7TAD7x3hLWc93jZ+JEv0K9vrOWE0NJp7pYOSfr6jKwZJmQ1
qyy0IFuti6AYz07qX09bLbBglqQVU1czxTKK5507QChhXjaXNskOZAS/ZIJhxjER94HbY2EQXXZq
OosusjbOhcl4mjBOchxMJ3WkDYtxx8x2+Eb/2jWixl/pNtNAyArF0ZBCf2nzW42R8GfIJdtpwRD8
BtsoNa5FLalJ7KSak3FXwZ2jc5nqAIJXVmuvLqVit6C4gYI+GURssAjgyJd1thoF/azf9aO7uckB
WSrbHI7OjUzL3zrCfNBnZFhf7cgC83r0g+fsOEZD/JcOurD7d1J6hbOKKRpTpKzC80nX9Tm351yJ
wRyhIHLGl3krOJDiNUUxFOsG/SlX2qZ5NBbvR7l9rDECvDEYh3XYYlPdUzbq+qwXwNDB8E80xIyG
MrdRZ3gZnAKyXTDNc//7hZb8kx+YWY0jjDhXBdnPP4V1V2Vd2RN67N7Kfcxe4o7hbrKYkBAR5KOU
4c3x8CMzMFYXBSLlvUbvmpckwL/OIKpsVCsV5k07y2hzJZvjuc/HWzqLVz5PGMB20fLTGO0dCSBB
puFN85tf1rKA8W008OyR2p9ftb1GFKCHePrKJ5PHVOtgyCVO4BDnGuAyEnfI/Wvb0gKlUt8qzhOn
9qRBAYmWVjtx2+Rpg+C6vCsDbH03YOOqafjB8ruGqRt9LsWK3pJAG6QxGIxmSwC8B+XFfZLS/7xv
0dpepB6viGy4jCdR4RPleam4xrrtYCxrHZgWOm7GiiD20ftWac7jkORFwIXqbZUq7u6Ug/gq00cq
ow0aAO7u4q5HOQ30c0rz1tnwBkSHjm5wENf+3w2o7ccCr2SUaZxhoBLCZyFV9XjixH/HKmkSlYq3
mJyg0Ef9ZD/RVJJft8f58adOhaVlIdyS6EXwojNaC1G/bvTj0/Rt0H3A0+DtW8rp8LjCdlFROhiM
xJmEi/LgMNZeKUugQjed0lBlrXk6bbXkd2ykjM/NTxgtIOE4xE/YpjNg8TCIZF84wBuWlqrQGRaA
d3oDVgkk2Ei6HJTSRESXOj2IgcNfsRFj44majk4wNkG2OivEwqeVs9IuNlFJ6NpE3SSPuRV4/nxw
7nChADM2kR/DxyaikHRtD/wN05Z7qEPTCe9Da3N+ACwjQpB3RB6HcVVdGyhjcoFizaJDU8or/Xnz
8Mv+AaQbaQd4bTT5fTXhyz6P/ul0NTuRrA6ppkioxji1D5GAib6vYv2m8eRQp2VNOdaIB/ANUXeo
vCBJIjycFFHt6/orCRcPXbhHOFMQjpiSEmsuOr/edufzIzBdxhdagW5ZZV4vARHHJLe/PiDZF1Uv
vgU16PHqPN7oabiofDBBRhreYyp95+NGZMIOkeaNdL/rRZ2gJw0QWz8bgWMGgCMbcBJAQ6if7sCo
w73pTciPAtX7YCnRA9lLoU3I2PuAoNzIS0xOuO/CcRI1LZ2cFqEvmWuHxtvP84myrulAuB2bHkaR
0AwL99huFL2ClguVtqPuHXlyWfR9ARFxslhrOgJLTvREQ///wbyrh105hdWGCle4BpotQD+qT3Om
NLO6Zd//LmUtumVNBps31QfIJfSJ42C0dgl1ytDIf7EhzSeKuMkaXbFEQrQEABtZtc2mA6nE4gF9
bgxaD+4ENf67EdrujfDCit3bsZUkHmwM6Qwk/i/5rVkiGQglnUuAKoB0e6T4sd2Bqsx6enVXnLsO
PmDKS1Ahlt81OhlXBnpFD+qTILH52FZ+ej0S2RhQroO8LF0vfgToLfNVLkWtG6IRMTTtC25F+lqX
1JtXlKaWekC3J+vgqhqCfF0tfXn7BPD7OuqshSMHwx++gTiSRRDqi+Apl/sAhMLUdBOgfVBb7afz
OlTWO9DCAQ+djuEDhIIjmQ3CcpFeC+jFvigJ68MrVx5Y7rrOLv6X4zzU5VX89AdIdbPiuxYQcZhS
7Po/pfTkI8CfpDKk8CTwWfVEVjfBYNnFlbPe/OC3Wj4b/6tyhETnI6VRgXmd5tzMjhbz/qd+mOSo
nBvhApk5RSwjNKyNnx0Teavvay+EgKM12+Nw3AYtyPoFK4T/2fBdtUPcvFPZm+8PFg+lSTTQDE8F
KHWfHH/mHJmP5sEEpqDqPa+z6aWuQA2xP61mI0bWAWWoCgUHHPZfp5NM8tsefffjvhbDvxxMjNYP
YsYFaUb+r02ZJLqmL4pnFvHXM1sRkmR8KxtEp/t2MSV1cwmxMKEpaaz+e3wVInnG+/DHpju/+sU1
SUXN7NXfhqED1YCIu/Z6uKKbYH5JtUpnQYcYvhcvpU6hRReMXickJtbk3DP1LKJmAD+QthSfvfyr
gfB9W4Eo2/2MasxenHwMvhNoJKdXevLGNfVkgAQvis7y8MRQt6DqRz8WQp2gBfQkbjAaQf3TVtEm
whRyUYHOe9VctYJTBCKQlQ5BjIJsRGL4+8PYdHV7OhbJyoKfF4o/Z4Gw2j/8VgFHKZUrYw2Z8K3L
/BsFJNMeRxtNf9x8bW9YNkAZaHw4hWn9CcBVpBG9AhIlbmXSCPQoejzWBrSqhahJNHI/QDUkdnS2
W3d4djMWie8iYOg7t4PknkPCDu4UXvBM1kw/YNwI8fV2dibogBk9bmBJ3onZLPuFpKTnuk1XZqJP
Fm1HZP0lAF83VAKzKD+LaNJnwCk62OnG9xKMapZ0OF9y6ei/RX7F+PYlx69+PkOgTv4XN4bQ3LZB
i70js6aKK5VydjVIkx4t9OKGjvtWnqTInrLRb0sqRwNJk16fl/xSGOTx3yav0UOqPmCuW8T1oT+l
VQOtt4sGXJ+t5k5l4Sdyg03daRUk5chtfISSCvy9/Iwx8lyo9LOyROpMjuMvP8PZqwaixed8PTtJ
gCycHDemVs7V4rNflvS/jB53I0uaA6VbP6JzX4xaOPUFn8yXFMHST2zvwgL7LFtJ5QHL+cwHFYQr
yioAxNSiKV8retvWvIOYDxuFjnT5Vqn437b59EJ/bhLoMmR3syAuXGlXnnTxF62esWEhAD/bOAkI
4dwFsVgOxGqYL9UX1BzJ+Q/oyIX7oYuZg8wN8xlVc7LXmRtncEkBdzoAUMFaMtXI9+LvxAbOsg0j
q44V+8F5QWE5JesXRADOGFj/jBd9/zget1hsOKUawEEDVTHg+WEb6kmNKRbEKHl5uVDBKuAHEfWK
hpPdVN2oi9zJorm139dcHicPncT0AMbblSXyhfD17r3w32GaS6Ymfs5oTX9reFVnhEueZ2AUcDyW
p/Pav0uTXytFPFzAJVtJSAMljTUWam6D2oe551hzhaAB1RRE4iWUENLV4WrH+rePWhOz2b3WyfYF
Trra3dKYi0mCCxyiPrAfuh9cuTZG0U2O8rslRZzobW9/HxNKVRKXJ2DlXvSNA0xax3oJPJ2XMsVh
h9t2RcgUawoaz8wq3Z64IJALw+ttLdflGSopJZ9s8qtZWX2N700L+2BbhP+avlLoIBypybbhOB0f
Iu7euVVvNUGnj9eoVR0hg8H7y/DxQ/38XmEp41MLroHQg+blCvfq84wMzlr+i5P+4uwnQdTdB1xl
MhikNN+Bybmas6d9afpln3dEpZjnUEFMgs3rX1+WlyUho0srMZ9NtCfZRJOdrwY9pwhtnWVzu4dQ
zzJAyewl5bjc5ylS4qkRFY5qoD0P8ivynY6GoHx6bG0dV170O1cKI4whets3csOGFXF83/5b9AaK
p/TQJjagnoXixTWT8FaTsoXqp+NlXOJ4pi+t3etI80k/tuLDYd1+RlqyUcv/j39FiqrcqQ3QBdaG
Q0qfgGh2Za/gMr2FWX2GBB3mN7/bCBG5TyLvUjLL5PmfkeVPyEgawM42nlE4fO6JVSJ0Rl3hZW3o
+rxJyvLaTR86jUyvG/FPD2khonHIDdGDlqiVG4NrPUwYlHZ94mEXXmmDewMlBUv7Az9DjksNNjxT
vcgqkl30VUeqVnz2JsshoxZv9CMwVgf9c4uKdzFFSFJIxYlL2gSiCHBPQSEHPAK0s/XDGnZlK9Y/
zG95Tl3WEAN2XltM0T0d66VHa8CMJ6bWLEBtZ4taDugbLGC1RdPjexMV7Mu/W+BLcC5RaXYpJN0d
HVvYBVwwbPuTsKLzfhTaBM8hvwWlTR/37mXv6liorp04pMhWL7px/ISwlsP3iyAdhzvCCQfR6fnk
Uw+IpdCXWtn3EJNah2T5MNYbe+3uyImuTdtOICvbwcCGIHC8sVHO4WGc4zDeTFdDK88VBKvzQ3X8
jIUNAY4HRw4Yv41+SfPM/VgM5i1eeObNSyrRmAbR8GZ9GDxQ79s1viT0nmSBl4rNlo7Fls/BGvEB
GYM5erY0/J4lVPsnNef0zkzU+UD1vpN8L3E/ffjzCDOcXYdk5uBKsSz1drFRgGjRvGrEq75LM/TQ
P6TfviDVoSH9480m5eI3DWzF9Bj9mnXUBnXJSAHe0EpjHtLZuQisGWn/g2zi/JiDpKTba4JIerb0
XZd2hF86zQ6f3PBS5tvXQWmp4Z4xApmsYwP66vTd5mhMbxwJ+pTWtD4HsOfgkxfh+jDUY4F2QVXf
zb8gI3xQ5DlvtrhrfJ73oJl4WVFzWoGxKMfpdv6ApeOubrHf9svwfKx6xVNjOp/ASyTYiYlGG29I
kOXSxUGuL92Rn67+phTBKEIC81eSyiWEpjaLJ9tTUHkzdP53cIK9s07soB/NCTDEEwD7r709rSiw
DyddcEmiCnLADoqHXwbxpRQAA6pqCQuqeatMIQpbIKwKLFKbT3AX5oTQdJWRGxYBz8yO6D4slSy7
sAWwWPlH8D1pBTNmsumuuUvENJM0/dt5/goOzQSiLLXGxF5tpAj89yITLPmxrw0Oe9+++jLDQcbU
K9szIgYrc5tACnADqhZOezqGqF8mi8NZxV/G1DMPM/D/jdIa+kffUaq6taTuBGLKetl1YWC2h4gY
MX6ay7j6uHuK13gugIgP1Ig/C8+8WOIIJ9jI4U1kjNzfoyjsdTIV9nyr8Ono5heGzmvwDOYeJiH0
MX72iXS8pBq8tlfw3A4YXQ7/llftbjtcTFUtzrOzImp7x9kConG+OrkKUfjmJNgH68SXcceJTjcl
/N2Z8Em3SVb0PAcTtyMKFKP0VZiwadlAvkk7YkMIt1zuVTu+zTB9vXcPj35DOJlTbeDuHR1lwpEC
GxvWb+78+I6cD1sIeRmsR8x9EClEOerlWv+oEk7t29sxGDGCGwZKxrqFdEgUIvAR9L9J53jQ3fLw
uwbZGGG4Wp+H/8bIq/Xf1wxNOFwb/zFsOZ4vpFWALE5/nI8vNY7/NRWSS/nUBpMlzrbU7Zca/upo
G2Gg1Kq+w2uG4x9aKEFuuQibc92lKsBH+ApEd6MT2LPGbd4GulK1LoW9wSiFbhhEaDDLCLbSBMTP
0tBFDvqtv4pFfF/aAq4TemmpRW3lXC8Qbm+ndI7KnGnfRZBKC46hK9zS4cCiDnoGDdcsk4FH9jKx
JuexyIykbsL6xO7KoFTR3/rqCtPFu7A8+c0NLRmdFGUQ1LndTv5ekG6pSqhj2e6PBPsa4tiuf8bQ
flu/QVAIg6D7ylLDShA2wwaIs+ZxroKq88eQbvfWrUmzaooXCgZvjM/Wwm4hEUsbJV8AZKx0a/TM
Sogp+BeH+WBdn3IJfJtHLIURFgkamUB8SfgGwmINYQIga5ou0SRDnGJyLlZ6Ll78faFkt2Wa5Vri
koOUg1KZkqf0yvBPL27bxC8BHXsF5IPdR1ObAyP1KNsTFS5YNK193mzJNlusyKOCzisbF4pZr/vk
yEyoJ16+rTLjmAKXH+rKk7DarF40MlEvUJXHBMUA1ls8ZUQ06lU7DSFdekx7pDDbaJXHw+tSfQlc
W2vo8R7d8RQH9zywJau7N42VtU06PHiDCJN8SAGo/z3kUCDz7qsfFmBumy3HwFv/qPV9M5sqn0LX
Z4VTBsa5rqYbb6eF+N8r8Mi1cUquZGqSF9fl6bWbUMonP4VEzSsNYa5tvUQNQRqkaauM8omDZGhR
gXdVQ/cnBIxM6p9huCx2eVxxVMvfbFTmgodttDckpiyhK/G9dYhgQrkGuiRC06FyMdsoBKkbMjxl
uCxpWLRC7yeUwmela0+LBEo37VeiOeUiO8+OupHfH73zrOXoP3haTyensHwLSuXzDW3hqkH49fNV
/6CxT6bEOTZQIVgPCOfWQ0yG6PrYvxialmFh5dK5AjnNEnN1fBY2NuPHId+IyGLFHos2WTStDdvi
yCmKxaWTMjzyJOYHVupdEzi+LAWr2RxmCndUL06RjfuzEYVMXaTLtbIC2EiYIYKLAJVRSFozx4BT
4EJwFdKhkywBpsCtyZr4NjRvb7H+erCC/we6gAQHFjwuWUKZDF6+MIbiABJk2OHWaAXlgkzseCXD
/f6phluEZo+GEGKNqvW4F1lxWeqjJI/qC1B9IuB9gz1ZmOYp3f872qTzRdwR3MbXiQd1D+l1ijuH
c1Jy+LGV6S4l0h9HXqGy1rqJtEx3ZkuyeBV+UC9kf1oq3QVCWYsz1eQKMrD/nhQEVD8IdhCJKI8I
QA51pKsKE8JHS7wxtjnSApscTUE/4gRG559t6wc7U0FhVTZp/ggR5Fq7opNX81ViA5S6/Jp2ILA7
BUwpuA4omoAS6WB8BOtk/gpACwO8EYMIPK2YYuoU8rzTdv3D/nKDGxVXk0JXSSznMg01GW0KLbLQ
6YNCfn4zMA3Wck2tCAD1t1mH83OICE1YsXVXylsLbyhwoNdAd/ayqTAMgTglAsOV4JNjU67iXWt/
sJ5RIaNrClEePwPkUcUcu/zygZBHJXRVIBUAeXJga43hocFymvBy9FqwLiSZ4XI9jQU+2T4YsAtP
oU15Wf2uLtNHrD0KNOo80ZeXtzhPKWFnsFSjnavwGSX+vuIx9rrqcuDGpKqexH61FXGcEuU5dZcv
WMkWnGbEXzj7APfSlgcHUtQSoQCTwTjPb9JAoPIS+6nPoto4XMJzV4peWL2sEBTV8rWBksPOTIfA
AcPsvunJeMOywZDLSqclIu6ysVyZRgsRgdCDcMpkfFvZjODIBQf6InnoNHW1wjpgDx4HBztemtir
HbNm7eYjsmHknjnuVO9ivXsAgNUItPOTm7l4h+P4CI+fJ0UzDX6IM7ZuVjZCj2zjAtQMVVTcVVQb
cnw4gYamHdyLp885C2z42jAr7j9jFnDcAGgWmeDUOpXBW1+apYCaKIcVC6BbnNhfLsTESDqabTh/
kCPJNOniuYLZDoxy3d+WDLz6glXgg5XWmJZNXE7NdEDEAcddwzEIUgIrUtM18Z7sDw2RhxvIa/yX
V1EUM1QrEsu0UEcUMXvvjFStvz7RPBG7pGs3Co0HASB/lIXixKXDwViQ96snGH3W0b7rnGYkvYaz
Bm5Pt/jf91XMPOxSIkjKcH9b+y6eKRrgelW6yHqtYbjDccSK8m5ElCiK3ww/WBCYtEkgJVjP68s9
Y24hnd4AIxmcaCVeiFNVZNJENE9oir06v3nPsjvwlGc3wv2BnptCicVL8TtKVuIBOun8iLr70LUS
jg3TmbMDT3hGTHpE3GBfYyRij2Y+AC/T8OOcV1k1VbRzA79WVVS0UeObNw9bsOwsnSK53Hjki5wh
RGpqQEm9oDoXQ4j6xtEsoXS3+5izcbuAc9D0Fr/oed8dxHd+k+8uTzoW/QqW7dqUC/eKpadHiBzL
nJgjnhqo0chpq4nlPpjAxrjGQqLen+qSS6c8p8kMtUADBtBt25eii7cB9QZCrjq074ZOtmYUMSMg
hVL1fx73rdLn5j7LIYAmjPftwoHnsOhNNIoUZyK/+PgkOGpbxxDsCJRswiljtzHqGyNCa8F7T3L/
lzuJu8b3ZsNWqgS5NsQrOVFbT9iUOUVSQnwiD41J4ebduzY2PLKeGVFlffiAoha+t3YkEueFrgl+
E2mQOqfp3jAamNCP6Ev6Uj8lyK0Ep7EBB2668ioDhffy/lzs3bHriGp2c3iRgBgwLMyS00k2T3MG
yVCyoGNISsfK2kFaMFrd7NJ0/iDe40lr1hNDGN4anKTSW1XJyFtWfW44TYfcXjxXfgAMNc52aJbE
izQu8hg/W7+J84QsPHEKhMempruxzmC61A8hXDwd4kqpUDoti1kwHmneWaktXp3tGGQ0FjEKzDTY
28pkznUcUMghPRGX86yrJ2ZDx+LdHrWxDwgykNvKtW5N88UpTdV53c5rUvQMwhEBduLT1aFwDL6W
18Zp2EbuHvDUxq5igfwE2Vq9cndGMCs4c+2OT6lzk4shtoQvPOUBp48niDEsKAQgmF/wKl446kIh
rQrtwVx75pgwJd627+vZt/k1MQ2TW7ji4Zou2zKbk1KGpjz2MNKUdFdUfi3rDb/8m8FQX8zDGD2d
DwC6ED7SDT0euN18TxI07/OplNWM2CFzi1IU6p9Hf07vsuaCOEVn9d+tWDLncdz8QnjvrAZhjikV
pZYMM3u6Kwn4XJSWiT+x2unGoFlRtqMukKspmnBDw3Ei0F9/nlgafHk+oyhfGj/Zq7PkV0GmGppk
29X3jq9NM7E9d8MuATw8AY/8HUd3TQHlz6TH4A0ExE3HYZ1oNTyI7ZqLmi/0m2eSvDFer3qwCsQv
LLeQfJdedvQMYVZNIqLcJPsoW1vKoeCUNe/FACAq16zifEcDgi8W737soa05e5ZMmoi+Ogt3uDpZ
sCbhRswCyRKnnqyPnLAblOeeiGOyAZTy8C+idg1B6kjIZYyVRF84eDjy2fXciKd4uTtrsZf7jH5t
9o7Kf2+nfUfYp9GOd+oJJpFCOj3ln5U8o4wPjY/v4pb8Jjuz6UZf2myPrwC2cBVGKn2/SjQsq4Z3
trdWJZAhg9GCm42mMrXGtoMin6cXxUDSUDJOtxtOahUvjDCTn+CHr7HxX7XNx3G9F7lpBhKhXsJu
tqLFezsPKGipitJhZPjuoxoMm5UsAmvcYsK8mBJNiAMXXhnsmcqXCRl/BMz753Hzl/9gkh6VD2ER
rTP8r+PHiCMpoMmSxAfi9Uffd7ItYq0JMB0GbwGjyrMv+gTjAMmGhiJOKxiVCAGJvDpCQ/jj4TpM
A77Gp1jsmyZlV6+5vKMNY1loXCmm1yvFLex3ehA6SNWMq424O4tq1fS7JbfN1rvA+H973hG3FbJe
B0cCwyaQDRJrFPTj+iuSOHzHmnonUiHFyaWQ/p86R05M+qjo/lPXbDTCnkR3Al8mQwBSVD8DQpFy
SBW8mG0SnGbayF0yxK79WSwWKhEAsps8WDmDhhWY7r3Zg0hz9lyWiSePrWEpgHwkx4CyLuHQS5h4
JImNPwFRNmpEqehR5na6un9C43Ien6f1fno+2VxF8LG0SoeJ1ZyQxj96y9Cc4sKS2pbGvgOcY9wj
AfiqqpKIdLAcrHpN5QgT79PVEkP5/gFNXcgO+A3KtsDbrF5cz3Yvu/8DesNsGkl4WxXgnvywBjM/
sglJGrBpeEANApdh61p2a/AWYj8qkSXrbw3F0N0ULQwg3BR2ZKfPEneMl7Jij6diBvbVq5sQoDr3
8hr5gWC/MYhhnjHf0a8w5AFCNW24oxHNomKNH9Tb+QiumPWPHstcgenROeFNhpAjXhrVk93iDiIb
cVmzDm6oHifHwhBsab6UJSt/t3bVNeufj8jPswZ5de3KSTRBTUUXzBxMgUrPgRhUkneAYUbGu3Cw
SjDpOD5C82vz1Hmqc4g/eLk8F8pCDjz9dxKb+vsCz2xuwgkKG6nk8K0Z9WvpVz8hvCjEtMkt7eWl
rfX/x5LNLT8qApZfos5PsrhnbcAwtra0Gf3tDLVKap49DJnaPd8sHdAmTKDy7mjqTdMiMjK0TQfP
owsPDI8kJAWvKP9aLlwhrV+cooELbYEDc4DslU/QCpYyWlmZXnTWrgSt4TrOkLjgW+Z+fwYextSc
JUrVBtC1gYa3g3WHZ97Zq45kHmPd2WE6zD/86vnmicCw2GwkogoINOqKFBcWsmOeUYcJxYR+TN3M
7Ey3AMSZnftumGGfB/r+dL63nOQ1LnBzx5RJvqsQ0HQeD4X4Tt26f+hpXY6AyGzwx7ZARmCgLH/j
jzIQCZ/Jj32AnRgOSU8ZWCAC11OXTX/x84+gXREUY7AZrEka1r1hHQ1l0bIo2PXdSd/RzKPeaiSj
v1Ix7ZczrnWPcdwzpYSOrkE4le+IREYVvpI6p214Hqzyj6iWYoGRzCn/LaZCdMHJcSIacciBJYAm
sNsoqdeCsjpEP81efsU08i7E7RdkWjb48Fjj9dOi4EkuXWbOtFaW/L/SVbQgVlL6dUGJbHxlEo2I
ilx0d8Hqyq7PW7mD7ElqH54iNP9EDWIM5yc97DonzFe4lOsy/TCn2zlThnagJKnznNsKY5uegTfb
yBTG2ZJWn4apRMhTtishoLjEwpl/7/h2/w5mX08wdIRHxxrUdl58qPRjme4eTwP9sa0z5LqlavvH
bv+Z1J+/Ti1SxekdBEjkCxXUrpRBldgaSWJlPkbmfsDdWER16aw9GD3NurqS1+jc5cuKC+wuQlfB
oNSoZsVcNCvTgQJAHMLo2MZttIS84e27T2Z8mWFueRShJoALToJiYtOI24HjGjfnW4pqrBaFt0p/
nmcE5g3ED1eoqImhiwpJDkRjplp6xo6azT++cqumaf61Xh8WCmgirrAO4ovkR1eJybJPDNhCaAuw
qeMxYS5F48FCHZxfs6fjF22pL1cFFNTNR2YwCCt9j85Iwtmj5lWZbY0K1wYlHEx0FuPj4oKuDec+
m9cYttLzJuAReBPXQ6MOParjegFk16KCk3ildjA/pOrG8GJrN2MNIx1S+K0KQai0KvK1dTaF8f1z
18iI1BhVEuIQkVRht7lFlkful046AnaWh89qIlTKMYFD1pD5uwsFGVjp3tiWzA30rDsI5FfR33vm
plc96mj7axJI+YGzSg87BieXgugFwichtU99Add0O4I9nVU+xqkZBHSKJi6yD1nakGaU3/zY/JZl
il0l1r6s86KjdoHVhhYfCAekKfKax7Y+TU45hD8sruNWo97oQEIXOGGMzwg8T//CLXy85dF+wphB
r95c4l+ueLGpdpie3xQXWVQv6yn2TT3q8oYCzvnoGeSaarGEe2t7I+IkCtQs8UfNngG9UL9nTE0y
mxH+FROi0OWn7niPwYxuKmJu8G7SAJM85oxwiB25bAncq+z6XzQagu3pQbyumR+HErv34OVajQoo
I4VjX4m2FMKIK9AEQkukbNCCqCDLfFsCJCRFGryn594X18S+aaBIIpmlm+0Xv7d+jZ4yf0LL/zP3
55wR3Z7oOW7gfKJtwyYRok7mOM7iiqGuXZ11mo/p4HQl2KqeTVm377l0Ud7O+3nLGpGzGRceSO7W
P34KjRaFsij4NIkNem+mzqPF0a8Xq18/QmarIQTWaiUgrVQ3KsZhaMKpZyyvISLpRVcJx3a6K/9H
kZpygCin7y34k8KM0B6ctqbSskLPNHue9Bb1d7AaBn6Vrhc3t7yL+PbDHlEXDDGDvv2U+HxlZWnh
aem5oBeWfgGmq+jUArhQsd851/SDWfZqckNEyBnY7AqrzTvW0CDPeY/A6Z5i3kQHY8Z+VRTcPgEW
C1AvQiGe6u7fCjpx69PWFZrBlGkXI3z13rDqoEU+w/u83fa/buFnQkx8HEGtrXIsjXMeVw56khLQ
hYny01wwlp6ltOBl6k2mepex7+eQ4jkAJt5/rs2l2WwejZVrMjyP35/pCSGWKEIrv4acFWi5MOt+
1zQ4xTTdIh0Q4/0aT8gM+N0DX6ukmsjgrucaRqtAcqlT+HWVz/KRNB0dyuzCA7YYlHJwKhYqP0c3
ilUzTNF+eA+VSbZPV6KjV4oZLzDy+zhA386sxfnSSCr8MAXDNYlVP6d+5eut92fx120xjnw131M5
vNK1Ukv6h6RsSZEMe/6hNOjAeWFL7ypmKVqBgeesp1GXLlwXuJbHY4f9PcRPyMRVwqkmDlU0q7OI
4hYdSarRsz/FEFW4edd0eIz7F58s2cy9dnzjJtFKvNSYsk+cc2vniQCOI8T9LXOQeSLcmmfq+e1k
kLCVDmYi0vLqp5UJdLOUxtPxHJdPuGTeg8Er2oyHOrP/8mxd/wgayd+mRxGeH1+PyOxQ6AHiBChV
7VeCpVjBfl7hesH6xZk9igE8P4uo63wc87hb4f/Nc1zm1DJI930864G2qaNPUCgD2bz6IaWqNk9r
wNMj64oSoDwFD0DFeNVp4horcoNvU5AKvqbsmRCJpvfIWimDq7SEg8NSSQzY1IFfHUUDjTEu1XZW
zfiF1XtDo/dWfzUJk7xfUWcR+eTBm7gtx5ENqhAFiyjKU9ws27tV7gEd/KUnRsViY0Wkc3dP0Vb9
UFsgMmx1aBRjAWUodB1rvYJhSWX/+W0RARC/mzf8SPHVA4f/kMP+J9HOCYhfx5DC6MC1Bwpqok4C
6aEm3O/W5yU0vSMiFzMQsv+v0iij6kkSYdCcTXBVXDvjYq/YskABDo7sW0yOrkFMLbX3p+6KEFb6
xykCt/NiHM1+zx8+eKZU48/IBLyQJ8fe5YCLH5q4VlTulF2cdbMVA9CtAkgXdpI82aU7oOpwiLuA
loy4CIqn1OLg9hnLwXTgt90VfmnZegA3Cwbb/XdQYKJlAkBPXTEsfjrhET5oqY8FlEC6RbcWacha
Oy+ZrEpbZFv6wMro6IXS2MjB6+f2mw6ASDd4ttUHlj74NPyfdZtoVM3XuRQk3LbysH6EnO9FQOju
UU18RksJd0N5EK8758o5h/vzsPJUVYePKE4F2TCJvI5YAdDKzhHDVMc/4VmAqvvnric3cKfeybba
Jg+XEkc8JIsyCce9INVvR5Ng6h8o8gQndBVDCeZouDpyjgNhSW2/41Jgsc8awfqf1Tnn5TfaZU3y
RUjCaVR9sbhAcEdfBAFgYD26KhhNRuczvtutr+eTjMF31Z3TnVuyid1KTgKP/JlAJI1dLydilKJ2
Id+JFCSje3oNGlQ7suZUr+brMFktibeV8wRfszYUP4xGTnv5PB7KUiy3P2pQmDl/7t+L1/21ETbb
tELX5tbU0M2918ZjPf/VtjJaVImDyAYk8zmtQi1S8VkYQcQsj6qa/JR20b/5jEsRg2Kx5rRlDZye
dgailNrMEjNXUbC0jeW92aHMs8Zsi4J3BUaatTDApKG8CNcJdhHE6I93eIyaarHQbeqE+j8kKknU
ocUKbKk1m7/Kf0afePSi9iJk4bi7urDeS3Wtu2aoPjEYenZTBZbKo0r/ovIJo8NF5JzsBeMtdgg7
XjJZdOTYknH7UhguGyOsLbZuIvhSwTOFpYSOQURKGxrtgwgbxtj3d9OYIR1bbJD9+3u+kHDYB14W
n3+yhv1LjFeTZLeRINI6gRT/VRnFrefL8dPZ7yEsi/cjejSwYfYcm7p0DVtY6b3y7WFRfdF+L5In
kpgKbLEYhW1kP9pb2yIxZiWNwRU98d1ojiAsVfLiv8tJbXv68Q+GJ5PeKcgvm77kIKWaYANuhQr1
D3L6UPLWnTtCrGoq3axVsQmx0JtnWSBuGADRLV7xM7JjTNTgLgMleAHhih3TxICQygIcf3RzIoCu
Kk0pI4VnDyiQkkh1os7ybZL8HwivqMBUdsCpRbRGX0wO5csrxQePHV35f58dLbKZ9jFIFKxiqm/t
8pEa+PO+2gszmJr3GG3sHRCBpKVptKSWm0ng5Y1oZJa34jd2zW3i0CBmP78qHG6HYIHUVH3Yd7zp
tjNXoZiQ/bodw+Y+I5L4oy8N0ohfOVt9mz6aRVoO2nvK/Ivkgs8+AozLM1vmbRGs24zwFiYZCz0B
Lg6dWV+nmYLdGB5vx8jdrQs0RZP4Gdj4VIGtWnupYJolIh5VlYi85VqoFXJQhmVKdrUkWchHDHNA
rF1Zc6TBr9g5hSDeiEkO3B9KL5r9V3drM6Cfi4IiVA1HqnQXCIPSx7kLfKD8aLGpP7BIbh6RB7N0
+BHxXZb85ePll9fc5gmwgBWgMb8hQGxNradOF7GryCZ1dseUsgR6nqG6uS5UNZpa8a2ZsZsvIrrQ
YOIbrUlREGXjUyrqcYbGM+60Lk7YSYFgoqTsADF7sdK0jPw5I3+IYvfmJZdvpjV8Ag3PU4OgolXv
WwORdKBXpgKvwIac1hatTHw4cLFM8HPAW1GnxGr13Kiwa9YK0nyXZqXCXGjVdh0tCC/7Dx9/pHNB
gG3wPXY91OmSRVANE3wTxMYuX+O2ZS9g9qVkF6lQ3qLkbd8pPEUATSFpD10jp/ADXfHhcoDSFzqp
xHf370Tk5ZUyO0xsfUxJeK7fHB+xHKn7huFFu1Dl4vcZ94DiCeV9A4zxzTScygz+6E4TcdPu22KG
PCD2jXlgI8XTdcNwhgEiKR+0UCSVYFG5/SL0QQMwc61W/gAZxG6yiHPEZaYMFB2HGseVhlkcW+N+
p/aYUsf3+227t9+SXtH/RKInxb3RZus2YDTX9spcdhZvAF6ZGHF9yEaiaKXhu1BCDfRRkFK7UZbh
DdSH488fX6qd0WX7YySjc4tvXAK2ZTrP9PK9NTjIhOOw+ij1GbNqJf3VpZJJqxRVN5VyEivEcKnu
6uoHSyPsMnEZv1nxDc1V5UtZDtVQt0wHt3g8/xdqSLlR9gRBKupW7bjRupZFzhwwTyKbj+kVxf1I
/ZADHsTpz4btxzty+wad0R3Nrbb4oz5lVANm+/r2Jtu+F5nhJdPoQi9ge1cKmUinvzH7EV1MNf7z
q0T7E5W+lpPjYEczib/vC3turMxOnU2rtiqpmmIKRCtAUHf0zJiVqKmU2x0KebZFrbfhO/bl/Hzu
KCpxILFOgHssk34XteRSqDiNP6y4R9Bz5bHn/q/Yu5RnZdYAouA50cIldIZmPwTFUdGk8wCFuaRs
VFahFktYRQZr04S7I77DKR9xkvdrcTc3aXN6teST3WJPrSm27kf4l8CVvHrFYlFcPqfH4X5TSTC2
ijW6ehsXRXG8wT6V1NziL1XdY6NEVRB1qk/FmZDD+V79veMUTX9EnjMrSv5SkNUlQ3yCX/hd8net
Rs2FTaoKsbWkZMNz1YzFf0+88wpSL/TkVXTrxD68KNwY3TnT3KZBeWTRqWkGKtLAtnW3V0lz64qU
h2BDbwgufbczCEVcieGsQmhK1GnGZP6mo2Wnu6peaGvGYWVQqSNOAk9vJw+HCZcWyaWTt7GYPJv6
rlu2yBLUKGV/c2nLPmq2HqDfbIx08QMfvmdYhC+CeKn+YAnzt2vyLQBXfDGa5MW4cwiaJUg6NZmc
KK4H7AgT9plNOdC/2XgzvqCwawRlKpO29nG8PMDrtebXyhQnHwANdRSQ7z/pPgCpPbCF8N4IqZXU
ssESf+Lv9fYbOI39vwdVMJsrd3n178GlE4q3TEhnJYClpiNZcn7+hEOK8hOB653B/glfWIWQvatX
TK557SRB/ie7apnkju94QUiYy6v+E4x8bagkQLjAqqJQm2DHOOJpcEFrSkN5h26rWSUBYNGeHqnS
+jnTOuF1R1Hces5zC1FVGF/lZlw6vpDGxnTtmowmQToosIJrMdjx6q5NfisStORlm5d9WPfI1cK3
b9X1RweONsRn5jCjfqUn1RgqpiQwoDHQQ6HALkv73QkMRbXbBRfnhBvpQwAU0FhkLx2ftI0VKALv
XYXPcMR4UN7gt8mbWqFERKOLbfKwMOUYRbRSyCxiv5OGUSH78QiPBxE4DcvjI+IggRmY86d2S266
NSfmmltnvYM3xq3iLHGP0wNraVvPvH4UONmfsHcQ5Xer4mhx9GEejfs7tpP46aLNb+gdWyMGy2ec
oOptsXwdLc+aFweT5xVuJeE8PTUfwKhl1g6DpwVp+kksgelCUsUMlVanMhox8ogOC9ySYMxcGjsP
RcsjZWUit2bCEQoPrmZ8w8Tw44xrDVUgeajp6tny48HfekXvzb7KAju0Oh+sNAzN+F6VBnKWWRPN
WeBd4l/L/KYyCVryvfYjcvEQlVfquyXUF8kbSgzAnwfmhq467ZEV4G+KOE2UZxBms2J+1r67C52z
kgE2LfgsN/QlHSnA+ENFcAsSMIdYLtQhiyiobKfm1t2tIqgQJXhBsdNfqYKyVLrKPgQe3pJDwf5i
KHuUjBGEztgODzKGrIdGaOJkVCM/hfYRpNRdnAwALfhFehRT4L70MiodfNihKG+FuNIQIHKKYyS7
PxB2jQpT8Pjvip+QiV5gfcD+UKltWOAJ3yD2/inFqHUHXY5FKkntHm6mvUBOEwUEvX8eziWa/i4n
lSnBQj/CFF4Atv2TaiS9Wy/dVOYvxPCFyjAVE6q9ybuMxZTTRXIhcyDA/nhugulrB+sRSsvJB70I
IXrB/ukeDnLCU5H0YVFudfCtfR9M7cMc/zEU2heabag29itYsIUsKgIWCTVNKVEsCu4pcA8GMQhv
f7dXqEKHINXcpvsvsE0ExvSlJmjlUDO7jHvT9v2HeSI48n6hQXEp1zvUR7w1mZRu/vybbdhn8Lom
kkEWVCZbeVdsnBGHnZRJuy+qq9zWJTLprOdvbgHKfQKKpoqLx9BZ68UyUwDtFIoqwn6f/N4kIrZr
zFrszkGU0qz0CcrSijpU3tjSBaydjXm42zbhcadt/sUSSjLYFEhwwpKIJO2LR4XmifG0/DM5n+Av
UbqpnNQXtrBf2BW85+uVV8zt+1/M9X928DDCskyEn/VxIhZesn0alR0tLRO41cxhuQK4Op7p9A9c
rBCRV6RA3xZfXP6Yp3BZ5YffZAZWSNf39NlbQH7owxTxrt+SKqsdZCiRzJLMtCGm0k4oBp+tbF/c
Fos1lqMqm3/GMeXFVtH+WoLqA3pNArG/epMzm5o0WEVYfUJrMnejdQHBfbF7Jeqr+sqa70xmOExV
VDrWlXugXGuBc1WXF3J7x+V/B8HvI+THUmVLTTWPx+Hdh5lDHQePkFYQJWwbkTs6ILok1JjVqITD
h2iprsenoAvMQQEpYsRX5vyfePbXcnlcHJiSqmgDubg9liE1T125Hpq8FVAPoMzPnxSu+N3hjEag
DGnoOcYv2PixBjh6L0CxLsqZTSdI3fYqYde1Q9AoXUGdN4RgqnPLU8EniCHXmszYfaQ7K9dee8WX
84vGfbeQsd+7Fr2R+r16ZCiJqUGJRzS9Elnnibf8z60XonqjlKezgJBhO0i3HUcr7EJrbluNnlXS
18corjElBF3Pad8ZA91MPZKgzbVvRrZLnp5WZUu7hH3t+bHAf0mJTfUsrRHWHSg2RaRgIUaGhi3w
XKd2oJWUrEGLbs4Jnp6Q2bQaydvgsMnhRMuvR4RmsLWZ0KNx/YtZOQs/tbba2f+bEg37ABuaJt2M
JJtYzwsdZN1u4/2jLC3U2OLI/VGBeAhGX4WZXidYKVijr5TD28GNrsQyIdF73DQjTTyBwb5TU89Z
JrIju+f60/IlGExCX9Da/4MgoyjNhPvLPM7IXy6Fgi3NNXjlkqBKSl4dI7jOadQRMi82wV3u3z5O
0Cj+sNUTCkjWHrSveJ6asrMxuyG44du++EFXUjEObP0zk5WTqX38btj9BKm2b63LO8MuORI7uTA2
jOcrh+VCQmJwCBp+XFRJZDuCOUxRSRpJONRMMQif3jrOZyqIkGwolzB5cJnegKeyStzpUij3VYwx
qjbf2GxYpkei/GPZOTTkxRdnQngGEmwdApB3iYKLpVneXA3s/heOVI9aylDED8iN55QpQXNDT5gZ
3UXNyQ4StrM2bodU6WQ/uSAz0BFIl7ZE434eU6QiPUCmRO1V05uG0OYW3ly/cL6M6lqOSw2cyFZH
qzqc50c77fSAuPXYg3kxl7Za7sQHJO+Lxx+twJLrXalnOjMDWMbYqJXVtA4tkl4AVHz7EEnT2zuN
1nHZywsoRUEw+aRVYbCHqdVM7qkGLcvmuKAyeJzXjNE65e2L/2d39fapSYOuudUQXSm5LzVdBFyi
GL2qJDkSRtMJMArp4l/S2+yqqbjdYNcuoRIRiI7mDT201uriuPah+8wbn926ty/OOvSEMGThWjUW
PGlqtgxSQbXNNlr4O5AwKiUFYpP3xAn78WO8jqlLEkcj6ak4qL0mxhMbHCHCerNFcfd3tA/ReDXQ
MoZ3tLcVlJLdDBi0OQebfd8/DyEHVaLhtxIHI/5uejV7Zuw+eDcDtqIzscLP9NgOG8txNaDmKnKY
yWUqqrtLKf2s6SLhiK/qw2WEZYu2gAOYhJx7LxUSerKk3dUVjKI5AZPgH33qZPzgIwk964jWN0i4
aJZ02uZLjY0s1GW8dUVzPk+9l1U7vkXGodemvvj+aMVH2/j59XhrtNb973w0xavVzJ4VVSf5NO39
YjyHVrOb8FSZyGySMCGLWjYEIR/ugj1RTu4SSotZY8NiGkz5IbWOq5fBkpU0e+l2+DEQvnHLbEir
fenpU60OtB6OTlUVKvls54B9jqPq0BrxDvQZG1ydD//hx0GrqZjEb2lXsUdRgKkPCXinOhqrgBqg
APUd/C6A5uE1jEBbpdv+Q6HF0GJOlrOrL7P13reFlu/CRozWSEhs5jcB2BKHajnjDTuZ+g9X+nR8
YWc5+fZMk6KAmdJrd2u5taYOribcIS1qYdehL972tsISyJOrTDM6SxniIsq2bS2b8LQwLhHgXAOY
CFpl+0WX7j2M1FmJ1WK+vBJ+Zslgb1lyx5L4WqT0np7Q8Q1khqq8sWYUVG5ggGCZmkhCZTnAMtnG
O19PS2nKwdOonuysNzfY5eMOEsBB0DoH+gWBqBkUwin1ve3R/Jxa+IWHzTNq6wSDT5c4r6qyJ/nt
CS/bM/pEP1+0i1Rc2fxb4EDTZnKeKEc5TXOc9fQKnnNt5Deg4TLLxWCcp83aUcKMzwjzHzPp24e4
66RKw0nBNNP99CvN65wUT4H7bMIUwTXzuSbVp1mkf+zzsNYHRIAY0xAdoQrkssDFnGgOmXij0LBe
3NfRAux6qgkfoZFAaz0KpCC7PKLECG8pVr2iJ/+qWndepyCNvNs9MoFEKm+2uWFR4Mxzp4Z8DV+z
DGsaptDk/TuYyw0BDPIOzgs+XayybYbDjJAKW2AJJZdUC0fciNpn2T11ZkFgSrReOuqcCUR3cFYt
585+DicOizoF1yssxgOolRcJxntGDE0e7UqRQ/ZIyE95SGtf2XJfTIZ2Ijjvah1djFZyQeN0Oh9y
Ok/aOwVcAc2pTiB9AePpzfvRS5dKxX+Muku2CL3R1KtA5FrCxk5hbZ2aUEH6ZwBFO4ffynkmyGbl
4nEZF+J8/Tzklsy4AF1QaJtis0o3bTjLXG/3LUMpU0XB271oIjH96acKGjX0tPpWZHH8hIzPT0y9
A3LdG5WQsqceMSMWAuaZIO7Dwuqzhub93eTFxvcgMbIv0WqWMu2JubcozRILnA2b0o2cMeLzqT0C
+FT+qaYUfMP0ciaqNsNcOWsGdafUUgFVawVbyxL2ZyCgHu86xbFhpSW2Q388VlTB4oXKB3fX0pLF
a0S8JIHHseZWMuFxMbbka0Nc4hZkKZI0TqTEz2lhakl3uJdxWyOGLT/02GcKSwyMFlmC83DEW1Bf
4VTs0j7frCexgX1FvynCD96D1ggO2JeoqaUV3WdqODvY4gn/303kbUObm8YOBJs+JuTb0FVjaWnI
2FA5VB3uMFr0hMm21F0yuRC90yTUXONzcprHaA01WXBsDmkbLd/P7j7ObacA7/bep0ivZUofcHFU
lDq70sLWRbGEOuN4u60soZWBxjX5SJN4/m+PVojOFfTPOQjICr0b2/mcaDaVG1bWgBpZq4bIop/A
6tCX4MT6NJ82jSs8TypRfcJCGQxcc2iaqO3+68DoeKSHZeFNpmmoKJONztrByCmEvHR7WnNhh+RN
Q6o0KBSMHIdNaYcoY1qZOssB+L6ioRJTSWvrJjQ4jGig8RD5s7zL8Bb/M/ZoUzV3/5+hKC8iCcHB
hwECvpMkXJ97+g+X5uQTQEMv/kLKIPDR+ge7hMbJ2GiwtwGJFGdq2vBCPe8eRxK9a61E/pg1roX7
RU2SH6G9kTVZOuWEMuAsn7Tic8zU0l9iWmqpT/uorjIxW4wQOwnfigSc8rxwQeXaLzRavk6Ee6RG
1W9vHC7rKo9fkBkHqOmMzrOeNR5PqTLy12SeGYv8TvURDsTi0KJu0brX05gNCT1Pd49Yf5JIy9ux
38IV4cHKdvQvrk3Xi1mrAblmZLEIWyyCDG+++3OeTe64bPxDSavK8/5Kl9PwjMtMY1YKlYJAaw4O
5uVh6K68sTC9VePckq/N7tP+vRnkT5aFk9OYe9z6+KFPYuX4UeIiRkILaOkwtdBW8o4VrWp2Z08v
sqoRMS/N7ZWUWCB7yJznHQx8tf37RO6t7CwdRo4srJRhez7hxoY8lUw/uZCyFDPNVB81bRR3TVCG
Vi0Zn3vqNl9iTNSp3aS9pK9CPy/2l5JOxCsa7fPoVN1SO6uc9yp3z84S+ecaCxfv1nlbrrEpzhnc
yj+iy5wb+azLnEOhECV7sKbTfY/n+GK9tTr1A8XGINZ6Z8zrRwd4JsiwtjPP/tywYX08YXz+tKFU
Jj33/WYlcKcw3yGzGpKlnENevz3vvQamnS5TE4ueO55zzPpjTJUtYlsjxJ/+zK6ZjTfA8qw3QB01
UCg9dECIpo4hoxwipGNVE5E9IJblrM0PhBcvXrYeaT5suXuvo/92lUTNNKwakfM8IZmAQAqNKf/o
vLJumWKNWVI76YRjqSCSIdYPxqRd5OPK1XzjPNzl44bDZfWqCNDD6m7q6bO/ugv2J/LmRlmIkt9g
/8xdSQRRfjSufNjreP1+IwAylnMNqNgd/j191DxsGi7g8zp0h2W7eVZjXgkyRkEXoFe0NA8pEKeE
uFzjijgmBVy165e6w6uNS0HTasmPkT9sd/10i684BKAG0exUdCRHSJXBTWP1wTkvq764fwVrONrh
rCJaV4MT2yFcC6WEx9iNskDfPQg55YZ54b7RAfKHxmW5fKpTxuQozuhXhrM0MpsDgJef90w6yKtS
82ILDMyWoWHdVwuGzU3czfH70t6KhcUfgmf1cuvxeTB4i1cX4ZkitzVZImpv5Cxs6HKfBCKikO3c
Fr7/852oVmmt/6b2hn8s9GWQIalgQNAzQn5/+2BjbvvIBvuddBOzhOJxGJV63EFpddYk1OZzzOrr
KxZPF0PcTl0tGnE1TzuIet4N8UdPnkgzLjvGDIrIVbC90aUzPX/yYe10mSHWUYHPfhapG4x+pXND
5IYIjziGibPcEEK+gGDbqrtadRc2zHdYE6EyEeEQ4KZehen9bCW4sED8n9F+UqwKIK7hqc9Ok7lp
rrlWrkKs8emE4SPyMY4QN1LcWTsz4Sw4XbqUr3a0kTtVmz4xPqXNo7EvqURnhQUUHxLLQuptQy7m
lnfuZO56Yh5OeId+i9LRp/p3Th/cS1OqXBU+1UM13D99CynADrsy/wAw2DrkrvHtSv3GMF2x2GuI
YR8DCi91Lfqb16fLwKECLlUV1vHHgPEV2RMuxLCSeyQZKp7GM7Hsfmip5EMu8Mq0fIGv1V+zDlbC
/RZtlEZ2jV/JJG5hd2/KJ8E6mpOPJaUszeaLWRZTNIqK61/KqbO5IC3DBtXRu4WthdSnz5A/3w0T
JvxFd93fSPH6Dmu5gpOewyI775KYKB9lqTHhzquoFO0bIGKszBQobb9eYgQAwOygawD9Ey+LMIgc
Tb2vJBgl8z0fOWG2jpU3amMoEQr+Tor76XKeNXw0aQrbm4wBty1PITp1fKCTRdcQDW6B7jsUGjF/
yqZa6nVGahJEatBM3+YIEGCNvzvRZyckQvb0oxRjlFkutKtuh3vkdWeg4a5k2h7Nvo77WIUJnZDy
dQnFalyWRpjfb426xQ9frBpL2wdkaLZCQkziHVgxu1Giut6MJ9+Zce6Y4HJQQPZwgvT18taDEOKe
wdvrsuLMJd/XPIec0pwrUNjZeaZ6vOh0t6aG5V1/erZyjQrzDqDti6RB9RfRw8Gz6B6GlKVEsnG4
LjNiaVcIh+AwN7eyXzYW/YUT6S4J2YD7nlMZffhCiMNt5Z4J/NK6868cpfswxeLOy79BSPXniQ64
tL1QgUYHUNODwxCrlsNsWLdoPGIiXfXgpj57KuWIx8P7xoe5MSgPnl8iKNNbXAy4QTUKHbxlkoyQ
bT3y9vRORIq8rla6nXAOmm223Y2Srd/+Kl3s4D141W14odhGDV/AjZxKezdIdeq3ytXGUxgAe5gg
Luxwry692kkNsTYNlY3Rn/z1+eASadnBNEVWqJcE3oMNiPZsp75WmhH2fJbRAszMXv2MYIkJu1rm
TWhK07GFq7vIlG/Eiel+lCEQKXjKsSHV6PuW+746VoBe36uiElnLMIs0D27At2a+l5enfO4viN5b
mbhRqWgZJdarxlxnND4ayIxn27jR7SZWvkFDo1wUwaQaOHcoQtnl9H625O7POmDzCtem/j2iP0Ed
HwIT12ojjtKfhZEiaNo3/3DXUCmer326dMUdaxAnJFsYWTxOHq0oNz4bEofXqj5ZgTs0K2sDSaW+
9K1D5p5yoZYaohm014ebmXrPtiDbnNVr8LLAuOPUQ4ez5Oyn4Jc8HXkOFlKGwHGZdddtkhsEautN
s0+8zmyRCQYLuLyfjZtcE1DW+ZgK0omNYB2+lHS4XPMVdlhtrxiFM5mfrgBrcM0UZlZceoak55q9
hk9Y2HJY8tzQd2pgwsoQjbRTs0bn/YHFDCRHVRl9rnyfJjEdDjPtSddRDKnA4lQEuNUSl2AKdLZh
gVLv6Pbm/Gs60a776ResEMmQgFdqoQbP2/BxW/PgP2VryovA2n726hZ3iXebP40pFmp4Wifbv+uu
3L0Iy8q6NRqAoo5ky8T5fS/WWHj95OL6XlOpdAw+fsff7sBsYERw5uSQbOK3uleMNjzoxJ2sBqg0
nuL9ee6i9L4D0DdhnB7uDwk23uCm8GPfldc4qnSZQAJKs4vB0UAD0bp+8JyIuXNj7SHVi0W2Nlef
fd37tz3q/R6mJyinqDf0D1533Ix9251NjdFukNpt0H9pfQAlGj09ePW/SxISZiraB/QaEGTOih4+
yx8buFPpmoo/bVuR4TlFka5XL1SWgWg39m7WvDeuM7w6qfjVWWBO7e2r9mb3kafCvUkkikSJHVNR
vJMQKQWQ/lR4d2rYqNO7e/cg9Xs3d9x1D0XlcrH6UYiEmaPFE7bvYAzBQ/tthYZhDB9n3Ztk9dR2
S2CAyJmHIWZzpdqyPa38GrMS/311Bh2TI81XS7MpBEsTjS5De2wPWMv0YU3rEhIXpkwgwhWHXG+e
6DdHPkvjWENs+f+ZJYfD9H1JSHCy0Kh/xY6ZFn0MC+Idj6z85hQEq2CNRrf6bGI28UVSsUFt1V6z
TlMEcgZYbkSpRNUou2n+QR8/Eg+x45/V350pFag0vjjYVlUiu1axW4/gjEF9zhXhByLtl5GPZvNy
VBMfRzfGcNO72hXl0gxIBwQjdL/XjfbMF5NMFrC8xum40Y/BiwKEpI+GpakvTtDvJapkT0kIrLUO
tJ3JUUMKsq4XFFnAy7T1tVs7AgEDtEtuteEyrgGPdRdYbcC08S+TLIsSj7ovKM3E8tTPrSMj6xfA
HsKddq/ijeE/O7D443x+06U1IFRXnUJxo1z3vqKLxirRcKJNA4Jw1Ks/86WVDGxXRfYGFKY8PjY+
9LKTtrBo26I29+C8bvOZI+VlDClSxgTYnYAaa34MCImyCC8udCAwP+II1ej+C31Gh7NCYa1F4pZ5
rJC9UIIwGQpVAAkQFVFgGtv6U2zrodrAWN5w+Dke2/DGhHBKBZRqDt1NSD/5XNb/StJsX77/bEye
sWOEOqqnEbmVXHWXIYp0UGnS1MtxXlkZddo5m+FypeZAM0uvJpuzOUmrJOX2wYekFjjkL2f6nU5R
roiM97b2g06iE0KvvbFdL0AHS8SEjHrgw/6Ef6MrTvPnUG1MzQQ/RQMnkWNmOBJLKl1339tNhcxA
Zdz53d+TPasBG9K9eFBxvPm3KKgk0IQNGLRMP75XtvcX+H1IybXPyWZqngu4D3+DeV4Vk64WMrbH
5EG+EZVQmg3CBTxmdM4ovA9SO/TXvdT3GEmQun8tSJGk9aySqh7ylVRn8A3kdYHPYwMJarKc26s+
6JkjgsuWVWM15GW8nRlJVLVKzFD4qVSQOaFdzCfs8QvgvdjiXPVQcPprCnUUgw5RvSJqFgpvz1Hw
5HDt4xhkBftADk9d++raCiNk/oIEqUAxR+7qcgsDxOYcYCDTp+2wCSDPj0593sezhitC2Lagt4kb
vLBkECEiU7VmzddUmMaP8ZX8ht3S02EduNiFUZJ1oW0tudLVhWlI8OMo4W79Z59/XZIgFD75eE2L
ZabZjQI0ZQLOnH+6Qmw/RmXMqcGmghI7xEHpRLQU8IIfu4OZQyqUlj2RzetOUoCKqpW0XrBzgRs+
d+2+3tuMrGH4fXo9PKoSiNBGv1XG5otvQYox61pHzaLEqVPX3mY/i/J7fB26/URdgzYxVZFkeRNX
d9ZMaTSFh+5cugeUY0gpta1gp4cjDtb80UrSJKBImYGw9KgmtCI7jGhKcuwEnxL3642GJNw3XJiJ
cT+EuvpZU+fxJ2pJG/r+ih5b5SuGNO2qFevQ0FQAGj3aoe4MV19XpDwTCL/HVEkm4zkqG8JJgN7K
CzwtsEc8XBImAY8ryUIz+P6JO+GarFeFwuuFtFmafw73Bg058FEsAYVzTw5tLIv8fuU/WN4avFyr
NdoNRywCbFWKFFhKp429MngnCcJuv+LthzsbfebG1BYkkgxHjO/hZrQ4n5i0DQPmFDFVeWsNXymB
Gh0QscA94z0NwHlpJ4CMsx1NGemsaT0ORpWty58iTjSaeqUfj2W3dxZYuddcFfekQdMUPAHfKY33
DkVX0klgO1hKjqDlteWYbMTim/em/Vqmc1y5zfysTjdd0HSDHZ/61Xvb8q7YRwJ1VH4pHbnGLl+g
BQ8w+KeSrBoatTaxQI/f9O+hwnIvcdHXOdsu1nqeTCVE4FeQmuW23SKEbSJKNGLOzn+vvwOdwQjl
QbJxjiRzHT0Gkv1/sOSK8JZS3kxPCMo091dOvxsgx8gp0x94WcIZDxLVXz5FiWu9c4jVOXeFxHK3
3bxhGikK6nsx7iLSkttOF7ecNycRdLX1Ct2b5sLILl4RAqTOkTO7FxYZ+ZuKX3FDPRuYVp4OkOdy
37DGLZL2uQ3zNISoYGm9fAhFUSEkV6pORAWE+/087mYMqIvI4IAPoWstd+n2rdYaAsEwFnSnWzay
5eQqALBdWP6JF50Z+w7T1YzQmedO6MVuk+TZHNgi5Ia7KnH3DPDX/ocvPMKvAOovRe4VnUy1IqHm
+hiWdu4clo47UJFgacHVlAa/C8qTau2GHAPAI7mJWl0AS3B571zAqLkBCtsRbSQ+BLIyOsAVZDDC
8jS9Fx/LFB8qzUAfJjBT9ijS4CkxbcyriYyUhrOzmVsuStWeKYopwJ2Mvmi82tZib7D78UsNdGaa
B5+qdoBaTo9twc6MFQOpWBl3feR95COlfqP/9J1N1FxyHJ8Dal7eclpb/D6T5/lWw0TaLNes2bL8
CQ0KeUtrBX/+rNAk4lX1I2VlGPrcE8eE5niyBh5d6KWJoL//ryBwerYOwxawZJJa5wHPIzoqjYWI
D7aiBDYoi281Z96pIlDa3u59/UryQ653RYVvaPF7ttn+ava1q767+kQ9MvjSiGvLvzoV4A5FuPLQ
kru3jhq2M+JAMJOFtudVqyqaxEdlpTq2m+H7BtAkNfZ4/M6eL4Jz1FZmfwUNlwiU3JwBzJ2Oi/D1
0EtdkxTYBF5j3jAP1cyEl/M/T4VTx5zj1aeg9nop/ZcM+62lBDY86C181DSDbW9oxAPwBYRS6/Mx
Fgva5juAs8WJ2//0yss+b8m6eApZkxBwnou/NCKxPHb5X3oUPqHB39G/PWDsVTczTit63il4Wu9A
FOj9p43eofmaTAzHpXsGrA00tgS1Ma/+Dg7vpB893moVyI8uZfgRnl86wM7ZArQyG8rCBA9cI9QF
4iQ/xe+wv7QmCepXxKUOKPYCVVhv+josCoJPZG8oe843FWrLd9ARGCAGMDbUXEsIGLW1xLyZS/Bm
0U2O3PbzNQVc5hUl6znWy2hM7+XevV6qwWazHn/jCOo6Uy3NKQkqO7B+g72toABcxdvrQW5jlp6l
hSUZjowdGVxYt6DeVCfe2X1bLX7KKbsE8GqOy32AvtdXoIZDMhEmah65C4Z0/t6RqZCq5dY9RUEA
37BuMSVQ+bKEgrM7ebtSGng1+acrzNWnYJH7MkBv2kmw7OW2BCpNntTI07lB7aHk79s1dTwmGDTk
eJsPl9+xBJc4Ox/EgJ+x9vwBGdX1P37K/ofCIc1FSH066ZGImDSrUWqw1OyX8OUaxcijNEUPgerx
i2QPHuYn5KiqbVTnaC9alNFA1pT1pyMlwDdzsTy84hhUlxp1SXcHs4OtTHCxf7BV0/NRUdSMKdVv
ZJh/6gX09HFLQZgA0k7EPwuisz5djMPq5g8BozgJh4t/gs1bRA3+c+y99P9i2KQVj1gFqfFWBbJK
g3iiW8ysxo2hZ+b9sEf7q/l0PQXFWjW92I26Z4JMWoiz02avDceCC0mii6D62Jb4ipmY5Ndvgn4N
HLuVRyyJ7oC/WWkBoCw5IDcPiXQes6rs5p0utv1F8xSy5BrL6yFYLzBMMToPdU7Fn86Zfg3RDGD9
ssYwBp2CZUSXDilp/yTzCPIWn06FRpn/qipzhnECqOFF53Tr+Be/AjT6bgg+rBccc2OpDT0bt8nd
q41lSf3LHBPmWsLi5myqNurCtehGcVt5HmlVyXgmhypJ3nSGfTZ1dIlcIsdJMaAsIXs1Y/YdjXeE
g/AwIq3323g0GEsvzfozJhcPM8ANrpPVPSvSGGghLFf9SlnPvi+S1iu/p4xArXVGhO/bcx+dFE+h
blX2ToQRbiaHdaPU5hE9rOvyH1AqIGjv8AiV7DcY1VdhPfdmIIkKk942sGsqke8b6m+eXksW7twi
cbxHpZUCVFWDEvNAG7CQDx3D2aqxE0nOpSQz5CptufszyybKv5RwSuIaw/LCx4X8g7YsOhMXMoux
AbKNykx9gZX9CYDi3FNoARLPrkyUPe4aqgSwWMb+cNPXfdsJa3+vkyDkw9j+yMLCOAh165dh4Rtf
cvdik1RPFGdAPlqVHsGXZUxQn/Ji+44yYMa5jXhwkS4S9x155dWOMnCENeoK+bFLC3wwUccNgOa2
OPi8fuGrFloHg82WZV5iWGufW1VdfacOjyqXspIROIvpEMdKi6lRAXCHT1lJtMoYBKJLbVH04+16
LgJJ783xAoW0lCsSa3V94laRf3Og5V+dSuFc8JW4e4p7qFe4Oj8i1P9QeyZ+4QMt5xHDtgS2p90v
ykKc8aE9spxqMCqjQuJOvkOz/tj4KuI80Ot8igKK8QgW22JcusZxleePsCO7+ce3bcfwExxRdmav
xwVNr0R8QlqDs7JMwe+u3bRooM7Et+nBCcZQ4oTyvDwpBY2YS5Kkz5MlXZBSnUN1GgRa4peoH29m
QE9kkEMIZwFGj+e00948p491CIPSDBPeazXDQtnyiP3p1+x4FQNXHvT+yfTBwGoJfUAWfyNFNIOv
cUje3/sMdbF1DduqYM6upO4nci0O4ejZfFqnbP41bt7v9JN7N/wRlvGWWuNOkq56LKcB8IlshaqT
aWZAau+oavuEMbocu1k50ZEAV4YoA1uJL0duqjtqt1jMMEwBWSIu63C35BvB7Yg7I2Jp53I4rf+d
Jwe7UGvz6oX+UfvutbrvmX0bDu9ItToAa6cByvjkwadQPqE+xjq8ImQgdwIavQWjV5jUxayouJeR
8SgAw6hI7Y1oijvRMW17sOj5V+8uVsU1+heSpbl8bJacufB73xf3fE4g9kZ28JfecDhlCQT8dB9J
VA7ERCTWJu0a13d91HiiJUs/JRSStCHlw/PTPgLqtHXJwPmd05km9owLunO1I4BfiCriIZbHG9kZ
f+nm3G9pmOfS3flADxnp79Pt6TkGuxHCRgSC36gKUERFT4pj9rZqX123jqh6ESOhv7ysxaHewSIb
h5I0mA52SGdvzZ5gj7O4BH2q588Hc1WMbLJYhcDdzwPYJhks5nhl7jjLWjV1ebEGIF54EBWtcXez
gYGqtG2hMWbRLj7olggD0gWBFifU+ApYDfaoo/gsrz24XEyW4/emd6jAUQG5G07ecmWy/Lb85wJl
1hMicdYFT7X3AmeyNjXPUNact+7Xzk7X8Dq8u0xuz+V9vNf1pE5WqWDKDbf042N+6QiD6UhGudPE
qzzUIpxX/2Uivzopxee+9agAj5inOBWfgo+Yb8bt49rijHPaNJCAayYCSxugAJa+DXPR80+faFf2
KKBWtmZ1NGx70/s5BpmNx7C1PY/+tVdz8szNv1eex3GnPOF6wTocvT7o9Ex0tvwB6/C/796I0LaR
H+oAns8IhMFpVt3obzAT6Z7K2/ZCcrtSpXUMSQVdSZ17dEEvDWQ33B5DuADBHhbOpAUUKo1uBGwn
CG2LnJmqiqAVcTZSwR7VvBn4kk5jXmUDYomIZ5Xwo4DXDJ54XznhSzwTAFijyX831JjBj6R8ls/3
Y3In/1PeH7gAbHDLkJ5r2UATGZMDhTW1MKvRq/PPaPOgfOctN02w6RpUoeCJETDf9ZXmo6nZbOC4
pISJ4anmU7T42tc3OGlVQL0LwCxsW0VpZpKjuq67tUzaU4qH99E40ODTAfkvE+k3ODX1v1I6iVvr
DvvzL+gMaJJdaKJsgJlw3aDPX3QElnOHfk8drpW/E4KdmIRWLy/ARJSaFoCTQtJVouWegW3/tECD
i8GdUDFvnMcFiSHh+FDwUraMXbvpSbklbHUQB325RiTKWLlihhlZPHB+jgnL427ECzLiC2B5zSNk
UuLEz6spGUnha44w+TZw2A1stwgX8iOH4zL4gKW6lur30pCdDhwQInqcx0htGyvZYBcdEXrbJUyl
sayK6u7BcCiGHfyacLINYz+Ju8mUKNXynD/t5d3q1vfidhprMWEag7ubx8ltmSSzDwAcgUfeIx8D
cO/pS4YkL5l820uFS+Q0DKh2v8nbyymAea39/sREhiYFw1EwkGlgAT0VeUU9AvQ8/0gWUb05FZ4Z
ekursXuP+Pra1FUK02G17KO6UroOTIeUNVQHYo53QsbMLg1naiwUZA50XroDU8lnkhnYHbsiDD3W
6mPqj45vCqqb4CMPD7Ewx8GsZRXgdrhgxj3HU4zb6uH1KpUeaqxQSrUSrkAvFtNHuEXJgKaI4BnV
YNR2xDPhrNpHlCJgXcYEUogFTbQDux1qenlZIVbPCrEAJaunaTVLjCA3VN8O+uczZUazMmR3hmzS
TFZAyY1oO0l2KB1nUTDG/wx9yqF6g1fNPOm0JCgCtpbqorIiS6W99Oq8B/FIb9NprcNFZQgwk3YT
2BYPeM3ilq4hYs6Ks4rktKwdtIMmuJnMFd9ruKQaSUDQ9tRgeW7GIks5wDXd76jE9Sg5U96XNG9a
YkKCTJ4haxnZaqzN36G2Y+W2ExYw54cBJMxl7VY9GDKmJXA5yAOsO5tPABQCO0Zw2MLcX1DoREPp
L3wCgNvdpqIqApUp9ON7bAVB2n/XFh/THP2yGvN9Rv3zSJS206cfroAPPmfFMBcqUqzwF8xVrRkH
lqmDEZBCRf8u0Ty/0mpBzA2swoYSNbDTHSXrk83cB6KKzZIqjG0kvBdzqIlQiNqBybNucxLYptA3
I0QANn0IqzwhltcXO0w6zC/EdvOgBsK9rnhJF+HEoiXRvqFLrUO5cIn6S8Ojm0GGMyKUSUh9bH6c
5vpMLDJeDr2j5xQksrSTLEYuJqvnxGSDujGHYq8VIld5Y1lWmifGjb+f2Z7K4H7n6a+9eXLJ7jB0
WWRvU9wthOvppQXqgavUtBWTtnbnbEBItMc9fYBbD/kU7K1M1i35yoc/fWZNU38PTVJK7N5Ym9VQ
waLvA58n/WHYujALTPAwRQcrKF2rljlnvHXBKygWvr8wDVAhzmM9e4EW5ZSN3NlGhCwxBOf/VFWl
x2ceRlDJRBxd5ol1MW1u/yBtdxiBgZIZLIlm/ZEQNNKW/uGhSll08WMpiN8KlET3S1SIWqj2Mt+L
SeoKGzeFGaW1MdBDY2X7jbJL2zQ9AFDS67Puu22F4cGoElvOuLKOaLBrBGYKmbRWVePSg8K/enzh
HNt8lby392MANBcGzVqaH0NQJC0YYVJX2xAMC1/AQsPVn4YjN8ZAJPO2HBeyaFbyAZ3SEvWqP2V0
7XLX1fpaiQHEmmLvS7wt/F1v5qPwmoXIPG8llqK7ngjL6hWAYnt1gOJQMfv7eX5RPylmq3ilGkBK
V/jngYRdL7BXXrVLzQehp5aXO+thXblBfemq1gYgrLWIp4T+KCQ2KhEjWeCgiRWtNnqa6jC3hw6r
9BHFZPToWGYQFBDMXQUfhRoVbYysZyQBSmWTBsdLLjGc44ffC5YX9ZPOh068UHTthrZc43NJv8EY
gafR0zMHvjCJvJlT6KP1dDfkECaCliEyO1vJZHq2f4CV6a46Kv2Uj3jEGZrPTohoc5a2THhxQf55
t5cCJlb00/JK4mJKOlVAmybxUczZHnwdO5uG+zBL+9A9X9CN0dntN+VbZatY7FjGB+tiaYTK8TSC
kFELhlp7Mp3lpMZghCHDEO4RV/4rVqx/8VPUK82ocO6SsVhcXElu5iIbD3/RsVU228TYps71ZNpu
ybhgQUY2P6wDrsFOHAtH7Nt5bHCixh/TKpwpWaZ+5DjROaJ59yTlCH76gowjglzWZjjSMScpTWfk
Pfoy7N+Qey/6urE6xw3Z+n6RX0XC/UP84ZA6dFXQpi5hLNFZaHx1lfkjoiWq+RLvRW31hK6L21ng
tM0f3nfw9hv589I2c03JTHqNWJicxY9jtAuPzn3+emK6BUmAi7R6p1TqqPbCk71646paryrbMrtP
Zm9imgjEvHE7W/6V76uMF+2b2Xj6zJzmR/kPd/02zY4ti3gi2EvN9EkfTNOKKBtC3FYQUOT8N3Jo
3IwClaiW4Aa/I0Du/MWI5o7CcDzFMpmTILWsfsJjp0DI11+uWYTSxxDZKyQsRdWAzL2/o86tej6m
LXJ0++AOoiUk3w7k6hHkVfq0LG5bKZ3ydAd3RL0c/d2zdoPKziANCyVQ6KKedryO7oNdag2IVgor
0PvIFtC/NjJLjIOoDrOywmjSDJ/sS0STkzof4uEKMGDpsEsbz7C8lnx/9WRtqrwVRn7kDNjsiDU2
J47iso9NrZSMroc2NKWeKfNg3WvW4LPwwp43joJEuIFwepDB/+NY43SXZzItT3iTdfsO3WsA1PVS
OjX+h5noC57xaAeMdLyE4VDEDT8hPY2+ATy7tfdqmf39E7RDa1anptWEcIdfh5XlM6mZPoQWarRr
qlTusA5rvQRW5pBK+QKr1zWK0Aut98jXgEZHn7HA1tomHXuZg0czbKwO8nUC6IxpH0IG6bkgv9YZ
YqZHcUdLYGLWVNwKG7kf94VbZoqsp2vShvN37VQSSfkWXBtEmIRU5gk1URr3Km2iCFKjd6MYdFbh
DI+B1PrgLCQStbJoz2aE6TpQKNOfoJMaoUC5rq4L1GUoZ3mI96eSi7KoReUkKs+J7uTuLwH1Gkfr
dRoMp3fn7d+3rYvs08mt/9+qm+vjDE4eqr+pQUpoWV0FoN2hY7Vfj8Azlb3h1qdBk7ZfgUWld+W+
12rOcZFzQr6MUJ0D903A8IeTI0ZwyQnKRihVQ2+5mK/8/uohGs/C+jNjcwscWxXFhQyoCU3vrsXU
yL4HfuQ6xY/G1xUnl/npkHim6Cd93h1YvK5+stxMqaVCtqGR67inkct10hkwsCPeCMjAZdCWx8qO
IW2X17eHTx1jMcuYey5h808FeNsQ9ADy9vK3u8DO26iJgeudFlFvTDjeY/LdNi5KM8g+vP6mDl6t
dkwxNRO5M/OvaQe0HoDBdPuQiG7QigcL3fQr99dcx7ouVBgJMxBrIc0ZC22e5y3X1w9UO7oCVXgt
aSWZhwTxYlfVitkeot3JoOj1QdJTjT1gyExzOA+ldt3qPdXAAz2GY1nhtKcfM0dU88xyX779Q2Fe
IwW9g0BUvfum1/s3WqLAhh88wcjBQ4jkPrZla670wTkq21p6qKn0nWS+VBCYTFxSijeEo6admd/w
HmBnLbNGJmxQ6COoHCTP5qet/fA0HzB6u88WerJW3wPOKo90w3grwJnM3LwhWI1/XNvM/kgyAi89
oXylNm4K3dpO/HQCV6SYOO3B17lPt9Wfp3UZIj5rc0JEVf7/TXkes8P02MVrTbHKSu8HfBCH8NF6
GYP+lW/35Nh7AyYwD0q2dEk5WVmOgwX5yG3DccDXxrKQOE4x43kyoYjWKTQQdsEe6STLET4+gvEQ
yN3YqjZj5CInZDn4uWgJdwIESRUra7XBiwrBstfj73g2YcRAsgGHiBZxLPw+LxbKnLnocJWZFUcy
ZI6QG2sOEQIEAvAIyHJtE6OwkPTfGRQfvWGXHJ6loWt8Mk2djs+K5/c5AlpztV5qaZy5ybruOAm+
+9rJbC/g/lQx/nPlqiMByIS/i59mdtHCGxUg/gogowBdpceFk+3ivm/BONrOtWl466zoVr0vr1HH
DqUxeFh5e9PsQ6ImB9hhR7MAT8SUXnC/BrwwPvZZEBaJ1cZ+19eYmVxVXWQXJPSfXOygmoE1vjRO
rVFjOltEYQhxkptw+WQXcgr2jrXTtoQoo+bsgdv+ibBpEEV/eaY6U6Q3PtBd/vcCt2fkc/5QSkD0
LGG3OlSigDCZj47p0EnfZ9BEGbxwB2P4ZA8RvgzQAQYrxOR0bvl3RqoBbYDdf3iZcI59see5bT6g
jqQ5dSkZr8gleCM68pG2Jf4OQt2E09mLZTyrQKioVRaqO6Ear6SR3rR0K6nBmQJCSHkiwBb3SdZ1
4vBEnB4y/KjwB5dhwSBq7lViCAlGJH0S3H6paNy/dZm6HcqSaX4bL3rQN9m57/AMvgxLby7PSfHN
YjOO0Au6XnLcN/k9ePF7kG3IPLJ8gC3R3qSHX0v290fye3LRgWMONi8MMnaxwkDZO59rD14B5k6m
gkg4cmgjI1BhtqqKRI27Xk/dns6WTowJr5bmpOsxF4R7pq4lA6dfgGd86Xz7L3hvxAgXjbvq1LBF
pMlVRtmOAW2lBcoDELznKo06uZoRg6Xz0PSItSqzcGGxjUITi2yATi9GpieJK46/UTQLQrHVNNEy
7NRpe/IpplyxI4jRh9gQzfNS77TpwuMR/eMY2DzJH+dmHdPzU1BY5izGChrk0AKAZzL5tBtKDbXL
naq59BgCTER7MmEVxMfuSio2rpWNn01lAwcmKz+e3+o9W15KXHQ4ZA6gb99oKOriZsR6dYSHWstQ
RUSQq8HZPAhgbSDc0sFVzR4l0zVrKfeb+EMTxKhTx7qkiEzQIaTld/EheyKegLZfjQwGCaNrKv6t
9UklQ2uFvqqCC5O02IH2s8DHVsC2Z6XKnYnHxBKNGbeyg1nS+dAKdh1rbJinPO8EyYkyH2x2IA5V
1Q6nkgUiDCR5tc9OuAgN9pcX8Z9DjrjUsJs6ckGnWQL9r2inX6ruYfMb3QCdClABe2P5V1Q48FPP
4riGYPVnoovHC3BZsgtjX9axKU9LA+FqfB9HhVdLRBPz9WM4K6egzIjoKWyPnl9uKAWwaNnOZkj8
mDTX984n22WdssQC6z6tfP4MD2Cg8vFlHOg0DNdSRRmDhbFuJdBzNAhUYwlmpO1Ro1MgkjFLA39z
8s6vx72MjzG2h7bs6JKuorqVR1JotOd4ByTFusBddEELq8RtzUYPjKVQzPxtRwDGFJgowbhD4Ik8
asGgjQhEEefLAkfVGs1mC6IyVHYgFUWfN2u1YzCy+TCWe6MQf17zUpWxKqBGnO34R7boVaTBUvNc
qloFEQFtB6fCvdA5QAeTMZBGf+4htl4QBm1eS6kIW2Z75QK5bYj/TrQau6UxHvaL7YGuTGemUg8+
vIPDnGXlhnNCcmvQ6aLpnPserUrA6duj6K5Da//PZTDqYIudz/FUr1L47XOY7YPidLwMuPZcX7vu
34HRY8MHsmMvLteJaGbJCQvSL6sTw34cNa40ZOxmrlRqTTPuwuE5pI1tJhVyCw5TgCdrExugUpi0
HK0kZcKw6F14mIt6oUkQjaS30/RgCqqkSYPippN/qIBoOEV8zGGBlBjmngk5zP9JO0gkUBE19G4S
eiQxIiZdR80RgdXfpdf8tSlzPUaAsA7e7Ac5swNciFBdZkl5pa8hAv4W1DKtmtHAylmVDR3s2wlN
WBfvwtKtsorV3cDHEnFVfJiH1dCkAgqVcGPi8KXeWprwqB4//+Jp+9SPImvRz+QECNsGKZyUErYi
yEG8fMmCXNIY8lCwvJcM56TvOPnydQ5ThnDffgpXwY/bDFVvargmjp2lCnCjTSCW4I1Q6w1Nrb+8
qcOoyRh7w5DKJRt4lAPID1PQNZ21wn6F3tfnr4srI/mb2iBdqrLZot8ZWC7r184nM+zwnrXUdpXn
9xW+E0+d9IiC7xCJY4MLW4fETRTwcX0O42VmkPreoh+N/ewcVNS+Uzn9Y4E6dqId//XtXoAwv/pn
xVL2fRvbn4qGXCpk+KTRpuTDMlxD/KSTk2hewIO/KamvLv9PT4yycl5TsmcvCeeTOaiGvm3PZL1E
+TRZBp78GzO9+ypt+Fi9XJrxpt8Rry8uD6vQsb2y50HFgxkwdjOzJ3EIkj8RF/7gDqNjP5vkP4om
+iu/DuNeQ5jkVFDhzMJWYrUt82RU6ehxPWJlzNZQlZpVRWUZLRhU35eEPLbYEOkc5WMLL7/lMq3k
xdfImFlNfQk/OYmfP5875bzz0qhvt2nsBKdhwZEwCadag2Sl7m/vYQNNcRRGY/jNI1H6lPVr3yTX
qa6FmguIVnddbLhFAIx00DQYnphWedbqCHSWyScgFdYSD0CCNa0XR8EQRKoFBke872PzFVisqFgy
SLP8xwM7jtmAAxxlP9ier6kAbIiH1R60RwMjNc2SxgsX2AG6e4fqjkHM7iNWX8n6BMEqTP49le0r
DwnzR5bUakvqKfSHqTmlE3+/YsPgGylMc8Ny5+bBpxVujer4ivcxeLREnLOC535FBldW7Q7yYzFU
TLluvQup+pmpUOW/MILfpuWFr/w1AKA/WOEXl12Hwl7LUpP0fonIfgDtTtUAzY3friorZBFM/uDr
W38LH8pPlwWK6nl142TeyVHpQ4luiowZltz2IE83wPwEeNcac5VwPKrJY10SB0xqAo8eCOie6YAD
XcHbe6dEAjjelKvcHAY5FHWiKhl9YoRbO3u3OWAzifgi512BWDXXaKw+77YMA9w9ppMxfFk0jRGI
V5FwwTYs2GEeknZTgET3TwbAN9jVmXDQiPBK7EICtvBkq+0QjVrMS8qK1kSGJhHF82tafIUUoIaK
jBbabJ6bw/JvKGie7yjzPOrjZfSGGF7R2jEv3bfxuxQBDiZ5uMOUjGlgOiOI7EvP86ZO6KxmqAQw
OA92rCkfC/5Ovlpu1ZYIuTeKrfpbRkFfxBUoj5ZigtnLUF/kQlx0ZCS9dd6it0V4gkyuPmS9QDQY
mZ3jpmMe0PVxamXVpUM+KPeqiZC3LwiJIb2mDcPOkRvHoCclmun+gww3FpQkUUtYS38oT1dfvjg7
aXDvto8ktiZ42ssZGKRn215OkQ1TGvPg3d9MUxBeDUC136+gJOToRX2qqgtuRS/pBZkiJ2cy4kKW
RkYlHEPFrvruWnfMiNGgrv7mUv7hMw4ML1Vd8lk1YnoADF+m5GLkR/uiFa94Fpcaixbcy5A8ndwZ
R+3EGx7vP97xo8FF1RWfQ0IODwqN17P5MTR67Wnaq3NjeeV+wK28SMK7wTzzkMabQm28R2HaIE2A
L+7uVQ1bAFvY14zVrJTTDvWU2zuKhOJE4ZC3GQxirLkdjcCW2wxAi7gLxHEJaHL25FM5t0eKezeX
6DAwUWUYCfhIGncn8NpehxXtNVux3zw4NJB+KfmVPA5bGLhe5bYaCE7bOl9+QFqxgqMPt783Aopp
Hck7h6X9exycKUbMcNsagDxHQ/yNZh4FCEWKTkQNGXnwxLj6iujUM+kbC9YAyNVqrb2/Ahn2qQqv
OTVsMVb9smz36vt39MMwU7OWZttYPo8uAO99s7YMcjf3fVFRMuflxHYEIeEAJHKhtFkn7KSw3Uhk
zU1ZOYFqC+PmnMS9+9XQ5E+OtmODUCgUDoMd6CdreF2uV6KAYmqQ7U1BvJjTLg0ZQlsZ1C4NG8pK
MDHqqghn4fa8BYosAlhYmd2lf8voYHjydAKV6hFaDOOu9CHBMKrZktJj+KyqUZ0eSVpqNdl31rpE
nHCh7RPXZXV554Qn9RN+TfuKK3orzHf0GLPeUmbjZkno++xgMTdWrdaTmvYdZ4/z/nvOopfHz0ML
DJKx4mJUo1fqQm5+vcbeWZqZe3UZDn4qiFoXy4A9Ldwno6UvUCRwrUvdtqq2U7oOBQiwv+c3eawH
RbIF6A70bebqIr4H6HWes3lA1feEPB+xbZ/5ADrkZbtS+kzsiE7yyl88/YuAj6+wAifXLbMSu42o
0Q+0zzY8wxDKSNER7QbOH7krzuYF1+0a48OIvprx4oFsFinTUPneui8Puya+GbDjZIkRs7ed6teo
XwzRvnD6cypFvjtlnHqtpTIgB9PQHza/TFWPnOI7xsJb9JEUvQ4TqvNLFxM+Bzdpf5lZnrV14LiQ
mCsftb1ZRjXjD1w+Qn0d9cLvBEqFK2OZpdCfqmmPAHcwgxyiK/KpjBNltwZ8hdgOreOw/MB9Y0Vg
nww3mPIohGtEEHomqjtcxTu3K9EYknFy9CrtY8o/pfop1+xboWuNNfbjyQT4p8XRab2lcq3DgPB/
r5/QE2IXQiS0Bh0o5CjCcEAeyUdr62eVNfbMxvtsS3pnd7ml+zCwZh4QtA+xNZsn+jCeVzXuWyNV
vjk9LM1SrlSpR4RkSd69cpXBlWGuY/WeMxtY0PrnsO5Vjm1XePQUQNttcJy1SgNp+yPuLXw9VVov
eYzLYHTo47+gYzhhnHuD0aTcB6DVL+bnxUoLz+weTZMWKs5jZVg8EIF8DdW3HUWUBgvfOqfw1ZkJ
0xkN8qi1T6+Qij0aj4V+tsUb0wGAZHfNnsfJYCBoxidWuT6zvndvN8Z8bEAbTrdmxGZPMzLeoi4C
oQ9e+OcoPcKkzmf+FBKO/A2pxN7xhmSDer4eUi/kuWRt2C6tpKrhFOjbD1hPP4DxnLZTYuJ2GwRF
vNS3Htkj+xlnOJ5gJa4l6fACrNIcYgtrbtrYSRyICkgxTIrxIH2ITP53yHjZogEa3eto8qyVEBRD
plVCxFdPpDmGLApGnPe9Z2cBsjTJsDS9OVJHdGGW1X/3T103r9s/EGlR3p6SLDflEH8c0tbZmQE6
/wxSYjrb1bCQktbwk2OP+zPkMXQGhNlIQc3Q84uONkA72LcrANsoLMYkL3LQ1iTMpWF2ff2AM1h2
gWKoQRdgrdEpt/AVSqrbxN2RddpuqHLwiyz4GlS6hH7WKFjMpsOqiFt1q3/dOr+bTmE+Z/1Xtb6F
Rfb24sT5/Q2SVjFgQtzTdXH3G9T7K0tqGESIDE6Si5YX3FySS2YOS9fUcOVLVuTOo1+sixhvfDag
EbA/E8RnEb7Wpsh4XgaRiuOmEeaUvK4rcstqDkI7PreIbE8ywEqe9iJB7/TNhnWDjjH76ceHqgW+
HC1wKruU6lc/6XNFSlJ4kFjeEXeVQWGo8xeLicmwNeLLmzvPgJgvTP4BQ/1m8oobyTJ5Rg7eNfP8
cSIq0UJdatG8XZbcYF9jkC35Rg+SyujqaiNpim7OQjKtgT4fbk5R3YJpRLgvu2ypD9Z0yIg6VZfD
yKaC2xgRRqvUmrZcHvMzpzc8FDH2J9VRO0pXCt/BVICoNEzwoDm9xju467e73J6ZIkUl6tBTOMnd
kDcnsEUMdrLaAMvS8Zqqj7gBYELsrn59aK8qdBymM/7SRF0kqNU4CQY2nuCCR1uDx5Z3nn++ZhvO
1qCcRP5RVsZyO8Jx4V4MpXEubK5ex8+QC/CRpyAkcO/CHuz8frxJVkXzu1Asd4eQuCIEXY53n8ko
b0fxysms1yINntGOUU2/hwAOX01964tnOHyEofJRJHQKUOYY7DGPFKXufu28PT8SVw5qMFvplkyI
vzuNKNTYRwmoMlMMQlvv0FyxCNB5bl8mQt6ffAEMSBeZZm62fzW0Q7q0FRCt7YAH+RXD+yozBG9M
jMqzMAM8iJftzhPM4DbUGVxTYB+IH1GoGHZ4wXkUZpcEUI2KGbYJ+cv5hO1AqMYmuyyYNIUaTuys
TeY42k2AZKGr64esjY+lx9uxhK/WCsDJBZBraoybjsAk5ZKFA3s4UmAzFlRZHfFwLUBr1cKjCZay
hFJDvh76mG90VxFVk6qa9QFLu1IitTsTqir7eDp8BRIA3vwvuuEa/IJ7WDZjfvgaCEhV+XmQ/54q
DGrYYVe8OadtH4zPWRZLKdpM9W353YHFeU2/uNcs4PU8FnSuRvMU+s/MOdwYsmirOIu/pLNde/8H
BBJhMqE2H05i/A7w1hLeuLb1zsgS1Sxm0L63HZqYuOuudy1DZ9SCDuOvdMCWwt0348E1zUPTPDJx
sqECJsKpjwBf8O6JamHhSOMUl+L3QA3Q1H3T372TvVwCOY3hX8KxrQSVdRrtkxVMupUsG9vvUYUM
dsFq/J5zpID7oivx8QAWz+kItWALSt+WtURrU2qo70vbPTTY0neUEiUmCDGC572uK+XvugHI+w79
2YU/q7VkpaCSKN3n5n6pbXYA2lUgyfUmB1A+VfCMEvRGP8e0O85HEGDFjc560nkKmuX9pUf7TGHY
TG2SXmt6p7YvjSva3OIBECf0DAUY/CiSIObP6DLm7vNz3/QEVRxjc+gznIIjm8f9WRpxVpLFUyhq
Efh2gjXlar86qyVxfTtS9duWoaYJAaZiCN74DahnxQBpqXHydRkaao669cwSq9K36kvqoEIA8ncD
NsoTSQePaRVf6/MxUXuRtzY0iuVgTOLk6DMwZcT2pqZDic68eYvS/uHnvTGN8ZP4Gjg1EKN6nHR0
FmIzMzfCgFBhxPsDstF6tZZga57SgU+W5zoa6+VSMjZpyAGZZeE8ES261VPMCynSD3GyxK+3dnfh
Rv3KSRd2FmXlI11n7RCnrK0ANwoM1Ct16ngVi5XxxwkDfcNZzzmsDqSFqiazubIcEqYseZzG7eCP
/tpYn55xQhyZNYyRC3kpk7HKpxFCyc9NkbKyzoL38rMvifMEt/giFcCjRTkEb4hpECWdxSJiugnt
zWrGj/1VnF3hqUiiEhsvg8+jaL9yZ/qTMg/vxYbw7WD/FTt2A6GD9nEyT77weudkNvy8zqitpdWU
DFs9N9ccrrzl/AZRktkAHn2Hr1E5GH/sICacjvCfF4X9l76dJOkJTSfwbaeiTcgxenGrLizH6wI4
hrUSrhEWbH4SkdeA8wSlQX0KHqaWHa6kS5EwRy8d0gzNecN0rTFjAxyXKK1P5vCGl5gA7NAs6lSx
NWr70OHuIglj0VAnZO8HHSzux8LHCW6HWat385KkSlNG/Ou19cfgjPc7kophXS3B3w8YMxnNm09C
cBdVQ5qMvgrVy9NcHInIWOd5p2cSL/725H5msognt7r5BhcjYibny0EfPg7S5TGzXEnx7jZ3guEn
TGPFD8ZvP/3E/kBtaBIOPGDjKCCsUH9e83GDUQPbnCvdj4Oup7Xdmz1BlMRSljnBFU/nBrZSdZO4
PBM5lar7g726mBvAO79pl+ehqF8Zt4LsP5KJMruib9+/KzVPrszmP855lmCB2B7/txCp8IZuI3Cx
0vXhCTWTH/aEfzKEc7HvtJnDdJmp/oLFlhvnCA1bGYmqxOd9QO/Oy0oexLOQXAp+6Hhj5xzqYvPm
TQjbPmsllnfHmHIx9tt1oZ75bHLOfggXTFQcg9zNb0mgNdokj66eeKHeeM/UTgxbmWz3i4ZFI9nn
DJGi68oHirx38o8JvO75SBLeEY/BqT+Jxr31x6mRT+ArOHVrByp1mrJbVDZQJrYyQ4NYU6RTLpfa
GqqKg3DODuZ2xMYmNZMt34drwpvNyN3U6D/k7GFTExV8VTKYkGsbKMZc+t7qzABo8bWLcgMZ629U
uFSHiVH9bRaWjiqwhuO0i53GJ2+Uk2lT20gnjagrdHGHoCQSlll3xqcL+Ce7vWYvKGoKAi0y9pC3
ATddOzJ/EBtn9lnXbitlqnOO2SrWRFvvdQcFA1fIiFhc43J2CZ3vXHgG2elJbCXbs6XhAlBADovV
HFcRb+YSDLurTJylD2WsblG+sGKmC+l869ixaoibkekajcarDF3RIganENvP8tmrrZBAYfjXOJWN
ANi3Xj1xjHHckz0E/gt9EHDXDkKOzMQK0HprBw1KltmAMFanyDmVVnmfA1sY/8JHgP7UcWfoqAGt
pLbmuVHea2Swz1xvFBziVCZ3s7YJfH1QulMMi+oUiO6hCm9TL9TBcv17D9Tms5JLBt5EfJfyJ8EQ
bgxgH1gLQnjjohEzcfIPbBMwEXeqrPqlX5480eVFR00GZSoJdltnY4281z7vvifBmkCbo3HaJN2t
gLblXgdQM5VQsbO6QjTWWRh1CxwehT0IOonpUS/Ed1Xl7kuDZ84zi/mvRFOi7sLNETEC3YSFya/0
cJnoRib9PE8GUL9k4R97uFs0QbcleycjRtorP8wry7M8YdWokpCnjVeksZwnljAPzEAY+VGFcmgk
YXGHibAtVFEUifwD5Us/+8bjqMofBJzT3t7saZSuGWb182J4LXxUy8n1/ze8aaqiRQWMLv4KoWs4
/e45XXL7HBZ4z1yDMr5aU/eaJOiYKwgrNScNOHOqNU5pHliURL3HKtIbxUfCma5L7BwEZMR7axvO
cLz/qrYkWYHG5KmA4XvDL7Hk9yQI7OfjxUa01d/it1LHZP+2KjqGe/fQImmVwHJbsK2I31oq4kCx
2SEmMY9CKPm75eGy++gBqyoi2kS7ldOUDLTdfm1xNsox5SQOIRt+l8BBkaReRAF8TjJ67+r9zp6C
AMzkLq/SnA64QmJ22DNQ7q0yTkf3A8wqrRBGF0NJrLszy6ebLREDvztiX9ikNw9GzkJR19lUP1da
Y4cwYPWbl/YZ1kt1XUaEgiaowoXShn2rSl74oLQpVl2J3sSd0NncRhpHBKyR9gXaxqlJTGTy+oM1
dqdw2Ls6SQ8URmJ9P6WncUMGLrU5QHl+PtHbBpbcASa35dsGbpHwTtmNRcffMZbe/++RX5oGBfy3
EElp8TyKI5lVa93zaohG7aWHoXjcelSlrVXIQV7P3Y2XLYlfCa1ny82R2B7KwRQuTfzWucZ3b4Fs
g1q3JVtCwh6fua2AohnN+Sng5rdYJ+Z0l0UmzysS/MIUG8ZL38/SSZ7qIA895FWIX4+G7mjWhLNI
Q8BVwq4jHlbAF+qfzQf7Px5+Jx/l/BhrSkakyqvNEB5NlFC8y4jLgUzSbWUhi6BmzOH1ktI+Og4K
cQpqYr0yEq9awClH0IiA02OLVTethXUeTODHhyK4orDQSjAM2ixW0g8puBJYSMip15bOrr9F5c6A
QNGSgt0QsEVmuIBpmVDSkklCsYlE2YGvdIwZTKRJf2x4adRqeAFyQmYrelEvA4c8JNWuwHDdOVkW
SUaeSYmUZwB77Ax1XhvNzc08wY5+e6NGJJXcErTtiTOmS8RcikGjD6NWc5baqLCL1rjANpgu59Zh
BdfQZynae7a7aWH6ndiNGXU3nmf1m3/+hO8+T5Uew4ZmEgOetBT4cTKeRC89ELIYKsZ8RV9eMUfh
SKotJLYD/NULQpiGu56yFNnvATlhD1ykPc05EDus8HHDQQaK34HGIY/djwNiv1Nj3jbOpw/jDej3
Ssdj5ipbGayatU2iOxPnUz+8/jbkYBpbkvzwfogz0OwswOqIfinsKGXZ/oMlBGRWlcuGNVGvAdMj
ctHI1dkW/GjOA2LkggDnXp7xWh65QBkLfsc3IMRy3i4H4C/MN+Q1XcVZh1C44xPfYAM9pZDfhwEn
fV55GUu7ujsiGADCcnu59cdRnk+6UQeau05V01OCqyeXZ9YCLmdpuXOtSsSFeejmR2osZ1ridyqr
gbySjsGQO47K/5UAwrZQtRw5Ua59r973j4A2tFz3h7L2c1JmRH2Lc9NyANTF37I2evgpZX/hPNrM
vRFcve3WtYfpgTlgD5TGpT+fNeDUVUpRXxvc+70jF4KHwe7+UwSBvmnUaEESNctN97EHrZ3BiE5Q
AunF3H7uLVA/GN5HTN3X6F2q7I6Mzbblu3tvafWy8yxrex0tu0kRmSsDyio0M0T5wT4Sas+CU7Iq
KKiY02j8wXwh0CXlThfBTyaT4iSl0Hr/Czpci9rHH9LjjrGfNdPn5djS5NkYjL/P4zEXIwfXGsGl
q6xt0LzAN5qag9IH48hhE2wDM5+wNY2WbKLVuVpPLd+z1YR0JJB0YL1nfwGVfR+tuuCFFGYe19B4
N2EEV2g5YCRDHVsjCYfyo89Wn9Qc4VwIltnj3VL8asQs5wGLteDIwc3SM8DBtUazaiSKj5xlboMs
F3KS737Is8AMjdHhE9HQn2R0xMww4h7zWYqCNorm0fgl2r22camtTmJ3QBo3+h3bP809lZp3ktGE
S4jAT9SQa63lOEjc1xltfjn1aigzPfI8KoqqH5pOSV8nZeWVa3NOWpS32SHCCmtz09naSoMzZlnM
uWG+P/UAvW0DDjLhn6REjz86LRS42b/smd51FlHGQTgIJIoEBA2Er5rTEQdRu7gp50uq74s2iFn0
lNS1TrFs1RzH3jV2U0WE85hHeB9+YY+W+caUe9+RkavOTQtYKnM61biPNKuvVCvwYCNm59SZtJj9
eMuF6cxs0r+scAUpr++5xZ76mZZIkEcWD0KiF6Y0RJP1ctoLQRMo3cZVYmgKQgHtHhdzFcU4lyqZ
tw7515S/HLOWA3H9SoxiPFXd/poPkOiu83vAtPlkYt4UBR8qLkoN9lAr5o1qGo4IleeJSploXtno
xIHe2t7Ix531/1mm6K5GbekoKDHBXUpJnrgMC1UcwY6GtODzgNUqQSqDlDoPGjHIci1HfCxmeHsx
bWmeLRMJkTNtVliz2urCO9itKdKZRsqKutbaA1b4FveUw4SnXA0HFi/gdFAeb+RRHrpFt6ftPIDj
a8wqICKjr15AcNMS/eT+zAFljlpGyhfzIQmByyy0pUJi1ayh6nqxBlYdCXi4qbT17oV+XS+KFs/t
ipselM+J/jdpRTRQJeJq8hyTsE1aP7kpGfolnwgouT6ua1rn3zwMIZ3X90nWPxi7o4321tzs1mXI
cLmJU3x1r4Nf6xm7V7nBCKof0a1od9DrxT4A4HSOwoDfSgEbXx8gK5Kz6ZkCHclgUfr8RO3WYabY
FSb03+GUHaYxft5BqHdy9g/g4XBvmZ995hCF/cnl5vjx6rB/M9LvvCFSetRUYIaVBxkJ4PT4vgGD
dC9//n9eMbaF6WsnEcJCzDczTFH0tzeI5JQx5XbpAInWnwrPqjwZPehIUnFuFMVQV3Vfo4DLjH4d
/4Mw29Zg1ako97pYXNZBBLNpIx1o227aGBIoYGrcPDta+ZzpZ8Gu5LyniyFeTJ/uPZPLqmAn0qLQ
Xl3ftHiRlwp3wjg4LMIrVz+IdTOe/OKDlETvSnNuSRKFDXePrUB5wNzgbwDrmHxID2wXPp+618+z
IrHGLClfUZTxCmG7FCRWEFz3E6pB+Tg1pjsmq23B7WnVlxmuaVoepEGjxvH7TefqKC0srkBWuq7O
9qXmDEUMS5Ux1D27kP/OharlwVarPQirzEk6Gde4C6ITBJuhFUP+dtAkrpZFnk4tlaqwbppQrVYC
lx5SXJE/4SG8HoH5nLm1pWK+a2+9tM0eYo4ttv/HVo6GY2aDJfgZAhD3wUmkXWKOjDQfWpZmJMU6
yy3sM7cFUjbBWZn8DY5auldRlinqGVyMtNAucgOGzmkc+S0qOPngSXqpEu5kwlSRvKsUheP+GItU
l+Y8w8kCPilt7uxbvjfQyc48ckBRlVv54/xOnCO8dfIZPKoAXiLGhihcLJ/r0bqD6l3JsL2uP6Rw
jhypU0R6dP7PPO7o8rer1Us46od4EjHAxqnld4HAvjt5yRTFToZq3p2HnH/K73/9GxdwXYNTsupF
osLA/HBRA+SiO2SW4KFCVb3lKD8i2unxPnJzykyUZS8NjkP2DY8G/0+/7rl+n5qOb/Oau98Q6Xu+
dA9IbQmWaDBPPTdpiAzwNwv9Reus5TLWtozLOr8R8kAsaNi301Hcjbkermck1UcqzzDQf/kQNYVc
WtIlB5A24OwhpvVHJLiNOmteNSv/von1Frhq11qriQzp8/Crfx7JY9ByJpy+6qhPNWoZ058ZkB8F
lCRtUI+EmOHdjbc+Mae0WtmH1A0piotXpSz0iG7GNWHnksGt4lGz6Ypo9XZPJx8rGsvtaPkXOv+d
FnXNjUzACi1vyOSVb8TUU7HCgAZjwbVlBvaY3gqE7KUfMjuXk64nphPPI8aELftc/GA8ffQF/hh4
ah6PcoGAJo0fY45UHQ2dJFsxyHlwNv+MSRp4sGJSG5YdYNnBz03OqNlvKyi0SM+Ydt6dnQB9c1II
k412F+L8OU9c1ii20RidiHa8sPD7C5Wb0qtWpG38EanK/9OIYYOEcgI6Q2bkSDGRQoc/Aiy8aSxj
GUgHNhBI8pwy5EyHflajH+SFhYl41LTc5fGAvBXMPEE/BVpLRSRU2j/iPVMGODbe0Ny93Vrtg8Eg
UAR2iQCzrnfPng17bupgzOeNA4ih2LNn9fytYyhbbKo2hmhVlNZ5foASNKTU8A9IAXUbF4WrXbi4
LZ9FiGfsgJ292Lzl1SGZ9wREbf2hDDMYZAhUWOoOOGOZu0yXnObd9I2Beb5UO2+bxpieKMYcpsL5
YlUFdvai/15/s/WAn+Hf53zhywves3PftYO3+WHTEHEaZ9o8yfPVKanXKa+cvsZFu/N6xTRxo8b6
t5udnOe3Ljpevz+Inv4g+07N/EuhC4TAMQxAI/WGdsB39kzWdXF/2cbeFx+ANrGP8TXStF9Gh4AY
M1WHen3LNAhpnpeMbIKBP/eM1lypQjt7T1UUnh7WWSIRmUnEtZzXfRJGoGPYofdl6ZFjiBrVTA7n
TlLcn0XgXeuHSkauAfX/8Z1RavQpX3GWBKg4xjTeYAeh13I2GAB6+qkyaqtTP8AhCO0vcRTaezSj
G7N7hJ0Lq5pWZKi9Bj/0w+yYkVf6scLnkuM3IKTWoC1TRvR+qeno/aPvbIccBPzGCxaA4Kc8gTmx
bsNjGAzRH0PfpVGzdnoPyM544YxkJp+r81zkVhqC0rGZKOYLiIr114GX7KqpIhI8uQm7ej5xYmWg
4paeZktafv43lQRTztF2bxtdq2VDYqe9K1wfgjm2o8Z0wBIfOIx0WZH4m/v6BvMSWi44zF6FKApV
OaXPADc0EuxOu9sWrSnsjQ5oqiRitVbk1p5f7iC84dwpVN76Xpl2jsl9DPooyGuzhqFIUl6c1eXs
7sXf9hAbdMlkxiDvcb922KppMaNdSJJ7gknl9bphgt0w7wUQMj/dQcbD+akLic8e6iRT6nWSLmgF
VJZAsWNUtpKiEBQ5kjphPhl+NYqIMcFZiUe7I2wry5v5EIK7OnhSz6zys5yDZQj1SXAjZcyyzk0k
K9/voWisSNvcFJPzohD1a/5R54UERzXHWiKC86DRDkJZFj23YoFjA0vV43NkLYKjwgLCHDlSM6wc
PtahymIiebNewcwEYS1u3aLwwDws5LibZDoDG9bEMEwVRi6jMEcvNAL4gGAvBfw08XbC4dKWzeF5
NhHZKv3vw29f8tX4CQ0sh/B/RYZhkfxv80m1uHjlNXycn1MgubMzkn8pb6Us60xzOa3T+wB4CGwS
j8YCy/ZqlFICG9TVuScJ64HDSeKiV+Asc1dLv67/kbwOQ4f00/3Vb+s5/YTnfQUAImQjcQJHDF8i
d0Z2rtAUWTWk9IqebtUrNbygxCK253vunHYzWAiV37n8y+iDEYZ7vU8knX8qYN4cN7RjchFR2F6O
87fFItOvAcJCQwS7s8IxdWTMnz44AZQeugKtMnTiYu2P636qda3M82jBmn71+pdBhragKn1cqnVQ
XaPXQ5zzbrEkaM44XkmYWua3IU0bOuuBo1o4ie5H4rim2M50CLYxSKBkmQhPvaSRcTwgADhI6wBK
F2cdTGatptEkAZ6puU4sN5D4SlaG5JasyqsGFl+pyoQ44fNkeK8+lsR7euoTcsFapsOE54/KKu24
DFFJwmrqyzL/GL6CkV/kezQOpTjy6Eh6Cj+5UN3y4+jhW2dP+6M8UDdc1vYPG/OEN6U9HEMdkJFa
JMe7/reL/8VrLDtUJkHaNViiZCI5Ni1xM1Lg2QgN/jNxhX2EOpKMm+T1jDjA+4SsFBfhhoJgTm0D
/vxxR6KclsSQ0/SMdUBb7yuA3n1NjGFRnkPlogku9wSSsUYXB27dNR/MPY2gecaSvbLQqh5TjZ1i
mOm+aY/q4HfQ1RwBwqdZu6daeCJZGwdYKjbho2ohrznjrHCzRHkXr3cy/3t8YxaazGk2++VLync3
l09biPqX5PcCTvc0TjqlEIc6WsDTw/15z60w+l31O3ByRVPws2mjmHcnIM4hmRcvBv95+vrepfP7
pL9IBejvh3FkD6qQUWrdGdAafClIv0F818GYcfV0y1EBV4MHKTnz+PbWMp9YRhKKglQRGuER8dL5
E7k/hrG/y+vBjzyE0rxjKF+EatByWDxy+vhPFK67jQO3OiTmT5D27Qll/yynrj1b/doRowUjzQ26
zFCTqQYz355921RFSU8J0qZUh0ASIxZbYJctYWKI7cfDUvQZWwUnQ6E+7LzN7vsNPVKRaaRooDaJ
3aBHLw423vNp7Cl++6ZMrsxBycZGelYa9MyGoGAoBNminH1Hw3iABG8GJZBma5uzloJXfF9l5LcX
yX2czisQQE3VrPVXFzbu7qdphQG8NArOMDmnwlFiY/p3yg+ZWSUZT+htz9uxWFtBU6lJCM6XqO5H
aqi1XzBj8xDUgM9wtrKU/BsDlC5d37qG5XGnktyVfbvtC97MNE6x1VFo8Irhee5s7Vp0w77Z4xSH
/TfayodWwjqN0Vv2kUhjbIateUwKWBSA7B0LE/LISUX8XbycYve5/TywN5BvCwh00+2jM30MeBlL
HLnU2s5LNX4amv8GfA0uNVWocafbBN7gt63nZcCpfzQD94soow9czk6TidQZFbLG1f2oKlsrb3CM
BUeDiWa9Cp+emsh+1shJuAMr90/eSgPq0TEfuVrD2TH1XZ0D2Ag92zutK3+HyYawldYIiArMuRTj
SAdzNdOP/7YSCAQfwxQC5JhzblXAlgGGeSxJdCOSFqjJkAn4ssi+goMjuDagOVaww+KEGC/6is+v
MsPj70usIzQ6AVShX2uIGHiey17F++w51ZCVGk3RSJfu6c0UtZCsAzkTvDMwTcOnLQFZ4cGTa7gP
FBwX4euMfwMDZC9gxcXkJE5GI/Rs/SpoDVHKTFHlDZYmNRLw1kkEruH9sqVdfKO5rSXJ4wYsDKYj
c1l6c6RpL4O6tGqoC7TvEgMdzTGt/lwlOCV3ar1EFrOLHQOPYqVmvjSKYLDLJma1VHHLAzW9gRYs
YyyUtkDCeQ6smgXMOVBIzz+i1Pa/zGT/fZwzkyrVb5JQZF/JNo/+cqgprO0UXtx1M5sqyXpE1Aur
V3i1WTVEXpi1dnJPIPR+5SUclWKgRaxOvUlaungT8iXvMJnMxKFCKhTJNJdMg6Q7DYJ32K1amsaO
ANtfH0zRxNBBv0lMZrYKl3Cf/iFQHKqyqeo8TDOE52eVA6JDx+mGnukHM3v0xwbJ9+YelJ0GMSF9
upJRnmhkdRdoCtw6bV81DrSQls3zLVoW6lO4V0Z6LfKbHj+JqZLt94mDSTOetLbmr5ssSQVRxLxf
+L5wm+c4pYaU+nQ6xYKs/ir4Yvy4BUkvcaKvrFfai56l1cGDYB2Uxghu3irMaOjTwVYMBWZ8MU1I
Izl9YEaE/G7Hm/Zl1PxrNzgRS3yURjXNwxuHd9p6oQp+ePR0vGhb53RBf7rRNHZ46jgEc1i5Q60Y
TgIkgtdJkeV71CbEkYs3hteacpNKssFcn5u0M5Xm+ddhgw93ZMaEB9ezmSLJi3se9YrWMLUTu8O3
bVJyQ0zxEQAM0hkJauWEwDwyitm4WeFkQQdGlQahyTiYVWWR7X8WJLAONWeVGWZBqqmKrvAxm93V
wupLMyCKI8gT0rB1NOVL9F0v7AuAAURR6KR3LFtq4Llj6sBZD1gu3N1VCIU0fHSgtSAZRz1ZDIz+
DxQXkXsJ65uZPmSPd4ApXG6PBxRjvyliqiktgmbWdq0ypzoXNL8BKGWaJa+cGqd0DiyeIIvv99Df
XqbR4m7rIqIpW57JQZ+4/eFtub1OfigAtK/AShouZzQkNXtB01GeZhUk0eGyf0R3gQ6wX+HYrgY1
c2ueOv0ZJbI8wKBndinm0WPsMspSO8fnV9yK2qo2c0+b3HQk1+tDO4Au2SHGAqyOKlgubEM4kOoR
0ZnOdeNoYbNbSFBzVGHB2eMNi1wmYvoIbBwxKFyceAKKjz5k84FikqwMx64f3P53M6lopVCnbtY4
0NCzXsFCa3rnUUhkEwKlWR5m+GekkNBGEel2Qk6Ykx7fxwrbzmeDZ08O7KRq5bjXURYqQMf4ybi4
qZ6bvTXk6A28gbCAyHOkvZsW+TGgi2SNfNy1mqhDlME4Rp2m8nqwMbjIbLqyPPJailFY4k5rzalj
+XZj704TEZgEPz3QwoJXrGSTCP02YACx6I5wk11BBsZlRxyYWgx4LJxl50B/fE3+PfwyjFl9nHvW
XWmhxJlNBVOJQOm2amHW6Lcvkx77zXmlT8au6jA4i6PlPMsUhtdMrovYYeZrtmg4o34fkC6QoyU7
k+3ylERC57tXqms717tQm1r83KnF3zabIwQF05wTpW87ib3mhhZMECMiQpZoyEKx8LljuA1sVHhc
PCOC8+DLanLDpmswuAnzvvfRLIibe5HMQ7udO7TL3Xs7J9run4fKSNUbAUqUs+PcXdfbtflySQ6V
h5o1QCEi5PqXNItdBMYe46MKe9FkfTEvA5+yV5vC+i4BtiDrWkjD/qerzDADYxgv8CJmLWfSORE3
Tj8I2nAom40RRS6pyS1DJukCgqDj4IEX+Vb1YXQD9THljgdxErb5TSsm+/0Me/PbGZ9W9t1woLQR
jWkVePRjHHS3qJlGFT5BvBuifRLEqlXmi0qivlBEeaJqh2Nn8r2ptyIaoqzWIEpKvwjixJMS4RhX
vZa3EQibLvmMQJ4bOSyDMvvdPhPUxyToHYGjOxRb8gsBFiQXhlwxrrrMZMYK286otOfYy08kGVjC
2Wh+Ok3p3xJ71Jg1rKmBna5B65IuWHCvP5Cza6a6JRhJ5HckIma1fyQtOk1FSNzxZTewlDx3VGba
W0TX9LmVGypOe0QDo6KZNwbZVZl6WkRrHr4bU8BEkirpfUP0JLH+RrVbbEFZgdTTUNS9UwuKLIjq
mYmnCNvBybIJuR+5OgTt2o2/VtHXZ7Qie/iZlgGm1YbWeMdzPqXg2slUU3bUg+7lh9DCjsg1gLJE
HeTqdX61SLpNOCX931B9+/B4iVVRuwtegulTs5pupqATdxMzNM1ECnzyrs5K7FRd8I8XKIVxzZ4u
J6pT8zaB5+M3+cw7mJ+LAhChwNYtBmROmes4I7TLXHRUQi3/HYGD23TZmXzuxF5+BlkaSt/N/nIP
cXQs5+wksIObhagZAvmJ6n253SDb5uHHr+96iONL26gd9l8xxIFhb07nj71V8tIw/4apJ8+TW552
G0eB7zh3dq1WifMyyI7wFpC1d0UKMneZ+F8EqPH9p3gPA0mhTozb/YYbcxR5xcG+NNBDCDcqJg4W
AUmYhJ6mcwR1f5gfS5FdVp2TWXqsDO9msQhHbUeBnFdeAiFBYlgx40UgVqeeY7SJJguAPUnvOQpq
tG6DkjWBp2s5bgtqcdnBmaef+dCv2xoxHrHkUBbGF7KKEjSY0E5nwCw4thOR7j33Dx4MxRLgImlC
TnEV2PqrLlbZ2B2JpTyiooF+jgwsbiB8k24XqOksZPCdHdC5kW2NEwUYDGJhJWY5FAjTEzHT0p7C
eslmxs4+cddSXzL/W8cO7GEbtNo7QqjSoqZp38cP1mRH6pltZoKUYXsFgI3EPzRmF4xjnOtD3noL
7vlokmMp/8Xu0byAIYbZNdAM+ww3OxilvW+qid4iX1cjiOFvWCEIvYLkFh4q81uA9qMA8u/xgZb0
Vyq5CuR1iIIEdZpfYu3ZUH6Gfv6n2OR2b1/Q89tRTRTPn24dAd2OV4mteXEfDQdoO/4hgRIJDuue
FyGOuQpQrNtGjETTfqEyfnviOsYitQvtF9PQFaJy+ylMTmru+H8k2J2Cn3XwjbRKGz/HCDwQkcpc
48eE25GPj+4MWB9rGJxX6sPiJmcI0v5j6ZIuvrP6ums/nLM++PjfzU/5a/65xqgmYK4bIR86HK/H
6Djc5qXFx7/u1fxUtnmcMvoZzoOHZPVYnbHqOPctAMexFPqolB60qE5cvmAyMU1I45qEdqltWLxI
EM5ZeouHsnP5E76KAyRXvpuyjTX20eG7EyFU7FF3F3MAnXcciptI8SQ86x5V+cZ8GNXcAsF1dPND
67M4Lh3BFGSTWuJ/7m9nO68f058RKxhWxWwfVxtyKZMKEb32K8NumSQBsV1IgXXCCGDWt104Qx6T
GcjueG8LMes9HGRQiKRwjd63El/UgOxfJmlxujARnKsRwJuf7Y3305CefogPnHB2dB4S6UVi8GvX
fsg3wKzd426j4dtwvxOLAQOqdyblh5P77J36HVh6HRABcRGqbEo72iqmsINgiu6JeiKu7pJLwJa9
itgjI3rCxjewZgWhd+cHKr9X9m0ASyqfK/GjgWV2lauPq0x3iINop/AxJoC2SIhfHb5IOAZCiprK
ge1l2havD0mSVxMuqzgny5VNm7XX8rQe6yca36yujsL5R9ICFBxk7qhL3dnPYfx7QU6+sP7+PB5f
tLUVnM1SlBFCV41/whYRbnMe4BYRYIZKwcSrHWSdQ1+wtuBK8ExUt58n2bH0YzmTHS0IT+TU09lG
v7+AVu4ZdmhSghvpoCB4Lbz90ISDcW/3N9EgPM8wxSvXlxADupY9wp3i+mnu/UWs/GD3Omi7iFH6
Kpf1/n/itXMhbT8aeE7nKIlAIUt9Vw24wklVR7z+XHA5BlL4KSS8QmObf3fmtwzXLp0TEdOVkv7Y
03N+G8Hrfr/TSbO5oGm1fFvHEvS7KkMZCdC0MAryY6XfMcVH7lExOnkBZPq48KevfIzILYXSTGlo
s/2nHTyirA3BumgNKEBKw0BlycBEHc9Q33EW1DIWQY4xWVEn+lkVKBYyi51VsZuYP3ySiCNkd0sq
9w2t6g5mbAbEd9aRg6en8/oEXun8N32PbHpwQ2foyye8WgNIQaRzNF52fFU9zTlD48mpO8r4b9wm
Nx0yIdhm0UDSE2leRtWfqdQWYXJSDH2x0vEscSBw3xP3nRGS8mNL0bPTvh/VRdGc9TRMk7bZogPE
l+7dDXoYZUXnAe1dbzSNATwyth8C156pi+FViFSdjiD7roU8a+xL0XVmFKwBShid02mlB9lpelQA
OgKD2ah8JKtp8kN0J9un5VvAug2pnI3oze2rh6HQCaGusTvIbDpXuuq6NNFZXXS25ORHJJ6yZV4M
TRdQBZgSHBazyimcGq316x/V6IwjQIfNK7yGKR+QD28KAMjTpy5tRx7OITb637QmX8T60ZRUttq8
sbWGvCApZxb5oTOwAaa9tVwcyXD3xtHFRSMfVhgjLxM6j/xZMH/q6Az4VgsHRuieWzFvIS1KVhOU
mHzJPvS5Pgbgm91DUfhy7/EtrlJW/xPwO+PQ92SXj+4eYWWGUUVnzDT1KBNLduy+SNrYHz8KHlY3
4fYVT6TGBlt3hc5DDxMmHUiaZpqBsZ9/w+DvcHDIbx95CpJyHg2FQkhJlNa5VLINDLUP+rmnBHev
rQfeidIuXgeRot+Z100+HUIYLEeV487xL0mvFggpG+IOU1UuBz7XIRU82BOreJYhMXhFpKAfq1q5
ryeOsTdQ9Cq8gDkEEBd7pw1v//vZy6GNyW/g8XdzgiEzAoxvyt03pypsVHCctDDjICYthhwk+a0B
mTo+AJfzDGmHmSyba4W9mWRGoN9ri0BFQwtvGOzv7chaa77RYTiZWxz8/QX+O9RqqAlQ40dxorRB
oyU3dIyFymny+/yDcNjzE618WfeAbLK8mz7tHD+VJmp6b+4rxMiDBQQnkZmDRAj/ZntX+s7FStUH
ulpBpU2l1P3DFCYoufN/Ny3OCgYvQmMEqQvDQxi57vzL42BTan18MHjSckKcQWlywmhUe39Au3cs
SSoVv6oO17Oh67VWtROHYSARrI169ppI4BL8uudXF879vqkzDveXyXlxqUkeTjnqXi3vJDKI5rnG
DtLMBt0xW36Nx87fICqSgL5f+I2i9ADOPMkqN3/qYr8ZKuEEw95T+B8PsUbNBWTIdA6E9d3j12Dw
EBm6q0mjnz4okXUc9yQc4CCyk4a95Gy32kH9Do6jxQBt2VsorFrsD8OmPlqQAUFxy1hCjKkbXmrS
TGQD6gkDHz7whud8pkuhv49sD2b+00WLSwxsZZX3e39bA0nBPRfmET5Ysh8u5jnoLJu1bZDrNO8M
ZStQxGwQ7oETy0CrKTW15YInqD9fzxqD7Hgafehl/IPxb7HgZLSmWFGOd1tndgs3Y71+GfB/MUqF
+0872d4q3nG8HfG73PYuvIDZNPU85msS1vR2+AR+Xkop8YEJUzuLQZpq/RbTJrg6AhxH/F+kZsxT
xDWVwPVE3uC18r/h6/yZEPzFj0r5GBILydQDxWR690w2Bwt20WSIbpAga946utGvi5yegcAw45St
AGalUUIGE2DCAtDWrtarM84UTnj6Py0muyFy8JtLSKxnGQxGiMcTgTiCEk2DZpqXaWgKeRXfmU/5
D68srAqcw1A3wtUizs45C5OeDgInCCX2DkK/sjlxF9xsxbV13z+x6Vx38T7PUPOpgknwlEvus38G
xxu+Zi+gnmGONXgvbxdNfB5nrh/c41vdZFKzk//BMbC+wrtq1z0ei/dXl3xJVvQYj7yfYCqPTtF3
UbRKcEaDbHWHSEOXDujFA3p+mqcU6uQxaYwgcr/F0z4Yup8a56JeaAY5Fe7dWrrnivgZs94G7j4K
cmOlrxSYXzNxzXM5h9Oa9StW1moJvBKrYRxvFMk0yS7kgYxAZcJraa9DeQMP5bqwyqCvvnERDWZI
IZDfaqOvgsMPiTp6Pz/B4EIUJRfmlddTwQ75Ou7NyQJVYli6JFcR/e3TFoWij7TWyrssEwRf5oE/
mG6hGvmU5C75Q1OLwucrsqyqHY0Ozzmy+mrcry89seNxExmx7Z86T1l4oBM4hF6C/Fw3M1B+APyr
uCYSH0EZxBYlOd6Ujz4qqTPK+GEEhay31JefUuzob/WYh3BCecUta9hg/HmlUg3Qe0e20UnRBItr
kqQzbD5jQ4Ky0fQfPO3vzupWYFUOo6p2lu0YTx2m5tclwpk72meKCd2HVVSFGn9prErBgrhvkTh2
kxhQjP5JA8VU4NRde1aJP/rc1i2Fzyp5TambkHFxCmL6SKDWxGBe9HEFh7u9ElZy9v66SEz+rnBz
67GXIcL9QDpPR/8hdh722kzFznDTuuvMXLq2Up5KSQR6806Y5oi2AUzkEsQcmaSvDOg72kn11FlB
FayaEiya8mFpx3ccMnEYS/+m4/TiPSx/mbzq/5ExCawBsQEP0+mOvFN3gYUCyFm4Bbhp7spC1I/D
nhpLs0VDM4fpRIYQ9d0X409+OP1mubnZ5GD8w4+CEJXvBuY0SgIgJUwM1MlX4zX6lk8svZ+OMjai
tI4U7eQp0pC+NKcdY1EJROrT0etP5VjhW7nAuXJ0PvgyLxQcCvbsDh4czFrC61VSYN6zcobn/bVs
k6MxfUfFVg/m+m/a2fBJ6ZITwOWcydk2Z+J73D2jZFa+6w99qKVF8OOo6O+U3YGCGDh/tGubN6qm
2AZRVtTQskGghtzGW39fzjlfO0hVcuFMUSQ/pdgAd8iQIyMpJf+ngWOchoQhi+3cB0c6v0JrEKjj
UNIjArHTEEPN1fr3ePGTkR32psN2IdJ1bm5EZ7Tif6yVxbXOLAvQsAWB35lv6oUSYHTOHPYbT0JC
GOi6BMpiyURxCA5Gm07+8yRMJsizLNGQ/HKAjZjMxKrKFaxyu8gwcI++KnLortcC7JIhWYNrvh2m
62Oi1HwQSd/3nz6z01xoGc4StrCq4fDBh+3+3+Q5GtIGCukCdlsuRu8b6neKh0nqtA6Pqcf7Mio2
UjFBkQfJaIImKVaqlti18ryuMI9x/N/uMi6E15owq0TPVeGuQWfePA8Ar6ye6d2K0SSUrOZhrf+1
nE5JBzitMyz/mglb3l6tWUBkBsdop3fA7/k6DR0y9Q+mp75wqttxjyQQD91C8ijAWUpblc5Klwbq
8Yae+7Sezem2PdSeA60BPfTdALzjaIBgBUAeEuTHb/IbPDO42Xoxp84f8kN34Eik5xLlAC3lMzVt
gtwyVVTpbrgp3JNi6E7DmF9T+pW0O32bp/e4XfejeizuhuTH3c78ya9ZiG4reF35UvVeKF43hbqT
J/IUxgzLH241lZlUllbsEprZ87D7eAg1eLXt8fymYDfKLG5jQtXVTei+ZGe9c9reG50vCjgrqcY8
DDeSnKTpnHzS0EyppZjOqkH0NhQDeD4mtA4zLqQPhrDSwb6sTqT0cCEZbqZoPvOhDuvJADFRmv5S
jo7mCMoFsLlQUwAXF+NtAaXt2dfcpVkb4ymETsLclE4pmyNkwvS26Y9l3FGnMlxRGjpjcX85cVhI
R+iNb5fq7utvhonLmX/eReQuCjLl1pSkKuY9qrHB/9UAgfhIuUpy0jQ2YDJlyPi7DewAX+kXtYdF
o3aZ2Uy51wJuRv8iD7mZyWjilo4TB2q8OnEkBgK7o0O/J0kyLGLlxaA6XpvP6Mmy/B3TXxUYdmB5
RvHBtQxrMsTIZ84vqYbMj00KfN6xJESbO8gLDfdzH+j+JwqBRCAtrxZJcHl1MCcg9HoB7EZYoTBU
EyW/+6XD9pE0FYqzEMdvIJnvsLsMsxGDfXjFbTy6iFc0EzU3uqiicLIj12fw7wfua8++m2yfvZbW
HTHxg5K8plPz31lIICwKY4Qg+zwP37MBOggaL+JixdZbr6dGw3e6OsUfzpXNsIOX8GED/tLF5CBB
4sNz2kYdVbnaINZCRjyA3CF3oowqTypkZ4ThWt6mMnfK/hmyAbVZ6TGF/ku8dIyOE+1U+6gS69vY
PSYir5/1n1eVeDHs0cu73uKluYvKZD+smyfkP1ghyd7c0NSjG3cqllB+WIPqITUnhlw157xqwIZY
BGRjHI5UaJrAEHbPPya3ymKRF8zVzM/8RB4E+8LqwOtxsHSNAuA8OkZ0zAxNYw1uRNpp6AEpXtMS
646npCpdcC/H3DW0PgrKtrRFdBwbtG85/DMT3KJFD5q3sQ9T0bzFlN8ypvV6OkoKNoKTAjC7nHsk
sFAz/QzYky+fXW/A3qP9pudQ1jw0obKfgyJfmkKyEfQrkPyIhQvDRj/24UqCL3Vg6zUlHggUo1jD
JBtISZGxZ7ZEJbdM4aR0C/mfGXulsBnMgUaey+U7+eV2h2Ba9J7hfpOKhOOcK52ZEW8R0kbt6e2Q
lpXz1bXBsMDoVE5nIDkjt/leHkjxnUxD0zcQug09fmGGyHjdHLh8/19AW1gCNTK7If4ssaxIS4ko
rKu5AgFzRjU2zSF6U4o0rHCYqrIw75FQysM6hGA3Zc+PyBnrV2YPBfLD9JuJOxK7koSRclMG1dse
SJ4whI7Pkh/g/T86DOLLnmE0J8zI2fjvehQw+xOvE8TSSWIzlVLAhRTuurErkp4c7Nwh315saI0Z
y0neCBCKnhTh5rGpxM2hoIcz729r7jhnjm9xl69qC6TGOZVj0SkHUpp6ToDNWCbmGSIhCOltcDB4
vblq3dft1gWc4A1ZacMuqMKknt3vig3VuxtKQqQxcmy2lKpmng/a0uF2sM2xj5BSXjXEe13hGcYy
aZGHCyZ1kT86dnOAKFtxkFhyWYwQfqbMuH0f6s6Su/BokPK+GOAScXxSQ8/g8AUrtyOJLbTyXN42
nbp2WkKIsoePcoXgGT04zjMillx2QkWq8gLOnECON9CUOkccZnJ4Yqq0wSiWxX9xGme5uz8jC1XC
imvJ1ewugu+ApqUGXpG20uglVCmGrtMroQO1eQmKcKAUBrdN/e0VqvhomiTaIkhqf228er3G5bIa
ni1bRA5V3PU64ikm7gonzvvzJ0KHWEIr+r//ugcR8UJMgnA+8VUXDEw501vLbCGedD5XHtbpHH+t
jlh1qd6Bep8pS0LNq2SkudwU3Byng016gXqV+PywCWoMXM3Q8zCF7IuCB9MLYVdJoIsw3Q157+5x
blWfsIBBCzpcnPGzENOr5nyu73QI56Bgw/a9yFL534DdAjzHSkam6ijo9TyCqQ2A6h/iD3EfV9Nz
rUWVWK/0L5p+uvL5GvaFmP8L7zh15lLG/wd3b0s2lCyF84I/Z6n7tMpADRtI8nm3EwtuyQVQTmyt
FX0D6DsRjbEIx8g2TToB2n/AUX2IMHaDmes3kM61z4w0PpjjpRRuMa6dbxK1JrK923OXfnnhUKSb
+EcaeDtRS+3+/RhUrQjp+8g0Yd4DBXGiZE3LWYYQ8WXoOyNxxhbI9D1o6bVBprXjqnOeTPQ4kzKJ
kMJSCLKDtwi7ckZIpYv079l94wkJpJJjNsdaq4woHfw6XNmJ6j5ViCF3CBu+r5N3OaUG4V65GE6o
GFZo2LGgLnp2nLhQoZwQSNbARUuvkzcSZZF8lEvUij+T8HjcY9byGGUvJk7FzCL0x7YRHiQgKUfM
Rm4YDT04F1cdhzjDcy2nkjPYg3AuKsYiY7Cv4tA312+VgzLRDVg/T4aCSdI9t2fJN78pq5cPc7zj
k8VCbF6OpoLQSCqj4wDE6BFXKFIGtBCUokP/MncmkahlykthkuWemlHnKVP4HS6HYTM/uzUviQkU
EWX8/jhYAhwWwM5EMoR+Qyl9hQj1ypJwfS6MYrnjFnEg4SOGYk8SjAPqhzTT6TJ6pIFU1hYZ4f0p
0K0MSXxrIZlzyBa14Dbg3B1A2bo0jOIpM1+qtt1/i1d8vs2g7wWe0jlZk31J4TzDHd7WyFs9o5he
3lC7uhdimn9dO1OeyHLtWicbOkzmwA2nG++usp7Xpcj9pgzB31iqhmbOX591cgRjpcSEwAg3Uz2x
6KAPJ3Z3jzPhM7Zq8bS4aRID3MVinMS9AsoXmcTHdYh+V5iZ7mbInGliNJ380/pH4XUpyu76ApAH
d7t62Y43DUJLhKvIrHWMO5+Roa6INsNT44uj5Uoc92gI/uaZmzv0mcj2JlbxC194Wo+qU5vaxNkq
Las8No/Pi6YVWVWtU0BDPDO/e1z4QHTW4FLoEJxa2QkZM1hMbB337oQtKQzrooUJ9sXZewkT1B/C
uxIQMNBAB0PdsCNEtqq+TPMwFtl+r237BtgWG228fFjlaf6SMrzD3uwgvflRZ9LEs7u1GRM5GWBF
GPug3vPV74YOds+EkikniGHln/PAMVoPHRZPpNbGGo5H/8k/SNCcKgghi2A5ZFnqLiX9QrtC+FU0
asWXaHHs6sUh3VS4veaqdXhb9iXIkSo42hgrVQn9CM2RTZbq/Vo7YY20HSq7Tf8wHGZGc8tAsa5Q
IhnxEDDLWtKnzOwarf+2wqtdZvyaaN9ka2z+9Tg685mBDXBRu8ffdYncx1nEx35N6TklxumtNKET
NIll7uYqliCddRSDaSGA6vusaX7Sx061D5YUL9+tzv3DhFN+Fg5st9ktehgPaWauo/sWMwSP+fbF
2jR7RJI3G5ZS4iVRUTN+UWNa5j/nljI9M9NcVGxOGRsQgvMAIjkApF/Sz7cslRrbfWpqFVMa2uM7
4D5d5e5Fz6kuyeoC2ASiKBWiDuFPkKPdei8EUdgVHS43Zg8zCZ1uNd/HHNuavXwlynKb6e58KmWe
ChcW9SjMtDh1lVLxCJKgm9ZGelfiE8luyxRxlzlVdGFtGkTMkiJWAIip1xINc7hXdVyfdzUkp1fp
mcMFn0x8et0jrNP+KTlQ10U4V/RoJ/6+xKX12OprXEekm7Cr7PeDGp6OJZc0H+TMP598QcEfon7t
VycKcH14RpnieyytO/XouPgVbnEQZr31oSJElQPutvn3xWkeUOr4jnmntu4St0eRMwnhkgMWoxIE
7uNKIYa2mOU3d2lkhh0MMPHxyCqM7fI+Ug9JC/Aq9I5NxlXaF8Kynsa0KygdifUDWSQcXe0aGkRz
B/dO9DMgmU8EakVmWcotMmPAAE6M6VylrfHFQF75Nd+3JuEztsCMQaAvtLt/QZYARkQLHKNCSFMI
uk4pcbHzm8mfyrXAQwwY+U+5JlY2jbKmlq8TL7sDSw28bI+3/gVtlmqRpQfZuX8ijeUm3JNvvw2D
2F/LnNypgEAtPOXwXoernuDYzJ8ZhIn0TZDGmH6mTVwNswbhIeEB6B4mzHIpCEbhSYccWMmbiypv
aHQuGTt8cb7JCqXHRAIl+jlShvvnI+9i8p4ie9rVMrSdqX+MxiPf6Kvh2dukiCXpaS9lzf3+qf/S
wFj7huW/byxKKEMwXAEj2MXTDQscDuMfSDKmKDIIITbBkI4LbnRttSd2NK1czNqAtiu9Mw+bE4r5
kIlhgFn30IxenZaqsEz8pHmFMbSbvRHAOuUTt9P7h8J5IIML3N7fJo5/7pmbGV2pM3rsEkgehZsH
AnHmz0YkhGZ4AEKRKSc02lQBVn/UZm+EcXb7gXwHmHsPQEd4FD51VhjptvQFxEq5zKHLD+I5IO5i
H12uZrC2UdFfNurtnj5bSs1o9yzEpJqI9EjnhVTxkXIMN26go6Lcyd0ZPvXq1/dve6M9GKVVAAJp
DXHU1CzHGhzbWhivKq/e/HEhoDyWEdjJTY+9Bu7OSik7++CBGxqw85/5xGpdnq9qO/f1jNGrZM4q
piCeTIAshQeU7MQ1anGnmor7der6mCOhC2XYFnO26uuRhdUA9PsL3scxErxK4Nyp4J9KNmGULCNX
aMUFRREDl7wwc4yL/3dGpCfOQKsKfHEL1VB+7E3AvZC4BGTXm9ghVa+bOq02ygKeM2kMuRYqZvnK
NaTD/T58kjFfxvnNZUuCfiudiTT3yvAFh4eUsktDMCodCDsZoWXfa16H2RcIXz8+MpmbkTMp5VNX
jcpZ9d4OfkTR10vXPLxRfeo8UDXRrQW48Gf0wtrNGwpgngP5z5mx9HVZKwwah/oIog6jhwJtdgtB
tIUxVPKcp8uBcaXEzyVVuqdDnLDZdoVlwI+wVNdfV6VC1jqpKLeb6b0UA7+DnGTXD/U6ToXlf9qw
hOUzY2bHNEvqR6+99yXeBJfgGb/NrnXP8H/naK1tjpCu4TRPuB+/HEGDiS8b2CWKINwEWwt3AYG9
DAx4gJfNhXCFE1ZzcW9F9cfOgl4b6PqJu3UJvAsmiZobRnWb51WPNwF4UTEJ3lNGV3lcimCsIP4j
tMsYwpxaAivDAqZSPuMrCRp1fKld7gvOfHG4Nc9KnrQUqngjUCmyyAl6yT46dxNaCZYNhpWVD5TV
82bbsiLTk3FAUdZ7YeHPm9y3u1aZ6QiLaSgTvR7o697rXr+h580RcSbIpBeNUXr6jccP3YLl4Cjf
M3gDHUHwj8F9ZSAfXhg1sAPk65KZB8mCZC0tbLiyLQgaxQir52wm5I6o/NzAwAxDFLZfx+SzgvA6
dHIE0nZ63GKM9JSB9qAM9ktA0fvnCia3WCRbiKMr3AywmGVXgvHirxMAg5MvAxvMws5i6Lw8fXgm
FUEtnWZOpVKSeB5eK6uA+q/YRWaDh+A1dkwCfxiKw/UZLz0UjvotRMzPiN3tK1bYopQgAKYscyeY
tZfcsNyeZ/n3faqU4BrHw2uWoaqlTZQQivyRJ8ivnGT86mI91wJAgt/IAqwAlcetW7ZHZzbtWUY8
BlLVxPkmUXKWvuZvtopCe9wZPqGv7QS3ncwdHD6BjeMEti536VsyOL/5zJLz9e/ucU84IRcMwNZF
L/KB9uUii9jnFoHZPDkAk8J5dU9CIn0v/9IqRMEV+OKwSnpdFlYEna/L4+e2vLNpVV0peoNVY32r
+yBgx761RqCN6tCBe9E2cGM2BzvQ9IeyVN323javv9i1frOX4MelDhE9hix2ld9Odsh8g5fjE/sG
r9a2/GpCI0rZvHhI96sRrA9wUF3dGWVW46vHwuHfGfZPGebV0rQsZM1ptI3IH2xV/Fagby6ps11E
G7K0X7qCK68X2Wu/8inKQf94BNgIdHJ6g7Z2iM0RDvd2SoQgN9iRtZWO7k28lQkoSMje9XBc5LP2
Fl0BDw84zZGjYe1MxobMB3mcbxeKLr/17ZrcasYzi/dfS/6uJ6CGGBiczHIhUQuY+tU1REED5G75
qFpJ5atg9RDnTszNmw938cENjK+k9U1KJliLjXTmA3+pi+F7IB3xTfx74MVj42FZ7QMoC49rsqUr
eaoaJjxKlqz++RQ7xSqHOtImmCVtRtfTjtWB4lmdVjlOSHAzvkhoWI8yw7M64axqL1oWh04CRQtp
vvQ4vcBRtOFTNILzqkoMDZa7CO6n9uvx97T+VfkoIfK2t+UFOXwtVSVQp0p0TOlWTZvraGZVtb2l
fBxX7bFIC5XQV4nIFTtubEPKnGKc6jVTnXiDMuuPIOaGjkbdGvIJmW+3rAK/eaUd90R4x9Z2ZdnP
QaMTkZQp2Mc8netLs3qfaenV9eK2xmrH7fvVomlzjUw3PaCeskSZeMvebuacTA480zn48LTWabTs
3IfaEoU4l2CyMzGsXty6VJowMHjoEKRTX1remhYeRnaaHCoWd2kF4RQJrRtVx2/EG/A5HPA3hVHs
ykeWPxFChfgszbl8ghY0sm6cLK/AQWZTSb6GjByEuB16N88DZIYNVqr60+vrpx7ixqGIW4aTgQSS
npuU7xqYyBf4o7ZPO3m8IrFT+yvi29Tq4w+FX9l6VY1LRngWz6idFCS0HMMkBtyFOgoKG2zHBl6/
LGmPsV5JooVdSwqnjjsmo3kdv4r/F9Iy0XMtJWNOfEZ1cQCD9vyLpP1mtdp+73cEaacfU72PlDer
ewGda3npktBNyFyd5+Sqnoh+Lqf84F5SYiTb0NrjFE/DuAjp9vmI4wwpVsNoRdit9q1ijM8QomMr
UoDTJz8gbxNFCz6c4sVIHsfs42jEjdERYpimHG4lrlqGM0CL40Gm6dyMAreXnbSYgW4q0dwINJ1V
aqIXebVo5XToqMBTg5qrue/9SCkRz9M+6/sZr3VA97HucUDv7Uarqpd8R+atnvEe3/Dk20F6BKkJ
5LiMcNYcTPWokwZHlP9cjQR98UyRxr/kSoqBDshvw6JEPmAbKYxTWx9o7ZxO/o9MnyiXug2jrn9Y
Jnh1lCSO9UeNeYv42NlRmVyHeTw2IcHQX6LLAnw2Ni/4LhMhsW++S1G+J8lYscJx/UI8DZ516Xe6
ytFIgSqFFvB3wu378R+rjO7LEJuXaKdQq7wsJrvRAJGb+lRK6dT6JeDPMnz0IhWrIReBypHG7Y46
XZwYMVfx71QuhKOUJdygsENuweULPtBZY75Ik3pUYIatWHAS4pJ1gpGeKodGDJSpTfPWWs3BOiD+
EN51WePjG06DwJdocyCDNFVZBIQNH/YEnvJDMQ79RChGUfhRkp14eERfqHLJG0RgNDtpHDK+LaIl
FsdFEBmu7o2FdfVap3YyLZ0H0P7vwseLbJG2fEiFf7nPW2xEwSJOsXhtNR3wASBKInFzzegaVwlj
p0QF9F3fwAAHi5tA1osN9O704nOmn1q3kI1I+HNeo6FC9KYZ0b3nigkc4CMMafJ93536l7Q7C9Zu
J8gqoxh5Grp0tVasrYuj/u7VXTcI5/7KfgZwVwts50OrGbCspHwxnQDx7EI5/tUHtxh9eA1vmTrN
gx01wDIZ/3hRtF0y70YPuwMwqx9jHrBSbAjTwQw8Ksgx6leqMA57Fmx8xlG6Ixi6fNk5wXTSI/Hc
dTDAPFH0L8S6nFz9d/gTtgfrKPziJoH7d1xP/DBUCcOUKU3I3XsPgm7UFGp9GSEhT9sPFsMsOArG
iqPv7TG3gNkNqaONQnEz38p2T1ESI6tm0NQK8ABLswsd468hRM3dmrwHB/MAyepKcNIamY+wSh5H
XjUpZyx1LOnLKUgNGHm8aNg9GdargqK/PFDVS3K4MJwH0NxhkFMVYSw1lNuN5mvF1vVNN+uM/osI
v4UuUHHj/CnCTNn5hQN+FW5f3el0LH3ukeaRGZ8KsYEwWvrwv5YVDEyrOGfZ0dW66EMwnE1E5jqc
HtQPrlzs6hk72nUZHFe6MfhFjRX0RlTLe1bpl7Ml4e2PhoVNMvAr19TYGcLmT4S0quj3Ry3fqtnD
sMmu5D1vF0xPnPPvLBgwbShZeqQ+ZkysBpBeBoxhyOkucJpfktLHZKw9NZjfTqlXISpzAVwnpN5X
4pIjABI/HmogMe3tOjxmN/XAN6irQlWInokhD0ggXebD16dOPlXu14Z3ZW8a7bukHiUOv1idtdq/
8SuG7fJFLXnbZBws4zwIkpYRai4w9U/s3VrxZIkKyz9SNMxedVZW3+BTN/HpsHaD+FOYqEw1rnUd
vwbduTU6jDCbeiwX445Q80eikmEwb97zX3Bw0sgtnERhqbIVV3n/aHBcy50BKq8pv49yYJYgRZ/W
CUyHF8Y/CLoFqGwDL0QwVVi6LHr3wEljZhwuW7Pw2W00ymlfSUIznk6FJtT+aN2aifLFG1iCnDJ+
Ndeidt7WlqswngJ7AdjBz3p3PTZaPRzNtPkr+66zrtIWNEB8nFQeaZw+sBXhoZUQKz81uWUfOS/Y
NQKqEbyo8HwldjbEUF8Pj3W62skFps0AA8e4xLlCuykHKj1cW4BoXPaeaX/CfejC5LxHmk5+V/gn
7yavib8mLvP/52AjzeGTSjzOfJ/o3T7FXbkM6hfdwbXQ/JvGZ0tZ6FrjTEQRs9stQruBahqiWzhP
XORbHlpOZPK/LQaTGt8zWnbmieCheCneTbP3gD9gOeOM5mQMVoBFbvBEz/5WXHmbbLwm+lKdgGlt
GbsWU3mb5MYtIcHMfoAIKN40Ff/Pq1JShB5uu2IVf7gALNFhBycOhHIG/CcGC0a0Q7PvydYDqCSx
Q+HBkA/qhCpL+gv693srktJhLKl4gpluEdglNZogXNw61aGF8D7vqv8UWpH/Y/6dnzuRIrSf+3XP
dLw1xiDbde3uuX6vzuUvLyOYuDTNA0CiUPPD+bl/YEX5xU8kSRzuBnUVLA4Pmosw1PEYbSQm2nSq
ac7L0CKi0pwKK/BZeAIPWDcWqtsO7GgDenFz7GIzHQhObjjwvyk5asLoHMtlj7flFbVvtp2uKuuy
cDpAMAZyb6N0ov5tvmDRz+AL0dj3VBxqYdxrxRURWa/2fnlSFXRwNKPb9fkD/H/aIeefb17XUELZ
KrZUbHKngcPXehSFOIh6MslUysObCwiPFTP5OD7epxGBxNxiHpgi0O6Z+hmoFdhOr2CfHzd5hK9L
fHDyxoxZNKOiWdGneLpwN4B4bR/+2RxO9BChP9L9MpJ/KhEE0rW+q2osAPftp6v2NvRDbgsl+FDz
/GR9rN60NNbTVNrhHKn9TTWbNuYSLCKZa5aXIN0DBLQ0AULX6zwdY1S8z5rSNRKF6igyZTIkb6qF
w/ECQgGZtm9nR/WPxfc3Lw1oDMgVVn3StOfTZyXxPM3xQqJYP6JzgWrgpg+nnDEDrusx8ViiuHN2
QVdlWWMNqJ3B/hpnlZHSGiv8VIpJgEq+q39Xq5fAZNwbFHULcIR4rEjUJbtx8Rs8AWiL5ycDJ868
TMBGqFVlj73Ah7JdH4J/DKw74y6yGEx3zRii1nF/H0SVmSef5DRAs0K3/jcIkh2cib3FNJEFW3O/
kRMFSuXAneRd7SSSiktO5jAbSmgfbXHqZcG3cThF88fHA1wCsLjLhiWN/6Qj86pYM7vDmWP0X3Sf
6XbJm2c0Vtn6zSir2cHkF67sp0f7ie0DfVTBZjxvpLmla2xPIK0VKOFgdJURPkFCwOa8MourtvYe
96o7tPIUxsdyZbvBiOBbxeOBPR5c8P3GV1eKrleKeXmMVxjBRiC5uN1p+MLzNONGd5SHO7/p4HFS
OXn7fkym2DFZuCEhQ89Bf6dyklxIPPdeIzuUK1UmMrGLcKKu7NnVxCSmduU4vpa/bUwUj5tZo6jP
EpCgwRPqUGy2pjTS9H5SBuFdWHpvbzj4JPAcANf1+wq+55IQIoaDAaWNrmtIpmW5UIxRqobEEm2X
3RRRKHBOkBL7QUnDWuy4Gjby0uIff0p/TZinIT07Sge01yTr0nCAe1OubBEYJASEQizNszIG/7JF
4jYgzVO84ISWHunTLS/pr7MvHPXu3GKS4kAJ1WXl8ljtfruVWNQ13VJEXXq8/r+Ii61ciLIpTeVN
l4F4TMYXqyONxuwmYUA9MYmqi2d2Cs/cP67qa9N4bM5bnnMwju0ow4UxvRxP/vP9n1CH4BFN5/LE
Q3vAZtAkLAhKI+hq8AH2cLRWYgAJEXU0OH9wwRdbYX6hzEqqN+sAgrMFg5JGvZeaLQqqC8+xA2oW
USa7HMj7EvTy55baAO/0kYGvaRr+kliBD+rEEXYC3nRnRta0vD0f6PbhQ2Ncv0e4JZGcG/IisqW6
m9wiwqny9dUbOVXnhJKzn0fzGBq41N5YDDQYMDiHLBA2FZyDoCVbCJ9VBHNsyo4yaX/SGeHr02Wf
NV0mJ2mYnCtvL/CN2t/17avSa3Vrrukr4n6+9z6xNQJFqVxN4lJFHEc4Pk7HTnk7jZ8igBNupyxx
MFeAA6kCXtCDE/eprKqK3R2joTv7/JE9Y94lurbvpwtKzbHxDqKVXg80Poewb6P8wgo678+TlMOl
NRfpumr7B+XK1bvKqAvgYohpDN9fqBxO6/u3/XgX8gu5ZAPpqZkJosoPpCjs3rjvVDRw2IQ9CR0c
l0qPBb3GTius3uUdj8jpVULJXTrnIAAnTg2tIO61lWm8nyjxgxK0jYBk7FfN4/bDzJvxa0O3A/qS
qqkI7n6ELyP/GJd+/Rr0i2z3VZs8Ccc22RK2h8GNS0peGs9KjrY4eD4DWGHO2f5OUjOCPeCj5QRP
NtOYSx4/oZ6lj9r2DIy+qoiCcugcISoMytNzcVzEsOr1iiuIXDJMYUCBm6P3Pl0zSspDnBkU4hVG
1xIPC1tNWeqrWOriXNx1f7m/k880OMtcsKIjHIk3gJITaJSc0BgOTcKXieqUFsxj+o7ZQqBQrKh3
2rzwerGApSFSD0TF6j/OH8IXGjb81BgD/C+uBU+ZG01IeL+aPAIl/Fp9Q26yq93XwUr8ZH59pXNu
Y56NwIavFOZlxQDC6TXZUIG7soswZJZhxXgz2PcLxMYLH0nLF3lCY+7WIKbUB8sENy66+pfXMOgJ
XqRr+EOQOe2Ao9s9/G3yDfqAvytesEbDcuhVEk9vzHMbqfJ2IFb0UDQaQpigUNCGcklNvf60xg3x
penck6uDTLNGf5mgI6zeSzoeeOJY0wvnZfnZsnfMXXLQXjm3KkRT71odogfrdieIKVWh5NORNz4J
onfsPOXeeZdO9BhGj185QNheHJ72dH/jP8Qb4LCXv1NDhSdAIRqA7Uc/irJJsg0ig1+Cp/7dg3oy
4kVajLvPTD4bhB7Q3H+RUVN9tOykYqsap1ZqfCLZqj3wTFvIzJs0ZbEMbvQFjJL62RKOJvRcWeqa
LzdM5GutqWBg/kVrJ5OpXkMeI0AOCayL1hnPCLLq2ErrHL7RD9qBtPlts0l+lj/bt4hbLwa7GGa5
AtIWgftyF8zY/+ysvdoH+7ch1JCqaxijaN0pPn3PiAY8qJnUihpbF2KRAnZXObStUQOcVCQ0TY/H
pxRl7ru68A28qRX+LwoowyniP3yEz9lJttPjHdEyT7bJQAZNLCdtKxEFRh3wRkZds/qK80OdmwLm
NMAEIHQjJD9kEjGP5Em9h2amymvHRIOMdqfSttqdZp8mKKrUQMNnvq8AR/EyNfaqz6kP6zwXqPQe
4XwlRyRRbl9wlaGak37Djzekn0ErBj9GDpMy+1aYhyR4LSh4oHDrmJ12R1rIt8qWgUNC7/yxu+K6
BRCo+niUqgc4QHvcPV0TQHXHNgkkoNQSp52maGicy6A4gFXPt8rtcXy2P8ECa/V0nH+fLcnk8Uma
Yzvyowvc6ShAx0p2LZnu7C3iU58aM7sfTSMPvXnIUCKstLlDKMtTig0Y9gSjmgdWaTU5bHN/daHq
j1DR7tWqcOFiakZzBZTFpHIJh8yuG3DWBLtkMdIk07605UC5USVnWSVOfouBOyPfDEQ7PcAX8ozy
OAUFxfqRhxRSFf/1cDign1+IBeyklP+TQ0qmQacM3LWs6Gv7NMkl4DDrCG4/HrdQzR+B5LOjaR17
sXom5dXvgKyQJWLnl4KgcZ5pmnR3MxuoafxkABUHzSuZkI+qDaChbal0EZUk1HdeKEdudjCBIV/a
kkE8FtJ4h4WfHp66WGBKpPK8U313uqaTrnSVH3Ta1qrDMxPNOqH7Ijk0ewg3kvVk8AxNprexE3Xk
NgZOmCuonVRl8mQgWUoj+qU6CFyQ206e2o6+LZyiFmEaS/QJ7cqYDSLOt9zqTnasCErgvhk0jxk8
XL+cPp/rc93S8JM/jXx4ALnh8jkxA9VLaHTyQ3gCkIWkD6VLe+Xklineck3NpUxOblpcxKJ9Q0ph
0gDz67PSowg4BU8eiF7zsyHd2+9TdBZqvGu1Q7HhAlM7MO3qAZuht+6nCPLlismavw8mskV/XBvl
62KMhGs0RcHZ/eVIjny33EhQ2m5XV7q9aAMXjGmWsytGuaonCqE3cFcXPQb2MY8EH3+fZoPu0zq7
OVNDUm6QZUjllsnlvKHZfIYJtzrpVpnUuKYZVObmQcalODI0V35easTfmheXv050Mf4FAhHNo3oC
BPFuPhn1A0IisEKBqp0YokafkPLFNN92ewH2ir/8PnckrB0tjsdNlRpFycUW9T1A0BvI0HAcnqns
s/Df0w22RmiZ01w2T6n9uxkC2mJHtzZdEXt9iCLKA1sE5vvxPojpydwK7XtPzXLLEmd8KRjMJQvT
CIUA+DwfcFhJyU4KnRKkxexuLGxDCXYjFq9k+EDI1Lw8RxqwrovTsCUmq/XWvJ5gRSy26vSPlUfm
dhWy0n9UiItYu+JIcdFwR2y5jG/m8opLOKqzxnC08asdj7m5xk1PnmqSqgeaaT79E8AoDN8Moaeb
1OHxErs40De61dJooesaHeerDJ5mOzUTt+TvEHdLhtf45XXlFNqMmHnCCpdlUW4xtQbyTnY4Sjtu
IZRA/4Lr+OkiCTLxKTgSKBT4elx8cX/Pdwj1AVm3+bsqLVpJH0XZ73kShdIeIE92qYNh48x/3CH6
VveZ3q23ZsXJddJ7D/VcDXk88AmeqYflMcGGi/vpymwwP65sg5vBf8diJfsp2qrK7KVzxFaDd29r
C7UieJcEIPUo/Z2cwg3j3f2Cth6sRNdTfc1ywNxWc7ECgiOnbr1FkFg9jChENxHCXgQ0GPt6IC3W
ZVETOPuj5BNr94We22hmXjaSI0Dq5HiWPb+ZDALd9eAYZS587nUV6oJvG+nufVuN2KFwjUdNvuk6
s/+fxSttF/eVbtPpwI2TO9ZC5orU7+H5j6PEIeXkezU5ZhbHX5UDEpW1EN+Ah7yxAOJF1UufRSnH
ZlmO9jF3GL/BoBS/NKaMmsC/XnTI/gtluPU3lpYnHZpA8BRSmtgAAp+V6icBQo85RS2ynmn5GAPz
ZkaKSALy6ZTQwyYcFUvVyzMu4Yf9quBgwMe5OM/37nsLMqBgP7eG9Qt2kTQCjj+dx0KmT9wLAg7Y
KDQOSIwhp9IeGRjK8RXu5twn8cmh4WIVpCbrhCgoQHOTTpogK8NzxoBWCLL24Qnee2SUpOjfDM5T
Z/m5y2xCOPfiBV2ULsGTUQcwTe1Q8QCr7kshEXkeaqUpFmzVUgxKF0S2XsuvP4glNs4q96NfnfYX
/tpJWqmL+Y3lKaXLyGPLd7FBQMVzss34Qojv4dHEkFG/aIgAPzHUMxtZhsVkJQERC22/BrNIYWqs
sa/SZboMcgBd67UbQEc8sxoS9+fv1V32pfTN/YsjpHVkFkha9OH45nQfqsTDQxCCsjpSVzQtQqDS
bDbbh3RHTXzUQYIG5WJ8OpfoQRZfOr3J3V8IElQIj9jtHO7lYUD+PO3czITCtnLMerk/4pgUGqv1
xExqMYEJ78Wg9Tnw/Ho4yf0oCKuhiaWGMkiHS91gn+buuPYic3MYSbo82eUfmBaJAokXOX8yER7K
EaMxflHP4Lv4OfCa8vHLmDu3PqxTwejKbNp2tov4hWqZftmEQmpyqTMPjgZkBKR6mP91DH9qbwi+
oRsW/ZZ99uy3V595oBSZddsK0yJYB5MwbJhlJk4CJgoP7bc2UFHGzOp3FrDfevNYY3hGvGDqoCmJ
tZCZoG+AwfTjv8ZeI3np9qrLVIvn9kJ+W/x/aUaemZ7VYFlnrfo3gobYFmgk7rQ3hIGhtRJuBUvY
+VcMVtxPDEmTiw78EZkmMsgg9T5abVPVqLnUCESn6kpbsb1bJ3fCqEV/lqAgBFJ/NNpVaaphDKMt
P3h3rdGPAOBzra4DMQduxiz8zHK3T2JnG6Dolgdn1+165bg0rlaCbnxoayI7PBTAUkn4gE4vkX4w
xvXvuBPBBybUxMw+i24UcY1UNwEAgGnCigvOBikLNrW8hm6hsa4MZmqfWD3Mf5mEaijquAWLPU8I
3SdAGvCCTP9BSAdHEYDL+71dLtJ7ya4P4ybWZKliA/XnhSGfWgNT+MicKk/4Eqzon6txFwj6+eY2
oJL4Q6WiPnC8idGosqXwNaTwBk+nxLs1M81DEqzotpwV2Y40lE1fPovFQTLgK5sJddhWbF4d1W3m
NIV29675JUHWJQNEJkaFvULmjo4NECiV2QcrJs0Ooq9GvFgOe6bZcbwbV482OL2VindJT1xjmemx
ny7usPj61bHmpD0ihJe84qPMG5AlKtdnN68uN3Ys5Jkb2dtvINkwuiKL7M8SjHWK1Co2Lo/021T9
hvFcF4tLWc4STXkaV06qQCukpAU5o6dJFOuMAm7puZsdlzNX1ARlHLUR37LMFhckHIRjPufSrpwY
3H2rUYxnK/UxcAwel+vf5lUQJpEUxZXfN7GSUPoXh8KLgQPwPwRU9Y6YfANCQHx1zTYoPzQVHFrN
Y2BBdCdl+8rlxpAOuZvdPmVX1GCGLFJzZ3MzYspHtkzqmj3zA2SIzq08fgD3YQAKovAobiWu1pqe
iWN7qWsYhgdzH60Ua4/C64TFNbDNnEoy6WPY91t6Ac7I/KtGqrkkhOh77xfh1xrASouQj+VCdpnM
weL4A8NXTg+uSM60PU3AuNC3oD9xrEE6GdB+wQd44kyuTUcV63Mpb4gVLLNzu3xINMno0tvuB++f
GFcAQwc+5/tjtToJukdsY8b1PGzDqwXb99hT1lVC1u167WNfDA2M+kQkKzNIEyP4THGIolhVTqyl
zeCCBldsOCwKGpvvG2XaeaCdokADtnHMwfUbaWQHbdyuBsQ0vz1tL48QIfL8zD7VtWPp5u4p9Bg1
sdMqtLOyQizoRqiRsq8KMclnoGiLcGKTdfXECbg5VlGdCxa2L/1GbV7DqS2zJnrSTYZ7TTLGYinK
ebrQgp0lmfwYLf40E/2vCglf1cGJXrA4t6mgPFMw/zFBRp/WLSqIJQETbDuC7o7YHyLz6ftPonCI
zji2CivM6tKmeFMGxsQPU0IlJnZw3A/7JObHXdvCLVIysGUTBh1rNVkAUumVW2Z8AJTdxGQ7VPov
/O/qTc4Aw54A39wjmkS/Z7UV+tw6GoyblxRthhYsuKQD0XYM4Sx3QcPB3arB4GurPLI2HR/gM+nN
QISy6zr7eIE9wTjlSsehl1/DqdqDTbJoHaALRzgI64AVbyhQxL1UE4smWcjmhvPcL/+2Ja/wZG8u
Y1gt6KP+8dQTWOtOztLHy3D2Hvg2Zsa+4rAFQ9dHn1W0Fp4XDpPyIP0h5hrV4I4L37l4UR3mKQWN
4oPeBEngi9eYuONr5S5LhHLryv0FHOVxxwsddCCJ39XljhzlmDQpVD7Ha6d9hv/GeFtg5+VXzCbm
MM+OQG0PGamkukVFQFDZ2SOdTxyhcuo83CEGxZ0ZLNVa2ErzFGHKGSLRGk08Kev9swog9cfmHsog
dz3MnbZ742s5ViOc9tLkrHZUZTJMwwheUdsnXvYt+ZTQbVVBaaDKf1je7J3O5ISuLmPh7rJk78k8
0Jt2oheKQEC2mlmhL6dUnh4dFiW4Fp6W8fxhQW6P1eGm2d7u12B60fO8cowCsYdijcLSOCroSRn1
lvScs548SpoiYL0yKIVLLWNn5fInlXcsaYEOCR6rsgkMJGYRUkX22enQoknzu5j/uQzxn7apu1sN
n4kb+NLSEaUi34ptr7sWTQGVjKT4ApnTUKvcTFDwtiJL/v7ADdVhBcWuHh3ybtfgawpo7ciCWhzp
IvnzwfVaaVTjYSuTiLqvhXINDFhNDh6EFnPyCkdBe0yKNywzYQ0nSmGS6yOhL4HMXG13jQ0FCgkC
MUPYnkpLynwGux6THjMJJqR+L5pLua8eJQnUBtUuvdqYkUNyy735zVyMj7i6yCLrg3DO3VAnwGue
yRpMCAiLUBWi/DBQ3+8rLGfsU4kPMVEYV0aK/cyHOAUVm3JijmTy92bjg9bhimp3AQXKjbKlXypn
RcdkYefyMY1k/alXuv/v7nsv3V65cl/uVF/6tqLDrkpP9BJsVMQaoHkwRw4uWBKKAk51yerffN8z
DYmfViz63gxv31SYMidRBHPq15Joo/XJalvX5eVhcJpC/8uhjP18Ya4sx3dIDk0NkpSink4oUZfO
0wty1zq3BOVkbeRxdGl6Hao61x54Dmrq2779gGM5pqzUwMufitodhzeRfyOqz40qxHQhQRlbZ0K7
dMs7pNKYNw7/A9Fwm1eU8N6NOS9mOJNzW8/g6RPY1bpLL9h4jvcYZRfSh/U3LkZY4u6y8dfeJKVJ
VJa3M6YUjtnKKZ3ciOx64hIzORTuXBENhTUFgQJEIhtaYR+KKW9gzqO4q+k+SDuXo4N4aHtDl4fP
B0J7xDlBnL8FHhvJaYZXp63vunYPFrCsJmaIJ6gghWC/S189IdB5hZsBgtO6Np72R9SLNcnefedt
9vSW5/Axcak0MHDrWkGdHAxo+aaub5EoRk7pfWiN1sERvaC6Qww4kbDYNC3F6RQjoduiyEwoJjj9
bc+p8czEBGsDCdlCA1siZTOSp9XVnd7jHNK5zBuvPO4RHhLW/Hw+jpbT7Ke+5Ouq9C7zAC7ECWOu
Wz0cDX/bmcPtylJ3+0VdRrbVB35UuN3FmxrlIk6Qcxb72zmShn2YvZtfsfeXXW82J7Y74Rr/zAXA
J1WtxtvUm/TgXQK/exjGgy8PDeBJxYIVCsbOV2osZKBbDrrPhprD8aIHRjuLk6s5AfyK41MtjNx9
dvosh7ZLYoWtXU65ZxJNTnREMmuH8GE13HOJMa2yFclsc4ky+lg6C/esog624qkCjSiPEF7biGFC
3i9cJJVtmSMg9TFH3Uw4kNasoOHtt3FsrXIMtMLYaZdMXANHA/JWUNXfnnJnbRdEZD1CrB59Lzk/
HsK6OJb3cQQgSSep4UqkL/g5ELPnqKtRKiruP92+WRkXHdTTUdS2RhCx/u8KC9Oq7tss0mc5Xyiz
novDm8QfqyFAhLWHsdXV/0cPkkAFVET0NmlmoE3xoavt4TV/NZEzePConcLGpHnjStyItusgv4vB
JFY9jd8u+6F+evZLL4/xFtXNXIXQiVVs761YZOjTPoFf8EwnbEEyhhKR7iD7EtYtRauYLXfvRtwP
PWxxP3yC7QxWxWeKuXUA8bw+C0GwfIfoA5+VsNsRtHZtf/oG2UODsniENn2ywXy+/p876ipOjcv/
LTXMXSknuyBxLPmL6QAcLX+CHhN+2J4so+mLomQIWyQEC/CuECQl2fhuM4p85oZyx5diiA336tC5
+35uFCa16enhCCI8nHVeB0jMcUcdnf8lfgOnle1ILWHLQS+ga5S/D7jjgCIRSaDY6KX9rWFYYQQc
Cgh3craRUYs8XfC2EGm7uqe77PBa4Byz6AZQfhQuISDfp/M5qRcJPZQeQ5H57Sr5p2tN6kmidI3C
bLxU5tAocLTXKG5Fk9xIE3qIUAVbvHnXof7BIxzsnPw1IoqkhRvXETmVuEEZa4c4VgJ7d06+fK01
yC7iMdH/ZIq2x+ni4dS5WDNWIyQwrgBwW9+ZpmCxcsmcmbWpD9V5/lUuaUTBcImDIxOtR7rgLnY5
utY4sIWzHRfDMWyw6J6WzF5KxbOzIE+W+xt/cnMT+ltvKHXbyko7izCiTAEUaWheC+ZQiLXCcA/b
mq0mTUQT6ru1vwcb1OFuVVCWplkAN0LUS7yH5WhJ2zlSlL/WV+VOTDuh3pflbodMPBtVPF8DV52/
1T4XgoU6BmOT/LYsl4FnkOkMLoLCPbYKgyK4feUvwUmvGQ76qW0nm19v0QbH1BgZz/eh0BDbE0HT
axFqVPOE76gMh0gPeso31UH1rFbwsGYVLoyHIhCZxbbRhEnnKUFiezTwr4nMndryZS/dF7n48prL
6ajGIlq8+oYfrWkP9a1MzRG/hZsOHtOsNX4IkjxYZgAESTK5jZRjOLD4Kp0LAJkN/Dyi/tefhbsI
oVKh4TVHhsUBNOzmoWCY2rO4iz3ofIhyRfvNUq92Skfm6uhcInN0oBYfCxsGwbKQZqY++lbtFJt4
/evcU5koSgF8ZhDDwcotExlB1ooLL66sqSUkPWl3QutW2NJl411XQFUpjYM89A5XeUzlyKPmx5GH
G50VXKaDgZpe+suM22cDxxr5xK2J+nSPTRNHnSBJERKAxoZpfEBYN0/l6ExrFqOV146w/VVz2KYF
+bKAXzIBbp1CId2M3sKjco5RYocmMonrtacOzQR8TV9cPNanGkA59C318NX5tGRB2uXH9ZRlHkWb
3Wb6K4dJXeo+WNPbnrjs8YRUAl8wiVqtx2FQ3ekg5CCPlrLKdTKEFXbCkPPqa3jwa1i82AA1tvLT
mUOMyxOPiaPzU0RbEJ+Yemi4nwlf+RrAm1fnlVc25eFW7gkiPXFSZmgjW8MTfjeR2qyat/BKDIIg
wPpQQXAow072YtV8TSe4SOVM05qp5HH8OXZRma7PxPjv7coa/F+4Rowg/AMXM+o/UpjhHmyJtd9N
PzP6TlCcF748NGmdwbEOcHEAexpoYidrIho5s4+N/+IuS0s8CeaYxyBnqwgoW6vrtdncGbRa0EJu
NazVU8V66yXCxeQ2i3Q+7DqgK6zp08E01PTPCZFxBzrSFYy45gwQ+Xwyle5n9B/45kbk7qBPGF3X
00VouyuYXA4c5fmyLUm6iWTqQXBgIwZRIh5Q5+EbrGINozUIJnhAu/+kMFC58xTpU0P+Jh8m8AES
CkonDj7842aFraOrPP59LvXWYkPJwoFraG6avQl+7TOMudCP2Q+xIzgidJh5h+5ovG0wvfR8jFZh
Zj+zTvJLpWCRzX68c4XS0DKvi6g7FcIQyZrQqVKOcnKb9XEnwyzej1Ks4BE0qPN2LWxeay7lC8/a
o56CTybUpmySDA46HNNU45AxVETNu5LAHpH2l2aAQa0bhouuUB+n6lm4biEGPlaqUPWMTb32d8ak
55hPAnp2itxT4fv63QxYOxhOCNZNAWyW5kfA0hRdzHD79miUQbizs/gpZ8BtQV7q0jLfyByficeJ
V7gTv7X4kQBrDFrysgKb/hwAVch1HG6PTFmsYWHJEdcobEka8LAHNCwb+7u1bIFQzgKJOS/FG2yl
OH6Tx6+cubPaGPWOtuVRlqDF2UtMPUYT2JhLV7IaiwveRJlEQQEceoJQmqRvsE5l6NFpiazE7LTH
HJI0Cy4us4FV9FjeyEdUMxm0GXqZEvXsNBWKo5IboPpJGPEk9qOLrfy91IAFcnOY7tWq+Iy4vKtN
maF40UhpXJi37v+ngsE66TKTcZigGEDtjvowa2EA0g8q0x4Gb49HkwBdRP71tp1OmuQEKbIu9fYg
dOxtHAoECqjXIlJ0bdqs4/94QTuFKTZBC0udd0De5LoVVs1//eG2gqvr6SezjL3JZBMSRThShckb
7jkn1iNudc8AJ+tU3MjwTzfltB0fqnDiSAbImcpD0R6z8+mWKrfempqslD97g6FdDvEgVf6D2FyF
d/hYRcSQj5S+qAKN5NCcCjluvV1Hw5EqIKEYIkENUG1vUDXn+lLXxOzjDHgCmovk867EM6rBZ9DQ
UAz5CZZwSIawFYAtD5GSkJ55A9HFLdsGT6EW9486gZcPX73Yh1BoTplEDXsti515V8sHQBix1Tpz
TU2jOP70oGxFz07iQzZljTO8V07OgNrIsA+MjlPTcIFnyNee8RZhmqEutIcEPwiRFbby+K7xiA2S
3f2wDDiqH+Y3g/MGooe7oQtb/aP/o1oSkD4Bt26eWv/ZDzB2WNyNqNab9EGLD6TulY5ARD3SIczE
FTpd0DSTcBgdWjdbWnmZTv0qtCLUxd/qUeBZfUrPk7uwdHbJRASs/kzLIUl2llNHpRz5/5UEI7Kj
ECncrZhtIjA/NcUR3ljjJ8zUS8fLhHYN8s7nxOJuyz2JzXzqO+bPOmBLmaL+Bw5JqSFFvOvjtZzP
jYCPzGVgNNRf1XQAH0WQnAXRKVvOU+9I2PqJFwIg6ssoxbyLAh3AoawuN5cS5VM5zPLCR2UAGGWs
gXlgdw7Kd9k7YIAAOS+OY/xpXCFZxw5dcjyPxI7xPq21F7e2ulenRhLiQtp9kn919uF8ATrNpp+F
VtD+Z1Rdlizjjcoy28Mjcgojf/39v9uWrPBWDkYX0q2u2kxUP4fWsfPusWnvaQvG964STmBraTJk
Tb2ieaieNUumuVh4U2qRY9oSaDs4gqjR+C3xPKZz7EhYrw2DDOuHxVUDeXQ/msyZb2U4RGgA5OYZ
Trr6Hr63tuIaymHlg2f7yw69+ovqvtpfTFA1XoRNUUhLZtEI/2uCMaHat0E61taX1txUh5JqT2nm
xX9hMk+5M6X5Dj5JHIKjiwcy3Wt+4e0GqyXfAJkUU538Egs5X/th6/nUk+R6vJ4gLeKQG7Dskydk
nK7NrfxTZ/pn9oRXRY1JFmm1P9LwRC3od+fLBa6q8laU4jgNipv+2WJ/62mwhonIL/EUJ6W2UNMC
kt5fTPuLcpvbqGWY8Xz4MT4/C5qMUEwlAX3bG4Lbo0u4odp8vyeAMlyZ4JpGoSPz+3tc96UX9smp
GxZ4hWM1KgWj/67tWNSgRdf8vmeHlYcOI8av8qe1Ayr8YP4NWNYGMvSWWHsFv7sceanPvTE2mjCl
RDuu/DfJPBcqsRmFDaKqhXzpyyGwtKj+w7v5ngEYyqOe8as/CF8OOtjHwYSxPL9EUsz7LKoIoTCC
fAttushoLCmYiLO8A1YT4nlxaRDdFdhszFBTxH4CNzgESQocbf+5UT4LeEXb5H3B32eqD171aYZo
rwlGDd34DamA2EjV08TN5oGlfPlG4fH12MvQVkOF4etpjpWt72PhYLEH+VM55v6Nrma0yzriS/td
khxJAw3JsxKsce9f2NuJXqOvhXUGmDVq367YHGEJTeIyNe6wtUshwt/GbR2bku3fwDGTJkxoxUfq
3X33Ak3jpDvUHsGw8RXk06fneGeocjxh8W0/j0MabchLOjSaBZr7mD+YqciU3EOTCgfycmpHdrCK
ek9LVgBCZrWB6dH7yqrlFpTOaoyFADIB2dEhui0JwHdRn4z5MmQ0rP/1SyU8jcqCX18F7yUrkFTl
fMEqnQ4bCDMYKnukxOpWwxT3VRvPWjWUOTDLGw8UMbBU9mtEpuRCIMpoBcafh+Dt96c8ydhO7bZo
iR/ijSe8Q7zSmBzsf8SCwfQBh1aUrwhYdj4gxWR+gP+u0clpzXP+T071qBb/Cm7DCAaDcWu7wk7H
FFrS+rYB04FmMDROinlt4ocJrUvfbJ25NmFiH7bQjDYJQWQEjV6N13aWmROsJrnSQDajiK/nGQy5
r7M2eDL1/BiPRHrXeXMVjH/TweXGpg1/Gl/ozTDb51reNRvUGiKDjdOywfUF0vRNgb2WZLmyTyBf
TS3NOUU0mQPRQjz2SP/m6Z7Rgi2SUmtacZIywlimkUXmvZcjUCYY3BqjpfsNgA61gtuMahaLkWvJ
76iJvqGBDT7cjPEd2Wo8xKZYztx/y89N8FnMp6zWHpX5ir/cQJVvhYzSAYYC7HLGO3kszS3dwHKo
c9+NJ7aFcYuAIp5W+GZJsqRpcpZZwNDTOBeTFHOH2f26g31O8Jz4dpHAHIC6tuN80UptQ4EzL0ur
BsDnUL9WZzocpk0sAsjwyZ0Oc8g5SakZipIBkU/GbhXQgC9VVpCGaAQSdHDoVcXvcrKw/Ttd+H1i
yJi9L5L199LWXaoCoFgbGEz2o/BZd6F5yUx9FskVivWxFYKl7tbELm71WBQmWtZMyDYomubWReJw
kCJjjt5h/KoUq3r7wllTKMJ2qVMM/QoeQkMVTYvqrCbmMl7PLZQc7JhZUmTJEPxpmIEg7kduJyCZ
WHV6w4RgjG1/WUnw4PQj7P5YQVGzPTirNmQN/jrfAWEL9bdSauNpT9S3hzbdRTrWoDX7WLb5xll8
bfugj33CotQpV+Frfn+eKKTAAnfoV3OD0wqoN+DxIhsIPVC7sprrN2OlDIO5oR23Qdb90B1JqD1b
cMPKo+BSfrULcheZ2FVCaZO6yYuVL7IxiFP4PB9YSqn+xL3yasJ/pN0QIWRzLC5s+pyva2O/y6D/
oKDw2lHHw73FzJFIDx1qPscS17VpK+wfXUAPoBXPNE7fdpsd3qMcepE3l7i30Xdej51L7m5/D74z
btzNnVNB5XJUIGSPrZipph5dFgM+D7uZ8O7zLEitAwvJZ0i1gTpV07uxH0P+7XOWQZhpYwY67U+S
8MVg+cyQ8v//iidvIu0Ogcuy2cjjqNrC+8v7o0BD4/QRaDgdZsy0oC3EEGXt663tqirfilflbo7H
sHXLzTx109rbkXCXcRe+gfJ0PVlFEnkN5sOslmpeYV2vwa110vhbnI7hhKeX/goiw2yRlf3zPpaK
IilmtDFAlYyg0zqBl/J58gOSVkN3rIS5HhoTyt7dXQoWBJB/u9X2cS8r+WaUxgHQB2UnbkN6QTsg
sXq8fKnOl7XQZ3MOGfnDm8RFq5DsSNjAbwRY256bIIOPr2Kq/DK5Y77GWkfw0RKyBbzk7YNr4/Ks
BQjj8TYxj/altX/0CQFxr2hSmUM7MeMaO6Gma+VFcnR7nszkL5S00eJm2iX5yyW5ntKP2LW6Kf/Y
VIEEUCJQ+Lo0r8xGveCo7pwKlpJGCbeJ+xt5wck4UhBNkzPGaOHfF9yK2cxqboBhthf+KM449ps/
0WdjXuTBgZi8MjJ2Uzd0HHrejTe66WKZjqucezxjwVJLrVWcUUbjmG0+zBDJMbOC5LCpzity1GcU
8hBQaTYX28BHIj+C9M2YZqh0c5xos02t7lzjRHbb75WxtbZ/8GkdXT98SJIDfSoqtiOWEShmm+We
KBoiDyEDpDE7E/0xdrY8e8ySrl88C5N5oeEjl99jWct9qHXx7xC09+6HWhIRzxby9UfrwQcYEX/3
AyR+ccDP48FvkwfJRTAYUoqjeUqWuWEEOa9WF1CPg+35c3ukQOhIdo0SY7dDEaA8reUe7LI/VNH9
WfPiLIulxwHbnLwAIkgCr9qmh5Q57KAx8WAVPgK/HtiX1GstmC6nErXD7oPr1R6N9/jkrphmRF+A
xFWeB5tTuesgYb4+JrYuMkqhgYZqgZuf5e5SYwHxA5bBza+kacrMRnlTZI0q09gWyHE5sNz73OWl
zX20DxdVrL22pCOfq2tB95fF1s2BVSwBT46hOttOZHcMMzHT1mUhP393244Om1ivXyRDnuN2t0xC
UepyzJuMszii9LejkVqyJzrTo/eo9wqMM9ajXkmUqtVJMCmAoVTJr+bRFkker2hhfpOhk6+zighB
7zckItCotBCtxu/mqT06r0zIhGCyrgDkYiJgJngrKSUF9TPGHKFMb58MrIeXQCSuq0IlUm5qzmaD
HrlqrTNIp96jEZ3uQQCl7oSjW3ub3Nj8sQ6i32VLgw8X2Rxy3mzqKRoM+9BDdW9Fzlq3hnuiCzI5
EVmb92V4IQnPXNG+eH2Hpj2AcTvskAAyEEHuSA2yXuHjclhcXucfKApnV4uM8scXqS4Jj49mcjW6
yNpQvI7wuo/ABg9Fm8lkfdQPLsH+Hk/BPCh/pXfY/gVBP6OQzrzjS9rMotMXcGdUhNlLSU5zJTu8
VrTnUHS2XdhpQ0ciCPFqBvjWtxjSxcUpP5l+fWBS14Sv/opp3WoWCuJYN7TFko+SjQmR79XZySoW
e1HT+hSW0uKZv/Oc/OXro8JO4AVoqAGU+p1JJWb+DhyC/AJDpyABjtwblQYe5nSyWTdPuFix0UlJ
9PgYLAWF+YrzT98s8aW4zNU3chkfy5mqpaIico/vfyWoYcTXCiEuIVlY75qqTcbXHU9GPuab1iiw
n61N/eNRzFEtdnLiYW/jHcHq5rbVBnEayrssaUrfsjjPHxZ5GB5AuDd6Tf3bLzMdVBX1NK8p5QQf
x7OadQ6AaHQbUjPNeDA4Yq51LACirZFrUCqjzF3adssE3RfsPD5/XBfKV4Yq/+ZGXhYmrVmZxGQA
GlRjAMlCvbRJsVq0/LFBVw0wqS2dAZTXbEVaxrGKqlELxrDuZfbyjW4DcdgGoV+JemHpRVMmgi5N
qSwvBWAgExg+WjsRWuch53QcBniJtq5+BjeedR7BPF8au+rPdAOtzMo++m2xSn5PcT+vH1Gay69t
YIICy6Kjn+GRnunuiajTyNtmMphNIecAmd81LzYyxSkS/H5j+lU9swznIXg/OWaofp9fj5xZl0Wd
jq+wLkHIGAfw/CAHob4dAXvLgjOtY9jRj5+RhiO9EF7E6hdGHMBemSiP5cGF20qBqcxomkiBPTYU
HcNZkAdnAC+uDrVwH0NDtwKDfIv2b0rvmMrgFkA1DfeTa3G1Mz0zbHZNmvb32tEky47Tf1WeR8OA
1rBWxpUZyNY/0PxXBZuP4bxU7CSdi8vPsVW6xijRzYtYlVhJML33WsbWcUVOsYpwpGSR5MSbCnv8
uSqoOctldORUpQv4Z+ONvviIXwnL5OTSNE4+DbLDsq8IXuXCX5BoBw9CcLtUWIaoDTLIhOd6Vz4t
SgUEpPILWIFe7RLIfHOjX46qJXE43Cig3PdxDzs4n+aoVt/vuREU5TF/hQqkc9iTZMeq8FxKSZEJ
DVf3D2lsw3Up5v5dlsJVSaVWvoqZ4GYaWt33v9Jbr1KPYFY6E3URrTeJMT22o7vFYWE06RrmkHge
582CrllzIc9VcdpJHyxKPIer1jLp+PveW8n4CNqQGtHGaSLowXzY4Dux6aH1Zqz5Kh8jaH3Qvh3F
xVS54hyOs//bDjji+rAIeKMex/jYpxrQ0ivg7F46YW58/2tbcam/qbNGkSXmpokvmPRjhScf02Wo
LjXrqguERalLSXxba3Qeru4198HeBQugGvmfoaZ04+R5pWBLG5csNYnV6vz9UitoRc2EnjA1j7Sm
LnD4xsFWe2KAxbJgffA05+cH/8q1pxvdpbFBIQpmTJRLol6ofK0IPj3sdN2+phiP9T9ut9XUmXj/
JDDQFP9y7saV3OwAQej9CS5I6FuJi+KKV6uL8+LLdgMDCdDfJnNda4Y1rKcBX5UTn40Boq2UPbYV
qKCPQqPs/GyXGpclp2DLBI1waPwYc+B6aOsUrFk0+A+D2pOjLV84OnFzaE8I2M1mOL/D6XJ4/aSO
ymLp/XBKHMxzHz8EQwwlNkqVBL0po+3zqVNkUY1hyBEToU7ttsXzivyhamVCakkSxQ/pKO9AweLK
9E0tDeL2euvSBj/1ys/YD2GlIPqM3K7xne5HTuz+QuSKgob+I8q6fLm5/n6gQVxKLUxMI5m5hi5f
vn4kNQbi6wHAA8k3w5LkA4ev9Km6vPlG9rp54zhX3KKAakds/77hgXeg2LUaGtm5xAMlUJBgB3us
a2ORDX2E0sMB3/2EscUg9ttjQJHxb2AxiQYME5xwJmFs11roR+WeSkJvwW42GmlMgXPw0fAtiZi7
ClgnxMf/l9RKSqB9N2h+zezP3pRTfrprEwc8alGTYgdAHLU+CLEUCeKm6VTuYCHDip7E1UKtiu7i
EFnTCQ1WQkannCn+jf2Hlq237WB8Cs1nGAAHIpeVqX22wE62OxMIRimW71pjoCwf0rGqEZwuL93x
K51TMs8ixTSaK26hXxwrWWsbyezTJrtFP3l55H61J6Ov0hRResknEmNIq5MYkNsOCSLwtSfdeJMM
CKjr+6Kh4a4cK9/MOAm1bbeqv3k34ZuC0vGwuAc/2/JnCMJ+Adcq8hbx9aztNyrgCT/JdVpfLOxh
6Mp0SDEBKaNzJDmdk0RjvLA+dXBGvsxRuzR/9jRL6l51wmzlZlxDDcBarZhJzqGP6u89c5J+VAMC
Rz60tqxM/8ch1T3zH9cyFg6W7wqr/wuGrWEhJ+DkdKxiZ/JSeBPdfeWq/xaXrNvMvM1c4/nEdl0V
g9+7oQHM6E518e6ibnx63RdPMEEF6uGYEcseKabb8BJpO8GC3LOIGt4JgY86S8yhEOgx40Zm86AS
VAdW0rIlQDiQ8E3SO6gmDPMGLeFE1klouSqOXOf9W5eA2eaIYkbt0kea7ENhggf0nX5Sg8p9hTu1
TQWh7R1+2GgGvkpzvONfrCdkoYjhRFEpTaiL3RLMtsv+YnSbXPOMPxrXimNjfROqALTECXM2/sT3
4qpIovaznrvCCegCgJ6ou5QnGbyBk0VQ6895qiXAfwaJFIx/faNkbVsDBSbyLXMY+UuJrTRWAoVj
QECDvLDVW42sZy35rMBfwr9Rt6biLxXLLIK4MuWOfIIyC3BhJ7pv9RBSRGl0Iux6cPpSXeJ9/MfQ
3hKDR3Kea+TALJGRG8gbWuPnCYOlXolnSqvTHLaAdoRY9ipIkspLPhtCXokBK9wxEAq0TDRrlr3B
d2CPfHfX8NxhNMrXPbcCUomiiH481lLMsqg/6o1TOLgO3CM/kRyf/FFTgYH4BNxfmXnG2jkRji6C
+khllNWYtDzVn1TWJwuxxWB0unF/yJ4c/+pq6uKRqzmGOGB7bdk4m+JPekAVeSj4ylJb9ri8RALI
q+1202aKZ23vw3t6FAWuxsuVhAGehuiHSiC/MD4ikzdVhMK74sXgn1ZgRvKPv4TS28B1NXs+qkMb
MRwldAFZIFGRgnacnJAbj7totIPsPewNRUl69cPQ8O8EuPGbfeU/r2xcUDr9VYqWBjvfYoMqIs2G
Go7gZHwDum2WMUN4VYeGVKeL7mQXA2RUAl9567XLiXgeRH6Tx5qTxh4ygJcGPswnFTUNV/2qf01W
Wb/iWFCGglNm9uxPp9YiOTWmmeD7Y2E9ABFhSXPPqW4Qf2DMTNPLmpVMPhatIHUVamnEu8Vm9mR4
KUOaUbPzsv1Cy6+DAiXKpEu3YargJgq3aUZjTlIi5R98758hwH1zWkFkFmvrpdcYU2/mmH0PUQmm
j4MrxiPi7CdyCGHctMCSXJ07B4tGHvH4aWubww167gBn30RgGqEe0ALLSJ4FKgUdvQ0kG3FtUqM2
cqk9qshpl3pSVVChmZsY3ceiP73euEK24ZL01FcvZ43Ypnz/WqvRqxRZFcD8Or/hxZZcXnyIvKG8
veH28PaHPDJOg5FL/I5uqlMmG06CkWiZFrID29/RdQePs/gVIHq1oSRHKTJuZlzGLZQjW5UV9Thn
ACMrBw5cUX/IaKLfrsYqsQoO0/pj8JGbGELmpQWbhzA5MnqMtkYcUp+WrnhCCWDVctS64AkBgwk3
n01VfrmlmNVawkDol0HZUndxUX51rGDoxt/6ciK0jv49/7K1+bzropKcG08xSlQ/IedqCnJDuX6D
zJAY20hjD+GBS7E1E7zkM+PY9YpvINnFGIyclJFpnUsnAVVD/O0TW/15a7cT7h7H7pCfQ90vxj4Q
YYIw0RVBU+JD2yB5FWD1V/Hpna634hN+syMyokixVrumb4R0FbypOQrQ/AnNW4OKow87EzHKLhAQ
rbtuMNTE5Il+DmR2JSTZ73qoGJPOlFKzt80L7NqSrbmg4f61LLYCHwLNuh3mQaZ5YOPvuqYCcG9l
8sYrulZXFlcT9KDMeW+7e4FjF13a+q3Sbzvw66cIV3lUeGf59Z2LVZVWtEfDYirvGA6kQKiyv7F7
GvoOVh42LdYn7+f56aMCODSweFhj3c52b5vD7nUmihsRChI7hjO7Cqkemr8pZapd85u5id9VpoJw
EILe4miqopC2lFJjb2HT1V3DLf25HHW9GKrQHMaaNSP3Tnch6BN28UGbgcRMEIeezr0uk0ou//BE
xb3ceEgd24NYTW1G0uuQ+7XPKRTMZVsiqudlUeFRnlEDB5MVDigyhg9yXZOwFfKpdhUBQhpXkMSE
v2lmx29EKNIPRkXj6bY5QOJqw9InbqFkUuNA3pS57W1lrTW2ewMGQSBds7rcDFgpA1w7d/5PPLt5
UqHHnFCJ3s0i7Nkc965dYLTmJbJ/uF0lm1zV6T96SeeDQCAvl3fc5+ES9lWBi+Gqyu1H5njceX0c
XzXUcsvXGkfR4GbANmt6dYYj+fBp1hn5KTHc6Zl00TXJhAeDdkMVd2PezTB7+pg4uR882Si3GJ2b
d9NePKvoMhtk0xHR0g9/BI/BwFziS3DPOY+Rn9p67Lk3SrtBSlSBLhW4Vd1ErOR1t5JEdVpirfxz
Xr+ujiOHK6q9tFFA2xstSIkGKQGc9FJIU8dy8neS9vog70p0kdyZsGhzPkFJ4rKEq0UQSCOvz/HM
i/YPnBQOET+3tKK7d7g0FxHpCPWVSehB4yEuizefCoe+fFNDDTm3uWrt1X2rgIDPJ40Chq27tV06
UQ9apnjzBXMogklkoweZSCRNUsNPF5cb3CGAqr1SF0G+bPee/jY/amukxR/B6NaQS5+YAZ+Tjnep
qVG2lDJwxogKV0pxYu3kAspk+v6YyAI/f5x7MnR+xQkurtsNgA5ELmjwOkrQTtFBX+x3saRcitdZ
O22211JpYxqx06eDahHd/GO/gmf5HL73CwxsfehccvPyhCEsQaNWZGFk3KJENFM8t7JNV3S/5YwD
OPHhOu3tbZB9L7/I3fs6OeBDVFBI5LO8XHUvzS1DK+urYGIu9kmX9hx72Zz6iKyGw2fncfU9XIG7
S3MgytAIbOf7PWELD1YMLMzGuhKQBRvbjBDkYwtp6EMRvQsRdkVgej+uGMxpbOwmVJ0pYs4/+EL9
/ZfdUcEnBWjyk2FChlCFp/TuGEI7TT5webJI+lbZ9M1VgH2Xg2bCZX6iP/9bU3UzMo8EBxwXYdKA
UiW9EsGenB280GNCrL8F/6KxInVo8h3dVSksy1sX3vqLFL1tsVJTztmO0TZyt3p/Z6P1j8zUEdkg
zp+uR3wBfCAg/ciHjzDk4Hej8X2oFaoAp2rJZhQASEc9Cd1PaXz97suQv3/cIOUuESlsRlIqg0jK
j+QLeB9+OvRZGIW/9pH83qcyMTalmziGMdNcLznov6ii/ZyQVS0f2S5L+Mw/0Rni/5yHcGXhqZ8R
F91sTb9TviVbwcsd0pO9fvKmCu7Yx6PFUWTjR1S7Mu2i6MGtbo+vAjsZhuNisqgf6q8l8ePZwOHJ
l4CnZI7xwo9cXsYDFP/QWd/vCEbH9mmhBf/0nOH+93btLJADw1i0/P0kYZn+Oo3AmS6lbSCS/sjZ
Z4p6ckSjbE5Cqz+b0oWQMjO7uNRA3zu51AeMVUZIn2NLTL1rTnmUkHAqjR1FVyq+xscDU/Pq+qT9
71jIuZjJNxJj47wTKqCUPeecgZqSiDnw5sFLi+KI+OoNco4zhAJWEj6QKW2N2uWEgiHX0aaOmr1f
3gOCPjmz07EicDclCz4vjYZqkzeyy1wZJ4gfEprOOH0QPu03m3aFMv5vvZ3wAso7M+SON821720Y
GCk4AnPXaqOf74T7JGYyt8wXzkW25bVXOK/QydPnxLMjJizjLa+/+7VYwFsB0Fv1BPWrJb4B3cxG
ejQn1vOpdZK91UnbD1DpImusxCku67WIPsjpkaBp1xCPr/Lb01r7lY5uGALDyyw2Xp1LTPe+ew7m
74emGFi88ajSNXEIUMXin3EoxZnUDSZkSYW8BfjGUpqqdnBpb/G1y3jxTzb1qn5k4cnFLe+u8eZS
YGUZR4GDmX2CyMR7qfNavRUwjoMqUj76+szt3rm4KKukLsISR5rC4Pz3J2lQrB9FY6UU9ALvpWUM
HDfp4F0gV2BPTKN0tkHpn8FDOS4ulVezytDV2bfaUfLqOKhlCDCI9GOpesliBslzCk0TKvUUXxwF
3Zwvyj7dehLY7qHoAFXrl9WlPsGqxODRAA/GTydX7BCCeJYUZaGDcKanp0YVPoEeif7MXAlug94S
cXkz8t5SQmvsT63fTip89bmxy/XZe7AmP2kTTq5kwAmV0YhGlT9XBLmJvn0nDFna0HP6adTsX0Y+
nUvrNITU75nymGh1Rat8LldZKZf9tKUaJea+SRwW7aqkBE8bG2aeTkcs7nHuUGB1VoYQzKffFzMV
uSweG9pS02nVvYgxenNdFaXJZw3Wr73LHixwoPmI02fHhOaPiDRJTaZ/Mnugtq3EIPqYf/zPSUT0
7MbRko77Vb+JAHpP0BQ+eCL8m9UxSe8G3AK1cbbQI1i6OdWj0nY4SRRjZsVh7zNs9ze1UF/Do6Ri
TOHGxOXhY2m5i/4TCs/b423M6MWemrwPBStV5Xd+8N/QxlwqWSNs9stYp9EdoUlVwJHS6zIM5MdC
uBWI927nv2akI1ZKRgVIN9/yooJ5XUToRXDAFVkTziOJu+5EvQrvwhV+m7WXFsieowWZzpZLCc59
65nqKPzezUGAg+M6h0BoUHlbsmPYY1R592cs1RrKl7VE4+87xvteHlQulxyjBoc7IzJgIHSIsHqB
mviOGB3hMp6DTQJpEhqeinloZP+IZIbLiv25vrYapqjQ3RhLW6/xmTW396If9yQLIzQGJ2+LK9NU
ERsM854ae+lVO9+e+46bzBYM4bdvbyuMzpVw+7s3th5qRkoT56vOnScvEC9NWiyCk3PyelWxMqOK
oM9dcGOLHrYFwhVKLGWfo0VrmOJqP41AOLiBKXhu7X3wlv98OMjou3eoTg9GIHQYk9nLACg4Pegy
+asKOaRqVsJODh3IXpZrm6L7pcqaiVbmZw00Aa72T0jolEbplJIvuHvpO2XlMnavIdv6po/Ka1Qd
Bslefiv22/mJGKGYJxeD3xAv0SkkcEoRbw2VNv6wHTBNuK2NllosfFxkk1V+kvqK42BA8SSFxUXK
Do/XK0Js7NFRkaEmgzDfwAae30aRs8X3J+fGZ4bb/pz0+KWnSEFDIFFjw1iaOaL+pdo1DBtBv1hP
LveRw9BCFAZ1XPKZFhQWsKSvWeTCIash2k7a94y8p8/+iRoL8CBoXPZBQPQ49z3Ow7cYlmcNubRI
yLaQl5ArCcKrUZlMfzBzqSCcrp2JptP6xyXssksHIHLlcAqG+ZFuvwWsQv0pcqoQ3tZfkAcPzdLv
fCfSJR4oJazksPzDusI2NyytlEiF6dffgygF5ObCcVE+pqGgvDSnZAFLqdiCebgwqyiyM0zYmlQY
XZy61dk/19tRUBM+NknTxGNn09pImilkSv1dQFFQMRnM6XbndJJN1h/ZHmZfEAQhVwr+HHkEloeV
o1ixYvPGof/7cEiz/HG4UVOlPOjQfvxQGY+XUCa8duJpOhG2sJFLdCkZmvI3Vbq/teZYxtkzTzM3
tlh4YRKw2qwd38HZYjzf2Ll2hfAkZ2YaehhqzfoJQ7t++QdwwKENQfmdJ8G48yZ/oqcOzhBWOpJ2
SFiTX5abdAtkd/RALemcPXmKYzc9lnv0jxWz82f6FMoDDnrKVKYPXlwsNco0xxpgaZenEetD+wRb
LObNlDgqq2ZjC8jlvuFpPZCgWXFFu4zSvQpCmUkgf9d/w7/QQXxp7rNfQgoDmuskK8KnspBoMo7W
warrizEldmeJ3YyjaSsvmlG0C4Vq+GEIMKEqoTHnRjhxIknEJvY825IejEnXaVrueJvI/ClAWEHA
NJCOUaYwJoteX6psTKWe6JK7Of9MBNIMlZ8agOyC2dQe+8tyE1Sgs/R66mpenfPTKGEp50+51R+U
aplbIGP0VdCQm9sRrPizqbb8cbtzFJhml/qFOY6FadbfO7DDxaVzndGXAAsfssR97UDFhal+Xc9B
klONvba0hryFJBpnH7scG44OE8uONYYHs9rTgv0IP+aRyeExl89iAwHsNKiP1qsLTMbo0i44/FCl
8PT5eaL01wpXPjyKOjwadUcWlLtMvOJobAbzEq4c8FJ7EPMzO+cGe8d79st8jjLqjUK/HNjnh4XG
xPWU+aW/Ds9rk6T0sJiIePw8r9XYXSFNJzF6q9/GjTUpRm3GdXPjOTdRJDWp9QjNeLpx55NUsgoB
tbFMPbUIDT0sRs3YyIHYqDmHtvD8dPZtEqEdOIFAy52KBgByxpSyU3mX3wmG/PKrQ6w8ifQd/pSx
YstA2SguH8cjQF17TPz1krbpiuOozrYJp/gcKqAm4SGmlvjq7r8O5hQA5nx8/xQdLQgrONEsE/Fe
bEED26R25pkM3cHG8YE3xwYfxWVYGUS1Y+NGq3IJyX06MIv78a/UoBY+jPJ4fwBJhu2QOgaXeHjI
E7dcMrn6BI9GevY/b9lTP1+CyoMFDmWbMZF4v0NGjoPQOjUBNj3H7Ieh4WvBxsLR5tWtXL7GDsQj
ECOeGKnjArA6963ImkjcQronArOUqrtDagyC+PaWnXoCkKCb+8Fu029n0+GjiuMz7UhI10Ap1TdP
FGjbIbWOvtGk6eqjBef7+uFbq6ftke+NfYrSA+PG/5owK2TVg+ZHJDDz5nI8Fa2SIG5jyRq4qVr8
An0L/vvj8PSWHrQs7QGO5Rp4CdBcn3aAqJ6Ni1MYPVSrjDcecVM/abrPcuajSJP/QMphWwU/ISt1
0Moc9wruvHt9Wu2AwkdneHtqhIAW7DdUBPXbGcodWcc+9VEia6C14bqdtyPiv3vV6LJMFoK/wp1c
EgbOsZ+RLNIA+XoPcV8JixPWBkzcC1KW1cCGkCX2QJuphZWMii7O9hkCAqhaaSTqSLVE0qxoQxUZ
6OzDb57AZMnOUkKbMiqvWcVXv2slmyMlI9YQTAY4KBbCE+wN2CHyYfTwp33sfYNEh/38y46ygIqS
Zj5AgYM3ZigDp4tt5nIFmTzsn8JChGEwGKwYPtfsD3Xjikdklvit8TA05cTVEeWopeuVRo1W/dVJ
AHIji0wd0uFFrnG0MMHnzEDQMj6iK+de4VzJtJUCNwM3cLcfZ7C3zS9DBa/421JDm3udehjUsKok
iyemgASjQ5HJ/QV4sNF3ThdS5ZFYXOZ35c6yEUcPalU2H+wvaMaaujDgftnEP1J+TfI1bJYKC/97
QniMWoQh3znk8+Y/XUcs0kqJLjDf7PNOIJaFEUwV6Ch/dVaH9yA6qwjO8fQ7TzZD/Rap7cXKlL24
x6vwWQyWqyh+CbADxoyvZUqdczmTbexvZUjkqTXtw4AbWkPKbkYClUPfPHXg/eBGvmLuA1cqBodS
R4W1zyTGGBcPIAMRiz6a7xw+AGMt2Md69SUk9mSC9s03Jh6IqCDcNr78j1V3UmiJwOHyZWFw8gOj
OKIc/j68bVO2RoAh4i9FPWCca6nFI/BhA/Eq9a1YXc8g+DltEfZUW9zJDSSKUJzgX4ocfkMQN2hx
Gog886zFLhCsEDLaVN3WfJSRGX/Gl/endJwu6dNt4118dPEpegvzptx2GgiLc9IWph5iXqQQ1SMc
SROmudQI8n42FviClZlKBbRc+u/ZJXMf+/GzWjEk0ZmkUbcXnbT9rgN1WbZBXogkgUZ4zU0v0drZ
9vBZAF6qmiB9F+pqec6Mpzqz2EMdAkCimqeJA1Rp1n0/iSccX3cpY4qVdbEx1r8DY4moWAaYXsDB
9vL96Z5VhxOjvgwM26TnVqtH62L1snIPM2N6tKrTgpTCXcTGisqG+SRRcJEEeCvJ1Cf2rWFBYp7B
3AWL+fDZ0XmWJsnjbM2G0NF3BKg+R7E+yKASCfj7fM2Cs6tqx/GODr3eKHI4d4nOyOl7a1lPdzii
jTq7BkcCdu0D3o3jOTJzPl9awcEZU6NLi/XAjhEGmug/drt2cOnCW23Vsewf0Ykgiwvf1YpYF6g9
8xJMUe4DhOaDV6Y6kG7s/xA7Dp6URCcg3BwbVBp9vHuBw/hESaGkl6J3YwLhhvXPRYjty3vAH7ZS
i1ynh9dg0ZYXw2jm86S4dYGYs5wXgQLNAXDGAvgFAoxmP7rj8yj9cN6Q9VfCi2/QbSmF/hrfGH97
9tbFOHb5hrVZmVYRY+UKij6gato5AFxA8raO7qbNjfogf5/Oal+dVEK8MEO3VrjCxvN3HiR2JMRI
2qCKDtxaW/9prCousir9/Ahrt5m4wDZ+M12VyCgdlWv9EZJRadrFIgQn8Z3bzbZy/7lvnYCWetXe
OKOziy8hkkuaMXfI11ESjMzQkhE7/JIv91SRRns0h8zIdw4BeoeTP8NknfZcrUUH4b5SEFtqpE2X
+HJ4xrBCusDw/FQpLnOROiDrYHh3HSeCg9razHg1krYZ2GsbH6c6dNlwAThHbQAPiNWxmcWIgU4F
IDqoe+8/IPLxj8VHyDK2NMOaMKwaIyvoiqXfFbs0hajNFBLsQjTsdpuh/OqgPHkDfDAGud5yHUa8
jmkKUx6hFohTq/ER40Sk1Pm63Jh75VV+jreLpgpfj/FwDOAsGPVxYKTRPp47Wtool2YCtAe3U1vg
w398NKD83Qd/lkTUjFpfIjqT1fJDBe6zd2IqVgzgBFjREZVUMYuu7TzNr3eySbN43Fdd3zjowK0j
gKHgvona1Uaqvi5RgXS94+/cM9HPZx5ZJmEY7NP4Z3ZxaLhpS6R+hxiTAnIsEdu/uN4M5hue7kwq
MWNYeYWF99KFchxv3SfRny6nZHVtVWLjw7x+plaKbi2Trc/VTWeJV5thVhS1M+U6TEfZ0BoHPqlr
YbOI9xGUXB9SMAfDZOKHuD84ZTlUjeqLIkxnAiaB+Z+/e9wR9CWFr+oXMsAlIi09SbEKGdFOVDKK
w3m42ZkU3iyUpYM+4FotgYLhiaHbmfXNLul1JUTPdUoMLfl/TXYtvhpfXSGlq7EddcPAnheRqBq0
KxNltEubfsZJU1crXvrAenKO5eg6FK574pOdPb5jjwZ0SnGXmqfh427gHpUjcjKwUaljrfCf/F2H
xUU0dSelq7SASHEAK6RKFxgXk8dNG80h4m6jpQXwzPXYW4YIBCNLt0/JPD3LB3GQgjr2l8Glrx5K
WyRsFhv8XVL8jYikT+r5RvOjmehRtADM9wD7J30diueif5+/WWWUsxku30jkSoWlJC89/ghpXWJH
EiGuoer66fGUkH+qVxSypjIexiS6Dj5UPIZkXMGe9UIhbtWkufhUWTGTiyhEkMEwvpSLzZ7+dXrm
Rk0lJUwKRCagKWxjcxFOFgU3/HutoCwOEIxExaW4UYBv1C2mVRRyDWP02ak6+N4qOM4X6uFrLqpC
5DAszBCnfTyFephzpISAftqeMYIkvIcPkkeALD43XP/Tz6DUOKWh0KbJijjvZ6gtvLJ4be5aTn4P
TjHAWl2cs2qjIyfFRJ/kSs7Gd7VU8znL/zMWvARs3ge8ZZTmbQqG42cv8/0t9WAJorV0sRJPomvs
yotzFZgucfF7RPzi2rKilksxUfLw7qHKlymTf+5U9cDSuDcPoMsBiiDOW8tf3JRq70+52lZPG6QH
T6NZa9glthRy2Kh32yUPzMDaqwNYpjLBocVql0OvoZYPlcX2GLWRsxh187xUZeNwMP+YfYr6LpKd
8auNj3Bcy38hqq/kw7PBT/YtFLFdMnZv0vKmExCfzbHGhi+FNcTPN1Kw/al4MuF7hS/iKCJRSY9j
Y8ykmz4oO31mRV1Vt0Ggj6+sDbMqljsCjMleeOJT3woazBi0MXREi9v3gekofyEINsLnWpw3B6Bq
mCq4ZLOeV7amsrOIQNjs/eW2Um3OSGGAanWogHE0tIWqwsbyMH9BpI7N7DLctupbDyszlj4xDUtx
L+HYJE9IhofqxMkT9L0K1I/1+VxbL9SoN/GVEw6PbEFmplVectdp2+UvJZIEf+XiX+ymWsm38Dmi
gkoERzzqEEcNxt1rQwug3XYwlKLcT8m8+7/b6FOtPTNjwiBIzJRaHP6ncfZAbo0vpj5wdVgPnGq2
vEXgcj9zdvisIAyzXQMv6e/AeDVKVELRlWFNc6c5WHqqFqoMcGXaKe+CjnsthXDngrpMc43VGcJ0
M8HrmfV4I5pKJCTSRtEn27/h3HUBYr3z/Fsgt1SCVM4H4RGqUDtRR3pqoY8laQ8xszVZ4PZK2a44
xcDZdaZuP1k3nxzXVgV0o2kMAngMThZehLlOujmwAUG7pFEFQdcIhtHaauxLt5LQHMBcMESo1zRe
5FzHelPtDwCBn+CybyHgWZAep0fFpTs02Vgr4Jwbc49G6B/XjkZ9/p5qKFI2V1tcD9b9EqjfeACm
CfA7LMEMh5XFEkjcWndUjA/QZji8co4/RPJ+JjU/Cncg+eGu9XlWwFbnUD7xTMUs5V5BzMvZFOio
lWiwcAusOgWsfmi9Qq2nwCH18nrrs4nfqiwmhlB2Y5lKMF45GH7xiR8f/ZutDkMsDJjbsPHje1l/
DwSCgxetOqXcz+xKNFV2j2ui2w8XTPAMDUBmZRl7kmk8Tv3zBN58CKNJ/FlhQYk1OxJ8YewecFib
OvsLzgGb5cEgzBETLTdsemNlWDBNJg/jKShNWuaYwRhwnVPHp25viPzqnMe0/aw71FnwF3JaIT7g
kAty09dQpB7KUY/jzXoUTuvUmI0eS6EF+3hB8ID4DbB8vEI54KpE4molBcibiBVZtoF4nL3+MbUg
Qb0EYKYnaVctv3Ctb96ATV+t0a89JyV3oVzdc2lLcTT0rBguMS6aGpHC5U3Q6I09P4COliWrWcyw
rXknsS9vPZH5pClQWBuJSfptBamtZaEBC5UURudkEWQU7Gd2ZCjpvRogob3FNRSwFRg+Mi13EHlu
mOjOZ3Tu441hKBHXd4srTRoVb8bmXFTQcCCbTdoIf5JD/9tMYtRWbt16rmnr7sSkG8qwqOoOktpm
HFKdG2J0xFDkKxyzAM1fochgy8wBENUKkcsU+bmj9eesyJ/s9F3TjmhHjFHwS67p7AknshvdNSv4
LVaD/yEm4wXs8Dtdpsh5ehj9BNKUpoWii60qEknFremQK+TW2QE6TZExcQvVTw4w3SKIpOG0cIrq
CWh2+v3FQmAIU4suVgYKv4+Fm39OD1ncc5RtPOz/kB3uLrR+hgDdLQbcK74YVhzXDHHQXVfmVKYD
a9cpvsSIkq5bcjyWYInJM3vBx8Kb3s2ZhZzLlCLmqZbED3aP6oYC3G2MyN0RfQn2T/A3OBe4+DIC
FPcmWLCzBVHHWrNnWnEsWFdqTZUcPfv5OWGTjYYGDfZ5P72Ix5xwk7MMYGSTXimVN2uDVLTVudUz
rwx/Rv5NXRSFPrWr18g+UxDmBEgdK2zo7Zfc6cXtYk3VujOh6KQE3J3CI7oTz93O+ABoOFFowLPB
e21YJ7qcIXhyAWaMfZDRRbqIB7XRb/qWY4FXvUrEiZM9ShI/k7EXvx1dK9L85O0wwvN7PcOvPafH
PFOIELbWypXfoMzWPWztTuHwPI6rLfTunwZuQJUFUT6nMmYXGqUBhYu9tbPgAsBC7s+/For5H+En
pVlHWAQaDCDCggXjDpkGQ+bGTLn/m+GBA/U74kAHsoqzw82JRTLSajq73IR3jhy7tWoF6+dity26
626KwMRGbRvk7zF4582Kzb4nfUTKgG/0JQiTKhhf1O8Z+oU6gtPc86CZBKqTaN89xW8+x+Plc1dI
jW5nQ/wTi0YqaPrG5dCixnViDBMm4G8Yv0YANpG3w24O4n+SO3qD8/ThzrIngrRwDGLgDimDm8zo
7LwVMTkKI7Lu+l1ssR5+ZW88VTk/7BJkIpqAMkSSJKstziv93eI+dFFUHWLvCNZ/xEEF/q9Xiu7B
eCZfmazV25xFUAmaGsMCH7cMqfQEuIrfvi1nPeDMexoFXK2o4v1hs6QN4g+VzKdD8FSVcv3RVRdR
K3Eb+ddCBu0M6NZ4mQVcVy7ZfLSz+bJWdVr5wFMHtGw0MqLJ546YZQjYN2gOl9yJF6JRgT6fsP7w
TNN+bxtIoLraKJct4wJVmz1H+tW9p5o7AKaDag6kz8/QVq23SWusm86tH83g0I5KJ4F0cECSEaxI
Hn1PLPswEPHnALfR2kEdeKsDVdPSWSHRsX+BIdW+5MxqdA0ZSksa3M8gyTL0KXXihg2JbOY6uEpU
vWJP+M3nnuOZSkVVrWdpc7cx4bdnHtksBGzC/gm0kCPZYkj4g6IFaG8QFOEZ6HmNWS6E8CEUHWbR
L14Ow4JTrTJfzc/7BAiuyEIOO3YyU6uswkCe/SsoY74dLzUZSN/fpq4bFweVAEN2LgBDFTJ9OqDj
5hfXAL4zDqBg3JkWpl7DkKVq2Uo4+GHlfilUABBe3CxY+Du5FY4xLMPp1clhfj8dfPf1nVfPdavp
7dPttMODnTR6Tiuq7w51eFlMrYVbtUgEE63PtRmP/bEXdogAWRZbQfVXRD3XHIxQax+OWqV+238h
IUKVTgvw3SV0yqmfoRe/mj9rR+nPf0HZWPrV0NL1EOsRiYbreSUZmErHtovTt7eCdxj6qosc+WwA
LUUVzDSAcmpnivOwizsIhqS0ySj9/C3XyPx0ilD94HKvYq4R7SdfM0sAlrmguu0bs+bHhiMjQYgc
U+AA8IFw6NKrDJtoexUQvhKgs7WsJBw86GekZTZRid6jIl09lpcRRDEmuBoiUvRd7GRpdq3pU1y1
nxjf9WxQgWL7MhrppDteOjaZD2bTj6hRVWvdo6/pI6BqHvxc+y9FgYEbUXJl3r6ReFBAKHt1JWQJ
zqte7kKBJsKHELNP+5HSK4JJ0NJB2vGYmvCyLn/TMptvzoFkDxVPLCYvUk2wS0MLgyoIeyJOMoh7
iFFMKGP0C2BZXJl0OA3B5TisV/D8CFGnajU51qY6fs6GbDyIxNR5QtXZlRV05uCQ1MTDRjL7fG/P
Vp1JAEcXolkJYLe0jiAIpFjhpjMzzm90+bvRaR+boJETOCPYE4iGrW/S9jQTxw4qOFCtdJ8DAsaj
SF03wqJVu1lDfD0XUiYqL2h0ygM/Vr/N5u33bzkFWr3g8xvazKC/OGd3I9BDJWOSd+7MRBdpmZXQ
S/TpFMphJmj7T2c+ewmspcdwxPyESkEu4uG5sGld/izjXDC+GQio9CwZunVdXO10Am5Kz3szaADD
B/zcJ93pF6mdijt7sZtkpTc4rAFfVjMvVch2HEJdFt5I4uX1g3ko7sXPic6zU35Lq5aBZYqZ3wEw
USeAVDnVnNgZ0zGDPp+cLV956usAN6RJ39BzcuvS2UVarEdNX3sJGQe7VnaXIT7dFehG3+wG6SYH
tzBngZhYT5lDwQGYLyywaUnkPHsLQT8Da7Y3c4wv4W4EocoKB3mL8vS82lLLlw6FCMGzRDap2Fys
zz/yvoDMt++ZOboFprK3a4pehpS9H+pEOj0iBuoirQXwN99nv4nRxDxhVFb0FQCXnbudInepU4k3
DO5MTDJGcfMnlt2TWiNPq2FeAYYuO6/VHCn/BLr8gGr66BEKltLVXcyGAIKztDunP0LSKUVRDIfe
a6Mb6yXvl6HzIkDL43Meoy7gxUWttk5Gomov4sFYgRJe8N7UpzR9Ej0Hzsd8yFlysDl3ck+TvFX4
xZt3RYcn2DQ3FR/TaXjPyZRGbdR2RANb7icllV8lTX2Px8P9y/6oJiKqsOP/LVVcv/6dr4miYlyq
NtoYw3EFe+7ca/3MMo4sIyN1y5Io7RwlDqsiazqMWnCqMV+lOJngMgL2WBpdjTx2GyVGzbXfaMBO
mvCGRQR3YIhTrQBA3PVpCr5Jw23OjqzCLveqLHp21A1UDcwtfi5jWVYg2Yc+jsYhWIIZYXdURDRK
wOHMnLQGymn8nVTzzzHzOyq8R1lkRdpS9+ZiyJFhDUDP8cbmgzK1klFm+KRX0LvAkSVQ043VHdUU
wNCsdeHFt902LxeSZhdnk4isEODxHE0qe7Ge0Bdk4pE0pMGDhdRfQDFCxYY9HpBZ7bP6jHh+C1nK
p9HonsZe3kXe7RHOg3MmUZ4JFo5oDYk9Z9IT4bYvyNMs6spdn3QiJShnwCulDiEvPsQxaUV8oJIu
UO5ylc+MfTffVWVI3ufA0oTveiNRr4Xd6bVTFBETsu5k3aoHaA/jGe4kJyfCCYGLpWaXoKSvl4kH
TvU/agjEvg5oQMxUpuYzHmuFWz1d8jjEt+T5+oQ6UNLE3ZlHvstEsgvC8AsDUunmTSdK2LJHRAyJ
m6spqiTqg2y9+P7N9AzC+NDVuHVxSDl1NI5750bhZU26iIYOzD2nkN+eax5luaVaTXjxSwjnOfbD
YEqM32yMjVSk0trUMyA1hnvJ8GPgwKXUImdN1vGJ/jZnkokT+s+lNrQdJI/6kAe5RSNOzf5e3tGt
oR07jACWhWFUr9MzkjVvbQJLgMlBEtCijkcHSE/sJ2bEvk1x2SGjrp/Z/V8IS3ppb/rgFjANOVjx
Xv0ZoZLFvm02adRS8IR/WoezDH1B1VZrLEOka2G9E2yxdZaBaiqQLyLZOFpt/J8hzNi5aeR8d4mX
Zv5nXQCXwPlAM8jX/njIR/8PyINIIPl/EWK7LWCWh7oSCx+geDRDuEKLNsjEFGk1zWrTJLodMz9o
FFvfkLVwxmC+9/e85U191UBE382Zunw5fT2D19P6plzZvoidwdQe9+QDEW0XpcysbhyWoCiXaTmu
QqVhq1ojhMycBRiFGpWUUVtXMbKLDDPp8g7fjr0ad8yhmOmItsgf9SlOEA/YmZM7bLRIaiEwIGIE
ZColHugo/xlrbxkFqafGvcbIagNsnyAilRTHPeuMWcasAdRu0++1/1OEg4p0V8EqLuMW6TGZMepf
vTz5LCdCQm90gYGZy7elRuaJquw1O6Db4nxVXZpL87MCsyo3G0gIO4n5fMd63J9j3s/vZoRfjwO4
NzGhT2vFmY0vXE5p73Z8xhav5Khler61+J8i+AF/0ZzHX2MGHx720nsBdlSTu0e9viX3A1u6mkIw
LtcuhcOxmUAxv6ktJrzzBt09UwhU1FA1f2D8tEgGql+230YSrtpDqNoKAZ5Wj7grTY/iuMPjIVWA
PPFvP3ZTIf4667EzUmKFMy9y2enAQpAXqIfl0gsatXP+9lWrXgN6FXsiUnLS5YhGXRMjH03Rhm5N
4LwsVnlLd4rFliAcm1rV54FIKV8cZzaFSHZF1EAVPw2odHEBkHGMQw9WeXdbLTY6eaJUypvnbffZ
a0jEOJ72k8aIt6V1D/EOtbHIGLzUlF+yuF/cu5BuAC7ABuk0QpfpNyMau0K0BsuNLrBuyDr3VN/u
Zr1Tw4hUY3CE5oIQxbp2eq8dz0CUIiwwkRNGH5SuB5XlRMeo41kswrVmDiWJOtpmdutrGI16n6PF
g7YcYoc4NXEZ4RcTYW3F0gyWN0l+rw7al1DTWMLKJpxPCYNSvRh1051OABGa/5FgNMEd63c2rzVw
GnhzXjUL9kp+Ycm9/hJ33n+CW3xE4Hk/0rBGUAjaGeAQy4ZwlJBZI7wJ5yZNSkgfdDogFuWJKoJZ
HvwWME0kaLVyIqCLIk70VAGIGSRX00Uc77PmS/Raes0Hxbo2ua5z0QJksOX83xz0qF0Ey+MVeWdv
yzXU8BfP+droFOHJfjGPGwUiHmt0lU36YUs1lTOJMOfaRzrmFaVUXI8KHr7vhkKIGTMRBYHAnz5r
YJTOAgGt0bCSdYq6vgmrCS9TzzYhGdMsx//LXTLVIo9wp1VSnLyCXh2YSRx6SleWwYilnmxIbaPt
fzNg8u2wzwWrpNMMDIYBcvAUAynzVr0TYbdMf1BMl/3ldqj2yQE/O64VILRYNBQABpmI8v1p8xUQ
QEKfFOtzVX4gaxs8zN8vb0ppa/FCo+ohT6rOjMw1lmDkueMIzJZMTc/is8M8yvf2UkTKWoPYuxH3
/BVWlAAkLDYgeKkI0+YCZoYkklnlLumX9x2R4OZDKgmg66JqaMv6jKEI9lLaAbRIB9TVewcgiXIb
xTKkEwcTsogRvzax4bhWoW2X+c/Xn3mYnyBH5FMRIAYV8fmzbVvbSg6tZ5B93yGIbxiKw3RocMrZ
oK2PzAObrBoTnVVRkiIcx5bX+0RbvCXzotkAeE0Ho7KrE+OD6t4/PckzgCv0TfxlmZcdUbK6L0KO
O7xnfolzswwW3Buzenek1oNE2BPm2YZHyz0Qrww//y+g7ldSxTPzquffYV+6pxLmXSXEI3+g1OZx
WPo7cDoIxfwKmfwLyE2EBScZ2H9VbGJDxMtAes0IISGTlSoMw2dxAc0Fd46/VRFdy088oRX+dkCc
hrc1PiPi1eIZV9wQ823mJahUSib7Jb7RBvINftEFQJcZ+/J3NB6A461iRMRxBbKMyu3GLPv2TqfJ
XxLXAQqXJ8e6YjN/qbkQRc1TKVv2jVajqRu6BbuSlQ7HgzbN+/5yrlR9FReqRChHlrBmiAoUjGkm
dYtToHOE7RDpmH9WidAqomY3OOXyFgkQmGN3ZE7j0peVVie2sQ415nGbD2GJ27ZVJ1r+0hFEntx3
HRp7AL7tjR0uvncLv0wfpMX0auHPOqL9GzDMrFCyBUp1NY/3G1WV/ZARobTJrRyNoHfjN6RdStxP
9pMason6j5P3RNW5v1GaGXzBqKSMgV2iAVL9ACCbU9t5sIg259u0Et+sNJiMXlCVaixKRnIGpPUL
2AUhgb66Hgvl9t+3YDi4IcoRxbkBKLcGIC/fr1r36aw3JUh4rRrlHtDU6dnZPFRF4kjvMYzj44yG
jXrl5BdbMpr5If0wTzXRfQ/4MZEAX4f5io3IlWdlfhXG3o8ZDLEXBGNcw7bVbxhSJEHcI0RGL4Vy
0QSnADoezAJ1NLQVSKReatrsdHEiNblS9cIOP7isT9j06qq/oVZsoH2L01rw31iapdFlb3dM94pf
3iKr8XOFkyfCuT38mEanM9RpB8DFakisPfzyqVS38GkxwVeLnlXu9IfZw9SOJ36FuapIsn58Jn4H
EDIE40eVLkwyYke4ENOlPuu7y5vTYGh5QTTeSQDvttIh+YzT8w4hpdDF+7fK0OLdpR3ATzhp6MmS
Wyg+zwHy+U6ltEf1yy0LAN0HVPOjNwGfKIEftNt0c/6lcqX+DTQW2dpo5OJgrOAk8ZswNiUwl3ux
w6PtneKPI50Aqz1o0tSATsRhcNQLflAaNHiblvpTsxVEIcsPRQzvirtPAVRWo5Dv6RtgMGHIqy3W
cWTQHpaj+nFlgdqoVVdN3VJ2oFQDjwhDcN6dl9a3rPmynjTHghw7Wq+kbiDh6NDDiifaJnaOBygQ
ctRMtonlcttN9R18l0SYzcs5H3PzePXIqRh9G9GHFL8iqlC3P5ocBC9vp2CSMuyKb9bi0MAZ7/Kk
MtoukPDemGKSg1TB5i+HRSdCRy79k+jZhUlPRv/AGWYC0JeF3OlaXFZquQNQQPqzaxNbUQBBMpqO
tAXhFFAiJss4nburkVyDlOVTQnea3it10gruJk+ByUThp9svuGp6/hrHiwX0UIbYjYVAuVbgJjQK
kJbUvqpZAv1mcM/EhM6ysNNy0NhRv1Zz9jYdPjwxjqYn6RoDQalx5fbAE0y72zr4Bj0n1FO7QATp
ZdE770D/UKTA221JagxC1einmStcJDmNWzZk6BVjx2I08T/+kKq9BZWxPhkOohjDebv82PmiE+DT
ghD54yHV0TM7xH+/8TEoDo2bJa/ZLtEKq7F6hDKBrOGc8VAKSBfa3YuW1Dr9luYCZxpdFRPBfNws
HuSD7qoyczmiRC5/DmpW8VvSN66CHriF3yMnebkNcY9ePPQvXWuPHn3cBaCvFzYWEwTFGCHg+/Pv
9S1clghdygn4m4Cq+A39n3ExrCP/40OiaRZba/+CclrJxkv84/JGu+okl23wKCLoJgOHSPQMya0H
CKbcCfArGbivSoH0Gnnsk4Wp783lXyPPtCWDX2DQ6L+8I1fkfmifAiqZV7HsNuroZeS+D/DPNarF
piybueWO5jyySekHks0sy/cFeDYA6JGouR8iN5ti+dqxJgzMP7rJ74zXUvCxJzRn96Wk8sUCjQfw
oYny9yEPpXW75lGF42VpzxNuZwzUcTnAmQ3PAtPXFFnaTjbN4XdXQI9EEWjFAG+/tJrms6TGf8hO
8gOXp7FIQU26Ue2sTxDou2qKhtQQcEfJT3TTrC0ztDbKBbAEmC825CvAQMDTpcqvd4DO39eH7s9V
atJkm9kSifEFzP7yvooVHvj9aux+CEJDYSxLHuxLkNpNzu1ueunxIUzomF2EIAr3YnX12gJTziER
l2OgiTzgbTdzJGEsbHG+qmLSECd3zPlJxhBat84bOMukpFP+nKbq6XMACo0thY41T8BbU0htbSxy
nBbWUJWfuLSOelZkAiA2aCOGDFj8avrqiPqhr4/aEq0VijECvph+1Gvds05EeSlp5jKmV8S9LqL+
cHJBBSbUfAiY3Z4llycsdbw5w5Fcc92EI1t2amnfdVLRMDEWMnCd7zfC0X1u7XuOIwKvjo4ezaNJ
7E89gUtmjUXWAIJMbquNtAyVHj6m3WPzpNZ4t1WtMF5O9jpQmKohO7D4IUMRCFDdMfoOCzhI8KtA
GFa5Nw4YdjRYH2lppif0P/D7zOzPDpptdJFV5wgief7YMtZGbHMDKTiSAVqDc3KG6CztJ2tEeHzX
TpOCodx9gir2tzg5C2neJQok2De59PrEfQ5TkoHV/lG++owTFkLbwL+M23Vb52XgPLDftGcdNxMC
yDla54QPty63F9d/anwf1A654hzCFzQTsjPAXQXAWWu3ZOUjKj7gR6S2c6uWC1rZSTTljqAWQBRg
7koGV4oYJ+2v5p5bj4yvysI6hOyvgUavsPWyljtijIxstLnsYShGG40KuQzpeWUajj3OTHlYQkNf
OyzcOP+7Ffrfm8G25YwLfqQDWVOFBNDKy2czIv0FIAPNauFe2mbWuF5tq5hi/mWWzgItKyD4Rmhi
Eo+hpVb+3BWdtcNkutVumLx7VYzj/Ms3iPxS4iYtifrYL1YfLGhn3K8no6iozO+FCTrcKHoXrkKQ
rEwqxhx5EsVEJRYoEKuldmMF1EhJPKbfHYxbDfdhl3W2rW0PtLoNpMhPIpsiF6YBJX3OgazDdjjE
FqXYFVrDwuCm39poRr38BDuF/cNpUTKFTihZaogzbWw/H6g5QnA1CtxETSwkl4mtfjc7JBYu9Reh
Xg4QJRmNUz4H4SABO+qAJEBYgTeszh1/kRiKBSNLCF1l+XmEx8xfQfw+jwrQJA6hfCmmIVxHG35t
MPoenVn0QrQuEcpiGLlvfKWRjNtDvgHpTu/2Ret53vJ7IumjXIIx6WRQhuV4v2n85N3VZzExa4OH
y/bIZpPXcb5WD1pc13G0hbe6fmyBUYUc8M99afyj3/UPUbp/U7oSMn6zPVdKjajU83ot1YYcayDp
UDVMZgJpR/iubUz1Vry88fukTGbGUajO1R+VROvCyXIBBRHJqyWkmvDRMFem54txb80MR1vHgpIe
fBeOB6PnXBaFirt+lkvYK+R5Bg2vsIMgrTuF/4W4ud/FderoMtceWddvA8sb1VwYcnDtO5NxrBcx
/xxDb+oTsZvjUiT73+KDKBYfQOCeqnfWcUNy3wWp7lrRlDznpzkFcnZyETfItFQslcXBCT4aW6et
PYyz056unThq/5whjOurJUSIClNxeeB10d0vEVzgWkb6DfwjhYtlMfyA2REIQ9ytf0IiXR2/i5HM
fbvpRNbDaJ+gn3sXTft/l3iZFCitmz3nBBVy5YMpRJasUzXGKg+X0UrX7kLsJx6Ir+NeXEQBgegR
2XTuU3t3L961p2k5Feoc63MqMc/ADGWqyBqoJ2XWZWVFLrKzBJ+XhSgHMjn3FOLRqMqZaUCSbMMt
ODrP/lJcnd5hu0y6iIs5UobYjgOU9dJS1M+0SApFFhT72tmlPzkkmK89lS5XaU6SfvJQw1QDaE/p
CetQo/+jhqh94G8mII1mluZoiRTRP7SYpD6oD2JoDId3fdMrvcT1gvi7iOi/9SGJ5s5NKC6hxOBU
3hj0l9bN2NK5Ow0a67WFGqIhKqDRALdT8ZBR1S7lQCnnfAu9beWO9LCoddE/qkrj6o3+4mzqHBpi
Mc3Hfk9kJFiZIhMFSd2UPvXJQ9bvzMRXFiG7bB5C31I2QfG+sZHJdIXpwHAoP9dmCht5v5/2o8Qm
o/H7wQ72WvxW++kKngXh0H69g9+9XnGipPoT/GcgJjdOwbPUA1Yr/rrGYdEot5N7uZmJ77Vr14P+
1fOSKzJxf2pmYW3HpPAe64RCTVv3wYGtp/0f8PZAoidlWsC8ao+gWDgwlebQfjetDpzmhvKxfzP1
NwyWoJIdU9kRUbZknvWmUuAhDQzJIQ4znxZxke0+csaPMl/XPc0PKQoEJgNc2QwZqQ+uD2O2XUeG
Xltp35aNxL65wWs0rmstRj0aTac6qwDtbPTLsNrMLvx/hJwIHJT4kZ4PdUfONbJxZ/7GVbMhCU5D
flyzDJxLBdfb9xbeqwoaRAGEUiXmRYT6YlHgiwBxED5HpkZVz3v50QGGWD1+6h3Oj60X/3KdvBW7
jMmf1d6DcNAC/FB5yVhdbAfQVaIJLq6kqwRppK7TVLZuJ2ix/KnctRokvKpwxL5LKAVl0/vo8PHm
N0uEH8OwQ9x6Giyz41QT0gw/ioX9YTYlp4RO/XrYY+UaNKf05Gw5A4IT+SnZ0+cR72HFfWF4qXTV
FxZNBQoBbbp/lyJVY1rycytrv5k7CxfXHdyVs9Q7HnDtCQtvOZHrsA7u2bRwhA65GQ1GsvESXWr0
F3+LZCPtw7i/ATcfT52mAvy1c6QXXIU8CDB0uLAvCX+x8lJjplqUrtFAhajElwUI6V2n30EjqZuf
2QFw3jOLTNs0h080fCYOBPnyGvWJyOet7b4F8gKIRKsO1TgdZChIssTBZX44Yv1+Lxjrhm9Z4DXm
zwukmcZCWZAiE8S0AYQ3WrHPHYScqF/6e0exkK2XaYjRU7M3B6c5g07R26qUINPP2qkP8CP9birW
qAraqW/cUZUOGiPHOnjzPbFcsIUreLeEoSuHItOzM8WeHOL/LRnier8UPSHM6NpcCAvAucIegsWV
7t3kf1mn6GgkzJ9TlXtmddMj02y/CfHExsjsJvvxHgTzkS0CfAMb/RXV4HpBjkq04eU/tZ9a0BKc
0cd2KwtJ0DhxFj08c4THHbslsZ+JETtV6/W1yREiXrKOLJO8JFjLh3OhNlVAiX3NB1FZ0HssGMPj
YhWGtKoK3HGzqaXQMfqbi4St4ipO00JiEO+UOnZwgUnLlSnR/G1pAm82LQNngnUZkQDeW+cPopnW
eGLWFcjqZ/ej0vzMc4jKLmoQQV4q4fPhE+CfqWecU4WuWpF4EN/q66oVGYo0p9/WkyUnk89FwdR+
aWkh0kqcwBi9aoBkHVBLli/+AvibpB86ABzBYNAkI0DlkJlpPQEpeesrTeiOFfAzDQXd7XABVNQD
d/6ENcB5Hvit7fTY6liGYRS//jk8KKDxM3oIS49j+H9dAVdVPHO0x14aQJGHr6bf2drDjldY6kom
+4dRZ0CDxcMZY1ykD1azGsz8lk8rB+BgopC6a4IjNV90izXgF6J/Cl1arpEG9UTX2Yob7D49r1YQ
QVDnGYXyrMw3HMlf2n54DYVoMCZc3UeW4ZEvRGG6p+rqJpTWEUKx41EioiEcS5QUezKDIQOueE3Z
X95pS3RgMBocLPOKrco0/+I6VvlQFouBbwKGDsNqY6rFm8IkfvVvfWYsiQicMNPJQ9FOsJ0JpDS+
O6nNqzUgTBzp3NxHDsOFAEsIMHtRIuL24WH10jFjusHgBCLQsr2BJQLRIvv4iAITP9uNI30I0X99
FC7TLNqX2tgcAnfSwYJCkpKQy7ZFDeIBXsXZt3d81w7kRbcak46gIqHEOqDupBx/HiZEqTSBTeNO
w/fbtKRWLm6lsKsWVR9WCuQX4kCaUOPYCOBvW2J4ks9tnpTtbXm6tuRgIPtNcZVYS1dclZ3u6w+H
RJvogGlK2EyojFzEA6gFhBuwNJ122DQ+WiUz/y9XxK+agCjVcRdZAeNVIcrN5guPOkTBmky2BsDD
gMqdRFqFFSzVPxB6Goc544F8lIaz3XG/r57vMwKX2Sk8ou5+HBP+3Ks8WFTUqeS3FZsGCaD/mo87
0QCglX2oZvskc5lyP+xM00RYSEfknqn1+WS+cjjtBQXsgo2rPgkV3bZSCWenOWNHZFI5GehHN9AK
OACSEeoW8QMX8lZfiqG92gUTl06GqiJWeO8y12Pj4/HhgxgCp4Cv880nZla4pl5Ha/6UZA0Is6BK
g4Y/Kh2Y170ActsPeFu9Wkz6Pd8G82fACrTtU7d9wlq//L8EQuL+R4UkxBDm6wllbis6HzGduRlq
lm5Lg8nEjFBTCeq3z8w6cmWMqbytPitAYo6hjZ4/1F1OaMeB6w53UXws3gTc8QyFG/kB6Dvb1yc3
SR/YQhuPgA9r/cDM3Gs09z8UBTcxmHeBCBpgQOIARGlp/fC4+qfiYYboprzzn1H34jXXPGOGdByc
5Z+I4KlmfQ51Mvr2I+oOueGFGSIj6KVPtrcV3dkn9Mcp6SbcHnFPDQqJtesj/CmLrvTjt5yerWUP
6hcihNFf6g5+2XQeJklJRAACDoYxXgUIqoAK4h50QqMziZCctjAm270vwTPSXY8jnpFIhHhxmuUw
BDssf2inzGYkQnyn9dBnpBr5p8BuAjAAArmTH1UGJSagtrrVB44vUkKtzY6ZNRqrJwtaT8I1RRMX
X8cOUayr8FrA79g0hPra5t3S/e/bSHVJI0v9T4DkmOI3GxbFtXPdkUfQ7ZzEjbSa3D9uFndR4Sdx
iET8mYal5dNmaqThUAuQoadi+XC/FysPuZx2HSd/QMcQz5ADGXE8wIjZS3evbgy5nDkWQYzpdSEP
Icu5QN2yOY2dB8Y80WtjcGaozv9Y1PHB/SOzsK9ccgJFotT/q/NLL37FNTfatjIB4YpLI7Pjn0yx
FWHa6kbzDh/y/e9YTbW4ozFTitGxA/GzijI3yCx2NhYOVGqeEqIO1x9XaEMF5vVpmWkCd40ahSJ4
nPghxPaheawUUxUgKacjpE8+FfmIje8HOx/TDrfiF1O95x+swvqdGn1HHZdXhbaDJPF+49X/3qTh
2JDoVK2HFJ0K/UulVFEvHWbbRZw6HT/jXlThabZZKuGHzHkE5aRwGgVlBt9UaBW0BuKvdV1bbKvt
mSOD29F150SkyNBBfvYRj8icoEQAqe6iBOopTvJ0Z01if76NyRtW9ngTyOJ+GpIajwaSeAU3nGkO
J+j2TAYhVKqxsGGCZgGkOCLhUx4zeQLEsODreLB2EL3j9jYMYA5LNlnfzNFtWa02fCsPka2jO+L3
TDCNfZWKX1+3BV9QUwJkq31bjGkPnFzCOR/8MWPGWo/dTLobzBxEcJuXEGGSSeIod9BZlSa2QmRn
SvsR/SEbHitH9aPBDOgw/MxdoL9AoipxX1dYwLRaWgxWr8Znd1aTo42BGfoxWED16O0IjXxicNEr
cZS/taR0WcTNC7J1uA4Kv3194hR3tWoQOFyrLKwzVG7csot+XrqY14D63hx7GC0haA1Xh1RHQfFV
0gnwCYf9SfEGK/i21v1/5+MWsFFEQlnLWtaSxHsuQZttXJxwHUZyTq5FLEEelIeTMi99TAnVVVlZ
r+RasmXawTuxPYu/sLFWOJZ2dWCfacaha6xGsrNP12spSjduwW0HD0HlL1HhRKINiyq15rlw66/M
Guzd4IGIqkOf5kQcTr8Zwt2dQtfdAEbZWM8j+DDXleJC3VaIdDTEM0dp78MY6qPNeL9S+uYWwLS9
xooS1OyI2+jMZ/pcFqfojKLBWsBqupCr6hw6N2Lu7v90flYXwnRb8QhQvPbWa8EJuYQ1TNVkC7hs
Jt7W7wXhHj3L9ZwbpjL4n74Edju9rNnT8p+FxYe+a9NtLPyPgAPdtxZNMVhS6UgXxHr3iBKYv9KA
T0mj6jjiRAc9IoFP7C5q/CnIzyRzYAU7rA7jCWxBX+Dooj68sYEbTEolH+veuk91JlaSw88+1aVI
O2Rnj0smwYNs7cgpVkfEQSfWundETgHW9wiFq4V99s7LH7x80GNRo/yHFJ5Bc92ODyaUqO2SIRrl
+6b8+dkKoCdtdP4kyxOmRQ3mMjHcGLLj0aZ8z/WCh4D7FkMid0C7zM39cJJslVRomwMO5F37nOt1
scl1WO4RGOwD7cHZkhKDnE8OhaTHQ9t5YkcaDnYKdtxIm24lvouPXAsOKc2rx7v9rrKuRZB0LzVX
hCwuZWfTQa0HdxJ02844UTSXNUugh2lj+qpGQsMF9CZFNKj/Hg/IPqzc7mpP4I1G/hSYt2Cqf43K
sa5XmqD08qN46mUwQOK1Q981gBQsOZ0IA/1YMmIdVu/H/rrevhOJvmMW77HbeBnULapZLP9ZmsXF
0SbfEGrMw06obZIFMbnsXDP0dlJZw4geo7O/anELVgHptWM6jCPgVOmhsbrlRmd1FVXGwZ80m8NP
12LCKNiK/yDEjP/HOHL8Jjfs9vI9Q/ImRZpFpyBHW/xDPR8gbLDR2dNVNno+uEn1rQIxkLSEM2/1
tEdiNV+I+cTzt36WeUTgGY/QwHEnCYDI9EgRTSBuy05GFLiWpLOY2+Ke7tCz3DryodmbhheO4MGY
BAiSf947JrGXTH1NM82UD/gi9O1Ef9jkRwf9lv/HaXvOwnGb52vc+YGFLn5ZR6ctF+1Ti0BcT8aD
pCyZvt3cTHTMVZ7Lu5yjVIf25gdGZUvXiCNPOzCLDcWst9l4QXMdSY5fP/sr+xlmHbBLR+JDAME1
Wcg8G/zMXlVmwHW+sdjgxrmAUgHkpkvvT8W0R0FWPw+OeMqxUXXRKsF9E9bSM03Z2qKgM5VyBSwK
0+LnxM8+LqerZ3QYPXXITvP+PYlK5p4Bi/sP/aOeTYwwczEn0LtaNAbMszQyucmDCMdEnbmCgcTx
ddtzt7aIIshUIV2I6SM+kkCbxUcANE8P4uIWoXPd5yhwL4enKJbYGXqaJr2aZCXjHdkQCymVmPYA
44e09/ATL6l7rb3f28LyowLc3A/ZRc7YHQnhxendanMMSqmelacK4RDD4up1+5noVOfXYjr5Vdl1
eHqz46SzvIE2xREZiXY/mISRsNwnOGL9yQuqTTGGPpWPKfg6+fAFnFW/B0ac3V32uJfEDQd08M+u
yrsJA4+EPSb5GIarhUSgSqP827Kg5TdNg9/NER86v7T5igcdfYYnAI2neKDaP3QcA+UcA+C2G4Xc
W2yOlq5sCDjN9mpkacBxYYTXfhoTVOC7/NyPx2G8yTBBIYmEPohydP+efcSHlJHgg+Bh39Ktrfhq
Sa9teDUSpWIOUcsK2yutRUCFfV1L0eahbyqOQM+tlgSGO8t3hDukeOPp7J8ZXaSg2MZ5tpRxc9t2
R9X9nDdRLOL1lSqFbGnuihZmJp1UqtnHtErPMsGrcskfPjJrJrPHs8qhmst+6wO+iLFcQSN7dS0l
0te2CbrgH/+psO6yAArtyNiu2O4HYvTElxLjrbZKQBiuoFlsvJqA4/JDub37+fPhgVAyl8fMaBWW
5eVJYWUaX501r4WLf2PODofpgDTxzQZa6bqqSBKSWkO+lvtjZXCJj+2G8GoapBUD3EQCUQQf/GhN
dRjV30y4cM0AZAqNE1qRyBqj8VCzpKIAXVjMRKY5E3MleObS8igK5wkxoAeKBWUWIeBvoF46RDh6
Bll4G/cifpKz/ROtst3ZGHeSUoQ9ROX+KfNqYr6cp9aEOoQyW7Y6FA42PFi+XDzCs2O7FxRUj9y4
IWGJUCtJO2XZnqWjiPLNXD7lYfLtq8OjbxV7ZqG6a5ffg15bmGXRcQA5SKUIJ4G+TCyqU2zPMZbg
ZoErQy/8c8ImVBYGus7VhIFx+PQiHzifi5L2IssUOitb+lIUe5/T51v5XCehjY+t5t2lEcN51+O9
ttQxR/DRgvYkuh5iHS8Ist0ZN9hg/vqmzlrf3+HNcSlh9m/wPuLqT2hdY+R/euXD4p6yBzXJ8d/X
GCIbHenGuFaBnQrVyOup73anlEUcRba6TVMnmkZzFgk+0ElaMEB769F4PZQ3ifhTk+PrnEl7MnKa
XCJwcb5Nv72rfMnH6py472jjt1CquYkwiHGM6/HdetL8t52uIzNfaWmkFj2btA3ig0szIaEOgA4W
dfCYvxw9gHlt1UJKIG/KtGw5RAVpZFq3dD6NGU/OywnyTdeMe2AMAa4JDZ/XbwQZKmy5/Ye4Qp+l
N1c4teKFFrbPo3oXV8JEk0MsVpXxr80+WI7Zxj4Vf6d08qfno+NYOA/UPTIeUw4+japQkNeALo2y
upNLhwdfswWyH7EhDogQhFcbKZdCByYDYcn2fars5Sl2jPQev1LfoMJh0RcTaw3spBdEAWgJHuu5
nmAZElG10hYqNTC/K7sAafSne2JIUz3cCAxHwkrAqteq4edruRFtS2Wj7l1+JecwhnUmSYuOB4Du
XvqyjQUJk8eEWxwpYAbxuZbSiuB7jUPoZaJpb0F8cpOfhdl9/KHEIkbJIwBO7bqxtHUIlmO9e65M
E3rJLglwIyj+pefa8Hnec1AHMVcAO1Vfi35nUBKe/ytMsjwSbr1VZ3iQNJ9f29vN4vUU6GFt5yKI
rnJv/65yXk1UHip64Zm7uaXafayxk7+sUcVLxQB7EDRZdv84x6juNIJRsdrTvOL/ffPpLCgzGJj4
Ospd5MtmZ4nEpl3oAUK2rSg0SMJoPmGpxCrFuuQPEQk0ufDUQgb9j12wF3F02e+t6wBwpUwFY8eD
iLFnt7SY3rrPs8vt8yIX968RGpwAtcBOcj9me+g1DwHhMytgMGbB2M4GYhssEBNueb9MplvDXnib
12hdEH+Vx2wwJCSFnkFpFxIhWIsBRbEGrq0xMLFJ8/V1yR0luW6lEF1f17+/TKWyOI3Ikhv82Bx8
ZYYe+ZxvFKVPBGmTxbxR01Dy6QnqLtclie9WJ/6uKlvTqOSZtxBapPxGYBjaicmzf69csgKgoshj
gq/H36QFr1yiTBhkWd1wZDU3AvTa/Ee/8UHYJmbkFf2ws88L0G7L5pR8IvaTQhWRSvR++xx5pLC4
hLueL3lUPxDVtzh5jsUXEhZmT0jr1X0Z34vOt1wFyIeiMyLR2dcHJh2dW3t4bD89WxtCoVKdtbSv
48DmUPa++eeG6S6xBoLSzIkQMHjedoMdocO+/5sYDR8MALxxTvPnBJ0+XTZRrz6Mhv11u+KOSOJA
SzBHlSfbwOc1Vi8af6asveduh6pzH00xM+HoLqO7XGfBhhHmNl7VCCOGAwHWCxNNyQrSC6mLXqqv
ZiLW6WIMno70IxMqlx8KaIvmxv5EhlwAHFv6H2DMqUwTfQaxjLBBY4yyUCDGq9IA081LyUe9gvW9
NXk5wxY2sHm+rHwikAPVGXPF5+51sSBGn0+51Q+YtivzEtiWELBP0omJDW7gEz3Tj9eqYih2yflL
oTf/wM3dlW8A/U9vzOJU7tbrPuk8yz26Xkvr/M+GYCV8cVP6XgGkkgUSII0QEuIMQMycMNI1jk4g
0bRETJygvFnYHu9NBRlcPi8q+MSIbFTwOXunWNvQLzXDlIjNU0Y7YURdCKK7fkJ/9+YlJlKke7OX
3lPfymRgr3W5KWdoGTpGPkLxh7/Ne43kJg8r34RaS5th8gSHoYI6TqedF4SypDkdQp8iKSy9YEeX
EKXdWmj3+SD2klpnQPoh+e2rTB3V+J2sbxFpiDQsZkHDYyOGri4SgoUedldRaH27mfK3v/+yNv0c
Be8Aqe5UCpsudQbHBI4oNvfGNkdTx+nYqnoDGbUHalWcK+7DQEVj8yBS/6biocpAjblhRbKDiJ8B
gXEfmbVqRneN/QTXKdFewoWvN5Qy+z9/T66jT0jPDWrIIzunTmh0sBXSW0SkzFAdsZ+wwYcUeuUI
eL7VuKRmdJdjf7qL0pjf6XLIIi7h6ohKBEvn7rGfhjSQ3Pnp+d9K9LQWabfY7VnAtPXGCdsuAdjM
aWS4GjzKuRdLWepH3a3db5UCfVhu99cchn32tAu5Ia6Af2ZkVI4K7WLaotvkwnJusxiwboVnRNeN
NGq9fbPpBxus6wB3QoQbrmwaR5bsY5a5flGimQq4BErXYcZwkqbgSOhYD5uzDpaG9g3MDUQou3Qm
SzHxrK3JqUPuY1HA32+/AlLK1te1+zkxneiikCQtcTvwS5ehOsym4cE2pZGg/17ZXJLyvzcvx21M
UK83Tmb1KhflmpLoWVVO7yEX414CIAv5xmvENOFy9an4mX/Brm7wtXoPFKAit7+beyGdEiFvuaIp
RY38IY4i+0oxM4ezZdsMr39HO0Jf12OmXqmLryaLNKqsJWY/qi/FakHY2w2XXFozdT815MXfybR/
pOTbEC3KlxGu9vI0zbyMTtGMloqChdZsBiDZCNN1plB79+sPZGC4vLpnwUsxhoinzfHramY1tEsS
YKJLC0jzOrenKrvnHUz4mDPJmCvgG80G8WnaY9sgPuI/Wck1wSPMFVgPj1TG6nohGFhHPw/gTi72
AE97r2IByFcXkHvaR8mp52Dz7qktUlDWmea+AJnvPZSdc0o4k7VyTtiCaofQrHTX0LWJ4cRIXYU0
Zj7VJOgrYLMIf96r7wqCgHihjX3fFvYuzimC5V/XpXiDpVMDSY9dxsq5GcOKDumIz+gIVuLUs1oG
TEi5rUjSuHpcO/v1w1utTIxwjCvGKv60/SRw5RMnkIXFL315nYZXWj+XFG1T0lSFMEev4Dm+3GRb
aiBVXhxMUADKY8JTNIikcMHjIwPMW6eZ4hZMScZ7eDCSenzwGVfd+8GwkHidRXUU8jAdoK8JpK/x
g62OeakLEzKcNbjp0xoUaEfwq8jED5URFAekDQ5xZaqP0yWSi5dmxCCkGcqBwKLcO/rzYPkntvgU
c2BSt1j1DgqgFwRwB9I9vBfgb3KIiHY7cDcVPkPNYbuMTtCU21etWwvvhYBVbfy4r8MZ3eCLw2s4
0shGU9zTuuZyWNcoNs2S6uwWx+Bpyp+zNS/Xs1FJQcljBeXPMoIivOHbHCzMfBmNSU2m0gatuv1p
AT3D7+DQvlMybfXEyaEsoSoXTCg2hNfX+zltyx84R5pXhuXBK/v39nbMCPxamlj6/Tm2dlQZ4zDJ
CL4qFIFBYVrU5Mpmw55G2Kg/P3nIrKfBcP+DIByL9Ehnh8tSaqm91RTO7Py+pybgrobwIjz7OP6O
4I1GSu1rZDY2hJGerizgpuG+Xs2iZ6DDZZZvlqZRGmKH/UGyQVCAYZ7OMckr3NmawbIRYdaGwCR6
yXgFhOBDl/41tmWA0G0y+35zIFfNBg25upJlVvZnRgn/GNqvLNbmTJtgHjXubkVOEINf/3+vuPuN
ao6p4+6dVE8ZeAW+3LQ/UjMqq8IJovUDHzxAaGuwLYhaYZjTyoge0xMTZTnlyaDKyHPi/dC4c9tX
5SfkaU7mYBC05+u5n4pimDyAD+4Wt9jJ3qis4rPb93ucSZs++QBZCwMXNEZH9wSR703kg7iC7QRQ
Prz/o0zpEQf9lFeHTGtz+ZYptCVDXNaZa0o67/+HB2N9UjOe38tFjKp+qeDMoovPL5x1c/DCJQNn
XY5/DJgtgvMgAq+d93BxioBYrpZ7jB52yUrCVWI+7/igy59tMOCrmJEq7rOIcrXs+KJ+tofnH7Zd
QzejD7d5tXovub6o2Bfe22dbM2FVPGHNox+T8L8jLwpeV2rSn8sjMReVIO0HCdZb9+zCnxMgYW3d
iCcEgB3ekJDvd5eitso9TXCOwUyLlTIi5oB+aCqdI8Tai7cjufZeoU4h3riNJfQs5N0GqIBmkt0Z
lfw5VTaGqawjeHOn9f/2/hgyno3+sYJ/eir2VSrfrIqrjQBWjzhbS80qJ1artLb1vf3vQ2xcOZPR
tW6LWL/Ce6fVmnWRD4aw6oo7E2O6QiqYGp2JbOehUSKQIXRgJ1E1N5AVgEr04LR/mclhDynX9/52
Ch1JvWWkOsUZbiVVrPbqOFWAci1dUKyNlHVn8165clM7DDrtETwXNAX3LKm7wIXmrlzSOsDOh9f+
sM+mtQ0J54W5XGU4XongURflFqNs8+t0NsWJL4J36cUq+Ff5pLfU69iUrp1Ub5GuF4cYcoYXo43J
/2bqyAeJ8GfpIgPCyu69fG4Fh6E6eMuuPNhUcHv1lL0kJ0LZq5ku6d2wXApwYJliabGCGuExgbfC
gEV1Kqdtv5AP9GDpyYOfubRLVc/uVIBxT+s6nwfk7vxE7LiSG6EBl6Vmi/CWtkbNFFvro6thKPll
uOHCE1F7BWNYkHy7LW4Jbez9kaSPTnAs1c1WPrIxd3MDoo0LI7rBOVcxHm+X2INPvc36HcnybbNP
az/1QB8rJ1hWjK9OvHDyg/Aq3TK17JjX+5PNxleTAU+c/LG31JUBx0SlGGWv74ytdvK6RL9PkXY1
XTQktDOBt+9mmSYN06cNL+5djVXAUGlXbbsf2pE/DmvylyUJiOEH9SOXJ/XCyzStWhIbD/0kKPlE
XvPWDzSPT3yePuuSOnaqumZPCnTTbvbyqVtnc+cUy3qA5BSoybN0G54+bJm1LpUhIqQrnwY1zb/a
7V0nVCwCcSPEnMuP7f0Mk5WtG5uXfcItoHWiSwVWfeDGQzt5/K2OwaphlTkSqe2FgNZ0xaKcCMxA
+VO61WeVcHpmuG5Z5Cx/n9WLtgAhuT97EJU6NrETG2oW9x5j6sBx1SF2QhL1ivVS7RfOreq+JgBl
ZeMzCwPrebJO/uRUVWZ4LCOLudYBvrldNllrTWekEei0p165Cvl+/yqKJibS+Y7Kr/PTZ2HfeTkw
T+3T+ZOVJl+/T8eGG294wVWyayJziEHj1fNKmJUNbTm+SF87fvsAqP+gQPjfxmLFQ60aeQk0ufHJ
tQIgPSuVNJPsXmkcp8lm8RDIpCrCQsxgcuKBWz9qXkHATw1l/sZsC+l2iAX+FnM5KcsG55q3cVjz
5rLIfDlWozwZrizyaSNQnmvFSu+nYNb7fFM5Pd5iCR9HLM61GVXzAHmBKccWbeY8bbyIsN45D1R1
Zxz2HaUJNYSRM1BNlx7tQ16eiW3btzJTEfLPWQCdmk0Klx7CQB5XqZTrGLLGsEqu2TksOosFQGIt
x129q6m09X/XIRXbUtMU1RwZfmXK9FkTbzRVWpX6a9QcUOyw//pHOUkrOBHMSjUgHIZ1mD/qNiYy
m/OSRr2hQeWQ8ZmBPJqs8bxt+cDjt2Uo129tjWfzy5JPvdFyLbnD6TdMwz4Qj6x1RVnClsRPZjjV
0Hq/QWdGnw8FsF8/UT6Lb2ivGmBFmbpXtWXNwbGy9ZdJ0Za3xm/RoLOHd11QrJnOa58nLPdL5sJF
FcerLG5EvZWWLA8SR8ukzjcAnMYYJiLY73BGPmWoPrAJSuAWIGDCGLtzN9zeW/oIouOO/53l9MgF
e3cJCbxx6Avd2hv9PDkJPqb6rwMs8jrbAjlf6uGejcMd8fT9+vcN+nbvhPBd09Mdc80gstXOfL7F
yt3pcdTuGLZes64pKsne2o4GTGmv3JjHW0J2BvlPbrJXry/bf5vpn+rDtPrM+aGLZoLsOcfx7z6u
zDOmaNvKC4WF6O1Z8pXHu2mSoXFPayPOPNVcWkLm8uF9YzTBiEWhw+k5iR0sU5Bdm63TXIGlywQq
UqeM6ZxhzyQCJ5fNErHgcxgHaDQCDyTkLrohQ/YiKVg0pu9FxUdahny9z7g7wBz5lJnsews9s+Vp
BE4jp0spHzWd3A++MRTT23OxITKX1fuojMApHtE76vQM2rDv4fzKtvHPgu2uY35kzbmB6Iftacf2
yeHLGZz/55XYJ6MC48daUh/x645CrJ42i450gTbLo7/81heu1V6y6bfHtyOaN1cr4URZfzh5TjyD
JsqaqCHTgXhYZreZBmeSCa1T/meOiy7sb1RbvYFEGA/FBS7NyRHTWBNjJGPfKpW2+37Wm8U51cjP
6Z8tgQtAPnO6fD3d0s+udGTzx4h8ssLJA/6jsb3PDg01pSrxYZmDUOpWND7d+uxLwG+7yXPNuodn
ryPig8H7DHl/1X8omK0iBovUkNE2Ft5zCz6KB2iO+9VLn5pGnJxZS5AihvecO5wEZzIlCe67qUkz
ZcL4FvB41QVjInBDFpokLT/qf2TcI+WhGgIVT7tjFxpM0sbWtqsPc1N/vk8yAPTFVCp9CbhehsvU
Ip+6oxoIzU25U4khWDuaJo+dTLWCUDb2iI9QOwJPexkMFh8kUP9cpZaZGEwbAHAY4TakELvZiusa
WPPEsO+M5rxD2BKJ+k/kYxWwPPgDSUCpKE7q+9k058UTQgPH8sCXTajaZnsCBGxIa4M4TJB8CdEX
+Yd89nGDjEiUgu1OoUOLBT92EiILtpgcf7dwZ/bg4sJNIrppdh9vekCjQlL2+dVJ/TCllMKdogO1
WV+ZJ/X9RQWW8IKq68jXEMb/CL1LoRBtO0DUHmyLNnTJx2EZhkf1RIrOZfN8baZl9mnIuC92lWyz
tm9+4gyR0Wl3zlz2flJv5FWSd3wohuHu5e/FWWyr07X4FlaRtIPZANxvUysTPXn0ekGQJ2pnnRMF
Qhk44KMJLwCMzS5aO0Xu8riJUuK39IlbSdho2/GnmSnFDmTFA/Gj6bTPvoUv4MhIHxsiYBV9HKJM
m9wUBghs1mxpkm3XY0ySzRONXkF9eTWCdbKynV5iH4vhiB+G40eNWW1/twyWrbakNm/6NYYeBcNN
EaQCCx88g3kdbt2USfch1XSGG6S0DcQ6B1+J+qMQzo2+uB+SmlV4R087FKlQX3rgVPH8I068IjZs
euurgfbtk6hFwhVZGMKO2Waw9pB86sz6F7tju2s2Jh06WaYzfCJAp/9vDK4tWZzFGfXrQ0lwMDBv
uKYlpBtUUKjBAaB/Zwj9Ks3PcNvwnTvV34cVVaq/WCg81Jq2gZ3zMLv5RRD+9b+7t7cwPX/VkJwZ
rCDde42wevlEuldnX8MLyyyjun535W3A4mWH8O0Oa3Xvd6G8ehGcIwrtRzK/Zm0rRwDtRP/Z1H0y
RkRvZdIMpacQ0ySNjfaCEDC6UMr5ClOGlY6CzB0ONBMXg9B6ZG6jlLCw/YJlKHltuiNkLTXjFjO0
LRBCK1CqX3By1OI9aTo6DgneX31uPFty6EjcjOeWAkdH8ShbZug/rHaPDd97TinHZjrHh2/Ugx/Y
07nFdq94lVYOULs1ezXxfH9UkvCljprT9jK8hqZM/pFYQRUiakLMBf6Tp/kyuLJJmwko6eOgBfEn
aPb6LHWxM0I60lSSG+anRf45xrGu8LtLDkyFyTFcA/7524HfrjlkpDik/qqzZyYX/9X/Q3gJLVwl
3VJQe6rwSH3txPXRz8OCcXYHCCcF1NKXDG3fWGIsn7Yy91PYkqvSuaLPbZ/e6Bvxe4S9RawRgDL8
cHJsBKfpNCigGvIEs9jF0P9fU1WbnKcOr6cBlPn8DcHxVmWePiO+a43hbxjYT5k1N4SfQxIJk6na
aVEWYmASKFOJFOew0sxMrSMK8XTTTuepCOpkhD0zADsVPSbsRLwFIHw4zuPxz3ZMBKrkLIUBXScs
muRsKm9UxWS1ss2veekF2jX9fE2Zgr6SaF6eJBmij4dlBtKPC2iUZIhRptqG74w1AAgNrT0NxVrh
2qihTnWX95J/jmCeYkON87Hcqow1EvFDh0Mtfb3dDTMqdRVDym+itPJv71Vpfbp3etgiT4Kd41af
GKBn6BUL+AiVuq4NMtXG8CrH9nMRMVUohvqWvpDnlSu5qmigyiXhniesiT/lJTc23YX9FZ/qz1Of
dkgwYjDcE2jwp/9U8IBjc+ftmlP8l6yfl/FAetfEzwHhHWWakyunTH0HuXt40GzdB0cHh7nO8gJJ
HBa/bBfadIp7IuNFkarrrEoWjnVrKhXS1oxlTwsXYxyrmqlgns3woAJOPnDb0JLKpa/OS1O48+yr
C5KcjWs+2fRh2AM+IJJ3nob3sJzOn2VZT4NcpQp6VQOVvXOmPw9vXd23jqbvVywmC22tVvGmKm5b
S7gAV9uz7LF2fMGJaLodBM04JSnBUmQyHhJh+UdVWLulZYO6rB/nZ7qpRqlJVN0HPQ9lQTXTTLTh
fovItYNJ62Ceha1Jt+SBIKGdRjd/tT9Tz/dBw46tZ8J75SEG5mNc6CjneOOIuIgf4kcgZW+uuq6C
dewy5f7AiXsQ7rO+1OVaLBPLfVgfSSMchTSzgPFlyd1yCkIsKOWJ/zi99CJWQvgwDmvYFEZ+X/nG
ilaqd79Qv2Qjz3XF4ofcmG5PQ+oRwQe4wPLkYQZGMqtmDbc+W0UlaLUyNAuw+15I1qrwqnzN/JKT
fjdKq7onqNhp7JPJRfDq6pskmni6rV4knzN3PlPzrjkFVm+W/LbZ3u7RPe/q7QYFYvKFYXZpVsdc
PXjwDQ4lfFIsSl41GomG1Rkp5JEnOoHqpYsBETm9K9B+gvK9HA9GaoZJMC7LpYSaO/djjfZ0kKDF
2BbLRK9W0hBCgEQtvYUhtBkBQtNQn5NIDQCOdl/hFMpuHg6ENQcXnySuE4I/RQtmmVuu6LLjE65A
knrVHkSPEJGwNYjTFuUT63aJJWzPGKMTM6vsG+QhWzkI234ZKnRqpROFuNEvN2Ms8zqHEPvs4Mox
SUToew9a/9ZKdz6NMhsvc47MBO6HHnXBeqP0fzAn7u38TpMddHAA53q03VrRrmL5EKk17zGpAyU4
pZHpG6/hKS5GqKORQNX4ph/U8XNweaLtZ8GUsDtfd9lmXYanH1gcwvc/ytPg30zDC/1iymTBR92I
usM1cH5eHJZ876I2W8MfbYQKYTwW9gwocXKcHYFu0WopfW2CPII42Qbwp7zzQOrdyy1A9WBKVudy
j4LZP/sEsN5GEh2ra6QtFRur2MGKmxzctfHjYHT55NntsOrj0gER5M9qPzzckcMN5tdR0MDiWQvO
R13xTLWBF0IfRzB7XTagIvM96+HzN8YlIxogrRR2cn6x1idGLM68d/M/oQYuiJATPe4ktOf1yxLJ
od3x90BUI+0L4Gj8RdwiLEuWEqMYKvgStswjsHiOgQ8VW6oegr5JXtVqfwPEA28bzGpiCCYoD7Z0
9cIOm94puucnUCB0ueusgIsDm6v3gMlX85FxyA+wbR13q1zd+Mvi/eUQzS4SP+6ubVc3QafIsMCc
suUZVQEd/vPxJ7Oej9uyNwaqq0XmWKxJofBDK3UeEi3+W5i8FHvdOlNWUezDILFEY8yErmpzaP4G
lemnq/cfk0HOmoOrRUpLHgleji6Y2XrviohHM4GvNkwGDs4WBhoXHaTeojgZom78iiJlJGlbZ1vO
D0/bm35SLLKJ9Anw9JHEKt+ZaFzjIxSM1RGt1OQG9SIxNl+OOoQyAt1DhTBQVxqqNE3bgTGvjxEL
vFa514wUcy4OKMZy5nivAtdq72mgbz/GNL+NSUOn/uTkZ6TUcSkbreDH6CCSpsppgIOqiZ6h+Zyq
XzmtkCNw8uYactP6gg/Bixbx7fASbgbxuog9l4ROOfgWF3uOU7lkePKa9mNjkAJ0iv5CACcXy2oV
TYyz8FK04YK4sOO+X7s6IcadACgoTmKUgYo8pwYiOGy3YmRtGoCt51qxmflFnKLD5KImaqHTMxTi
i+uK7rmeu/ttGRn18GBfqB9PsyR2Kn2AsIh6FQ4vxgUe3ZiO2fJ3bIidAp06iflrCnbR+SZF4AuK
BMIVGPnRZEYxSz8yhV5gzC5HammY41hQYw2fNCmCPmu4WvSfzB0Y2NgCtOckj5F+O//BssF0wZKv
Mw3EKCBoWmfkbsoziMYzTjUvi9eFQ2nYXfrYO5PaVSOPRLY9TxIHlYj/IGDB0iSSemBm0KisiPZW
BcEk4TsFTMZJjKZCBMdD1IWw38EBTGuI6bPkH46zv7G+DxI4PogG5kRFmRwmmfdFhLenZ77ncMYL
px36TYPtCT26zUMCi3Ba3y9+Cz8ENuvQxq+L+TEOpR0Qyph62BZFI3LNqI+kV7a1VgEn8yQUbSS7
mK7uRvZRSAOHujvlc7bsWwdhdGjG9O/GFIr5YZVCTryHwsGtd2yqFmv0jdBNoqrN4CEthJ+BkTRI
QSCklZV3gKkY2rED8EBZe8q43LJTC8XmNwqJzUop3DmxIq77SUgX6zClF4YN2hYZXY/B6300Vkje
BeBlWB5YvNrNrY8rL8pZnjtvhKiTfBeV7liMkeh3Nx8/xyyhoUIo5R9tlmgIbiOdMm3hQQbp4bYf
ZZdMUSAPX3bgXEGS92e0ULCX8miomRZH/E73oN47NwxryYrl9BKnYbpJekWiQejYTfpjCpXfmAQ/
rEtB7gN4QCpe3RnbqIlBrQNidMNqcFBM3AEHljDxa9B9fJ03/meSiolGC8Kg8GpuIGL7t55Iamxn
rAPtAfJwFiThXXoVrEwzaco5oYOeY+DbCza2CUIQxgve5nqJc5jZ/yIRIzhHCVoMegoC6TVT3maY
1nNoHJhd5aLfuXyHYfWcz5zCZiovitHoBJx4coRTXD2GqnAUdTs7jKKlroso7IaW1PJTcG6Htk9p
p9LIbBsiuSYvWmRDHzyxo0uP/4Z4tcsqm0EvqAxBLIeBzd+1+ktKxeXGOG6qgZ/fjR9HTXiPOKcn
K0x50DzWQzGgA0gKrUS8239PTGDAproGmVzuNv8xNXelBuovI+dmPzQ/PaKjMdAmUWvJm7aC4aq3
8gf1/awEKpAjxTJLFKVquu3kAx/F7Ser3bUcjUVnJRHj1gTPAPgLQEVKQBsSC5Anih9UCMUQT8uJ
jxoMA+vTK/gLuCovKRFazwcXWvka6Ycv5deL8009BPp9wY/oDHjYGkC6NEr2cWVTSnZA2uLHQZBu
U3JkMQzdH8mNamg7Xwq2i2nhsQCf0FSAqhhMD1hwT+rimzlan63oRh8HbQfHSzBWVGPcu9oUACJ/
vxSd/w8pzpZoBAxs7O/qDzZxG4F+iCXq+6HXYHQb/uHU3KDy3210S1LfW/EzfgTcTSqQ9cqr07up
p3FuLsVWNwme7WldUjiLC98tCzkfVrKkoicqeKgFun1fbsekJKyMIcTOftUFeUVoi+xEpacfalCY
NNklKxcZ24mtPZkxhf8CXosnI4WHqpcjB6ZVVbQSSsdUHU7OhTdGSgY9qvPoGdtEyWKZyHWcQ8fh
E2wlrB3mYo1DEijDrv3vv3PdiwTza+JI1LUlANdavwJzlldRyDY82fj7YQFqktit7pQ9Y15O/BIf
O/Ns7LYiRaLwVVlfWLjOtol3HJ9JSLSCxuoMNkDUmNe1v2B4rOeDh3i8+yxjXtdXysbtiv0zqzx6
gHpLX8fplYNWJNYt24t2IECPhJR2069oAORJn1KqJlkfcBKiJVVcfD0n6or/GsUYb8rWhcFJD/NU
KlFx3WcQ95LbXopQRd0UKB7PZlZ7sT8lULLO7WagW0ivoblrR1LTY8pVKUN8wQKtgeBnuzUCVQ/Y
Sq1s2y7K3ttQcalNR2DZu8Az+c1KhjnHO4lUtqdxShVwIczseQ/zenEmR/4Awqw3MyMouqEJF3Zv
c2hZ62mYEoXzgAaW9T33IPOMe/MF+vjdyuDoqYQzz8Jh0sfMgJfDYsQ5DG2V9Syyo8PVmjsDmx4z
BZH1/jpt15FNxUJxKrFwmo+4HPvoUWtaVXdtNRGgzdT5s10pMFxF1VORUIjLozC59w3kQ4rKb3s5
UUZHJdMMl89cC2MT1p/gYVQK54fC6sc979GSyViX5RvS7XRkbOjs2YAO/JJEAE5Z+sOAnTM1iCK6
9lnycx9/Og9KjzhfmlEGyRZZggic+W6yJaTg3AmRmySio326G1INxMmlwGzaJnYLizq7LFHxKy/p
9BYX/5+fRjFi7s0fYgyjnEwDeu6xwKijINNmg5N5P6ITLjGWvSabq/DSmvAZVWlM22CI5Kvju73y
+H2u2f5A7c3MEG4wLFwIPfi4PZ9eOSk8b0OpWrcu/nLYQH/RtIotb4Qe6+RPOSr+KiQYBomcThyj
Zr5mo92nh2E1csHF5whXfuKMsiPcWibVNaGoDnpzvYQ17LyKqhX1Iq5QqlNnyKZ93CI62foRNNmt
gYbWLN5O850gikpETo3o9yZQ887uSX1GgZb5NvrMd7fUwKTgLGhHITS3YWFh6rkup7V1kUjnvpw/
DFEF1mHlNLlo1rFG9o0eJvkyho0TRdYkvsbr2p1fW5gNi6+odI2WJXh9tooUakrYmDX+n2VNOU51
s/iRX64F5pZRrCMx/JljnbrI4adNp5FshIjD4Ccdt4Oe+CRyHjOOcQjlmMxr2p0+UstJICf9FWCU
3TXLb7DhyIbrgyR76SiB94bVpBl3vnvI7cqY9UXE/a5IaDrYFEAZP7ovpq5iFwg2gz4nU1Fyp6IF
wa5aQnLxyeuPWhpn6/RQLugrJQQObOLLcaB2po9jc4B+udpHl8MMdm1tkMsKx3je52KFsnokiOD+
VY76FG30gclX5olhiIpDCV1/F/LJCl4fJi2nAIh82Y9La2WVPxwmvnEEQg5beKO2rTJqGShXhG7/
abRjGLk+Lld1Wy6AIV0p7oVH16uYzJ+zfDiJA6m89RrLqnQ9ZrNQmOpewGD9mRnSV4T9sFhzRnlk
iDMMMnnC+iiZvQl1MPIe5S5nkQgtuJGpuuCIvLEE9rQd7O2Blr/9YYqw7iTenivUy9ZOLJTTp6Re
UFFRmKwRFYfLQBYaiqo6EBXe6iujip00ike3v58jGoQLhWnX9Mz8pW0Oh2F3kIwS94RygwzHV+hV
13SC9lhKQ9w11MUCRcei1oaS5d6VO5fSITgOt7ylOPAikBFgCtjpw1Ky5KHcp4gd/uAnzIO6Kd+X
H1XOPQOyjh9hjFhy1PGn45bEzljrOExzaxYbLxCLQl2+eT3HhpwsbhjPAXhbHhOr2eQyPczaOfUH
mi2S9VSIiwI+438656Aiokx/1gYqX3bZ4wtcJLP0+SpppeY/yQ9uACa7dDIC0o7mAp1PIseyftDf
pwwViLkFGKxzJDHcLy5Q2/a4VF4cV1V+0E6FGgZLBG9NyG60QXuvzGy/GhV7CFSuVO8jCwVgMjh9
UrUqXnCWlSXzW2SUNnJQzeFMtAtklLxx5muFbcTgy+6/Ni+I95FFAXbbXOTBvqa7xfncJoxJxCHC
7Jd/Ph0LXRQZKOyvNBZh/ZSgMy/rl8RpStdOfL3h1LZQzq03IASA2ki1AGCSbNYMlR5o3zo5Cmmo
7d8Z+c/m5ZUjY6TBBhp+22qtzFK29PAvS/IyZh33689QcrZ2MHsZT4T85IVuc9NEG0SqOURieDQe
WAj9CoPSh6UXGQ5riVzJ/LANzlNlnRbTp7PNapjBIrTm7+mOT1l412//B+ssuqLvR6uIThjdq6aB
Mpwu6/p791cu7LeaNd0FoRlGN0lmlh7GkTe7oi25842u9P09Owc934CH0aroeFrV2KjdAtc/yhTE
dmAzBkmptG5qczHLmxpM+wVsKETs1UrBSFeifWHMTGTvkzFlFkupumfYx9J83iS50hEhIzJfV4mA
HRMkzXM5RG0LXaQTzqZ5EjT9PDQmX/svQtxqaFuTbqNePVTVyV/2tCs9tsHnEwtCeIyRqYrP22eU
mxf/pxfpcoWJI6HLXJGN122wNskGC9ceCC2RDs2SOlNRgDtiDiJNaLBx6BFafnyFS8YmoZ3M51O5
lOV7Zz3qprCgfGIi6/dsxGUmd2z2C5dyg5PhxFt7m7BKWHIQh8M+WJxfDh97q6brna1Ym3AFAG4x
EzsY92LTzmBqt87Fddl4MXYpZQxhzG7jw22SZgy/qPV0gAHQ5r/PqpQaNDiz9VXGeZoxI0P9cGUu
duczYYnGssXLC7jyKrBSVCDEgJCa5wNkeW37Y7Hub6Da+npx7U9GqyMP0olEq7z7JTz9zH1xmn6f
iNMQ7LQ0ueP6BRfJZU0IprdmxhepO+bS3CflSOEobLKHaPDzu4LVbgKxSSbzia5MkZaazqKjih7w
GlP69SX8PQ6siQPaN9X2YbK0xwvyRHqAibrgvCXGOd7uELOV7qI6jBF18l7S4bRpVPhXomBHVRsO
Tdsa8zl7gXXIKYeC6OrubEZX618gHuTo5yZBmoVMCdxBGJFRxuplBvtxKA67QqMNQFkpcPuDwbz1
vh3IBJGD2j1pNKOGp2hbQblF9cncbMk3o/tJgNFER0Hsjvtt6QUoUT9MV1yyv+SlBqpT96VP+rbd
xuVWEJSA1I+sJ9DcxBvgEYFw8zT3OeEDht4HMGWGkBnXVWNxd6zK3zgSibCiRQtLVJ8C3/WexRzU
ywNqqIfVtF6xIt80yJx2UiAHkeupW8f33OPk8JMl99pBk2JmK87KyWXeoIkS79kaxUWPeqMLjx0d
qvHyLQqjd/0TMn4Vc3oQ5YsVZn6gNvIMQEZznpUk0A9hceanN62sJIIhIxgSTqwoKmUatFXhklaw
Hv5dyeqhF/zt1eDozk2ZLxlxKtlluOcxUfodf7J4utxK6JQtKxaLMnbwrdJx8yQrMJV0PGeENQXw
vv6qWTIcHKTnS34QoqOZMmQYwexwICo8Cwy4SjB3b6IUu5JgQigHTz92/nnlqLw4fyorxMjvkDly
iZfraXEN2xrmWCbd3AWjWSw+IhIGk5Ylo7vpt4snHg7/PyG4Fku1/yybLbJFcWiCOd9okhkcqIKC
y5K5d3UERItNK0kNvlsSCo+t/RAtCidiYalJBsZ0ZZbzqcz66y3ICnsFhQV4VsZPefsxTvLbnou0
LA7DN10UePBNwXov3HitefPZlA7aKAc+guwqLwqnuPnfxKW4Jd8oz1PpgXmh2kA8L4GL+QKbmr+1
uGmr+lqp4ic7cq+a6cyObvWmX7E9JAEmh8r82jbar/A/KEAHHJxr3qQi60lY9RSZxBsTJ/+Ozr1n
bqBlxK7bHQ5mTNxYUbZ2apml5KQWC3l7QqQNJLzeUzLKQjCVC8I0uzoRu3uFQgws/F6PQTS7PjdQ
6I0GLImwXn0+6g2cEI7Sb5SaDzJuDgx8n9tjYYGCGKxJVThbytWdgsDrutnWdJjr9t0Dr5xzk3oN
JH3eVbx3AUi6KBqk5xtBo0wtwB3mQvBuaWrjafWKPogGw7GpqCo+zRh8ojP5jy+kXbIonBtZWGCR
LbsetQokNiaRpg3/vNKNCA7Kb5Jse5z3hIYbSBuh9nhq/9RD09XUqgem//5ZziJgWyMtQCD35snh
ObO3LXGKrQ8Z8+gpNLL2JY0Eqxcp64kg0RZTPWpFJV6d4pKv4EjQwfbTTCC3WseQU0Jn9nfRj6Z7
JNA+Z42jPHjlAkQHUlxRUbrYWSw5YFvuckaTx6hIKkM4HJLtyQq8mg4lYcBoYDUO4fBMAWMHbFI3
zbhL6ulf30RHO/x5Nd98A6yK+UEKXo3VlS3yypCaOGnm5BvX7CxxClrFzK6BD978vCGU6h7scbo2
v0qvyPmWM2UUejApalaVXgv5zIFdjmb33oUlc0NpzlZtUfPT+HbzRW0kqbuMWrGCdGwP1J6h++Tz
zmxGLtsoyxBhUi2yi4Cf9dt8ZbOc/BQSiqbG3w9jPQUegZV33iex4SZh6jB+8xh4Pwx9XfjCzfxc
dOmV2xYR2KiT+KaA9iroiVvmQJZ2HAIXUTo1AAGLWinBu1kdaXCddyBZoKdBPSJ5s8u8dN726sHm
lOBNkihlRdzdo5fRW4+qQi1oZIN9zAnN4wCykFEHGRIBSLrp1yLjCCDwBuZi1GRY7xc4ISZNC2JN
FbVxQuiVPOVntRcTyjvFsJHZt0xTEWz051uH4hAZHtpoFatxI9e3F9eTQUHOlo4CS9cKj5oY1lZe
OLPr58ZzGoy7DN7jdjfgCfIxihp93d6brZjbYI/1S3Z2J0SE+3ecwrc+cgqKSEBcP0GC1XqDxvKZ
7vPFfD7UgMrKZOVGRMZl4OOEOmjFm8aJFTXxIukjrxpzyJGWezIFGl60y/eXwaA3lrj9MtkyT204
wvP1DNbJ6wBmc45qQo44XacKEJE5mlsLTsYOMdmFE18koJV0275U2GaK7UFWXp4FAqKnxYFxob9E
x9+HOTQJVRAlbg9/+123kTYWFTINmUfSw4DwS/yCzH9vwSKVthX3qW4QKzwpuGX31AISQOemphdM
Nww7d5j/l7bJcPCbGabL5StaTdei3zgwHWn1U/PppCp8l6dot7f6r5Upx5uYQX6Cte7+HQwixhBZ
LDD06L3V7JtEXVa7zH5+RPAiO+CvymPBhcRcBx5CPqA/arHzQt9yLecy9eWnBWU/HewRBJ7FlJ9x
mC2bxjjFKJA05r7KcuoNdUAzKUlX0jhGGUQJHTx7HxEgGSaseL/XhgvxiHXke2s9W6OcJ9ch/VFG
L+aGBI0IdykgQCz+imFUqablEN5WXoP02h+2YKRtlw7ZsazJZCltygtyWv/tLnhbUvYWLwZzhqLz
9GIPyGw+iAiqVTQ7oaKQzwQDGk3gDPlgyFasa+atikO2LVIwK0mAyVPWk5CEHn3EatOje0tQa6wI
7peei9v8tF/twzJDt2Bq2hAPYkfXei/8ygecvn03lOfJ3lblSoOa//iGVkCCsaKSSExNpJ8BjZQa
CC4SfDrFGH1x9afQExyb2O0sotIw49sa72dOBINZX+G60cbu62IEREjlSAtoEcWT/lTUEbq3bKUe
4QU5EGIrU/RszxLrvOPeSiHSYWBsg65a91WDM3UeNc6+RB3gJYKFlKHt1lp25ikDoGTvj8VBX21v
dylGDabJT8M8xAU8SK/Ns2s7FHpMODZquOWjFtodr3DiFC719yUaSZseiz1o0cDDYzVoqg0YnGNx
ku0ZZBonn/clUzirJ4+Fe3UPc71sKlONPjj30XEXw3WbonDWPIiwhHSw0IX07UEA5KduGqTqzhTr
3rKJWNnSd6CF9n6CNoO0zyGD0j66LtRLDqG4bpGQV3aDIrBASS+2GTOulyGjnzX2e6TokOAHisWp
duOFX/bmknf4E13JjQ+jpaJNOuZlmsrfqhkp9/RFZ/pBsIHq14ZGS+Cv6CCcGJuaUlDE2yB1Ao3d
Y8j6kswieHaGd2kjhGto1GNVYBORf5kZthRG0Mw8khMYqiv3dKwS9LWaF0ThTh0ehmOhYiF3Zq10
lrjw6rD6FizoTqRhVXgTgJqwpV9Lq5Qb8kehc3eqmunbEDJvOSeb9WxiKcZjtoISZpv+CV9WNaT3
wHemjOailQinVMpNBXIhnrxAh5J+HhFcYcJpg+RZWgqhmwdgDpJIsmHwnlj4/tKilwGrSpdQkgkK
oc0f5mrhNYbdbJqAumVrj5UjYdsZ5nXgHLE0HpvHnI66j00uXGpmEdTne6waiz8eGvBr6CQF5hxL
dISUJ1YQEW+x/uLyNtaoXDH4cOeXIZPb5EO7ZMCslJUqRvC8XGxDWKbeysjoWBFHY2BOjgRtm/rm
e6EyxWumvCaWPtoUVtD2NOiOlpFnuW3Rp7WtmmThjPZXBSixNOScdXA5djT6yXZUH5UcHu44dwe1
/WpK/vt/48RhSTpFfnnj/+OEiJXfMrqVb73No22dRuIrxrf6a78nzp2iJ08ooB7zpYh1BJKa3iVB
9107K5zvIfAE39w1IXdwn586JTUgl5QlxGwMd2oHBZi02WuliS5uI9no8+YJ/6Tkx0BseKnFauBL
v6MV6hZRS7nXZHhUtP7yW01SUFcBrxSZ8g0uXDlR8htviWeJ7hH7qCnQ0wNMz89Ql5Bh9rzCV99e
ZXIWYjR1rAL9QPadrWqkkCjSWvOPtG6GrjE92PvGLT04njyJaQrR149QsW5g81ZzC+ZXzY4uIxv4
iye1uIaz5/NYATjBOVDJcalRvslDyqC9fTFIuGXFghrIrBBC8CuAacY5J5BFrbWp95MPn0hVV/yB
TE0Y9pM6CRAaUm2al0Ktdce4SroF9wNDmkZ3wqPCA3Bwwax6UI9RXrIviQ5TFf+a56Qgcfl0QQxz
4QX/0lHZGek2kJ43ba1fTTSndca6/bJtMvOTfMDcYSzQhzLeU5CXynoK9QNEWf9bUFDUrRlqmt+4
TLFkx9GCVE2IJi+H94Hw6QrgYXXkYM40M122K9ygyjS3GBUyHkI+nkR0fFbXNf6r5cPxPU51ING6
HeqdJE3cOBLz8Zxq8ElYDSBdNaT1q503phEFdBKoXTJhfG/T/ZH2wgV9S/DBlTiMctY1GBaHncOD
5aV7DMuI0L4LfhXGXbr4ptXRQFmh1z7SYX3ygqlh1rXyDL2QoJ/C/43NiYw2jHERzSDB0B+smkwa
zVsDdC0L8b1ax+aGVd0gVjddYuE2fNRiPd74HUk+70qmhBOBSjysm9SFh/RNotP8DDEXgHexdxA4
uTCBhJPzePPuwB0WTGkZfewJwQHD3GMdECq6rdFA0SEyAzyBuB6SQPOu7AWpAZiWSt4NgLAZSCS5
htN3DZMMEzBWlxVgziwVRUGYHV37B1+DbMjeoK1aLPP2bgU55ju6eqfK78/sH8ir5IhQP2T8kINE
L96PWrAGsm3YIx0MyGrdFlJdsVvxUl1oJtCFvemzKQiPmwmvSwfohbjzs3bdjugpTpF9Lvk6pPhD
v5cxZaijTunlHgXoCCsokF3ip1UUWCjJbKSCF7VoDZje/6c5XA64SjUZsblzmvaINxufjrAi5nme
ynd1FX+s+4xQ+WXvsX9FyZSPjkgeKOiQCc1CSMQP1UxfJ4Wf6/hCCnzZfo2krw6R7JguGRwIVHd9
R7E58hH8A69G5oF4pAFc4Y/VrVlPmeBqrO4IHgu3I10Jp1bN5IJ527QKPj73ak+/DJhsMdDKPpN+
3w8umYw5ZxAF6pMm/VH1GaiG2/5DMDt3LcmPZkFH+jhOOE4X3p27T2SCvmHihmSI6TjnSntf5E1I
qSE2VibUluLc2+bP1Xu5qlwo7NxuQH/7NFQKp6kKk0oBzcc16OH65C3Nt/YZDsB7v65OCFHzYpnO
KizbFVIQOgeFfVwZ6ZTH+0N6pd0m2Cu9yshFfDyzOiXJhUTJ+yl5WiQnjPRFAn1fL5Rm4LZvCLbv
87A/yAIvKlDNFWDKP/a3JouflcGKJHWIiH+d32yyaTzBGQlVTMlk5BZuuakwdhs+dag63g9uAPjN
Lsac4K+8RyyAJwyTzk7vqaX5xo3MChEXC5T3DhO/6XesWPnOwPe3Fi4zUqFSltiCnA/H5fFs9Sji
XBcS/zmEP5Tp4KE+fjfgkiWyn/ZkaHCTuYO+fmypLdkT4EwDdzAEZA2Kd2ZN0aqC+ZSQs73lL8T2
bs5OFUydRV3Dryeu7G+y6WaDnjASLzdUbJX3m8S4l90C/GsnrhCROFCX7t91CT/5Z1CJzHzh/HmH
vK9Cymtw/bpbW9yGOOr3TP6DK7ujSo0I6uhy6xBDrbmQOK1j7d48EkAcrvuxaemtfZd7m83VmVrr
pRvC7hlmcWMoQwtTyOhq1pEN04I3DCfknovAfWix7Tigt5ACkj8znW4vaSyIyJc5855MhKqSAuuf
uSe56ltoqLUzFiaqz0v6vOEjjldoqcAWQwQYFI133xlvdoSHvrfjpfJT7bJF4GI9uMPfNYj0mwav
I47oeTK2y4XL/LW+WJmBOi90QTYivDdcL49+y+RljCulfDU+veg+BvAWHilPQ2BSsV1L1hj0byxy
cjQjfIK03nE0WVdLq3SfwicHbIhzQd+l015ne8tob+n7cYzflYMMLL2NkjBGGFQLniRrsEENyNy1
70ZJtdQxTASl85bvwCHj9RxbHiZ4LGVoaJXnFPOQrR6WhhHJ4GY349n+DcNM4tKWSWL6IraPQn3g
JQTLfx5ySGDKg8d+Y5GyvEmFXeN1phNqtC933ZImAAlhz6OXBP82/qrCqxRRXbyxaPHbRBahYY53
PZJKWSdRllMesFHjFea+myD4jxg6ZI1M+MnY/WGLRpTftOaV5c99ZS2VWP33sh5zIt8gz8x2mdTy
Qpu29M+lkZmHEy1B2uS87Nza4hBuEv5spvA05rd32LDqsNB8PfmGwCyjuNjhf8wx8+7VypGDD6Qt
cTFM/fuR6tozcVrqjt04F06xG5rzt5U1S32PuyYhKA9YBKFeCsVB3dedFY8gKLCia1DAclSFwW8n
kwZR5/+tlRPbrzfwrMJYAuWe6UBedFGb1tnsIwrr7ObaPbVJS2/Zhesg8BmSY2qDHtqBFlhYGgdf
9ohJmygXdNTBommTl1fEImo1sFcqEbiyyjdZ+RyxbVeV9o2ABdGldiiBKRRyDt+NpWr6HR0o2xy0
QhybY3jA9JXmUKfHuMBPnNBDqN6Nou2kb0yKL2HIqAirb+vYDmOsD90Qavk6aUsv4u7wiJXupRoQ
u7I0RjS9c2COXYbPJw4dxRvxaZrcS+VM/3UCZrf78rxBLENR/kiArPM1zes32a8OiRibh5/ndBQV
pNYMzjC5xfmzIoXxy1T/N/9LEi3slMOlOlow2BJqFx7nkfkxILw12qlBvvYavOHBoeuKzCu6bvlQ
8JxFsidwvuEhEf0MgVPPvCTQeJviDhXRpgo018XY3JjczEBvAQNyRRRq7ixiqdeeFm0/9jUDWJ3g
MCQuZvFzJqzlNekFyC1fsGOrvN5EZJGMfKCeiSIeQoJWMkmc+g56kXbS0VfH0ZtPwXcy3nxSoCH5
6BCoM4D1OVQqD6DCgpQYAp16+CoHcMu1cZsQvct3K4rE0AL8tJEMRa20t/rwBThWYe3fL9VgPvt1
sr/SslzVnRnNZdWdFjQ61EnyKeoSG7Ozbs/l/V8eJ78Q+CCALKj81DZ9C4OT4e+MRvg/MYBAgwwV
vPRbxQMn8jMHa1tsRhL+VN1RQFPlusAuZaPS9My8En+Xo8atsnlVbhtbMZyxd/q3Iy4xP4G2Ed4l
SCsj5wpLVAHHagTEKoeZvU9KP7TVp4Lrt7+UjpXZT7LQDLLu3g64mTa1PGPeXTZcjnAQmirAbvz4
7YOZs8EGWDhQhadW08xYHmM26q1W5oPnfHy2HTAzDxoGNQrmM3qvt/ZlenuVWGe8bsAofhAV5mLh
//4cfNO9D+ogd0y7eFdfbpvDRO/YzsiA0OKHlJy/sbwCF076fJeypEEsrg2v8bjxySvecHYo0IOs
2GSx8NCfnRGOHfREA0VyvyyeZzUgqnh3CV07yw122zd+t/hCjGz50d8tgAGMmpz2r0C7qYLsqU0Z
dxTtpdwT5COdHHPNxY+lp8honw3442Kou7MQVwsDQXvai0GkVl0ts3SR1D2F7fsODkMGmqypq3BC
lsqWIM1YxmOhmguQEwSKHLftgipq4a0pwpkAlJ3bUqngwuu9XA5cUNHp7r08GbbikKXBTTHIMyWv
kS6uujPyL4ub8GYu/M0x5Kk7rrG1LHNBL4PjH2ze/OOkP6umw5DlaB6IgfNvrJTfUOHDGDVvA6Z3
OB4HcZqs2qktwsB2sfFH5W9pr0ViZSRlFQaotzTEwrUjuQ9/BRZiiuKkuiD5ZBH+fwfuEx3CrXPX
PYSQ9jWApRJjwyJjcAdBFmgzuhcj0dkFMhfWw7SyMuG4wMXbqy5iWClNPjy+YS81s7ZC5tWAfzLU
D/n+Q1c2CZ8d+GNkXxROB2nR9ljkYLktElY6wxGfybJ/N+YC3mcCXl+SQKX7M4goJJm4MQ/yX46b
asRLatfrrf9wIo3AOTcrdGSS3CwVZScEIepNhHDNm0USzvt6n0vxNv3dTPapQ4Ve7+nXPirRGRZp
WETpiFkYGyygQgHQ2aFp/e6D/dJqEpKEAPzPBVWN0KyvUrVDjKoFwdchOkrZ1WRaW2lSM1Gqnf90
hW7+fzrSVo36ZXQRkHkSnq8lhX4TdYWoMBDpIvb8jegEltLJYPnPyzUF0z6CQynn6x0iJdaScGLF
oSFRzvFk7AQKyPWEyEyqnVHCzGpX29ais9cMNfqCtP6xQPKVUtnGu89u7fegXA+jzKCMbzQ4HLUU
F45r5PPEJhhh3zYz5zfIXnJC9qYXzU3dHvD0ANFp0//wI43PQRKU4K2IqsWF0fe2O5hUoLTKtqJ6
+zySJi+koI100D2Dl68iBTXeeiHuGwqI4yGg4pi6CIEzW61lxsgvjFg+Llal70jmM+klJSseBMLx
JH6s5RjHxSOsNlIL8MEYiOXM1mB2/HjA/et6tD3Rvu37gb/PDMczqZ5WLicr5LnX9vqPlOA6hynI
lRMpA3yy/S+ad3oaYYa37lWghGZn8BV187B+XmooERmxbfj3je73FTTXAayVgVCbhOOc6g2HfBmF
/BYilM6IfOE0JkVw1L6V+PbL73qqomH2y90UaRw0sI/McCJqeeZWes916+cpyMO7kca0ZUVTsHOF
t48knX8BAy8RWjiMHpZB2xPSlfInhLO8s+J1GFxZRur5NTLUncATTgSPlWQQE0GExwJwCjO7X6Lv
5SAl/Q1mG5nW/KUpfMAgzvvqoBlD5Fz9sHej8KF8RV+pUtgWjFW699VIXDJbry+lQUp6PderTHHZ
fKAiRLRXeinB4FcoSgaz6169KHXNOBxPC0k0eBd//nqdIfqp9Meu/6d8UmhvuJfVg3nyr2B4OoLT
YdYinfLvZQPaaTWXhw/GJ6JD/WrLwrtlSzSORstl0z6ukuG2Nsk4ezGx3aFUJqCpVnDOxqO04Moi
xall2eKU2vT7mquImY7mxGSlM16WqFT5VZZoxxPFb9kxD57qokunSZYT0HL8jiopDs+B+nxJ6/Sn
iSIFUHZ3MEX2bfV2aQjb9fapun1yJQZd9VAvnA4MvV2wM4UXAt8tsjFEwA/gHVgZWkjHXcgmqBNu
nHSZdVAauhIe4/l/mYZAEv1k6kNwQ4iV4gV3hus90Iavl5nmG2PcnunMWqpZyBUNW9Yh0p93sTwf
GuKJRHBwNn+FQMEdGbwH8WBnq4Q6xSvcpoIMhW/izgeCNvybd89Cl3eJkzIkyK65IMIqbVfBu79K
2bU4MIjAvBJLYdSFFdCkCMH5gojeglT/RAzLtFusrGa2kU6HNiKwnX0N7fWcBhvyAZCmzVKr/uPN
YVv8xSe+07lvHsJ2nR5Wd9SOwCQR3SiCfpIJhttGYRPvPqeq/Czi7qdS9wnDxegeFyHFHEDAymJt
9RRvak+LvGkoKgRvxD2RHaMP5S/NlekyX37gpump4ffHYttd/I21yfQWOwhaTx/mey/4DnlhKSgK
biSxcGQFGxsCeFFeoPeQvOwNJxT4Hl///1uIN0FwAbgAy9ex2NyOlZ+oZfpd5hYjIDPytqtmhkso
jdoZxaW3kx4YcE41Dr0iZJFFSebBKiTseB9Dv4PdgMLIAeppFNYWhfYKjEAvogvc9ksh9Eq4lztH
GZoawhYuGBRkJo8CiW/aqcLGqPgqVjQK6JiAMfEmZ6fu9bzfpoGOcECX6QTgSIwoRmk+byMEnfQy
v1gkpQHeezTSKc7easn5yucdhnRQG2MnUZDhO7bl2Hu4Zn2x5FsFU4LOHYgOKD3KrCliR/1z6aWV
pf/GnQIMWqfWJ9PF+VBeKEhZbOlQnWo1qvnuPs6dxbcYROc0u1ZPouFF5TTq6kVw3O4ic2EObTVt
PScRsaWQDxn1L8cF+gbALP01MYyDXS3pL/DFRsr+kMnM0USbsp6qeRCAPzM4iXTdv3swMFikIrFQ
F3PlXGTWYek7TdXfQ10A/sPYmE7HoquklVfdljGUH1VgKEdvidH4FH6GZ4cy5b9segn/pGbOL7XN
Iq1WRbxHhfI0m7rA6rNT3mmGcjmQRMaOg/8sPxX2IhSnCHBRpBu3OBfgTFx67n+nEWy1YGHGBzcs
o2HoPyX3S6vUfB2fjkKnqqo1QhPJ2fazTBp0gE0dfZhBvKP/MldfjT9QTKZ5jtvQwGkUYdCg9+9W
FOCi1q+K2FvoVaycEtqy42KPc9unHEVTKCXc7puh4sdTFKTjKG4fWpNtfz5T9T1A2CXP+BJibxYy
S8NBw6J1ZIARmTWhuNUD5YDE4f9NOYgWL6VFEuPDKOUWanrMC2ez+JXL2tcwgyEGi2tbAXgb/mkN
vB9H/BB7r7ccZk7DLuixPnAkdGUyxuCxli2uJjhZcmaREUcmzykPYj7EG/5NsLV+OX575vRzpdTH
6zsyf0G3oJDRV9/XpaYHootQviSJkOiqAxkEFXgmxae1K72XMIqsvMFpWnIJudL/k7O6vlQXaYZK
oC8OWShwNPHzKmx7vBlXH1NVSLMSGeD0jNA6Mnm3dK71ojn8h88CRT4LDmlgVZSjdHj0q+Nk3J/S
SqyDDa1lYd+VN2itTcaM/xJ2f5pHtv8vVH2KWLaq1bUndECFkSwnwtZmz+wuWT7cFwjxiKknMhMF
v7fIc3ud00t3dlkDeEzT28cmJJ+xEOld4BZsh23LDqmc/kYzJlQRCRl0IjQTsQi2d5ZYrVTfjfFZ
3/PL3GAt5cETrrbqoSbBEVuKQGWDpnNfTg7XUwuv2wEWczhf2kch6wTiTpcpEahFtOdWNnKL2V9n
jtv5+DEcFwPPa4eqRTKK/AJ0TL+3Ey5/vTMAIOwAlkUINcTnWM4W4CAaSJZDndcMIHIL1GaTDK9j
pGCuOzkyDzSdcEndd0GJ/GgQX11nt4uKiijmmACqxKX3MeB2nMbech2Jh17MfLAb9kmjDzf7hspn
kyujSgUMmV4cZVaiJ/9sVPXrkrRxtGyqG94XaIrAwMNRTVERKmOZq7aEHFxk2ygGo48yvYI3zECG
agFVVodZuj89vAK8WEnqs5A+SZgkGvzR0AJuo8ZUURFBp8Jf+WTWm1zs6k468NsReDiKiam7V0GM
MHQ05ZpZI39K1m9MxQA6QzXNAAhUrUjdjxS7eWXlrWcSVV77yLvphN4SPM9ceAZDAklGoWstatY8
RnYRdlW5n/oi/GWrjLA+6GrCfEfEcA2FCeHD4qYjMGq5xYiJKlh7IK+GKhMKyV2nEmhWYLOsmDls
RPj20hvm3rQzhmTnE9qkF30Pw6CG3w2B4TkejV6j6ns/Qr6QMaa2kCFdJKdrzUoX5h3G2nTT85qH
4mYnhs32Qwh6s3GppTbvWsryo26prnubYcfzHc4QGf5ruuzcLuUEdgKhFcvEw4JloXQ9vXbJpqn6
DtEpy2K7Ddts+jyYU4uMgumgRdmKKeqjF8fNNshRl+Wda5L2UxvG2rIlWor3mNRHsEsMyunc4GmR
FnoYwypNttNWaU6q5osuVVIPbt0b5yWvzvBsq4L8QK09rBZpJ4ZAH4mwmdK0MjPoAINiJTTJVFN4
N5XCVA0RdQdZuz3yv16PcaF7BvI+sMJ7aeboQThwFkhEmuFDTLsZYbiYD6EANMub/120WO5U7sCb
pL7xt3fvMPjoQQ7AdQg9y3DIAsclq6ZxzxfzAvLJ/5+NVDM+nO1rEpX/URubsG24UcQlFPW3cV9q
rPafrYMiNWm6xo2lQnGlnbuK+U4OSnK5QMAn/eGPdXKhiErdxNk3ssNBim+XxL93+DLEmJ7CYhXW
Ov3GERHlUkeLZg5g/xt8uxyoSa9R0OxlD2XRh07Gt/FfF6tWR/+90zovK0mSKk92Z/NUvqtWQ0IE
aCg+znK8yNsZnOFHlOsM0KEpX/wV2Qc9204Eo2Axm6NVj7O7b+X7TEm4ApsHLjaI9dseMOUCadVL
4dxtdE9Zrz5wBUd63pFtsWDXwOAglkgsVpEJN7x599VbvOYTRj6tl9qlLEU+QoQs0Ps60e3xkbrH
A0KfA/X62zjWFFetswRkLVOb1P2a6zFDJmzylRIcTVmA5XpKdG7EvrSLutPYlQBBDc30mGtNA7kB
9tLHQSo2m6ADCb46ote3EDZfWEScIgOAbFXv+K9HmCURI9JjlZOPtGRjcKwE2a/Zv16kGop8nEJY
IeYuIuxkfnzIwsC69D/NVMLlq5lyOH0/UbdNEiv7WzGF4jPUOAizUvftjjVzwSPjJQbM0cJgYeLr
DcJHh06Q9k6tgiYjYTV7JpMWbhILot0VqjtDZ88/2x7o6qBXHG3naIWaDgini7RRAhYCnSx9JARE
I5z/IE/YDo5eIQnMNVcCYv3Cpx/7EUUGCd2RSFAakc0r9Xgi08BCzrhrIJ+Iy5R7InWhiZsKA6o7
CZvDBdyBq4FHUrdq/dOhrZ5flLB7P4XTAby+wr+LckKXqBbKGny/SRiz3cdIgGSkT6CEQVUcmYpW
yY4AH0Vci1mkDOK1IOLxBBwk8p1+fveu+8cO+NeKX+9717GlvTpOECnDKeLuvQp/KvLG5J2kWqoW
DXVYGSROVd8U872AD2WkAqKlqzlCkrqeutXGbzFXJ8YSxxOu4WXBnfpNUIzfCISXwBQ55VjM2+vm
QA85UP8RWrdCaJk7+Q1Z4PzHBwgDMPHHW170nFR0Y/kkMd3G9rtsCNC1tO7f7upXUk+wp3HQpmCg
0FOS0h6ev2Ft9pLc9vdNddDF9E6x0sL6ykWm2IB9iEKmnZYTflC7kRMnRWv8kR2wFK0hBNDjxMq2
VGtn4hCLmdAy7W8qo1b+IfnKkJXToNl45jFn+CBdN7vE3R6fhmzdrK9iz21PwnwJMVrw4cxXcXqt
oinhd9OIGPf3QSNeORYPt7C8ueIC1+nWW6dhdTONdN58Ft7wBwK0l+YMfCVjO+BGAV3wckfjxjzI
2tbNsXC+ys4Ov9LnSEpdvTqWCCRcvpVTy0EoF0NSuK8YnU+tdgb3bIqED16VwMxa0rjf0BteLbDW
EC7elsrh1VJlLAasIIGMYS2HvsFDs999UbRmmqf/XIyuRFCVsiteriTO3pd3Q4AfduJPpFztYW4r
nRqqWmsAUOUoMtUyl+5h7cyxN5uZ9cWIKak2Hn/EkVoQBpJ6U+PAVdrRdxKlaYug1arYkWF3V0Vr
4sltvQlcDC+M9QsxDvEQHYwQcp7fAUsFqzzl2uXUzjwNJBkH44ie72H3m8MKl8dYtOfbToUII+N2
JilJswCRM3ZpUJBEixYsbtZ5PqYG9eX4bz04wSXmURHK1MD0GyT9zPk5afWM8sLG4ZVU+zFBMagT
BVoIuFOJ65eDLTFthHjzyvrH70EoP8AUjzf436g7QuuoMjKOrN4Cxt+10zb4oHpNcDYCAimev2vG
xlnWnbzlXmXDedbrBsD1d+beqgrhgFn5436G+S6lBVm42CT7tkBFK3X/XfqANe3M4Qqf8SYXzCYb
4RCwWI9/YEBaDgpTu6uXTElPcqlIyMRjQ3IWiJRnQGdOZOIl2j5mUBg8ERkDtZfoHggm4E1s/szT
jfx9s2ZLyBrqcg249UR2ZDL8NYqW7v5KA1bLzbCaRhTEivhC9SjFhEOjrcBtg4iPAf5t0QLsLVfb
JDkL2fzQ+SQ1uluYl7chkeRHgyxGyESM9mZ0RPDvTsUT+ZPzfXTSNyTwAVTz4nzH+Slz92jin/y4
JkD8dcmv73xffnag/69lXy0qRcCx3dSkbTEAFTH2rtExYI2WbPKafsK0ckG38tE7eV5DJ5H+ArMf
N3E7PcqnUq6dvryFoWW8QkDnCGWRI0w0g/xPamZ2qytcfBo9d+UvQAIO/+B6bmF3/UvJ0ZrRRXNH
ApP0TGBqgqR7omdOv1hUPsG6gP30rrjwndd2R6wVwNxnE5c5+p4ApWlH2KMPHM+8FWMwj37YOky9
gOvkc0j664UKK39U3/fxNwnd0e5bCP+n//jBR9DyxmPslovKhblaDns67LtrBdlzI/0EVdQ+qkX8
0Szu0Fsu1Afaun/59sBw1fL60G0M05vfzQupTXgt8TkADX3hqGOgzueIht7FffmZxb6459ZfKRgl
F14Sixolj6/EhbGWW06GY57j1Uf7dKMj+E52623n7khVXh7EZcdyIxO7SqW1IxPdOQ79lXQ49cVw
koTzqWLlyeV89cIHf9HpIZBJSD6OCoBlKWDTQUiejH7RMVe8PqjVlUsEcF+VUGnID8QcQ0FilPz0
Gp7oCmaznp8xAsAWioCgD0wbHYhyQzcjvCDmLSJP80if99dGiVrtKHQzCzHeqczz1hfIWFvDfYfE
Z9Ns+Wh9rissQ4ap4qavezHJd8IHr3ImpvZ6Z03Y39MsQNTvzOph78wgAnCz6d1IcLZC4A04bAop
nCQZYS9zkufvyvghtv6+m4ANsSIG7lNUQ78SzlFpN55dpmvjR904uP0ZoFC3wtDLmLWwoEN5Z16C
Xk7WBwjQtb6UlNyT5wWpMEBZMCVUQ5iHOJosqSYC/OkRCDE+0F7JPVEu/m06zwjC5X1YpiFVRrEv
Gmf2CJ0JRfk/R7U1jsyGUk3ZJLfXibEUrKKgDNO0WeL+TUv4x0leR9LdCWdf3eSZ9OEz5FFUGJsL
9M+52d52U7qrEIeVa0eQQ5ccMMQkJNc+KEnx2cZ8I1Pyv7lFsIoXtM3F23VpUu69GO2eoo66j/YJ
RVyANbxBtiT9Yy8pxmYsuMnYFRJVKatiaezPvIUn+yXtw8MTE94L1f4triDoOJWlzJXNp/zHup+o
kW40sltkEctPbbbkvlRqp1fA/aLIiMNRcOuqJzPbJwnOQm/Ps0jEyryzoQZGIa2qnPi1vGfhki7N
0Ywm31Stj7qg8qmVmhf4yemeWGNU85Gi3EJc+x7yvZj4HY+RgkLXMj2klfTHCxus95he0uscxUix
yXWZo+YChONypZYu+ZQJ1R63WfFrus5pA7823BQODVc/jbU8pnwrdXERt38Yeky8XUBaZ3iFjAqw
/hgW4sARAtfVuoPfkMDUiXfeqqEjzhYjiTOLfuiH4wXinVYQutv7h73mgy0APb0Ma34pEtJ7604h
IvHNGo/Vd1d8X0S0qYpi6gcUcwY16sCjUKqbUNHL+3Egeu9/K6UN4Fem6FJnT/eGVq5/s3sW3jpb
TiL65SP7hLE0+4NFhCTuNZYm9FGNZaXghgeJqiWeOzWOpxWrT99uGMEfSDWKO1Hy/XcVRicUcLcu
BfSV4XWvwo7K1w5QzBYgs+sbz3CauMYtD4AMqtF/mWCq5Y9oMBl2TMmN3cEuuADWzgimtWXScTzY
pb+QHkKkEqxtT4UeoOtuhRrIwFifq8sSJLVNgV7HJHjKagDG2gEGP272CN5DpYRCKUKr6Llgya2S
LXvsLgaEbynShhsd8/J8TKJQhbgv12YW/Btr2lPteSNi4u+8UZQ/bq9rUXu/TuYkjU/iWWrsHULh
UvtpELas78L2ApP+ndM6Dh7GTEdFnZbKvVT81WDezfqCFcUN3KOY7OhVNBVWHlLjBjDxIu8Aaqi9
7rL0aK+giMMTrJ086VY3ro5m67Vy2QD+p4morW39/RvAoC8sVgdqUFCkxoehvsnddBiOXHBzChKe
Cdct3vEuKorFUY7fiEmWbcxkLhnqrot+1q3kqD1rLOhsvUjoN1hLGrgjpD3FOmbSKIiR/YMbw1EA
pxApgK8bR09GB3QQ4+sYZhjLE8BtRpU8ZpjfbNKY4SoIsCe2o/HOnKgaAwC/51drIndW0MrG4u9Z
XDx5OlKEBOhptzSsqZKrmZN/6spQZOBBgu1PerjRl8PRjXFex1M8fxeL+Ya3S4xk3SQjEAw8oJiM
siH+RlWpIH/yFCQs4p749RTDH0lg+7cu3d8tFH4RMWzNVv7jljV7bwhIEX+8vER2TbuQawcsRG1H
x8HHSusLVZGKY7EDgufEFq3JhvYvHBk7VDGc72fSoivR5Zk+/v7rvCa0Jx+nb1GmEPBcWJ3mMqZR
Fr93AyYybjZTMCqr6g7/3xhzPr0wpQRnSThi8rCh+NnNRScH0C8oLFqSedVdrayTvB/IsPi+toGo
wP7yNhsZWxk1b52l+BrXDL0jb9JSw94WdabwdCGSc40GAOdblVr/3fD5PIUScxjDBlOkGsL9EElQ
GD7Pv4EfKCY2EAQT1t7wYH9aw02Cjzkq6sjBctyAGxr9q3Y7kvhBO2ef8kqYqTW9qy/J3KS7u6b9
TR/LZj/0KqQSpi4h8zQOnxAQDHI49jtzFI2jZas5KuJsGWQQdK8uYt5xTAVuKIO7W7D1UtUTKdxK
Q46JWhNuJMzWXamnhUlSlgXIBsRPQKMXmotOPpuXtYLnR4D565m4Ft6aEX+KrgVlYkQ3lwxn4R1c
f6ifpF1xshEpmapTPaABtNEwGDM/nq0G588LpFRF/AX1BBURPuZ/iQOitLk5tSfJABXffGZrnH2y
lnXpCRC7/FkIYPxyHD+1Hd6fi4sVII23m35IqrdVSbdlIMx9IE3tnxfoBMPOGOUD25Z3kh84v0uG
dK+ov+gxrNDKTmn3Aqu8C0Rr+eqawCmGbQP+WFAU6y1qar6ZNjD7/qUEvvNzcgCgIGjiNEIYke/c
diFTTWg7+0tnOQ8XP2wyYPxviFYHbHyLREQruRBTRdyIXcNXdtPAKJw0RObwygZMLDNLzrdnxJrh
2IUn1KCXSYaqyvflZUL0hLIDwrK3ySZdQx724WPv3Sc5AH0N/EsKUa4sstluHwvMsiz8AjLibBBt
3i2FSCB+l/ByTjEgqT0i/PZyAb9gBgVHvdsNcQLOCGlBld3EVmVXQtbpNkA2E8GPJSz69b8nRYJ0
ez8mxXGF/ryv4tWcvdw3E9nH6lKjHAbZNBeGVRXyy8AnT4Idvg+edHSkbyWP/Idhl5XizDHETA5s
y8pz2/W15nr6aytYiP+9ai/po5/rh2OVYgovymQRjL5kxtHNY1YVnSbLEGLad+mIvpXB+7VJDUzh
50VL6XnqsZVka+Yz9QyfdqaDYoi6dTpIaWzX8BNwNFYjc468jF37bo/75wF4e+Gni/oyxcXe/mDX
190MKJb8UCETa/zr0/1Me83H7t483su153WuHAny/0xIDKbDssnx2Le25krrQM2uM2+/Cd3vE0A0
PXNIOIWdK6yirV7Js9gNo9ww4Yep0renomXz9+U/oPN4NIKecSZu0mKNAQQHWYDGuBb7kF91vRNA
2lzY5uMPkj6cNlh6PAMpVlA/4PYuNnC4hKH77THwd6bmonYEB+rBMagCr/YHSn+N3ZtGpAb04mRv
7sJ7v9LKgs8gw4xzUU2q5QTYdy0K+gHG/HXNhZZ+iDfYD2h81U+COgxi3IsO/Fyt9VnN6SW1Dg1C
9kb1f7d4t0S+KfB3x35k3oCyGTM5amHWm1r2JgB65R5b2YwyogyWKT+JC6UPchCRFgyxcOPZ35NV
GucZJNA6quzTHqUzpa6GqRbO/B4FTYDljmhD1pSN1o2B/kwP3fRpPTmEpDfYkfxFBNReQgK+MClb
hjk1+FmV9Bq1gfbnNjavQWF3xeYWtJxmhsNih1GKIKXq9v8NMtcqat0P7qINPvb38QqhR4djWtiQ
7Q0ZDB8lOKaIdiFee8MOkokJKWidDpMQ/uMfOs7d0IA0abITKpZZruPCdV9z9F21d/3IFSF7ObG6
aDDgoHJsAHUKyy7H3c+AGKPshQSMz/J7cvfUKNstF9w8BmgfNw12Ncx8enOD4uGu5awuPLpV3gj+
GVsF40O43Q8HpiboxzLxCVwVIkT9aUdf4HmlEJG3hw/ZGNB0fitlCTDm8/oM9TSEWtAlck5YCpgb
qzkXvZFtHFbiAe/qK+pKBMwlunAbk9l/GTa4wlg2pott6AIGwBiZIPwbiIea7JG56vtDOq3AkjkA
qmpr8KKuumsrlYvQyaGObtvN+R/mLo9g7FHWdl7dkG+93C4PvzJv9KjapKvi8RKwINUty5dBbWQJ
qt7ERW6NeMCiz06zmn0EBKgSiUVtkZPCdMCrHCkqbWW042mBs4dwvdPtypJmWExwuVBJEc07VaIQ
poEn3ogUOhZ8lyly7C8crA+8vHEqdT91SbERO1yJ7xoEbNz4u7/0Tskh6LbXTzLHVFgdPyPDFJmL
/XX6JlH/Bj8Iqrfx6rMMolOG7vvgzXONSSb8RB6ItH7kHXSq7ExKLOYEai6KoQV2LJTEYX48PVpC
wbhOmAYLaNPiji6a+71XAls/Jy1TSP3eLyOXriGPNetO3+yv9Aa5CjowBK+SbRwi7Fzi7gWIXxPM
dXQd/nePrf0yppvi/qCR+VK88A2hcwh9sHORLJO1LHKdZnZ6xM3LTLqko/REEMuoPvbMTZ8bWiNP
Nee1YOR9AM70wJsRa6QDgOofmKfg8OuDwVNzwyBnpJYphZ+aeuDvUug0FoQ3NR2Wc0VTObV4AKdr
EBTbd0MFdj1g9LxhTV4Tjd93AVtmS5zDroHcHGWOyMsVaHFEQ/2XCT9XU+sR/PBpHUddwj4zgyBU
wga3jMWzxvFFVVob0yiLuig9WI5532SwKsi2p63ZztFpw9oIHhrp+8k2ibRPjjUK/fHZAa6nHsyi
lOPWVW8GPBooR+Q/cp81MS+4Q65KGulJYOXuUYUG8uCkRLKZbS1jf9JOPOYOfaYJmvDNW7GP+VtS
Rf5XfMdZ3gx9rLeYVGH+vg04xGiI00eYWDE4RAwc6CpVYYORgrqjgv/Ai8Ep7NQwLGG/ftlHVAh6
SfraSUiXIMAAvA/owScOY2j5uCXYwWTF7pyjNAnEiBy8BE9fbLWfy3V4ef0kciXP1kQKbLaiJdNx
mIS7OtgFhvn17BRduduR3zA9c7/CBxpCUCYVKzYxDO5TSY9NPIGeOenAko6FqFn5/XJ+ZNnlyOvi
UDC001pddrWH914e1CwrYy65Ls0vpp0c9kBZO2QyyJVyOyHQusbl7+NF0CgX4l9EAMze84mUyqCu
osztY/1ct/sReVietlY0tmnighDhrsUt0bUK27X3U8a+iiLdD8IutOu8Q+Gk0DAMagOYdTOWt1xS
fGURuYoH+f7WuEQX/r7dVJUPF1enkS21Y2KSOXnBrAQTYM2qj65uBcja8ETp8XEcf9T/eoZLvexM
dv6aNXqGELHSbb3O/i84nQVSiUWiqYo6cp4Qnr2pEiyudUJTXw/ERwr7bYZIvCx75sBeF3kD2eaY
NaZI7ByPdOzCE3cfWipcDoasRw1gSulCcPX4l9KnmAyZ4woH4n/WVLqp0K/UjU3wTlzBHH8QyugM
jKk07s1eJvXAUvdJGtOAfwerw6X3eJJCQEkwSuJ6ikPyPuerIsuY/Ikdjg39gPYNkbNl+hIl2332
kgezWhTGFjLAtTjw5WKf6n8hDO9+Nt/wfA3k/xT5XAIneYID6zyKRPlYe6f3wcv0yORyGyZEtm2d
ynu0EqAAgWaHyO5PVJ+qDGsJUpv+SOkx+C8FfXGK6er2cN+6rFCXQTALB49YpgPLw5s3Pd7QOHun
MamdspdqOOklZGdrwN1KYqxjdu621RrD3QJ/ASxYQsmYomN6uOv18ZggNqTG/3zx5ssyw0R21Nnw
ozmWF6qgWFTIDPhVTxYPQ/p/LehErk681ZKaVtqnCJGM5pqNPaHlRRVhYbT6kdTf25Jf18fafu0w
OSOs1aVFe3eqaBuf5QJ/w4fCr8Bu6emMQckxorDiBnBBKKPG4Ou+i6PQuPI0I9TNCintpjLmap9H
SeFcNNff/UiVPNeiik79sE6nBOhyCTDaBVrmuj4hs83psxUDpc/+ZgiceQOLqOWT2ynoAWU3bYXl
v6hCOGjECkK89ZAVo00D/ceG4h84BA50cqHSYcnTQFamHUhy+Z7EcqVZXDqs4E1W4w2rLPsdvuaN
o82qHQO44VUJtr0EBfvhI27Fp79zPH3H+P/Z4Ld5kJPgFYz4sjMXr6Rh272tYCAj55nH1PNXuYlg
abSvZlfrwIkIXrRx0omX9PAzVljLeoDmcSMJKk1NZ4v26chROHY9Q0zMDqEarU0yQafeOSdv8Ov+
nq6BViccAM17+kTvEQB8u9fzeRAB/JkD89/a4pdg7TEcDPTjw2ubJ+cXGNe5OFFfHgp/mikOY/bi
c/IdS/KmvYhZFInIAhMjCQ6LSfwIWWaWLMuAqNDR/2Zv6X5S09rbs3j2kG8J4hBLxTX1SegplpCW
H9ricqKp6wyJ0/KRDfrnOTq+DzQOmXNWNgC68dF7xMnoBHHc7BdGtjav0CHEoY4Rmk6tU7yITnvQ
DmNvhlM/QWY6AkaTXns9cbcwQemEsYw+YDwO238OR7Rj5v8E/XqHSAMe5z480xllQEqLWDqzsYs4
cYKz0RmH02soe6oUoyYJuUFP5YiZxU66k3Q2GW2WKGxLiG0p7m9XH8oXgp/O0QpNw8UJsCcZkr6I
zJp5pLDgrySV2uk/5px8D/46o+ti5027tvo4KtUsWLypmz8ga60eYtL+ZlngYbQyMrZXognCPIX/
Fl6O6bCFYKwelbhKcA8JPjPkDF7HXMLD+R5J1WikFxVXHkYNpAbLgdvg34qY9bvpbV88ywEDDXRe
RHL8dJ4gTIQ1460upg1OB/SWVpn3+JWb70OSB0RFxMPBg28772GsECjQO/JeldoWH3Je9fBLQdxb
8+h+XbkLpWTjz4aqMpcEmGz7uoCOWAdegjCaGbq3izPME2xmL/3QWFo5eyF6tAJ23JAVAlTzfGhs
Tg0JQfjHJ/COPUWhNM9TQOAJ4s6yO4uWLAU/Pd7scyTBG6hMK/vrYQ/bZIPt2LzQrHRtu2K7YLHR
XaqADaSQau0Q2dg6isNcLxsHm8XE/1TUuIf6mZfnGgEeUeo+/I9v/kpbhxKM7vbmPKQIYSSyRxLh
Batyktk65JU2FlTarzjCbOLtp/C082S6vF7e1zx4xUX1feAn+739tu3UeVkqKpvycfjFPfRpqcSk
KFKmRj6gOa4uecJ3T+EFOWMPx8kiFNfekNgofnWAsAOFzqa7yXzJIb0YUJjd05zOKy55Lk+dfUal
r6zQwtskaAC2gXZMTyFxs8JkKjxLI5hPSyrHmKPsxR/Q5aeYgvM+hWJuqhnc3wnZHRtMzuoEVAaw
p39yVRd8k89dlWQWkxozNcBNzfQ4DVNSB+OaSYJ4qlz37Tb5hFkhFeu/5sddqia6VF2KSg3sJ/ny
bBnu/XwxiTidAYGgcXFwENHd1Zkx7u8BtBZvY5rIPzntmvjICbxdNK5gy0dX1kKX2rEC+bBa9kyw
J44C4Cc2YkEMqJUzbvhvnSYtMcmBIO6cEZcu3uqWQLCYmlHSOX7knzMpbRWcuzg5eGwmmkKhhU0N
GQHLUZNMyVMhjRTxP90/HuTaXzZdA9GMF8CKwkPz0YIdbX0MnGkSEM0RHWMTvDjuv5mqSx0p/45E
NGNlWULtE7VFdTzDdkeI5AYfZKGhezeyvqT1y0REICYnO5isxehzQI6/Moc/kMBvF2lychFUE8tS
FwsAWZWDEksExIOoccB06SG0sXNNpZ45pTmTAXyyBPd53C+2cGfX65/6HsPA8g8qTnHFWAAD1qy2
chPCR+z1nuneqZF77vS5w3j1PcN31NrNANm2EVm58aCzQNN8i7XLQSAAU+EtRr8eCrLbjwEVITKP
GUgmjqVajUxaKiiPZ9GXJkxTrh1BKeRNNGMuG8Dv82PbdpVE7nZEn/dmIR822ArVg6CrQ1Lx/NkZ
G4G+/NnWITE0BCp/lHr/dd6+nTQzGx3XiJoF8T45fOWBBPT1X99BObiiK+yCsZYwMCw96WOQBk+L
5V1UaHeAMPuLdykNbsM7v2UXQVOQedlx6Sc8BhNxlPnsZz567X3ph8eR9Fr9y3bMz/p8DNDZbqt4
z4EWdwC9Cgvu+977DiOXl3NfZTKG3ww7hcmLwRZovZTGL6Vc+58kINNHMYKmGcIkd4VFffgcsbxJ
t56TE7pexsL4FvQk8ABJOgzQADp0TH+iuQsLF/aiTwpqKd546Ob7r12+OY7ld4xL0dK6MfzRNA2N
g70OCaQv4NBrEOwi4qZY7af3WfDfvCop47NIRGgj8BaTqal40iTUzFXz8FL986hDXu39LiV6ey5g
5MvB8nOt68hgGhTv38rSrA+H/zztoUK7Z9aqbXJGOfz5SudmERbdNH01YDJ7/imM4n3sW8LuDtkE
wOq44NUQQql+XFq21uV+Rh91cfugOc7UgpnHgjwefsYvhW3Nbc74qpo2dPRu0Ek/HUnzPmtHpzKV
cN/ll9zByJ/+2/ZKbfmqzWsFavo4F1JSjIWUIccFDP9APyBrhSp7p1zGqq27Pyubkx/8sY77fvFo
y+R6oRVOHyOkHxFTF3/H18yBG/pif+2OqiJRNXlYYPM/dVCj/d9AHWGj+2LActv5wpu2XfHBGWC9
gp12xy3SjbmtAG2VlFIwgBF0VRrSNZXX1z8g47pHxnYG4J741iQ6UtvBql//kuyiBnyIcif2CYxt
gFEL/zfsyCOpcGG3HtYoxe1wbMsx+jSkqDgk8YhgxE+cVXTk6F55djKASTpRqUsdM8Ax8mYcuDsP
v+btosnjfypoHYovrPvKenawqwFt64s6iOxy1CiNVLUY8s2yg0e7cSItinpQw6lqtn6ui2NHBekW
GEOwxsC1LyR+yJgElfCQix7pPi7KsyML2zqw8v/AT6bF4xVyTOOobtDVUMqGyp8/KhqjVUbx8Xmc
EGUmo2MrpGMTgjefujW8dItGvZA6JFDwRuVSRStgOjKqrkqAud6n4/2fX353SxboBJCfNsJuhOJG
2RgOcW8qQwhJuP7WGG47Xo/1ALNVCXPrm/ZlXDm+zNw6Q0+87GnCuYh6LLyZOraQJjN24X/SXSAk
Gm2jk8ohBnluYLecNpk67Xvk8zERbUM2dhTRg4fruUljJvGtT0SYfMbIDKPYOadMpVbnBJ6wKek+
Iw37XQekn4SD+728cRVenUq+YSqjGnpr1/CvZQiRJvr4MGK+rNYMWHzlNbeOBGb2dwIBFrX8bkBc
wU2w/25zi5vVCr0rkq/gepPNZmfNwtt2g8ANcYgxQbHDXZFGKHHKNb3BJY1aUXNPmhbRF8R6axOP
7panFzmyMngDhC8tQVjf3TcG0TozrvZt2ZqsBz/KR4E6nmPTt796u5mjOKm3eDN0+cKy5cJaIo3h
r/1ARWGXgWw2Nydgj3lbOU3wT48ywgdWqoSXb6fmH/JuaOY8W65XhFIwVzS7OkG4pjur+ePL7bkD
gnKvgswW2M62093xpngHqUPR+2nTz3zM+9haHBa9cz5cm1Sao79ZFM14pPhNI3iWh4YgXNEtIV16
/47U7M5ghbpo6W8VLbu7C4speGS2jZdg63LFzpx3bixToDuTpuBOQDfoA0qwg1AbBxfX4Ok4Yr5A
C+9Atj8UM2iGUM5O1l+BPs3EOyTuOfC/QJ41RskQHnJYdbhJ6PrGYwplDF0Ctb/PeQNu8DtskNYE
AM0Iauq6fjWwGEGE1l8AwQV1ojMcq28tfc+IAuRtgo3KVMcheU6i6mAOLrjVgmWAEzyv48VG/PNb
xA5aWb+iOFzDKaWIHa6RYpwSFHVH5xKylZNYZuMGgNuALAwm7jBPxZ/faWUA9QnFS7BXaHb1/Iu+
gW4yOe2ZFJ4pFHmk2VRV6/ANeqNu9WcSLWRCiVQmWc9baZ+gL4fKN+pXwTjar7646C8oGj1JZiUj
gQvdZbBYvRi9y7MwVS6W3GBvjvvCYLkS7pQey5r+HrPZAW9756NnJmVx49nepea4BLK81dUPA9hd
Znlx3DLu4VFVfVy4gHAoEuBpgjbf41lNB5l//U/eDHBueiBltFeuT/BKlnnP1EAC4fAwAkiJ80nJ
//Eb0Y9NhDWdpxKypWI9M/OVppXNysQ3L0sikgB6OliB5A1U6UsQr04eC3GDToP/iCEOvvm/NrUZ
jiHXTZcQy5I+K7p7GZi2vyCWTtU8U8EdqzKBSxFIOk4njCbLpdxjhp1vxRcwFjCmfUqw4QBIGk/N
Iq+QhR3iz9JZY2Y3hpsd7+aiDxLGe6cGzQA286iixExl0e//dgOp9YFu2cPNZF3L6YUyQdswZH9m
sxql8YG/UifdyokFdYtiL1QvqYHA/mqv26rime6hG+67Rntm5MrFb3Y/13d4OaOtAvtYn1Y7l4MY
5qw905XckEi4rDk3R7bx6mWD3yf9bYxgOONNsFyTasGQNqTyzPGX6vXvJ6wMfkEWaO0uDjGy8WyD
fYlsHatayTgUQ/lxs6IrHRn04GrFwPuWE4ErIzxVaPnffGgKRHEMCqC2TH4abekZR4oHbzIRoX8O
1kw77fKu7J98PLAyalpYnAClJW76GEjD79J9v0uW178E/7I9f2Hgo4NgqDnRQoL8O1nSACe1wJGM
8rT5sKUCggbOOx67Uqf/N6At9UFrtXKD5LR2KBJKILLwvmNijn5d6c5bst2QyeRdl+xOcYCaRlrw
Vbtxg5UG/gSeB9ozKe6dAMya8bHBvTGHXgjSJTvOX7CyKI7ljaNwut1pZuuZOIGfIkRnaMSkMyXb
idvQ6ra+GKF47e+hPyQ5ZPJwfJGaKAt9ZVojejkuiPFvTtQRbKX/GBxD09xpi8Ac4+KD1MPl5xMJ
tsTfEUAGnqaC5aHoylGOsdkJaK5l86tapjq9tIbON/F82LRMiJfLNpV/8xOpf6z4Z5/i/gfFXsUq
s6VfazeETgYVcquiYQkl1ZlfmAH/C9xgVhzVgomc4VVv9FHdaPxEdrPNwGcgatsMms2rw3lh4UR/
b93qIpj5gK/VZZR6sKWEdPqeQj6JAxYiEdOS2AGPITGjU0mT6TGGMdvKXkUSmeJMfka87F5+uENY
T3SomiaXV4CJtlGJpf3xg9vuvF0bn0L0QPXM8NNPuTOhOEtZOclJxOp0c7qyxaq4UTPRtFw2PJYE
B7NZiwmFc7cPTgDyd5VN3PtKidl9jbJ3qAhWSP1HjXVhQXMI0sI3ww+xZjbwvOM5LTV0OrgC47M4
cmzmfCjRIIeNVWu6cSuV733ZxT/FRLGCSeoChpa17cqC9KwQ8quvuzRRzZl9O1QU4rxBdg4jKXp6
drCZdEaoup26gN3GCDt0ztPsiB8+D15VFJZaBUSiRwabj0Ds0/uI3t3BYNh68vokoRNpvagye72N
cgH8n0rWa0jP44IgzDjv9s4N6v/Jlz4nUb5+6JqgOko0rmbLtQ+Qp8ZAIX9C6jhYBjYOGGFneIzi
ni9sNHGTy3RvXfUgaMIYTnjfEKuhAWIqKWp2IsEf0OfinmfaPE/e0z1MRgqoupvpnIzyVz4WxpJu
qAntkvJub94N+GQUB0bQEAJ7hFyAm2lVWt3w8p+X2Z2GTEOAjTx3cwfjmcHFvfpNXtFaynpblDDn
fJi8NVAGpLBGV/IUWgMuo0GdcuOPliJfY3QZ9LyN+boAwJ7xZv//rs0tV9YamiIY/aW/PaGik54U
MAJR70HgWWJAa2SYCRC9kzYclHp6qWWczvEerPYrMgPQdCweaXaQctNxDsGeBYB1fvseiptZ2t/G
1qh1sjk9wUyrEvmj77AkUoqVe81NwCusVO/7XMDTHp9g03o+WjzLZR/mO6TtYaQ374ykbG4l8VGA
WhwE66FCEX1dfPw3M9/H03DyvgDPyaEseNdfnXu+5rdMxB+CVGbU92sCil7ppXgbgdvhAVkGKVet
z+tPacgO17YiRrPRVPgsYo0p3FjlkahshFS4K+QoLBbC7Y76JwRgnKcpXBmJLrLgdZG0wgoNHG+G
U+qNz+HtbAtqYGOWPHDY6nUV7W6ej3ZWugI5hjqkA3uxSPUKNqHccyrAPP5K6sOHWHgPobCiNe12
N36Q0SrOpsX4KEN/tqIfumk6wpA+zbdqHjKjTPXjun9KJ8s97klu+vZcCYbx2RFNWEaPDDHEVJZy
lKsNY+AsASkFJpDZocnzPskNvceZn5lnIa4F5Oz03we5F6J5rwW8tocNQnIFAZnkrSeWX8QK2jlL
ANsW5k8krv1onQ6Rsgix7y0QhlKUPQCgT5P/6blncYtYv26xIyqYvdc1znnLJQHo1mFMFR6aYdx0
niplNcD6OCr8OBZ9u0B7MyBgjVFm+JH0YKrTP7dYUUhyaIpU6NICTILqVR14GSXDchw6CsWRR5RQ
Ov7AeTR7Ni8lgViwBZei90MHwU8Rx3jhL94Ex2SEFnLkUWuIkiHD8hqw8clh003uVTJy6QkBoYLw
dxeQnPOpGkcczV8bBePuqt/nEHjYyf+0A27FaFF4tTqrH4v1C8WhuJBxuVtWObIzHLahwMblbuXG
e6LaZwz5Z6CQUif2GxzKVLy88zt88PlY9Nao+2AUL2rw9ijtiiHiosfBZbs2JVv0/t+JnEORfhQT
/8k8PhCwsL8Wb9LxeJYUtAKF+zzMvXW1JBp8ndvxxZMXK5qUHho7S8ATPTUhYQ5WVzhooAIUaqY+
PniUjL1u4RGmfKfRDGsoum5gXhp/q+Czj8txhlHyYRV+2M0l8q07PiYlcjXfj/j+jJpabAwbyP3V
M06UHHXcymAQF7tN5VxWk3si3UAUF5ZFnk9N0BiSAJNfC8tVCg3O9It2gYXzMN4IGxk5S7Ktzpbw
F8dp9U7jHXGyVUO+fGgHZ+w/Bf6aui60dswlTdYw6/6CGhCqL8OhDtTfY4WM/TNWh2kwJR6bi5S6
eID8JmVI6bnuQgyt+LBGAuSJxrLtmBa9MkmU06YXQPjJVES+MJJrqFYhe70yl4hrzwY7BQoa0CoD
1L7AGaKq7Jvm3UjEHNvD7lA9a6/QZAxG4mqNLx4hxu3v8bG7X0vSFAu4HgD4YXxBLS21rLyBCjTW
NRWayAShVxVAGLTle9Oyr/rjAKGNvju4zzleFN/mmKq0o8aYQ0Hn9PDT/1fML0xv4cmYY8sGvAoA
3/MLbyo2uAurMWBCU7RpNQb5acJ09dkfKJjlb2HI9/32pYuBxfbq4InP824PVEVn4+I85Dul74ym
26CMRaWoJkDhWzoO+UJMcebVTxNJRfDmA2pbdOF4CNlRbLPlW9DJNEj6CUYq2ttXgAkcm+vjdojT
TlgN4Z6Kdn35gtoVyyNVVVUfZKW6lXGDIJAl59IGJRgKqigQNfcZTWaI2uBqR6NBSvdyLSc8Kce4
xJyYAE3CLkqg6XQMh0q07Xs/vIhz4SZ3bf4rMao1G8PbLRo2aGz02g0vu1zM5pDpcs4YW7XTfO0W
s+zGa5JqTQEtiYnwh2bp3AiZ6jJoxYrLWmz01F6WIHMJ666d2/XC4nuWNbhiRRnojicEC3ZRNu7B
R+8mKlen+w1m7J+UhKa9Z0Vm6bMpoufN58yXKZMB51+b/XeMgXf8tk7NmTtiyJm6Da2JZUA+z3O+
XotBJGaE8/H4cQ4PN9XOWqTKs1n9fPL6P66OBAnikR3UMU4Xdt2Kf50q34MvinA/3GKykfYZfiwZ
msEdfx82wPVjbMSsR2zYObjAy+bmfrG/4yi4THQyRXZLz/3bUCCQpAvm93tvKfdZlSaNm7QpCjKv
bTi6vhho6fMBHe2DThTxblc+eAS/53d80o7QGxdnyuiB24N5eL5LcDvVUPPECQvrNN8gKtbBFJ1y
1KMhOsDHYLBjvoo7dLNyCpF31XFSEF9wQjbRI9ash8YdXbe1upIW0wkvSnUYVcDOhjal388cJsmi
+gxZKyaSszsmp4EWvzF7jzYaEk2ED5p6zBKRbtqvtAEvzFXvqp8dkL26JzfSI+LpuNxV4mgknWUM
OIO9mKaI7HyG8H5MLp5e0gfjJzBDYCSNdOVpuvSFI3F8pZ55XUrcsRmCC52e+Vp8R/flBkthb2TO
rlAWZknX0kA7tYFE6fc/HVL7KZIfsAQTKg4qr+rW/pmdwoXW12E7GcuG4z66IIrvgPXnBuMGJKd3
7Y8gmwaqEeQ08HkZz/9JUAkwDTQ/gVwemTvpED2ylZ9zj2VvgMJDEA7RsMOXe8uIpXULsKluV0jB
aIdG6wgHJwUGLHzaTlX/rZGJOnvEiVsB0UoRCbIraZC2Eip7a+xSgjpZzYMyRJ/NH46wQakqG4Jc
9zbKVho4ilWJpfo5aaKIsmT3WyiUaZOlPaFY7w2gqxXfYIt+XAq63mfWwM2+ArctkHvEUIq4Lwtf
URugm+BqaG23E1UgHMTBC30sCEHu0+T/Ow7vca9q3hr/XmJbOEwFXKndCXmp/dJYL4uRSRg7lqft
B6Haj9sU4uny5IIxR+6TwEFO744cx2azRGVAGkmSWFQ0pZ1Jck4J6PhdOYpQUB3MZVAhZpIK71J3
PutFVZfgjMa5qfcjqWQmveZig/O482pvik8ErRwUIuS2V3Rz+7xzafo8wzWCbiql3gE8+CJ/WHMC
TF2ZxyrVIbCHOSuD87yMlt0T56bRijAvI6QsWGu2iP9zxqCtU9KsxKhFLa+y9UoIkTNzzmrajZBn
EQJRcOCLrVpuuNVUg9L6QyXGv/g0Am7spGSEbTXWnI125cGDfhnj5Mch572EwcVVz3R7VHOT0TSb
n/gjA+V5EYAoM0Ih+auPlNV6C9boa144mkaRdurOXjcXdj4NLbqli3SE/bn2cDHGVyJHPqUfKli6
9gEXb7KVTYSJRe0oFcyE0UhEYR7QKEvsrY3S0ERDYmBA4XuZH2ykhKaR+bqTNFCgfQ9NpNGspwfX
Hmlxbl53tdiCi5tR2J6z+uj4Gy4ciFzIFTdBMQ9JR5dFYzSs8zAW+YhxqQFxuRpJMazEHudUqepb
kLu8mAM+tnDpQAKHbZO+f2vik8jjDPF7WEoh3gP/RxPRFXdlB0KIWcg8gZQrfiKGIYz4IP1xjlUM
JlBwcwLWZYzWdoJuaSZoG1JGvXUwQi2Vsl9aBfqPmTZcHytLzWMmKGcadbw2Q0uGp84lxaXkIzOd
pMnmOwEqkzhNYzs4tDJp05LyPyLEMgZ23VEXoajM80BS2Z3d1utBz9bUEItR1RMcrU+0CA7iXWrK
tsiy1zYaV+2jHM69swSAb2V0LKcuh67jfuamFIR0xMlzDDqP5/JjnF4SqpscOLyRpHGnfbTpO5mQ
p/vjLuUKPCBfmxwTepskq/gXx7XddNnj8MUS8+FzXNEKNbnZxSAXtda6V6v0bZjaI42d3NUHFiuG
JBjwbcX40PjhGlfsgM+HdwOICD3jBO13IEAffYVvNGjvsdFiZ8unqRSaTSlhR4nx+mmd5kIUCXW7
QThetRPBKnb+2QJNIa/FBhhxAMTc4krl2C6tSU4UkA2TNrH6Ur2vZ2yhHda4uabQxoDTWSHEe/3e
jCh2FNj8EtMwndEu/DZhAZDzRdLpFF5QcHJUvcxyLZij2Rx3jOs6gZZrJB2lloea3obh4TYMTE6j
r5KpMjSNToBq8G1MKMDNvLyy9+r/TQybSez9OQLkrHfbKzwniYDo9rog1vv6HSz8nvCHcytRVvrm
vLBbtLZl64y2QlJz3S81m6zXmHBPS7cFjUt7EoeAgb0ZT8X3zg2Fo3X9RgZD4dG5h6lUbZwtERcx
TW5jaIHQsOWBzib9s5yZaWu707aJk9UYGhC4HEOGMn2V4/KG5gXSH7sWjlugiUahBzmtvccu3+Cq
2S0TnhtBdKrDKOLe122Eck16NlN2Suc1b5l6gzZVuikIABzF40j3tYyO9nmm7Q9ZJRXWT+JjOHJg
4QhB2ia4zHXSCHu+HYYo8iG0cPFkizmxoodQ/dXIoK6JBccWFkgUIdJ+WwfhF6BVFM40smDy3PEm
c73gtyQ1CiE7Vlb5K3/oTm1x+ACPvniyH55AIe97z0fcvMbEu+eI11zvvNcavChzOqv1/Tvowx0O
XncHnEMiOhok+uv79M5nYSAecBmbJYqijcGVy1ibunk5muPjm3hwaYy1cdHUocngoT4xUwcS9fxA
Vcz6FzQWQXKJpDbcOTnaAXZXLPO87z+va/eZ2nA7BLNQ8T3UkopB8xv1uZYHNi0ZYiP8s1kvd9wa
2InTVfGbnB4HhcgUOYZkwfavLDhTLyB4kaWsH6nt8TILRpgyE5Ub8tKRQrLmX817DEas3tnTSIDF
5+IA3pHFIQi7tkOi1xAqk6kYxkJQUU9p1k4I9FZIQOxEVTxwj9Q+leh2KFbTnakoncWcTNIaFZv/
U+3fMulnocU5BOIts+HANDYlkTVAiRt5hU7GGP3GWg6fqVtm5nkFGNMtN3ZdGmK5PX4a7ePq39aQ
37aodHxN0R8fdDbCsRoZ0IKwVwVvaEJUXgLW7h+LLY4+chceHaf+gquhClUQ/NnwSZoh09vZqW4i
QyWxCmei+qqqzsrfLbYB13r8dctQ6mBXtXVkBD8Ir9gk1NsPhf50PdydPn9lP9aIQCMfEbWKwlT2
ViicMDYfnfcvil/WydS/SL32GlxH3p9IaSo1tUvT3LXtVGpknonFbUYi5ahKt/AecLQEh4t1w4ax
woVRB4ZfRsnM+jlqH7TLCAbtP9j34t/CUANi7Y4HuBzTKIYDNRidW7jd8g92Ir2k5dv3IAXE+uwD
cmA0WOwif0Z0AIvE5IDMbftRHptKzV+2xJtb6SdzpjfIYi9NQM1ik5ePvzgqyNqUpRjZywTWMgWq
6E0YnthjEKA0XQKmjrt4AX9VG7o4rKzJA49eaxJzgy8wHn1jxZVggiX+/ZFX2oocASMVSlDH4im1
y5YpmwioiHTNcE1Na7cf9VViPbot3mTnmFc2OXyv3q1pHEVrVUj7JiayTnA1uiJjdXa25FwvH3Mm
TyNO6VrBoB1TTnsu/zBEzbyVAzoS6eV5aY1qnq9AVBaGoUztzHKd6akrNm2kpvRJFOOCVdJtU4OI
bDP2ybaH/xuIJQmKnlgMfG3GCdh/jR2xlUXXsTH7egOcYmNlXt43apFplVbBeQ/l5FFxo/QsVYHu
7yRMW4Rvtucx4HlrRel3CWCrVYvuaUjLqJRstkJknaM5a6lhj8RlBAgB/Z3+eoIXIxPuujBM0mHM
0z+2o1KXQrYN9GHwJvwVwp6goEcZJK1DK81DKOCcpbXNobmT+RnZXwLjDp59c6EkhREqKknsU8Sf
Nn+qAewXcX0EYDamiJpoYeVIte7qDwTsYYjoheBEGKOGDmxZDiBphIZ5S+3j5GPg1OlZ9yNFxmXP
vfdl8ISauo7or8KCrtKgb9vfHu6TgrTZzsfmaNR5SXsFeGiZOmQaVZj/6PD1lhs2mY0l5ms+lc6J
SlT60T1ySgwBF+RTfqR0bY53dIxkO8TUbiSOLDclUi723MMTWkpaI3EfaBRnGg3NBXOp6OkxTV9d
oP3QgnqVdzxYbNoiQTDeJzFb94t4BW/umsa8iDE3u1L8l3fYhoDkP8KP8T0uLBKnTCobE3BgyGyZ
JK1CP29r3Bw+0UzmMkB9496m4mGr2TpgBIRnG65crZ9499WY76lEGpH6sRLyYPhe1ur33bVEuhhh
kL/g3RMgXNM0Ew937sHeXv7barTd1sVh7M61v/bF0Tcguoe/dZgxc/bRITbmDTd2qy5jLquKGXNF
Wwd1Xgc/MifA/PL5pvsydxdTLjoO9haAA6mCoxKWcvFURpBRzQeqRg5DQbuFJpnaBtKdp66aB/bg
nE56pTsMHKe310CAnLdJ3/y86WR/ctLaAMALt095yQcVhrWjnxksY46w+AR43AdX94ulOwAG//tK
pgKylJOdxoWQmuSXCn8Xn4Lvm1KRnZZ56TmYDQklNVQ4FIi6hUhANOr3BReQ8MDK+YH6ouVqvzLY
xYrUqQ3bOL9K+RyWqf7GdHqijvprugyPuIcI2kqeQytU8DElV8klZpwu2sJ3ni+A7tyPpP2gL/Vc
akS0DIccqbI9deDBOQEeZillwFS5dGzKqWcC728ejyDDtL/zTBwkb0sc4REQxtEF0UGTcaQkjzrs
XPFaK7d9xyaLB2L219LAwOH2KIf+/ayFuFQUkQry7K2NRvDMSVt3GsQsKFtLjcpZLAT4MSIi8N7Q
T8+YRmAZ3SAphhAuOHsKs6sAYEqd46p0yti6m3K8GTj3bYketqNMVWFaybHktqXfkzHhBOzPBTF9
iUasm+Gy4pyu5OaYi2o9oUuYH1Z6698qV4/GGFQPjIoK9scNXMznjlZgVEZE+MlVCOFq+Wa+fb9B
/ywgJhsUh+AcnWYCBXFXYQTExQVLbOtu8Rx8v6L4avpqK6jVxfvO5xtDg8D+2L+mbl5FLVfssANF
2CoNymr3cFSDlnzFQhdRsTDOmsuQhZQnBNnuCKqwvnr6228FqK+KGX1Tf/bv7ibi5I3DyGt1oKHg
1iEaVku62NlZG4EhTnHA13+N9CFGS40LzVNRJsKRT7VkhFK6E/Y7vUNtP2ddlkS5EfpYehJhdTD/
6xnZCrmtmyw8j/3aZBOrF5CNkehyXk8QkiiuLOa0WExL3QjR6nllWJo/h60acGWq0PO8rPZW9v+R
DyfC42rrmzFhZZWiK2V/8zfHMj1RU8Bezip6ku3tlT89l/vUGKz7LxTT016/7Yh4x7e2m1BCrKgH
W8gOV83xzPVJ5cJ9IcTmCpjzeSDFumNCt01WIjlCaSIpn2D9lVJdwH8B1NEU6ZZD9RPUeD37eHDq
LhSsvMWOZKjzzN/3+wZd/eyUg/yRMnxE6u5D+gmhPdfD6/y/CkiAD/87oyYtdefbcx+Px0AbGNMU
ZZuEuewDAAsksF7SRh2PrU0Nz7fYx5E3qqjMsIstxVsMsdLC3A22IpaDIWntag/gAw1LkH0phprT
XVFJ7tPAwvv6WaVcsbbPHnhDBlrbOYQiDMoiW4UMIo9i6lATecnSTaGPwVeeVuvMlmrvFuOdQAJF
XyTGW6SCV57C5RSjuHvqSKvUwOOzBwTOzaGvaQHsHZg8HkUTW0xMs1mSCX7O12azucL7QxginCKV
ViVS99/JFVXQ92VM5NOpqOsDfvvTcHyd/3mJRFNJroDAbVDPl8n7FJk3oBbIsGRJlAF30OGikjva
zKt9d5JDbqPhArUXQCVP0M8+SkD7xoC8OVCTp1gH7p0umJSLPrdGGAERVd6ZcbdU+dbBJY0s8dZ0
MqhKo0uIuft6fsMWKRKhcQnmjh7wg922ZclOUJogk2kNobKXzXQkDM/pWDI30ETV/uDEZO6l+5ZT
N9dJwQmMyRUt+DD/AehYnW5qrDfHXX15PlqWM1GrClKj4AaAqP0/t2c1gSNZ9JzVaaqGvfSNs51h
I5b5GdFW4hcjz9k58h3NGlA0kRq2zEP147QcfCQ3iRZTdGM0XK1jrMJvfeiQfONO23x/llDxDAJz
NHet6FkFn2FfHRZ/Gv7+xSwMGEOwW3kGrawT6OqTa5OKkxBQUEYCL08MpbvcC5AV6oOX0Pq81PCt
d21qoRsvQAEwlXvsnkYPXJFdVB9jOeJEq3Et/Jue29a7R06WSIYQxcyuR7MuS8wY1Ocrkc3GRbpg
9N/0DTQUmbpdpreBzXf1aylVoFVjSLAuXfL8d77IC/DdVUWsxc3RfZ/F1Lo1vWcvvEyh+WNb3SmO
TxgB3LOu4GNKvz/JMLlX2Pn8/YeMosJajo2qJEnx3+g25cAvx0IQ69Mi1ZIFIK4dt2XWpaFQXE+3
/KtLj9MOQI+lgwjQZEOKxNZcT7nfEiCaqQuESIijU0idgg3F9jP8cckevSbvd6kGVdf3caZq0GPV
wQeVTRxoVVII56RAPGoWT9vC1Ow79siTKvxTM8S91aES5kz78R5KbSb/7MruYETJYGfX8925tgBI
LL7EGsyCaEYlx/XiQmwj762HkGn1TP4SiZVP8UXvjAacv3liq16lfA8SQK+Fo8bkFqcN+7hE2GOF
IaRy7rrJR1xbhR2HDqiUQ5d9XZEu0GzSyUZqWevvq8hhzSqxgwvrXzpQPzdKoe/Sr4ScHRkLfEmW
s6nnp7SD69Boa4/Fapz7YrKksaa8w/+ZTrk+mMR1d/y8VBtRorjoWi1X2UxQtPNKIP0sTu1et8kh
Pltf0rIXhSjGWeLEAKjRj5/AvgA8a/8KB89qHN/ejh50S+4h5igs9yBJUnZytgCRwxhdtZLqZApW
hogb8YalFATV+DrQTW3xQ9busUP07uAFesG6USKWng5NDisTHYenCFORLh0wioT96WSZ3fJHJkrW
f+V3uIQ4sGYqjP3++rTZPjIRPZbqDrwC4GvlH5JEY+WvEw2jaZis1aIpL+/03iAuXSe9JKuvaXWP
8UfjlcZuX/8cnxhrW/2UJ7KcGaaj18nC4FZOUe241THSYZRQVB71+CcnRGCYIWqaQKzgWal++8m6
uitI5EcSpu+0lqr105HcO8DtGKUCffqOceFwLYMf5ab8xx88am2kPaR7gSh9UnZToOpcaFE5W+rQ
ovn5bb23viREFr4lM+diSxZ2LxyMmqSo9d6wTcQf/XG5uhfUoo7Rkvg9KSD0LC2MwIplE1q9Xvyw
jBNdD4EWY7jEjQPfUTf8rxoR/+daw+0SbzAdxPcpdy/ZKoT0QxK9+77Kx2D3HTdZO2IIuWJcI23F
5kU29WGJ8lmaf5B3GhdfbZJwvxrnvkqNCGJiJ+SM5Jhr+HIuN7N2I2SVnxQkhY3goiJZWUe7sFch
6Cj2YdTxb8974KO8EF9Np9nSjjbHEnlVVDd1BuNGBAtEt1O+hyQWO9c15418n3x+cHWDDpgk+4/d
vR1JW1Q6u9vuuufsmFAMxNjI81Ih/q7ozSImpArtH9p8kppsfNZFuAYwuY5m+gWv9sFmndKwHp4s
2Wu5K3/RSsBDVoRvE+mSzS0AtsORGR0MQKbVhKxU92YNcFH9OKod7tYUlIa3z2dUF5EVD+RQ4hFy
CukbzU/+uui8Ysh2GEs6o8JrsfV10wQ5nZHjEM8kFuz5q/f68iulBMxRQ8uhUGhOaO9DF/dyfmmB
PFxmnTxf792jzqHVlkwLzFO9qbsLO7207BjnNbvct/1vzFJqglC0Fbv+PKWfiwEFwWsGrL54U6yA
ClSlevAPR2+y5dlpduALPcNOokA17eW6UgWXzmnmrAPwicqpc7QymhgHp11LBKOK1xDdkYez15OM
0WoQ4BVq0a+g15XYXbHMoGejDBCJen7Ky4uWXZ9TJAluSYqo5AFNnL8WxUCTdMrAuO94aA/G6u6B
on/HUs6SoBnomfIEvKcv508xK7lWaXa7zJO6HnWuk/6QvQCe1UQf+EoDSBCBJMiQPR4uEL2UHyzK
4iZjSrnW0WnLSw7GbuLADWD3QVCt/hsFod4OyZMcejrV/jFZkATsHkuMStIUfbajA74rLNt7dgSH
ffCSxshByNjFQTDv+ksxSEfDtrszq9dCl72fJWVYPeldG9Utcdv6RcLXpJKmPCFHYFkmZlIu89HQ
m8VvwfaURftPreAzZWwbSuapnwMgWDpQ7y3b9nHUB8An59WzQU29wQTo7zFiEL44tdWJqv6ntV+Z
lqouFKAJ7Y3Tra4dRpOP4hpUQRAWXdcViqdwiHFSYcum1agnt9R2UnZ3ihnKgtHTygDHTRf/OSJA
Kk4QG5MwPeuC6qAEjTJB32GqiC8Vk8oJjdViNbHVvLol7sSy/43EDGk7t+WWcG3WXcMw2IzKDmsC
5yuRakrfHjQqYBR3qTJvjLp+q5WUbxmsqJIZybrwBl4WhbvBTQT8wkM6nQejCHBq5wrC5pNRWOnU
/8Vd44tnV0o50sIPCubGTTZaNWJxUoKsy3SdMZp99mcrzw2MP9hrCwZqA4xLl+go3RFCcHOhxKTO
68c9CzFs5enfZFgc+CUdgLwmwxn/Utd3gNhPpE4uVxRrU4giBVEqh8M2tNMH74Zth5I+qpMQy8R1
RTLSBUoeKLLhg5oxCtzlCj0RLNp5BG5bLmlUZVu4V48EPBNYVcRya+41S46Sn5x6zmdYgvmunTqa
OyE2wWk8r+U4c76ZV0kU8NddVwE7ELK+b0BkpIfS5iqkj2axwX1j969twvAL7ZQD9/mfj9McisYO
AL4L2C4uY6PRw8rU7A7Qct4d/pG/C+VdFfLTewMpHua0W3uHnJ6zU3KWaOupXZdOJaoxESGxwtq8
foReSmPjjyphXrbRwiPV1y6hy2pO2ggKaEFn1hBEzQcIac3zgGWliSJnZQzphujjIrtVf2xOXBtb
OqcaDp1LPZIHOA4wbORLd5b1iSH2DVLwp02iL2izfYAw4o2paDLyhmu3ZTnCYHzwpo+3jURyEfmF
k8JPsY6IFQG8i0v+K7ErqnpiFQyTqN59j6qJcE+obzwZ5fdb/tbx05M8qfkrPFAw4rchIGW09L0F
2wDqSHYyLffZQfR9xqITi7Q6u64qhFVUsCUyfWJiKk7OublzahCmKMuV9I/YSQU3CvMQ4Gqme5+E
EfBwiIYTNkjtigadtQF8npcAe7im+GbyNsVgrxeTgllbgOX/rr5MhoxQMZ0m+yDTwHHZXWtlROVz
UZTY0l9KwLkzYCSndXFpArP5tXNqHUE4BxaJSebicVZ75rXoJqtK3YF84JiIf393RhwQCknbkd4i
qXMJqL5koNRTzVQ+u22nNdQltWhQjJ49IMKWWJdD/aiOaDQKT1UyteeDF/Sl+3aUpj2Juu/Z4/AQ
RCT1lsg9bl9vW7d1WJB534dUKWVnVg97HMNVCfF3jgtZuIAerNs2wmdlZO4CHSpV5hECZ2QbW/WK
4q+h7GsBcfks7mzs1XiMg5De7sEg5nPZGJ+38aVI5TZsORB7ekVeMrC9OSDMYnIF5DGA08VZYaQS
Bmq1bMYEkOHYso+0CU3h8NEbgLEk4oCsgfEQflHC3qMqSbW/vIA+/84FTZtrBKi3Fra0/nOkgFSa
NTTjXcql4lzjFFLUxG1Vg9AMUyFaCkTDMgZM2lUh6Ud7J+BHDwI+1qRGnTb/E2bmMZp77dcpfrzA
shTI4CU63ycE3OLlNPZlKgq2FS3Gy7ZNvxppR7HMwOzu+7IGaFk08eWsudzCavCIv0eYt4opxtZK
9IF5VdyCKZoUN5vROqc7n0FIWNIhj5Ja+SGuW8UxkDnz5V4O1gBRZP2L3mw4qicb/Z9izZD/R1W1
yjKlpJWWVbLSkgXybNNBu+2j7fvuhOge9b63DUO0RDOvvgOU5GAsE6qUhX+4702ZT+eq6H4VDUCG
oRO3deTgb2eaoUXxTpR7wCtplMjCRfWQWwdvs+EPz3g2Krg5yVh6djzEZVEbNAKJPDeiIhcObh1q
l8AKlOvYa8VwZ52P3wiCrvkV19chubtsW+ZQHM9FnOHaFXJxiQdu1da4BItygkbf4oizYQlt5RAe
QtiN4H5zvlCbF1XuWvX44H0qH7v/0X/Oa4kedS7tuWOOWfhAJ3v981FCMhVWYslfGBaogg3O3U3T
yRyp4KQhziyWLhVX+Q1Uovtu5hTGPfsIq4sZc7y6RhY8nDPD3nSTm0XIBJ+HciuX5GmfcGTjr1BH
p7HBL4YiVCZcOR4AsUGY5brNDiytHDQmDAkHk9Y7XUsKETNMZSN75jAlgdKYl1P9JJ6D2sD9pQKs
7/Om1nw8Qk+8WPH9umWzVya0Fkyimq+8L7juWzWe7gSBgVMY6zEB6tz/DiM6bJc7ZMEDWFP9jg0L
fryr0j5nIDQGeJkZap91AjoTUb6j/VqwZrsUpzmTj/uzEagqRngJ0j3ifwAicZO5ebMzInwzOZgG
9j8j7bPrSUMePh+mG5gUd070jGrEtlKorZqqcHSbRI6Dm9WhRK3B+wdNu97vzyMfvz9o9FLwgJa6
vs5ZoiRnMApe+WxrpCvRYACHw44e6qEq9SoLTnps7GG1P8Af7kXhPmjms5rU1nKUZq/HPpPwCOP/
akgrSNm4zJjJgVdwNPYEy0AeDwNiDtPZQ9vPPgGTwG7ReVBhtuGsb2N4sQnIWcfVrW7nClvxRe5l
cbru7x09ecLSYgzHzJfIiASdmSUWpEW1VIidOOoTk7HXgbAquOzAIptM3aRNJhHzpzDldt2NW2vF
KRTx2IbSqzthIPSoyEikDlBBqxH7GzpwNB/fhyZLIUhjiGGrpw1nwQrl0FjadRZTV4M2Y+EepkDx
W+EHkNY7xF37aU5TMDH8LkyqZSeaKeqvUE9JnvRg1Fg5tC1l8j4X1PX04CTrh6ZJBOcd9IMvtp3j
OfLPi/OlSB1Oh493lBjtVCkwwqHAL78c2VidAxWAnlLv+kiVvTa0xVKrsxjWXaK035WsUgckFG3c
ODyzIlSyGGveBc2KKy5hDfq64NqSczR2hhVv5BeblEXRNK5ZZ/789y337CFLUJRJPrCjWuhF/lIW
fvGJNjIFYY25x8zvkbqYOUq6YvEGzvB5wEP/bPX88pjwnA5qP/AWZVAcleDAGh4oC9XpGsAnrWPy
EsSknm6EE9g8tjcYSR3582aSe/FOUpjy7R4sGHHWuV4lM473IaXQtLusrYJnNNvuvI5nJ7uYQRzK
Jq1fofG9w9K3/IwZzNvbqcmYqHa5LU5XkOViKrxfNAW40N8J48MY9KDcszCi7aRwN5KcvpxAmRP5
/C6+3M+lc7/SuMTIbs8GkepnohPcbFnQRrfPwvSglS/tFYywiF2tRYgEqJa/yUQN1ZCSJXi/bOzQ
GC0W7ay4GuSYpOKrLckTyD93qFAFArTk6OKCDRrQo84zYYl7D88v9Uy2P6J53e8wucnsWLwLq4bi
T2npH5F9QtggGm+lmrXK1bx1pHnNhzhWKHT0Cd38lp8l3FcgCjNVYyYuswIX/lxJmHnO4HZi7xGy
CQSDXHg7fRmBr+6VoZ9dDGBhEGgtNNNmL9L2zjNj+BYyfxW8DvWJd4GpgxaORWpCH7Ll93d4M0dL
rpWJFtTfj+iSKNop5Er5xabL2bMxmRwWZNy8jz611My0gki5CMKlrXFzdSGvZ8JpDFSB3DpcBtXJ
uNyZ2eaSs/jWjjMyBDRhYP6wLKkNAi2OlL+2O9xpAS+8NllloQlyNs0FZrE3pCDzbthWzkt1dw2A
b30toDCxV3Jqi3qLkew7R9HWGNJ45It1ppMF4lCmRcxRq6YKPvZ6XnZYGIyFIn3HqAjgqxonB4kL
sg12sODklG6QWDzaEBy5KYcOeZLuqnJ8PLXQs0UFPytz96D/GCMa+GIfEEcSX2RKJ4uACe/IZvql
UrYnnGCKgyuKOh/zBQ1MmJsC4gd/zWI2phGEeq6w14zvfpf8h6RCaYGmEJQUSawCA2LAz936/dFo
jcAPfsbwnOWvcudmm2XFwmrbBuTrpazB8KsgPU5mwlxrP0RpwPhbUI//JMn/z+nTxLXN0LPrXfvc
n62Fl9hKj0R5nQviO3Ii2L1cBbaaqU6j1VtIUlyMc6EuXRAD0WFK7WGEMRLGNK9dbHURRSuHp0Xa
e7O/B7oLhEhmTeuBtO9xTA67gG9YEEGb28QMx8mVO6a/E4IBIT+IfY7m13jA6RZle/6HB2QCuTWF
OEzQgGdq3GCSaYsrgh0H7PB/wsMAwlOj3ExkPR7pCa3tsPHhjIk8pIWbtIFCIcKHse5ux/0urk0b
NNsbfXaBhc8WK2/V0Y3pIjWTAieIlbh6BPXX5Ln9vU3i5xw0P9HIe+/j4XN8RZeXNfW+ltjMmpQ2
ew9ENLIa0zp80q5SnQGCrturHO8YKyu5J5SB4/JH7jz3ahM1CRJwARBPSpNbb0+8jHDudinfuLlA
8qAqY4CAnTjS3LxKLxcFsHWj19mC8iAgttVYd75tNfouY039AP14hZWTX4JVnN84U1UYDMtFeF9p
mNjwtKCH2yrXctq7hnvPjINDxBUAeUsDhpGbpwyhrDS5r1c7kxZ+uBu0OSoIfQCeYhgRg1b+fyXR
29NFdcHyPheUrjY51OLzQjLxoenjiZGfEuzmGG7iqaFfPkCbV5Z5I73jdyoGJYnb8xXWPihtwZzt
IEdM0cY0wJM46zH7Dlmzt433Fsizhhzg6vXrsiGG8+6CeSSUqhQ33qA7500DZUVNw1zPH80LAqF5
GxL5HVDPjQ+89TUpnZjPon8hLAVCA1oIEmknd9LHxK3767H6bx0KpKKK6h90leCgvKfQss0ibqij
KmEdSIhBARN1N3GOQW/mw8FAEjkunS4E9clNrtcCG7a/kboKZ+68WKgHTyWbdTUCwTRvX1ADddwU
7/9Ama4+M3fB/G2GLVaZ5rJzfRw/CKhomoSTbJwQeo0IHaaxH/PjfBRx2+jwZ6gdMgF/WNovLxgy
pPhmKbbEbcUQsPEWEynQS2jEtrqTAAjsr4KwE6Wjexfu0qk9AeTZMbBA/D0SUzTCwiednvc/7PYb
68Ap+E5KffItYaZdUUDDmD6RUntcmjVAL5WdxnvRqNtpDPJ0PTNqQ1kC0C3b17WKi0wcRNVL7ZyF
lhqrK6d3jM0gtrltyTYHpphD1o28t3cYjerceT0JLL9oJ19FB8fPda7RZSwFElEB+G1SRyvI0dNX
unBs+F/jph7pK2bKYVLXQSBoLD9YkTFt1zn/WQzloUY636vHhyhvQUUs/XJf0wT4V9U3cOiSdSik
3Rvs9T7G/JdXwh25h8Q0U8IPKtH19HfDOwMqf3lWyD1bEmXOnllBGMbIYnQvQ9IxMSwB2eIsDS0E
7x5F9N87nE+EXa6OvQELNqI3YPI2v7+Q6Vso3FtFw9xpQH5tPrfSnS42phhP9S659uCWKCeJCYFy
SjsIh8ptxB3/hZ19Enb0fG3K6iI2mCBn04oKrb9TL7k03NRHgX4YhWU6xVvlJoSMLhNhcgI5zB//
4xSWfQUJwDrlEEr3RNQk5IfJg9frSHHEAWipPXQ4Mzz/1yw8+BVAxbFyos/NHQ4J0fE9CWZFAozx
kPeyJP1caTYZk9cms9GRVFXutF6tToDaoQ3xs/q8saLv5QFJmU69jhCMTPrVMVc02l7jJD/C45uY
r8KS/+F4qFhrT39Srgp6Ah3I5M9w8y2/iFUzvDf4xTxsKq/rKRqPBZ0SYA5be8UlHMsMjxhBVTjP
ZltFGvpBLw8pQBtaCxqSktpRKk8OABLtXFbdbqZHfzK6vYDo8yBUiM2M8CgnvpwnvRS6WdI8W7Gw
KEk6VNA/Ecax6KrQryNKng0ElNEsa/SpRQJjUBZXE/cz0AKXYEWTn2IP3YLQZ/wivG2c949sP3Qw
ZKR9+o4GUa41VIbdjP2efUSjdAim5ZGLyFOhOlmh0DcLAScWaLBFsfN9dproir+9P7Tv4kUTv3Ah
kgEI7fmqMmB5o1F4zbeGvDMbZLmtc7HkjuRK0nD+I6lfKPxEClAcSwLBd35nqIIsQ46ddOUjOQ7P
3V/9b1UVBwPy326AyYlvr1jYevBVrup3qg8R+pHKHxR59n11oYMdzyxT9Y2WOfpEVgPf+d//he2Q
tPZNDaZbmdAVnrAdNWYflF/N9LGVVk64csuhVogNgIj2SV4XdnK1yAYUEx4gYkX3LWkDHN6wZ8kQ
lDp6/fT7+ERVjGhJRQOhOU7SBObCBvGGir4yjizWp0yz3PFbQMfN1vFWUm9SBW1ZY/c7Phui43+R
2ch3L5CBAQO69dhKmxXY5Rxxm09aVhXho1y45TvIrNjL/MIY886QqeSsaeNCgpuhudc7fJFpcrqt
PC7xE3bd6CDUZ6taiQTchgBAbIY+1n/KoE7fPuoxv5alR6Fvv/m4+YulZ6v9UqqrvvUAoreCCrEQ
hA2NlHkrXzOZ/z3/cOkd2SdcPhMBIXyTiLW6ePijrlQi2jOBk48uxe7AKfVPakawwRV5YBqSVU9a
F8Yqd7dTSH2iN2jZL9wbX3AoRBIhnTj3dyeQ+fO4VpMA4DlHM5bcj6wXHZ/2Zhnkk6+YJPljTymT
e4xMEZRaWt0qD+rcojkvEgZxShQA5uvDr6dH9IRqEY1WdElTaj3JTCu+i+/2LJO5/OrGGn1FuF7e
qJFM3YQd3Bhiy3XjLL6t0STCfm93khLCp+HufwVDR/GFM/tDV7h9xPcGEcgjCvrnyTqre9MI0f0G
zJg4opmiml4FzxZlnDWWisdv7dU+EianGScybQHuQyugrdn59dmj+RwIUtgu1ycgx99cGOUfl0oz
Zc1kpifJmFik8q6NusYh6i6koHSqoqRaMohSz7neN9J5OuZpoid+yNPMYCXUkSnDwRORtINZY6PK
oGgFe+CNXh3shy85SOl7QrY6jh8brtf0pBCCuo7DNfSS4XVpHzDw1CuHV0XfGgO8PUCksRCrr5hl
74qxmb4l7tDZWrbcPPcq9WZgnsl55HcmEnThzDPk848yooDrHjwzeEkGDgzb/lGpzqQFrCkTetuC
5jjjQ4gzkTW/wGjt+pZ4YudZeecflvt3ZYly4E9lNJQFL67VkC1P/mFoRA/VnQ3gQSO517j9hYX3
i3SclprTJlcnQqROUePpHRIgr1AtRFrlRdMNCNbKocBMwXYLJajCZGF6/v4GkiAfyqNlTAeRpD2y
Tle8+CB0ghBCD9u+x3PgGP+BsRF8JDRmWebC+HKNENJpgQ8KkWC67ewAMtOKhBiss+Jyd4Wyj+2o
TZhK5Ur/qb6Ei/smM6bMxpnwaXWspui3T3qdwvXHJwiBi+tK0gh8gP4oFG/bmil/Nto5YAJumv54
cOR1BmX8X9luiPxbypJemqvfTTFPHRue5RnQ+DYazQEfRJ0ZpX17JIZf3RInHRWt/5WnF5+N5ckf
ZL6vd/o84VDykC3iyDkddDe2YJXUwY2IwuUeOkpYq3+h+AgPzQj+7o1PUTfe9tq5Ymf5QwkhKJNT
kvSPKrOtG/hYPJTKFbr80JvFev/lMlCPYaWrvUQO3ebp0IlfcgY2UWd9V6DBdj7wpwN+FGaVpKdD
h8REg2p61vSCXjzGcMi5IIdqUCEXifMeWj2hzOz9rPwhOr3VWp+T5a+cSUaCdWksugYIWUk1MrlR
focWVL9VvITtM+PKGklYKbiFJVPSJYEaFaWkT17pa5erAh4291bjt1XQB1Si15YX6hsh+4mFjJM5
QCLZHcfVOOj6ZSJjL/4WIf25gE9iAMQfSuCw8zDO++NbeicBdoBQNSjNMx5AqU4tD1Tfu5LH8r87
EROtLkxjJO6IcQrweWhYQgNOxW0zYSWIozOV/A5cdfA7jwWY7UCYgtexP8sDJvTNXrnw3DMPxH2K
piAURu8ZrjCUwW3bjNThtrRGRJgC/+wG7DiQ6IltWALw0iPdRiRS+DLblyQhXNM8ehruIc8xaJl4
Bj58Rn2GQKSvJE6N1GBSaL4x8z80iisL88Lb/LAuCFnhtbr3Fi1rESFi47m6HfowYKErILXZh0Td
EI4279eb59AVSVhaSQIfs4CheKOu8H4MULocZihgW+VtmMf69jF75l1bc6tjvfyUaMGzMAvKMO9V
E2c91RHo+aoNzbQceELrY41MYe+3uQ97uVzwmhS8IVyaUYexwQF/U7xhFfsNfE7uI6T368nF66EO
zwbQT2eYxtNs9ExYAIs6G0dXW8g6MjfuU7mvBF1XUsjPHnHrVdRnbafUBYndlqeaevb/JR3yA8VQ
dC53bpDKwPU0CewBV7QMDZkZoCkaxQVWyugFe8gowUBVfb5g7knNFo/82d98hm47qX0R8EEMJHjL
5bsAb95j/dGxsYntnntRmYS6fAsPdiXD9c5spTxT0LKx//nNGbQcYrOH6bFK0NpJJfzMFzrSiFtZ
VtqJuZaesxiAIbgmr0Z8De3TsfDpC7IIjhiBb1mbQVCwbFctxWVg++Kldq+QYOYdZclOqiPMnbaK
ELDOdPr04d1+OLTSVMe7MQ0lOHVtEiTi5EcoFU9igqY7g8zmoaFnoJ1jqI9UMSSTarVA9eHoDksc
++MqYorqZK1MQTHX+OPh33VFxW12Ud6PkCidqP5KaNMZ8TqLaOij97Z0ENTy5kscZTmYKeQ1TIpv
Zt+H0s4HfZSR37OT/+arktmqbTyGWcQt9eUw4fAvEVHCT9ke0QUmf7xe4cDAJP8IBOk66P3OVkP3
JXuwmh1a9z8gwi8R5kIUamareJgo0F9fUmvsXGkfq2f4GBhbdcX00KRakWKQ+8uWh0YmJ5zZ+N6H
+OHd1pCbsrkvAPdpfsiHwQaqdPUUTfLe1wLo88bOyucnGqF0LUXh1lHrqfosV+ijGvKuQ4srzCv8
EswYjMf0a2aXfbvYxtPDVD/VFTmvzjY3G5mNZBC3EjrG/fsJViVXUX1GpFnYWVDULnnGQBHMQq+/
ZNTaiZuyfzDfAl+VsH5rksOED+n8GR3fxmvfU4ZA6dCj4Z2TJDp+8QR7TbqCHBUKZIn0V0LlGnPa
VEfsVEfqptFIcyYWr49qCXwkHf04eNPFSC47GrSveIGK2EQVdM7Naj6HGP14Lk4hiM9iJBHKDo5g
fSjzDG+eRlm8fLCubywKULQ3AjRGpnz/1L87gSHwVWvE275xr4hICTDDkgnJg7hFCgDE65fCTYYr
Z41y2YvcNaXHwJ0X3YjT4eBUak1P1P27MZN6ig6lmRUgYldWp9kOOEyOEgh4QWdO1W0WVwPSEdgm
TgQfNjEHWDLy+V8JkxTUGLrKaSeoV7QMD5rJstHDcKDPqkbjRXsz+v71SGuvOV/EHG/EMZaJfkbR
BKpupItaLixUVw8i+72s1Sz1JC0SrHzX+yJ7SJ19iTz4AgPmYyrUuKrylL8gqZpdMuPdOA+/1RhA
dwPXY2PgqBpiSjH3omL29NjyLOGE/pfby4Kd7ps9sMNCtCTX3E1ggt0GXgW1YT9ckHmVpxCFrx6Q
/Ihy7UTo+IfpbdN4G5El1u3vWsEKnOAF9w9xXr6SyM4g04wTS/W5o5QLlgX9GBz7OkvPvdOmFVbN
jB6RrvoO3sCtDs3tcVhiMGUbZR1MRiyAyPN611Ur8KN+IoOksTjJreCzVawj6X81ZNVpwqgtmetA
XylV3HEGKY5WpXjKfS/BomtfmCzQwbjKeQdo0coo+fizjJ+AItWzBfXDmvcJWHBU0nBk9WmIc9u2
YA9fqYbpy/7g7nDbujiOxmF8ZlgV9wHLJNl+pRQnwmYkMQtDmKSFUvLu+0j+txBQ8Cs2HE4PGN3y
rLJ9H7vbS2TuZ7WcFN9TGSc9UNcgLUoNHvkVEHrcs75fEK+jk5gd/BTXikaKmChLIYCJVmylQPgz
Rs1cS8qtRh3+wOPghm3QJUI+8dmd+trR+eTMvra3XxUK2ZuWhadm23PbAy17lqbjXB86s3cCCnSF
pjBXyFij6hv/k5YtuDJXbQKLsmzD57WZpMOaGewPsWybe27S6boDGbBm40PhISAmebsjB4Gspis4
tP/yajBjJjbshHTkLWYHoxvss6nQgssdVv78NbobH7lT1v0Z8T/vNOmJIolh6Hgxs5FwjOlo9rix
jnouifFgvK98lIgKgwyTmAELXddnCuGmhdaQkje+CXhMLQY+H8H5cJ84Pic6zs5KoVX5P/5/ue3D
P2qouDIdbfQKOxUHpG/fcRN+f1ULFMZz9mlASg8WOaRBNHvZ9qsRzLvs97E2wwnCndxWH5pJGtkH
TbF1tEC7KTNxYkfkCyq3YyKzbwZbZ7jBMqL8FGO5u2MMcVbLZG7eePZAh1JthVs2idX1tdf5m29v
w0FoxUVOtwTpUIaD4BeBFZWHMpX2Rg2ugLSabL2VvtkWEh/T9gHKSjUPgNgeVc74xj1p18+ZawFX
JYAqBhViYxrKBT9yCfXCJTSf3f5KnIyvECy/+y+Q1LoONXaIj70heAY+ioxL9uBMuL4HXeHuazIt
v6hYQVbzwHb7wyvizz05F6P9+ejktbqZF6UQSvUyxINjIhlxxGek/ZXMhFYQdZ/7ynla1VNY1zXQ
Wi+9cDXNSPpuTfXf/a7aux1FUC+baaZEJQPbFKEZ1oBjUrpuQC0dFidLEWXopWM6roWd6QUPM5Sl
T70rMtZhVBGqq/9tc0fmjaAZdny4t76YQP7yPCECIQB5OlwzmkTUcsP6FOjQSW2aBUJPjYS98Y9i
DB207AZfIEk2UibSn8j0EwOtzNwMmUrlMS6Cer7I/Ikn6xS2fLuRwz/mzTNYrxkvGWa/pQZSsgSk
XuO8mr9CuFd0ujgBmZfHlX3p1czx3+64qtTzM1YTgzsXORFBGXTbfOVQphYmd6Ymoux3nDxDmh/d
/iG/raOm/vNF3bkwGiQHHTqKYb0PEU5RwcaVtkDrPpL60gBu7Xz56ZDOMhvYHGO3fSU4b0RgTKRx
50qYg4fFvDmyMOz2xA0oTU8QatOtj2mm3fgt61LKx3AazHZMHIV+gTYeIxD5ed2EXyXg1SFRajag
ZgDQWM+uGDdWUiRJ4ANa4Bsky4NH4WQWtLWWWFkkIVG/uxRDfGX6nkHpSd/QmLomSHFagNH7S7Rz
al7y8cGkfMnff6gLNNWrAMeBn9j5E/XjIXoma7G3xg0aUDYmAZ2Kjh6DEpHo1XjUyKiTjDFzKDhd
aFKz6gzmlu+7upLlLF6dC/3K54qW4I6Z01NQmSrl3pUdNBKLSUWE4VhkqoyyO2TwIKrIGETQyIKq
Vjn4sXhOpMhDsRa8jSuGyKQGyAIuDxxT2gxxFvvXh1fCxT1vn36mXyGw6T7YBXj1Sdh0kDuBUVIZ
Mh+89lTm0yUphfgqnQbIzNeLqPCtPcCCO4xUl4WpY6Y5CVglzl2MUqaRatF9Ku7gxfLf9hSFP9Kz
kka4rXbtYd3BAE9K8dKKXvfdYsG1WwosROtaPaO9elAtlHhyF+LIJgFsSiW4c+tzkYLe7m5CqBtB
fVq7cjs/ihUo/4bEL752tAz/x+0fx+PbgrZ+lexVYny7wVfxPm5QLdnWMStJRoodG8pmNpRIaWz4
ck+GguDSDwU+pYaMxLS4aXhlzK6GS+dJHwxHdPTUTy5VTSCQQdb6fQYXeKmiTUan4JRg1ZQ0ANAi
J/YvMrjizumPJO4Lg44JNpXucph5sDIeXOIqeMwkkTVIU8UfZAnVVy+cFbT/CGBx+BqqzCQp6/QF
EaJdPJopiJ8kSvbB6o4zmoCzCWRCnpbRoTC1FrvfWICzCa5r9v/dpgzygzK1HTPVylaiDGfvttN9
u7qCE1CRb1G8zPz2fUJwyU5ecIR3UEjtcm5jabWKAw8X/YyZbSn3cohTWi7ydeMYKIFWJl8E1nPg
7fFQ388CoB095ioQh8ZeoDf6wsBQV/bhvpqfLSnEYOzNip9wQGCd/uPJMcpuykoy6pX8Kib1T5Ja
ahFoJpXWH1CX2iapgFL2XDi02EYU+DS3kckgA0Eyx0qrwcIX6JxzQ5LYh4WreNLFtUXP4UTmnF6c
JoQvN/z/1BqnRcsbXslB/fnKUGDatc2XJcb+7oycyxyblpXeI6J6flwz4T+QDKw6Kqkpc3KQ7pdr
3c6FMU/oyPig0QEbZD3yV9lJbZZp8DFGkJ0XvyIZcTz02KyRG74BeOEkyBuiuA0XiWFi6C3Qp2iq
HRY0JorblCQxIUjPODwmY993bFVgrvcNXZJniBlQo2S5m7dvwkpWYjcjqTvM6c6c30QOF9D5YcRG
oWGE4dunU2NZPbYztTwFhLMstGTJH4vmcLwDNVfPN+52veqDEmYrt4eSfFV6W6DlIsFPvr1iGXAs
Dtf9bHGgvpTnWhCidc8P+PQN4++XG5CYSBEkRP9ijENyLtmPzPKxFiU8w3sjOvfKSZeqB7cvkkrz
r5neZtBfs/msozhluX7IXkEWQWWcWIsDrRkiwCue6wxhJ9+Vo28Ya8Ush9bLkW2nzC37fDAnALH9
3PayzasOpA/o9c8R6iVCOCeGeu+OijuSWMYFd0wtBOx7qUFMVcHeIVu+FOrUYjjbxVp5dg4AbIOS
GJ6ude9vH+0TfT+8ScbCHQGNjjCdFV5S4EjvF5+xRgN2VXpWWlnjR+xwrifsGth+2So7htLm1a71
/px+SAmdU2RSQ3Ug5vGPUIrjPS+H0AbI881ZWGOKVL43RqjpR+Dvzf33ErwmHNU8Vhgs53w26VD/
DdwyndzsQ5u08wnNX5hCn1KgsSxO4AiI3YEw5ZGyJgUkeRp8IuKXPZGf4cOKifBuThfIRoVcRxW1
JCE1YrMIFpga/S537O7nbKWTrFDPqXfWHeFBcr8Z6E7kJ+cvLE9FtY/5qUtvlzZcwuae/xv8xLOp
ErlsVx0bpYPEW7vR96Dj6WRC63A7B5+tQwvca0BGML5ZeS4kze3p0ox9J55X4x/yGVHsVmcEAUai
ukxm7NpFcbkJ/fHsC14lb5d1frSVozRVol77bQlIysdfjlzIoRFdvIH/6b7hlkOmnOUlcCD/wJep
RgFhLZuq86Z+ZoscFwfa4g6Z/3oHzfuSpC765i6HjH061FWQtypEWsdFxoB9sDBYOMqBFEUI/Nv4
mi6ZFwuG6Q/4I9e1lPdJV4OUxMVwE8m7ziyvz5fyv7x3pq+RyOrJpWJpIODfNnffVCuZVmmeF00M
3ajRlZtdZqPs2njL/XRy+usJj7MeYppxq+A36emX+HcA4aA9VZN2sSAsI42KNkuxGTYmBjiMxjPC
R2K9udOYJG8BTFKjyzqRq+3hD8SRVgrRKeeVEl9cPyNtuJd7yrxao7zPqn7ijrEfZqYceaDm7D9M
fiJ0nCZFl7DSYSUPUZowmxWxts7g0VOTzuM1DJdmmZaLTXaTQzk7a3bK5Tkb2B4O8H/lAuty7Ipa
0x2scqPr49X3uJCbkYmrJU19bUec0c0WtWtZm9tm+PwkvMwppmdJBeCbccPXqfdd2wlpYzqbPO8+
F6vmbKXVXbCq/9SIDf2q4JsSCcLCbsBIo0WHCYT4Wv9WFxBPFD10g45A1ESCXRp+0GMae9uEj8sU
ZRO3OSVwKGCoTLiTjbpJeWYFsf4WwL24ms4iwfPbPRsWr1jpVrj0Eg33SHqR9HJu60E99gFBD73A
8A3BJUNRub0InoUgrzyjhqAd3a0n4eF6dclNgmMhKcPSVPb9MlxjUSsSUeyFs3FD52/6U/zCcl3G
wDFJwXf6NZ1PyDjKwO/iUo/3xexINjrcSRrCERLUzd8TvuY45SUbp6C8C4iHFv3KwrJqP6hN9nL4
tT9MEtoMh8Rk9pfHoWa24IUZ9YWXP5ypcN87mQlvIzeLqWpnoU/xYGh7uz0DYzxkifSx9yjZhdSB
9e7zUMKf0PIj1A1HB8cjxQdBdmED/CjJRTcZA3y1hk44un5q2IOjUpz2BM2OqaNaEDKe2P6B9sD7
Yw1AZZDFp60ORTAVB4A98/PIQLKzrTt2kzOEwrG9g+Vcxi3UYSPqkRh9gv8ogXyvVHhLcPS+JMtz
CUQiUs1KFoAr2hRDWNAvRWfstAIzt/S6Q0JoZXtdEhBPnU+u6DmZ1gFdsd0wnMAygdIbYzGo8dNj
wFMAVxPfa+4gkLgmCf1/O4TZwbe/R3b/m2TprIne6KXnw9euWG2i69MLmun+qR7GzwXTGErwVd5X
YC7L0uDhfrBe6LKXS9I1KYiixoTvbhW4/psFVuKN4VsANE0ns2Noa3IR5GcC+kP5G9Ytl3KvIcko
dwyalc/pxhUxVIXdiTHsGRNO7JPVtVKTpkSkCtF7UC1RWJFZOEITUkVx6eMNovNPLFs1xVIfdofe
tz+8GbZVR+p1zeUJazz7ptAz+Rarty/+zgBwn3p+0u+y/Cfn/fe76y7MPipQrAz4LSbVodTwyOfH
iFlXiW9xsviPn6WgVKd5GcY2pOnZCJdqIvwRiwoXLIM3mFaM6EZtGwc8Z29GMgoD8lFzXSQ4COmt
PycpvsW++LUCxzpTkNjNh3X4tCx3fM3Eadqx65hyF7SoSNb7cvx6vla6QFIYKDNZbJOt9abwjdpp
O6HjG5u89cDVXva6KwmtUxOXvK5Dcs6mr8C4VqBejGc6CS/YzPaZ7gKHNRnyIvuDec1Ett5WmBsO
Ybi9ae2CITIfkq9ULoAErG8CXzGcbUMb3jG7mpP+/3m5diM8+duqbwIGMFPFe8znVIlsW1/YuMJL
azBxJtS5REveF4FlM2YKq40foZW2MCXl0l7HqRnxNcW3f5xfu6fRVUmSzioDVKhlG7DqiBy0kMRC
oeyic+12MoQE9wRDoVu8ri+y4HKWY8R38FO850deWEEv93HHGqbfxU6kJ9nx48fjj/AE9UC9CDFA
Jk+txAB54dsjKtaSj98acYsqUArFlUfmCkwJC2C4b5tpTvdGmufLYtZVN8Xusdy52CZo4MZ83cvW
VcNX5yNvEZLR0CT0qddqfl6pI8ot0DxqHnDmI1wvazKoj+Za0Kp6Cyfga0aJfAIbd0GqJuEy3F7W
ufpIBI1kzgFp78tdFzksKtDcjsUc1JWIZ4ih377beOwoOxvdpqY8t++Eyb9CWShIKB+59MEy8Rz4
SEmrEKQ7S4EOR6+sKSifai9hDdyrpiTcvdcHHhQmpYDjy+pUHYrs8uQWbGZKN1GW5usKO1RVECA7
Qw6Vz2S6ceegnYxpvz93PC2VTfyLfT8kuvMwaWCiNz0IX0JrihF4qcDHViimDjN9m6U5ZBHBt8Xv
hHfLZJbDJ/GlKrFUYuaLOeplyamWCnJbqpBCvbz+88gNEDH1/6M1r5I7iLDo397wlwNvTqSBfhfG
lBHf4cv1gW1JL3gKd9itzdm5M1N6jW1ynJxS3tJqx6cMVkrUREdXZ3eJw8w/k+khu5aqGNOtgxQH
bDGfqexaze3/F5pjpRs16lZJJeyxnul5Ae1edH+gbzbjfHz7oPgumWsTwDcYc9kLzmXn9JPtbEbm
qAW1erZJVZrzmS/3CW9JFHjDUamFMxuJmZPDkoXpn6fUABsKVL1cSAOrptZqRZY2+ZMoOvbKx6Lo
wDffE1y1bDlVN/vfAmIHIqdwhQMZSvba2x/pC0YSikA4zwAiuwalIjelEAdghm/kHXWpLgAZkFjg
UOx5w+x1f7in1NmNWm2JcnRhnzaz2Ixy8pbpszm2vDKy5G8tYO9rDqocdK8T0bOfAoONdZSnLPHy
IMRTeSAht2eaSqAxrqSj0YnTwZATyFknsKIbLDs1FIs3tfHE+B16KvW7pqJc4jjdtZlx0CESIlGs
2mfd7g0SnFbWw3/+nGfBDMmDrhYAMdEy9stuVbgchmLQEFCT8BvQ1Ew43NIpFS0gDLYtiRuM+NWV
1od1A71U593lR9VNzAdgx7gQuO/zyRrGiM21KpfqwEH1OdqkiLhxmrv2p4qnIcrGhgNte/TPgvf9
gHSuXlEJO3yhjt+yWwdsD79YN5VamsSk7DmquEEeUXf8JP/so3PMmFwCJlaBwww9jx1MbWvC6LdG
2bX62Dioti+jvyJz2laI3c4jy1me2rbSBka4qkTAEk56eRBB87QBtDDg6ed1i1aMQL3Ksj5O1pJL
dnIcQV8jMzWtm1bDj+k13yKxim+BX2yfiFm2AFFGWAJp1LxCShy1HJN2jOyhrElXFw1Vl3wrvKcv
6x8oJiawD1xYVnYm9pnk3SykIeUThOHUYZzzhSL8mcTlCTGrbBqiEIE8eyWuRUMAYzbyWvBxzP+3
zGeF9yXuGKkSGDfFWX7+qim03iZK5F8sFKvA/oXfYmwjj1CQaYTnkjvfTJePZNxGRApDgKaM921T
5qzeNHeGHbMLbiVqPGDWApv3R8GmR0uLyX1hCYgNwrgs0bZCVASSXIIz/acjgT5vzVVyiYLkB/eL
cFoK7D8HuIBDn5UDvbOZDLQ8iupWMPzimN0HRGnjN804E5txf42V4sk/Es3jfnN/wegXKfr9TsPA
0xVBf0/deyYsukhmBQoPAlZ+wP4n96f4Cj58l08DAND3ODXsAjPEGZuLJ/z9WOnt9h00SS+pwpCr
rixg1fU8d6Ah4N90FhIXRLaNqL5mUUJ6cj85mPUZonCIFg+moHpwqA/HIA7YQ2xdo2wc+U0LxbJY
uPMsFm8oX+3LNnMyTdg14ZC1wvJRoHc++e/fljt1WlOiKgbOhB57jRWPbCAzuOS7cRJMa0FuLV6r
NcrZfZmi412JnEFAlXs4Qc0v8VhsVuHHYQuckn/dZbBKdk/ARzHFRBLjKcRef/aCffhR4ZhV3UL3
1bXgN5kbYnfFVhr3Si2ZVW0XwXB6hWWC2K2PAIv0cmub1A9YZzEeFkzr2XwHC7f0vw3ukkzSvNtN
ejdoOnx7mpJYrlaneDyDp7JSkTSigxHVfGtPnUMZ/05xwOCFRBjB9EqbTbXTzyO19DGQAqGOaqXq
o+CBxfyrFROGgq++lMGtyDK3CPvBynpFUtA4CdSgJiNslIumY7kPXDTj1rfrroH/paeHJZVxE5Ix
5ciwEkaYdGSq2XrbLJuQtwuIIMOaXdBEr8YgKL93LMyH7Kmu7lZSZGxDkcCmsr4Nukxy0bsAuORM
Ylco2ypfbUaMGDvn63u2ijRjQxDoqhZJsrU3qdioBM+T3DEjUSuhQ+mDK7mp01K4xIAQ4Pna7Zma
mIT5T7/56kIWIlq3dZWiiU2pup9IVscJLZS7U4pI1xs94Y2/kvoSiIIqfaBCmh5hyIeJMC8xv9kB
mX7iYZA1XgKAmLmw2kLMmH6c7vm7Tk6Hr6q8mDw1TPk5HYPA4TwW/CviSh9X/jOdWfWXWD7B0x9O
vhMTD+eSd96SlpEQP3lLu0PB4NdII9tacBXxQSxMuGtDYMAMliPJ8ms1HQV42Oz5FNYNIAia7vqC
qR6Lug3KfU9Eyt69q4HXfJ+PpjqL+IJbDBLvMZjPYwILUUtU6zKLBWSBEz1EceGcj7Vb/ZBgjDJr
X5m9rRkrY0B1bPgNgcGpuPgkZ2TmoQ0gCjzLADm6V8Ca1bBTWFwuyn5aEB19xTqw8ZhWflCndoPA
0XO2ExXdP6yp/dDFJBPrZyuifN6uyxsJXp7cpl8ILK7mLiLE2bZuqSfWShkeChqHlx6yln8qbfVt
H3IWRiWdNz6bG3hyChiKBfqcS/u4PCjJl67XipRvdmHNH3Q4/nOYxL0Ex8J57Ps27X9khQrB5oAm
FkyFwSLjVS0fLktDhV3npk9w66/bU1NP/RDLlDk8dQb43baOLX8OC85Z3nzq5brSq4PFVWDwYOd1
rcqr/oXFEBZtolc2axx+zq9+kN6Ac8epzYZaO/zlHuTzIAEx2QyFBTGJuGTc/3pmO3z5ZGJ7BMjk
SJE16J+ToxylRE0vhdkTgPYiKy64AXxa9YxtEL3ZKI0C/6lkefPhQpaeM9K4zsp3Hsgbk/aLB+gR
56eDisIVrc54d+YB9ipYjbyxflohnfKEAfBDSdXllwXHHGs5oSn1Et3+DJfkN1QU8cbBjGeWlhNN
4katdc3mPlnscpvK1PYODHCnf5N882TCjpERk3HnO2estFOhd5Z11hJKuzM/Xl4JSsmHPCbqkT40
fbyd1QZEpECb1m0bxFtSPBUn6C9YUUopmuLZF8EqnDFT0S2/9JFx4DQs2H+sLS83qyYPZrmS3rMv
Y1yMdZa5q1hKEA4S19zLrKceSQE26JazE0RCqLK6UOQDjQCmtToQDzQyn83Re6JUahieLowiYg3Z
eIqdTU3sCNsQtCXQB5WcUOzik/1wMmhInCox0ovj3RhmRLxv4C3ylhoJGdpj05z5DbP1egms4bNJ
ePQWSoSc+qYnyzHPckRmrPyhXxVB9h6fDS0r3xs5rOhtm95PqkMXEDtWi0y4NK7tTi8CBJX/3WJX
wwCgCEoo3hkhjlzxGNpZxGQf3/1nwrFvGHj1iPx2A8dO9TlGwkybDy9cg7MzE3s6ObqTOLDn2CgP
zBP+rLvffPbxXbdaueOa07JCCh5CPOiQHuB4FNE6pBP+0NOspErTMifLVrx1z4LStDl07UqYFbnV
tcUU2dT+RwbdjTQxAe4WQy17nLYeTWHlhZwWfULC7n2LbwKjW182wTuC7lG5a2H0j4k85g3Tv945
bAnVShMSgmi5BTCLCzGB1S7xRsk6v2QQvRGdVdnQd3qY0Dciy+uZ0W/AddE4ZDLbM54rAJ71Ls5y
oj0Lpg1sWuH4zBxOOMz9MfrM8ujHXIQQKyw2QXmAzYwlXguBLvF5TwBLRgY5opvujTAb6mtCCeTM
0QnQwEZa6NhunGT+Awi5ckw7WbH4McxiiomiBZPmNin2Sy3rpD3uXhBGpmo/Nvp4ugxe/qFusMsb
F2LHZrtQ88ZKTsOeY+Fq2cytVdyeYv+MhHjHA/Jso71CBl0Yi6HOjVMuonGlmelbzVblrQ2pg6yP
S1YrkFlVgp3aGQ+XC2SftLo3CctRqhL9rNxZYpn1Weo48e+TBmSR1egHSVk5BrbXUPyPiEBqGBc5
Pev3eEisq/lBwNTzzs1kI2igqmAeD5dDsH4PRxFTtsrrcVrK8XleMFVCsg9EdDW3koAiiu85hg3S
3NdIYO/2MQdWDf8VltKYfzcAITxX0TEFzbpnm9wgbEpiJLHOtuneGMEdTUewprs/myLR4hmfXFYm
XFnrUUyeQ4+kv4U51+Z3GhjE6XrMvyFkefg49yFZptRThss0D4gzV3YI1G8mWH/k5WqgVlgLdJgj
YIXWgK8iayRI2okHW9eVQ8WDu8JjCbgFsfMHDrp28+eeN5G+995+vn2+/fU3s66leCzEKzHbAmSd
94Qc3VSEeBZwRfg9YOY8qk5h2TzS42yeqLS0LgCB0GOVMaEn3bi3tk4Ryi9KbU0+LBeKTfpgHICW
sVw9qIeJKjaBi/xrSMh/m6B1fMg0FcWQqiUo5J6iXqtwXFzbsW9qU/aGDmg9Rrh+IoEExiilgPKT
zI4+4T2vc9bSexdNGC5UTE0JwCrtJbxZKJLKmx3mXhqZSIXQ7fTidRJPjlsWd5F974PjIxciq6wF
tI4t3qmSKOeKp90RKyAwLSpyoTVXElHI4rZXAEennZxMagmDXd9z97iiRI72i9G2v/ooz5wuAS4g
jVONi4Muw1RE7jax5UgAUeLpK0UkCaIUOTR59VmZgFE74seOOuOu55s9ZBVeUBQ5ahx93Omjo2Mw
sOFNvK6DrRpNLXLum53DChUINlr3UEB/Lqc+GfRpsecOfIg6Zit5UzvW17OrGoO0P69GAke3tvtI
ZhTkRGqKFIsBBAFWAnUWjWKDw6zsf1LbIikig75RSuLRs7HFkmlIfOROHpkG6g5gO/tvYOdP1soK
ghkbAwwKpOqcyBW6db/u1uEjhLNnRWbhtzGACOX81OAIEKkUzpBone4KNYogTvnfPYt+Szw597XQ
cVDk+Hk8yAniWGNciNPE0yloISweYqLs7DlSaL/uaOvlGwcMNS48UZLky1BT+nz4Ki1oeszg00YG
1zEtnai1b2F8FtZZnAOiK/hK1oPLVgZqCcF6XWb6l3cqIn/8ANVD+CPNM5F7yxcSKQntdG/190DF
5OY8wCcQKSI1h9xDmSlws6Zyjq8GmDFqGyVoEbXrafLT6fBpIGkQy4/ZxoPCw03WFnzwO8g4Ersf
V+wSbYFFWh78yucW7CNin7pp4TA2HrFuVJ/PICMVbuFSkoBMox66neLguXOrvRoRa+wPcPVi8U8p
0/e+1YR3+Jv9B1OiRpHNiD0l0qw+URQIjTXG6qiKhi6pBd4rPfKRTXw7WiSJngH1g0gLhaViNfID
mnr+SedPiMDGHQONQ8hg29UM9Ma1dicfHHrgmqfs4AEgF7EKWE7pvdMSKRpy8+sLiObLmLtOc4RO
5k1LVgQz91IC4FWRsjYLnPZa6tCvL9/ZQKPODeZU2hd4lg1bsdGTSKwgiW5E6beIdf3+ssljbbNk
SDhWP+/I10OvtltSf1mIh2U7UKAhVrzNZWy/hm6KigbZgcZaG3u2dch14xvdFXmyzMG/6TN4LQHi
aFAfSj7suwmfyt0sMxG3wcd4HpDPDfvyChNrSsIV7TSoslETS1y3MngHZPj0dRtZg18mF2wnK4qv
MGYFYgz6gm+BfK5FQ/TIe9QMib2B2DUljJ7KkAlt56292KdTleEI6Uybd7e+OrcWgPn8cUEztFY4
YKTHS2uw2qZTrfiFZNlk1C4hocO7mbYJf9zi0ZT5A+xarDzOjygFPyw1GKTPRFrpWwVU09iU08bj
YkQkE6xzPOmjhnOA+bKlfTWA9oNQeO/xYWR7Wi8J+uzjOc7oA91knp6/MaYTo1MFMLwllBsjspG7
LI1MBHsVrs4gmPR8uJF7eg7EZZKC8pNslzpPVuQbbMo+vCvebxbu939QHjZxPev3pG6Lame0VsiC
YuUbvzAaCjSVDz/jpNRZKG05IAEjBEPTjIKQvdXKJ91JreQjSdPx0QnrRlky3ROmq8xz9Pyrtl3n
vACdA//sxnbmUINKJP1WdfxOvFIyl2ObibowvAQ/Rj1X2fixDrRKSTmpcDtR5bNaHvO3PJDufK3W
zAIaBucG/gbw4EiK1SkAtftZLOSq14n6FfPySbG2qmIntF29heMoRFLejEfG+6mqeOOfrsPt7whv
ujTLPXIvnuJ5Y8BDCPuAwFpBPLkF05/Ypu448tARh/NrEoaCxFrNxOGDUA15rG2rzhgIeOvPMW9M
B0iXL8Slzl9Uc8yiFcXkQV7RMi1WlUVfsEf/QsgDlyqhWAEFKvFvYojBCM26ZeCWnrBjiKDcvEBC
jHNyvU2gbNpxN08WO1saumxylDy3ql1u1sKi/39OLR/AN1NI5X8xr5FRPljKudBTD95ZB7Ga1I6b
0n95n5DFRdBX1/AA1e8t/+DhYrnJ1tf0sayTU+wcTiC/pyyeAz5KZ/ul0tJnr+ztd6sfJU9l1QJu
dBGPATk870JdxZYfsnVNSNPYD4zzuJxI2Qk/Bl884Eo2qrkMWJLNM1dirX9JCiJm/SDFk/4T26Uc
W9sN0m/6vgIZIcdFSCSxrJ2QUemeUZ76eSxdn2Nw8CDrfHXEpXeP0B8ynt/zGDqx98iemnoi0ev3
WnUPxe2DNU1yRIIpjXcO3rEsVXY+dciG6OLlXhktToSgGyj7lnDitCNzGOxz4Ik3nOaiE3pzNRbE
vrkOO36sKK5k+8WeG9C2Rnfb5Rwr1idLPkpJPl8tVmu7HFPc2LzI1Yitok2hrEwB7qw2mwlNqO89
DUMa2Xe4ROMP/XIixqPJuDbRYaiX+moMizOpD7aRqb+wqqKRVyrhirryZdSfjq+JRiQ7+E3pZxLy
bDI3Qbukov1w5xeDormiWwCwVmmgQPLIeaigCq3k5PAS0z9SeIkdWPldtevsZITenPeMHAvJLTyD
wT59r8SKsnlCHAgA+ZpyWL/witSEDbS2qGWPaab2N860V+AJUmBwsgafDjSZg/G0u7w/UNfyGx2T
SvDASvicGbEUFJWqE8rYCVKfjOOsb77F6GbiH4sNXMs2M8ox4ebFNkfabz5BEsH6oairpBbmydth
tr8LycivAhERfp31hYj22KSr8ny5HTqrxgiQnByKt+bdlZ10QLf2bS1ScvqAwcJa11gNo4DNZs4p
GWxYfKTNf/OdOzgVxtzyyEMNg0DTf5Z5XUfcyKs10JVwSgXdUmCKpnPrPFtso423b58MvuyRg9t1
iO6BiZKvp6pTCw7nMQaG0NHuBtiw8dYo7xS1edvN82peFT2m77Smd8fT1mKiuXDII0S+Tq/WVb+0
kLZzUszPe9frnyH74sO3V9hH5+nH3GGhjDGX+Dye48W3slGOuXvxmLaRPCNEqoL+YNlggduxS75v
8e8sU68swavO8Z0Cq85+HElikgxJQfGg2sxvHizxm//ywoN/sFQIL1LtcCGbG5X8iMXrceo3WpMk
EYXuacJEkFLwXgZKzAdCp3rl+TWyq68fvMpsCfqNODRsFayQPhMWN6nG88F1tfrlTMP9KoHwb29/
1uuWjfh0hXAplVbptKVdesYB/g3xK2sF+7xNQjHlTkFHxhcWXpHU1t4GoRP8Fc6LHI2LdRMFYYLT
oCFJpIIuj9aIStOopilMaqc/CNoOz3JxP4auafIgPfate2mqgHM+ldgIUioM5jo1dm7aGBrDOP3R
kx5qk/tLkyQgoXbDmdozlhmE5NKZs/58YHgaWiNo9/x7CPvYGzJsD35s0lD+diNXt2NRMmTPrhrv
WlTl+X/JIepgjYSALALoZzg6pVD56nGFa+RHU/wFru1tuworTqUU7bNgOGLqOqr/P6enfj7w7Y/t
GQplt24Ex+U1mZCcha7mI8N8ndf14ulf9dRRozPZMl01iGLvq6NbBj+5KBIfGDaDBAfQ9tiJmMKd
0Hc57d540IzbCbwhOuEkV5eAwH0tDmX4SzYfUe0tRc1BB8uR6giBMElOXP6jCfC/RD/eMeMnT56U
fZzgLi3cECuMlyU5AtPRIZoapG1RFdeLUg+YQ1fitxieai+xFehhADR4Ro/YEKULNdYfVqfVjikQ
7k5dHlGaQAZvTDFmSlYXbcKP8jVw7Hq7tzZtXfopJxy1W7s4yUFT0eASm4Xxwgci2IvwqURA8La4
IvEVSIY/+MjcME98Lqla9cYMsunw2cOlKTOl14wiaiLw5TQTngP+QKdrqPdT3hwHyrMp1reB6+Vj
0tBg6h3oTFFt0AMN2g11Oq9/Q5VuNfRL25PEVZvSe3CDz0twtogv2HcB0YMjqMQclMsjn0nr/GBl
6kb+MV59hOKB8pUx6eP0BtGtBm2jLtRF5Au06xG3biax7tktV8HhWwwCZ/xssMgsTE5VcsodcN4H
7P2NGLRS0mAVGuDDWNrIALkWlATaBLk7AowlliKUywbGh55AOiE2ZCrpAwgIS6861yzElP2dySiB
iSxJgvZNL7x8ZtrIUvGjPfjKSioPVqTSJiYJ5UH4jWgp6w/Pku0L8yeIOQydecGwzEEfWNcyQcAd
X+6Ed54cSSFfJ+KFtH7filHDwUWKmTh7EgEE/PgOBNN8mtw7oHLNxV+qqkm88/5DQNqpuTC8t3/k
gT3Be22CXZfKIDJ49x0I3VAeav8BCbfAoCyRxxH35g630bwtjWshWQQXlL90wSrG3A4cbSXnABC1
2ZWu7bFA4R5nDlxQjlrtaT3/+eu3jhwaLgKZqyB9ROVBJNQrTphWuD22LenVkxRVSOWT+2HlAJX1
X38V8LJ/YtcWyz2P4kFzvF0LGwil6agYhtoycOjqOobCVnBTU00sbRHudX/G+GChOpmaDbLeF+iN
Nijg1Jfpl3tk/Gz00fA49P1EZLQWgeoFFRIeLe7eboOndBRNXJ1macmiw9/PBl5uUF42S8F+t9s9
d5aOA/l1rBfL5JC0WGjMbRwBIzFv+nDHUeyI1A2m33MGBy+s//NMY+8elbOG45Jbgof+1Xk/SWoQ
X09xecUJ+APkV7/9yggxGk4MJegYBhF7FEbSzwhHjcKSyxUvUGD3ECxB/ommqsqxHBPchEFLCVYV
k9T9M0O8hEjlmCigShboSXRO++SRewRexMavJrepZmTSfoNNq8SXLZ5JQJU2weXcmfVoBmu354qm
O1WSnLLm2vqlje6QhXPBF9GZodeSVB3946c4aSVjW3OkhrHymWlb7LLzdGoVxsmCfMFU/x6hCul8
nz0mIv3pARdGhz5YJzgzaQFPRYxStjbd1eVNU8BgAnEn8ej8Be8/cdiavc4sBAsQqs2BuNnk6Byz
oin+SKrz7/bHJ2kaU3lHoWDvpG5IVVxOumlAik0bGeCAt8ZwiPnHNoqWCHEiSJhbLpJtMMWaBLAf
aUEtipHX5fcqo1FrukxfyRf/NDxvvL94F5zD6+zNhDyQAVjj74uQmkCZOT6UdUuUdJURcPKcbUxF
YbxBD8p1nMPwtTNNsxrCUcriKHQ/ux/GtURN2aMqWXCk/u8IxH6mZruyfQyvmmD4N05NcCoposC2
XHJo8hf5fAbJYVNcasft4xMFX6JRy137nuIi+cwROpEBPD0oequu/M4jDytAxPDaS/v6RP/j5p4Z
qGc4R8zko2THNOkJCHSsGBzRVDCOO26GRNl2fyTOIfKWQ3puvsyefKbIiX1/Uu6FbWUkDbHjEeTN
w0ttN1O89crBXWOOG0af0RuDW3yYwEc+DusZra7S/GwL5YZ2es+wmKcQgCnDl/3kMEQaWQD65ntO
NUl97+1YXmOg7N0vo8Vt1MwkgSFANZmKmeOxl/t34aWuhpFpLENsu9MKzQeeO0/sYxH1q1Ic13qK
axJvAUkIEr/HUyHP8/22ploy/I4lIpN+GDjnKYER543Q+BnMs6r6JJ16AtxTsyU8oTjcQcIMidnz
aTEgw3wbOYzjD3LGc19yNAngUmMugsMiGT+mdx5q9xQxIqxaOYcAckT+yAImMoiYH8LGK4O6jU4T
RWS4yP9WP7tnvUOX/+5ZGCQj/lgKHjt04sWwRL3xuGWap4m+6C8cmi4c7y0GYWw7FLEkPc5PSOcl
YyPB3aVnKahIQ+XMqZ3cDi0/HVCVaD5WHl9jk6uLuTShmaAyh3osE0C9QrWSijoAsOe62apDlkjv
RRjgvmiaSnanUzN1bO5Ys2UKMa4CuDX584HbJeS2sVAgD0TEj9gmtOmE/1bdUSGu0K4MkVZm64/s
v5FKhOiK1CCFdjZKLEEjiExs76SXOGs1YOsvsVEazrqfnQKH/LwHrF5lcpNhYnpgivZcPHocH/Dp
AneamSNt2EyPKBTVNjZbbHTxLjUPZB7RmQxQaZjbdWd+tOcw9mfZMvbIl5RdW7p6AWn4FZajq64e
wtUws7XEQ/lpA01jfqF73UdLyFZSRxjnSpq5SXirE0H40rvi9yUbPDoI8OdeBe/cwbOLZDn25ZBL
28EPYO4heU/AS47wDjz+69HIWXdDhW9L40aKN4Wo+StUTQCEKRymAV58ZelcQ7X0w1FPcLP9ZOzz
HYmmczyWMm742TtVYOj2SEFo695syRXfcKCqlnosLuXUt74IOUIP9PfkaxHWePTEyXBoGWxzYquj
fc1kt5A6cYUceCmYCC4nsaaYVfGQ8JuiPO/1bTDi4dXuO+s0eFBuBn0l/WpJRD/hChS9qgVcaEX5
MvNBAhcXvKoiJic00DBZlb5HsGJSoIeO48PSKqepAtghkCz9KiKbiYfWfjPOzDIGwdS8liE2fjZS
ZFlORXruKHReQ/I+dIqW+QYIXdnAGIXGSu2xUBIgq0MQO2eRpmt8Ea6En+4YBuszSGDP0wTpOV/j
2DUSIErjrTi5j3lZ80xyyoJDR+BdIDApxlIBDjISx/hriJPMYE2/93mEbA0bx180HwBvlBjs+wPE
4rh9NsXmyCWZzPiDH9188HASM6WXtXwjr2TV89JiSjaIJ4+K504UI3r9LrTYmWZShfa4ET2dop8F
nFr+uPN7sjTOJ/YSfhHKdCTmlqUOH33K8oA6vE8TCFvMCLlMTUg7H011xCi4oib0bOCIWW4oZfbO
EWhZ0bc1LYag3gsCIbPpK/AajPajfs35d5X7F9eQ3DvVlJ93voehlfOBKPaotpz/UKHOoABBr4/c
Tq9V1b8iAIcgRHWws3YNKpuiHZIT+GznQHyYVA545x5UbsJ2UVL/tuA0ZA3oszpWJaaCkUZVQxnO
oWF6MPdsTmJnzc02OtaHomE3VEmCdgISvzCUAJKK61ye6qbPAXxvYru92G7pce0mX1GLTc1XySZO
JiAebOZ3JKkHYKdh+lNeNmYWIOm2Etqxq961M8O+R17p3Mvm9jSh5EfzGkgIvewQhPwvx3sykYNT
PjIn7hNTVlDPkeJY13/LP2eZptLd4DtJrRhpOOS2dZ+7bSm+JQRRSYWV/oOCckA0CJKDJBc5V6IR
XpMakjJaP2EqcFsksEZIWJfi3zUHarqEmN2n5uWS6pYoIGQ9UoRlssfwM1U/9E8pjThrqS664gUA
Be/dzmQpD3PPh6BkHdmXkmWcOR5D2/ARh7dri0UXYfBrZ7l9MEi9bT9ngx7pp5U9QQkc08dZbQWR
t/VCuO8MX1SnTOft86a0O5FbE75YIzaw0CQL1VqP8/fMq8WYUclmvxMY/98UHGn7PtTZzwfgXVQn
yvifgByoWhGIy0/GnNzPqTuEKNierK7zkR+Tqo5Kmwtc+HitZBP3NOEHHBJRqalN3Du9fagrY+g+
xdEUmci2OqYsPUUMlfmeUs71v7jS5VGwI6fQTT83JEYA5kep33jg1rNvp7E9tOTF0dLq1a5ULxp2
l8BwA9tWva5N0yxiBTspqkM/o3tTEPKSp7FsLnuKk6beUYA2P9WGflRFHaSHbkvL0b0cdj6x87wO
wnIPFSSBTtDo/EKTAllUWN4+fbvl2LuuMaUD2KrrL0sCgcsoKA9ZlpZ6p87UV6M1AP8K1v3O9qBo
E4Xtkco7kErih82pmiohQdS8ogSE3uNELedank8LRZUNaCyUq4uuu6Psfm6GjCx8StGpE7kT0mA0
HetXPoO1fzyCvqcq9XolSfpaNwBrg1ygpfuIQwXRKLFwgcGqE8SJ5feyfv4N26VHPiXNXnmIkv9U
6radPFtVatLkhm6t1dPRtR+QFAdmHBWXjJ58GWSh/WEoyV3rtaLMyrgYziN2zq6FKbjaywduoRTb
m1Qt9uYW1w3UQPHy8WE7xS8xIgxqqcb0GAm0qX0g9kIDrHRkDAkTm9cmrZaZ/MhErZiPBCkhyBHL
M8TrCfGmZ7VkGAEb9IjNtH4Kiv12zEwh8afUD/Lzd/xyPqEW6bgrKnMxlYMdBdxPbknMCOCz+N5E
SmlkIsNKscB4GaAfWth5VV0324xTSQQ5QhFr2zRZruH7DElyQVccgvDlN0imNlGjPAPZvuNeh38e
YHfyODWbaUv/vHeBUgNmLyGDf7kBJSeSFuLMmrVrdiiNVIHAGhjWwpgl3aYAV7ZiL52V5+Vs2Gwy
KOn8QGMEHTgObLaCpj16WKvvEjkCBdK9yyd1HSq/b5f54kBlGwiG1pYV+7xLmU8nOP5MbCxoCKK2
IGkELrhwJ2t261LaqNin+VvSHB4p3p11rgYCLDfufxLmFRWpiAvUbMbNwfZ45c5gvZKKnbkxDl5z
aGKY3nj39OZ4VuB+xJC+ta5vKOza6+gJZjXpLaizJ6Lu7Kzo3fvTsfSRvIemnZCW3faG+BLpd70z
4MZ80uRmB20P2tFbr7oJ5ewi1vkSp8dixqPc0qHQIShElP7lrI/SvND74X7qe7vjhwGp9rwPNWEu
xqAVWd3t5YasoS+GC7r3TC+2K2OQ8rUiI6ReaE2iwBWyf3cH41NJoR2JdQ4wp3eD8i/sKj0FzXdG
MIlvxiO3DxyX4ebAKajxlCXIjCtC0MQ18yQjZWiEhexKI+0TAEa5IY8jjBydHDNYb4yqmIhJeTJf
ANloF3VCB8WhXpnNa8fZs9xWLMmWhiXPvhYds5J663hVLdh4lEHnpGXcyoX3hkKijU9pmS8m0KMc
7Ykst9AnVOc0bkrya5JTZZhOtzWGoWdyhjPdQFB8YgOJfECByGgsXcp+aabRb7wYBFZA4n2+eSbt
vkCslq6GAOKaLDHfPm5y3DE5iVjkszOvpV5tcsIsG2tQqmfuNOtwM6rXHZbAnufLpN/cSGCZY7pw
y5E5Ep5+9lU6MXIASbPZ2ci8VNLBupYIJTeKENHgwkMPcZY3u3Ay/0rrtQFxO2sjc9iToic6YtV8
BNZRTobfOF23zoRB4FMbJ1RUiLLfelxodsBdmJmBCiILfpCPNqfjD91kFawUsB44cYvCPbZ1EHHG
Sb1mcxzpzrm/WvU26kVGiM2SwY4Z7gNKrPpGzF+GFOZ3/sAP0RGTgzfbbZKfsC2VHo8jHVSy3jSB
NWk4pmoRxgn/mLkZc2fHohs228po5ZKlXsNBR7UoX/jf52bY33NsWRBrdONcVjvkIrWeD5gZve1m
whknxeaPvvrafulkeFnbUZKS5YS82jBJN+wyfyPjHSe49cZQyzIcNuDyWt6h8hdrFdhogskICf+L
V/o4zVNCDqKc+sHhJyapHk0nnWB4LRzB0A3WRyuJRdiDNn+CzlMB98d/+u9HrmEpcYUshRTeZ0AH
jUefGEP7IxSIEHYibvNqvhITAh53nqaPd62iX4UAIfbgdCiK30OYVx3532IfH4PPNVzdPK0+5JJO
MX2UG0ksJ2aR1jHwHEkT6nfv9dAQddI3ZL57b91TlTLQmfbeFg/bjjX1nmRj0VsD9Xdvp5VqwRKN
qxHdzBmgtsl1z+EeFXqt0ZiZslnb1XoA389pLzaImuKj9EYQUCvVCpcGKQ6AdkJg61eOjvHNjL44
Cam/xL/iWJ94rd8ItgloJk0cTOphnkXqRUkWttlHptpnJ6ueWMIJVjv9zH5h7i13iLv8pjlDJW5l
4/4qJxLHWgNWLPALxxAkxmKF+OTbV1Q6ut0CRteHVs5jlceIzomaQ3ORoPpimcPRIcJR8y9kkRo4
o0TY0av2GNaE8ioo6LIdyo8t2mJfVlmMP/R8ThkP6NXsx1U7v+V80aDJNj9lMgz0YqmM8YxUFYn3
+fTDhmySyLFPEAKXwyK1DBtaKXbXIPYptTcHZhxLS6sk1GmMoRdprmuiy35TrYbr7Mvg6elmn4zr
Hh437uUMqiyeMSkC3DY3N5o+4iRz1wm0Nu3PV+TYP7HLT35GG3ebeDptqt6QMFd33bB+Gjd9evDQ
r2Z3Rcr/FwW0++YYXk6f4cd7My/jBi519QO09y5+Lw+q9xpReena+bKic2z3y19uZNV9XrowrNZL
iqOfdOFzzo/4PjjlWKV4+NA47Je9MIxU0DlpwXJEJNjYasdQLKy6Kpv6rBrk4wt7GY1flwa8oKk6
zsqUATKe0X/1DR/PyLGF0fEWTXHKo7WWxPdBFSNDxMC0q8DRx5ZS5hhIecDvDDdqojx8TVsFl4IW
zmdF7sJMfKZq2OenoiwSW5fYfC5cGl2xXQSKUwcpZa0sazjHFVKK4J5bQs7ENCDyIkZI+U5F0/yo
MInGyXwy8DAjBip7Kub3CCT2/AYpoaFf2jQYj17dnafZGsC0ZPJhNiTj1iYtSVnCA81tHGyYMzZ5
2GpzbJJfShDxoI+dF9xqPLwSGr0TGFHA8Tfjjv8jIjRca63ZQI8sXv5x54SlfT21Zy7zUiXZA+Ns
UTKNJpuTzKF4Ajpbov6Bf9m02BVacIHJ5+yXkGrfdcEf6biTVUoeKCNFegELrLLXtGypGWeXGQMx
xtvs4/KXEUabpgrIjLjlD5G+RanLWmWw1ukF/fVRa+YawZ7xDMmNo35wtE+YhmeaiRuwlf1a0ZrU
GFrqSD8RodwS96iQiJxqJM6dX+vORb/Ru2Hup7/BfSYhATsvyhz+wgx62Hn1gIWgOcGcqFoaCwDX
VDaFOwFLXwc4wpJ+GJxvcztx29B6J1DhhmvbDo2HzE/6vf91atclwWSBkfC5ggq2XvcLwcV27N11
pubwMSsXwLItWyVl4KQfzAJnmNJHIWmUHUbjj4emjBLpjWgf+3z8vY150VFdVaBW7Hh3ccTWmfx7
t1jOSZaTczFP87iAK7xPAt9uZvsdytAildSX0USyE1xYRW6SlHG4U5dO6wtb00A7zdFBIEa9dllI
Gff8azof5gpLMAvSffEqu7oWhOt9SRUUIxfyvfqRtRDkgTuJ3NCrKuF8BuB1+ERXZuWNxCwfgraz
UZAl+Oq9JUbAdLZ2Hpksvum0+wqpZU+5T0AwUuK/ZtJ9WMrCR97lOn6AFNQcugVN6zXT0XeX8dh7
JRLXvdRIiNo9P/o4HayVVQZO8CLFycXBFSfJSJ9KmUNVwI22ktgK5VkRyysbYA+Q3SqtXQv2+Mq+
iycTAv5SdOVaHM9s0qbxCR9fV3TC2dJkEsnA6iqpqLuklRJbE1lDhkUGCUVodm/g5WLRpvoymJha
8ehfSqT0EKx886wQre57RR4aiisy6x1PhjV/rlRKrciXOL3hGq0WnsoaRiO8p04RaTZxp/ATcZuO
Y8V+DlqzawQUaek1w8avfdAdJdnky+flwnNDoFo4gnY7IjIEJidvCwW2jAIL5R7vKwME3JlaXStt
J9Azcet11JbzhYvA3hxOteB1NVBahJB7/AiJwY78W2sfBhjFogtqhWd9uymd/OnyUKuG/1YTCXMS
ci8fUg4GlAkJkwADqhlxJPxVYczPm0+ZD5ChIcj/9ypegpJ3fe7QghfQuWeqFTpyf2D8K6334qWm
01ywrDH3fnAdUZVkSo+ZMRtDeQgUkcDgy2shPtJnjTn/9+aaeEEz7hI+ZyaMgL4eJmm7X1FcI+Wx
eEy4Mh9bZ7Ev0+F6jj6KeKA5CjdlN/HysiIPUI+MKe1Uk+vb947vGGAZNsovpYYO1ZenBR14HysL
rXg9kOeMaaCyssbR9Tq5xCSbXYh6e9I4FqSvLhnVnnBIcBuQFSF8IhGeX9uaGn0Y6a62EB/b5Fw4
dFJ7em2iFj4l0IKcJDIcOnKVGVZkaNxc7bsTws77eCPvKBXMS7gCTIP7pCTVtciI9l067QSY/6Hf
Lzdw95cgQS1kHxDKbLO3ar0Yizxq1dUIQMn4J17VAHxVKrM4GqjIYNymMcKESM7RqgekWgtjxShV
g7gIXIrOix+WH52RK8QsTZPkNmG5m3ymxni4dGiyw4/F79aBIdUMvDhmBhEThEjrrlty6ci9xnW3
5sU3t3zjaMNVa0UuWDrzcYSstqO+HA6Msj+EjgPyPqaghnsUDH/Esb5WCeso+SUo2DMpE0pW4ywS
b1mO3ylo9M5m29j0ZMj6jPg5KTgFpgVCxqQq7SuSssMXD11QCMMjlPFn7D/yVfP0Rmr2nAX1bS9K
h6kQDc4lBD6mW6W47vumZwle7nJxagCfBlhweBDQmTvDOU+rDlShYUkCeL1ETQJ6oupauvkFqgf5
pm22W14ruzYJwAFq1RokgyKgx9iRiYaDcxdShqIHpStjyi9eK+nQIiHTJ97Xen5zjpthCKBTCAw6
ZPfJfF+Ox5U2iAaXul2g71TWi7todg4pNbXs6oP46Kg0rI74Vpsln8peQXG5KLay6hg+cqjwlngq
KXupGK4YJDXfqyH1RS3vb5HlveGwkFXG7PyyL9dSNLlRoh+knxF48hbLXnDst3X7bc6qx2zstce9
kx/zC+Ff8i/T+CO6kSaZSeWLciLg3aT3QRyAPNUbmmk6S1UnVvCRvvLhhSRytd6FKzYx6axNOVQ+
uuHcCpXHueP9n/vdEh8DeEMSn7hsVcmre/aszBLmqkkaAKZnTa4ZaENgDLLahFRRZ3TI5XXkkYC8
qrqwAC5DqB5hr+l0K7lZhrjmbXAxwjplHoOJyhky8msstU2+hk16jLZkTkyhEnFDR29kpmonaBmu
b25GEnVRWxoQ4g5Vw0NnV8DZy1zTJpbiA04KMlttyzycOhTzVI/jD2QFI6y4kY1e1CW0qKVMskS3
iVrFAhVpxGcarHygy1tYBgz7V4vLGVmcKyJkY0J5+ZmjEycGgArFAPQINn/qjop5OGvUZ8AZdvrB
yx4rnkjhePRDnonIAhTyuU1VnXm6kHyiXOwxZC2uyMMas1rDDH9fmAPdbaWO5EHOxYw39Qc1EMvz
PvuUuL1LrLTbwXqWM2PAw0V+qvD2aamOt/Amd1WOiMRsw7kv65caF3dvpMvpJOicX3ZcfNyAvQVl
WqK3u9BFTjsQ6waURtbdWymZ05p0RK21jstkuRH8FBX6sICVkZXwZbyYJiOb8y6IJlVq2Av9MZYY
t8kFEgGIFOUiteNXN/KgmORfIGmC4jNqiHSGD6UGtoFg1193cPDzrfcnwDMzcozeT6v1VAu2FQJb
MGuQB1F8LWmzTppNCLoi1YPnZLmPExKi8wn403om77stzywpDf8y7y+OybXzRuhI43bggPU/OURY
iM8lkRhbqMTWakIKBtGxQVHfmwtnnY2vrEvPAGYmdDO+20sBYFHlSLwcGukGmKMB5jpj4+onJkuy
WgvrWShEzwemsyIcsOJgxWQVTF1kHDQ3iJBEhysqRZLehO4ByO0UpSLb54TUrIWMTPZvHRGedh7K
fyWkieYjsjzOLaPKuc9E79HfplvnYlfUkqAelxjRxSLpzS72unjQ8LNkbP3bBZSORf0nd63D43D2
SdK5y/nIisGtvIx/sK8zBMkwrHSGc/OBh/N3o8maYQxWPFO8lVqmsnjzBVweVVTHFp4nstk9jVYu
4crpKdo/rQHwxbtSYaldyRtqjm4wTTkkGbsQ/cEZJAEs8BMm2z+q+D0Sp7qXv3iWsC0BEwBiiHUY
behYmpWpDpzCVA6mCs56KQk0i73ohnwYnFJuQIhhAWklIU8xdnc86awyESx3Vha9LVK12K4GcKQ4
N8AjSrOZLLsb7JohKJCgi2Y4kLKafg1Twe+B2dk3+KJMFUbKO97tx2gxWQtxt403yNqNSjPLIbs2
IBPO5Pmrc0c+RypXkcg3CYc54y+NGr0fHRwIfS2omBWxFoV2qv3zoInZIs3olX358OrUxcBqVPFN
2+idddocmaZTp+iHtycH8ZFd7lfnqbEvOD7KUbfGQ+C7vh9gU1B6y6u1Zs/FKdrSBF5rD+rDAOd/
OYUgPKONSURXgQ1y0a+BXzbj+2mbKHq613WspoP0DJsvUKsS9aq1wP9tew4t7MioSnm5vSa6a8fK
RUU5urnJwu6LewKiOssY90uRXMy8hzB4wgQyL2FltLry6Jd26/nz2KiBZcqCXwP8AgjnaQ/DtZsc
T5w7+xd/TQbaJloJnYE20NyMaEUSNwoE0kVXtUG5xbjkhFk4YKa8iw2toeEmOYivy8iaonQ4x5CL
ss+Fe+YcBjsSzmya7i9W3Kkktv/5LmEfBy9cOzq0i0CnqU6eae6ow/3KSymxjrIVpWrEPecjkBVp
5dpblsWqHSnPBBABJj8pN//YliKta9ASWkXCNm0S9ary+yRhzcePktVzPl4JBTEpsP54Wh09BiTD
cfjrRQ24njk9lvgdnJyAkDknbKRrg+PezHG798GlQJAby81pg70+I45PWZ7Zz23jPWC8B9oieW8t
XN+Gu/E85eDBIU+CQutv05Qr9ixjsynLGDTEEuk/Iebj2k9GeFL8bHX+ssfBfSk+Mv2E3UMOThT7
3SovCpTM15glMbVfQqfgXA0wGflxmVsguPgOmC1ObvscDT5iAmH4SP74AmVBlop+1UWvpn80iakP
stM7NlRaa7HtLctB7/EmxYa1Uaye+tTgR4Off0w25fypnerPh6eLIeA/lsISsn1V4GSpDAOD0A89
C7Dfr9MQYvfTqNntjKlSqKp+KcOjPYCJH7pOIS0Uqj22UupGahL4o4Vd/QCD8qhp+W+EYrppnkVm
P5PIrKa/qni3VdM7i0HpQK6tJrlN9dHYciGMzdIocR3slB24gNiQuP1bPR3E8LYMlnavPbL0C6HM
MXesdt8Hi+ov/tTbMi4KCYSJytEkGcOGOfczFHWeAUq0ZnYzSX14vuZWY28bYqv8LBx/plR09OvR
5bTtwchpWI4HJwUMxJ4Lc38oG+bGrB+HVG/l4dVLPfHz3CPrYEQiHnx3R9M2WTDn7kxDUWDK+tSX
Bc0JFLIcL1CyR6kvdNCOYVlFslsWYeilcOLb0NBbFIeh3lSnDDduFq26iv1Ysj73zVznaawGyfD0
WMiKfNH1hYPiBChTPKkYreda98nL5p/J1kHwZ2aQNWLja7Xeesv/uEtEPc6E9nMqz6uFj4RNmmA9
HGalfiqPdqa3/xPKoJFYHNLpqED9Js/zVmBTDNAHuXj3gTe1FtfaIXu7r1kVkgNriMIR8/uWLQ/E
GygzINVKroNBIP8xjTHaEzvl3O3XQHfov5W3cJK6fe6DcX/6w+kmXspPUMmwsrToX0CAE4U4+XZA
Ll9baajqR8Yd3vto9EkvxF4rVlc5J/0MEKWc4HL277gP+mcKodbGMkZ8sedb/Yrmh4TyifvhE81/
D1EMCl4U6o6+TYirt/+2566uoEh9nmWooFhytjvQBv9trG52LZSjCkQlKwCE/jOTq/BQER0hnNHn
7lTknCqIIISBuXxVj4gS8ekah1Y+31A1EDwO0+zjDYxCaoP0ypl8p4A8vS2A7a/NqjjbccCWJh+s
f1r5F672fJNbtUD28DSee13GXkTYgw8AjzAvZIjMs8JhlP6hMK46VEETW3j11hPFMAamZobWT+Q6
TPXIgOOc6j2gx7DeFx1T2a8lEcTWYEXANhqPeMSkfmjbfF6HFz7Jv+mh1z6fiU1rmsxEzW5azB/d
3w2LSsAjIKNhGWu7ibX5hduKoavxXfCAUj35ZxzGOxTG8zmpG838d7LpHJwx+3yNq4SenGap+2wg
w3CytfpsFQm1wDjHpq5ZEIS4FGKzfEf8tLmSvb/5TO7+JiO9Ey6m9UmgAkulOdIGeMK1JkxuSSlH
HHv+FxAzsHczjDiuWJ1QD3L+v00w+RxMEcbzqSsJjAb67Rt9wFsc9elLPDzMb3yDzuagoyaKRm2D
zziN1y+cuP5IIrTG/0y/qDxriapvxEPqGDZy2LjuebUal7zvcfjpR7UXpFGmuqMOuAliuig/seGK
gU9ydn3my+Ly1ZX0bStA3OTS5L7JFuegOnxdBddFmJldQRq7fmhnqXw3ng6Eoq6hVZjrw0shUuB6
H0mYru7mFFxFHp3jpSMoIr7yVkHQrpD/+RMueUT3n7uyRB04IrmrRRp6Rhsz16mlw/Xvv0k+3409
eRvF5iMQeTrQXMJ+rV+AuZ55w+e+PVotO9yUbDY33GGeQE2RwPeNxIVao+D8irj7QvykG/DcTHTB
f8OKQirRSFdEZy5o9OClLgcoBxnktg/5/ng3laxlR9vEPF2on2J9CNh9RxOmeiJ9LXaP2wX1m/9M
VGTiTL+9+ynfxDJBp7350rfxRteUYhohXnbT00Di5mM7AD0c9jTesRQiXeEXQl/+aCm+OmoBlyVa
cHibhlFbQy/xONHIBAF4tLzF6W/4zMjj4CZ1cBcaRKDIxPcdhW4EFQWmQCcLjCu9s/TA6uhMhlhq
lOIsDwF5BDRKVoXvKt5707OSgZnSpTN3bflSmskbl29yc8ciS0wS9hfPC+auD7h6PV9va1UEWVE3
KT79Z3awSv5Y8OY4Qa5Sx1/6WtkX312ZIdyV8EawQK//EH8F2Wqhz4MsYTZoxI1h+bS1XULnADwj
9ZftdfCSFmOZKL0EsQRamJ5wxPexonfcxoc+i7rvVyV9LIUCXxptWyNQEIO9y4mAvpeUfI9//lFR
6xcPAhGdqRey8gz3iCVpExCulnAPZhQZ5IbC7e9D2kWYugTCQCkcpQ3FgyTpEZHTMbEEdO6dSlEI
tn/IIPSlbeTttrOZxrHPA3sIe2u32oEEiUmWd8s7LKZjyRvREwRFmcjbXoOjHFCjoqTsP4D4PAfN
gmrxLQeUaBDWyl5WlXwrReGVjz7lzTLI9dTubnEgVgL+LC86H8P0sG/iZ2NW+qgTJIQPyKC93c+I
MO8eTTLpebai90v+ramH2uFN0+SjrZSHcRITmcGEdRlfPqyp/PEZnwBvrnGIXX0T+d5iL4mIivPW
N7eqgSa67T5uCqVKKY8dPp5VQ0pDG/chLamWaWQ8M8PofzhXwlQW9Mbc+5CYbPWPpAzNz8NH6ZCf
GlOrtS+ecd1MSIvhMXWl203RtFgYwzCrFuBLoipRpqeZF0oT4fj8P2CfyLm3oM78hxB23FZ0yx9l
4EvGDO3sEa3CAbpV4ixRBzYxb83PAIGuzLrClQaGqI6VoZyoI1faGSqrm2liXMfvy0VY1ukDA7cJ
HokYDzrl+AxG8N4mt5bZPyQlBc/aR9h4MZjh5Nd/At5m1aKW14+1EWFO2m4xNnzVLfsYsb+x15il
CG8AT0eWWLpMAPI8zannNaBn1FyIKdAlO8NpuieRxw2kSlhGQIsgQh8PxcxgU1PRvRznklSlGrPP
6c65Hogqhrz5h445IiDOPO9gSriTb/9N0Gxk4a4ruOlQG/hfwRL9tUtGjbZoWny4H+TWDi8aiLPk
eHSsPimpUBPElf+2uZxzmv4yVekFSDtQSRDan8cQ6FiYy77uvZWCuoSW24lJVbxk1zYgZx4oeR2b
DpP1ATPgCInkC33by5nu8os3pmw1F2ssLwhMooGZeYyVo5CD/vUylt+W0f5Xui/C8o6rlKfSPV55
yghFpgr6RUX0Z2ALdX/cpnEnPMtrqE6rhZmXtc7akVaRCuhnG1bZiaHfFoPqlhbNAWyD8YnNGCan
kp0/Os0SHXWN8pipAgfaGz36dBsIewq+nA09aJQZh7NJvobWlMuXSGdnqgfdpGvsXkeFYNMTreTp
oU/LaruUsanYdB4AoZZ1Lk/evjN0hO/gQOoga6dR24p07FZQw6l7TGc8+xaOTaZpwNqip7/0PUvK
ZCogN5XD8X7iM3jwQRIZzk/T6HuBSyHeiEqi3K6e9TlQv597v/OF8VXOYexnq0S016I0eJ6xSZ7j
tCb2xSiyen35Ej2nbQatVpmL/v06Yt6DeY5M1MU7Qh641SNfmfqHLBpqKmSQPRSKNHoQgZ2E74Jm
PzoaCnAuCuFJszCOiAv9mz9/ewrmHWNxpCc1Y26mfvs9LbWtH4p0dbW037dIXl454U0ghccsWg0w
j0qYe7g5lg46MjZr8pmK97nZq7/rDMfvFvzSwno3/Feh1zJ1y4TAJqhqFFY4QbKNa188ZZR1Y7V/
aMfLG6nBJmaz6dazkIw7ZoxkpAZD3uBsszhZozVfO4BPOwb+ESzHx2zk3xXL9C+5T8csmQQ/1gtk
B3UIEl77H+Fy3qJ9idet8vu2MG9OZ9WcReAnFFMzqb1UkfQEPt0Cvc6n2IIstyXccbDjycdK20LO
UOhK3j8/2imai6X4NFUCbWJT3b1qT8QuWV++AN5vCj6peZy1IJOky/fvk5BjmH/FuZzdRay/Nj/a
VEpXIMx3E1qnJvtOzx3dUT+MZhv3UItLmUYY011T+kL7UTuczXK5kMJVc0nUja19RX7NBL27iZ4V
mqbM5n73YKduSqj88oFrZinXQD4YQk4Ox2CmqIuXNCITwYHNeicIKPgUhfK7l66aJjeA1CXRzzzL
6g4JHnbZ2Qk1VfMYkqtanUupqdB3wkHTDgG93enRfjdUaJbrKH+xAfobRWbco0EHB4nn7+aAt2vb
fvK99M84Tx0vopkIaMaJM2zoAc9vXTNPNswd0wYuwK5PxTr3vbpP3DWc093kDqULU+wmbR8RJA0V
/4SzC/3aMnCrvxWk/VV5kPOTXAdQh9h/c9pwXFp5cq/adwquNpJmZyaWUjyKyojj/WGyPEnjqmJH
5wBPQnllj0X04mQ+mnbzRLyLB+9TWmqpUgS6S0qHmz6ziRxZIyZpxLF+tp70SMsCHYSCw68YFZzL
GDpFCqnFaAa85LbPlNIbw99L+snA0TBt+tJlXgRzxR3ymSoHNTIa20W7yJ5Sj72w4tZ811gBtimw
cemLD0Z0orDrq8umHXFIbRjfNVQfUaJHWCuME/94zBpvt3BoiJodvkHUTTpllV/XxOh2J7zZMq8h
o7Z6813WvEpFGEdkb7CIui7GC9xpoZDTMXRBTpbcnBCr15oOCLMiXD5it+Yewm3b/7H7cC0j1yi0
U1+DeQ5wDLbiJoV2J1K1Wz83h+ul5E3EnyPqnLesj2tTwz2zVbP28nneAdkKhn/kiWIBOBsqncU1
C78ZjEpVld0in+dKlOyJ8Dq3PtbddtGp5dlUTd4LTBvnVnwHkJ2vlYecq/pePU28oHU7zj2aQViJ
7poDu95fxI7acO2T2OrdLxt6my32AMUoeqR6EZJU0SJ/ECdhfUxFgWZpWTZtLlkjti48eUc9LIk4
pdIRXWnjCx+OXnizMVUF1Y/nbECbVE1VBgFE0IbOqAK+87Su4Kxofc6Mq5wNr0eMx5BtXDD2Ywwd
cuhG0sgyHqJPYfBv7MDIkWkAWclniUEl6tqJOSnPZzlR9JBz9YdFPa+Sgdo2wExUNjXp/Qc0jMCw
UYN9ys7n5lGwQzPIieZd2WH4uCGqHJtRhIR1b0zsjgROfd+QNew8RGTBQwdbr64Ki2x8l7SBQTKy
19eIfCeWR0xoyh48i1w9PufZMbwFvB0tBcNq2Uw1hm2bVl8aHMmMSnyFdiHEJCDcOpDPWvrmvr/3
BXpQoHBhVvGjPFl4HdccLWt4ETOzQtXO4Yv5bM4eegylEmIv281KTvURO0JQzHpyz6zAMtY0DyMM
+wHsGUMrfmoDEycEtrMNhHvitu32UcSoqbNxf92AzgPS9F2i3vpq/nB5nssS1pt96p91kxoN6DfV
IpzMf/X7j3BcRQg9QWl0GINWdKVx6yZTovcUcVWxYc8MpmHj0tmY6OVeTMOkVHH0zyR8Ah3ey7IH
PgyL6wnS+vBoCF8Nj+8YcbiD0oetddDybtMUI7wLV4gUrY8faVMnShTdbnyu4RoZTKiK8Lph0DCl
hN7DQcJuXjfvAL/ngEDCdfjLvcdUWQ16N/ZsihYmKfpCIJx7Y5vEebueA4zkWVro2tbajn60hqk6
bAKbdPIGFFHYAEBATPuA26yOCtujGBTZQhaHbno5DjhYgnmtZ6O2CapZsClUP1iSRMqSG0pNLStR
5tBjKUbC8/I0CQOvcjvjDUl+2P9Wv01z2rmVflppb32N3t2ywtC8thgA1RgIAAxDQmDSUPTnFuyA
WzfOlXXnFPmVsTagaUEsUGY0d/Lbfcx561jzX3YwsF/jXIvvmW7XyG3DVvDGNhyXB2M7BzxwH+kx
KcJnSHsGnELJNjG+D3W7KJYeBWkQEdSei+x3bO7n5fMx3pdu8n6ryobDsF4dhZHHOZ3p2h7CrghR
/G5kuWdECkrKf6QZqttn+pvZVfKF5sXv/Q9SOQHla9AGDaij23zYMFzpQ8MxerG1qR+2ACSjBMgm
/A9Y4AeqrdNlCzlLT8D5sDDF0VfysfVW8pcVDbOzNumh03w9UQSEV5nLDhRfNAi/aqz/iS8HOSpa
239DNHdTpMnJIOl1QppowTZBZOcnUELXhfnYJR7S5PZnZjiw/9ehfAaGxVsZEL4EnAeoasq1IB6r
4UdEV1KRq4NItFfz4LzvK//zmTEehKFA9v1xMwqqcP3C5Hb8eSXJOZOiHw3+JOEMubrLmDu42/8w
J6LYn8FvT1KEzN1F2mY9X6hrvk63tYNSnhue2g3sqUsk3LdIL+xdK5rSiXDNVozjLXrvF5XxkYbI
R3g+M2nSYBjg2a30FsE7AlcjDaXQB2jGLimcP54yHAlWnpnHbsTF4V9Z1U0/7xCbbvRLDH0FOMhj
dF5wHWM7ndSqqF64TLAahvFmIl104DTQqtXRZp3ZsQV0cGOiHjL3azlDgWFRTjnlI+uYTC+3U7mP
oGDHPby28/l/ML6WdbfUZap68frptbS+2KIwlnQL2/ShH/mzRetgNx3q6V8qR/hsF4rREPen+nXR
yG/BHpooIQKH0l4Hh6w4GM+s9psl7nBaPJEYOG9FM2RPTv/IhdeP346QyVHoojtcbY1X4LXg4EQ0
1lcfUap4vtdo2hTD4ivTF//0v0HUYghhSqcISfu9LUvXZggTb18pzAChZwOK4bHh1MPTwt9N6Orc
10ow1+viicNIDSVBtowZgHGayY+jqd63dMZ5mfQULww9K90mksEjd7cyXNa/ci9NFI4hv1HIP8ls
CNXTiskiVYF4DH0Fm20Yv5vQKMCuoKlJu+/PsJEYZJadPcIso89uz0tus7leK1lvphfTTrIj+AqQ
eK1KiEnaDlB4nsDlfRyGiub/77ibPAZfmUw0s3queY1UqeI4AMcN+hadkgLMuEbtJCIe4Po1TeyV
ZI8p7t5gzM+uh+NR30998guGw5vkU+IxY7lvd6OXI97uu1q0pbFEkooAQgVAXpgMtHGxZBWKhEj3
hbMq30/c4G/Ppk9uYPIMgW0GoS/Zuk1iVGoWvMKvPMgyXpoXJH0OifaQC+h+ByTK+jgm8KtbZZv0
8X7BUOTBj5l9WvF/OGuZTdzzWD3Uyx0aGeFvDFR5XaYufW/BCFFGPVRHWR3ATrshbDfaKPyoQw3N
Zm9k7Vv4EathJBJkq0SK94Vy+zMLJmWxsgMHeKj5thftAXDmvtXoWQmjm+M+ATYY8nQPWJqgwvZx
K91kQXY4engGwL3Q9p/j4WCbASVgHA69qNaNIhM4gLD/Gwzn2Mv+d+BsTicw2dL5PgL7//Pvdm+z
XYkV6vSPaA0ZFtCdygNjVJ6ewEhfCIVIs9iCV2QaYjC32d6j78Nfo0QBCGRwRRKK06QVhHYs1Msx
Vno9t6GZStLS+qjj1DhrljBPFFxvoJV5TCnvAkIW5YWSrvyym7+W+RcJ53jaZ9/I6u5GzXuRwTcB
YhJ0wL+bLpyZ41Zcqe7Zy/lV1HdHapsTnxINBbjDlEga62LPh+p6I0fMVFNJc5E3cN2FrWk5qsVa
GH99SUzl7shYwOkT/20S3utL2BKUeI9Z3emt2U9UHM4PxLW0b9FGW8DpQQ78tVOBGf08QlI47Bb3
deRQau8bIX8KyEEIBhU5B11ioPgMCWVVS4ppii381a/iCrMcdLq2+mozaTtyFoGewp0oq2yX+BOl
U4+MqNbuvvfj4Fey4JSUZeovERQf9j7hK5WWuE2qqKQbuYyIIoNtdvhTSZMJCYSH3lBxfofGrBn1
Va1M6TlnoaEeE7HBaA4VIy/9UhN7iEA86RYGcqCAiIlGiEJ4EaJA+StldIRQrXkcX6ZfEziA/NIY
Hbw6s8dCAejC/ggDoq+LN298RXrLZysz/dBMhecEFyhKoApCXHSE2VX94LUV1UQWm74e8zsP6CYa
5tXwxIDwpCWG73RUrxocn+Cr9UMezHS0QpRP6XP6tHWgkH5eqCdO1wHKSJsU0NwIZqGsFuKvnrr9
dSoBOYf+fz94Cteh29xp5FYUWeI3KDveF65w4/knXiCNZu4gpb1DmxYYKkkibVxwadYJs4LATS85
ppaRaju1s4CEML5NdJKrBH0IYl2C3E/kNwhkCwegnFSvAWWnc/ki5BbdjbtlvUJV4Qfm7PRsEyP2
c08OOoJpmTabOtT8Jr/tSPwChbBnQOJyqVK3roniGJcSuz4U8kAD5TLg5bunMa9CuCMdWLmjHgxI
6v3Rv6UmuJtzBbsl7ZNE5FE1+bErB70++R9Qt5YgVi6jGaOTYd9Tw7GyNPlbNKbmdqAtrNReNNEB
SIsfoOzELblfSpT8290aLIRjVXjFnsZTyRM8THLyPq29AP0BWzqj1j0wsXiMQlRVxNEvbDGPmnCi
is7Tl0HSLPnHlPILVUPsNI7JHJ1drfYQ3aYPQCIv1j0sGD7ymTeGYaMI/64pYMjRj23OAqownh/g
/p8h1HPPRtqJNrtpd9WXS/IS7P4o+PZk6trU7Q70B9EeBW1qytrcdPGtNZbusR79SqMsBIgFNxRs
W0j63CTxtuRd8QJfEvSBwKS4dFwwTc1gj2LtsNyAPWuVVejTibFwhjRlIJwb9vEFTDBVHzt4MlNt
mq/3Fj2AJa95HhD3leQxzECAgG0NU5Hc2v7Pm0EWVGzGHI2JpOk6wV0Rx58Fr9kUhnFKjcnjBfMa
IBl8jafA6xBEsdhI/Uvkj/AFhh7aFUery4FVwFJHz1O09bTm7EmGyK8Zo9AvOj1mqScfhz0kNqhR
+q26N2MYo5cM7owj6x6HvzaqzXBskUMwEiRlsdGfHEH28WQARWWFXAcb1bVAaQf7yJJlK4AvMUby
WLGEGpCeEBVspmnoX9GyMZUPTHpkxrQaCt7VGdiT8xy/oEEP1rgEF50GEDBIBDB2Q9nYPI4Qg5l7
m0gZOGTGoPiTIQVj6tDs2fnobOy+r92i57BPQiMd8yEQwf/nxCpxl/cUkMVYaak9jes29l8ijxYS
X6U4cdt8uSgztxxjsag5k5c8E2i8J8EcIP1c1VioG3eCUHlDQJvjY+0+/peWtT9DKuSBLf011kKd
lZzDVkJ0YZ5Zv7NshbydNYVcX8m+hKXiQqrLR+tqIPVQMMvkUZUJt7Dd4VUZ3BvM7SN3jkASsskt
yCTlG9P2UgSOJs0JLuBXMSHXGi6jdfVYx25fBprmIuB0gJmQ9JkcCCvz/XJfVZQa3bxpuYaD//7x
9cUMKPC3IFnCyYyB0vEQqfBBNUtcRfDKZVIWoIXOo9ibOZnalsZ4q5TsHOuDeaJ5tTa9e1udrI/9
wZ0YZS8tAJjjuhN5q21kwK0r5/YlbPMJZCPaRd+cdy22BnirdBQhhbQUOZ2cuHqEfUQUlNYbjL6D
Sc10l0nWG+hcXweLgRLCTqA7g9woxEuDRbE3lolWKWDh2z3LHq8CcHQmj3P7iGbhnul/+rWr/oOB
V47f8nWTif0+kULqNLWVOPO9eejfSmFkIdZ/gHuFmNanZHoqm73FLZww5a2B0/asB4l4Dec/6GBT
cX75l0dZ3XlpOgc4hj3ig4rucKwhOCdZgc8i/3K5ksTG7k3v+oSasrOpFFS/p1GTemJf2OYLIIyb
5JXtwbZmHp/C94o+nZYL2XSfrSzcAcg1Ijq1QFLWkD8J2Wemzv4MbdmojNE1btSURmfjEcTJHs3e
wos0BDzpsC51nsaClimkSeDEx9KYhhrmYURKrYZ0Wc7CQr3DC2hR8Sz1qjTvLnYqemQuUceRJ04U
Jp0B2m1RRArhZJ7G1DSNjmSoheH5YDEe3MVnucrmyRTl9MFDTgAZVpV6lFh6P0XdmSmG9RjJHrs0
pr8k3Yqnfs1EMJ3gHqPiakHnZGnaBWHUhBG33Abe3mJ/xLQQBBoHfvZ7f0Wb62miKARYgNA0cevN
ttBWfT8c3xZvX90XuLHUG5zsFHk3Zt9JbsRIfydAoD6i+EyN7jhUym32gVMnWCzGGnZvhLtWFggf
5x8OITD5tHxUfZcANZ9Xg1s3xdIR7Eg3vDWd1gpcO8rj6QQwh1gbGTeR4Nj/jxexHobpEBN6sOwV
lBGFdG2ExU79wwfqdZ4bVNJxWrP/l/AABqREiUtWphESbIo7s4sSQILUW86/UuS22QNGG9uKjnsE
oq/nrKet2LbXsH3PWUB8YiOGaX7lZA+I/nnDsHV/SNTcQEQAiuQQh73ChnASEaKgoDmrwYULrMfx
MG1NBTs6DSAl0URIoBbcyCwi4JAHdeJicSW62/SVs0J7Xh3leukXwra82XRwrh8HBrkusgzHwbWW
2lZDwKHIuiNgiW/RUApHK6X9+ruwIVSnpfBJdI1V5fUIlu4W7pvmXQBEMd9tUU0irDjGqBO7n7Jp
VERIPhs/VlJLwLenrPWj/3QYLA2z0g9zY2BatOqes97ReRF3LCbBk3Vry8Sr3CGaRF09Bn6pU+7W
tyioNZrNaLcasnBgWEzetmcPZyGR/n2usnEIHIpdJF07RwRo1S7xwMyBZuThkKV88V0jQk4Yxvm0
mla1JPG4Fc6+MyC/yKtw1nvpTFNLRC4cSMXHA5gYjwOfD5xEKErD7kXBVOJREczp4+ErOSNPfThg
v40nMKSadNbEOO8a2hIrmH5fV1Smo/EjKFH9utcV5sQW0Q02EmZ53WcfBCW/9asi6F2RDmzIRdjf
8dRx1vv0oHZJa3wXp4yBWpDY7+/SsePkiOmzji6d8dZ13cztgv1hWTfxLGLPHlzbXK0gXpvzrRVr
PGtr9zj40bs3tKOJPt8vHsigoJaUsG6mIXkO7NSeEhUXAER7P3afgIzas08lwJXk4PnFeG35Gc8l
+CWCCPscFDpA6YaoIxZOgI27N0hwZRG5P0IbQ1rWH/YhXndPGbTuqJ7aIeO2fMQH7OfyClYYadlW
7g7n3utsAZBh8J47sctd9G0HDKYVriV2AgRAJbWG4ay2ePH88dj1ov+5QHn9S+s2Sff0fz+bq7rM
KevvdpcmOLHWTVbjJQxJBRpP/igW1rK+c/zOyDKmiClvMuI0kNl4vqFHa4SnpgpUa0NvTdNqOH9v
AHCdbAT/jSTYB9aUb1IgWu/ISlsjCX+sBaerNP5ZHSRSxlHK5fZsmOok6rodu3cDQ6Oo7172leQf
MMC1BKK0ppu9K3BLnHsFDCQf3hqe6msTnbU/IQiIqRZNEguWWEhMKC51XE4tKHUygfLP/rN+O/KA
T6tnjBqsJSo5Pq3xS/iV6tSDfTJwhg/S6rKoyc36YzmI/QCGf+MghnFvbHdgmGpk04ZyjJVG+85M
tbfONV1BMwYxFzRRYG2PRRTkrCWaTPy8IKoFStaYJfgHA/qDR/W4qVM0lSnPrPDMocb9sgw3wQtc
jkZ7xvCSGL4t0foq+OVOR/pW3MWpFEqm8D+M/j9yJvybkRlmN7HJ+E2S0pvQ7lWBaHlP6vQ3hug4
/EvCX3YZcqrFZNqj4BmY4VInEu5Xlchfi7VQrBTaIMD5Hyrs+LikJjZTqbLwMw1pmLjRLj0QMUh0
izg8PLL4JwThw/cxfPmy/GwE6NcGLavZnkYq8TUpoIYZpArj/1ufx5zviPjMyPhhigSOSdunO4i0
WkJ8HooPBeUV8wklDtD5wuqHMUOcKDxG5RxMcuhH9WRMjseSwKXEsqPMvHMEcqII77CQSZliXL+E
XnSeUX168MQ8dO17O0GER26rvYrcnerKPNkoZ9bRKXfFYr/MxJ9nqPasFqx8PSj77mIHRNHph2Q8
2T91cz57l+uhr/axSndcwY7rUTh3CHSeM2TwNz7YmJG+Xm31N3pYPQTkDPl5lY+uS5o2Ce1dLNsf
4/gzPoviWKVTacnq0iqVg05Jcq/b3P8PC1S9hpnYmg3E7htJeICkWfiLzkqWauzrdnK0eenzEYpE
gy/gIS3LjPI6gdHlaBrFqZ+aOYb9hOUOSi2btIkAbgypUPcOvG0jLZwFJy1Cr+aLzX2bymnTH5eD
Xhx2hTVf3XaeIuIbVDVUAhwhV5UPjTAP0H3zUADck1nuffyv13PkHYi+1flkt13stGZ5F02JgRij
Yei6DLY1VsxPYZHvtOcfeMMF/HgFbpdjsdo2BEVpi8/WBcMjhqX9iZ5zxcPlSJI87N8GJiEEzNc9
zTwsp7rcgcOL/PEKISG12b/DsyaYBvSbaeaQS98EQsJcQXi1ZhpZBbWuvZmo48uieScor0i8EW8z
JqopsEAExeh4OIwcYLUR2dM6/xeaOzI3WwlhaykMUp2WPGaVCmGT54/JCzgxgW2GhT02JCHc4AgS
J1kKdcPNaxJvz4EGZS/fN+ZrC4Pbrsv+AIRwLA0zbIT110lGInuyCxroGZ/79IiBWTSxS10rJH1e
1nGcDcKNUnFUAvJ3c+w6d5CyX6o924dVr+VXp1FPGEVAI6DqaVMy8kzfg+ATwC0jgWbWStJRhLeS
WwEgDswNACudkocJquYcUVih3ARNBPGG5n1FdlegR+nr3ti1nQIldLT1VrMeffbYJxLBHOQg6MMQ
V6SoDEZa5FkzzudD4w6dDih7bF9vzSKYCd1X1/1VB9FbDOfnPOOJJtWCKjYG4DqkwkPZj2Vqerpl
aDaaDrXqE1bXYZBOwAKojw2InwCBjFAQAWj2uzHBSaWCOqfHLUbbC4dKphoptE1yTCpKdoI4Afep
tSAa51u67UA5AkTCahw//zudi7PIU/iklgKLEEDGSmeJZTfEEOeBhp3+0/kD+9J4Zn7xEOUCPPsb
uwi8cpvw6EShVCHncaZJW6WhijzoV3C/btH1T2ZokQT5ypyj9QSCJXlTxxo1dVX++NQ6vw+082lm
KLtqrUF+AcPDolWXSe1NualTqRxdLrj88vVm36hU+P2JR15S9zZfjx89M2lpNALRTwVRoyvOoeFn
NExjKBrq/D184GqzROwIroP+GlK+DXu7D+UZFX+iU9mM8rfPHyUAsaarktxxXY5aTTS1ZrgymTpi
0Pi/V3GkD8LZEsHL0pFLn0QhO66KISrsh70BOTrunZEcYLjnrAVjUmPS4P0jtQYHQMzQ65nxYdin
S5+aNZlOHdFY0u80Z/heUzuLt5lhwk9TAxBKjBfT1yAX2qmroEyk2E/3OapqNj1ujfYKfIQog85G
T7qlIAzU8V48lVELCmj0433OP3VnDjdB7e/qVhHARq0pCfAiWgrv2M1sh6ZygKqQXGEqSe73BE4v
Kv5+k4ahiuvtkQGwhgMO1cLEPAHIJXtIEewASt0lXNoFRzxO5LkCa3boB9F91KnA9ax+RzBa5EB8
gGx3eO7xK0nutPAmWgAWlMyrCWsagmLju4YFVxl/QEjA4S3TBB+My+JQCHClPsml07eSEsDMm+ve
XafvzeJ9iqFbGbwu1GhCkFRHBTT1xhH/U55Zw3h8+BfNkDnOexqJcWyQ5qGcDixUGFEVfW/uo2TZ
7lIsY9Is07XOE98kee4IEzow8PrCXJYE/0JBX0XJ5qKXonvalqDAvpl3rz4E6Hh03IaJt2CQxhqB
1JXv7cEg9PtNUUfV7b+Qu60md9bBCFJhf2I879OttYvwtbpzvl62CRVt4ql6BkWQ+pKGWly2uSiQ
kfFMSY8P3MEFnKdo+d6B6JLz+tujI1Pe/9Bx4lJxGYn/l2Y67MQD4t47WTBHLeCGTlb+mcpqUhiX
Bg7nblxpKrHTTyYZVOdox1Qex3JvByh5cdh6ItfyXICcHGePvPO//xe4KKVGbdwutGGCMIN1ZfrV
VSitPtNM5KWTLD5X43cURhcN6ZQEJnZdFiI6jvJOxyp/cRB8we+LDysG1r+kJqTlK8nglsL7tGvD
VEqTxUV8deN+WHmLaK7YZM38YUv5+1lkO8tGTprmKeFTDrz1w8xIlj1NGdE4rqcNTBzWUJ7FO4Iq
hoaOaLFf8KlG4NuI0gwb5wBX0ZGcpWXfYW0I3XXG0NYHEjg6d+LB2jgeb+6AEOW3ck8Kzk86PWXe
0W8YAZ+02nkkHCyzw4pzyS5KMZPqrfb10wyZmAg651ARjsJkVj92EEpkKDtWzoGRXvEr1ObFZDHV
GbwpYstMkvg3JfhFo4z/OURb55HC4navDbceh1X0VKH0aIHRiN2fKrQCAp9F4Gl2niSIJdWTEqZB
7g4ro86BPZGfmcRui5KBk0GOHhsAd9YZvBqa+VxSeg3KzEtmTBm5DCyfNDXo54WKeTziJxcENM14
40rVqbMSPCn2Sy9/s77IpliKCsrgImUM4M5jLpwDxysWuzB/cMCC4HupDKQ2MhFiB9rAzZWa8N8h
YfbhrxXPmbncNtlE7+trzC2Ve/tR6BmfcSwTtz7ZQy0laKzy8KqAGHYMZIKRPH5QKbT8J7CZs/NZ
tKuOpYP7dc5iRuiDTrhZeHp0kxTiPXWatmHRy0J0LXQYBorCFyXweDhgeqx015KcWMgXthj1mF7y
F4U66Z3INPEfPw7NUkesLSF9ohYlsEG/GCIbFpcXFj6aYd1BpVB9Y/IfnrMHo8rrIquXLaS1L8fY
0Vj5lTrPGuUDaImxJhlMKaKgY81RJaJdx3uUrIzmhWjIop2mYewXgZAelrEUn4uKnSZSo1xuXPrW
xknHGLCRSEPl81hs4i2+a1dVwALol27Biuf90bFLKZj/NZcGgWvk31a59fg8v8+CF9xyi3oek228
1Ig0jLTkezFUk2GiiLaMj3uiUtu2M+GHupDu+X0/okq2qu9bnu2Vkw1pkwA2erMF2jTkVSznQp7W
ZpOlMzHoIvKTqDVF8Wf9DB1r8TEKTdk8omDf/R7IOVq2Xx4uulIYAo2USqcnc9kRe5gCoJW5hCiM
4A1jsF5qHXvzpjREM/9cRPKfUSnK8LYw0NEjQkxt7bmmQZ8BMQBvB+q3SRgKt0TJgdzRSWlZiipG
zjM6aGXnTRQTNGB2H51ncM113stvfY8kmO3cYY6JFHQlwWLirqp8IDXKWPy2rGH/c+L30djw7f0q
r/S9JRbeZXc4cfX6m1zgnWXKc5N9YTInuO4CbgPysGaeohiQQ17oZtiMIn2P0bNuOqVBQTkDRCfK
HvuIkNanhSzwVgFLBXJT6y186yCdjLo0uOhhsNaH98WAUKe92bQO26TUd0avkyU5GYUE3jvEjb16
Kt4sXDp22sTqc9bp551ovsmAeVlxA4Rt0lnK98k2I0JD3tJZ9zICK0RwDNf+fJI6zif27wdRGNPA
h08FL6iYD/AZ2tAqsQSid1j0bX0wZ/VaW/x5XRWw06J1lgQ5KojgbSNIO9cxU83i+GHz+n7/hxcj
2+zzgtWsm/O96E+rmMqX5WNhV5Mn47nBWAs+AkKHBiYRQCg/zRMTnTkUbdXFsKDp++qC8Zf6Cmcc
Q/USioYtCZ1UkruOFyJ0owgsLF5PsnutmkDL89H+TjHi2yoxND7wlhXO+64W73wff0Y/laerkYvU
BXZ5aSIsOXpkxkvuq7mfAuFxz6oB3Irj+6WIHbkEN1kCQiwOsnNxC3m4fPpze22QGCgjEfBQ2Qeo
nt/E8KmJlKHfsNAOLmZaTEPfyzeKyro6H7IExd1rXJ6hPokPXH0iQq4rKusbWuLhsvU+Lp25Xoi5
D0bJSgVqIPV+t3tnekrKXWhW/dE9W+SWy00UeVxnG8FkysJ4v5E6U4FY6ag2OfUy6soDUWe9cvc2
P1YPHZJ2we87twy5e/U+Gshq4mZRmDE2hJLvyr7/bzj9hSEuZaYWXNu28EvKRdPD7KMMY4U4rExX
IxCa14pGj4/zEWXpYLGaqEpHg2BXxE8TWMFQ1ZysYNKWcxyrWTYwYBXyh8iwTitk6VbcAAGzz5Ij
2y373TShHXyr02V3mAcRVjbRMrAtWmBUezajiJIVlHatQCurQ01TaPbIF5k4DyO+cWJMYhCAVdPp
m77rAAqcwAtKr92ROw6SCb7JBQzZ5I8QSoKO1j0jil10oGoeYrklFRSCFwgRYAUSJqIngqN54mqV
Pl+l67q7mtla6DJzlhFM2YX05SE8KqYNLEDxDmjp0vZFH5TJ4t2qcMuG7GjzJ7HsfmuaUeac2wg2
JkQJekMJBXWuF8rxQ8WUi5taT200WMeLA4xZvzS20Y6dSIZ8LacN0cijTvp3tzDDCpEqtF2QN5qX
dlvwSHW3q32klTY2WwiRAySltywoiz0aJFwb37qANRiLwOQLauZQzPXOhFfZXaGJWm+naO+q+OYZ
K/pmQYSRUvt6ze8t64VJ1TAIQ3MCssD7Sg03MmwUyuXl6c83hQJnCDNWE5IqhHJ8K6JA06lxiSBB
rYkVXc+DPZvNx4iCKJ9v5N1kjer3usTnvVL8qDdIBbzu7U1nYgRb813WsjN+NgjjLJENbsKRaRZq
OYYhhbqnLa15wXJCGenNkEWnIRxspR7BD6iPvwZlgC5nNfN5tDKY7U/bExpqrc6zqcLEIpBf9Vmk
yrPbCx+MOyIST5RRNJhVz25k2x9+o7VMj0ikjxOwUr0SF66+QmImqWaFIrsdCEEGvLkclfEO/5uZ
QId5jGBjz6DCVWllUKEUJUgSwey52Dqv1VrcgDwbqG+ZbuxlucsT4713Pg/EgwXel5t0DAafmD87
Hi9vzbkm/9UhlhEIn1IECx6s5KAsAmimkCm/1trCZKXWBBCSUUgyvGmxXOmFcQJ/PJjpF39w8XZz
NsMvUMpknAzDS+psF2O951jIjGsBOpKYjNyhJOGdfHawGOXGgnuLyOImfPtIZvKYEjARJ6ZKa2CB
n8g8x5MKPN5hb+WLAj8gp5YHT8vV3KV/OavS575s9l2Cu4z6C9YRgzCCIuiMADkIPocdQ++1zJYz
nGsi9PvRsQEEg+4BPo2Gj7oxdAgJ7YOHEeQnwrMMbYmxdF8CqqSWmSo13uJSkf/93wfxWRwPyXWs
oq8uiguDvVIs2Wz6fEyTIgVgjxVSsohv77HU5vUoWJPfjmUIBxNmlHsBjQtkHsUtm2e8LubLdXxG
3JKrPZQutrWSj74M3RSVE+PD08xXR2kpFs4Z6xqAL4MWGykz1bJzadEM8d68ySombolsD9knm3nM
NrrXfPrG5GGCSpQdZ5PenEzsdwsid2fCePUfKfV1DLbQleBimxvfn0bukQSbLigayXgG7ClZ34oe
PaVfVMAK1RfGGVlp3Ze0Eup/ATvPe3QNFb5EEYb2CLm+kgg1DWfZBakNP8gtZzJ1GLkqoJvkKjzD
bLfIhVHDwBLuKI1rqdmelZ/KiWHvK7OFbXnysWkmAPUJeO6ZuuV+A5zrTboX4GP6tcFCDmvrOuI4
je8N4CQ6tP2Ccc1k/7tVcuIfcgeASftyevwZWapoB/JdgnybSAQRMQjDmXtuHbL/+v9qf/qjZ/EJ
3w8t5/gbYurvCf4QHeQ0RUh7ejiOkOZKbamtsDwqDUmtM8bN7W0MJZ9ZhRFpa39z7y2u4v59Ws+4
2Qhplxvj2yshuk+U6Ka0tqRxRgufPVFwicmDfX5achUOx5hXVvksGpWqaGsc3kVBCyektzdnXzPY
YvsWWUxoXQLlzZAcbbRGk9pP6PDxHDEvO69yP3CQb47uPzk0LBQ0sqvlQk/yO+XcpXYKQkeEO1w2
Qs55J9vv5ym5IEeryII49BTMRM6ajVVrfQIHMoQo58taYfJLPYyaQeM0TVyNC/V1ADXs0jsMc/MW
0/tp0E7UZIrlBvI2YZczl1SaMnygKaZlv2r79As6aqkhXJ9bP0aRfajDJpi4AoTio6wWVXMRX4Xg
X6JWjAz0Z2s+6Kwv4RM2+KtkiYv1Fzs/ke59D3049g2abGvwdPRAiqwhhH0fHcxPtHqLN088HTU9
5xah2QzRMZViipWKjMt51W1uFv5rTnroPcD++/NaHJoO6d6GJ6U6rhU0956PY8tzBjTzQQ2P8ij8
yvjq5XCDorr/cTm74kMkHozoRC3f680t9g1kFwfxWjKQ5gVsbrGB6/YfSA2jAVnPhoWwkd0b6m9l
xJXQviOt6V8sUhfZ4RDmNVhGj+WyHnhsDCZ7vTpv7g7SIyBL9xFEfftWdLjaZ9E8e6zgZ2lmgzPW
bLe/blFyw/dn1HVtL2ljsKaeWNkZzcO3OWkT4thQj84fpwcf0LTA+Jmi/Mkvsf5s998KIs0SCKTe
bbgOK+M5HBYhZGJN24sEdCmRwmIJ6B+oeviMgSEiQ0BrF/Ay+e0e7HWC+9s63QawAC+SljUb6rLP
MoJMFlFdI7PC2wIS/q59XHozjtsVbNNUj19ODRslp+liyDjskcZLbDfAnLO0uUf/LcLpBBgGL1h6
qUfPEdG+UzKT88vZrsu1FJSn6F87K7szeFv6F6j7RAW5B0K2YGowKMu6rKUSce196eDxTbzvxGvd
vozAqI8BM/P242/E9hhE2g+b4qF17VuC1RlH//Tho4xDrBEhFGBpZ/O+TcrK5t9uprG214zzAOcl
8xP0Btm4tYI834/s7StFYlVfYZnLldHcOx0IH/MhPLp/5PIsDeXKaitrShVsoGZz9ezsJShnRf9G
ZMMBpdnlyewInvBRRNh7+m4RggzBEFUPhTVxcMOJNhj0uVTvNFwuLIhXajF1ZEbWibKl622jGadL
CQzHUpx0YzfDePLduJu0LeHCY00mVlQtHJxRBuvKrQEcxAzZujh9AAhBxg5+JRRGaSUVfKqbCQG8
f0i1lbcsrzLi1AvNh2aQRLL0HcUAL3uzqN95+WRYC3PvT+JTz4PcSHBlJzPQWvgTJq4c7H5O1+c+
/vmyzrbVrELdRmZl59CsADBmZRgsI/DxLkLMJC/sOIPrwIClKVkgUZaSD+l5NgmZle8v0Qdmg0rt
14STjxgUOjsEYthEeKCx2QVoZuMQ5HrE5tVfLTJ9bk0E0kviFlDtmab9zVPWb+by4Eh8ogFC+uBI
JcStF4OMdmbFcZkueoyDiXEHJAaSVuqf34hg+6N3UHi2RHGQT4fxVogZBQ/l4dh4VDAzSuN2/PvV
9TiPfUw8mpkt8WImHjmzZNGUvvGep+13pAgAHYvhAdivrYbBl2Eio61Esc3DgsDzBz+dQigulM2W
zTr9Poqx6eLoZf5fXLiloD3EqrwFNEQmdDLty/c5+SA9giSm3W5agH1LE8Sa1HYGpp2pcdbNMkIR
SbFWnninLBWn2rVS2YkiBVo6MSaEwN1yFQt/0KkKKXUI7JwHZu2rghzPy3tLlJFEHVvl/1JmZqwy
1kNg8SNY1gJ65k7xDS82XJjYHL3i1fl/L9jRyoDXHf4+Tij1xxNZGWmm4fCPAlG4jNgzeaFRt6f9
ktIntoPPri+LTmwW64EdLtAdvAtV8u3c353XwaZWrzTw8wFs7FfulxC8NjwmkyiHFdY8ywSd5G7L
Tk1/pLI0r6DQgCB3nR1fzq+Z9UFmAU7iI0kc+yOoupOfnEl6ecZkwB7eWozMjDApJLLSbGHjmq/t
IzKMSELvfz+IYygCuSHF4gHdEqibta8w2N6qF0saSvWO5zbK7EVOnXkJEN18aqtuUkKHddO7Np2m
S2h1kFlUPYaC+wOEpKw6RDTD/yPctIly0vJYNL71qHZydnLA5sL8ClUNjbogdtEUm/7zCoz23B48
7VY4j/iLjGnyhrXEi3R99XcvH8ptxlgWjkAgjA/FgXLfRQQawcomRaFJHlMeLFv1sibRekYdNA3s
0C9l+3JrNvdi+WPIlA8Tfs2sxL3AEb9FYGycpkF+fCKYvXsSYfrYVp+POwX5ED4h18S34N++0/Dp
LCw0ZAL8THhNHF8nAK7qemAzF4bWKb03IdO3PWy7dEeajHTRi70KwoBqAO1KHemfevd6ZJFMbxr+
8Q6Pn7MAUm2a16x6Z/tqeO2/O6J0jKs2vw5pprHn5Ce1Q/6oQO+CAarUnLDscaHpob7Bfh/gOwDT
is7Vq7leQqKuo3FSXdJp+d3ZWJXnCKsLiu0drGHwQqBqnyDrXhO9ChlNpCjUBfz6GCbNLGPIG3pP
SquH3WN7bZy/PTNyjLqhut2bvX0YS60+uDSckAxObgip8JXnO1ct3ppf3V/gbzL8EiG0Bw/oHJbk
crYXfs+7AC5odEx70T0bPx4/LWmUt81RYQpuoKytoOoyOHxPVQitUF27j9z7X6+LCHLKE57SUi+l
VQL74mHz75qNGILujhEtHoRhOJlmZs78EJaCaaMLvKLd8A8I2j4UlLrj46wmO0fl5KfD2eo01sjp
DCnJGjcCX17A1nZylwF4zOvm3oc7c8sCOb4p6nABQTg7FPgoy6exd2bR9Q2K5iY8TMbaze5OJBPl
KaXrDJRQwXRXLcQDJN0PdtOyegnliuvxWn7hhSbPVkw4a1F1lwN9tu0tyBuF2+uQhD2UaSdq9k6Q
nrXNJC9bHVLotw8nSRgZt2SjdPCSARWR67YxW10CI9N6cdloprAabK5YIM9o8tGOPc6XZ/S6GqJ+
oFIOH0VkoCrxpYCjd5y+wKSgCymIJzFzzhrFictfpgQ9ldighb0zJE6J2PNayoEQ2UGltpxu2xwQ
6jTzNDGVZTv3MZHvDFPDbgU8bjnzJNu02MwVE1cC7g7I7ohyj3zSm9MOhzn58Q+g24vZghYoSaA6
2wxiaP9ccPzo3BysMPT7H1j5onPemkr9ybYrmOdcqmgXUaCI1LCPyuJxxHfntLGGkUNhRkV9V5gJ
b4HWB/DPIT9oqRtiAsY9F5WZUL5XQe2IxiSU5WnVwx0SiSCvBgss35qmn2ShxH6+frBtUYH2Oa5i
AXDNFffKgNVFrNfjST8zxSUytJWDXVkhUvlhlebrROQ17olDnuK/Tbea2wtB8AEIwa+k8DxQShov
3NuUftp6QHEAlYEVn+mLamJPP+EjXkqN0z8PGpWIsUP9X0CqdEn2WZ5OOyNu5xR3pei9PtTMg4Bg
UdQsEF50yIXpjBN/U5u3hs58jheYxUOBS7M5XD1G1GWwRSiDMk3idVSwB8g+FccZIrXN0wsjogEH
gVXpTbPjV0ab7g01+l0/Xj5E8A9wVnuIZQWQipV/Jm5dJGplKR5iHuHhE3g1C3xopMhHpjaJqpfD
zNKYkQA6O/IR1H7bReL4swYwrYxiJBz9eNUpbbUwQu3MaKnI2mZ/T7y+KJwxjtCwgOyxHRoz+xCm
jw85y2xoPN83Ell+C1y/4t5jGcdjcvzVK0slWXqn3cj5yX1ca2HI0g9f049RoC3j+JNJXZ4Ggxpv
NTrz5seTOWSRfz1papk0J0zfZEEg5iBoLrirLG5aSlXr224gfkLnpJ7/xW9pdHKTkwz/jJCy8PtF
u27uxLunTVsqY6rD2Fw3f5N4yCnuTAFxqkLS/f5CeRRu/9zEezhVhL7Ph13nShjonsMSQFDBr9ML
yWILkPIIoaoNZ81MFvn313oGMD6D4l5OhuGfPLxra9mlUcziFY8MF8n/ecowOyNA9oaZFNHX9N1N
lHflRq2ijEQTr5Kq5Sruq6spz4cSqQ9yuElBJsehqlO/XUNcURldq58Bm3BKY0Jf7DbGOZaLq5po
aGxVphnwCA/su0Ib/RDDCpW0r89qT/OOzosdtSdKTyaPyWuZ17xHCbB2/jN3XvTDxa5CRbzagIdZ
7Arf3DtONuWESM6ZnY4+yqmJJACCR6eKegob95HUyCHIMi6dAwjBvEqNm35FHLTuFWAHB6yMUHZT
iM7e67sBVPKTI1ckLFP3TavG3csSNLMc8kOIMOWHke9/T3CBIMfBHLOb4CZyxxwQyMAg7vr/QG84
gSuoHotUtcmpw62LOOmJ7lcEOfGMjq2sfAPTnU11YTp9mHEmZRPgn4O3CQsFs5a3NHR6tu3zlJFZ
cz3N0A1wA5feslSz47Iva+71VOkaGkwUQdNu8cE78bkwZA6fp2SChRrMDJ1N2+pEoISda6tq44fp
Zxu2zY/oL5duNrPhoIwFwNDg7fxscF7x/139acCp9rRJ+nFasx9LLCrPwlTm23yKeDZ6kF7nQZk2
2K0J0vpqO05ACK+D7WCLm+SUbPnTSyK84srkanFhdlsbh0Ajl/gvInI88+2c5fzXrJ0SuXPu9KVZ
gCCJQFGwU9ugMRQCS8k6AZvIt2JtmF4Fig5JKonPkAxrH45vBYFyKWP2ypyaaINtMQNyZUuKt9K1
hE0yzqNrLoAlmhaFU642mLGoSn0lec+tjwVc69SpLadxv8iKxjk/WTddK3DZs2TueWFvNnZsKIPI
kvd1Q7mL5LABz97cTlcA21icYkmunrGxGn+oilhLUWIDyWlOfz5KfUVCTKUyNtrwQ+zECDbxp2hT
VBA+e+NTQD/eOQFRmhBidTSrtAFuGRBVeP5B7ftzP6VQj79yLIUYwuqLcKpWGLCXK+JjA7H4zhNI
fFA+ZgMGfSue+tw2e55MbHfnp9lM6IdFItMECLVjhF9S7HnJn9QbAZPjeggPzNFzV5NRPVuiK+A0
njUsXAXWSEXB5ti4kbBMl+6858HZNxVnYwauH753RA8nz2jbDk0un2ESVqyCkSEPz/B9Yx7a6+UA
JoMxm/MQtFcvMGCGpXLsW2hED2n/KppHViGRO0z55cacQUWh2PYfAXpLHi96WbW4muyA1+LOMVS4
SHxMixJrwvnZb4NzvUxb52ErIiNFtp2vxyXp+0NEcopdApAAWVyN9SsgEH1IiqvZcpirO4sig8By
EnbzMVdZFeqJL9yhuCIWXkTftW2GdgEaU5+5yfJFnLCg8GT/V0TecAraEIsIric5PgKgm6i3pWBh
yfPvcbO080nG43b3EuR/ZPJ19NSJvad28PyGjFjYLw4iCkBV506FVO3JldBecP1NKj6oBM6Nm+dV
QNwU7LNt1719+XFC+0sYtUdS8D/gGJ+kUG91O3z8Iq5zvHdWj//QZvHut+VOtmfyqtHtnA619D5W
yXhhK14F4ceBewUweBHpd6Gxof7ZRnowyibJP5f8OpKxytcU1STE9zuMGlHKDlmSntFrbxaE9zmb
IQZXITtbBpeaXoTIheJGE7M/j3WEndnukvD585byRzPNc5F7JThjqh9Dj9vKJDDLPsFB9Pd1cFAa
TCIMCz3w3sicLeFdIGOcwP8jzqRwaoG3t2IlZzG2pXE4sEtIs/6yBX/VQFB12FJ6zZkN7OOMporv
RIEOaE43ujeLInPqbFpcTA837+8J32m5nuZe8smAxpW6Ez4d82ov/92ch93Z3Um0Hbse+IAk7oru
J7Q0+vKu3ZuNcSA/qYLp8dKYYENMYb6c0SE0GOEzOUtBx+d6/YnHTagowa0H1Q7RDPHS02H5i1ia
BXMjWLNqKpcp4A9EMgQ32JrYRPTnCTY2QnAswl35CwgMU3pcxJY00raTN5/+wry3XdFTs7ZMHGkv
iXXczRZbNdyjQG9MmCrCCwnrtnv76cm388PAyFzCc8BPtUrbBBKrwibuwmKfNSFf83bRxMIw477I
O6u3Y8FyZvlSq/cUGA2rxOrdymuo64pPpcXYvP++yO12waBobeYGfuKRAqEZhE5hjC6rGMmc7bYc
v2C9bz+kBSIYjac2RgxG/kxhkswh2fmW/0QQKuTboBHsvMdox2asL+Sufuu5BXoGPQM6LWSDBc6N
oWDCzM4KT+MHloJyuV0EkD0/yCw/L+g8eyU4hCuo0+P6BwFfqwN+v/yuP/9VEJjwFVhgq+gKcL96
bEFJvOtr99gRoG0gYtvu5lRDZ0q9KvE5gG2ZwbWvBZYufnk+/iy8AONU3Q0nU1oviDHK5bwnvuzU
IFFLupFpszEwnZrYMi0JpWmYApAqd0I6Kvvaa8vmGvJpsopJsJ44ZOexUT8lPfgumdVpW9cKxinv
Wf5EL1vxo9sy+cb1rTB3opvK1p1uiWz569xTICSKOl6hvzuRMVYeRtNGA1lWDn5/SLHBJb2akYaf
ovpQfEbeh+cWmqZMkom3YjNBTksAUZWkGqO57e8kQ8tn9SzRqXeuE709Cxi+gQVbJSXy9rwfcElZ
t8xtogbalfWQ4r7FLxYiy+YYI8vKaGNppFXS7yvG6cGaz9JlWgz24J/Hgak6LgfqF6exfoxq2ewH
1J87oJuHopWnExLzLCx532jUpMR1AInzbQDAZ7WNU7+7dLK2/AfNmcjgvtC9+9U8UOmwygu70XgC
5rgXAjjExBB5o82val7cl5g5cHxMgBNU65kGeE2q81EitT0GaZXSBYcSBTiiyI4eIx6WdR7SZ1uS
K+Qym9hKhQJyoTgcBiqQGzkZHAgkvyVeGe3dk8GUa+J/dj1naU6o11jih3ZiGD1FrsRDqoPuNeSu
fI7ffNdFZVpj18LSwEiByKy83V1T2cM08ZGzJAZEtLOMWXDqklKGUIQuI2il11TP0rfLbt09f6O7
1bssVP/Fu4ZL2LWlYVhzR79j2La2rsVaZUoi9FQtgNV3Iejq/2R1GDMvrfryUOwCjKQuxGPX2Ma3
E6JL9SJx1llzKSXpv359LjLxObX7Tp3O712Ts7H4jXLOs8zpVeH7dGpywHS5/hPJ7O+jxu7jhBUP
l3QsxObXxtaR+w4ygsLcuNldLXAWSNEycZpvy6eCevk46S/jZyCJ4vXIafGKQWCPc9GXB5qoM70Z
WyVal6nT43pm/QdyKfRpB6n4b9FdeL+6jncje0jdoUtl3NcdOKkKW9Ncer5+4Iw1kuvKl6n7GhPM
2RBazf28LYeQ87prCBti2CDBDdc+urB+fwx/WB0MCnZq2uz+THqqddOeZTXet1m9ZU9TUtrlSa8f
cW+KbcAWsnEsPVahB6Ap2t6xTPQa6WvITIOwcjHlaaJffHJ+PGAc+RawCXDjFMftlNS15UnRQAFY
xG4VM9txSulPZkxUomc8Yd0zHb/UF89uQkIxA9XCHZnYQudBEb/EgWuRXTdkj8MG59C/e5LlEAos
Tw1VMyPv5/KrIh1W4axFyiLCWa75iaSLVem8rV8x9Kv9OOnf5UO89UwlxnIxmbP4fQtyplEpx0r3
GTfpRcOebEUnbn203cjb7TskNH+ShBbcCQsSbgM1DnMMcGb7uNDHrdkY46z+rDp7MwyAhj2UwIfm
PxQa/93j1/zFBch6Qznv4Tz1bk51TnVmVXveam8g+qMki9DD94IA6ipe3sMFki+aegS3x0JszZ3+
wV6k8hRNwstSTVovyKknXXeqmwTQIIhX9+79jW2ARIKSp8mqjRy2/gUEZ5KizfQV5PG3LDtm5U7e
zoBp47EIv9rZJYwVVBsuqFUa47qLnHTNxRmky1w+sFtiHV7wD0QNkeh/JwhokShPiSyk7SKeM8co
ysNfoggJbKrDn4WnUavTx2ABzvAGh1TK2cxz9vqe1rm8GuxNflnaonFTydqgSSlLKpeGbl+saAo8
zOovFx+JTNLy1vIBycwSsp9K2wHlNF4gGVZQlKq0DVLOJ3Cz7atKs82zfcPI5EEIA3UDx6HDDQLU
nvEpbU5QDd62hKc6WNtq6Ex/woJSTpuS6EKX4hI+hrc2pWWX8gZ8Hp76+K/1rf1RqJ8gTI8iZKsS
WciKU3lZamgT3HbmBw+Mv5tuf6DF2jsWL5sMx6n2YkrSxIVQYFR4kZ/FmH0CO3u0JjMzqJPYtOLE
oewjYDXNTrrkOu1WyEDbsYvLJkeWedkDBkEqSqTT+HYp1edoZ0A3f4z+txEqt6hTNFeLriBFoPq+
gaT9dZdf7Cwjw0m/qr56OdrH1Y+Vmd0NZo63qmeyVRgady+COwtYM92+UUgv57OMgJ2NX/svt5zC
aYVR9EMFDzM0cyiiG3w0FzmvZV75nKoW8orYUpaDWxYsxTQJ4c/k2qgT62E4heyLbvFbjkPxB81y
/hshOVCchfgFARx+NZZP6x6FariuiJqoLvHXMoXXBiV0PYogFpB9MQrk/dYmyjBsYgNkfQbsxn3e
CtsghmQD2nqzYMOTGvM61d8YrYwR4emfbsjsr6xN52QE4VSMSOfX1mW+MOPAltmzq/GgYq704AEx
ezAqCCYfSrRzm3SwIDVnwNbU1NcKIT3rYbzi8ucP/PiPokYJ6/m/knOnCD3oUIBmous/A31Tc5Wr
giGwTt2Z6PIxTSpnd8Pcp2avIEKnN6wg6fsGV28XXn6qCATsIOsD2S85x3wrK3XkoBu8VsC3eqZ9
pdhXqrSsUbFZbcc5e/iIvyKh7u2d3RtE+mMWPIPg78ZZGc33VV4E3OPUNHpCqCOfeyOrLyQN7HcT
fVeQBSpnZ7vDNKzMbRAq4c24OmOg8yU9RuouTLk2DT4D5RGWnxFmH7MQFmu3y/WsZc6NAp0TCxr6
Cwt6rKTMpHr47KeL9tcsGkqEIf+SZDueTFul42W1OXvhQN0Ju47nNDzFeSonAOjt/f+gcxftrZd4
ZWnk/ddwS21q4Bw53hmF6njcg6wAtkSdgJ0dQt2bSNjdTX2iJ/xJ6nckIM1MxiXb05a4kJxYy9iL
V7CmNOodsbERsh938jQtjCwzgrg+V0xlV1kkaVXHchYk1hXpZ9Bzx4o+VA2xXX3HHUdNtLIa2juf
HyOPci5sZnOXk0T7Dt9t5zxoWkxQjLffVoW5BtfeME3O+hqSTZbHgnKdBCOP+9ts21qSd4HNK428
mu1rtdQ37b2ODbBZJukE3WLVJIHbp4n3N4FH1yTD94CqXeAOxnw/Eghp90X75pRJq15tbaZCaq86
Hlv0fUP/wEhQB2fQSBv9502P1z61GLU+f51T40oBAna9L/wXk9TOQX1mGkFIovPh6gqOOiZty/IC
a7NoYF2abiYYzNTviKtDOq3VNa7A6CYtfod9tiEIJV8y7/VAIZIMyY23Q+m++7qNgJWcIh/SOjaq
i+z+EcBlzZEfCyCofPvZv1T7cBUDUox68yyHV5roMAHimqOIe3wNc6HCGcWE4md+f9Xlhb2qlCh1
PX6LSF4LhCYamv5aDiJ0fEY9n75rdsyuwF3wg6E7B6qYbMfZF4aqbqnDPEkPxR+q+JG9enDIyGmY
Qsj2yRpEo9VioY+bewlbCoDASAyms9E2w26RNC/W+FuVg95/D513bAhBknB0GLiBvJMGHfZHlnyS
Lw71MHmH4SDJOqMu/1dlyYJ4WgpN4hh5hcn3j1mMYt2plLpSzPYk/G2DynmFjlr2vUmBxLPpoo51
6wDoBbnUWkqshfQ/aVRvyDOi3c44OxeePhgrJCC0z4lB8rJG7r4lwmFtJy0gxIckD50vlPPD1mKy
O3dCV0QjI51A+HHL3ncCv9a6TwoutxCv1BkUo3vExTjwFIWbhEfYhi4qVrEb1r228CG2oVi8ZRIp
3BGuhNITTbl3+1ZFCdUa7WomIoMU6Wpgee12Mo+HacDNGfafSjezaHPzl7WJy34lLZGV7T48ReeK
TzSI/pcxh//EQo74ASmKZAHgBqVoYle+iOiM8LJlB08XWylUuNu4vvLfzmE6Xp84mzZ4ttkxw5JR
5d5FE98siD1EEmXtMXsHzOcEkEUvcHuLqA62sk9agt0REiLJq/mU+E7WXQWw9q8oJq5dF2E/Azi5
RyrEH8aKTtNVAEqNTOe91phefaEOODjpVfrEIlo4ZI69kiwrsYfsojKCPAbOImi8rT5BzpUgmjLY
o2ECj7GANLyf6ENgn0jlvW1WUatz2LpZ5HAdATs4VrVhyrftVoW1wBuwEOBpCwKruC5jTaeYinb4
h41Oqw/SzTyQae/TtZByEL/2u8RJ5cRjMbj3Zu/EmWiGcGff2/mP/6v9tFbImL7TC78JEqPxlwHA
+mwIWiQp3GvHHyooDtFp32mXJLl7HACNO9o9W46weRtxv8enjf7lWXw8VjrYe6o1x2HgYZfmOhnT
CbH/emIiXeQG7GkTBsqKbxJTwbpyTAeTm2VTQsmhRK1l8yvW0vfoAvgK1uu15nr6f/AeBVk6B7B2
QK74d76PvLrK6tPnTLPNHIIZAqLMowqecrCp29fdM4tblyWMxm4Nxk4AehIjKkWclQkMgwshhr2E
4noPw5I47xRJq8wy873crg2Of9cA0wkulKEws0Uud+gGUYUzg2ZUG/DSlq84GF8YEGiRAUIM5i30
d6rQKqEvKBvSs27IVVIUXML9qxUScGOhcnq+lnjEtb0TsuLDhtChD8m4yfAN64fxKlsxwhhPXFv3
v9Zi9g8Q9tlKTFAHftKc5maTPO/4bhbFE/ldvNocUaJPogFhbLVzWvoe8Rdb7gu1+qJOxRNKmZn0
b8cxjsEEv44Lg5E5i2oK9eN5JO2lCke0zG4EcsLS1xraBBzefCEPhuyKp0a+8EJry79BGRY19zuy
wUdnmHmyQlNkFjSjyTYrzg+b8yyqFH6MrSqoCwEQyxjL1+Xlb/VUHQtxwwmFEUrXfwgTPCcbsEsg
pHcslVz8l+13BVsv4EKa2YwEub9i38zRoH0iGcF11mRZrXYZIu6zlTcb3TdpdasZBA5ucyoWPthJ
GMHjQlbI9Yq0bD6WD5YfnW0vbtWvr0ecRP6I5PKSvJaX0LzkzFoH8E14CDoZ9ZG4tlVWQCcLlfWJ
v5q3QPgsv6pTn4cARH5sExStMVUDzeGRqc6pp7DXAy5YwIp5j9hYA6djtOr5sTBjV9w+MDRtQBLL
NL66hStkV+RDWSRW/mtvnj6blq4dADq8pelDChwifPm7YEKsbYsOT28f6fsuZBSzzSiwW76Gpw2r
jvtZkfrYy9cmnulLR5AEkAu0ASG0zrkciuF/M7cU7gXcuK6iJG8I4SW9NNNK0GLWMN5jAkC4V8wN
OJ+R+DFkev/YkMlB9t0Re0D+50dY3EPLnNuNB83U20ilfy8x+RFgWGXHnPda3PiScPPc02MVRgQh
CkwjpHJsCI9yHhCBU02PA1ZG/kyAV2iHVs5xf8qQVDudb/QKdoFbnolkSuoA6XaFSA0sZWM3EC94
4XUSL5Bqq1BiICn+cRz0DpnubuzEJOKyWvQjbXUetAhsppG87+FZ+o6i8//7qY9U8/EDc0G1QL3T
aohJYux3l4ufHklE9mSxE/oYdd4mEFLNIHVx/tRmqWDxEmzBNhngiGq0mIJ4emRmPm2NJIr5e+iX
4lDxGz+gqo0qCENR5TygMG+dYCyS9X7jtQbxQj7UOUXuuU+HMSv6QWxp/tKCze9X7ih7tlTMLXio
aGikc6tZmtHUqoZfLNnA/n0OnlPk67ddL4rqm9rA2x2MW91CJnktVHqHhntb77lZKHl7SiG2EWQU
I1qgIi5ubyBQZx7+ErH4mdsaKVld099DKjNrB0xNrFMNBvTAzPSPUUqIrhp3Pr6q8gb/SqB3jLm2
qhcnhj9llnCnsm1X4iPpq7tbfWS9nVcToaCrJHBk0EQGnj6ZoRfjD937ILIZdmPZKME0j6sdqW6E
UZjqz4KZJDQXfCQMaW9Klt4CCwwtE0ee9wHNI7JqAm0Qh7kWDripdJtiLebI9GEYp7HMijMgiLI/
U5snfyyDtuDIJxYRdrWi9lJPKg4QcsmQapX5GSnf4vSAo3fW0pN1yhPuISUxXKvrgsTpTHaj0KWI
p/Gebj6lIQvxsXdketM+LFhoNxtUbuZfmir5fTmXa0hSksaEq/iFQXAAdrSTtM2oPEy3GvC0qDIV
UyO7fjlGXciI5KZ6ulhYWzEIogQEpGaQqgqLJrmm0t8Jp+n/Tx0KksWKAxuoc3Mrcc/VEF5P6RJa
WbfCnBOZerm0LxnO338z0D3+Hxn10KIpjrF2D/xbhKLVTtFEuA/Oo7ltWzbi7bPWZ2M/HmiqGyiE
rPspKnKCsE0dCE3KVuZ/xTzoedjDyjcMbkl2KWGive9NxfUAQp7I3aQVVP12olVHYhnLSUHAE5t5
xKyajSjl4ZxvXi0RW3gTEAZYo5lZ5YXICfXY6QgvSJ28kUeF/2FECC20pGI8tNogTxkJfseK21Sk
cL1EVmo0LJuEB7XAdENBMAu+NKahkF1nYI7rH7MQsCC073pOia8a0pjeCFUjh5jgcHm3FJfReIMC
jMeo8Rz7g5ZtFy/U2km90Raw7TWEzm4C0FGog02t8adik71wWZdKiP/FLfwu7YuXACTPWTR2uPfv
BaPxqOHTd7EhMOwIJ0c8XNBxUfM/7Zo3aueThqI3XmT2oXTURBXJ1eHlrNjN07p3vVumwSMK1dcY
qxoW1GXEXgaqYrfdWZTPfcJAUwkP9WdZ2kO8tYgA9nebwSBAVTGGYmlM+dKIGLA0dpPw6xTSpoom
yq5bdur1DYNfknKwTlM8yTqEsvQOYIpoP00oiTd8u3eZGXd6cLOyrpnMydQ6Ce9cjVtifRpzNJyc
XpdgCyUzzT7RBXQOuHsfXo0jg2+rte+ECye7VpeluKpqQkvJ6N6w6NtY8DvwxjwbJqihTHcpclCB
jhrS51GrrGPuOnoeM+pYxB4bCNGLOPJYB8YDOjSRqK+oY4eVUYroSLqWFALDUF9hJHuL21JHepy2
qoxMU84Im/cWQwR0nf/qVRvdGCaRIeC1+tHeVeXT1rUpGxOIvqcq1v1PaW7mZ7NiKc6MU0mZJD1Y
Eg+1qkTwwK/txklREa1RDbfQL/4R2CMTYt5612wVgoEC8pZCvFxzYk/XKsKGpInAKg3wVPKDSZPM
xB5fMvGSoagikZQX9LIEysCAf9HojtLIi9NfDPw4OJH43JsqUBQmS0gY6vJEzC9yjxRiHswSPlGa
RleMl/Kt11P6AC5qoxp9LavUHjhqujZL4q0gdzXPydlhkX5VK0PK4PXGJCfekwgFKMXQEWalJVIu
tVBPOnxlVmP2akJxkNE9oH0KT15WZqo2onurYbnT0sbwRcNj3K08DFSE81Hmq21ZSP5gVn0M11Lf
47dW+dTzOoc5yv8qaZK4bQulQ5ZG4RUCWt+RcBbWMi2n+pRa749nyR6qoOqT6+fYL64HTZF6Auu/
WX+3g/q5vR8n3M+Gye3QC+W4RYrd9l0ifg2lMPuy+rnjOdh8l+tt6GfXL2XXZg4v3yvdq4nLb6LY
q5SRvyUBvXbDAjJhX0oOL9KZ4/lFToJ/9mXWK/70FK48UzJriePlqUxnc0R/4Mmmalym13Oe0C6/
o4x0QqBGQwRNvOggpz0NLqZnITnu4ki+TjwRzmh5HULdaHpeZ320E0N1lrFbGndI5B1OEtJqaRTp
3LZii5LIsNpZUqAcNdxbTh/QDTLJ/+jjhn3CIOM5kPS+PEUPTqipXqk2s3S9LfviifbbVcA1qwWn
qcYGXinI/az9jtY+2D9xNFlwz29v2UzrkqCQa5sTb58FLHzD6rRdKRXMueSkxgSyyJctoa+hzQqk
yjZQBmiznChDiRAz7o2lRgxRzJrxiChaKLcc92tMJyod7jZohjtkcpr3R8ZYvezzlx82eZ35aLns
ZkZp0Z0Jar7Nhcq3kxmot0Khcm9wufn4oD1SaDLDqVAmsoPs5wggxMma+/FEAv1rrolr7G71g8H0
HoRR7Q74ZdXWReXWjoYeFsDgQtTY9Is1aXJrJyhstKcDhKAETV56WQtI3XazDQE2Euic6wnu3oyA
0nBFlm9t8JFETyg0vGfDuKM3hDePorvqbzq2tVooygIUJ/T76hy6hKT/WbLqbq1GHSyuXq0aqzUv
d0zJuWsrY7SzdCI+fW3NWaurJVKhSh1dABRz2U2yizMauVoqUW0Mw63kiY2QGRZlrO2Gv0vt2pHb
aCBpL5bjtvyHu4n29Qb2qqfsHlJb8dHngmDCcmW4A+lKdqt6dbtxKO31T4THrDoaSO6i7ZAUxjlw
PuMenEY8kVMVWcoXcPTkbaBaQSUBTmPChAbAG5NH/9jWtDJySDPk3IQeO6d5N1xvvPyus3E2ntOb
bN/abeyJk3suPXomHgCl38NvCHRNE0uVcDQSnmp/xV7JVoZINowj9Yq9lOEQmSqSk/O/QJdfzBVJ
/ZvydnldxNwnbE2GHxFCWss1FiBFj38fY4FNpIK8h09KETPTVq259M1JgA60gQ3+yMF3OmQBz1Ee
M+kskbY8aBl84I7h6KA6CczM69oS4xnbH9o7RxH2LgY3HKrPfb1uT6Uj+0uQh3t8zizJNWr6FVgB
v4NXgK+FcAs9ME7mw9ZPtYSVOIZrnd6GTOeXCV/MmzU3FM2vrky8Jxi/ya1T+rosz1np6D0G8via
c4MyA2U5xS2p9ffxBhocanY+gmvQlxgnPMdGTCSMeG/Tp77SlMFJef95tZJvROKlbWp8w2N101ZY
QmKlFHR6WdiPseThXXJgX7nenYa4Aigl6r09ItslOZ4ZYvD5NXqy7sHQV20JIRiqBCFNRputkzbP
vPigqXFC1k9cslbNLVK0YmxOxlu9m1kLiyVLj1SNh3XMmsoxkOmaGUTq4By0V/ySUyweydRnZZai
g7O0doXOjECOj/Fd1rHhlVvyWcyyQSGAoGIIpNh9TCM+Z2nzxKz8b2/9jwcQw1jAYtxuUU46qAJc
nhvky5jBYtQllubpTbMot0y8tQ49Eu+OYpZoCi+mnrckzZGSTYpjHSYZ8oU3uzsAGDi+dNMlByoG
FlinSkagPL+daRqJNW7hZF3Ddl4dT1G6m8S8N5FSGSB0Yw5l0E4G1rk2bTJxfVGunBYeYKvL9EUo
Rh/qwAHDN+pG8QZDhe4TXXtHD3yjsUpsKjKUsW8wyLNwH2O+BCiAElLwvN4k0sp17hzzmFuvp2Qm
aDeL9+gsrNUFbky4K7rUjgi75w1ybMWbA6lrOfMXoa5BywpP0Jh1/gv1aqXjK+EvYhC8j5d053Bf
FTtizSV0/Bcqakaesn2AoHFzQTMwGlfzZjmxWWxbCX5j1k+EJSvKxDOoN2jlJmHTD4+Eg8IoV4G1
56rZFSPiFt3BCIJwGDd3tJD81rZB3J4pjkJSiSc+JeaSENe/YsUNraiTzxx0Fo9I0i1VofklVUAg
a90SeRXkioQE43K5dI+4MUGP7+gRX/mM88zAvEJAc5s+sDlNgkex0SomXDB92CXwuF4aAdM5piz2
pb5En9RfYw2f1hSIOzifEU/87UxtvV/msZKpoIgHM7x1h1bWjPlLBd5PPp7n0BOoLNMlG4Mz4k3G
3Lr5+XFtQAp+umHUmJMGcTcncTinRtPw2egGe+zOsYqYE02nkgi/XG1buk2QWbf9Zdpr6UecIuVh
7w3SrZBriZFhnJ7jy42n5wde023BgdEZFTAgUzMrIi0PmJ0r1MUDR1VgO8/UUcEp3RiQ15E5HEWx
YJVYLAt+DVlgNKEVXbK89VJFm6q7Aevg783KkmWQCVcbOKzV9JaPR1jfq+nlLdBh/mc0p3jXYdZe
ppiy3ILbLZakiIDnJ6b1c3SIFQovoNzznr2wPp5FUKHqJZJDlk0V0rfsyi4OrTzCIu5QHZHS19kB
6YQeIr4BaKzbFUqwOpWZ/6YbiYZoDqbQcbg9PkWy3Dz363p+OZqkuGYfPmJPkQbkb/1aXhDkInhz
7d2c/bP/WBzcx9JammC7UMvWhCTAtLvzrXQ5vMwpEHW7xQoqIXV1g6pRmomMO8cXP1+Aw4irT5N6
bLx3PVVVKapsbQXXXpksVhrF9MzBx30NupdMS9cfzGfFgc7loHwxOQ7T9hKeRs8KfFq4CTAnL+je
0FPUPrtyBlcu2oJD3xBV4uSUdeQaubsqFZdph/aYQAVzoVk+ctHzpJWnTi9KwIkPg3VY9nPtILx6
2tfnRKEcrbeva60Tb0B3Z918GAzUnKAeadVzJFUPfBxmBvpyFpML7dk2sNX32P4YHiCoI+/U2Txl
VLm2N+HWUUrtuz98qYdRh2QrT4DSAAvYayJEAIqjdlXa5SlAckfm7Y5kl8/yoZs3pqdq1TndO2ll
KqqAPK0wsmZB8ePoPrBKwGMxVerCtgnUnfzoR3hNFO4Ru9SzpCpPCXQTdiqv9ceRUESCifKZ36Ml
rdJiJj7MhGdFTsKmPYyhhvupPAA/Rz80BIwlgnf9WHtD71T759hwuzW9tVVNWtUsW6GzU7ACf5Fi
ltPYAmiW6KTKXqlHdNl99T2dAoorpIiERprUY0LUGZ1Zrs/PpRfcXoyQ7NH+H+crVwQJrP6sP/4S
cAjLKdDjPqaaDdvNYJyD395Dc4i/x3L0LtSNvh4IrdjcrwHiOE01ilwtMu1gHKcNSRbwlO4ldx3B
kanunRzxa5Mmf9eqGsLBRkB0yy9yCCce9KCBY3XwAjpzynV0MU73tqumaPS5XPlUKRac4JnhtR6U
rn9X9AygmZJ7KYbmof964i1pBMeZj4k9GjpvE4/iBqwp0GJ49treq7gYMeaRj++hD8P+LkAEQsbJ
Kp0FkEXzcNzseredCw0t+klP2a6EgSbCRG/FaMCG8g4WyYO0mzkVxL3PDri4HzmGgdLbIAxGX4dl
NlKS4dEEbNaitN1rLd+ehp+tvDkoOee2wxYxPFqhy9WvLuD7bvkU2Y8kvLF89gsytWMHwMNOwm6m
J5kYwQG8P1bceEAKKZ5QinR+m6NWbWw2yHywd5PS1hlhMh0rCKmqb4KqMGGMyWoudD7npycBjyab
5d25sJ58K2/cMsD07APijKa8tnhLMi7KJJz9BHfwV7hKr8c6abEaQmVcMvof42uMqp0StfYkbUub
Qfg1A8G3u5nY970b6h4T/g6VDUPmSYvnYfSiIpBvkqwIGStkkSMhPD/MF7UU6yK+QhBXrLxhJJqh
P6p9bqetAZjI30/GhkOZANx1I4qX14zmOX5NX1+20N/xIxd1kex8SgidLp5XZNdna0QZeiH1Yonh
rb28SMicjrpOruKzLq4Tr0QWXUfs8qAbyRIJKIj+mnJus5kDAdMoKCabIw+b9MUGeGYdhj5pyGjY
whp+oHgJ1F5sTK3RmujS3oBqvHXWntJDx1gxn+aRgAX7gzEoa0C4fmCFphJZFJ2/y8xQLQrWpSWT
n8Z7xbepm4aaE3SMpeLhPsYcyDmL/b5ntBf2r7GFv1gGNY8RIrd5mSlE0ELl1K2uTI+qqPfwLerG
EoC67VT3MIveagRKI+yod6FPsr+i2F4ZXMFAXIh78KZZW2Bjam8Zyboj5iqMuA3oUfRc5myI39wJ
/rQYZscZb8NlbgtEk/4jSQuBE7oENRi4F1lfhbV3MoK9GtoS0p9EhYbftj78D8YXKA8mdl8bLJFM
jemM7guu0gG7OKlRocwvRd+ZVDNHP3jsIllJzgeMzjsd89/E6f9UmLwWWr8apRiHtYDb1bl5tQTL
/v3YkNTZeinkZwNI5wy3Vt3KV3EuqROVGDypDS0iGpzXhU/CulK/F5Awa+cFhqcp8moOpkqWs7Xg
rkqUFawh4ZDZG7LH+t+mY7wgJ5Smq7V8zY7yqynG4oRYnJIMlYuwS7L88dIBgf3n1srogZVoMY7u
DFWc4MKzI4UtZOuX29C7X1I10crzHAPYhwongXAy1Gs5Jkg+80jDdr4oE/MMLHBCBn2tjdxuAyCb
VCKOfBVX8pXv0yjthB83lk7CoxePLpflDWxN0/mdRXyObrz+77LNuJ4ViSc06SxsWJZx7axJ7rpb
th5GlC67MFfaEvlHhv3hKI9tjpQ6tonR//gQqT46otaE8tf+EHXOg4XOnC4B94v7xWmiBz3lfb5E
MpKiOKtHUZ+GA9OyGZgnVWdR21iYsH2k/BGtNTI1/caZ6KZebeJUe/6CKa0K+iJmzX3F0ka/GMSe
WjA9Tpyw7qhOEB85m2nJxqY0SSBhIk5w4wa/4Nb0iAQQNmbEftoCKzTFWF7e+mdEt5HTgJDZKvtB
NsTrrFY3S0NcquE744p1XmhuuABtZ4HukDNOQMJJBKZn41hvc5NGTNUdDwpZGbNkqwUltfS1Igtr
kZ8MOlIzpO0LKczR1Zq6QqImpfOwA9GgqIIEYGFsfnevR9SQ++4c5x4zoh8zmlLrNUulNGZpkj3t
wKmFtveXZpYsMXhd8FLdJypPTWxGxVn02W14exlg2vew12DEq4RMZDppgXukkSXycWC16N0glwYA
hiRF7zaWfi3N3X07WjmTNaK8eX2t4Q9V4+YPJh7y46aI032xGI6AZJMPXifH5ibI4b0+M7EvIoNg
M+MqIvYL6yeViwAOtpJ46C15bIk1S5QIjFqLoR7sGyAuNC0f8CtziniXr8dtoOESu5XprL0R8mf1
1F5W+4jdcm/LAtWlitTDX7srYLnSUpUoA3S/ZWxe27GHVRxN3f8qL55L4ylrxpkQfLrcHyNLjMaZ
yA8qa+AgCn2OLYkmqyNn0KB55KbGjWsCSDPhA7y/UyuC2i8auHoQHlrUGa3jXySVnwt5WyGohxGm
YkaD22QfywzsQ4XzeCQqPwJg8pf4BrtAK3qkYo0205msjzmK80dRAKN6r0Pe34j51ZgVBBPZIkze
WBFhXQ7AfiCi9ZQllB6frAyhP2Uk2nJLaTLUcSa36fs/FkSufWCjdN7fNiPhidWufN64hQ2d3wfZ
WBLOTctQm/9mS71/E4YFFx1MshT0DvkgTxedyvBpWKiXSC2sV6i/hz6CTEg6TiwX6phCeG9yv3KG
cpOC8QG+MKQbpff607dmdseh0d/BEjUD2/fgmMO1YOkx3yDCnw3RuQYx5xSjKD+l7QCnV3DoD/bl
AUzaXXFssJKdPFstkHbmX/RokeTEJ/lABkjbQ0Iy9Xu/zqJp+xQLCj4Qi8SWNAyFxXNBjZB6fJD/
RboB8uDX/pDr1uhaOUkAyBW4kRR8KR3+5PHhZ/9O+aPMK/Cv5eAx3pGKlvuijWTDg8o90RTGEMUS
RCa6Ewf1eIK8gDJYsCIXbRtYI9zvdjh6bIg3AU/SKfJ7nstZobs6cgcJ0bSdrulowi5NdOozbsl8
Cswzxe6Wpbi8EeeIYXGcnC/lLas3VIoMjYQbsV6VZIiHlM64zzWvCEUz50JGkxgnqS4OKz75UZFe
wBof0Joh+nu2niIu4Buphai1tniffOksSvOuouvUlNzLJbqiaO2N1hCGppL+wPXdAZo7Su7wVZjS
LeMuFHwFLilGYAPzpleDgD+C5aw8TbFW0Fh4sAmbp8pCW4EKind6bm4GSnHU8HUjwGf0hnd5xkBH
i2qYYPkDMHd4httQDSJwjFJDeYtfNslbsToWke/7dIU4qLe7xzlFvZ8Zll8rb/V7J92dAZnEgwfu
feDrLddymhbm8xJ+ZusPYS4jrL07WUJSRifASmzXHge3/5XkJmSMOZMryMo46lCQbv5OtmtHTlLS
5Hw+zR+6Jl9hxdaRGwbgMZI8w13/4wlmNs8HCaM+7wgozBgfq9QpDGEhRMCPz5IZCPAQAlBW3e/8
fHIzt0VVoJmUfEVZJYbr7SJTFETo0Lh3w9zaushMwDCaRcIskZikTvLyBC6WtU8mK12AUGbO3l87
l/U5HCaKuzM7fisGZl/DLvA1RTQt6nBeAS+ZuMGSamkbE7WthGqXYG64I1wT3E/RouR5AvxQgLjZ
R8dQdsXyF0phxoYHGvTi4T29KIJ5WfAdelhmk1o/UXrkqt+zugnlgIoan78Rj9zHYWj9k3fih8A8
C0wgOtUdTTjh3Gc75BfUMFqzVD3nSv3EpIshUC1ZeOB2ANq/McV0hvekSaZ1xLjwjC9RrVikZe5l
mX2yWyRCaXNYgbHHWbLBj/Webo1rjQHgw8Xv9yqCeivr8dopLD8xz9bnfmfQQpmseW5wbH33hS6w
KkvaugZSOTPvrSSfKWv8Ecc3HGFb3WtM7sRM5E/goJPYi8e+dQO78gkDEOpCVNYSyz2Ld6F02zCE
wDAq2ffi5p21qGZz9MOWXyc6iJnFHBs/bhnsesq3qqhNAySYxgO2B/cTlEzHJPMRxE76wH2FMW9F
bsh5zJyFFs9VkoNtGo9eia2r7ytmqPhVrMpYYMg761FSzYlzLzxgHn1B8EhqqwYY1oYg99flKZ5s
7vDUBPzGBOdzDbvjCp+SYnzxay0qh1zV5qTzRNIaPClwZ5Nzxn0yKohToW583Rh0A6PTmR7E1ZS2
rbFasOODvSFDeg1h1OavHZIzM4HoRo6rL9xh9j8rFSC89hduzQwKr/0VihqjERF48SgkXW1UAOg8
ZsjFBr8AFE9YNmfmuWt8weVBGiZQlq2NSQpvs1QNajUB23H3OFmhwTG3XImGh8HHUNqthCtGTKpt
06wEgnzJT5xjX2TonXM3BG3XDFf1mH2itrXexSY0E/YIkI521+3gd+3Ky0uqSdp6/JUam0VnuTwO
xmdHJ643wwMV43ByK0nz9h9EUv6y+N0LV7NXz4yAbyF7FfOvIBLhwqF/lJ1cErH6JHUK6M+mBD8D
MP0IA2vFc9gjkM/97QZBo2j1NAKrm2+oz/WcHXqlFCQtxdhBeUCAW620nbNDu87/CZ+bc9Ck4TuZ
v0hcD04eH/UffOknflIaL4SL3sTZMw0Czaztab2PUg9Tc9dYq25t16stlpsqmoXPnDw4eOpYky3P
frb+TZyFnKO+VVTtZ1FQWQTorya80Ws4ASiktNrklU0SV2j2kFlToaXuoqp+u/+RQfRXQ+hEh8Wf
3zRTPjQRidFSqYUuBWXCd7UetTms6lK4nejqmpAQg8xOIWYgDDwY4wea9tC3QvBJJh89L6uQL1yN
jCWzvMJbKbbP5iNFt5l2b0/2FENuFo3l4qmJ6G780qMQ1yxED+KnCRhvdxQaDQBxV0HQZexxrC5d
bZ2o/BVMCC5W01tsp6SNxU9Xp8JfttWJyatMFMt4nYy3BcPdDYJx2CbhfFB1UwCHKrfb0N7sH43z
N6/UIBbBR3SF9AZHGU27p/gQqmzYdW3XGL2VtBuH2JSBnyr0Q9yJutv7lqg84gXL4gLOLZcj9b6a
NCzPTtZtYkvSVuNZwt/f4mAezVXAJt29wxr56EaIKgxnTPaRBRBjT03k7jvpQjpY5qlGgt3Td8s8
Q2TdpeLpaqktQDcO/jvMDqtoXXUKMW81Q6FQ9VfpjGsu3Q9R/3hvJQyeGUGLUa1LeAhCVO2gqQaz
tc86fEzsfrQvtWpDNiulwqaS/3/3eOAwksDfrTRkv+CqeS3ML2Rg5OlaS8xWWvx607rVmEpTQitB
oHIROP+wCSzf12ZUdEn9YLleQOwJW9jttVJqpoASK7BZuI3QS3/hy7agl+0Yv3rjvfY3dfBS/er6
N8e2lrP+TMDg1v/aUZgxbzt5PFW5hYMhArlCMksPFmQB2/3ryApcc1iK7kND0LrtgkNayyKPcaqy
45BRQOxDgliLBCw55CudV+H4xX9REjs1YX2JVIDbJauZSHDY9OdUVT+wxlll36qhSFXLc79ga98S
UlykeeAvgmkfm1gTsshYP0JHjTNvSkhi1Z28l4XiIQnWFceIQvIDRA4wl/9W16MMR9ik9Hej7lKz
gD8novRrshJAxV24Qi3gYtFFMPpikXClgVTNapTmphWxgS1fU4XH74S3n0Zv6xMpK2b9oDWnA8+C
eNgebFXbnUNr71SmkmGAZwE0jV8s+Oa1F4csz80F7YIDWVbbPwgNEPeKDT2sOb8jcGi+fqek/WQn
FKIdzTwn5IfnaMWKg54ziCTSm6s5R+GbaZHSX9KKF59WygB5jTFKnIf9nCRFpRkMUXiRzPerIsIq
66NIWTs6FMkT1QvowtTdoNuQZBTpoTtr6S3dNhGQX0Ct5nppBjcRBhvA4IaVseV8qanRbcumH5dg
0kG9ARbNugOnVh6b22/AtTcOj+G/vduc1ZNS9eiNnrfuhq5WqqG/jD2MqAV5gJcYn/MnhR/Ilp4S
H5T6ltqcO1Rc5kOY7X+yINsI3+zMJ6v3QQ/yKyiuldJdVB5tAtAdISH3pKsyYdGzpbiZpQnUGW9P
kKGagoEXVvCigcBjelGPHfdpmdsRQdYyNRDBdbhq0eeUy/aPaBpLVAAmBmWqWexk0MhBNekUt1AZ
4NJVi15+KRHXB4L79IrUjPIpxGWAU6OaPJqBoMcNeTvE1Y/JN/rrb3BwFI+GOuw7It/2nLI2N/bG
nVXTxsMS1JIpcYCd4sY93aGVxOo1zi0jlfh36hqL/9SAvRE+aOgRzPHNsWuRNIf9gVfTreKc9+Zx
l3Ywj1LxEXR+GvDn/u0ufZNj4Q/Y8heQpxb8IGPzWbvXdr4YeOqmNjtrlcu38SUBffH5+NfVkqOl
GSfk+meHtGne28jSfOptQtfSzBPE6sKconVdDM8OLNEy3RhAWYsoqZiVKdDyaB3Oc5BnZWrKk6bF
eqjCTu77QgWfDxtZMY6hqJI8TxTZExzBNeyXo3o7l1RRYZtIWUsI60R7NmW6toCvssTm1CC/84l8
NBZkke62LxFOAaha3/e8uCo1YJfFb+Z4ENqcv+o7VlBCW/B0reevGTDnJZgvFCa+NrlYAVtV/67K
5vkPrJ2d2oszafZnOvVMkOQfwmFgJKygCTzZ15kFOEMcI4QcvCoFu8O2vBbpeTa1vdazJ9SYBQrT
qsj4gqlTpruouVFVfr76p51HyxJV1glJsvEPdKWyY4Yw3EFTZwFhfIl0djGF8wOGTfe/r8qXQVWT
VdoW8MMOrHolm8bOTs/qouEjIB+sDPeiAvKMOqrQixi1QMWLTuDLh+3I8AWzBKcs9gLQLJmawfMK
0sIO68mBkWgJTLKk/CgsBA4jjfpopKkA879PH9NT/kG9KYqYQZZkotGZc585tX7lmJRWuOMLJF+2
iika2J1YGkZSIszGjqXNz7x/qt0Sk0BJ/AuyPWUOsMAl868GqAyRCLAFf2zbFF5XekLVSBwmTQXj
Tsc7JXvrvtgG7VDLi8Kx2w0P7RSpBbtQVDSjDls96+tZYmX2rvjU+OpFSWyPGlUrp/XXb2gDlawu
zrCLZgalgcWlBJHQvrnvIR34K7mRyIEn5SJhjbv57oXBXhDyNmRaifaMAjhF+lQ8WOqqp68Ye9Zo
Yd7l6MaLW+6qjX6BiGojavSja/gIgrWuXrTNwaIs0PJwRptMiOZJEdWvYeLTO35jY7F8H6Q1thKk
45/lS9vGr1hfhudJRxuUyQiP7MLn8RIxdj29dm+IkFH/r4+5RtSttwv2Q1tGmjwwqyKPd6VIxXkt
DJVKtRmvGvltseJq8VquSifzzd4teZgEIACtk2mvRGVjWza9kCf2CPPAr4irH7ApnLF12gao3lVS
g2VgrFCz9prSRGT3O0Fn/c8CKEnuFJCKLbJ2i02Orf1qs6ctS1x/K7+IumGusL8uL4J2EGKoFXFv
H/aVe56ko2C8OSKV+alwiFgksIxEZGqH0ULCwb0UIug3XMULWQrZWxtaD7TGNG5iTsL2wbgGza6C
AaICMhVbRjo3mlBNJhfckbJlC8Zwbd+O2l47WXwRMfgPO+PdilMpbphkotlCzmaZ+zClHfDQ3Cnw
aLUL0EcxArD6jDikTBc3/LylRzimQKd6j0cr+YNVb42P/9iDcYV+tUamcTxnaVa5D6RBZUBQcF0D
fH1UkImYMy5Yv5FaAiYKrstepseO5B6krhCzDxK5YyRqhDBNnAyJitZgak4RguGuVliznwPuWhu4
Q+T2BXk7NC+1pRVrd5FLBp7h2vX2sVinofxpkT1bXu5SRjse+xyS4EB/nbSMbBdhqLzV1d7Endjv
plsnjiC29Vmx8D0VS3p/Sp1s9PK2saLM6b+SnAiB7xWRCgCJiGNXvRY9yAiwHl0Pv23n0XFVySko
HAd3BP0e/yPJtEy5ZtVYwzZ1U7sgytYlertr+l14OtKyGj6BuOtv1enfwTBV+UIyz3Ar4qHkov5y
Y8zR9fjUmBb9gbKxVPRWgQzPzp7i80U+4yzqAsPUnLBZZD+1Xl+Hnds4NBJCleTxMWDxx6+9eaM0
EgA+SGfIEUfcVCxSoIlJomUmieCPoig8RRB4W4wdZKzCySIRJP/mxad5AtvnpIHhQqkWBXD2KjdJ
4p4BPnYBISU1iNM1Cq7QRMyrp6OsBQ6kmD1XL6VmWPuPmL4XY2hfSQTpVWuKdMG9PkUx3gomj19i
/5zWOYBzTUTDuvir6seKJaDRkx8sA/Fja/nddhRlNo7oQt7gAG1AW5px6ciT38lXfIc1KOmS6aG1
X4gScH/T2Um7ccNdSeIjchdW95QfjuBEO0lrNsoXweHTSvPBCP3hdsqfWbJ9dJf3K9J9iupqd1CG
J8EDUtWBrhXtN6ST88hNav6NorA54uha/voqVAttvL9lAosRzhtdnVX5NpZbiS1i1NZal/Hll5Nn
Iqp0/l0HzDki2kRXfulNpvmO2gCTrjSukDI1YAHhcIKDAGL8Ayc24KFcC+T8KAM5altZfKQoySYC
4EbdQ/KHZbIzR2oB8Nqz4VvHDQbUaxK53MXSSWgp28gofaxw09ishA8WvOdBMmO893FnIWbs6zAw
MOmz0sqhY4SS/91z1BwChExzszipo/yVrQ7rGWF+XvSnVhPPGfLNx8QLscj8LcNOlt5tWfqCwZxx
40jfJXEu0Tl/3Mb/TGyLGilvdGOepQg4LwBg51bm7LiRdmka6ADvj8ZSjJRcKAmVJPbGi1/kIb0q
lyJVWQmh91aaRumjDYO6FowQW5M+nbLxDkvN074AkXTeZs9MfQajetOHsjbF1HKMM+j1nxyiQGnq
cYKZRlUibUhy33Ex8U3wMSf19IoWfv5HwWGJxQGUEOtFPJUxZMejLh+da1EqlNwm/jHfgb9d9+I1
Ii6VYGPAwkOazS7M38BY+XSU0riqH5aT/WpvD4UV/oSTw40Mlu/c+s3dlcEEZq816ZEq7YYDaRfS
BSXJcB8QB01L00Ayzdcoe4X3meanKrYQv11CFxguwJynhRkJam/z2AMc50kB0DRB4J1nXP2pIesD
JYPSYKexOV2dkqLWckJalxidXx7IwkSw71yNASFELNCCoJXprADUOM/mHLFY9/Jy+zzkMyHS1aVA
PB6y8lP/B72+UQ5fEqblTdXCMGyIMycv2/aa7+0XiFQsqjZxaPL87TNV/HcqogtLHyYf0AOdB/lF
S473NL39/c4TptcdFGuURnqXN3luP4tx3581jdmrpo68A0OOlqPbjRniatsg9UCXr3NSpDWZL0d7
eO4A2WDfqfb34m2t7TsV17QnHgImSy8S+/MYuWMTDx1wXFM1Dt7pgR+DS8XAE35O7hVlDlkcm8VA
ILy45qvjEs0O7KgWUjerDcQQRoFAd4VoYlBeEtlRFbzCKZgU26A1YUUqd7oN7uVjd8Rw8vb6xW9s
/gzlBmX3JABNe4gwHG6rraTlldCS6s6MmzyaNnCwFafxMVFxs0sObzstyaB02sB5d7uC9mb6p5Fh
YJAwnwTVuldgipJ1+FALIujqEORhhw6BJS9jfipxHGvUKYttt1PyuIvCpdo5MLRcluNAbPBf2X/l
a4dao/v+Qi2P+f6N5FldVwVawAUA9AhF/6b1sFp/shrtaPDAWMd516bT323G6jdUKpVJSg/+kbrG
XsQki61LHYxXPjsJlZKVt/1qtzmdcev57zGCgebk69IRP9h+87V6vLYJLpqQK3jCU8gTVXSbyWkb
iOcq4R1g95Go1zGGVb6Hn8UTpLwuSUiZ6Pw5+btxibIe3fayZrxgGEc2COFrtznH2aICjshU3kx3
SIZQ3QWUfgDupklknEqyTTzmOyiK3REkDRYMhmgNYjX6GJu85li4Pmr0Rsz0K0Zao3ZrMhC5VaM9
qY4+zfvk5oCWumoWQw42fOv+wSFadYXcLud3jfZ5A9Mw0i4rNHTTORHT++Bi8GdzKYqZdFoR2HUB
CfrPWWsSG3B9c9L4dfbiJIZ/vRZLbEE/y4fBVjWhAy+ZLRwme3jCtD+wwV9hwBQuc7lv6KbGlPkE
6R9Q1tJrZfirtStaJ8r7EOQeWa88+WGHWyonNSAWlVX4R0jbRDATT0AsVhTYgFESZihSWj7qB574
aUM3EWQeP6xZSZETXerBP/xAfZ4DLLqmKKl2YC1NA4WW8G7a09LRQ0UlFJV9GYY42wcE0XoE7DFX
ACf+nF4Zr69rZPNMCxi7s6/tbvQFgMYz+7YMe/0wfvXO2ehGLf3/aa70EPhUULkrFFslIVmJYXDk
Ud4lzP3dnI16Y+iZlysv2l3/jrOy8+S4X5ykPS/1YRexLnPtNEoBMQ3nZRm8amhzoJmlysnPy7CW
IKM50HIQp+mRiJlDG3lBJXxAnusu4Zc2Tv3wQO26Kj53xAIhxA9V3I252FmbVHs5l4h94mc2Ojdt
iSUIQAJfiQAiAoFNyCEO+ripfbIEwJHme6Yc2B9DcCDBb/8uJAccMcc30FZP5tnN6SqZbr0acPhF
Doe0zMS+pQyJ2R6SI5C/oaVQJEVK/zUhkZAINX1WnnFr468CgyCiLyXyCWhkT+gKxNlL/vsXHAea
IblBfbFkwq4ls5mgYiIHLkvUAa73fzoI8YeQCw+G+ULNgFZ9Zl16ToPGgp+R8EKMGk5JEIUbGMdT
O6R3jnppbFy1DpsJUnUXdzsiF/YBWW0gne4zs4UKt6eqg2XoZhuK76Jr1YukshVuAhDb/eAjtMMe
fX91KLibKbA+WrKNAr7y0wnjOfs3Hm1SWWAy3tsnDYWnsnePl50042R7Y1oM75yaWJQm4m23TkRj
MRNr6vK1SEPrk3l4ETiPMLK0wUEmOeWV5zMCCG1mLl3NqHtDJif3SFe4UsyuCZC4YpLgWKwnrByf
AzHsGmn7+oIVeTFjtlQlTUW1U6klgcDJpUISOlm278OJXNlK1f5ahdfztkdvmzZEI6k/3wTcnviR
/T96WKmrsbZp4v9Ly04ay937No7BMX1rb5HqqW4dZql01eirOkfZ22S27JI26NxLQShV/19o7ZvI
Te8/znwJr4JxrafoaeyIeP3P/Un9Wf5veTun8KhWbk5leK6AegjB9u30Tlhlo9deP2OUHW8bmn2B
acU7Cr2n4Lt0gqoSDHQfhpJ3gTz/NkLzuVClaytym1xdogqoG54HKKQobAeBtdjxwoSPw4Y9ehjZ
DAQ9uLXqDuPYcU2Ln71J/3wvTp6DhqUlp4W2xLEbuxdtRS2zUF7X2nEGt6+JxzPWoVXWqlq+VjOp
krPiYAot/1vOOWkT/IirD9GyHfL2D2V0J48oc+Paze22qjYiCnmHM1GKDYc+vAq4SLoaifZ+OrUV
f2UKBOEiVHbCP5RqAZv/RCAOOSJFG4IXuDUQNnM+nk1g1V/az6SA7ZcE5/ijBC+9LixO+OgV8uG/
PUh07ObPZJvaS71PJMiD5OWjN1iXIPIyOEGYBzxCbNIkdbPUNxtdjzRjsmB4StJ40640zvwl+Gf6
g8/Hw+GcOLTBwz7Nbd6AIgvG1r4+/xJ+Jnw6JsO74L/3sgLH3m2+gGh9Cab2CQVtgvG6oI+JfINO
eanyX/sOYLwSt0iHaKJUaCuyqpv0XrHeFktmtlpD8wMSf7XQwYoVtaNVsY4/A93+mFfbYbeyzg9s
OMQ/I+5OAEA/74uPbdffX4Q1XNHOe2/yFraPT/Gy80c7lEQV719V5CAEiVopkrQXQqy70cza0jS+
cnPZGrk7PceieG/HcnEBzKqRRMUkFSUf6OHboZxfBiIJuKnW+40QC64zSyjyhJ3SHIZQ7Woe2NBa
MSh1X7hi8mXKj8X++IMzdwraD7YSfmYmT+x8IzSVkOgPKFk7Se6wSXyNh5kwE5OlCDYZVolosUHI
yfa6qGdhFHWrzNU+mgSRhYeLjD/7BKOvNswE8UHfyqhlCUUlBz0AemRn85MHNwRcu5aE21N0+g/D
7jl3yuH4G4+U8r9IAJFtyZOk6KLng+6qK9NszBF0X4aYvhh+NlfgFcxxlMnulTHreJyuc0ZwqbMW
Rpa40Y87HNzvE7qDe3OUgio9MEXcP6/4guIjlw/5gsJ+5ekH1ykOBLsSkJED92iM4omAzbnYzCnz
TeeXyqOSD4/TfD/N4H61YeKLJEQUbsakavqSRR05COcL5D5MB9B03Tpn0JatMK9CMfriTcQ6Wf6X
qbtMWmBIZlvaB/fgAC+x+5mkkwSSd/S2CcdOABh1KToD0aGSFnYvTbD5c/nVu0xa11wteaOV6ZKq
PwFDhdTrnN1L8ls7lq32ZW1gviP1GfL60pLf9Rw76PCAEiQS0aGTrdp1NqEMORxFdQVksiUbUL1o
vKSGr4uu8hbhbDI/8H3mUVpfYLbnWN3/3FlMpKpq6k2J0s4J+PGss/UUlRyNsJPOt3q0wcjopJyd
n6UcUO/KAWHDEfxwOXF/UgZCVHNo2kJ/MJ/j5zhhQk+8jAAQ9K1B4h9paBwidpdvVMGWVeWZe72C
Tc87t+LtEcU1DatqsPiZ1QnZONKbrWRz+FSQ0b3UHUz9lnDj4qIK8V5B0jzOgK5j/obf164nAorc
7O0n/E4Rwc9QyrLxFu6+K1GImTRleNZcRQETeXX14bvaKcLVpjuH3FthZ5w05MAMf/ygFmDN0nmP
QF1M0f/f4d1HBepi2BpfnwRHjl6qhGOT2YGE4WpZOKxqJBEc6HAGMUDHIwXgkOsjhpu2oIYaZPUD
dnnj3oJIVYi+OKa6J677vARbkpKb5NmsgNRhzqpZ1/RjbmFmyHrMzzFIpo5rxwuYz7M/8sEc+9wQ
YLaJT/qbABj4mYVqe5/T3wuhBCMtjRx2TQoyoSbVlHrtbdJBAQpLM2VGXF3NqpgK7+vxVZP0uYwE
ZjARWFuCH5HVkIAiswYn+0314hKMeSNfCXHp9yapTTXGPz5+YzlHSxrmX1Kh1DbGkCEvfeX5Luo+
MpgJsyIWWNgcWST7dF0zT/CH8ZZK2Nf5n0gCs1lg/lpPwKnPfW126oOiTcTgiFf/Lsgmi86XUtRA
T5lp1k/istlSmOzDM0/0WoNI0BQE0UEmFrPUmt4tXmvDQNf1yTRzG1sMKck5VYhbFqXgMUANM7qh
ORuZvQ2de5zSSQIctKJ5zkexB/IovOtgOsAOCfpf8REubHt2pLNvT4kZRILAWquTEYwqBtZbWbGN
kBOjLpFwa+PjwedB5NaoPu47qBYKMU62CyS4oYnh+raX7eH9Tl/6zRu0xQOjqs03ujiEymHmZ96t
E4NMfqicqwm5i7xBIRYwyNYaaq4SuvspJ5F0RCXQ95Czkkiq/12rvW8Xj2sntjpxSyqKKg5fD3bU
NlDyI6C1avKCsfajWBNv9zEDlGWnga9M3q1xh8zSXb3CglxR2eGO65C0DSmd0DW6qqXi9wLjS3Sb
aeP9WolpFHkZDuhPrkfFLfZr1Mm2rXzwZXM4KDhTlZ5MfVNpDwiDCO5ixgUakgY3sDqfbMnPDKAs
BPlYXc/VUTPbuZv1YyaduoH9aOUH6qUIzLTXmD8sqUw5lFvBpObWCjeM87etcjH1WkRpApWL2JbX
PNNqsPOA5Apb5HgGcdR6mKixLyO+De9vyoi2UAnbgDnw/0uNOpjJGkldIZI/u9MsTiFihBAIYkRX
yOyssZJXHAluOsnonRX8wc65HaoCa07efrC14qPmoNJ85AreeNyTWNzOWtqC5sXnxfPbBDp/r+rk
/gM++hcXiJZLTjVb2JaY9SlZpicrXX30BtL2+emL34hgUdEvE+E97DxxxAGVYqVfEVObWJsjVGlY
ioJEQqW7vhtUf25LyEZwectJdKj/+sAFS3KIAhLFmVVQQKOXGLMaPSF5ALfRF/GMOj7tvbPgG1NQ
/h7DFgebM/G2LZ4yueUU4q4YR7jgqDLQta3zo/PsErCRdDXh+2Ai/H29uaSCldVmTtvrmpxreIYP
1tsVUgg8vjUoYmOsBREwQE5Pr8VqI/NxDJX0RxOhiZUD2oTm/0UKNaqB5vOSztKWARo8cTWe2Cty
VqacUz6R6HA8Zls6yzDX+51keh0XRTMUZc2tNZkOY8L+tloE51zmBc6Ob2g4QKnoqlHNfz+S9C+q
qV7nCcFDnVzK022HMuJvwP0Ue60tLbOmxoBKTJrZoKaifiu07ROnYSFyrREbgl7+k21Qn0D7jKS2
m0sQr8dMq9ZmJe+1f5gPdjf0u/2wU5Zc0Pw4nAJyXlM7v+taQ+jzvjKmKVmQlrgt+oRhJxbS7e5n
B4mC9nDJ6vNqp9TCueq+eNFBzw2rk+r5/zlWIhgQeMh4rmo+EctFcUh/hg9oqQPt1gbUQUBjiGyG
SC8zFIrjERBZKWu2qGV5fLTfZSCzptLoX6Vmmx7QGJEoGtRvn20pXFRL9Ua6WCDMXK7oP0Y5nvkz
cd6N7xuTRvz1pq2jOurN+AOmd9Da9Y8LRc5xs+2DnJskNaev8LDIxDPgXjJIQ0rakZOwyN37vVOn
IWTrRinxrqHImvyUNCdN9IH3lOhIcLNjFugW1odGPY0BO04hBV1xkM51PmS5cGgPWAMNpsboxhnP
ZnIHHY1jccDhwP7In9Xr8cEDJd3ZDJH3JKROUqiKZ7NOZDXhoybHvChcT7JCXoARoQIKaBylxjEZ
tI4jrTClP+K+QB55c7ilv5f3ZT/xxPbWUCoJ6mB26c3puTxg4VWiBRAeZ7B4NkVQH7QTHV2l7mdm
MCfJaE7YZbFrhvGGyMeN2qKbPFSKhZgyJsr5OcanWxanMd9zqMk5ofByBnFIXZWo9nbL3zzDlH9a
cLQplKm/ZJ6vbtS2Zf9S06Iww1g/bTbAuNhk4RlR4DaUujFCfaJuBkZPjuEsoLTJPT/Z5tqJnNfU
SyUrgsPv8nbK3lOmGL7oa4p1EA69ihBIDLrAgbZ1XgLq6XIBlCrbUxVn+Mtqe+ZYVz28bFBbSuVU
ok2TW02T7y2BIqzgkLWfG+nylagV/oxAtAX3/pKJuhf+6Nb5n9wPQk5JNT0lxflcBwE5D1kwDrQI
JgDpgMrVCjAGgUwgI2hnmuKHgUlIDhhQVK3NVB7CBX5h+QNZxCG4bv5rsXHuHDRQErJoeS4X3pfk
lokZWhLAaVv56scPGlAPNbDVq8shGXX2nJtfPSDQ49Jvs5LBL7BdM7IXUghM8RmJb5+Dcs7/M8V6
+OJ6QLAcRfFMySnlOgkSkMX3yj427gPAWGlIzdJ8Bje1I8ODKbQFH3hIbryerljLW7mJ/8DVnBWE
IFu3EAzPNMqnJ62CwDIfLX2wU0J/4GpjaM1f8Sgjt2QZ1XY+40es39ptUq6BNR6brjccJxilArmw
43nv6sCl4GTnaggfF12MQF9zHZZK5j5FPqXYiMRCkLBeSlZFGP+qFmCxRPB9+q7X5Jih8U2SPxy/
WnfKBVleXhwSt+xCPtyzTf551cEMsfdWodod9Z04I8iyxC24TuB0CLSwSqJV7TeQRuTk1R5qZ8lG
zh+7tJwlVWl59usugzs82qL0QgGrd9qcYxuuH0gawHmcsR2Me/tcCg/wQVCJBk76t7a+Jxdi8rlk
FmnAyFcq7RHv6t4OYakMusegL4y5TNYc7f+GDJmKVNDNkZTvxPSRX0BYNPMRMXQMGwKV1VNpmfR0
3fQ2IoTZoyRTo5z5k1keQuj6pLH/ffKYxsWz6BYoAEq8yxfBPms68lQCvgRrsIhJB4kg1z2cPK0H
K0Upe3+U5kYHiG92eglKUk7sQyGNbn36+9hFXIJzAK5m9Pl0CRRGymB/GPZ5mWRN2ehY9N22Kgx4
jC+yqNBrnF3Mz/IRGcBdTg1RMj+NMkN621hmkwvs2X1/FPlgplOf+aE9ufZD32oFXBuVtYGZD4rh
tM75xM454LAND91GTmtXxW00M13tmJjQPX+c4OtcTp9Z0DOoDAMcy/Y9Q3zEJ+NoRe0IelUjBs5d
RUYgN85wQSfSRWydszMEOCE/+Ief2dzFJp5RDrtwvdZ21R/zLz2dzSZVRDka1oPvSU/hbe9OzwOu
HJTc4o5gGpYOepptCkFo98kkcSi5t8001IGu1QP4coglvdMfMKgbumg3lf+YQ63KjpV3ZJY6kQya
DHQBNrF79jM4TM9RbosZNQP0TXVR1AX7obRsN5XG8oS3MlNuyVq+t/SC6iA0uGe94+I1jJIUJ++4
dgEkMR8cwZVMzqhBnr7l8DFL82bZ9rZtPJiibnGw3jYLLs41O4958Y5xiPXQYTTY17o63RLDkYq7
HP6+PnntTDUEnOt2KV1z68KWSHscvbB14NmOqtoX1hFm9x4QIcae0cpvGXrpkR/njQ2Vlh9ZLeS6
6QB6ezVsuJ1PfwTNKO7AAj1lf7r0ezrwH6E4nWhlvqpHojMkVfgtCcv3HiZvF7+jAJnxR1JUxyUB
ieIZ0iwx9vL2QhpNImsvbSkxgrqGleWTw2u4ZHE7ADerMvLRDgdHDxZK+a7xQkE6IhkG+63Ak6lo
zhNdw2T8xHg9riDkLFhkFbhn3QzYf9Vp5XTjHzakW6CE6g6GS01gbJ1vG5HvzyTeuUwa/aBmYjmr
YykaTIzXP+kZwV+q+G/FFyUoTvNSiy40o5O2reym1tY9XztQ4pRsQ6SIex2IRGpgArFN6nuY2rZY
RkfjMVpgZZju7vZIAlwAz/bIGDTLuUHpvksDvMmQ+6KfXAOaMuSqW4uiqH1263BdOTai1QHEFSvC
asPD/ykyCsIF33IT/qtDaet0ghX+XoNEkzFbQZwKpze2+/hE9RS9u2/Qq7otwao09ofFBv1anE+0
VMCJgfoVMdCx9QXpmb/8xNLix56X/mQotY1denIkjOyabp4l63G6A5zfYgy4PhdrJjRpCuIR2cyT
h6daD81DKX7tx2TyIwEAFCN7Zx+ljIca+TR/rf+TlSZ+syeObIU8drwOIf6vzhyB38KW/vyeLHL1
QFZ+xHdBgTyxIBZS2c847H0H5vAZq0M8MD/EEeSIm1pEC4c41MBG4jap2EVOS5MVjpr6AowwbJIy
4wx4tTlsaBFgHb2r/iz5Nx+kt6W8aKQ0lhQNHrssap3K5zHKjKppbHp4mexnTIhQGc5ZTjyDLnJn
+vn+rviKfE0H05FAMa+qytuyZG++ZNHgyR7jUtNYWpcIHVu2Pbpui+SWjOTcWrCbikl2jgHxWU5N
Zw2bKnJG4HsvFAwEWSbbH0+CPje7I6L4tUDKyBvu7+YMwc7KQTNJN7ZE91JPcdocvwWo4wcNUTTW
u2JQXEL88dZI3+odMtvSMOrqWsxQIS8qb9si+LeKlqKFzdXfzTMninjLyngq63u4bZgx63DM7/hv
72klxWXHm+A7QIACb7682grUDuq/alzxEMfMQkZLTpKD+B/E8s+Ae6a93LJcUH1WgZBghdUd1WwF
YpV969Av74A5IMex6quur79Ocq4eWx64L/oA28PATA0pA/18mfrSf+e94p6pDEI1jN4aF8412Vcg
rIKLPE3UaMaorMK7KxgcsP1LvoAJeSfnl2lAy5NvgC3zjDvRgOan29Hyaz+8/zIxgwvOOx0NZZ4D
rvCHm4ebaTB4Erd53STMjs2G56e9QV5hGU1QgrNnQ9ssqmYc+JmKeJNWURuuWKyxtrvRXB4RJR8r
uBKzjwtF2BMPoWMCDslOgZT9Prm/oI6LBbqwBLTxk9DBwlEZ1MXzwogBvyvGFEI9oWJnHPgNFkqe
gs9X1imHaADiMeYXBUzMjSnBnAq3dDgiiya0kOI4xRZXSqvx7FMyTUgrGasMhE8XFi1wXfCrJST+
KFi+ensCBi6CdtIlVGAthQe+GWVKg9k3xNcBdYOY62kKJBGS4zfU79FUZWwnu6WbJTodxGqPRRHQ
Qsw1n+3dvf4m2pqGfNcKNJiEeM4SxJTtwDlnrJ+8HBpYeESYgob1uw0JmJ5ND0vYKQBx1uIc8t/Q
LYkJrHaYz8ZpjuwRsw4/IAfIJAa3ONRBAgzaYzj34wwmG0fAwoQMfc1ANxB888Vty3Msg8d8burj
eCromCcZ3M660BmnGAcnVoIT5Cf1YKb/a8jOWvNaDYusrnU7RGElXTpUgyPiPZnKVOnu2Jmmuc41
MR50823edea8eA5xGbQnkczQQg01NhYjfnO9nLiH8kDqPqE/vveCCLvhawljMbIBS2NAwAig8w1P
i3VBJ0RXrJCyiAFefI6OxzRHVTiF/ZCg88/YLKQc1yHWjknD4L0cIYljoVmGRUNqtblxmdHrS96i
9Ab5ap9InOrScm6N/6sNW75+uDdaWmlZefbNrp1FevUv3XctUEwavcdcrgQEwp4L7djarF9f4hCp
527EGZZZKeEm4ae89B8wPF3GoVdAYjLvpqRQk3Uwc3iKc+4Yzs+tdD9bBJafAI3CzndyNZiQygoc
6NoZ4l9G+Lxub5SeosPwIrvkRGkIGSzM1LfH0lMKNI0vzSobz6Rm1VPU3E4L3oTVTye9wBI/vWUk
TGLoavCFTyCEpJNRxjuKSYCJjuDva7cgq/6rzWA5zBOU2paEZBd8dexZ4d2Edr2kIH4ipalFwbBJ
co4Q/qT6gKtGdjGZy2gxB/4vA9ZGmD2c4Vy5zUGIFWt7tq60wkbPew/4sAmIydXVj8ayZjigtiwR
31zGGnU4mp4+n4WdVDf7LOH4Kq9vAbXNVCoKkj2LPiAX2gRb0qYfkJ/glF12tFzQAU++p83YHYHr
SrF3QruM/7IFUZTHREKNqpVKZ1uZ9J55FoDPh+lE0qhRTK5qVqmUyqassnMS3u9QsQdkniS9uajy
ghcwxJ2t0jro7QRHVGm0H3TKHw86+sbyawK66JByWjgmVwZhvGcwlpVtq7dUGs4GX+JyKRFrIYEG
cFhdn6lhSRLQw4SzMJHHX7PTKN2C/Kl1PUBwkOPb7EnRbXNtusOy9puSzGl21SqR6IaNQmvZ+Be2
VOwgVW6ARp/Ikg7YrWaB32BuTnERhVOl0Fvu/GZIozwi+CKpzB9kVacldXehzzj+bhN/9R6lJoHv
fFlsuaKFnDSrYXoLh3f6hny0YAcIBXKDA36TTaCBIySHtdc7dK1SMr/MR6daWprK9Zl+STm8Uw1g
1AliRuTfE33tl0hHggLMy28xUaQ4gPm7h7BqwXHp9yjDVHSwKOwpeK9O0NaA1mOooWhjnFVEQbOo
+lJInarLbyuLGg4l4PU4fvh1eBY5waFyWreJmFiSwFsPTRFkoartHXxfsvThlD0d3RAX1VxeoeFk
6JiKFPvAYjMcRsQOKUB0K1l//tNcVIOwsxefsdF7L7xAbaMnK4ZC0rw5rQfF+uHsFi9bzZG/x04n
3zQJ4q0hJlwVMRVbYAo09x0Ugk7jmJeG17zAG15EqqaDPc0iXNbvKQqPybYhadldjmmZ76+sCUib
THxYnOK5ylHqBViD58e0OtLCgfq9IaLjO1FDot26/fsBGHLHo1wgvSlRt4r3PrmQaCattncowHnx
ubkge4SkmAmil9+ak+r3W0VIQlaYSvxvRfnI93rIJ+GaFX5i8uRafe108B+MgbWh3qYiqnPxm2+E
EH3uah0okeXzUwvQeAZHu0EV5cyfVL5NqIrg+M2UxVinPWSsJmUsWg/ICUsBNbKPMNSSEbWQ0s7r
dbbjsWVVUrbrfmYzSAoVfYvPv8ZanT1dm5Wn5fTBvJh1ykg34VuHov8hvGMybnw5Ccpvlliz4Kqv
Zov0X4W6k+lOaP1JErfu647E/xvqd7mz6RAbBVOTkrDEyud8PNS0K+m1HTipd47qUisTnsVR7ZhL
W2ssxvrCffrWIrXcMtIJ/FJ+IzsVcnRjpWUmKICGBoxpYjyazH48J2IfnQeP6O9EC6ZVpVBwgxvJ
sYB9RWkMvnxVa8Yq/1pF2wTfjBoBxHQ/08xZGrjU30VlnFMZPIjvkYN+zR8nm9G5va4iPorwSIcr
npSh0T8VSAjpPwGlln6bISJ49MULGCzUmWTGfVqqwcrojzDxtgGVY5xSZpYzoLvVkyqg37kkVVpp
t9COrhnSr5GIuZ+QsNrrg5SNqh2OBChy7Ek0FBmmRv7Q0rOZRZLHNjQ6hy+x5WbLGqJaHGJQH2tu
Cjf96IUkAKqGy/4a1GHGNgx/8bZhJIrkbAYAhQc3hEo8/g3pkv5FTLcFkTJZyEIvQsqWNhKj+P3T
E4NQV5ASYPq9Og+UWIObMg8zvwGz4tEvf1mCysbYgENMGfTPUhGPxiZv7Ar0/qs2di2JQavNCJRB
2tfUQxLnNRTWvdYxUKxJLdEUaoqBrgBT7Qcp3vty4Fps0wV4SUDSqok2MShfVmjW0dE3jrn8BZPL
ErQow7RGExDhkCuwIq0uxJGU00toAbKIAMB0/YOw0PQRStxguQHn6g5xJv+LvjHstE9/7b122e1m
ucjr2xIJbdeDUlF+ieGVx1UGwNVq1cF+8Zccu8zeUDmgR8bx1twjJXt8Jvh1BXtJBRc3ZVtjXKWi
TcshRs13OWl8TrI+OCf2cvTKV/w3iH4dGJgUQiWh2DL8mcvh7cFAMkz95SSb0PHXZ63de8RNTZRb
Ic8rncKTipnl4sUbJUQ5egWw/sRDcFz3hufKnMGYFhgL5OxtuRxf/Eca66Lkeq/qevzBXivPF0qg
jOgtSd6kPfWdYAD9ggdSXGOziU9pI0h+ChjWOp7tcKjwYixueOfS4OzkeuYDxMAwgN8uKNZVF5hx
H0MY0z4UIZJUcjkz+8w4bNdxDzJDHoXcGYHaGO1EZxK27xjczDEdbu15J2Y4nfZO54mVfhHGCBm7
MIiVuSQp1pMXQmScvzSsHZ50zDCJoNCE/+DEAHSLOhedGrxSpN7wzv8Gfa7jyJhq+hYw8GrvxYcR
aAh2KFlW/l8vQU49roDMNUtemly9dRiwGxUmVobqTdYy52401MVctnjTTd1ak/Tm1mFF8NJlM3Ul
dxChaXR2oQD0sINm7b1qj6BHKshqKWfZUl+Rbjs0M5pW5JPYnSRhZ8VkE+IVoPRStEQZqZQ2AtGv
EEREscUgE5PrOSJdr33D6sup1GzyO1dRENmtMjjeuljqOqWS6fWMXviTPGwnmkk6OruBgz1REdzo
yzWGAU1Ihj/uJHhlEddfizxVDFWoPnKS2vn9LxpaHroAx5mhdy3qpaDH9jHfp4Trbv5MB3ukJX8W
nQn9d6m0oi49QE9ZU/FC3tHlJCfVazRdyHdLXRVQf7G1pXTSnow5Kd9NGXO1NUKy8E5XhMm/OE+5
Z6hLgE/DaLZ2KPvIJZ7OP/1N10NbfwmU5RigR/GIwwDQcW1WxmmPh5VD9ltexM2fPtaE6r6k/mXQ
l1Yf57sl1Xc5hfFIMBZK8SHh67asRVDqdnXBiiFcMp3M0EjNLGzwmvDtd5LRva5n7wxzJdxrkFOX
Foo8MjmlL7czQ8HbW3trPoqxZVJCVCiF2cWiM0SqSFlzu6rqpQDc1+4M66aQufTxcK0c0z8FgAYv
WTQKBJ9Y+zJOLoMG6tEtxIwEWOqsZKa5z1lBQPIlRmZz86f30kWqCw+JTyEd9Jxx8MukMfHtb3wR
7MEWAPcnKEJBjKwj1WqrUiWGhTWUn3TdBbNy8gIq9YgFwDVJg8Xxzg+3L9bOayMA60z1IEr1xyXo
4Iar3WHuzmIRAYR+VL2mvLGu96wi7To9uNA57DcPKpNbeyZvgljM3sqIGlJ0GGY2OPUVBWv0O3vh
xDmjoCeLs8byprEBkNXJoSzKjJvT+AsJUQ98We/j0bDA6rnP/KXqg566+a32fkw+67FZv65c3vXH
QkfyvYEnFsv566u0lCxpVPvkbe9uTLHs4emAZ4k3WXbKOtswoIE+HpKutR3rur9GRbIGalJrrU0a
Aylc47zn7D2RhCC5mN+bSPJTPMo7tSw4F5m6ZEXuo+gRrY/5EQA5YL3aH2n2TcyGyfxW651zleTy
cybM77GrwRqmpggsI/vpWGz2nlEc1BbSntipv8nz1HhKICRZxwewbpMYGRmYBL/2TkxqZXMR/fgs
leX+CAZlGPTwpGx7MAET8ftXMGp+/hXbKzYbYRVkPCIk23RQkumvAe22kZUB94ZqllwCkqh3yyrS
ZYjDpD0rSIAHrpWDeSsN0ofdCdGAK+HzQ82wqUuueIwEglLvGvMxSaEgBAdvYj85+oj5V1e/4FQx
VTelnXbyna07CRardmjfkRoUQRVEe7FjzFRdOrYzWJJTvmDs28zlgetlwl47ZFB7BPBzTyJ9Pfge
VZmb/7tt1IAqEv63kXBn4bKcgRiDkCPnDrD6rGwe6wJph9D/ei4WOSRQrO+JDPOQfTkvcMJZVPAG
6cVTehFxsMW06oXLS6pRf1vlBYeKhs4XqydQXFp65bEaQKtk+hP64ss3nqSBIUiqCtTON1ST57GH
X46JPJtk8nmiyfzMY7fuO5uUuh/a+q/KZ/RgHo3cBnEq1/S0rI9uIGsooHBMHVcAirgS1HgdEcaq
DYHwwBxYr49eUpYQETfjH2skZc4qFnCjyH77mDJRlOyUIGy2xWfGlt6lX+EzUHsChc64KPsYy8Yq
61j88u3xehxeboInOy3tdui7Gw258vME4zRFcbFmKGbJr0CLvD2p+W/t6Z0WUZaT6x7CTJ+sryb7
Cs6ngktnUR4ICyRX7Z53aXq/uovkYmuZpcMb+oslHHks7EPF2IRHY9d1EKJiPMfNw8apqihmlnuA
PWzuo5YptJDIqt8+RecrWdQh6GNwhEAMzsBLf6ILXqAbj/PfZdE3xpR5P/9hdiUtIsZrh8PAfyIg
09dXjlSIDt99j4dyPyDtmD5evLYdfCm9XuzNgi7otBI5AczV22fSZj3e3mT1VVUBH1TUcSgjAvX+
GrzVjUrCM9gDqT41bGmj5bTfuHDf3O+TC9yMOSb3O3XJtygoki3ZpqMqgVTvXmbOxGU8IrFqCQMq
kK6CeHwllhB0GojKlzKml1GgyQ4fWBaZLF6wwRAIrEXqaoeDDV7Twipp6TLlB4Rc0aGWJAPkmsnR
ne/RJpguw2eQShP74SKUBIUN29sg2F5r3mZSvaScanpOfHc8K54ziDsKXz7qKbGqOaBdoQQC7e4g
fNU3TxoWUMTkvdfY5HRUtlkjAfLuWdrVTx5ycMrHcll9cg6YMd+w1mw+FKWUbAayDw+DDsMbBXNq
ZoZtU+hlSfyHAQFtSsQ+IuC6YXTVIDcoU/fzfivZRuKakvlhm7C70eQanv5ajzh9GrmjiJuPHzyu
mE4wee5BrGDKrJKf4flS4sfIrAYhCVIZ+xovi9YAzR/t6tXf+SFql0RuQMmGms9Q2f6fvqwgSyW0
992cYej9qWzH8QtlIsvQsf7SfmLPMH4qnpPPC1WwnEvaAEdeEd7ca01rIhbqSs6xis36sBA0TlWd
/bErsczCK27ZMJ1Uqdl11Src2DErFCqVUC4K4JOd5ygp65dpzuKcPjQUMdWWFqvuO80QdEatq/ib
zimcJ+HSxm/CwTTx5Zil4//4xSm7YHLkXBtnMyNr9JAAlugdjnzbgzig1BjxEP+EG469JKbUJOtZ
a3Ii3gwloCF3a0zonqpoPIYKu3x8H8q/iAUnfB3uuWSpQuUu3YtybBM1S3qrXnZ9gr9iVJizAhzA
H73KjGAJQBLw4LLqngBaU2/0/MO2egiwvA1wSzsiaazxbxO86QxriJSBxcPt8Cc/Dc8STKZFrIaN
JsnkCojbEj4AMyXtdo2wuxI6oV1VFGBNVHZQZGpFxQ4W21rkUA4P9Eh1xeu36D0mNkE7GrLEpe9d
dwZkbo/IXtKHWQF56v28ky7mhT39Ufn9DacNVA3Dz2HhVC1e83kvLGoGwAWJnBOHH6xFbMLN8Jc9
7fuvKkrQTGK/aNgplPaPPj4gvWdR2EwmIQLbUKRokiSSxjZVuG4+9fm+xy7mHmruHMr5dtoE+SE3
q4I4CZL1RYXmL1kkrWD08mlGCBadFKiFq7BaCxArfpBIwL0Vez7OGGnzbujNPVdpTNohtvfOZKyw
Yj9THv0D9a2vnAY6G9I7ty4Bjk/CxVGcOWUE5eIePVXATDZ7PbJnkamGxdgd9SCtEqBQ3j0m1OtV
t3VkAc8ivcShkiTeeg192/tosYsB1bnVhgqpAiI2ihknx0ENbP+Codb/4ciPWHILip8g9RsHlVyi
wMxr789f7xfkmSfMBkLA0rtVIEg5NaW46xMJ4Cr29NrcXSAxOdI65AxtI84MtLl6hAopSAl5dg8X
oUOaQtpkzWvXBzkI6yesQUKS5qmxdcM2iMqUwwWFXPASnMuGB7AyRjuhN44mMfk2C2GFp1aQJ2KM
URZ0EasLP/BDCBeQbRZ0Eqv34vCN4toyyzoBTR6Hpp5CUT0YZcv5MMfiDbDTcbYAUg3y+ixtXeOM
GjSUWkZv8oekNZpIpbo3mO0xbY3dxlSLN7Bhl4/qaSyJLWx6efi6TpgL/B1QTIqfyijFH/RTEHPy
wt6EYYRzoipacJgiN5AJNWYeXqFJl+1ciWbezWBOhP+H7izDKv4SErhGlRYEW9M9lQaIH5FAkO41
N2cVOw2zcn34COvlmnfrZmCDPSXbMT3i3Ov+4kEBu1bQifJ0tYEqMrfi2I4QUX6ym7WFGj6TyKn/
SiTw+M6btVr+KQMmcbvtVEb5nnaJa6WlXftdOPcBsqy99xpd7XHifxhfzfIWgZ8HuFz6TV/X3hCm
j02GMJUIeuLGEbxQMl4ZOIHw7aBdZPEOc03CZruMFngBboqlDkHpICPJ+Y2Uf/HjOKipUPF4gamZ
WZe6IGoCoDvqSzKQkNCbkqYJNAZTaMJBt9OaTfrgzStrNphhRFSrfYgVOaVGYbw/yZzWtEbRX7vs
oCL45aesY1N+ZxALvJVrdcaBWp4G0hOs3/ygP6ZrZzTbprZSdsJJ76cSoKm9/y/7mhaCDkJr3TvR
1k5fC3cCZCNKNCNdcGCTcCeQKBqr8QDNfd1fFu3dGZdyzr5VqRPCn1w3jCOm2HVzgNskBX0JIvRL
oizEW49cpCdGF4UO67iwNMWu8o2HjSugJDT8HhddJcd0G/okgtPrG4K+/HLnm5bwyQcRHuGaayog
aSSzDqZk9gus5dnsksJePNyuD3nTUfZlQOaTLxvNjXLEsOMuxiBZ429EdWE3d+w0foBErIPtYCPT
2xGTnXVuROSvynSP64Mp+0Xy0tBcxtGs8arRT3ASNhNLe74JzYhjkCCd+tEuOlD34oCN/stp5ibG
hh22xPfhHVQmAMJdStz0KpWv8oCwOn+18XUdRrQQ4YjOPhX1sChfK9Wi6IjGS2aKx4c+LD8Ycqv2
msy5jQg4r1L0dkDMHoI0AhcDwmC5YilkC3iHznAujA3q7aB6Fx8vTPEkGNwgb96Cft/4E9SKCqd8
KpGnQ7JQSub6cNLKNYiRYLRTqTEqr9Q75ckvEb2wLugo303JhMjrFL6JJohQXscMTxdo6h8D/aYp
zGjZoZfpd1Q6MwIfb7wAJ2JYtAOEMCooL1mrHeJceKwJr1tXJJ9pUz3YXZdfgbN0d6TEkPBK++Mf
Z4KzGhifS6YzjQs+5V/FJ9VWIP3QebJzyhGDkUfIPJMsM1n7A0j4VRk2UIBzxPa0d99zeszz1Ado
82aVwDcFPJ98zJ0euxo0KbV1/J3MQrzgHM2/uCVqZFOsgrX8jQN/fUE0gS3xy224YZBRRk0C+yM/
aKeBW79P2N5gYoapHIx4pNBQth8cDXDin6L1LOlIY88yvV3G6XzL/BVUXt5k4aMnry6Z5LY3JHhg
/4fWRJmHy46UREVmjeCy+CSkXA2Ip1Hme/k0x2Y8e9BsOXHPNTAEP+CbORm1wd7jvqcZ5NhePxSB
kwMJVcJWKapXtf7UNy+xUMiSIMHn7mKGt4H4WzTaGiJPWYnvqzfGtKm16BgDxW4sWoDOx8rtB0Jo
kxyexlSnC+KDaKrJOF0e1aoywgsPAUPIahRt4ZnxUksym7nXF/ZVAiqK6xUSmJB3HAsidZTuQ/3I
aU3jjLRuMz7QjcQzjp2l/yS//13uN6UHjysf8XW6vTzuIG3uIxcnMoM8BMtwxqbb/GjtjEulikrN
hfO8ulTi2Apiho3VFrPX+YOZi+16fm2fqVtW4WiVTZOUCTRQ65tH00V2ZpjQif4vUEbYKCmjDOz1
PXcWH5waFmn3iV7mi4IT5gOHxRnlttPemGvZFxYcCn8DqP9UDFMm0NkwYqmOdpXrQlsna73maOAs
9hdsuux1pozBzk4R1e9kxC9Y92dk9fF58jhQ8tYcJNkAiSWi3sODvGbLG9GhIANZadUfUkWa6o56
7szWCo5UFqcoGDtHlN0+qnlbBdC7bgdCgwp+59Cu4LZ3UDFjN2yM977qFbIOfzAkBD/LXZZ4/vyF
HmwwjWul0i46bsVUHnbtPZuUnPLC4wKGPHEjbhHolHPZHYQx1XKRjR/Zu/uh/QQMYD05c5ezEEAb
6sWqc7U9nmsj1Wkk69MCJakhgqzKTD2710kJ7F7TDu0hONvhr1bWR3iplZGpc8dneeTX6VQGRxmo
04RGXHKBgrHfSk6VzYHV7/+Zfrs4YFmrgCj7saa1u8z/nDeQa6K8sQPO5O9C28TGhXBFg540flf0
SLnoazYGfWQpT2QhIVtGCpLzDeeB2PXGQZORv0lZgAoWtp+qOmqpRKiIwSercz6KzgzZXh78pm8L
wdFGmFt4kF3K68FO/WcCIhZJsl7zjngKenRd8hURxReTI/C8T9V12S9Vqes8YDJVu8fQ70yA6oXv
YEpWByKb4D1S1QLGsb6CUvBCsbp32UD6FprrCVpVjTtCtJTQNhpqYK2ujlrkblojq5k0z8WQSrMU
apCI9BkI/wc6uiwbjlTVOjtyblvW2q66ynZtvahWX0GD5ou8nt2/TpJqJL5R7Cg/1CKyUHLaxKhq
rY3MhLms54gxMzSOWVfs25RhEXaaoAd5ZcAel8KfVf6Fi8Hf2/+gX7KhYEOLVXaRZfAkMeGvjaUB
QnudiEqSRTHzl7NxIvial5OYvLS+2whtbwvB9CuC8Dmz1aE23riVh0t4UAiSlFaaFyXLQBeT7Iwa
KjVtppRS+jpv+cpxZxiq2LCO+Xs0ofzyD2LXp8U3drRp8NH5gscJd1RlHPqwXAvEsIUTNqANRiyD
qMs88tZXhSfOI+P1Rm+k0mo6/d69P2+IhYdwml89RpfLViqm5kWq9wNvzRmlXahjzMsr/DuVUUJd
G/SitgshtJFAR3rWtIFc4pJlmiy0g3M2v1dl9EK1n5iW/j3ByW5qvED0u7F3gZbfNXz9qcG/zK/u
hijujnZHadXkxNt9uPY03ovRwlbzZwIVxQikAgk74t2+JQDDlMHQ0du1ACaalHIL/wwOQ1hQQ84T
dGdwl6IDiyaIGq6RqiQ8M8NfEWVNAIcVVbky21815uTkX9+tjm0RSqUQV6SsOxpirFt/dd3AvKZo
DSIgCikpKIRzYGRgioGy2mV3V4foAyPff3a+2KJZqx749Pc8jNAf6M877b/YWcXtoRJxdxHgHyGM
BceydbzcEWJc6YqBRptOTKI9GIZgJpP1rkMZmwB5SCGtK4iFSnBiKcWSwRrLKGoHrqNQuAZGIcWX
lPUHOvWa2DjmAMnK6koMxEliADZ7P8YAqesUtVvI87094eRLF3sbrA4zSO9kHN+/j2mMCxxuZ3Be
B9jjABK0WeOSCmDNQOS99CQX6Q/IQVuIJhHYIoUgn+gdNKcdRCwmdqnh9t1hnBeNQsBRrUkD5bK9
xhhfBsBrP1w4wPO+4MYWUHbrtDr+02e10+Bl+0rf9IUrUrOzVJTqj+zy8XtYEWDTHOU6FOzCznYK
lGrl3oYTpQPYcisiL99h9NN+ig2dOVGaEoxrIAmrNnqexaXN5voEAMeVZnor94z/FTMDXQrNjUNd
QQ6qCJSw+8AQjUySw789GQOw0a/N7DRi/H+PiCeB0gjAQbbTIMOAFbfJ81FYOIKGOl51cvoAy3Wc
+zqOPLjFGmUZyLXfMFtXgMqk25lhH4qLHlfYcIIDvqRthEsm+Diu8IYx1Wfgeom/OHkCKGEyjd6G
T7wUhGJLp52NfDt0p8KU1kNGLxqpM+4Ly+hw/xRclFZLcSjw78PVi18luDULRK7fN+Huzr/do68j
S1DsGKBJlJL8h/KRDfh37Vv6qSO8uAUN4+SfwPOEh0ShGhWjpwMBeRfePK0tm/bNCgzOtg9VVB7Z
09hmrRzB1qWMIHfgfSzPNggskIw/U1TEIQZhpQHzNyGabBw45N/DVfqV5bsm/kMM5+Hb9diqCK4U
j1OY3z6qbisWWhNZtF9Il2JLQ6uKkrrLGjNzHI+CRjaXZhVRBUuhTMfsgw5II0hJciw7VfnEBzvN
bsf3TAPG1v2Vv6RtbSSd/xHC/Qax11GxepotfAQtsksbrM8x+j6F9BZbbwEojWMxohYAuUkK0ua2
E6BAQd2uSPNDeliaC0ouL9A6o142wxt6Qm4GLM+vJRRg27XnOptQabqi6XqM7EYzz5KqISrIrOkn
Dm9mqkOlhXlb9ZdlQ9hFVo+AKnfPrskCndjJEjUfn28Ie4SDozqKM6fjBAoWQyITVpAM51Mj8cbj
0XyaOlRXSVi5rP15EQBHcLr3mXIDHWf4dHmTZiqNk9hHblju7cmdcc6CCvoyiKTP52V8euaj4jwI
5ygmb130sFEqnhTlRsWRUajYF3Go644xjNoGB2LtkivxfPLUZPOd7+tusyemKT4TiqaiF9aSDaZv
m+pEave3InNMXAcRfR8otr8DABWdcvmz3olUmAHZyFgCtN2k3YxgtbZAAgqr7aLMTFpIZBaV5V2o
dsxvU0j51TR26BD1r9ZTgk2LgW86rcz6Qvs1RsuV4+C1ZqlTK6U+UbSPPp+D6ap68Lu9qHdwyfLq
5cyXeO1EysPsr9LgcpHaONfuokbfmKUuC0g+LIqS0TUMVjELI+Y4n6BLX0a+jDFyGiThl5wEnXmM
eBMZq41KxlJHb7Pww4inqiRU3QI4aPI87M9nz6TO3bhgEQ0TAAI/XBVb2zW00GRdmoL90R1+BW/S
J9+8a9Cc/hQRxIsmfoRYXub0JTGZc0JF4jKE6hKkE2k2gaJlXu+15EEW/jGcNJYcISQklXPqdR9y
jNhdKlCpyigS2YeBtPUW94JgO1+ypynMDQ+zoSPVHfqm68jVDIQv35HodILVZyCO+UYUYzVF1a4a
mPc3c4/CT3hR1xEv9z5NGFIm/Z7isd2qTuyVQWHeyA4N9yfmU0disRPxyloD3qqTGn2fL//kVxjY
gb3/9YIF97WKqjy1TOonsGGIMxAqJho10RrYMY1IIuFIV0s+VWlZgVGFysIk1z8+Ea482dVPjK+J
tLTSWVyaYpKMxaBSZk1H0bCAR8+4GXBwSbvzOmPQE6ihBLOxhEONb/yUJwvIX2MhYOB8Fl42GaTt
wMRbMcbs5oGDZZ579BNwMLvZNnRWRNrthxenBkSorj8IK/Y4ObhcGPoetG8tmPuBwSw+gyaRZB4F
dSmptaEV2BTsqjHT557HWAbsP08eNTdOfwqmu2dyNpngmCunDWkpPaR0UImgqga0mWh440azSRU5
phqRHODV5Tb6VBG4X4TgL5PmVouO2T0VpcCPoEM9efnVarqWBzyMgKaXPTIXUQHgz44UYijhQEgh
HQgt5jtjB2XtZ2xXZ4L07jLGklOBydbvYwKR0z0MtqSJCmAmo0E0oYh2YzYYkf9jAnEgjnrys9JH
3LK8CGXZJt+lFeG1UdLRwzsLNG97Mpjjuf0BENxYUKQKfWqbgnX4sM3HiTpkm0Pm2wAw/3ZV8PYu
UB7vzuny7yBVA6OFdfJGc5z/OT0DdKIv7KYdgNF5J8FC5z3PxEB3AfEfnHlwA+IPKYM7wv/SqhBA
Gpjflz7JhgOPgkl6TKx8zDK7RtKbvqhbjITHaKNoH5FS7MZ+N5R2w48qQfeQXYbyf24jdRX7OyuK
cT3hjid5Nw7TwmUa7y0Y9dJ5WBINI2uZvsvO8Y8I9oN+nC4fhb3zg22M+N/YJkgJnRN0Rr78rPFd
Ofh6ftNv9wu2Vmi+FTfj5zczXdD5NQmi96KQxjVXsYH4Md1oLq777uULGtVRtapBI2w7XxsgOCS1
Ph07mDNQGPL4azOxMEi/jkN4r5yBhn5y5aUCHkSPKzJRT5fKSjv9jWJQB7I2/kOw6pH4mLG/TIdC
/74sjZZmlWNaoFuoYbW5XVicN8GDP5iedfANoeZqPuudzI3gnQgOVcihrB5KV9ek5/5NU9wsewPb
ISm//Sr91/XaZ5sPPeiIFys8yKnx8CouygmrN44+Q9nY0b9qZpSHOnAGMb3jnIw48z9AbwZaHOJU
6G6xC+8QL4uMUeW3opeHvv3WroUiDpCQDqGlEwrWZY7JPDSgMEIgyGZU1k/A/F445dc5o/MeKvtb
R0G9PbxGkTLjHr7oDzziNfBZUXUpaeUt5ulA7tYcK30mdB5x854K+CDp2oO38O2EIViE6UL7vXeG
xnX3nt5LpAWWSCbdM4yDXTW4GZ4UTrDEvW1fd7w9OMUnVTjJNc63RrBLiKtG92A4ozUpVNph8PDv
cYkQDcnO7OGYTVk8YIQvvrUMxw6Ui5rK+sdARP8kksWgQRRvh5jXBUxQJpHvduBAu3QB/1YJ6rVF
h0mE9CzZH87BgBPrlATFqMCRIElF47jX1kdaJRNDnaBdSRwjQBf1p6UgH8ZTA0wRp4ZFj5ukOYnJ
pGH77WX3hW73olxLKOTXr7OTEfGwofiQtTi0FW7ArcdmS84xlgd8F71kqoyYaIXu4bJ+Dc4yrW05
071ph3O/tyHyeILo/BGmT1AEAywX5v4Jlj2i6m6OlpIPBcwKs2JUGGPXfInYdkL2EE+ywBi5L/sC
UonpXzt4lQPEwYbw7WuTT1IIE84d9/AImBXHAGiSnXI5j2opBOYAM2eSrTOSbgSmgWMwDXXV9sVs
4cO85j0bDRBRWqpIfF/a/mokMTG4wZvvge+TyfNoXwCnNWrnn2o1hBPuNaXtNfFgbGP/kUCiaCW2
Am4HDJyW0p3NieFv5nKNp1aqPy7RPdR+jIVIFwCRxmFga6N5uo1uU/st9S3LhmaRo6HQw+Zqcq0o
vMkdX+Sy4nWFQOTqzmV62DIoycDSfqksgvUKPZhpC8uzehFzQ/R91jyOh8tsiAJ3Cz7sB7K1EUYW
XoyWeC4AUtKaJ/V4AOgrEQ557bnWXHAzKVQkPEI3cbalseMChAJQGq5iFYAUasuWzM/qmPXfYwJk
mZ2wHDAFFr1p3R0NLwmeMRXIdV8rhLsCrSAaLFJuKrJxi9cag3KhIZT/tlGNwVMxWKtnJ8HfPNN1
B2JO7EnWPzHbQ8oRW5Rcrl3HfMB6/8yEbZ2FGCcxYn/2F4qWA1Nv14gnvMTtCk1+ZH92foG9x5pH
CiBHAAyQuLefGVE/F9pCEKxnJvFrSctptb74hSkBBFLHhnEBhJ3jnlRyQsp9q6o8HBO6pjHA+Log
P6mBd3EdcdFqNhbOvqrhJH/pqvDSSC6TLjjY6dGfRgf+wHkQNVn5cxlcSm8TD/epyv+nD1qQObEm
/z72ExU1UelBNk32GFw/zIjHbsCh+3rR65RRbqWR4QMjQKv2X8AO8IVew2GkzAoRUvX9iEI8bC7W
iTZjUqehE6l072XaaD8xqL5JhsCW31SjM2h4+ntd+nC9kOxyhNkF6PBeuby4FWa3lkPjaf1yhaES
pgUPYPWA6Jed+ij1+97+OD6GLcBIUjkbLHcaalhzJE/KIILj7bnINIfknVnHtO1wi+opFuZ+EdtB
okuDQn/70tCsqHAqX4iEd0xOZYU80yWeKXn1+Ilv/JRjEKDQWwgBdHWh6cf5CkpOlNZcPUZ38vDF
BF0KRBJ2L+KnSJBNcoIwe+W7DB2TC2EPhYUA01aQiF4wi5R9FzMygx6w3L8xSuhKlDGq5qVjBMt0
xk74NUmMD8l27oMFkvnzsSeljRtWa4ga614Hm5/w8m3EfKpyxc3QcdZo/ZEFnVsvXhhmbY8FidFs
hzlm/H6CDz2sSLVbpg4eeTqRP5mVDD+AORuOEuSyx+izDTmZSTsCrQxfLXpFqQPwoINvszDCkFnI
f3gU0IcTQQRl9A586ZQo42fa/SbN9jySrbBFNzZdRUUTUKsU/0tcBI+y9C/AMQdu40RJCGSIuQM9
Ltczorj3aS668Eh21vjmZQ2p7IeTyVUqkBSbLdJ9r13aFBK7q1OPFL5LHy3EpS7c8l1Pg3ujvCZy
CBmzTwE/t0wc39jg76vLpXhIKpBsXZGsofttTFZChLswKjyF8jp/1QJUi/HMB7RbX8kHHUCMLPuV
Ruh/dmk1ueKyvA8fLZbGl6wYDRbg0boDMqmtF+motYrRMp2Ry1iuSeHnjcfUu2UWmoq2p7g5TK8l
0dlLp9OVv6KFc1wHOoe3qsjVao/S7LDy7bWjxzrI4/QrCffuhGeVakxCJrhfejtAJnGe5bm6xDPx
1plDTp/7rZVFbrdTZDIfTVBk/QTJCeDVtbD2px9VHnN9uqjzeD+vS8nD37ucGWNkCuoeJVoWEeYb
iHbVGkh1QAxqwETGmVMEHBJp4PryN7rCI7Npq6ctECvLyqRM6peKrhoE03tPI+7OiVShrHZqt7J4
QuRFCjgNQ4dOvQpF97cNuyiS85869JAawnwtt8UZCV+Ffo16d1HxyWMQ7PEBjkE3SrqlmfIEy0K3
jOuYbGs3HrwAoE/3W5lUVAYhUFZVJtNDIhn2dePcafwxheOyKYI7OI/nCs5LYmvZIYmdZecvF7Gd
JWtYUpFihDjfMi4Tyofb02Q56h1tYDFxl4lLsEU1q2CP23+SR8PYXEmFMq3i28rwxS1eZvhS40Dn
8Sp7EgZXK0nUIgjxe9C3fSgYLGHxxykc61jmcPOcniH45sW/GTKbLRiNhQmk2eIk8KJyy1FU2PcC
b+Bx94QDWI0lG0MjD+E+FioMn/t+tMkD8FOv3sBPK+mG/DpmXg7wx48SyLLPIPK/F9g/hq9v3XY5
5Z7m9fCH1oR/HUsKrS+gFSizC/SKGB9YZ7jYfNs2oaLljxCRviTf+1I0xGbpA1EAlbRH430gIpiU
9vhRQvY6AVdHNZRLiPTdCZOr3BbN2iNF/r65A3gcK0pSW1ZYmCj///hPWO9AbWfbvZBNfWAwULyC
Ot1uKCN4A76ji0hqDcbV4AaTOn++5jlnACRHULTQ/8mVjl468Vf6SnwbRXc4RNZm9NpwNV3QAGPi
n3Woi87mDgLvWHroHYKC3nJoIPIKcuTZdMu4Y4/MTQ8Pyre3ncYGL2Vd3adBsHaPQ2gwDQvXNWeu
FCGCLNMtAi1gbFeRX1G/FY9r5CK3YKTUwRaEH/120pzkN7wzTB/exFYuqpR+chwJGddikNXesPRz
kEL+MiuAi/YQao/bOwhK9E0zNMb0rqYRiyHN1MbUomEf1nPis6A78hMqZj7XvarYo6k4PFMCxZnc
XPjmuVNpHxkEJFl0K6HNTkTayuQAeZJbMsoWZg7zFq0xs7m0JUrj5V0s+hcR8BFiLdJCeGjcDgyr
NTON6R4Yyb59lIbw5XgQu9Zyy0Wtm8z+9iIdB2wx2KSXADGRxZQH8d6S3xf47CufJ6zSF6YR34GY
v6muJGOm3uQp5n5VcFfKTvAq+MV8mbx/vB8rAcwGNX5pqGOW9yYXYy0p5iT0V9V3sQ8BzMKb39dq
HZ+HOQ4GI9YWBZP+Ih0c7seG4y45rUOWbuNUhpptruHtWY2bVqRjp4p53NnZK363bjaE9aJcg/xL
/wDW9IBdebqWjaRK8hgER6TyzloKvUA/BykiR5yN467Xa9Hb8pTOd1wC9wDRxGxlp64r7ceypXpa
kymFF1d8eGh1k/q3OtCAAA/oYL4CM/Egx3HWS9BkSwyTZ6DsoqESsHidtBM8BO8LKw913sHwARQV
ReLzfwK6DuNtVXxr+n4rSW2JKzW8XxkRXrnbcyxM5H3gYDjOVgcpkIlK7UCiG9WeWUqggeDMtr3T
YzMfPryeQugqiYNiIEMn/kPdkV8PaYKHt2cg47RBrp3AeXGU+LidOIYhYi10acJHeg11NQzcEMdZ
B0AsD2iyZmmhtx9ho1RUgeRrTF5cWOytYysIl6RTLrYTP/AzI1jT8h7I/UjUrBL3aJGwJTH2Jjac
kS1XA3UA0WiJUsSXZUAhdK9RSpA+Kw//eYwtckFkCVIhzACrWJ/dE7W/a8lrZTckC2BrBkAkoyMk
7eQTK8ft8a96p0ymwYQN0+L7hOmtbdMdXPwbAYF2NJqMEGQ0+7PPP5CkPgV/L1o/8nKwJ+4wIJLj
Oy1TAE/2qx3ypmIRBooZ5VptvU585ZWJ5i7aQ15Gio51XzzngxenpXjbZIdGlzVrPILpcBIb1nb2
w9CaGVQxGsU+rIsO8JLupTJoD6+lz7G4GBvn7AXcYI3lUQWX394hVp5SLCCX7c1EXZZP9PXTfQaV
AoUYih+iEFxL1xgZsEFtlC+4zmeqOvS3aTG/zGGrM72d1NH5g6Dwi2f5MhvnFIPvUyHmShEHQvjn
iYzyTArgLOdooMr4DMrcV5mxrvPMxFoRnLQjKmM825RsGKWXryQGUfwCqS5H1zM+CvQ3D48KksZ6
CkVIyEle11Ud1l2zz4SNIALz/OrX3yyb97VyF8Ha0eRp2yd74bNLY4HapuETvvT2htoJhOiOPOyF
RvoendSP/boJvRSSn3XfIliW0ghbX6r9JXQ3V1Z8Uz9kYLBfnfyN/kY/X8eVhRD1B3iFKNnxFgC7
Iqs2ukphFzUmptgh5xBf/TFr2106D4938UOWy2cJ8ydEAM00F9fAe1z7YIDfqmIFACDTc2+iqcH2
EYNQC/9GOsU9vuU1souIjBm5k/42yDBJ0axid16bwk1+tYdr3JSFlYS+jZQTKq6IYhHv8+pSquyj
+Driy1TPLkLVfoyqmfzwgZoGxLQXmzi6KQqQ9odyg/DDkEJS4oVYmHhzXBJrVSHj0M9ml3smHg+C
iRW7UVTtS5EXelKJySZMZK7A6pCaQnI4lJNvkci0ntxG6vvMHlMv6y4+in6sTp8jUWjjJ/2Zj9gW
yemnc4F5i2KQwUDeNZ91KLLrbpHjR9BQE5E/OSLRs2zffgjJEhXJpTDJU/T7O/ip/6puCIy2tU3+
7v9N9GYPE+qJoW6MfZtfrJ8i4QHAJWbvpuj1C8sTBTQTxhgejcWteV9Ixi8jPgvl665L/xE5FI8N
A6Di+8kURne2Kg1mRfqtVybvqOOHQOoi03k5uGu/SiPupaxJBslIUnDdeH96EljsDaxkMR90Hzu8
NpbhBGtMNa6O1l7+VYEEJTCT9lKxM7bLDhxPfsrNwCuE1qYRfrdK26Y0iBklsCk2QemnqJ9Y/XKA
Y8u6ReVM8/2NKTC5C+i0EkxXPT18b5EBrr6PKl60oOcUtTi194JDqF8tQ/9DY4yMONGGT3TEZy9g
IOyJs7O5bmXxggdyuiBCY7BEjIXcI28d3dALmKMKZvhi/eIpT85ocBZulhYgaS3c3hjc3oRaF/yp
GVQEgyPPjOOIgJ5th99B7lavrCVzT3Lolos2zdWfsFOe+pe7YuAjp0zM5EL3ECQyL6G92OtK7634
3vHeuevYaJspwMX55qo2tgML/Q7BH/WzsRTksWNjJYHyqCHckKLuxIZAAeVe7/JSUzYhDBL1vKm5
qMzbn7/tOPYFMfbNV/Vlq6ovukFIOfWOuGB2VNicSSlkxD1SgPcNLnS3bgLLadtie4Nk4nzoleMG
zAB9IzxqkJX4oMMJdESlgrUY0mroi6ofKc8WXs0edgnAHAlX6aE1j9IUlfN+pjHuijtyMHxVo41O
Fq1inNht126Cy1lBICUsvuMvavgIUOMVzL+TEi/L69Z4tBTimcGQ8I0XJQqALWOt4cnU+g+nAsU2
udpp8palVjzfGhvw6HKBj7vJvV9cEZ4cbFiGxPjeJu6+6Do/3MoJl5tjg8Cwesq3NfoEdJUXyZuC
lvIzxsRW+7lRu1CriTdHIbUFAQyHXe1SeWJf6tq6np+6EUVzot63mf7l3ASNs9rbVdrYeGsmXrAF
Vf/bxwa13bMoJha+3BynS0qdZOWNigSPebQaHVP8ZnReOFbFqS3XWN2m+93UBSoSMRdwAiuCM0jx
BBpv7pZ0557ucEd0BcTS54U6NX9XAh/JMoMI/14Vl9zUHVPpiCd1ppHV0fpoHRXjQ1xoG/OKbE3t
bGfNg7WvaOydZiQ7UTFhS37UhBMsUH9jwtLYksPG/3e2vM6iRmzioOo/t4UsTJT4bcCVeHOarNAY
Vlaef2WHR0GGMIhVkFem/xcleZvRCFXrJdJ+qH0gzMJ8jGd99T6HfQYU4/sz3L7inMGg/8YAOQOC
h1g0fsNMI0BmOA6TI7Um0rN8bW3KnJ+i7tIycJLYMVvOdSrgZCypEskfHdjL5YDmMDl14TXDUZSi
PtCzWurZpWRRggz7ITe/TD5G6lUVDAAqy5x2iA4zHu4J0c5A+1+hPKt7vOLDWBumAAknI4PMX3Av
02jIfkUJwRC/H6Pc84uc18f0Z/HUOmb84lGf4Af9r1O/PLtF1nnr+mRwmY8+kyfkXRwcnga6pB3u
dxj6O15c5pYHLutSdWbdsW8I2FbeQ1XKbW+z7rVg1M4oIVii3a/ozw+DGPo0yuLEJ4NOU1x1/nL5
fxAM7iJBZNzO33FmTAJQEtERJn61cibIBm3aiVxk/hB+5vPuWuf9dnqixYzGGVnBTd5MyYy4JDCl
PPA1BcpJAaMaDm2xJmUfUAtOJTeAu5TRGWNN2Mz+SGuvo9pvPnQ+ydzSWUeGM8HVbCeFBO4X1Jfn
m+dkC/BcEPtU6j0OKQt2ey13sxNuDRwi/xCT3iqlaPyO+qlw5Auf093U4jqnsx4hq56PZQ7RC6DF
nQGtQZTwQtON5lujOpnNY3troyqb0nnUjklNZMAcP8KCs/han/CsANxdE3Yn9/TzvINgZkSVOvWh
qVkN1OE3hWd1v2EeOV4UMRi1+RJC4AHGOLHKQJkGw7EGcfIRJ8YEPTBaIUVdcJsJ6G+z3ZijnWwY
5HUP4QIHukF7yoG7zyGUelDzMWu0BfrNMqs/He04Cyr2cUoBMUgALe/hOuxtjC0gffcbmDlGDNUf
pno2YdHNyFfN3FxYS/ES7jEteAow+WI5UdT0qb9NUjdiOtKAWhPMQB0OqrPU3Mn2KmU6YCIZY2df
UZRcGJh5Gg6274sJjRrXRkecHbx+Is/sj+JGqiE41/1KzwrYsk1gtI1rb5Wn5fFg4Rx8n5W+1mQS
a0v8CmI41Ih3+rYTPNml3XWZ+dTpyH8nm8iuP69b9uJGp34R6PcTINNPnnO83xrlh9Jj25XazMGk
6m8T+LaW6wNZQBIdWC2QILfqw+CE2Ons6wUtYC4hJYsX++ZwvboDtft8KbRL71/Qyx4Drx5wR3FG
kH3O2lITZvtA/7xyyW1+vXtxdfA7i5VI4AGbpr0JpI5FjXLVbC9iLIyBnp2ZBrMig3Sp/k2OvZBE
yyjXZVbTBRh1pPwHGR2fT3AupS4/YKBC78LS/MHHnjkTFl/jlYjhpCPi5+2iYh/CIySwXVqRKJAV
1nt/BXzdCFplBlgewPqoZT+q1P4QNy7It7PDgBsjIEJvvOhzlxcawh2MmlZF/0OpuZJCLcSBRhVX
fkMfvR604GlN+ny4SXU8ygYsFe00kzk13/TJDGRgsy2H54QH2r06ospJU8ONmUCqqGUUs138QGie
w8zyG/Jd7g5e98lmlm0wDAKMdSipI3DMSGX/ZCN3yQEKb8zf38q1CXdxI4ywgx3uQqbTIpoLZ7Kg
p+BTjoe5VlbO4e1/0vwceHDArtL2p6iORHMSr9+P4c/8W739FNos+U/hxYmMGNiBE1/UbFZcSQKq
8PKBcU7WJ0iMtrmrGdI1dAQmCMEStM6Ew+UxdhLmhYBrLYRnduQozqBgDFVALJiBZFzusIxfA8Gf
LUX5gBmcmvaa8GmbVpPSqx5w3IxlWfdn7fCMXUjZYBRsXr0LMGWgNDSG78tx9B0sdRbBzDfHi+8e
4SJABw+69nQJenWZunLwmVQU1L1SechsuF2Qw/Aflg3PVc19iyw0OgFX5c5on8/MOu6mJILIMy8B
5sqg3IdS9CVlTF1LudIMqQj1CBi4umertyVKkXu6oRBLr5zlojjF8zUDuxGRVeIZcDLda6zat2rv
nNQejtMV+wzFz0RJjNZ2rhhfVbv2GBp2+zAVyx0zaQLtdYly/qMAu4B4oDKaqBwbZze2jMAvNqgA
OIBFSaucgtSTagGwA3hfQI1PmD237ZSxjfEUGhIhpSPYV1CugjpcPq5hxSvClMLJ6/XQM9f+nA0G
cTlQw8Rb71vvr+T/7ul8p7usXi145bPR2eooPLZX+Jq4HIw792QnYGNezZl28xy9Y0Imoj3do/oN
8C+SCAUWSgEto7Mtuq2x3Z+1KCHa5QpYHEvm7LewpeAesqZKx0O8HHWcQQFmLVwoiTbUU2s7CIUq
vr0UyDJT1VtIXiCEghNRTsNkXqHj6ScNtDq1dq5Th8cVNd0I9GqHmFBXk+FPTUrEyZRwN/Cn3Qud
2AGKVYrVhicfUKXBc8D5zaadPIK0CWTYag6ofyh1fWacVcaeru4WfNYBTZH5dkqCnmujpq7cFO4B
qLRCAHz9Dm3bmYidQ5vR/HBVcE13LBqBqMw9Po3iru74JbeZBvLwLJTluYEWloKYCSBitePjH9sX
zquwg79VFQozu+4x1kf14LHxpP88B2X64Gib+nZxfBa696VsTtTJpQSWBTZRdj8QZZEim6KrC1UA
u9orilZxGArPnrLUpno8l9y1dnPqZUAOuP4M/5MsrNvQL/OPQCgkjDWB4RTcROpVoxgXovz9AqyN
y/CpqxGuN9x1k6teBexad+X2QtFmVxq42ZCp5m+flnNnWpOXM6AZKyvIAKjqIjaBMYTz0xlqTZQB
+hEUfY/m59N0STuEye6RC/6DnN48YOn8JhNPYxm5wLD3usdC1mvSJhZkbEctfKdKds49MOomGrtI
42ZIGQHuoOyzTPg383BcLSrjpM9KL4nXdqm8iC7rrr7GmI3zFzBI/VI/QO28ogUmiXF51M65D1qo
56k18xRbVo8CQZOwT+qIZ329Kq+fzBW02jI/a/Pq4e/qauRr5gDPF5iG1Pu2s1o3aLxwJTM7cPTL
s89HsCCadGBdii6QujyNUiKMnE8askTYWZ+8dEseJM8Onv4WXG5zpgCunzLdtwX0maxMcYjDvhfz
HAIpWJflzd5K2G91pYk056BvDMNdR6EUnDRu5GS/8CO16P9n2QfYYNEjZixlvDcIimnSp9SJnHxn
Pj+XfuBQ33aDlPWRFY6VkW6nEafQmSQwWY8V8vyjLRaYNgXdZ0f1ZWFM9m1CqKmPptPX80vY3l6A
leeRZOLPXAgp6Kk8YPo4ylnARdMNIRAye8Cauj7kW05DnSNmmQEXwH4aTzvAbOAYqDUwofW7oX4V
8+SoiG2PiZ6/hdQ7kY8D6c4Aoue05+PEip1vadszN0hc1kBPGAJaEUp29pk8gSlEP9M2aJbPiAKM
jy0DlMO6WBnETHQGcper5kssyE1Km21XhRYbnjDMAHb4xr+QddNII3v6SuCoV+tIoD8UU4t4wZ1+
kMGlvlbHBvFwpqM5CGcnF+aq727I5N8QdbyxMTRWPMulLM0FqY6dfIVAPWmMRdQb2HLLG0TQxFEU
KMx2DtJKFlIgosZoIccz6Vpc8AgcFs/8GN1SOrEn6t7Wd/mhKjZKFG88/VKkAdHCVwjVLZI2k9WU
/0T3+hTdG1dlXkRtZqZcMxuSdoSjLebSQgDLp1p/JND4GI4Z3aaA6R09NcTqbrTsyZAIQxcMa5S1
sbHryTmH1gN4uucYCRaYJjnxChEOu04Sgz5fRRnKSALn4lgcHOOsp4ets8zBNpsQTclDrj8unCIY
IhtsVdmSyyoLmHyUOQFoKes684NIXFsVgubEIOpyABYlWwXqqXZriMAUVWXg6NxkDvbFjvHyfRmO
6Oa7zrvaa100NAc53qvEwgqYvwVPREBsQo37ovrq9iz9+Bvt8nxV4VDm2G8O7USa+WgOMNvVeRTp
QLh4TPwjl6AE8mc/f88Yea1sW230b/0OaJ5CO02XBRzAG4S5n7TBnw1sE+Y153LwgagcnGPbCXYv
PUMWv+2ujc22KIg/27AM/CwrNHkOhUK/8XhHcEe9k+TZ76Ka71VaduLhhpdTXTzxk/RsGE+zs/+p
bAD15XlC33vUMhGB/SIZD8mX5hUdJddEhb9zu3T91lAm7ldAubuSw73KVa448VS48+tp794Zw0Ky
CsVg9IbTwYyu5SOo0vSTQ4oII1L9QQyNXw980OU8eAAFSxwZLqAHRm7TQtxCzaB2Hb0woD4szVDT
YLK1l+P0UpEntDDTlqM9uhV18uF3eoAsrB9Fv/SEZ/IJ5WyOlsUzgZlfV52uwsNmx6VNVwp0VMUv
zlLJ2ZPV1B7f+amg/50YJzMZo0nWeUBuklR0NsgTd4mWVItaf4K2y5scrl04ZqXUbzwFdQEsrKo6
zc4KLZP5UsjccfMhL5DciMfKUWu0t9xjbYXVvE7y3N1NLnUbUdGx5fnwA1A/3Q80irnlK9zAMuc/
JlKzAm720oMpRSqDNaFB1Qe/VvUhrOYgUm8+KBZEWgeZc6HZL/zferhQVUzhZ1DhwkYM5VYukKhr
PkCwKFNnm9B1LOXkvfiFcCenfqm1DOAh+5vBxGmvjK0nJrvDgF0fMYlmjyUNBCw5DxrmeVK+SUc4
B8EiCm79mD0c4ba99ZQhBox2K8Z58x2jP5f6heoyY5XvKqjcgBlyTfD+J7uiftYo9UVmaboQ05tY
VOPuqtL0PNB+YFtKwHFoq/vvCE+boxPPwt01U7K5edIq7USyQty9N4JyEX4MU5fO95Lz2mGeupG8
sFShDl5YprfzXCaH+GQehcvwcz3TqK2b/m7B3OpKvRA9jfVxWVMTbkaZFwKx1aBQA7oXAV58gUeu
/FMEFEftMe8VRwFO8Afl8930f9ka5eUeywQkriaCI44rsXOWIXWO4Xpb48S8Ec8mbGf8P5K/B4+K
xRbNR/N+GsCE4s3nnBe024gtRm/dMCV6VFEjzqGSXpxyyuZfU3sjZJ0xxMtKsQIRigpBnwW5L6aZ
Sa7/mcQ9fQWve5hRDB6dqJIyO2CwCNRuuiXKEHV0CpNQ7lcTiINIlfjGSkuRHq3SXcHK4ghvje2v
4oxV0mahYSvhbDVsVwTu+k1lZbY3+mmHpTq5NQt0VTDroFs/6hCYqQWw5TOzqf0E9KMVKKxQKXUy
9O2718pRUlX6NGcJrABnzva3N3Q5+8cMrG5LoTORwn9ALbR9kV0EK2mmfBMeI1ON3apI/HUKnp0R
5sO/O5bs4/42Qwvsz4FcJf1W4GzGITmKn/uip2fl+H3TqP3aP5jNNbZk13oLdfYg5ERQu7IZ8AEv
DQsIdu/xb1F4dAKmuiEZo5YnvP5m7RyamcxkaN8BJyWnTibiBYNXsnab0pZasaT29FEzpaVvl7xa
bakbAcOnRy10sEVhcG0YTH7FuITbuPfPBGgKvEMnvjWCGH/fixATqi+Nm3w7ugR7CKy9hqjGObFO
UFip4ySdaRjIEh9XxIdLDyaRiGH3jdik/wTSTzJ0KoELUB3y8A1ws85vXM6D6dTb4QEZJwC/C+BY
QSAk8lsQXK39SQpAfZx3s06t00y8t1tcXAbqZMQBXPkHrQ2qkb7HkzgCAGectfEyGGni2kVHY3D6
Ua7YXP0MGsHWuQ7d8+aKzY9KgB2yeJKWJePwGsZIqmNr6DYGUlndm1e+q+62gfQkFSZACNDNr2Rz
UMBS14XNUiQXDSHosObP5VuuZWiqIo2FC1Rb87rUpcYWtOnZT9rTZNB6IIaMnbDlkaXCSebOUIRd
vtl4909xO64UlIgYHiBqfdnIZnFcWXG5oZtDA9kSB+hIvNPDPCWA7UMUKb4bCIoSanIgOsbBANLU
Om86NVwxCK/D+4x7W6BGDM2h8TgKrJY3Wh2SztSxn6hXycZ4+6spx9H11azv2/8zqdVgPaaddTco
3D8rn8hxvtjGbATEVFBtIa/+bOQascWgYyy8JV19+EydazzHaNLdwYKkAOj3RpoG4LAo/F5KLRb5
1WikuX16x7IWPCpMXUhtKOdNJPWGrSezjxramPvg5LBd5j7gdYH86ZPHNrjdqnSDX61uebvdWlsU
02OF2O/ryH7KqJyirpw2hcjmU/Z3jubqmfGiovsv3+nRWJNhrFIu+heQW5oZQgGZxhS8GN9G/jNz
wRFkI0luC40jWZ2P1BDJtLZxPFYDGKzq8NNhcctjG4uOQ/JSCUkn+uEeh8P5zU2iWlLmbwE9c9NX
VdPWX0STk/kGQBPehCnZlFWmDwHXCtGn8a68fDmSW4ogUKUMMne2JeXS737hxgK34JjAmAwHpa+l
9l3l+QVr2zz9ib8AK/E2P1H/03vTWItikMoJ/HXOv7F/pEPB6HNFlk1GrszYXu1T6ek7H9cODal+
NrUp8t6vSKY2czlaV9NMc4hNAioXAiltjk2bbMq8mx1fWs4KHHIa+jds4S1oAhG55iQXVxadKSII
6K8PVcSFuKeQGBmgll4idnVvPy1Ll4dmit4x2ShZ2QVntxZ/QMv6L2qe07ORJUAD+a2tqz/I6lk5
xEcG8TRTKoGhQvwBmr7XorCAoXWmYjar2vo5NNEpOQur8yK7uA9FlIBSHemrKX8g5ZmqvvmBAU1h
luCDzxl5K8D55+yGqLuWi+jFl48za5NanpZgZRFRoUj00QAoxYldqeqaCDTukylQqCyjvt1vvs7/
cs5tPVzURoCrzAv3Qdbzg4xtQvepjjByYWHOvNH99YXc9uq6PbNaBFNJnLPWM+9ZBkfvOa9xKjkP
gsJWTK7Bg1BuA/nFqjeWEv/SPzHeKShwzGdVcK/8MKlaOOpb1+NHwr/gqMofB9QstzrWqIfQocRh
MkJzu3i69wlFW+CcdIjQSAaxZwVRYNXjSVoFda2ymrAKXx4v+HdxQOKyBNyz2HJ4HVUPCOyHbNe1
arKUXH8oGHhI4+xB3Tnc8SoT/unrsJJags5ZJlQ0qWmqNbzBieMgsENhTLeB2norTBSIGhUrvMia
TANnBD2Bwj08Va/aPaht2Txt5AIGfIoithuFSVWAQ1gd3xNHvTA6mP5TvD0+k78IYP+USDsWDfT/
tZb+Ho073riD1pxh3uHmLqgCwBTWBs0YCizaSMgvnfc7MoktYKXfizjmrYRVgGbZ46mV/WSsR0dz
rWeuKhfiRZUEg2lavq0MvKi4OmfBmunwkCWyFDWHBasKBpVdLr0mA5yj/7Omw5U5wGOjJFKILlrk
Fix0c7N0MFHfbsLQJ5aN1HCPVFSyeuwLGzn/TzMaTDEm+dWbUcRIE7gXzE5IV9iGoCzzUN1q/yAU
rQ2V05rtVG7Vij8vMINzhf9HonFefeeISKS/NktPsfjBGq6+u8Wamcv0vTul2upbovsGLQF0wgq0
Lac8oaqciLYOqNesOqe6fcmMBx/Cd0UuI5A1ISs6q1xWxY6UZH4IbUlf278SYmBCuMsvaW0Qx9b9
YOvJPEnxtk7mc5xyLN2sOvf4Vq/TM2UVNmskrZT1OrQ8A4qLmAb5f/KmDwYZGgddaeK4rENIfzny
bTfKJKnpazYWwJltB20R43xyvOV5lTMyExFrrSwm4uyOURieo3pTcRvm4IeYIWkc91+OZEoIEGVQ
rB9hiNnm27sRKdgVGOqsEApuThc40u7toIaEhQUIj6WIZmq4kqdG80fHF90ymNqv/VbHXqY0dk67
9EUe9hChqMlgk/AITRD/hoiSJ2Z2bkt5fpEXq17Dquz8bvdRbSA5aEUTxIcSQGaqFcEOTm0L4Okj
7+uQotS6HIEv7XrF0U7FATw8N7+LbZycVCRrRB4NUT7XXVaO0azmEcX7J1WgwaczMgTEiBfN0yKi
CqxrWpLrSDTqzeIBUy2BpWAsOy0HAOeRN+lhZZqFEsAQyc1eshSZPWOvqPRD+ivnvdU7ESRbw/6W
18QloUFf7w0jViv43VH/lEbsFlGWehWXmwBJGfx7Grc42P4ZlaoQRSeskgp02E71+xUyOAvD1Pgd
XMYFSic8kneBAXGRqlVBnAjjkb3g6WOkmE9ikUUeT8iO4TFmieFQucEwJbPXatR5jrfeDYNNiNow
3O9g49Om/8hGo7Fwg6q/x7lx/SortXDt4g7fYxYl20EfgxBG1Lr2PmQQfNqckn7xK/0s5Mu7eIFz
vhmHWbc3XKOiBVDZRS2ajvJvvzxIs+FqtxQf1oJ4P6Lb+iyxjQ2QLAnDLMWvWC25ygIKbil6khlA
pjmuASgfQZBV3gvAY0sBrR3ufE8QthTiANdoMFlymXShvu1MC+X8yxua0zZC2zz/ixDzdNqEF6GQ
puN+3F81FOJLKapU2JByOljfvf1CNT7N3KKg9Pgee/Bq3JDA5u7cXbKbYyfbDhf+nVv2v6J9gGgV
oXxrpII7asGX+vsErzjhdxVbs2aA5ZYyNvr923Bn+aK53rMpb6bZtGsvxpymAdfBlOgrf6tgpRrC
bf83eqiTg53XnsVGRg2NkugJv3cY2itA6YOed89vxcWobDm5qsG0fp8UIt4vd9J8TARh/SNWkFqn
Da3gHOKCsLVxkSbpoTDrwT5Myks4CcVowNhpWuHuzo9GkShgv6KuVNNE+8fblD9DwwxFxbpViVdB
s/OtfLYkF9eq6nmThvVS1ahP+vYVy1YKqRB4IwGAAQvmuwruFp2A4Ww8j2du/01zeSirpIjnJrps
1J2UrKYc7k5Z1KP+Gbp3AbCNcaI9BzTVA/ommLeNd1M3pr4Vf8LvRDcRS0wSUJMvlGgn/Rp6iD1o
EjQGj8LWqgZ+Jb53RVl3cY4l4FG6mp3lnThd3/s9gazmhJEqo1emlKWxZ96ob0WkXVQBLGd0mSdb
prqc/Cr0fsTbPUOa43qy7caOKhxaar8Of2I6qPIbdbDtIv3XhAigcV4Nf9UTdh1DbsCI2kQu9nJV
2eZcFSVxJATLYYMLzszZhRiR3Gj2A+LaHabBsugvX1is3Aq0D3h09iiy2a2bpCnlhCE2Kw4HjbXC
wtID0ymB+WDwGSj7mcx2us21JPSZpWXM6eIGiyaEzYstAlli+ZgE7i4+B4yMTebcYWVdTyek1E9h
MJ3YyIQsDD/XVdVlYFzlLKJpidC4wUqffqA217jfW8Pu+DUAITJAviLl5ctzVu2IiZJok9hJcrsr
W0N1oOx/haRK1pRiyvGpAlzY1a7vmVjAdAgS4Twc7s8so/1KLXF9vZ9oGzd85B6p66DCC9kYWtAu
dJeG0iOajvTEfJeTKk7E2KYeX14lKEkTT1XbP8G4MrRKjTm4acve/v0W1OnRxLCuwN9hLBHmO1FL
CIBlii2SNisY6B4n7VmFVQ5warZdQkL3YeQAGkWAz+hEmiWNOq2wailOG8YDzx/R2Wn/nx4qt2LG
4EfLmjhMCBJLDMq3gtCigh3E8TQeZYCOp+mnNfMhF/t56BHuABcSDBSk8BZRVnLGHxKzRcIUw9Sq
oCK9HTv6TjwznMrs/Qyhuti+huHFGXrCqklYCP24rMzHyOFePhgwe3N59jdlrKL4rbXN5KKrrs4d
6DPC0JQ9Db0NsNoBeJJ2CykXbqfEUnf5jifOxaytPtMKWelJppdGRrGOetMtO958AMIeZsQwSqWW
1b61HVeNoRNMEh9dsB+XYEKeUXI02yB6RpI34S1F+cadCxrv+0/BA+Ajzgu3I475e9c89d/nogNK
noFKx4o6kieq31NuBTvvIM9ha+/jMplqhAce8Vvndj7g1zQo/lZnmPy9TGPFo6ONXOSt/m57JgnU
ScFGe4DI7PN4A/cYT9N0H8A96WNsya+1qT6SoT9aK2bYCfZ6S4KDpMcKckEmxAmQSAOyYCvOezLe
37nkixvuatREm/G26C7sXqmmZpEIIlXFU/4yVZHhAJ+vN6cVxS3eAo7G6Z3P4uov5emuBntfdaCw
Z6JsG95KUfZCk9Y28tQShqecKoQQlOq++EVAXUKdwXNhxIH9kjpujHSrAJdDKRGyl4ryhw6jcfJB
5dbqInWLJAxsgW+lQQIWr41C4tiOS9V50yrzaP64vH404Of75nim+Woq2HWdrnHCyZGeDkXG0ru/
4x4CD4ZbRAQ+cOHd27kcwzPJ1n2xPzll7b3o8hRAZktd3Mt7/dGLSijWNmBR7zCTPfqUx5WLIhX8
Olxcff3zoRGeAp5cPJbN5iem9cNSR/5UJBb+reI98lFIYrmYs8dH9JjN4zXlxLdteAjS+m0qc1G+
QyI14dLr9lCJAJdye+yynxLztE6kJjW5QCfyweOYDrNtEFqghM2SD9JQczmo4jwDw/jCL5neY1lT
8aPp7SZuCWe/6GLqS/GEXwP1Irfbso71Q5NnG9ApzOqmqhZpWIuElzn7/MetBR9jXlqtPfR+4FnE
ikho0/CC7ENgn5nZOAK6Vy6DKMK+DwKaaGQiGmKiAVpgJJoaVnJPWl9pvyJnCw9isF/gF9dQ/gqU
7e58VE0y6PLVzHAf9OIL7feFNchsvSPB9FF60GCAvqwK+yrbT5YIaXC3Z2+BOH4I5XEEVYFO+I2r
sEbjx9ihUbFB05BSO60+OFHtuwwzfGO92tJ1bsOqMC52l9EMwws8iPmoZTUCp2jPp1OGQKv1HWVG
1uHKa2lmrqHiE3sQxjiRN4yP5kmLbDNgN/WbLg/fK/KPDUw7qW0zmIrTcmWNraPE6oAZb3DetTfE
H6LZGl9Lt2Qgl4iuhyNzOOjMraNov00OMpZQau63eREJutxFye0EGlM6N5uo8ih/5n3klRMOZ73u
dco0Ule0NobeIEFpumoZFQmWOTaqZCpofcsPjlGdJeo9Ht2oaZg5hBf6mOdId0otI3zzZq1AlK6H
8IRgYrr6k1r8Cno9h0OWAApeK/mc2XzvxRKs37+Ai7y7tiU/5la2Kq0hK/wv89aWdwuILcl3Ezw+
W1javvkyVsDWBMoKKeadmcA+OY72ByH2vvA2xzFYIZ2/PcQB21grKKlRgTTRbxyv77oTfRSl3kFh
WfsECIx54Ac98RMoOTA1jAz46TcdF9kG20Mu6pArqohzbLA1XO801m+rXG7Rk5UqDIL5fH8uV7St
HujEZEpDfjdJhK4ZFE66/RwPEAEqwZ9jbFDIxXl4I4GWPERcicrWWe84CfOSn2/CxAoJ/5C7tKFE
nrNFiZkw2nmdf3fA31YhYK9RO8h59y9jKTPFiVbKSQTxCJDzPTmgkoNBJDk3TeuOmLVqifiWUY+r
SH97iQmFaS+ItJC2QI5kTFWsT3225+CVMv12x6dxKFPMheEz6sisfnaSJ8XwSiUUtW3WRSxqgGV8
B3STVOgA60lykkSYOEZRumQeeJiNr5zwB9NQNpw4Ga+Lvvm9oOWfXprl74plNkgHPBit69v9trUI
d+j7bS4S6aDi34TlLGuIdiB460lKtfxMazBV8oV9N4YoT3SyOETh6yLRwxPDuNI/1VdE3AR8v7sl
BnBxPxgPznZ+LMYjl7qVFz3t3E73LmoMNvLz1j+GkOlka1bjWea1TzYtAcgeo2B2djXp1+TNySOk
RSNKtELJFsN3IVEIH0IAC+utGi9o1XQDm4IVLNeT6u4ZRQcw6dNi/BsBobr0Kl6nWWBh+apMF7+i
EtgvrCOZJS3Rl/c8nGvXdeYWwiEIlwAwy8qYbNzAjS7moNoajO/49zPkdL88U70LFdhu+CHrFKK5
yezlEangnlM43IVPCslMluQjEKL5emuDKXLeqUilSDHDRVo2YDwln0eK1na4O69vIAzB6onDtvu+
oU77pNWgQjMhOwGzOtRJcrYP3zt27OnLvz19kpYKMmY0HFrWaRzLSwXJC9nmPKLJqA/WADpcXKBH
LsT7oM7akbBEfNIRCFZqiskbMXrrLuANuey6Yqe39eG9dxa65s4WLli/zLeyToKENIeJB42lxUgE
mJ3DFK6Xmclsv2ukHDftE2s/sbWPB7Lb4Ijy5/a835iVQoj/9KMoFhDt56cWI0j1KmjKfOWJpaEo
pEFjI0SJ2TXMY4/6/zy8Tr7BuEiJZjTc3baVVuaYiOHZWEBW1QWW+fo8bKNqApsLXj0CH1Uz7Zi9
3Ssike8OVD3uZSOCKBDiw8siSXvSPYQB+9oZP5S/dSlO690rsXD/0du+b7Y7a7NNLGonWdWI70vK
OTueunD/vuYbnkxULW821JUUH0NfprCV/D15j5T7avknnRRLb7PdC7HN8q5Mke4aktSwpCpcofdA
v5yTnks0X0Z+/KiF+nmhx0Bm13cVOSP1cdHLsCdr9e6raWarB6EQu2D9/Y8JAPvwf7kKKtIoe1vn
CFAvL4iZP9ytEs5jNv6TVT8bI9Rl0/NVCt4zEied8CLrU1rt4AvgVsxV66jM1JpFX3q4KDHA0TiS
rMwGcB4wgBOUTPsjhfIaGY0V2LTrHPoAmWJAO/EGsBAAS4VQ8DAq3P1+hSYnBvWToh8yPRoNDMiA
OypoVOgiisziRnj1ke8NC8nujGz08SoKjoJmDdbq/DcveQ2Lz/3KTMWGGoT90aCyOMLtXDVQ3hUB
/D/gw9aznrrXPmdumLFDTL4P6CJaeQIjRBs/FdsFgru20O11Nqu1lSQdM3sFbqh5clwyhhJgpwYw
39riaLOLvzk1vTDidO0mqgFnVFcZa7eLRyTlxOe+CV3gt20hzKWcHT7aUbiTUf3Ys7p2vZtX9Dip
Zw/2ydO3WAlmZRwA/aP/YceShN9wilOq3jHOnOH4T0P+EW/tT2DDWsRbYk3U+rk77BZFlr6f3l83
GTLvy+2vqZqRAEVzGw/tFlq5c7FDwdm5eUjtzF1Z/Y3d6AqkmHlSuU9SrbUZ7sYOqmE+M5Fs3MRb
bWnZUiZWgCRVt9XHpv5nCSaNapJtvT7vEaJoDDCn0qFAC+OP9xqljwariCOq4di642fN9c1sxh4h
ym2MAw21TeDBHJKT9/Z8gCAs0gx/Pj+pcWI+/pBhHgJwQYpi/Zr0p0jCJzHz3OWbN+MkLzSPcKwP
i2bYLji0s+XIr9o/0VO5ZGLbcaQn0bOBJRFAPc88jot81eUTZ0sdt4W6ovtLXjTI/Q7MPJLA7ISp
QaIAe3ffTIoSiHEpyQ84cqCqSA4Q+kZ5791mkDzKflZnT7x9IlBRVb2Z8sxrlILFjDfQMSPXeaKu
Jl8pbvrYtsCx7PlFwHdYzichDCRsJw369LGbMS5tPxC76V/yI1y81U1iWBgLK9cyaLczYfHH5CIk
weULPGaMEH04fTUaUrrnAA9lX8L30i0PUwK1Im2bO2XE3V6X53IfrUckOE3VmekM+jGHMYLgO+rp
OwSRLK4MkRe+iipFF4uYTCXrFRx2rlPSGZ47bEDfjiVy4mSiM7DzTh0nFaVu1stQoFSDPqv/6wpf
FntNCmfXHJFFvrKbRIDYCN9jZpPPCpugToebJmTpNiUfvmgUrNqQfeKnfQ1wlUDc4UmCvo+RSP/6
EAhYWpWU/hpyqZZC6oHOw8b97YazZ4WlgCcaiqeC/5BQdx0Zf8VLy3TkYAs95Tm4LBC7ekPtpOk8
lf8i/nEtT+pMiR1tWJqEsZJb9RHfG631KsYZAIw7xl4wDtMvQXICH8Ntepc0LHMMOzTshHaezUHL
llLh3Fz/5iWe3q9nWlNUs56XUqxgV/NkPkxcs5AWIbIbaUJCO8hXQuzYlmJ9/q789qZ0VdO+1D02
uDt+yrIeuVHmKWDmsoxnecJLPtP1sWTwC9aZb8BTNFi6lqHASZgDk8MUv9e6uVVEb4LAoBOCqpL7
De/JXdtAboVwotQ3cnZex9T1jR0NViLqT43Kt1YYub1zccCbeO7Cpihv5YDprFqsGd363uMabUaM
S/QXvabBIWjgKuJzXFN0BvXY7o64aCfsgm1HCZSImxPtpYiXgkpGroNcMoBGEXaW4zAk7FUrWzbF
w9Cvpt4AfoCkX1ZmrrugGdbgHuxlRlTAtNo9wj+7oC2mROMwXJkq6Qxs2PMskJZOjOkg0gLTXxVd
tH8sfu4nnEb2kVp4sPA43lyc/K+bd6bSVNa59RJNc9MGc9wYMlEEYor5LTkvgSsWSHKhq5FRY3+W
nc9tHPKShvbLv9VsHQb1XRDpLIBJ6MEOInzKqYjWfz3Ew+i9oDX6S56W5QZDuC0pdztBognn91d1
8c8VZwJw3wLSo+5JGYff+AI4iYtbRp23YALBWrH6lCojHaYRwogdkNWC5YCgeR2BiwLZAkZMjAa3
WxsPa/gSL8FaYtTkt0ptBUqeZrM3u2WpR8N05xkRm28rpIzdvQOOv/NJnTzPzWTl+g8lSRiMCA7x
vrHXsz3qZfJf8MzQ4MXBQv+cjSebG4Twmh5zWcUPmf/L+FeAW6m+vDpvybOZoYKveeHfA2PYwH3U
QtLU5c4rKRwpLUa4zE/ScD+0qvnkCYOftMat8mxC5iBKytu+mtq+9Yhs0LA8wt3Dho3sTfGixwqw
eu/NDw1NFjIWBlHucAm6/FLiD1C21tcODEU+/o7/6nAejJ3dECmAudsz5nyxo5d9wnsYLpaiuFfB
XFWhUBF6r0cYCpfRnJt731y+F6vZa7X3oX7h26/OhexTqabs+BV5rmFLeTdilt0L2yovQKDphJhT
MIxStWd8yS8CqofS1Jzg3RvZoys5GfVHCwi3AiuA1bzgAccpNXhexBlJN+jOeB+ii5pDjuMPcPN0
zsLW3pjqcX8BpLH2Gq08D1aMMkeffinliaiXWpzeD+XFQp2kiwwU/bIRh72iKUTA9s+dARLTkdxE
+fmfWtn7JucxFs9EDejqHEePqk7EblVRtXy7roJxeab4y/o3wuJDmp2hYGdBY5w9PMd7FYHUzmNo
NOZQoS6mPRTScD2hxbeRn0ht+iaSjHRRG2IOylFHe8i+UZheXKA/vGMnYJFKmjYu5J92w25OTxZB
twcE0F9e1bAROp8WFfS/xCUlaUYUmEEbPLEikneorNeg0Q4ARPusUNVZ0xZDfkWnCbHLWZ0m/8zL
Kus/H0VKWBtXYTXOqNSgWI/qjxojLww4iVgtr2oLrtoR6WFWnjs2UK7Wm0irvdAos8bZ6rpTMa7r
VTyYz6pGOk+YrgN8i77MncBKW2N/2+UzIMIh0myxw6gHaUzOcwgPcmV6rRcrDC9C+SmEvkZXbogj
/lpcA8DuBy4D5kzupRl39C+6lGMrsgj9MYqC6eXwCVzyA8gVlpSzvgi9Q8aPhB4HpiQI2soH4qLS
QWE48ue4HMvBJy20UtfF5GK4JjP+SIiS///sCFWePGLR5UZ2EaQYaka1Mp8eHmh3VYwJaUmZPkWv
tMXi60forMJnvXdZyIgR5MRd5Ur5cmBi+lPiLBZ1w2m6xF/cvtRCdaEBvU57Qwr5lXPGD2Mk/NkE
XTAQgDVEN0jqUuaie0Nw52hYEFaTfD/dm9pLk9Ead7JFh33NtOPC29BpfP0osazugxhmPzdvRrTk
J/0S7mfMW1NNu4m3AYAHkhjxtfIlQWHE/jcgzjok0IqUHQDVCAPX4nbaKPTRbcVn11o7IP0wwxcV
fDIRpq+0pLvc45fa/ur93XySHk3KvfSHlKXbE0SnZu1QaNqUrageKVYfbozizYwJ7eeLuT9VeN7y
HInX7GCZrXksUiM0KMFI3i4uW7Q8o+ysDJq3qUYczhrt5R7oDHIu0oN19VAJSydDEmArPLrBQzj7
IvFcq7CzOZ6Uj6K4L8JJeXIMOWG1KcRD5osIqNNb19x+vmEtdcEySZLFhY/Amt/kFxwQqf4A9Q82
B0QExk4VZJOEPXpOZkDNipdUiK5fqJozVYeTJQa/8Afdm6r1rLo/xMLkJ/OoLUC5HXiVNwBsTOOh
p23HhjoPMzwBIFjWoh/PE6HabDaEVMJYBYdNCXp9WQwooTMLAK7HmYBgrTHeasIqfCiYr3UF3/he
tNTBD1PfFIYVpFeXbcIeTzXB+kJlOsX/Ghnps9jwYqgmgc6z5Hv3qVYE5lytZtTzIc/EtJE5yEqA
1sBWyPXvLXyNT+ftBFVcA5MSgmojNwbAOqEkrt+r7fLI+xc00QAY8tICPv+kl0D7SqOB3aqIZSok
wTJzoYCTAqOfqqo43kddtA7O94uT24Fl8k1gq2eWchbl4SH/ZDstYX58LZ7bBrE+rylOK69KA8bl
Gj0q/OIjKJ7M/iRRtfi7PI696uPlpWDqXu5xph8IzGHzFxbYEVzom8N4F87yGtFGCONF38fFdcoZ
wogzBUoKJWx/OkD60lAV4AoS72713ii5TcJjviZ3C/iWp/h7PaxYF1ZV7foaB0yi7yGmx4fcG/q/
PaxLva4Hl2tAHaojgBsa5OI0eJ3NQ0xTNFDSXp6yHSNpMC8oVMzBRHq1mLOFH0dDfubdJ0G6yFvM
Ee4KZ4kyQuEIuMV0Zmh2izSyIdApQJiFXVHUtixYxcGuktzj6Zsg6JUDOTj+ZmHZXoZ3SA8MmpcD
3Upf2WA5LY6sTlzXFuzoGBjCMofZIR/rZ7u+abRwO12eOC4JTQvLxQ1GQzj9eE2Pv3H+c6VLl5QG
U5N4M/NxvFt2ek6/PyvqSxlvLhyQ6BxW+o1vN19k9m/BnG0hclY2LZtgywKi92EPNNQLwFagAlod
/aWVL6qDInzSgZzHDA1xGX/Z+ZZKYREtAlDyZcmePMEVlkyrGBbsjLdqzY6QGe5Huw7yWAWb+YBD
YeyFZZGKekwQTFdXVak6ao5jT0e+L8i+ycn5pjyPYec7UHOyTHW2AwihxUBirPHlh91rCk2y7d7N
70p8MfTZZtxLChJUHQI5EFMKjhScEsShQXWXOleGYfVU9EeP7BNf5PgS+4KYjCSPuXotGC2FyTES
tzpn/1+r2IjXmJyMFelDIsZszRtiOoBWWRWUyXOh3gpWVRiUopgwdZh0p/+gxM5TFtkY3I0RVBGR
KNRV82oOekp5Z50R3z8nY+aLD5uc/ROqEzXTTt7rf0ZMe1UgSK2yYxOltNVqIG9G+9nN7xJJ/fUr
AJRMxGzt3Ta3Lx9tgmHsPZBqTc4k/yBL5TXs9KFulTYquMCyf9aylNIo/mxwZCw+cX7qklPsK6Dh
EpplrADP4Xm+APx/rIxPU8seyCqx3qlWzPw50I7/v0jTygmfvZ0SanL6bzMiylphmPT6GQ6sHqCI
hQGLO9Qq49P/D1w3bynoK1AgMWxqC15C0GbEHzJGsy9twZdBvOB/yeLOZXWrpRehaNl3z4BsFYBh
pAj1gUU44BtMi4bLsbRoM/t1Hcm8n2Bivvuez+pyWsWnmT0K8GlZYCPCr2T1ZlZTj+CVJQI9ibUK
vax+jUG6okkfNdayspr/fjTlE0ePbR2gpVvYAbHcZBrKPGYEuqyF69HG/53uUxv9D3qI4e/LYgOk
XWof+oMl1SrzHmBUYC+2VO2FJVEluz9O40+Iozcrs8VDWz4Y6JEbU/fh3dgy5SJw0xQS+UQvh4iY
UdqRVzxN/JgOhLAq5YI2wRDdqFLgOC2Q36wda5ckJ1DvmQqgVlWInxra685y77AEuKge2UlEIcxF
75f1+CEnWnGsHsa4UFAo/WKx+R4/722eGKNJ+66eK0ZtvctLpPQDJ0JSGh+QtI7xdnCi6NFqxXB9
Qtclw4dvJSdAsvbpYy8PIqb0eDhNsdvIYTOvWuqEAC+4mtWHWWk2nT5OYHQy3beSP11m+WY8kcA5
DjtuqNwxdTTBUbK7f6A4jrSQ8wBrozrCRAlcB1FWAyaevetg7v3vlbQhvkHsWwHAJ+hvRfjkpl5G
2XaJXgdS25LEP5gC0DSjR5rBZAUPEorM9Z0Q6nMAbEzuN2X+Y28qGxKM6SaqY6QXJDPXKnKqHyJ0
tKX4PnYgfLUsPmKUgBxVRdoq24Vhigx9BfYuG1QVYJeuopq9HgaCpFGJcIOa1nKUVEYn82PkjWsa
ungP7b1Ht4+JjUoF/R6iNBQEIkwU204djkHZ9mpDjTEepf1LC8eq0gotZveSeggASWz8ANpVObjs
cW6B+R0WgaJj79vuBtJ7afHP9glIWrX08IZ8Z4mGzHfUi95ZNJY+Z+DpUO0sTx0SWt1DrQPhltRs
xwbqxFjqenf9SMUcClN53HOTAuxX6QDdKfhU/3Or1hgM2+raqO0QFJZJnXoHq3XKrbuSRNAHER+1
58PHnPBPGrHPnysjB2IBjSxEi0lgeQG8sOrrvsLk8XPGXzhfdR3FHoMFbBn6ezEC0eGwjZouAocZ
2rYmwWXl7BOnGtmC2fLo3rEtWyWomVja4AFnVpEaygbpGOrFdaDKGdmCkPnYsoK5bEmyXIOtJoz2
mlu1mfQRG9Ffv1PMsq5Mok8heo3d8rXF1z193mMqkV+jNfq62qMhPCwMnRqbiGHaiVy8JZpZG2fk
euB1ktT4MqWE54gO2ChkDCeTNNFiuSJhM0jYqPF/2PmggzuoYl40zgd9dIU/um17I5I3xTIQqENb
C/pP7pujyQMWCz9v0khYkXnJANZP77h48Ro9fjKx+u3PqcxldOEGqOL3E//ppWbo9UOp/DzwZQ7e
l7V5hktUCPyO7sTTkxoVE0eGWoLg0/DZVgNxfI4Q+T2lcsGAa6pFjnCL7doySMz34GpcwcTshseF
l5Gmkavtc/KBtPKcG/oxO7uDvpi5lzEXByzsZ/IlqIjNymErOXnkv59FSe//mP0Mls2H6hM51OLu
gvubOVbidVmcNRFoQXgqmZIxR55PINWApJEi8PsR6wUNkHx6Nh19mZGfhcbUFgQWcDxRDYSLfHWS
3sma7fcxew3fqC6VHkxh161+SMa4udOXW+I9f8lkUgIUxNRzcTWfhkCL5tUCTxmm7nuYzX5IQaR+
123fEnz96/d0tee9SmBtJnTcaOWJA1897Rjc2mSLgmy+4/f0Q+YIWitCOgXf5m6KYXROjzbrbA2A
jlRLElJ1TkxffWCREY76wTuObrkrqF+bgI9eRJIsaOsoIpwJ9vLpcAqyV9D0z02/piVJhWrD54NB
mgouJdMLemY658lqUjih/YfjOubQtjNGzliov5FSQh5vDcT9an04NG72bizUK78nq/61oYZ0sY7T
EUYumTMCLYjUkkxvuv/1siQVk8nEhCzBFSTlaZJxTr9skCShFdVavPJu+Y7aZxOwsvXIi5QfmDfm
jx5qji2x1GkMWcYPKB6dX8Sbya/oTt8RN9ovbqppP9wqWLF2bEXsXGaMMQovq8CwMAdXF0q+BP3Q
kQMICputuN+hi/ZKLnglCfqW/pDdvruGtFCzMU/+lSeVfe/YYBmsTeMubELsjz7tXKw89CEJwTmb
aUe9lOz6n9XKW5qleuEWeFEFnNOPIXrXkSljbwzfcd9oHGGgoOYkxHTiaGZHFv43MR6R1aDXtRcU
N0wqpfaEl2m75CPwYoNZPvy49/f5dPRbZT66nlRnop8k9mn4od8GhtO5kRgzn+sYZVG+EY/vJEET
Jk4A7IzOcVpyyGw5zUsU4ZVjybVmHysycAt5+aPMmiblhRDnaKa7YAW3Cvk8GY2YIq1eri27LFb/
bWLdY2x99MwfpWqQz2vera3XBvy+9U32DBVIjRW+SfCu2y5ZPx0EI7SDpYHvMokTLXcUhT3anJ4B
f7W720FDBVlAd3+82L0tNnWu5rF0IXnVThj+H6074e4iI5CpIyLRY84ZCAhDcpYReQV0K8cx2H2T
b6hVbTZtff7waWhtn+ErUCDTsDf8ptamCRL8JtJcEoNQkcEvcnqjluduz9BeSCnb6oNabkW6o/yM
2B8UDE4DkZ4L0LRfqF4sbPCb1F9BhK7idN1gwin4neNu1ybcKDNXStP7BPHUB2KHy7lQxQ6W0ort
yJYMZZo3d3I+ji0pVx5wuWGmW5rNi508vGAK40K9J2lfJ3S/2UYHViLOYt+2W/LCh3bM7dZOltGA
sPw0sMkorqcwoMg0GTirn4O6/4kLvQ91uXHrczBLOuZcnzCO9uNIY3ke34ajTJvopDeRopMLmr/i
6hYw7rEltD3ULBOJsSqq3NMC1mmkgi0mG50RQ6b1Sw0G3Zk2CmlgpckqDVoE2wScYpGzREEHaPuS
MU045AkryxRYRqW7+zrIL0heZlhD9IN+I+MHgQFJHAv9MHstvw7tpi10n/20MuXrD32DQyuo7X/9
rlB4v9GKIc6yvTp0wDasXYJwwQY6MxcrSwOHeKsl+zbBBU908PYRPRcNdARc4m++Nt9xuM1jpp2B
3jsy/Vkd54Mr0i8+E4pUoAD74EsKazDXKZ0pT6rs4502T4wT3VyG0WUSiqlIktrcd2ttt7iNXdia
OVazTMPOKjWBam7kE41/kCBLZXVZjZ1rdtVNDoHUVhx0NAYkPUnfsCkENRPlHIW2jYTvfm5Uzlht
Et3tboYTF5ukCk1hbP8WnqOgKlrQAneYcEVIp4knYhSCjTH+JYQhQIuFBtwLzakig/t6kBaiIzad
Y+vyf3s6XxG1ZQLy/wDdz2ynOQoExmjJUKYchtRm32xqby38GAL0zdEXy2qENYzwpAQ/O776ttTt
TDAzQGPeXpL6MSRfG0quwd0ffc/AFtgM7qECYTkYnjBjEFEhd/kB5de5Rd5KMcYuLl9Jf8a7QWb8
+f8ys5EW17KsOiOMcWEFedDF2JpF7pWWFt5zz4vPKcPWFEK2nvPnyPVB3S1j2/JPRYHDfyW/h32Z
+yKgoFb/TPCmddfGbfR07/dTff9MIDIOYTbvltJWn33zNlW1pgbKSpzJEPZINOFOOvrPmqhvuR0I
TvMf12K3Lo6dSaFmDNDef7d5qa9B8mkmN3or2HPV2A58HQwgrg0h40nKG7pvoeM7ZmSxi2mo7y8R
j1a8TW4VxFSmADiilYDJiH/Cg6dJscMkb/tbnVrbXfpulMVDrKhlcZxS6Hb87GbZbYuI1roBBdfK
pl8HBRUf3N2csM8HYKP6C+aZiYZl+3TuGviB1P5jdyaBN+PZPOZijIuZysbgy+GsUg28t4FmUPCr
v9lQ+ZKGYfDNkwPSZuq122ulNTf6ZyZfbXxw1bBVyJfV7j/2s4AYeK0kRCdTGm1CkrXitr381f3O
abX3djhocREoo11vo8e4yZVrhkOQVThG6l6fcJxycidXGiE8SRi9+eFGSjECkrh1Xx2A3PShduB+
50X3+Lk1BlbCZO/8XbAy+sI4Kwuau5pOm3CiI5DPNfuoEb5x71KWqJhAsUwJlObvHTZ2ZlccvPKp
PgkYCjjj574o2KCILC7cx/rRd/3jc3ouTuKgOxYxWLWpc9SQlAwMHbfKqVBbZaAekDqzkwYj2vbF
GXQ5hI277ZW3/qWQ0lkShJjahE9+FyJ1vi+G8uUXjQNYwSPnuRkqCGl2GPiiuw9W0Pwvw9VkRo3I
Bd7dL4fyoKHmfqMdzhgsqqfYlmoNq2D5zlPrFh8p196EzsJKOietdULE+XEqW7u3f6+8t8WNqpT5
Zo9/lgtEf1iknPlhJHzI4P71SyF6fAlZq0GK558tsBIjZN2uYpMSefs/Ue1EkFOFI/RocwQqf/Fv
pHG6nNvQHZFYb8dK26DgM8qs7ROE+Kk3uRLEC9JoJSetAg7ATtF/Zq+HjqlwGnFAhDHOXk9Ao98M
cNHWMx7umFWE2yJbaGr/F5E9u1ixD1uYJcrb63KamwDGKmWFZg5SpiPTsLDW6+rw283+0KbWsCEl
LwY8iFG/iFeXN55n66dzdFa3f9XEN4X5JsR3XxiEq6nib6cIGQogjXsyBKdoe7vJk2+hudWLDXY9
Cfz39JjB3zpZ0jCU+pEMCBZAY2WD5aOyseKJGMe1YNj9RfQWQX/8CCRw0yKJdLE0cQ0fAsMuLa/f
9j6BsdJubjEaG3ZapwxNgbah8f4Q+C/4oGbMmlvnzO4F7uApCCW+euUxBhT9kBij817Uy1Mm/0fm
ICAym84dpKY7OHmrEhWEnGLAoiRa+7TtALxZxgZ2cU2mIXgZ2Mt4JcFc0JuLZB3QHnpDgYBW7Wjb
wK72vWXmt5dSdZIr72M6ra03WuT6iPs8qPfkozxxl9fqPCfb65xXqvIRhlmhMpbD8ref+5PQ94H3
a83WG2A8kr9SMq7Tmtu/84JGbZqZzHc0PxTZpHmXRPn+M0WgfyazDPCd0RPejM++mySEU3mD2Vhq
T1dAzHRG6RS61h/VL/aQAoVOStp8icqMsJg5hftYn3KwgaqGvlnGBh+Co4aDM+JoyyJfCTaC7ASw
fH5zILT32b5MUSgfMsglXKqd/zSypnZL3DADg0b7eMoE0zNmmNgDs268h6CYgp+J8Tessy0/iC9Q
5oiS7PPk9nAuqymHbdBTcaKyGwFLg68UewSGs4lRq3gx1FThdyrrVh+3WgqCl+3WB8JvB2WzEhMg
GUI6qI9qt7e8tmO6Lafa5Z+eDF2XDvO9Too8ZQZScAv9JHub3UJhyD4QWu9S5Uj0fiJlWl8b4FJj
s+4YVmXcBFuHE4sW3FHZRfytp9x0xrtoEfUjN4fW0ICp7+ynAJANxRmWeJ1dotyQTFU0AcWvAW1Q
5IC2LXDNfA/+0zhNQNI+K+KbnOj/kYAiksd59KgiwXh5YvJ3INvdT/7G+mDo/0RHT2an/SsZpTnm
zlzsgLBAb6JB6KMt3ehJvbEli9kH1QD/+Y/Ti64yEA8eFpRtwuHOBCSW16PIw/sARLwmK+tl3MGn
WLzykD+WmjBr51SbU49xHTgbbzIDOzuq0IUPRX5bMVywtuL7SWIxsP17JpMXImCtte2IFDU343GH
Mvo2mxz7rS0IvFS/D8QVr765Xmd0vJBIplZYPfb7UnacL6TyLhZypgvF1zXdq8rTSA0u3JSwGwSJ
3S1zdbK4uUyotH2VhOyHI9xg6z9G4Spj7ICCVBpZSKg5n4wukSwPQAsAQI/bFfW2ptGaFni/YHo3
njfyA0umfJRgxnRVDTe+KRlcHihM/572D8aYkg4zWkwIqRSQMQ7shMnWAt9tP1MzxP0SWPKp6lFE
94NlFa4BgDYzCxGF77RjKM1TEDashD7xowneBzgGyY3bUaGmXNPEFYY0U7bnhm1IiJpVb/LQZ4La
0Z+xM2KYUNygjNe5AQpPO+sApvlwS8QYVunjL1UlzSpS5x09YR79jD6OP4ux1iqWyneOYFp4w7xc
QeKRkVcNglHPlTJ9R+TuJliqR0Z/oQsaiP4at2xCSweALYahrYSORGl1LxzMRU1fUT+NrH9633Oz
Kt39ABgf0xtfTVYuwze1VDxg+v417UauCFSdvNgilZxklIf/2chZCOhUSP5OVz164i4lGvVUCZ0c
OafI7xZob/AXRQUNWnFzL5uLMxznDkPtiGby2EXOwwJEULpmcncj69Wzgpg6TZsjImS+Wcc32yyE
1U84uXbCh99iyFja653Z/swgHlVASxdwTm2b29et63cmh7ObJdDGevQAZpDYR2wYo+2Y1h/e41O1
H2VkObNSuQQoWrtHWfw/sFTVWsDH6gKhEHuVZFon7YtGjqH0jUWqRzd8Bu5zt4o8K6gPOTXdBhYY
y5uXLNJrbf+4mHuuLnldXx7EPU2kDLhZFLGnD4fj8LlNEawrKVJq66t8V2W6essGjP1/05V7A4iS
+O+LwRFAg+FvtIqW35lBkmjZ+xIUySfx8tZKWeNnCpQDCaXVqw7ZEigb792f0I0saHyBOuGeBb05
JRLK1EIh+Hixuv4nnUHA+hUoY3T178k3LlJWZAbNsh28eBdFYBnr3qJFW4GfFX68JnPvydF6A+kt
dEhkInKGOm5f7PlKxH31ZyAYqaOxzShKGp6mj/A0SwJACTcxFF0LPcV20uhfSKBOhIRdth+jLjvE
8bck+ZJAMDjTLm1vtvclbPG31GL5yRFqfmuct0JqR6x1Y4ABgfXscTpR64t2KbKRk56kfbR8I7bG
PSUIhcjYoXWkQFLhvMTYM30j+vVKD7bAZAZoRbJf38HLyI7zkc8nKoEogDNRkcmARZFg7dEwQdbf
XNee4mjzwlmybxSSNamS/5pgMbytIRycGRr14L1tH6TjfibJyqdW35g9RlLxDSs+OzISM3fExI39
ZKuY5XV3NbwCe2KjrrKoetojcmepL4VbD16JqnE7Gj42hJ7BpfFkX1i8wyHHRcAZZ7xB0phYhoh+
2rajC1/wwN3oPXZ3g+BlFokRy7QcN7NGncUZ9NZF3y3CsAepjTlZw8BpuG+9lEjWt6K1CEYydfas
YDeFsZmAD1018LDxKdLadYeNHNdh5i17D74UnYrHAfG0IBe4mGRP3E1tS6wxjjXUBZ6eoPlfOmb4
7KNf0/Yg7gzLQMlIFA4OKA5EeYY0MoHGRPoqzW4rxGZ8co67M663zWKbNwbuDUnWOvOoh1dqw4ED
Ymu/16eH/93tdyouvyaTXVjxYhEpFuNbnENU4kiRQ/GH+YymOZfZuKC3ikeVg6UteCSmU4oFPyfj
b7TUDtvp20NyzWgm3u0/OjBk7TrKIARZo/xDeRkefpC8F9eHymCQF3XBLk8ImSIp+l4jQoSjPL/U
1Y3LMng56WJBCvyLBHSYfFcjZxF7p7N9QFLz0IGxMkd5B4UMsfCzFZRyJarhB7LbiLAKbrp9k1hc
SQoHTqeL/1/0MU8TkRVJNlXAHYGrdA4hQn/OsT+sHORQJacKFgFNM8u5OWIi0gNivzP3atAl8vTV
07k0hUVZ9sCAtTyl/0swMN2wGbLZhQ6gK7UnvhZ5aQWX5ElRccofEqEMO1I29JPkmJO3wUoAoUSK
dGFMSQM7nDvDvKmp+V/SAsmZlUpCWKxAexU1jAb2NFjBxqDCzMtbMc2UQIRuusz8uC1OIFOn04t8
WEiRBqLoFB3EK9fz0tKH/b+XfwA030ROPleE/GhBmdO42Tqjxk4LWD1kLEVCWLwqu7jBD7evqvZ+
RsSwpJuCUwcKECmUdij3zIYMhETViuYsSP5CJjZVhQGDhh9i+pubvPphhmOzSsHkfV9QMsd+gACe
7YVDWVIj+JtfY5S6YgCXc0em8gKc0f4CHazCHdJLOUrMdRp0Uy4IJuSUHQpnK8zV6ugx8BZYhDcS
RmYBBMH4bufL90v6xrMjG9xlOxQVfwz/VvayrkZZYnm5dk0gW/MaiEfIr63bh7tVqM9quL51rvfa
jpcuCT29zEYJpHqXj0+gvwQrrHUA10unO5qZZ/98jjtrHgmNUnu5jrpPpIK2e475L2hRdzjNIQHL
nIn0EklusE520SBnQx4vH82vkzo3CNDqSxCRBPbmwZ3DtnAXnsLU9A8VxIbf6I1krvcvxhDp5waz
lM5DxsyBXTqha0iW7grbWmVOmnAgKg6MlQiw92aP5WJ0FFpg47Jb7uO/9XQaaF7X/yv9WKIqjxBA
swPmtezZRbptD35NArpwpHE5B8y5sZDnIUbk77LVrkPm9BH8/mx8/WbTCuqi9Kfx0ddGdlJAy/qA
7xzAD1ghTzzhbLJbbnR1lT2T8zOPEECmyE8mDn2Yuh/GcVSVdG9LQUw2zSqOxL/ms9zkp0fgsFMF
TXa7mqMyM3DcodTtu30G77/7FGac8scAoZD2kBHEQ+Ul58SERTPR2wweHB4gC49TpCZbOPEiL+Eb
ZIm3ocLxMW8wpzqiO2xns6cNPLwQrIbVKQmD2l9F5HPQyqU364/S1s0U/cN8NlPpONFzv9Xk5dyN
wNBkVrwyLpU/lqL4bPafxGNMn93x14pzBKewF/Zt6kXcC9fnJZnCKaHiXQ6qYxezpZFNo/0g1hRQ
kgwSMVm5Rph025bEykOa691u2Y12de1KiHVixSnTQiSS7oiXTt3AZy78cGhJEcTok8aUZD+SsKTc
huNEbXKUjS4FJGgvJTRNBV2vgKKKvOPcxKZi8P2Wo26EdSaTXLHUyoBCWVT2v1Hf8lAg4yD1h8d7
g6GnJYwi/NrebmopmuYpDM15HscRK0USHlkW7URCuWqluwbFstU2ji2xMTA/I87vOWYFFUQV5htt
FePMcIJnDTy0/6IhreyZ7sytO/PwAKdXSRI6O9+rkdxWuZvQB+07ceTiyHW6bJK+ZES3NpHkWn/S
bseYy6L6F56U5O+1NLD+znl2TJZyU+p3q4VjjX9p4QKs170t2/FSY0qo7ccqoOo6o+bIAAU3BUEG
JkmUldtaA3/UVs409bZkxwoVs3rW/vPxWD0CV8q8sGljasV+MVBY/VboaWPpJqi0XdI/gG4K7H8k
ijcQSC0yXg9oY6wOuSHQ6pEZa3qopzUfhpCtmmnODM4AoWSerWwV8N3I0UpUWH6in5OpLJVWL/qM
GYj8VR1ayOsmaZPJO9nBSyh3+wipYLUsLD3fv8P9RSB3JH0m4l84iK7RNRY97NAs2t/x9fWARUSP
GFaGxUsKepSeN9ZQwSsalg6++Rp8hyo0E7+OnmAemlbJy4qSgbzawqr5K26SKyMacRAduBoxozem
dAGhEct7GrfI2oaIyQtdQF5a/uWGgnipJaVXsHkDFh42nZrSD0xCXHKF9g4hBeTQ+BFwU/Sii/8O
c0/0KvpYBOgyQFoAckpcGk52cCNu5TZ9WMD4pYWxFJM1P6RxzEN1jr6b3zkwgD4yV0XNZS3wRIXR
nnsLEicL5DXNkDANwcKW5uVTGnp70bQeUO5fwPQ6/fsAuJjx3n25AN5VHuDaNKMfu8TpgGD4vmpq
4mDq3/6qI7xp+PmUUQ+QZu1ozu3Gr8SM4w5LVHeuChsScfRqV/qw/BjTLwJJHeJFdNw51p4K7DVy
u7bRWhbNev1PB/lVVNSw5qi/6CAXzFB9iIcJJRVCKmza0qG9NSCENtIL43SRbQOT2sL4CkxTs18G
+blcqZ4DMmtc7J6P+boL03gCUUeUbbwoRpCvu8gV+fcZXIH+UjRO5fOhVFhSLs/cBk4OFP5njOJK
oDA1fz8sHYgZ/y1q5ygql/gtPLYKOujlAAmsaxf84zlg//uhbS/9K9icen5BlcGqg4Yyv4VgEyMn
0YOZcKnwyDQ5xemb5NZbI+1SsQpFvMhUIDGU9N4oz98dWuS1Kxr1ABy5NAnmuRTgpPO7eWC/Fu//
7d+3yYPGRuSUEKJ8WH9FZVBLEtMUnjpwSlsCz/iGreaCKNhPLAB1m+xCy19db4gqk8PEX38NWRmX
4Rg+6M5r3mfYDs3tZQXfBs8cN6O9L1o2UlZOIR/+2wIt5SrLk8Sr3xzRwzDG8zzS7f/R75Eqt0tV
cFpuyNb4EdBsPGNZ9V6BgINnDWWL6KXoRf4r1TQuqkHMju7Rf0s8wmgYcic3xHJo15J631kbgafq
n/Nrq4RZIfE+Y6jzRRhvCYbAhYESscvOGzngzS0WtLzlbOAkRTJ5Dt5KHnZ5+8keduPVgxiyWcDC
wnrVQHTn/mv6tQ4J8ClKWSp2nnEmzMyvP3TSAboezcI0wyMjVqWqAPJdRMxN14OdvDy+eA0OQIjJ
MkxvgTlm+X0XN0FYnVSe0OPc9y36Kvgru4YjUgigCO1wr4QE06Bauds2hzbKBtSWg99N3hsKTpQu
jR0NigGhP+PSWISS30vBGmCz5RdqSQStfrRXjIaOq56GCwKSACKpJ7oV0gzG8qRLVOvluAsMdrwD
KHtTpYABzQRUwZ5nU74N0bHEF6LT4Ey42KeoHJZg+hyzZFgwlnBx9vtUfcs71wJYg4T5kdhT5deR
2GOv2OBn9Suhd7R+fzKZTy2yAcd5aJDRn4kUFWr9gQ8T6lz66oQs7dpIIDmX0BE5FD8GrLH/7sQt
YKnrICLhhycRIajg2/eb3scp+BjRKLm56mVzj3QuwcRTBGR5T6I9RoCziw3fwonODkLJ8ri9d/SP
WSB9rJPQdJelcYHCO3ddtM96ay+RQPt5qT0MHsj3N6YxMzcCfz3+Geqj7YLyFHcNtm84DoiA2hnj
cyM3XwVMhlWEwrB6jWEfPCTiIJauMURsI4XVyIXToE1Uj8KXDFgz0ehWglMjByExVR/aPMk8RBBt
vXtKuRsfjpkSrcK3FvfztoPFRN5i6j+OSsLh1rMokn8wx12ZKBCCWApLrdlXuWGoTwK7TLK8yYSp
FroHLHwU8767b+a5riU74tC9Ve50m0zrhUHGyD3C8/AdD6pkO+0993vcH+Rwy/L2pnwIgTfWUogP
QTpJWrYRDJoi71o8RSD2qxbm81hRk0iZjMUFNkYyW8wARqehgGxkBnqCkx8p/E1nyAZuBFOWfJjD
XyyCmN4PI5ZO0DynJJzJPEzmL9gBCEkcGwGtIFXEmPWV3wRy7iskpUawFUW0XSR5Q5plvxo+ZAgi
mpZd/WvQNcLZ/BhlPr3vGGywfHUOmQ3cXzQSpnApXiTLOUWNuGZX7WS0DfME8oADiNoQ07abrsxp
xECSU47RzafKYK8sSahwE/RMXilDv2sJwnWY6DVv/3TLm6rBJJQe1RL3JYPZ9s07WujphLiGa/nc
BQmZELKL2Uz4vNsCpml4V3eGAGlkMKfdSscylvDsENoAbfjneT96Kqvc3WQYivYvYlqJilXSEzW7
YIE/dOR4+ttDLCtMYvKn7iinkMZa/f4a5iV9vuiwwuYKk5Wlt1v54ACD6i2Bm2IL2oYJWi+yyUju
JkQ0AXPB/ZauABtebFU9yIHmdHJ4fej/4Cs2HuryGME9gkfLxYHd+T6HFmeOjmGrFnACI38ITJkK
8l9OSOmDfKKLB2TCnvbtov69NXr0v41ZwGxxignIJD4eehKkJvh10+o9HfNmFNZ/iBVBcZuKbQfX
qBEi+wocDh+PMBqkUebYu54fj+YpXUpr2bmdF1X51zmR5KQRWKqquLsbe+HFxIAbiAoZrXdDco4s
PpIrXyVw2QfQdRhJec4dHadM3TbFxtWWMIw9QdSyMSL9BG+WT65W2qRr/gh7/rJsDzkDTAc9wgxU
BURdStUh8XCTxfz1MQ+3xtzJp+Oxh9NCS0etaU9hAj87PiDsKQ/I5CJlq6/W+UOMzuKkFFtY4VgO
G4QXKWKYIfugd/1k4ieDFQIhR/l7ewo/D/0TxVF+ZmtktW8mtWyNmS0aEWZzGT15xOLPdb97bZHp
pEtSb0o+7WBK+Nm5/VJQWZ8Lge9QN3pGA+vt0Y0Y7m7l1m4dzCBf9/i7qM22RjdKN32zvekkoApK
ePFpuOEC1DNlZqrmpLZsEZ/s9uqHdFXJufaSWDD9U1TeezweGnAt2T/SkpqUk5/X1tBDY47WmkRC
MKGM/qlK7cB2tfK8Tclu3A1m552BvJJN8tZTvHQuae0xf5xuzYD5b/pZXp6eJMSDCOcaoFoLVG5s
ouvqxATIhBvwn1uXL3aYcHcrJSfca9ZaH7hqLS02/3x7A606EknGjaLAi/kgWtUJL97OKPARUIeB
tV4JhLnymEogoUA96b0H4OkAYCMSQDrixCTncIxJJ2o581F2ZTD0kS8H1fESsSwGGnf8bWx0WYkq
8MWHn3LEnim7CLLiH+fvVKGoDQPWrR1+HDlE8GbuA/wsMf181nCn227g1a7xTidf2H/5jL4JWt10
p8aSY0xkZ/2xc/MqP4BJFaY90rlaY0Pw8dczYBViRbgo1kwtckXSgdMsNGppQxHGmV+Eclmya9rs
VTvKsM9T926CncjxRbX99IUTTc4UwQynWGpbV1UXPGIgWUoXvJPC0KwW7+04z4t02nxGrmHylxOQ
g1IGbaczOzvSBxa8jp+8hUNuVslDAjSC/cBhkENX6NzU7sKPjO96x0kobK8x2Yxpbpp+6rHEdnZo
zn5tX4dVFtL9PFgbcVnRoXMuPPvDUvCxGR3ccNow1WRmEOS4g1hpDBEytd0TzROYYC9fj2XkXVhv
uzFcbLG/xUByYJCU394sshGiv1bQh+NszIGyEirv+1MusfVCzw+CZLyVOz/AR6pKDoRZ6OsADvQy
lFqoldkMvFHQ+uTdDDBP9e0DvJcCN1PWGiYHhVOkya5/YefuSRdalEIVAVw0+VmAzldhS40kKTPa
xTRT0Ya+96hxO6R7UAb7cSZXykjg3KyBqxCdPW/SxAMSGSCGIPR/KaJwW3VtUlx6ux9WMof+ARXI
KC9gALw5P9uANdXpRR8hQljlZkGhsoSc9epLtZEe+Plj0VmNniX9n62fPGgVCk2zJVeFvEp4sIJO
hAncdx7eEH66gxGnLGcHg41CEzvQOpdv60u3jkHqjSN2xKdXbJWX8m82TyDkDUcKypuhOMeP3NEh
2U05bqLkKjADcmM4UGS14eWsFucZl4mSKdPCdB4SPqIZOgDQtEfIxhXMqNw/5upNYOVnxmUdGnf8
EKfRsMx0AOjzifCJuYWUDbJDHibp0QR6U1ow7YXrIoHGSW0bYhNWSfVnh4x09HBvq+G41ALoQJjU
zUqAHb1ICFoI5+bwHzujhLCb14pzK5Z1I+6dBBqCZ+NPKxa5yIuNVnVqH7LL+T8/barX7S6ZMi19
9b19QwPaY8GY696k8WZGwxu8ml6K5uL6avXrc5EMvjagdkn5o9cEEe42cEEavdOytUXtM0YQbHiv
goas/CI7N4atm393DCpgX6TAtKWl6LNHefwz6UI+XD5JIrP3WmveXu/ZJKqZu861wqtc9uaBvrdE
oxOHUQYItULuc8CKxut7QFxi6RkxiTYg9dAT7f309PIEg+zGABwSvYP05jeZIRYqMlmzKtcYvDC3
JzplPhLL/oPZ5M6acb83sro4yAAem6iUEBf3OIM2sleC9f0a6BU+4PGYMsYLSS0WFG/wmCceKwlR
hObEoyGeE08n8V8LPu8UbLYscYA2hgdoXg3B5VlSUtcDH2JK85R9cgN8cISTAADxyekNOPc0uhXW
6kJHWDXkAqtB5CLWGrOhBJYLHASiM2CpqRu6ZyQpo46+/JE2UcqLYFRS1TVfIjxjF6xFckEZiR5p
B+Qc5jRwgXIdJnqjk6mdwkyVSsnA2gSP5ujtQU1eA7CcQb6mwMwV/F3f2tCoF9h1iFcdcG4ulAPh
2iYKTJGiFfuaSCh5JI1f/PJd8Rs4r0cP+H9FIL6GXVVNeBy/WfERodu4S17qWEeyMokVWHltXX0p
+E3u7E3z+eu+I89Lc95KO0yROWCy3XcG8AL5F6IWqbISianpsX2zRIgHHFG4Auxuo426n77exhUo
bugWbFD1y8j2E2VDnnHdoXIBggeYDbfLyA+tzk9jZBoq2c623EbhRgwuKu3MbJZuUD9vAepUMy9t
HyOYo8ugodGBcl2jqtJENbgC7umlLtuHKztMOlDYkPmBIoU94wb8NUa8PInMkMc/62KasPxv2f9Z
251OajeqT5XN3UsEJvOpC8V5ne0CmVUAwNax2QazF1egFFQZ/kgBcWFaMrrcVQSXELjZd/cEQ965
HOKIe1spA36lV7uYvosnFDzafTr6CweRo/lWXHIcUrfANX1VmCOD4L/M8ZYGXFyXZd6KM/JZyLb7
RJ5ql0RoiVq1c2tcPQ6kVMS5d7Qx0T+hUjr4K8LdDhbR+cmyCdoMialMMY8s+ByAF5Fb+7BdbQQp
PfMTCTPj+rwZjt1PzCZ6yWe8l3BPwh0KdcobrSUsWPIpMQxWGcQUadeRGmMynjslGYT4yUCl3DVS
jiOHjIKek2/7FKS2EGATuqloAaX4ntmAqhFnUWa+y2hhesAMTTSjAuHcwM5zbv4K05ACzGRaSzgN
AaZBmWnm0LaYvth5ffCAYGyvaIskmktMf5naJaleMQ46IFy90BMwBaXeEANzelDT7H99FtSF3WgP
+Lj9S7SbJfYPNp/c+Z8P6IBWhirWW9JxbpTFwC10jBJlGm9s0FSDvX2g1eketrnl3SuMKN1SuUeD
T1Iu2rll300hEgDbhfa2iEuM4Ym2F+orhNaENJGQ29ceqCRnYcKwo3YoIOROAY/tAx81sFDnbg29
j3GvSGf3tRAl9bCRqWqG0zXmP9HMtlP55d8djvNQIHUKQdasKdJuRWxnSX+fJZXBEn4ngEMhqgxu
gK9yBpAggDbF8JwwQOlDTTDtFJ0ukpA8HHRfyGeOoKEfmmVYAfQ6nqysVMDyySYKd2FGr6SbFSbA
Q0zECJSLtJmoCIX0leEIM98ndgg+aVrV0/k4XKGSGc2I8/BLsPJ/a6TFnRi7YQd78vuZwoB5QNQA
ai+UnM368zGtcInpgZF57+qh5tAzQprm/AwrdvrxlnYmxfyXf9tkUW6Qxn99zml25vq2lF3RiwbN
WInlp31YDkqf6kDmDJGUq4K1lAWqKSKkI3wGMLRHgdwn5qGxfBcM2qQw+PC+SRC0VkA76tcAf3v7
fiDHar2svyXUbF7Z4qGj8A6G8h8lNEAxQnQYYs09ZrpQnY3ZUPu4KmXmvGeb2rY5Fqdd08g43A6I
H5/wiXWfLl2Dl3rEPcAV9x0IBx+MxRV7D58I1huvmn/FA/uZiOfooTHwv62AyhHda+fN9ZWakeb1
dR2ptfcnbOIwv7PnffD2cuaTiRNtyHn3rTf0Lz2SFirxsIzajam4De/bzyfXN6IM6nITgcE3mJvn
7jGqrMxBA8gQd+Z3dY3mAujIusuY8aSnPyDodkSZPZ6AghRjHFtXjAZ1X1gfUI+sy8KaHjVl347j
TEqbVUFJCy6FMJSO2dgv+ll10E98B7sq34zhSJmlkpVsrJpZN1bPpk9DOT7QjCF+dQ2fTeBGFOy5
HBAMV+ICTP1rpimq+l31viSHo32IQlFNEAX/ZU+OO8K/wB/c/SBm9IlT7KxDX60/sDu2RjfLPTxX
Bpc95aP4rtVwFSVznwrCo0I9nCFVBoXf/qq5EfZhqspVCamJ/1NgmNbHavcEvlzUdOUpchF1ducq
5gyps4IJvhc3IVNl9BKJp6Ctrn9oSckL3IvJ+TTPsT1K9TtDWvOJVqQRRe/FgdksX+xA0WbaMzPS
HOcIHhV3ktxZuRPIEYKBkUJPGWYCCzV2s95ig4tSnx8KQ0zkzorSmlO5DE+oJa1EgYtJm0bZjQOx
Rhl/lbT0kJI/bNzagyCJWV7TEAPAi0YfRCn8NmpIP3jPy2w/sE2+i4u3oAm3Yv3FTvYurddT+DuH
3utceV2uSXyiTrbkIWg4aXikVVqUjGDrMqGIQumA+OfSBTS/zdTFYKbccjvpnQ9l1FgrjElolS3I
7lAIMZd8lqnRB+LW0FdHo7xY4WUDvOC8nSpdM/8JzgFKUEYaq7+O5FVqmTzf7YOx0IyKqciSPIod
0X49/W+AulbutVu4Gl5Ek1Tp9XGer/BC79FzmUlUeF3vjVkxzePXNftJgx+qRVN6LRF1rGVJcarg
uMu5QmalF5EGo4oSDaupyzIFV1hIhYITUHtZXuuJEw4VEvyXBf4SbrhiHanrdPtt6dkZ0SPd83LV
ARYI4ki0kGaXky/IQIlS4sb8acGB81oSLT5jPPKkRetG/c2WYh+3MXEWxNAGIW/KPCo0sHdSrvXS
ZP0FSeIjF5v5wxq0o6+Iy5TP1+HDdUxiicZe1upMUDoMBjymZdNoYGblxNsZuQARbZgCAAjayXqZ
bHi8IVqDYbCCXiod0REQQwcLbvzenP9Z9by+X2qxYr3xn+9Z69Q087NXgK+YovDORU5qviuIbjOI
ei/qjaj1NEUWrZxqrys58xNQ0J8hJVyJqDv8wBD/jpDJYw6R8DLRT3cKqIHQcwX0X/cknu9vgiUt
LXF5F3oDt7VS2k1n+KD9BrGVEvRTp0OTBHzZGHB5l4KYp53xtfQcaotPz3W7T9jHzOMN8S854dsF
fmzRyeT1nafnQT2rByR7QtZ2TvKVulYTBShvA9qizTr6oKK4EvGhqciyWxlDTCpUGynSEop2T4RL
/1tThhHw4wi4zbu1npORS/lUKl7GnMKPRA8Gsqz6qTTh9YSX3rlblEV651ncBU5i840ysRF93UU8
d7nBtcv1NRdu2mWnCDfUdV3eAVEyqaFyMvQswhJaKXMKej7IdeWve2pEp/Gg6cfeD7InIXRE1tCz
6tc44BHkNvMjQ3w0pKlQEcds4dBr0lVxkJD/2tfX9MWLNUsJfoUBTejCDhCxae3HeuFpc6wjnFxI
EKma5vqi7yVrzphVsw9qMtu6P+UASIoPHStWXxruBvoZZuD0++JgLurtuD80FD3KBSpkh2nvem/y
df/2nypXPVQnYdoYzxzHObIgfflOkqgqhuFHZXv7TsLEOrVkgd3zEB2a/IO9f+EugDOzDi7dhbGZ
iPWeR/bcQTGaTu5GPYqENSrDfuagbiZAPEFwV+PQCXil3NY5ZVfIjHFJysQUltlLZ8OrEDT5seHe
FwxHSd3xg0vvEW+H24XozDyHJ+XMubgAzUbRN09I/a/v5H6tuYNOMCi2j69pXtwXmJnYZOmb4oVh
AXeD5woq4chS06wOoIYkjrVkKxC6G2C7HjjFAt8RaNkatZU9EJ5RSTIiDVM9Cix/aWOgF1eVXz0/
8ihGHrQapuE099y8zwDj1CcRTCMBPzNl1kVgXvBtMPBm3Xfs4XJjXCzPNpT0tNxbxr/7ZBOD2Bin
Bf+oUlrVHtLtE5IsIiwyTpiPE1MgKt3D1cBW2Y64Q88E9OAFX4qJK0/KPX5fZ8xd1vqYzWK2X5IG
t08X/6lZkWdiqdZ8v9YH3/FZVJ2ton9sYyrYfx6fOpmz4GZV3jlta1WjqKAOekUv0KAE6F/nFaI7
6BrAi1u/vrrCF2I5R4k704BdJz4EqWa6b7RDied8VhHoQE5YSjv2QiTJ9edo0k+12GamevrnpMK5
nAcc+si5APnnWQy9TX0IYT1jlk6CG03s4qmZ4OOMf5CgxlzWaVXjiGwj/mNGcjIobCVufH5t0rBq
m+ocR8H6KbSHinEvloQXPNUlMrrTgWtVlp1PPlwKtI/9BAUEc/ejiFPSf8tHGOtL066H6Ar84lEP
GLoD5Fvdvo+Wwfcx/83jEPc7pyFJaF4m9Z3qVcAxuGBQCXleD+ZwNBMdCY4yBVh3J5n+zvHILJRQ
LwccmZag7m4A5vLpx4VZwIDUQXdAA87xjO/m/2xthsxrWphb8iAaiOfjCy/SA8vrsq3uJBq16StQ
dPbQn/+Szy0xWP97XMG/qt/UQQ2LLrNTvIO7vbsBEOSkLvXTYrggeSYxK+vwiTp0U8/bdvXVGApQ
QQXrY3/S7PRmPxO1KZxINX32rlOQJYHktpIPV8RgfMj9kw7ZdvxiqkTlbqnv1e7yx+Fn67IlyL+j
bMh8qA/6UbuQxoIXCaBxKbahYjk/dF7WtPSHS4PdsDWskqkqk05lfa3OhymxrJf2xLcorv+PbzPN
glSc9zHu9TJnhFt5knt4M1dAwLAV5y8vCTDuMYLhRrtgrlJUhDIE4dT0yoc7CZK8v9/HGYXr9Y8z
4lO614DjgVMssQKje/VCas7tQTwluWGdMoC7lzQPSHmVVcYzibHzYR/stZ5/z+WGahrPLsIvN3xK
x8yaHtp/+08YCqUpW2sO7S9oTGujn8wRRDPtYXXFA5KZ1zSUBaPWjb4VyshFfT+5YElKKGCvlXOL
hJF1vHCYb8oUdPmt2yfQXmGn3hTMKGK29mQI6lvA/Zf51j3fdihM0UohtkSx89jbhr+Jbt+WQOQ5
MvDP6CVsrIxxopfNR9kIbSxw48To3GIOAxyHbAm1jkA++B5e2BXJ43hLpOlS7jCwFdAYQFQZJVNx
T0Ay7Bm/QeSmin/qQ0QGVxMsflOdlwlMO/FTrIrbs343spJ5DTn3ypbP6e7Zn/fMxvK4EmW87s0U
QBpeh00FbXDlOsr5NCxkQ7ROVBzAIDndzLd9qNBF15RrlG8ZTSW62m1nwdUzuuhO0YJ9fdkBBS3L
ECi/lo2RBN3y1kEx0SzOmMZbuxwm8u5S12S1Egm3lUb6fatS12vhuhXpsSGoNncxUsdvYfy1fCqP
w4Yu8FOHLdSiB9ihp4ywSfFkoEv7Pp+B3HNhP5cB+dtn81YoJbWkP3SNz+1k1gn8V2mnQ+AyfXsx
NgU3lKRYy6Ne5j1LfQo6KAWUkRe4oAhkglCNu2P7cI0djzJbrfU+LX4Gqq7zJCLwXbu68X3lRB6v
5l756vbgtda7GCZql9VxNnEfWXG0TFafXAhF/dOkTE5aoRidvv46DT+RVA44um9I9x+H+BbqkQkg
h1hHFPtALB6dKMJEA1D4jUDHvDOAw1Rj4p3Ca99RWLBzsY1xEtSDdInikgayzCUk2fms6bezA28F
bfqYoJ1nPsr03wf+fFVvPwUD6aJbhYhG4m9xWewVWK6TCOnohgkpIxthTCZn6CbpPALN5Y0A9vs9
5RHCbMgKP2T1k8IyulSsA7LEOUr8riFZ/mogGuid5ZnrVdKcrvqaFfZc2QlzEcuTynv7ChkFeaed
3pvL0CFjEZGCbIUMkoH7xX0UpxXTi/lINzPYuF+R2Jvx6OIBsJAcvmEP8lLB4cxnBVDz0WvYE8Q2
rv4xYzdSo0iu0Yr0VWJBcnFah8w2VJWq+uv4OYEEYdqVkBXtV1cTdMpTX1lCj5DGlb4ouHCwUZRr
HwL/a9W8omJIvGmOui53inM436o6wnAZTUVluF5x4qlp0136vYMldW/7i+HfWOKf5PP2hA9ts8Ea
YjlIKJr/ebwDUYyj0DfnzrSDnCtzLgCSqosvNgDbTpJdTwPObLvmxbLOLo9gH1yn62F8OI/wtKYe
Aa72iSajT94q8HTZ3VLjCiFs+hkmkkYoGj3QFx90q5JKRY92dpwK0APWDcQNzdmWkVbNiCeQFUdc
URlcsb9rUURjZprEFtHFWlQIxo+2TvrY7PPl8+GI4tfgvZX74ifHTPjAqPomWc/88OgmVE2gX1N/
Jch5iX0Gy7QFQFFbADxO2L9RygPKHEq9CMuvaLSFCH0NSag/HjW9b38wt0QBS9y5UmVaG68/NLmq
F+uAtdDl5E/jOFm/tUzKObvFM/JaN3ZQhxM3pJinN9O9Xs69SSZk074S11A1NQkYygHbZXUUIDRJ
4Sn3gg1nzEJRq/cpFr9NaFTesvx0wrPsqlThGhGQRwZJ7e+QpawBbrhQf6HQFtzXO+h2P3Z0rWDY
MG7wWP4GZptH84EY3VClpIEiZFzxlDiiGbAPnanConk7XJPzkyxk7rBIC33s5SAG3RKwihVGOIlu
LncNGc7mcl+KDudXqRNZmk+XdbHLUh63U6DSrpmp+eYRdiumYMf8HBahWGbB+XG5t1NF9ZJFNhf7
qsh0gzSh895jyUPvAwbvAuINI/zc7Gc6Z3nWZXWsGdxH7K9XCI8hJMEFq8BixT02t4eGBeEJrK/8
iqICCOHItKIP5O/LyhqxPMmLYeErIxFQjac6qBjHofJktq2Nh/2wL9ConwVBXQOl4+oGmrcnyql5
YaEDxZXVYxd9VxvfraJfk1pZDDKNiAxHbnUyVGQoNtiY47B7JuNhhvC5mh3pxr0/pPly3oLhIvf3
2FJeEsfstbfVxjJ2qrLYL5LjtPba081jM9dd+Ru20ahVuJFS/01IJxLEMdBVqZ+WI1gRHHQ34PxP
K/n6JY+E5eU0LGXTA0HBCmlI4/NsGy3prLqjpKd3epFQlygs1yRj/DOaW8qFb3/FQPa8g51a2pzB
CF0WSfOwu+9ov5Sybbw4zDVhUtbj+Ay1h9Cn+vwH1RP8W3529BkFQiftbE0vK/WFdb361VXRf2j2
DmSlCwKx4WauR0pwE1cvfMKQ2RM6UD+mMtvJwt5ZyOwJkOFk0t5C6zANinRI48G3bzWv9BLHYLqZ
udRy5UBVxu8Y68ToijoG7WdLDppsHHOkLMEi8h/y/Dl7njj4oIGkPbwsqlR5uZNy1qKX95bQEPvj
KSpal2DCXXPTvOAVQhrPA1bHKJie3MWNaW/QRM89AUaR5No3qrrD+4i+dckJKdyFwKlvHD2XVJnx
OIdbYHqirYzj17c0nQ/iUGnEImHY+0FK2umU+3ph/apFtmt3Vz7xdCpJwVdCNpvOdv7eIuFBj7LH
CNd+I1Uk03CmGTcyBGlgu6Dr6nf/G3alEJ3PhUCYF43w3j061EEqSOAOo0eIDDMmpsUnRPDXXrVq
P0VLponRdh2x4BZwpRmB1gl6ub8UerXI1dg3wCfCkYFYWZ/D2oBG8aVxRYWQJRNRiIbUCiKX4k5x
ZvlWy/Sm/6dtxY1lPLOiLFX4lVNBQ0OZYJqAoK1+y/DOyq2ZNixQ3On65A+CNYW9Mqte2FD53WOF
opzdDgwBj/p3icT8RwWOqT0sc4KeQR7haKlx+jRzwkuaYzUV1eMlNSv7gDpdT4M+ZZdF+Rlxx9qv
U/VrcQ4Elga79YPieLTUODTHuPKhTXlwcnA52IPZ2P59+1bt3qnfB/klC8nZj6U5av1hvoaXxY02
1SLAGVPCnTgMAx8oZKktuzOsd4EpNgi4rhIWjS9SalE8M99/S5/mEn98PwyXwruuFX2CdQH+sDkc
Axni2IizXD5/IpcmCd2HSxEugTDam7TjnQR5OzwI9AWlsg6rZ0r50U5M0TYOfGas+fTgofrH2oOb
CSesJ3IAfRqumizIiTLO9YDjYmmTKvOjEAottGkr43lKgT9Q9R+kbAiCeDF+j+QoP6upfmIql7CH
aebEywypsZIKo8CnJXEvqSLW6W710KRJ4XoQiQh1UFBg9TODq/aDoQmkZRM19eutWGE9/gEhthkT
JNGid0BAb7VeAKVny4a87bDToFHi/VA26DF3fEvdxhdfVUZFo7Ylco5dxpulwcm2UqlZGkcz3Qe9
tyfWpDR3ZAZlK3DL1cmnheZ/ed9tipYcHMFzTL1fwvcc4D14yeUEUpbRR3FeH4PbAedPRiFYA+of
goim1kz6yevwVNQec1AZgzo74hD3iCYV9Z9D6vtqq4UlNjbEvo/3RGOEcxb/2PJ44Fa8WK35Fhbn
7ClzD5aoFvqir0Pp/+1pYj7R39w9jW6QSlp1R5nP4mJWC4p/KAxMezwhoYq+oVvisdXWTAp9aRJE
0bUD86N0TSkUGNxfG+QN/D7De4fHOOKmhgVatY6y3W+ILl+kd250f/ArO6znjtgVkloL4Wjgrc1r
bpo3uP0BWoz+llFw4N5FD31Q5DrGhFQiYfbV+S5XT7bW6uTF4Eb4rX3GakRPtAZCTaj0EfmLV4qL
bN7RcjF2ud60JF+dCMakZrhJCULJRBJKlcAzC9ngm+Ccdv2J3iKha3CWVKIM4nqPLjbGuSSd1WjH
lp//FaqwTB+HEU3tMpSwmoQqq3xduRk5ZwtAuIGtC90rPKsmTEv9ISMA1OK1GlMtyBJPQgs+cwjp
iNe360uNTmEQCYrjiXy2P5F8jCNYk5LVIxWjvT/6ePHvOforBCfSKX9pYyxDQ8NOI3/1CGLbAP4w
i9aJg7bC4bghM0I4q/CVPsWo9UAGrj6Vw63CaQc+zbobS4zc/tYMDFvsEpr8tnVJ/NNJn6gJiHnR
S9qGGBe6AH8mWscZWGwfH9gDucyqsjgUVAm+WCdQLTuSSFXu00O4Os8RlzYJI+Fqyi4VZpL0wpjF
gmCccw2MRNx4M0fAqzkFb3X0kmzv5IDt8b0pPT3pONJoaW5aMqYFY2i1QXGKLeylxPCwPih5cNyo
BHr3VQy2J4U0w0qu1SAtDvaW6zPwPJHWM69zEHqGBYIrUZBLgrVtdDOVxjysU7u9Tp+X/Ddx9eb2
WsDwgCVXh5+WtA1YQLrMeZl/nJKAQyCNxpwnZsDOjOl7KmJ08MaVE+Y3Ja+9APIBVFUGScswLA6v
Cw25rDkBywGl2MiBaYQJ+f2D60slyhDh2bk8BrFxxlWkzJTvfmnfm/GUF0J1D7GPd8GAowJR0kLJ
yZDmqjf9k7g7tREzrO4mTNmcP0hd+NBsCIAWqpU9ID5ayUxrrao6M6ctXdCcjjA1zNEUGmVDVVI0
vsYefFllEBys03P8gdF5sEg6FEgmWzKejpSLFdxF/1/FJgBDHmuZkGvvZ70/bROZZJpYWV6VpTCM
TzdaW4EU7a03XIgJ7XXFqqC29LnGuZSYgyfaIM59xt1qnI26KnUmwG3LgImr9NLBJ51AX2JEkQg1
MUcxvxrWH6YLhyIpUcegmT6eUH9H8jL6wpm30tptJNZ36jkODMpTXJM9PS6lzS7gIctrwMi1IXD+
l4QRRhClIszNXqfqYfm/mLkwhgLnBUlcNtBkhwGBd3V0jsHVMrWlbXaL3IZOLVzJ9qYz32UyyImi
84fjBR1oAFD89ivzWaUVq/td3rnXEz5CfTtJZbZhZVRynIV3AqZT5EF1Jmbz0pmCONroEIRUnfoh
GOn3uuFL1W8Ieix+y51n1NDVGapUaPrk3H+7nFMGaLMjSwIZbVoZrTgSFqwvnhKrDtCCFEsG2SLW
e90vJbERXn0W52LozqTsafg8hJxBoI0655PuPKHWUDqaW8gVdGirZMdUqdtWTw5DRgRxhI6BaTVO
7QhdlMuU7eZ8KC2ScN/o1xWrMAkuCA+2unpQ7PYyIl/gnh4rkTEWePNyLmN6nLVP5PSZcE+ZeQ9D
OqeiZ8vQmuQpgXkhLgKJaCc9IKdlVwJJDqETE9JIbgsZoKtzx9vO3ZTLXKbFU5OHm9YDxHyGbu2H
SJy6qocgDQw+n+mp9FW9gfvC9iGrPqh1E8z6wWv+es1/4UXZpMu/GWaTCQiwUMEcMWlH7NghH7sF
Vznx0VTrQSE/r1Vr7Rk7+w4Trb3ZJ4lLYi67DnAsG83D+xzh/Z4XC+KXtkGiAB+3jdVY7uAm13DB
+OYOndpdyDlNCucaR1PH990xkunExqOcZTMUzz20X0LE+1mhIUnUJOvsEvab5ucVEvI8+MVF2wfN
f+OvBkK1QaFbSTVQxqq6hAqMWUWu6XMagrxE1jsZx/68/WpNcHLdmBqHMzw0doEamai3P7uMHoI8
bN49RXTHTU+owNO2eTUgxYb9ly+XecU26891M3/vZqLtKw8U/Zbs2QeVsEXksQVW6u3FVDMhD60k
dtEnN6M59Ku5j2N4enZp+aI14Saqooet6UYeuSL4G1RQ0qIoO5iD+k8ReJkdc9ixaf+j8xIZSCd3
YEUvqvZ4VuiZxl0z9uquuYqCZy2Wyn+QYJiVAYE2ommnenNZ0nsPKX8aBqIRK0tORO/zRjfVJugt
SG2CF40vsLCGFBDX+0DHCJFgtqknex9wHP4oeqcJly5/7cvjAUMz9JTfJGBK6gwCUTKFkSH1TcS/
e6M+4FFvM+gGvx5ZVSm9RUzGF2oljUGlymH686lxKc4qqp3vP4RlEmlkWvFxJ283G5TGzkXwxi05
Zk3dRRDJRvfCAtUaA9knzzYidH2IGRgrw5c+r6RU8Paie/g+noHbb05Cwjgb9WqyGQ7Zhpe2mGUR
9v+/FBP/bUgjj+zm8YrKRl4uelTNMYNr1O6Wp/25PUImKY7bJjT1c/uMZfejDsiBBIMKG+dYtI8m
oeKEDgFYawSQe4zzESIf43p6GngvyvLh4wH4F11qYz1bOJS242YMg/hTUFeco566737fcGbNeaHQ
qp7RyD+UfwXH744bXC/45vGUlS+BioJai86rsXp7XtPajNQoa2dj4UARpwfGM7sZonZaRb8WYQoG
95BvNY5QWOZ0yNf10nMjzZ6vH/b12D/1+w9xv1sdL3U0KRYqWlpNE4YS+bBqF/3kfe9vVkVgNd1A
ay/OyLE+O6KjKNUagx9nkTb+bEb0YJX0iCCrpxoRp6hQDdbgrZeQ7dBuzIyeyzI5i2G58HNSMktP
1P8rpJqDW0KcSctvPyClrOieNygJWTczsIlYg4811JOFdlhcLm2xLX+vwWSnRFkSOnl7ud+za1Wt
F5qO4Ynq8hvBxayNNMlnVarYmmxGrAjYAgdP6+GEXBbnRBiW2xLkhhpcNIcg+MuQXXD11fMtMbuE
eGdRImqLgFosD85PRbriWK1gQQtGH0oOgA8hl14zph5SijUBogwLr7jVaMlA21Rxzidn3+OvfuRR
lnmlvzMj2y0pq7FwiGTVbuV7jC4KxLMl6foEJhG6dig/ROfPzIl9LVLzimE1unsj9FsXQa0kogJP
x2oIgyK9m2iWT/ydVpJL8PXHz2UXSaq/HVINc5t8sRUYxfPuhMUsHvIvXcbRK+H9jBT4lpSFf+R2
RuWBix1IlFAChWQh04hmuA9pb8MtNt/SLwWyBV+0DjbYq2KFebFJ8BVdUmNyM/fD2ZJRezF6SikZ
1Qd3HTyJMTga+q+GQoDvbfAhmP1Lz0ZB0TpsOy1R6W4DeH29Bg+JXToVX7z6oHjBb5yT4tU3912+
64qq4xRHGpnzg4HtrzSvRX8u443WAoL9h5iUPvnkivF9mmZ+6+ZI/unu54evx0wK7cRIrJqTc/40
CAu3LYO3DXdqFQ82lWZav69Xkm4lD49XyJ1Or6x3vOmYMnTutD7aWeX/rn/xLO0MWYi7JubJawXH
zR+qlRJMwJ7mFMNg4yPrgy/ybep/cbfwAlfMDDZ32znuDrH/b5HLQBoP3IBqrR5emC+fliAzJRLx
YjI2gLJyLTKyVRBai7hJtdzkJVlH2eaQSYpMSIBzUvY3Aw2YWt/SdnoXiIzj4ORyYULgp5GTWXlX
t1ZeE2nBeNno1b8zyEj+BNG/Qa2g7ebTtG/6JMrvFXeRiez9PkBc1aGJraPXZ+ATmHXucfy+f9Dh
+mV04BTErPJ4yhUIQhxnMjlzd1xsn2GkB13me9m9ruZML8WDqqdOVGSchCv9UKehwrtkCGCEJ5v8
NgBK/FwF9QL1/ucdEjxzpmGbg3xoMQ8WbPwtwMphPgFh3AXe+BvSIE1iu2VRVcYxfv5gJW1Ea6mY
gmVt/tnre9zo3TyvCC4EzoYff67zViBJ2o4vymXbNiw28tDzG80rwqcPlL9CpQv9Yzn8rMwIcAhi
FhZr6Jd2i5Lp8DUMWDbJKLhNGhI4ETNFyEdQvf+A5A4+/8RIpIXg5xpmSWKLinyhoFhgDLplnCbt
6ff2TPaFJFIZIm/XVvqdqwVu1FFJwD89AKlVs19WFWe6de8BE3rHzk3lUgZ8bwri/RBTucZ08UEb
zSSKTxZIccX+MBuYnRhkeGH3qAbzUNNiHAX/E0ZoCmANU4vDLQM2Mbg8abI9tKuDbQ9jgpSsjhPN
ckDzAPFPorlLNGKI6817LqTcO+pZ7NqnCFkERvv04fi6AV74iZTNgPYWcNxNWpmbUaCwQy3wnRp3
eYyHhCQMAYMe0d8ebpV4UXPqMSx04diEKNe+LvExN3bZG9yD8wEoRzVrhLE7AusDlKfMUL7P2sPr
qTe6oQgOx03dTOYwUIkb2FhLyBi8plCpISKJGfeD1aRxZryI4ERwWoMvFeE+lITSrlWPho4VQ4xV
hXtuizvYtzfw+Q5wJ7MXs1s8w7hUyoAYrr30T+5WWxz0FaYRrJSYW3nmgF9gYKfK+PGnO0NPiyYr
oaeTGJ1CYWr3LkkiZ7XNitoTfIye+dNhWrZSdH7bZUvDN6bb4RFpmBm2Xp/E2EiHsfq4qGZJZv2i
XlcWmVmzJqapKLzFz1/A0PWR/gLt79hrfDTMGvLvJWH55xQXtJKZCtcb4FIpFEBqF12u5/Gugn0L
bNfZd+Uj0LiFAkFu+R1hDjnsxrDe6Xugi662CKB8ziKjmpZksW3uVL9wcL0XFj6TbByjFQcHnruS
tcaEjQhwRPthuIcUQvOcLpLrGf9hp5IF+XhGxdJtEOQw2aupsmQRCwGpKF9zjnk2mtQesUtweWVf
9k1poeaJSvN2AUmmRvzWNavPcTmfxp8j/nuyIHcR82/uG4aX08ALOOC0wCtMfxQ9klMPr5n6xCBR
M3zysaxjJKyRo+9DL1eoDC3yMbvPq+LP50kB1a7sOdqiavdvd2bQOTQs6+0sHM9cQ4a7ehss7lgG
WpA/mUB+YrA2IVSOamofEmjFl5HvDi7pQS/67lKRiGPIqTbCKmuGFOPPTR590rPcCKFMGKfA1V6I
cxICnqUDjE7LHILIRRbdnuPVQ/tewsQ+y+V+brhzT7bb1BoFlaf7mbRtpnDu8UU0X+KL0XEkyG2/
8pO6cgRVO5on4C3bLKfaUMNGEc7c9sTc2pkksSt7WCRQJCBwB80Eb2z4uGTeL4pEiaRAxblZo2f3
IRRrXUIbSsXrQbWBgqFuPnIM6zwWi7Iyv1bea2d8Fl8udzbA6Iu+GKQs+vFnQys05hpzDMdrl/tG
ZSs/rkj2Ho2IRK8maJOWgQgBNf6rc3mSpgbII/OlH5Mm6KTPyeoAJyv1m53GqQ8dPp/Yuh8EWmua
1ntkpEjUoH1p6USXIOCkTCKn50FOyiULRHC48lkik0FRq7MQKHbHapo2LHSnB/KSx07qsyl508wJ
RitJfTasnkH1Q3StE80KBF/ddFB9vg8A0Q82jhPeZZ7yFyw9oEWPGl2/2GbfOXzHWM3tbELcFs1F
MkVCR51XR+2xUKmy0qWz4MO2i4MdTszln4lPSM3Dw2aibjVqNdEInB5bq5QhyRJsFA+61qv9cmyU
p9J/t/eeS0jGEPL2BJ136wtYehokoW6wzpTUN2LuXeLNBun8vfFoEk/X+4E2nPhzDpJBnZdHckRo
i/u+GP6iYllTV7zjMSug9gqRYuBpzs09u1L6krtIJg8DStPJf44iDGKYMkP6S9qiVwFmf00a1uI/
0v/V0UDUGBt7GlHWaIkiWKpu5L0xUGauNEbroGW0H5mf6wK3Xlw7cQoQBynxeFe4xQhOj4OE6Bu8
dcdCiEYTgvXGybYHj+DCc3AJ5FNjte/0RdnGrhwipwikzspBulV9tIJEr6OVH2Vpald1JEXwS2K5
Ynoebir7bxvAh1AhS7+nY+v9XkGMVCQ19Jv5smZxt1r1C2ocSWlQFY5SlHgOJUs7r4f/YoNp/edW
9c5vR9km6tT1r5hDXg4bvHn2xU+EocMFXWVsshv5SR7LAFRAhYPf9sIPhvQh+jYsIKtsO6dL+lYb
OFaXqdwCHWYl0Vxew5TNxejJbdnaPvpNoqkvNS+TaU7B4LqSeVpB3OC2OyXHQ5HwxAztdafXHyDn
f++BO7TEOn/7HzVMHFicoZ07B/+q/BBpErq/jX3szIah7G9w3WPUFLUeRm0oAcJn+sXm7hZkqEuZ
bxJpWvMITDT4qe33OIeXRoetAPypxNPAll4qLQIoXZm8fMTAa/Cww+h05JZvwzncDlDkbILAf4yF
LNXVa3GIPO9nVBlk0neSpt2uiRyDzknfT7NwfMhD8YMHdXGEv/ag37Hi5yqpRKrkfqzlE2UEe16X
6BtkMIHm3Kod09+ybnwHvvTHbDaRpjvOWUu5iLLnxNLyf9+gVvkMg366SGP1ILtKJHs4O96lEYUR
99+7g8iD7rH+bnlmp+rfvNJzQliOrg4qgrWDqnUYquKopa5p1Nd3M/dbWVuf5bAbSz8RUHrTlXTe
hnQ+N/vJn/8wl8gX9B3blwt0FyhbqariYikkKIaeYIqBSbVH/IeZsp9A/7UL7Smnw3RF+JK2u6IT
lRgUW8Mgi35v4vRwwcRxpRq3BJsp16nmBeGEC8MihHPOv/rbljng0oHp3MFEMMrWg4QFZ++rA2fJ
NIXvWTOr9ZxWpL2qd8LBb2/8fiOAdsTJO8YqpwcAoWUgV1xclECWNtPo7WH4VRDwQrme1+KER8Cz
SLcrt/l8gqlRMxSgLv7OKgAlFeOg4Lm1jXOEY5Y8hqhcIMxixezW7m4deImjnBY8KAmI3lrvSliE
8Hui7WZRfLOUsawwEh0CPwJA9I8friZNaqMND97gBlkIrOJBo8G1rxwXxYhcAX8nS50dnRva2lFQ
w8GSqFgXxlnxyYRvbnKgRyaDa8GhAYIgK2Asd2RXP1kDI4I96fNXn+AourT5OKLEwKrA3oFvek01
UIS5h4FVqd2uFNm4hEXvGMsq3XW+6UuJSkEU/vHp/rz1+JofnAyHz/L/PByONjGw8eGR59Aj5P9Z
V0DXnub1brvXbVVbKj6S5t2/S33rW2+upYDy9lAYAk7Ja13Ngnq+7xD899vaxq4KzrFujnv4sJNj
mXvBU/XjkgEp0ydatLO2a861D2CU5MCXsWpZ4Qm1xHD3WY15NoHfuM/IbGnfK1XnEJ2mmGzQcVwo
6C60f2Q70N/ee/3tGj+zYuQEMFBYkx+LF3APDY+I/c6Y/TSN2i+N4LCrv2JjPgp+B0n4qNfdxcwi
xL79MN0S1ul9b5PxmDA3HIKxDdWJ5DDu5OHHjbmgKnphamVZu1u0K7JjypPWqxccPNFhgbXi36I8
Ux7T8N20nQlQSOxkyypUcpnqgnfMo5X1zfF12F8tgFb7HTUmo9G09xPXQgEe9uY8YPDJt24JjOGz
NWKJ87iAbdOUuxwAASv5/+wB9w5St5cWfHzEj+BV8IiCNedNWsqMHUIxuvXiauMdONBRYT9PSs2b
qdaS2lKKdL93mCXKHHGfOSQUuhl7gzgn+gBp9JSwzGEspjGO/ws2wVp8NroqTGMbO8VxRGI9WRWH
MViO5fonpQg1l8+DNk4jKQADSCYgs6j6pLSwpuYD8Oe2LSI+4R9PhJMteU6rrFrh6ztc91fk6XJw
FBduw3LcaYRRH9YiOxo58RMehtzqqPOnP1Qyltp/m3AE5YJdlOgtmVMADe+MwuR8QJPinLTFIGTq
HBcy+vAzlCiWvQMenWqp7jThr5qg9d3Z4+ObsNdLr8QZA9VUmXjPAoTUoVkGuWVaNFJl+DDoKLr8
ImFq5iAOh2OJStQ10XeJWGNqKQoDZtRDkkySeri6jX3UBJto8WaedoYP9zteRvQAKSCRljNk+19n
8euSJA980RTQSQJi+Cxvz3AgBMvTdtT59OPgFZslb1meVNACJgqULimDYFxhvpzgEsqtdwtmgWYm
HGrdCgDKweEAxrAyCYjMPg862dVpJchUos6WqRiNVxawCHK6d0fGyg9Z9tE94A7hKlQSLm9WTVXL
qP3dLk/Hy03yf+g287AyxWLYcHe80vIojPsGX5re7JtakMd5PFp/sr2I5jfksO8caji8L6hjtuVI
kAUKngyymcsG3Jx6mK6Dfk5xAosYVQ9SHEsLowF500UHhdsAj0fDNawCYWcBX4y/WNrwJc2dqNyP
SG61tU2Jb4EAwwdGIidGLXYljtxRA5sJhgezw02RW+1IGGAqedjYtyCPPigo1APu9R37X7Su3OUN
zFZq4P4FfBM2ePt35o6tS+l5IaXWmzPXuwZu9TCKF0a8ugin7rrcMiNaDi1FVek5vPhEyB0dB7IN
QorLz8wH5Z+6IvGVmm0CIjrthIf0A8rUSiiGkwxLTkFN384P2ZN29cp34ZD6y/HptNuvjlhQgxB2
ulMV1vAE2J02zkTdVsIxreLCHcmuKhxwGN60mS1kQ3xlQ6wjoskVlWYMdFQYJQAF6tuxDT+tD0jv
2GBdaQSNATLEc3+ESMIimfEfBKtAXXMuhodxk6VbhsFigE9FFfj+1cz5LShyGy2a6lP0GMbZCsIU
ELKyhvu8tII1h8hUO1VtI2rGaEwObel62DZD7INlFgVFNQKRxrk59IoTBforU3ue3aFUarLez4nj
xzPg/UOP+ZYmF7XpnPRDK5CA9MWorKWvI0wTmVUf/jQWdsjEIy174BmTbNdoVgxrXljNo4UfyV9a
C7MccAEzB/V2GR9t4nkXDUcl49PutTanoyKWDXsn7dw6NPeD1It+8wSYkCOtuQ27/Me4U/S0iTCE
b4LDQ2dFmqTO8b9yDKLiGMb+2g2xyAZMiC37kil3QaLYb+8U/0ZeDJinRu2/t9LfqIuNHz2nMjsW
HOQfvM/XfYVEmLfyseJ3pc9BYwtP6KhYvHj8og0Xi1geBPOGKxrg3aXWeRYyNXcbGr392h5VApYZ
aa/L7itWIVQVpaZ/p42dm18+sBvW55XTfS0vMOrnVJIK7JmImq3IKgJ4wEbdGBFGd7eQfVl0k8IL
zL0j11CmAEdOquxFrm1CWHDV9MVcCHIcOoLB94DjgyrQedvdX/qzElA9FOtodYpzqRVEIczPEGog
uG8qa3W881C1CUK4atJZC+Qcr4NleANGz4uwRLslmtqsmUv4wZo0wkPe1JmJ3RHo/Gld1b8Bp+DP
WK/ItbhXNJyhoboGWinWGYsmNDvohyxPvG7TLCE2tDIfOfTlGpBAwzFNQ1VTOupCanZzWzJHaCih
3sVkzJxTyIBnkn0Cv5LxM5zu0HkDecGNaywUum0MQHhKA15GViQfVMCHDpa027mFUBGxqr77xLzc
IPMWFbncxHCQ6qaEU+mhaFPIItGOCPSYsEx0MEaIzkXujZpNdZryyc6LN9ljEqwdg4Z2w9sv1ccs
rqhGIAKa7RyWcJzrPq8yvcwSbpo1UBV2DCSKejomzHFtEhMf/lny6sReOzFw0sLk0/ce5SpExYFj
sKiDIGaWq0EA+GJpCfmg5Hf5ZwfCGA8VMTfFEEiy4BcJu7UmIvtCjK0VuAtTs4n7ICo/YhN5OmKE
xR+iiDbbZmzJbhxsMWziwtYRERMUdwQUwRV2ocaqR6gWMw00LhsnDYKSI1EO7HUuD0/1gULw4fhe
o1Lagj0dwI+fzOnCeEFfyk+jJCNTxHSCo1xe4yCT23IZso+MvL/ttUWn44CSmb3jBerTbTsKxm7G
EDkNJBuumRLopIdX8prl4B3eW27F4wOvHEVEZt7fdfVqXoZStZCZjWwTVt8+YM9WC+0VkcFqF6si
iRTuiv1GkjfwIjoNVysGnWwBT8zf6vCGVVwt1DzvKJWSJt2c9iE6dcOqO6UKVNe75/lhZ/irfQmE
1MemQiF54uSEVwgOtzCZvUUEFAM1lCOSfQCmIXTVMvvfQR0L42FUU/B1su4uIEIgYfMr94ouvtZx
uUE8QjfDhahGDGJ8+Bf0U0RVz94YT8pQW61X+BlTvTH7xDsrcG4Ye4JTOJvAXgpmfeal1lLu9Jpp
yR+fzzlWpGB4BGbmpjOdQzWKNmN2TxM/nOYKxwU4RHGmWPFrWq7KqV+A48iT7Fjocbotsssgsa43
qCiiiXG+H7nF7lc/AGXq6EMzfIvPlesNlU/A0hXYjafza441NPBqNLAiQ6FwBvuNg+FloX+AF9M4
kc3hBF3MwN5Lq0vLSxIak0I67vpQicwc7+xZCCQjCsBvl+QIorUUWpTTM1MKoa03R75DKR8H2eqb
ZNY4qBuxXXPm6XxrFQ021Yp3WXLCWncRlztflr7veDEtaQlx6TONQyzIAgollEhZv2GDIAj00/tc
8REcDvrKJIoI0ycLC27IGElsbumGHKZ8VvPQsfi7A0wO6gkmAnvzz2TKMfplf32PGqrXzpU4NiXm
IhhnD0IdXuWD/wN2b7aByTC/NZP+RyYkl8E3i/t8vzEQRgiYX+asK9OIb7GTTo+DbQlzuq988HrU
6ILoUpzqdqhhw5aCyGZWJfRFYsuFyDSWC0/0jX6/B0vIvIA+uy7NT536RMOjhQfVh0C1jo7wtJCw
AKUtMjksSpA8BjzDUnnPlyHDHLfxZhook0DVYwqap2WP0RBZrWLFZv+w9gRLfPpqutN2CqLjQ7aZ
n+bFNU3sB4Ne1xpoAdjvMaFrzfR+EPTcIG4bE3FPlHDyNhPdwceSXyYuyg+YKQD1mVvhbkZ7rYu8
0cQto0bvzzBhUc+nSh1eQt4mvgI7pcWfTQQxgT1W1epMV2V6MhIBoOGCV7BtCshlG0AaY8ztqEjC
tgGNJE6GwbZRJ+Z5+6y6865+DGceRRtdnWjzzcenliAheJK1QlEMczuwqgb1aNSDps+u5NwNu2n7
5q7yv07ySVpcCbHJlEBfsEagEvSX1S72oC+rsIKXmkQ/hiY1lqNINyMoPyo+LM+fBD5sZZ5u395c
xdSCUwVJaGh48bcQMedSUUCWa/4avmDlReON1wkKsbl4sEITvM8VWgavcDhYNx4lmgc15jjizEMR
DE3AW9GvwryQa/3+I49TLPilTi017bqNGjjFxt0wcn3bW69LOrWH+ZkxQIKKBp2htYTZZfWK61YW
fErcQDm0inHLC0c2ffNVrSIT1IxK+cGPiM9C2w9pkRj+HZdGexHflAVxrZw4iNkDiLGfqKF+QJbF
zn9y3XKegvCHz/i5Rj/J0iwkpaOL+BNRikam17AEou2iL0pj5ttWpKScnNa2p2lZHLKU7JaXtjhl
6dh8lWnjh/zHMe1vtrdqBoGEIMF+4u4bZGPa5+mYbb9I1uiBQZ0ktjTv5eZYDnzbPiB8NSs2qwBk
rPqvWwKHinWilhRrm7f9WVXKvyh8zAqobZFfhf6nSFOvhaDhQ1KQUCizgL5tmTXnL8pOsNtw4SYl
nNyoR1tnF494goH5Th/GMRQMSjuOJv/47uKLF2pPuihD50NgleQjnGkpg5npTyogsAWrjjn6jJ/s
xyBF++r/tdLo7kNdi6JYnABlDwTeVP3X+NeuwKrTHPDH7gomK05oYna5kKVn7yvbY0lHva9kCF9D
wMPwStGUgpvpxhT6ulBAjevchmJOXG+oQO8mN97wV+fyEPutIc02gWebmkrRldaLAjOtIv2pkJrq
03CH3zaal1pvKFIKQomKUWpXt+p6YQEw0GJeCrmWxuaOJwwYLtgEsyDnh1VXW8H75YBqJpT7uu4z
7Yw2dnJFlFwXVkwZm26Zgq+XmPl8JmHScFo+H5nDK0K8xF6u3Es6/GKQUTA6nv7zn1pEzCMCRLjn
ZChefR1f3gAfcLu9HjrqHTBi1zvFXw6m98hddf4q5lsDENs8Ou6RVEsRN8MOY5y4s2qYespTue5z
k+lLLzs6Jcj/Hh4CT+NPXz/t9+/gRAGhfA1/Z8dRg+3FmQtT5lHRKxHIdVF99ypvt8SezKzVsnCi
Lo5rMIcKaXC5aX15i859Pb67VGyARDyQCgjencClLJlYiYhzGKLk80M/myEG3FaJVNIqB+DmaTe6
pJeRJ6/RLzzPBO+xLTDfi5Ql0HIU5kasttOczai9iv2uKRxr1hnVvu3D7M9fVmZY0KANREpXPADb
gQS2p2JT2bYAsi0Rk5m3hJ7oF080Rue/DQvbwpB/XPzQwpZf/H76BlWv033GkSzYg5RvnhYrMCV5
I3iX4498jSLEBfrGNLVl1SkfnNxYPGqqJjlIobWj01j7Ky3BC2TOOIQf0xnqMYEmimV5DUygjUDG
8vQzsI8FIc/QEexWopwuQCupyCyLsee6z99NwC9SJWxdYZxecjOBR+XBMw5GMFwrigU6lMXBTAFU
vMHqSwjm8j1B0OpMiwB6C/a1gW385eh1l+KHjwBTnR2W3Ed4fvCXArVGUM6f/DMOsdpxsdVQdpSy
Q4EcxR+XdoWWju3Q3z9q/h4QXL2Jdb0RkCxRpk14+8NqRA8uIPn/KSlTaJNT4j6qDOE5DhBDpwAi
Ex0rVdzPKUKK9B4a8Lj6xn18oOKJ7tOqdJAbf9ttck8CArbZW+f/b7ky6+7PXAcF3AmLBJI9qP3E
gGtZgSofcN0X8tr5YHq8hoE5v2Bl1OIP79sNB+bzv1hAfgpCs8tVeSEet+USGXPKFKB31+LsfN5t
clqn5oXDqFmNI3H1H4h3DfDbLIJXnQoqlmfOdTQjhy+7RJyqZcTDQuram+6dcUzgaY8/K/ddnLgu
1+CX+6wbQjl5V3YZdwZ/ct7h0/MXQPGOc7hjS+4DX2LySKPKmIpwoTbPSroCg1YVMw9F/z4p+thR
gnljJPOBzjl0F0LEAKxFLUXUy0jzBroaWGrEIyWrM5r9pka9czZ0/V1qpcTGmFLVhmvOZ3i+Yf67
U5Etocxt1an9we/jyBF3WZTvysoTIV/xd1OtBCdA8ZonUhotVLuFZtJp7H05kvkJdhEkOS/IswnA
xRoyvz/3Z2xnIQT8H3294DmJIDNAaZgmpPdBNCGkipk5TH1WwBp6fj8+LhCKBwfHGBco8WWGyy2Q
SDbLE4lCI1fW9/GiWFVARVdpwk2tyir6MvMV7UBLRrIzu7SFk2/+UaCR5y787HTXt4r5f51uOBQo
Qy2AXYnhhNrT5Xkdv1Gw6Kg1rDzon62B5IWaBXxN+YEgVz4Pj8+UeQ+qp0CAkXZ7FN6shoM2ewwT
Bqd1ToDa+glF30QWKJgWYgc6OkvbVk5VgPwp1EKwEPlIpXRXCreGsDwNPUWUMcWtwtuNXY5GlwKm
psgd9UFm/NGHy9ie51tXEMNEpKj1MLKj2SlZC7kbrvg3Y8TOCMC0xgnoizV/4Q9zjXLThxBz8IL9
1lU/a0WyikslgbUwP2zmWQoAX98WKS849vs0/ePg34wxD+W5FpBp7sAvJ07sEf+M4NFDQCtO8Wqi
spaq657z2wAAUb3bB3TUu3f6n2MYMLeqtRJhKdupsoSfDw/C0H30x+6o6LhaSGMJyhG6FmzzGEun
7yt5cIwFnO50TyOO61cymah3KdE15RAT5EZd/748wKt/yeGzHKuIU2kk6jloyD9JU3CprichweAm
ZPisZcAZznUmHuRVCc1QPgaxVLOCrsFMz4ZSF9bxkaoaI6xuUUtO/ZFsgMAvsaWPAIWxMpMN8u5C
Kc5Sg3J9gBk0eW9dlau4200B3bigYCUyBXSZBdkdzTne5f47zSnkRFqaOT+LgX9hs4SOTgfv8uqk
zNDZmHtag/+8JhIqoIP3t/hvwv9YODUZJ2rU7pbas0RTZhD9DcEty2lcMZaP2GcX+9r8a7kb4yJv
+09zSOv0iVxttm3FBMso4lAqzN+kbuHkCldgnNJH4+usBwlgN4a/E/VtB976efYgEnfb2n6t4a6M
+f7jsfLWc1VyJmeJ30zECPB2Q+UTBtDhXlTnloH2oY1OD7Hpcpb3ybYUb3raoL7tIxnuupiozLnJ
z7TUupxG0wxX8Kl99EKvbFwBCV5NLg2RlrnwLbAFcuFHc41YV+3PRcFJoT8BEKmcrqzdD3VticmV
PShfGiw0w1dmFHvVHMPjKjholQL71D+iEM5D94DQKYdgfuCcLaSn/tybmJbHJrqwvKe0cKRpw2Gv
TvvT04WMKMk48vQrOXsPSv9GyJXOrmhPY8U/rWknujOd8G4LFOaV5U6Eidzc180wZ0P1WxyJxZne
9bAJjNZ0sbKgURf/602zjT/iQwtZqQdip7L8yAIhovbwYzoCuOJ5ooMxgZJq00ywQH7OwGfF+oN0
vbOhifpZrKg6ZVvu34iJu2tWuGNA7duC6avl/1O2sV2DW27qmIW6iDE5rjSpX1Zz8GEs5A6jfLuR
1aAyCgLKqSgIYQcELuuTqOfq6lAmhu23BNIRzYmmCIxKjOySqcEXjBEB8je3lnVRExCPFZeEjQAS
3I6aBmC/3aesS7Za9lrQ60oyme2o5z1wQAU/MP53VqZUafpOCPvbYM/xuo20M9yjYfUeXRuR4j6D
5w2z3PoAB2Lsto8V/EuY8pqv01UeTK7F2rm/t/XF9+dxU4TFRqu4loOOXmxhj9Fvo4S0EgwerUNg
On0xxcjqItVVlg2WGBIr71r0zEBdSWSc05A42t0iimHtm65hIvi0tw+wOsV+/+Fvx5q5J5+sq8vk
5usZ6pIS83FGDWZRi2WEOqUGRN/rqgbRAhAfRu7NzCUujLb8EkUQmAakCTvu+lro+BFpHihGxoOH
iIce0KisZXyaELMPLd5wL09BHmltIM+omOLIthzpOEcPwuJYkxr1/OAblEAKBa4ZJiNPeapzcrlS
nk6+k1Eyust6iOWZZhv72CNpRf7Nm6xLyG+80EJDUb3ay+HQNoycNUEg5quFe4MGGE4RROpBxbB9
gKe62S/MKLNEKgdYqZEIvfvPuoYQ4mGRGtG8Vb9JYFoUM7f883TpITBEoOdvb72u3bDJMrP+JDrD
D2hUZdAG0QSzfXmg6NmDF/i+r9hjvs/gJN2HAvZi7Rr3Z59sRkJvzUYmaK9Q9f+hFvy144gE+QtW
0yON4GWohpJDqqBvld9mQTAu7Dvhmi4CzfRW/pHoMi9Xu/XbXwfEpTWoPgJjRRpTNLklGKIehx9F
tBGiI4ihAllXzcH0vRke8cRP1JLiYBIfuly85xP/p6j0Koh1YW/G2C63Hf1/9k7vJGuieQGz5dsf
1GwHgN3E86ar69o7rIiGbpNFqvimQyl6YqaDAdK1vbya3qBzJQZgLckZyD0mwyESHpMhPg9pTpDb
NHqHJoTvgnu21rNzWjrz17dBpOPZXgrpd1CcgE0LYa4RLr5SCNhOIi3R8aDpry/Rbgr3rO1D/3IT
Dd79ykH97Zuux1fM1W/gwYh168yxRim218/4w9HmK4MVNPMcBbeGMUubvWcSymWZJO9iJ6lnflSh
p++yDfWG/mbtojsoahuGDULPRC0HQ3aQATEN6Agvb+A6HBpYZ+OhqjeIotZkARDdC2ni/UV/78sm
CMc4COrX7RdWAcLkw91XTODk0Os2tYWypMo9LzQ8031SI96MP08AAivDT8erM3/P2tJQ8raDZP1Q
W1Y3pbaWfGww4f4OWxzZnAYAEG3NlDsAXExY9LtNMDR01cC4HupxKMPcZyZyjnt0M0YUMUvwPYOH
wq1WoCIzO3GId9GfEEZTf2BJGSfIeCTbsleCOGZBMuCO5fKVsF6uDhBkF2wKnDeEhS3/1gIe7JAw
1ty9mX34M8za730Ns7us1mcCcjs4ITLq2s5rCBcci/pae3y0sQgyBSuKFNvqXcSovZkdgs/rAEjg
gWCgREqXuz88k5TH5yFFoHeCyR8vV1SwCwxaAykTgaZNVoZqF5SC64LkeXzPg+a4xbtkaNeLnVOX
GOEeDVkDp+eHASr84V9te0mVNA1TtgYmQgylWzbsaLGhmx+h+oPXIts5CK+WQAZPOrjV9hidAE2l
ZgTJQqUpou+01RO3M+AnubeAAbkME9xg00LqGMH34qI+tCqOblSCd506JeSDsXhDuDhrwPn6QsZ1
SjzPMkzTDiH/oD7//4lQhdC/B0Qp1Xb59Isl5wkfDl1+gtDVymIzBvj68KeXTZHkYOmwppIULn0d
SssAQhvOdhU6N/7vzdiD7dCPbb2wqH2r/0rpnCEvScK7rOZOlY6qkMambp8DDfhfPFPpfcXc7x+R
20TBBdvZKxZH24EV5KmF6ab12SFPe9g7rubVBQfoSliVGpPZoctp1rc6MQ/HrO2altyS5Nctld1d
l2dvv1kSVWymsvhkR8+pqNCWZ8BtOCpDN29JgFcSjrPd0JrycypFvD+ICpTv8oFpVvv+WLYPyuxg
eVwE605gRamOycD9TSjtzDrz+ElH35K1BAE+JL12KeYBhmg/9Nv9q6mxLoJxxKoId0zj80gsHUUY
Uz8TAxmiz2qlwEESWTOS/8kvSN1Ey65Hk2j45jwZN0HBKfJPdddrvO12Dp62kBU8/d3VL7glFJZ1
s3Jix7tKv9zieYZN1QF2eetjjwH/KYVpVoSKIVIaGfGXw4DAVfrIaDB3I+DN6ACFkPXh3k+3pfG/
dT/tKs3Nl0VJBZmIXw51vg97Fm5PCyGxtzt+cRBz71FUrM8SEsWm86UzzT6vDPzrIdIAkplJmFWm
nll/sRnSeA+zJD15h0A7m2lo1h1ItYsOX+eRBBY4OVMC4f++XJjN5Y3ipiIMPQeseGpUbFEe6pY4
1t0nFDqmHXMMOiZY9MITYSYYyuIcA3ftAsBpI5ii81Sp24v7gYSEQuyTtMND7EBASHlN3Z1S2MJJ
o+ZaK2YnF2mLfQcnwfZLRr6p+1hFMriI58PLxA276yHYuA2joINpc77aiWGnJzi12rVyc4ejFYPU
KcmbFEKERzcfQzfYCqAg76IPBWe+ToFvtfRQisS+J96jI5Ag/eluhbyvYCKMxHcH6Qx5ADR3bE14
mAkc9Y7yVWpQaWLtrmn2RSwdiWQIDSg3wgvxA+pMQplub6g/4J2a5q1Gt/hc+x6cipGvqtrPKaaT
MMfeps2sMGT1NPAsi3PJE3HxZ15kscNx1v8oynsQYc7Zmn1vSF0dh3T5OJpAVPl7TWORMH1S1Dtc
GM7YMdsJOHDRpa+QkQSiMii3DRifqgBWBJgci+NoPFIfpZ6ZvMxOMQS6Ay1sUr2Z/GxDMKMAkntd
1rCxFlytQeVkN0zcIj7QLlm/ushB2XjrwWXXFRuSZSlKrD6TEOKmca8WjRDPbtBOeWj44yb0sbaZ
pXYq4bF9e+LJngemvHKs2wnkP1tLR4xzgHiIEim6CrSjk5wd0pW77HECNr+/Jy4gGjUv4LxoXLYA
UcazgwNQGznjwvMa58hQ7sQrmGE/7sDy20yut7+L/dDMqsd8KbdSbH75IeYofQlvFDly2xeu6NS7
JZ1MWwVc3w0kRcKwqUY+RZ9JCNoBUhEEYV6/L38dNbFRJ7C49xRTln/fB7rky4vwhepMUWmHygXV
yTcjpCZt0whAYyebFZ236bWLiI3SNqm6WzjjYXz+IBHme7OajvYgVS395zgTJHVbwyrMbQPFPCD/
/PYNv1Tq+2bI9yaZzvOkdWMS0k7nHMrMsB7L/zx1ezlgUPXxQwuxUGcPWYJXMMAjD0U+K3uQrAVe
av55Lv9xly1yyEwIIABe9yo3DskAduPzgx30ARgpMJ1s49/P+oxX2EHSAgNPS9TddeuRD9WNoAyY
K3VNh+uJTCeo6+EYrn5mLhTm1RMYxl18uXkxCZ7aR5tyOjp7uQF6pw8dWLpeEQJB9O6BpYDzHU7x
4tKXUF0uAW1pWbJYU3kXxHjSM/zT/nxTP3nNvbLYkRd8hvlU6iBA6xgVobLCTjxvzVV9VLpzuxUO
KRlzdH3yYy3eTigCpnm+lDjQkVgOkWWXh0DlC74gF+gk2PrqK+330dwpxBp62ly114sN2gs9EuME
LTgYNv4Jl6kZEwSn7ADVAEkUu5B+/9QUgHpNECMY4H3k62foJjF8MsivjKeoFA9gv69AZEX5J40h
oEU6qrpH79Zuql+FEU1ZmTQTcFb0ryK0Gpj2Toxy4VUuFlqsgSCw8r/6UlkhUSJOfDKrb8Y6so0N
gJg9MZ458ePrJQj9BOI+MTcSIunZ85Rg5UxAz0GgLVlgG78OdTxjEYyRfEsB6Ouaz0FG88jzWelR
ZPAnuShaFD3ejMw9kquYQ65//GGw80icHgam1uyKrwXribzWiuMrh7ts4ebBNvgR9B08R6b1iVwl
JP/+G7jhs+qda06pHm8CpEbJ62ScU+ZqV2jUZ4K/LIP2XGXUZpeYRUThDhbQ5KlaVYdtuAuehZwU
AhfBjpYf+f6+v2QHXpL9ha+pmpxx8VsVuw5rQVB4es6ichSNxxkirc+9VFoXEoZGgrP7gcCslC1D
pCiOGQPU28FuCFdT/1mb6/ASd8wFE+8Z7p5ytlYy3Q20aAoKaSvBwHSMFeatTKGJYZFRiF/ciVf3
3nQhE++2nnJKiW1DCth7Bx9UfcIvt6Z8prjVi7accYzUQFJ5N1UBWdOYh9ov3I7ptcf3h7KxgSAl
dm3z1kUhPj4JSVAISJIMgincJzZwW0JlVJbkhXyTjCQgd9YNNf/C8ieQ+F9znc1FAJdY1zLrl+4f
S07oysTbD2M9fH9mdyKf9CschD5P4/h14UIx2VXM3B7xzH9oNxLJzAESYxbmLtJkEdwtISsWE0Md
6FTBePNpUMqVqlgK1rkYGAklTT8yFWLJCgJ2zRXExfTmeDPEOUmkETcmt4KX2ZF6V36cmEdIFB8D
jPFpzl58QRP98HaJjYXysWnVnz2WS9Uc4uUva3bFhz4jjeR//TJHqUvd7wwP2LqkfKVSuBDbdbrz
qTVCSr320R+3Gs2OG7t2LxijAkUai8WPzCY2bQu/CNZYKoqVWtuhdI2NsQjju5CIUfp2QbGTFU86
VKc1aNekLPh5V03pqyNFV1xjtZsERMRJKW/zE6XHJmyYXJGNSqnU5lMNdlPNNnE622tpJxG5EeAc
HMFB+KU55X5sz75bvLXKejYoYiwe8zRhcQgf1zOJAMJUQ8q47d36PaGrk/Gbzzo7aOEY2hExHgBz
xIFSis7dMJZaMGt7GGd0ewCbFxYmZzJcvgyEuexrTNavaCIp9z2tCiZC+RfpDDBe92dOIGMaJRL7
J5bc+0yeWd1Ix4RsqHGZ84bRjvWGGCTEKAoAI/ZQkVYOQpbRvYw2or/6igVphuYMFvkRjlbTrvSd
KxBgY1YjL877keCuUTYbxSGbItkw+8GF4qthBw3Ka+RUtq9GWn31CUIFyOK7R9RxhS3hjWe25J3k
uI153EfvrOXJL1LST+tAf5GqYQe/WRPKbrotiTGvcifQzH1YYzt6AkLVhHilPNwrcirIAh2AjF7a
ZiXZPJUnsTh80eupYVtjK0IPbLroH9p5+wQTibOt/QXmCeEkgszYxvf9POvoZHW+E3D33psZs3/S
aqFW60ek4qEONtLmrBRJNHiOc8BH1cLJANRulLcpHDfJXrUNynDEi+un1QMC6Y8K8eG+5OW1yMac
2YuTI1vxlUaTvg0Vu9BdxdM99aWQwP0dEZPXNmCst5n9GDEMn08Blv4w8w8svY+3ugXxP4IEIJMx
ufZx5KZT9pWTH2fe4AiWQbsiAP4hxP7yjjGiQaIVt8P8wA68nK9V2GaWghlm46GhM37g7s38Ob0q
tzXYF5BdHuew3lWFcaeYqLd+YfgRvQSuCD+W4hE7omJdFs27+cnMrRqC/qciHUJZWP2i8T2VCGkJ
8Wkt9d7l9Jaav0JlcDcBl2KibhT9Ew5PcUGIDltk78CYqOOjzTdjvkfdotyySpl8urwFyiSSNdEy
fF7EuU+XHuo0rkix4foVt+Q7aYlLVcGJQhKTEFt1PE9bv6B1rD9r/Wm1MhqTZ6B3plOki9T8+0Lw
FoAlIijue1I11hdZta3ZIARdNHCk16CPC8RU7KXYl6TXiBpYb9MnlXP+sUpUG8BNEnEO4nf6IDGI
xMEi8V94di2l4CxFYzsZ2mR034haxrP3vUtb3fZq42ZKblk+6FfI/ZRlYQ6EThiRM9wr42e4xqbV
RKFfKU6wvhLV6iIVujIW4sRnvjGml1ez0MqvjpQVS/i+oQCoag4853d563udnD4Z+uDYQjl7CWEp
O0hnZDUGWw6sFeL3YuXqDT+zPmvJ/liewbH5VpMi0rT9x5x6+DubTeRzW39lGFXSH+0sCNvIjHzp
6mZjncrqhn7V27xzxXHHrR0Qn3k4W+Eu5/4NWPnyZ/0wd0rOaxHvVwZdxpi6eAKVE7iplkfTZaEZ
hapmFt9pZufVAUtO7n5OKhuDhdoRY6B78DkipybGUT4+/zNxOnA9t17HGp+bs4dO+lIgMKV0gjLI
KIDK2YvK3yGon2zInaAD6lWvIHIX1dFel9aa2tJW87N8IxDsip/rvT+dbqsqEE9R0dhvgPGVQ9vI
za/3cbjiXX+lncerEnNV3X6fFo4HeNRrP/eqiL7F4ZBOmWcFNe+yw+q6Bf+UoyoqjtyK2FkwPu7/
dv6hO5mXhitOPnWrZgdp5RJRVr0eCU5UX6dRz7Ani1/owCiuNXthZFO1Mb0o53F24SwY52jQlg95
N8rxXgDP5seCEnRu4dchF5fGkGzlez/nAFPCRRy7+xE2XH+89wH7HXmrSszq8WyopjEhjt4MPgi1
+GNTJgnblX8V/HJFjUGpua7KISLakkF5yaz9AWkOTMIwTd+bT/rZUppIOP7lA7kdnH+5VVOsPluz
dPh48wrX711Km/jijnfB2s5sYduY3Qg+YxXhVIsp0PjJnjAg683lrN/ffgOg1XeECiUSprilSoD2
5L2V/J2GoQ+BlcnXHFI9C5R6MZKwegGC9rJWygM559SEbUJepG2pkDDpiqNnxAP2aa3mtynfpGbT
kOxPWLLjVyKhy16r9nZzFn6dS2TudhJvSdk3GSLnIWjiCl+DikX+Ge4avHqtCOZ/Dxy/gzdu7MGp
20jxobGT8sTtTI2Mm9oJJIEkk09h2/c0Pjqw/GEjW/Po++Ow1G4NlxYABcVjuhibew+ZZNs/pT/j
hFGkScKheGedWesB2lTgnxPEfZI1woDNDOsqlzoKn3vvC7ahq03J/b6p7SQiqbYu0ZcB4qzakHsY
csdskjut+1Q/dxIWhqW+ft3TjLdzOdv/EKB2qdEuLhmycAxW9TmT0TceXm3odbpE6Y8vbZOiyaTh
mid5W03yBLXHeOncNXDZdOTErBj5Pz9VC+rsI8r0uWzejunuT1UZrpOAOH5LJB1NhS/3oKsrFeFc
QQsdAxRUAizzIu1R2g89qepqSmaeXIP+kWzp4OMkBK9IdjIDMSaMDO1WhMQVM9VpVGMkLIEER9DY
fh8sHzAGlUPnxAjvZuM2+akVxPCs5pdp1GlMQ9Og+qH0Zvy4ydcPcaiPrQpPW9Jd3VzWokbh+XZ2
r7JzJRHfcMmvvcp4wVkFbCpmv/VatK1MjM7adV83Nmd6BeZ8BA9wHvJNxQ5jiK8hcWZPRYdXds5L
hsPnBrM/KbplAobGnbNdq7OYtiFDQXJl6GIZFqVQRBTtGlOdBd3u2z0f1wFLcmjdBqEgUy/a9Zxj
s9mIuRzGJW3eOmGs0PSQ2v6gQ3672CWAJjoAZ7kn9w5EjejBmvznHkfyYK4WhlgdC0sVRTaGLMuM
LpZnrVDrwYAHz11Wh+NnvWy8TpGICPhismtm280Q2w5QrCzWyK2pj9WOvZeeFyPceJJc5GTlfz/O
qkenRqVtkwjah6h6f0rjeaBNONzheO+YhnzZe7x2dbV/X0SPGupv5R39M9i9lPmVQ0IUbxkmf4XL
RBW1VxNpnkR3CZZpA4VB1qVrzl84AyeluuqhQGsen6RzMTYEEqGLS7hTYdLVVcm97wLjXLBVtxH5
HrCk/suHiettRy4uPwONoCpeyUt3ftsO6qk/CD95G8/y5/7gBxDw4y8ZxRKeYoy12htECNPaBXiz
rI6UegJSQ70L1EmsUUr/dVYfG5TWA347pRdaMSeNrsx+LtSEqEEEzkXKpLH6ArHkIAdwBh++d1BN
xRIxoE38mYdkIPgUq+cTuIyKqxZ/EL2WZAzDNJnlbcoPdE04DsuaLPfL3KntF6cRADkWt2e0QTsG
Dj4X7Ckt1AgaxuK2dsDalIu3zbFT7rMe3Zu8NCEKKE7B51KvMkJ/2ZJvzPgwbIymRNfvMB6mjPf4
fJw5Q5kQVOfN6kLwG7zP5z0hvnd+h74YlH29TyWDgq6l+9NxnuBp6Y8Gi4E2loiJb+B78OWPYc0F
lIWOzsi1ypC3JCnIeThJQ3ify8RDAHTVxD6IeoaNzAvtQoZfpV+4Hg3rVN9FvEeqr7p7wHnS8bCq
sxKP3Ig1ZVRWIqfz6kBoGiV1bvl6sijbLVlqcPI46Le+iYiOvMTmbKQu6sVDWPNJkQ8CdkX8kUYG
j/pjkoM1fq9mr2H5R/6907vYF/XvHxWs49SD4/kJ1agUgyFMTrULEctW81IMOpflH/lFXTae7sVl
NAA6UFWbep1vul5tPzaJkRSdhvO+M6IVXY14PE2c1LYbkbfMvefXK7vJdwbZhCDxIUh8ZANGJWmO
P+jaqZwjpZQ2rH9ymBqfkBt3sUcHGr1x/mim1d56razxR1fl1Ehuj6cdx7/+qVK7g8Lu1uXNiccq
qUJD6nH/qJVXIUVZL+77PauDfYBRzXlJdL8PdpKT6MxMMW9kn4015wjv48CDJyWXYzDy+7cbADeF
vt4N8hjqe2Tj/ZBhJku/THHWO8w0eWx60Nbg1Y2wsFeT1K8oU1VbaiUceDSpf175zj/XIs2pGaem
+Z7+RaFFMKGjz4UtGxDaBuYUP/U5RCR+qHwVeIHrKiQGzYRm7TeQ/PeOzzlAbIVk3h7sd0LLvEIi
9t0X9Xm/IBhoViVjZ3n85e5eKxaCKyJ0I/p901CIpDbL+q5g/gp5IIOtF3U7kmvd1rf9BmxORuXC
iegSIu/uWt3D+By8HvaHEmYaCEPEEQ48nQu75YkpA2hYRukmgnHIWeIuh1KklgmxqI2mR3+TgHZC
sp6xYadmVbbEYE2+I8RIqX22oKyImYCFBdGVrzzg6vazSVEaFWbzYVqVfb5F1ud/uLHbT6zgEJjB
pMgH3fviZYDrxQB6LNZaGN2bWozn9XNnWkSzevzeviwjlYBo9NO6Q3DN8mjmc29LnLQPSM8SJedU
IHBLjLFFJ5zLbJ3BUYDUPkbNVFavgRVquqK4ZtptBPOctTlAlVuWi5LTxClFt16BCBGaBDCxjNAF
5bIJ46s3hjmvDMldNL1hxXp/ZXDP8BDRaWCf+pgEUvPV0G7Fp4N1L2Y7Mtb/0jkHkZKcBjbeo464
jNcZG2rbjx+yvaCmjpXch8LfnftmvahKC5BSmJqy21gczC8VGL+UXM2nRaOhWvj2LYwd+lFWV1dh
N33CjMP9ZSyHSYezoK+P0++Vcj44ivlvG6j3CtAF421ce+tI/5FG7Q6ua35eHiog+TPweuKwBu8x
vnS2qDPQSkPkOSCgILCOxEwDOJlDA+VtLwG9cT6T5KL9zHgyjhuLxFW0BUTqnEc6WBdFW4y8m47D
eGddI3XoLDsDm0ZDd//8XHjO/d1KbVdh+nD/ntsTb5bnLUhZnHXc7zwbX9mvM2/sfHgYaxlDPArR
j9kqGB68vKVGOERdEo3MHrRud2/bnfGYszNAAeJWeXyb01Uq51Yzzerj6JyWqGsvEJfPbW0umeJ9
yqzjC3CSs+MjPyeBxsPgYNHhrW0gkRwF0c6Hw9u8IjZaa/k1xYRm184FrFj2AL+EL8ogqn8z+3Wz
vY4B/fucj2IughyboswheTZ5rfy7ScjaFQS5BmYM2x7tqaT46RVVHT1pCDUpAVBbXzpHhXGMHlhI
K6zYAJYCffX0XsCt99Pv2/RubFN3JZvX/Otx72r1wnCEihpmSQOqyoFu09RtfYpWu7g1lweyxBM4
gZBx6+aja8qUjNfgJ0m8B3vKOfDmmygOGU90vYknBa3XTOQAYdQppfJpSs7KpnKN13W/D/+z4rqr
ZjeIYKAE8T1BKTcVaeYHl/znrG3STKKPsiUk4KQOZ59TL15GhNZC1juWL28giFcJYf9we9HXHeZF
ZgUOll/oq2y4F/wtCSkL4cjK/xF/hjwZcA+ldIrXdMgfu+zwCR26KaCvYRiGG5Q5bGKhcrd3pkfp
Qi0zcnw8Vu985pwJG83FcN5IEETWSBvNbaWSnwvt7zMnzSJ2+noQeJ1247A/fZQA6UX6T3th1JHr
9pwOfQ0iAtvEfJp0lJVRtaaY6eUF+rVC+ZDYjuadH8OKH4ZtwzVrGVc+2CWQXZuhVkKV766lAJz0
A+8CSvBEmefBkC3bTFYOnHQwypNTWkXV3NdTPb9urNdmsA44tQrEynCAXS/lfip7cI3Fk9+BhTsT
dx/l0EImnavYbBQmf41wWX/SphkVYeD091mbG46VCQ8gfHUmJ4Lax8iuWfROGFOS4SZebqRzYP4g
pWxqZsNaoz0FQpkxHxVUWqqnlK54lrPbOAJ536A0sWMRrYxot1PxzT7Zdp9dDUHkhlzG12RJ4yqF
gbmuOQgsDF0uuqrKq3iE65CWaLmUD9+TvpWPnjy9YhPsckEqugzwTCncBo9KxK6S6ADKs7trBBdP
qbnnWdANg4GBXSYzoZvInqWULCSY0QAbp11zFb83dSCfq5MlNNZjBaOSDHvV7vIDaK0k02OlH78V
yxqkWtmjjRRgrDf2teYiWessTJ/ejXMnYU9OfTSAUhCsJ6UcpTethWuRT1TjVVM2UuOXbVxKYM05
lMJXHeHGBvFvoCPvWVC8w4dBwGJCqR+mDqlb8TgaSs1IoahKdi10Fqy9kXczTad32SiYzdumJ1Kz
nhIy/n8RxvLHMG+YepWFgYbsNlqSeYLtc1v0wIkH7/+YgVm9Fms9pXZJ+iJdhHQawb3z2rKpZvjD
ibYCX0TmeeBI1F1ZMzKn7Z6DNtK5VDq36Q9STslauUDC0omkGszM23gTSwEBY5BvdboDZ85/thLb
mqoQw8V881PQSdxWxoF9tgfc3p/J8dLcWrKpTnxWfWnTS619/zBZIe7ygafXOs4gPFaJ06Yj2OMH
2sKwcO4s8ScvCCIWCC+D836zmNtXrPsPLdrQdoqIMd+KA7r8Ds0Luy6Xnj2Nl+2OdWvIaroaF6kw
1urDzvre/G3B9tPJmVRj9SmGFfWuLZhNsMQlpaVGGXRv6Nlt+rWyDokKMRrD/YYXivj/G/QNmwfJ
eBrSf517Zx6zNrv6+ABOXosO5pjaFaFO/v5rduVqVkxZ8WgGjAeJfoLQVsLX+cc/8PmK9tfiCsT9
1fVx8zxK18masPN5ChMfLiQY0bswKMS7LAyU9OIgD+W4S5EqVfZE0v03QfG0CuZAG23d3y5vqxc9
uyXFK5gp2vgzfEt1wzlSFnhIfeZGjLhDliGKDS58BUflEp8n5gO3hQNMOAqk3SQgV4/hOQuv78q5
t1ikvyMLWke33ZyrTHGArSdNMcMb2d6T5+yqE3xki3tsN2lQ/4RAKJfDAxtlDlbCqdW8vcSzXN3O
HuecDfw9lI1KgZGTwOM02gWnDNwVaz0Mi9o+SbocnkHp1tnJu1BUCwrSn7TuQbr4NuMdoT+yuupQ
XYGAhSbo3OIo+i0E7fXZtBa/Jd9IBXUeOHq224NuCO4ylE9hmhunK/X6s3B0iFt0tneGAblh5XsH
ATgJL7yVPOQM2/XglDF27uTjtcrCbNPTrRoTXkamFnxaDpVICH6jCIQeeKt35aOh6Bj9PmOae5qC
X845HobsRHfxA2IGdATib1navhUxlm2YBYq9IfnlGeD/1VFV3d3fVedKQ1kvyB2O5pTHmW66YIfr
5xru2sh7A7Ql6yRLpn4OelH9BGlvAFOMzv491C9ZJaLFxknSTbeYICawDVAPII1HanV0CFM6/vaX
BvqYpEWrpTzaaRiQm8UuVGHUTtQyMJHPpI1gTa26nPGT6zDHFupJKDIl+tEGRMUsNDIdDPaFVAfo
e1iG8I133zm9/BNRs9rEJZRdOSB89Xoezord2oyi63V1qFYY46KjFuUy/NCAH3WHkj4XzdxjutwM
HMDyG+RZ04FdSJ1QXClp5/ZFk+R4NccinGeO+vdFmxsQF9smS4mDkl2M46AnO0ukRM0jHMc0CrVK
mBc2gfPCS39MJSyFW0YvuwqOF7m2lT67KIZ3EShxqcz4H8LgiK4veYSrqwqvEXX4ecVuuL2FmdiW
G+ATGt2mhJFRS06fijD16an2U7VLbNpFp1fqPcVPDU2UApUdEVJWQEffmqp5NTOZOJSeISNG0nwI
sBCcREbBD3Wt9uVYHzjOZ9dfr6QVBAulx82pPXlOJ2F+LcT5i++JwhFAiS2pRvNOP/q1IQW7vE1Z
sYbXYxx+SBZ32k7PYZlYVM+OyM//SpEQd1/rStT7gvlBhJzJ2iGXDzDgVuU/yYmAOpZOIV20FGvT
z+DVtdJYKw0BlWrxbEvmhvk6ln5l/AZUcnUFbBFVJpZMzE+yP/GmprRdRmZD1a5OPUCUFt/1/q4N
YqLmxXd9fPrTIUaJ93JUwqBj05t+rMDyg8jONNdxKlDbHkmzo1B723EbWJG09MmJWcvptTun+Pqs
rYin0UG4NhcTHowsQROdxYF6WTjksjXwkgvY1cgKsbL9xERa+0+jZ/8WHEMpZZN9UI/i4PvCIxmR
PdkGIlUZFxKIDY4kfxjDrlL6jtfLP+8d15jVBxVIBt/pGVPodYwteBDYixWkI1x3acGAlHpDNFd6
TeDmysQHYnJtiyTAHt9iba5NFp29iCQyrUdZViiPDsT4C2Tuxfv0eOS6mZ4MQhhtd5NQiR5vvWd2
0P0T4oDQtA6jzmLZf+WJpm/SyFPv74xlto5UpvQh4CY4+lU5UsNmGlFge+qyJgd7TeWL6eHdxp9j
TtxE+gug5EA3ItE/3QrTJKvz2hjCTPn5Mdgcf5PioGa+vbkhNdNb+O08k+0Xwp7Qy5ITAT5orB3x
vD8qzAs6ou9a9R6+wG7pvOKZwpZk2oZyZzJyotl/P30yIyS/tZc8yJXUvFN0fD3qoJ6djO0/2cjt
m36z9+JwuQR+h+j50Kgij2j+dnnSqSxOOmh5NLya/RHUOsJAbyESOYcjPBWDzWJBmsMYaPCNw23q
Kp0cp1yiFpL6qFaMbto5MJ8GOHsyQ+UDvswbO0mgmjENQH8LPVz+kzqoE3PT1VU1fBpPNUmAAqmL
6xwdMR5fyFcqGPQqIBbIbAwJ8R6z4qwa4iytz/XeQ1q0QuBs2cDAyCrZtY4VTWqjmlnoHkb6sr2x
0qabNFvW5shKSyf41vVj/e3jNjfA65+lYpYeTpZQcR4UHFQFnfX1gQm8vhv1Dno22zRKjC9g2/Er
WYdkAui066ONgOkJz0sgchd7SvcLGtayifPprTFDY52cM6ca2hZGl7vwjx6AtqCwNXWdVGaLh05A
uTzujB8DJaOMC3SwxCgf1Uf8mwhrKDkWq/SI+mznNZWghPrTX5vPPSW/t4tawxVpA2t/gULfZoOZ
Joif+aFUtmSN9UhIcIxi5IBwqDZZaBkBZyMAxbKMiQBYNSYmVb16hs9u+xP9MU7mmNpEXM1U7hOp
ZDDGylZ8KkOqiu79HHAuF1ntbVzQgqQ8pjLtLaR+h2m3ZmdxA7OqvTkP+UR5uiYPBnjPl4KoTSOj
r9u25mCGLIWqkxEoxPh0YiqWMuEry7syWDIcREq4X62kkAMMg9bFmgxfQIxot3WXeiLh4PsDE0TP
JsGVrF3Lnhy+FOqQID7aLK824XwLLP0F1d4Vn/GaxyKuvqSas/W+Mj4h4yMNgCKKP/C5xlw7lbj7
VOuurF0/oPITl68VjPB80s83eWPJ2qW9AjcIozxc6XXriw4/UbmYTlWd38Gon2Ngz2SjTeSFvmQ9
YD3qnI60gVXG1HpmUR0Co8RGvwx/E5Cfb0tNHAALqI6MVZ9p7hWSyLk7V7te9Pv1MUjtcvI1TjG3
kNuLNMyXphggGlcZ7VKWJ6S9Zw1iUyjGpV6km6FT1WjRM9G8aKk5KAkYZh+CouY7lICMfdnan5mQ
O6hKMlKsEHPxpkmaeeNDXzY5Q+OA36GX2pqFOz5hH9USNgGWT3stAbbPFI7LeRa6cQD0yyhS1DlH
SDyUOdSLEoQHinJEaF739rzHFJF7NV4aVGtLhxjTZF3UmK4Nk7pU4/KgkpW5//2xpm4JuRPnNhJH
O3uBhdcTwP8mKKrrxdw0toqp1lE2q+GdpqlIJ5k00nP9Nlc8gB5yMGxQMrr/6PV8tBIdM4R6TWvX
DQ6/u2ZhXlQmMhF3C3DYWOIm6C7tBYpzECKpTwtcV6aJTIxCkbJfM1ukeFMFOBNPg2kH7vzGgOhM
Pm+mcDcCzQig/A0kBcWYP9LGN576LMp6wKiCvzqUK794ALXbvTAzCj2a9ikVgdh25Yt569yoi++f
+HlfzjrMnFOcBRxn3tAJ66xOIal445dn7KuQ7nYE5oKLfA+wI6B/PS2AjcziRMsBcXDdPmOT3MkA
CCX7xmhM62Z64uqsTUTNAFJVE6kaoT/W3JpJFePqpJAMYx4Wwgf4ke4eZpT7H9nnf7RczFyBLkRA
qyKKi/13yaLWfKQK7fylS2mkIJpF6jml+1QnsF5IB9VHRRoF2pZXV8GM7uNDeqrpGNmsjwsj8nNr
NlGOAJSKtorfvYJV8IDt3ugmxeJgXbzJnd2zknPx0UnlW3tWORnT9I8VUo9bRGEJevfROQu2NkUs
Z4jxIl9GH9WKiup3WqvOCJk8pA4Zw0sjLW/AcLixASv3chOxDfcBILns/BoYdVgJthPKYij4/slx
3wl0xm2jhmu0QgGXzNqM1mO+lN8arMWGFD8BtoX3tNBgBiZWobSZnoInZTAgVzsyvaNnXoVRUrbN
7NqiHB3IKBfHb9hpdQD6a74VePKZyp45RoQEEaln8qDMa4JvOkYB1O4c3YcdTWH2Yf3+vCidzFBF
C4YuVlI71GFfMn3SNQnNxZWe28MUo7hP7OLQyOaSC/xrm9IB89xZiCcNkMs70LGTOmQ+HR5cnWTc
VvA+m9HyF5Avbs3pvRHYshYffTzu+Buul/OtQHdgXaOLNa2IL7Mf3msak17K/0mYVQmPzwXA+4xP
1WlXn/w8M2xY7BeooRY20F7Ive45oCUkJaOn0XNS15U6PEHFcCitUdyfhGflAJznKcoVEE1iyaus
6Ihue7JNApLY0NibgbPe2A6+9vJJ17VQQBhmlnfmnpf6gz1HbC7V0PKJX4ZPSaAboyD17hmGAe1m
pdJxSNq2TWSYkkmO9WBKlgk8d9Dj5rHKJf+2kL781utGAjvBVNqSnd1UCuxyP7+gKK7qU3P319+c
DI9+6trDKyon/3872sotdvE6oDqh43Qu92M4alAaCyC8mFgGoZdtRWDaX+guC8YebjSSLUemPE8Y
cjJlNkQafrKIe19DfKaVyULN26ioNM9GlIrfwYF1d51u+PTZMEL2z8bV22OPtUoDjHqbXUprdQXW
u4KUhNhD7jee32wIO+QB+R21WqV7wfnIz9RxwojSz84HD6Yz6ZraHxZuXDPbA1fpJ1R6g7dxVBOy
tiuOGSlfyaxDUsaayD4Vns3/59M32kp1lGyiNmYXuj7KOVOqal4B7Ora1ndGEESj4rKHOUhXRxi1
zd5LoEPuLPpymM3+S03kkI/CI/rY9MyzZqUBodSCi3IsRrgeUuWZg6uBntaCuBx7upZMZuUnPcrm
hDu+NnYFxH9a3j/BwbfYKaO5/2OTq5hciH5MYe2TTdwOQzNNYsjOl76YmE7mFkiwhQG3npqPwdla
sa2prCfania6GlxdZuTmaisfzTVda3ndwAjt5jCNST2CgBIjxYA2Od/axHpLtLdiON/O4ellCvFf
R+HBM8PEIO+MEPxAgs8gUbi1xdFQ78KglCaRpjV3YCr4SuAX5Ewqs/BghaQqnJws7MqLDn5X9VMJ
slFn5pSpEfwUDxOllkW7Mn14nsBs68JMI1fDCLXnGrbv/0wk+Pza9q2zWcefkquhEyfwyUggkwBk
AKvv6AC1GzZ9VPxj2+QJ2H/Feaw+8Jp6KaCgpXnFIiyrcxh65sc2g1BQjSVK39iAWWnNl3Me3CRu
joyyYDYG1wWi+ka93EDjwb9mOlR3eObuEeAqrR358vKJxBCJtzxa+HipbQwfiBe3RU7us2+M+27t
m68mFsjb5xe+WuY6uMsKbTb5/j3Ft0Lcwr4oDJ/UWi7G59z5jyOb2RYnP/NfGaweiqN/my0D54SI
Y+jrrlDQiZ5/i4sqZtYGtrtwaf+KaDjnCVev3lbJguOPCI/S/QWPbb4PxFRhyw/ggJ7kI+EUo0B3
BX4OjFV4uA+zYr8SuBMt5TJKMKU9E5JSpU6mwSNUca9faEnERmyW9lRHR4hLzCZI/oCZI3VtMivA
uvn3nEyKXoXc2XL4bvcpW24q5tuA9yn2Muqfs7hrtHXETBaYzd9byEvZQuBk8ye+4isXyFkO+943
FPIyNh6PJpxLsinjG6QA2gPGQbwuGNCtPrXWlVXeNqbxKje6N4hgJinLZ1BMLZxwClFTXnVP5lIV
07EiiooOt+jp9NINRBukJwM3Gn9fLEhxQniD4bjL8KOCpQ/9MCI5TZPgP3RpDjVORKqiqdIK0Zo3
aY1rh02uxMqoOs1UnASQ9fpLxGrRTtsxdqpBCwu8zpBM3vh9bTzRWLNTLnztWZv82xSExVzEVzpd
hLtvP1KXYPI/sfVtZC+h+Myv6i3SIRfRDn7ut+ZzZseXhpzjzk28TnIlFW2yYv7OxBr/WDMbv1rO
kmidbuG2iEtnhIOD6TNoVBvEWHwg+a0Rgl8tgBimKgOE7GF+Ni8G/bqimmO9zDwxpUu8uABOif+E
jFItTGkhozhWGfBPe1M5SlQ/xKurn3QEBK+CjQ1WiNmC7RwBYZOnGFxp/hhbdPViNyKiai9qdPwk
AaV3Hk09V8gX4Nreq+YjcWU95mNACVB2jk2u2Il8/LgiYAAjT55j+CJnHP2EG/we0ssBLZmHajKJ
4Escx9UPHsfYRgQqz7KHropx072WiTwo9P8OmMdt6dT7n58oXlccDRqDEiOZyPdKeKrE0Nrp5jo1
Zc9Fut+urpeozOR+VzVNio/z+1tLuZeCAkYJZ9GRnK3qBGB4GDNjSmBAx4+RpeU5xt8jDYXm/kYJ
QhaKp/g2b3KnVNG5VopW9GXZ11FW0fdREydltsddpVl5BQQWxNDesZPILljHTknvewjctSCGMxnz
CsU54wY165qgxI8DQFS6QStROpbq3NIhMWCt1nQEhUcmlfZVvNdUGiUt6wD/c8ET5ilwmSNNuDaI
a7l2ERI86/qHdi1Pyx58GV5rMaO8p367lRYd1vI1GUm9bIgBWoQLPmOXRFyghw+xtTnCCKZ5GW1u
AJMz3c3Lv2okm0cxMfMj48o2ImFVbu/XHpWpUKSif7QDGBR3QwmNk6HkzOr2SAbGYkhdjutrCJvH
uFYJDsTKD1po1qpADzAleHf1xoyOTPClU4O6w1z2C2nO+zGjVbGNi84Yg6LGj8N/ZWOa0a46nX3+
K5yWmhuGAqdC21hJYBjh6I247aLCuAJUPFdchGBI9BzYVmIOe3myIXnER2omXme7Pv5hG7NogMH8
yt1DHpc8u1isLuMHCCBqhWax2ffxbqS5QqiYo+lIaftQxlQDVFiNAhAnv6p+HMMkSVUBXEvhGbhB
0Lomx2ikoZt9wUO0DSpOCRlJic+PLNmvTf9jm71Pycz/Gyazo6zdqv00yCXOgJpxhcNmdFei1/a5
s2nE7XNsG1xTjMfxCZKJJe3bISrRYFTYFgo1IJwtw/miF0thQacx7nrFz76KgOP7OPE9kSioOYrF
JHC1SPAZlipA7aVw0oFty6/Ma6mHKrUyMhN3n+CkI9InfSwyOqRj6q5WgnKIaKSUyZAsCX4J7/a3
/U8XlGCJy++75adoaprFTkVtnePvrruw43nRni8bzzc7zreXh5rLsDYcgbv1bbmJ+5w0PHlj8xWC
1inlT4+yQ6ggO9HGDV5/+EK8xa6lMPBZYXy/C5kkKDK99fA7q0Wjhpaf59ap8J+SRd/SIdKrcISF
tg5VXywNNgGdHXTuC1zDFHIgfT5HOsnbwiD5+C8hkJTqlH6Yq54QlRpxwBTVLaKHIP2+fK1tIn9g
DsZFACsNcb7A985+eoVIhsFv+LD9qANiqrYA1JmheopIcPPDgqmweMcusaWPgNyYUb6sYNaozVnC
1qYUokIt9aTbkHbB755jmKg/W2L/HGMfh4DdUOC7/BUFe3ltmgP8r0pxhD3WrtFa8TQH++o3szIV
V5YU81WeV7WpfXUDwilBK0iYBwtzFIGTps8Hil7NpA0SZ4Ejob7MVNVZ6iKuxXsekELhwJ04KeD+
ENmfcasxVGWIwIw+zYRfqVR+34fKSBKqVK/eljB098f/xi/SmuJ0Vkd8VxHoB6U93i53o2X/YrIn
0iU9S7/fuV2i6qWuzRaymWXbTL2Zig8pW74ZCg7LhQ+C7DkWjyh8wr4+ENXPkeUxaF1USTQZMVUN
hRTwnvVkurl+PBrPuT3kgqm05CBzzqzzuymtu8qTNdAFpFVkcTEHC8g6ervGlTWjBevY0/ovlvfY
Y3VPOSRLP+mepbd1wqs1lS7rNvJuLrsSgXXSUlocBps1ad/y5ps0+/AcqIQ29BStKwKb6dCMF6WH
1YmQ992Or+cUyVSz9C9dJTtohs3hssDpl0jPW9rAmvw3pMqVZ/aqLd/qkR1KTs/OWnZlDUOzRitF
wtcpB6immbivj4om2f0CYPFcGE3sIFrOiW35uC1Suh3Q+NzZDP27NFwfqIcJImor8U/hqsyPxGkC
rjYu4pWlQr5FlSJaUfz7Gjn9dDva5noQS/SOlHjBkPhIudynMkUo1HBrAuWFBKqbrCIAyGBDDEQD
Mdw58aaBZ8bvJjngJIjoKO2W1oOgRUiXkCvqAiks3v4nvE0ZNcwsc5ImT37mkGvQyhtBSK5ez/Ot
uGWFSCy7afocgBrDlU2QL0prgmGc6bJw04TIlwxLNLtoeaw1TDe2GEvFkz1lMLwvUW7FdOBGkVJd
DYJZONi1+BcX/93AdxH0k8mXzS3jIWnKRSdisyL18oxptlbFTHOeeYvgtj7n0C3fzDhfQCrrN6I0
Hn3Ma0ZC8R8ZsEx5UxW2VWI49hnpdOhCfQzUfm7POd9KRfb1RdiYylXdFlW4+UIMAn932xKgIjzi
TDSj1wpan8l+YWsBkwXNbuEUgndot9o8ezfeS0J66NFDugS/3MgnXW5KMG8+9VbG+qaWw2C2cB31
dhRkO9Vy+4mTb8uNyDYy5ASRPCo9y74f/ovnbXc+TPIF+t56FEiSbxvE+EVhiGHkPgpbp2tKOapm
vEDJ/XWCARw67+E+Sc6Jwl/KhPtJ4PrrpA20jVAZNfMIuROOPfzwqLfGm9YHH35BQ8cmymIdNRZ3
Y0LwaoMKFsszdDzbLyV1++Kn7hw9EDJIJj57eDvU2ASoTZObBtStjIfGquBxAVp8HpbfgSsnIoMl
/l/LndSNdxNvHQzZeiN6RUCCljWpvnXRUKYH3ZwOQcLBhYJwIGA56LGTeq+trE+1phWxz+AnLiTz
MhM28qxgm7yiFzvBRis2xTE73DSug5SUyfX8H9STkwplpQID/pKo0mwzp+MXyz5CMljwrsZl2AoU
sXzKuQ0zZjPegg+kfD1qfp2GZeBc67OfiLEX7nJdpZHDAl6H0XIoWh2tLgcSipeU1bWT8luCAKpD
3IqE64c4aiW1VhkJ2HH8Tyx4W62rOTRxFnQHbe/vGm91/I0zrjdJBxu2kwznu857ZHjMz9PeK3Ld
3JD5gZQ8wgoJiEmt88ZT2A49xD1KNaJpwrQWxqh1YGc7mrehWavY5mGh4iSFLFZ6NioOzNl5f8g5
w1iKOodAh/IXdlpFOJ1j9N1QtBCisHaAFqCdpm008ewaTaNeS+RhH7ZHgV3oiQ8Royf+QP3I7quL
i1IWs5vBasU8z6F7QJkqqfAwR2dbUiuIP5/XxYF/rbr/ckGJoBMSqmAglVsJ8KFKK12EEow80zrl
fcweWlFVI2Lf6gJaoXJP8vd/dZ9TLAtsgF4dgB3WYqXJaFuA5DVvoWuytXq72EJvgGmx4PGLZ61W
S9wGSuUlYJLA4eiTxYy9GaFz5D30G+It58qN2yYVnWxAiPPgl9o35aifjFzlkAhOJGXy2my6LDft
pb6wFa8r4VnmZJPVVrcuS4vM54tyM09qbgbzPauE7lAb7j1zoFOLhjduM2gJdeWOhDFh6SPjO+NY
kMYCyYjVp4h++CJnglUXsPx/DY9N4eUoXnQWhd7KTwKdhvHrjJ9S4kdlm9Cp3zDFKJB1jk2Iug3t
lBQ7q9Z7aH6cweGK699ZcrVUC/9giefKCzPNMzmjENtjw9GmHxH8jVa/N1WISSA3NPIRoJDm27M3
Z3Z0Gd3RNdTTNRPccAXIUAJTrlXJT3CYgeL0OXhiZQzauxwmlsXhHepGXgfRCA4DXP76F5ufdS0q
MxnplqQb+bFvAIgVWHLRjQl8MeT6wchYjG0w4CtCC1hpkHBqxqeCTVFeP0Knlp4d0GGxcq+AA6xS
jezGZ4/sx+9bI3vbcBazHRJefEpwKL94pKLNuosv1xIUSxgOr6l8D3RzVGkyDCTESseAaFPOreeJ
xqIulkk/wacpPcUnOFNDc4SMbtoxKlymTrwVArqQJ9MXTWrDJ+p0vmy0mf4485gBtBVnmitE4xwi
r50UWu3nc0fb2dCr9gew4M1VVs0tpX92KmglCYoJCHcnR+r7tG7vumXKx/jVcCWoheJQbso6Xxkq
8FNa3WHnS+5y8LVpNbo6nVgzw57LZAFKdL9UCR5Pt/JIHE0Irkfs53WXPEXiHELhZltUh5U1qu7n
TnSDB4aAo3nPzaAgLl+69okDViEe2GRIdzg30z4+/LwIIiRqNcTVkEaKwZbvwbvMKPaH3lrgi/Zr
qRneF9Fi1vTIxqEggWj1E/eOduaH19ogYBpNmYLZgnGUrdGVvcmU9k4SdJXvH2Nq9ffiziqlND29
IBLoZXZJNZJic0M0N1s8I4/F0fGpzswXehS/vXe8MAeFy+r7c9yX7FkWfQ/RRAanDtRrQzjbW2FR
p4SrYn4WUil2cqTNy9A/EIBWZRmvXb1gcNV+k23HTqTRjmt56Id42cYSSN2UWtV524KegtVrfY5p
KvDGqq8zTZKjEbWKvnO0qtZeSkOLKmesoI4+KTFRb8x581Mwue0PWRjrA36hBxd5lQyJMCHD21Ze
dc5ucXd84VmCEjnPludKP12adEcTyVB0lOe3FyVB3/vM7NsU9jEuIBw0cfcaLDJiE5wprZbuZzhq
dHB74B+3cb6cP7rhoeOx6YBFTZ1FaJmOv6STEspUBX+Trg9UELsxxtaOh9uciBvBc/eM/i+wa0R4
J3rHZ0sepUkp2jBwd4BkMEOj531DeJ18Je21uEf2bfO7BajshM0Y+jN1ty1repWwhqo8nGOdVnxz
yKKhvkSwLfyMqCD310RF7/tiNIdoDrYFQA6zf+yBsVE5ICShezl5msOLG7FmMiO8WLNjR0XiztKK
RvZZ/FroKI2cNjp6jFuUFIerkTdR2ky7U69TEB0r5fkEY6n2JvdXlScl9q+Xysb1puR72oeDSk8C
KdkBHILPVUP2pHB4Ta/F+6W8075d//EBeT8aTBbj/wmlEmci/UOuvV4Ta8C2Bsbq1aADyxeQ0mS0
S9sl46kd1Fd7I89DMCVhgVn6HAbhESgJvtkFfS0eT4ntvq7F7gLnrvicRmpe66z0mmUk5WLziTCA
frmBlff4SIex7V2Ah2DAhszY9GV7ohlTA4vhMUKSq6UqamIi22Hnc6T2flauzIMgeTNmLtXs6S3M
MA/fUiLF0h3nT9/VZFXY78M02ybEe8PT0pobU83BJGS/nOKCGGs61o8ddBDO8WCr6OrxpPbJ1zGO
sR6zGqAbK9RDuZRm5COB2+1G6GX/HbRXXF9O95PQBpM+7UwLIbmSzSt6k0HFCLvNo1Lb4ZgvjgHz
oxU//Nh94ZF8+NWMAEm6P/aSmU+7QulTkC/vb5Cz/LJWnE+KAQ4XFqRi6gLJb56pcgv8fpEfhKnu
h8IGSAGRXHOv/YX487jUoGjVSWzE+0TI8mjgOgVIvXmCjvoFAjQojeAT6JpSIy5fKQzZGC5SsRnw
PsOZJKnXKjByHtodiGcS5tyGwK9xSkvJ18SJvjQjlWVNsicpMNm6tRRq1zNN/KiZWDZXUKnnBT9v
SpU0FFEc4SVA6oIBwuekAUVU7VTwl3MnlvuBt6p30kBBbHxI7IF+v9S5zcqyKTlXcvMXDOJ9mHWv
hUHtzxE4ytig8JwMfub/dYMORyu8pdieOHWhBiIMsFaQu/JwZynyKiBx4aaMQhFGmaeHdxwnNuOV
wVWMPgoqijW4N+dJzrMcwxQRZl2H9ngBR1FvkPL6iYbpjArox/8AG0EE43oJEUOYZAiZ8s5RMIs9
idJqJkJ7Wdfk0T4OBeBcNe9Rw64YORity+gTqrxTrwIxCN1AeZs+yt4KMjcAkBJto20G/vhlNdS7
8M3wMw96HFxrfutCUDejSHB6gGSWMCyXgJHe706TQAe7LSjWMXoGdD/eoFioL4+dfN7uJOZAzXJF
SC2gubhOqzDFSplTfbdVXzLQjAq12fAcIff1WvwhJ/w0id0Q1rvT7qgBvQX8WzD2ChhgSnehtG8p
1GVi5ciGbXzxpWAdAVRP/RDV1FPemtTIZdV+9fl2jnoq6gJzUG9p+OkVYeB3nOoZ/OYtlCjsbYA+
N3krsNJ1h86XMgU/LMFTdAiF1Z2EonvYEvC3K/7T7r5/tyrQeuFG2j3+2M9rXiMX5Yxzs3KF6qTj
doih+9AEEcRnI2LD2wg+S8/fBKSZMGX4qiSVFcaw+ETtNISaBnho+uYCavL+t2Mc7jsqSeNG5Knh
RyzDuqeV9QKhb6UlSFx7VfXqqqENtGQeIyKzaibqJ4MlEqEBSrDqa4rUneAI15l/ShN5Lb6cJKZq
uILhyzekYPsvUDGiL6FN3OQniD8nFLlrRQHnyPnAOH8A2zWwIkEzlj3ui7tc9AydJeEKsySG0IXN
HM1kE7uTtpXWowYQNV2sQIn/vG9RknJr5LMGjg5ek0rQ4jaKZDUuU8H+VpLLuxehoiMhTA24mdzl
9/txV/8+Yko6zfbOvNWeuwgZec8tiLAGeb+jSUH9bHMySFfdALOa6eK+s3Z1ytPjmFPwfGxfKckv
Ut/TUb4lKFVq56HRYrRsi9kGniEkGuVl5FAoh61Q8zZxE2qYC2oKylXO7iMatlIFMtGQykvzB1GL
QgW6p+XLeQAKvH64R/La1GztOR1Jv6nwK13QQuDCjsSS+aP7dm1U044LCSgAQNwK50ubrMyuh4cy
YcP46cBhV38g+eEQD2Akdifzkw9OKNWChCAkxKUL+tnee9PG571x8Ky9xp6SRxMKf+9FWt+NuCA/
1zVADT/KOeCgE1b9fy+d3YTX9K35e5Tz4yoOZ5jwyUseMw3KsTizmxV+j5JL3/p5AcUozerLl9Ez
uIIW5C/ZYVFuwiEx3Sya4v7ezHCl2W99Kj7PA84rJrgCfSbVIb+CMeo5KTgxZTbg4mseIWcaGIw5
uDn63puVmFiB9t/Wk5IeXZ9mJAXzPfxtRB/GrsOy9lxBqnIft0866ReMVRQJJEPToRsEC4dedukr
3r3SPgNIs0UTAUF1sLcRtl2mUfXRbhYkfCxtcsiZQSy0wgtV0HJcYetPSqou/0FFeBCEXPGoiP4K
MPCP6rubNYKTJJGrK6UsUu/39ZnZkwktucgZco7dp5GDsmCZi95iVkLwo+q4n4sr/PfqIMu/b+0x
lGCO+QVXsuFchmxGzI80KkGUlxmWmr+k++/0KkUIzosnJwMBZb5d2eMUHcX291jUTvcNV8ifttQ5
Cbd7DrV96AJfpsEHo5Y/AyxFSKEFjQ78Z1l0P+y/RvH4Vw71lvgqljb3ItNoTiwQCZ/2Z+VOefWk
p5BLWmvttW4Vb352hYXLVghL80HvdtUQCpCsVa+rvt6rDAxozcCLHgJgCnD//3dWAGhRsOL6aEyX
aITfsMApZdjqJ0/3KGzak+WZ0lZb8WbrDZwoO93MTaC/lAuSwDJgKXacVfD8nj/wEXu9TYkWIz0f
0QSk41dZ3soORfrIRCVb1wD2BafmGKKQ57I0tR8ZEGl3HwJnQ9kquX6lqusJwgHrkSe1miTLE8Xo
173PQiCMB69kZdk4g0dabK3haumjO1zverm92cSHQsaXh9cJBmTIk3rzL/iUs4min8DS011+yvpN
kxKdEd3LW3dWnszgVRgUOwFcVzZ0NyC1Ei97lYofKwuX8HOq1YUDdg/HkEaCGuj4yI3xJUu8bqQC
KOZnALZR8wQ6q/tLHoq/Nbf3jqI7ziY9VGpevIg92fOu6t7xu/oKS7+/WslTP67xpdmq+L9VwZOa
xNgSLEn2EcS669tZ/lDCW6auAWIUIiOlNmR66Hp08SP6iRiqLFg2qiKc0GvoOJRJYFvsYZPvvvG+
XXJYH8fU+puP0d3iOM+lfV1A6jbv+Hk31Gu8Q039uq/CgdPJN3KnJYnicidKj8MsA3GwMPJerkmy
G1sbURPzm2K8hMdN9OqsHaTQEYpvemo/6yNG0vQPl88SL9XBoZPO1MBQb5E5ODsJosXxJ0yxskdi
ESssee/uaVwqwGULM6lhNxLtNPKBLBaofSuUHc8d/ZZ2uCbTzSamKnJkXxTqpZ++JhK5DSm5VYIg
YHcv0Uu2wELBj0K0OwduD9AiQ2YGRGAczpwLKCGSVtjAAzzn6wzZAj40GNqoKwINK0QjFl65hN1t
K2KJOsnigbdlHc8PbhbM0djy/TWatz3bie9B1ydblORYqX4VeOsXl5XwdKgvuBEyuWmJol50gqig
n+XxxUwk/3ck1YjexnOtRJC0fMRWMmLeqplkEVfdKU6zwZgoyLB9vXapSV5wjV8erj9xdNQCbBGM
PC9v4VgjvqQe0de0Pzc35wJMyCoyeMHUb1Bg6ZeWZjY3w5uIk/70GQqxz6rpFSXarRGD39I+agaE
y3hvZDQAg4DsI5XFbwjAGMHi+YjkvOTg+QGofE9MvgAC7HMs7orvpF/QEGrEkLukJ43yh5971cm4
5o83l0wHzUrJ+Bm2WaiDc09JxIBhpUe93IegHJSlojgXKoPxtgs7q4yBTtr91R3G/FdDErDydMyl
h3BFbCXwOrG2GAXnfjs6RxlLTXa8XMyRalZDLlR4D75toLJpVYqZUigB2wLQekrORqaBSeq+rioy
PL1LwAW19jXzAkvFN5JRegb7WsgKgAOV6m5uzvWzOw06EOSvIqo75WCxft4bOfIt5H8djZjnfmvL
Yg9B/t9x9D0rQVaxWiDqMX8S6AWZLTqK4O9bMYcFSqkamNlIcOkf2SI56fHAOjVhlIXhA8PtSbmQ
2rooby4dw7KPC0ckuyBmWwgXeW3JHCzzfrNqsluY4VdzucEBv/vKy2HnCJL1+1HhFiYxLFQ20eLd
J0VSJq7S4rsx50Wkhho1TQIpSjUeCJTgLc76N+CR1bkB7nhZsZXIVpoy4FbSrepKk61MkDoc9Lp7
zPvXhvQorDrRbPqrLHNrZdLvLGU0JobpOkea5xNkHCaAvMPjwSc3WHFiz38Q47sL/v+jgSoV8fIC
vbqq5q+B6knR2swi47rJreLy1nROVHzLUgvtUunFzYM7HWR0zMLvQosCmgV8dJc3v+NpEwYnTe+x
kaVKZCehJQOloLB5vLgncJVVjcNigk6wrKKqEC7MtU73MLS0ns7KPMA+I0OspOhOVt3xeYKuabIs
QeojTsj0m0fU8dlQz8v6fjXHsClhwB1jUVwHS6z5V1C3wU2bhycVYiudNWD92rt4dc1CFYWwxe+W
XuIv+LKekvuQQh0ZzxiPBg5EqH0J5CxzMPo7TZIQjCK1d5WB7N22iPBXJU6ywObozBwyycte6NoU
CoeTEyGBc/g1tCWlCfVkMSgmDyGow9fmFX3eVF/KShVWY7VWiDHpZbOHQ4FwL3SL3gxj6bARo5/0
tGH6B4c5CJieN0TQEIW2HBhYj8POASoZER6pA2lAGgz1rfIvzcsIrZClEod6Bav3AvqcTadbD7P4
q0UpiBPJRwzKA8I925bHLcoT0zq6+PGWENsZL1vns8WPpWin9ajFbMv7bYqSLYeP3JiG5v/04jer
qt2209GdtOM6hAsRVa4N+hhNUgVaxcOlVxDh15BbS2KzKMv6Hfox/10khzCnb8sqk92ytFqtpzz0
ZWoy/uRBIrRJGhcCC2cF7Bmbrq9agtuqaOQpscf5/O/KS3fvyrZfAWRf2LXv3KHp622QfwX3Yo0f
gPAdThRtiE2V91a7qPBTvuvTISS9v4fFaV8yAtO7C2VcgoLlaWrQoXurl9CRZiYeottRgDmBtUml
hfUfEHtqxQ9l2B8YtR1af83YJNESxnnm21lCf4kMqwaCaoYgTOa+F3n3z+gFu9Gn34JHckM0LYCZ
OH6hNnCI9gj9C9V/0V4p7ABwb3XYfbV8GTT1jbs3fJeAx5oX4htZtaon0LXxHkcz+c23wOIBW9xT
zhM7fM2OosLI9LDB0lCTMrLhrSn8Yi8ORChihCIPLXfQ4z9OaCBUx893XANJQ0n2Cf6lSrsp8EZ7
JyziRX4/dYN+e+ZSnyFghFHenxCp01SzgW9WlLOhPFAgegkmon/eGACu6j703Osk/wQ7ujL8hCFg
nhEIm7y6ud1+G2/PE9MjYuMN3D/MtvxHnGhtXN3d8Whgf8EUWonzTRn3gfeX1Cce9E4RbNihu5uq
aCqJdidGQpTaAcY4tmkxGCv4Rq6zfloADbbLh9oWNHQrCYVZjndIB0BQqbgBDAHxHFs67E1PIXsu
Kokbczz4bLZN8BDFZDsstIZBlao64fk1PwXaWiq/YnmLXzQC24fGG5z+QFV/NHQHUCyuTttdjmWJ
4x21qo/ODSCfHADcaf+c93Dyr/cFO8RWE33f3n00yt1waqP03cuboemw005ybFAglyuwIyS2h9de
bEbaYuzraPDEZedHPyL+98wLpVF+MboQpg1id+Wsimsqdp3Pn0REDglHT6oQ8PzP5+p5Bqz5uptA
Ewl2RFDbA4U0ZaP4zSAwTWkX9A4H13soZDzgqLMY5qqwM2/yePDJ6fYACxWwuzH2XJA715ztKAzo
FRkdI2FlJVwEXFcGOvBPkncwqvHJUOxi10XRPDnjGH448n6Ak5zXaBKVqCWrwXssHvVvYgwIs2hS
3vg+e+yzmOi3v/VfGgbpJzEFFdS+TpKJ/ROvihHHEyD1ZP0RdwX6rlYoe3bb3UznR9v38775Bz4x
o4AyoV+L1y2kDlsMkLvDUylWwGx+9RxtA+SAV/JXy9+p/tUXUnPYq0vOVzwHwALKd/TKNFpq7j6W
bBwz74sVQMoQc4wfrHw5IMoe5Ah0xnOQPVAtdv9NnHaNj+wzEeCOJ8xs8dTIS4dstoTGUlkmuyif
jUy07r3jrHnX39lzPSBANw/PNBvpggarA1GnGISrcXEM/iBkg44JEWUep+MwNH7T1Y/zmz+g6QGY
Q3Mq5ELWAaPRFsumQUc9ntS88dpBDiXDQ3QVgSmGJB+LGrrcKvP/z0BoimhA93NnCTmFCKhSRXrE
glnmrU6/spnB25mAeYPHcotcQPQXPIWMEa/Kk/NN+aYhh+RnRFJKP7Jr/U443CQ4let6b3AMV1eN
u+5uZXfrl97ZiZz5GblGVGEY2/BB5tuSdQY05e0ai0nyxEiM7Z7bxPEUvzrvSAX7Umt97ptq02BD
8wVP5DDDlAXmXaUmbHC3h4OGHb/jGi0JhLi2oNNT9MSCKvZJBqJkgisTxHoapfk6voJtpU9sqkx5
TUuZkNvdqUrRUPymFqsHFjNr4wsn1CLEG8lghBAywLCtVsKong+yRNx3ZjW4ya4KkIgYJNVHhIpK
YzyRMLb2wrXQekBXKYCCq+6YiOuRkF7XEW6jJK8WJCOvJdbcPltwzoUFF/ZBbQJrEaxDGH9WEVaE
vd1x7l4KOot9Tj1EaBATVHXXR4KPy1YXcICwY5wXlQd+yDuBCRa+/jwd8tcMxvgOl9HwpMmhjOFA
7ErkRv0rrcETERE5TEFakNAErIb5JkXMmPn3rn2Qcuk55ZUtZWd7SF2E1x5wNI19mMKmoJ3L+N8b
HOCIfU+s9LOkRzPhL2a0v76Ut/BsuOYS7n1oM+7nSh15ZhLDGBI1j0zhRZ84QKMEO9dLSVAX2EPO
gq4ewgzzFkgWhAB+qvyzzZ8UbpMzBDU0o4oX/+iUVB7ON/fPQo2+luuJe08+1/5xaSq9aaSK8s9B
veoNsjE05mJV0YSmukDNRaQKf+3DAkIgtM6CqfHVTh8YF1Lb3ACB5TcKGaZ2dPqpwJl8hkrk2xIL
yonwe4+OaafFaUFoX3saN8auXz14PXGM2ldTjSUgp1WMKnvrdS2i0eFjOO0J30v1Hh5pcsSV3HpX
kFgu/LDaOEmD3Hy4vpqEV6K9fWazE5A5DfMiy60ttK9FuWDDDU76EJ/qy+Ax70IsgizwkorYZuWB
O9lynKnm5r69D4kEfXJM9fuJPI+zy+WgZAqtM5Y2kDiYE0+6LPbudBrtwDYoT6Habv93vRBkR6dB
TjwtvfDpTxxVQ8o6UKrG72xmRqUSbwCk3pn/WQs9r6q4kr1TTLXAXimdUI7pxxuZzKyr/y8Fwlmt
7R6BkDpcfOr30QAbTRBp1F7Cs4+nLqoimRdznhAHm8hGX+YGdqifobM/BI2IRmuD9TqXzbQqYpVR
AuyEVELNZQY1l/NyLuuYpsCWJ/xE8qe8zudTev2mV0nxvBmK2jmn0itMSeANYMf6H1JlsD0DfdUh
lkk0LykGWlrslB+m2K1cdZ6noR72R4QDaz31nPHWFV8X17fMAf0fTU/NTW2KaH35J31m2ahobUe9
p4gwlRLi6oU8Xk8+S0tDurG9gve0Aaxlj0xMn/IFNnjWj4UIKUNNWnMq2YzdiAyhHfnf0jjsLfVF
SB7J0CJdl0S9rmpTSIQK8qITAz1dlNpv1yBsV/VjalMg+5P/RgUM95w6jUhcPX3dml9ahjA03akU
+V/3Hr798I/ZtSBAJOwhln7vuZf/G7RneYxT4N1fV68mvafxytHU1DwBVx50SboTaGBgQ3K2bE3o
CosZgcF8Pmp9FSgBeo0zP4dpaUbNrsOfWJ7Lb9KzWB0Pc2Qq53swsUQkjx6QWWthwawLwcbS92Dt
9VJx+xPIUOWjOTNzdNP3l/52V3RNzHocSnXEcYZWzwf48dSdvl1p0JPbu7xJGpP1NzuBdSAuOyuN
UPavS2sYFVgWxKiXAF32JOPbRFptBnkjuwP9kfSsyq9tocXBQFbLwlP3QkdRsSRU08iWCT3Hsfj9
tRVmQ55x7YC5ptYov0aJdGT+YacvzWca5mqLkUls1pBAZkbdeg6kCjHxVwGpXHV+1BF8wrfjke43
Dyjb2E+5TPOMpv1cMLKwKqX78kYxUcXJ+pJEMSx+7x8PxY7ywfSpqymRdWxnNfVmB9JJ1N4hwjfm
xBwdavCFK8PgioXpnVJv1SqV7xIBGrt/mTXMvwHHU90SwKQ12f5u8Hfm3P4wGydEQO8bZ+c04lJY
iOib9fGZFrGhK2QD7rX2jRbHr1+XA9Nt52QYhZ4pNN5dEF9/WAVIA612x2+uw8U3Qb0lOqgVRIid
SRsAETd+5RUdbPGC7qo3FsdPjm2W3DeJdScjmoO0EHYVSjN82YvMWecfXULh3sN4ZZZhDOVq8cNw
15FPsW3r8gJe60mrHu3fEDw2ywUH+p86de/Tvh91c6CXWRCloQOp6lid20yh+r6najtJgQfIMlGe
tM6ZjWfztbPsY0DtC1JuIiKMPCRghwcpgPUlAiJngooZLy2O1Zr6qhByvsnf4+Xrj3gMvrA3oCJx
jWjdMc7Ru8mVPEDOS0Xgo9cWdWJwZceKN7n9fdqkKXlaEmj1HdFJ86PmFdw7kTNV370T/7fTOOdx
stQ3r9ZgPY9K2ab1msi80+qAgWZoSo39lei1nBec0sM8HhxkddA1zssJXgGNEGnbv7iZJ2qcz8EV
yDCEm5dHXVlF9xU0VK3kiyCYFQzZjAmY5IqZ3iMUvwpfjkIl9gLQb4SF34ZtEYi207CB6r6UuZmg
QNOgnzLM3MUN/6dEThukE3y/d2h9qUPAN5Xa2b/hI6Icu5piL+G4O7qSrGPaSJvhAu4qXpIJldmx
slWvaaOllwb7LtEkrFIfceK4V7BJFVHElUGQGGPIQ6W7ZKcHuonlD3SqYMfCfGk+8MLW6huB2xDH
ABPQNMSIQKWYiKc7omNJ2BHHiZ10JoKzdXA5MDipS7cudM9q6O/rqvrKCciYwBSJH/pTw7fbbEMB
E8PynQMdVc39ebX6WFldc+dkR3EdGXAnb3dVdRPgrH23aQZTCnrscssR0iFFm19LrhkyOOjid+3N
SJ1iitiVGteo+mDuL5TtYiZ+VEYTx6H8ZIxABucEP63Pq3htjhVoadmx+6EBUly8/3TimugYzt0k
cWu0dinIzPrR0CuRAPLiYiNIQTA17piiWZq7fjl+a3qa8KIUSzmcq29a2ghHGx4vLoxs62HJEL09
IEBqMkMkqW0QSRNC80d1m0sxAVP6P173la9vo/c5OPR5lJ0qXMm640fNhZ9HdFOw+3nIZRz7+Jir
QsKn3dXOZNBHzh5hA26gJhAM6Q3JSbMwii86GkAzIdCkv810L8Z44x7hOYKjocL2kk0hNyBmpxCq
8+UTPIJID15YewqCHJPErmEuhdtLhB4Mhm+tn3g26vTfFXHPqt3Vjpm62IyqIwL/PaKbTuzm0djN
ut+uwV4D4fT0qgZ4gDbafhCgaEgF2oYaVe4LVpsvF99lzvBOPE1x8dcpOQUJaQgIZ2h28jcrGNRL
CNtmxtmgKFQMRIEA5j3SyrAz+65Ge1+U5+tqvuqOb5Fb6NUVDAvKSqliZN7SafOZf1WRCvV3BVFu
OYlRBhZBx0pLnYVTc9ZF3PSFiSya68p/8O0zIc+naVEvg7voVY5wkoFce8uRFU4agwkt247KArci
n1XMBQpouJnNiUuVAVgRanEPFdEJ0m9VI1DYVyv/6BsmvWAGWqsfE4DUZQAtpsYLh7l07SQARTQ1
s87i+zayNR25DNR0dxvnShLgygi0RrfjMPzbQAmES52T/m9d0IKS//2W62BPr09EHB4van2T2mZL
nYWrAJyNZP17/eiZez7JxFpB3gGrOoQag6iS4XLnMwM4JH99tws596UAi150nHJKZLreCtQ7sJPR
fSSHziH+et04VGfLxJx8eeGq5Ju395ktN0EA95f2ttSEsIJR3Iz3LDiMFarB0l4EmXwVY05Ydc1m
4BOnZJe39DoxRi0gPPwOgydWwG9Sskrm0SkzMV4+7PYHofr9SpRwRwl8ePfXqi7HFU65ExJtuHNt
QNJ+5GrGh6If+zxFmxNgZId8j106ZOl/uLvXUG0HnOswKKXISp5xFgxyVe/XOauU5eyjo2QKRQ/d
Wq8iyp7bwEnPM0vWpZ/jg/Jm4snwfOu9wPv8CnwK9SsIom6AHmBZ+sBjNdKqlDwHAwAFq1z1NXSc
ggsm0FgB7jDiYCh7xZJeUrxJf6HU8AbcMtVb5mqgQfScltgn5NuI80V5iCOV6G7T0KkB3kEFogW4
wknLjGbBFK3/G8nJSKNouOJ3d4k6+h/vpK/mt6glwIm5/BC+zF7olTBTeF/b8R6YV21Lt3nh05j9
wDW1IAr/ChSqQoQl6tHjyCmZa85bZp5bL9Z1+i+JzI4D9THBrBUU9o+Jz+h3xuMXtcpuomDBAuY+
E/RROCmpUJTVLXdg9r5bkqDHzsFToBDYzllLVGBSev8rS3CpRnUJ+RsOo7uQWujDGXddi63Qhnsn
PbsrB1dN2VD+4JYhE/IjO9RUPwMq+slmkH+rdz+sl5HLuGq1MRW4b+2cwmFi6mduIX/wiS30mFxd
QIWGs1GhTSbbFhNJ4PdsVXHT7eSrxXFZAvvp7DxlKqteuvfON6q6HzNNZIlVoCz2lfu5Hr81OdKd
cCdzJh7aAhZxoFG9tchBmvGK0wKgkNbispCSx1ZP5qANts6jpHOyDs5WVLgwaAIOM8lrJIOz4BIA
cXhg86kBC1vNEWWDRg1FxDgATIjpcY8KcuvSoW4YlCuG8RTG9q9WluJjH2j1c0F88UEydbeY7f9L
PDrrwY2pErr3eVLHHSiKBcBApUlEl/kaHMr8FN8pLsVgnYwiMh5s6xFlpKua1ttsaD2OEWmKuzGz
xin33ymEpW6U94FxQUvmYZalPZZunCc5GOY+0p+Waj6HFZl1xVh1FFyeswJqqdmxVBfyrA+TSvdl
w+H7iwvoDY0nv9j21/UzKJj/e+Q+eKU7RN6nyZGjCehoZPj+oUj184cwBirwiYARejrUN6BVQwdx
SYGXC473+rCF2LKHJpSY1YG5f7w0Wsx8raHbzx1Nwtogbh8nFndNJ13eWaTL8es3OvRnHkiBOCgs
YDhJLs6krd4oF7XZJoQxdAx10xGSWa9HBvM0NnrwjNpkeOmpf4qgpy1kGNCnQFGYZd9YOjT4OEyz
0GK8aLdOdpxfF3a4ebN2lkhEf8gdEarIch2NKMaNRakmPYjX50M4g9Jf/vbNO/E1PFYwrO9hcg13
v+lDSJ/jeFx2N51wq7n1grc1oKQhuKnMO7ZVuH3oG1QqJRCrNoyen8ZujbwiBFu+CQzu4b7V7K0C
YAkYBedaeB9BMLR3ikWmxE+YKF41uMJQdXx0OmN4uX+B2FcerUqfZfVKC18h69PcSn9mWevmZe2o
2unKD/gLo2eU1NNvbqKpL62ZHkZkIjL4Mu9iTUq2TAES2+tG+LTe150uMRveAorRUpI7h6mwFR9W
D/zWy7+Ms7B/pYLdNAltEccM4syn8UVjPLWPRxXNRDkjgG6vtbJDVU60yHy78kulv8GZGwcLdL2S
5rVCy9jWbU532Lhrz0QslbDjZwSulDZViRIt/Xb7nRay5gy6l9ihh875Q7fs+ykBxY7ffH+zE7As
Y1635do0KO30J9si3oL3su+tKbGjVsdIHiuDHQQcL2HQ/tZ1wUdFRuLPvtUaD05aF/gGcpZVjK1j
GXCE2vxJkHI31J4HcPg5EcgZJazz+VNxORpERZrJwxpWYTV0CoZaj2nRw5zLr/o3nMIzxojeL8Ce
FrhMWVV8uuVRvFuUaaU8jc1TVQcB+3W99nSM8EKEUfttHuFpSmyyLcbuFQWihEshHCwbe50zylod
YY1CwMsoNdymtre1Tw81juMnmRqzOGprbAEFsOYP9G52B+HOJLKlHr1pbY9TTwpS4MQz4aj1xeUP
ck8Np4dQ0CLtp5tJsz84lgIRtcb4KK3d88gGKkwSolpR3MwE2aBx3WS+70ylSXeHiS41LQZnU3F+
0ydxMcqsFtR+LSklFyCCn/6gaY2ms1s3th0EY0Ra9iL7Ue+COLzLzIBOhq3k063jSzxZDEpuRiEF
cgivJ5ArCUfwHv9GyA3eqi0ib2HLtkpM70a28xTeL1G/yWrQIWPNvx3frGpvrzuQyOaWbfYdLTVC
hhZyPRzHAgnroAy1C7Wr6JQDofRz9e/CmEt7PnaXiW6iHaWteBJqQTNkJlcIYusYxfLlxkyPzLM4
qtogeYyTFKiOpXinIvHas2aJ9+J1iBPNs0Gg0wjes84U+b0LSLdvakLlvW1JhsrA414PchcRJMHK
z9JrjSkbmx9Ugktb8tea+SOrTOHZVX1YzGTKXrse5ultfyl6e6PaIpASdxsJIVPXOtX8njWlusLM
0NYlZgjnHDRpbXXNMGiNZk/I9/FzOLuB6FwSlzn32j3W6Toqgh/JSIkrJbg2ivWcj7R0zVA2mf6M
ks5xmBMZrvE2BwXTPxLfzVoRH30UaFv3Alhz6utMzzcklNP1oufDxpIuxaCblFr1+wkxn9Etd/my
xYbVdq8mxJMm5cHEjjyDTXa2LR52tgG8CE6tDad52ryBdfUhOhBqL0U3x5qThu9Zmzp0CzWKF5++
5MS6MBPAGIZoiU/WEa6Gl1VFjZJsX2bTd2x7PZZy4o4JIC3pIZF1NTllIANN2KlCNxIy/bxKE3ld
u7tNcTbtAhV79oCEQWzlD7BiTcRLRFSz443rjFJ+ZlsNTNxFHidqHl2HQITq7HfQfj9nkgZ2ZPnw
yRjs8IqnUiVELc7nf2lVDoNfSuHF3OPzBwmm+C1XoP539hS5taDNfptflu5Z+tCqePn6KgC3yzmG
mJDMW24MbCp/7tVZVCsZGNvpSeVHfxbtrQCGNqF7LC7znUWqcLgWJl8WViwVSD+KiyGxrgqpxZiB
hm2DDrIFL0DPJWr74kQMFpbl7aX2ACOLFsykuB2IpJZTiuw/X6UKf/Kf77nvlnNt8/narn3djZ5j
QMSXUF7LPzhwmpwXeWiksHr6IBLnPBi7Q5TvH/FD3Bu4kdV9ZP/PNfIAA05l6+ocKuBzN2ES8nBT
IhyfRqTf+LvBrD8THBYi9laQzhWlUGs0HQtCqfrGQBQ08c/wEtsSgCXGt1BpoUBGQ19cy/HNdsle
41NTQycW8Es1mnR7d3/1AjeKOwE4Ef9PwIFU1ag2cgAJbAn/yvPN/xzHrqpw04YUYS8Mc8sNLMPI
ec/obMlMczBLMTe+kD6LqBiR589PrTX76NweYEtj7oXO+wtgae2xxRMJcCO5fXJUdRVANv9NkWgr
i0refR7TmsphnImimevVvbIoABli3X7AjC6VwQI26mgwAZ0pIGIP2TPEThuOdYUK/qSnGyWpGNzM
XNFSOg7OfJp+F9CW547HQx7vEiRq+oT4w/vT9sORb47MV2QcMvHCKLboVDK+1akqQb0LSvldfY1c
4OJ0xuC/g4oq9au/jjXB/B9RDud40RpLLdci3uv+dhGw+CBh+sxQ2PXdQd7hSQXjL4HBaDs97CAx
sHHT9K9OiQUnbyxSNiG8o6db05bnzC7C/TQsYkEEtewN4Xvhs/23h8n6VEBbMzHUWmAj1AaKgqxS
NNa/dxEPd6HhY3GUWh+8DmA5cKjHgKq4iAlNzJjZSIkK9THQHKNLffrIhkyrW8H1E7TLazUpV7mv
ZQKxZNBPbPLphsPDGP8JXs7F+5xwiOgBcD7EzaKtCjL0e5HXMqgjxbksFTzICWKAAwixLRVw+dxj
9uqufk5HNtjYdD6FxtJ6t3/DRgGtQWwF4W9mlJOYezj43DJeung4oz8c7FW3f0rI0Psv5iJDKijs
ZdvqvVan8cerHmr5IHKpfKzcVEo5wFgaHVynGNLSz1+S4ElsyBAKiTYZqagbSt2SX+uFPvNOvUQE
kGNsmwq87NxCRYCc1vp1t50PnhdAJiVqi+pXJ1vDaUqZybb49GVp7lF6fHi/CGD6aPCv3dCciq/+
c2tVgOVGiytxJ6aKqnDxpcw1aTZf+Ysr3ulnmNaaT7aQ0BJXosI23uGncmMlvt4mkVHnVtBpYjkZ
xzQCjYl1bBpwbGZPhbQqYJaNcM4DoQSrNQmIh6XUb1GawdngybwdtWFOi41t3sHr6vM+VaDukDKU
SKljX+qRBc4v/YFCHaYl4/sI4Ip768tJzTmNGVmURVze9nvZ4QIYLanJxORJV5dL+f2Ol1b4bE5o
OR2+b3sbaSK1jqpjTRRWJYDfjfzmtovLKDCB6zxzrlWMm1ebRxd31/UaHSE7QrXKPS+jwrOa0aO4
61ohsicdnvK/jNwuhe38cPDxRhxAH/q1hcJUleo8cxcLjaINqfJSq2xPWV0zHb82asL2dQsb5hxG
x8yNXpGv+t6cd7P8E+BVmKXbuWtDXWQL3eiUZvw2cgo2SSvkxXtYGZE9oAqMG4BSXNBIqjzUgddg
1H2i/PppJc8VgUUoPgmrVB4oSkh3hCHuHu9d6mHONOt87HnKn7ZKiUyfTMuUm4CppJeBSJSHMCPd
M9LVVH/Bjmavp9vlyrYVaV+2+3C22aPikyclsNSUN5NiQKn722IL+vkesC+Mo6yMu0wtF/6o++gr
vYE1JTCma6rI3Q837bv3zqQTRdLy18rxwz1rV53pS9sjdUMH7r/6zmWGIeLQ3Bnr7JVe70nXAAVl
7/UhhxHB4/MvHh7plzDjF/SkCifMlTP7nDhjxMN5+LX8EZB3WgkxiE9i+8Izo7kEBmiJeqrOn5mi
GwJg7e/Jf17FWsHDz612B9yYOpYo3ROE4QFSZQ/2A/1Ud4uXD6BmSwBe5aKl8QcITnFPginZamoJ
gOv7qPIqHSDITeFnMGTZ8alE7D1yw4Q8KbTUtwJtsaStBbUiUup2TfNfc5FlHmXn6L44qhYBDNgj
4EN+ZLQJZ57ClwkFY5SWpyT6UnRDgTxzl1ShdNz+NOTRUVTMzUeTa+AP1hGvaxBP32UK1xCyrXrG
5amehfun1sgJiNhmaOi6Al3PLGZfqmrDzjKtnKz2Qr09K50hXG7VZr5tlycF3WeIniBZS7hrFlO7
jc8EaYeJZrBcnnslGKX+ojWkzE+dXfTMONh0pjTEdYpObwIgDrvrOccYaw/1MU9PYqHxftD7ZzL/
TqGcEyaiFbuHK9Pbc3kQnO5vV7Fa4ljdvtOBWS5VV/e2Ezcshv5+HgUkfyAvqcfKlWOlkhuw3Dqm
XDLvTXp0lA8S/qMDO7v+YkwmyCe7gnghafqMOqy5wvFopgyaf3TlVx5DO7rmICD95e/zxxXq2bld
mQ5sZ65PLsfjaB4IyJW6lk/BSWBXLTh4GSioYnchg83UKqozUMvn6TEE8ml5kVTF6MmSvnJzOW+g
6eIK0pYudDUd+/uh/P/VGRmsuIuCVXQhWTVp2z9/lzytDiqiotkD40/daT38ShS1Yayrx9AaMlmU
MoQS2q6HJpdoM59h0uTgzkU4fldWtIr0KSdq/2wtsi9dE6VoIBM4KNLDNHzwqEYKK/Zees9DzQUa
OeVtdBXr8tYb0X7uQMoGLq9rWUzTsZUWbt7Mu8lMWQFTL+be3LKg137RlEe3+W0DR/6iKrmjlD7e
n7nztAzw5pKWVdOXQcCWDZI/777oCzHEr1N2HB/ny0sTMpY1StKvIgt0ioZ6BK9iDuljo6NfxNaX
dwqqdehCnb3S8VhAwgozs/g8vlrLHECaho3X1Qqvqpbdsl14SUVRuhlzUZTM80oqk+3FuvO4jmvc
7AQN4EfLAbOcOKYa+OsNEIUrp52NIHmRHn5HeIH3oavbucL53/7xK8TM/lQ8DHwUZw7EjXooE2iF
5ievUV/kWfbPqbUyaHHKXmlZy6gFzcS7SJAkSRMDJnHRlqSjt4mDugVzYC6YqMGcmfudxcrU+JTe
IdJ0S3knFBiblkDW68ylfFNVKxv7OLsBXItG8TOBj8/+FQ8Ptxw/KiPJ9Bcc2j9Glf16CiBE2etx
5hkh4zwO4BZvg3m2/Vvi+D2B8XVpkHPA7lQJRr8z0DxoRVto2oDz/vmfvkl2769xo0d4zgXrGTn+
N7hRfUFNcG/xejYwy5xHh7/zZYKz8PfhrDnO9RErgCXNNNVCFPY7a/gjYpyb8WbGN7wZJqAlHc8L
qHsuhXYOsvJhXotmNicsslKkK54Airjf1nYkGrgR4De7D3xnDbP65CmSd1rmTcifSG7vK5uJF2UZ
orY5cxMNqOsAX0z5ZKBP6yWNiM7HPXdP/A9DfOo7WGSbOD/OcFpz+sqq3P1wsHxfkBn6q0z6+CVI
OOjoURGRiSGF7hZ3B0MOmZYiHztykYsvyR/y4r8OISftJXU6DsCpS3y60rJSyqCCrTi4bSXjPBYt
SZUN1Zx82aUV8//EKEjGmV48ioI7gt/mVUSxX9fsFLwRfJEBLQwALxaW+Gbe6V6dUsvMDn6juFDY
IsbnnugXy5C9a+QomryCieQwwZPCeAgiDwRqDLe0cSpc7RnEJ5gs0LGVo8eikXfSYegCNhl6BXs1
tU+j8XNSrN8E1mUjENaJMfhAN0nEKKr8hXiUatB7MRRibd73Zr0XZkxTR5i4BjPRJn7BpxzjpR1A
rssKK//TX8wG/n2e53bn3bwKuiT6xArt6BjkI1PB/xH1KuljME3nPJWZM3Hwt6Kq+hyhm3gsQvVc
uG5gps/DOAK5ZH0Q4aeCQLMFujQp7m9qYA0X+kUQh+r6e8GPJmQgheEA+Fr2Qs5cZCjFaYrQTqRu
eEcQadOam1ZY/6CYgWcgKuiUzwsUJeaIMTWgDG/PIFYUz3nnDSOB/UCjLG/vR8ex48QdFX1BZ2L2
+vYpQY8k5KVI9AVT43pgk7w2ZJdFi08LA59KpSQYnpzzxHRojc4m8UJNjqBAk31ymdnnXd5oE9fw
APJ+iYpq1Mn8oNOVxmHgYerfbvLIANUa6aXN2VN6Nqbp7ygBcdl67lfuzuuthESplGRmYHUZk4RH
Ia9clz1rmQB5X3RGlsQKex/1F0NzJY1x6IHFcW65MDRSQ5REeSIaCxjotUL5ABwAcKzp527vQ0yk
TW2yb83AdSK01KQeQ7Od2yncvz6HtHry0gNo3xprF9rg6j5eWaJi/ddlIa9764s4H7bXTtpauHE7
JS9ei66h/7mepOkVcm3OI271mCbd2OJusKIIDwvTckKDwdKP0fANAWtgcr9O9by1oVAqewcKeWji
DMcdx9itOPq4niu4208k8WuSHiWHkUVBW9Byepxr0r10gMawYmaa5fYLA/1P5HvFWO3qhsLwuYaD
w2+w9YbZHC3KSMibwOoFAmh5UmZQZCBX7umqJ9oynIXpFudTnpkJEOwsVkAmp7iPH73ZYKLob/Hq
FwzPl68uNXRedcZkrBo09tskShSkWtJTz/agQfzvwP+q6FJOGROwYbou9vkGed9sWcIlvub1I6ff
5ne5jkLBYRZSlCIbpk1QbnyxbjsWxTSTzYwcIZuv+oIjK1f1VtufZ/WHafmR9Dxah0TsHrbwk09J
wLkjZxRrdl1mRBl0YkK58DlIIC7rJ0Rb3o5/tTzrMiqzuFC+ffXcmT5goywZUC56zy+a2rVK6u1u
1AbjQOf1eozXjt36LV+rQfEqt8CX5MOikh17xR3C5P+6B0aqS5aab8vCy7Q6JrRKxMyXkTCTGeQ8
z2MiFxH4XjuTyusX8FZoyq8qCEg2D3lL8JKtvbEV++uNM4TNIWw3ENP2ZZevI5NYccGRGNwmbcc5
H3j9rIVRMl+/B9w+dd152jen+3JRs9ekXdnEq1QtnXj9Z1pdR9uRMW2QNWz7BobrsTV+13VLxBDu
oO+m2pApzci1nwYr1oZ4AYdh/N/DMEMkstHMeKJBr93Qh6XteXZ7MyEBaTO4iv1OG0gaYeuWZL81
2M1F/RbbGGvy48m2v4Gh2mGCbt6sz+ttlflAVfLE28jScOLolnAkLQ3C+mBwopWZh+3i95+AMRdC
8+K9iTTg1XqSeejDwwGw+Eyx4MGU3INh9XCXL7fU9rXUeKdAG50odFfnL8e5z8BGL2UlttKaVUEp
2LGICWkR2wfG5aplHTW4jseEDLMFHuMWtwRpgubXkh3wZ/ZnZc8S2pnWvslpnbg0fy3qcDYAtckj
MmWs56lmSyJp8wK74zgKZNFrYX8NuQiNm2o/Mf+D9yN8Pdv1Lg0FBZq5de8Cn+mgn+vFd1sUBA4k
zqpY5lU5TtGlcrg5z7t1U9A0I1PLSTwFib8CPKy3Bcqo9634Dg1+eWU3k4xRPB74wBYVZwR271PN
lLR6+lqDDt7lF+ES4H7eGQlDTWncqrcW/YSi7Kf5187sOKgfi/QRKJVxDk6zNkBrDmzvENi7kD7x
w55DpS/oid25a6tyk6KDDtcypZUyYSwJpOgswcGI1rlRZTviTgt3QsOn7iZ0OXvxiP4hyjus0XiS
QlRFJBBtc9rp9vv5Mp2QoriR1E8CEh9JHuHmy0+1W3ZTGSwiElYhJY1dhLXrP+PWrBDm8HdXuQcd
VDYPX9suetQ0G6EKccYbj0w4ONrUHiNO73EDyV+2xWoTHzEMfittsL2tX+q6PjGbxkFjnlsW5bi2
pemkSF5B/3q5oUcbAA6G6TLzxQEkrfo/GAfG7n/hgMAVe9bPGD9VMf6ptLM9T0SfW1edKMV0hXYk
rtayw9/0zT7PWIgHS6sirWopx8taIkvoKEkwKV1p3B8sO/9cztUEorIiSmXm6QMTpk7cUWxwaJ5d
+c2nraWP+sWtLxpAWR3ykBbHXiakXp+lsaPYtZkg6nKl2FFpjjLXdu6xoIGQpNDNLEldVEOcLvjB
dS4V2hD19B+ve+GYkSIdDgFURZEqoWMMi1HXva8FIhsrtS1ZR3vOBhvM/rb7XxiyGrcmxELOKMZM
2bTIPPKB4I5sxOcPXOIWxL5xXUekyzYkmRX+XhwQtaF8ikL7Ozhx+iGxjVOLVP2udyaTOSjFkRzW
dhtRZdUyOQ2E5al97z0n8INjKDus4vGbNZOc0omoIGTI6QyM3X0va8DKcikhRJFuaVOWve+dv2A3
Gqu2bgy0gRifYSXx0n7Agspb8LYmSZL8pWIHDIVr5Hnrjqm3SKNt1MlfeMHs7RX/X+EDguqX3y2Q
J2nr3UuCNvkRvU4PRW7GsB7afQDZYXpt+kfBLD9MHzGRtg5QGfNG4OcrqdTBqKzPjf/xCxQfHID8
LoajEIsYZLzbP6iDHZnFO+5iLkze6/JW22unBX44BXRcCiGmUArHPf1vFlzOOcXEhHq81Tnz8M6X
RYeF2bV6Dn+AScBqgsh4NOXiSaXL7yxmNR4/23jJqISGHGY+zxJH3vpGmx0p8qdXomY0lt0wPlW6
1X/VTa7n4oeP01avfeFxclpoMc0gsz4pe34mIic5nkXfzgkOGxe+yp0gKkohx6QdrMxQceCobIOn
m3xKi68enDjWkUCypDDMOyuiq1lUrH1oiNeUHW1cTgE0rJhVKFvl+zC2IryqYjCqaLDXHlXS4JOu
4XhIKDm1LhyvWrHrGLwT6iknrHc54PqQC2ZimYsq+ytb0lSaK4k/PjpHEH1WWEEHKmHZQ8AkDgPx
monba3OxJ8U91Pf6l96nhcGCwRnieMhuRE4SGFgzB8XPY52Dh4TJXk4EeZBzlJ1njY2yUzvG0vHD
N3rzsTj3jeAlYU1fQzdKo1QwUtn1G//pP9AQ1MoSs+tT9mCLrsFp5kyOR3aBUaFBbFdkvjoXbFcS
XMxR6+OT3hiTOv2SgUpnfToeiKjaovVX1bITnxI2HDSYDpKfyoq0Kn8hP09RhoPUtNjiWXKiXfm6
JCVcb7gVwAMbjjn6W5Kd7Zjq/bpHCX0EJB7aWTejuD8F9c1DEMKDVUdjytAmKhCt4F1NDEMwAsAh
aqc7Gf7qUDC0EjbqR9C+kJvX1tJJUURzqc9yfthD7c76SM1kfNA/Vr7GtKkLCi7z7ayq52KBJa/e
WgXWWKpaQpl+4qE1XvemSvF6jS40rvenidjSZyEzvyePTVVtKVzdupWL10hEFr7oTANRc5RRqfj0
lUJWSwdwzDtwI/0NHUtbYdDhvcGLsyzwQqCMg2Q/cR70WlaICfm25pWh+SqQsChUWBLX77POZJKu
5oLzPAtnpBVpPFnXXfweZ/TA0s9hzcdLfsa5J82++kFQOcAYGgkvPu3RNq6ykHf2Pyx8IAXsk6UQ
+t+U42z1nsFvPuZD4GsEiPo3WsJIHN2IA+LXnWw47YglduTIOc9kLg2l7jR01NsvxzPsNBazgGak
hKs2wIUfkPcq6GrRA9FAC24XjHrK4pocNQ04MhyxTRj6j1N8Z2tUVhB2dThFbWUSLwn7txoFmIab
e8R7XsmLh5osKVyvjS/Ch4wluO0rzY5MpBX0qH7jB/Cn77hUUiABBLqoZZ0I0O6hk86iq9giBlX5
vbkTk3rwK+RfLyLp7Gp//y8izXCBuxY6wj+yx75k2PBCpPxqQDqKr/bWWIPz6pfCCNdGR6rB5aWh
iJ44t3bz642v4Z7S3sfO6Svd+EPL8fUlP5P+K/YTxRwY2ePHgW8KEvkPcDjcr/hFy+MR2QSML/cY
we3vt+c6ClppvVOLFovpVsDueWmDTAGsGiPqn2VwDqZS0Ik4ANXR899RH8f3F33Ohr5Dh4ePPa2+
9WbIkup20Jow+O91YPrJ4QePoV/u2EOAzEkKNmar9vx+1Po40j77OUc3lfyVBq7FZaWECTApmsXy
HwgaWG+CMbMT4gGqGYXdCw1748GesIqGpHASVXHgaX2NmiD/WbyWkTBVj0r6jb9DgxfoQ8/aksQr
fMXqyXfACGYnXl2hQY+zltEB4gEvE6rWCr1F7OrQVcQ5P7vjMn/aNPzZrlyj1E/oBLZsPRqiJRLp
1V/rEBrahO7LVIjHIWefGonmaeMBsLd/wFzXexeVC13zP4Uq5dX863rzXW8gdBwzVMvIfo2F79xd
1OnFQRpGAIg1Yeq1r2El16/B9IUHJqcEvQf44uzLHsTWUFwl1ecXRWt4jX5yFg8kRJOTu1WfkJms
ECYwgBvylTk1VNh/g8JScItk8oocy70o5JGz49qFomYgXcBkuo3YeJKPi+ZdKD5aVPA25oOlsZrw
U7yQoGs0S3xDSWejZ8T+HWdGzASN5SgZHhW92nuG5CiGjRtQUKGL415frQFjeXG8h3MX5njzBfCb
A918du3Lv9Qz//8u9VCwAzyvVCMQ+fYqpc53M+0pDT8PFt/6KBMTiy67nnPX6t1vW01XCUWoC/7u
MRL7e7Yh+i3TLP5VnWIxZ5UwXzORHMIr78URfC/hW2ximhLRwe7wP1F0ZBSHYVZAMRIELhTxqzjA
J+XfnxF5nhldvChyc5aC+XvIZRkqT/4cYiHJB51D8Lkgv3RBuH0poc1aUK7U31rluIhCUWAMqNgU
uKd5wALFY4f+yFKWm1QXTrmBG6z2O4N7A1tcKVztzSciVcxwdktvfS0Dt+lK5AuaP3kx/OQEiiqN
lH5vecK78dzl/veogzOS2Y3HGJu2I0Hw8NUVbg6xRemzDjLGwrPMfPNlF2B1g7wQAhzvKm7k5o9J
aCHqBKpgNii4S9GRShLw9ytvJi9dsIqIIshBgrQ3YLWNYmLTESg2D1dG9mU9BE2GUG4PzowkSeys
nfj2YCFmv3qW1Z933US4fBNjmeBtNlcXEZaYMyOUfB2PIJNcPdatbF09RyYdCNuCc1rAmtNkq+i8
+MgasTSamLl6yG++bIosph521/I6VMGvx1cP9/nl5H3hKMaAMTK9cxszswS7hbv5tt6VaLhdhI5+
2titZnmdEx66n75Yd7X+RKVE3oXCJmJi0LMmrKQJlfm0gHDPAiWJfgfThiCG+ZOaLKBMp7FYNc8Z
ZiY2lIYcKgU0S0Y7SxJtPJyt6Y5n+a6WtrjmZSWmbSHVCsl5dVnUJIXaK6yyDHdshjwXvnbKoJKv
THXjeI7kVrEJvWw3JI+kRr33Ne+M7634l3A+CnSa2945Swdrxz2jEjPI3r3okZi4hBgvjfe6d9Uw
isN8TOnrOa/P2xPszHiSm0lSyhcumCEgoUgDK/HPQmWi0Y9iCtvnu46gOmC6ZfbI2Exz1ZBbapvt
W0dnypPpjPM5bStoz3TwuOJZJ5zFCggeSDzJj5Jsg4BeJuZ0sx4IimDsRbp/8fYGK4TGMS70f6yr
21GE8wT9fDF86WQ2MpcpbhG/fbU4p8/yz0wpn3uVTAsp3JZK8d3jIoSEiTHYXImvC+wsXYBvPPE1
ewj8YZJA0YAHzOwUdxgeidnSBKUrD/jJhhz1ztk9HkuaF2Gg9OAPQaUR9MrwftZcNO6OKT3xgQIb
tZzrJxm3LxMNJeRc9hqB8te4tTLFAeSdqQbB8qbcnmsMrCr9E78V6XioBuNYQJGOaJJlDh77zn3n
DQApBwL6RAfwviVSyEM863gWx7t9n2Na6aTjfBaGfQvb1ss/ffPwi9LhYlN/aMshX1cCse2VfYAq
TmOhnJsMLd8aEA7gGnUcurslBGK4rZRFcR0TOX9EEm25qDYB3DoL0U61KuWN+Jhvh9D6l8pXF08f
e1xSmUHPg9xqdhG/mOKQ3O/Yk8B/FRIKCyNns0Vqqo9NcSoekuozxfdm8F4xn2q4wZ5CYSKbcaWN
8Ucw2EST9OP5Y9/D2A9hS+WR6D2bqnO7mSfb8+ntrT2avUGqVWfX+n60l9PJd2U1CUKK9vnscnrq
Z3RmvkWI+vP5/kri84NUmeqcCV/76S/gkLInMDBrAsaNQ3CIh55l2Yqr7ZV8KBskzFm/SHSSbZa8
9K5W9mBCMG4xMyJjYbqosv+jZ0YribzX8h9A0sebQeF4seDZJOYwfjLOZA953AUOyf9ibINeg1+o
UNMbfU7/KR1Oml2SWHf3aIanHZEAMjSoqgAqMDYuVzHKiOaT0fMzNnrfIsi5OfVRETtvEQEfZAFj
JZt+u/GRCS7lXc7WnTnVPnqtQOfn17udgnOClhFtwjN57Qd/zhfBTLYTH4Jxf5LAjtqJDot/dsfK
pcPUBiWwqD/e11cmu1YXdwIy11GqiYn919XrTrms5aqQmtICaf/1+Nv9EQGuHFwewQC6dczW1qZA
scb3eBeWo8fknFmpiJZwEbhWHdWsIh5/4JyiHKJeCN3ZV0bNA6x5+lBtZeaV6Zh4gdpMifT1y2oI
LCBR+irK4dK2k06gS5Av6PZFbvii1nO0R3V0YhGYoEjkP4FIKpAL3Z2L0XUHdRKEFxYPYUD9d2Mt
HBpgmJt402sCCtjGqMl2Y+uVxYci1/ZJwANSxONplIkm2fYJydFt98qYGAmC8XG3LXBtO/RCePtQ
jdPYOGunqehYBxtANVNz+5Y9jOVTROfShHuG9FE0kDdPxuK64xHmCCVBT8MRFbr6ZRAyqA/kYvpV
mQFd6jBTL+9klHUAIfO5wVMbsoAlAnPBC9e5nk+hIodCWHm7RbI722mc3570i7yXP58S1lROF3Kp
vJcVwU1brrl8o3WImLGSyKlu7EQBTndWfUWrxjtAVeh1quEmq+Iw7E4dWkSDxO5POOI5+yWnmWoU
uAlVVVXK5OitD/abU5NTcBRIDfqyqUFCzeI2lZxh0RDgojtaGqtp2SK12HDMRBnh8VxO5WW2M8n3
boa1R6upcoQYfRWnGNqfHfSpxjzkVwsHKjft2p99aAJjr+6V+DhFA478NqrykqgYmkFyzM2FHebd
Pkvzez/U8AdnRKd6WHUntlxZTRKRKeydMMTbdsiw6L0ON9Jatimijk4kH3Wo/D3mgYokDcPvMTz4
9vsyZrOrnxraQr7tL7HiJmgbkoSEXkbNfLm4NMeq5FQHdrVNXWGI7ANjhB5HnDy+/vRFc+mZHsi+
7BCFI1HFEjY9deiwN1Dag481njbwnEetRNtsMxv9bq4jL3bTSUZnAaA6bQzrCBD8x8DcNbwdQ4ew
JYIwCCYfywnWTM3QTl3Q6+TA+4Sg1ZeYea9uuuuMeevxAiLFDQzbKR5VfByMPUY1Qp0u4yqvOp3R
Sk/Blx49Af+ISbBK/CrIkA/n9pa2doiZr5zXKEua4p8usR9qcvLnW0/6Cspz/SGrzClfSHY61ZFm
xlLoHZr6hcTmOCY4VbKetOHKAS0D1eu6Bu7byBR3u4xLDe+iMkzQ+9KrrwXoZwUpHFlH2rGtWTyS
A0nJvj3An2QzyE5zEQrjasHx/KP7MJbXYSTD4qfBg53+9ruc1ZT2jV2He72y6Ez0iXPFHL9Qc6a2
5/DydWJjdjWIQ8AkF5gj+EgGhHQoSpMcewbzRsM63TrRJuknnfEUr/WZ4fuBBY9fSlQhcn8f4pdu
4k6MMmDEjo6YCm1YPYRvPq8fcc2vQx4Kv1cdfLAHUWCrj7cZyDD6tSUoLLmCBm1bwcC0v3OIYhHX
haKRZyNtBe58UdGE3vW+k+BRK6v0EqT2YYX9MlNmbBSQ2nbCe3OmDeUEwa6XT8L2n2j7Na+SXmGY
ZZkmI3R14jcBQ/fcIGnDOeG4GFh2tBPA/4l7bdReiyczjp1ySQpvY9dE8Mt9da3x0jJfyxuDMim0
DGEvMKIlC6B8qJsEW8Q/DUhd/Xfslwc62M/W/NGJ4j3sSGOjvJKotVAX0SQW+lyeK0CsYh0xasKD
XWGoXrPd5UEPVW/SEtl7K0VELDOWBj2lWyf0+fNndozKV2gCXyHaTcWStvSJNR1mu5L1yHpfngkb
Jl5WRkFAg6MpijTOZ0RY/rj+Aqk/7sL6UDsrQKNILHVXgsbYOiuqs8avG1s7oYJK/kmFoSkIYkD4
Dp6VArTqQtUad+gZcjCcbkRdh5EzhXmv32qMAOdsSfbPojy7rkXBseVdLePLpuIl9HltGtAgwG7H
/QtvXvnkKA0o31zeg3JO1u26xrdiJXFjQ+Y0ErYsMUfUAR1h0LNTnGzxDwNE62UzVx3yUfugUUf9
EHjd+iYAZMk0v7uV/2E98+QUMF6K+jLt+bKalj6XP9Z+Y45S9Dbw+fhchFSJGx1b/aSUSXHA9L1Y
0DF47VRUJ2dc5klFN1DwJVJxg+A/MsE9NvW/ryKf/CVt0c8139ZKyUqEbm/R1YeCQtQPVPFILSYS
jCQ2TOc8vQwF3BWUid0geYsnTjqzggzp9sOSYGF6lHxrFMiYx6GM97I8VzbJ6Ippf7UhdvRp9Bt2
fjxGZrljnBTh9JwmFQSfN80efmdjZokxXPweuzdWUazDQaIr3EK/RB3cJtUez5hYLXbOquK0TX7F
jCBIozmtCU6yMEQH3R7q11cMVC9zPeyaVgLAWn5VNLzWH50EX2x9dUfkPDojC90V9/r7G5sbSqwj
XNV/kM32yTiS7cu8qlOy7+eFDTXVLyttG4gSN+tc8CpPoRXr+QeLJW9mR/KQ3Att+tIg7ayPOaVZ
/ij7dJGgFrJ5ho3JA+f0OdW0uL+3kqMeuWIHzpUISrKKWhdUe79uij+Df0vC0jCCIbh2a46h2f7R
saZB3sFn9Vs2ai7zNo35sSGCrUi8mane6b0zlmd6niWbjkYiKi4zIQczHKX3+5j6OIkGdHxtO2Pw
X6LK5rmqsTFiv67TDWT2r7cQqv3T8yPyKInE0k1obKjohWEaUYfK4L0pVLBavb9I0HWac2hqDdtE
Ki65j1nU9Zm7JzM3fTRlURvBulNaHvTFtCiR4U6Nhqj429g+YYHtRY0zy2WuRv7rxCu1GxFr7rq8
Lns4tdQVaOTHe8oYgRRi4VjUdP2aqH7/LaXCT7TSnUGwbNVv2PoW4n+m6+6aeeJ6m2Zj5HJcLPkk
Dnq+++jEkdBD
`protect end_protected
