// the following constant contains the activation code value.
`define C_DRM_ACTIVATION_CODE 128'h91B3A2DF14A8707103420CAE246D3F43
