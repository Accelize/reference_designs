------------------------------------------------------------------------
----
---- This file has been generated the 2021/11/22 - 15:46:18.
---- This file can be used with modelsim tools.
---- This file is not synthesizable and does not target any FPGAs.
---- DRM HDK VERSION 7.0.0.0.
---- DRM VERSION 7.0.0.
----
------------------------------------------------------------------------

`protect begin_protected
`protect version=1
`protect encrypt_agent="Synplify encryptP1735.pl"
`protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`protect encoding=(enctype="base64", line_length=76, bytes=128)
`protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`protect key_block
DlDKYdLCOo8E/iLFdp4m6IO2zBd+8u9ZsKBXK9smRj1iHJnHdGhDGkoltBzNY9kwNcFIcdyPPvuq
+4Iho8E7x+nq0VzsQ9RA9a1kzsEGKaL+XNDLCx5KwUvo1DEypTpaftWk8laimD/XUR1dq1FvKe7Z
78Wj7YlVtnIn1gytg2E=

`protect encoding=(enctype="base64", line_length=76, bytes=906752)
`protect data_method="aes128-cbc"
`protect data_block
U6S8/vPuad0wfc9gQVWL4fXpQZjKXvFI2QzHyPRksWVw/DlYtQvIx8CC3FOI8VijZtFsq1MaTed5
UY8d2jbrNj4iqvjHDbz74FzMr17z78B9G6yCjPN87mtHRxxEHwsV4epsHJ33riwZ6TM9dl30xICM
bzeFJ6KXjbfjKRsZETkybQjVmHl3Pi2sI299SgWT21PIF196PdYdZc03rXZSmLevfdG6u4CdjDxn
Uai4IynelGdxGvA2ruTdLzUnOxzodI3AABTzDpleptB+hNecOfY/4uNqkd7HL4hxSR/EgzleOk6x
pPWyMtK2PVelHMs9zxhHwMqP84yJD9kqBrAM6MT3sxxyGcHtNRFZC8caoqzfG0HpNQR8MmAzulOT
Ub1nUtMtjuLUv5aoJfXxODMD+9cIj+M2VTKPeR8TEWew3oEkEd+Em9PSR0pAHUbHNef6qcQ7zcSf
bKRSjiNkKXJmk6lERqj7k32mR9TTLzRh41dPyD7oFCNUaFQcYMpD6NaKfEnZZH/lv3RPEzpOQK9n
C+rjENHLo9/JxoIMOvnkOSK6SkYm9MBdJKDkduXX46DYvamb84ba2jAD9U3BlSULEZvkVvxF/Edp
D6DuVK/EqxdcTzYV52p++s3UCTAxOZi1SyQsXrWt0njty1IxQBHm8tDj9rrKNTbtZsRLQGikjzyS
PTExuqdrJom9iLztICcdgTKFaONkhTrjd6S/eYTMjRjblKsTiGYVFoumcHkIevrYlFVk+A/pN40h
YQDo14mWke7MiE9CD5b7PTXEyQeMyW8RW11ZB83he0ex7NHmePVHw1a44uh+UtZi9361XNkXGX4A
qiS9dnxon1uRtTeDsg6WqxSdh+cdxEP2EoBKeRi6xQ1pzwB69w590XBuKxp7spHMfmleDx0Ic35/
rlET5ktNssZN0/jy/zPB4WmECQhKMkbp9j0fmc42ABPnla0K2rrXdoIrtLJodiiaNyw4EQJXmAO3
pEDbBclBIe1l1TItMVIMunk3KoY2ZYTcaUyFHKQV5ktKDX7M/tTfnIQT9XBzqa3WVC4qu+hbdmDQ
88w/yuZfdevC94XiqdIPDvYQYKND3QsHn5+ogN9TZuPDq/1TTW9Gqp5xumLvESsw+gyw9agcUPTF
CfUhMPQd2AUS3g+XcgOINs9zQQqTswr6hTwBVf6sTKV8Fplyjr9DX8kfXR6CkYKIgClQJhzKVzRU
VGeRU0H33SpEVed59dKqzoEWW/64X31F5B2L/e7pUdRPlxOxYyNmbW2mNxoYI0Jmw0RIH2N/YQGk
l90KlODSqeCuQIICB8nRhWXh8YZfHGp+5j9xfVFPL1oqaAKIq29H/FwCG79lqAeOeKZE6d1xTZVJ
cycm2UonsdWZ1M6RYQIB81UB77jkqA8HHzB5RVzyAMvxSgy3G8t+gK4V7Yz3NPY8OxdVjxYFtPpK
z+y7/LEymL+N3EiYFu9FyMjlLROYpGf4WvfN910mIqe2a0LCk8KrRsVfFMYODN41sXLyeU7iU6af
g7vYetrwdYe8MuY+0YObbyDfmCDzoc5kmfFhh3SJtAQz3IkuUgCIQAOrcnkSn1+XV6mQXE22gFu7
xeGx1f6TxU1veKuaZ8CpAp+LlHz6nKCSuzA/uwDxuQOEPuQ19F+pXTIWl8pWHbd8b0KZ57G2dWYt
ossQq3nSXVkQkDhSLcnNouVQLW8G10YovbEZvs0iiN/atN8Fi6E50v9VB4PZRLGOu9xxdBt/HTo+
ip81sxRG0UuEgcglbVYyw9eYcl+rPsFCrNKatUfYfZW36RGtHGrN6mQn9kpDDwDPRe6L+R1CXJev
Ve3oH8JjwKp5mjCli7cRG2hkmfSVN3ThdyVdy3WyjTnsFOT7lXgz3aRBU1BkYhqJsKSPWT7lQ4Zs
p+CiowXNKFt6Eg3Ge7sRpby6vIirP5EJFIT7dsBvICBo7Tb8kCtsMYqTcn9qoPuGER7/70PZ91nu
hSkd1Aw4RCLz7X4cLurJoO1TPNTSiuEV49zWRXkFrA7+VSHJ7yGw+uffVN1ZXhglbK1uBI9+yono
FmEACfAogQap1T9oQV18kjaegl+jm9nFnWinKuofdMdYLHCoEd/HBsSpPDK3JIkczlA3YYUL33uO
CgSGmspjbb4S0n5wQ6J4bufHiwkW5IGg/eaTMUkNMPwS9MHErrO2jXH3/EyufOh6N1IQxLb1EjGk
NsqSVNL6VJdM1OZHDybrtGVEkxKJayWNdwRh3eHe5frN8GrvB8009jtXA5EX1JT36gnHYXDFNyXn
2vkS/kJALVLBa5+OVIONj7B++BtRfpNRc7Fe6UeAuuFp5Ku8RIdGa94SHzBpS01eNCuFLyzcazOJ
j1E5XEzq3Gr0GUfpytCn1vp97XWg10ywc1vK+xfUkv3w+lBM5+mYy4SoRy9rZ34PBselbLdiQ6HC
dDy6DDvutWohTR6FlStzwTVIafKBkg9r/qNbu1nqdZ0LIc4iDl5vsqlAJH7HZkTLaSO3QtadZM7P
Ikqrq6LE3Sb030kA95ofkPJ8FT3FhlmiphsGe5yN7gbtaP/6/syd6i9p+p0oChJlNP2fhGgRurGs
ElXI9qijRPbGKj3kSCodRuR4SQkMyAtmimg3MgNtUFngFoMXkYLqtSxRqUi+Sc0HwzNUA02LPyXr
65n+j9nNPO+4cdvOpc6YRZrPfLdvaKtO88YHbjaVgq0/JcM8BX2O0vU3tHMnrAvM+s1GnC7gX6//
1b/1zDmrDX89NLHI6pXgCJ+Dt/S+8btpHH36goaE2r28ib0uUJeNDUEgBetUvKD9Oc3+z/rxlZni
hq474TdZS8CsU5HxFyAhM96DW7ZR5VbaqJotUNaKLPP1IMT1Q0bz+h2wtmpIijgnFVf1Wj+1or4r
krUX+kBWyI0OvzvGKqLJ+8fH/WbSP0URd9j7A6rsH9kyIAubZO38vEWCKzyatApyG0zJadz5uWoy
An+uB+ZT+zo5B2eeE3QXW7oLQ3a2bqQMWgnS/0SLTvzX8ia7A5DQVN/MaqCRMiwE+dMmcmMAF5bE
PC0gGo7+230ZdNoHRhWp9lvakH31oITQuLE0foK/wV7EnAtmM64aOrBftxEs/ltIib/rRbqsz9lX
SImy4p8ZnhH02CbMYirtpJHscTrIxu9Lkfjht9FTJyHAzq3bcko/Z0j0GzqJw/UI4uZIdCjJu1EH
IF4eKS0StKoiKO0tn1ebksQGOtXwrSgGrIAI87YraJ5nGYI3ioAhzauNjeEamtZOaRcPrPUxMP/M
I5SD2LR6ZoKN0WYWjGy8NCtSsaAeJ3rnndHUoVKppYJ6h6Z7Ei93CRihQHgCUCk2teZMXjixC1cr
fril5DpxPcUOZyceKlsWti21pg71Sd8/IZOrf1n1xbljXVExLCBe9so/fUFFYgfSp5WG20qxC8LQ
KGuDBn1GECp5lyIrMMCNGxtLKs9JWRDYjYcSjPHOY8KGCpEwMQM80u6D94m5SGzL2GZDr7ErP+71
gOG3aaCHu/8HudfKPykwIZQizMr/YHVkf8To9Y8MCENuvZpyG6RfZYiGasq5FBD3KtdjMZhJZN0/
Zecsd6OzHTY/9SrCOjTBm6XkPNQeHp/11iJTjzMqiJ+S74k+ATLBgNvZUMI5KddsIb6liCIUjlJX
SgHJyqY7a8LGaxpazKg2u/Vnfq6Ox1tZJzKpR++u/B/LmLHKtA1JjSUqJsUB5J/z7wWMrk2riwJO
O8ZUSZVBbND8XusPidhKh0GAEzWx8Eyf7w4oTAo8j4Rncngm7LvBsUgs+iGLjb3Sv5ehtVIs5SCv
NymUowiqaWOiKzimjOsHqhOU6hnLVGZiOkGCbX7ltmPQn5UceCXfzL7BC8Mif3Otx9b9qlBt/lpB
IHjn2fuYXoI9HkD4dFwZl7mNXRpDSabOlAnAhFwSlL54TGnNe1q9Yxkh2G0WG9kky2nw6ur8CrDi
IiS9du8e07mHBxbAtMBe80kvQmMbFSnm6lU8RjgsMTDhEToXvjURzI0nknZ5OQ6tTE9HpMTrBLmW
h11aMdwr/Ug3zp+STCzSBhesmzp4eQK057l5pYxyyjfj6BLDmb4HmrVtykZnwhtqRADoyZw/vePG
/xJju+3BnAPsCe52Dq++TebmgDNSLa1UYcS1JBqNx7STxVLSSxxMg4O+gYauWpTBCURkMs7CQw4Z
IIpzMSRbPrL9iER8AoAP6Si3vuv78bq1bUH8hTshtEF9xK/Big4rf1Cw0voCOamVlZuO11mq+c9D
eN+RnSrBUPFfOmneJJyx5Cb0TyjnJRJ3xq8zFw5YlSMiR/hZsXugHJONZZI9+8gdDt8PTu27C6dE
MKsmgiG5KcrewaHFV33RhYrnVwLQKscZ2xB1sqJzYtpYcVzSQrhCj9dIoapMgdYRPFZuCKA0RUkf
8JScyNv5aFNqleSWbiWpE6MnrRmdcD4kLUGsJgGRdSmn42O0pBlM01C5uzzIp2xs8b2nGe1aa/wM
AeOaPURqsjz0B3zgWY5aSBZzEugoRKI9YdWPy62uceLtutoM+65gGAWiZkLkgkJpGzUpoRP8+lya
E+qAhxmJlFA9E40XzPxgMvcIfmgaPHmIN+pP1MCYPUKvub/z7wGRdnDAtad0iQzum3YrMVqporCY
5c+ttm77m78qcxTHcbMz53G3xxSTTnbj41Y7BERq6FaKUrK8uwgzYik0CNAWRFdg8rbccfDIGZRA
//6dLqk778jcq9hkkmgAaOfY9w23D3bBNsf75/qdYMEZ8vqIv5j9W82L4UCIpUaj19ktE/rNYJD7
n75SsjlF4rG4ISdQ/j89Dcqzbs+pObOQwuQ1kVklHYE+3Em4xYYXfralS0JLP66h2r/im45zyvFC
o1M7KKnoItLGupHByYJjIhROvXHO9oqKrqSDTIf/LHWHj/4UCKNvLctOWyLVrKsJ1dtR5VuViOTO
evN2dnSgs7UiY/gsk7mXxsr+1xkuBH6b69d7RLicMwGUCNbagoQELHbmRWdt9Q6OTIuDS9kRwY67
qP3lQbhDfa+gIK1P6s3V9rIBfq9W9+Lh8RHckiMzF10SYlbrVBat4U75NYGJ2Z/YzyHjm5103o8u
0ewft5wPcWGjN8LsbFUSd51cNCF0nMx6TxUnURYjoxzMm8HJW2qCGdizHrzVBGq4XUbgbZfBxlzk
tUGO4jNP0EKlWZ289rk3oig3eQY96D5I4SxyCN9yFLjvp9jqgGL69g9QIuMZoviNZB1/7xAbfyX9
D/bO3IzdlPCEqqieOvPmImwNhJdulHXvrjLaSxJEF+ApT6Y5rYvzY6GN9d61kBhQ8Gfdw3zouHlg
he2BK1dcWW20NFLG++vQzyHB3dHCGVKPTk/QlxggYVnFvx+9naTbJ8BsBtYUvOKg/6zevAzaxsv7
ScVIJmbzBWZQFc5D5Kmo0atDmjBFzWn7i360Xtcvi8dqpbDSDQiorAWIK9eMciatoD1JEIlHRpPl
I5fstK+xgKKmIsZInc3I6GFEhKsMQAPG6z6chtLTv1sI3grjBSl1EtLNMwk8SKsUIeLJfmHKv5Ef
zqngWgsZRjpukah9DWu0ORMK6LwGW2ZIDzCRl8O7v+/CHe+9l34MKW7ZHrNvTLsFPU1iMy6ySlP/
V50gTITcT1zGEm9RUIEw5LbAbZnClES+Zdfx1gzC0OBUeGPdkeHlkwHNRywwjp36LWO6Pa+E2kcr
ngI1CjtFbv7VsGhPmL+bE7NhmxRwPXlhcl5dfSFWmSGFuglPGyQQUIPLAy/an5/EFMW8QHn+VayU
6NnbAGZ2wH7cUKQ9/zusH7/GwBF7KX052+gmH8ugZUUFdOhjTN3dzZ0g3CpySoLZpn2yY7bsCKbn
eDyWDD/axzgbdcHHy3we5hGZhiRf7hcqYnonaPjRt/PVauGv4qF04Ce5qLqlma5nCYbuMd0myO/a
/VEQLO/VPBECwG826ASx6xueDa+BqS0xmBbbZJeTd9D9fmEtYWYoSvq2LKXYGEYxUqAi7fePZRmE
8e4+7hB1Tksx2RZ/FtbMLYUFsUJ3kC9/xvh1HRHwAIMDgombywWgi/ozvIM2r6ZlnHYcrTLvtntR
HbQmaPxbedhKIcs6vWY4+tU0/+7z4o7GV/ZvwRLNCeowGMhikFgBbtglMVwTRizxPVhtJPIGht+I
Aw0JrmS3sylRZKeCQ5BlijU4iP5nkWkWIN+d4DPGSabIEssMLt3EDml0Ke9YInclB4/pE7vmDI65
THoD4+kWp89XhP8R402BsceQup8CiW18m1H11j4lzOJaXXPtYvzKTyqPtE32mCrdpfQSztySFVmN
I+bzxCZVPbWn5FirflbYOcRc5QWJ1w20kOB+c4oVNwIxep5FXjU+R1LXp0PB7S57OVevOBUX1Zmh
QzYKz18umKrleHUY2yUv8ekQ8BEk80dwfzVoOp+uR+Axq+CaH8Y6jKNHfIqz/Ug0EKkbi2DKGT7q
UFSWvZR/hyrkYSu7iJZln+jQn69ZaLomrSDgaBM4bycjU+9v6jJLc30eR5Hcs5/chU19VhCfiRV/
UNDSJIdhlHGSETjkJJevfM0DtSSeYkhORE8juKPaGi4vPbsRJ0YX3If742Mp+xjCdcptQKSBTMLj
Tuf4KUm/VqB+qboMuzQWK22vdkwqyGAm/TF4I3oLY8nieQfpVHtdzMBgeAOnIgI0DVPD3hK/iWQ3
VTpYS0VWjcLT5zK5lmWjRydZylUF5rLCR5NeBa9Tsb3/Y13nssqB/egdIIJJ8ciRx/UG3t25nnLZ
eb6aBrXZ9/XtTTujrHODD2xN28Vs92Um5m5IXefW/ilXQYXFSW52RtwDdqe69QZMiUl8FL7dhUBr
b191m064++1oMfHq38+2w+HAKMa6c3pvUg/NOvU+O5Rd47LlyIIhg9S5qczjEBSub9wrWYqIlexm
Lrxaq/KkTpreW/JdcA+4TgFC+/3FdXPqT7hURtFqmbiCIrR3SQucSWYA6syfWa0V53tcLLasrN3p
tSZo5ssSK8m2pQcGW+WQCfWkGmda5WdGgz1m66wuqC8sjuuJl00vpr9TyOx5SBLJxnlV/3v4C7oP
+lgDehANolc0j9OZ7+YZxl59x1rsPEvWTVbiAWCoqEBECVOnZcPU0WTf/XnrdlQFdOqfuKfDBr68
18kqnZ7/ivJSzmy8LnHnUt0dtDhmLwOC/h0LvqH7YiH74Qf7//7KItcyxlEZp9ARd49af3mjyj00
2DriUgPQHNdhhts0vhYqa2g3zu9fgPTrEq26ZzhrjCZlfc2s94NvOZDaxdrk9dvDYK6ztX23eoh/
diVTkijv3WO4fnuHtq51/VQafokqzd0VMX7dGcIBYZEKBT61CIraXxVgPqFZTqbEn2KBdXNj8iDv
4DSwwhYRfWmyQJWX3yQHBH3M7zarhp6IEOAv3OU7k2kQ7VDdqGr1Q/uwUrG0FPod3Jv08npMtB7F
DrKhY472uhCOrXFu0NWLLyYVqvEdQWnBVck5c4I1esXmZw8WEg7Eb9VGHTTPwLO7DLuA8QQg/fxF
tBip7vYyrwC/VtcOEH8eNwq/KvRPdxDC082QKyei3UJYoqFqJGggimYY9JtsmwjiSvShZw5nwdMo
ARIulBNPsJVB0vAre2P5WRh0ApnkAppz7+z7GOOZ97oFa8y1x3EFUphJLI3QppwPcFKcxQC1UGKj
jEJTjh5noBDCVqDyKENYIDdYpaVc16WvLznCSwXaChRg4mbKaR5o53nXBb3gLqC1VYGnz3uJOCCJ
sy+nJhEaKb8bLtEcA7ilRRLHl1difAmw7gHqGe+2Mm2rnAvu7nTJAwI6eRYDTsFrLpU6c6dQkxFx
dnme6fTA3Sod4rrO3gL2OsafiiGmRALu6NxKi7+5IIHmgBWRKIg/c8VK4HuBVYjrfp7Sncl5PNCd
/WdGdNQaNy5T706iosWwP8WXGxiJp7Dpm0L07SSQ95ZoZ9kAtzrx8dmHQnzzXX19vfJRqveWrnin
xI3bSWDRCOZJY7hlPU8fDy9ODuUimPXwiuMVmKEDVEJTmyFYO0tk/OMTJWAdEQZ5OKDPkMnIs038
LbT4O1+/7+xlUbhJPukIezSGiE/H9luNde0MQyN/j+UOQrAuIwaLsdaUBru/CnNgG7kAEeCGI9+Q
50IlvUFnN4L+5kgGAaAzpI3gdR6q+w9BnNbbLvUaygamySFNqks+w2WV1BHik7hBOYFnhUYSrhe/
gUdxIcl+lW9B/V3IORnGeUfiI1GeqZKSn2RYHLs/ytcGrldwptTWbOnp6H6Nb8Dd4BmT9dI+08RQ
pQ2vSaLfEp+SJ6rLslhmaaU1DMnZGIC4Qcy88VPAOihzZVFj1qF6K6ybuyBHiwfwH2qfU9EEI9ot
3tT1+LkDw+mH7eH/R3kZb1VYF1X03BOEdabCwc8aFCvnw3cogSjiIjdhgsXacsXHoLDehKevbI5x
nHNNe7Uw7H8NquTG0vwdllzdrs1yNuBLwa308nn72va/EKEiEXVwv7QlbpMg/b+8X6tm5nWqVVnD
PNjuJWiic014f2CdgQcPcjsgZTV/MUf1SFQ3FTqyvpJJgSDl3VU7mujWv9gXrNZCjTRUp5taonrt
VXIN/wtKldTz4eCNHj8yDVMP2AvJRGyDzFxn5Moj5pDQNox6SI4z+LQNr6inm+5Mvnt4KpTh97ZC
Auvf8SpJgSK+wihdAp2T2EqHDARHpLl9GWPVkfk9+f4qNq46gKg+tfCSvtDz4iz1tEajAGIEkGv7
n1LeU8HeNxMd+8D/QlMvQ6ikJh1f81zuUjZpRtf2fwKIwqIVsFM5mAAcbewOmUcTR8J+2iGooY+A
H55b8quPLX6L6GmPgswS42o+wB7gJYBP2i/Zs9Xsoco3kAzj649/YBH1Jd0uYjd+FKdFBa05KJfu
JGZ0NlnhYrOTjFDhClC2wZ3rV72TVuwW0IDlGg/pBd4Ei9pr/A/9Vt9idgnUpemAWsYtU29CHyB9
PFjDBRXmMlpnitjAc8N8BwgYTZYCuIVE2jhRQhKnoXV3hsgyRSgVNcZUE0dcnrDC/mLCK0wXmJ+r
IcT5ntRvKUPCXy2c5MJznCZcTGW9hts0WvfcSF/eZdIdcS5hLfdjuSLJvhrfVvFhu52pl/UUWTld
3fLghh1e3gyN0SZzviufMPH3kU8dqY21HVwf4Ca8dxq/wYUslAl9rxoRjLQQxdc0JWb11PGLrBbI
4R2YUz7qKtbZvt0CEPCs/az5jLhMGhbUoKPpoxVpDaXiUw/WePJPtu267rYDhgaMV0JdLTCr6kim
IocBUanr0A/7goKEQkKN228xgvhNc2rC+mD4sHgG4tdOELMxG08ecGq7Nj5HlMZ18USMViQurOm/
IvtQnS3j0OkyeMIGDwALWHOa1HBo2+UOiLZeji9zDpsd/SNSaOj4SoqIkWY6zPT6oYAcfNssYZk1
oSSR41Pz4GtzaniTWabToUKEcXrPkiez+3twZwB5ZuGVJRry8ZmnE0iPCi19NFxqrip78HtWscKy
ZVEw+UnPlC/gLPF3ih8qC0FBwBa1R7eVJBt6uC+AwKBGimbQKtnA8RV9QVox1AQ6b4DQtktb4iwf
2pxQ02IoNib+3vjLJPvjL+rksXApjeGMpCGhlAyzGDcU699vHRWcIHmzjRIIfg6v/xVUQLjr5jDc
2OEFlDp8i/w32PkWFH6aGG/xSOBWWA+VcbQTHdzYLJ3NRAcZUeclQO+ToN8PqlELuLSS0hj1ogL2
wtr+qaH/vBLfJpGAvNMmRecTKdUGm4KUTqgrnMgRZCKFz+9/97zdaIciuuQZYVlXWRJFPDN8GNxd
Dr06hL8aXU+c4nhbxvDNl6iLSHH6Pcx0FjOcFkmjXspA9wHZCXeOoAZS56ymod6t1n6h74cCM3gA
abIK0tLmG+lLCjZdcNkOe3q1RdWiLE4JhaPes0MxFC+3v0zOQwsHcQQhfRX79jrDUNdraxpGFBO0
fbZtTnp2OSoZBRn4nKt57ybI4ENV+p2DTMZzWV9FXVsvc/Dfs9b/yMX4py33mZd2716o4i5wd8eq
zalFUpy7Tf1JKPVXermsCXKVtQK4paQ3TdS3ye2Fju9HwOlCT+i8Au+OPkJISxsGg/8sutgpXxeu
6ZESi2OCtdzbL+tuSYAMzwVZSEN6v9IZs37xzsPeByl9IpEqb+9Z0vEh/N4YGwgDyOzcwrLJMIVM
/uSVL1/wH79kO+nmVslVCGJ1ymlxR1UFFuyRHN3LGTcJ+zRb0U9dlxHqappPec7qVY0WUxMCGnkj
wIx3hptpfNlT+wM36Sd+gqZK+eWzio7CGHCDPsgpjYzzaLY0coY6GiRrTKvbDMOf83jwk8jGMuBQ
brZCSmluhXdmlA2fgkoh44Rm3qsIcUvioETTPmirQtQqIsf2ZySacbxESbM65ydNYpO+we85ZdGo
dgba00tJdg25rkOLhU9rPo6ouZ2pnloe89iGV37ugFDtfN14dSA+fjdnnfbWPHmsHx6GpVPoF8Yt
mhyNkFuBqQwq4+OiSSB+AnPs0fXpKpAE8Hk5NQkKE14kXVaJ/2yjvqfMPRN/U4982ANXpfQo2ugt
ocBeq/QQ3usmr4If+pBHNilGXKwD9RB3KVM9SXU6ZgMDnQWkZ8G4lRjZeX5SLwLIoY10HrmSGAMl
fzuf3ObjHuV6S9rakk7T0Aj5h7sIWAIgob7kA8I89PH7WHjOzFh5ZS8c1vGve1VgD0HG/z2uQCK9
VBkrW9W0Sp2D8qSXV1ublw2Wnkdk/f5Z5cL+IaCQiz8ga3BACyLrifdDMv/IllHP0ndJH7EiSSgG
AUpAcmXEjoCN2gvifJjZD8NADBQ0yYTR7aT3/jMWn+LR46R9DlYKzk48ECXob8xuRrNoxbKdMqSz
hrcK1gEwjLZDgw4PxivvxkeP71o51JojYMyQ20jWeR5Yep/1p3EK4R2N1+zDX6scW4jEVBwkg8ip
0XGfXM2b7qNX2R00Ja4GYPKUeHOxZ77/4/QXRPlpvarcM0UABGU+JldGNKJFfk+BR8zUsr9p8EDO
dYWAPIbKNUnhG90n+h6mWnAHGDg278fgcqruzsIGn4F9zOBpv2N6ww+oznPD1MZPTNVauxpWWqU7
uojR7xCdnBEFGFjhvuFxNJ/GdboCyrOBYulTNSI7677VWKjEAUA3mfXq8ZfOLPPNrOWlvu2MsR7t
xEnls1aMKpERap/8HKpYa5lwR1i9sGGn5F1EZAk6Sy8ZchObvTtF8ZllE0HzgtC1miImaKXr4XF/
slQL3HwU8R6GL+OLnYyBL1IavkJ+1L7kLslNdmFlWSES6EBTfI8Z3y5VJtzZJk5OikXkSiVZx51F
pOPmhcbK8yAw+dFXeP30BppjTDHZNaoiRxTycKIk54CBDbOk75Isohcoqw8RqnoFPSQy0TkHV8qZ
Oplfjil0uI0/l6jXqQsR6lQdXFit0Y4/O6sb304WScLyTwNBFHP8WPtXXxWbDdGd21JgXSpMswD9
EHGJuGXYW9dNCzRqBQN6ynZ5n/lr8H1HXhcQ/kGpVJYewY5FJHy22mptvtS9KBTWr/o1v9RB9+v+
AKDcHeSN8E8ynCku4RKNdE0630I3+JxObmcrwoGKnJi190v9QvAv09fRrNkDLjxP6jFRkHwFTQLr
5UC2C2rfIL+Uc79eZ2tvvcxLrMW4e1F8zWFNt3gv/SzZU1tE94syfHAo3iM/IDhal04kLJeYZyuN
yj0UFYJAn9KZFJO7JScx4z48b0+iTLYY332EUGNuzrufrzllaO3I7c2ngedeTf1JI1teoT3emwFE
lg94hmO3cZITVsG7ESjEizBTgkPKX+U45EJzgtimN6AgNJJs3V/YYM2OZKdIWcC6Zcg/L1sJflQR
cgMj12vkd05mutEMvyrtu5kXXyl0PQGUMAvDl4NuJPFBYzWTc559snkFTKI+XphjKpy+X9UgUpH4
cxJENmFesFtTRhy0kVFbmV6HbdrYiWzq1Kr77/gfhrQC1bAOOIPn/5Y/xfpG6nWxPzONa+ubxtGM
hxOWSSeR1BdaDasbVriwgvTTvLSf9GTA2N9VAo21vog1DrFCWlX62eNHlmiNPLwDSDqfHg69IR1A
KI5fhpeYSsHsyPTouQnw2bJ8TKFHJwf5tTqUA05IiqqNVPpnXKQHpUNBNdzea/FSqRFPT1otQL7/
HIkXzDk7Y03uw190qo/Pr9rrcoQcT/GXNNAFPrUyKEzoIy0FgjbNRSYV0gg7yUuIALHmZzUMzv1a
UCoFTshss3pVmHEoRByDtUb4FejcfhbUjeFeN7t9d+Y/36qaAk+Af2YQXD5C/HY0CsjFwfQZDVTt
3yG+yISDPv6kQx6C/VAXjkd6ZNwY1svuFpa1v70EtQ/7kK8igXmQJfsx7UmuFRyT8b8pJtFGmqym
RXTSzpJCNdT4HT8BFGXvA+NETYA5/CTAFIcn9qzrBwDBi290g36yiYGo3aA7uJt23MhVQtNyU/Cb
znNcWd71ORABcI8kYCEEX1qoxY1IRNTbUZExk46Td77giYXZtmfU84qY2lRs0GenQSJQ+rPjf3lX
vucwEMB5P1A+QPNJVphMZH5M0Aegh3VPQhgf3ZAxAlE5/cGqdAGhqTTlt36FGD3Xi64igaixz9Ze
fhT8dvMuywP2jjcGOg+FReFRllFEwFXxj1t/dqfII+NKFHHWxKmI0+BSJ5CMA4c9RBlJpOeUqSb0
OvwqBhvSuvpIhTVpW+wHvEzjLmF9M25aDpUMMZuRQGeMXDNnkOfaLi2ANHtSk7mmn/ZtStw76R5Y
d6VKO5R6c/ret54WTc9hpWW47PeULUiScW2IBTigUEVC9elmOPSVi8H/syNq1XsQoC5CuaOuie0G
IAUjVgFGz83yozpyq8O28JMdkT58gsAhGWTwZbMSh/g6Mby5ektID04TENwp6IFu6/G3kHM4ohsB
XWRqdLJnUGtZEDfwC7nvcLikPAMBbX6FjMB13uS8QM+Fs0QuFxoZG4A//DAfvWWEuuPnljewqrZy
m70PZVxSyE90AMwfURCOgA2NH4RHc2IInaOQrJY/20S9VkvqGDMXFb0AjH2u1EgK2FAkl01Tsmct
oJ5WfxVvDJh1eQxthGlRgPi56MzBfD0PRs+fFT2CiTetYxQK75LNp6lTQzSoLL9Bqui85HSrhc+d
mrkafry0/QtSyxLhmctVuH/HiaZOQDRpMxtjM/4LAvx/Qp9mhUiqFB09xN4XiyzOWOWxryIZodJS
4TdXS+5EAuHQKl0rbkbF4BcOFe2/VJYt4FJuxmPhs3ZtQRt+QadDL5Aib90Wan9bjfQ4rQ28qE3e
21qbIS8JvXSRAJ69tjKqQxmjt2QnckeyCZgp/YqRtMqzfmyearJN7EZ2LMHkLTFs1flbOAiLLhYZ
IA0c+PoBkqJpFFQOZWlv87FNADJpIq8qtVnwm9X7nkoZ8WkAvQ3lKCPPgiKbQsYH+r3SkuyHKgYi
4+eFwUEy9B+aKq2XjIWCIXLQZ+YrL+PDvO/HZoB1GivZ2lg/kCFWL+vnuwtwx+fJfqhUjXpEwDlY
+L5EeoOPkzzOQkGzfEhZLO4eZJ5asJ3/zWOMtcv3tZHlw8fWTUSLpaGOTBJ0qRYCHmOvK21mHRGz
KA0YHIvFy6jGk+u+9tRxgzNccmHwztNFLKkNS3kVaeiL7K+g5rw19+PGxOToIv10lJ+6BCXqh9mC
7FsoRmWdDl9lrx/TOzqhn29KIgImhoNzkIZmFF718/HmmXq/dktEoMyZQWlgerBVbdgMt7i81zA/
d4GSBd0qzt01sjx7t5SC1xzHUq3RTSzBedalHhMSzRQXXcwiIAnKFq+ibi7uB77I6XTqGCFpcT9Y
IHI4zniUdqWr7oq3MeM/eGahvcU3MUeh/3vdEz5a8hhQ56/3+75gzEOrL/OfjYk2rDpFsI84y3HT
nFirl0DsVOEA8W/O+aouOyGzb+RQ/jGQmxVe8Tr1yMCJ+ZGZGrR8GJcwb/xNpU6Epr1gKuoktAly
HXzYxDMbS2Ul5g2jQyrzLfg00pP9q0wHy3oEMfP6opgCgUZ8KBeJesl7OmxYuI3xs/g+NGvs+YoF
pDV3IwZ3ufRVtAe9i2DtfVneTNBEnkWseyfLVg0wnVHJKZX32qFlycfUbOsDzHFcwdhsUEYQqwsW
77MD+NgILy2pMYeOOPkiqUuAoc6q3opoe2MgJdEu31tgwkRVHeiK3SfB64RTmS+OiWXxF4r2v7O7
PeQ76YBsGv1lhhXQeVL0zWJ+N7FiVr4OJHhYiGCmKkJ5FDirVkOGuACjMN/u77Jbl5uWF6bxbkr/
A0Ce5P3UL7xrOsQ+rFq3Kh8sHNO4MUu9ElKsuksDEHSmZmc6rT0r2WB+pyNjy4aD3fscOQ4S1Pu7
9QBKUJZNtOklnX1LVOkkWqwUVDUiBc+EUJ2fmqFSIWBfnXTUQb5X78bx0m+T4FF2mgyrFQdZ1Cxj
0kJc424y0NZO62kVEl9cj8RABPiGzxCD2ZVTiEBJbBgc9+LWrbi0JPcXze93kk0BTnOr3YJbinWO
fhkJARHvs5Ir/RFuV2Rr7O5tzw/xyILHF5F8kTg1MufpmM0X5afJebrbSQGOMSGlSEZ6ozuBg7D8
ld2iRlW3NzyHXok7cIpU/1OnVjYDsR5leJLXPKZwyXkFHg4WRVH93eqPnpslEUQ6mrUvt3MfBzUb
p0S7s830j2LI66fErxwUFzeBWjch8/kv7P2BkskZis1OveSQR8cYr66p225IBbzYCYCOzObzBk+a
joAWwECRHlUwlaho1gtj4+jK9Tp8u/D11hchgsB7X5rBKdSN9XfSv+5pbi3o1xQedVEOJb9lGovF
eQEudEPhIRDQXsGUEShbML7EjpQKOx7QDFyl9Jl7OquU+JkjI5Xgxs/yPepktDUIustiAnREQR9n
4HXpZfj1bX80hhd7sNUm9WStSVnldG6aZCPlVWxeTQ51fgTvd+gAAXE82T7EFCowrjFXeKxfr22R
juNyJnnR4wL38YWs23SuBDd5PMreLb1/Vtkzg1833S+kHGFBolyeRMFJ3SSQB1SGoiG9PsSMjWNG
z72BMK3MdVB/AeUWJAn+Mv7uMfj7Mbw2Xg5OgTruilaRRSbIRxa+20/jfxJ3s+daF4K7z8z1j7v6
KXS4uvKz0Rqb3YEoR1ROlF5KChAEOFeweEeCXjjjxdNyIPBgpeH0X2Fs9vPO7xQLBmcgJtVV7P8z
UtjqmDb1pnwDNaHO3n3wnsOHFd+GTOtMzwsA7l7QCOmbCXktCQp+QlfD3+bIV9ZY4xVk5IFhdu7z
8dt+Q1zr7u7RsZs7ZGdcVDgu6yqw0nUqpmLQwDkTSjRKYyuHltlOeTVzmDAb8A2PuIkFD6lJd+Ou
/Gq1wvc9p3q+oYJh1arnc2lw4zhQm57AgnE1Rr5Dh+tvU5q7jFvKbQA6WUgc0AvcAf382AFluYXZ
FPNSqg9XkBsPvYBQjDcDc6FY0Q4pnUvOqpRfq8kSD14krnU7b85yDVlJIRj7CfT2KA32C6kksmvP
NuHEcrppjfy0vcUzB4/EORrRUWVG6yhGnknmP4DNIsLkPA4xATbyeBcM1cwQ9Bx0TUqDfyoeIbJw
nr4LbV5Tlg7hMtBmHCGAV6RoD9W7qRacWzP5cugf1t3trBuVEn+KTA0N9vs77RMg4xCyCT8rfzCx
H3Vs28U8YC/L/I6nJyfzjSyBxoC3oYcufoIltJKOT8BzQpszb6tBqTyNw4FSrPrfphwt54qnNOXl
GJVdtKD4+Y3+6ycI73bAMpaeUShTxQ+bK0e6xpXzRDOSZPi16vqrBkORsv779airGAlEIzkP2Gyg
ESjx9f4pWCp33AOtRc0zCPXcibyi/bp3aj+wwOTe0UFDT8o2u4cjU+86J7aUInCvdNcEmoesAwC5
J+/vr+4dX8fhiaBZTFfO2sjsVX9VAwydIctXocnO3ACcctcDY67+FbyPXXILxewYOrP+tSQbVoTL
TnLk6Mnk47Ej85VHbJkYbAS6qGRHX7cwUKtr9KpHYeEeBojZvq8X30odIubWi/ywsarGNwbRH4Zq
xfk8WsP85kq5pCozaen7798bSNn6pSX1CYZjT39RWL6BXh8+V9DjV30VByQzc95E16QTDkhbbcvJ
M2lzO7BAJwkyFPxEWCOhuserUVsjK4ppZl2Q6idtjSlPLwx3T/kRz59BVLsWL1uEfeQ9FtGVi8jj
ys7C38sKDMLgoFo6t8X03k0d9lEp4SEVN12wOA1jsM0vVc0TwlPy+dvUAInPf9nFa2jdt+Eo/uZI
oT4hu08iB8uFYVvpMd0/HYLPPLuKJcj6u4Pl+PzpIRYnQQWVLCveCDxYi9OGoVtEdMbVQ5eXpW4S
EnYiKqFou3Bt4S6QDhF7AAfjeueH69UqIsIN4XQAPHrCcf5kW02yH6PZj8SESL9pclFUqrnhd+qK
e5DB2XTJH9t4drAWlZm+SA/Qjs7qikg8h+lqZfvO19x4+9DdToyOWB6vrr5KtZp5DOsusCDcJxaB
3X2L5aRrq7DpOuqpZxt+KDUVDKTkb9xURHc9E0+B5sTDHD9VtM/B7QuuaToHoWi9oQu3rYM8fPLN
7WZAhJMplgg+fr86rCPsbl1ssE8VuO/8gOhO+3KVqwP57cEFrWlxcF65wOAednwAdJGVdtYzmaqV
V1l0H70WnL6BeKPHC6zyto/0b8fYRLapWlPViSk6U2aQUBnLbHFqrGsyf/Vt7kTbsBqpoClZQoZJ
H9tI2bg7snIRIRw3NsaTrZNjlWTdS7itnF233sv/Ijxdr9W9hOzMsBglfiwbSQzcfeGU+G86nRuP
DRRqE5R7qQIsq4qdC+On6vBRTabdaxB/osIjErhyBpdIzJLecr+zZtA0/e6t+yIUMrLTFC2ig5ju
A6T6gcX1iCar6Vm6jVScCgw91HZJeRcXVOWiiyQs/pWzddoTfMPu+KcJle425GzCLBWnnKES4tfs
lX46lxB9FHKMH60lPwBjootruCz+kfKM6J8lCn3yllwmVqbuWOb6PrE4uG+nNaGhkTcI7KAa8V0I
HzKQeU+tKxBzlXRTBKQ+H5db2bA5MQLECfMMdHiv1laGEIJaeOkxqZjDYtSkNV9H+mGL2ebMD5p+
DpU9d35zflwR3dm4QSQEbNPGurKNdq3DaUgyyCYLaGToJGDpGsEjOzUjs9c8Torz6ZyzGsZmznL9
Aw3r3uqj8rg9Yfy1IOcqdsepsq4qQupFHns1rsSxs0ch4NDUsHBH+QKqXO3mS/46KUYUJDQyDNdV
rvohwwSNBOQcCtnxSn3DdOLcD2Yaapp6ew9huBkMc4KQh1J/qyrQ7MGv3EySW5xs0LgIkdKhrQNW
xX1OOswqC83mSE/y3w2GDzyK8doHAyVbTLcUl0XzNoHrk/oNbjYWf8rWgQUZIVDHSYRW8PmwRZz8
HXq90CN9geeOQsWwQxkAAhiEcRt1SCQMjGKNAC30UOWqLmANZre5msv2W5eLpHDx+JOcMKIEiWEY
ZQagPdK/y876Ebd+fhI7Rh9FPMpL1gRsyoqufRkAs1tZVPUKwvCmwpoS9Py8Y84fkRJU8r3DfzFn
XuslwLizhq3dydn0NeJqvR8n+rHoPMskNGUAGM9tTGwPswc93Rk65XyKTbXJ6fgyNQtJAyTTnXSG
qTm5B5fClFg28unb/TkCNXXwruGNahEhfwLy/h+X9CouIJBS6RlmOCeFm6Hz05NwfkPORNPziO38
kI27nOaA4CoiULdUhBnehTF9oukooOtY/wGZT2NYnpU3Zf1unaA+JDroyjJ069iTNVa0CPPBFvIB
DwvlO5reXuDpoHn9dKINnIniB6+O02kV3q0p/iKMJ7w1lcIRPUpNs/Lu5qvzyBc+t0uaRsuRfbJu
YVBjJnH1AkwK57janOyfIVH8EYfsiPM6yHPyfy1opDabVL1C5V0yS8UOj8oD9HYHPH00fz2rZjvv
fWr0+UifxPaqmQLitmrre5T2wukebTo/nWy1bKscus/XJGnRSgK9EHQCuKLBFQmc4ohrCVPAwsQv
5BUb9ptlyBnB+qAKAiMMDxszQXgSS2wCwhLI+d5D90W76q2AIttMoZtEwpHfsDZVUlvmdZNqTh5K
LvvPmWVi+TdNtNGOav9OrcItKnkZSJWx5GN3Gxm8ND9IuTKHezWdmlUwwlr97kG3HTR8+izCBS/B
8I89APAlMMVxiUByRuQUs80WhSdnx3NV7UGqJdnUl5ADea714AhwasWvxB7tMliVCDk+nRHnUTz+
kFtA6132eiZ2gio2F2l1uIGK8kqXXXuVeDQrwa4awQDtd3I0sqRj8Z88Tci7SH3FGoLYlOw0+HeV
yjyF33FxFduh8GKSqLeVWFQ83NG2+nBtlIEmBnZyhd+ZT1BtWK4petrxH7l9x1nojEVR1aCgwGSv
rIyHacQo4qfulhbXQ4il45b5SRIXx8ZY/j2920ohV+xa52ypnosfYPJAXDX9nENprncyuUHfOmT5
n988tmLo0sE9bTk9VLeOHqL53e+0nYea2fAta3DkLslhksfROnuP9RL/32biQrmwgLk5O2xnJQXo
4NaSFBFGlCZ1bN92XoBcZv3X5Um9LPLqPvdyb8wcQ2rfO7EFxyWjyPoEpZyhJdlv4Z9FpuiGlygN
j9/IjA8QqcgU597aOCq5vzhN8IoaZtAkuf0lcgs6KN88F7ZdkBOmdjf8869ZbFjaUHzH8FOE74ss
0wPPp2Lae2XExheHUEm1Ri7NUzsg7gXWnk/SR6kH+NarKtUHe5OUyxucsyegdlm5FoHpygQJBESR
xTJ42bpu5V5LjLcsUtdaueFjDIV+7ExPWuINHa0pKe9r4AZTMC8Tg+p86PH3L0pFWLZR8Y9Np7c7
rRyhAXrzR/lw2BBvfqAByUmZvAOkEXWP5hNaYTL2o6Z3a1x3zzCStNdtsoUmnB4YPIrDkbL1/Fxo
NJNJoCNTRK5EcaDYo6dfh0PaiOqSgdzIztJSFbQfcpSBUk16/SUUgulNq4k9A3J2DZNPB3e0MAib
IIr42SWrJKHckLURdPL/IWyTxfWp/anbsGm3essBVAs8mpKcmyT2OcgK1hu+D+XlI8JnevBfgGcY
t2RrqOZigGLQCnzhqtIkN7sGoFnOegzNJIhbtCXD2bmtzaDGHgNH8py9zG9LIe/kBhEP9z1jxhfD
hOrMqu7tM09OmJkaEAdmVdHDqwLm7FZ4oqLQMlV16ULTHjwefHGPa7JBcIq288pZSLuPYc80ojB1
e32j+DSLWI+9TbaSGWSaYlkyhSDyKN3UOo4anWoR4AKmO1Pv5OQRGrKOypfifwSkEXki1tPdlERL
P9d3K6dbx2oZshMdxHoC4jixZYLyBvlNzh/vnuyet+x9Agzvzat+xtRGgQ9Q16K5NhKsNt0D/XEi
DlrvuG6kO2AZOSo7bZqImS+2JdVl42Ads/4skBgpU3Zfwc7qaOEECLDkWVtRqVxjxaqBbcgjy2UU
RaXKF9WECLhEgx9YbGdM1S5+t2C68XOx7LiEu6Uj9i+tTKzSod7dljwqJYPEU2th2LefZrGh6gei
PdnemnvIbThH7DhvvGOO0E9dK+iUcOtH9qWRm44C5eNlIaK/bSHER6FzmuMwQVzBQumcCdEWhFj+
dJV9MBKpItkkTAkTeoXAa+pVF+mHDgws1cdPylCBLjCQDKltWxN0H/2/w/wifi313vcaYdrz+KG+
euVIJXcW4wAnssPISqyg2i08Kb4iYon+ecOCJk5BleImBMsiKWADj6V3safD2SQeB18852WOK668
t3BYUJpmUWDBre44chsl6xQ5mkXC6Rh2feIpRNtjb7tBbxwEGfTPgVwq8+mnv9UXiToJ5YvORjLO
WWkjQ3eIAoajLBg4T7QGtSX5VBRpH+YnsFmtwEnynE8BHxrtPXupk6tAfRbT21Mh8xsDWDK8K+4j
5UoEc+mBci44j1Ant4/zj0WKlPvzQpqsd+zEhnuwRniILVToOpRpnTZPHCi3Awt/jxtRN2tXl3gd
sS7Lmkhbops4X5p40oFSNxrMKr76jBjfeo3wZAGHnvXvv8w1Uu0EpAYVEOG7piQcaJu2yMg440sE
yd7+FkO0iwe5e4Jwq8gi0HQFoakAuMlnmLy+/MaXep1Raffi7iG2Fs41ZN6dE5X6UW2stEK1SrDq
2QTJSfZ8NJvIFrRT5/m87X5styU60RB/Q4NZEOF35dnaEB+1FYnA6XrhkhCI+LYJoMImiFQRhKdt
KydyithzBbVO1+rE5kFFvhoCxXV3r7jK9S0CFRpg69dH7hgEZ45U9LGEf9t3SgBzWP+WTCP90lPz
1055LmlLcyMq1lIBfGhLfP89LVpJIXi4fP/FbHq0N9isJ3kRbGK/TbtSxqK71ykvsPbKLeMMVJyQ
awiB++xf012AC+XuGCzgHVzVRpt3oyF1aFADd34zD2q2TINCs4BF7U2ojwRj3fAagLB9DrTuZrqG
5LpaR7It+Z8Hp1gdGdUDtZj03Sb7aIEun2zj/eiWxNBIKxEMBJuzwuhUr91nT0b+tx8UBK9FzJch
hueMHJ8BHePxhugrDHHwjEY21/Mg2O5AHfRw8vOXd+CQQdxpRlq0+Tcd72ifLyCG5oGyWm3NNQOs
cWBOpFUHBgyIi+qymSwBOu8I39y++yTXXCoev5VliAuyLPbJevgHkumQoCAnEwgslqrceOdVdDIH
BlPOwDn9pbl4BTO92ht0vV35ETaNfb6bZrgIbSSnEk1GXN+JtSLZhJYnYS8qbP3p5Hq9lvNJcsQd
syAQpyJ3pozz8t8mZnxt9mQPg9TUNEKk5NhuhYxfpwTHHwYRgv+Vvt5tVxee23TQcmw7svVx3ppt
Nm14bD2Ox6BYWwvLeYnIFxIUnoKQZir6S2h7u1YvrfUX1Cij0G2ZJU+opgWIiEHZtRwWrHS2Sxvv
9gr900RHZTWsc8o5FLBbUKXrEO02DfSs1brRvmTDrYwqNLjQm3+40S3ZOni4s0Z1jpoOPojdVu8U
jTaDWm2b7a/577H5nq4CY/rY9kBmcNmRm1ygxpFMz6rlMftb/ua+uNeKLDdxcAKAGswPigO/evwH
GxL6dG64CsVAWp0FLDxGmie6wW7ZeFsjMLcNVipKw4kv2P5h/Pa0Ume1MwemU2emQTHyvEYQyCU5
+Z7GBvwO6zwsb3bzyKpYoM/rBrXyBYcGbkEnHRmqZNyYjJRsRXO+f+iYhaK69bkpnQToIdQ9oLvX
vyQjunQdiopMbw4w0tbG5pTXQfrCZrspgA3sPVorG20y42iTYX2cUB2HySvMFfY6SoF3RCBJpSd/
5KswAtSOjUV2LMzQBtyqnW8+K6MhnqtQUhhuRcK8BnEXxamHtW3Fk1BCPotocR15hUjgtLh31NDh
FbobY3MKQw7Ahhyuuvsxl0cXvwawQZh1sRXMsoRi47V9AXyc5JDOcJ4IgkrSVuBFEvhAIHFkZhqq
X5989o5Lcgwcx6H7vsv1MBLz0O3CeekL723DyAGb12FgEWCaes+WCLoa3F8kXX4JyX1BA3FR9+Tz
oefogC7qhXtPbcL6N1Sd+EkohDLBYsK4BQ+M/xW4Lef2QTrUKyUudjbcfNv0EZioh9wgp7Rh0rNc
VrVpVwNWqp058PO3NDcRsmwZ6WEjxVyeFBBy7E8PZ265BF5vFNrXtJzJJbFfVwSMMVwneFs6R1ib
ORb7GjfFf49DCZiz4SuWRbqse54oI0fjZcG4evynbF1ibkk51OJVUQT2nRZ337vPX0NEwh7Zg/Oq
QachiA8n+dEi2Va3ah5MO0xgIeV3l0flNwyutzhFEgJk1oobsNaBpoSsl+FQcvt3cyTsrWaBcRpK
TZJIabltD5AjMFpORkQVN1K42La5isZzLPW5L0S3gkD0DaX1eaNKG/vbt9UKqvlg+A40cKPLE2hI
qCrYHUulQ6fQ1gnTT3c+LxN1zKrSHwR1FRTe4R6plVC3nJ7/O2GyhFYotIlX6y20g81SHo1LJrD3
pWxkTKunz0Iz3x95BiyuTlgsvpGgTHD1h487OZI5lCMm6VXTi5EvpvdJckm7Ly7CoJl7N/GOQOhY
ahksZ7/IxcQZTl80kfF7IEgf/12FTE6GcRzsv1tihmajysXcvVKc0nvErCnBpVSMsfNZfm8jZhSi
7e0LAv+4Rg5KAdWa6r1CGVpERPUPZo2dQErCBi/009J+6P8vz0MYv2aMuNvCLpIbFyUUdXfzgkMP
rTvSarOYkKW0BqgDLR14/eTeLgU0vN2CihPdQG4FkWUL+Zx5jnrj978bkE2YfGFX5l8d9kwBBdnE
WdCUIY5729u5Mc2uM57bGc6zAqK9OTpOEroNLa5cPHCw81/vw0q4J1LNG+yE3aiekOdOuHCmmmXO
yTOq1NT96TIqFhA9jFndM0V/lH4dm3a/rIoLX+bAE5rzxOov3c6MMdTFc1b4R+gJ45n5Pxzt2SNM
uVAHFcNmiKJqzepG5Ckp9XgiQscU3A8h27vN7Tb8XEkGp24p3PfcDrceo390CTF6BX01rQ/eT59B
DqVXX5v1PHSQZr5hTMTlM/onkrWB3HFaVp9dp50MJ8roQuH5u2gs/VeMyRJbXI9OpLgLMnksj0WA
/TPOQG81w0Og7IMMBlTlMCgT3teonN0/SEMmsRRHqV/SpdD9ClDqE6cXWkoT+aPYz+IZZTqyxahV
QGFiYQsq/bB/CzNHG0ODjTBZxUykwJ3S/pVvknhdllCriOH+aF7QR4LzcHPlAXwSyMdcS0nB9l14
FqWWv8NtjvZp2ZyT2XjxlfOreGMQJhRlW92UblK0bWwmc0xGuvALyoK0Uj0kog45XqC4aEyJOWxx
kEK7DP9q9PJSkI4QYHvGFCooQoKQ/Bx4o+7olPHmUHcNATofe1kie3iQSt1CQTp46H5IN8DI0pvU
UWmwSymErayOaB2NOrppS+F5p2Hzkh0Jy/Zr0I28hMPGDpgfcg0Ofit1QRKACLxnwSTri+QDL175
B7sVg+/D+vKp047fhK9Ze18nif8dlrbemRzQzxZzOqwqq6ZZZ6yOg7hI8L9+eoCKe/dOH0+W843w
umHLTYvjgquuYt245QvEQ4STHeXRKNYJxTjPMUPVWsF2PIoDDZHmZEcJzwnxQlvw2a2rStEmfmH7
rch+byYbIvajBQcvxrN8mm0Wp303qdDNnCwcO8LUqXH9YpJfpz+EEQVeU7nl+5Ck/2e5s9nYuLws
YAW18QiSStUNZgx2NlDpXi3AMBSGOrKnbksCzM/kH1JbJeqzbPLVx3vIAwTbDS+QjQywizR0Ftmx
wp9fAc3cOg1KIgd2M5nBGMO3JP9TLwLRQQn5UMbMXSvdZYx19Rkk/2WVC3r120PdM2fuhF+xq3dJ
xNtzPmZsDrr7QHCilQFi4Vvf7dUinHR9SoVBEGK2nBPZzX0PVLxdxUsxy09yPDKcstywpwB5L0fY
khsY3DxX88XD7OPTQjmge/6IXdRm62wPQrnCt/szXou2hxnK+2ml94mK4kckpESqV7f9d4xjz0Ur
Pe+j0gCrVGlB91QLZAfiR4gRhLu3ejTaqOfnsrfQVKxXUwpmZvKC1Tv5CyRjl3n5j4x12fd5Rf9Y
AG7aZH7J3+oVlQw7c2ML+zh5bwB+T0bbfg/LujzhndOKCeVGeu7EfI0wrHY5h2HVgB154j2J5Px9
/kJmI7wyPC9I7U6Wl3RHPWK8qq7Gd0MQ5TMtMjuIyzQvyrJeg7qHMWRdxYCCk+15a3WJMLhMTjIi
L/Hdgivw+2ViWD7w+Py03qVAEmmCT3Ru0sDBtcni1/ts2vnhqfYCgEhLdKwwK8WoPdhKxh9puat6
VLB+iREnEMEC0X82kHGDPfhxFnXgIykNZlSGMfVgoBUsZXNVeoe73JqqGHGIPKEgVnEE1G6FSJSk
f6nWc3RTSnTHgjmOXfAKE3PyoKz8SJQTdnsu2i8NPDN5FzSOY86L0HWt0I+WhYB5OmFvQRu7Aaoj
3dAjLN2jXzR0McHLvs+jtENSWd340PgaMUsVvzKhpOHR5LDcM+GQWwUcAO9wwtjFc1XILyHf1zWM
zoJTIxV1L1pGsKrgi9ZA9jmF+7fECD3PV8oxpjh2Ws22SCQsekJIn9tWrPvZbae6RZXuv3YiMgzb
+S52fRyg1tCfyGZBKMUjqf3QffnTgNJp9IayKTqKjT9oeRA2MFgUV/q6+gAoysLihCUFAvf7x8xB
of57LUFNEJqaDm6k1EEvOuUmGLhVu9oa1bxZCG0ARo1235d/63qT0iuOwunZdtgLVJgKkUGvHleO
KGFQDiBuyik6rqvJAdmxkfLIapWRF7P7t3cmL8EmliMYsWXUOj09nyGS9nm9WwI9QiYylMEiNgoV
YWqH6FaA3xPsN3hSrWO/39wqOLEaqUa9nKOhjWZEW+Gt5rA+5QXFGprkkS0RCunrj0gHWQKhyqFA
i6AkvntyCPqV3do+lUJGTmnHlhz6ttQZ8JdlKNJaEtn9givtQLW22P6KhEy4U48VzTTav8AlVDQM
ugZagy+tOp8E09OWtlYSX2nR4844lzTayjwJcJozc/tTrCFxluj1XxQepd1z2MrQcu7aQi43KrlW
vMHeeQeFHJdTX6CEClpPnLTHcFm1klQ4YdcWPBF4E5ZoMdzmmvbDbAGABHT1Q3ZVUEz5rhWeDpvn
9S734GXrK2LoK48gAi/L/t5tU+Dcy9/PFs/CMZtol79nKmqYqtgZP5PrS7FjkLQV+f7p5jnLLd1M
paVzSxYdI8iEKS6A3Px4jlrvr1xl27wAy/QSVSo63migtoY//+3gWsZ9Muxppqasqtw+h/qs0kkn
iHKjNzBk1xUoFX4NImdgHVSZSWZVnlrWPM9rez3tSTP986O2NL4SKXrUP4nB37Atkissi/i2mUGe
hOdZeVrd6pf/e9X1qhsUbAAfR9YNSTqefiBhPHJtoyY8xMIzwgwoWbd43CVxbUZUp59hm0ElcsbL
qEjVEiYUSduztDtC32NmJJ/h7u8rdfF6dkn3IpevuSgV4COdw4Vz/co+UvpUH5aCZJNRt17g9c1n
WFR7fBhPh12pSZ1um90UFJdt/9It6l5qTMoJjvSadI3K2MQrGweeVlbFcncVmfngx7uXpac659ne
jR/jl/gWuCPZ505+Im9MXiPaa7nJKyi0svg2N1sHnKuEzEVBJbMjU2B1gv3r/N+3S8TNVqIFJzaL
haBzbo32OuMDSSAqLcPO8oXs7bsSf1SR8765mqYi18vKPgcAOFb5WrI/454wcAhz3NVvohCG25x0
P7rP4nHj1wYkNAshSB5wBtJo+Im8rLqbg/j81E97jddrirott987egldsaMga+4oot4y3RrGm7fp
Sty1NN9HB1GwkP24Ihj28hc5zaPweTHiN8Zf0E0VGTdNSfaLl3v1kbe/z0J52YjX3rzZPq24diFa
KZo8tcW7fKYqweB+HTlDTPpj37iaaqqwW2ObBsCWAfMIIlzhBmGoboIcM0A5u7oJOrNDyo1d20Bf
eCVCYLTH5Vtf6LHzyK4+1SLtSEgUQBkrHopQaEB/y8t/gsQwDhJWp96vt3b1rQ3TaqwupAFjcM25
X0186tFWNCX9jqVu903hP7t8vA3dI3uqA/+pN3q/LKUeuDxkqOE9s3xTMF0Ywufaq1a7PGLvDbxL
NLSgJs/akDNXxWlQTg5djCUmRvs2kK8nPAs9yEd5zOw8fFjut4DGvC4pRdBbhhny7xbY6bvBHVws
TTx+o12Bv32UAHdykChYQnZksJ6fLE/htQrgM2GSewRUjdib4tZaQE9ZCpuQr8AqdNq/1F4lm3Rg
8gjDfKYby0zAE5+Xp9s7woZUMMVZMM2YB/GAyvh6HaS0KH8Ljn/XRe2cfoIcfCPbtvAcGhnbaFWy
YNpC00kre9NUvE0mJY3jJTbMaKEe7W4BoBn0kRLwpDNnxnkyHbmF0Q0nZomBMcxq78Fr7zK0LiDo
ivrUjpi4r2mrRiodQ50HObf3e4LLHrEWSH7s9tWmo+1+5ekgrKy81o5SOuNl3zRO9BtVmXLVk1UY
BfPyRgwRZWyx5C/9YxCKVUzGVlJrIG3AD1PdtIk6auj/y3Wu+4vksLWS5cga5U8KdQUhc88QIQCm
STZvMkWNJt7ExNFHZYYH+cE/XOIulIXKcQCisAYWwJevaWOE1tZLA/O6a4FsqtMo6aCw+j+X3dgv
posS8vfE7tXuKmGW2X5wf9PZRd1jQwU0iuo1SrCKARI0PUp6iyuuatZ22aw3yyLO0KUPJYt4MwYn
rgAIVl8mRy3lGhF3TumfXUa82Y0SVpvfSqg5GsDX2sV9ykowCd/yYUYwAz41AEIWBW8Q5kN/A/DU
Tn9/Xq75YTGSsIJriwtSGSoeOt1XXcHTI4aQY9UIRVKa3H0Ll9fVmawBJamlO/RHhCD7wwjJHyYW
YcM6wpXuDSf/gnuy0iHz8BQRiUfq6LjWbGh70tV+uTE2SQWyYRLwYytUoBrQjnHgpscLGb1e+Opl
RWWTOsBYhDnKwI9bbjQpVpjUqUr3tgoymmJBLcf8aQZtEtGfSoENai5dhUX0/ddzyytc/ypsGjQk
Nii8AYZNlPJtWJKRxzr8YvoUlzjTHLyJVqGY4PKbd2R1fsH8k4ePioHR6UGqzdTR7RLYvnzHEnww
E0vsDqnzI7tyJCfPn80ASgMZGsIftwMSoT4M5DqnXGsIu1yO8cQoR3x2qYigJP3MrkP99gRkQ3Fo
muPpPsGX4/LjPvnQB7BWsJPA1kGYcw0nkVmZ6QXeQFt6KICAUNUz9CoRSO678k218tqPm5UrC2Ft
bP1k5DtkIrXdRPSSa0z2+ZLjNykry9V4Lsu8ZZkFic0D0obUlAeCqZXzHgh3O/mkIEcySFMyIJ+4
gnzNx2bGXGZ4BhQmMjGdaff3xuZbOHXgj0GUyFtMhLjNgJLbhfmoJ8/fiKvFTxdOJSJNBk87xzsy
KxHW7pW0nln6+GJlHRD/K+GlaCjCZaU+4QZynO3RWk5X0yn3wccPNf3kE6S1hfzjHicAyZ0HWRLv
8ubgqIpUp40gWlZslwIVD+U/WViT2RW8OtYUfc4YDvI9Rlmk+UZNw71/iNa1dM+iP+6pvFifIcKS
iq5NB6reOW5ywDfHPIhzfQG/twFYemBmgio3c+Wiglqa+qRfYd/8Uhhu+lrN8UpZJ7CCKq8udjTZ
wuAXFwTjB5chzGNSMQgIzeFD8JnlTQQoWqWOFLykSvLFRnwEU+X728Mn1yPPsVC+aGDRy0vH9Gf3
JmgIJ6BHMX2kGZOml/dQ+GEhdVIGp7UohcJ9cONe/vvRJT6+naNBGvmW10tEaS9VjZK/3QN3uOXC
UtpQN0nMByu4oXOXWr2nZA3ZF8GkiKmGhrJn2Mdu8sMTw0nOXI0+GlJGxl0Nl+a0/2lTlEb2lcx8
R9VImYkn2pptzHaj2d1q++44s4XEaka2N7fZE4hqaV5ZB4PGTnn/x15gYsCPH9Yx/e9P/NSJ3Iv/
3fk/LahGJdmSTzLXT0JSVnUv1PHZWDCs6bypHLvOVUMD7rgB9RooIPzLTTlsgvx/yLR8G2GZw7oX
BojnB9PXMaUfGLWvWETlV/eHJJos7cStZ/rZDyd/bMdBPmFyEFrTWORDmf63rO8JVoJQ2+qBNSez
BLUASshwkXBE2FWskmhR2xArqkFRIx9HCFuedLutW41xzIbPHz6D9A5zBkOpqSrPfA3U0Dpooh/g
3lfnfWCfIQ0JvKtmhkTE02GYnHIOKKlAte/R1DcqnW5khaljJKla95z3St0LeSFNhh9lRkz8tdC6
L4Q6ukvM0vaefOGTOgZP057vawEYac29WkEU5w9avqBIHD+JrCf8X+AP4T5BL2vCBm18V8QZ37B1
TPsf76ydR1+IjoRe4Mc66fK41STxyv3FMuGF5lc6ZbwXCY2h9y/RHRMvc7uY5ESKPAfXPTx4EcJe
Lws4aBL83lDth7W/hYrFeGZx4v3sfXaeuEXTKL+n885jJUkFJdiSqbKIj8pW9D0VyXNIxbrTwa6+
uVAC+upnPfAu4wXi6Wh3qxY9eWXDL2i/B6L+4eTZDKrR97LXhsHPPywjlkWfjSEgSRFTcM8X1hEE
iYgR5Yi5hG4526IpbQUVDmH9YpOLGTKthFV/P7LYqi7VbMPz3qO5xrqi1Ai+caf4FUYttwE0Ia0M
1Q7Q4OKL7FJEcBx2IrlbZwsuYPTgm2xCJ/GvrJ0zaTbsXw3oTW/whrQyxB/zFO1jJGD0Miry0v0X
i62+YXqxyPsCnFeGVrMiaznVIVUjtDzhjsdWqj74LGnmpz8oaeqHARz4LGALA4mTmNAI6bUr+9S0
QZApNzj0C4GKus3hJ0jOSIPS9pf7iTEIEciZ7i/nUxWRAvn2sG43z5U/b9Wk0EO9YQDAUAAVvKQ3
Cb6q/GJtZxyt5azuO9OB0M0tWov13ONCpUedtVwXF2ojQAIY4auGM0puwm6U8zpfo/Fds/gss/eZ
Fw/xZP2l8Rt4253WVYDLor1+qxyN+iYY47I1EA20fAcUbBxWDzStgqOsYMmAzuGIWShv2R+QTtnG
D9OctolY1quQ9JcB3tzt45W9Cb8OmvHKr4VRugokS/DNSpvkLWMnvrb/JQV6VYYmBTp1eWI6fDXU
ZxJfpox/YKH3ttbJtA2fflraxB9NViBF1BWFxwUizt7vDa1gj5RxOEeC7wRR9MPKT3+ougViCp1h
h7F1TMkKfCJ2q97ug4Dey8B9f6Tol9JPBrcdfM7ha/LXL/oOM0sM2D3o9eFd0LZ3+07uM2Wis6w+
Bc6Jl3YLbUaV3iCcEb0wPK3B4Nn28OEyxluSlUgH6zEy3i9zSPi+PPKsLFyMrzObeut1dPm70oMu
U+0PXujpHOl8wsr6zepDoasj3xG+JSd62nnWYD1F7oWogVKhqqgbsa7G8jMAK9G6jtMoZtr81aDH
L5WAaPY9zDSxkuLZvqoCJOzCGGS+718iBS/c86oso07i+S8go2KbiySEEmIaMa3fQj3ttp+//aKn
4YsLGOPTPkHXq/qv73qIplpwHCS7Rnlbv+/UppF08sluktBOuIZ2+ViLxHDrgq9jo2jePWu88tfc
U7vinWMOJ0aNOwyqcxhxvZyi6PxbEF3lgakqJ2wIhIxm/j2K6hkVx0ZqkfnS+t2ERp9dC8CDQaxG
ImzsdRL9GoRWv+KA3869lSo+8CaUBbntyWEqcfrTxGWgmZg4d8NKTPf/bs1XdSmtDiPTjiUwE7dJ
wS5RnNlnL3/qHPh3jvCtCOg0OnWHJz3xcRAOiMFiUXMvq9EBJ62a0IM+upA9JiFQkUYAZOgCt+0V
3dWKIcThMWeoNrGcRmVE14CVAqRTvut3KFBamDe8RuRo9dEEgNWxg9N/fLz1vOvTRcyJ7dDdtTIZ
L96/7fSNysnQoPwdzKdIwUMUpT4JxqjzumwMqcWSmmf5xXxlGYEnH2IQuKVrOvreAKEWNYfcsYmP
yqMqSQLM+l5SPb4x+S/JO8DYP79rZyMHTldfNNfSCdznJYvPZdLCkTMUqSJeK+oa52MmXdBmkW+z
RG2I8ogZFaAQ3xSx+gXDzLUDIMraUc2j9c9ekcYZreF4MEG7AzuKBqTQyNjupYs5qB1YedLM8RN8
rwrLh9ddqcsX0I1qIflLZGJDU1HUUO6ed/9HSYubj9DRttrxL/gLkrO3X8qTkCKhVBGoQMaEc/Qj
jegjWNZuLoiHOek2M+VoShWdqwaGUpzyLv7M/VO+AInM5oy68B4bO3oBaFQXPg3jeHbSCMBzn7Gs
w3Low+/OLDXukwRe+haBNCkSAHp8ZUITs0IAHpFavHpBFReD80pB4m0q830gKOU4O+IPNPFM7B1s
MY1ztT2lLMWaK8ipOypty9eaDBvloTvw6WY6rPwjJslYrMfG3aA6XobYhMUQv2RDUYBSeTQj7gTr
AA6er3BlkabIidsBGwfMU79T19rQfV6iIbDnB1YXuZahA2jr0WheHBq8fPHhw8/9W79b3jF8ZYEf
Gxn4g1/18XbcPD+Hj7Elbi+VJrU95yJwNz7x1eu3fZ0VWgVqMTcPcVPkca2qDSWAyhx9Auo0vP7x
SWIgOcIZrSbOYm11cixP2Qqs/CZZkzqShW2xhx+zms1Y318aHsEmuhuV+WiMVNCNnTKAMKD7E/mt
44mcRWkWGbexnCpZKResZpw+XsB6rXgiPh/Hau+v0tRBnxVqdEvTtRk/tYxgabcNMOnxBdIFcjXW
iX50chYvUgD4Soj6KbFlz8F1O0UAaqNZZ+4aMCfdmiJleZkr7IJ6pWoOnZSTljOW0nZDYn1fBAIO
0YVugbVYs29tBT5F1wN0yywbG/9N6nck+HMZeSFojv6h4fYU5WobmzDsTfpc5P8ItPKTKpUyb0Ef
E6UjQthGqE/ooPc+9tHf6fX72gkA+e+0GUPAPlN+uOtSUhkUWwdM4E6JDkjP0beU9eiIV/igzBdl
/gsItEFWRxiLB5M8AofBIr5kMTks8jx+wNTy6Z1OzqFa06vBPT9bppcmWi19H0SWqYM/rxBoG38J
9Z1UlTab7jcnPYhT4DDw7YdpgzVUvG0bndFGvets++sh077tk4kosElQzFKBK5zEIvG4aRIhkgtn
ffmcAZIUkBpeNSOT0Bak1/g75ERyqO2eIZB/WTlicD5fxhrlLI+SwZXdWLBeEkxLRnAvfFso6tRW
I47J5UXa37P0g/jivWW5VjMxZ4sZnd/tqTLsuADdr4Vz2vUxGTHfgsF8gXuR8bY0/4Jo/d1ivIKW
KOQ843qIRFSlqdv272YsDufO6+dH1hxDiIsSbDGasOD5B6e4P+/II9j37icW69/KKV4DLb80P9Dn
MzmL6PhNBydZU5j9PRK6sQa5JMT0REZRwkkrY/Hg393GW90tsyiPX+WZiKDR7LsGwd51XL610qnR
h4M8ro9OXJHvL9JHOuvCfQa/8J0DcYzosinpYkprGRdcB+r4EVg1SHUyKvGX2y+WFDFjXdOaSHGV
Uq2Hw82ybOK9FsHM8A0o9tkbvB4OFK8DU+b2mH2Nz8+gmkv12FxnU04XfiakDqfMzOfeSVDKFboZ
3BR4TicM/+EaDXTLiMbwYHtGqwCOUTX43czBYPbGB9tN2qxyd0CMz33C51P48eHThImUN5ZBDhVm
G2yuNALPRwIlV1mDBGE4cYcaEDvN6WgN5CDrjJ6P5IH2gFqz0XMhBkBOy6KPc0EMCqsYteK4X9IL
Uf/CgnmZM3B5XIW2Q5WV0HtpIL7EvK6rgs3DYCp3xaHRkj2VXiBgPKuQlcBy85oORSjzOjEnPJxh
6n1w53EdfSjP7WQkMGIxifj3QxVR6KfIXwZciLguuMWqrkEeqVfqqtDETv7IAIYrb6m4vr5NWvIV
ZAd0k1sv48+7WUAuwEg+j49b6Xeq3nJNAFAMzcKDqAzS0G2/1+BvyetYaYYxkCmgR4mGnW25kAAI
0MLlYud+pW1FqETXqU5eegssGXFKbHFYhuNw6C6gBiR8iPY72te2a3Khguh4Ca7MrYixQ7Ouz/WF
D/TXvhe4VGwOPS7W3p9YXmN8fPDJxIUP2QO6s4vD+uqrMZK6VAvf04UYUDtaEFkJuds+3B11ok2A
kXFwZVRcM0YfNyyXMzZqJ/AIm+5a5/KxiQcoYcaMn/ki7Se1YTgGw01cVCv7Nq6uxuGmUELXSSxk
RF9xslwyYy1l1ws+c07f1+5cpucgEnwHarkaH1pt1R19po8Rys0AUZZAEPQone71NC+H8pc/sFmn
llLV3krY9HGS59NGgah7soucju8n1gMEORPqdbRAWm/qVax7yvbuKFXINn9KaQspHfkCWVeUS8cD
tHgoHbjpVOOkAxiH8fvANcXKTVzwngliz+3xio5/x4yVXR4bNxgpKJBsLk3kucxSFeR+L8bOmCAT
fCIQluVLRXo8wX8Wq3VR1FcvDGmIktaizR5G7ZrwMWjLlVaz1H7Rz9d2Y/9cKHay3UiRMPuqlZrS
MzFGb1bm7B4zK60lkhhfUS2fWXTswAbtYuCnJHPqaIhcaj/L4/AraM4KHH4OofN+xr/J3IyURX+S
fuyAjigKxkZBjVl7ZrGC8ewc46OZ7LPSZbkqK751RLRhXocykhRpnQhpvoS+SzJkGxJRyyVEL1Ne
Wfh67vVCeZ6VOsccoTEQjzPwO/Wsg1VKsQodLons9x4Xu6fJC5llmS1JUdutP/wa5mBwVzqkJbn5
0TRBNkAp2l8kLvOnkQBbFL+y3O8w1+m1kR+0hUueHmLzzOZ6V3Ib1kEjJcRgCPzXls4hRgQqdraK
rWMUkuUrS0XZB/d7v5q8YNpBZ761nkqHrNTJmW6GSvrBXfXANXOtgCGh+R4ytrvPzHfBuKYYl0eq
sFXZRVjPKyuE9uWw65vIH060c7iC6IS4nse+57tohZhHs5KfFbcKfdO1do3vu4J5TWIELhMfu837
FAojrj1UYVtcP1OemYFuMYhTI8HVK6TrVAVStGuZ04N6H5Iq1O9W2A3Qbz4NIJ6u57ZLNlYLc/OT
9MWeWAoDCKopFEAWf9g/JGgnA+oOSf9ndEQDX9o2gtW3WbHBcOaFqUz1YEq0OE7aIdwY3VqeACt1
Aogn6QsVaSIZeQ0lns7oalWQUoh0/Dxlzbr9hlOjcSEqafhIBF5+QtANJ6iRgnxyecQDFmAgLGWs
vvEBMGSIo40UxygtLJjRF30fILF7c7JdCI7BmiQQ6+UVDW9xui6nyn4xgml0xhF5Z7C0USkQsJog
DIAQHCCI/nwqiN8CNNdxGlpRV7IMB5MruJtPayJFXqfEeEkmLwa/2Yq3aQJQ1uowjdAB3xpCh4le
OOT+WpBfsyZufHbcAyRsG/RAAhYYSIxF3ZZPJuP94f0H137DDgViBJG/NFgWhp5zX6h1JkIc5dTK
sC+rfjU/yJrmELTQEoPtf6QbYh0itHORdfU6qdtCgLtI9AFLa81CIMx/AbqRmc8WSMUfftyX4JUO
0TUS858JQyIWF9ftUyAYUrVVS8MTe/Pps/E9bKr4J+vYC7+eNfel5n4msmG9zZfqLVD7NsJyj5wq
0wwKOnPkHi7YTqguPrbdAWW4MCZPvq3iRL3OPj5NMSUjC0tMUUXYygvrPmZYSbmffoOEv+QcyLRg
fnh6pVmdTLZjT6JXWVDisFuwjWzvHhN+zBJjF5FFbSdg13D5IeDFULoh6PxmqoUtG6KTvQvKub1+
FBzmyMrrPwcfMBqSOCiaG369M/YznYkdEP38H3gI4KFKKYXkJq9HQiaRBAfJhfGmb7qXBVPtGAII
EYbShtXcLVU3QGhEJM/cL3KT/vaaUt8QAJhb7c77ZvydIWueE87hpVQtWdMfPDTskj7gheS9DIFA
jVxHMzs3+PivrSGZqVAJyAI4dGiO+pmtLlHjjiwxWpxkKFtQy28y8l2cK07DZ6FVqT/RF0AJhRjU
j/4n1FESRd82ZmEF8WMaQrVCOQMGJCONShDHz2zZ0KDD0t1vXDUDV/hxIT3dR83ydg63bJvRGMbs
zsLI73UpJMfdcovtPzDv3lWkCpeTZSGJdwgsaMcxeDqMDzeB5/MzCJnyp8wOoUH+jiJRU+NA6NTr
tD4CoN0c4ea9mt5S7g021KENJEHOT3h0FqXFbU7A5QQS1tT5gsrA1G1jGlbbHWctCwR0VXcwoFQ7
alH9L15XgoI5ryUuXag943v4+LRocz5Vz/6z7n8rakcoQVrxytrelQaWI76eY2vA/unmCigQgANa
Pn18P9qDir4YrsMpqUHkw3B3WFPT3ofCkLLyweamH556ltynzqX4zhgGYQ5RYeYelgIpRIC061+d
mlZ2TnSbcQYniSnS8zr3fvhnb0DBwW0rsPVlPxiaHVaQkwoehNv1r0dlDmtDHjEIoRb+LmrIjbYQ
L8cQ6gbmvTAIpTsCp5INor7T9Y8FVYTskV8MBk2JUC+SQTFp49yk/BwUCYkOdawZExMMAzpVO8ir
Y9pYB51ArSVabvcVNe9LAQLsHBixdqr4ajuuQoaA9wUA8Bu0pMK/Ety660LlxIYN3hkRUZAiIjtW
BDIiyJf/70LStA5V49Rye/ASaad6pO5ITeAk94tUGJd+h2x4L3W5p0hSyasKP5+rbqEfRAf3G6yr
07nRc7fTl68iEXfboaK07iCk99AeB6p/GL5FDrmqiPWruVK+OTUVlrL/jfTnysUq8hBFw9nDiNpS
IdKNJR3SNJpQrTFG+0K0zo8RUx7ND11qH8qsStMKDndxssdrGJmD4NnKtSw8riU5h5sapMMxjxoZ
v+6xmOhRUhBQnS6ahtq+XBFc8Y7rLHKBz9LoP0AGZES+geW5lO5qFRys3IYd4RkzIeMfa0TQsgNI
/ixEG86+kwc/GSH6XpgAa44SE6oVWqAba1LDkdvPE7cfOk3E6hMfLn/ATW3ERvId2BVryjlzHol7
eEJI9mb9Qr93E1Vu5kIE9wOus5+QWu8bwma+3cho8ag2pL95Bwdopqt6YvhuXPSD54zA6tcQq6kE
FrOdjNbmvjb1LMPsepAe1zxop9kH32u2Pa4esNGF9tL7qe3AyrB/JisOV05SiKYUDOybTLHp+F9V
HRSYTT4ubrc67/fFddUnmRXz3jAhGYi5cQVJJ0KTvZidkPRo+WSgSO/bmSrLT0YrX+JHwJCz94e3
aCvsG3ztLaJDx8hmkqiTgwBzkc58lfNFijA6uuFPF9LFJ/8b9oHaSKy2Zj97hulyGuFPcS3UKCE9
01uk1LcvjDaQtuW/HdsvYZ9Z8tUNyL/KT66uBoQlmBBYCcm9gHDL/DiRAuCj8QJ/K+qSnURDSJcc
nZPVXyyL3zv9IJ2ykjrpj0inBnIye5QC8rlgepHEvvD2qIEljU9exOmMGmdoead4NhdL3q5b1WaN
KLtVqCkgKcFcLrF0gchZespvK/CUdDAQO2E9AIz7wX01H4NgB/WPRHDpPNyFSXipbFAdD8Gf+V34
u9CKg6Bb+cCfCZ8Ju/KItAb9IYVImL9AB5ZagU8gRAz0E2wJLYcxzTXcvhxqVyJtnBIdIiWNCQBR
HIJUu7zv9A//K2Gj68W64tK22NpbvUoFCMOCHLXNrpNPjNKN2wy8R2nak9ZctG/8DYV7srZW92oQ
jsceVx+hnoHRdb+6QIr3WOjIiKyYik+NZz3JIAPWN5oz8B2fNODSzjLcgSK+99qi52d4M964Q+AO
O+gmxFdW6yP84cX15ElsNsmW3fUlhMMHClDyunQvwlKj+SVoMD5afsaxJFXFuptvvHT6uRsVBO9a
Mtk1TQeDaxw/uCWCXlnxW/EEZNcLW8kqBILs2jJIr+IiMekIiB/vDTtegcx3LSiCmgTeSNOUfLpl
Dw2LSITZDGPaXFF0Hg3nCTYzjh2RUe1NUS1RcEXeZTBDh9/aFllzihceko3heSHtOq0tOu5UJ+JQ
x4kqxVNZTrpltXizdZTQ6Pc3cKucprWX/0uchkJAl9iA8lYxI3IXJowZCpbe0//3Xpb+txDLbXOf
d6st7DciDTVWE5BKF1w5hVxskzoZfGYsMNYrI85Mr3x712Eti5F9db46DDUX81DZxyPqH8pQbyTf
w9msnM7jwJwDRAmHbsJCIIs/4EmzmCX6ST+GkUXEIo4szFF8WDAxAC8CP6bf4WKYEwIR/PF+NsKr
XjNZlU2bKk2cLr9+iwsnSIkDuiZE99M9N4euTVIii/xjM0KvLbE6NxTFHXNM2Kw8eJKMo8qTReQg
CSJva38NEafHZPEx6ITmM0Zt4Q3LJssSdKcK7vOsCinEcm8pNMAIOlYd0+QBWBfHaQm7Z9zfc30o
0wu5PpvYriWseoITad3qpoUsGa0f+vC3izMfFh5bhgntORU6DiHnlsEE9ylC1Z9bUx60Oz/5vGB2
WIMi2IPHM4x9CVCPic+P0m96+roIzpI7pQerq+AAJw0MyUuwz45Zmbq3edsUIZXhQ+HniUsl6lr9
THjYxpIpy5f73nCW+b7eKYss1X+E9YyNAjY6Q3EHcbrdGsyduJAoynZ4auDhpNBzOeU+L5bLRrz0
j1GUcYPncj7OPN733HAObL7E9NVNjmRAz/P3szON2FpL7a/qX7DO8AkakfE2Rf5BAJuLM+hg9yXW
SQn/26fWhNgPT4yjIq21BBCqGTFCuFr1j9UCse5FPWcMOoiPzybabt6K5c5XJCgqMBV81plXhYEL
WHqNtD24F73CO9ZYVS6AcD21duTECP2tW8P0ylS7Dj/Pk+S/Y1s7WB/XeMOJYkDf72MzTzJaisCl
ZBEPOjEjHrMFV3yQorAdhJqg/2va8Fr0oKvnUJvz6RIWkU2LdieYkaIFtRnso47jWctwPHng1tk8
EH+Zrl3Re9qV95ndxvoSd7pTXN5ohy/KVpga2KC6EgiLa5ED1pRRjT3k47rmGiGGZRWSKg4U/lAs
aKWNhFQS5O5Bm83VYBuTYxQqR8QEqn6V3PtbUAZUbznXBYOVAxDHRZ8NbDpS8hE6FfH8TAsAq9kS
ME3B6kX1GijXfGbCY1Yq5DkzP4P9jcFg92/cQ6uTvwtrihCBZw/IqMac7CN61VUyuyWjgq7JqKrs
8wSOtsLY9axyQlz/l5e6i+bD3DZbOmpJEboQ8KwglAeNF6e3kvw6uVoUn+resuedvo5TBMTTP2bG
lrSpVjanC2edWSotDBt6d+H09xxu/Bg5xyHemYFc6936WPTbJXbi91JciDxvB5tNN22WgLk4IRGD
DyaDNNDD2QAd31LM3OQiQOi8co8TqwhzIZMtNIYfk+BEp1PmwFvAO+8NFcyRJb4kbk2gmAUPNuEU
mw4YNjyhrPaKykjmcY6QmqnmbtGSX9+5DmEemMw87Cwjhu0EzHGbGl1UCKSKwMfx3hlAfDew5A8d
z56HxNdRxX+IZZK3JMe0Tnj3wMmL/w5B4o0ieGQM/1FRO4qyjrTwV+GPsHSuOxeWn7Tka9L+9apH
I75xztNhWjYcw3SYCMzDhdi+DTi576/nK2u73uurOliHL9wWnE0y3ajxMRtWPk0l/ts0/BwfwLC5
mrL8KwK4rS0vP0WfGgimakSvpF/QD2h0QeWyhuK3jGmwUWgsN2n+GyoAotsGI7c3mzygjU5BMuxk
MKGYl+WUShRCJ4gKtzTfFp1TQXPe3Xth2H/nHxU66oJNYiT9UmQXBe2gOYRu8NjH97i9EdZDTMSN
n6gpZi4CCK0sKQG03HB9Ijt8U+YaCR1n8hMAhKFvQlOm2ISUQ0QJWnLE/IL7MpSndZJxUStEpros
n39R1i3u0sj2WTd6eMBZpuIUQbZNPolnsVoNIdTUDWqMmHdA07V/CCx9h0uI5e2BqcvOhFrnnZ4S
b6XFVT+jeM4OBpR1/tWBJVa25PPM9OLzguDO4f1CaxxGiZbk9X2WUNnvbh0kCeLIpujihmqu27z0
ouPcodu/jH4inswt7yog+hPpHr3aWNKGKeZhRvz/jD9rKHYj25/C1vK4LS1wHdYNYefltJ9E1Yoe
DHWJomb6/4aszFw5jgv6XDcx9Rz+p5pf0PfUTXmKVwDruoqhIWbEmIc2LzpbvTrlqnYf82ZNYFcl
wspqwnPscAUW+0VvqmqYr2ae0ywvUhpDxCoeUfVfcUNHR5/dtMC/+PNSV11OhNykfgiDiwWG9CoC
hPd8GpauK+HOiiMtqRaB6XZER2iVGd9ZeJL27JMwEHfk3XSq3FPfxiBq/WOnD7D9MAL3vnpTQwQr
Il2C+yygJK2GjxT3gfHPc2yTlHxa6okS2K0lGoBdSR1x3e9dkHed/ee4mwmFeSYcP72OVFLemibM
pmDTiJ4lGjr06TMqU8MmljotIg78U/gFxpt+4jwnnj4dJmCux6ieJ8OzG5B6ixDA8IBqk4gwmYFd
zlqANYQAfLpOHifzQ3gPpM8QXWzdM2Vvrmt89VSdB1SjN2jAXd5iKs9KSH640mzYbu7TN6nYK0Xs
SgbYKCczWZFcGGyiKipTjGKE2WJaF1v9dXzM+7FTG2LX3H3R3PkHpKpkfIRYk+Ngm9V8pbdEckv4
RTWeCTgYBWPDnLv6mRIvQq6F4EszqEvvGyIgL4uthJievJT2qlAQego6kyybgLWvU790fojLkFZ1
Sp0AOJTMmGTmJ90VzhdhcCR+tFsv0g7oeZbWlz49nsfDgaBXfsZaPDpPonogyect8kqehZlacrrj
dHEhNQCWf7LIlimI3FGJ2y0m7LXLkpdOJScgThxiQKjKe25BRgfp2EOc9P6yM8/yc/8qE0w3y0je
rqno/k3kfcBacagp4bxuFG2JwxXmtLjDkA2qYMt1i+YEbRB7bzHEoX/FuvFQBLTJKUY93uzkP3jP
HXSotB0xnn/FdTv0rt3v0lMTMIg7m/meCI7Svmr+KBg04dHZwSFQA5uqgaYT5rCXnaW5FiratUHs
vRlhUDLwFZ7JIGBKENSztey2kMVfZPiFziWfwKPiulhM4oTHIy1bAf+QNaGDdUbt/2W1B/4nBUF3
zhQSsDQIGKqjdl1KhwKjHRd3jrCbhUoIfzEvm4Xno1E8529gBfOb+adHmrnEnGf0utw4afxVHr8t
+pZCRsG+YJz4O/pBlwO0KQleJ4ybOnSHOWJ4yGsc0ec1qQObwcfU0W77LcKCBVt8bAGUR/DvDo9G
WzKL4NTFU/mT8cL29uykT4JWycyYEQ4I/nVYBTkRDC1Ak9xLv5tqn5CpqZ+RVenz4oZbbAlF9vMf
oQMAtFLtymP/QJnJbqWHVf+keRk3xnibLMuXO+FAcexmP0RiD2vCCfvtbewmFbg2/2/GBdVGQ+Yn
DAElGqflnPMsz9Z3ZXbx7YgoU7Gc+HskliT26DTKxXkCsRvJWLFYMMXSgZJAmUo8fVdLSe+egNR8
Q2L6ZofKapZaqpJ40e6DOlEetMInJ9UXFYI74wkkVYs6eXiSNQ9JdkKaHIat14E6ezBXXwxWBtDc
bceeCzomtPd3Eqp0AoAXdz3w5npAiD9LX1U2Oi4Bw4qAUfgspWI0A2ftDPHNGIl8q991Plbvelaf
Pegko0FNj7KujpI17xARKHduzQfgaZ+ffcDawHvn/Nr8I6ay7YI1UA84YrkDJXkcIKq9Yncsm/Oc
J1/DH2gkY2xJO6ppneRMD8U/Bu0Vvejr/tYMgKo1EiYB4VvfTE1s/hBV6ZNbQmX+KtmDlssTK08e
yotKPhFpWCi1TigFKBAewgimYTNgq4IWjUHU7VVsujxO689nvwolad8myGGKrfSpESS79YVfdAa/
ex3Lxrb7ifRrKf1em5kAfnHPoUmzNdOrBKkOd5oIv1ttf6UvXwCJRtNbCT0hoqCp7LnYzcoE9oDp
+SKYLZxV3h7XOqPY2Cxml01a6sAcvgOv3dxF4c+B+mA38wa3VLdmmqmlL05yUdRBiwtJ27iX4bqT
E87OkaXNN1jsGdDfgTI/9yrhbhpAqL47PpJVVEy0yHbPA/H7fdNYdgnstOWm2qZTdwJIfd6WvzCj
ylmkCiMb/m64yPDtuXJ0cBwPNdEmLZjVdMqZbJElpSTdmgyM1JqY3riF5lkfyvPx0Xz1LeT8bsy+
hlJrv33/xSmuj6/eSrfkqgXKKM0fjEslI8MAGhlWuNffv2rLOKIzsSbeNunZgvS3qMWJrbDqAvVS
8jx35NhnTpUw5yR9KmWrI2vZ1bfjaZOIYLaNeviydzN1TCGnMd/wqE6yTknXUfTzvfzujoXph5ci
F7AfTEKQWu/dlDj4wR3IpheMAh/t9R22F/or2Rbgj50DDGCl3EPGLWGia0r/+rFWu/6ho7tWCkUO
2K1rZguqiov2a9pHDLKqEBy/CssN8XELGINgKKiYR9+Bt0cwze5av1SYbp3PwM4lBV/ODulBUcIW
iOu6LTIeemEeTpgGyVZm3kh9c0UDmBA6HILvod2y6pacoX7tVCta6J2kCNFj2F417Y+fRuxyXCH9
3JHFZZUb78aZotJz+HdtbyusIM0QpdaxFoVUy/W7V4C1GVhlUvzS5uHAPhP2K0aN5HcMzupD/Iwd
136CiQxuj+1rXV6dq2fp//Vww7Vd2cngZN/jRxE03/cyXNqi/mchzneZxQ89jCkxKvmtXKMAKsGn
M54cJrOlPTBKaUywFaqM7WQR7fEJK8MNHvoXoySPfy1L88Cra48o21j2y9rALOUGQ3eV/Qw6i3VR
cpqsss9mlVOlOkBcuDgfvA88HnAnCjv2u04kFDQI7p0f68VuDUbLJcMZYBhdep0gEh6DH6PM6Vrf
XNf0ykc4mtHrGinWp/0+LZYKfUTH2QaOFPRaJUH9lxdt4iHUmFOlBnkZgvQreTQ/f/ZeJYIRBsw9
zno8xmXrO7ecFfAF1Pg6Iwc2yT2KC/LkatD9eI32R1/5UIg4DcScxOoyb3aSgObeLyjZhPo/aSXZ
pRHANgs+uRVlqfah9TvpsbEqgUucaT8ugY81yfmxe7FH9ghuIiCgCayRTg3lYKt1LAJXh5eIyXwM
3FWYdH49HX3NLNV+xlX2e9ujpyhz32orEMXJYKGtBTeLl5Oxj/zZV3er3HX0j6o4AuA4pQ+RmaMa
UQQLkw0pvLPnLrx8u7ORf2cmrnjV/SxfevcKf4DoxQU7h8nr7ATSEVanfI0uhNMcmNMERd5RcwH8
kYx9db/IRt98nmGoEWWPLeKL30ukdhp/B4nAFWouqJlup2/1m1XvtTz01luogyrrO4JCaPLnRMW1
T7gHabLkUxcVUbcDtq2OZrPXao4Xm8h+Yy3WzJOHS2AFTKiliI4uv9eq898JXslWzohS8VVp91mm
P0pTOe0j+YmmO4eLvIVjZE96uoKO9rK8WlS59FlxakVDzSwCGVZC7ISAO65XZ6d3czZmkULVBX+R
wbsHZs0lybvXP4STYhNhI0nhAGUjO+HZta/2p4Zukz0icShcH5l6cBjpU2fbd2ax6YV4fu7uBaGA
k7yqCVzIhVarOcotiEsnq1AC7Dx4VwEstymSwOOorL7bKm6uW//88DMNQopJuqaW3weF+BjrSMex
aITF5CRLwN1ZLbfmnHhPFP/DczmmCzOgn7nb16J7nQPIT+W21AZ7YEWqGzc/igwXPa2elrXFSQGx
VfxliiwnL4nEA2sL+aNszQIoXmo6g4C7mzYydIcf4y5y+hqhJmNSSolfG3A8a7KIx385tHum89jQ
Y5dfkcE5CKVA6C6+Edbxo1MswGHrjH2k+wA1mbf1SQYIEtCoofTTfHKQygG4ROzk8TI6My9/XPZB
dnwNMKDowptAduxoGCFP0XXyxR0c7HdKCSRjVW8nmHtRknvyCOStjj6XyiaEV/9pzwEmGV6iZOAX
qtDR7X5F5D+DvJfD9Kb4k+Ui7JOFKX0Kgicm7Zj0UQLpyA1UGh3XvmdyyHMTyoUhO0F7KxLsRt31
Dkp3lO0Dms6rnuLbCQhu8kv6ZpToYsznZ33N9ioIEhCDw/iLkYGoAkUi85DAQEUCf1EUBWkjwyIS
5Gld/7B3ul32j+knJZtj00V8otmPywn/ZE0RcXBYtQDIedEZD3rgFFA8gejJWYkwrM1odN7XzhiH
MCNBb7MYXskTwp9I7D3IzFUZsBr7CAoLCM4n9ELRkvx90Isvdxo+E6lytx97q5m6n1XgUN1sa8ce
y/V1cSA2dgwoRxbcmJfuGED5p+3MAtznk9nBZA5/0jQwptRxn/bHKRz8BRKIB/OqqaoaEOgjl9Ry
3RHk6c8uj0iNTV6284faxodca/NkHRoxtp1BGU+VR+4PlQYi9PgaIqDIy25hS6QCgutbEcq59bGG
Skyrh3plKtami37pEBhcD0UmqRJNwQoT6Ya/qiscXDyTa6RCiBjiYPzkUL6C4XboiajAAvhv47UT
LVssei2KD9QZnn7lrqg+l6mkftG16AZ7e2UX0Q0nf7890RnwRCL3/6WWA7dch6PHCmlaI9LFk2QK
iY6OVA2UxrhvqdkrpWmyinxB9jnCl0Cii9RARBYkQ2D2QH5sNPk2Q3TqWZGMlt03M9bZ4OOf+zph
pm3E4bD6vNjxp42A1IlHcZRx7V7nH6mZbMWQKbEvDmWhK+e6TsxYcvN+b+YYp0LUi2v7J2FkOPyp
lyY41WJj7W2+ecT1vkI6O4dug6YM2EukBXiBjudXBiCHZdDHophyGj2THc+xv6QvoMCW2i2sTjW/
VETJLKU5m4Iyoc6M/gGvcIZLkkbKrSkpsCfZP3ZGbHf01nyUTf9wjFvaVA8hyGiRAer/84BWgvTC
UviToZLZH0DAkQqgKQguPNi8kUMFO30Jbc/pVzkkB8YSfk9OsRhKODKIOZAywA+nIeFnH0mWageL
gad30f99XwwwqBmSVwKDOCMrff1I79/WHYTIAe/oiwpVY6JhzRI5N6CFcxY2I0hZzS9WxE3oNgk2
4dS6oV8RVPTvMQQ6EWfyduEV32A/gNv6PUVSa4gxZ9sK3w+uDWU28yqmm9SHYf0DkYh00dy1q8vN
lYPOY05fPKXVx2FISGEc9ZBqcZABayPM12cX5/n9wkIqZyyRyTDG0fRdYQEFd5vAWRoOUk93msxm
WISpEUH6ReK+77H+/XZzq1+aXHIhsPxayWQIHr2TfxdHMD9CgwkOgYLvggGWL9p9rVfBimRJoiuL
QL/WLe80nYkqn76s3p9g51qVX0x5D0r+ejQVld1zyl2a2dkUKU+YFm9djFwHE77f4BntpYRqIY7q
O/1yXEfYq4sq6fJfwmNt1VauE+WoeajaoA3WziqQCojrowGUgBZ0nNWyrHRQIA26Ii2GdlyV26tH
ZlZNQz2mbO9BZZaJO1+ljFrfnZFnbuZa8NM2bLDjkMSV6iv/sO/w+wgxdUJV87teoxrdTaL4P61Y
nq++xiVyxpB72J3n/M7hLa3M8IdxzGsq6u1SKvnWM/kKpAWEbBbS6YIJhpRJU5Fnk7Y6x9UWN1/R
jaWjtaxQrV6qdSxe0HTXGLKxF5M5Qj6XJLlkEpNsG5tFPS/OhpGrfwZR3wpVI+i0oPE+YtB3GE9a
XloxiFBHVtup4EDu4QevKimmh15Ap/STWE1XEtPPIhQP6mbEGv6y7krORds4puP8W27Bx+QF6/Du
1osxSlHv8/q6gjN6x/S27edD+rjM1UjGbKFcb4moBWDOW7/ol9GfXW6o4fN24IKZPqG2sCqC2K0G
9f2BwFcTpquBAbDPELeU8R8PCBErnJAc8rWVo/p/L0dyM6yjiGetKXiIyRcch5dhvPgS/foNvRoY
8gd9sGdGhFDERRe+34V3lS15JDKvMrswD8SLdyiMDtx245+ZXqMpqvFRErtk44NvmDo9vi6U8h4V
KVpGC4KhzEb4zuQ886mzNd7LYV2eJQw//LcJErNIn255nPM9rg4d2iaa/Yjmpb9sG29tzssaW4cm
B280kgWCQ7qgmeV6S6WolcAB7rZfUr/CI6L2vSp5su1VvKU7kXr/xE8urgs8RiDnX1BwrjKgvqjU
8lX3F2/2cxsu30ljZgQw2sFIcvCFgN3wXjkye0TdIxPsszIHIin+OyTUIj+ZVTJDTKJmld/r80E5
5QFPxLR266KCwxYXaSN+rs8a45YQIm+5HEejtjxn75DMqwg7Xo0PRJdfsDJtwxCDKUqimRUs/w54
YPXaqVORsbKZPUxUKjjphTzi8tC6RhxJxRN9fhu/MvR8fkMtsZQ3732mYW8KvGqoKJdZoDiZsIan
lWLbUDFxf5IjBOn80gGy/PbYYy0u1u95ArSkN7dXmkjk/7471Ps4SwIdv3K5HWtAePMiS8dcQPQz
nDxZmq+uSilpY3vXyV2roK8CTjhMCZfM6gYVCujQoHAUOgdJ8Oqt7FGVI9X0920LAlssFrL4d/yr
IUqNfpYlQBDc0/uuDGe8Gd3twWaIYJJZ+SlNZDGVawTcMmUPIuHx7+XeJ3VEjey03tuw6YC/j4X7
eiCv9PsnJsC1sryQhbO29u2WfCCgKNXnc3XWrKqV8sPQ3N+/YxhLD1Vh1hUJWvPluXEYB1Lq9bPm
elqZa9mVV6vcp+ogzd33P1eZ+tDgB4Xueaz4jYdef6EO8qVqw4R8r4IwYtUgg3pAvD9MA2fG0iU3
H1juTxnLaKyCDl0b9Yv6v5jN0+aopefUTHXKNpa3/aAC6+80uYzCz6YOBV52eJzlA++MbMK+2OwF
6Mjig8HJaqh7Emrebgul5QCkHg62hz4ZT84bswViDWpAnpwXNtt8uEjy0jxV89CvEkNIVbKnNKN3
44zQoSpO7hfuy4rNDmu0dp0nEv5SW742mHTz8W0qhTMFWYzQt2OsbMJnYCSxfiPyOqnRc03UcgjQ
Tu33Ph9+vYHdGVRjsYHqFpXuReSbqgisgWTJ1IhJw5c28KpCjdkQUDKwqf5RP51Geq4LvKfHagBv
WJqjsv4qNPZ2HOz2SODEV2XHyGf4ESngnK0RscceEwYM43BrinBJGdCEBYFWv4jdpKIQlsFxJyH5
2ZomvXaxANanpqkceqWgmhbIhY5VRmZ05MobVtlL1LP1XvdW2y1mtHwQvJ2VT2GkBwNKgwmgVvWg
QPTLv9CRcde7/P2j+GEq4nUmg+oY8hRA7lOFRz+MMCl/mVomskgEnkN087XRo1zp90et6ZZYvh4C
+JuvxF8yJL814xOUvmBAnRHdnDOKxn1/GbT3fAnrK997hT2Gk90igpeJ6pcr9xZuJnEFm/Ek4ZGx
bReWjt+HFfythOn9GoQVYdgkb/ATquptHEo/PJaAo+78Tnif4tOKyFfHr866CQCP4PjV0wAK6Gxv
XCtqpHmn0zH3gTOanJf8JTxxi12iCWWbJtZfCj+8wCB9siwy8O+jkvnNrrTUhyhAehrz+oj5zuzq
pMVUPVFTRxa8ZrsNfoONUwxPuIWTkpC4xQashGO5T9YAluyR428Ntl4Om87moxbIlWMIZBNrOHWj
64AIpVRpMGHNqMw6ric7/bd1kxsrguoZ11VBeb4UQ5neo8+FfcGjfLjDc3CK8tJmV5dNAJARfKf4
p51N/juje+ZJnuKtXQyn8bL05oOozp5OJaXx7L7h5+aetxcSK+l5jOCuOmDdCILVIkN1pZreE4ba
7A/Ka48nTa0CsfJU6BHFHDIxW8ioVf6L4/GB3qZufRcBB11J297ausENqY7MdJKFafCaz3n3WcKo
KiHPs0BGGoohnDsiqtsS/sSrrX2bDL8YXG9Xqks42xh5YAkxeSXc+dUj9d10af7KBIE2U1c7ApM7
AaKigpMWA1a9fKi7w6bKCBqA4t9sy+dm4GWwcQDIsgioPT4ENunbgOEfSHRwL/1DD9NiSt8dCjFV
Pl7k8RZ2V/cyNN1cWikMQaXY8+kxGZlF5ogKB6oJAk1n2fYkD2C8rqWBl8gzeBn3V7Bj2yfBbgYk
mYC1llI2BLgRWH8HgF6jP0GVBBHNqG7sey6EzH5nGLTMmjqQeDJn88taHfvXApSajqKnDz6HkZPb
SIBmZj+9QlGm69k5Zuaz6mIJihdyqE4qvH6VnVdTuet3ZHrh1T+gm/eWONUNulPLbK8V6i1ECF7x
6vwawPyscYlU2jCUdY2Y0uApnAZtPBSNK3p4npwgbvgyng66ukHbLupB2AXLUYPIRATYANtVTZfH
ivfCu1signTir/Xu42pAqw1bf8QckeMuH135GpdmZr12cPDy80roPo3HSh9zFWRnliuOq/RhdC5k
xFp5W7lhaukIRB9UKWCV0685LN9isMB36dOTdF23angoWKR1q9BH7xOFl0uELpakyi+KJok0X103
bg+Q+gj3h0pOx4KV9akf9HkIITl4Qlg68mBoNwyjIlbQe79pmZEbu5BFmB1m1n86zgvaGmAzax8y
qk+nbcFiFTrvn+fVol027hFpedsxiSRb8hI7vakLaf4klp50WWJCMvNj3oHLRFzFXFQwuWvP7jmU
ejMfFm9biezE/tbfXfjgL4JiZBtX96Jqe/xtdZUjOB7MKGznD3h341c0oCE1IDns0/g6EFiGq3tY
f6+HlEL5znB9Xf3wcFvIxu/u9jAFPaVZHIyV7Dav0h/eWXKsGHEmvpeAgM5J2dgQnJ0EBb6VG6gl
WhKLJGsUPWnwTKKxX3OCUfX5NnJ6xDSPYIqg9tm5LMDTHUrHHlfcBxCGZBgU4oGGDJu0uiV9W3wh
66Dt4QV9vXf2xDVkfBnzQZ5q1CdrQ0ucViBbxHR5L97lF8qDZYPomr8Ug2LEaJ7zGokxSZhALrth
L0Sp28hdJTndWI/AEAIwE/3AI4IaYkqA9jX8YJrCxfeys+dxWFnPVf0/K5uWs1oLHBcuuqnbj36R
MEqzvz1/CmdErQMWgw4WvWhxjlk2FmXUDMh3vVRehdfLIAv0ish8sNWUd+EK0O955zVFlZl1m1wT
4iHg7+Y7vp7zj+BQ0YvLOamvDBkU0vpP9rBRP7dqmCkYE5y43Uu9/CJVnaxBRmcomhVPaiRSniQd
moooUdz9CV5qqsOzXUmvvHpOcjXyd0kmS314O+KiMXox/0VOxIHCyOhQPJL5RiDMxTwwFn7iPNr7
KNIMtWEVNh6G86Hnh1oJy+0uqs28Ja9Aa+vgaosPWi/scX0hPxb/1JLNBfFfVjtFILChrM3RfL39
Gvxb9cJ1b16DN+zPPv4Tb4NzNq8DYvBGCgKD3q2ZncMoH8lwr39bmtHuUhi0t2Sw+pn6TWu9zack
5CKfNtVJN15aC80RrwR7+8jjvpnWLRtF4tqkaiptHlWaRnu7DtxqNO4pAM1oIvYXpvvHpMeeCjCi
CyVH75ZFMS5HE15dQClpqbhDTSJT4291s/3toiEdEtL4zwGthzyYIrAlSpYF/klZlXRp6CvmVVYB
voQqR3biSm3cr7pAaSWzYxtVj1V9s8aJV8H1FMoVKSL8Pjr9aJ6FvLwwzqui/85K6j3xvHFiO/bM
zWLMYh7HkNDGANydC+d8jMYTyM0FD0RZrlhTDSsnOxSpWyCcUIDxsTThnVhnqrol0GM7QN0kvAq1
2/YRcbhi8N8JCaRVjTnmnFEJf4nBofNQROmcHRcncdblrTmoMIIbHa3XTpNvw1bvGO3gtx5fWKc/
4vHVZG9mZx882FX/DVQsoonWvcH+D4o9x9f7R+dSp2SGeO1rh3C4ohDvTcyTq3WAIitgia1kCGu5
neroeBCRBNhTGEipW6o2Z7J6O+8YLi32n1peG0Nqtwck8wo1uANH1vms5jxVtyxU8dqeyWRfiFuH
2cnXOJlDN9Etf1wbxFK0yIMNfkdpbGtkaYTiez45GXU9jPffNwfy9XuYMAAdI+NduHGOklMEjd52
uSq6tGzLip29ie2l6TOnheCsywW1JHOA2Qce8olNVtkYB2alPpGMbrgErOe3EaRyj8PK6PSBhKlA
v+U3EEYppkg87tIH/Q7ru56tYwZRyOEdp7ZLN3YFn7cskUzKDNu2KJ4QYhblxY9eu0fNPLlR9Wbu
343eWXPgpqpEh6akxUOKRx6xXk9JefqM7YQzoe/ru2sL7uyZrTLi8oPSxizFspevjksu6TBXvEgd
GRrznhiUkzj14meVd1z88K90b496kosRFSJLcTFDU03arU7IvKgmF9d3GinPYlV0VkD2oS4balSd
VQlUQBU40EPOUtTUXs+W9ZidI/Of/dejWX7Aicg+MvOwVtl0At0X1X3cqOZARUO/aS+Fg/yStwXQ
J2uBjecrAkeXbvLdfb6bLdC/nNdo3cnLA58rQrL+K5Taf0pyVHUBbJpHTYCYNV57Q2UviLvghwf2
UlKDgSaB7JGn+9KybQjo13eJeSYtJ7WhKQeQBuQ7rik7+1YkyRlamXtWEONaoUi01+fd8YWNv+Qo
01KSn2cSAfMsI2hiqaRvxlSVJJTGdCcNO9wVNFL1Kgl+IPwOlSNTgNSZWZ7/z9ytJCemXY5NUeKn
46LWpA2eaBTtMYgsMRJOVtP3eMMrLl2xY2un8Ckin09pw71ZiUqze0t5NXuBINMmdLTB6vosP8Ef
KOyYjTme0M2mgrfPZd21b2RoQsln5Bt2mK5gThY+cxWzHmeNbhiuAHxO98HjjdMnE7cbNKDhlzyG
2RdYgjrk9DJUwVnKeQXeBzCUQdWa+HECb2aEhjeJnuhbP0Q88EsceviLOPOBkSfD/tHqgmbtQ7wr
TR471vQuaR72UyH0rz8qa5RcHt01y9lzVBSo2JSt69G2a/U99ZG6u6SdFPWpgNEFDfrm/ddRCpvU
N9Q0EAgQxNdAtoiC5XuSUJffM4kytOBMIko+1ngm3tQW7Hdv1NtjbkvXdPsJT0utLowcWd9xrgcy
e2rb+f6VLN9yuF5htitBA4i1joouoPApLfg+oeXFarqq6+KJzZu88NKqmGvziL7zJPbzdhV9Srop
aizmjMhurKBtz2xvya1sQOMFqeqAt0QWQ2eIvXfAhotf396Repcd4e1+/kSu/6aIrElhim7q2/R+
FaekYhcOoyA0fC+fPJyo9tMUvJ+b6IYTWcGsS8CKtNma1G38MLOQ6dASXLcfHJcj2DftJm3Sg1oD
yDkwT4/8fNVNGGJanmqD3C8QYhw7q9s7nNxjjge9WUjytOUTC2wMef8CUZORNd20LOfhNVssYElI
4I4z6Heo8NSeHVdwbQD9++hQgY/ezd5oKCMfV4DmmuLdnQqlCT5yPPQ6xhEUw0z/52IFgos+zaTR
Wo8XrKlnvLgN14M6DtxKDDJDjgaHipg3qqrM0ziAs4g+kckRQ1KUL05q78f8p8LaQlv/3L8bLnpU
GRkKIDT3hN9I6Yh7v9ji6u9CoaRchm/C+NDrNObmnI7RTLXaz7F+KHfcnzG9fO9Z/T0RiCa3+AHt
zd4pn5SHLfV4gMdNwUFBy1KHUE5b+Qu1AHiXaEJszB4iLLOmlTCces82NI1HomYOTBPvz2B8xIQq
vDpKubx0+1I+VVOuoSgu8+EqqhTECZyiIu+m9//S9S80dyJDO5ipY3Va9iErB8JtC8+JjqedoX0Z
txfBpVVlv6/+Ap8jKpyLXbrs4Xz1AaPTF5Bn0w9qGa/NG8WJejJjCX+ClfMYOpnVYulTiwQHugnI
//aEzXTurMdZ/SaIvK/fxx34lsBEFV4nGtZOrpJH2+7WPM/ifNxNkQuOqSQ84RSPGes+kjAQFqiH
yKPsDy6wmZ0zQ95stX+2t+OZnxiHkLHlRwJ8XhGx4MUC3uoU/K6Ww8mXbimUrK0G1iFUB5QdlYiV
ld8c+AV9TwYy7c5P7nhx2jYpLxmEoZgrXykqv1SfabXD3LlmO2urKL+KmbuGiH5u/VpYnCc1BHZF
sSmhnJEbA7Hu9okMS0CvyhrQi1XQIg5ueUxr4dIeWFQDdjw3EyZDjlCSgYOi5CbPZqYdhnc2ykd2
2YitIgbzQTOuDrHsHEKBqtahEwnAZJmglQ+IqJW3c90oKGHF4xvAfRqRJZPKbHvwDiYLvkGbN5kx
+SUhPN3PcG5dw2RmMOEcbWpwXw8BawM/nGEeoNbIzraHP9zWd6Fe0ByO26HLyPogLS2rWHJmYhOL
6jAUKnr9HDjQu6GM/G83AxM2UdPtLAR5hmlKwIFDsziWZs4aerwnzqR/Zb1Sr/7+vYi0BmQ/IbsV
YelLQQFsnQBIqHYicussWlnguHqxj11CkfgCsrQf/YXVujDX4LxhsatjiJJK61EpJzsZ8/TwAnz2
6ATZNR3oGjwhrFc4CJQ0meYxiRGK8C4w79//H6cQqPwfxuX7h5FSRgtli3TgfUABDECqH8k7sToM
JmK7MqgCVXWz8PjmmvEj8uCxRoJ9PXEdClmr46gkYgW/MBmp7mkYy0AjePVeiQEd5dspql6MIff1
61NHfleWnoRX3m4vy3QVbVm5fqk75wVUVRIc6Jbc3pSX/YZFGGY0qhsZYASfUM12EEqdYmKrBKxB
7+e4SbtqirG57HtqepHzZEL754eYc3qIlSSToCvw2Zd5smWLAgFZI0xpqmwkuOpPI5vSBlFnQrHa
xnvMeXYI+C32Mer2Hz/FRLXlEGKvRWJWkD3/K4UZ/eaXdNXQBoeP1R3HLFE9JDRDzgDyzHksgzxG
dSDqwYM2ezTUGHKabgcoupMqG7L1fwDioJKhmqmgd4Wa019SGPcdYLaZ/E7kmwBzS2DtzuuF9tlW
i0mdRXtCir27GCHBD46SsemTBTEBBtGPHa9RWfMiChWV95OefQ0qO0WgTK5g2t2TM42fjtrLPzGi
lU59GaaCCYeApgsDMwHb+mSQHymDizMKg/ii8+0O4YxH588CP+QAdlExpYEhzwdv0epC/1+8QO2b
LJSW41Rx9n6ox1Kfqxc+qmAgtpiEZWoplo7V+tq8RCeGjA6lKe08/japA5spi+hDBUaol7N50r26
BDnLkfqv5ZjFsU3uRg9JpOki4bcsfkvvCij3i0bGmEpYZkW/ArFqRoxtwByKb46Tl9ZRUb1/EPSL
wymFwXnI0GttaveFcfjc97FvoQ7dDkXrzQumb31gK5Rk8Wb3c26Q8sDOhAQ+E6kwULOzLhRtwq4x
6nqpYcRCHlRNb4gYxkSNOvyV2nVAeaF3a1zxpAxgufKexkH+3OMni46EJUfihagZSqL+7jU8l1oD
0prV7PtcfzFNPf3FdcHKV040kri78xw+9C1y19xaKSP54t2pas1n1HKjE3k7jeq/8VSZzNKOqmiT
GY315exxNqC89orygJMs7oqami83hj+ISsrIIY06XkaZKL65pqhvKjyXlSHRTDXkBU6O0mKHtE4S
8o4X/Sfn1oUQMzY8upEUQh7fXDh9BgTl4Lm00RFDZj47cbrgYQ1Kig/Sso8jG63hdw8fa3xMixoZ
f4QJPb/Kzrz8wAiogqyVfYPP8c3bMhqBrn/3KGE54aV5r0tXv+SIJi7nLtLjyBDIqshqa3RXWv6Q
y0fnEhm08BapY/q1u0Ni8EwEAkvBvaLBWNxG++9pPiQs1ANa9p1mX9mkfHqaZ7LduoF79QRudJsA
onP8xcVdZuq/WNpFUMjxvcwVu2NyCnU8QGfUSoEH0DjVnN00y1D06FFXyhHWfHlUBd6RczjE6PYC
W5Y1I65T4E+smC4OyrnETlMvwdh5sMHeN9Op4ljyLLyqxOusZoBo6gHyicR9/La+gFqdIzjyjExY
2CwWqjtp/LZYftTWGdrD1gPj/SEZpPKE37Hosq32OhbWxjbGFAo7QhPF+fiVqcW408OyS+gPiEiq
UIQOI21qFNLWbk/X6KNyTh1mRbBMC7SyDnt7X8Uees6O0WqTglrAlKf3e+WV8IXrm0hRy2sSBj3Y
Ce3quNZiYINyFMPEI/DXHZIsdm6d/mK64hecoTgRBcgxP1OstBhKQVPPqXJ2qo6GDo68b6dylrhf
Wbr3UO/F6NcDpY3olkfbazH7ZfPcBkpKJJ/883dmpsfPz1AiTOxgYYBu2a05EQHcMe6ys7Mg3ZOM
rF82t1ofa8be74D/4m9PLJZd3dea4tq9O33wwLSPMQ7nUWjEpaR6xPH5/ghYIweIUo4xgWi9pdVV
8jvo2xJs+2Z8uM0Z5bjtI3HHjwyxgKMcdl4Jy8/GtPQ9iOPqwGEsvlDP1aZo/Zv7K63Zp2E1cn7i
a7yxZ+/3NXWkqAjZWGdVfZ8QDjKw7AngQSP7Ck6+7643iLHRuVkR/kAOjcqbs5QkeM/YDUlLxyqv
6QXKNrHFMRpPoOyY8ddkcMB9KutMqTw4UmgMriWOfFEdtIgi2/SEX6hgG6f3/2hgCV5fAM/arMCT
HHLfx91aiF804lXhJ2WIP6OpInxxaVyPu9n2ePaEtRLdreQ9s3i8cltHA3XY9ofJpO7ks3k7g/yN
SCwO0+OZFIgXPO9fRNpwxhIoERZpgN5Uao8O4eR0IUq7ZKD/Yy7TwoGyQs2Nm0v2mAukRMvSF9AN
0RO1gRde6sndMq1RsbvXAy8a+GfnMJWeTYdDSOEE/jiAVdaXbEbXKmGYijbV5zobVrnb1xZd1hM4
8lPDWZL0BjG7+5MZ6dJ3J4uhdxDr/P5tAEmjAvmRHpu0U1JEP1SyQuuGmDpsFoeoSMkbV8nA/IWb
I7Dli1DnhEs8BC8TecPKWwlE9lvQ0HCCb/Uev5HW6QaICAdIuxxvgDn783oQogAxK9U2CtISK/y1
ZUDXCADuZFmtBJ9AjKb5I1hl0kUkGf40IX9X7sS9fpsXBjiMnFyivbNrpY9POcRsR0DYFOywEFbn
BiRWq9OpR8wu9F0GqmYevt7yCca8DCV4oAANYJQ0AiQyv+BmAv/2Z0kCd2KpyVk4YjP+mOE+8QL8
P1bo0l1e8IEY4PnjSM1BDJgXYd9gVQGiH7kVPRIuvtO//1f4I0gyQfq3ljl8eex0pCWAZaWf+uWi
1cubgCrBvg6vO0hOjWEAmiAtX+Eo84yV1Ezs8wgVZMBvaBdJ28XwjDOM3WVjYp6FItNaPptjTPiQ
isx8XKoYvZN3UMiy7AW52e8HTKkjze41McP8l6BFIsOFrxOzPqvY1KgglDlQkBItSA+CT8eeQ95X
/YQZSzVA4CtwROVrD1vEYVLnufj1+vnWsBV0Vq1ErbNnRRIaZ8ByQedoh7EiY0sXfFzOAWsPx7HT
gfME4TgezwiEYWX2iu/fQd3dxzP/tlgImFsEjsOy9oY+M/+YQAO1m/7P8R9GUhiEDhIlkre3pE2l
1DvBFSLICuiwf5sWr8U2bjpSXK6ASGBXS5UbdTUGDUtpfDetxNYbeHp6vgA2BgCIo+hEzKFBjVmp
sW7JkTxh9AvNH8+F0Mp/Qtump4pcIJeO02bz6mqax2+3m7v0ygYFzHkHdBzyP6NTi4/GAtXsDxus
qUUX0/4ZZZBWn2zQw6vZrF0QyFRnLT/qDey0V+1AU2DbpNprqaBpzYtYJdP8Woos9Mkk/DbWYWbh
rQncX/qxIyAiXJZ4oukRPesExEmM/xcRHeZ1TG9KMXm2XqBM0kJrYb58qtd+ABptp5cI+iRcnQhQ
pb8ATloGsMqcpogsLqvggnLG4nKI2yQ2jB+1Z83ww2YOxcdLsRf1p/lwUA8Oz791/DwfyheifNGS
SRL1WXAmX7a9SbZuuzlPl7zB42hZXyxHBYuK2xxBNS3kontAWAwz4u0/q958EKCDPXTY+BOCBiqe
fDyMpiXuZCMjqYced46bA8zKAERLVPqnwBHfTOw4h/XTqmj8yoB7QTLaBWen7o2ozhbA+q2rxIZz
uiwRfU/fFD5Pu6dUb/OSdk1fI5TaDl+e/4c9T31YojC2WYUu27Yrg8jbxwMKCS6SMN6w4DNpUePp
B3AzMrDZe1G5D5GB0VXikrv3PphRGZNuCmoOJrnleKmilEaSd08Egqhzv2RHyncjzQV8xJxT7Cuw
c/DFl9dtKZtnPHQZ98ywP/2TnSzbavC3l1yN0T+HY0utrP9uFc5yGI0oLBGp+D5XGXSJNhiwgk0A
ZLoUu2qXYLIWbHYiXnTPd4X3GV0YLh9voaG8QZgCPjMtLN2Li8s8uSQv5FeC+9F5/IEUONchGlVg
RoRPv/P4fBxvixdRly4FTEFdR0sxjyIJ4IxFcb6aarPXL22iwZksH993HEXXFu9vPIamyqIQ0eBA
EsJiqgysBq0+WTxntSnG1mCPANvp39ITgnLvCdKWCGeqhpaifY5EMK3qCb8OiawJLSo5sSF3JmjA
JbaYOvtDAc3NBbJDGYbjKUq+r1zoyU9rNchRaOrrvQutEriEETQL0BoWWqdNTmdO1fOArXWQxO1f
6Nc+i4puWZwCT2bV9uLqGBXPvV8Qn7ct8IC+G2fu3JarrzpQ471Qaq2WA09i5aG40es+xwJ0U4Mp
Eq8AOmgyToTqEdLLowlWkaefFtlWiL+48QrQneDw2ZNfs1chxecQ9GDrCExt6Kokbhp7hbv/en4i
MTsoowoQ0yzJwv6A5CQRyZvq9R/A8Sv9shWTHQXv5nGpcP0k8847eR+5O1D6vSOOpBieblxdppwn
85uN60PnmTLdpyM7X0i29vrmmMjM/6hDXUO912CE51pX89NgJACK7Opi9EHaDyqTqemqxRo9BFpS
s7WKgqEnh2l6ytqgONOY98hEqOOvW2hELlOY19EPjyes0F0qg4MfJZI4YqmX6lK3Ej/d5V+X7u06
W9WRQv8ggVSdFfxZX1dcRDp8fGFVYnHZheBkdTOo0ce0wO4+s804hW5uDW8f0dYc81gw7z6B3ayV
PQ4lsvfpHLZzAXruKlNzvXOBITagDakUeOFpmvBqd865NbBCkUxXYHTfVb6uuAVap9DDfOL0GJzd
16LmSINEHci7HQr0eAc59rR72E3/4J8w39hwOvzqF/A1gkUZrtRhruYML1or1E1FdC0xWpFDqeI8
D3TGktOYH+azUI0fevF93n5Bfy3tXOouR/5t162hoNk6w9qpu2LIcJ+OdeSSWjmwlI3QSi6/bAFC
/3/23mW2gMa6ooeOmPWVJh/mUeDu8DkrdIq4A8qanB5kTlDZZBNmeQ+BXaRnn0dg2zrJAGnPvj8+
1CWn5yFAv9RLloPv77oWJ1AwPN87V+4GPxKCgNebmI1DeGJmH02vMB70L4JqYzEWUtiYZcH1Rm98
vQm8ly3iHDMLkYoY8UxQtHV4/PVqO8/Y6488I6Io4O+b8M0E+RPMDU4rwyHpJ6CtbloTC/d+SbLZ
6LwyhO3oTmkIpzyV5AoONCSlG/Z/15Z9O4LLVA7ueUA50NLjva/osBRNmB/ZeWILWpVAQVNuOQQg
OfOjSPjDERA20UXhiLKOO5NIyfvk/7g8KR2vTyEoNteS+3bJ/BMmVAHNEd1NCXOQSOwiYqucyFDq
iiik9TeA2B2H6HC+pwCq5ybXLVX3Ef+jQXtu4alhIPLFjhEhYukFfmYtGCOdSkr49ic+1SaG8D0o
lwkp9MqrQbk/jKAuRNbWCac9EVOpNB66LJ6mYlYLMK+V2y++ufTnQe+msmiUbAjJBL4+jA/rQAHg
KWlVn7LortEqdTjGRm7kog41zs1ho14Qxby/mQBrbnQkSfbTrVyj3kJIvsyn6NOTvawGBunOzzdU
nn8trXVbaY1EL2nI1DLxWhoGcYNNuOeR/wSJnVniKzKN9miXb/fyrLPn7sQafrlUJv3fAn5pOMB9
c/BnFbnOwHNja8C+fpgoY3eazELC0aLcs+vK/P10xb4uGllKAMluTmOG3FhKY04prEcrqh/E0L4K
Y1KM6G/palr9UvgPOsjs4//xMD8uUSWa6kfFAcdLi/OFmzMgx9WYcKwzTaOnZHNnnuYiumkfjXnz
BagF+LYgOAgRhTXLwDOWHQXVv1gKS4xqSJpsYTj9kJwmGnbl97uDc9wnQCvXmCW3iy951TGWMiBs
LyJ8cHu+AcGvsKzf28Dyff+HP5DfrbVuPQRnQvvxuQi0b2PqdY5CJY0EngF3EFLdH6+84MyJGIu0
/DCAODTTsCDMbT0uzVakN+/GSZa5bRSUtNa7HBZii8i07ZttF6tXE7PqMliqlYbZf6OrE+W9xT/G
Eq70si2VYpn6LkruOxdOcLfvCYIqZEEdkb4DuH3V99nu+rhHk+uhfK9fmqByBLYqXF82z5JAVtfZ
pAObM0oMx4t1TaKugCFNUZRR7bBoA+Tcsc8Wu6Qda8blWKhpFl2h7D89oXJi7U3rGfMAO8Ryznui
GYI9hpoK4Q8+8pvtwv9Lmc6JOUX6Ak7DMyH2xUqtMN1gVAjDGDBTC8go96YVphAKkIqZYgXlmU4O
axo6ubNF5osZfZBBzyVosX4OlQBoSBsFnd5dyw4YT9KMbRLFZ9h92TsGm6TKEinuN0DWnMW0guZr
jQcIKNpoKEzbtpOHlzlY+zX9K/Wb25dacXBcv0YYOC8HfnIQ5upalxV9smFD9BwsPlQBFLDQCm3j
Rxvye43s0Dh283clCDoDfjuYZBJqBgjfQaLxF+hup9PtKJBetjubYk23ueruDJwJz63eDjtT8WSL
+2dtMOXQK23i7uwNjlL+bRsfUHq8mPpEK5yh9+LG9p9hda0psLKB3G1K9V+O3KMhckap8PuGNMZ4
B9jaX7zTOO8TDndtm1cg70hRxchWJlEg9X2rKYPA56ZIGEw0SVbBjecUVhS9Wt0yHQ8j5PtHuaIW
9LJZHltzQlxbo8ydjg1uoccjHkPI5ZVc1LqGruA4DWgy6fMyYBeAd9oAT/UCYYbIRlNWkg5Z4won
o+8cZ31Ss+veBzVJ+ycHplsqPxKVZU1v3lAeqPmzkxdq2v+Si2E14BvhrItOYbCUZrruaN/QKUDY
BAzhdEj9djkniWUJK1V05ZPWVWx4UCYiDtlQlhqxq9m04+457oElnbR5bFPFL8g/RGE+ahYUPr0S
2L10XMyC+NNwglRGYzkbpS7c1U0yD/dFKPYwp+de2yX/wQBSVdupAZr6BxH4cTYaFiLexS+s0+/8
kp0kAhYu931z2fx0TfDE18B+UdOSGvXP2cYEIaZLC4yNkzWAIxRqmhlkc2/4Sqgr5geD6HdqrvYL
PFRaKn4Jv51T7/wSfHIEhXCUMUFOhq2BjWAkDBB7jYmnjbr5fWsaPZIk5Lk4JuGn06wLW6jk5ZIX
O0mysBRiNCIMQmW+ZoUSsGnbGjzfmV7M6Llcgi95ab1xV0OGTBwh204O+wQmi4iVh2UAkRRABmnG
kS0E1isHtPEqk0IaRn26pAXg1pkXoLoQCqnQ2yhsdkjvsqxEun+2E1eeK0owQcM2RDn5uAl8Bg2c
/t7txiwLtVFZAHyFrUcqKZ4AFG1Gv959/sw087Iz4WHaS+WcbG7T8soq+Fc34OlZlbbGzTN6bvP9
ZlRAiQnrSbtBU1OVxGBgOh5QRoV6VFRzZpGtr2TBlz9SOUm1wgzuDbAUhG1ZE72GA8jbHu5bqzDS
+1nqqAkR2L2HhmD49S/mY4zUaRtp1cS4WI2knh7DNBUeXLNysRjSmP++YpKrmfZoF69Rh41I5tv0
HfgCBrjh/PHPcmoSYtFH1e+/e+0kO8uSmo1rar79AykRiqnIoz3Bj1lUs1C2zC6b/sWS4exGhQFf
rFdurVPcAJwgf8rsrufCmAVh3nhci+nGSMxoKvPcsL0ttYnA3NN7oZQ002KNNX8lpLDEKCroqz2f
Zq1diFOWjYK2vh1Z+fSzSYiqRdeuNR127SekJsxHzbltbAC7UC8RCm/ilVUoMKdmtgCYDJJMZoxO
sE/od4dyVj0KMMftSm7zAi4T/B65rU53DSgxCO0HIS2igO8V1VyVUi8wZBmgWiiEuc/dY9EAFQdg
qPb874ueBf+XMTo0zMiU6lEWXxDOUiHYrO+VpmsuoMl3NKgoVBzKdaDa9nTjm6VhOnBQwRwlcldn
BHnfeVpA+5MADpdb+DGAR0j68DPSZ1Eer1V4S8wa9e6QRjuvu0h8qf6zkfJ0nlL5/LUiBTrS6eQh
/WNy+DHqW4Zb4pIZ1oqVDQWtuuHAp7UjOJ2oPVbj3tubDP+GipCHcg4povTIb3YfXiVrSVOX1siY
yovJU5htsmRfOXXixD7I4ysjW1gwEiV/Wh0EVRJW6/ZDAeKzQA0CBCI0iV9KA90gw8E6Nokt4vBi
qzAFa9nvoVqjfOPJokbrDtOoT921vSsSrprri5uH5707Jw7enmI7U0xtlEjU0D4P6gbnEYmA3dxH
7a9SEpmQNV4w6sKiA/BiIFry4vtA0T3nanEyrwF6ky97vUiwMZ+VG/kHZBJQ75q9qaCcnQhJ73z/
Z7sz5gvjx31YM8A/4KoBiLYOKW6dryY6pMU5dIktDJnzPFH72MCpQsS84kxjCxZtNC4QwhYzevhn
lzOZDwlYOAgD+aFGkI9Ydy1beOlVst7Xac0P67c/z2dxZ1ncCTbbtaRt3SZQ0N0l6aS8C49bqgYj
Ei7eQnAB5bTyTbqrhCIsyFkIShBxk/cu5AT4Vct14lNngoXXgBTZisBgQdIfR605mBiEXnyOz3Xn
KEfM+4qGrnoAYga6BOLfHBPiVXCcaZg4Mgk9AtPKB0ODTCNR92lgjbzaVX1gXDLtrP/BT7XRyoyZ
pNz9mJyYI/PYR3HfgkwR8J9k5uumyiyUHn55KW8+ZACJ3qeuZ/77ShPoFof+W6qW8MF7Z0LtI9EM
F9mjQbXDuhrJVUo1bYMM86xcelH31AmVWN6xtT99VL+Bx9+AMi2o0QJCEY9oo3f1L9TpoDzcuvgJ
EkyWF9+Fk2CqCR4O+1jh6+DscKB3zgkxEa6Sdyxzbdjto0k9g/Fs23zQdbJhFr/4AOmuWJ8PdELi
xj0BgBd7376yEBSsE5vUxGOt1X8Y+PHmS1uucbtp67au6Urk/bxMmoqyyONHZk17Tjl7PiNYyrLE
OGahmlS7LD2SRkZnnV9qjy73h6a9ypAQuarpKk1P38ZDsa3px0n5hyTIq7u1tCgdf7HD15GLiCk1
pcsdh8NRHYmcQrhvodK6yE1MXIyYQknJuECQAprzyKq8I71q32sRVVL8e2psOmhmXuymff3HhIJW
Q47PpT194Gh+FFy0uO0f5KoLz/yQbA8DWh+z0U3kNqYBYCiIQJMFU71wDpdZFioQAmY7px4SmTOR
GIREYg+fFu4ozMergassW2tyOpAVB8JoX99SPsS+fuTT7kLmXiy8LEnTMRM/PIa7zNL4SuTj1Ogj
qcyQ4CGGwK+7m8SWPnFLXvSEbt9tPN5OiOlTO4WPaoX29MW+UysZLFIXLG5/cpv4tCvYho8i2lWl
Tj6V6fwyJndjJRhP6d0S3XbZAyxmmCNcMMKWh1dI3ekQ0B/7MKalCZHJb/EJWJB3o7LQeElefBYs
0bTEmXHwPM/5YQqS2EVhl04Wr3l770ZIjAQCC0ONXmZXwJlfVXwwwY68e+WY4qry3uCqwL2W4NJ9
bO6oHFaaZJVuQyzUg9Emn9KtD/B044cBfcpD90i73WKdT9/R5G31V4Q7ZgvZL3e79F//5+1CM9Z7
R/r6AdrUjjDCO2wt2G4SBGnM4XdryTmV3qM2uvn6deoiR8Rw6QRREXzIHQZouuTLhTCS1mDDCyzA
3Di3Utvv6Bkjxff0htlSrtVICsxqxBn1qtPQjlXVhzr0lS0Am+dOFmDsfYyiKfURE85XVM/YqL8D
KFn+v5ud3nae4aax7Ky4wrFppnkM4ZLN5mn2/5W6BAbNdauuOFDlGeNmaGwAN2jzZX2ExuEJTNb5
1uje76cAsQMfjT/I/1DK1l8848EwvLRtXvwW9D009DtupAOGT+Ty1ILV4Vb4kzVZEtDohIkdZMut
Sz8T0suCpnpEa8FaQGTkborWX1BPIrOLDQLVd5fjEO3MGh8D3F2p3h8ngnfhLZJqKfDdeukTtUKA
IIZkm0daKvfYlCbeRVtQv9CLY/Xbf6rZkr4v/onZNUQWaV1RaobHsOeEEYWDMuhCPWWpT4/7WMRM
jmxmOnp/S1XA4H817NKhWYI7YMweFM8HLd3Z4aSzC+ZxS/CaXxhL/mospF5OeDICAPRrn47U9F3d
baAthxyIynEnL47US7gyftDHMuVMEV72vcBOR5NBkM2JTv3RS56Bo/5zP3F8Lc7mYvGR4GMiC5k+
5+qWkRF8TNb54IeOQgwuSDPsahzCXCrjvdWt18abco9sgdcZX3/jCKo10yABR6DH6ya3fC+txNu/
SLkw0iqXprIllcTNdGpOMDqJc+jcO8uAsgCuNFsme30GFz5ilMyvwRq93HUu9hVhdUDC5DU3QIgi
gMlr3ZOgJSzh+a/kf6zL1iBIj2JbCA03IDpaAjOswa8tFU2F1B/lZflDddnJm55T0gULUxP2hmNX
f3KiYVWwt/30f14yCOFt4vWVi7+hMfwRvKLmWWIPrKZRKuD29kJDtXoIFHqW4SLU/reMjOCM5aV+
tzQoEnnfhpb7f//bj3rM4IRSFt8ALatX0wRygJtG6hnLvaNsqG6mik5x0zoCKiEKL1hEOl98HyQc
ZFcdD6Xa7JKosE7cI9k4Do8oib8g+qO2LEGvctdYLxwLDWEyiP7HcRnPsJtF7EVPmX+mD00nx2HY
vmBmEqLd7OMkkql19yztFJD0jxGwTJXMTft7OlL/mZyV4Gse9LlixB4ut36xFZEAyWnIIvK+PUwI
bYlid3OXlYKHWHlk24NbDJWaRnIyXnjemb3PUsTpcGqfL48y3eanLBJIua6mjFrLqiid/Jzbsau8
hlVuMNlWgm+U2Jyg+cnERPxrVK6deqcqEJ/ZnLs0oebdRcBRwGS9fxdgxOe3y8Ohm5Lw0yvztzn7
thvkqcdYY+HDNtXJ7PNuJCXNUuucZwVID5720iO9ybkugJ3Fe4KDRv7NsfNf7JhsRJGooPnwbWL3
Mo1ptjQKPRsQ5MPB2uZ8IyXcEO5CwPoGoLYOgh9tOF2cYsONz+VAtDU9IOS61iNI5xRTUAGnrvr3
AF0jufqXY7AVL2W3lzfAyCcXYyNAFo+2c+pcf/etGU3zCA3JKNoSDQqMR1VirU0vaQ8SYQ+19j37
uhjnf1TkMR2jXU7YwF2nh5ewHT+FBSez4CX7YkZhICtk413sqXJAAFrbd+hqD4FCCAum4jOna+BL
sAYUw/AOkDnU0JE3RIZXfI5ZaX2xXExDMewev3uaKdwN90cKnHkFHl7AWnAaD7EIA19py7ay0uCX
QFAPTTb7gYCysgyLKYyDPXAw9lhV0N40AQp01oSbMZAC8Or9JY9f7ABNti2gnRsopfCgXTb+KJXm
p5KYfXG3H7ak793KCQmOdPVMOkMS6DEXa2PwgkUTsBC1IjL3rWdVrsbIeR0j316upD/F2Wu+JNvv
Y1gkhEc1C17AzGHUXIgHlzn2Nnz9MKx2yauMDROFYUjm6JKrjm6mRCFTt0ITElEtPVmsen/AodDC
PF8JPJZLZXZ7QcNqGSK/Qx57fGg9OM/p+FdwZZfZxuyVWunDnsba1dTprolb6BecXGHpIYthEmR6
MkYkMPrTddVnneIJQgJR0PNwy97BLg85fxhmVfxPH7lc5TGntIFp0UvM94HhhPIqs/AUm4JB4EMI
Nqs91VpwfBkd8Oh34qfGQsfL10r4D4HF/cZsNrPD5eyz2SUrzVdwE1259uvy/chZiZ+cxyltdXnY
0i03mIHkIc9guit2lII4BAqibV1+G0DZvaKyNu4rjnuFGKZDEaBXuZCAs7AncDSx0gjvUhfwN48s
UFg7gThBpOGCr/OnEIm4Ts284XZtPUiGIbf0w0Y2fGtZkFTSs4XF9B4ZrIzQgqk5vT8LDMZlwtMH
F6us4tWW0W8Ic8y2X9wP+RQ5YXAtLnBQOmzRzjs9JxlbnH6p/LLd+rHtXMawc3OSBuDP+NGGMp2E
KN1Lo0Qh2v6ET58tyVRgBFteiSlsMNGDg8EZIzOz5jsFTxqfHfVovmyYhimuh3PQLD81GU//PJPQ
TU58LksiYSLigwaS0t4QLmL2FbagoHvzLOmtUR9y5yyU1xjLUpwI3EZjOW7gaeAGjChvklF1n2PV
RW7yUqLnAMq5AU1EKGwRhiCLse51NmOKKTly3nkkiA8cMgY07auJEosBHDoFqFDjIMzPwfHr9G7G
3bPwBBNfHNmGwk3BRuJXu0ClXzhO+zekyn2SIew6+XWS+9V5uEvOUx+O/igWpm3Yxmp58NVgDfcd
XBRZfYNlLlDW6Wp3SXqjgYl8YxOYrjF/jqdeUnyRR0sDmOvV4vAmTjqQHx5DoEoxsrxMOzETl1SA
UcNAT8uHqIR5X52GFXzfIeP53EmXgxO2mNkeE27fmT6tvQjgm96AaRpCcy7AAKgSaDnHnPCZRAgG
s6tVafWeUx5TcvUBBqQe/yxyDXRgK4j683F1f1xtx6AoCoL2d6qhSgynFoohC4xJeu+pqkU8bgx2
c1b7JqX7vHAHW8hBnvdOLZ8syo4ruMo5FbF4sYGpBDWBrm0djh6A2sJNQLMYIauUGppOZ9BJAOoM
gFrGLjZ6jbNCvoekc3Zj5KtEq3iyhSilTTfUG2kkE9zOqhFTl6ZBWxBhxuIWfE+47aoT97XwUye8
W+foEjeViNhR+xg/GDwaPNlkAywi/J1d3QmaIRJQuo8eC0jhnCu3An/hRaREBlcIo0A9EdGQH7o0
caFRPLhv1RinICQ6WW0UP3Ghe69tcnwumoKIt49rx+zyQM1++ActGdycJBbG5DRdGI0wIvr4oWD0
yofY9/nrbtqrOaiEDHjNC9Q3AuuSK84BW1h6bfNbNqWRd2RgfwREwmL1H3FXfgOaQU1DeFZHt0b4
QnSWMUsIYSHKwA7V+C1GZkDzuSHIo1j+mR35/K6nuXGEWiUEwuEzVvogaqlufSaS/QgVBkqdNgdd
QUSfwrBT8m+s4pYqbC007X+qGH+kAuMiTLummlm4s7sZ8FDudqgYkUUiCX4hfXvU++DtwtlppX3S
1PnblENoX6sQdLX7K7/LBWCD2zeRRSTQbuzQuUwABEnWrAHmv9o0XTNM97+WuBIDf4d4h6Xcv4lA
OHGv0rSWMtDiG7QOBejpz9St6Amh24tNcRLEqQiyBFUtnReKaiPwkuuPTavQfNgc8cqmJw8q3onf
I+0yjv3E8IEjCTjUhRFhHcYJHEAYyTjacOogqRDR6mnBuws9sXARV6LYoHW38qYtX98tfvnY5p+0
oAGtAV9m/ElF3aRczj817TLAHiwn/EHyR4PA3kiLhdmwcLt/TGCRA+ZPKoxdYOzunpWTZ2INRjUW
mzy36gUJ6gTSdhLaDDVJUUpzmBls0i1c/44hXpSeFNuHjsIcLHsdX6xbCTcRkW9dXsQTk2vr2GpY
jf8hBtq0yjK8Hf7kg2YBDsk1MwaDMbuO1hXteCF4cvE4r3mN9v2egoJn8dRKwl3r79rTx3RPxxnS
NMfRHVfpGIJ+G+rCeMPSXWlXAVwt5ylSMa6J9tGsaiznU0+lyVK5jbF4u7xSfaHLZ1ahMjXtR0KY
VARMQILjmDgVU+l9oXgMsLMh4WB/XFSx2JT52mXShu6sY3J8UF7eixqawcLGWvfUJPTHeHVhqAX8
r2qH6ha2lTlhO3j70zHdfCRTNfs7AAf6M1MoN0nl6767jj5+/MfQgHnDI6l2432cEu7xn+hAMCWo
JWVXj5T4waP1W2ivhcBj0AzK0nOb97FZ5XYdw24bS7VrtXUjJdwQFkDE3JHmxK2t4tZDkyr2oc+B
uO8/rz8zHoxKchNQQW6PsTGEoa/ksg1BoR4lIT8Itqwgo4/TPfMuyIAaqZ61HVsqwn1NPjj0/Led
PpGTZTxhmlo61l7fOMbeOr/GdwEIpeWuXC0yVMBB9pMWBaRl1omNSAgKhuIqUzIpAaDBoq0etzPB
M31VVjDhPqE95aZjXdRYghPgvl6gX8cBY40fZyTaCgF3zx/EWCX3yZOSwWaB9BstziJJHbID0ZDw
DnDe/NJQwUrJddh2JjjGQ9c+tgohXM0Tjez/Qx8wwHoJSpsv3RKmX2BC1B4jon92fkwFXaH3pHi5
loVqSW9g10VW0JhOARS0c3TJcezaRR/BVlzFCJSCSn5ktcTFrxiSqKV6HGUL0wr4e6/CdYftJSQD
Kvq9bHhuQufA+Gb2/U29bLh8NJZokEvHJf9Wrb6lDV0o3Uu86jl+/fgUYrkDl6pwel/WuYuYWOSQ
zFkrTEKl9VX5KMgRgyJQuxK4ULZs8lh7iqNdFfShIxv2TSrXzUEiQKJgdTQFQqe8uPcw0kAL6fik
/Ts9QKw7tUno2WQnx47RuFrJ5l2mIQVrUCiNxIt8/TDGf64EwyRJj6RCtxso0qWULb05ho3T+xls
w3GsPFEkLGHaAmpadhcVSLrrl9YG0Gf+stFjWoOuzfKhXlGIJDCQHhrTnhcReFzslirbmVU3LMTx
aDOntFopJlWpd/RqSv/OkfoyzSDwQGUdEtKSalCEJWya1J14vjcvtVI9dA7QIH6Xm7+bOBZF/ZBl
x3vsez5GnIaq6Y2jk5ojQknYU1BSY9eyr6yWG2+MoSax2xvtKuLL2RHL/B6Z59MYunEzxsacVxgZ
y8YlXW6pvT8G15Z8rxSvWm/AGiWgPzyPoepGJmJE4fqN7cv2iV+iPbNJb7UtSaYVydB7Fpedmzta
x6CDLhADDoArajefGoI+qeRHGOlkj5XIiK9Ke7s+FvoeK6GNXYFXPT/AIFLTsLjus0YsW0ElGHsQ
dCk/qzWDmLsJY6kz3fimEk4aWgGkNtcJykfddDHvZu5F/u0Iy5QxIeF8OQ5HLGYtbVq9YZJmsjPq
YNb8J9G7+sVZ4ZWGhiLL0trW39bYjGn0CwyoUldoSpAYH1F7qnJJS+WKLo46B23pwX5eHHppcTR/
8XUpGbS+R2a3C6f1QTdcteScMETqfEJxuVIn1aujvseGNU6i4lmQFG9H+3xxaOFFFtdh8ByAW38S
H/iCQhz/9fUkT9LpG9or7hUkOm6+vzhp5zIDo0gYZzng8Oz+kezmz34LhIYtaVI25MQ8gw5lh8VF
yIGuP3JVdVRRSqZQSD8MHXsdgFAmQVYOjLrAylKpk3N9+qMZaNqEsvTpnFJRFJ5DFs7vLadBIv/q
MxNeswTzU3kaI41jNBvMJFd7PyJjKpwXr7PJuS7G4MUzE/tPrsuduxTN2V0qk7nIMt45/nsVNpUL
Q7A1Mdbb3qBjtIQXMec056Ower2bcL4NV563GN72rOqASiJvsUz9R7q62XT+h7xUzKxZ3rQM/XGg
Pa+Yv7ov4eC/Z6fRiAXVxcaTE6TtTOVtcOWZjqkc6U2xkHzvhEB0XOuTZwBMPZDLZU1HkgWyN0ZS
x/ZT9HyTZ2K33uiRQoFfdGWSHPKKz2MWxZeTRpruO37DoS1aOgkSJI+KxBECjwgarNwWsvJff/7l
E7RdcQY2IN8Nz+pcNnjzPWkGHm4ywk1ZMv4hy1i+coO4Pn6QwkmPaZ0MITo4wQqdjKxZmYhp3rxH
NdlzlymLkj8Nl2AMdhjDbt4UVWne4G7ErLVIBI/72+82Ta3f6kI1jjpCI0Gzo92S3GIKTigGmJXa
P2NO9oISqUzPa6tflpZU9fx9XlVGzmJGSYUlvBu6CSja2I4uTVj8LXUzfkX9Yra1Z/KSA/qxfnJn
ChbMArRfk0Cna1OB9eMNv9oULPh/nQxTXGyi64q3fAPowsVFumHXZTswgv/f9S7GSMZB8D/F7Zbj
J9sidVn3SsP0JDvkvYdLFGaQx8X1M8i9u8+4kZe3j2ziSS4cfj1aPsdPyf2wtPqPK2NWai2WIMcL
Uw+uho2L3z6+XARsnWHNKccJJ5m910+33NKPK4LB+nrG3VJ7D1s2jtiwkh2p99lf/cB100JlSgcE
aSubRiNI2r9bwwPvK0SKVJK6T8dqG9yTxlkRtwIs5dRzHJF7TbmlStHQvVncB6U1aJdZhYnK4vxK
f8y4uv+tfTi9vh3tq75xItcsRe3DGSrzih/mEe0hX8lJ7dyMw8K29DjhymSlSmFTj+YHn+v92j/8
c1qdH2icY2SwSgzdMVh8npwz4rKROC70FDPqStEENUNLYRZ3Kwr072mttFDGFdU0MjsSdPdX50Zn
qeF6WEytjHvsYa1EzaAo27tJhErTDFSYa5/arnQoJ843hlesmdAsXSlIFxCiEw1+iYMYXKlm0aQN
5Rv7PXDv0oJmaEwDLM7g/407liPULAL+xEQU3561IpnmQxhJdcWX0x7b+XRMsbECRuZ1XpB+SNdW
5FY2KfwOk5u0l4vkX/W96GuGU4KbN3dptXY9bUwVjGvUiZhJdM8YKU46TRlV3HkniK1TT/pqxgYa
+kCmfEn/aYDPquf7TuddpGFOaG2J70HJ1YhsfiI0FRi88T/MMonH2FZGavhVC7EoSHtoFRNAiQ/Y
QIaaesGjL1lKDYVL754kYlaLiol/xXKc3K+HnkSfdm5SDJCrq4QAjs/3p1PQloQYLsuvYXeN0EfB
IURzkRX0Pe0xOcY028K7yhcwEAaC9jTMS6NEL5Y0M8rHO4b4e2oiZf7nqMoM4BIxcvl19mniFgf6
EXD+ffdrkNixf60eVVoBTbL3WlNOEBzt604hRdfTl+dhBz+OR2TiN5wdPQv2WX+FMlNQYvByoGJ4
8LXBM0c4wedhSWm15VPwy78xrEzf+3LYueGN3TsxxTDzo4W7DMDmV8ehUPZCnkW+JfOJiv+IkgPu
/HQYUbD8szR2eoMqsPsr433Pqi4c3TUMRtYz6+pKZs1dFQSCAhrzPwHNhAL88Z/HXrj1lK1dv5oM
XtDMHOwWPnx63OtfD0aeaAqUOkpQ9KJhFd0ZlZ0/ZfjJVTEJUbW+lSKx6zrDfdzbW0izzQSw/mK/
cmqV6WOZiO7TiE9yVbWguJ1jsNkuvF+6ZOBJGw4c79/ueWtjPXnCHKQigBogF+pDr++cng9tJ6bc
ukB47taalWqG7cBAT/OWhZZOQW+KWrL4gt7Mg2r1hKPBm3EWHDqMNTZ7ef0XTAySFhkCyLYSwJV3
O5/CAwDP8mD/6aNP/5tQjP4hXV1O67glZsCpGIIPafgsNftXM7axQqUSTWYEUk0yRy+Ev+FCVNkK
LC1NqrjyH1J3yWzHvLWC2RmQSTifhNk/JjH0O0sLkZYV4ctmoSKILTForn4YyOj3zoLvIHKu+uRY
M80bXxTXiNEiIgCw/rdN30wFzKFvVXh1aFBhP6K4aNRfTllhiirC5X02EDT0zEGOwy6G/OJUV43p
xjAv9l7SGYDhnJXg0GswrpFAAp4v/0oLpziTwebYtzgRutXVshZlExeAcepl1Z3mKVU6tJMjokT4
j7M8hrSvECgRV8crb+42UY0fbPurblB86Qr2Fg6gkTvCKgvPj7hIKi0G95RxeNYjtb206uCbkHv3
380kBowQntgsapguUTQCix9zXIM1gK5ScIIjxUJAUcFNoWTaM8brb1StZL6D6sd67YCYREdgqHh7
IM151SrzqcxmBeG0Xbcd2BLZPCPB9GkRmeqJIiK0p/ruvxsSESNI/5IDjxuS9zXFqSpVAi+TXD2w
AKIfJ4LaSokWzUhhXMhDBrqfefzxNq/iqLT/eeOO0x1xFJ3s7CQ+OdF7I0sAqEp0AT8EV9nHrnm7
4vcgHP1PlOwAi2w56/SgllhqspgrF0wNBgpzqlu7PZtmTG9/cGI7RB3VNgIfLaCIPoeu6H+O+Z7q
Da0EdKCAbEVWOfSWa68gUG1U2tuQGyy5vJJ9M2oeL9fqBgOyotQgSUEmr9brz+rYCOi7LpvZ0O40
Yu51Ad/e9xRdj9RLy7xtizIIRE+mp2V7qPH/KEg15YpZiayYYADDnLZI8tKj0WTHy3bfeKuJzN2J
Lzgb1Gu7LVDbgBaIavFnQdXo/tWiSAtJ4VKSWjSkGQ3/GYisAu7+NF+H3/DRec5mf+RCBoVn5m/n
9Uf/gB3ULE6s4VmwI/ejCvjORZdmnG1LCp3oJD4PsQLEPbTyr5ZO68DCIKq4LyfvRtrFT7U0PTJ6
OPRk5m5A4HMCtvQLa3P9fepyRPP2Wfg2adGuqzDDeMiB59Tg8Hb7hILHKNdRjfq6Lpya+29J3irj
uHopt8PKOHzhsTNAQh2/4VxfY8jTLpp3BuYuFXTyja6Q6tlsTin0BsiqW3TjvJ19BE5kpJqsb4rT
77uiPWld2TVJLkoFYS/NdJG45pb8LJAgXdlZuk630cloNowBSmzmo358zHXDw/ZQ6nQc9u7xNWOc
eMmdN6TWpPw8oSKCfXdiXwF1/30oEBRjqj8pyXylmX7Y1zNu7XSPc3qnXXCURq8ZrYFiRlAvKtzr
HB0T+6VZIq4ZRn/R2tKySgAdlPw4WMhk+MYl3WgQkvihKTahXSg557UqPgcl7EOChGWgFV8Dt4i0
+HtajVMoiqv1Vpaib4k23tvkZov84c7yJK3q0CRU2//5QEgw4t0NV0oJ0+N1nKfybOV53zKvt27f
mp4ZxdfhV7YuLoLxm6s3N1Z9Jxb3HyXRx9h8ph6K1/CDP5DIUX04kqLmwOv8Be9AhKIMt6Rloxji
NuCEkRnZm3NXqmz7focyeU0nos93m9Ilxn0uDE8HhMdYDZiB4DkYfhiH19WuMLq25yca+LTjZTOm
1RQqfQnxOSDAieAqz9i+Vfl0UQb5OfFBtFMSYNwxW/3iGg+G8BAQ5cgoL/i6KcQpsMIrX1lyIea1
wCThgjmnLdZ/VkLSGfdIbHDUuG+aEx5OaRbE0+/5a9Osd/D2dq9xwSHXyDhqJCcUCq70mn4aRlb0
EJbc+8w1N42dtdAHVm91fq2i3IjIbWd77rf85nKEyASxDATRkDTSD+wTHr9i98MXL9w6Ke7Y3H7B
TB5CfRi8dNDrgK/O0uWpP/q8eXs77Jy0Le54rVUDpH9aWsAaHivoVQySlVhYqROOKf9WCj13Jbbu
S22EZeDqsnP9C0zcNISPZJJoCA0XTRFgOiD+sqvxiRxCvPlFo8VwSuE4LYkzds+jBnAQcFE0mfbC
I7XPNVNnCKx+g1+3mnv5o7cx+FXDDYYs7iDLqV7r1QcZmnZmfeRqZSAv9VOa/1GjnGcaRQZa7cxI
NW8gekTB9tU//ecrD016geN1j1jP+DbzsrznXuA0hclSrJ7dQq91qrk871UqOWfhgOgB/tUB64oB
QrCjkvsvWQtiOKgsEiI4C40hsJLPenVIcsf9vTQ+F6kgqDvXLuGcphdD6rxLFwo0xD5Al1M3vcRt
E6bVpgqSfEUCLeYzHg+8ULBTkgEX9TxWw+J3YapBqoBUqxfbEUMkjaNTP66oIsZbNdIfURJmHSSY
B9X+tIGRVRG0vIY+kmIHjqpEBcXcNJjk/jeA7n0rpiJRF0asAWWAhd7CxcDblglUS1FXholNSdLq
FKvW8OxTQxJgYGcMwTyW5ZwVY57cxxpBf0vLHAtyqkJ94KIveRghJ5jpgRHwXdoN/bNlsK0vmO9r
wWnQzT1R2jBWdgPH2mDipaXNPPtjNyTqygKCjzoATJ/eOM4dqErb4vPXd3DT8PsitK/jCEgI1SwN
EsRrQ2zLSO2ZYuBAeDD4K5V/P9XdsoJcC9SDXVtPWZ/NxqZx2tAEnPU/948200TIcuqA9ievqPl/
IkUyRQbJLaogKII/yYz+O9z0p7p9/uSSO/tTtgwRngFAGxv9jaI6Yt6/gxNW1g248ajeOCRRgY2u
8DQKn+CEYaCome0zdNWGMztllsVcOvF/FNL0z7j8eZX9Gt3DJ7/ppxG4NDcODTUR4uPdBNb/rwmg
Z8ksmdvekicwDib76kW6b+OkKej+vzCxuV29e5xJ4ooYb1zwJgDYUnk28rcneB1IOylysTRbybUo
fzE1aSA8xIOW8sWKcbYPLLnJhOQNxApJqDl3ZXXhXPtaBQ+niBKb22HeOOTdpgsmLVRuiGIvjpZK
3qjNA170hpwZqgUOudlNNofLgXHOeB05Rl0eAg4qR8pFq6utWsdKGlCKTrFCzE6/QMY4iCqUBB1C
ImFxeAqMpfJaB31WqRwmItsNwpJQcLObl1YvAz6yFdU0MG3EuwWsK8JkQf4YPzdW9hU9Jx5WOpsU
9nUadpyB+5NCB2tArYI9TVMiTrjOp1b9CZSma3aDmAId5M3m9jD2go+y8IpiqYgPVBCYQfijSAEk
0J9hoC3AERqwgDuqadAWScoNchIC0tLU7z9YzN+epjciITxjZBnsTOOWc2Mh0yMD+gRnpt50jORe
y4MmnFlgVj6pwA69sIE1+QDr0qdnbnIo0xa2N9wlPXwf1H+TR7Vvxgz9s9PV0aC9QUC6asRbA0Ms
ZxtcPm0C6J3cjxVDzWT3Ml3cFzl/HjmfCv2KHqeeTxW4Eko+GRckp+FZxh1bXVIYqeGGpbx0e6U+
Chtm0sDz5bX0XammV5JvpCXwdo62flUcAunZeTPKdOgJapmcrzvcbvu7g3qUq3ei0wcvwuMSRbSI
t7pPRahD5Yq+46ry9Vh4Uk+URNQPTz4UwRvdmFWO0a6WgbEzQZrIY4zde2u7gGUS/7J+ZYAIwwsl
4XdhiWYRQS6CFkF28GwA1BJ4buLlmX3SONnmC/rAx1vttXuRV5FEh4ignUG5IjjGliswhHPRLioo
Xu+KZg4IMipyGsqGQbfWAvh6WxRb4ZMlOqz7+yfacvDrVEvWhB0cu1rw5OQJWdwm3ypVc2ougxsi
FuD5AQKohoFgFXPcncq9aP5Rz6843pox1yxPWOARkoJItv1x6pT94eexOMVp7z8P+xzsGPswbMOq
4coHVv3EDnQkHt/uNcjTiOanqREwa22WINTF8TYhD8f4UKtKyElrgAo01qmMVuBTZwnlX8kVIW+t
Fbv6kP8yy/LIQkogYooDmcOjzsRoo04hAVIePBPmE5fDXfp5xS7r/+uFr1c7yhYGo6SgIRHGl7ck
B58imVyqVGlEmP5Cn3fIFpjr5y9d6drBNUv3tTpVv4MQ6yN0kRkvJGnSgT4pcHq++Cbn7pSTUVsk
PChHH3ladCwEOXheOW9Ee9fUt8XjmLUPPxgfs+bV7dK5nmF9NCROjFJRUS42IWKr5H5CEi3y2X8c
BmUI7E8Zn2w57hDh1x8Lr61q0cgABMrZ0DI7d4U0ZNVTUgskTNnDsuuWwCWLel1jpWWvVnpkUVud
Y6dYnYobG4+2L7F0dP8cS6dL1CI/6Dr8+loH9n+K7KVI5BDteWG6fE7pjK+M7hURWc5AEWO/gLF1
5pHMgPPjzhKLea6Kafew2fCVXNS2102IT/L0MUZa5A2eQf8jTuYogzeKx2h69b8bATxcUxVNIkDY
jXH20HMonp2I6gx3gMf6SNZRDUai4RzHAGAP+sGIxB0iQFwZ4h0VSNp7IY0/23X0ZOdgkvMw7JuJ
wBpbHTgUBIotW0DFr7bReaUFyidhH6O5A7X2cW26Cssb2lQitfm1VCcefmiJ+KncJZMfa3BbwGpP
YI+YXx0FRpf21h9M0fbikWFw9LltOd9UCyvLr2ksNvr4lyXhJcJXM2HfpZ8O126tuYtNhBoJ7Jx9
F0bVzW3ayalhIuBPA1c61g1P+07ESEX885tthk5XB0ouTBylSjvm3bUq0ysoudstUmndfgsSBfcC
yyZNQglMSX3ewMKp8cavT8ONE45eD1So2syTj63Zv4X+EFFaGPJ3zS+vQ70kG9i4gz7fSoyIs83F
vIFi/ctFzzXV0h2+pUrDenvoToiizp0N3HsZ1TA+m/7h2tI+SJKyMO7gYGdO161fdq/QmWKZ8hVt
0+rFJtj/rMsEuyRL7jH+WOEwrkJenDg2bKs/KEkKKAUIcpWlDCfKrecjHIcPmzicMyLZNt+lO/oe
BosVGAunAnqvJD/GRG3TeSgTW1hOjuuj8Z0277/aB6i3Rmq/eXwMQuRFZ6W0c60F8Qp9t2cBcGb0
ILjcj5LZJY74AKaZGpp06eXfq7FPuplm5UOVQcspkFewZJ04PCagRb80TK9AIfIeD5dkemyPzMsP
Z8U39LIQeMb/7G+0A64YzfIVT32D/WqgEyN6Y2Y3ueVsTJ2SddlsSE0WgYnFFsI4afE9gMkTS/fg
2GcSYsqt436ta1pjdMb/z5pc665iHBZGNeBtWeC3Ojx+S7AtHgxfLknCAe2Z3WbqFsoA2sLXIH9+
wu5JR+X5ReOEBKsXI9rD91I4Q8nSvzZ4Y27Rx+rVvXWwv91BHRViX6SoMeSWc0AQa1ggTcqd+0Qp
x5zSqCm7CiruWCn+xpSUM500W3nA7YKIHy1Fgu2x4wv0SkliYJhJfKG+VpdieLoNX6Su9Tvy9N4r
PqPulOU11AXmEiWLkJJav6RjcxXjWwQXchFzX0ujAkQOb3F9H/mzrNz69qnX5VCdMZHy83sIdYDf
nNEG9BAO9jKBpLWiaA+CCB6tSgWHyRQdl4f+X8LLr/cEprf8Om5G+VlyXbZTMJiDz7/IFODt9sTX
Lshw/JqCI2Lp3hdZc26WQhBSuC99Wki4A91eUOPZlCAMk/6R2FzsOP+2K1/ZDmsnXadXZ+79dM8k
m/jr3Fw91ht+r/gO0Y6MlUNPxnq74oO2sGPLWARbSaOoriXSGxlvTcs3ulZVKQhRkzjwIhNBJ6c+
019TLSpUv5oOleRtWbF25jlLU6AMxXQRJ4EEWTh1Jt/9xB4S2XTZKlzxQhSbxAxru3pRMPcbGQjM
JibaI4la5tXAZuweHamDf7sHPJHLmUrThUoHJ7uOGy5rzZeEPgS6117ErQhBChoJpMPSbt/k0JAV
/2NaSgpYL/178SCYFPGxTp/W5Oj5RJfWYDCZnscOxmo6VF71c5Y4bNrhczWgn2h/O1JhaeQnYCdr
Vf/rSduYWa94OVZ31vtKgE+JI48MkkRg/YeIQxTBejvQHzJSEDHfZcikSIml8P1Ksn2HDS3Mx1r2
QWzzKsJExmLmU/DEwWe3BAmJ6D4TUZ186x16B4u4j178sINfYYE9rluO2nVpNQMh0j0uHODdJPz2
rg+nrswrVhZWuh0s4ZzqDm3RZ2uD6RzHBvq6aU0yTZYyHez30ces51TGZLLuba+DxWEqlKtaHDv4
WJkyCeXfuBA9NRH4IqqZWgfuzLKduwMHycRPaH/N9zvlemBsoKonDJJPH2AFotB4lxaLDUm2RYjZ
EcOlDF/crSYAvYZZOI7VZ4oAYoQ1y7mg44WLtQYZ/cU1LeyKqHeEiEdmmT6pYuRQh1FJkUmtWhEC
uD3v+5KudmtS034+bYsFxzNnbScYf8303jiph56rwWNp2S4NmbgEByMC2Y435nW2WMsBa37j4kGF
IqpXvkuEjxGSMwhLuyR7MyxB8PhiLvLgRIrAkUVmeCqCWF9RO+illeWQWxjD0hfaR7snuCegzfrO
Hf8onnjJ2CtZ3fWqYaROCDbx6LXYRddEHUxG2RhnSTfxH8MVihQt3J84wTmI3m4PaID9viWKk0Dr
rCsgRliIpJm1+GLQe2GR8MFj/bMqUFDqaQojBb4oZPFp5SBOC8HcI0r2QV6Z8dksv6oRuwHfzYSc
yR5tnUG0/yEWOISCMAqlGnX4ES2W/xeWshFnlWjY8GzR3WifRlbEuYdKzJCMOtzjsDUNgVJ4M+iW
xQ9ZFAtG3En3vvMK+EmhxwZ5ETNTAfA1tVYQ5Q4FWHbXShcjaMhpJbzA3ja6Bom38hFe4MIesxU8
nYDNUNq2G4QkHEtL0SkatbVo6/gFeixuhoiqEWNhSdWntNQk1QYb13w5dvl2oPOiWgEL5LQh1jlk
GpBvVnS4XWqSMsOxcCj7t78RCA0V2sLs2ppUHT6DnXIAsbOkcgOjH0oFJjLurw+wATi43u4Mw5Qa
1VDWO6tg7+RuuBsuT8MeZvLkKdSrBPT9MDh1Wt7tM+okK6Row1oUSfwKLEcGhTnUYaS2xhUzVrAl
hFRSbEaWNYFbspxEbu8it+sw+l3DGH3vLJIy/7z+My7SedzbDzknHpAUn79zDGbO86yTCMEI++mZ
esyu3pITBtzhnWPuBXznoUPmGOwWNMksVNPtosYwUtC+fxT8Zvv79wY3ask7N1CBafYW8CKANCHo
RLDUAhJc5LdsDDF87wsX6q9O7IjOqq4Jd65W4NhoSv2jRzyulv4ClQZwc3o+qC5y4gt5iqBVd/r7
v7Mhytrm7dVWEVRUe1uYq3/IseiW6wcfPSAqEKObDriS5YX68BVbRfPZg/oQ/BVKsFacftmRIuZi
I46oWAhDpCiymdqAtH9srtBUz7L8OxuBBP5hb3F4xVBC7+iI3z3txyxeZYnDxp0uTtnEdKD50h7Z
M/7EalZLX1g9gzv3SQiEnvGu+6WriO0eW8lnEuK2yo7lMgyE2IXR9dNAFfT4dhLYf4LMSJdxU0jR
sRY0H137/fKck0scxIbGJSECE9zbhQ6fimNw2Ii1kDl6iQGbuT58X7UvWqhIDORnYhksBma4k0u4
AO5r9jWOC12lolw5iCNN+ZBc3Gr/oHETz4E+JegtAD4U7itFIKM6y9M7++FGzvUaHkPYlWrWY7LT
em6MiyQ9oV6wNfx5SiIvc9qPzwNpqgpQv+TJr5WxDaeh+oGnrxCOAfyM19hrthNZ8yQAYO6LJeZJ
5Q3qvyfiUbIuS3230j1jFzzh2NruOR/pJzA7CsrsDZVmtLwLXG96vN4q20z008V4T5Bv08wF1dFT
DA5gduQPvPho3SBL6D75Wf1DhkXixvkSuW2+U4670DUX+cA2kT/WHowfSQL0syBJ/j6rw1r2WEwe
NSHtNmsI15csOgQ9WnMPlw4qk4uvwIVcXa9Gqs+JxJv5u1Qs2piOTo8UAPXQiFm9TFXo6iPxFBlJ
hV/0qfbHMZSXT+nMLvVLgsNxBRCiLUi+vdGi7x6DZWh2UlQKsVSCvgDXHlvInhqmPwpta674Tk0M
WjZePi6EOxe8WAGhaKhMTjonbepYpdnUWYyRyTkZwSpqP/Z7Ok/LpLB5JYafeAxtPo87T8rgQsyE
O7gFwiu3YEr1zcbjJNnE+lweZ6DNenuyjEkc7NMDB2xG+Hkwt+dCu+YOG53vZjYQauobRmX2FBXS
yCsnduN3aJ/oPX5NW1ScDEsQR97CVdoeM1j3W0c7vcknDTJo+0jBtwfuoE1Y+OVzCHQ6GEK+eLK/
U4SixCS4xO0Ya+m9oU/8L8WdYCvj040x2Ba+PKw3m03ZljPTvi3EPydU+KnB1fROQnSklaHX3Pec
RnO+AgE9hTvjE7d9gJs9RKbA0rY7XZxCwmiqSAQLW6xHEv7jaodWbCekwE76JQQBOf6iD4BRKDqk
kGoiLMq4WWoQrDE0y9L5Tnhrra7dB2llQJQWMefIjDjZkAxHL0Rja9HZhS19uxESpt8zbFh1EIFS
DtkVvQ1JPNklbtrG4ftNu4t6LkDhHtdtrSJN+8FMif6IwgtZa/pudmEsUw9YtpTwbnaiGjIKbn/v
NsFrv2k7H4MFXmTwlOJD+k3EZWKLNpeZoxVJH6eUCrETVJUvagQsZTaDWg/DkViXs+9EZfgebzX7
iDsboYX4S8G1KGHO1kZX8E7q3i4oW3FpPrgUx9pRoQUTcyAJXs0nFVxmUjCMtpgkrPfa+eJ4siSV
BbsJFCh1fKGJb8rnZfbvzEkIwMmAa1v8HN8jAjBXzevuE56YHGdxD/rUAcKUjVCvIXho8O3tMX1B
rvI3PDRnleWoTZZ/uVpCd4nwXuA92HzySGuJP+Dscpd83Pt+9Ns93r4a0mv4dX6DYldXjFYZk6Qh
Mw5tQjCM91q8UfSdkgGYTA5IDPPG61lO6uOPnUfhX5J51tmffyr3oZPcJUG28DYDqv/s4xXPQmk0
KMnPh3Lx1sdRl/cEeTotW5/6JaKk/y4dMJjpoPoPLwpl5/jsl6dno8IbtavY6XSP1Vw5mKkCKIMK
uqJFxGu93N/r2fqLc7aJvaYlZyyVgXHKoXA2TWmYht6463rZk92VoR3YoyABpRcuCOtb7UR4amav
xZhMsIJTXLaOviSEUM91sKmpFWKelCIzIesSJ0H3IS1dpyppqHeMX6R4jKGPJm1jRhCiLAB/zwQF
Dnr8iRZtyuMS6UGZZWnC5lmjGUUsjWoBX8xUmGj6CWDE/e2Rp8nbmAZJi8OUc6dpfXaw3Y+6a91k
FPnIu9kq8lB9VDxUthZ9AEbBQPB1UHuMPBo6xIN6qH7lsrdkmLQG0od5rpc/F56gQX0DiGoE8V5k
5w+gbQ0Y4//EqV9C2U+eB1eR22qPHe9fqrvvY+mO/GCqn1rc2xVD+S8fVwt3puFVtoWnwE9wh2tl
QMxU+eQuLK3R1D1gOuoZxdJxH5gvb2Enw1z/jxWB10WWJBRMCCr4sXcQ8Ngz5x9XYrSuhOb9vO+v
tlsf+EQQBVFvXsY49soE13VUBK+Ujp+kFHJS0L12qbnbLQFG+ERAvczMRiQSGcpvDWtIMtQnVqdr
IlIA4bN9LTqsbZEQQRSKMy8rTEW3+9mAeCrGX4GS1jp7ZupTSwvpaA314NVoClhFmPn4PV9dA4d6
jdcnZ1jvOvj+F6z6yQ2sJ46BXD7fHk0Puj6sW7dkODuACTBJwnZio0cEDjP3yfdws3k/3xZmDCZj
yp3ZTSkxvQLkPX2aD59mtTsTSff7MZAkRcwWUUkPBSb6y90Fwa/10Rf/lnYY/KfLDUONil3LEt3+
1gW4eB3LDi+dluYHPdqdPr12tcggdZo9wpx2xvdB5pRgM5U06jsvx9JXOwtYZD5lNasvpyjJSVQT
wkmte2Q3FRnOGpO8usMEWVdLj7FOPz4iz/KX3FUV2Hd8HV3ZMtpIqAsEpPlRk7FCvNHdlaXKKH/K
AsetCPjIJM1Z/TEc1X4kDQGwk3DdJ8LDXgp+lEhl8fxHyuTZYZ+UdgvW66GdcZv+JiaduRro0n6S
1bqm+zhZqs+CHTNR+lrT/hzOpZpmpHXbCCahkVyM2LbP+jXOhGsUgTojMqDR9jHJeW6UaQamnz8Y
yLIxAXpAI1gENNBKR46N9mafgCdcOYzykD36PlVWvFvKo3FfmJuaxKTZi3QcBe16CRDkEbK5Wq95
O0PYkSXw7c7pQ1cQ/QlHUxkNEZGLwBaLk7wZ1GiCgZkzsCDDR4biOj9Yjo6WKBChAEi829ox5WTz
H0oHk31NHt15xMKvYvXsQmQNYkbRjSchAYBZ3lDl4RxXlbE3plJcXIJDpZm5gZK6y6SBFWUIYuXS
ugZi57aCIj6xcuGQKMAoNMzslKOYnlUjzEYuaEK+JJ7OaA3y9BwC4SDPWN/zjHF+lLf0vmy9EfGV
EAhJ46CTj2qqxhuCHkPZOfXoMGlleDwVsXMPx6Pbr0JX1PBX6tjugEdSMlBxtvfpFmYrGgeyhgef
wcfE5Sx0eMc0IvT9gPRcPu37PLBxU2HZBf9xzgUW5AJectNPgEGbVcl6X0TFs8opyKHaaErgo5dI
/eIC/1HZRgU51a0UJbFvohzmnikJVAwxSh8mPxH+4avymgMB5RTCNvGUpN9lteK7m0KWlyfkoQUE
6o97hTCMfMtEcipyfnsCIx/c3+5t3Nz++xaxch0WHnVg9yaN/2Zb5Rzmt/Jd0vluGDX82VhkpY3M
5hH8vw2RVNhr18hx1yvwAyXd7y4MFYTns6a9u9rCWy6I6YMuEe/KIQy487XyWapA7ecIvdPD9UFG
bjGFoe/1ZVwyd/75O8gUavpG/Uu1yfxKq6XYKWuDD/XRzy5M2dPGOCZG2gTEz4Z4DUy9TaG7VDqA
JSGk2uo4ng4Xbm71+dd4ivYJ/giwvC39aCehVW2mqVBC36gdeIac1FPwPiYUtx5ihlUsRzRxaL2+
C0SBnB5bO96qv4CtLpJCK6Dzi0rVmPaA+f/7C5+TH/haG4SBAueIQoDOOW1ZjscdIf1uQoD4fgeJ
dUwLb4U1djCWgjuDkDaaSLmpj1nr9PGWa4W3nYUtlZ3gFn28vRd67Wos/dfuI1v8a4eKv3XG1aBa
PlKJYt1LC8IpM1JvXEEJlm0vZYPaylF2OS00z9QrptIVQMoKkoAGiQceVv6r3PkqZ5g21OB7nLSn
gcT1QRTtumOMmKHb+hzH/M72euSLEKzVM+ampePcDQFnrcuJA5dFtILUZH7CWTUxYWVx8t+UGCE/
/FqHwGseWL9/6aOGZOp+q6nVhmY/lwClXKIXcfEXBSpfxAYfQyH2iOgEeSHphHqtzoaYgAsE9uWx
jLh4/1PkQgzRN6NbnQJSYZHvSy4ZUFyfdL55FjxKEVIDQWYJ6LHpQRjsLnZ+eMqcZIVNqlecA2x9
Q2avBkxAOWRm3VTBtoYJIDuxsKfekAMsYgPcdgJ8iV4ASQNJhc2FW+pCplt6uYV7Go5CCRuDgxz+
JgQZ1EjqmFJvkve2LYnMOv1piln9ao7KBDyySfSL/+7ZPDGI3MzLlgxn4iYpNBLtNqdcNFMtqf8P
6OUp/Ves/l2XyjUuudAscA40xtrCWnEGUIkP7OkQGZWyHrH3JmviuSGydyaOfUOnc89QX59B2yjN
Xa1OHmeaYvUzkcyXvQPR7mDbyUqIRbvZT266mglI4g5QtoWPe8XJqWG3rHWr4liYbO7BJMl0/HQo
01J+1hzTdqlcxPzWeKLbz2nYDkrRj6M4gTNYC80HmmggqNpIFhhDGcpEsHAOHPkVcyqDXCvBq3Cn
GaNkkE2ETZPTGmXPyrgtuy/LyL0v9fYypBJBgBjjgJf1phBtCnc6fAWSXYQtg6C4vlUXlce5av32
ClFJMglbH4ztv97ag5zNLimwFN+SvvRr2f9Z49fIEP/gu4p9Axfk+6aGty3mlx2i/QyKaJokRJAA
v6T+zFUUjDNrS1kU3Z1a0CCS5sCyLyFPdzxmRvUxgA5YjZYmyxqhbbpl89yiclqOfGIPPh6W92lQ
ZZZt+tgeytg5BRhW7fkc1/7WL3N0YQjdTLnFkQo57UR/BcMX/OsLMOz8YXl4vZh5j8jeA/2D16qM
94MvzlYnCtEVnqxmeoCQKywyBwuZvps44998Qm6Nnc0Wji5veDgdzTMe0Z33XExoRR2KfkGHCfMU
6Ns5VkX/iuV67ojmJ0B0hpz+yolfYEf9WRuvrk9OJAfkXG9MazeNnIhYlzC5NkrCknjlsuPOBQK3
acukufgUsp6MT0fqrqMwROreV3q77Cx6L3OYu6iUqWxK+l88XrRkW2f/a+8SetmZUNNhIyzvhgNt
HPgGihe2n8xUwrNDqQD4D5bPoiGbEm3JkZrsxXGZhUlaYwA+2DYZsT8tm1V46b76iKVT9YM/g87u
FFPMq6TGqi/W4QQMMXmVXt1D5Tp12q/AQg+9EXoioGcXLHijNbZI6ajRoz2QNXL8FH35fH+iinio
tXYwiBKC9efT7TMlqLJ3zooRmyltR30ob+p+eUTJn74Y4Jt4O5djo1+VSOIoXAR0AaWxCYwePp07
8xjg7I548KrbiNGKoCYmiE95hlNA8RaZqYhi55YS4X1+rXtLSteHMxLtrXsIhdrO5vloE6ntgyZq
Il3q+hdbHunGV1efiq7QxkfTrW/jLgNesjPKRh5U60gdMIKxtXWFrwv4asqMMfusUJMBsxIdQ4vd
9WVYkVtQuxD/O4RUFy5cy+WpA2mSd0UlRLqsfl4mKASkfmKkAV2HUimwtoPwPmQ6dUgraNHp6mGr
owDpQAvAVOTwEHGI3hpT9MuxDIBXOtHjtRGCYxciCayfqfZi9BPpIopnIPyroK+3VRPpFCx3zb5S
5ckRzxOzxmRqlIC/SZCjU26exq4Fu+p3LBC1NFmhUmNGy6GsHwnCik1DAdmMDWMoAp62VsXAA9q9
VZEBXa67dy1zohmqcbw40nKG/wProFin7rzU8TN6LQT55jxWKzCnI9C3nfzRRyDE2kEdmfk/KtmT
IPJ+O39Sgkc/Cqd76SMIbuCfu8kG4p2RLMXOdcHmCFedhZ/1TMZu0/yo9q0GwbJHEehkyC7itYIF
hbsTNV6IIC6DqIV4iyQWjUJcPSTBa0MKZZP5UccFSn2tJjnSTq+HLZeyu/nBkj5X4yqmoy7zdJJS
zLjYGwsA/o7vYQ5MHWVym+bHXjoXNEx7wolN/i2eNpt0jNGbJfhTZz6D80mknjJLxW0isJa8aqP1
aGiPPGh76YtTY47cwtMQMohd7Xig8dqfECUPFvk8AbzTKXDhupkXLziMjAeV+sC2cciJVfTDX9cl
c3xjf+Mo3kvn1jKyaWi0hhqwofBPvIq3HKX+qNa7OfP8820ddmdW4MknzZ2Rp5ufNfox7rt3PMJu
t2qoFIDQeoJpUae9pEAp4HUWjd2PcwdNTVfVQVd7hbvqNtSMVzDGRoy+yd0N+Z9nwXTJLZ/95wAm
ozZ/A5gWTtjH0947Gw7ucX+cUQBSLjaCxnoAEFMrV58KIFTSTIoBdfrb46DqpVUNAKc94+nGJIvI
db9zw5WDjxsGboDZZ0G4BhZ8ZOIHEqoX7shX8zLgWZOsN/up469Isp1W+0B/eFQ5bcASGgH7dv4G
02+F8IoS0mBNjCv0pIgluFoseLYe78F5IefK5ulWH45OcpSYlrRr29T1acL/GrHXqZ9eSdTfKJYL
FOApozYeuGNbmh4efSnBmQXLOFG9t6DJpQ2qiQVV+WqQaybL6H/h/cEiS44M8l4qj4i/2VewUHX8
+Rk+LO8mK1C8ehSUKUhX6eIpdsz0hOuG5SCD/X6uISiSUuSgk4Ga4fDPNnV5z89KI0NfTiPqLSA3
2KStjKjkziVe7drETzB/VtjNtuBDqJ1I0Y0T27m2Qwnt4+dIEehnkiLUYEfZ7+q3UTq1MF67I2Eh
23Ya3QSVGUTZJ4jBx0js+xaKn7zagVF7JQ7Q/z3bBp0h5S8B2sVyDdiMmctL701YiaIz68Y4caFt
AyuBO+NRiiXydpdNLyKQy+xBaGMLng1EZPd775YCBqi1N5werC0tqnHKKE5QwitqKda4ODpf8h2I
seXhIBuOX+P0VtZ2RHCl1IvpefRwRH7baQNznNWIZxY9b51QSTyEIhb9HEiTpG2BqHxlSf4Ym/UH
7dqCGrLZTHb+s1diCRXgO1PEwvSVUPBnjPOooYy7Mu213AMHWDkX8DRc9RLCjHqsctIZSpw0CVev
SUM/iVQSJvhqjAMzihioDMyDmHo7IS9Ig35iXS8EdsupzI4jm7ZJfDA8tPnH45pWi7OarEAMBY2N
cfBMMh7eoctQr7OusESKPe12JaKpIl5Brta1uolYOCv/dzX7Lc+a72HE2D/MOeliGNJkShVuCzdd
V3D44UJ1ZlGrk+h0rSQswt/4iFYEekmGXjQI4MjawbUxBJsdJg3exsmbJt7knR0PhBPYW9liYqyH
bl0JpHOmrqQcjNflnbNZKEtVoVtCM14iJm/tXWVH3MlMbrYeJyxYOzCXcA6N13SDSawIMxFatfMW
9m6NjuV3ED6H5QVtBbKnhXVylDX2re55c0A4yRqT0PKoikF2spHU6PqqIpibgi7ulG7BZT5Nh/i3
UPDMtacP2gWKLvwIVo15SGqUNnNZyJp1mmUWPnMMSy85CCmTsSu29B8fKuIxs+4sjkCbLR2DdanC
ZeSVTl/bngio3D6qW9+o0rc34f6YXJeZJ33DtqAh/nviGi9WSHJtBGVPMmYCafPct+TN8ulf9hRF
mAvEhHcYiuXG+KbLTXAogtfxPD7Sn1MMC5nxAGYrk/2y71Cl/QAb1xZSsvPu9Crc4tzV4lVlA9zs
C1adHlAFBEuVstPaPbh+TUYWr6NJ9ZTKNz+X5Ffdt7zxnkPh12WWheCdTHQ7T0KhWiR0Qe7Q3ur2
RLg/nVMCxFCbvRee7zjQt6v0NSIreu9HYkpdgNt2+IA2O65dXV2QZGOViH33J8SJg3gV4qNhaCJQ
nHFfo4pijBRYChWBg/GMSD9yFXaDFk9qE8k1QqmN1Z00Sh2D7YVAEUqzm4R09MbtvbF5s5iymAZC
btMXnlZuwTE342dVUVgnrTT3iRExBXZLERloRglLbHVK3RoLTGaBnn6/2hcWgln+LouJJbkfwYSg
iAtkvmUdiZ+qFFjJX+bgi37Go5Q2XXNsBZhwHHOYSskc4D0qpIWvT3e7SbyC1VAvUxaY1ALvrZl8
J3D2hIflw7bnOySGILfLH2NPc+WhGT9unKKlN6qLTpPW9ZnsJkpShNH2QkGVZfRkj1hGlEFvRW2b
2cbo16tKo3Fj1t2P89R2qxWwxgVKsUVIbscBiA2Cm6MtcxSDvusqc5Bj09BB9DE4BDO8sIw3viPU
EbqTBP7qNWRCikNJvXVk+jdmeSMuUBPdUfMw8b/iJIQeLmdhrxV7En+qki43PyagOlWnHU9aTOWx
YGfVAFX7wYQ2Zxjunbz5jB9KQ4n5yvB1xPo5+qpARwbQn/gjSm+0AH8ab32ztRYaQDDzu4MIHIq/
DzRwRrgX+Z8Ewq3m6zs6SbAZKilQmyjt34B4H0OSUeuEefzQ6oxyJQbPxOxd7zTVQsl6vuCVYlMQ
eqp/4JVNgQmuQyib+93KBt+VcBMqNMI0IZGl9BwBzEuSLvMOg3OP3avfZC6nSzH4JsKszfaQQibG
tupu8s5P5CIAEzsnDrND7vo7rxBh1tm4m76oxaMwiIG5/wxzVq1iaVqfNzB8E1jKZhhpsX1y3LNq
LmaopipXWTJC/S35MBKkeQLvm56FLINyAOOxNGccXXRvERkJBDyWF7Cu2Sd+YGFDKydCalPFsJ2r
Bod1jre8U9vg/LndHmzLClYR3+gGgCCeVO6EiuBu7dYtPgS2+7Q6Jhopa2Vo0jrytAAr4Kja1apA
/erRsmebWcNBhKgHxXeVD4kQA+eiJlEXF32ubfYwVsoh5FMMswNHnPMgYP6c3bN098xNVoi/qqu8
8Qlxn7xLkjPSKAC0JnIIerq7d6iYAZVuAM5XIcvoTm6W85yGL/GphiXKGXbZ+XtWV5VeJ3blu5d+
m29t3It8uswKQoy3fWHpiu2MV/w+TqgR6W3OdM31/tpIObbMNHYmmRIUK9h5Z0xX+8cvj4JHwM9d
aaCsK7jC8z2kLRVS8gaqkjxH2xytQzz79YMjm0NzKwzBPWB2BO3bzZgnqh/M3R+DhhBVoXAYZ4JO
LqVOAYmvLiLosW2C0NBoM4WoaD4lK4ja+Ua7r2iQzxFT5g7Guse0aCHVySrH7ZDA3mkaDsVcQpcH
5scv4M7i3Fhs7Epk13wSF2WMOzVv74oS5P+2YaqYauAW7Pfe/XVnuGZZTazOmlIdL2KNUdnAR5NN
mVvEjBIxnG3Oe/v0HDqCjS5QXF3z+1v3HpPS55gjp2E1zx6uk9lA6Mh5BaWlhYkOslIMgI2YmAgL
X4R8azUbPr3Zcakd+4mPJL8JQ+9O/B+Ezrs+MWeaPUqZOMEEf4a1XIBYJ/K3+gZGwPwVY8OMH1os
Q1BuWAVREhkTtyanwRvLowYJIQGrO1rdc2nzWTMXfHCFYuPKD54dswsEdkxvobul1mK8ybO0q6nq
qwxvUb3KpXYWtefx+u4bu9gbMcMXbDSuEOvFoCVvmEjtBWOKG99SG9jTfy3Afkk3PD3pRaOQ/XZp
IZsBMcGV9YEFet/AZxHm+E5F9EPboPWWS7doczFFzkyzCNNU+gj4IKlkcL07AUhigvS+8cR5YZqm
5N25s/We5OonsttJj5sVj3U5Sc8OtMkWdwu1q6dtIZBFoDUzSFD+B+crMElDonqXgaEHboU/PbOD
tEghNyLlPvZt0D79lpxe8cY1I9GKrUFFD5cgrQn+VUqSpylZJ6nslIckS3B5Npy+a131yGxztd0j
wpQv9C9cWgzEQ7sNkM1crmOT/8mYRpneujZ9Hf84L1K7kTclCBs6KH5lfnbeU6pBcT+0rmk0gkdt
uITcweaYQs8FDwQ2yBsJskrEVQAlX5cWUVAtO1ZATz7OEDtJe8tVUMM12IAgzABKgZPv6825OH2E
7SywKG2joJsreXQrC9fyEArB3KhNtYhTZb1sCii3EBt46wmgQtWE57558iJeKsgdxkOZgtd0AvMw
fpHR7RqtMZzQkkJa0M0qJdBP+yMhdEjddehVlqVWEAf9xXMlus3gjLOiJsBID9df7kM7YT/P4Po9
n0p+86HDNxxQ583oCLb/jVlCLT4CCxIN9qujHc7X++OBzGcwdWbErJTg9srWNDmwFqORjHtRiVU3
AThD7rVsMWrzEyxlRUOLiuOEBZq+nfpoXKTnHC93Q+2tq4JFws4HWvh/sjQh+zcCgtR+nPlNESU0
VwnU6oEbtrAtqPX0cbvFrAeuB+bU8CvZL/mSWzq/KrNahBFuTlW6MUBYXDCm/7qMKi6CcVbz0x0m
r0GfTrmdzTLcGcKU/bQ2YPInacmwp1C1rPP/RvRmLaHI4BCq7VtjexkorINwT7Kgq4lagD3oqh2b
i4P2b621jWguYVCkteYVs1/xW90VAEj3b0iF14Ttrwss4x9DkAW2cn7moBDZCLzaOBrOPmb0W+83
FvTJTdef1rZAPvzLyLH3dezL5CSZXNN8McpWz/dJ1TbqFc6tFFCpGSB5nMPcuYuKh8qGguFXpXj2
bcDWGkZ7x4cKFFQw62OE0OPT9bMFUi5Dxrvoa1TXbznP4OMXLoFg5b4/z5jiSgZx/IGoxkdEaAl7
OT2+udqX0GPX+vUizgNBrul6hncumdrKBoGGvDy/RaycR9QPSWa3yu7UGo/7p2enLvgOYK+Ow+lD
VsTPmPgExp/vFFF7MwkPKPev4uwDpu7E8gZGunw2g2SiN0yh2/SPU7DeRKpoZSebWuSgCWYA2cWJ
ltd7GAp/y7VzTUBKvZnawwAsluB/pqKE4ewJ7P2j/A6FqjaYNU8emb/F9cSr4XQwrXM7C6geBGmp
jHH1QZDplelXmJVsNqU8reFLROkONVHht1SxMzQwtuItQkMdCCDupiB65+eRHPL0NpnxEWoAd2lj
mCa3bJPRcXi0+1/BHha8SN3xQ7iiVZi3D5NJjA28Z2Jv1kYcVe2R5vnLYdWi+OHou/JQOnZYmm4V
vVYUS/6KJ3Y21164p7cItbZB8oxKkLJ4xJ8TgmBqLJDlixj4b2Vsqfi1QOi6rKdqkO9PONN6D9No
8T8iQM1iPO38ekaOptiWGosGIV5qIN04f6HElwR3BMiHTRFd1cV6xfVLUHIhEMKTSvUjeC+OC9al
f2b+R0P5vrqr7jfOCVz3+9UD5zhOHQpKF47YxnDPVylgzflrFw9ftcDR1aF/FB4ux5dStfwRCX/4
NNHVKmHWIg4YpeoAaL5sWtpCFnSo53YY9MKZz4/wrp95a0zgSOsa2UnV8ggL7OQi+wQaev0TvKsE
+FiIZ6AGoBasZ/4yCvFbT7lgAc6D9bOHX0vlewO2VRsTAEvYHu0tx8OGqW9BUnPZT5zQGI0ea1+3
0O3ev5MLNKlISZ9VMdcYI6ibFwK4TRhViSyqvCSrD2rxzTjGU3mCArkzkSEzjchBlPTa7biqk27l
VKJl33K6J+sBEBktN2ToFHJUheEewYFAP2C//nBSHGjeNOG+1jvUqykSjor3/Q/Sdj+YkzEY3hlx
1GOUDhuaOahg2CVjP1gdieG27ogT+tZ/hvbiFEUSBXEZIq+Y8/iYC5dEk6HR372hH1LAuQBzLrQm
by7+x5EwsXRGxJy+RCjFzIKlgKu/nElOVZI1DkE2OprLGVu0FY/kUEIjzoCOPYvjbrF3GUIafn86
0Q6iKRoP3WivO4kBkv6z9rEq2AOJAy6t1s0cbdrwLR0j3e2x1M74xqE2iyk/Gn5njLTXX4cg6NtI
FrdHoNxBkmAnRlbPyVWfgi34B4X6bhFtUMRsPX8cpGUTfE/jvviDBIbOZa/a6YaCwh8Foc5gPQkw
Ps4FPRkZjQ60uTxiGp+2reM6LzkIfzd/rJ6BkL8Jdri4HPNspkv8ij7b2kj4dkjfSfrerunw5EkW
nfC4f1GfiPY+xWpLS68sjS7pD/4dv2ZSwIRKx2ZmTuvKOtvzquzc9/7yzBtF4pgOTDQzxyhPjbas
hSAEjPdU0IWIg5Xdsyep01s9F4kpierc9YlVIkzjaF+R7cM9GVXdzUQiyimq1CuSD84fWFkfYwZl
SPio9Ont7OFrjOs/I1fz6WKZ3PbvkcPOYDyeY1P+jE/wdFdLXzdvb0QQxzFMmESorDOloH2fPj4m
8Vjh8Hk/26g3dmnM4tS3lipxT9RqmQyal+nkuKGsNQ5GDcqivx1tKM8Nz+uu/yuymVQm4bSm23LF
DAKW4HCqtnb0PdikIMfeQTbq+q6SYUh2A/y4kdeSGH/u4yXN1/Lp4DYmKzVmY/gpl7FBuPDTU1L/
AB+ld1iOuHxHupBrzEBhPNZf1TTDeuaWRgki9CmQ2U7poPp/HmXMH3UjLfarltXcCfw3kDuYluUc
KKuD0u9R+2bQgjOwRRNYV8KNJdSgfHAWm9vm4Kf6UGa0XUpTtMKsDfTjHQLxaP9NxqaMFtwXzxDG
estmXLGckkvuOGmpB+TKOW+k7NlSsFCYzklI0exdH4Tc+Y0Pfhtyb5nq8ULjZHZEESEvDquO5Oxg
rC9DoA/gkdc2kwN0aTCHLX1KzJoyImpSbxXocUcupEzoNS/27TLKFYI5y/Er3NNdF3iXzPVz5avc
Lu4EFsGBpjRibw9sSX2Ui56EKn8RqaXTzpNlVlwVg9T8Okp3aAmpzwJaVRB5SyDWUiqDlrmEibiU
hbrL1yVoTbRD94paLJNEPsrvw+8YgzeeVsB99aZ3/VSRyOf1TBUbh11XrLZ6AP7fpiPqohV6QqD9
thQtDYjKzvL2O9FL65TXnALjcRyE9w0TBY88MrOdr6lZ9pDCW9TtM1mAlqla3u7V+R13HVMFzcSH
vQaVQsL1QGuWZjtNI2K+LOyrNswZU0aVzsrGjh/sNy6M3hxQv2GvHqfAbxn8Lb1u+opUUj0ATNpK
iOooR+J3M5G5ROv1Ds+RpMzzJa1sHLtl3Oj8jtJV/+/Rl77lVaumSZGRcmCFmJWM7qs8E1Xa2Dzo
HHjWS5jduy+7qQBxR829uXTSPKxAfy9Nv+Q2GcCJYKBC1g40mP8/wQBg8i690ajgfL16FffMBFPK
y4Bnn8vRYg8Qaf0y21Lvyd695nu8L+eIkalP9BU7mnQ6pUWc1eufdg9y+x0lTbx5fs8i2uSSHOgb
gvQI4JjzA8vQqsAD8lK54ZIbBS3U24kbYLRLCA15aey11NarJJBRIJhgAC4R9X1qr3a8cyf7WjDk
PZmd5MB6xaI5jIRGUc1/4VbGPuXPWagkzcNXnZAANtOtsS9G+/B4LvDMr1iRj9ucQ/CJWBNxRFrB
yiLAY81WSHemqkQIYCaJJfABV1yAOoUsn70b9hilPbGY/JgOKG3bB+VPyun4edg+CLthrBdkHLsN
AJGNY/Wpv9jjZ6SW/r/g0kshp2K1suR1jYUYaj/kygWo4qbRE+5y5xoAs03SpI48VQBQCYno1SyT
SDn49wwQwW5XxBgta9IMPCNC11BEvuqRfIrPY72z5BzldSVliPajYhANpnXKQKDPYn0nuh8RJhyh
0BV6sEiOW02/jymdH1gI9hZYmhRQ1zf8UMZ6dUmLaASWasfd1xp8sFRwFvncngrvdR1ZgeBU3BJ1
2gb8+15JbgeIkKDV9JrjZRB0y2CGFSA/U4h4MztrYfuO5aGD0gzM4dWokZe6P0ogVZE8rKSH0Bb7
p+PUNnu3JbWIlYPCNZI2TnTrEshrpz6q+9u0lRox7fjmhBwkjx5pWUMiqN9HbggYyc6nvlGbzRo2
ChA7pwyVqUtC4rQ6kEpx5ElLZaNDH+TEum/JiaBKAVsH08dXyvmE5iZsZNvd7oAv7F8TJN32QG86
0iROFuW/CcfiQvjnIUhSzxQPWGzSKPuD0cGq2ad3QlnM/2ri3ggFdkFgmAeKaaoOH7QuN1V+Eo35
duEnRJahVtS20gDHAep0HtTQZVDcaYHp81Nim9/D0BDnshzZDFBlmHTyDCd/oIkkvYK8kZ7BN3EF
aVSlKPG5VRZV1lXBdredquS+s+mA1r0D9fvmpmFz0+hI3esfqA4ZicGB4uVSmEWU4YFmWRi+Re65
js+CgdW88NVpSEWlseI593rYSHMPkPpmN2RUM5iUw3ni6Ebm3Wh0Zhb0RdbQCmFzzAKo75mLNtDu
M60qsVQcMTJ//IxB7/eQAem07vwDFTH4JGnUcLiue4sWQx8otH5ZIdIhaM9pw2JnHpgXzGry4H+v
OGUyvrW3hVavIW/7DvGNBVq5ikp1UOATLxSmfvRfXMXu9pP1DCKiWR9Qh8ZGBb3V5IiNLEaG+3qL
0aty8b2KYb4WGdxiu369R5p3TZFtzIbqv2YXqMoDu7HPwvJid5gQrviyUksafFKnDEUMjih8VHZS
M84GZxdKPDr5g0sV60KEnGDcZLFpBNuqh/I/Bx7uU7PI6H8jarsmUd4l+/QcaibUM+FYzBk+H2k4
prLxzqxTl7xLAYOr/WLRWQp7hyvxdopoSZsoAfJfJOlwLnATqtNxy9/3qsAeav04rb99cGNoZrkY
l3bDbo9bGF/HtFr009l3BrZ1Jmml8Z9z9IUPo+hwCnIFxTwSCvmiZoJXbsQjzujXr+nb3S3S+gDy
vASKtuNOJdfzPhjhRXqtutnd/1ZsJ43yTmXrWBHV2s5TrmoeYOiQ2MV2YMIV40Zz4K2lVtTVsXDB
FMwLs5nzLUHMZ+Tev62I7NsCkY9qUGJYqnR4JUBRaAVwMNP+Kkei9XQgHRd5gC2ptErjO374KLBS
se+hPvbb0gq3LBLefrvnu7PDDrRrEY9LT+7X8jJ0cOqMHMu7OgruQNwyNsP2ENsKXVQl0f+lb+tM
WCCblT1hfjYVnr7UqNqZTgElCdXiXGfYck4pCxytKpiEBeHff1hu5792BNfJR4MqN+lK4awBmWwi
MqYI/4d4bDWIXyM79S89ZPHBew0eDK7jq2TW0a+QWIueEBv14fsvRYvnnjA/i/c+8zw/SKpZOkW8
mA8wzT3mhW5V9OPfUw5EZ70s6vhbE5JrTQN1W4TR23CDks3WpExzp9+aOb06jUorgH8W7pY0YpJ6
h+HHcbebkZ2GsZamOow0nlU+X61TsvynAFDUGXFi1XscS5O3fFNE24OCHoen340Q5w5FJyd8X+3i
MuZ514UWFvu+AFVcxwkiqu4Jo5KsqSUdPyKeR19Kl/2G3uXwNiLOma0q5hRU9sshKP00bzMF+p4t
xeQDY/ftPe5hj/wYxnd1CFoQ70wbMkeMpnC5n/pISJ15cN5iWH6EzjI/qWc2Ol6lmUUzoe54K1z7
rdNWjw8+Ec7O4X8XTx8+eaqW5MrLuTftYyKJkPJbRhHV1kWH7DVYIdgXf0UGM7Z3wYH0N5AgfjTj
nwU8sTeXvEIRpT4de71PghtdpBG9UBTTsVDQ2O6PExPbXGO8nsCCyWze0hocUFatFjdqeRIoRO51
BJsyIDL//pd4c2jHMXR2TH+I3K/esj4tv5QX9HkBfZmgtuYBSVTQDznnYYO7VMP1EfDquULoN1wY
E9pAdhT1ngTZXIOe5PgO//Vq+Wt2alYhWQBIXYv20d30gai9OGiMW4PBg2Od9SnqLq+AzjYnaf3S
shKJMmImHczqWR4wuonjI0wDWgLXPuiEfdWYtzDuahpkLSiNsB/n9GMm7Q0OQVMc17vYbMQyQL9R
L79IYrdizR79isc8bmmoMhUcW9/P/qTkPIaSYMkfasbsp+Qt4xBUdoIjJddt57ooXM7zlhogrlu7
Ts1FIbfL21ycqfSt4UDzCg0+K/X9rqNpbC/UFR6fEY0b9CqZISDNFtyazzsZlaGTwNW3XISDmWgE
LG3AlUWK6JBOSMPLmxfyPRpEnSuNrPVcJdkmfiEnpDH1EbTSX2uFFT3i/WSk3BBllX4sziLroZ6q
CVjan+lq4cHHZebhm5Pfub05Sbf8I8JXFn/iAQILDbPkj97QiqzVLtxQEAoGV127O7lU/v5k4eQV
4HFXQMJUeYa5wouv7D/tBX7o6ZLXn1G6QTcT8IenFjDQeF28r7Zon7Xneny67xmmIin80lDuquJ6
zVEehhPfE/Zd4MV5Q5jj3XpoKaOZlZJcL8ERU0ERS8EQUlnB4bGHYqZDBjJMoiKax5I1W4ZRSeRJ
s+j2xLhe+3CEFmVTb9ozNkYKm2mb432Ys5z1vNvCQ/o0E1yaZoeG2h98uqzwknU5OuOIomFc0Jcq
akMz/DzJWOR7tzHht+kKrpjoMj0CnnP2XJSiXYeOqaSglsaHyTuwcL7zS/rgp0WlK55wOdxN/HPJ
PEDkrWgapaoWwv8xvxMa6SapBC8e9cOhDFReMWh3Sw8LfqTdsLg4zQ2tCI2zcM2hiRlsyGMIIKiL
hKZxOXXkY7zb1WeXBzc67Z1X0AAfvKpppmM1rkQSOf57Qq7FAU6Tazub+Dw+KXtIhwSNz7qhekE2
am/FgnKUBbs5LKbSNBPQcQwGhwvQz8MNMwg1ApbC5i+4FOS9QUIA+4K+1pcDoEplYcfvr/rc2E7r
8sSg6dXNWf8zOkasGh7/WxEU5fylETYrYDnbulw1quk8hB7fYb+Q9FQ6YMkRoZiAcT2nITFCcnxL
22Rl+F4DXgOPHMU24JfJA82ZXttofe23Kzw0Su4dB5Xmky9fU8hgU9wZxkD2NSXAMyVm0ET2tmTZ
kCm2pYE7yvDMNEKY0bLsyg0jBiNlNLaHx75PUQUb0wOxqoNLUVa2bG6asy0VFxCC6+gUECrTG8L2
X5etmOF4LkFdkph4cWMIior6HWcnvQ1k4z0cffULb6o0qxBWUsXlyHW7zIhN/MscYhEBo5m9NvtO
oRp5joSyyxHWva3pyH0Fks6lTC6x6jSm9Bwg+ajuSsKNJrXtwZsR62/K8E4bVXLZLNE19z1PGJTc
7lK692IeOqq43l2A+5GVHYAY+xJ665Qtmx+FFbAfd3CboKg6COi1mUP5GMUgj10qt97XefNWTmBR
8N7b/HOVhS16IzjREj8fsG5N0iwUHVCwTiD8SyRB0h7q5enwSyO+grZ/RQjZoT/ZFjJqIRFxCOjb
FKU0jpv6Vu8UnbvU9CceLaIud2YW3oO3AI6TsD5g587XN8qvZhm+wmWuiwp0H9PBVQgBINu5U0m+
vi0zdAHmWhpDany7a2F/mHkQPo5DaLOLRMFI1nwLZG+8SOeqvb5EWa5ouOgfi+NV0rI4TBdshqi3
qUNQsJaGoci2Ic6PXzpyxTWnLMPpF8/JKcV7K1Sc9yR661VJxoir2+Cg4Ugjxmu2lgcV3vYobyb1
rsyowV7dXHiASieD9r8QMR4yvgepY8dGG3Lby4TvxgvAgktUSBJqjAptUOvv5yyEZqI/e6B8gp32
rdKEUJWSMIX8ayy7IJBWmD1O7FEAVZirL+vdIFVNlbClzmsbl0JTMHOu/HNC7lzuGF205XeETYz+
X4bo7wJG1Xzb3J6Z/hmKNskjBfNM8DoF8QysLD5gZuV6gXH276zavuwTfW1NoN7s75NmYNWCciHu
jotm63PuWzsapBAHmePavSYiGQioelBESJEfE0Fu+d1WW0YwnZcB64xYStMlqdZhdmHcI3VEn8jj
NOHmyRVTuRPMp0ORogXgwAklgOZQ+idDPxmQdjStrvZGKknmQTfte2e/IVwOqIbOS2j812y4pm49
i2m9dYxp72bM8euznTGXCKO+CaiYv530lbhALfWOpi/ACewgtvUPRIoN9ieH1wsUsLTG6pm91iKu
JU7ZH+mNsniw/k0tnYV5fwH1Gwf87Ejh+ZGuIeXkrmil8Whe6+nrC39PEmV1cLGkR1L6B8iZwnKj
JtiVay+63CXhAqogleoOUgzKxPeaqoDuBhIFWMvRrKu5q9YARyPr4RIuo36F4CvzrupZvXyWdLbl
zdptzxhtugd2VC8WkGrk0RyYeqHDm9Nk97+yGte1wSRft2+DpOUfXn5awnbNSRyC6KttjS8Dn9v5
U9OGYJlYHslNcjboJLOMeN4dDjPFc+v3Nn7HOA52SGurncRCpLlcdxfXat6RN21Px5PuQyEIhknI
AdqHzTBnL5YjZkOLa/PWiTHYHNvjJ5ynMmyNFQ2bBqHvgZ1Q+wtbCRvqijQQ7Mvi/BP8RBOWRxOw
3pN2cRGPOY6WlPRvXoBX6Ft0wicN4bEAA5gPbOrxDBvAF/jojeRUy0xrpnEW2Dk4cKPjD2Wbdd2p
L2nf7T64q0/SFtBq4HhFEOBCVfRVmSbhKXSsGtlT9cPH2qARpMiyMV6sXdOTH8Xo+jK8Qx/uGHzv
rfuzpzUcSFB43Pj/dSMITMm3jTZ//1iFqlFS63fN+X7pGvCYWh8ZqeMGaLowqjNpIaRAIodqEftK
BRaxxq9HPrOe3PKOA79JdBB+7pOXt/TXSdRqYqrbGa1u4vTKS0dJNIiv4h7enoF8O3dJGNEsBEtr
SYoQHDQF/zqRFlhoZ5qGVoizWoDERySPkNBf7Xp1tUqGBAZ/Tq5hFVGkDt5cp5ipJBa3HdzcNLRX
6JkjjqRMkIZn3BTTz1RVbxy5Mt43W8qddlo2qiBKInITr1G0WRjDBN7WTn5qRr5Hr7w5qZUfsYxg
M9aRUMTaqE61xNM9Pbcl0e2O/HyaMllIAtq+CQRy3CEfyKupyWHcaKM4TsedB1VdqsGFkHbG4aS1
PcwbQ0LzCma9ELaanyS9Sprp7GYyFWPpRXEXfZ2LYU+vHYdxTUpPCH62TWXpQGHUEldEYejNs2PL
DUXQ3CC9uWlnX+XXBg5h/DbXeYTf5PN1Lbkem+Yx5wxdMb8nGEVWsIUT5VEZnlTS8N3QwnWi1wjB
quXtCpSgArDdMcaf5B9hN4C2BlC3B8viAEflg3bm8UM7odVLBwDnNz7j7dYc8e2m/ypOMkm34U9R
tz7+HC2kMJa0Esjk6wQYqdyIDSFALa9KMTiyQzoV3aRZrWLVDi9B6V+tpfRE5tTBQ4NRvqf7Puf2
Ub7clDpTHrB0Ee5Zcw4cpUWMb6aWlXWzOXrpcLqaIWnatodf3rMpc8dyujriIO8J90ZxxbBhHIoi
qrdfBraMie8qiynDvJbdhrQCKBvedlL1eGzhq4l+9pfTDGxhJmgGHG6IkYnNPEcuC9jW4RUexyGa
Czgy7ysIO8xE9NhzpOL9xxcqTRkTb/PifiSpVrCvVppN/CZVAHt8KirBHvoCQ12Gee6kpGg4wQ9y
y7U60BOdA2Hvq0ADbwQpDrBmYP7Avbgzl/1A/Z/9N3j6em6e6cyE1gl/HMngJa3J1UOXF8uS6UZP
5tSRt8XEMf558xBBL/diuXuvOoIhUNn1r0uNCYu5jZGqHxyq6rQeQGHwWMhgQrKIlP3VoCLpw/Vi
C7leaekP9tfEWX3OFFxtoa8O3K880Zmr+JNQNUk5Gf4AR4NoN8Pmj6Q2sms25FOhgrqva4WEWa3k
I/EWIJ1PbcNV91iF8qdtpdeGajcS+wzEHs9DIK8isJGlzE71ZWGmc7ukPMsInmzVvp4NvGPTbvLl
ppCbhrfJ0Mk2qj6ao640Y2Ouj/6ZqjM98fIuH4OQi2b/gWlnv4HyzhAxXk7DC6pE2sme7y93T1KV
uSzqXARCdNxfku2ffOGC4WzQWVQUWI3wMb+mQ1X3DIRgApqr3uArXjaEh2uh1ohynO0X5d2w4Eu5
6rz2sxwJg/s24qBxWlJIRmchsSnwcy5d4vkiG9zuily7n3AuUT7H4edccb1+JQVkJ/z9O1xvn3UT
0t3TiGEAw2O2wfWW7oxXz7yS7+QBIrMWSK1HdklykfYE18YHNiA7MZJ5zxtLMeQNUBHcd3pkcsrN
tNnPxYyv/ekMXa9P8V6h1zWoHIdnV9OltT205I3784XMEMb2NfnjeepGqOjeLOWxSq+mADQVujqV
zRUrC2Dgoeb4OrIt4aEHocULsPDSefHJIpWfu2C8bWpVJvawnYeae+j3BYGaWHMh5+eUgVMYLBtq
4dW+I7Y/C6fsX/4jvjHzYqlO2NpQ+jsXTbtfkagkUWO5NUfpcMUPzUg79ZgNgac/V4OMbX8qGp/2
axY0GgPm02oPloKnCNIytxG9cBsA2d5NLyMo6m7fVAuDm7Q6lqfdI72qb50L9PLjSUYv5h18Z+yd
7F80vlNT0S5T4kTdRECT6qlW/tv5jw3qUmGvSlZaaE/uC+8Zv6i/HC+PfSbvsEl/+l2GMPjpm/h2
h30qMTgqES882r3i1NNsE8f4D4Fkbtd44L0p+RSwWU2892EDwIH2Pp5aijxPc6iLH4Sg8eUqoD/7
XNWQZVUiG8XJTIv1B8lDsVJakyepsstMx7oJDrQh+P4y4xgUEiVF9PSKcSJJbK0peVCR42iuF4GG
ktrpz8FDyJJVyvtPZxhIGq+FO3CiN114InnqBdcAGxvZjxcamPODuWIyEB4mB9a4zfEueUt5T4Ta
U2ubAnamxuyYPfBocqB+o67H/JNh++Hx3w1QDPTKFDeYlmKodmqSQ38iaQ7XO7zVkwHrVb2+EWnU
ZDR6GC9idkRblqyZrvgmZ07AZ64cmV1JDg38Snz/gxLMDhRiLzErnWTE751fhiV95iea7fEVTnOx
50Jp3zwyVFJZughDmOBsM6hwm+tPIadBA87YO5Ip+XzqlfFOG70OQo0VulxFE5C8HspWWOz8Jp9Y
bvrYPtpL8u4CvND4U7vA0k4b6y1tN2HUWne1gYRdArmNfM0G4I/m8+McNN/SzqhpOX3ITLlPATke
Vpzv6xCOan/FHZdrVW+sQ31g/frpTPbP0Xj2zVWYqJBAMrtcO/EbVQZC1TEPjCUmOBPTtv3gtbo/
AvqrAGyPaUk2pq4meuib2QpnxL1ka8o5hXjScIsgfmStYcQrXMNlQzaVxcWsaKfdrdyjDbNOj7eP
sUlUYMkxuyeUY5KYaur5yYl0vMKUnZ0BUWPTm35LT48q3qHA+powKXTRIcHVJytCiHXxFlOe9Tjb
kTcgTXyeEtLWnpvp8ts4wWVDxnWg+x8W5XPn7svWWo7ymORLYz69wSEPNXA6s5h1uDrUArA4fGZg
wrO3IbhC6Mg5uftYE177ytaQhQr0gqO+GNeSY0Z/XabdvLtaLiUH6yJjYSbrVJwvFmyxFmeZ1BF+
zCHIXv23piji/YVmoY/7sCBKu2FDSR/BHRVBDO3P+ZQh/rpQl0h8YYrR6PkcRLuWtFWi65gGXynx
+YHAKmiEG2zhNIPOdKwr/oI8Tz/iw8H0jrLINx6HQUT0NRwazReoHmkbR2i80VUwla68OCXl5U0h
Ig1lpSX210/lnDRu1qI7NFwt3vbeQqG34PQjoUjMWXNPbHrSEwB1jPAMIpnZy9HWhSjTSB6QxCxd
fTUexrKpOXIAe39/ugBeFPm5LvUtbuf7S9sgMcGgrIHH02SQuqqqGKmFmfKdaMuK5/8qzhKhrGna
ykXTPKYkL27VC/pbQDe6/9ZVVjQyCKvohYWlTP0k9Z9avdT6Knq9Z0n8rnd1kzXXpJ6ZR0vmSttp
2Ha+DnEJU9mR4zHkfR3F8dOBcGyghXtMdHrblJRen2BN88nkiOWUxrYs/q0UM11lxk0BxEJXuPFj
34b4zCmM/f/YxvDCDKikURIuDc7FJXPJNKNFl2Al5z7eSF0vv5fADV6hs68kouyzBg2FEG7HS1EE
oYgHLXqaYGIIfMYGeIdTecW2qXzwA2E9ELaiYJVyg5MGMSH6aqRPWIHzpUaO1u8ebtb5KnhDmAs9
/uYkkjuqYyPun2t3sBp5ykvin8vh8SgyTqr3JBPbRxqYH4mQWrr6xjVISIWnOJjH7D8FJBTMAoKE
P32moc2QIQaXz0NUeSXQKSsEUeybRe1D8rf3JOdIzj8rZzlFtV403184lOxLmEaY0Rz9lrpqlPke
8a+xwvgqmcOdt+lMpss5ml4ZDakWIpIJwBeRmqnpLg1bW8MurN4WtOTWU9QDxdK28H2HUK7lxFbF
7mzqQyY182Y04aiv2HJHTW5ZVcKq/7yEdUaAm5Ru2IYPrScDIKJ1Bz7XbD6YGbD32LMBABkiBsCh
3rXi5w3cEOTg9ACGzThxA84w7+ajHQ3ZTCPJqA6WGA1n1SpE9pUveI9fvB1b0PE5bey/ifiWD4wq
e0+MrcQeuxKp6HRqykm0ZpV/l0/TTk09y/nOX6R1QIflwuH2Op/q1svxv69ZdlYsLrGAkV3nIZWO
qUcgm3KnQFg/VtYriKR+Fq6adRY629jqcf9FcGsO4locj1KxzvOEBEOVZBAzFMXb0XV8TqvtUYHZ
Fl05h7dTS5WztEb9avFES54+4vtL8epJbm8+Od3DUkGlmoyQogB2ztC5wDcfGzwmV6DWENIYai26
VSC2NIWKg5pTmkypf/zD15eyCi926bxLaFrSGC924jp4UV6pZD6mrN15qC7Vh7gotwuqDHGSZhpp
kDD17WdUj1fk/hirQm3s5YEA0WtJ8xPFF7RJtxvVuRAOS8DocT3K31jysvhQjXcpXbNJZXRI28Cr
aDSnae8yUYk3CHGrJJbwir+Hr4vdkaoZU2vZQZLzzrOI7Vtg63xlicB0rrI2bKZvRzf8094MceKZ
bAi7IHQ6jFatJoThsArGRqDgea8CUd5f3Uh6wFtWFtWLR0+ZHqgPKtrkFCBRhbWWlp7RWhbwxlJI
uAM+lBPL5PciF3di/2UnKKGvRA5C6hmUGNFzx9vRXg+kNli7vPeuOXBS4rjp3FzZvBOY85z+l03y
egdolfbwsg6hfKqWE+TI8ybHNr+SnuArjnhTc/xtSRLRLUXWrdvlyZNUWVyMx+/wQ3WspnN95OXj
8+23lI/a+d8cGzhuib+vDAtW8tdEYXyrK3cl8LYe/tShghgYK1jD6LrHh6I8l7vbBzRTmEkoMD5j
TppbLkfzflcqtoDHSZbJ48/oCWspmPRj0A8NdLz5WKVIgLinHKXf/Ozzqaj6U/k6ZAD4DXYPdoZO
HGdAEOAvT7mHVP1ODSsNR2Lo0yo2no987T+oAZ4rvcyzgVnK5YEAtZHV7VYQotG6gjnKi3mdeczU
OM8J5vNwen10tq4+tJtUH0TBpZIiwpYZvCIMhLRTqduBmn0pBwBnynZnadIcEIo05V2SjM6txVqL
iwOQqYaXRY4toxe53WLLpTBZsOZU7/C5UsiTK8ArcTfV97ENM1ee3uY2xkwzMzk+7XX5D4LNHNLv
sfMbA4Mphev6auDwBKyHtu9DHv5RxbzVRohyp/D3JovDyPSOTve+ZM4s/UabutCC4eGjaAymQY4I
k0R4GSJBSa5z/nbGg9N/7Cz4pE8fKgrMzwRE0vJXkpBHGmz9Lwuh/H/VlNAM8x8OVfCQeJ78fmDe
3GmKOlljVOepdYU3kOdqREyNRWkM4Lq2b+PReb1zO84AgXbgcCREMvoZrnBdXK6ioFASVDvY0rn4
0osp8SsSQs+e72jo3muQDdqCYuh93MaqSfZd8a2DS2wKwSDx594l5PAAPd/L1d9wcwaIEPS1uxIM
bYzeNw7OLJAjgSjuOVRUgtkDgpAg/ERjlkUH+ULyHZtmPdiAr1l8R7+Wj5O2JAdKPpsER86v+sfk
0sbJ20GvI6QH0kt8KH1UJy4gJ7d45+8gZSYkPKk7992tHj431yKnSrWmYCLNJlF4YEU3q+TfXC/6
SS4Cdc7Zwb4KXVszue/8HtAdUqPl7kBFLCiS3GjZUyzJTXQEzsWTmvzfQfc8wyu7hkXJHHYn2BBE
+kV8HvyoSFg1t9n7My6kBWGqrvAkoBIqTB7muCiT00I3DP6ozckp9Jy0+nPb/0CzAoivXB76mC7P
HhTb0G3eANcVKKUlDBxDIRdGHzT7cjk/jidyDnXTDZyNEFMQur8BQJtoUb2fXn+3Qle7liYSd3jE
bf9U09S2uVNVqCrkcgnV3/lLsDLW6osO7MV/MM5Vinqm7uS+onL3gVZNMLAQ6ajNd1UfOpOoaMsL
ei7h7WmAAOdnalSEWzCJnHL+2JinhD0sH19KQUVJ8doTES1SKIFKofMdzzS3upSNq0VxTy83mAz9
YrXzms/OEOwxaK1ieoGpYUrfhacT9fNSremU2uF7OGyGz82j1g0flO/CjZOO3myiKzWn0fr8p7qP
EIo/KXhySiURg3f75MnX1En91qLAWpZ/UqWRxeUA23ExpQcXxri1kPOD43wD/VY4nAgR9rO/iqe8
FWe3/G3GP5+aUZRD7MjoVn0eIIYrDhO1mx42y7xLZKsUd4zfp/P/qJ8M2RQQcTCtu+pTavcoutwD
Xdh658Yqyrfpa0RoX0dLJPeDAo9U3iwxFe3hqK7zy021Lc6e8KO9jIRfU431YZlO9htXJQQcV8Q5
cwr0E5jEOx6inqEeCCA8gM/lKaOtOwEwyswP8VxJAusLot0GZYiPZFJXoZlRGZvBcDN0KNqxkqeM
k4OVtshn5tXnZnvygIr0Lt0ycyBb1IVBPg2EdEERO7hl5Bf6DltS0r3RlPJ4Wa0X+yo7c54zNZn3
70S7mJoO5QRUXuWlFpZJfIBrsyzCQNUPPbLr/6cOL3xdEv4RqD6sd69cjRbUfpceN4jk4F3lV97K
bDDOxc9FP654avMfUUJQosG29+h9NKqI4svUu+TJ9IS0tfkJhW1NHKgfCG/2TCopubrHZeEWfsyo
IXBYaP/FIcUVC//2NxCDDEMymeagJjNug3aByMh/xuEqIdBBjFbKzlHw3ouuSOhlw+E5B3w7ljjl
t1y9ODonKueMH5BcC6cdcSCv353Ks317npkG6/V3GC29RVpFWvvYoxFl40v0eA0mmOtMWs6eb26F
UZ0ylsf+my/zg6N030cMy2woTBegXg1brKK6UaJht28NhfeQg0lMm1GMiHjklo0NrJ/evk7VtCOt
FH1FJG1IHcpVsjykedhLG1fsqw6bxESNEFbZnX69pJY8538I2PQFzi5DaRzqNnnIakt2/hyLyDoM
s5k8CUYupyp1HpDnzh1/mery7SXQqWiPQIzgxgNKhutWmwdop74tEi397srILUbbd1ahg+hLW1WM
/mBQ1YZH8/FySwS9HqeeQQEHHNhCQv40mgNGGqJHt8wPS7PwjN/AZ+Kmz5V0gSW9H2tr1MbVLAfF
zCrwfeOwGOd7SCdiAgNAbceO/6WBQIpOLWMXRbP/LRfJCl8Q+k64Ce/UTXPVfiJB9MGvaCqiOwqY
h9mPBCbS315ZudL5ReliGQ2j3NmozP2e/6POI5of9Pe/sKyrFVjU0m1O/Yucepo0QHDrzeW99HqD
StXAMjfjsFTXDOIwe0eInQ7zLHdSxKKbs6F20+szJ6m7ENbCSOoYWbWiYAEm4W5BN2QW81a4kvrB
AfOz2qLqT1cKkdIRpJIX9E1IEaG4oosl/1kPcEr9M3XRyGQ7acfzZ9fJOA1E+XA7Bt9LCH0MiNqU
fwXVwQB+V0kA7im9ca5+Kc9pX472wBjldnM3wRRnu/Xz5o2gswKlINgtFBKCnl8ljw4newW4FScM
Lmyxl9hbNJ0RCBf/38EqJtRsX8E5jOzrmDCipKBZtvG0Pe//ZNRBx0j09OGBtI0MzCkxgLITQoV9
5T59BtSEpLOApEa5KmmyUGuoFI8edorQCMz/kdCyU6XR5t8AeIwrpEVopV2ZTihqJOsdT7Jx0NiX
1qEdfTnzZ2RoLfjTp35xjYSh4YE9ue1k0SKDR1Smh+H5xxUyGrMGW+D66LwBPK+hSGVFp/D5YGwV
cy7nfWY5P9SD+m8BhCQiS0dZsAsgEzcN7cs7jh5FnUBABvpN+QfjpxTK5NpOBDB6lkpXVNfUrvjD
ipSIuz6O5WMishc6AaCUr27E6Ni1DiNSCpgOKxVvaq7Oqq1JKQ6qJBcA0N4sMT+jjrg2ie8D63r8
ofUAV7LnOr6cVpD3DbKfc4UwjFTs98oUO+Sk0FQ3QR8tSvUJldn/T/FGLoYdKqc9wawqojE0XDZP
rpCfT5GztK0k37qxlLikChe6dF/nuiBaCdcYKE47kBIF0cA3RVWJovJNcZ6QdfhbnejTtWsHF46I
V4eNQLM3I2aE1CqfKCpQ0EkBBZKGKe+UTElJ9sSZmzepYTySLzAAMjawuoad0oEg44bm4MhxfTOl
ckeH/YTzv3ahLmWNw7/1we0TZRPu9OoXV1lgL0rdG4QWxYxwekWtAGv55VByA55PQLHeErloNBTb
I72UBoVe53JEFrz/Stmuf5i9g15w4124ssZFJ35cRlvXE1GZyArSvDAtaFDzFERwb+0FV85i7WMf
9cMQETmn0NygANLOw9zwCsdkdhlfIU439UExztKE9plnLByIYY+J+8MbOKB6of6vNuCy+avUIVjx
CrMDonUZs/6IlFPmxdziDAGYA++qqzFntrItzy5/+aIScoC0EbUeJ+37291F0k/416G+Zvbdeyf1
RuubDx4Z9p3JCb5dmqtyUVsH9ioe6o8aB80GWvWqdOOGofwtOCFRmbZZcOHnbuTovUSwLtaHodbE
cH1orXNVQ9ab980Qc0nl1CKuql0iMbboXteSfXnzo897goSRAobhe1YsqIRBTqp53Ba9cLYDOkCw
mbtPvdC2N+ytyO40T9qHULJoGCAdhTb9letBuRLkUOlnzcHiJwPihvFW8wk2ssJrNgx3hEkHSvBe
Lx7vibMZOElZJs4nWvilye6KoQABe9fdvIYTCNKLgHAI9uDKCD9Kqyy24roWFvjjWk3Ua5DEzBW/
cE7ohJ0932GP8kw8Em0tkQciVF9HIyw5IussQT4yatAbZRi0PCJDxBGXIVBl2lGHNXMi6rdny3Bg
SPX7eX4tuJqwKH4jsX1KQWZJAsYpiU8PhoYEboaNebhxP/17wih9KAaC2LXOpLvs2XHiCW9zEh0U
1HM5jadKqkAtayfv5B+Vm0h5/1SQQvV+PRiWieG9I0e+DX/mFs/hKRi3rOzMoz5zptnV9pIO8vhL
54LbTKwk/MaJx/gr8u2anudoLwd6pmvugdiISBfiLcH6WAmL2f7wJmVX9oUid2Ud3pLPG6tnBS+E
OVyiaK6mQepNY6L/04AyO9ycSTVAtMgbMl6nwY0/LRemD3gnEJHMlsHw04QWS+jcm+C6pxuZI2Sj
GCOCSiMfFufDVzI88JryuiGLyhMjKZcpkaCF11KGIqShGVVPARJAxSraYrs+wXN9//i4RTnFNM1L
a3oC9J1FZwzuDciuVo2RD10xqru/jdmbSdNYGei/aPbHGATcuyp6hFD5t1/ZubG4+lheFQ1qv6RQ
9XmNU4drPfmExseK2tbDUZreOjXx1nIDJseBvZt1H9Uplj5/GEsKh+rM6YFU+ZOHY1E1giWWIMeE
qCE520ks2YguJO6QJjnHsYc6ymSyFHqpl2xq0wpWFKCDvAhX+BzgZjs0dmKQesMjrkvz1WLfHjiF
TxF444ayrNO5nyKGawqLwqPZUgd39Up/GEvnYv9sKRGWxkGO3s+jX7p+OniOVkxX1obqzB9eg5Jo
UcP0x10DjG5gv7bw7M2fJ6iiUYiwPJzE5aBK/0xxTBnC8jr0K+B+lEIPsPwzY3TnYUzIqlfDqb5c
rmNXrZLnOlwPQ7ly9V2L62vi5kmVQWLDYOEHJaBXRJSaiGMpPZ6z3IxgYJ7/bLxJ1NSnjzS5YVze
qqmjS4F4cBRlgiCpxCdJ0EOVRZuVPiJNmemve4R8VUGBHSDUspcCosP+VDq0Y7+/4+SakN59S9ir
ny7J79vZMJrhNE0aQFwxqIpf9h9rBXy2LD8yqIBsPI/PUSknKWIGMbJC19+pAURJQuPrtBY8LQlR
gRFCCgd6DSJkz1c8mC+dzRCF+6oWbqufh3ljCAOqmE1+8650wgaZdI3KWAcFSErSYP2QLLDYWNe/
1SQdpPzhn+NP50xlCht7psBIv15f9t4ATHCABAXo3XhlyR+7/6sqJvO0t+4bulaT6353swH3jdMY
4AnTF+7h1VrnGImozfdGZ594tzQoTu+FOtYbJ8rQc+XdJ3WRIkpG6v/JiHBQLJkYU8EKt+oW9Y5l
ijJErmwB9H6gn5Qm1yL/X71/iojFPC/mTHInbSSCG4uq+Zlypbt4uAHdxrpP/qRJb//4L55OLcRY
A38Jjgk9niIXlrQbN8nTgB7Zy60rIMKOZKqbI+DuJKkfuHbvVHbWrShLMHZBfDMGuu8LB5XV8T/o
Onh8FIwOx2WNzEYToGpFPhlPR1mXiOFCSHYM6D4zeI9yThcsF+JibRfiN8AI7cvVBeDtXofRlSbM
fRsASZHR78/YVbp3rOvflrLE3TWyXbZee6Iu0is3Xt9KykCQzGtQySGxOj+6A1gQbbPP1mBWsz47
GzHR26vQfIBMWLeCpRKxZL6Y+4jy23sQioR0TmswN6nR27wSK43/rmGDgbwYetMjpK9njPIsDCcP
TW+2Q4TVg5AQCDYcIz/3gFrR6Z8HkMTSBJ5oqodwU2dcdTc6K188n914Tq6daQ8ZCylVdNL8PmNb
RcQ25T5JPwjshwXW9b5KQcIRfUIkYC/QkM4kF+7ZfPqijjpR92G1IuRSWwNnxCQMrRjNy8ajd8gN
P3GOFKAmdlNktlahqDmnTmLObd/cJAkJA5oWdEq4kfRjZXOPY8kGWIhet7cvROikQ7jokcBaMbcg
RB5+ZvowbX98XOWhW8mKZ6P3ttgm1oVyIYqajJb5Htx+VwTahZiSO7ev8Yr4AVmIKDH+Lr2PWjpp
35mrmOheMiUawGWxQ6jSkYoZEW54qq71TlcIJbrHhznFF1pwHiRMDtzsu3d6ZVaXZLv1UKXH2HMZ
xygLcHDAmKLSmTndFm105l23mrdd8gFIOFSnu02G5Uo5wtY+hHlLxn3lhbEqDA7fKuRTUnJBiuCP
5zjJQ4uiVc3de9KKh4Szl9Jr7TKDZgSOqULjJQR4XLx7ZEZ+zG0BGPXDUoBww7Uf4YykGPuS3nsD
uJedrNhyRvpn1EhBW+TsPuJ4VbkT5lNeH3Nk6ctmgHujIM621U8bovXfJeKaYQxs+d8dvJCQ5QTm
x5QNnWTykZtVMyTEX/rv0bZRDMIUTnNflwRqM4EfoYHj9L9QwnGaAXgIbnjB0U204smxzw5Ewr4I
H0UopJo4Ry0zQtsZmC1yHbv19BzBAzRYJrPkZC32KDu58/PWm3nJCi8gWTdok1eqmkSuJX3UDfYB
ZpM+jtLg/eeYzN45aqe08U+6I3nR6C2I41VrQF0wwGN/VOruqkFf3/Rp6M2GIVwgCqhwoAc4tg60
/kJHFLPz6nbwryiMj9bWzox58x3e3IrZeAMhf6z+wtttuPN+cLo7ku2ZQmThFlEDAiOW7wi01mHJ
m8DhSsADUj7LSHBE2S6k2+wqFBGyIbwfWM0YTZKyMp8ocWVQSDA4+3kHBN24aHjkMzAKB/3r8nQ1
wym7fyMNwWUzD7a0BZ7GrBCYytNTcyyAVKhGwFhoWAFLN4LYGOKBojE55R8rnhD5jfRb/qbPTG7E
EWS1vO7wwH95mj9cB0Dbv5vFcfvHIyA1uE0jgHt2JBEqtB3NxJY3F+LK2ncouadgYu1uZ6PDFwFb
QjKJCqo4dd9O2sHE0weUNHSwuc1bSxPGvnkyzuZwlSnwDP2j712Cu6glXYBpX6xGrcuvMv/LnPzq
3x+/rttZ7Z4Em8/PVez/IxlvMgMA5ostr3voIFiO+Q+n62SrUZ51yAedpM585TyWslGRsZ+o+h9u
Se4ahnrK4nIiv1SEq3pB45wwjIGseT+kA6Pbi8THTAg1YBVdAspf89oG32KhOkezLvbZuIau1drA
ETn8GrW8SD+ppA+bJukVBdBOufsjSXGw1m/8dXcmK+y5MqqI4yTQ499QsWYuTeY8E0WsnqRdQztb
auIJJMejbh54jpE3+HEUAq7eVOMCbv3W/wygtyiAYx1R7rlVxZ55kV2idzARYEuGOo0gz6XDNw5W
uuUXUPwTBzpC6+Rj6UKGnBfmtNQPtn3flazfXattPwdgtl9zkY3DGQ1GZoz6ckTev5s9Whn5ltOG
mu0Bcv6r+wk8do9IPHeGboP4MnC77+JfLZ0uqQFosPpTj0rpdlLNLhgFNC7dvqz/I5fWDuROTtjJ
WULU2WB70bHEoYj1dLwNqmS5r62bvJ4xedLUJZ0q+I3osJgxNqprhjtsE3TmnB5H0S9wM5BAQIhp
sCWgEkBzm5nMxc0Gdpzo+p1cKv7lAQh+GZl5xp+LeqSs5SXHInD1iwyilJg/Fe1dBwZz4bGXMLI+
Ac1Gs3dB5jLoEGi7LAjXfvpZa90PAXB5DGg57fkeqanixWhiqYUHZj88kSFvSXIjvO959P5TRZXt
MvK59mbaBdG1f2xykZPGGL3dYpxgjVQJRpCCU0WjavvP4azRBh32gV8d0FI8/DzsHKd5BHRSqpoH
eW7LXbEh14sEChaTfjyGEGHUMWQ8YVKLwXwZ2NT9dhPvKKakVRAyvPis/SXY3+xsZso1ReizrPYF
PLnGWHyM6ZKMVqFkEdp5sYRRWqofPhD8Bi/YhzivaKcAy92DrlqHIbHPr7QWmCnq8h1zgewn7y0u
5J9wS+FDPVHI21SjALJZU0qABlLaBAugjJn75Oya6tYHz9kQnW23wN2FgLikOKx755g0Hsq/HO9c
hjUbqiT9cC0+sX1n3SbtCQlaB3jIu+bnwtckTO13d+UCT0H4Ldr+NoF4E7jmhdhw0vUg3ubjWccx
5bqd8YYa/vu5DpkeN7a4xC2fEs1PMT9Xa8SEZJhCgbeKhYKYWOlnbSTPhWKjijd2qqztYK8jrv82
17afMYTkUtpQiDgcQ3TnPFTpIkp6CCAyTKipjadnd9c9V0aslpHcUE4HMYPk1w9NUesYKnsssI8T
gwo9IWF0ACLX0g65ls3cPRkk9ltWafOBo15jx1kOoIPXmwOS3Cav1qpokq9VsTXjNf6NQCZhd87y
OAySi3sWJ8OFB2DZ2fGZ5I2UvMD92Z9M+NQTSuUMdvneV7zMFt1abB9oYFS1ZFYjBp5GE1KRNTqQ
nanKY4TzAjQhzabohF+WDF7Bv/nkhlOUCUft9C6AUgdOPFzGNWQz6tJiVlo7wudSZgIBnJEpaWNO
wQcD9mLCP8sOScuDjUC6tEeNoxAMa71PqFmfR1iBq2yoMpPRA1Lug+4JtYSKJGnqKSlMuQmyEAIc
ns1Xt+Y6EE5E18DZzFsvfYO25GnHPkm7rfMQ/rB8dG8gzgcOFQSPjtfrMkI/07UnC6tvDAOTfjuE
KTg0hmXYAfaCnzJFmFX5/gFcp6TpBavyHYMdwYWeJNG2GXvqUC/t1ZeNuODLzLS7n7r3cikPwVle
qyDClG5rphMNDQrnrS1KrxxinV4cBqkcqrf2YDdP6m+cG8JKykxvSzpf1cevJr1D5wub1et3oaWu
oT9jpbNVfVGwF94oBWayYKkEdyIh5TX9z7SwHR58U+OoU1PKaRXXxh6ANYWbnAUQRurBiAVlVHEx
iShf/2QhjR0prZiNaMxLAxfW+l5IWRI4taGJe3wTrKJGAZCRFtWTsrOH5sAjRMOHcVr0rHgtpCGa
6YsAHryrAJKv5P1S8k74nTEQgFUK6V5QWIx7vEaV/AB7Wrx8Ishhor1TuvxwENJinPBz8McAeWB+
3S6az3hmufgE3NNWL7uppBvHxoMYsUo0AWpblLbWVs3d910saOJ4ESoVolySsrEauFnOwnGPTHdv
6jKYWUx0REzUyA6uTEPWudbhodhDrN+LfuNrQUBEpxin15t2jFGrkOo4a4udUwDbl1WM4wrYI3Rs
+PP9fwfvBAED9ryttUGSIImAFijynHyEDAhhfLH63tWXhg5qvkLpbKSXEAqodKQ1ne9+tFbOLmL7
jALT9rDxKhNTqj5fmqRdBjkNiKbGq6oZRKrfgI+2K8Uz21Btv9AN0hGs90fHoiOTFe+VmApoSUhQ
3URBeX9vD897gRPxSABV8EE7PF3jaSApvIxFxv/ftvq6OV7jOOYcP2nu+iTkJpwZ04oQLK9ANTvf
kBYiVazS7xDi9lcukLtrwQMt88w+PZ1ELZQcwq7vahz5D2zpSu/CcH1nvARhkkU/E1zkHiNdb+8h
HgApu4FmsDOGBpf0P296O7zY/oI0U4DGT3avPlKdC5KIoxP4VVwO3N4nEh1NxuSCWX+p+7+AmwsC
X9pPMt1QkHrmEu36UEqr/ibe6//zi1MbkN8+WROFIWexZ7F6Y2rLTF77Mbxq/uZwCQcU1COR0oND
iTQgefwL/FtGrPmMI5Mgm5QtnbcmgaVTrZ8j2P3/5K7VsV0yxY/E339BUkjj6tkWMYwSY1KQbT9z
M1E+WN77O/WExJXCvJmvY2fkccGxHaMe0E1jl9iC2yR80SC7Ah7QXRGyUF7iq2xadvZ8PDcjp3JR
FXUEhAkTMD9xBa6pzyS5z9JwlBCdEZNYpjlZlZSvZjG5S0UvxYUn/SoWmjnDDx3lvJHlZB9Yp26V
NRQv4xmOlcvZnzRWa6aXX8E4gbX688Tx5GDdiZN/GNSEAJ85mJUnQYXZa39bGSxphEbnjoRfJX7G
XnL/RQxgNZNkO3Cu05IQbR3x/STpPPmiIw7hZ9ggOsE7Dlnft1YQS/DD2PuYNksnicFi6hc1SdXw
Qo7vEfo1Pr/x6/8Un+arXI1ReJRHWa9TeCef5s1W1pw44A4QESR6Xjpn33R9Q1g/x1Os+2Sq3w2s
G//atnHDuZo6QxD9QWbtYN0GtL1RILp0Ti/ul0v9LUuufMl0wRImGiL1sXIHkMH2XKQI2nQSmSV0
qZ4/sOgT6GeozF9wYM8GTj2WAcuwwbAo0+B5K/vWeulzr6Xkg6uinYdbO9f1BO8yM88UrssP6bz/
h2qQfHIwCLvcUs3vcoK/7zPzj+zofamt0ZeV/o7kiupdHYrX4rSUjjUanzKZLHEMO98pAA6Ea0Mz
9JUEl1JQEaAhkpY2QeVQlWs1OWyzcsi2SBBqMInjIDrjsQycf7v4sW5aSimroIQoc6WoTmhFXWoL
N5NNDlZu6sqyqP3CtkuoW7taDEGIEGx24SJLn+iAsGUQzRD7tN5cm4qB/VMZz0+6FXffXU7xv0mA
PlkJdhmhzppXGWiKMYhtyC219HIF/yaJS2BCnb0Aamn83qtl0QxmOCyZ+SiPzUItvkU0O5Rn7pVD
Z484UiCSjfbdeU7F+LNAOyLZQUkDsL0CjPzYeSImquHXfKlNm3LHGoCI9rdaRq7D7vzY3FTu+ra3
YL+yScJNYRemyXA89jO/WX1gbVUqohXwHI8wO2OKl5LIS1VdsnJD7GyC0isUbLOZ00i3SDkKvrG4
9Gwf8JfJ268HUmIrhYpit1GxodaZxjjOQB73nJVrjkxyIYv7qR8n6Vn85Vpyk9WTtrZdDLH15kis
iiB0XRDf3RxhfgfGamg2uRmA9LVsJd90351Ty3CLHYv7AkBxHeW0aINMhoFAOpnehBGDb8A7SHHa
u3al6aJc73oMqaZS8G9TpfjG+uf/dkt+658NRgDajQzQt4b8RwOH9UIuTMR7A8q5rt8lq04tAFis
0a6JH8YrXrLr+oiqRVIDAQlLhoD/DpxTZ1RjZcip1iog3A4w/4Sr7L/xVW3yme3epscHhYLeX2wZ
regQm8Ku9fBtAXxgh6qODjv09waHEC0w4yoAp2L3/YsiBOagQhjZ7kSHTyhDUYgqc/5bAUa0VUQC
MB0PGlKNchNHt2pkwSCZgrfVVDdkStgsAk2ttsTbX9bcpNCee8EDc/NrDfbl82YPQR9wmNMMM1p1
xyBi5awVx75wUyd4sfsKKV40QgSo5qSudMAKBe5ZIdgSAQuMMak6KKlWeCSEmnmnAtnrrfnx2FTn
DbrYN1GtPb0Wg4g8N8PEH6bcn9BuDy3MadLZaoh32awAupUVDt0w8Wc5oHW6tDHKyVLT5DhUe7kv
6uC+6i7dO386Rgwvbi6J+Puc2jRIHlzcCjezL6yT4a4nf1PoOjZ2yi0sQaCK4thZMF0OJI26J7oj
rmC9OWQXZCkLooYihKqILqa+QUK1VaHRqov98zwRS3+KpOmhUV1yFcB8u6XIi3aGWyIbBVgMLsdU
2wx7q/ejAok0lLu+eVBpIl5u2IV6Dd/ex9+Fdyq8cnPz7uFPRb5I5e8RtZGM32DRr1K48QFeYLC4
2pCf8i9e3YussHCkEmbyUefbIqD7QUiQgUo7QIQOH7SMIuRLCUatiIJWcFO9s1Cqr8tp/+3z7HeU
xepHMMjyXc2qyiuHgB/H8L2zCxg4RvQ+ze0vDSyJsD2mICeVxRPbAGJmDFqwrDJuZugZybARCdXk
7BRgte4vobVh9RCAU/xUo0gvxmT1p6WjWMAZ1r6wHl7VEkc0b03YZ8jnhUASs3Wl8wO3TvKHfx0z
p7hrydvoQyDGJ2IdSsOmayLUupSJ7Rul9H/eoGiZslP0cbmKvzV6tDixTA8wPTK7VplKkZ8cOlJx
oyU1ZwqcAFn/y40uxG09qAKWFr/Nx0ml4Z91FxqLoFmFblGkI9oMwGAkYCJerDLyJpcWZi4qlRTC
n61fQIv5sHgW+6ev2gtoJ1t73tsMsSDxsw0XGEMtEW3v4OUEGXG6wh5DsQEDRhLWKoYCnYo9yhFL
fr+1ZJ2JTxFJfLIumYAeHh3lKxs2uWhKhq7TsvF+Q4Tmob9PxXA6XwNmhcfEUUB9YjYAgWmpJBh0
NhsSd1RK2swZbTmkwGGUIFfdBUICQAjxu6dXgW2N3ArNlePHXId9T/kUr4PQYyyGqGMHxCHJFQKY
g0Ef7Hd+tL2Zy54ZcMWQJJ2adbudZ1WG03sDvR6vyMZaUBcy00tCePSNjlb1uBi5cySlFdWRcmkk
qt3stC0aMBvIFyT8uHgyGqrmHUlwCb+xJG35/wNsXxOb7EtwEEVRDE+cIySDmlEb3MGO6SmdXtNE
XJ2Y3+Lo/NzdYwuLCtXpCj+F6eAhgAjkora0O/4aGaIBYVbGQZR5cXeRcl3d9wgLhtE6JKwyx+0d
osaXL81iQgujlIJEWrCONSb9cJmhQSzQRf50/Uta1n1avpoFnRiflvOcCNlSmJ7p3kRnBZ/VDnf8
c1mRXws+pVSZLUhGvPJJrI3AsPwEAxyAv1dXoMGCLqq+SbUSl3F0/hXMcN9MLwI9zawEWppOA9dr
VxBZmmFo2/U9nn7P1fCp+Ajzxf52DJ0lhVSagi3ejkZ/D3iglqZh8/1oAYGfqdTA9FFXHYzsiksu
oZFtQ/7/4EcprO7oqmOEnOTimL4FkjyCe+pBPW0zhFJLuvQ6NnCm5ZzorXawYxnC6Dz3363evJgA
TUrZTLKhn64n2RC70Xxo4D14n0HHFebqobR8ktZ7Na+hZoA4KbP7Fr8Fwq4Pb5UyyqcnMjDZOIHQ
6kgi6jp0e1w7vlVHzc8o8dsZGvXHO1ZBzdDkcIdL4cWeLVGIsD8+3fZ7NPKZ+DnT7NsQlk9MvPi7
qx6tBzAbO2ahe6I5SPOtRrYbofg1vZg7FYFQsm7aW69Zrqgmj6wmp4oMAvCSBUGs+K/6XubA3BN8
t9pJUV3VjvwmUDHIecsd3p/oAV2CqmgMj8wD5+sql+PGFW1HgzdrTX9FQU5UjSo3YrIOcJmD93qv
Vsttr7lvQ0dtwzozI7d8z7wrtJ2QRkbNp7zy9+/NMzcTRc7V8rDdhvTSOEhzP2sj3FaEWUsGGEOn
iCcXvrrJ/vxZCoepyPX2vQBqPaEav5bTwqK+TqkNWSsQKKm4wckBm1PNbon5VWILU3z6KfnyoKbk
0p4ZFbyqeVdQw3STKoFq/N6rnwiIkLLzN6kucr8/WXfgCRCJG/OHuNQFhbxV/X03q4tIN890n/0l
O3npDsKSByXQFnEN6hJ8diKjhwjfjznKWiAhEJYf3/QsGIt3AxwYcLu+fQQ3TiREGZuILakjqmRK
deuG+4UPBCPlqGfBLviE9HnQZnTHEbrgm1sXQdZh4PvYlEovx+eVYnm8O1ipNkoDfQAEqIkB0v1X
sDurIYaW/uErYy1lOKx/6avW86Jhv7tIcEUQ8X7KWYC4clgMGt3NoXXIa9iINa1BdqNIh8Nf24Jx
JfMNO91oza4n46QFlyDMtPywMwH0PcAJ5QaaQp9dQsaBdViVaoaq/DQBc8uOrToLfqFoY0Dhmivh
QpnV1ZP/Axh9SO5TjvS4ZmL5+HZ/F9meoJuLaKLxg0p6DYTnxxDruBy+MMpkGRF9yWUhKwY9x6qS
3yQIdkPefZRNjtUITl/EyMrtBvCr3aWzMtc/fd/bo45UFPIfuEUuTtUvL0c/SB/INkgJV66uAWLN
GRixnl+K/2vJfB6K0d64/wkO44jdLuNTErVtPwPtw9mvexSGK5ItVwBA2Z+NiJhmtfXuYiORQBdX
YMHvo3wwI3E6fcxRvNlN+SoseJ0P7m8obRXQuLcI7yj+3EafBy6d96twJHryiyO7hXE6AxdMpxK0
63VzCPHPic/dPMHNx+rBYPHoVMVwh7lZvwbgrO/Le9D5Vp1rm67Deplo0g1OplrSgZNtYPmHau/W
owifcTrXFEKOa/JG7cxn5ekvHwcuo3pojXK2S2n7rDEMbnrq/HADz86dqTRGqGzOwFS/DpUAkpet
NZOnXQ+o28ToB+8A398TmrIDf6lwvU2xSllRzIIQp7i9d8iePRqX+tGV5Tqg01CkXU5xX28ZzIoJ
nlI57Y5tbmLw9qKkT6K7WKyTuJmvNZz5xHbC4HNkql7+Crj2YJbq0UC97sIDzPoTdIF18Pn3X9NK
A+Y/utNzZZXQXjwmtMlj3m9W9df3gY9nFJB+fpy7ys7o8DytpcKHa3v7wISUMIQ/wC7Bm5IBvs6h
eq2RxmSyzBtJxk0cup+lP3tGoKqqsXeZYNxO9u4BovP7xgJ8hARKPSsTF1s5rgHiend9o31Hr3ML
Ej68bJqogurTZeMWFD7rosL8TnfN4U6g2OkLLBugi4ZXZ3fLSdQsoRftN3ITGzfZGfEU/N/lqUXA
CRpTzhewGweQ06HjXdVVcn/fwSxSPMOGo5a3RzHU9DDCC8JYDV4YpfWJg70pEnAZp3CdwP1Xecow
gTSwFajC5bceHSe9aTZSwj/GaugXvXytOkHtaGZc0BpNBHmyKcmKFrDOmeUtTRW0S9SQgNcMqJAP
jmR6ZMGuZq4N4CivJHbY7ydW62nc8q3Nlmw+Q28UxozbKWI9OiVBVy/TIDm59zjf7xXMNzilFLUL
OFHLKHYP1jdernvvF/XOpqxnlwqHS6bzpxobigv/6XO0qHXT6sjC3Dj1GlIXsJo42xGPxtOY5HiW
MYoj5xiuT33XW1UEOBQAjoCYyIUaQgQxM4cNU2wxLfrnGCgs/11W1maH891aQRR5pg9xVckwmv0i
w4xl0xAmgVQcwkBDgMphPIEClA1bU0YEtmGrGjzWQnYDoZ1AQJWWEevU+rZpCJGZi9FV77X0NFKs
zFxjOqoyk4/b0RayS0qUg3QEZzk7mA7W9t72GDRcIMmDkHMThx9KI1emUI3v+x40/Z214TiULgOL
TBjg3uyyD3rywWp9AtGZG6hVCZAJ0RFUalci7kIGZH2JxcKtwW8ZlJKBUZsgxwywOS78Yh7k0V/y
Du4YeJLT0AAIJo9WHVZ8EmkQGH8P6vBuHhgkDKl5M6gpCRjuhDfDmuHRu6U0UaIJxlhHxI1nMhwa
8j7K2jjcGvYxz9645GQZrPy1kva37F/IutQImvs4WxNbFwMV94nrZ5orRrcssg6cmO7YiuPPpZwP
9526Ocf2qPk5y6Lq/O+G0CKaljOPt/zH/LmgCxWQMYwa0hZJQt0DYlYmEyb/c8yGawdQbqaPQUA3
l9XWmewI0xNFgOy0mSDLUcRpOI9ldT6KxqFjC4xy26bDPb19YFuT66Ce08RR0O3r9EJGIlwSzyQD
0ZjhGNsx0Iyda5n8nA1FhVYOf7bk345PKo/XLHQTeIQN/KGQoUvKsJecdx2aO4uEDgd/YuDeWxP8
KIiu2O3tLEJ2KjUcS99R03b/co0LSMDQFxnTCeuyjR4VQduAlJrVFkgcUlkRTFpGLv0Uoxvc9lAu
Qofnem7O5wSjXOK9LVHVhfVlaa7U79RUyO5sNLO8rN/+DzWKe7AgRKmVk9EfhtPucIMwK4s7KL9U
ltdj6aBzoQRg0f0948d24udqFgc6NahrqLjlBdan2FsOCxQAuEhVbW0EF+xdij+b58Zqf1nVs1sx
h+81yLWFSB4/kX8PisS8z9QJ2SvT0keLTwm0g12A1lNJjctciK997c0JO1X8Iog8Fm4pKyprAjqE
3jL14ZOuLIv/Qnb+UYYXslqSvOUIWJOanQv8Ty53iyjZ6KnDDan1dQMy8EvaVoCgthU2p7uJPKDn
tyRQUP688cVQ/ttsqTXeQYXbsLr5iOBvrlcTsmv9WZIFl7b3sggkjtyiXhU8U7Ptke6xdtKXCEUJ
2QtzCUe6XEJI5+YVq+QZz4zB95bUH3lSt9lKzqvYfeESV4x8tF+evZBCOLWDK6G+2FaDTmVzDVuA
6b4qohOY2Tv8t1B8y2+2BYk+NpUQqiQ4MktxWs9WgjCxAFf/eiZ7WWECe3khV/qnCKYuXhor/7k/
FS4gsZQgUdosVJP16+EHuTUAMjZYdWBoazKv9MJbbEYoZDKVLdjsH4fE2FsYWXu8t6VcZfaYaMK/
cieQsIqVWmCg4q4qnqjWGYGmD/IDRLPj6xWWv/Br0tqq1L7W/xRcCfHkCTk4vG0OFzd9vvQqmdk+
mH1Lf7vagEy/vNbfos+M8SuroEQiERJoXvcs2fAwaaY3F+YMRo7yKc5yPLR2KKyejkGIETcZtPKX
vsrq+Ezw2RZ3QBDKPlFjet6RSkfD7NdkxYVQkELKXmhXH8fffdQUWQ9ytiOLGx+ZCFgfaioaiTrD
V1kT+SI0xBaLQnX3gAC6kQg6UM9RGKUOmynYmHzjQuCR1Kpoq1nfPj7DvhhuZU0LLI27Jwlbx1yW
Uw2b3avTbTlpcHx++yE3w4VJpdxzm8+aKn7bleVbQGAbmWAKaM04RuANWPdoTesHKU+0viaacign
eP8FHcgKL48AqzlaR/608CpWOpDRVlRydVo3+JS8qyi4/LyYd/sC4/M0t0Xix8n35Ouum84yDfA6
qrcMdxiH0e5iLLKpiYMdXoI+95/cBd/YaW9PlgmoGvnvIV6FOL3dmd0mTbjVgM4NDw4VuEfXLjLZ
0FbwEfL52qCQmMsAOv4LgB/618wAmh+ilfUMeSiC1M8dF+sCozN+NDvAewC+sRJ6RlhZu+D03xgz
2SP/VB5ACkNJvbThKmKLI+cj67rslqFuiN+IDVZIunIs4H4Qi/ZfpY95+YO9nsiJl3bazHAlVJF+
3sC0/OxbXTRn3drlAD8gWZbtGM2E06QGC4/xarqk9LxPZp9bDHkRahNUGd6ADXi3AmhtXgc+KYdZ
3GKp/NB2vas6cSfe7kNRWQk0LMB6SWbgKjiu0BVb4wH8N+O/SZv9khor3pyqv8APEOOnbet/s3Oe
iTwD6+1Ohw7+rJGyo1QC4PJ9vvrNvd86uOEMF/VxtMAjLyfQAiKVLQJPS4uzaoCqcXL0b4aCnn9M
jGXfAmGXuz2MHUxp7iGMjdIS1H186e/e7KeDciYEj2Y0LJVb1fQ1l9n/w8HsNvKufxpQ6hoiYwFa
In6CQr6FzBmM+/rDvgBMB56PhKs6WXiHxTOMm8v44enZHpbKa6zDuht4yQIHityM7gJ+L6EtecMt
RCJ1OJttCxCROL7ua6V2bAjXYoaOhk9yTk+X8zP0Vt45kFhKwyRZPjaY0up0dRsroimg+77Xgoav
BAB1OgTXg9dGhDR5iDMNPTscl2hwNSzwfiCUMbOhpabk3mSBixqsMZnFPE1aIA99U34QRvGfns/P
zO5xO6rmomMJJcmVYAqpve6Y82qVQ7g9915RJaoAlvCmJ7g7/ZJahGYmDacYnRIRf+sBpHSqgNl/
nYJdz4ZHeiIoeWx+Erbs7KGZhobj/Y+jZd4EmDpjPxohdA30kLUzGSuFTnLduG3LkrAKY62eHo01
0JnzoFAn9NLN59CsRcy15DPpGYqtWnsyeD1GQGhZlnCHbQE2lHXe2CMt1R99kqo7haYJMrFQL/my
PJwklMfDTnV6LboZ0W2+/JGr+/Pa+uPCk7tX1VKIWVCJze1B1ldfTSNjBYtTbENfXy/7c1XXKCyO
YW0ixhcd7s0+AQLPppkFbdd+gBsukdSkmZAhfxHEnhTWRoENQ3ZxWPOBL9RMRaeKIUP2CWPab1Ri
CCRqrs4gOe/Hw7zEhMt6oOwEMpOmbUcfvWDjOBEMiQ5BUJkk093gsCuHBdA48dNOwqDctdkJwq1/
enby8auVpOsDZxS8MNTkoinRspEcE4oIN6wol7nJpxFUhfULA0wFwsZQN//8+f0pOUngaf1RuLlR
1jC81eIjMO7b4RNP0nLA8C2vfR+4Oo0pHVrgkAkjGW9/KGLNxpOYbdIMf6itkac3cXVZps8NNyRS
hwngbr9T/3eRPes+Ouou6OEYuKrGWlEZbCJmz7sbPHbcGsWDITJNQllR2mbjMrWUfNMNx+vUS3d9
xsg8JihOSn/5e2+/uxFU6WcDiDc8iARGh4q4QiYOiG04lAN5T+EgsMeTIdy8Sm1OQ3+gcOhTeowc
0vf3KAwsJiWZpayagVvdCqsStPLqOkseA6pyRy49EpUoswubcPmQu64/WMzBMfwORwWqmIwQuv4y
PO+7plHnkaSapoC0cTwZ3/mwLRofT3napIKGw1WI8EnxfB1gD2L4yn0DKLeDuAZxOLYMRGkRHBwa
DO5pHq7gMrIf3h3HXDOkoJBG2L8ij10q+MWVkyanbrmsCpjH68KPwNVgvqBKTJtr03uvwDflzJWp
4tjsMt+2L/uvYH49NxmJ0ihxbBRSTFYE8PA9yCUFiE2kBFdV+eUrvcrFwi4T4RLPDDqf0TxyKS6T
+hMo92pIK3BKTV5JEksnbatAslug5Ov2b7Q8/OkMD5IEVw8jJxJZpDxssKhbmE+/ZD7YAkwlHH7/
neBG1pbzQR4tQtrzA4/0Uhy3y8hCHRrLIovncgfYv65L9HhksYCwYspB5swIVebf/O4vYt8YY8hI
FEqlHdMwQ9hxyPhbWkGKHeyRTD9Jvelw/ke42aqK71nrso+scOdWXDqF+jK7lGHvgKTwo55QHnRv
5EuU1CE2vwGfzCRq/Ng1N2F34X/jrsN440qNmNqpLdzRVDF/lzFo0CpxxKyPVr5Q8OvWFUmrzCK+
Ixnjbp7PTRhb3HuwyDQcycYpeicP0C3BxVmZYDQsSu0MyF3pA8HIrw845QOLp98ZaFGgEClfiF1q
w6JMVxUInm+WEGE5SquoWUA4ADY3ReXTZO7CMa64Y3A0C5+9xp8+WBNv9r1kKfN3sPDx3uLeZUJn
G2I1FaVfrp5htUTRFWO1cl95BDoZuUR7UrWGtMriReiMg3Ro4uzU7RjuPBeTw+yU+m2OlVunFhZR
Np+qnGW57y+mAoPJv1z+teoI1rIPnVZuttWkySCog/0gCx/LbXRnFzNL6T2/bJ+OTOneIee2CEsF
SB8tRApdAAMVvPXMYk+YEvkARqOaPqrAjBs4ktBP1mYnRr2GkDwGBX/HYovX0TuDj01ejCPcI2mq
4HHW6xmWOHA90G4i7TaLqgWy6hxD59S8UTu11DMTYP9ZR8MuVTp1+EjR6V/bULtEV/y2Dbsyfx6Y
e/hcJr6WE2wz9Zzg3mEHyLQUuQJCmwsspnodU/BdpMXYK3eu4pitluN5otoWwgrFPM6g6rIvfSOg
iaZJJKxPMRGd2nqGnXa2jCNTum4B1Er8QEjmyZowbziSoc3OhAcvQiLKk17t8c0yXR2vgNPscrUI
RTNZf66Rb7uNeRUbxWrmQsB/jLM3sOmKHGER1YpV5rg96Cviqtp+2se2PljjvsGQfQlrA3u6UkhP
eGcO24w8XbQ/m+72lPsLfcUFDy7OHUbdN4yUugzQyRihS7vYOfSUp9gjv0lQXWFTWYctbU9bnlYT
k/QSegog7QK+1KunBC/Ozx6zHqg0YuaDMbe+l13XUJm63lPlyXJ+RZXLnb1FVKY9ER46JQzxW6IY
Y6iSxkaWrIqG/jMr/2j0jZ4nqupw6VnWbcqVS9EI4NHXxsTtI06DVWW5aL+lFk/yCFnVMPAA98lP
5bUm7jZ2E5EGDzpnl9pQE8rAm2LMWFv6DsTG6JBDrx5Oo0XW9N/3zCkBVgmWqdNWqvKwFyXH088v
TkkG7Uh4UeMxZey6JPG9i/YB99RaMFh2uG6HSbm5F27IKI2gsxMO+U4dpm2+cx6zFlq+hNFU3lMZ
UYHAbyBpYILcsQPx4xW1mkYaQ1citVwKcx2g44z0VJM2MvBhWhmvTyNPd6CpHoRZIB+fB/GKq8tk
ZDhmfZ3rktUymZ3P0/a+h/mAgmABmmCmpffxy0BtraM6sMR7EbEIuLpr9TVnrcGrtEuaP92oGcnL
Y1/7aeBY6zSh5ymn+TmNGsy7QzpUKiLBm9NamS1YEFIPH9449iKR2OX7V2FHBr4QGKXkVACcEeKO
Kv65/SMTwrfI6zfBnaOfvz5vN53vpN66k4Tdvh6IUNqb08vlWFE1GVNyihtoz4oMc8UXoh8avk3S
oS/FPuQ+t4D0yPmPXdxGds9/JeWj80F/+yKi/I1hoVfzocnGNJsjU2ca7GDcRXQoO8UpQReyrSSh
kVuxJeBf0Tnc3x01VzV0WToP5NZPHsJk6P7fgYsbyjS7DrsGAw52c8MZwHRvoGEtEInoSUb7iqFt
6BCXJKk60V6RFKIQtOG5Xs973GJMPX6SzbScvEYayDRa6xnufeNIKJqwcc8fJFOGIxkT6Qa6c9nY
Db/IdtT18tyQTwsg3YOg6j0fxHhnvQjkGBsFS9Yjs95HdpwqoKyI3GOHXTWwpro39SfPpBYVaFaZ
WyLS0n0vhu3eLO7tb/zKq8E6xc7KjCZqCEAyS5fYBlw1QBBU/fZF4WurwMaJcMbm1AhN2Kh4wSxy
SXhr5c31NmpEFPadxe04iwhPA64SdfvRSjPa6pjHPI/1fru7YlEuAznkdHZ2+AQQcPq51hiFXfg+
2r66lHoWjinPdyF/QI8JUP82Iu1Vs60UaCt5BxFf2YEcWwcutQmSKgeoqaiu3dMP9dVuuvE2180r
Sd3ONzydxyG8uFCfSfNH+r7zWDfbKExfrBzXPiIoAG9uu5EFgNBwkyzZSrtE3zZX7JWNIQnEJ3rv
4KSo9gx3QlRAI+QUZpI2jvp3aWnEwdSGxHV7+DF6ZhW1UXI6Rdpcrmrsbajag8zAMWIwwGr3iWIL
mWqizJkEoqgd6bRL9N3drShZo9bj8ct117p1SqkFE7vIkmIevptkSScsmnvt+zIqLFyKQRZLEqn+
OVGlqkYs8wruCJxRa6zshGNoQfvn2KfE8tiTSURXi6Dtgs7FUQIr8qijDEghiwOvyekvCvCQ7c8+
EOqH56jObQgtD/LdI23kyYnheY9Ak0cL1H9An9ByppnVLvznSgN+2N5kR32H7WUvQrZsJuZT3Y6N
g/lB4Q2A/KHiKy7JKOxYcx+vnGOlpCbPKvN7MLw4F9Y3KrhVV8n1cFo3spLdQ9X0zyHSzOCpxK7e
6qVwy5LMEHKjWSCz4dC5n3HDNir7TB2geCY237kUM1uWF5W3pDs9huvESUFJQJ+ZuKVWIR5LCOFM
B7oWHxkUDvBbxZAsyK7FjePLQhZAr0d0ptujw0qPbAt8/ZzWf825YxrpiMW4ebQ5a/PY2Gvx5u/u
nM9bjrxK+jYNUeOowsmEMND03UmgW0+a/nwakl9WDf+MlREtMUJrnQ2zNMot4u60doterfBR/b+p
d/WJzXJWHVcBbGrI2pRkZyMhZsbjO4lAMYWraZi2ge6UzpNXtdwgVnpADRwbfsIQVr4Wy1P1SVRI
Voxq5CzPcwokg1c29j6fl8tL+j8ri8LhSt9S3c+79+6Er84Eh+mOxZS/1KfRLbSAp2omqISdU1aG
hrjhSX5A6fO8GL8C3IYQvseEjO3i1kQmkZKSrSslJcWFiSEPRDFFAmdPN5Mj0mu/cQbPfyLtlyh2
JXbkXhectgL5dTmigRoPUfQqHgSu8Z3P4Fd8u04WB7M4OXy8VHhzD0+ho8kMd6i7VXNUoV60XEzX
sOc3YH/XvsK7iQfLkvGYSPzl71ICc1Bz2enfEACN4zo6/ofz030I+w0bjQWJYR6SkSe9X/s2Wqv+
SNEavhgTvDuZLGk4yGfy6kpsNGgnFqlFh0gf8mwXbaRXSSmoCIO0jDY/vTuwmyLC0xpg7CzzESJh
gcIQfOCrv2b7r249A963W1eHqgBc+Pw/Un6thfr7oBC6dEX6tgVyBmYT11cGLw4fwhghV9WldDRp
+SCoSn9PML3gB3Kk0kunLrleG+7fOosJ28L4lOaFE4MA4TxyXReXcLZ3IWCBpDUSIFaQuC4yi/h5
nFwF2z7TNryaX7dn7bPcjCJJtZKxuu4GwjljCxKwo4tnD1nospZm5cgYfFufzofZPN1Q/r/rVXzJ
2LngJXw5nkW3jpU/1HLtvKD2jGwJEESeOD3/DYI2xchglltzV/ERmhleIETo59EeZ4XL8pSIpdTg
XB/b+dO5MSU1lXoBlDRANT1omb7075rCP5M0iFu1alQRstjG2jxfaiE1MMyYq157SpToVI+CiGs0
8wvcauFdyg5Yr8JJh+hkOgwQMXJRO00gZvrOnF7OYK9Z+pSTv9nHyElmqCDqYVed/hc4qhDumR78
KIvKWmVWcqjyGfBcq0EeWkwtjQhjRI8QfWidYEKheY+ocWbt/VVrD7qtSRQrZ1bgGPX5iRFEBaJ7
gjkcAixxF07l2ePJziCC/GL0cJcA66LWcGCaBg3GrBvWiadbgA6urQzdkl2RewQbGts01HBvzTO4
E4OGVZbk32FynEQwblDEzusDW6eEH6vGm0Prxkr+17s1Lxi1/3JJ/MN/fmLIo5KYPH7Obr2xeRlD
jpmGu0XAGH/eCY6qXc7ApXLK/mzUrxVuzNKcHM/SNH5OFv9iQyoav+E6bDYkxHywgCF9QAS8SfP9
wgs/2u2VoMuZT/0cAtDsT0FI8I6621zpHdvAHkUCCiFXlduylAJVGRR0TbavA8THUCgSQleDHSn9
Ylcxwd6QH+8CBTwKd38A2eDcGUuV4m8aGx7B8q4ocy/3P0TVzM97OYvPjsRCnt5jeqj2iUviRhHG
s/lCwrJRBxVzQEXDliMCZ1/vldhimLpcA7DuWhPX8zimZWbXEVH2JxjMEOQwcKen7NXahbMw4MZ9
vLUK0flwhNJq2TPsGi/oEua22sN895uET+m22UeSC0FCGbuZ12BmeUsaiY37G7tmqsct9aHV/sTA
7TU3Y33e4F9oBdpQ6LPslZnlK/XJwZy1vnIgNmNBoAK25kPJBe7/3KxmezuVFTavK97sWh88XtrU
TdwFN7df+Qi9JR1Eb7vdah+E2vn0G/jmJ/0p4uZu9Zn0JbB0rIDUBsHsID40CioyZdKLtIjsIhZ0
crLak6vEE+7WHKTLaq/+9rW8xlre+aVt0dOS8+HhYT9XskcvOF2nDChpilYbSm1dpSvW043CbT+W
W653CkjX9BgcdcHSeQWQY9Ew6XaDlhjH+U2pgyEmJKG3b3banMxmc8j0WTStqmeRnVJMu8WybhN7
jkIpRDN5YZZHPMG3l/VQl4+k1uaA+7e/Q0zc6vbQzOqfLE1oRFzJ9yKbXa+K956p0Glxt3V6UBUB
xMIL05fbLYjaTqHB1v7HhTqA//wH7sZ5ANcqDM+RQZglXobJAd7lfkJHOeBQqvjoetyoNxRynBBU
WreAjpfcJS60BVwtYWWBvqPgVKhYNbt9JCE+8JYalCsg5EhSHwtQf8NGgi8vKHXWGvtaFupkdvFo
T/jeNgMWgfrZiQM7nDEHr7wpiGdlnaoP81WcFpkVJAcqs3HzBDlUbrcbVePOcLtK+4gtMvhZHMwl
2Y1d3oORt3+r+x9e8neCyzzcwVAOGTHFIRJtcKU4OrzHbdmwOCOH4P3OrwtxPoX1QsdvEmXSsomQ
NpD7py9T8QAJunN/UMRA6ZvDOkmEtojS+ZvA0/6mgsTBkwb20s9m5OaCa6dt+lsJXXRFKTBbqqba
rG66MtiRDpSunK5MmGk3zLa3iTrTNLts3sOpwux83voOoNn1j2/B29rQpvdn7bLaNM412kFDSuyB
oUFrMZbMqknPHFhCgYsd5ihMUD4zRuxiIBAJJBRr20i3A1yzdv9RJTKD+QDOh7Liy1PuPrxgSNck
7MTpHU/ScilOdafF7uSX7OfMOZW4/858Pc1cxtUkjiBV2TqUAv/JgJy7MgpXGqzLyOgDB4yOxnc/
4+gNGYNdGtd/N1wavwFMicae732OpHhO32zwokcFQNTOoKUs6TLuRabDATiBIUwznRqxV0yrfxha
jSZWAj77lfjKOvdPIIdftpDqb7cj3gBzzFQaE2jg4VXYumjGiBvdUUvd0XA1SkFnctsfowtJ6Szm
FjvgG8s6Xr33tIhvv/gpje722LyyfH68Fibkjo1O6m5KwD3HhQgaWkGOKIv00FcU3iCWHAyF4WHQ
q4xzHm1ueBIJIm8eXXKCl9i7SAY27khOyiAwdkUHNgjtignBsJLaLnd3OvRBR4d1rmrOoXe6VviB
yWBWexiYXnXsdI1Kns3auS5bJCYm8o+l34u7cwQK17h0aGR+0fo/KcMwopk9+c+3Be6jaOeGvhCk
haBl5LRIbz2zVEqpcizp5zATwPGqf6mSf3qycC+nmPhKNwxq3rCommc46njzfJgnSr2Evy44G3PL
84ZzWVyZqOO/fWHxGlEPapjoAtuaPZU5GzcZd2NRwEOGn+wzSZDl7Dk9mH4LK45LKyyDOkm+Apyk
BvSzjw1+u8tr2y/LLuJAtQnsIxjnqikB6W379+2y2QgkDTQGzw89rfusLp43g5aKQgnTCxP8F5+d
4DbmgUjqSNZyXBem3ac/ISKeyo0lHo2NA8hVQUXyLYdO+EQ2cfHg8akmZMfjl8Z8TA/CNmmFDrgJ
HUOoO5cEv2VIdXirM62/RU01exMj9i1zb8xgc2jQlTBRVCOJx+P9UgBgtk+4z2+bkQaF9JHIdZJM
0ijng8jmR+bs8HDVILb9/Kp93HbRnfTZPFmM3MR3hO1sbw2OJPrqLtL3ccuLqoAJCKJ+tvOoFYOx
qnwN+fml3XPM1OIizHVRNDNZfD9ENZ3PdLuasHQSDyggwlDsCJp0PvAA6f1sIedxn7OVDATuq+Iy
WyrsBe1AwVqMfNdhuZ0AWLwn264apVQSIzK9ogQATqHwDI0eH81aNhNEfWW66Edp5ERqnrEZPvCB
KA0qowgJ35Nhtuf1V+Rn9bXBS5viohMAP2O0otlIWUDnSRS4Mm9MVh9isBBdeqkgj9nOvmxxFWfr
npFDocj3pAknx3QYL91L4NQ+VQrolHJU6IJQAqX8zI+GsObIIuWtvFd+9jtaUrhUEkqm+a/SVe2G
OeZVijSmM4cJayRoALGT9Gxgxj2IIWZLUE8NoNWJGnUabMgXS7YvLwWNOMrU4jU+9e9GSMHG6pfh
U5pRS1wU/iNmM/kic8thaJbZjBvRMp916ghOZZ846+A3Fd7bBAV5QgbvoKe1gdrP4koRCMs+GDgo
zCuFsZW6w8RqpolvlgUwkFHbEpZRg3t9YAHNtiBQy/lChle/HOUkLNDmgi4SkdUFH+qPBusdfYWj
u45zY4kkJAIin8psda3BYtW8hBO+7mjak9DPoL4QXGkkDaFNuDdh0feriugtpLLtVRJzJStBI6T7
9/Y+H3iaW9kVA350LV4ivsCddCWCvrCotXCps7z95ch7idNubrmbhJWDv3aDOamb8ebsqQzrkwbe
Pp5F/hE2QG0ZP9D1GshWBZTiIKick2stY2oqkeCdGx93OtlKhou01DrEG0o3qqdO/VvZex31Yk9f
YCD7HWXfpGa2Mmg6BVRFiarTUjhp+9oK4zTEJTVB+N38cWWqjN87TnAS6AAL/F8/o31YcURPiqUy
0btncp6VYRw5mJDLglqkIk2hH4BoSuiNnE5fZG+76zHZY9bS4dENs8FmdD8oydHf5YZa/gqvIY/E
wjIpuG86eUCzy5mbtJpsY6G2oaROpSlKkrWaynpaUTx3Nk8GvrlV+iD+m07daaPIpByfaPmw1Q1e
xMacO5Dnn4prNB2mK6XXFo/fpAPUP1rcZMFg0LdX4qYbxtSI8uEUx95JzxIGHtPS7iG2PcXw5YUf
8sVLqLduDhOVqxvQmKHyPd/9c8DD4q+5X3HTnROVa90v9h4X2idfbEO1kmEUFj0dF7592lXOdzne
1wkf4wOddCe92Kk1YpQmXDwfjDhMWM95IBh/0z0eJ3J13PaJJLf6WZwLOa30KPkseP9dgHnQwAMl
JjQtgXmEb0RBTKk3BaOSwTu7RvLV6yZrNglwrn6C3HjCAdbZCaNfskNf1GTqPVmDUO0Kp3rdqEdA
GwESNkeQaqr1K3tKhbUGttikXZLr8OnuJT5leQOadJFHipOp5fFZJw1CQ5MNZp8/NBdknS5enF62
D8wKFxUZ3ZywSpR19qgspkHUVjOa9zGnZq3Fm6DWctQ2UfqBrhmV83FEH1zWY6Z0x4D2OGl12GuO
zeO0daO8mj77Og8DEuZPH75ttDinwqmZSPNBMvtkRKosUt2AFF61recmkRIejtldyoMN6UFhcdSq
IuoxzxvPq1peqcVJ2K/usZ4cUpt57wSgjIDpT8V2cKeLix5IDnil0E4lpmMGTzyudvesgTnp4ds7
qy6WXQmkj6LL8BjALtN/kH0kTI32RYvablm4yExwIk4u9vd0eDkyYyRSVAdkkx3xQ34+pdO22M4P
t9jGMFaFnf/8+x8bCf5FvyIdAsYPkTS8IPqQYRoiCxgksmCsyPZ6Hpj90Mupwj07ATeCYZuGLCbs
E2NbCEnIcpxNZ7LksnRBKbv7GJ1aE1cHlZ4jWV8Nxg7Xv3cQpE7oCvQJRFjVkNA1m82lS8QYiX5W
FwamFrRScuW0kGMrcHObhuqTx0cuV+8fQ6/Gt6AWe/Idusgv5uf5WOIa8tZhNOWKdyW5c8evIgzq
m55YX3UQW5U1G8L/V+Qhs6actz9Yemra13iPUOoVTDovKHwDtqkg7dhxq3mWPnwx8lyPCzDrLzqu
IA4p8Q3CQ9avPoEqh7NsOOcZfEssgNt9HpRjLtqjozKM8LJ+hmcgI4x6OnehQ2RqpfZ1NcJqdXZp
0yD0TuRrO7+21JMpnaRRIYVRoXJ5mmVmt0127Y2ijGbg/FIHtAsPETyc3TH+j1iPIq7gLIn6YbDp
kSxqd4Ch1gb9Mi+RQ1tLa383LOKYLeU/EzLbZiue6c5Z16DXtBXPRvk+KMApMl1kRNlUDB+stcNa
JOGlRlU/vouDyx1DVkZ/dx1ASjIwmckXw8EG/qZctkdlvHhkQGJO7FOg9GDARPSH3086ru43q4go
p9GIvKEPpsHuePO8J/RjraZSTUHp2ruMsnyqfgatYbhkGIxxdnmnpPtbKYzzFTMCbdSkyaiM+b4m
Mf9iZQ3tA9H9GaNekKfc4Chz/4011Yg4RM/THJ1djB7xCU5KsLO6lkMwffOYxY5kRvG3DZw5Cw/h
GqU0HYl59FkfX3boJ7lmyudNeYHWxp32wlx8ohq/G2XslzjJbXIeAetG7zvc9zJeeq5yNuzHjIA+
/IUDyxiiWWSP9Z2k8FjCWDML50KiQJAdVDaqjWVHZR7KJHEsWtlk8j828J2frwphvNIYZXRWlyVk
UoEaRvcwtI3dan5jXBZNZSAlr3lkVoQYcPi22DbzQVeVw3mS1qBpBo5hN+JEk/SiTcdKxSLik0U4
TJCf2D+xa+8xjoNnByXWIHbCWkDPBBBBfQ5s6+7nAo4/dodPbzGweR0xQaqaVBfTALshmlCmyqnr
UTwCa/i6aUa+HPbSx/5bZuy+6LcFSycVsW97V8DOXGSMQHMmuOOhZgnwLWPPC0bVY8VdyDywJsGT
Cy1MK9Md3pt6AS04gkn3mgbEJKOhWnhZZObkrmcjwvO3yuJ2sSvBmlfvvTLBJY7LXsikD0rT8br0
H996cA9dRl1R+wwJicaULvwDJyvKzVsiMTTayFrsM8cuQITaoYT0w3CuNrI5JPLX3T92zqLq1tNG
y1bzEfkDD6cBfiIplg0vVZv3E2EenvacmT5pr+CT1nV8CXMaj764L+WfcF4w18Zm7ZF7YaAuVa76
MhwrLO4RK+sjzbPePN7+m4WyrwAR3glISFz/MUoyrTbtQfaKm3VXDvqSLlas7uCzYGYCCjdTRNcB
5t301YPtZZ+c8+1q7vws3ZKUe6iUp57HWSXM+IMWd7axkOffQZhaDq9L3xZkx/wVNUMJJkTDTFgU
GIGpwTyfWb2ZEsE5TI286O6mdzLIN7b/ANypl9Q6qBe8rFKtdjKM+KpTKM2vWcvBVCAnMHSNRLU+
OVPBiytuY5Gck/wmxMmLUM3I+Ev5kd0X/EAu36woLRQKEp58Pm22dYesOUvH6I4YC0jlgWhfu5Lh
7tkSKhmTrhRKeLAugJq+IUp1qEDUjJvJGfa5ru7/GpyBmZu4+n8/5v0rM8ebz7jeTuENQxp2ZyEh
RwDVd9ZEnUZgTGioqJVbB/oiUjUdkcaF17rS1SjjRJJ3F+uWEcTrfmLjgMCxnDbb0YpSpjBIREz7
/HY9sC4pmKWQbg+8a5/JwFQdI2//G7xGQZuYzk7ii9SASgFhWKMHDwnJmt2BAxKeea4wu5ICfnkh
JCt/FmHtgfifdS3lF51PxzNPD41tECsHLf/q9RENpJn4z32Gc5YhELNf5ATpY+6hLRB8YPLiVSUq
j/YwRue6nEN0L36twURn9E4J2WXiqWWDDPlax6AK22bDrdbTRunL9hrgrXnQ4yjpU5n9r/6hSGIx
pieVa1D5y2ILlPIvLISEJEo6XslqVt5FNU9TcUx4knvOK9Wy4OMz1SE48J8QX5sqboGZqtrOCguT
j+g8podZ4rUXn4Q7/yH4tlZrmgq66ENzZ2Ix1cJTDtMMvgA2QuOHxaiEkkaND1bb6Y7W5f7/BLIa
oBC6WN0VMwJCN2JPbs9vTThoYOxRkO588TSoGHcAOKEDeeAaC5vwDuLJFVyt7e3INxcUVm9und3f
gj/v1EuryPbuehkXAXNmgHOnUkSlQUgslIHRCdDIHCvqpIcqdX7ipsC0tqbtviP2MXRwYMez7C9a
2NHXiGNwQxq70uoqGFnGlvdar4br+i+qRyY01cCYIQVoRN2ZkzJuDH8l+Tk3PJw6ozOd1LeR2k+C
bJQpi0/NabvmaDBCNdhxMnRHonCuLKyfP8BqQ5/HTaXiAIcyQrLEu6X9kY+WPY34gO8jXEpvZ6WI
1JYqkaU3OFlvjc8vmT9iU1qFQ8/r3IqDiyCSGizyQ/vQaSSKb8d0K+ar/Tdxg8Gr8w//sqzl4+za
Ag5QGB4JntogoZfMa6VtvnJ+SOgYBESLtLV7FDQ6wcQhD0opFtz2aZA8h8U8MK1UzBpG4H94uDm/
RcV78voq39yjFanNLZdLm5ybnm05wNT1WJZMd+4e2oCTlcwJ/oSt+dU4a+1V9J50zarJyIUJ1r3o
UT4OHOpUAoCTvQfdHrA5Wzb0diEheckIJzn8Zw26c5tTkPGf8jxsyp/uZz+ZnsQj/JTtBWjmIAwZ
lV+wzVtTtU3WjTb2G1MueCakdCPMYKd/kluR1+IPLYT7wqV5pI3wv3YG16D7t4MgY2qMioc0Ff8q
rAdNhSLgbdo4RCy6Jr782iGoWPBh4iSvBQ2kZZv9mGrUtM7EFtzZ7vuJDWUbYad7wIqYfnCIqp2b
oImIcfl3GTkeKmKi8RT1G5Ess1L6oJh9XMtJYPPx+n7yrYUk7e0URyZy893R0VMUAW0UNpksQGmv
NndRDTj+xvvgSZxQC+hj5Upaa/7/oUxVAWgk+MGce79NJIFdbIKR2xlIx20NJ+WpaDr/II9goI4x
wENaKq6U6Q9lw8OH3wda9t5sS9qo/PQG7PbguK1ZeCHCmzZ0nQavVH9PGKDY7er31XqC+BO5zbLt
U1oZ3kBg2oMKzYAta9CLnfaufZnfwz2jOxKaiywJk06TgT9QZ0MgB0kIGE995euNfgmACVvm7S6J
LJJBpqHfOu7X1i3xefSU0n+/Dt+fSJY9hdP9/8eRrKsTQV0UsQOCvR5Blo0Vzfpx8nPqosTcVGRm
EoV/SjlZn48OwxkjOXQupNsGJppITjtzTzM9o43Mnqq8VCMuW+7pxbsS87iDiMUozPaMlVw0ZotH
teP65/7m9uJktuva4+QHxufx4HusrGgXUHjcdQyFi86e8UoDkrZRO2jLaDi3+QDqWjCJgmoCPdww
8ZtuDHpkjZKlUhFTJZps2KPRZVQtfzvtuTZEIV7YpLGhH14wGd7+gTf+7KKG1OIIY6S9abESbNFO
02jqKA41ORBsuzZrgEo4Ecmvf6kie6Hr3K7TIo39830BADsQwFm+AbyX8vXBDFO98xcsM5C61ZOY
FZ1dNxGQGbVPJO86Rq9iyVXL3AVVwLBFD4ymXNTSxB0LR2dlGy+rzrHln8923CFrCYfL8fG3Zuom
xYc6+7G6XRAMM9xcqvkODd/ATJFeEMESCVU3ROyItza6iIh1ZNvEVKtlVGRV20F1MLRnslswmYYl
0MVLZs2qADZbT4iMD/DUKFKidiaqHKSlGBIdsI4bycxIBIm6tfJF30bWrsVJBBjIkIfdOTojTf52
6fEEuGYBIHVhzvHU0oC4TbnK1yq+JJdOW7oIQJXOOeJTyTK92t8/4TYclo2wL85bxnDSW9Ts5Tz7
UqrOLrxbLD2+efIY8NcpBgGAfZa7Z2TROqHrzpJ54xVU+Rj30S/2Pa5Wd+ftM8V7fhHCkrBybtM2
0qaDZGpG2Nqgr141oSAzHn1PsHCXEB1TLc/ax3dnffUNvkM/Bqm+oBxpUm3vnbu1jTvikjJqVyFQ
y7CGqJa0TX7R7S8aRv1Jz6EPxLzmbx0HtA9DJDViTE/1g1J3NSft49tcOzHKSakDs8osbwUAqVLy
Kcqh+NGX+rCV+X8jbyl6v+JmHtWW9/f8shb/CJlR1neCUrgQbMhcDYNnBRNZU5pAklO93FZVlxsa
BFBEO0Po/FjCWEFs/jwmW3YqKPUk3nAWr++FAxQC0lQv0UMXRBfx5VWA1cjlZBRmqs6AA66kK9R7
0DYVS1NMrWYNFPAfRG5fwOGkWTSY4BsPmVcdBFzSi08pimMSscJjqe11hHpq1PuC1a/U+DfgM2FX
XGSpX6XNRS1OP8P5S1HZ1XDblCWR1KQUutUWg3MAvx08rsLuER9YK8euTto81L0RUFKP5hipRTSZ
PYevp8nBB13t2s+AZzeKFIgDGNYW2L/RvxGZ24FIyT2rQIOm3qN7iE8t9P44B5u7g0V+xPCETqFv
gI9ou+pKMRzy4od7AN3Su8LumOoFvvb/JrJyGGcvm+ITtiEoCsM891HJ57+TLls7PtkO8W29hVH5
+unFXUmGqLWZYqlklCDmpIWn2KGwSMsemqY6elVbxqwD9lNY3H7lnwzE4oLXXI90PR/ee5N7n0gx
vkiwOXZVqCa/W2XDtir4RALypC6rGfHxqSjrwmQMcCH2C73J0gMF6yTmrEt4VmP/Nr7G6IkBr3VR
irqmPwqhutzXmkpZ3dxEsLlla38qm9R+5SsoyXuyK2aYeRqWrKettdoHjlIymD/swDH7bFr5Mb7t
y3FcZB32w6wSkhPLYotIgTW0gexZsaIIie/lfncPcDA80VwJfVJLelFFjkMDyGJGHjHo26oI8p2J
b2xlAkjCiAPZj74kEwyTsMMOvAMuL6A0nOS5W3b2/pFRj/YQalsZdjssYaAOoyFjMUWbFensy0kL
2bcKNh7MMv/Zd9T1j9jCU06asafK4bLP32qBvbniqeImZBlTr8y2xL2isAbGYjgk/z/udZhB3VAi
nl2M8BFN9WNVCzMARFjMSUAJwyq8wQhdkR97hGCdBnSTHujAe6M7oHtdAsyQEE3oBwga5ElhcrKC
4ftomyfaBBgzfLtGgJRCvVe3rIzRhWXftFRKk83/oqr1rPs8VtDkBavP7yCtKDJ/lPS1egEsGcnI
THJg9Y+JDsC38nujpsRQ6EhTQv+6afpGIjCHikfnlY/weWxsmy2B41Rv1dndnuxwxNSoMKi+xoCD
zyRzf3lJSRCDQxAW1yFks1JFl0x+CSOOb+UcSgLLxudnX/fJdmTDt6VjmkIymw0Hn2yUtwZ8c/Iy
uMTRzN525Zpd+T1NQM8Rr0vn74CMzt384cryUUQXWTh8Cce8h7sMgZZg4MDaRW2rBeKujbLp4kl/
9fuIIrBmmBCEuLu7RAvtpQXLqYTh44qORJ92jLA52mTrc2cmwj5BTLZZHLY7WzS33A+TcRs6va20
hQiQ7vnkSaCTm+Fhdl7EhPOhEjWGo2ZdPJfQM0Jdz2DKcgqpG5okJcsTLEO8EQu2giWFtC8hK/wz
tOw2Fk+usXXshNRVlvldgkICDuAf8NI62hyr2aGJFdl//Vu9Pi5amwtiSMbnm5Ot2USU9910/D5s
rALGmNQEHiAdyiKjddWQfTy6jbcGHBnimLJBv/2RIJz9ujjxfAR0uXWxpWhC7sYNIWXuAsvMtn3G
OwL92xXOWcQuq0SwbvY07yvXu4qaQYKBXelqaKuknweT5VQnw4fCkeVYDmGdkk+L8/lOe8VAQ/5c
LYUrD0mXY3OPoeHia2wK7O9GCWECiRo8iIlJkEn/k05yoMQAxafxjRiytkzfYqAEGIptm84YpP8U
SvLkm82JKLS0m3ZHtHKMT9kn7CDnCOq0Ezz2GGyJKHaezbC/vCd6+p0d3B73vxaZyAkasi/5uCAm
yN4ij3IldDEAOSSHnXRFMkYK4HRh2dWn7KAs8vn6biNHz19N3vVUFJp1FrnruPW4N28L7AQYn/mG
UHXc0ZvbjnYbyBZpIJwlMeQaq3GLcONMB+8tVvbELKg5u5UOYB4/XKJ2hG/L5aEh6Csh80dT0/Lm
GObOQlkQebc1XI3nKE7Xbv9wDBqLYt1GTSDAoqOkH8OmZ0q2bafMBuu4kzhuf6n6HE6gBUcWWiQa
hj6gSnE+YE2MrA/b7EjfooE72OW7m5rxknpwJXPf63ozg6E9Snana5wNOZ2mzvZmKEbb2Qvf65+J
jikDr1rpjRQmd23I+C4YYQS5WWb/2Ot0UInnDi3bhqk4ysDIAz/UL4rex2Oe4ZZved4HFG9Y1C6a
4U7HWgg9lW1LO3Uk3cqxadJv5LQpjcPEfURmwuyGbhDGnHKSaK2uWFO4jIVvNKHQkg0nVz0Bo0/6
i4BhGICOqelEE3ndIl57LKIi1ceDQqZCXW9KNiMul+5Bo/GiiCeL8kSkr0MKH0S905GhFzR4OAvM
UVXG28TP3Ehpw65nkFdlSHg/FR8U2hfhAT7kQim960GNx/38xHh79zWIjxqErcpr5tdapdEe0Z8S
QRSJMS8gbQzMZP4ktmcDV/Mvk/d3dtGbBeDaSz6I4eK3FASouLSugxKZkbUw0SsGSbsE5Zyb1glG
aZ68YrIDtQ7fLFYXrbmHYb83oCDfCv4oOMMNJysx/U0CXNKJcQGKHwkeGtIT9qk6TSN47dijCn/p
RPnq4irqWHzcnv5k62bl9Zx5fI4F7eZeQTUszv/b0Zvdn3efLATCFwK2UoSJqbWD05nsxfuu2tvW
RMlfGBiFqFXk/UWH94rk33v6AhPBUa4+f2mG/S54uGwQys2yVx241sYX8W8xHVwRf738DASMVD+X
AX1C27nu6jjkF25oNA4luucd/IdoXlKLAPIWoL2w1FEguCLw9zs/0gejOV/binrE6Lc4QV8d3QWf
yctO7kx3PpeEl4kRhVUL9L0y6Mm6lZytXBwBgL0xzg//BchWbkk4JC++fdLhV90KczMdOcVy0bIh
bftHlP0Y2ewLS5S4WSuyk9jiAcMZx5M2k63u00lvR259E1yc7nQjVbQ4H3rgJVgTgDjJ8zxye4Dy
7mIlAmOTn0Lf67nTUTj4RgLz+7ipwonaEI47cPeCyz1Z7cfJgCUzubkB0bUkqIP4TUCHo7my4Esv
p/Ma2F7MZhtrrZVcUrcYcjd0SPLPjJX8uYw3y+iCSVIKXQQrLBF7/c3XLRiqfvA7pP0FLsSErc52
F37R0oCc20j+qlnzrznT/BRm/MEvyMQAX/udea1vgobbzLmM+WnZeWG4vbBG5XjHyUOLyi0GWldj
DeqEtMI4AKElhMC1qkwkWg7maJjUFA4EmKbbet11Ca9pPQhXVqM7UO7fejK4e8kWH87BgbQxjBJ2
ZN788k4RQsr4xp//81xi6YSRGqUnULYTnoCCrH51YgEYg4LEm92183oBmeLLp0s2Fvv8KiQ0+ShE
aS5AUSbnp8aiIJ1hykUmEJWRq1ZWWged7SOq3NgJiO2PALF0/Loqeq/gkLqNiweaAynb0w3GJv8J
L5vKGsXYIkyCxTYQ/F4p4d+VqxeH0ub55KGBS9omutNg86o0AvhqH93w/kAqqyNCisdzdTZLyREE
38stgg3UxKdF+/Zg8IG/VCNE1VipnVB9z5fmPqPlDUD44QXqgoura2i3pUKTRCOBwm1u2gQn9Eyv
pODZ4mgYqqoTG1qCdhZS8OH/oesnpTc3z5JeMhjnIqt4S4g5cV8YAnXn3myZy+BFrd1YitxKtzJA
MZ4nCLDpAkroHaFctA4aDA/MQsFBjkYOHtAIQxd0kmze5Hu/H0Q/YEf9t/COxf6zDNhrQ6yTDOtI
XVoVxPPorTHmrkbgnPOGqjxwVrcfXxpbR+l0uIukTvOxcnEEvSJoOAok1h0x+oTnqcZxP0Pm+I87
jMmnDmv/o4v57VCo0JAq1SYGoQebmoxg4rLxHS+bUJnlMXDa/4ODzLKbCf7SuTyplhrUy5nGgdVD
Lj8yymwoLsh91egB0quQcNGnYQIwAwcLxxnjYInWJhRy6XRL6uTp1Jr2DST+iIMaoAmXvbP6b+a0
8rnWtM0v4VAkFj4pvTiKvHlnjUwDOCmIZu253Z4XJzJeF6BKi40rwB2E0tDxs6e5gt2yidX2D0xp
9StB6eDhhQAE47Rhz0yp85Imc/wBMJksYuq8rY5W+ZKZoqphMcUBPHMxMDPBPyBbNH3s5JERvHcO
JIyZJcFLcuCoCDsyuNGZsYXoGFHeF9Id2/yR2AqqLyMiF4QBGTv7L/lW0ha0s/peJgU3DVkNp7S7
sm+O/mUH5CqFtvjvzqDu6mppt5bK3vpoRlrQfmbqd8IAP7bwkpd19UVjJbKVleiyl4T1IL954nCL
g+hzzvqunF1MxUI75Vzc+MS+GvG+Q93cXsiaX706E4oQy3yCZSL8SF0g9PMGN47kqN0rYRkH70jC
VDqsAxh4hYfuK57qOlaMHrXQjGAJzXBf9n7XO5p6FCwxwIHT3u36nzUCTAcudQT6FkgMQlBCNfg7
JClV0FlSeW4m16wRsatJgdjXQZWi2eiJpQqQTPO8xtqlR6mN4hLC+8j2H3Q5nG+qlTifyvlVMoQu
bQqCucriwtezr1XlXNQUemWZ/jFoeZhG4ktBiTIHJYBd/g1w9L6y3XVmKrBw1a6GwBXstc8ZSC/A
gno5U5cqyLePpHjEU1+75yihQwbWQ2aCOq1Oyjxju7FFoeAwuQb0LgjwMxEYHJE7vfEztFgL3crY
zFBCx3SLSULmCYrvGgvSH5ZFD8YfDzMctlp0G3TaCTYFNrB0Pg67lfczPkiQnaMGdCtdK1gYQwQe
gvCv0DMssOn55Cx1mfkKT8to8bcBAJGmy+6ZJ1OBemKZdx083UVsfc0x4hSGieNsdQRvmhy+BNI7
9Z7ENisRCLclsyQI8RLLVDO97QL8kfJ41LIuhrY/mGegRBGVluL4iPHa+cok5rWHUmFFw3AQobh6
QkbV6bMlLHKJiFGr2+joFMm5+SFhWacDTwvCkRA5O33ef0W6uNSWRlK3RTMC4EUBGbMyRT6QqzUm
/ILhUHCNB0ZjxBiCHhPq/MzW6cmbq1ylvp6fCbTL1Lc2eFBPB+4xu8BKwsDYmkdghZRHJ17q1tQH
Qjz8EpdESTg6noiAy8TRumNj8np6BhDTkSLrG3eWO+0b1m42s0GR6dpfEp5c5OtC89QEYnGBzJj2
Ix+LPVgS1pN8USe3N54H772iCjOqYI2hiomP4wO6NxHHc2c2w31yJuvnJAkCqHGj5VTlFcuwMuH7
yvNDOhbQ5nTeNmAB//55D+KShkk99ePhKllMOPW25B49nIoKmQj2m0MzCkHCpd8NO7+MjTlkX+Zt
AOaC5xWJXs0qsf2aHrT1THzs1OVz03hytj8/B/p5fYFuyiliXDLdbi7oic9jylWQiII+kh1BOcQH
dA6KC/V5BzSkATqD6cFGj0BbV9qyDbNNnN0cQuzf2KxGy4aQ74oAv/IJ7iJU9YUjlXrOukx/1ZYG
zP16kKWrXk2nE/RRl9d8q9IzH2d1vNPiIxQXcdC0Re4KTzinmGf+Z8ObT3UUZfT/Ac1FnN+aKAAF
lsmFqFblHm2Rx5uMBNMs1q8I+nj0jaCH4JSwBGZ+Y7jvAq5zxzXG09Ea77KhiUvfhl/5ns5doj0/
tTMm4isqt+0y9W63J0IEpZqvEOsUhQruUi1TB4hc+NiHs0rkztnyB6jWgj/reJHfXtelLXrqrYh1
rJpmNK7TkGeEks7msQDsuCshJVlZMsfNU3RlU4aOsHDePQZqbTOhZnBEUO6D3NtzmtSiwyU3ylbE
JOhso6OyGeXe+8+YIiasbJadihZvUt29mcx0XDcyCU2K3JO0bMDdIiI4vxkUTPRHMTpQJgD7Qv0k
pv5vdVYLBivLzgI3NEnMkvo60jzDiOjLuP79NAg8j1lP2otqJCBOQlg91Ax0t4djXlqgHbhNOM7Q
cPpeFIS31a/dknT7lSl8adRQ9YTx+PkXETY1dS7eyngOhlXGyxQ0KM6ebsjN/C10/+7LVGnuPS4b
j7qK2RIhV3hAaU3t+Fdku/x5glciPiAXEUvygqLU7FrU1y+TfjvKaQ7lkWQG33qa24fMTELPFG5k
3TYPY7yE6YDgcRblG7fOdB0ral/09ICx/KBZCz/8AzA5sb2pAY7Cjj5VtGh8E0eaaDnJfXUHKPro
PgORkb2QHFUUIHDc5chxebIKfVcM7NDZVMSY9J7XnrSgBZSooTmFbGmF9r2MFMncccDT+kqtWEwN
5ENWTwwFfeEe0bkGWKsLKPNiUYEdwVWl/sUsGYKUNoTTBDvkAT1zPqrJvuihMfq8da/cOSHuwXad
ev9Lw8DQLewJ2mm/+aGOXkQDFkfdr1V3sDItT6FgPbQjILd/gCAIX1+84huNwKqrJQPi2bKMQI0P
0dJ4xFNn/ZrZgD0toVB9Dball3XNq64hpHtVNtAvd7gv7ZdXKACA/LvC9oqZ4SZ9xYZGojnlRClN
HrxbdUwgwwjrRmKoNUOvQdQHx8V4YWyTJuWO+jvsvqN1wUEPnHfgHuqcaQOvg5xvur66O+Z6MJxo
WIbmsuPuG7l2z4eVJSG++HVd+U/CtLuMYMhgguVA/ZrVk3GGS97UU6jROWaVAxDmwpwgHStdLGX9
XFOS6kmZCUc8KrjKcKtptzdfxhbp5HSsa0D6xfbvlnz238k8PaO640wwvsdTazz1moMJKgLqWJjD
uV/hRI2bhQi7EAaA/U5lkt5YnkkW6mV/EZQzAWU2/AqA+lhyZL1YAcM3DCZn1rh5pCMt1VQiEkDc
mSi86c0n8MjtsdKH3M9RKyTBXL/vjvLexlyndCUr65k73UUBzeHPpIJdgrkT88ucNr5fqoxh7364
vcxXbKbOT90objthBJ+oyeRQwi3OHSZknmrO8ZaC+qBwEF7v/ocGcmEAOEHyNDSXG4lkRlHxpNOo
XnvQGYjx6UqHZUZ4FE2Wu+GEOeVICZkEW7POxrdQJf4tiRSg1FUb9wAESUH4xaQuCzo78IissvwE
BaYXjDf4Mxuu3pfB05weuwJi73Em1wEaM5k73/M5EnPIF7vgRLoua0YodFuvH3Thw8u/NFbTFKw5
o8XiLPLJ4D1fFa4OKmbPpFZrhxYG/1WthXbCreXwTQ7BCHSu+XDvAW/2YU0dUpUy79HEQ5h7dlCY
L+ARFTEiYp7L1vY0MTJT9c57nRxgU7NncHWteZIvC1itlbuTUOhChxTO/OYcAwNbYvCDURWPttUk
PtB45e3hCriLrSge4O8b09WbXtYjJSCjvqft9Ddj5+5jV7FD28OiTvsGyZfSMUwyIZGkgaGhnq9m
NyPhIKSvykw/+ZoPUdv7w5QlJps950CHzTzaV6rUVQukeISvxMNv8ZjHVTQpbzerrZCbaHeni1lu
SMEVTzy2wNFXLvAF89qy7H5wV/mWZ8vfJsAlqYYh1itLZRvj/epxBt2Ypq/R+XOZwFENppNA4AKG
mcuYUmvoVu8wPzbJHKwdofadvotT8zZttYT72e07xGdN2NFh2myMm9CKRvp58DjBKpFRQiykvPlf
kZJ+Q9sZ6zxHZU57YPehTRsJP9pKtpIPqT7tdSD9+2e1M8ebnQ3oZQSv8ee6mCCNeBnH0htT2UCP
t8sn7CLv2lphE/i7j4C5QzBnRa8SVcmhjUxZSO7U6umikoYO83MUNQG1pIMTFMoBMAV5JWUb8kEy
q+z2leQFF2I5CnSlex1k1EufXzhfCkr8a02shW0whZtXcMnRDvrKohQ7JsVFn69GlTC1i7cMnzQt
TguO9lCIJFSF6HgkqYoaMa1zwgBpnJdHdFvdC6RmXUcl51bfVU0UrM2Lf2NRTcYNGEZEY7wbztvj
hYZ2IJSJmeMa2Rq3JNP7pqYtB8eYRZ8pmOUNFCfGVbxJ/G5h8hlRUWDMSqI5NZbznBiaER0I6QRf
f91rBMuZlNRStpMa0Wt61mk3T9yoltq/1jp/IZ+MkwqEskxamhbUYgPB5ixhqqRiIaGCSbf7XYdx
mBaZ221hoVmEnbHUzaskF/ssrbV3kFWIpB8FklBieYadZMhJJc9tYEM0wrFyIG7fu6fz+6oBXrUG
od889Pr8Np09Odqp8hT2NOrWbrTomTzN0hDmvlXYjLidnmGU2HXwZ48N3NGD2TLioASv7l8bNjA8
VWmYjT9gP2ErzBsdMdhVaAJfQRgnlSy2eovATv/3qg93L65epKV5cxTG8f1ZSVo2KvD4G3sycpSs
G/XrUlOqJhwwpu2G4ABF/ygyzHm2XurjCejfZSFDQm2X810KLissG2RIw3r/ZJLDgM5P15iIdba3
Y/CoHi/2D1HceYfpdI3inX6m5bAd8p2Vo1NiaeHa6g5cnAzoMJlUIV4soeDptN++HA+b8vVU2Qv2
yTCDSciPnxCifl6HFZ72PWzk8nENnMYGqjzoqQ+p9AuD8TZ6k4CH4TPdSLQYq838wYCFFyRQ5Q1g
AkwvZ8lvy3Y5/lZfR3dYbodd9dKNjqD4rGB/nByriGfMb/q27EWybFjLJ8VbmouNGoLyaEzle5sj
xYsfUnIZuCNRST+vegpPHp/fdg8E9UFJ5qI8QVmuuFZVN0yftmVei3s8qfscK13E5cWzycWrLjWQ
Zd/Fzys2Gri4WHh78H8oeXBKFe3c36/75sXuRVoSCuYjYYCnVNW9A8Hwn0HSb1Qc927mB2O0uzX5
aymgVtpYhxGZXh/8qdA0VLrr7j978mokdpA5Skjv8rYPru4ovCK7XZ/g28hLlVO5xY9pwMuXOvmE
eTfBKIYIhBVi7+SQxLdC5yOUpo84SGN8pTPc6pQf3pADoFb9Nyr29DQ00mL/BO6k3ywMOXosc3Yt
xgJnvolPNZLfwthsMjjkWKe60RRyHVbeFMX3qjSj7I/h+EdMchbYbC8NGVbNWe2Z3LcXA9AuR2O1
nAMxFDLtEF8tojBTb+24qXd+1h1smqz/82KASgjvd8zRFVsxB+CU/t5lhxEo1UOIhJXnTxuoEgnK
6I+l0hMzbB4VOMTLJ4BB7LeLhtbRR2+9Hf/nmhKXhNpIajP0s8ctJVJb8nO+P7o/NCDnMzu9P1BV
2HkS6jBWFQvbAQEOOe5hy+jH4J22iNZneqbRc0rZMOpLxpMeaJ1bojWvKSB30PM2Yu5H8aFSaGHR
rZfYHfNUZmT+X/0KqhawbFj6xH0wmX8F5yvGgKdjxuGVV3p+GvgmR1Ity0H/a30ycBMcOLsICep0
WjLmxC5Xczk1a8vT8BdUwP1tuvlcrOck/66mP1MJ88bWtAy2BwrWNoDZNRDPEXVICRtNIqWHxvO0
x8yfUagMeXR1cQ4Td3Ae52uSaKoDkvVDoFTa0THw9oEIXzenK7wdG7Nc6dzNAx6Y9GxhEZq0scGG
+L3c5V0hBwAMeOPcFq5biWuxKKyGVlGG7vbKnqGqyIVm2dGC2w4Vuc3kQu+uEHnhKQMFHyuyxCFe
SrKpk32C5PXpmwDsWPVkTWAlk0P5lgdRm1V4C3DEA59L/BYy07N+xYZq6B7nzQZO1vkLw68wmplo
qNfF/H+xYeEZsbe+gapTbBM7tQYx+fsryssQ0cbYYERIvUaIbQTZli8KzNQkC04bJZslqp9Km4FP
Vx5sU2Grg5nWYnMrg2wGOwkqJAuz9pqYobdQAiyMNE/98ecBz+6zeBK+6yQOejY9jwtPFF3KaU9C
p/ZMqMjbh4VGfOaZHCJrefYJj+Esj9vmEYfnCHEPLIwf35+CjwUtnmrldTt/yWsn4wWCAdOL2lam
TCTzAhzFfwcO21TH/48vLpuPJEZqYsR5XPGnkQAJDdigDVI5uWuKCUp/IXWd87cdRBWD04DRODD3
eiHw6YmDT10MvBjQY9q7apCA8qBcG+uzVSHMSyRoH9gmK9C62ZSx8DXy4SI9Il/N42LFYAJa/X8a
wTTvs7/4T+8R+3iU73JOXtbqVjH2Z1Zvom/xJcIseESUusZU/9VhI3dA4x36szcydFy3LNakokX3
/qdr/Ej94Puyd8Mb2XTr44IsfdCLhKLd3Q8UZ/FNyCpOGTFEkFGLUmZiIBtv43jE5itoeegIe7GI
opyTORqMrsdCwwMfYoFv0+xoxd9y2UlgSsBEEiW61VIE5uIEZzJXie+Trk330Ka6tGKOY8BiaoKt
MH5Yur8N8W7aaGkxkrjsl3FHIqvOzh3ns15f23N2puIz/M4kIiCDpNka2wdx85pRICUTPalFblBd
vlv/0yKvezdOzVnxyILHskV1v8fRxBzvM4319ZhmQoJ22W6wFCmpBr7bAIDVv2hljfiTQBQxANj0
unVaomNrvPrGVRjBUaxS02zBDIHejZUG617+rS9JUIZSNQN8/+75K4p2kY47n8B9NdT/ujuOVzAu
0NUkp2SwYkZ6brvJF8RPLdHYmIDoMdPzbxZXVabvJSpxRRCSH9qtnJq5Lk6JXf9DImoN0nBfCzIY
hFcrkn3xuIxabMb1KIwPaPZCeSrNZILGYmGyDTIPZGo75SAsUgX/lTCvltDhXbolp77a3dh2QRZr
W8OyRK2j40amqXSuUGZtC4vc9KBn229leZsiZLoojhLJgExJH4xkAwHHt4T/1B3VJaQITk2cBimE
F8lrkq1GQf5qrUP5tNSk23/zvBYZehXZqqSfJSxfC1hChxPZS7nh3li23BJ0b5OuEatEiZqYWxTz
X/QGFu64rVOqf9iVG8UCInG/d5BLZVgdNr0jzqObUop+hQ83paMstXFqfjvylTLnUqULJPWT7PS+
tAE+P1+B56kGesvbCBaZl1AzP5hgSgwtffYOEMIk3JYTzXsC1n7Z9HOVnCl2tGBhmmMapeuytGA1
5MA9Iwxdn2EJd3NorMoHl7OeYdBTpQZFzBamKvbKKQbvzvO6oAzuLMJ1A4jIgmiWBvQmSmtSM7tW
Cl++jPj4+DkumnFdGQbcX58j5HFngsJl0FfctkhheaviU2tvHXpfcfTjHjMF0OwBakpZC10vtu3B
Os4qSs3qHh9v2W0iaJepBr7YnwppS+5WJcGwEgMnqCtdoJnRvRlVmoyHWhrgX1aR+y/XIWwCAq9H
OIRhN9DhVurq9F6JWMtoqckGJku9bYSGpXxko+t7blEgy3Y3Kr21Jk5nXqqQSKNHQ/w2RCYnc80+
pqVKRRAkeOLuPvODeEwk8dPAP84rhmsmKB4YL43dzxL+gYmg2KI0764+nXHRlaM2xI6qOmJ+fPM4
YFWuMehKreQMHoTFA17XNZuHrInB2wHoQC0Mb/YnOJMCStdEaNNqpjH98HLxIhCSacJBtpgdpfUg
PDQ4aJc7ee3OCwfY36do3368siFiwUCf1Uw8E9OQr4shcfuV2hjP8D0bddjvPZ86EwxcoxeYyeJf
c492a2pwmRoUCr/EAATiKm7vQW3u6RZlXw+mNwthifPupXiOkmGu5coQheBi+41mDAeqr4GlGkSk
JBVIJcX/Gup8E3ao2m35QGuxvDXEW1rFAWya77gsER+G5PR54ljdnsMyCwB8nqDm6+5cphwW8xr0
0JvIbsacBLYLjzXPJeUhAc3FVThrfpA8tpiljLu1KQPTmS9VHeLNd8WRRAJDZcyWkeBe5tEQSkKL
1cZj+QJYlT/n9PVZvqInu0FwBRGpuHAmNDSRYhmnZTCsOzVQZiZoxrvXwC5RqvidndXQEM0GfpcE
GJpz3nGsxr0cq8bQ2mA+ENuG3pmS+vYQl1uVCv5uviaOzO6XxikFIc5rKzi4h+ZV6dTJTzYFE5sQ
8yafMSPiF8VqP9rvV3P3S3+IWVL1VInh14cHB4FSBQvuP6AQ/SyEuhDWker2QQhNQKkxKbaQQ9nS
EML69899Kx5YCbPYVmY6DOizqf5xLPAgmdOshBUmCSYJywEyXM+ySj+u1gJAkL6jxK6mXbwbcJpR
RD4BGuMNaFJDWww4UiD/0iiQ1hJVb7/MwguRL0rRVZTRsi12Z5VVT2dHMUARclYxJ3AJPinhWAqt
LUxksSuwWisqQ72ezs0mSP5FiqOC+iv4BVpgkj0D3t3JEEgWcqf9CMj+UTgfCSjess+oj6L1jk2/
o/gn9BL9cikmE9RaFVvP9VtK2cGOm9E8N7j9avYxDv4paw2aYSZOfOU+34mUPFLwfqsk0FBptTNG
6S4h1Ft6K3dgjhK1E2enimFhd1ZpNOnPGqbNn90ZC8Z8iCgWv0gcbOB+65DAf27C8HKJZH3jhrC3
fvUCFx5UReNZqXZnOfDEugpi1S0gLXRh1CpVghDq4nPtfB1aV5+yHXv7itKTS1mbAfAsmFC6dZRr
QcbHslZaVr9sNmpEZnUgim8I1GUIlkPhpwRveuqRy74y9fQtC34g23ozlJxRKUvml/foG7KV4aFL
UzVzxdzjwzsLLoHnai09Ofswf2pSuPBc+cUUEZaDnywMkjD6Lszo4bSK8TTb9/J5NKUla4gpXjPF
OPRyuXrJSGkXVXJxpfGDmuUt0nfPCXrythGCZmNGwIooinynv7DolgFk4INDdg8eP7+ZGS0JJTGE
Nl6UwuH86gV2jfoeSPr0uW8wcPsx8ZPuE0fZMMaDjDz9PGH05Cki0sx1v7N2iGRXQUdQSRFBzPKX
qL7xuaU/TZMUpp4neavuMI/6gE6WyC7svLXl/N7wm81dDGIpMR4DYFw9JL3UIXSG/FYispmcTLbe
953zXybx8VdsbInjMirUteaQ8j3j1qhTyRefzyoS3Jeaw5mznbXq2wSPgMRt0UJHKVBAM0QNABD4
s7xy5BKdnN7VgM6Qb+i2wRtHV4589wu6370SGTmvLjZiXTpti8BcMGvRvgPCdRAbozrnRcadVmzz
AKCQLBv2evxcpXP5/0bgJ1oQospZih6D29fPrk2luu0u+Pv2A8m7+u8jnuwlf/Bkmq8mA4c1Jds/
c8UtCBU9FRmavs0SkpBA96ybxaOit0e/Fu3UnzW0MpmmfppJ1DEmvZR61oIAmw8CcJ9jLmGrOizo
G9XUyjlyHqvvgD5h30eGFbiC8k5Z3S0GP5K+gltJzS5YjGp+nJo5Oo/nu4GAmYs0bNatMbadl4is
xuCKi9J2eMiPs99Zoz9hNF1nvfLnqXr6UQBhisJOp2dSzx1IuBn36v0mLpKahitswImA8X9FJSlY
8fosDoFyLIipOPESN2TXI4op5M7TQ+Cvjzug51Xk5CXsUadDRo9FZ/JsQ4pMlqi1CFoIoZzanxFL
6iJEA9Dh+rQcEN8+JDbwPfIzSQjwDWzQUdcRlqpzZ+7RR8qaOUX9o4jGN0ugTc1XLpeAJL3irDDs
E1MDBEfGW2Hw9dsIaJxwqapeBb7BOd3xsHAZKPLgle8tGS+pD/ZpfQi9yQBerGILN7I1p24LXIKu
WdeVL7eAdMobgA8zU6U27TC+4w+GWxBhPEdUv//pJLln2sw6Pm2ufFysMZVm6r2AlVTLoG/+96cG
66F9MpUBZTSybJkuj9T2ciZCiJRYw9wTBquC9/0S+1jkZgjriAspKSrVvXXECPYd5Q9gKuvd/wTA
oFb3hgXiHnLVNtzQhv0w8VJ1qTixrtYbpuqCQsLUEgsZQbQWHTA7qFOjvLvCwAx8vwim2Qo2Mvn1
8fXdjlQzicBt95kyUKoscVM7fc0X8DqgiedrPnnCUVnJXmaRu96BumdvDxi+BhKPFonr8/z3rguX
kL0geNL5gTmeCMfg9i5Vzhvg3Do/w6Lu3QRRdjtZynCpcwG58lxYRbw0CY1qa01PnV58Ej58m5nO
kuOgflSfj5Okgndv+0qledq11Tqxl30vKvvkc+WUikLeJgt9PhATyKJodudnn8t0sFwGjxttJt5/
fW89qmO3os58nehIh8ZgObpBP0rXyJIM9mfBIpG0PiEC9zPY0k8AsgEaN6gdTKbSC2FQJagjC/nu
qraSBRP2YoD+QN/qWTjfaEUCjLGm/SJa0BfUq301+zhHagNspbIWvUjsj8KfHxQ42jAu/0zNeXfn
WaYfArSesqxeL6wz6nuzRE60Ohm2tHbYybQVjNc2nB0pfT1gtWyAR/CII3QliYLXQykmUn88GeMz
9hcmdv+cVL3XN7LNT/ga34QZWPvMeLNOlofDo1Z3eDpvjTpuljhL4nNribS//wEt5vDofx4wzhb9
mRMziBIFpGYaAdK2CNjrzbyQ9/H12lquhgD8sOYGJRtSRDuaa4OhGlIOYkXHw28Z5eCstVNT4fbU
QzSqoBHgkVISz3OdpIaqcrNlPr9UKVcdrCwPLDjnRdlm0NT6CeZhUWfvMXm3RMISLuFW4r1tnYif
4TNLPARBNag9L5aLFKi5ogKdxfSVFX2jw8bQoY0XDCTtSQsI2CVAnL7BhzHnN9OEgGBnFhwf0UMP
s3erkw93y+8LUyFmz5CKTiVEwueblEIAE3dvmEXUDY9nSrOIm2wX+cnd2FqTfFTMjVZsGQJ49/Ic
D5uhtWdgMXC12cys0V53ybSs7RVrBPJHX65qqabmkkEN54Yd/8MOTQm8jiaZyLPB0YeVW3red+T5
pmWhs/4Ba8lOiBrZn6foFH1oPcQio9MWa5u+RPfZkb1XZGNTKu5COcHvKLthkcbcFSeL0GLV7tty
y0JjT7M/XHm4GGfe1rmRbJIkpGU44dkDS/rcsaByRHmENkvcGZCvIm7YZqsAskPkUgyZc+DBgjkN
QLYsxond249Z6N0+QZCfCruwZy1ZQp7kT4yacGKISCBXCmMXPCqucKykZwDzzhAALS/1XOSjO/5n
neGy5vPf5w7qxmcFKlODJcEnFiPMaG7Aovt5e8KVQqGaqhXfoz9ZH+nOUTCv3C1FwxtqtRzoZ8+Q
sw8ytineJIyaMvrxx0ZgpEVxO96PfRYawC4F0YlJ/oD7kT6QMOTUQv9erCP4DbI93o3Mr6AcPb38
62ruOdU43jJdS/37ocr9sCsvfd7eGWGQg0+IDxI5FKc4YHqsZnVLwHy22ce5n3bCO93/Ppcnta7S
lXcAY7ob73XUnD+h5hFPhYuQiO6OUeGLvl7QfPQ8Q/53TtJWzhzxb58fE8evm264T25QZN525zIS
QvDOyYyTH6zjmnIOwHlYJE35Y2wcFZP2zCkWuEzFRpcaayMp2udAtnUZ84VU/hk1/FjB2mlfTaTL
nyYhRLWUT9Ed+JfQKrNRgNYLfLNXxPQ4wffx838xFbgqZ6v7Q18w3UJnZDDFRDIusdoTI/lYARxu
x58fWHPm/diVaSs4BqiP2IDPV1Mg7l4Z/GPxnR+nwRVIEgx2jW+EL1lgVHxmtUVnxzVVnJR+hD3S
7c6VqWi7qD9HjKmjx1RquoFR/p5o7x4seJRNvv6d3ms91GGhs4X3jdzeKEEfHa2FkByxpPrx90/f
BoZS8NFUz5itNBqQSTR4ktY6IaWXobRgw9z7Rv04JzqmsXzTrB9dsaGVGk2pvUZcliRj7oBdrL1R
+JUBMl6eKbUL7onynv1N4EtUU6SK3g47xjNFhKXx3iiJXKtPfr1A420+eZtD1VWHocwjAFojx0Gj
d0BYB/A5itI+VYFiJnVno/B6Wt3xeLz9jr9GCac6Y/Wju3gebCX9SBjnd+r8ez/eRXtKk4VF1PQq
1AWu1ohqYWgNgXY+KZpTP28psW/VUDKpIIsvrECILZzr5ZEGfX3t8QL8pqy20GUTTjwbWYoKSi1n
YKs53WY6eKxWA2WvJsLArtmCOxz3HXjtEtMmuC5ovIQF1jtuoKO82GJw11+gkNAxqPSRc4aqmX18
umoivBp2QEunXSpThFmI/88kmEYIZoeK0hVRQUzLu+wez6OGb0Nps6Sc1bNdeaWvxxLdBR2UUeHK
iV1Ieo41FDvYOdbSg1uruf2TyIW93gaUnoVThloRAI6TBx3u6t2euTDnMFAafFiW5Ek7gJrKIS36
ZOO4x4O8gZUCGUVLrVAsDa5G8+pWsoEfsCM+pIpLxKbotcXQurTy1vYiJOHudg9KVd7P7oj9g7+k
EcrKAgHRZaKnxKPvbF/FVaLuEWqBzvImi9hjQMRbNW5OA6esT+Tyz9Qa8DoMzZgp0XbtB72LGgaP
jJnldJkL3+1u5EY8hMqRcd3YYNWoOZ+aPzqZCipPqz90x8jtPDgC1bB/raGwGJvfIHDwymTiMEOk
xKFolNYOztGh2RJs75s2eaH5lepm5L4sQIwBX86JaUcUhoMrNQDgX5uO7TNdyxXx1gBi0J9TAD01
E/Aa5E+JKDDfPU3vhOfJu70o2Z/YbVobfXzxDwqS+ngXsQRikmdsmrtpNg4EQ+kUg8zUGwCeJGe5
9MPQEne+UGzWq69Q+GhILinOQzxU1G/idnAPhrmFUOAtT3oQ07utrORq6rolcxdjY33PsZwMdjy/
ymwqEy3/nLzUMWLMjlxNtN0EqIeCBH0buqhdp3kJXJgEh57zMoi8p/vnRLS0PZIxyxiVxFtkHZ8R
OgWFU+2eBMtpwT8u+wzLRoA7xp+cXJpa4x3qHdfBYcBUj8DBVEsTBSz7ASGgoOeLdJfmBQBeVpXD
0XlsOOl3pgBVuLAgJMWRN4zIiJfHT0IhX9x/TX47GWpIosT2Q7C/oNHCZmoP3znwB2lYt4zpfo2r
mlpfDI7uiHejQix6b4+dDIslUs9zyC1nQzPQUuQmsgc+0ruSa2Cob5ekCE0fHzXGW/1GxK6MsiXf
7HF6e5grZxU8H6gi7bXqnq2iNpBJdgXrkn4cxW2bT+uSdZ9dUoEgT8nf5t/vbvKEXGGJE2TGU0hi
yFF15Tl0beBf2VvIc6mYb/Qkc4R3XBV4Cg+ECRtyYXEieZo1+ChCZTwExMWJpEtZn7lnbHO/X63o
eKcyLugy6PgC/bweVLDh6+aXY/DjiWKEDmiSbrxY2nmduJEUPScX1U7VDvJcDvgGadEG6ywq0jgi
UKQXidjCmCN9AW8cF5y8Zk+snxIyTj68W/5tRvlvL+izr14bIMwXpDYtXjGekIVmFEKh6PjllvsT
B8A7td+QKz4zq27QfPpGqJKiAdnKrB2e2uVsuH5miIo1kx1x4L3AIBVq9CR9bT7PHM4dxVa4zCVt
cy3ZUD7+/uKTFDq1LYkLoRWOTVOqnY0+ov11aD21JcWTKtHKNLjLyv6keZf1xiROmwix96FAC27+
TSScRtREw7DbhLuLrDIgITh+exgj1RztUdnXpePRb0P5KmgoxfeLaUf6fe5ETASe/+ar065AXeku
WevjO01NSlnjhgOKMeBiBSGg3hhV3ntVAB4iH+bD0dx3FJQGKN/b6CUToaLTdFag8SN1fvOHw4Dj
YMrPoL6R5GRUsHAsZsCksJ8WfaEc/D6XPNUU8cCsHxTGcCTYyBqADYgLrQgH737BNzuC1EAOepGp
77KqXvb4SipEgUMCVyImGmTuApEQIMueesLUKWO7ZyrmQpfoLFbCckMpTEQ9IYQlwCm7yVYY1vIB
nGjfT1LcfT/zR4YDxeI4V7uV46CWsJ4GMZNttwj7+zXL1htZrcTpo2I8HyIIAbOJpdY/o2y1+QuV
gB1Fen3F9hxbcGW8ohA/wOIJJ08OzT7S16ERPiOWXLRzp7mUQUFjJfAWGeXccv+0qQFsR0xg5WBp
CIqqAZJaW7kal1g7jxFXUR9j2eNmzTaQmXamGbjUCmKhyRWN7IzcvL0/USjUssJNOD6fGO+Q3jdu
HJ3pd8HaCIhuNsGEgeXmjSpDMV6Trn4hMzAOgaqUFHtp3g+Nx8OpODYublh8mGNBI4AGo8FRG40j
XgD7uNnzxQotkiXB3sy9jKZ3fQHSVOSZUOPaR5Qbmvw9ZqgYtywr/DBXKgWEXTLdDnIZpltzaQN9
g6Ynqwla8sAbLTeEVMt0IBWjeA6AFRcBmNRFQlkpnWJtIEn3CkvBzd6AGkOjZpYWcNYbVZvIoJDO
i9ggBOH0N5eMDYbO3GPFdXyhekLYZpUbm8u+yyGx4PPOWJqzQC6KdYpPdfeIZLfE29ssuo4zKgA9
QFiBVo68LEggcBRmh7xjeR7bYuDeygPrrwW8eGw4Ou7LmK43RB+JUCujJeqXlcV1ISfe+wQcqQEx
cWxA4biTv1BWCT7v3dupx37d2GNeKQIMEpXMT4OeK9rmyprjYQkUdvdPSsyy2GfWZ0ZUaiGTjpQX
fbyDm4ImRTxV/3+zQO5AKyUXGV5IL2hl/473XCVeorLlA1igB1zZYiSqoNpCo8ik8Rmn+149WcFE
ADe92z6soQI6qdHRtFBQwEeorVGeP5vzRUdoszDfG0bemXA8FBeV1KrflUpCR6dNR/jl3bWBkP2u
rdbuB24ezysUzrtf5rthWyqUHr0OCYXsThfBbDJVc++YRIxo6MrCyGDZSnV12B38zcL0MZN4Dr7X
nGPjatp8DO9Uh7KftrDIf9L81m0XBgPdKd7nCSxEWrcMpczGCXRHffe6fAqRMe6CynnPmsIiif5/
12t9HsZt/5zxlTnIu9OMU2yypt10I++ObmvUf0KQKE398FomLJMxMk26d0njfyGVtWGxnXU5P0sa
LPnUFHW9kQoYcdA1rDB368k7UE4xsCpMNxmLjbarBHV5Tc51QSpV4g+VPCF4n8xrrVtcuYV+hYcE
UMfv/vKgMRD4fIbIuKY0lv39gm7AwZ3U3gMxqulEBjyPFwQQ8y8Fy4Z4tcOiBccM18JGidQ5yCkf
cPzzxgzZJkftJHTGQ3e6Wp96Tt/aThFKx101DDQXPnC1MBOoVpsMzoBvaNsISaVXiDf4CyCYsOLw
ygiOGX9IpRro3B0ycBvPBgjF8RaPkj4dUR7fJQkhBWkSYSqSOpRenKyo2F8sxtQ8YHzagM93/1Yf
XVEQfK1pfC+DEmrhmoJC7oQ6ZAoCzvDtRt7IwHQlFWpu1gRgYcKPDguTNDgd0b13wXFR1LFaSCPl
UlhiRUDMmaXqJqiRY5DJoxOnDpVB15aQFtHb+yZDdV+JXOF4WuFL9vUy79DjVFjzOdNtPsNQWg4O
HWv45ZDvqb3WkItr9epTfuYhhTgv20CAZEq+SqvfGWfaCrq3J6J8FRrDS7nL9ZLqAeWb34Iwy+w8
WKvFvvXd7J7lpimFY+jPIrIHLPB5M/gyxNckzahvvn/HXD2JKbalt/CNP+g2lsXvCvIhAJr7dcvj
RJpyk8yAr4WMd+OTq/ODGRbDcZorvGgWvOjdqfTTBRpwOBaAsUl7dfl5wiGaYiLFtCFH4RDp1gND
AjIBgJG0XcYnO32v0C0y/2pRO3wXUQaJVWkuLQqL0imzdbil3tBXMYbrIwoEqL9CzKC3bhhswdUR
l5D3IgZLEQTGdgDo3njdKGGDaUKkHzrAq8SD7reEjXA4ZqAooJeHDHo/wwFScaFJgWOHQ5ST4TNV
ftOScJxKHh0N1y4C6VTNyi0vWKsGwK1vFlwepX5cGkJHNi1thkTFG5PhNoBSoX5TKUjcWCbNFgb1
SdOF89e4LADUHxJZCWiVlKv3jypSC5WSKS2cFSSFW3BZbDH3DclpCzkYeOuEKkW6t06tylisjH0c
w0RoouWNHKWsipyHYLuDPCubUgEtJk8TkfPcc7V9UALJs4l41mz5vac6lP05rMKYWNmdWd0quEMC
yEmJQ57+yKneVWCSd+7mGG2dVVGXTIyJ0N2S8TSfrGZcL1XGc35ZpAz9Jx/3Hr7HkwQ4NAUVwrW9
W8bR3LaH9luXIRi4XIUXyjqxeLEEim/tEPHUYjbTkh+U22inZT9ihUqFJ+4DG70Cb1W05oY2FTTI
p9iogb+qkUT14rZ3bE8n2EEAPlIDiTNu66JZE1IPWdU0WNAPDkpOGk3Dm9RV5+hmAd8hMl1L/WSS
lrhMrzL+ANf1rygBUIp4Fq17bzmT3jmgI2jcPaLxVuKPCLPsMH/HOmU0mtHnxu2m39/XgDGhFV4m
pgtn1iFzwdJMVumTwimQawcG45kwoRmWrOypKk+hISQlcWqpzUY6Prw8eBjY1qKekv9gXAGCZD7y
m0bVM+JKrJ0g8uYE2jiYwSz9gsh0gmM4M+he/hX0zUJD/JR9Ob+dIrNiztU2x/WKbIHGNu6lBnKc
Au+FnMPIfmY7rpsGGwy2XfWa2kb2BPqNw+0AXHf9TqWgWsy72Psjs6WwqsXxr+lpXglEu6NGpSdn
8OFxPrxmf9lKn6DOhA0ue+WjhLewKF/oS7Fn0qXOecAM66p4FqFHWyG80y/XrJWT9Ko8PoY19VG/
Ng0qoFOfBcmgyKk/zdEPHIRw/BGhRnCRmU1C7oO0EB6Fp5uo80/TOhM3nMazfeSHfxqJwRD5YmAW
TiuEt9J34Jt/a+w1UtZDFwlSvRbKP2j9pAFHptsTW46HlE8KOwm07+hniY6eRbe0I2aHDafcJKEd
Rs9j++Txd863D2R5sqrsTSReOpbTmoXUrEfN6drlPraIlUu7ITwXxGoeTaaQUdPB4vhiHt/bD7E7
Lc6/hMlYZCeApmaE0LBDds8r4+BHeysivSBkkJ3DteX6F2DdWaUci2gJjcZy9Wlh715NXbdicWH3
oYBZX0R6P3ghRb0LGrmIMp9n2VKtZYCjRC7Rfg1iFgBUpi65R1wRfwKNmYWprxrI535XGRMnoVrx
OMGq/1fKfRLPLfMJcyqZwHJedfdU7uFZbnJIJUFl6rGbmcjTpxEDYTny1HsxL40XIG1eFUOGdPyx
HfbRQg9U16KYYu6qwGJX7PzSghvDYK995HborFU7skwHQDiC5TTya0LGiP1oXixBn2nU0ilCEqwu
6hFr+VzMif47ROpbS9X17tHk6IDrenJjhGLi2CXUQIxbXqBg9/vjSSttp/Hk0ieVgn5TnkkBDY+A
hsYj285bbU6SzqOZ59DezlCiFiIgHgwxcczgfjFsBg7BGdBliRP4nUCaUO/B9PeiJPHlGQc39C/y
vhvTivFKHIZuVTzZtnwoBde4V1pBgE6jqocA4SD0YPLgSPTfvczgzcauPsaInbER86IhTVagFvpz
IZnbSZXYDf9UDVf6/O5MNTMWtJ7uaXJSdjNYFk7HJ6Cp+HQuYnV9TU6bIoyqsv6eQjl3kWT98COF
80HC3eWwPXPpb4rt65a32mTiwsh3AfKubVWg6F3bLQQld+g/DoHQLn9iKJsk2ZL7R6KsUgtfoUoG
8vLD95c1AxX9W4PMldr6ene6P/HRUv4hdniL8ZeLET0JIRPbC3PaxO6YkuA+1RPdA9DSSyUMxbC2
uO7drhiUPRWF8nqv92mS/KQjVIG9RxqLJX168pFFGN26ffM1mxoXEpi0XF5TnJ6bxFZPBVbYWQGJ
B9UW1FsoCZjhTXCPlEaJOHAFzYjWs6UfA4s2pgkCzUfw7dfmq6URGCjtpBxn9mFaCA4x9bcjJip1
I2rIkOOtxQTmyhuQVdhozAQ1EUejOREl+dRTUPErDi5f9fpdgEebiUleOmkiv8hWq2TiM5/fzp9Z
3hqEQ5PHdCqWokry3XxibfOGbx2whFubNCbBmYpgG2H/2rfgnJqVjNora848608Pjf6EfRtCJ0IX
0ro1QgFPdT1LuCm39XGkX7KOrHstHPijBqDpX//hc6ONdTYCHaOOPMMNms96FDWbxCfT5SOdCVj8
vdOQZxnah9ZtjWP2QVUH/eph6Bqe+U7QLy4+6LFkztEhurZEOHwkSY5VOhsezHRGVe9zKu4TqVe2
j66Zj5+bbnETu5vxUghL3plZxdyCCrGly1r5yiS8PnqPoK2cnmqk0fNtBte3STEFjVCo9lrv7+ju
8bxWRk+GNPSD68AiHIRTeEnkCTRM1+92U1fPrlnWEmCgLewkgGzcew6M4Xp4Yq9zw6vjp1ijPOWQ
ceV1046sufIwH/A56NauYM1K0gPapBKY+7OxI59bpEqP04/miyg/IW0RnX/8zwj/VgZrpi1OAUKf
0aDpMj2n3hc1G6SR7lO+3pSXvjIkCysRFHRSLsJ7aoAIcM3pPhl78Lfl7I6a00emw2+zBigfHIqy
UmvbM0QOb5CB+LRqHiGNcR+9ZFgQljqVLAhFKuxgPja72hBzi5h6OrqxyuNFnSWH5sea6XLOWjpe
Q6t7zzAeri9W5bpm7LgblnVoI3e8uM8UBrZP2qKMt8+ekzEKwl8Hrx0xUETJrD1+ra6QDCfO7x2r
bQ1yRJ5pTTOKC+0h3nidTdXnuCrVXoIAl+m+4n4tZhCqax9zQTFvWLS+ei/wyjvd0dU520COtt+f
0NDN4PPfP9s77godEVkrq27sXM5Mr0hyqBDgVC8quh9SYKO/DivDXGposMILYyKs9HV1jbbjV3/Q
u71GxYeMHw6Z70j6t+CQRA2kfpSYhqFhE6OEZOPQfA+1aXA4g9eJ9Hxhf1QN6JKrhAGORJ8h05q6
DrXlFBpEGXjgaB0eHO7n7jro+R+htnSfguOO68fZjjz/JyvZFBj7Ic+duIVTbICrihAWoReT6p9j
wVu4LSyLtCCIMIKPQOpl03vsR0sLaLGnOPaLJzVxEUWqj1fkDgtl45kCuH9CnAPaDn2Ab324As8A
yg880P5NShJD+oYtTc05a63QULeecVtP3+SoXmOT6jqYJG9taZ4N09ZC0XXM5E/rQmjaVBXW+gAa
V/aWIaE9LiXFOF5EUt1NDn8bSShAerXvq/yCS0fcI1oi0GBGHUNQlIwHOt9FYK1BcfwUyWDe9Epz
3hGlxmfU1aKlbzx3Oljn+O6YCr7j8act+yF86GBJ78kbappIbtZgR3ZcW/+gvuOeZyrWtSm916L+
evLjoDeelpSzuAh9Lw8fd55VX9dd4h7nhUJQvdQ0OfUNGr/tSanIqO4CpAF1mM1poQEPU3dJcWWk
rwLNSgkeXfebJgNTwxjdt4lzykyM8t2oBjRln8C9QI4ArtZrEwoUoDPOx9Vt4rHtSMb8hGhTU2zH
TbQR1jAO+361Y5rJaTEn8gfpH5v95EWGuuk9vKn9nM8gaTPgIz6Vx01KiNMVaxVj0hQ+YxnApcsI
aOJjckNXsnIaCsR6eqWBXUyApNOJ8ycAPzbX5Dgt5pV7y3jQVFdCv/+wN5Y52YBy6ecO+OeFo64D
Ixj1nS6kVpGeDOMtPHH20M2i070YT428xI248s24cFwPnc0Wxr7oN4969S/Ki+ORVjKqpJaCN1AO
O1gF2IeT/LlHmqcMwVGyt1l3b140y2HMVmQIB1bh+1WgvfzpOdvmMeEkVQa/e6FNen5ygdzk8DbE
1VBDok58i4cpt8jUeDeEN81SzrqGdwsKAso8fOz9TQbGL6B1SCJOFQLSeEtT4KjvCxmwk5PWvmGk
EQqRfpFeniyrICMojNZjPIxS0J/CJ2SA9p16VPgPZtIGDyaDCk2uslGRHQmcEwyChlc78/e1xTrb
/Bfpq2GhRs7RLXxMKLrIYJbFaz5+W1V34gEghMBdXF5VEptb7BFiwa9lNkNRjYNGAfZ6J8k4yL7I
1dH9F+JNai3R1nhhAnklWgaGEokpGAQafbP6zcscsv9m574Ss1DF+DaruJGgPfCt7zIfa0H1oo07
WhTUrY9Xrp+ZtKuUiR2siXGucTDYSh1ye914mutYfY2AuxdZAljeCbew0bLK77PqREf0bjQ17KXB
APIuCFjNmv7Fd8xMiUMgXseBgQM9t9K4Zr66Gr6oG95BjY1vJDjQVD/49yHBpiVmGEV8mWW7s+Fc
qND+XI0YMAycK8HvhfcQB+McRA/1ZhO4PtDjjHPslFzSExoFqKo+E29/niHrudRtplyHOJ5qRk/W
PYkTI7RAuChVmSGLdn8YhRor62hYcz00pGKYHU1fHO6vVxPR64/CVNsywqj8WcXpHC1blxJdBuHW
oEDxAugShfOETCUcGMCQo2OU9d5CCbLcEX0/WnYIwrTOBuOIQbTDsVxev0er6TODVPL07r+PHTjs
b5Jqwl5nz2MEd8aGSLb38ehJOfidTVrZpCZqE67o8zE5lmxatTru09cpNtp22uaQSWAic8g6Llxs
zJHPKFGaD1lTRXhaGAVGGyzT5vR9T2AeJSOzlHQjmSbYI2Tcw1l/j+tw7AWnVoup/a22VueMzoqY
Y7m43+bSnEv6yKCP9ORrGl7UabSz3GJVR0Ru1G3hgKhGDRqbU4Le6MDroFFLPkcZOdChJPIIWXTh
eg4tHABst5KEAJTdmQhBmAUG8bTYBikBIhF5L4DkDxzUQJ8Y/8282Cbnrc7asKz9FfFgawo1yaHz
w7H27pz1d8wzKvhNwj7zhEyeLDvyJyUSMI34l/LbmaKpuKPvpS9fAIE6IbKOOKfji9mEHR50WEFg
YpzdR7A4/G3VnA2wQ6i3ivmYfU3Uss/rhtuf+/VLfH+NntVlNHDoWvJWXjLeY4vVY3Kv5EUkEkil
rJf7PU6ifRvf6Ju688k5FJCe11iPkCLdvlXuQxBCAZuzNrFII9i2rP3g/lU5rWgub5kB7DbL1GgR
2mcTtFXgA3AbuoffLfJelR2vb5cZmIdXSlkIoAKxoCyOvNxSnjW1IAYPVjgkDyswIKJs8uQbT4wy
hMfdy6ZFggzTxSZ8EmvoEEMDnFnM8SM9Y3rmqeP0HKCbLiH6lNt9pwcD5+puSENgUI81pKXukPOX
xZ3ufci875WP3FcWz3nMSWXmiucD4RTomRFZFggD11FpIAeLyusmxncWgd+f+VFc+l7z4BZrzBaK
kTHdzOakphgIBuwuXuJJA4HjbLRP0BUgfYdoIaxX8tsWp8VtCOrkNMRpg+Qo2tdJ+W/oSduCwYRe
QYBbF8GM2yU8Dh9kTuqpWYN3CEVyTO8i2lZmZp9AL0+aMnl2RUXQcl0TaaViMBI+AaJLwkEUY5eD
VuGkjSl8Q8AOhWCH8BtmgGPwHsBSqKnPqekC555TqFeyHorqDogEvVbHUdC6cwxqtFTgruBW5BeJ
OTHsod8fJ52N2JVM8MEX8JJhAq7hxRe6lz1WtbouUOIv4gNArvOD/dPmCjnFFhAk9rGxjRp3t06H
uPUln+hUPB+AR849w44Z1yQPJdJ9NrnkwUVOrqkdvAMyMfMXIRLF5bE15veyc3e9ltxi85/M2Z8V
fCqHbeSxbarm/KJYhdmx9eTYfM/3OUaF6lpnDVRiLqCR9QrcrP+K8lsys4C1wP6euk0gHNltaLfY
D7y8tDbEb9l+3ynkJ1G44fIaaMfbXXfUBbeAQd3UC8t898yqd7Wiaz3QwGan3wpP5mH3CzCzDYFe
sKuxtbVhlqj17lAnZ7vqtUOrX4ztwnBv/5Gz+sv+52ylqgwWjD4wxlcQaX2HAFXo9aCGOR+NBmz8
s+NcFZ68IoEQ39+fvae5cDFyVWROUbovgLWSU6t++1Lp3RJtFnrH/6QcKKR4bXdBuvNjpp9N0Ob1
SKTJZwywqAqlWDCv9UlfJw09wogYHBZXy04yKdimNsK8mXRNqHx7yN2uxA/YJJdwoqiIcrg+T177
vgIPz4G114b61IUJ8UNZ0bIJ7IC+lo96v9ZL9AQFgImgH5lYLPwy0yR3hxa67paClQlkT9+3CJNf
SOtYTG4kVEz9YkOS1o5EnrJesu/moL7OT9VpdchLiJhFrfGJxcb0XBoKm7hgoK9d/jNQcmnyj+Sm
8+LsxYqo+GlMIvaMNcu4IV/YgGzgVOhjd2lGmygTOvCzjSCpmeUjP3bmkTcxy31eOP0IaIj3LHQf
5J/hH4AvHFi2MV+pMUF4ooGsPU4N2+JzpjaAIfiwmD6X88zH+q9PUFaX7/8NKQdptBmYIIbM3jEl
vT4J1YNr+Fdzf7fMXbjfbQmjyiY35uUB+2nVu2v7zx6nHiMZLQLl52ssJOn4cCtHsbTHIDbp1qkZ
f70ruYMVblzT/FZbHaMFu3n+zSfB26TeVHmIAGANz8U48Xl3+u7Oh5rSENTaHYP7GmAY1WxFheuY
2K9R9/e+7i/EhmXnJqKhq5zNnT5ETCTzIMELzfV/IQDWLGRZ3kZcUBIJyw/gxYxqslV5yIom9xuH
cR+q8DkNZKHWwnlcpcBzqhVUJclshvFaudjeaS91P+Xd19Vw3UfpxI1ybKt3Z7gBl2fRFWtv9O/p
OgkxG008z3v2XCnThDn8xx/OjAGvEBb/WpM1wZWEPmB8DEIT5z92uEH8Wjsu3oXVcDl9ichbiPiy
JN3G4ziMHALy17Zp4SSHj6gOcGe9NAqueMW9UVMcdjBkC8Pf/aOMaeGSrDKzg4DKPWxVI4o/kURD
1niqKPmKXuviKsKNaviaXudCe2LtNqsmo3pt+H7HyOkEI3iakzRU732eWae9HgmTvECwvEE04vEs
LZzErFyRQvgnWOMO/2zCFksVjKQJv3M3a/y6xFYPUrLMi4sfFOtpnVF4tHT5stR6WE921LXQmaAI
/RSEmUvfrkT9C5wDJHZ17OBMAE9PJ0k3Z1UiV7YnJKPTI87EIb8v1wM92mkTBDMgnkhEXN7oj8eJ
F4Kk+ch74dIX2B6T63/nOcHd9XUz8gCYePgrQSFsEGSQQw2JqyyGyrgLhAD3yMT96Tt9F4Fh5HzP
M4k2Uvq6xkZk8hi8zovSMtuZHrKev3bRWfslIblVf5ywIS3uC68B9ejQ5sS1ObMwMUxu9B7SDgmV
Z6i/5cHXt1C/WXtNLXreGh6xQhMfk+4bFT7XmIuCr7m35gora/RJkvdPwoEMbqSgJq7OE8565+OE
jBB48+623q5nbLqCP5mXFEU+g+GivhdbMlIzvaPkomfJSCaeyhtryYQSs+v0XEytOHUBs+GCSd/e
fn/AXI+C97U5HNuNT7QFuf4IeYmrtAbrjEtKFNCRjsEQ5OpPMFt7rs4bCU4rv67b+IypgVlKhKPm
XMVZwYb6unLP/9XxPS3XEbmYruJclyD/cZ9ss+TYOITrTzTzowGplXJwjkJ9tSQbCA9oTWijBGjL
slJ7WW5/le+rILY+Wm+ntY+8Sb53rTVuxnTDFEDcV40UWro+gYi1MosuVwaEGGwpbygCVpU2OcPS
xAXHy+boOu9aRAv+aA31IZdP9lCjquepMypVs6jLNZdsG4Nf5SUU1g4FI72i3NWhMcB/nIYLyDAG
RSkPFdOGRjSU0YgY73kwXdMqFJ/Hg1BHAKkueDsl9Dt8bfa8b7NeMiGIDtxp3I6vF66ZfVp1c41G
+ZOW+wFiBLCeyV6349hcmbs8UTbeYCupA+MhzlVyKYA82cGwPNHmEAr4uOsiNGxn0EK23pF/Wl2q
lxRngcPREHcN62jsLEJq/KybWlEq6l9GZmdKKZ5lf/SqDpIg7HQGYVbCrfIxRX+5yqmcKpBQ2XiO
4EeOWyP5AbxRYgHgTjItUQzVtp6MkT4LBRO0CPN5LNvAMMDBvH+mwGj3oC3H4gPwke07qeW3azIr
Si5/hQIZaS7zx2I+pdBOQ433nrceT2zjjgo8Tcl82y1xAs+jk49f6rcQm3Rm6sJyoIs8AqaLTSJe
PekJwKq5l4LD+9VGqTKknZOxdPjR1z2Mej7QIebBgtz5ECHUzlUIWwZKWxE+hcZXOgLPtEMOM59m
GVM51I9oYzArgU/pk2fjRUHLQCXsAnm1RjbPJD5BmYgjgptYcrvBpxDJCcgYZxTSgYIhjfs9C3CY
CY/7y8sa7rPO1QSQwFQwImYMGvS8QNwQHi5Mk4chbwb7DLWjTQvRU12Mjr8B4qYiNfo+5Kzt55Ts
3nqFvK0dsuZv5GeokcSjFwzS0FswdP6+B5p5GXmkit1+YNaiEM9WDicnNbr3BE3R6kbQ28LsiD+f
1CZ7I6MilPeva1cxLlQwdSWIXZaWCyYKzWKS4cAYzFMvTMbtegVnRLTLfJjC7E2hPpoAYgDa14Zo
bNhqmCto1UwOtI+DEOlin2ulaBVJuFYmJHGWURGFFtV0I6dEyVl8LEeH1KB7zfK4YFGJpJNnznMX
lxjlt0MPiLpLjl6pihViRpCMGVQVU2Ygm2K+r2RtmBs5rkYmV/9NfDrX8LJppHKcOtsc+/QdHjIG
84Ijp2CAH7b7YG0eQE/LGV/pZSYzgkDAOwjMxVERAA01+Ct5ZY1VpEQVqV8CISwFNOXxFmkv9Rma
fZT4RrV/FvUAGmqOjgHItyld9S8SpkmZnnTXjR/8n/Z7VuAyHu6MtxHkozrrxIGRleAslPo/USLF
rCNXydYXJDRhXRJLy+GK4RvhYIHbUx4sm/JhVWThLhKG3gtX4yf4uQEW78+mLjV6ObXjyC6Hr80X
gwzCLzEx12RxGzayh/JhXOaxwI7UMwAoOL4+s2pCozlY1VdCc9urMzPabrFLq2yg1lX7AS09BtLf
hV7lCtisK+MIOPAtiwsPJK2IvhxOjOPGK72v3f/xX9jl2+OfeH/c5msVJn0w+a9FTYzk4+2p1oa5
SGcIwFToSwUvqMV6SSg4aljgsLyPcLhePmTcmn/2EL/JYNYcX6OpEl8GO2yRgbUKY9rD8k3Gp3Wt
fre+WGYacM/Bqlj3Yb7rGVk8Twh35TnjRtNAM2oVD9xSFU9jKZSKNCzo1JI3JKUoPtBiKXXFl9Pq
D43zrPqrkYEdQzwNchjgy+7Py6VslCyvY5kThs7b8OrhDHIP9IHOiCnztPMWHxPrMMb3QqSIoMu0
qoMft2CRWramCSbPtnLGkrF16xXprWPjVu9ebelB3Ce4ZGDxckAiGaHXV9vRR0wsksAEDVspiyGg
2GAMEPNSSlf66qymu/cNOVZm0E4t4IH3ci/JaRU5HmikNnNalj3BJS2NOC4KEBfFjaO9ve+unpJY
i6e5x5TU7jfrwg0jk5LOA6kNdHpeTGChWv4+8R/ZUnlUu27fJvY+bMxqs+YA+mpRDIGOf2DcviS4
L0OJC+lbdRkqhL9lA4Yz3xLuOnBDDhJs1CtA9fD1m4xJpt9RpzoULA9KpQ2c1ytv8Q63/VlvFRIq
nuEzQkUpKlokOoOkFhUnoej30xu4WkL3GkxtB5O9C3wXsHu7uRfnRZ+qa+eAZL3YFNwGLDIPOi67
KYljKdZI6ZgK6cqTQaubQHBMvUNU7K/pVwCicn9+H1QZSKyaoO5C2I+AVGbrZaHt+0IVVpFYlGeY
lE6RDoaSkM+8hrxrMwJg/U0/Uf9DHW5l7jD63ecC8uic6nRg10YmHqXHuWda56Z5XCh/NWBQgeob
Tc2L45m4R/iAWp+tdS76+CGdWEhqz7m0L2H3jZLNVfj+9aq0QTrseRYq34daNj20l2sJM1p7L6FA
nPiK5j87o8yrjDwUTDiGye2JV7DBuBJwuc14aPpVoBfNjuE9S/4t1L3c1FjEjUe7KxbH7SEe/ey6
fMptuBS5WKVetaB0QySVQjor901zlDpACpPY+m36uNmPWUwmXYbyV77KUPI3z9ZtsSXptmGi0FSL
ZbrJkD110CL5BtTUzH2Y+3UWoyPWV0eatvMn+DYVTIYpSzM5FxbR1rk+2yPvPHLypGT/eH29u3tQ
ooYIjM/eOKGTlHiejzD4P/tOCuvLjphmPN7gm+ec3uX8e4Pf1YeAXiS3njbsYTFO4iidjobDcBeA
hWI5P0RHTR6hdhebvlXQNZLf0ZWS4UMUcDqGUyHTcV68tHle8tzcUh9MnAwwdriV+nAy06wjuilu
B8mc42GNvRBGk/JckmEyRzaJj2sn4fDKdsxexGf6GOeqfCX0tOkNWggk3ii9MFHhWbU9cHRfTps6
seDqcKJh4WWykPmBZd5U5+//FCamFVC5YEiPNcKh+8reEysT418GIV9qbVEclymmBeS4Gcv1/AOV
ZIZkxL2+zSIwvNP64mM1bpqDoYyAEa9Lir3Skf7WhZfWUIRiykU2KdSOVLy2Xfofy0VP8FJd1imw
OcBrvGEk7iFGg13riovo1fuoXc7VdTpgeJumMhFlEJIYsKL5chnTp+MdgF4KKJEwrZZqbvpHS8Ra
ZSYme54TJLX9avB10nuhAVzk6mIre70jK0PgbwSNx8XgaXJVVGUEfVWxQNmNMvuF7VWd8/QQYaBr
5yz/ziyfOOKCWvxPWjUObb9RtnUK89oyz/nju2FRyl3Al5bz2bgc5kt0+Tn0hTq0pcfVvV50BzzZ
0TSrEr6X9jWK5vo2WvTszjQLTUKT/KCULlN7kz21d+Nie+QnID6jZCXYyKgVDYpTqIQJSqRaCTi/
J/YqhQpvzeEWX0CN3j/TWC7G36n9gccc2w/tKoviB+Km3DFXDHyceL1sThYy4La2xg2a4+n8Nav0
Vih7+XOuZeaXJ1p4exaP/7D6xptKOP8qSgItkOMtpKCE6PFEIAMlj6QGv/OxpiQkqoK1p0btUlHH
jaGvoXJSUxu8Xhq/gXLbS9r/SPYg24B2TaOAn69dSfjwDISbVf5k8ByI3IsrMtZFK018xsm2ho/j
60aXvf9Xm3+JcPE+xrxJ1+8yD4lEPll3bQP/LdpdiSG9EbD6DZt6ilzmMBPgkqp9fUw3JlDMgxL3
1HV/0fbuumSmNaElaHajYjxNK0qwkiYq68HkjHXtD+u4akzxHRFiGFVeXzyi7XKuIcd40fAViPcf
yDLs5vwr9VWdwABpX/iVJ+ltf5veHkavWZXnIAYfe+1tuFwyL+Zqdy/gcjpvFN5od2/bAfY9482f
400Ri/3XDjtm3U3aqoJ9pHzkmVX6C47ZmNML9tWYsZ+G5UPaqNSvqXnRzJx/eE4c/UQYyWW+hEMx
LLvIc2EM/LKjB7j+/U+PB3XiLWnvAoVAypMvsG8KK2OOuicM8/gHLSrebsV9Fr6Pw8CgBLzegiYZ
gSnTZ6kqH0ZnnirEXX9/+cDpJEA9qJ9a9ejlbw2h8IFMq86c4RXolrdEtV2yHcd/2OJAG1ZBCMS5
vV2xN41n/DdnE/Rp8k/V99f48QR9NxR12krX2/GQr5sKmazO/9dSNUT8dLvs3Lw9axdTTvqgutpM
LqG4orYcMNvA6Gb8y9hMUPJIOjXdS6WR08xAZUHsunaxDSE+Oia2lWqf3HFJXqoxgUrZKtiJSQP8
OahF9vwSCn/X5wwPOCK7kjYN5hR47iWzl3EeHzVE/dbWFDRyPNT+gQwZSCKQTPgxHqxVw75VWXMN
MvZEdcpXyekH+fLF/Q0rCEh7JgUYi21H+5SGCijsfE/gKl193qtGJWGcNcy3LSDgIG7/9b+cW7eY
WDsD0n6g3TRhPRzsWdWYuvhLefj/qP96TIcAdreXmSln19/DniDUzzoK4WWUz834AsCBFCMa/W8x
C8CAMcNFYQNhnmQTBRvkOwqKHz/bECyNw3k7qNSS1Xlk94gE1Zv3MGM3GVWXxVHr5EalWHesbgip
xK+Wof/EkynnS7dZXhMRL0THLUoKciaMOHejkp/iBq0/c+lNf9+5/JGoQnacg4YwsddvVW04OXK2
LdImPM15b9p+r2gCbD238MTVIHbb0p4tmEvxexObRFWxdZyXcOAPM/w7h2lb95HngI35IgJuBAmJ
I7mStZiqVP/FUOnn9Pxn65iPgzww7g3j6WxUd5aTgmjmXL4BZBkuGm0DkardepcB6jpSTt/OggAk
P+PEdsFmRhyIESkna/102P3NpDCrN4F8Q1PXBrqy2/PF33+778aetVQjgg71nObbFg93HuKoHIU9
6GuxNG7gLfl49JVTIZKrMmYu3iHPeTrTafGA9x99DRbYx+WlItiFnS+KkBzGKkCN45OWvBd+1QwI
UOzfIhIzhMNBNcChBzQNFIdwVGa0sTvmIP6gIgQx7YSp/qtbkrkYUWx7fMgW71B/TDXRJj2fF/RW
BC2scj78xFXUHm78OjuZrzrADN5jtEP7qr+wix52O1En7xszRaTHdi5aJfEZGnW/jEMGuMnMHE+D
NXWYfUDb3n1314Z0zaO/hHw0wP1By/NpBgaLLvzLkCQLWlQiyredLKBUFr105XRCivFSrSRzfz1e
TLajOCjmjaf6aKsBFpLWF9XEzfiBv3kaCmpyczLs87mH4f0eEqx8cPo3Tq1LcGETJ8GRFBE80NBa
lVMyRkgI7gfu507PWmLThIsyf3XdJHTsRDQFWBNhJLPtRhZ/zX6qJVLTj9202+zl2+xeFLCa0nbn
THc5JXC+Cf6uLQ5Es/6LRJqIZeze8Ho7P4iZTVsD+wrDQ004qbpFW0H0oBzvK8WbE/g1iEBx28XV
w7LwGsiMNLt4Ai73feL0byv+paeDYw7noCuBTihpDAWBuW1JF6Dr0Kw+aFtG5KNwdTyWO+LGtfbl
udoVsTQTK+couw6OyH49FZVih9yofKCk360d+Fi9SWNgcvjBDzT+bMQOe+hGmgHIftQB/IzlsUuO
1nIh6wnDY58CSY9FXQKpp4gOlRqYbmi/YXCCH/kHL4W/Q6noflmKIm6v7saKPtH5NO3RKRukpjr0
ujB5PZgLtbnvhZoz6xZdMdUDk7eodG9uz92QFLUm4lvNlcZQ8KKBkHFcJR4N4DGi7SNCPozcbZ6N
jetPcvn2Pwbvjy+JvdtLlufUAtesxPz7xyNMTVkCDt0upI7MGZw8MfMMzAw7Au4M6L6iwPDlLhsf
KCL8yJUljczJo8TmTiZaLvOGNO/XJoTb/fLu9pLQFIWbdwZa7lahZwa0c4WNdc8wAkrCEpGkuPLN
B8JDHC1kD0i7WoSnr9UfaWZ5vo7I1jUkvIqvPzaUSykYJw5WM8rtrdPDxXe/gzWVxH2uVY9ZFhJX
jcadcokmUa5M4ZVTd4DnYrwh8KMvzoj8F+bjFfj8BsHAUMU/3J4mxejBUTE3PNax5j1YO4s1lK2z
SRLn4i61ku0rRg+UF4Hzpe7wufA9uKKYwwxIhX6ehLDIDR9Fe1nRbORWlCpj3GP9++MxCA4jLza/
MRbkrB6Js7yXQ882oSSatq3mhqJa3XfXY1+MpVv3m9wgt2AsHWH8RfnFj5RRMhkJltab6GO90OfZ
29Tb0MXMVREf+0pBCV7Y9GBlhR/rJr/Z27oY6OXOhNUfEmHselXPTmj2OGIKU0TIVx8T3PXUZH/A
PCARFs53/JmhVZ+TzXGsDXS+YPeg1GX2FwMkmdWbfT7OEYRnjD7U86Fjjpv/NVpYh/srz3GOukh4
rZQxaTqijA+ne6jWpVR0DzR+PIAM7Pb56si9NZjikxoj0QcH3xx4luFREmryLoYyhR6b/2x1FoZb
m9ax7sHoKGx+EfM29GKhBjQz6c1xJqZ2SUDzRDAXQ+MD+eASE4YDpaRNZk7Jdt7uW63H5QYbAwBB
yUZc2VP+Kna7EJqvG9ZO9PQtqqR5rn4yChFfeb4P6/7VPaucgRxe3VaDHroKE1mUkT7Euz6MDWOL
BH6+Mnv3nuAoXC0BEpVy4g1d5YSrd6KaYuLuxcyRLX1p3Kwhc+kGWBWbxHIAZFv7ugW8Euym/lxL
1nqLI/9eXmItdKjji2RPcCP/xPokGs6076+VTImbW5cfRdA0IYVPzMXpq83vS1qWwTFIRLDG+4E/
DdfLvmuUlyL5A0z1XRfcRluY/Bt5Atc4rlqKOmAaI1cCK1TXERvIUcnx1FCyo9zX8jGUKT0MzkS9
Xmcepj4CID+StbSS4/pbBMlrIGtk9PTrSdOleoMby5U1QO08GLtJJHhgMmTD9AxCXZ3rTU9KlXeX
ASlstlAYwsKzciDesIwW8YtVAMx9MemL+I+0abY5keErYOXcTMOkqAw4+V6ib66nTHIt3RRDWH1T
Yutbvxkrb1YglZN8ZsTC83HXy8Gc3s049C12PiaiqNQ+HD7F1Z0T8Dn0agcN7uHcAQnRiXzVnaUs
a0s8FKyIaO1Ib7b5rh/FN6nu5j819+tj/cFyPT7/nJEQnU4ufWdZzEoR+6psfQ/zF4eIcfWUAcpC
APu/3qlXz6ajYBHeoouLMCdlRalx/3qzMTOEyxZm+AyqwNLHZPN7yJW0eWJFofnOQ7kQmvklIgTg
c4dN8Uc6KUPZk5mew0SDqa7pUUNstBhWwkN81tS50pZjSrZWL+mAHmkzoYRiHGAZGRpDEKvaCErj
CXdmf0vZxjj1tpHQplwmgKZzmORUtY6qiRm3x5txpXBAKJMNLH9h24v7LLOp9Wgb4Qi2pCghwuiw
Cz7emyLlt7O4i2fBJTYYofUrWLxYY14jTlpunJxqPWIqadPk9bIqTFc/52892mn1VBZN2nJyo9ty
AE0QP4BpGpVk1rkjtOVnIDPi8POYFMvzHuFqCzTQOfntbJFo/PMeHRl1l6Oc17r6G2VX7kqm5XQT
Wp/VotDKBUYmPTlrUbonhmo+xvHFs1QzPsmsIfoygZqkhIyYa7aVmW+D/Z93wsxnSPpqs0is9GPk
ipEhohpMmlNyqwjyRbGd5GPsoYB8q6N1Hak2xT0kGxh41Ua2FZQZKZsZL0H9KyOq9KD5kPH15KKD
Ulh9VjkFHFLrxwAhkV8LVC2miONAb42y+eOMBlvDmVr7w6sINbPRLRcqfswauBPaZmMr0s7ives2
oRUbiNhcXv8/XhCEG3jpGV503pQRKoIsf7lZdtkVCjqMVQMHKbaVYmyj6Ca9Lc2mX+3vRilvYNU+
hSoa4Q0BkWfqBEEfSuMVrTOe3iTiYYcEME5S8xkMOadDUJ562V1DON9Z68eVPOswDn6DPeuZzpeZ
M5ftljeRdCEQv+5bJnG5gmnzRoMmFIUbJBi7fRyEiAUZJJu9hK5rPksOo/tLsOWsKhKcCiQZQXAm
PKDiib9kROpi/5f/drfSN/t/OM3uTlsscDg8NidzXCvaiD7//d9sNBBPy+6h4lPFLv9CoTSfpfPE
a9KMqLugK+/m6Oql6JtYFR4VngZKZ4RZy1wApcS/jk/uqzum1arpwkGUXBfik5k6R82j4CdzICz6
2pS/Xn2NhGnlofapnjp1a8A+KbkilDPKEnHkQud/u/tjzCLypzWv3wJaAPDCVIZ/fu0nac0bdfzT
9rQJv3/+wBAapSU8uKSgKh+HgtcshgyTvHNsONN2Gzahfo3Qu7VdCOKCYgvGEkpkqiQcDx2xjj3t
W8LC34sDTAG8ZZxKUURIBumuFNnckbypbVLbUkzymuCLLp0RGkLWpV+qLXWOBK4JvtRM5U6W9UfS
Zmd/gW+HTlHccW3aFe6e7F+ILrbaIyNeG4voiTVOB1/7xVxDXUcQsTeDVYNhsmn16eQ+CIzkAvLE
auINnz09zuy57I0iFaPRcGavWvgWaZ6oJftol8nMXA/vALZwB4r1mH73oF/hXFdMbuI8x+FHO82n
w1TdqR4bZBuu7ia2H+WdkKzcAE61j5pKq/3Fr0w+IFuR5vvAn0nKMKl+LnhaYXaI7T1Jas9bUfo/
asiC/isaE2gsCSISbyByjb7QVN8Ekl26Xb20bZB5+E8RfosGsfKN6Otlbdq7TETvSJfB7p8pGWcm
BwOLDblt6Dk+6qBJHR6bpEDXTGyVIAFD2YU722JMiI8HXTaj6X6JboaTM31hb6X50T0BABpfMxjA
TNcm5N6ZCt8FJAAIz7h1PT8aAFIcDpGJ8/fsWc+DvvRkvf7py32l3X56kDv7Qw/R/OnKyOAz7mym
Q+uG6OEPkQa1VOQGu5h+LycUHBCNY77TkFkHEM4d9/UKEjfZDNo96yNLadIFrwEDl5h6OqtgfPW4
gMyfizO2rGseYo5kqYuh2ocGxqGajuN+otF5T/MLyXcEVIUSVK2PFAma+bA39FQXCS2JuzezokJV
OgJDvHCNh0MVl4nj13pytYRyJp+VmchuW8TXykufLwnZmtHS8eRguIhor2oc4IiYoJC/3uNiYFgs
ff30vGkcRZQUcggcXN69krS1LmGmGkxBcINZg3z7dja+/ki+up9fdybSS1vLZVW9MezMP0de9BDx
zmvHXWsOIbMnxkSa5Tah4g27EmHSCiuN9vTUOJfT3DZ+vVAFMZAjzseyAvjszsai4iAQ1fdAta32
DSTm4IBOSVvhaE0mJmq4dB0gJVsut/RXGYuu7W1Xgt8dwWIWHqhbokA1AysLw4pyOJOx6AzhHrGM
pQpqsM7PxO0zzdDPDkC7JmCJhI5whRK8CrUEKTk/KKz98mZSbm5SIUqdUFRC2x4Q21Q9YT99SRyN
iwy1TPOsjBAzpi1peFRG4DYAsdrA8oca39QL66GixK/CdaAavwVGc1B38pfjESvgcHXDWtxlJms7
F8J0UP8sbGqSFU2emyCHTakQJEWZVYEQx5ltyZqIaa8jVUZG8xVxHyck1qDUuCA1B8MwatbXyI7e
578D2uy0mwHNqPqcFql1sUCVDU5ZvASu39jiggocqHb2phrosCPsKM3Gyw5WH4I7ulbc/VhXI8y6
yoKUf13RuiVwvCKkQpBI/E1oMmjkk6Sgta/UFOADZfq7TLBltoM6PBLcg5LZI6liFV3QB66dqjbW
qy/Oh06BykhVLjESKs0bNb2Vv74OJjHvPMDmh6IxC/kNxTue8VX58sjuTIjZJmsiXXkyogCe5qcG
4NNiVZRGANFq3wnjo4UCLuJ5gPbnrGC2ArWWtNSFv+IQtSbG55JK6KJBb7/qKVc1dQN4E6AxlIAW
h83mtCygJoDxXBkdlXNa99GmngkzoOzPSvJMeerXjsGiDzGwQmkutgynrCe9sOOhZtTQwC1L2NY9
BKbg2OYILxy8uxNGoArWhA7oJ6RopbZN9SxJcU4Ojv+X6BcRuOJaFbm8MTpWIfV7JsyRLr2F3nM7
YRvAPp1coSq+td9HKlXF9JizI1EgBLOjAw8dP8EtpxzSIgN0KECF4gdaLh8vkk2WjPi5UQcM4L//
vjepXtSlcayjRBrLFsjk4+OZjwr/pJqlQBGyF46gW2cy4gwCCnz7RNgUn/ojl+l3R2cjwC8jepIu
o/1JDzwKzjmwrfPidDB1bTeRdvZG4TA+ydzs/ZF2TGHO0tdRs4wfpXeSRpfvuBvk4PTNzFeuRZQi
aaUQu1trXiiaOlgj+Pmi4enmNkQvROMzNhlGyU8aPoVTJ341y9YfWtfSkU3y79tc/Dh/zfxAK9/r
teTb9XfjDRS2PbERJMfCuiZptMo6IlBd43u+IwHHnpxw5EsHu0BlVtIbGM5vo+Epamt6ItjD+LuA
Wzh+k9mPsR7yje0+HjFEL4GwIZLh/Mh2fzlpDShfyqo0GigsgO4Hj/e8IxpJiruSWsHi/fXIbGjy
ox7LQTPZLJ+qAlBsIScO1gIykaSE3lyhdEhuwXF1/fNA8A4sME7+DlrxDnJHGzkXylpAfmepvF9w
G5DmUuO2mYJxGDRJMHddaeCH1qIOpfK3iWh+Tpsmlu3yWJ1MbR1hLwjAXYgNfVn/TSMT/sNflPWv
pwmMl3TuCN71srZd/m2UZt0oomJEHyOMvDjviQYNOQTPCXhg93rsQxgbiwk42sKA1hrmISk0q0li
k3AsIM4GntpmXom07zS62BPGrONLDbH0u4G4YnK1eRAz3XKDIqQBkHXnwPdducSjX/4UAIKjb4Ew
+gX8uqEt+lvyilj2eM0a8i1YAZMEilSDqMpcgiEpNyt6K8Q/Z+0cPzjMGG41NMYi9U3xfnF5ZniH
diRJ8BJbIZwOXyQ6IC2vXQTIwS2DNAZNnT8lqJRcrZjzpr00xZpyTH4b1UJpwaQfmcigjf7O90zq
T2lbRB7kJ0P2cA4EeWdMfXnr8JPNGWcTtI7pCv8sggqOL/N99/s00cpcHtXBsD/Pqv+Htlob0PI5
JRTLjwEqlwtkyY86fZm3WXcprPQV/VZg03HcAaakljvoWM7CfWdknvImK3yKVzCE5LnUo9KLyRpd
J3Uc667DAfs1axw74iGG6Hz0RQvNi9nhQ/yt0Mc0E0e+wd1fdTjqP4EPTahzCLQOi3rJuzVmFRnH
jmArtjNBvS8i2M+Ri9f2kfT/WxnPHhy5BWLfptIg9fGMQ7sfN4QX8isjSOPkfNfyQXYrXsYt9yq8
rb1UwMiGsh1vCu5L3t3iBT3NgVwfZinHZMzUohDXwc6a6et39MHyxkEad81iQ3UHQd1eKno/1ZkS
ytMuQSc9uPjCA4jtwKvwfmGWTm8hNjPLe/06SW5MuwK71py+yqTaByYWpngI8zbye1zmD1CND2Cy
lQcNaJJksJ/1xYBL3tqsMo06sRA0l+pK7ZajmctR6o8cQ4heeGs4LtIjfg2Zf+y0yWzDSVNTgeZY
OxIqdOme+EzcKKzuVB+5wwJpICKKnamcVpXqHQvQcGIOtiveNoVgMj3TcfoIDnXrvy0BUTG/6pXm
txA9Q8W0yNDRIhItNsu1Tt4AdnSgUfL8iaPRBLcvpE2jostH4w+CQhjYagx7Lzasuh67duDFe/u0
a2mRP5dgsIHE2s3oJVlKtMW4LK5bkkk1LWAvrvuASWsjLH7A/J+UJBUEwxHPhM2KYZiy0xJQRwg8
CwZBihOCeJKHfRALZ9CbFUfTg1K6FoqZ0vkis2Lxm1yg2MO9aW/mBWfgJ9ry9EKNKjRc13jh0Eke
WZnmAEgd3cWzvze8vdq/WEG0KmUjzmPN3SU19uJFzyZwl5Qww6tOIFdMmSU6168LmSzk3VRjzhZ7
LzYORwtTT3TYuVAVGB5ruMmEj/9dIEPSq+TGk5+u3HqA/MkUkHHWJDd622RItXLygCBbb33NePWC
F6EA0ngqRsD9Ub1P2bT7m9hp3BA04FAhVbeXXzgbjN5Pyy4PqnVcDlSfW1Mdkm0WEitQKNRiQDH+
ZD+7VKgpA8HgFVec1DmNdFIxWkaQZeULrfIakb1Gvq0VkaZGYMV+rUKGlXKMlf42Eybsiqgz4fbV
ZDLSG2iP1SXoxmHsZ4l/tI3iEeK0tBCfW6NnAgvGIqQ8tp6j5UYBGlMQcXKCre/qBDMBstI6OXIK
KGMugEjZ3yaDOgyvYPzAVdlRqgrKAqiXUghtS+5k4HD2xhLruzzy3ayo2t9eHuDm5chvE7OqQAXt
Uec9fwrr47plBkHa2+hQcjDjUy0D9bx5RVIY3eNQGU35MZOwcb6qFZqXXz57a9QFp7JKCqsMx6yV
dBDAduWxENquk1+oS71lT1+fqYPiV28zZnH590svQ45gPM8HUn8smSUFWoOOlA/zy5iqc+fZ0gnY
OAPc1TXR6u/0+1jaF6KEcn6gyUawD/nDRH8c/UgTV3/W5uWc7HZyeK8p0Xgvr5ne56Zuh/ipCEFs
vALwrrPXGTcPb9ClAtQG/gIx496WT+Gwamu3Rvt2zzQ642Qf5GIpko7ZYEnl2JlEJKyZhGSl2PbL
mh72u1Gy+L+mtgu/GFH/wXOP2s5qVOPBiskbjwhbS0cu5iMJzbHFtBJBXuWHZX/m+7A12aR/8Idq
4J4/9u0CbyLtCKNsiPCZcAVEJT6Fw8Le93Oa1eEgGd1jrugZi17yp9VMBhlyk11A6Zokl/9mZXfV
ATp43Cy1GYPYo/+vpC1NYM+8uS4NNXEOr1/lrssk5Z/L6S6KAnne2XXVHDKACIEGUlhV5j9rMY/9
gGwzwxUhuUCvUZydA6lKVExWGfpgPenn77K+9ehVBiShRNY/tIC85MyYk/c9C2NiUO6nUx57cJcd
n89tHiV24jYVBE/Pu1CziMDK0z8EkLwax5fB1rB2vL+jKy9BaRHUR8iZm46Rj1bGBNhLv56ZTr+g
C2OdoVsVSaeSvCUS89CDGGcfgZ8o1ZLNxa/AsthVgZFz8WNJk0XRZa9bRtOMV9nhFFZjQA3rf1ae
r2yhyonI/wvNWPjLDM2/KLOwuYPsxQcCxSokwVQ8DpIspcyb5Jvc+HyjL15Bii7HilWtmHAIRUi1
6acFUdzo5e30jQ1UNG//52igI1qnMmTc54QNiFFYhmmS+TaDOFXDQF5rnZNdOIm4RD0HMjDs5Jov
62JlxwMLwjSpiSLcJoa4YeuxCldNJqivDkALnVguTNxXXRFj11pNlNcMXhSuHHCgVJSyrBubOqbh
pUqdJIzR1F/BcQ4fdsxBCs8FFkKiCOwFJIzXkWt1qOOq+/AL9rgvuWLuRJWIOpzdYugrxbEZ29iH
DEVvUfgYppbOFlZAq29tNAFdtJYCHbNLSeMCMCPQK1PFI2UKBdjLnxGid1NNMkTW+PTWeoHClikR
ZVq+u54AHzIBfJZ7onXDw6rb/5aQzB1LCUoeCetqu9jwv0/AdQe7NtZRjM6zcDYZiReZy52uKlHR
hoD1pd/i/7z2aPqvAvtLDpy8IeV4oRhcYfxQWL7U8xJWInwTcwfFkGsOLcY31xvZ041lTpYqlWIz
wKBEYvqya1WYghCClwps+4tSrHOUMYSfPuFQR8/XhQBAnyyoq7/4mqIgFfU1PVtxfb6KMsspWLJm
po8nwe0bwKKaLv+Cy6q1V+7oZoxvX/7y+tEiEEIMWVnMVo5bIxKkyMSl5Fn4IgnUzjpHkaJMCzj/
Z81muZZRzMvaiOyNMlicwHMTCHCemOnIKcmC6Byib/7PCf8xvH8zAmQqRRR1FitK/5WmF7qhtBK2
BUZRwJtUl1OwmoiTN3QfGWiEGOCaaXX7xH7zmPyxrJGCzizBSncVs6acaKcDUQeBJxz2v+/W5slc
rX76UjKMPMQ+iw0G/E3mhWQndAZA/0p5m8HfMLbORPgn8ymNF6ydASxkeEjiWOdKRO7qq0TN3OcC
Sjqu0qfm9HZ3hmNjE7u3xh05UQ0kbz0Q1rGN8JOXYhzeo0G0zU9Ox8TNNDQHoT4MS4gQ19LKiXA1
Ddu1TbspOzQQs8y6KBOhtrL5wdHI1dbvig0prexFYr/GvZp9DanEDLvn/HHGFtNRPzfiIMXUJmEg
TZwIWeliwCjw0iUZdenO1w2MlV9OntZGBTXMXLv3YZzEuw1SFsMJiiKSOaEeRJdZephQAbaq39E8
TkFS9Zuv5cGNbImwpmLWna9rQ/bqGQR2PUHwEH8woZP8UxlWeJGDGRj4KlTFnOmscgfpsJGgen/w
ZtBemODzvDY2ulX5nvlAuE0ZS0m7KRt/tvOnPSrk2cvr90LR7FecBxmWKYYCukFenV+38njcFcS/
qSvflJ1E/6NNP6HRjd/2nuqTY/aX0XjgApcz9ldSpeB+ZDIgS2WB1NZZ2pJA2vZ1ageKpyVZwNMo
Z3R164N/NMmoSL0pchR9FmmOo+F7qXumR99oT0C0mt2BdRAjFo7x3X8CTbHLAH+lwOMhz9YoE+VZ
CQFNcDVLqvXLMWPeWfgKtsPapoCpjnWRyKM46yD3UBfIZb0kP4x+7LyNe8Ja7NVJetd0B6qIVfNA
VdpSHSaEk+ik152ptXyv6zUvm2IIb2DeA/DALca6R3aoQLSO63k7Ob/73OuXXu4DfaccAVNksXHl
41scNiTngT5Dweb4D9XFR+b9tHzySpmayP+EdSvAaNK2saWIzpDLvNPCTGsvx3yjYrn0rBcXGn+m
hz6+iVVU/ipIerEXQpPaP8hh7P7Svz1ffKpjief3HRqJFCTRHqhXf60sW0syXm0Oki+fU94/C3z0
sSnP2BOdcDapDkk4oYEIAStGk393MIAHEDH5tFEDt4Wap9B4JPiLPJxms4VcPWMpOv8WZgSBdiWf
5Ik4Z+a0BgQnEtDLiAaq8dkA8TXRTxqFoedrjGT+9U/M7cP+cuV19ra0xTzVEnmJ/ti/69PeC7Or
c70r5Y8KGNx16eLcbiKEoDOkKcq9bMdpHkQORG6rBUFni+wY6SkzqogfLbucAFyeyAI50rzZqw7a
97evX6tIFyGJCanrF2395L1v1P5HFCVw8mGe5j9vuf36E5hOSyHUhlMDyPm2BL3AcE59czWl+dso
QitPiM7zn2S1EzbJurtttB6X3BhRU55a2hk9Mr28lOp38dUVriurIzP0ZWLhgkwP0a6AlR/wsoqB
yD/3un8GaVmhOEvGj0A553qSHsrMEHtqiuR9+6sUZO8D5pIJZ1/h3sD4JhHBs4CGLCOxiEpuugZs
kPjP00lCJcDBe4tDRkEVNsr+gqxEUn0oGB5Bd9+eczUtl8vErNuLYJ2jDSVrrfhLt7dK6p1vhK99
4a8BcrvODpZjthp0SYrDATEbheU8yGVne5WxBMkKk/C+auv4TjqD2zNCD0wnvKPXOaA496kWABAH
O440/GZ/aNVdyt5CNNvle9+beI5qnQJ8lIZXrOW9QJMz8c/Vk/+L56ueKjmTobIUsqBoLnf+X0o6
tPPtmayzkBXm4y2MNH4AkQgb0ngMgcyqFStXFiYJaFigTYgQfCPwOcX3lbj0IG6z5lebrneqOrtu
plN1oMwjD/Zs1qJrPOk1zfpLvXd3nk4GFZbCwPFQozB12eN9vBiROB3cwo04b+V+bBb9wePmUING
eJqto5JGTu108xysJkcntjmX/loXHpBi5z5cfaxiGZhqR4Kwf6fvGbOfUYUv5MlyFxafB7KP91ZX
e47MAw3/odD+oAOuN01VEfVYeUeHorRv6POYIoUQjEK5CUpefVQCNBmfgCi6bHGP6AZXXVvExBAK
s2CUt+pVMusbautVl0ZffjIEF67QeTZ382oDj8uDInclu8AR11rRqBJP66qdmBA/UdJt49G5Fs9W
Fpx2fYanYqlUe1tKw1XSTJmHqocQ4O1x4rrS+aUCpjipX1qwhPmbbbzWF115J+TL/SPVGktgqx07
Tf+oaYKmvy5HpL6mbabcEmn9X1IvERd1WGINK7oyx+V96zMVQ2sd0XEOSTt1FfMssUBzTiK+b5JK
2Xi9rjyP/AV7Al0jP1S2ewv9ov3XrGTFi54faapoIhhlR0Wr/uPwCwkcHJVD1XBKgwcn5O9PBxR3
EaTXTkadMw67UZmvkWyAmyggmcXsVpAzoq3RE3NrjK7gBciOOzzAYoXwXxC6QB/IMiFoT5EMCCBh
FdV8kYLyyXpkwp1l/RFMQQwlokiNwi+QUySl/m7z6H6mULWC+yaVbpGLIzcOtu/OpY9F14t1WY/1
l+rtojJNXDmuEGJOfXrRETOroSg61VV1PXf9cEuGfWwTa66ly03HzNmlIZ/F6kYZ4UG6MUXJ2OO8
/P647VVHUSd/4lyBEY2rtlxv10MY03rmWfSnn+4B/wtHh47dk08+WgZeoYwPQmmk02Vt1Ja79C90
9NGJfhiGzbC8KfwuvowRrHvWiNcmHswN5g4xUJcIjy1MI8MB9sv5gpl7Dd22qBwVhtiaMT9icdmD
vo8C94V8FMS0LlU97W2gGoetjd946k00vo/8Q1z6zdQloiGw5D7BPtvcrYn5oSwkApVcLQ6pKKht
c0RRew9XAbb5YH499aUdsc3MKi+nFYC1rNjcHuTcfafw07vRstLoWDxBNcO47j6PFELZTrU1H3Yo
hSdDd3Y3T/EUsGCH0Ctwrj37RHihSJEz2/60npFDjZuVLu+jHz3Juq6Bso5XDquzc2TVsauzcabe
sxRTJUxf15mdOqdQ4gszVRuWQDvYqVxNTxzwRna1OqepOTz3ueiFRNlt1LNVOCCcTlcFAjzfUv7O
b175NzfZz7s5NuYB/vXnIm2ctgkyTjT80tEl/NFDrTr4fx2E3ERoxMT76uktzOc5LfUG6zmveXK+
n0PnwQbs+K6FNRhrkFlR1l2Zj2h/1iha7JjjRW4vZhmAFCROrZOR+lWzP3ZlZheg3TnTvNEecPCt
WcS00vIK5/VdhxcE6pQNQky+5Ic7q1Uw9E1bGNb19zApWL7zkl4jtSiHIWJ1cFYpEPLn6OQubFm0
JBxUB/hCZkEtgiXE2K57wVuPynkUnJ3ybXqCgVJuX8IxGPrGUIB7AFCVbWo9j6RUVZH0oMOak5bE
Ux+DpU8hIXqm6ZREOXUtpxPypKwSGau4hLet8MTEbSn5OC2KpGdAXhqjpau5C2Dt7WoQrQ2KDrcK
8YAsTgMF9FZTPnhLCm2+glXS9oG0yIQwGhhYmFEPwwhw+SFWZHfufojOVj53KJp+46YV5bjtYVdd
eW0apxXog4doxEshWlyFsg5eoYWTg3FDqyGhJ1KKhsuch9eam9Nk1F3HXJyNE+FBhUwGv/CG8Idy
vvOYdd8RURuyBmeVVnNvXGmMRWxfkExrvdlo/n6D1NQG2eQukE1l3lUJ1WA527evtzoSgH4OuZI4
fJrf/Ad+CHRlUrDJr02WMoBDrDk1zSAHClru7PnD0y80qsUr+C6BrsP6Qkb8zRG/82dphtLFw9G6
EmgeArf4lZirvr90TF+tbFPa+sgUP8EPKwwUykU6vjmy63+MePmJxvZ2kxSXro57XKzvyHHRpSux
lEzsCdn4eGWRqgz1fQ94J7H/VezoVTrlFmk1Bu7/VcTBMvTgje/prv2FNdjCnVHWNOFa/UeDc0uv
f3Tfz8V4BC+HPAaCQzr51CBk2QOmpPyfm57py1tJ5tME51aNQpq6EIyEAMg2DGv8e72vhrDpFsa5
CpSVLrWvTwbkiY5s9yesHw83SLPLXusMRQGoY/J+NmnQ5PNiV6J4u8nrZnCsIM5nSm1s8K4C840Y
UwqAalQ84cfmX+rJ7q+v8iE06ZTN3DwqOeUsTsLspO9hjfBAI4ZRGwHL80EO2AGiEloIJRRdsy69
dDX9cm7wqjA9YZNiuscxLjh75nClMc9cmvqvH4ovO6PAD2L21GpF/OPxwqbYtE9wQX5CJn+0z/9e
aOkgT9snA6kSoF2BFIqmivBlGxR5hHK3ztLyRRXLw6Jyk0QdCmlVNgR8dSd/aT1NDtvBPpsUdmxJ
5ayUjVMPUl7YktLXYGPsyG0qExpUURqk7IklZR5AXKzleSvwjLB0mnknASxydah+Oedz9J6EzXhv
1LqQixodsmhaMaqQsg9DUExHjUf3jGpra4laf2cBv3VnTzY5a4me5G87rDm6PLe9OSb6ASQRb+xg
DAuoU/6Xu0dBPI8RO7XjbFIF/3H4ERtyrHH/WrupBKu7962MvqQ9SwzklN7ddxKBbE/3Roy0rWFI
7MnC5oPkkTKQWpAkNYNZ9VuqqMwxq3WxSWV2UnQawi9KvEL9nEdwWcSahihIfDwJds/VeH6KafIN
7cLUpTHTkPHpzm7d5I0ZemksNgtP10oWgLZVWgtxzIwZz5weRjWY5ih27dyS5mhr+mtDVq4q/woL
Xly+QdyqGsa9a2SQBFx5iga2wtBtipVKMcOfdR4I/3FyMMpU4R6eyUyndK7UCW48SFhKtAwot+rz
o5zM0bIggp91sSSPxVwptxJHVFkej8kTEJujlvKRjuhNmAx44q91jKTwSiyjXvn9Kyvugh2KQznf
D+kjC2Qsfp9YuMt4QRFCjYxvOtDmP2H1turJctcyaOp/5F+TOfGSFmNYiRaZtCX94+6g4E7IgCwO
JBJ2Iykmnrsk2SMWzhyMXv/H8XbEDcWIOXH0meqq+kGtMQ11XqRnRCPy1xa0H5OjJwvfQZ2ZFA/h
+6r1T4FdwqfHoEICnxDu8fUIEWqX+kQG1TYyWyhHhH8ciaB5JrfzIDtkKSdM6ByHqW3oQVTTdZFZ
dPFeztSw05UgjvcJNuUNOMggVRLWWlyUM60I1SRodKb0060IC8vqAdxOO0waoM/AkQdRHjgQzvvB
v3gCiWDrN0ewEEzy6Tr2GMC/iz5AEZ2y0E3plOl7LOWhYHA28athdbWpmMMSUvF0VDbjy06/k3Ml
CKtYckL+tkHZZF3KUUq7Ab74kvUbWqxIsDhPXaVXcb3c5+inFR8DiBo7ASET5W33ZLJmao1qydx4
FVhtUDDi6MvYK99E+zQs+QER0wOSuZNqLNd+AlPifODCP2yKbHRhoAjZVLDtotIPtnXQpTJ8sA3C
JYep0yvBpCJbC7+zizp3eCpoQEanbmsLRkL/vU8y9Xn0pjq4AgP49tpzJu4OL7suIsGC3AaSKAGW
7OnPF5EotK2j4X5W4MReS01CmoEf4Gr/KH1JXq1ZaDNRx9PNIRFrorVHkIuSFFxQqRPEPOCZP+mP
kf/arE+8GQaEcOczRsuv4m6uBui0vjUZtn4qV32hNxnmNhVBMPZSnRqb2NI4+mv1k4U3+LC2KuIk
D0tOwNYMWuAdoz5MBomPtLCRtNPGF4z0XtK0NUfAwOG/MCH16nGcFEvOpDT+BZugA7FdFN7+d/gH
wnYc/CI+girN4tsK1Pao/F6bxoq9aMrMkv7BfKtgCUlBMCguJ2VTJScwMD1Jr74rwaxXBNb964qR
dNqrR3rn+067SrEdRfvExay2qFARHUIsyvv1G5Y17cXsl7jxe0Q8nEKxnXncTpug7G0UVQmbVPp2
C4BlkWUt6vi2aYNr7XNFf/OsTmwLJ9sOK+GFgZaDzEOvTJnEgMKt+tsEn1XST17cE8yTowv9fQ4L
Nvc3J2itlVnSlDIZnOe2QuPzlbTuGNkD6ToKHOgv+PoqP9AF4a704EQHOpFDXHt6GZCaB7cA/R6i
R+MshxMKnVpomEecTHOlnSeIbT3w17585pavDt+2AphnVn3EACy1mMYkVQtAsSfnpk2LZtRp3hWF
yDcQKJXHGUXv0H8UYcnlT+1xsXIVU/fiH8kWor0zuC2BYBVIZLEE2b18BlQe4TBJFGRSDPhoj7+z
oJoYnveZXnoWR5lvwFRuUheZjJc1/NxrYSH6j0FBD3m1RxVl95dA0aofmLGXD6VLUQSupXojZvmG
SLWxqn/9QT3gUGZQ/c30XusxtQjS/EqO2B4+S914qdjkR/v5fBsdMSdm85Z69tCTiBeHwogBPPul
Xk/4N8Z0ypCdhjfXyVU14wz8+qgZpAr9Pk6gWhK2CyTlPk9Suk7rPpw0UK+8Zf04FSEN/O068ut7
0AxC0ISMvioP+fnlxmtZmXUWIsKQhHksvnpP9z9hYPauyPA3uLKg9Hn9VxVExHFhh47YN7RRbPjj
EiIPCBNb5eVaOG2MM8wU6sswnNDnFwZCDjPKFsxQnlgkOWks2sXfGpX7eY1shW9SKuUFTYDTru59
1vYOROl1etxmZcrgXb7vQfIx3UAo6I9lwbEO1qDOztdvKIfNeLb/gB7e9P6hHWzdYT6WUkQD4Tp9
ZXbvEuHlveKJ3DOpZfKhPLWsr9QNTpVRc645AX29By9GSLJDw7UGMxHXGyVCDlQzIXTApzUYpOEe
tnKwycXP7yHW6nxhw/p0b7TV8RV+2IZP3MBBWfROtO8zCj3HocGmDn4nkZscDMKSfd9zuhtLtT+M
X8n7PAzXcMarlzVYm2ciaAs4nb5fPB8dU1S76pYJHQJnYjZYzaoBhtXjvzYqWJRHdlxSKynrWuwb
iIC3sAmsuIJFYa0dTsW4UOR91vs80CKK2up3Wrloc1IlxvRhc6naJOcxfruUXLAToMkeRLjDETln
AXvpNFrfKMRsNxcbEhSLOPSbTiGqYLT0gy/+FTELOegbUUBUlps8KX3tMMeh9gEopJeoEo8tK8Qk
gSNfDcx9aGYRa7RKjxXaLX/o4VtOH2vvYQ5RjYDiH/QiEacWokvpVhgAvnz5cgS/XUjNMPAqri1+
FkNe8e3zhC+usCz0IRJT3UYc64rhoaa+z9+ZF+DCPyJZE49kJnvqxwXU+3bD0tOD1Mp3HJVJWsOB
2PcD/672OYAkcgieEq6DLjVXXivqAqAHdWD9SDWAdO2Lz5P7xSUVJfZmjBs8PSfLUt1CMCgCFJWy
0gaBlK4yW3qmYCjSZ2grwMUh5jCyLuouISIBdaAQ663p2M0AKupDz8u5fKh/ap4B5UQEvvJ+H2RV
1n2hxhSBwjwVAQKFw3vxYrK/hy71zXILiShTKJeV+eIy5KmrE8zGVmwIwBiTiTZgMmkhkLGpC2bQ
kiadCEiM8EHibMupKEdE7ylbtzA0NxhHfISop45+IfbOHDm3z/i+nknw2og0WTX/l1nId5VcvemJ
tfrvIrxlclPl/Gdb1Ho+PLNZJHNuWIFKsNfG/NDartHcRI/nb+FHQtwQEqt8yfQK0fbG2gzeP/HL
93Oe5DRVf+ApFhAZjM8rUx8FlamX0ufxjsUC8KJGdmM4prGiAEVayJaU9l38kOUIdCH6TPf+iXr3
CWsRCDxCG613Mk+0WYHT6kdUH0fLZOaq+u/FtgyDPzBePBYiZxk6C8Re6H3MfkpofpfDtmOoQ0pl
B0ZvAABRL6et7GW6znDyZ1LW06DQ9GaeXZD/KkpKwXE+SAmMlySzr2IobHMerYeTo5dRY8tfCyTU
XAikdtJArI8SH3V1RKCqpyNDczNmS4DSFtkyl2lb1EGJhP0C6zoGb0U7N2OF2LRk1CHvYc6qzkTO
u26bLnxnauIKLqOtnS6f7WsMso00iG97R19wshP1GVY0QIZ9+jNSN6xIkVs7DoFZouEz8myKqGVw
QZ3H5GRM32j+QJHGDXXPapYaq3b4i100sq4QctCf/7Recs2VN0ze5xYqsrCoXZUK9InJ7dUiyUun
d5GImE7lwqn2q7NvrOkIANtwJWXi+TkG9tu9pFIhQq/TjgWeUViEw/is0jhFZIzarvfRkucLg5wp
my8pOOxqQCd+abyqOV3FucgrlJmWTKoFLVXaYaeuVeMsnfx6J6q/HNJb82t8+RHexrz44B1WwQs7
rz02YaX6Rz6M3ihsBiuJ6PFuRh3yKuAVyLimEiOxz7b/1xiwJM8KUa3fuhJ4n+SNaPDZ0yfFi8Bx
/3wqSotlMbJZfUTIPZNYO14AU9+HJwtLeegh9rW/LMMm7jfJsU4I5f5BumA9bQ7KhsaV/zYyp7Ws
hM7SsEgHD0+bp1H/IEXJ5dhS3xisgV6F9Aaf8pvUa8uGsnZpULP/b4IcXnSqT35XaMcwS20FplSr
KDN+6LZ2ZfSbXIWVNII4X9YKs4eTul6jfj4MgfG/npyQ08DRfK7Mm3d0kFMTAJf+nzw9RIkE8cMb
kjHLqB02hlmdPfcaBIc6WzdtFXVgJuFNc5cRllYxqbUaKHwNz31XYSYQ5ln+jUM+uf++nV89pXX5
kFe4nc/kqGGHY+Eh7901lbIAjNhoVF1sHgk4HPi4CTH9HuzXJJ2369GUgv8ZVAvZBgAWBNRxJHzR
h83fKn31Ud5BAw2CK/55yh+Td2HoRbQajN4EBH8/bQ9/d/A9+fHdh//m5DPgmFD03KpNuthiCjPJ
wxA8/ufY59vSzNY+v9WMVDnPZLy6ImJkUJVesw1d4QenWVZTYQCEC0tlrYCW+xsW0qfgH5y9wIhW
m7yB8RQAwgYCHhgXkgeDxDsDDr1GJst4yVBnuspKTCDe3347F+mC/bmg5uuOaqRrs+lIRCefdhdS
DPAVWdtl7Sdm1G0/Vt08x330ZRCxkj3EGta5s+eoy4B5hnAn+B/uIUC9JLo2U88TKUNdKLg4CXMj
pYw0gDMi3g9KSiVoniD2qyv+0T6wp/T4G1jFCoAH5zVyqCBzkiKmxKv4+u2WmEDq8SGduWzvOzY1
kLmaLmHg9YbBtwnMmil/pxRDRTb/O3gBVPkmtGnp6X9s7Pb3jU7eNwFQH6GpAL2Uw5lKFZuHonB4
MengcOAnb6Q7OXFDz+M7l0EiyExEMvTCoYOuCEZ1lMdWKn52vm2vJoq/isBdJ7kR4Brx9p9HUHi+
2waMaG3phakeykAH+YtW+8AiWpW56a3/TiA/LvIOXVEjD/FloZa8g9HGaO5dr9egbXHv6PTcXACg
P5eJ9WqXLA3dNnV7IvUZwVzMb0BLLCaC9MzikZHdSpb4vhmNc2nItRDoi9ZN06AChW64HHYRUVof
RXuEhwesWUlCzIIu2/t1U2xY45/HVJGzJkzjhcRZYkEvBDta/QlWUEkARCN4VJvP+maP8I1rZW/I
H8FaW/hASF4yPJC9hRZ0nWRqnDcfuADE2gxnD+NTkO0btep2yAVmeGaGZ6dcIBI/yL07cs1Bck06
ruae1TLedMm799qoi8r4nVckm6F5lxUsceTMYMOnRLl7BRogaSkZwqwJGV6CHLDT6/qdFdPODXk3
IZh7ErFYRgdq2X/ukH3klsX46b42kr4/t2LNB7QwyWK+5M2vZ9CLVkS+dOezk9bNtYU3lD1adgBR
7QRbO0+k9wyUmDE9VBCyq0J6ggNkTQdMnk5GXNtzXmf16OUf5g6k3MtZ4gMfEAcU6ZDp3hRpnbnQ
uP+AiOmc9raYiYI7zW3x7x2zVRP8KsW98M9mmVlgDOEk8UXUz8pbJYAlBdMYYsfxrEJE8ceZ0+xa
tn+c4WMJUrBiKWnWZp/Ts60WX5ngTuxWUHjmiC13d0bhrpZ7Qf6XlvwsiBs+jRP9oEtaTw/RBRyq
JK87waRA04mb1NEIG9ThoNSiavuhyhz+FxTJtucxlaVIwjra3g7UL13TJauq88xlRmTGlTr7LeAa
kswORrdtQY++5+Oej6ApOqNAK92reqSn2BvfMpcgtMR6N6M65F2SfLkkZIVDOkPvGJiiqt5+42Zd
R1yOkJ0OhXC4eNz2aX2QbapeMWcQnMocJ2GtbWmxZMEgXEMzyBgpz8HTCVuzXsfx3I/d4CRzNd6V
asoznzzv2+cs2wdNiuGL/qFqZYZ630mThtp6w05toNV3PyuXMXblbQSvH1HThEEphxFsS1q4FlPO
VKX/jHhBqW5LZCCOvIlHzdQkTdIPT65PtSon+ZymYZ7Uc+tmxgFUjF7Skk3ZiIIRzNEMNuUNvkFe
XSNFAH+FbRssWpHkc4cadvXWAjypArKeEzWnSYcGuf6ZFDLYqNfKIjr9axXrajYhLxFmx7jFQ9ed
Hb5Byn7TQWFUt6b9e2FGiLUPld/t4a2MSErB9qFbF2UUBoXT1Kk/+QMJJn771g6qiHQ/qLkDlR1L
pO3G+rNWw8FJAkBpzcJ//m6BP7nmhWhZBHrn9guNSCMBiT10MHWpSVCOd5oAPq5qS/o71jDbZYS2
pRhCU2HwST/um+o7Bt1Dy1gKnG5lX6G1zyIVS6GTbdy7/q6H1AMN5n3HUui+N8GxKje2bPe1I50c
bTEp3x33zbQs66R8b3J/2z32U9SwREkgNAOfPB8mY9BAt7WE5VX9gt5WKpNAkVbzOUqYZ8+lhmFD
Ov8PYXaKCuZ26sK47KE0HkfXq84H3uXQLya+FSGWFB9scHBuTffUsk5zTb9SoLg1uQWUM+2MlaCW
JOjWQj781LY718Xi6cyhKWqbAo80WZ8sMSk62tQdGpM6UhGgrIMN2hQYYYBgAzvDUu7OSq1ejc/G
PRi5fPKdW0ktS1DkrcLYzMAX+6ciO3GQ6cdwus5LnedjdKAQQhyxL7O/2AgKhP8SYy5cUsYwZdyj
b+xfzz80XFvR5K7QZ5F96jAQU+V1Yt/Vfg1bpaIP/C9hAVSGVBi5pCgoNTMfzo3CVrgIo6b3S1uA
bsNIAUajKeKfp88kvxj3OPMgIFtGw1C1DEGbc9M/qVaztzEx8jpQZHXSz+TZvbKHQ8AEK81P0I9Y
6WXcchQog/g/VN2EGuv+4GhM4VVGao2JFC9/S021ObMjJB13Og7LOs1g506UwbNMfkM/eVoe/80Y
JeHo/Aom/GavyrlbdO+037RPcdsB3ZFvyRgNMz6zbByFJVE18kcSZ9HhZpdDH5veB0Sc7nQptzpr
V9cW07UZmdGGMTrctNllrgoAQ7Q73HNoT9XL8zY2ZpUsE7RJIKM7hp+BYYIK6X23HpRkqHeUHr5R
TVTIaY0ZJg9Gp1L6N4qnVlewxMCklxQwFR3Y+t+Z1mpbL6dTAUbk3IHqOZnk77bu+SyNLXS+Cuen
VwojgDt6U6yEXyGh0mJQRbEiBLSeJ2LKj/GtUvyUKjGUtaJ+IxTS6GO2Yum+XhNXEXXniAI9pYUx
gCpSvb8xKbm1mDciu+pL+9HWtcd3Zw1KRg+94GADNXOpIGMcKPfrvQGp7/K01Reut+eZ8X4/DicT
H3lIhlNLD6uDlrVEZsPY9kvb5F2leejgFjzFimW+CKuuSlhUytFSy8dte3/eetqSG2AamK2DWHaP
wSTVYm6d0Pys9dUZD8svV0j+/1RPAsxavHcF8fBh/Ndtt/Nyhf0snb0kByt6UeqT7MG7gVPCdqqF
FW1f2ZES6OJVZk26vhvljUekPG8rHJrwoVtq6fcDxS30UWHbUdGcp60PZG0d3tL6PNBjgo+EkLuc
SUDG67MgkDQk/VzwYCq3oc3FphnFoy3NeFZjstmBFuefiVgzkFKDxydk6EwBIINd0eu5QfbbwllX
JiRfRz8yHhxJabH61BUTOh4OeSVoDUmrOAMI2dhtqyl7b0ZGDDpPuIkHgRW+4NiIwUK//lkhxj7T
WsBrcESmkq8qyg29LmVNPuuaAb6jEmBy4sEQeh6A9QJpfaHduHpbi7az0slpl1NcH7NXL1/EVTff
XGsMewDkN7B/nDhozOX8pNRjEXyQuVVJR9iG2QElnh9ETKrxph9INUUAhYWRpS+XNYA2mYoaRwnf
qfssi8NR2MtI8rimEE4r7pZ3FHKtYzTYK0RZ8AhxHQkoEfH+xbLOajVY2YkcLwRuldc5UmFgJfYW
as/itBgKZx0F36GrdR0dYYpPxJitctqJCAsxM9q+i5qyuyi2W0BpKUCiGhtMbeLhkiuhHMgf9kZm
LKEDC/7m+lNAL7GnST55aLWAGInFawdtciSpffCFE07hkEUgdN4dgr0bAIroWVdyn60gp46Fov68
sxd8QqspbatAjSIhJ/n96wpjkmoRTAnlbf4xauINiy6IUILC4BQdmi0IkuNSWhHsEYkgyN2z0w7L
uxg0sUhq41YlhrntOdRI1peS1z3bV/e5StS8+tlLwbrtymeXqtaDpPEedAqBrmE6GOY5NnqfsgAj
LQ6y0kBS7wFsMgUV5QB8dciLfgJwFqu0uUs7mjyhlDeTpz53s6+9ap9BiOgnBZ4blTq41jj0jxkp
qtvhkOT2p0qLXVt588qEHC+iShGCK55RNBk3cv6Hd6qAKrkmvx/rmfdcfD7JQOvy5DKVSc1z2WDq
83qDYXnH/zPUjFMlbDqFEL1XvsHLqqB+2mP8UTDRLnPWnjdNV6ZbOqPQcFqv0q6me/gKMXcMZA60
X3YqT8OxZJid6k/TPoOFR/5qTAuOnYpF2web05jsBZhHqX7hUJ5TOyTCtxUBu70UkDBQXew3RcMQ
XcwF0PcC9k+bJlRxfIFqSw+Wv3JeOiX7e3TZMy2Vu4HpTBUOjk54Y3Jrze9X9KcQAutSsq47ebTB
fsUIe259pS0I9QsdSGaeSdxMsdBJ6/jp70ncGkm9DzMe9gdk2RrmjIaUAFwHk6CBP6agTTTKHCZs
fFFM/iSbRykfhVYg2jvw8NVBJlyVf6pI0Eaq8D0ObE8VeGarEIK7PvJUmnInKxoqHTm3oZuMRN6R
uhvhpH5IoS6XfVNX9ruZRFVp9mKv60bdZynaRJUaZnPmUdrMVaKPbiUZVlHytG6wnqouqXowJe6U
L89XgNxEBOJeF/YXYAWg+3rNbPjcK1OTnemZarTwK0ZkJFKAzZJvWFwK4I/CJXUXmLGljEu0QAXu
htcrLKHs43iCyjdLWaqviDzoXa3Rs7QQ+UEQST/eTOHwB6jskmktek0552kY5uSbAKo7bC0CgRoQ
aVcEFwmJUvYbx5YGAxkY5cHOfNDX8sA0tXiVfC9MK9bKxPrK2X7BL/GCjLjBPnG6L47LL298CF7H
f4aoJs+HcMXc9OVNq+jRlGGCyM6s7LI8ZDIwKNc/2xpfXHHoYElnA8m9oOd0799JYah0K6i4ObxL
sYvYfKLR3NwBLZlVUhXVPyzs8QquMzQjrOZOddmX7rxGMZ3l5FOZI73r0WBnsSGlZhNPM+ttTOBt
bFVH8+dDy3mB/oIh2QOrI0GqQRXyXFGn5arhsGQ8UkRIybrbaMMdWGfGx4jmtUJvwzs4Oxq4pWS6
4gsbuKCLgt7FZs4Jki1ASWOnvoHikO5OnKexFXXrQB+bT/6lfP/hCSYqE27Xq2PlxOKXAiFpi8DE
ilDjQBOzGmMQEtwWCxcxzYwgd+IkJm17COkBzawDNTLH3pKb/mpnVPMZLAj/LhxgoAuoT5YnIyOf
57jC5ihSoSeVgugPackaLVoQX7iMnYhV23ZfD41mQBqhhnoQvUki1SVIGKdqh1wZUSRWimqYWt+1
Vo7dCHbmfQRLedmLD0k1Ta1wxgdfkCWA7FkJTgh5/m2746NgI/PVHxn5UvlggaPsb0iPKh4Oj8s0
Xvl8fkC3xLa8qrPtkWoq3f2DnUK6sU9Tclhb/8l2HV0vsBYOssjwHd/ix/mhAdpzPmdvGJJJX20z
dm3sv/u5SxhyDGHjmbVi3oMsPO6zPzK2C4pu+6fScjOpvSaJqhIu5U06AgcoueoT8mVlFfn0JwDT
TnaFCBkhq0csAQ9fW4jH1yvclMPg+lPQJdz3dZVIp28+dV5iKer98Xu2QlszPR97TcF84yG3WpCr
RQcHhsid+pU9/DDL/N3WbUyrtEoBp5ZC/ez6zp8yMwsiLpbmsXruwCQsKlYVPg7FePq+xub8yn40
rSkkEcQgtqt5ajyDGDymG00trL6YAAAF3DWcpgZZsLM8Yp4MZIG17n8ojXUmlRn7swMB89r/ZMpa
jPVnlNAidEjsV+AKY2mnA7y9QemTB0FRsQO1AynkwywDjjIm0hBJmXrGtLdE9/W2xKSGzUvtrRDX
VXwsAryrVfASizZCRQzyxYw82tN5lGphnRC1h/0/4D9LNf3gV9P2jaP5r3xOes1khOtFwcvN0Ppi
y5dL9vyao6QwwNpNBz6j86YQPL6g31rfKt7uiGwcjgdNyUwhBe2zXlaMid5yoDHc/HwzN8qZE7UK
zXnd7KMGSOfGjGMf9fSBJAUayRhjhm3473PdCcagtCfaWq8ityBEpiR4abBiniKoUni94hJW+F9y
xDIh7vUbiJ0sJhVAbqtAK01bB7LsMuEvVVtj9cSnJO5IHkmhff7uSy3zv2FZqe+snl4IFKWyMpyu
PRAd5PJ+mh+SpOlA8MFsIKX81po/Wyx921bOvbKlnOy2GwVuWKS3W38IER2yFghpiR9oprICSw+x
EIZtSMWg/l/AA8GmACAxJ66UBnsbyvKKegaOpOdyg63fbBn2Fk6cBzC4nT2ejJuPHXUcUyQ8khQs
D3949bEm53nPO4uReLPfb0OOIuPk3SKBG/ZwP1GvHqTj5GQ+Xg42iqyYRAo6IiBMEF+Ku59KKMcn
m17pcbspeB3m/A5fc8IXGdLkfhVw+BhS7Nx/hW6fhHTqaR+ro31JhVrcFxZovUBeFZvk+n6nVQw0
082erg0RbTG1/am01gu1p2b+bvmX+7K81FWGj7hfh7mQq0ru0SdHCIDTzZXwV+a+SWfi0nmULt0P
iHLYkPdlENJS2RFBsYoq2oT0zZG1cxZWOjFKJJRwxFH+Kr+AUU02UDAtdiG4d7isYzQue8s+XYMg
UWltqem9kNqnnCeSZWvVt9ZZ3fg+QuJzLZ1redsrhlZq2UkfpFo5Jh8y7LF14K6LhvPbgB4zfnyG
B+SUlYG7+njZC1NMX4kVrEVRKq+RZTM5hpJAiygSYZP5pTpOsls1mgbdTwvaDjAsdEsWrEKHQCjo
2sabLB9VX1+3Sl3AroQ8RP9zRwvKhiU2dYeZ5sWAv5a2cnJT1DEiOYWQFFT/h6el1NS5cf+I6YOI
7C/OfHYIKF3CgzsPQb7ReGAZPvOJUSrApQf9o/UTiRQ7NTUKwE5EKCx8VN6RVVyJRsdxWrttTE22
atV7n93YJ9vRKUz4MA8QbaFCiQKcHoEX5xPrHH9DjQv9n1LZ0u16TKR1UmrU0pNw0tUEffCryZoA
eYaFwxyiXJNoCau47pAgLLb9Y5mLCvP5EWVqtWPnvYCKQc+g+lp/VPV6+c/g7EskL1qzfeTJ6Nni
hECygUm6x17x0OLuG+tA+pBijQYZiixXhedCscfVSCe2d7slLP3yClUCzbqD6QA5H1q/8OR9ptd6
nU+L68jtLBYHkRFa1GPUxJNogXAWO/z8FD0LApC+k3nX1FSylOZP8AGQIpyMaDtVJt4m6ne6LIOm
HlpPIQvWDRfn+aEAe97nxEl5vLmerrN4v60iqwlvp7xij8FMbtBgJ4A+y/jbHSJsdW20iPYcnAbq
LqFzuwIj8R05yanw8VfqtPxh7jDRlMZ0P/So0Hu62PEPOziy9gO8UQDOTKg+uazI1jbMrwhm0R5P
Itb/XgJ3hPTI5KsJnvrohLgj1sPQITEYoHXFg/4kVcN5nQo9doOyOIGHvQsvpEbcg78EJ1KoyDtp
ykyGbkrXAFBSHtglwJamY4LdccekCwTFF6GZoBuXkt979uxzaWLw25nRzjX7CqdUMTuiNo1ldL6v
Gq4SQ5I5oW8q4TqYH+NNpOpEwlRdF5jB+/BnWdHCjThfNIRTy9Izy3167HIT06pyhoQAEm8rTy+x
OAsNol3U4X8d40cC0aS0qs2ejqH/goy1O/YUCcamK/JlicAsNnyzKHisOjEqrGFErx0RbxAUJm26
NNo8+c7j3gJQZldAm8hxnydmM3XwYM5n8xP5JMzXNpm6fx9XWW931ezisnff7Kc1Z9oPj6/NbIrk
QeJdI/Vpu+prdfP97qdVfdVaB/hefwk1thLZxQrsk8DfSnwtvCbmrfZVN8eOhCJLvX38eJzpz8ab
BTdjdh1RnzWiyvHW5/237RqWfCxxf/kldIoJieu90deKS0NH4KKM+0Oh3nWgXHtTv+5DUM4B0KZV
n60D6y7pGIkl5fWbDMnMenX0o81Rn1/HSLHDmh+HHG22Tyl2MVk02EwYUAYtNnPkWk7eGGnNIcrO
fGYc9Spgv1Dhyo7NcVbFH+6inPiYnzwXjf2+qaxzNjEchWblgCq4kvI+5hFSb75uYJ8r17x0M1CD
44sVSsiQWLx8U+/JS5zjeQ0fISUdC8URJr5lA/+BrKSG24vpqRvrcLFbyUoxiyTkSLZ9DfiXH/qg
JBoyA7sEyN44Px8oGCpdYst3aR78wewKH48wZ4LIe3q17ahR6/DhKMLY5afd9ddCGneH5PL/LaOO
SEjAWaOT7NrnjqPSvOdm/mPOiDzw5ZRiA2dYvLeW6gWwuPaAnk8IpSQ5peEvb9aPFurtw/mXUw5f
AwtjTEjFUd0PjLJt2Rdc5Z11ynOPtoTie+QHfAcU1IAxPD6lFXMXsOs1hGY6rIUZIAz8EnuFJMdA
R1mi/2YUCnDA8UZvvVBBbGMM9Lzh6fBPugEXPOnUEPoqsP8vGr5WgcZ1e0by5DRwJrKlTEaIP1T/
JJ/g4lAm9RcNs5ng/amWx5nmpdMGuA0DPNCygRc5o2EGU12ej6/QF3YBShncvN4yrO8Re1YpGbeI
bsRhOVoyZrG+esonZdbY1weN83iG33ApI4LeKDLtv/lu4Pbkurld2icMhVdUjKEQvIbqoPkmgf7w
eARy+F/fxYLke41rLW+uT6/u0PaT9t41dfFoFfE5U10uei6msUmXq4vkl9XnDLj+sVXmQhIp2WnS
fndFFexNiTohHDWuo0KA/SWjF14d/GCXOetVUOwTwTw7+kEU4vtUdRR3YpiMaSlraQTNelvl2/7t
YpM2G8vjlLqcbYoa0BZqEFHz3TQRVIx+bih1F1Xcyxr+gxcv1IVjBT3PvqqxBn2obFGSZkODdadU
QmHWwRgwhrOO2n9wdBL3W+lr6igtiD4WbQKuA9sCaQ+izWX+nHubvJSYr1YPuZ1wCicnFIQNYl5j
T+f8Z2BV5AXFH3uL2iGyJcjgkHCTnEzujGxDLinsgN5NS0G+ZcX7SyFpJNoyOH+3zME/qEKEwzkO
1WcCKjwgCAG0eZixJF2YZrtf4OiyNuerQF95dMPuz8dhOyaaBDD/lczHw1XBgFrV1UVO3X2sfldT
fnry3ZoNucRcj+pbd5uSuhcQaZ99J1Ow7NQzzQPVaRPTIux95mH8Mr/6SQ7NNJ2bfKB5EOhpUyE6
B2GOMnxUT2EbLwdSpr9U5BLYGvfdDWo3u6/jUxdXnFqmUiqzlxQVnFAG9pnn5yx7zQocs2ARLFJN
+lYsj0c3KdorGNyJbgN870cwhqcNWq/rkLjIK+zK5aaO3MRuzztgXEmBF3FG9uITdhoF4dB2VRfG
nocjTxQJSwrKB7j4nPuKuacmzK5eWjjJxPTY1XEVT2PAqJzDMxpyW2XxC80lA0Q5ezk3TN0DuHNw
U/w5yBsnNDAqYSd7JKJS9glZZfDbHMcpqMxDImNgrsH4VvB01/YinDXjSsHI3dRtEMI1mBa2ApzQ
OtTRD/ZcAIBqUVxH86dL4CCMy3bDKxGDqfEGQIkAcOBcizeUlfVecj4jrP9J8OF5dDsLR8gCMwlZ
klUUGXJDlPRUPPjVT6SQKuGgReoGJarl6uY7Yc91vmZW+9AlXurJoiEIWdxQkX/+wVHpd5Fro0bM
115jOKbud0x7c7yyMh0KRJBTJ6kz/+f33ex+xgd9vJNDTiJQK+qnveWukb42mBoYn6tywbie4Bgz
TZhlYG7VFS3zWirFI1ypw7WhShT1Yq0BEPnL6fUfZ5GA2BhnMZ4pmkRXd6etpxIi4m/WkUU3n6qm
rpYyf6DV1MPsLjDGwvFxHwA54Vgdos0rtCXVTSJ8708Ax49V+DNkvMyQpE1Vferd9di8ZhJI0TYB
9kl6j4r73dXpdk1zGI09K8N0JAPESYB5p49XyPi7Pb9hGCZ5eZo1vAl5TnolxCAb+TJMJPRKoYNl
Eu/6OY12s74SUrP+ON8Jqs1mqzOkXWp6H5FYgswm/iC8ybnHdYIOXpEVaWzPe74xUxLNFYppJFOg
cx+D7Kqisga94uL2+HWnTTP/CrO4EzEVFbZQsUX6BzrQLaVAPglobqlwB+yiBr7Cg2g16iGi4yzc
UF2QdjuSYiVLQRLtPh/E/Onjkfbb3PNCwsVNFosrbLySZtpgNsNRzmL9/1X1FtXqADgBGM4f1e6C
ZYgwsAdM2ifWkVWs9xLF3eqjz/TW5cZWS+19TCuIgcnW5aoarC7EWxVQLcKimeoG4GzA/7Fd+cm/
btjgkK6zbI1wlV4Memrj7OhAIEdGtGcKvZrFkDnnft69wFXpWDmru3wBkFfD7pqXBv2LdZ5+2/ND
8LQ4RyMkG66bndeDaIrqgJ8SxqytYuymLBw9y8m50s4b1jFvQzD6u1ukySH8977q6JYivlZTn9i9
BZU7WwEiLkBNy/5rbH5dTdhsB10J9vu20rif6Y4PLojDpzaM8uLGZqCBH28OWOn+g6ez+feK+cGV
35rJI0+ovKReoCNtPdjbM5UoaphVrQ8H0xPHz+nAKQxOdPrrNH1ug0hJStuD3nYojrKd8aV0pjQW
h1BBQsCeRK/T8oGVQDywplncnoTmRet52mcIv7mcVA1wDHmcStzVdSyoTQIQ/rwhJXfXRPUk6NVx
352kUcFVST6wbhxeaucqWizjdzWI09ff3EmN/KP1eCD80E7WJTwUKcwy9nyShYr8MvLp4/xk5Lc/
B2tdqmtzcusErGxo0fKizxiZyv3P8tIMlysQe35Y2w2zDgo1iX/eadJm5FjaceL4i7RHZyJ5N1J2
Psiw2WSJW8l+kiv78KcPCLrS21n9mXJcpPKcTrq0iK8GITxL3lLxKawAyHpzvOSEWuSphrC0K2xv
AGYyM18mFe0ocROePFTNbE1oDKlVp1ODd5aOs5N2/JUDwZzzO6YAvp0ry3ivEoChkeInPgyFD702
eb2xsRNCraSx2CmIU/aNAX48J4oEnBup3sHfnSpasM9kDPjQ7xfy5jVvay7mMTodwkJ2A4UaKDcT
OxkLmEaGFtMVhW1CW9iPLcTO6mtUKN73zy0LZn0o6OcpNCTlsnb2VmBl7I95DfUwmGqACVU3IP+J
EybAddtc0WCVq1p8RER0+RepH4hF1uD51sc8B4NPHpllAjr6xOrdpzllO1k/qqZzI0iY4zlH7YIY
l77OQbmZwXt7yrx2/72zXHdqRwSTCKYjfLSrphu9Ul9fs51FWgummOJIRo6slSDJKXJXB3CgZ3mF
4IG3l4RjF+Xl05J3EdugFCQH8phvQ8nw1HGLv+TcLygNd2V25BUUIgoVuQAzqMCxKwY0RT7IIBoE
Ck4NwynFXz/qWj0xEgVFxecJX3Qma25DAD6ddxu63BHtyWQ6zGsr9Icx7XtPWS8YHE+xXYKTNM6l
3lu/RGTM4KGj48Ca0sz6l6Yo/6DgbREzBQ73wNC7tFMFUWvniPxbyLV3TRSPSu+jYNI5QuW9tOZW
9+XxNVr0t+qVC3yqIfabsSP7R8qL2Vcyzu/M428k1s6Pm7u2bzVlTSBZvpyUTk9hpSuq4nFKI0EH
bo95syaUyaQd0PYC5bmWzFlHCiJrAIVzwLTkbIrLoZV5v/vtwKjrdc73fbMqIvW52vjpl1FWbrKA
akpvmu0/xky8DCCMTJDrtIXqeF7np+Vl/PLwC78pRkeOhzlyY3NzSZYR7df04sJaqhkcn1btbCnw
IN1dpluHkQs5dAzfoa2ZnN8phxx99jKBH8Bpf1kSnuqAIFZFYy4npd+k+qTCUwjDA+fKrT7QA/VR
PVW5Q28drBvdIkHTPhNoWtbhQynoNgCTyDsR3DtHI2TbIDcak1hYBie4BlFiZdsWfHS+nt6ysL1u
WUrngx1EJ0oqntq2psWDGWGgO/7MPVIb17bbtnI97bheZUXiQ2EaCslyqeDJ76GrH8qg08pwM0Lu
tVGlUiC/pmDE+7HsyCjSV9MKsSAtH8vHctfGLVXGOdeKPSRcQ5ya6NYJvDWGxUdby2s2xCBqE71P
EJdnp41EGWEdgudtph+qjgjYAvx0MoQ15BtyB10hth9snsOADfidZb/SUv1i4ic5/HsFSuCtw+N5
DRe6USaDQeXSsQAlogSwIwsIMo2gsV+kQTAQEgS/3I/aT+HT4IlneSmV19CLvHM2HbWloouhwxAy
3JpSM/wzKQtL4P4pBCwAEKZBQk0SV/Y23jD/p44iONdy5Ixke37dVotNwuf6drQy1XHjYdSwKeyP
eoehPwEGATYQwwABYQHiVINnNacZzd/F+5/T8TRLnm7zvwQcfBQluZJqShvJX7Z6e7zLK/s6YOep
B6U+GLIg4b7n6jaqfBZ9r1OYTDc5W4oIVofbXWpbZcDOk+sh60QzZasnDdUy9E8lhEx3LSsEj1jE
yq2jRX09U98aRjeIH5QhqKa7f7gqswUOfhSDmtkOo4kxt/s8WaIE5cJ25HGFG/5oaNayFUZ/TYR6
+G0LBhnssi3TLmGpHzxwrFU2GR05RaDdJDjBpohEBpWLZixHb2u6PEb1MLTS0ks98Yh4KYxP4QOq
rlDkFncGzr9l7ZZ+uXgudN7eVgk9SoR3n5hFcROKfwYA9OFVaRghbnjUfAZwQLAwBsZ1IA/+M6/p
AWbXFhETxWhn23MpvK/Uyt3HjWNzO+pe98sfWrETRfCKAt/u4kE7xKREA6oZJFoewMnRoVmccQ49
932INjWIvpJ01uah7pp/tj9gAkLDavZyJY+MmRrpkKIgPvCi1FNZqasCf68U67nc29i1yQ/NhtSA
SIIUTfCznGU2N8dzjNB4j4QHpkI/uH7iCzfijJ8sq6vYyGS20SOp6tU0GB8A+3tpzf3zQ6iwzgv+
TedFEYn7OMuqRr1umDCLoHhZLbIis2KMga36ls+ByACwI/k+7cJzL8eJtaRvELzmisR/EOpzpyDH
btldhviygxbHLhQp8UfUCe7xByOGjWoEQK6ndLfKhwZL9KnenLMN10R5gS5KH06Evq7oJgcwhxHf
Mhd7h/QL8ZYJLMrUNy0MmnURHytCCByHAnp4ZDOjTSJJP43TzTK49Xjj9EKXnZXSPWFXmeukKkx0
TaXWK4Fdt5wLkbZ0EXavddaHMl+PaYUw71D5q+6GxOYLmE3KBoPeyBWGbiSoDVmpMWPJeXHj1Kym
gauJfIWHFX8T781cFB8FU3NQJM8Pw3v1eUOloTFegv/isvpCIGgrlWCBV/1Udz87fAXoDNEgXXPR
I/XAX2qXrmXLNIAg0GQrOG1bMaNt3Den2Xy79K8D4RNOT+nGQhc6TK9QMV8ILUMSwvLy/N5J5N86
fmO/mC7sxD5MT6qZ9MkIEwqC14VBPlTwZUCzQu2mhmYQqXIsMH31jzW9iNrPkOLpyyaZu4hyuXBr
uCdI8vDtTtvrVYDoQTOmYaEo3Kf0I2XJ4FzjkmSJncayxQgeCuXauTif/3t47N/N0usw1Gl0kj/5
KK126YbKeJDl6IdWNZMPDJpzdX63GmSDiUyc63VqSZVR9Lv853r4aKCUi9LbEnFRX93dUSFTfTwn
x9ebjj6o+JrvtlJy5HtFbA3OCAZAiOQBEzNx4xYX6sKncjuL6gAyoQDqDX/8D8+EU8UD+qv5x6gQ
M2nD3Vy7sLws6L8K2CaHDMs9KTg3y9YKQ7EOvHbuv6pDR705PEpbXpbPwBvneS3qgQ/T3qjKXJgP
xZjm3lOBuw9eY2V8TMYoxGaol340CAQHkVHfT7iNItWg5CDI1wzSCvTAQ/kbcxm8yqlxf3oRa9HV
8FSsEQXxeIKVgWqJPRBUX9BNkZfY3v31MbIpPbZNJjv6vODnyEYlWy20VhOlxaZWxpCNzUBwSZX8
1cKYOmYtSb7RUwHWtYPn77UPp4RSXTJCvZBPyg7BysY6MUk48MyHboGjmgdRLn2z2G7n7fVZMMO1
CwUwHGroG7Bf4qasPE1k+tnVI1c6y9rEeXiIqW21KLTupPXCCOEqFdKqYzptfqvoTOuaS95QNT0U
ZRtABrheOyYpSFlbpGsjWoxNkuruQbcMvyo4+aFQdd0bkhZSSigFMfQxpOg5dggRLXyNZYOtbSvZ
X7NtA0KNj+Yy/3xQZVhg76zVLr777sj3CqUNKOAa9Uzke3CdxdjgTkV2CLuSyBVPNUHyLGBZEDJA
ie3QhHdIhwqqTvVAo/8fO/EGF408xXUHat+oLBUT72u3QSNeszy9Djp8tbiJy1XT33Sg7P4FqP+M
RSJ5fYQDOmnG06mP+rC7vzosEO1wnu9HEi5/UHpiJC6FRNPabSUlR21M4af4H956SjXxP2syf3hq
xQ7MnC1K9Nn83NvHx9bMfd3jHVpXeD2x5YS4jYESRX5i83EbDc91mOm7ONdM7vw4bSn6gOwZarE3
W7B8cONTVzkiIi1uxjicHYrUcySwnMmEUzUb6HbRtTHBtRYJ7d39QZzJDrQKT6cOqVLeeijwRvT7
Sf3zheuU9qxtGt8n5X17TT7GMZRhjojmReP8r+gaFMPqxFMp0s582Oa7kgMlh9yMOCl2dm3W2kYK
a+N3z/G+cj0Be+xIxv0YIQFHeyXTjG7BTQA7j0k5yVb3TPnkFh4p9UkvhuDI3qT/Y3nHVw2QLVNJ
Gt46efrzVOxf8VN2xx8W0Bw2MP3ZyxKQ+dq2fUnMUmCsFJHyUwn/oSoEHLAFco6p7pyvriOfjGnW
d1oUhMQUOI6EU/85bTz/+liV7683igK8u1wekpeWQMu6ctnZ1M4M8tcJ01m6tGwOsgPardRyLeVO
07YD+37JN1pBwBoef1l+G4+igVuKBTlPEJiuSZsxbg2dYJkE2+Mnfzo4MpaJlsvQ5RLu9Vchq3n4
Q/BzZ3QaGz1fWVPo75vQ7rletyPs1nyRf0/kOHoZn3L7xKWqmwEWEux97aNWPFfT90yDp9ivfAFF
efCQ+ymQCfZY3MDIu2pJW8oYSOyRXgaWWcP3lX+We9C0qdWoUYobl8wCc2lfmp4zwstlmTNp7ftg
Pkj2SPQPc03mi1Sic12M6LGCAZLief1UfCrfhKb30CWi2ECrOxVj8DaODXPoUx6n0Ru91feb4XAo
Zf0NDjk2iPuyMSsiQdqzabDClHSgE0ZeQR00iYUDJI7nIax75oG7iXHCpAo97HpD7Dqw5GiK80ZV
hIhjUAPRiriaiOZA05f6iT5dppxypk1SoKB+Mdlcl24HJtQpB6+tBhlkr6ObpN9cpSCSLPmGprGm
apfWLDfAPeZhaklhpiWzz+KSQqKDt1RDnAs+qOG5IwGSygS2dGod5dcvwckEfWFemLoVbH3dwW4F
wJiroaAWfrUm5US0QfMDqK/E/8q7MNRBFcrgGSb/0EQmL2uEazfANilj+POEh2JhVwpmbk0m2c5u
XKbHxMk0MTqfRCbL5DOCiC6VTKEH/ocNlY7Hl0DgkQ7ABjngMOvpBn6znPrkgsuVAwpYlUbhDWO1
SsrVYi/ccCwGX56HP0LyqC38m/jiYBzM81xgrI1QA3eyQ9nebvukwLFWOUdPc4Ek1OIKqFOrn3wK
7iuLHZYk/3xalj0a38bL6nC0/475Hmqon29OTyCN/K/cITOefH5Vq21C7w+sKqLs6JTtwOJ09w6v
1hFEstAI44FRujiCF/mjOzZ7wz0CeSNF7hlvzkRK9bkRe9NAkTZc5J4iE35qVn/RZcnpODWCT/2F
+tVb6Z5jBvVCDxY3B3IUASKBx0ZH7GEG3xqRAMlpicgs0a78QAB0PI5ELPZsLlkN+bNF67MfWveu
VttV72bcba5a+0CvOggw6K4zaC24cafbwvchYlvsueoRmFQAwSg6np0mibjBlsQl6j+kbsBBOWUQ
bYiGXzb95Fv+Ke4/j12Bxb5qKjtRIauSa4/Qobd63YV7r+DqaDW6cgeZSzUVhE5JUh/8OAFHf3ek
tgdHewSv5HI7+/JD8H06onCX5LtKgoO8EJb3FCdOUe0E6nuNcqksAzSomKMmMo/f01LSOqLBmDO0
7yaEdvaJr+nVT/ljaQP9kjJFAwfKTBeZ3AqpODrjfy7JIBYw4KgBgpI8vp3heUEjlxz4ZBrv/nhh
obJM5fETyur3O2EwoqK1qRwcp1Sg046xkdH3vKF94Nmkvympup+7+xPeMD5Mdjp5v980JkfuC26Z
GMvyReoO7YgcnkP8EoSHLlf9cnoqqhm8aPgUjMktG3XG1ZoKid7r7KkDXZ+9feNGuLPfGaPh32uI
BWNA+G7xddJNM+h2DQYBXB4/r9nSkd9c/7ZYzsmMno77dFE5YAUP8UIGIIZtl4XI5OdZ3vcg6iq4
JfWBWd6pxap211p1F1SeV2XhBueNJbg45h7dUqu22AZ1oFpcDG2fD4s+A/zrw+8+Tvzl9smVnEpN
qrgYTfypNo/6r9KoByzBfilFHt4TC5BfSQN20ZF9FckIDWAw35vcSDgry2jEVnfMQQgOSqPpsi2h
MreStVtVFbqHCpmMVYIBMh5tw0ftA7R/veWhRsERtt1ISpVGPPOf1cRmsGj4rvx8xHO08KnZpQAa
vEn0pqd2f66KYCvFqFC3zxXIlnalzOmj7OVzXF9oh7Xmsc9R124t/6Wua/7lwvd7jwfpdyrtDkSd
HnraonNdNqdcOFjfFNzT2qNgX/OCKJFIxggVn8USNA1G68rruuv9dE5T4tzI6ht98iL3pQxFFBvI
zNxQcNXiYtInqyGWB6oRcUzepQIAkFr0czEPvk/mx2u8sSz/KWPgro5vhKIYNczO/PxhA1C0A6ql
KHoH8I+8awtuoMy9FouCXNHRJKXRpySU1kOwsKfZNUHtIS+fUzlwRbtAF2/EZAYLNqtbklGVWZmV
2tUbqddODJA+MOMJ7Bbh0AobxmVhPjyBqw+a1GUxaeAgROuCg98enaWFHDoU8M9uQ+5zFXvxd3Ls
O5+hRE/mxDMUXleDWO7TtZfR2+VKmoy50BVvS3LeTyVokH3Lv0Vk6CRBtoKcIMk5NAGzYrxPXn5N
I3bbt/QebQlSUGAe0zbbWTjEhSgwAHZ9PdbfKfo6Vfx3aTFcepD/zFWT3pfUqJo/LrQV4Yz+NrT9
ua+/Efnhv/v2eR+vfkYHx0C2HqutcE0ArudP0wYIeeLizSRPj7KP2kG6+wB6/nP/CskU7NckwEol
OGjoPJZ3PzqrSPqmQsTle6DMqZu81ZZ6qVMeS9S6ZWmsbO+fVCWzwyMTgNS2yhWOBpGW4MC7NjDY
lN2Io8FR/EbOnOEoAJGLUjDU2Zk8sZYTWJCPmJ3pPnkLv1OWGwWR1pA/7mgiFTn/p2YT9AQ9xxhD
msHcDQ02DZz8zlnebkpcy6MA44RbjZQpArM6DdTOE62tYIgOmyNnXYUm7lnGshWDNGCjVj0j+kQE
Ppv9wmFJcj7xtng/krm/JEmmIR28KANaZPwPfm/EbpJjNueg69WTT2s6wNbzdu6druFqtnahGt2e
2MABBuVxb45a8Bb6FX2HNV1gwFWD1OEfB42tjBYg2HpIafCgtB+22MYupY0kxunOX+oFttFynr+u
TxrcEIWQ+dWxGgBPB/t++YBa0wM5kGfZkSjPYRL9znrzsiL0iiqbKJFNCAQtMizMJa+3VwjP0i7D
VWR1XqthLBsfrZVdfCPvMM3GbKiAlwd5av9XLQ1HjuZVmNDhFSDnbnaB3lrDYSimrp79v8b7TzrS
yFSa4dVruBta7SQu+5r6M7z6Oxk8e8GOqnOCg2HBqIM71dqPzDrIO0jbzWz9Z94y9yMjjcXEf9PH
rFcAWt+MVt6qG1G7QtkQxiFY+q/XItF4p2yr2fx2/JDDeqLvwuRyB3g2U+lLV3YCVkILivQU9/YK
49yXF2wR+6ojSa8vitBBDq3v+hECXaK+inuXSekVi5JXIeSPZpKAMYG6LmX3yuKYn+tnRI8Pw+JX
75G6lsbLm5vOklsOB4DnU1OsuCLHBx1tvnttBw4FhqyNdOzHtLR6xbzq8GnbSUenVKJGryH3n7/N
cUSKSMRVTZqfEzHE/29kLZae6DjIdZaQ7kaPif8l7gWgLP2rv/coteFcZbhmAqGqys41HrGDVrWO
OEhr5Dkqzf/m8ObFZeIIA/n5SKPeX8eejsvZTTk5l0NqQfGuMA8sGswmjxszyULrSOFDPjSrdu81
btKF1Kq/QniERXzXQWkm0cqoRFWvh3eqtLNeNG1C6ZrtnQkHJ+UmhqeojV+gGN+J0hLJJV+WAEX8
GL64fw8AuRMOzjrmIp0mc9xIvSslt4KjsjdSyqDGx5VfLrjdmm09s3XnAF1UqHNbShtOozlUOW3W
uPx3WvsLd1RQmkYm7d9pyWRHLaI1LUYKBDHi9rqEaLTCW387kZjpkDGs9iMQhy9n3GDsEUqGnIje
3Ka/b6ox27G82wfdGmSSVJsbkRre4QDnm97+SqjdqkMBicd5ymIPNcx64nb23eK0e95WW+81FIOy
7hbzhbhFCEsF9wCEwmbJqW2eijo56tt/rLUAngo3xTj7Vx1KJr9Cas3nGmusYP7EcW2dqHXm5U0L
pZqQFlDkpD0mekaUj0X9GA4QqwzAp10P+zKZ6PYle5gV6CCNhEJAFuz8R0/XRnLs31xr+Qy27Dbv
h9zYMFh1s16Q3PVhiARCBkoMM1yb0Iqyri7p5EisjwQxJ9wnhk/i329K2FJbFE7DsUZTbEqNklCd
awUMKMEJtdx/4XJwJVbSjEy3pz6o8eLpt26kwpZVX4tI20sN/nF8KU5VyY91pkWVim9qVC9SYvH6
9jMIFPLvq9ZoRFOycG7KKvA72DEYaWSsmokRJoOzlpwsSn6B5BA7VDMQkag8k01rGRRUK1DHkYeh
XZtz03yYyR3pqlNUsN7y+Lq7mwgKZ0aGraJKoDA/utOYNnt+WsU+kwMvsQpAK29cB/OOqw5Grd5C
kRSl4arDfzZi5FPJBFdW3jqVYRX+e3KiZ+AcxyAQYKl8N7T7QYqZSxD4YClZfuKY862JmzTIVbUt
/L2o8bNeAAx/g2PKSFFnbZxrwMXwwU+6A6ese0YiKh+7Ei5AMWRMId5F+4brzoXGRYEJEnbOGyZs
yi9sYIibtDPaK+C5z8GisUmHrvP5P2Jb2y1k2W9a/G26+Qb8gU7SoHNpT4ajiqgW51i4xg4lbwJN
fBszS5BbE0+Y9UIQzhm1WyL9TK9ZsV/uy/i0+/3bRjUBY8wuB+QRsstdeRYNxDCCEHlvfW4CaQWP
PweNSQGZnOkclq6aH46TrtfpenOszosndfXp7Ui5rU7tzLNJtWvl9w07lVlTLxD39dR7l//wvKlY
JXgappsy1j1Eh6pmi+nZNK7vzKZPrqZPnRgeV83TcbwEn8O5XicvN1fLrm3QtBZNak8qTlsvwOa2
adSAjCNm+jOI0vTI89UisX04VxtMddvinlpWePA61iz4bV/Ju6Er1rt9HEeLLaisPlDl6i1EVcTC
ytwM0zBTR8kBL5ibtCttDOSZGF0kHcPF7aK1+Y3d/i0SykhorOKbZ+ij2jdlxXO/GN63fMXmns9l
eFy/6GBVK8bMWm65EbXeekQuUwtyHGW+neJ7qa6PdWlcdnvpbzOTdiSnD7tu/zOSGY9Y8FReeAjz
3M+CUq0kTUioYhSD45nPCKwvfro8O9iYg6yG9sUghogQgt0oe46gHJKxNVy0ZUZDkNbmgDYQjtIR
yUbE107pX2bWC6s0chpTiQVP+/iUA18hJNKadEoxNHhQHcVJDjDF2G2mNsVLnhDkwAtMSCsSwlx7
FjQ9nZCco5M756sMP9JJ5ItMm8oaNSyghr60VPwehmHcTNNgrXBxmcjbVwlu0VvFIUpH1mOp+S4w
h6cmVVn0mJsUZiK/WcNYULzb4La6juO+Oaq5s9z7DwQj+fr2BGDeVW9KEf962ECQZ1pFpVjl6SFt
zHlrxtf5qw6/FsI3KUXqIOhr2vWQrnCabCjDRUu870WRGPI9D2Q4vg2vxpNDTSSv/Amt3Vf1Ii46
oiBDNmbE3RxECcqUhEEUhvi3aHU0feHJ2C3CWUpLVJlycZfe5T8EeRc+7sMxnUDtq4Gdo+sju+Nu
p+xgA7qay5AZMk1kyk+ucE9b6cxwUEiP28Dd2iMdxyhck9GFgmCtAHSyGdbd+GEwQbPwOJSPePNp
1x2XcRaoa2qs3MI0EV1d6XONIKZnutISrHSrgSOWQToHT6oXAVCjd0IFkVXUwZJkMvrbi/2PXHX0
G+RpYRkvDOr6D7ZDW+G0yg8L4aZ9G/+f8SOOxJf6/1Mgd+LKsZUvOx6BcSDH8tloErV0GMzGBCJ7
wiF9a+2giha4WRpzIOWzCSKfifjSuVXLUNWvY/+4Gw1wuKKFcZ0/y1YFsaRNcAFZU3qumdZ3lFvd
GTc5VS7da6BngxWSZ9nWVcB2s3bDf8dpmWrwfa4fZX5iY3f3HlYT2EQXGztOQrZUFHFXMBj+kzBH
8oGF54qfuyzOQwq78UO1hvDm7jiZheMLdkcmZSSXa/Llq6O7fk9sIam3cBKPjZ/oMelkcnpHrUVo
jSnnkbnN6URN8TrczMpgjaADorgBaCZojnpRuhoB/ml263ENb4uPoZaLV/bob2ilJqYU5RC3bWBX
bImiOgiCG4qzPVMVlNVQxdFdih01BLpaVyIt1AWNv2lmTHXf37PWet0QCl8YVulib2o7al3Hbn/z
gTNk9QlwzYMkgIfue5CcIiFtkz4tMfMlk/FxnS2KavU9Vr/biygcbS5Bh5ao2I7iAh71AaD0zF8b
Bqb5vx1D41tkSr1Rrqta56mWKxv/XyDYiimnvdIvKnVp+qxXgoKyzUUFVe3+li8RczdeZeQJlhJt
hKl8jIlQscRpU4dynS7Oaq9/WCRUKEYV1m4LYJ+g2eEzuco/S2amPdJHBhF5NtgxmDywHahe7P+y
a5Gl1yStYEV0uvIICG4ts1gucZP4Ud+q4cH9D82sD9ssk0etfIQT3D8nFFgLwAv2a2+cPuGRHvVB
vcBlaOpOXtfGj2XXZZ04E719zEgOZZJu8dwFalzMdwd5/WWR8ntnEn67xFTt+6jcpWqZKo3kmbg6
Bi387NHjKr5Ayx6dLBS9YA2bH7/TYD9p68uMV3OQEg7izMjdcEDj6TKvKozqmexhxDu5bf9AA6Wr
4CDkP4G3NbNNSGIX4eEsazfv+TJdDK9+q/BeY4wgxPE/7puSya3muQJGfypBhs7TjODXEC/l3oML
puJtVJAWrcNVpbch7dwSTQwTWj/ShgfE7S6CaiVlDFYPSKhheE/tPdNCOstwnwJZ3Pi9BZIi2KHg
Q8yaxJcXXgWpB6zTWIjBNmLosY9N7YlJEbPd84JpE1BS/si043+pjIbjvQ7Cu4zoV2pC7oQpOwJ8
zDxAweh9sE/DhN6rUFPglFHr3kzeoFdKbDw+mbStbgU1043+FuPRWqaa+/Of7Gy3KvsTe36OY4kn
b0fZNtXJ00khpwZgbzf9nrbPZtb+UpFaN0rv15bvBXkX+SMtAgait/oJwxv1kIgrme+5VdlKv5Q3
FJYibZWJzBCj/tyrZYpR3a2s1bUCjt0HMHrPn/n5UK34TuM+LWSRNupktSalx+u9JMn0UKxWLT/C
4hEIsVcHmJsRlHD5baxz3KyJl8ZDc0Cnf0QZPZd/kaVNYhnsU6kzHn10k3DkVikc2gB7tFsKxHjZ
Tn8cXHCuK6SMejHckIBLVfz8L/j182x8xuTyWOf6jJTXNtGfR8ZGkUwwRB2h1jTrAuX/QLPXNncE
K3QsRQt+aKArcKX8QmzL4FMi4zF4Rpx+xWGm2XWZbcL0/0cF+GIt1A38ZIOiLg0ifLIL9VbeeehR
Yq5b/U92QhdCVx/jcRt3RDo+b7ckU68qO4QCI4Rubt5xrW7oy9l75x0boHr23x1otFl/EiTL8Nmj
7BvViDEcxlaHDHkD9JlMubzlDuV9+kk3uhcf5LXjBWfoQ+ltFOv+ja3spzbvf6yi1IKwk2ronYnx
2uXm9XM8156P3jPCfStXkE6hvLtkJ4/lDs7W/B8MZaKB2oBPacx2V9N7U5nAp5VhyL35tB/cXi3C
b+5kDix1BgstpQo6Jr6k4QhZW1cW6dgAhRG2GUK+vI4HqoYKeuRkYzz9OQtRv/xzNVu8PWiP6HbI
Zq6cYHjGV7bhdAt6pZo/yLAmLH9Vyt6dkyae66wEoHtEddul3EDgM4zoX6WyYuN0PH77uxSwdQ9l
6+uBPj/VFdYCYYHGxuNIqKHaY4D8at3Tgaca5sKyRQ8YqLmVnfrwlnpVIZ18D/K1Mo2RcdwByzRK
4IB9bXwOEOwDakC8MFWgR9pelA3RqTrKDn7mpP/FOTNnPej6Wcw1unQTvJwI7pmgDZ7IIV43cLUP
qBmaok7HI4GzJNmdmnzfLbAb5+HZKuqURlKMYkR3ZqfZHtBTUlSpom90jvttBLkp4+7ac45oCjMW
ibjDIpVbdFzoIlTfPc17+aYk1peAd9dKJhTKugTUD89nm7Olv2Jt8ep28Lelyq0KRNYzQEn4DKSZ
mNQNeaugvbYh48KCpEiyx6zQ+J9O5Y5PSesEba/KDqDtVOpHmwguYjg8tMfWEsb48cQ0RNG+ckLt
yZoOUxFFyVdNKqA3XQaUDE1OcMId5jGRFUJnCjSHlPvTqJhg1R98TCaDmcfs1FSQeIoh0SPlfGBk
tjpEtARXHo0tq5I8Bw5le9efcPn2SWCXiw40Ri/WSqeVquPYOQbh8i1C2CzrLLVjFMz4cvabRQCn
RfVnNhkkaldTbG1QfjsnfFt00Eby9bMWCXFbVkFwv0MPp88Q6BQq3fhMJGsmN7XoSDdzmEXVb75W
qm0YhKhhxl71D/tUL/4fQgLU+D4rsBJT+aOkSsx6ihoTljIFr7qe1yg4YyZbL1APMBYpasS+RK45
Nkkfm+tyN4PsilGHZedpxremC+10XHwnNAnfppUxwj4FUepnRnvmRWFE8/6xYv/2lopgwoy/gllp
GxtruHO5ZmVmywBz7ipBDBiJuwNuc+IcrboxDy8lC5TZS7VYkNlw7MMBb7o61WGe6f4fPkjQqwSg
Ion4JcjPHlm+/mO6ZiX5JUK+VgG+N72bLLQtuYK9zo2jo7zGhXKLNfWIDbMNoBw+1U5QAUOJyCm+
+7O7DJM9VR6RvvMLcVPf7uY6nFYNEIHy0HhmbmHqaj3IzZCSsd4Kv+NdGl0hTAi7WPHTK+dD6tFV
zDXANmZpTAO8OY0Jr3GurlNXxvLmihyArSOTsa+KNpLyXbqnwJWEocOLHXsYCIzAw1GnvIOREgTT
pT69slak5LcNjkR34qW0ohfODpdROb0o0dL6cih5aYImgEaXyQaXLvCCKA+Ab50FL+j93hbjoFI+
Ep/GYV0ozw6xSErPbeV970RR2sGuRinZmmfNpXM9F1wnMOuDmk0pzO47h1uWT2TvQFbNdhnjR88f
rc9Pe2Kh+2kNjnaR5QRN80Dbxnh8riaozFQdI8U4jZkw3bxHBLGrnQxEaZoiLmITjnJFIGIhk9oi
H87zKqkGKkp5d5ZvtdlENjN0HfMGDGs16tiFDMZdOQdWDYwraKvr4r3x3W5oEyZs+FrC5r/rYym1
nnBUPKdbAO6a1ztsHUIxHg5tTvjPudehGQ46rCIgAW/O6A1ZpGh7BPgpVjmnqDgsrgFlCyE4am+2
H9Z09k3Y0WTiiMNAM3DN9fet4juA5GTshk/PnZa9lwmVQsVEMFSXg8UAwu4qhdidfwsfDsWTFFaw
ArMDSR1PrPD0z2CWIXnV7s4tQC/IlFK/r3AJ2bAkn0/uXlmZSaRZnarjkvlSBeGXdMQk58LVyHDT
Korw342FUhFfXNu/2VkFqcGekPyQ8/yfNgQhn2UFzp8fW1aVk8sBAG10e73ZAj+KFg08789ocUCH
x4o4avnxoZvHH1TAHqnFHz2KCeAWjnYoDQB2MEWmzqG/53+18ax0R8kSIEYwVjybXYP/vN3NVYd6
Ch7/r9bbWrgOwbasytcHVEyXqBy2lk8XAHkJ6PIgRw0CAhf2GeuD/O2lrtwSon/fOZIJ1IfK9Y1u
j/uvaW+nJsR3eIhKya9dMvnAJvlxAHdSpDTateS8l2zWRZq4LnRCaDYGC9L6uZ41ef0HuAIPAikj
Bn4dYb5cImyHGS132CJEZyWgSNLcV6FXHFYF+kRaRwhSSw/Ghfu1zB/XQzYspcvbKSrsbCyDzkyd
ITM6CHVedwFo8Jcn7l6HwuSlg70rMRKw53xtsiOQ15C2sRmrDjq5QZ7SjwDN4LNZMU1OeZRetk3J
mzHh/zTcAhpr8G8pxPVxZE2NhoAaDPJoRsfd16wduLatZqO9d0atBIr1LcOgTKWYprrcyBF4H3rL
ovFb/V8qKmbhPacJLnuE7K8fDhiWbzVbxU+c9NsleNw/QkVGMroQi0WQCwD2sVsqDKGC/XQ+HhzH
89NJ6MobHr5hmJs6c4ZHsJcQ0KzbBq+r7bgwzbtKbW88dsLNS6ufeX+WWeom8eFy9Y3CEZOQnVHy
6hotgwaa1Wg1r9gBPSp5pr4QZPLws4tmF6E6bjqtne6T0sbP9GsyyNjOaZjtRB+i3guPW2NUSDKj
uTpi52iJcqEaGRi5NjVjnJtIuW8YbmDpPgOcSwOphDBQSCTlBmIvAmU3ZZgIrfKZ7qvR/lMNGRkY
HhPKliWNjOGYH8uBMMfajT+xofFFB9lmxSpZHwarbsHmIBseWbk7fG2YXYiSsImT9Tfr/9QAQsTo
VB8CZGa7jPVvd0aWZdHFORBc7zpt4kVA5lR94ftnFHOapQHCIntF3paqzTF3HAW7/DcqmYK5Mszx
nBCLgQI21IA4fC8RLC2EejgcZhoOdApOVKcGx56xvoXAoi9Pbo4w7AVkmSQgsAWrj9QCW6L2tWrG
cB+v/1+8roSHVz+a9R1K93QBr12nyWmUTO5Tu22eKcFwZM5o+z171NIa/RtWW+aNV3nEiSRdX2YF
bihdYPwKKCOEE+wBd0BZMgkVqVsAmUJdsDL6NEvGLBmH/j7TzHCzcdh4iVilz67wo9tcm2b550ku
ce3IhZNHBqKnnfGAAqGx0TFknn8LeOFlVkFXNG+6OjEnhXJMueWM3I7d4GdvilZ2dwENCH2eSal+
q3QNYvo1GvgsBca7SeL3BgGxOmZyBV0RCD5/5nD7Ry4pt0dlqt7HHSJoisJXaKcoUISwhAL71PAs
F2MDk50vpjHvq0W1tzjGBRDPmw5zT63VRJe2NrVGpXAUriye/xSi+Iy3AClNm30aYYmGxXzqTr3V
SlzqGzptxy7S6/Y7swbnY4U+PORnN9pKzaQC7c6CUc1ICvD2pKiIw2OU3tWxAkZxsl1+rtUOE/TA
EowWC46c30uSUZIuk7neprwuKv3xLJoMjTJyZMYN8RTBCxhVpTc3NNb9ZIWdEXXxJlcXMsxsoj8Q
0vLjmB+59SudgunULeY1EId1lG9fBQtB9O4ipG2mXWcdhXqliQPGTBSLWHwdWjBXLZ9qjx7cjASE
YJuBOQH8LVu3R8JB55Os6qypnafB2BhX+iqppZ9cMG6IKxG9srkQ6c1e1YJicK36zGoOJ3hJrHVF
diVY+Y6QXsjdcgPnCjPyiZZoiH1dSY/VmC/lzt8qTsDBssR4jSeaNIMJOG2uDJ9gQ+/jwnuhVlc+
RcU6ditJ3PJ3pB/J3CrwfEE5VZZRMijvUTEJEjwwX/cJL7xanNJB/7dkDqqMdthhHw8QABYXO3dI
LVtj8dtohnIvj0AcieJr+RvzFE3kNXfzcJ0Z5N7ZpvmYRxv9M5k997tFyk0fLI9iLHkC/+W4UWj5
9fBGfUUPpssoUTYQjozm+SOcUISyw1MKmSyZvGhoap2NxFVcVRYxqkDMsV4YlnDZvhcWrnSvSdP3
r4AgfoZ3wAGxNHpusL9a3OHs/tHImN//geyFHKQobDl2TG1vvTjTPRYMPxjUdXI0HUo6JYovbt55
e5vSqqpqTx7SoHEvhSMZNE6N+Js1By+iVv/3bhK0aWxFi7Xp0HiUfG2w1G8EWghPmCgiZqCHsY6a
RqjSatjHYZ1fsV1s4mh0IEsNs4WurEwp9VGilEKgwhZilxRze34oNszEaXr9nseE9jU5tj4aHPh4
T4GiD0RlhA73PtGoD5nWl4szm+FPgDV5ouoW3/7nKJ8/JPeoHi/P4IqnGFY4wXw4RFbxUrHTLmL1
twpdAHFTGqiQiFyLsfSeXlpYAGuws08M9+ymPQ3mjWvesa00QYXxwB0MuyM+VCALiwaQVniz+fq1
iLvA0JW48pJgVDuHXXGqEn+7vD8yJW9s9Xfb1atuCXy/EBDLJeqTJ8Fm7mJv/kb8F1vv31wBnARo
I05QALwDZKOexbGZMvwJuiyyd0rxiTGuTfsv1lM+XyWe82EZVcv5ZzFW7iFlI+9kDIPjdytV0ByQ
UDGfCIwdSRnQKBQAGyypDWMqDM0sG+/ipELNqpGadqdNIrK8EdRY1y8qbnL7dR4a9uhDWkAcSVO3
C0Du3WndeE9/5NNr962FDvTjdqfWLCe502MKqAcpZJBjx/5QjeJRipe6ONXyDi+79LO5mkJG0omW
X3/knjz51/C9y+hC14Ucfg9x3EPajF6LpdQCowYQxhCNDsVNoHqDc/VjtXb2o+W5/pdAGWaY8GgE
5WgT3ycu8yfz5Cyoi2IdTP6oTixsWRM8eMNaf/bNSzKEdOKpQXB89yF02ja60Cvxd2OBdhrAR/20
YrQhH9aTDkU9SKX8mrowGvLPhxub5mwO+aqJleWoSHPBHm3Gk3xIC9h4gRg1U1NKlgQSfXmxEfS6
TtMg30dVDY6AmSkefvH0lNrCmZaPANkbKDuoq8c86DepcEnwHjK16EQGG/440T1YbPId8TLKmzPA
UX4jcqIKG7gUxfQSx/VK/WmeWhtMIUu6TBaXk+MEen54rXEBKEyHN0g7/kUsAz/ttDEH7yGuW31j
WXBdpjNKCCe2AdQkNINtdoHsPcYepvG8xYV8w4rnFm/5xGQWLC5OLK6Wyc6v+dW9fJmXXMj9UzAe
jZz5hvNViddWwRt/HnDwgGVq4CtQN3kwa/EtKbjEasTOPrcv/xtb5OwLXC/PXGGZ/KDyeFpXE1GR
niGmN/tCXkdhK24rSMkjTiv0mMwa6BW8KGfoF5t8+er6udbtzaEPvtO2lzZ3pcyq1cdqIavbfJRK
KnJ4JW1x4Xb/UXEFsipFmVjsAWnI5/bboIDPJxvHdCClec/DAeICGDfLq6btC7i5ypiu40Bqmyby
twUxHY3aet34yU8oFOSsAKkKWqrIAN9moANBp0uALhZx8irfQPZcFRrY36tuxEzO5Bwg1xteWqIG
iGDCbtJufYpzOXaPbkScxFScidNSqmjcXWkqVpsW+56lmWEelcqThIVVueOv10rfw7tqOBTgAjJC
5igRHo2ICfvA3/PxgeuXTmtS1n6tS3Kt34yV9biArkgul0lKs0/9awT04PBdtkdLl+ki0WWifnid
PEM/bMRTQ4hjvPePFG6Rfs5+jn+tNR3PIeJhBQmytc6HhgWTUS0bCOt+h7zcRjIJm3wIIbho0s5u
6IbQsRAintsgeX47pV+pn/Qe6s+INPgEspzNW3bqK2DP84Ym8Jv5mvdQuDGaPwboLSgKf9UEFOgx
sBIyTwrTMr7c+otgK9vNskYJr083q85MlrZQ3ZiF2jdhwRxiKQmxDa88dAJfxS7EaQiBuinXkx/s
6O6rKz+AtDpMd4NPHWzt2BZVdRRRMsxOabn0+LBntAsHJ6vkRC/ZcTEM7OdT2p7EZYZHSzuuv368
qmWhp4Cb2vettN/NnBbEZ/8BZ8hmAflutkj17ANQozzxr5dt3RCuXvjw/A71uO+NJenGl19c6e4s
7/WEIVpabhArVwRg4k4xdhIDqCYuTpXS30hFbSDJ5Xrh+3HBbw/UDMvcPI9EDGGiP3xsdHbZgByi
UqBFi3FY0cKGb0UwN+YyJeNwYYwWybGO5AgEs20iWY5evXBDXEKQ+fvNq+Q+DsCxQEbgZi62YT+i
MucNl2ktixskVbY7w1jBqJE4orwek8NNWT1s1v/qNts2MwwUT8rmLS+cgGESqknjeppersLARzfi
K0nH/k76u00VfXQoxT4i3ocBtDj8JV4FzF/0IL/Q1tC7DJQ0sae55K50avqTKMuaXJNwCD/ESduv
eig4zQpgEjpXG2owHEsHXTG0HckmhOFYiSR5EO79LG10szETXundNqukE4l9qxJeB4oUS3ZQUlP0
naJ4aa6SC57ri0zW8KGhXpexDztvXgWSM6kOsN/hklsWHqe7gJTEuFQewD7mYMhPI4eUCjfEPIAv
41IihuDOgbrMeQD/2nj7gw3gSlF3kmHHS7t/PoyykBg3MyBLal3Qccbvw96U8tfm07aXbNKxS8od
Gfep+e837p+xLYSlg7addvGhPywZWIozXs6E3oPik9glLlFqYPhOapHD5xP+vfXhG2rb/U1H/x4F
tWGTgYZ5GRMNxUwo19VzPe9A4yCI65wgoFHkc/MeWQHkgVpRGSFONu8WfUlfGYf9vkVIOHic/W6+
3GCtD1Zg9pqf4vlen9glUQA5vCsuuGRtJJUwo/GwQc+VyeOfi4rzeEF4QL+JxgDNJitt0/UHm50P
5n5+Y3oLq91mVafDS5iAgacwfaAdciqo3VbnYpvhUlmfF76JSlNYHPeeg3UwPGsG8RtzV1prGkUz
kEKB4LrOTOwvpHYgUWQ+UVGIgT+Lkm6srgw3WAwwb67NG/WIxEZI4fPkg8LyIZJgmakVCClR8MkZ
kZ2IneYABav+u/DxMysZuRivbxPhmXYraisk9eTQNTXbvQkO9xJmCyD0ke4OOlaPG4l7jkqdWKxT
bRKXppq+d2rnG/28XiZaLcqPv1zBrtka46epKveNzbQMfmaJi6zhFSXvRR+M73OT7JLiwGAJnVvp
Ua65Nb4gCJKoO5pkdlpUDLW66SWm/RE2B2LO8+LGGCtaYQs8dnT8ojW0Hjw+V04mbyT6+nTozcvc
Q3U5M4wxlNf6fLl+YCSqllU/kSJfaWjl3+WJASwZsds+09NMr0W/23r7g4Fkxh+eMLLQtPtv+caz
8suC1ok1Z6PSNcBngfN9cgT4hqCUMLVCFwGrtjgC7ViYyg6eJh3nhBGK87zTorTZEQ6OQso73RI9
7qvfANdymK5FR2u8nXCHl7Y1qfcc4I2hhTRJ469Ey0Yng4wFC/6vE6yGsOlKySDUUDqkNTTqdvNu
9WIHHNDo1J9V45kjTH2kRTnc2Jeek8V9n1DOlKyfJOYOHt7AF2znSI9GyvBkD61UJjfqXTAyRbw8
0HRpmN7Cba5qGdh0oiMttZO8OBXtFgwE2YIUU25FXW5mjb6A7DbYW7tJPCxEES2DolVwHUQbnqfi
IXrxpTNF4EVN1gnSLsEbL2tsHwHh/YL0/bISmL+k0GHVPRMbF21R+ve3ojApYdhRjndbZaEgzq9v
98eJrPYEIfsEVIEB5IrwLGiYMWjYnFZ3pJnG7WPVWTofG6Pkkh1f7XP1ewEuMUHysGAy2cCbkTM6
r8vERZzwZsfJ8+xgDETh1OVQnXvaxpBAdd/K5bUIt1GtfjVJDkec1LmC2QZ2lz2ZB1ScKlBAAWgt
IyhS97EbC2l6uX0w4iJ8KUGw7WNbhlZz0z2iW54IJ6dsu1M0bVb1F2R9wf4Y6E7BrkCLVa+3rjLb
Sw6MNeOyw+jsXnkLpAAkkYFx5cU2KkMzykHsL0Kk1NhXkgpmT3xPOvs7jEjtrcI1b4b/9t4/MNr0
bvDEvchjdALo9NBuFr62xW4H5B2i7YyaQRSlXUcNwrpWGR5Og35TYYk9Z3LTo31s7DJWlrLBtbjT
RXBw0ap0IrOMvJcVxDeGC0Jf52d5r6NM9MGkP28R1Hv1qXrNKK/9BxWW/Z4HtkiMGWSCzcKBWvLB
lOLXOSArXyhqx123c28IX5Xk43rjMn8B3JGIlBi3cojYSM/mI05/zJfc2cBoYt5GtjIkU/7OXqOg
5d2CXH484JXF5RpHv1oQ0yuuKeE57ZadA/j9FXZCJ4QLPO48kyFBfRAzJcPtTRKlBC+8nNoVIiDo
UE/lCdKaUxQErk5yBr/4IfAiOZJktBdI9h1ITVsUlg9azeTzzDxBjdAoWo1t3Pp6ftZJVGF7P9Zb
Wv/wsQgvM6dsdPzjOBIIgK8vaA2SjjpsFBIFbNTa1L48t0PdcYxHtI7asJ7GEuo/43hsJnnAXCZ2
65aRPRIqkrKKZmOsR2EQjjsxCcdUG+chnTa5FrNak5HyUGF6tRLVCnsEEPsP0uUpbgrAmxPKe7Ez
aNgwAB2eb2Ft+NklKx8wU3cR/+T0p7LGKbGuh8OdXRNQJ67gbiT/5giu1sTKsLklawGbWCbfUUtY
TSxi4j4jF94lIiG2ATrHZiUUB5wBjoHfedfM2jJmjEtRnuDaxLpMxg/usg+iNFZ9PXmUMCATdd99
+peJcPdLCSXmdozczihjU4jU8D/R7vB0+BPn7tH6Pb4mbcgb7PtKAWdIChjBdP+g6iti6ZlID7It
17xG/YWmbmnsAGt4XHBsnO8qNclHKgkARy2ooc4RrNvrW4o4jdBPVi26aBW3FuyM50b0xfTX6EJb
u3OT2OE43sb2amki2htcZrxR5yqXYEZHh783WCfgq46KAddp2IgCDvLdzg8OA8gn4M8DovjrB+8D
N6/4QFD136/zfURaDVk7/VGizWXqMNEVObwxthB/JLxc0Tnw/huayBq6mJbNiuXmoAkYLQQ925f9
+Jqu2JodrtVO41ycp0Opvr7cD415ahtEUk/AJa6h51tpb50n0jDDaUZd0edFAGr89zPo75vJGGo5
9I6EopJ5wgepLmJAioH027KdPlvRf6GuCzrum2ODXtPY+RVl0RkzYhDtXc2ONmC9KabNGXycA7bh
9+KrJj8itYzgRhKfeLBUfnc13rLFebxUqmz80jbcbhRmG1y5RbCK9TQw6xYnNumOaf+vFh4ty0+y
ykWB7Pr9Ci4MBYJ07IPWQgwaEnk2iw5go4xXOMsgi1rmGumSbvSBefSjesm/CQgL/ci8QbYxtz9L
6xBlNoCytuQI0Ru4oPnSsnbf8FHg/AGtyVgCnluzFv0EotxFn+bNy6xTpu/O9ewZqrdxbUwiHOBL
34968vMgzsyxgwKHfPEdV1eGskdxWZd+MqaLPNKcIYyZ6ezCoIhNykoCma2EAYoQM59tykTE6bfV
Ko9B48uLVwD+KEJm0ebrztPTicRzQU7DGZEVabCapl/2l0jFvCoAqRgMTDO7S1nPq5/T/cKD9IS9
jJMiGxuvCGB7KUTpHNxcXVB628ujUsysmNj3JfjM2Fpwh7eOJ/Ysxu4kYWhYaGV5EFMF6GqkyVa8
Bt6OK0NRtGeX/4tUbJMrZw22oQCE3tF0pB2IlLd60yfNsKCf1dAPV+qCbQ5k/ulYQ6/+lE5or9lR
A9copL2IjxsNgDxJidPgk7iSAbVSNM6JvJgiyyFQhr6iXS0iTXZMy/H7C2lr2gLHmmGmeRdbcEK8
Y4b0y/BmGh0cEcx6+cieq0fcXohrXhQXmepwNlIQ4LkJg6CUkr59ZS1VYC77UhN7FmRlPe5ZP//C
HtLNPdpA4LBDRNbD0AQEACzGA5kuGeVJoKNPvGIHQKl4Ea6+xCERQoUrj1axrNpduhMCixAnl6Aw
FEKykByTW//LkF/p8lhQ36HBQLyabrO35Kfm6n7QbdopyXaZ4Zmt7Wl7Fz2QYLMmzYJFH7sH0gAU
+KwCDYUMJVl7nq+Ssw9fmQ9ggTiSkb8wZ34kBmknCUWJ122dWZUE+21M19f6XTp0OSjuQt8ZC1Tw
Av2rmPPJNbj0pY3qEO4xnMEhnU2hP5IFNpVLpoBTI3OtRORlm0SbYTU1VL7dEvNP4KX9qyMZruzS
rGf0hQuw4oiQfCLdUO1dwVADdKWVfnLV7+4D9Zezu+hj2qPH9GheHrJaFTQDiE/PCBo9ALfbktvr
9g7yqdVXYBToe1SoiPqDKyQFnxYtfgMZhO+hrbpCNXXdrR0O5Atd/WEFrtJTlflqbKIDpA3jvrP8
uTX19/oi4pQROoEqj9/reuMsuvd2txlhk5JG1FA3oJ1ArRhJPKLBR/WH+zKn76Qh2VS0SHCbzLi1
ZDqkqoluotaNtKFML4AzQHrIXqu+rUyDSF16WDGgbmhq4PBQoysE3ZTbBLqDyA0T1abTdd/AN+O4
v2tFi1UFbhA2J5qG8/3uHhO67ASrCkDdTLqYJN1clwPA49/csuRVoC0u/xqiSy5HC/ODclwQNghg
/tRxzIgvnc0EMewE2lG1BptFX8/+//X8OTIvaSz4/ZQvrFEeB42EuCK4gxlgjNNLiFLSvOrUivCJ
VdtaSeqzkYVR3V0KgrIo0yMiRfBjxMLsyVmX1UUy0EhisJ6MsWci/+Oa3E2/tQDQcaaJIr7A+zU6
psCukSrVBflyZ5+V7YsTYwar2jcEfpgSdsVrVxC3JRpia+OZzLATH8iER4DeAxxWJq/IYoL4AZI9
ISHhspUQnS9Xzh7uUaQ9JYlJ+XEe0MNzyOGFmCzmKhtyk7cRF001XH8Ch5boWn+nx19moAyaXwa6
arc8/fDVI11k7VMpl58fe75QS4QSU4pyknUj6EKS4MbM9GWSxfUw029Kv9wgB/eLR2LFAirQWCRA
gOJwYvWVOmbNM1ajFBw3ePJCAVZRiLCrelrj5866m2DphW6MO5CTaolI4qqFd/86v/mdc06dbHjK
AOEfNk1tfToAdia+TCcGA5V8u6NxEUaTsU0EYgM+EeFTdOn8q+QeUX+Ziw7SiZqDA5ydoX/J/k32
Fi9ygUMLu9x1PMAb3nybnE0rU75lShRVtyW0Hp3DJVP/VV6wGKL1gdXDkPrvSCt/LphOToK/9I7e
xx9KcdBASQSFRwmGhsCsBHoHh4RU62yaZ08bTymwyfVUJ+ef3qfpDtdyqHN0kJ38rhM4aw0weiAq
V63otrWx2Ne03tr+4mS4Q1VkrYdn1EMg9GRDWI7V2RrBRC0NV03nWknfzVWDbBsMpT4vhzAXjy8+
7nDRdOsID41yv3GtUZPtYNMGAzMeeLNXHTQEs5JLdojoTQYuvGZIV0/r9Qi+j6GAvFKynb1HHPzV
VRnvxrjjGEMa4/99ImSRiO2hRCd/nKX+FSYI/kIc2zZfiHjZFgo6Cq18nhbIlZarLLrhj2LqPpjZ
vzuO47hxBBCkJUvIzfpu8+sq+K8kaU/3DoYI5V7hcRBpomLC6lC5eX9UMbu89uj1KufFe+5DjOHS
N3zxk0NlCbsw/vsmhi9D3qpJ5eM/JVVUHty5NhlD59ld/x7TomGsdR/y3LVJqnmEvXvDeJsni7oT
dJHn6FbrZRmcmB2/gm5notbX4Q7EDrx+fCiYkasG0EQ5wu9Pa4DK6AJXt7ga/lh4U1rhYrJrmZbo
wcwhneTZnISq/UIk+mPj2OUQPsMGSJXeVTgFJgFB8iI8AznF53cyakiYBzUKM7QPuWhJYzloWsf0
T7Ymkv+OTqP1pkoAYYNwiVA5daZU8lCpf3F28vy9Y4LtOqZNTrgxtm9sJfx6hiJD6huhR1ZjmyHl
DEMWzgDexs9zMtGub5BmX5WHVuGtIpcvoiZqvbpHVd5pQ8qqLwVpRzheMtcpTEF5IaOsvXfWmRyY
NvC+S+JemcoqpV5fc+7iBd+zCC4ZrarUThJ+b3P++ZVn8rCP6scI53ucdiuOwrwIomYiQ1dN+jrt
9BMu5eIxmTc6ToTf8rbFhuxzH9SyMrwxQNnGuYo5itu6ygvZJNEhxyOzULS9r+KYrjR/dWiJ+TDo
ooDZiapZtSv8nC0bnHLeADustnXaZtG/GUNsMSSlqFvaHMHJMVNf3oi90dmypi2VlxBV8qhzKej7
u6hTZPyWS6E6DBR2VytdDvEQsNRo7uhPIzBRn5896VZuL6dRLG7Dm/C5wqTGo6lnhIb7yFhyiwOU
iu+1LW42foz4auRboj19ee67lOm+luBTV0zfkFe78dzYwuAJU2WJalmPR0ER1tiDJN+SbFLrt8AE
OadAj2FzVYpe72Y3U6MlMJo6jeguUPtbMZz4BnIfA+YF08gSqq8d3AHBMDzuCqRl59qMcGpHPzr0
BjCZmcXt677q6TQh3cSDci2E3E+7dALSE37Ys8ly91DK7Fm4RFGqB/yX2k2gLuPv1TQsVL21lNRg
Cpej8oKuiTHLaIUncvQYgvLhGwDMrNtRMpBj/Wh5cXp21/5f2+/cNtxmn7Ebx5iYGJfmv5bOIgpZ
F84tpcmuhJ27KIfB/9VTbsqrxE5JU8cYh8N5FN9MgbbByEvBqysJLseWKD3l3uvCU1vqiVbrfnMF
p3Gr9MIbf4GbG3lXmtzKBc2trm6VRzNPOEYRaR4wCiL3OOAMb6AFjUxq8OqzK9A7i+eG0QumduLp
jDrfQ8QPagozEPe/au/B0kL+sOt/8H3qm7O9Uztw0qrm988PdEelAukztenqcd7FqnadVcteVbDL
pezCGZW8PKoIY3glfwatVYbH4t7wISxoLyizF3+dKlgKo5uXSE1JeY/gqWLS0Wh+X1ndezSykkdf
+Wp6UdCIAsAlJX9Qfzy+rSMOpefJuv015O5XBw7jyOg6mlXfdAD06dcwMncmqcKQbauQv14YRQrD
6WZwOd9+giuFvmjTEKBDvHmcy6/wSnEaz+uU9oW2ppIhGs+I9I2P/rTK/wNC3X/bw6YixukTD56S
i74GuDSsjDThnMQiKgLFR5HeBHHoVScW3mYRizVbLlG7uXi0GFrBnZGn0GN3ccIYqTD+IAjDcDS7
bDPJbuFNb5fmNJfMGv+hMjs7hKFyoyEgdDZoU0fBWA7jRiL1XQ+Rs6MrD7ZWn81+EWMsOuokTDom
aAt5ETItAoNKTl/EkiJoFbUB2GzhQtFpmRT74NikMNhXuCenlbynxMub2z+PUlNc4SHGlhnvSetg
mUt9KM9CLnFRWsCt0xxM0Yi4HuctAuBF66ISYODxpAldjcenkLnf+qUHQOUf1fzTS+KMYEkyAjz2
vVDwdIo7INL+f6qUbl9HbfqvTO0Yx5BLVee6+hA+uE3/f5nj042qV1DSDv/Cv/Cj2V/gnJLobcGk
CVN/Z5DBiwfWO+ethGva6X+7Bdl4zqfuRIYU85EyExLLO50SFvZz59UNhGQISg9ohTdmIFD69Rmm
xM+pfu09EE80gnogP/h3XdTe+fFfDzXdkd/o8M4JsRvww7KcAMx75pXtKmhRZU9OFb4QBDxKvto8
7uT9EqWE5e6lLuJs6z2tw1l6no8nVHdzfkMWwLV0meF/2pIKsbrt28xT7mzCbN5eA7lbYUJ44FyF
MlzpWgjbQZGc20AKtlV9iAi82c+h4pkcu0wdK2dyxCuWf2GoqW1uluK34drKPURcZ3hUE0gBuhbC
wQIwzxS4+xLd2NWTMxBSa0o3OQBPnSqDV3CnEiihyRstdGof7uYdH5pU4KFv00sF0CwhPkacK+Td
Wh9Sb9yn71XlFVvUxw71PYhp1ibTni72Mwgh84Wj/Fwwwun6tadUva7Y5nvyXOVvQwO3SliqshbT
RpxR3jP6/RA9gGaDwI9KKqCOXu6vwGTsNyJVfpvHtCdaZTEFimNZ/EWM82P2ldAx0d+9H95QJaZW
cGHCYFP+GI8KFkkPhSwrbcABT9p7VvDhw5nzj8cqopIEtCHa4NCHrpPo3zjracOwCNbI17jApMHo
R13UfIXhcKckQy5GaYXb9aDfPn6O2ZHiQMfJrJsf4uITptLXi74miWANAaX3VxxOylnPQNE89KVG
A83A8xeXVnQxEcOJxhf3HlK1XK81cTpZTZQIk88EjvkcjWNa5Fegx2o1kdpOXr6rKReR0udrKpga
xzGoKFHQnzlQCo+sDVRtqtywEiuJahAeVWxTPEuGfvqdPbEB05JwoRES4yyAntwedohpIwKwuFhd
3BJ97ObXvACXinBEIA400s5g91v0YZMJXGC5UZ/DNYtcXP6JTveYKNSEdO4J/S8y82XDxWf3Z6N8
wQphe0mxOIfAIHE20Xga+a+VAPzVx5wwt9Mpx7CpmAtQJbjqQWiWNvxijGa3bRKAHSMRnzCe2gd3
IFjX+AmKmI3oCWIMqy6KcEd6Sh+CK0rPmzC1YoJtqq4Pgo5aulJeGKcfQZ+9Kx2vxPvdigU/uv2x
r69HbisjlbJ47ntTjlVFwK5QiQeSIT2iazOws/gkmwslfZVUNB6mFTLM4moNIfxmwhk++f1FyMOr
UzAkOBR6Re2odu6VXcDsZaI37zXGDfz+GTxNv+4pURpczc82JbpJV/n4In6hasxxqnwf3LuAeORt
b0lQJocNUR3ui6A8YdH2CA9mqRqLOQWCm1jaIjs/hJkNN06dIF+NVmWNsCD+ua0OCoeiM3skIE0F
EOfpjzM0gn0yNY7564Quz+LukWSx49PbPZmH0vRCSX8JGlDJVKi6aT/d73iJdhPq6btfCAEVJgdw
LXTKfjUZwPVxdd2OiZhYlxV8LiAEXuYLXYomBED+Gj/EHrX+u1w47T75+TDDELyyWu4L9gcb6Ozx
8HXX8QTqjMw1rhFFfXjX9vLAYvUMMeFn7hWyyPwg/1bUXTIpN8VfkLJNIwwz9X+WZ47FRL3r8+5p
YV+CwsN1yz2dqOp6fhwQFWl67+1V0cI/T23D1Gzq1g65GsccuJNDRObnRihbxYzb61mzegUWDcA0
1Ejd09/iJkhe7Ro3mDvO6Pn9QgUAd3RXGeGCRVgp0/t/DO6StZrn9QuIR4SZqT1WpF1oNi/uOHWC
bTd4baHuz8Cp1QBqJvvCUay6KIXQCCaDo8FKA4fM57FYg1iXDbV2FqYp6Ab0hePls0pUYShLUzq0
BrUgO+6ypu/T5R1BwMGcej787rEZCU7CaBxLW8XqE7Cxd150EB0F1LaITsrachcUzHbYvJ85mUGR
CUClwgGwV33SycMDV+BrwX4JOXDDtBUFQgzepDBn01f+0hNb8mDH1cHrxjoV9UpN3ObVrCyziJZZ
MnWOvgjFjcphBV6JcD1m3p3EOWY2l7zzJD6QU2vvUTNiJTC5TkN8mo9FMurJ+bCl7GNSSEbF89lA
zX6UOfsQ+144xTOSWUuw4TfEIB/mS2CGhWkzN6n/jRfLPZm1AD12n2J3qmWI0KZwPT+AyNg0jEsU
QxEuLPCwEQDRDjTFBCje6I8H7Y3MIcMSEoAlMEams8RHUKAeotxWls3lMfpFntFxZNsBR556Zu9H
RREBLZ3tooy5gW9JB2wxtPDhmka1WqSvH4e8ffifFRctH5bCEAvdGwgKOWak4/mzGmScDMb/9dsj
xNeoKLlNDtnbPwl/J02+2Q/AiX7KgFmkhD4frrJqIgqnQ++3r6ZcYGA+7nIfVS+siWI1D86fXQ+P
AAI56Obim5kWfXiCXZ8IOB2ny3pDvjQhy7k3zBa8OQWCAKrXhnkWbUB12G1M59M5wF5TMIE+MI9/
zy379HgZgUOSkvlgzDm+GsFSbXAHSF3guUu64vPknEUlXzyxYyLoMiAPxoG4jRo2lUr1bmVNQdDe
N+T0t6MO+IrWOWQ6oHSmqdbyhQLjc0nkuPorCDOnvJgD8IkstoasjYV9MauJNZjTYRFZxnJUFI3Y
ZEx8ngRR7usBTbVkrtrJ0awzW0k4ATXO9/XQQkOLdWz1PjJnibYq+inF/nBajXp8sjxwRJCB3fpi
6YR3U+5I+4W37ODwB+5JPiqOYW1qHUUvToAl3clwiYU6fqOKrc1q83kkkJ4zoEye22AmWd4MNj5q
kJ0838LfBkMDRQg/1z2UpNxkinE9sBJ1PVTP+6eGhreYBUuW5mzfpAVCxAZYxPac/dNaVX9lvnve
dbfchN5INIks07cs3A9YqaUP6EJcazzX8FgKY1FQd21klcf6GOMXa23c76k7pC2+oKmmu9izhESR
ucssnVvNu3IBx56VhWLNBsRS/9Xe2wrnOIz6TIq6idqM0js6ZPTvmmRO+h6QETyDFnjes5H9TniV
PxCId3XPODhlUffG96EOULJq2dKmB+Jwy2McQVlTNSN4Szx6lyvx51Dn5MWWq7u2N/3mecKik7zj
9C31au3OnCeeFk95ytyHHU1qQHILbG6pVOQbRc5Q58FN9EQXA3E4Nw/qCZirDu7nz6VPGgfN2kvZ
0LwHZnead6MAHz4K8gPuF8RoD/wOJ2Lc3eC2dwMzhQcaYRdftIGORMoZZ+kUZ/byHbGriyp5BMYH
sDJgbe/yifROY6gdTcjIOrXjI6/CetWQgS8DJ0otnQDQ8lNQTBwbG39Pz0ynvdRVkOsJ/kzoSWdb
W84ytuHf1Exkl1aifmu7kIVzFxsGnvpvk41s5daOkE4AMwJUWneoRsENZ6YLUBnCKqnPHVyqTZsS
D244NpctEqq3/B9RrSxPMiTIvCAlt02CQrm2TfxCLxw3rnAFeljBW/rwS7uy0WLvqEr9LXFYaFl8
QACoSttWLtuMEz+zncFFh873DtMjH/XagS7+PZ1T7wJzhRgFFkHa5RVfeSUNFRKcrAdPaxQgkVD4
w9bFb2CRBG6R2h8AZE8zOmgbLRj8E1B1+roLK2nIxHjVuoGn3G5SXjpuzxbyCktSk5XRzoACbP2J
1vUXjAngOXsADdGcmNQVpZHA1TBvVJFZb6tfSXEctbd2M0DG1P2aI/tmfITadW82609lxUnYziu2
AINlfGrWJ+Katt9TmnWKNnL+jwFMGkdtyv2CzmIM2WyKcfUm/vvRS5parJuatNKUysTnJQzN9n3p
iive38miYJuKnXq+Sy95s5nzoGZO2aQ2dym6Z5oi5/rWLtMKsfqUlsLIE9iGz0WZT6aoXYoWrnWu
RjvMiAXVlNAIL5MxA77J4s9HrmsDacvrs53JPMIerj+o6a5cl9aWRupKV6DsnQ5/pgl5YTW66k+a
WOj5hbl7tTMC96BGmoOpBmjHusjSMg7YEXKAFEAlqe8UGdTv13dSdF867AtWIHU25mDO/57rcMHA
rEIGIRpUKN+hGwoCM2oGEz10A/EIv6V95BDxoOOCw5z+yhWRplF5GjyOuYoFGqKQ0UTimqbLgyHc
ANYhSlvQaAMnx0WeKG7A77l26KDLMP2tlTn7mLUYNIjBQV6JPTJ1O6Zn44Gw8MuabS3AUAz5Wus2
crJtpDpSzjP+oxeLbhdsOUhTo4iKdbdxT25PatviqyaP9gyF7b9u1Q5UaQRb3N9BSMaWgh66/Yz5
1gXNOwduxqKI0jvLEUvYgzqb3iUznv5JW+nPNaSqJ63FzUj5UViqlwYsv3XXRRZ1XvMF/TCGwWHc
sfZMERNkb/nsKziTsMyzxluezdt17rZPlbCT6dMk9EBYuQ6SWC6qQbGntkyufbHj06XMbXIwX9I0
9QiXHmeHG0gukIDENnLgrpLiXJKUUfDThrI51jG0fGNPlf1J+tIKvLLCqbO1cw/SkYJ0U3HKmN6S
7lOx86zwEqCbHiHi3vEoY95CNiSD5KNBl3l0jwB2tzdCFP0NKeK7UYOCDJlpdZQWYP9pneDsetbu
WcSOfPIVT0muY2um7NCYmfg/04D+LhFqtnS0urPoK1UeQfb1IJ+O+Cdu6KyFp5dCE1h0Plztuo3J
+V6TBarzXcXj1bX5MLdqLQTylcx19uh26f7RYy4xzwCAov7U0rAjSq8fPGYj/FPRBIcJse2eo+o6
Vfx17dANCAc3cd+bQlFaWPb6jj1R9lhkNgikvnPJScRZdvJD0fGgH0tcmAHwwzcUmExtmI4bKyhq
0RiKqXo7r+tG4CY79x4VMk7yidfrw05SnP1pqFnjFp25c6qHS+7h5OdjOFqEdOPuMcBnMkTj/QEJ
TYVKv6TECrrNHcciDJrRRDf3a5awZnKwNnAA9ouUCO6hIkVo0Nkof8qQd/CW12XpczxJCmQl6fT9
B+PFuwzlDFexcfeI013Lzw2ZH7zU5j2NGtbkD48Z8/ThIwp5bJXEYgMr/VwI6tMPOhYiBcCK4gn0
HXb6kTRW8O+ZcWAXVlG3S54B8GrSmnHuLXmKdRX8yNHwnOIk8E6aE3IK7q31by5wgrOokpblr/V2
EV/vqDFMgDoi0nu/GOmHafo4rEs6P9jQo/oHL7DUpBTTG8Dt2YeEuvqZ2pm9Avl04N+7KM1KT8Jq
jD5BfIt4aazu4c7n7HguQlFqwewqtmw8JKXl9hyXcRvb4fO0imtzYf77GLTgJ3ssMGOBpXc1pJjO
z3W5UX3bvfYCOOLqdrqh0mOwN+75KV8e1EIwnCNFvYzQzeodVfk/UM0f7etpyXyxvzepkqP37wt1
6Nlka8AV1tfCTCcbKEiPhpPtCKY54s3iK2QWI8BOn7kd4asrzYBhDlSlbQ1soQ9Q9OMcfnAicJom
wpo/ih+XCzwiUauFN4hfu2OTXIq4xlWmlxGjBDGeKU4immms72dVavwMpcNHCGiEFw13zYbNnCAn
KyieWDYOeg2hiFX7BXJD+FJuy4MZGCPP5qpHfkTIS4k1si7qbrDwZelfWRXpg4RydmouQlPOVUuT
Dezsbt0v0HB+SdDabwtb+y0fOt1sfDDlb1U21Q9/ZSmjRrAbl6SlgvtvX83cKRl9pHLgYqqLuJvQ
4m0kbsEsUr3v4Ki2OBUMW1RAE5t2jJ5ITbN7W7Bcr0JcVBcQqnBE6aLrXH8MIOhAj9Ux6yKUooPj
vr+S4ZEJ6HVc2ACsxvaGBcX4+hYeWw9oEV+rs3frppAjKZ2noXHJ44GnAPKF/Jv1UBINu1vpKTTc
r8O1HsgdQuQiSfDegIJzYzM8cltMu5G/uLnhwvKrxAxkE7ajMr83OIaXgKaEU2qnTJOaYa4kMlLf
Ynra8HiImVbjdBtSUMIkV55twDbGhxfGd6yNLxRTVqfrDsOhM3a2I2g+HIF4AcpYJ+W/wXJHI+/J
Ob1FvhXHAWMwy02maljHVlATJYC2gShKCkOygvLCycdtosvf1Jdk/L23iWRwJrA26OkqiH7qfeSe
NHX2tIEGaP/3pWXVMAOFAd7GRnzC/DCZUy/ApoLip3kcYM9Wguwiq35vmLPeP6dIzJ3ZUi6scshn
cbztd0SvIs+ZnSQ+d31StnoTx7FyLJG9ncNOiadbzTJnZYdr+2zLm/7U+Dtu0Tll/DhcHTNAS2v5
WhfENkfyqLOmRDD13j2smd4FKjEnl54XTsUznjCdT5QVOG0CkO2+y8Il1Nfyvs3IQbSDERMTff+x
W0SNCkzFvfezRWbHUxwrVkIUcsl4LBGEJs526t1E3nNhKxzjN3i3N2GSOkYe/Hec3kMJ8NLnE/z6
eG5bUZU4rNlg7hix6VOKRqm7meAdmaD6yoXYNHDWXr6U/MQL1qfyvO6RChkdzQhc2RQRh1q7VnuU
tVn1pBDD9Yu0mCvqTnOLgqzG/PduFPK3Sb9Q5qAR2d3ZRk7FZ83stFUEcmUnVkYUIFZHsLw3EIlZ
WBgIkzaLT2J0YSnswwRLyEhDWNN9DFWnlWNfaucPo2KL6FZFqe2IedtURdArg/eK7Jrwk51wMMuC
SmTU2+PsgJGqATmlIuOTbbeQ7f3Mq5iw7EHSAriBpMXh5LFdo47vJWo4LHlXghz+L8jC2jT2Z0gm
+EwqP+nfHR0oHGVVwMT5/yQlF6++EdsIfWjhCJEquk68AKBf7kyy4xV9NCzrVrfYyGklpJJ25f9+
DyG9AoJ/MflgMvh5sin6/Hrh7zBXUuuD4MhPIgpaD0NisTIkIWjVfKNOvjPBW35cwhJ20EcGJbKn
PC0VBDeOqT4gpNLoN3Wl6IimFGzk63mSzaZwEE2QTNfFBfUdDuDk8pP1eziLGboyxFDyKG0rkT8Q
ngK9KZG7/bsPg1T2patqqEQFinaXZp2dQlS9E/YVVTYhfQm/wBDWudJkoLwfrTidk5F8M4y4pIqG
rgiIeK8kC+P/QZFq/SVPeOhL44b2nY63bnsOGBMa9Sq6sp5vvtpRWg4pU/xjhGK2eN+e7aJivgWA
4P01Jxpld8mrJRlHtuxUNIgRQQ3MsdKPGqUFRAut00fB8ZZIv6bWEQUdpmg32aSWDZGZ860c0Roo
qYK9lqfuX6W6CTaun4d4ZkkdwJelZ176m3Z7sZOp8BCKUmztukxi4c/0M4EzzV6Vv30v5VKmxwgW
GvR7RpcfoC2wv5Wbw34dwHqxPwpGU8dIcxG/Jb/qaJ0CCVgAuJsh8Fex3xmtQEuy7PflvGXGtfsL
mFWIsrohWAYLUm7LuaXXQefeB+Ii8Qm8WGeYRAaEo0OSCmgMY3p21BeVUVzQq0vWEbShyG2qdHFZ
D6raJgJTKEZ4nHfVPs/DsrBPkyFroBcuv8bdH8cRYklYcu8d4eKIEtA28Z0lVZdJcrQDWKv8Vsd0
gUkDYLxnEOUsFH3iFcVenoXZw7DC55IXgHRpQPpNPAxBOltMUVWVF4ErGmYQzvo+UgBqed6HT7AA
ERwtebIpP32wzjQFhXhFyDshVZZadFv2pKGmsROPIaL2CcFqSHGZ5kxiOrimthTaBrn8/+5q4oHb
7UidI3fh3V48iRSleq0IyHIJAzhy/UMoij7gRYT1hw/aQBoKOoidMwc5TS/g0LxoEXbs+ZDjJUKt
vTLJ7UaSqanNAItRyi0Uo15HLUx998jp+1znDBD47YBm1f/YjmipCn5t540dx2cwRbRH4qBhqHDB
046y69DzOTJo+q6uNhaSTRNQvfngWi/tBtOFUBhn5Uv1DUDkUmdhZS2i0s4Miwx8me9lzWwN77ZT
N4p3eykiGQuJUx9lM3a/4RIdeSwZ8U6DBbPvWrI7JqpvPcyOTRo3aFAElNubyeK2q+U38BFIoUyf
9lxw2b3+tC3KfS6qeyHfyfTK4I3btdxxNIJw/qq3HaetAUXW22pE6ituJ81Z2tzxNeCRv2iNH80B
iqc+YAn/j5ebkxiSfqT1gdv1hT4r1X1hukQEIR9S7ldKnLXlA3pfFrw9XZcPyK9b5q1pYgU/dZq8
oGH7q9WVqailzOmjxiWVh4v6Cf/tT3eUrNe4ehpTBttgjrAhY0Z5YRYWP5w8+ACRL0nOMe+XObmK
76JjFyE4onztT870+JGlBdO7TkcbB2Ce2JWvFLeSAjsOW6s1v6fIvWIjSzWJUWKgh8kR9PjF5FQz
LQGGMIHzvah+fuMrt5zPuCSF602/OUFkll566WhnSEeXO3Ec28thZ09N1HQyeDfz0xC49BZdXOoc
KwPLCODjhopZomU+aCe7jUPc1hQdF0Cqv540zvglqD/iehrh2fWKngms3jJyl/nkLUqy0pjuxeQM
000bqv148ss6WLeDIdt2KBThVeLWOWXCnT/c9x7fsIDXGyxSwMor/aV9uByXnNNzER24DC8QBI14
RvZKeE+HENKxpuB2mprbBI8OYc3cTZGsaZAk0WkZvP/dVY4FCBWRRZuuMwRzD89ZgWycJZP+70XH
pT6Mp3d4gBhygxy41iosMb8pWksuphJKhDtdPD4SMY7hw51viBt47e8JvgIM/xfvwNI/L47/Xhk5
4pk7xvLjCF3HALiamfvgtMxx6n3scMK37vc1YXsbkq4GLoAqxmhe+mFzf1ISrKcz3h9JGMW0SykS
jfXMC2c+9NcUAoJIske1XYOJofVsiSBQP/S1k5Rtyo5baoaJ+Iv+hmCdbfL/HyYM5QiwfyyyZD99
9w5Zyc6aR8kpj1oYOzcLAumXMgZcm/QAog+qUXEWQXwf/hfJpfGIXs7wOJNssLkxmV8x93IUWlH+
+t4kRcNPwwi6GBYoB7TwjfZ94KL5nEdWx0ZUG8KjG89KrBgIbisBtW6GnoDU/JFCmEdeSYNWyxzJ
YRxEAcfLCRNHgWv4vRkR1IUUfdCqAgT3VqxCbjjLI6JEs7PSU0mAYuskHvDrvBuy9g3SmRw1R2rr
1zPDywYAOUCX0+QBQPU+dSyhTfqDSyRzJowFox1wReSwJoY0o4lR+cjYd22Hd2cjBwxpA4aTrQ82
ffnGVqwj1G5KCG97OnTnonxb3Wy9KHfiKEDhOlTJW2O0hyglF+B3FgKUAQ4LJye8qmGnB7Q26Gw3
0QPB00Z2Mq6MR4yHglYlqRTqAckAWpO2na0p+7MwgvNFoO7jukzO+cwqQyhVZe+ZYchWGmnukGYG
GTwqc+efD8pfCqmWNOPDiUkk0u9kMKOHPzHm8/83hQxUTDqHZakszkhSvfeSfz5iWrp/Ye0meeV2
pkBCsRfhcoKQf6udak7J6lP1SWedGJn61h+v1nAHPf1VJ7JLiHUo5YpvbEKQ4EZZYU0mRjRQUGIc
arCYeWmq4pJFRhd2graI5FAhzvUDimn5CeKxrBcdRue8cJ3/+ghOny13T1ghjQapgZsvMzPrL+g0
RR1CyA8Ba8g/a7foda08ZW7vkkG02c791N5BGzp27H6U3mHjwOvNhG3CbIKz3qkoeQYWAZ5ZhBZG
3URZNkB/i0dq4NBYuSHVFuVVAz2nZ9+Ur0dE/mw++JHhIDkWaSz9bU+3IfybmlS9bo3c4/2S98nK
ge1nAoCWNpatwVtgMHdtAUdr3QuMRehd7oWNtznthYl5a4sQ2EHFj6VwbAoQTFu1tjzRNL8stitc
r199kD5MQw70tWKQLxWv9BZzpUkYTbrXpsXJ8lB9vc24gqBQ+uOgjm9DdxVCObhPb25VPqEa4EKA
0FCCRyUH4qN8GGJfqy3+5RmHAT0SYHu+99/rkswHbKe2qQs6TnkP6xoORTLkkw6F1tYun//VDqpT
D8G36MSvc2A3y0AjzT2y3Q9twU2DbHdwGPPEB5nBzg2eHHjFnHdVh+LgDaoZaOAmSBwpRegIA4lG
U4UWZGfuDBV1Zqfy57uI0/+jSeDZB+gg64QWfryDzvZucvqHgpoGlXRyVQTxlcJ2G6g6mNyxvULX
X4u7LepUD9zVOGxfhHV1NT+aE81FGEbgKsxvsO0Dsh5TrOKzO0CtqN5Fjo5QzDQ280iLXmBvpFKW
cYaUCbkDuQpveFl8h1SxzZlZm15ZI/U+YgNusXfO2yqHvCNBBhYcW33AN9ELii06ZVjilFyQFfB+
hr8sqv6Y9d7ckCdJAri1qc0a0B7z7x1N2MTQVO4yX8UqyMB1AeN82+uIRiHQQMqICQldnMRmr/Bc
TWnupRV5Fv984k/MKD4csnoZzYr+JHS/rzbINXVcxafqfPBtVixfIU87jPUK5zhJUFiuUDIlxDpL
z42NekEnS6LvLsy1h8BE9aE13KhjFtZQhfJYgoEteUVKJ8Lk4ozfD4Up61QSnFis9Os0Cg9VcTSZ
8hG/1faxntOCi1GJCRNSoEJffNfJY6XOpJlVOqHcFR/4yCn/Z+P/FCu86YeD7dxA53/v2zNbYGYE
46JqQTvIAk7Q6ujCgFZNiDI28IfICPyuvkllkTS5a+7bL+8fSGSC/xw9ZDAVEpudKbC6JxR/7Jfn
tb+yV3zulpR6HBImfCNZnujSse1I4udPUl/iXB0gDUPBPfPSYiOILGpDSOcsRq+PtmrsJF54qq1+
vY86D2TUtG070/TTVSpeW2TrN6BAgh4kchVIP8L7ngvTJ8xa+xBFq/RAuoMBiTZBospq5XBqiMHl
7JQkvtcecB6DJYMu+Cv+ZSzZMis1YpkIUylTGKspt3eaFb+t51Ew9Gm9Y4SBqYth+UTQ1c5tNJeo
i6Bi7J9dq9bT4YS3h6LIC7o5izOE4rPMo5IwZrgUA1RAoHeaOdv2MoMjb9JzdW/QQidOZcvWv7ZV
mx+Wm8GZOcdN0jQogLxMlJdtHLVgORQNPAhE5vdVIK2wcFzJyIr7Dxj3LPn1hIlbiDHgA7SiaNIj
uwYysf7yblkKI5BwxrNvhZ8EOBIdQfMjsl/442XIVmRO5q6EbSGnAl2C+6JRaOsTfuit8ziLhPtu
uBMJ75gjNj3HH4CK22PSShVhb5W+5N2iICX+OClm9tFaA9q3sHwEUFEB9gdKVogKhtibP2NLTw8o
lT3Fgy9RQBjyJl8j6qa3tYUmolHAUZy2aaTQdFv0uHyBCkMBs9EKFsGMzEBOohQ7VBo9Ch21TDV+
+KPMdfrGtlAHOP0BL5DZVPcZ3AhIPKv0QX8azjDYc+S0YgPOkvUJukJpCaIHkOAf6YZ3yrm8qOIw
HdUvV0WDsbIDs7liVvsYNxsVVxe/7HRPhN6IXUQBHpvexXcT7t/elksKKv3NmpWJDbplMc0jAL9j
7k+N9QG2nzcmDsNO/REzPf4KRmkFtGFhx4iZHSp+eYrYRkQiEdD1IGerCCidQGxZwxIClJ1k/kSR
WIgsZp/cmyo+Js2fk+Tkr/egPkutq/P1bNUVa/ppfVrK7GAY+g3tLUben1y+GELQfpkT71AMQ3xb
Tk7Z31lLtvYsPNmUvcJmc6u+VZC2tZwyEjTHmikQZMEOhxQodjX8+KGvvqv1PvheaZkl+fhEa8x7
p/ifWQaCvZr/oX7zL0wHnfb6CJr2t53KAE3ZYCWNlIke2Q5hYc5ssdPRMRhFVdPC30r2xQmVRrhO
GtOpvWQM2/VbE4CZLtdYjAolIOTM0CEMGHDjtx+FDsScd5SD38pktD/O355Z383IA5LDRnToBARO
t2oI37CvV5a+8FYySQ7pjmD2AdFo5a6/8US3SoyQGuq+tRqxkVLO0c9j6NVGy3jyzLqrNgdSuKfO
zwOiy0lXhxqDL9m9fYkR9R7wQkInxUkCRRomNaRjZNqcioRo6rV/2XRdlFVCtv9QOYlD4TfOv9fT
JopQkIwOZmhOUDooWI9iErCYX9ol+6IfyRe/PA0m+XtyqXsQFVivjn82j5YiGhw6gX3cVvxLVWGD
dQ3fMb9j0/mRLtWHQZDQhTxQXggLceli5mKYgvaSxaSQSEQCgkUwXwsKrixhFr7PFOky0GmYBE6Q
t5tiMgvxPFigpd37c4xhFGEX72f/vw2YPVIxThEZc/774i1Yr4PAX/9GQmdpmgrCZe+YsrlHqYI9
EQ0PbYXYfGEyAvAIwpeK5SMuvYPYOijqfpvc3uYWp1nZZE4uq9Bv5Ae/6OvuvFcDp62BfHP7ZBZL
NuOKIyxUt12+Gg1DuyYiBlp+wYeOfWtE66YnFETqAYSAecZxmBYmjtpbDPAq70HCW9fkDT96bIbx
bwNfrRY2si3MbTkdNiDgc8XBCgkO/rEG56TgE6S3m16b9ZZCMif/sqkRS4HY9nCD98mM5yKK3NV+
GDjbP4Fs4Dc11HSRbZRb5lsK1nNASja7zga7K+gMCjptUadCT3kSxS1ZdpfS86emIA/wm0EIgdrx
BQhGraWFHvkNDL6hkWgM6cXb7eyXgdH8vAp+Ae1YASGMWGobLeB6Py+c/9+xgFvZaaKwN3YhhFQ1
DBEvjFnf8NWT9JB5KAlrFv4/uTEtDyFJPDgKmJDYo9uYE1+MAyKSs3uNCYbpkQl2Myp2m9FDkM1A
/hI8IGGWMpyzVFVyTwpjHkaVJgZM2jzje7zQz4Hntanes/vfw4JBekekUXsZv6bLr+35qS5SVt+y
GOPac5J6nJP0GP3a1s87HGWZ2hYkStkeMrM55WF6eU0n9cSDKkv9XwME2PAIWzwftDfFiyY7T5s3
qyoethBmW2QAEKF8D4hOVgPggO7ZWbNBeIlHe9bTzYjD+agHJcigPpyK4aQQmu1PR16ldZIOaMWL
fQNumUfcmOnRJsfTAqKbRlIRvbhbEtDDJynxtAyVgdltkgl8SVsBWOBDvrKy57hWFBdrIDcnkv0M
O6osmSBSrtG0kawhJseeed0KYlRrwDsiOLnX18jAMIC7so7SB81Eg2GQZy+r/TxkoQMYSBC2JKgy
pDVRaWZtdqmA4r2HT3+CR3qaVz7bUQO3s/IAki4vJq/27YjyBiJUSKTDrufBtcog3fdJ2itFJMI4
KNMQ5EuJ2Eu/defpyFWnUyQKXdP/hdsU8uAgORNoiLZxt9xSZi2TMHOb2QkSz8VApvc/rmztlkhj
1yoJ8NT9msMAlb8Noxgadyga06nXNL6ZtcWIv1ch+R8+qc6AfFbBzOrW4BqQiCl5QDf7eK9+zDkF
aQK0DfPEw0DwybuHElar37meZF0gZ23+2rBAEF7/4JkvdglDm966n40/RZV4rHC1OMZMUwpoLUIT
VRkOwozpTzR3P39xHTk/VBv+ge+ztiyyvpsWne8N2K+EjW5bJbuCXyFYRF1zGXBpNhePttM/JAwT
PBxkXkL5MjUGXUPgH/VbqUPIcL6KWrDXNupwu3ISm/+qjjR+ERDgZzfO91ZcRvp8tnc0+OSNcaw0
ukRdY1T0O1dQg6qvrRBkFH828TUIAhlFSjjo8fxxuE9BFuw/J1n+1DHqvs/lsmgjiL46k1BjBG4n
aiyacyPI3fPxs43LjdyBtGlfdQQVENVxoyG3AVhjbDd1nVD7W4vfqKSNa6rKtPq46chgz3PfqpL4
AlQZolzs5ZTwCW4cGDszc6SzV6LGKhevzGnoQmYUbyzzQSJqQZwJkZezJUUWdB0XYS6WBiXERhsh
8c9LFdUM25R5NVCF0QJGt8E6jLccR4uILIkDPdDYmFXRHIRCs6+DKBGZl2CYUm/zdop4Zch5ol7v
iy0jZZo9Bkzy/i9punLwmY3nnT61gO00dilUu1EpzJt3bMlWQMz0NYPvTn+Jde6O0WcPuwiz7e7A
KlRXqwyIUgI2NnKGv1tBTadyyfRjC1JsgR6re2c1FVTJFuHmWrWl4pAJvyJbPu35qjRh43pN0nQr
A/88IzDgJzlVe4MTUkMW+8N7vPX2GF35XgYFuU8zHa+PA/5aCsEtcXkB/aGBRvfyeeN1lUkrmEa2
zqb1floD6dJ2NTb19Yv8469z7+q4TeA26qKpBxvjj9KsBiMoljyOTyhtAqh95iRwSuI8YMWnKxRc
HL2QDInM+KnF2JYM1Nq6DJJoYKi58E7C08wuW/DnuG9vQlKvf72O1p/NcYvJI+SU9ayeI2S4vpVh
8+4mJv4Q1gFFSYD7JyhSNgQQLnr9VxRqdmIjCyK8uD2lSYlFmzqCNi4EB8Oxfb5W4uuMSf2+8RpZ
UhXdqOM7iArv8IOlhSqYwk/puiu8XsuefkYfoHEz/XyjNv+5HPIXPo5rF6jQVzO2YE7utTht0Ztq
AnVb42IMAW2gkrm+T/ajHfpob6kRShEh4kLl53VhHUKnCkLGVzfpDIe83DIq99GacDKS4A5LcFqZ
weB77KTSC8gd9CJmGzD8Iq7m22pojgPHO/fUbd++hgDGmJPS7X/fB61aehcBd9H+qWr7WQjHUhqu
sGTZ9AFUWrGpIyZ03lSbGwQnSIrUFiirXLXGIBeknWGAyBR88JLaTsFSp61zTeKCPnDSCkhuoF/n
tWRB0ddBsA4XDCwuSpuwwsFICFKLCtUvVJdqYLxB0uwbkaE6W4AYATWTpb6k4Xvi1RqSC+k9fN4n
2RaI88RzP7FMabF2RtAslb9iEdkcn8F6VNfyJfxsZG8INFn/TojlZ6sWT8g+AeMKpnecidv+qsgm
tFkALBf0DRYFHSelEwfmIN7sTYNiVLyF5mcRBtpC/cptmkkDfvVA/KeRDDjYAPrjgCKQ79i1rR9J
EGYdLycxpQ9odM4eEaQHRhzNvESQHSbNIK/WO6CgcG2P7ILZNrGdYE8Wj4txrsyk1HeVNQ0Oe2qA
VDYyfC21LuyDFarbrvvds8cR83AtyrA288mWuyEIszPhozzzkFSgbw0+lBuwibhqi8HE9qX6G5sk
seMzFAFOY8qfwLjI1QfV4Ln9Wpv1+EmVuwht49ityOBp5PQA0B+r6EjWLwZ0ICkmYfg0eSNEdHf+
loDGwDwuM+TcoJUJp1TYynDUY/hoH6HDBuEE3nmEJgwt36aDRy4bdX95bX8BnWzAGkyBThPeb0r7
ruARTPTBBhUZUUgUqiVka1mG0CPazB+LgIuclgzj/x/k0LjinJIYL1K+l8BgLt9oYxeLKgAmIRA2
roa4mnvvdV/9f+BWA38W5N6S4ckQEcFSzB/JsEVQzxAEBU+rj3E5nqD/fWlRbCsRkHfROiuvUpBF
8N8CQI7zfziXx8EnVrrQqj/DvqX1skMaX9OFxR178NGWK8PoAxmU67qBNHPHKEhGMqfeQQ8ztZRY
xyb3pGaAYTRsZ6KY8PDlfbW8Brj1ESij3sU85JxsjiVl8nyqIHGf7CWWSWlchyfVgsXjZfBTkfSz
Vyp4MoQCYnv/9KOvHorwotNmqEpji4lKGa5OfWqBaI112xXC3QJRQJcUgDn/2ouuriEdM/VHilxy
4LF1ch1VTVl/nPmvQkD1cQqWxDWmdFCH69zmIwdr841a3I/uE4X62/uY4Y6LBbysIC+Vo3xIfmB4
sVgY6VvNHLB6JXRGLGucF+mwSPv4GYKhZGYIofnYVOZaJD/xRH1O6N/2sxJhO7GYjxebxqTu0uVG
8yj9d8HO69ANTmuLQ5NC8YeIaKtuFvkadkuPRe8dgHgZPi+gc4ERQs3gDAG0CStT2FSrErf693au
bPBEr8dI2mDflXjrCxbB/8HorVe7yHP3ELBUcZCS2fki+qU/xMl3fqTW6wqibzWI5U3JeV1jq4Pd
Bu5rZOWZs2Ys86ydgyYYBqIZMq1cwkKe+McrUL/kvz4scVVt1ks+hKjRg53BeA7445Omff/KEdAf
HWeph1ubGYzPM3ixt8T+51kMdXd5011iZno6SXhsxTI3Kq+sdumz0oCG4SgyuGjFl+FHfN5xxawc
yrfa0+fNwQ4mCZsNYtnqFsEcYeGcUIr7cZex2QziW+zQuitcRXA8Bgj9Idk7OAGRT1LFsdp6p6jC
rUKcNkdjY/D/8akInQEZhLaafJ7BJlf6ksEV3j+bBWPdM0lXV3i/te/lr6eoExdrRdWTCNfa/ZeK
eJDAfqZrvAxwB3KOQhYqmrOQv3zqjPBW4LwvjkW/dsVNS0X/UcXrhkP0RTgcK//Ap+cIlQUj0xhP
E/heosmmiRuGPUz1aB5BTIC5maQHPmFzk+dGzZ0r7ZbSHTH7SEYmasI6FnVvDB8Xh/Rn9mdtRHyN
acogxaboDyjCOyJgMTKiTCWM611fCDa8QoskGznZq9F5+LEBrlk6yOIBFWh1T9zqtGYCTcQRSyiO
E28YApQ8kceK4vop3lZE4VY2/Hb/tts8hw6fT0PePmjWEvnfCHG2v3nYpq/hKPZh69cuVLIlT0au
aPziJMAHjPZYgIFqQ1En2zlZZbLpUHuXB+hyJxsoxHRZDAkALr+LkLbwCUn/TIT1Cd+59P8AN45o
TyYwYGmwFnqBFM2C0pzbtsebayKK9CN+FBhY0Zhl+Ealhs6hbW7RxDx6P/4iIe//OngvARrsmw2R
BtgYyZ7SNxQrwZPgsLJG/4tmjT+dVYoENexcYPB1UDkEJQu/QaJmE79wsp7enTowSSJUqDD9F6Q8
b3N3JOQiL5B4VaelvYpB5sYk/+dmIbNDpMLHPc8E7X8Lkcql4CQJGWKHBPxtwK2VSTTYkjdOodlX
xIePVXGvnfZrJ9fotZbWHXrqs8q3ZJpj2r0DA7IJ1+BIWXSkgnXQrLIk2CRRUDa8tu4KdBy/Q/Ld
l/8mdk7FP/LvIhTpsCUNk8xW++H/CdlcQgjoBnwTL/JisksaDdvCbyxzpB7HW0S2pl7zV5HXaWy2
ua2chZVnaBxPRAPmDIW9Ys/FC95McZHdiVqiG8gmf8Z+FiWV9FEtb+2CnfgQ3er+/O1rV1qjyrgq
34NBfChlbqX5g/PaMBWKkRk92lCy69UVNmNZsGwhFqQM/A8sD/OwrqAiem11ufbh67M/O22wRCFU
bLLnAHtKgvnlbXDSzBLjVtOdrepwlubz3SwuTNyt5P+qneV9Rfj1bF6FqLJREXR2dK2CpfisIJdr
7x6w4wd30+q8COp3F3IF3cBLlqpB2zksSGmkU0yVMKHkXQfriR4yQjQFv2hHs/dIoVaedfjpug7K
QwuG7Zk/1XdQD24mqnvbOsXehF19jXPitz50UISHRHWS0TRJK2KKkZ03gqqrtJ3XfPtDJJNpGm2h
nqUaICLPG+O+BJg0JpV08xcQAg0gkdX0ITLA7ld4M71/wLaVzM9PGI3Csr+WWDZ+EdmZVGhmFAPQ
filLfX8EDud5bX6OJufj2YAzzWaLtnkvhyadxrrNoeCw8ArBHhSgNohG5GrpKXmbg+dOivI8bAGj
80GeqSsgJLFXc/Rz7udL0bXJEaVsxsm9wh26vseeBKvonWMscbqweEaovBoRJL+Z0IQMYr9xZGqY
m7Qcj/6sWmEShbsoprwCBXPIXpNa/xcaHD8/B/rv/1xGvB5ydn40rbemrz4rl221HzzSWWo0Sj8P
XZ7P0A0+fRORfH125VUPsYgY8L1UPskyf82AFkk9f9ERpeuAOfdtIuqHxkAfPaRR0HdAKNoSEX28
/tTEhBZIsOxChOvCgGGBisb3BdyhxagTNYAX2xw5q8N7hLxp++Z5P8rK3c0boazdB3mXfievJB8H
zh6XNq0s6Ty+Dj0zT3uCO/zLsHisrUFJXdkCgs6k8sNyRXSRJ6/EUQu8jj+GvbolWhAN8aJVSpS2
8RoIK/9D5wMIKNXgBRa5nHti0JHdezEWRGo5JiCQ0ReHa8dTlChvDuvQABK7kgsP6H3MpixLiDIL
oAFrFY99B9lfSE6ZSrfDZJ/a67qwEA5O/P9PInGOfwSkGbJjsyRyE7K6P3B/tE2jhJXLEPHFRjx6
LR0e3R4odoRRA+CheXBxKazjJNMelZaZpm3ftaSZofbtYaEIfrsE77Az88Rvp7oqGM1/ePGVLvxW
Psmizmc9uL/U7+MO+h8Dqtomzsz/y1yCq7yOg0J568iZUnYMQNRUP6vVpmdR7Sq7xmMe4hjf2aQc
VBYWgc81nb/WGq9dZibCnUjBNQmyDj/dsKc2UtfbK8sK2Ahu8Nl51Vcv++dVzpnrTw9mX1XnxvXa
X5d1vPpEKKduHq+8XplOqSKzYaKe4oj8hsBBdJprhocIu2nNf49Ky51JBBCqs+jZ+tH5sd7ZUHWI
YazjYHF3QtTO+88ODifW5bKPTiZ3Fff3ZxTKLy7DyJNSw20engXfouSBUaUNDKCDwUlkl6BUp5iO
ZC75ZwnfUa6bQwYpSV42CWHqQsMwi9HJG7FpTbU+VbPl50RN+V5b2Xf9zwF/S8p5xRYkQ/if5E63
ydO0uQ27wKEFYDSd9O2GnMSKbhFi+MLnuExpVglZhwlwSTTYh0ebpKJ8iN/+upsLaEZxGv59ArV1
jdInjeP7RxOTJSPreK4qNsoE6R7fnFixyl1HnhbK3HCYBZqRiSze2KV3OanFfaUYbjJHb1+PKF4D
2V3fWfmwNWzmMItPRSpstdGhwLl75himU3U4+jQsfd/h5FnYuCRIzCCebtbwK5J6g+S7Z1yDC02i
OqVdnEMcp/3DCGc65lrRFBeDMe1Va4u2MhrEIZAQ0fl8D7PDOhCGfadZ5Uy78B21l24lD7xmT93c
ee8Z7n6ltR/2yTkPeHkpaApfzSaDCcmvWVnDSj+B5jw4NpcF2bhSpVBz/kGhRk+p3c4tg2V+7bul
ipx5/SGQTRcTn7feAP9qGoD9SWyXrSBxeysjVZiaLTyaGfhEjA+VlLB9OjzQGqpdpfwPWTpjzP3I
VXAU1sPpfW6cT81F5wnodsHaGlCWJ1V6ALZ8qHMVT0jaWPJGlBRujbUyVIc39TpdOxpa32eS5Ked
qkB5taKsFUM3QxpqC8V5ZfR70VkMiTIMBJQv7PXMw/N3lRyLs9h7bYdJeGmftlK5LvHhQFIBfUM0
zGVGmkarKd46t0LLHTl8z9qIRayp53U6pto80++vL3fIB7x2CUGtN3/d0M8USdsBbqFv+GL93Ef4
qtDFc2UDh6G4+Z/nG1HV/5TcP1zlSfjgvnIT04EEYmwqDiOKHCxEI3OHEGBb/6s8OXF91aT8CfEv
AWbCv1ddY5nKW10tWWY0Y03HroIW5N1/bsKxEgjhXqi6Vbm2hrpmhHLyeu2RQJIT3V87fxfYRQ+f
1G64iz6jGqMDezHFs3efXZ4+UluZp5B+SWulbnMUTIgi8deaH6j5hBw2Tg4wfxLjMVczIXgg4ovw
FiHmCPcaPa2VUkm6Ig1FNHAputgyYvO7GBclsUfjusZMlwTbuY7MZmgMzP6icm+pz0BxB0BdpT1e
/0ZvbUL00Y9i8RkG1dKyx4OqHaAuFct86DzfgxjvQdiu8OipRMRYbff3uBoAXGP984nIEI82uNWt
F5jnUfO8KDMQmP99LuvvlEU5gEDYJRmhxZyHGk9shZxkBl2CZhWQsytKnq1HoEpteZ5ejtrLHFGO
m6h1FjGrhBQwph6nnSwLTTzSTJ435UjrsfI7i9EuCxaJvKhr3SZHIcCK11ZYMg1ES+IemV0b8DSk
Ll/+9BsSb3NVMjaels2AIMdAUdAwqm/jkzvozzR/klj+BaMcARmxsnLSURT5vqBO4EiAfxHoEMVa
V4U4yb7r6tUEoVUTM32CXzult0Boqx5EXXObxw42oGcZ41O4BmeFOAf6+G1xaMp09A+eby6c7+Dc
0KbfZerXcR5ClinfqOgF06zHkjdWyJUAp2xC+Ihtle9UjbFk19zV2dKn8f0bGqZ1Mn6Odpsv3b+K
yk85ZBGzwR6oUo0Q/tFNsJEVw5WYfG8mHz4Y196KcLJeeVF4cUQk+bJEqyMLGguuBRb5w/m7tUYl
vIQpX1vfIMqlNY5HsBQU2X2Syv6ZbAyGBMpG46k0RZZarEmcusSz1uG89X64GceJ25YtMF+9FRkU
DSY8hsyg0V59vLw5xfZPPYsBvzAzIWl+OM6iC7T6v51oRHZcz7WP0tkTaMEspvJLX7vBjDI5SGx7
t7c1KiR5igUdSrRuw/o84Rc9S5jRO/TdWsZefqcb4RoFdJIe5JZuBDQjplIBVYJy3Gz8m9I5WSEh
M+RfsfHUtdByfmpA+9lTfvFro9/uyLsm8sNmWhjacjhSIJh3Gf4m4BENBn/jqAv7FLU/98nTAIO5
l5iQpQkm/b8WOeiW1pQLd6Gqx5Lk9sg7gY5EmSXRA2Ydd3ur58MiOohLz6+sjWLcB0bkuWlIi1vm
OsuaTleTRHEvkvq+pHsCypuVyKRyXzIr/17sglEBb/t8BgJs08e++VDUUxxr+p8NFNsVuVkfa5eb
tbFBbB0ZwfIkQ69o2peOLG7a4ZQDbM8zzPgP+/SNQippTOez08gpTqANjFLDzCHYxLm9Z5cNhJTc
4PQFO1C/XAU6/Dn0BuIxPXDR+MImtVXEnACeBmhDyMJ+z5npcpDajX7mAOgiigjTXwuHwVVPXrGl
7J2y4rkri/BbH0GyDk4jD+6KyCQAGhqnxAYeLgNzTxEXdu/T2jrSH5pASfoHDtkc2kHEYOFjS5UG
myYGugaJ9bg4mWfNKCT1KxxAFFvgld4ltJctqyoZSFuHNV6fXUEO24HN9QdfhQ3NOD6fbm8Ju4oF
Du69u1MEC8xfzt6x3gDX2EmwqpL8/k2VqmNu6DyC+gf/N2IWln07MF1lSnhMYLHYaCUeZu3IxLVI
zhzW3zx2LBbTyVqQKXT8IZr2WTUPVVD7GshPL91O2ZSQGNm8jArI4R4AwlbGJ7SDtCMiBdvXzlSz
Rbgk1x2lcPhoKMthVPGVV2H0poWCQF9qwLvCUSbYWgdIChV8GxiI1quUWz9JJ9ETnyBM9jCjl34M
Y3uLMUtMsJQLeY39eAMs2cm4BYtWKMapmvaWetNHg0zCkd2vYNRzAqXSi99BrfPJVSqrMy1da4h7
+FTRGr3k2K/uDEnqoGwTo2NJ7+pdDVH4wxSPVlojUT7OWih+b40a87GTzfUm6nKNp9jzMuCuAQAo
0HNG7H0LzpW0wn2on+GvJ3/vluIR5ccst9mr+oFevebkavoOLspDEbv10I1cFEYBpbXCUms+QK9M
F/8qSjnXcLKdY/0U1qsPuwcXatt6YlcJWT3c+ByCxhWqvn9z244pXjEspZqp3BRWpXKHGZ5u4MAa
ElNsqw7aFG6Twd0rcG8k0lbmNcrZN3yCpFjiaUHki7Llpw+dm5poIqMyjxlYO4817ZvsYhzv2Of2
ufIqE92EeCU++xnAZpN4LeiNPDpP3AmhrKSd3Tj+0AtA38WuIfRCRhtM0Fn2QGq2D6c0iEhlA3mw
2Z8GUZjBBxtoM8bjS9UHQeb18AQDnhmwwTFWc0tteVvxz5/rXmRsm5yoISM2vdCAA0oaNj0zZtHz
qOqFvoo7wzvYyAXjyHRR8oZF8+kxG0LmaZXAYWrSFuRh+2hCLqpEeFmgTWFUjxW+xfnfDIbAUF2F
Iu+XtLRsEVcXb82nU+jTkBKAMlCZ31FVpO9AbwuEQLWpe3S9ThfHxCynBejfzRcRZnP0NNOeWNfS
hws3cge1v0i3zQLI2XJgwIfVAxpjVfZmjNSB2VSBhJ0Oruy4nuK6w/dpT3G2lO5tpG3jBNbUyMgl
8yMyeLwwsQUibfdUIonZxzB80z/OqJP2WM9KNYoq+/NaeXDOo9ofh2Y6AslDybj/i6G3sLPjTJrP
ttl2A0+NJ8/6Xso6GW8LXFJTB/r1UdMtEIIVavQ4JS948FNAnuaWxAlegMaKkzWpgVcU0mmD5q0E
GwcFibft7wOkOekwqJB1N2Bjsh+88zdlgdIVkyyDSC+zvwGAouQfEa7GD125Fr7ba5lFgGsqb46W
0gRAE1RgvWOlO8Qu/Iogyanpba0i+5RWp3kUUHGRYU5L5Na/WzmEmR+E/9atBt897XrDA0ux8534
vTeIbnb3YZ+tswDb7BrlhoILg/G1W/ef6S9oRf88mqJuA6P+IbkKjpLtRyZZ4goaCgY/IshEJpqV
iPjwPhCuqtzf5Wv+c/5wBOcDKtwHbudTFzmcyTmiDbaafehtPxliljM0SrzyIJuk0ES5FGtz52Fw
n4h/mXBERAelDIixEiT11TQ9oSLi6Qwccf787VGilXXaCo52VVrT/NRDJ+MgY++xFlt+P27W1IBo
3f7ScNr9kBhUT1q1ULkS0rUkrYwH+1IqhEqujrPb9sPDN6MxD5fIJNG0pPjMzQqaovc459pvlaxQ
ffUvnBTPolR2i+7qPedjNJKhbG59GzOqIUIGLlM+Oi6zNB+ziXcYBvMM0CCCYKbawN0c/4BB9iUE
uOhGE+klmi/uq754Ougt7batfOcDX/O5UC56tO4jaTAJFScNpe7mM28//MbCpk7y2evjoGXjlIBo
y25hspBwFfOasplC6UQa1LpOt5jHxncBS4jZasKRAvPc/KrnHj+EukVmSaEsbcBso+iDqV4kjyh4
36QAJraORPr6CzcVRhp91W9eG2D50YWftciEk7AS1ijcaxVq6uedYslno5NRPS2CiSGjOaiXlllr
0a2tkKAcg7WTNL+fpr287kNbEcT7YRXlsxtGRejQU7sX+t2KSqzetqp7xENydB6hP89TtAiTxPpC
zdIveZ5tDT6bO43yg8wbVm0YhdTCLPuMD+5K0ppXQpHZYgslvIWu86KKYAng/dO/Y5mZK8+c8iMH
CJd9DWxWD+1jgbjtOz3vrLeAPibQehTsG1JDfO93whpJrfuwibcfG3Uyo7LBM0r3FdGYfgMyxfdA
AAHw1yembyLgmVnWhiHl/oYbhnf0zZboQIjW6UaHbz42hKMlORmqTSADUpEAPkHseDG5OE+t+aMw
tbVvZDvJYBk48wG6iCt+8XcUKLHWkW3pLZSAO5MzurYSgi+qQSo65G5+jpXBUI138q9wSGspho43
Fg4pS7NBOgg/a5TkQz2mrsAAi2AlDBMg942AvKf2Q67sH36PdSU2+EsUHXsk6Af1hOgAFuNOVLX7
VOchjT/BdQ9jpHcB44Th46lGjrupdzpFWZzTP1vqTZyTpDAylLj7kXnG4i5UDcXPn15EQ+Zv+Wyu
awmXnz9KINjyzBU7x75UDKm0iP8MT8apf8t8YQdW6lYcYrcntb8t6sokKVyebDehJOLsiuwwxb/i
o+vpyTRpWjr72JiTrhHHfDGgu3zw+/Fps8CsUze4oq5s1QX5SroDcJq3bQySVmzKa8ZDTKMlxPxX
bqotPuqwDFp+BSovOQQfAu3w/JOWQSha5WMg7iNepg0GlP6guzUHXNq/z9CQVwBGQGa1B0sLUAYU
S9pvxlbex+IffnY9ps1Bn5Mz1XdV75+oGTwFBqU5S5pnjV5TmiXWwvNomBYd9Z9B2aI9uFTIp4AG
OroeUqTSRzQWQfrmiRAXtLaZCz2b08fYMjkOMZqhHOVnGxj4iHJph07svCiyhRaOXMWz7F/o3OKO
3I1vZKEMV7cwgp2zHxu0rDrAc8gJKhs7uxEtTadLn28EzNvH/RUHGqhsiAFe1UMaGVDxXkNTB6jy
bJRAEtKY5Owdc1K7D3ieBycIkFhIJYj8ur9lZ4xzK7KojguGVDkbQlKe9DZTA3jBv+6flSAPasDj
T7lMIpqhN+PIG+IJrPR16Cc4ifUnQNaMR1qa3tiObPjGO2ycBbsDvVrEsPit1v9vxi1qCo72rd++
NdoCdxna67vbulbafJbEagmyn8Sf7nDn59J4YwVaRIaUNM8FUXTIwClUX25GM7kYAKA4BS4utpTI
vX0+foYNj2JKwhq1RoLpoFDYRo5HFK5mFgpiccWUMH//Ik9lvBV55rcjDd15Ytxak2+jty30+X/o
uIMGY++r68oJm5NBl31mCZLMelaaqPt4i0MAHpaEiaiZ8xaBzHgo1Dlnz1Xptw7locJXEUlay0ni
mFu7te4X44JwgILLsgFivLolO+Ma/fuPN91fZhtiRzeELl2VmGHevCpcqTXafwFvuTSMPSAdv6Z7
boOLu7EgMvLrwReY3TX+94IiXjmAlOxMhYt9qtw6/nyb118LPMt/CvN3rlfzHijKpNwK3/G9SAD7
HUjQ11l26ABas7jwfntjER73aq7yf1nM+2+aw/Z8yQW7k5HCNTNjHpIbrQRwpAlWN4V4E5eeC4GK
IqiHeeBALc7tUEnd3jZw5x7QHBsd3YANY4j8Z7+9kaqyIaOew/VPCupaqC+kzLvZw1KB74L6+KlI
nnhy3ieRxkLSrzW6cguCIZLiMHXOnxn+E3sIY3B0cSCThp98lvse+erHVSNXH01ekR+J2rzLGj5p
hPA8aGOTH8T9qLy+Z3cjwuo6N3gdZHlHXGI4S5VGbTLmU5wTAPlhxGHo5tn8ka3JQEQbnzfIOySZ
aE2oGG1xipkT4pko95W3bHjuhYnboUA42z3a5RPfySUdCGuKIm/ewF8UcQ3mSYsBVQ5YNVrckHc9
wiGYo1dQR2XGiMXipKqhzpfBofCx0xaBF/YJll72lDf7JvOrDYnP/jLpKbi/MDSQ+IK16EdFOLqm
Dfhqpw2N/D1fz6WdXzMmEBDkUp/nm8f8GRLHzebc9KyfoMK3v5YlbV4NHOvClZIAn3tpFJP6rSBt
w0ZTaeoZiAxOxnDn14TL3ay/LjpRi3kZPBBC02w6nbjS3/+dvc89KXRJte4tM21hEMAvfboBVK3E
6XuKiF/HjFQT2LUzO+TjDIY5gVe8AS9JFkPcbfZBzPUI4uQFJy9ukB2HCuFCf2CumbYvs/Gxh3NB
EM4k35UzPMvHbhoZAs8bGn7p9qp6EmGBo7FgvpEP8bqdSyfHm7I7DsMvwg+rJyVrCel89rIaLiGZ
gI91fdMdejVs6mqt8ykV63TLeA5OcIL41GkFYYS1v2cBJRSw/zMDR97cAVQJF8lyJ26FaQ2YKkWP
oO2/ZnnecKZHx/MEQOL4nRVRUx9Fw/ma40sbWZx+yfhyi3q3XTK8D2POjPlWzP9LlVc6xEk7heb/
HVg89H5UeoYa3w1Bzk9ec0ILgW1HnmODKy/egtTLBf9/5J5UVxryrpWil/nhYIu6ZBFdBfnK0kAw
Aq3IyVDCG5O0jQrQ1Se4hSesZjdWaj3P0ByVwB77mEyr9IXYwD2F997YTOfOxuWXvfL+qa1ye4Sr
f+jKVUp4gv90ldG+LXcQoFnuuxbxOM19YgUThBzbHPc6x9uXXtnS6gkhnqZit+WRC9cTAtjh/hhJ
6UHla/ShWqxpVciZ5I0scirfjWfgG/uhVtseXrYiy8dUI3vZrZzpwuiha/1l9+QSg62lZRlHeH0e
xNd900PxFEsETyvFqtebmnYPiQm7KJAvZA41i1TPrq4HpCqJeAn5+j2LN2C64LWpJAJ8Dzx0LXb3
lqPS627ezToT1WpC0wv1wGBVXzqBYReKd2mquVvmIrKtAfkZECLRtUpn2uwMOsvoxOHQpkS3QLRb
d+wtcKtvzbwsvti6FZro1Y3bwjkqs2K++F5V8lZrHlAwnd6wUFwLUgPIXauLp58sTBV3OMUZoFM7
kGI8Gs/8qtF9G1n1DHQxzjzUs+NtUcly+4bWQj3Uogi1iHQUgIjxq9JXii5Y+TnDDdwqb3QxH0yZ
oyL5UjZCgRh0AhKZ6/yi5gLow42Mr5ryRjmkwQufNIpc8gvKsGALnBTqe2w3QBFcLPgfCbCDqEgs
5nj3vTbConj59jLkRRQr4DUWpUf3xkquqffBYTGUw7eLg2rEubBoSaXMos5+/2KwDxeNLopAqkuv
oy5Fft5EgbOjwzRveONyz+Jf7PNsg3xh59w1VWamu6ksWj3UNhNR6DWmh6Yn4vN4CWfEk8HP5ooH
ueXEjikX5Bn/oo7eSz83J1XmmATei8qRd8yLF22oJTYjOO+x9SMu6qKu+iZLoOsAyapoPXQu1ceo
LSnFirzNJBxp8IMpbbGfmNEHZ5xgo+908bhfCnPcWReAazYho3HE74DIdlkf4L0hLgAQ6fJIGflR
MgH7PzV6OGaIfiMawswQqfZdQgOT1zFPCQgtyGCRwi9afDQjOmS62grzmefDQJt8JrBK8iJGnwBA
ZKOC8qEgLW95p7y7ocRgZZfckwoB3UW15aYhO0KTjm0e+da591UdIaZUSd31BGauocFqtVBzpYuU
DW01o6wgL0SweE5p4fX+Pdtospzx1Agpl8xzSklg02MZSxSbZOLrV7GDULQYcIeyqmdfkE0xqMki
k908+Sps+Z4FKuNIFwi4pOQgTDMHv7eSE40OtBsYQ1/95pqzvXBtw8fhdf8hPZB2zbnatX+eR8Ns
eWgWtFBdovaaDZ03mN3vvzW9Jeso1TCagZ1cSTIweMWdXoWEQaSJSHYUgXGW6yylqJHcUhppzq7m
B6JQx8VIL/gohXTDcWAWdC7wLV8gUyX2RbP3tAojZXkAF7o+wSRB+1wodAUaw2ug+AEWJVLsHmw3
Z50cmQlgDJZx3wf4UcnslFccjauX6GygZkcAWVvvbMAd0pqCEZ8Dz2WErk0SFmNXsQNfuF2Sw3ra
uFRe4X1Db97S//pag7e+ltmkaxvCulSckv8W7A9NzgVvIu0g+E1Lt6/b2xtb1YMUvLTje2KyoYfp
n/3nIhqoPAkta1eFYCs1ocZJHrSEURI1JGX1OPddUJxQAsiN7QzCTnAhXd2nJBBAhTu61sYt5yWL
48ke6a+WCbKd9aHEFi6sTapn+ZZINeCp2rCpkHkLd3NqAQ78qZpgk8yV2vawcmOReYnVaCXUxNd5
XtwFLoFnNRogiSokYfhJxhQnBTpDN/Ct5lleWDIwsvZJmkmrAA2W/T4N/UTZmkiFq7uBcjdWuf8L
KZpaDcaR+IyzeJA+W9SaMZYI5RCx8EYxvbKraCjydDMOImva30QYLnarFFV9LDhg6Goqiwb8alRi
IgNEN2Y2PjWYv0mgqdLpD4qW1IpKCUT4gatSVVtIftFi3na0IG3hjxEvpafaon/dzxYoSHFxRiH1
SNdnjMZO362oGucr4a05teJ/ZrKY9aF5RjTASLeqakApkXSJmEjuw/M0S4FwEOmHAIl+yjmpvx9m
YrITlHiAqBR//01w0Wvm/D+fDXt9G1abvml5ZlmZoJBlwSOopOT+T8z5XDY/c4j2rHgptUjz3I4i
yZXhE7uhIi95WDFQ/PR9R9v1jBR+U9yfDvpoV17El6SJInTzygUWnIdWZ79vgB+qO0Mbmln0omxO
bQWkiFN0K590Bci14e38cxkJrvZgP8DabVt0vulDcCUhys1ggZUt4e6my+9kXsp/XAO/IJsm73oF
TbBEUYVoF2vZ1Pa3ETtecR9AlMiqV+ATG2BliQ2gw3h/i8O0bwqXqhEced0Avy2+LK6+aai/bxnC
VUORuyv7SR5Kn89gZ+VTx97p6xN30zV6f0AoqlGiF4AedrQay4Yl8Yh+WH420id6v2/Wpi/Ixppe
A90ghDBZo+DHp8llFAHvzKCOMGYLsmZaTQrsaXuIOLG1jfph80FYg9eJz7rRlrGov+0tsAlQ67Qy
pBiFDQ7Cby8tkFcJFdrghGsFXUwPyuP3GJHnNlrZs1ZMOkWsRmirTT3eN5Yg+hNqx/atCjs/Kj69
N3PXJzdMVtteSLUjMXffQGS+PoP54/lD2cLEBSJ+oaqUj8pXfI1OaObOhwy8r5oVxh70pa4RU2qR
qV0a8hDngHbB5V0eMn0/hM7ln3S+Rsp6gAkQLS14gYycP6IJno31Yv+yE+RUBL4m7lNkcKMvsFfE
Q15/fW7FWu+tAOsxlQBnoOz13H10g0htrBe5HQi5+YkVGOzq3Fq3e0qiwZjvryic4W2YlCmHGq9J
ffF/jeS9XPHG4LXS1O3jV/Rmg8VqgvObwfm5gKO1o7bEAgIrOInRm+GTMOQK3QRVP4TP5Ddzj6lp
OjgqPvwlVHs7ZiyvlNsar1+V/6aCd1AtBCF0WAM01DEK9e5b1QpOJqRCdtQ0NCq8TMFc8VcQkj2m
G1LfOl43971i6/bpT8rqWtE+rutIAiPpuLmCp9jyaNW6czbqFAiaP45ABvpnyK+bo0JqwcU9kd2G
th4fdgq0+9qixi9bxWsNZVk9d3AQzS1LBWVL8JRK+ud3jCEnVe3tmy2JkxoMKYVqcolfbrxHh6eE
KRl93Z84PpMAUpjh4ktHM3iOYEkbIPAPvzoqmsYT2jaVVzrtWjPLGi0dntj2cSJ1852iaYQa2aGc
5qU0FvLdzHWYENAZWALYV9rNIvLWyWkjGNjzzRlrjbBCk/dAQYiQpM94HzEqyOH8v89JNOlX/Agv
GnovMRTaRBYkjjwuKShQRAUyFCHAM43/II8o/qlTK7CMrKO1UfxFwFpPM8OvgFGfl+w/uIM68XlV
gw6xUyfOmJ5BY7t7bvzZ5xPllG1vC13I/MGmuZ1xdq1NRmviWVDovho3mpbWK6CcZQ8CFUrSDlwk
7SCaymX+A72531HSssvsOhqkVbtBaFMJkOrsR86igxj6xF4SrMHLZ/NfToED1RPEeVB8MijBl+y3
gFTbH8SBlJkNTy7IJW+dZr2a2K73XnNIBfwdOSXdiToewAvp/rNYCV/vj8ICHSDDI+45LBwrHHzw
aUhRj8mksI6bGxEMwrfzYGbCWWgq2Xp9A+R6nwzUbHR6wBI1cZqthPdmsb4Z1WVx8lOFLBIt80a7
y4FwlUR4gFD4N7Zmuq8RAW064nM7n1UKMo2bnF1oasaHgleJDKlpodjCOMfZi71UA3X19NXeSRaH
mUgVWr2MoU7X0UdOWERrT9hEAixmBQ4golpt9vjShS2cJc3yM83JZsykkpIpGqz4ki42G91tzJ4U
XDhP9/8H06bhSr43xnsre4jwQXgmJiSFPHJqPX3itGIgScWp/qKyikizCHfsRM9zVTzfHix2nfyr
J6swWN0DokXn7I7NQznR/h6A6DV6IkCB06iqL0LrrAl7a36Kz9FWN3tWVqbasoqj8BVpFthvu0eg
Mz/4RSBRJMl6aTjRv0c/7cy42tzC35hI4aczD1mWf6kbn288c+zruxuGCooDu6hZ/pXKANYUiNxp
bqWPz9RsyCKPdq9SIlj42kRp83EpwnUsfj2Pl1l99VGhJeDxWnEJjknVKGPuGDriSdLmEGmHfJot
h92i1eBQcxoEDhSVKbG8C5zygapCy6d9QvoI+WWQN8pHF4Y5XUp1r/mza3VjxUODw/QOAiooljNM
3Dc0Vv6bWFfxyWCrOZbaug981qZudwlSvF2/YdQFGbmMReDWqDZLk/T27TMQYdyLvK2loC7Vbj5/
91V8NqMhVoz8xF/fE4AEUe/AFpFxS0Kh0/5dH4cmOa87GZaLQrZCnQ5mzdcV8+rMx6FGyuOMD/MO
wK/Ch6U3LNbW6T2nZESpAbTQlmr4GOCvQ4uLbxSl6EKyzLRAbKWfNTZ64IPwFWBFfyISzI8Ul9Dd
aQAOQVfYVcAULQnGW5LQPqW0VgeUVT4SttlmNiJ2Ho6f9RT1Efrg8Tb0YKEPqgT6y4FT2vIuKvBO
empE59qw/IrLj5P2R7qRpALVBnd7uT75mGkmwl4HvJIqyWrr0XjwCEL830otnT1Uow0L8K6dCqWl
fJPO16VYtEP31yTc3iljbQ+oSbEQjaRFU6CgP52q+ZqsDo0XMwDHQ0H1gjsxyswCkF6WIYXcgjsq
dh0l3ou/acTOXtG25lYpPvoxJfMHpMB3fAq+/ZSziAsWoUKUQG63kgMT+TEXEetpYsvDg6NIsN/R
GGkhIxi1JDIqZxy+3sSYp7hsYJE9nBiUiaUhdCkmhGrNdwKy/0HNgrvMw9DlGSm0hq/g2HPEeJlU
rzcenCIyJdzSSmHkR54hKjgxrbE4M+7121fVFhJJWNOlMjUnvpuip5LMwvvrTRBsawqg6/j9qbZ/
Y1r/DcT3+FM5Wge0WKe7vQFo92YZgtGMSBT+jGrqBmuuCu2b7nmPvLBaKR1vjEhz9uUhxA4epD+2
FICOJhMF1dtF5O7b37Vino7+VhsPK5Q6qysx1+C2I7wM9X6xGBTKkoAZ+Ly9RHaHB8DwpX6X7lFZ
9ccjM4JHoY1eDcBxMeMlp5mYt0Nk/c/ifSebQKaRoNmB9tbhRTLktrKih2IxFobVAq27q/BOWj4k
0Mw2Lw+LeAi9qptpKy2D+QesQ4QqnrJX7gLfuXHDbH4loHrLfwCRXk1A5gKaJBUKLr1fumMl9Xr7
Pw1HSD/uUfuXRL2OaH1QeN+iUxX7bkvWqd22xeE9WMgBMI1m/H6rGYFbvadTFrGlBv/q48c5Q4rX
T8l3j3EU88+VkzvF4FLvncP5xnffKKa9MvXOnb7OcuZwJGCm+YJBm9D/KN3/0Q+51zZe3Z3J6ixa
+2nUbz0n5x3JFvV/B0W8Qb78t+rZzNbKGonTMocjDwjZ5l5NVo/rJsg1DT7jgMXv0rxhFiyBN1T6
klTzr3P98lw0gUwVWZL96liuAd9CuNQ+SUiSBkYma4dy5ZdNmq20RctynsHOl0lRjeQOyOEs6yI7
8SLAOaielUKpIOMQind5pxFGUM7PKYauwuRLTkgGjfqufAbZ22sQU4Q0U1/FhTal5+APkKk6Hb44
A90ASFzu9jSobYEjB0nSqAj0talALmRR6cP57ub5hM3b6h+A2vb6BQrmIr9RfoEnqrQpHgohrKQe
rYtCmtdUV5cfxRMIfOb4fJxyz7uUiZF4D2OaEKHyMoEH41FQ/tFgHJ9wtbEEzxLyCEfHa+pIq7L0
47carOSWu/hF9BZaM+MCvCtjCpw02sb8uOktBomYLXYxic8EyZ+zmAZkSSXqAw1xp/nvG4NXGtYp
ZylaZB/niJzLxDGTRwFQLCeWK2oceGeitB+D9FNBLioKZojOgkZ0yg/x5wvXnoeBJU48nVV4dSHp
Z+AMEX2MZSbzRehcJf5BNSwp2YsDREK94x4z9XhsvrmH3hMOwXrMJE9g+aJpUK2R+0D6+AUqhNlS
g4wnkkf4YizGJC8EUJPxov4bCtP8UXtTZsJS2yMlMrX6SeghcmPHM+nop7Ga5k5eSNeI1TXHWBDX
dNlx55BQ/RGI9062lGoXZDJWYXqpkPLGZ3DECmeJecpFxCdfmryGoNqpo3YsrB+omXUIJrttVk8Y
L5jQp2FKZQI4xKk1woWWatVck3jG5GUi8WPdxLolOAL79Uu/tWny9cvOzQxmssluOI+P1KZed1Sy
fWwXadSs6gxj1TlhkAU02lGAXQOgHujxMTrt7PEUbBoKNMEhKpcYg9jhetd0twZ+F9Ec5p2OFsfR
1Au06GKZknRSJi5edstj3w/f57HD+Gk8/HstiZWHEq3380rjic5NisVF9AUybnauY464eAXav9gP
B7fae2mtWcCgmF9PQHOzpLUtUHJpz98DBoPMzectAD+RNQvwPa2StTwxUetVrTzmwcilEE2ULTLX
LeixW8tj2OAA+kvu16ff3WJnBHxVuHR4/4gbt9xi4PelYmHvzClN4q6IRBLubFEOadU9CHuQ6BkB
Rf8QvywHxsZ22pvHychZlzWCH6s7L/7wK1y6wPgqfraAJQG1oaWLdNJksD16mgQnsw7Q1w25h9Kl
gpBk57QW1ZDVoQU0nHMfegRdcIWbJNstXPB0Nh86dhwskRqThfgr1fGjGnzc/TinC/KAtpvFaSkG
RK/DYiUDUhlpE5gCpZ4hfN915JAfBt8XpDeiQIRceGjp+iqpc9UCScV4cQgtCe4YCQ+2bk+nANdC
8CBATfgkTt3IEz19+DVOdp7CqLtEbnyCnT4iLjIXC5McS036U6owV/RUlsB39OOrYFrC3ggd7vbH
S8dsBIARINxQQqNvP2xQf6EB/hYiJkifOA8szp+78QAMg47RHOThFJBvMXlCDN9IJzi5vj4ie9TC
RfLlx+Ib3Y4BIOgVK7qI1EKZkkgz9L+k+EgGONPLhmEAgL7t3O9k1GSpSH7sYw7hfGMJ9q5SHSE3
ncrDC5OitCQ5GnBBjv3xGKqi7uU7I/Uo4iEaxmKIVTkfTukXl570cDVJhwTsckttO0Nihn3lWf3a
kiUpXMLiOK1KKd/zxILuhQ3ZX72otuf7LQlTi9XOM1prXVNQMJdTD05R+/yCGtEmA6DTKuOuK2yV
Fd0s1wlPqn+NvGsJ2HWDTPxfhC5GGGmTqWyOe6NpHkDl1pqDve+H2r3Z2CzCI9tehJ8iRvwoYX/r
obeqZuolVFQi9N8aBUDymOab2OoZrRvnJ+F9Mak0ID5vrOSyxlc7GEVoAqqvCoe3N9Ah2k0TcUi0
9RP7ugQ+PN15ZCS+2ABj1vVdTGkFvjXB6upaPVs5XjO9oy2mrjBS9tka3vL/+XCG01PWzxbo7l5h
DTi4Agr9jPpNnuJbI5FWRnqt063aNx9f4vkfvVfl+2vr/fJNTcOGpcCJaPGMV/zQ4dpzoMvhROfw
O+CrZIFReShFfnOh1EQUKVdonfaE5xCpZb1+l1CLzPKAjmyGbMiQqpOxpmz8g7IdJx8bF7R2PBAr
vK0O8Cmx2tLcw4ACVuMdgMBH2PddsrhghHazyeOP//soFs7lJ2PzwZJ9RHQnSAIHd3CCXPgBDsxV
fSVHM4U+Hi5yTKF0HmsO3hdwiUU6UouazDV347zMIMOpV1n0m7g5z94jcVIEOdUQNWjtjnQBkd5L
RKlfmGZW0NZGA0I/2H6IIKahwASNIxhSKbl6gH8bW0vz0TwtmTx0jYio3T8R4jT9SJuozD2eaSgg
kJtfg4gTvr1WHoW/oSoClZ3VpYWMN8gLrLoHzkQQLnUoidPslJaRIPxA95dj6XEBvOZ65Jyca6GA
iiw268GBJF1MzbgZHJ3bDgXtPLNczzmpYK5H635AeiOciqfRtBiHtng39QOnPuLj5ClNKh+I1kl4
+dtXNXF34bSkbGncNsarUhNyZ+pLebVvja+vXTk2NkWtTU40Pjwbn+HU9PMxlo+c4YzLpcmZNxED
is8usktNe6x0xYhiUtIsCvVA5lFN9fzJNU/l5BhDAzamVQf8fIuaHno8poTUwQuV42qxhXuaSXvi
hK0IK8YnJpnTuwL/2uc/xqk1x3iTfN0qvxmKF2zydfeOWxcVWEhFF2lj5YML7IkDe6T6lgGRvVFZ
0N2t0DFCBT/qnDf9MKKpNF/EpUc3umAXvSaIcfRrCMFbWg/nmGEk7qMtJ3sr/6exMp+H/XDzIU93
88m6LS4CUV3ByCCLqIF3S1sgswFmmInJl5t5pGPJGWMtiWeCukgHJkkPnRKlzW55ieQ9KtD/WX7W
FqUE53QTzhpZVVf+iICZap+/jiSjaJb+G9qiLRoOntd9KFu8kndtODHMhmVP+w8IKIYNRtEz7T8K
LKPHWc5sU856B6SX7GdBjHluZ0jlSnXpQH3ehTom7vDy3xCbI39nw3O6zw13DGPMMcG1uMqxclUC
40G5Vn+Kw6giDfoAhwVY5kmThxT3ICMFL39yz2F60YDyYa7A1nGL/7TJ3KQ8M2p0+a2sXgFASWGV
rNO8+bx1QEBvH1UBW/xwHjPCf+QKtqtSAzWpCC+6t7yzWCqskSIF1WnwjiFCtqNWrFad3Hk1ICZU
zi1Ni6zQEuAOSmwdsa35A5fqGkJKyweMjSfp3crZ6zabZC7HAtG+ijxqtffon7THC4Qr3sTPgfxl
xg9Fz5oLiOp3/YjE05ITkFrteuuKkNEGdrWVJ6aGCuE+QIPwdYKIS33a43mXjsNAN0poZvb75icO
878K+LgBqUwWaEy+r+e5iUpeO2Fd5UzJMveZsZGLEsPpj02XyQyhbq1sYODPZGIOWjhyHZhJ6vNA
ugwnOPmxrHd8y3i6VKXzVWQ0SWF+wEvrpK+lY1gSSz+xFEFX443zexHvQt9K8GZR9i07EtzDbZvY
vAPONf+g7NHko32r/QDqOokHlIESfXpYxqJ+aY7YpNadDiVHjvXFw3Hs1vJfwrdmK1Z2fTwQI74A
5JGl/ZdUjHomPfmbRIKcBTQUNwOgs3kpgCBXGnq/MibE+VoQUmex2aw8I7Xx/YgD8sabebboXyYu
gtSKzsrNDZ+y7LTZALJdIuI7mWtz558/2UFT2JLtr1tznRdlMrSGdjf1WO/FmZHb3ZpnMEgpZQFI
ml3ROTZ2izURPuvRjUym38QghiFHXY7kWcaA4ZJgTaiaWdbmQ/q4tAs2XpKXJ5xm/4UdwowyQ1Fx
usefB2NH6Y20wIbX3L6Px6tZowpDF5445CJ2Ud6t+DI7+fdzPs8vHXCjC5jRzGgNdeclasH+CzBH
E6di8sWxTmRi6AY1PvLXZtAmQ5wY0CaCW7YWxIqllakPeB/WavQE2OK40WItPRGivts7Evt50+iC
b7d1f+t0hAILoXYlH/npiwxNYCko5j6twJympOjhVwUVWKjzwHNVEVPMdJ3XAmLHCVcue9iRG35t
KHKY/y8SepD3ZJWtpIMBWKUpgZc5OSRPYPrWgPBNeaZ+By+H93ZZaiW9SqPb1TNdSYtWYPxbIwoQ
j+VM6+JnD7mVXhgzWEUkQZaF+A7L5zrcOVpH1Vk4uwpm2B1cpVt+b3T/iEP04gFmEi2fQBnh/9w9
w7iWAOH4YHgBG4x6QnQGlEjXJhRla34CxzxLcxhQWrqOWXlwSffyT3kwrRCiKJlx/HVe4V2TPMkR
LnqPXs1pVcQnWXlb3iJxu40s1ASgXM6qKV8ocxtmpcjp5Dn33PAe0KFaW/4ATWJwOx8rQzBwmhQg
zQJE28R7goApTlhn/choea4lOopeojS4eOxzv96qJCp2IN1Um92L4sEtBzEvYTFE+YYx/08zlZKq
RRVYaQl7afEm5FIhuLeAtmFQCCSK5Nt5B9eGtlJIk7viakscQWpVtUR78Z6qbkmUQ4/YEaWdS6vT
Omv9OUjLfW7Lad0ULl1Ef0n0gorVdEB7rED7A7Sug1YKyUqKlYf39kFNijsj7MW+8OwljsSHc7AW
DY8EV/O9PBJsOL2YToJ5U6/4eX80m/QH96/MRbg5bHr42N1OM8bbF0OkuFrUNwwetriM091x7mrj
CtH1Q4P6hNk3NkSd5g21Xr4DeCF0bEfL47XsI3B2Obcuo3DgR0yQRovCFT+NQLavhNZp/QC5Ku7x
wym2Mj8xjsRkxIGnERRcbuA1Rq01Mes4Ex0d6CU8nVJNvJ4ly6gSmWUQzuo8NK5b0FOhMpttJrLm
ssxZHaU+2wpT8komF4Lj4JHwjwcqyEJ7xu6WGalzHtY1AYOSI0Ode4SDk3PixHCRlYySW9DPlNzE
JyCIxYy5uE/pw6fATAcF3ChCYUO9b7tFcIH9gNwoQId8qZ62XgFz/YvVnsYx4vlIR4GnkEsOizAz
DL/U/1R7Wf0vOJY1A6fd/5cKuc8L9rO3MimrdPEUUedqg5vRz7493K0WWqbqzIGR2oLi9pVGITYV
L1tnSbOS22UkObrL+ytUNiyM72K5Zq/JH0Bkfiaj3f4Ro295KLTwTQ77BpCEXpOKrL+/Oq7812/4
xTFz9E1cJnrsykcXdvB5Zn5yH3+RkUdr2+BfNixFp+zkNRWsYR98+AzM0YFUHGIUTZ7CDWp1oqwO
4K/BzxHWKcAHs9oTMW9cviPvzXV+UV2gXRtsW5olkc/iDSrXoZYqtGRDTVkZMYWdA9gO4e7AD47W
ZONU7KsFHtgNmjnMof0bx70WqxRyTnttMh+qnTpNuziD7VoxwlTM8c32HX3BIMDmW0D25Crqqjo4
MHLIseRyYWWgWYogknpQPCsvhWqaC3lludPqbvFSw6DG01/bLkPzrvWBNt9eOSic5cV60m82WY8W
8uBoLADaaXdYQFl3J1AX54k5h4iGfDFpqGPXeJhgSdryaEmo6ZoV1FRUSdWqKzx8Cu8o1jt7roy9
Of0BTY8j2bLd9UKK4Kgk7fe2IHGwrk9wogaNo/f6GBKMc6VyEkCgOP3q7ey6ncvTsULd7MVrx+RC
lJZf7+PmEbqsOHc8VAm7MONc114JlX0LRe8iWxiUkOmR9Cm1bT4KIbGY7QJiVCUK0eP1bNdvfFZm
fGGyhr+4hpHXmZEwZKGHdYO2ZaKUoP6SsePn8jX1vfou54kwPph/RU4N22vOePw0NF40uSyC4gBu
/LYx4Z5ZUGcJkodB07I4EHfhk3yf8S2yYnd0dbjG7HFV4i9h/eJ9XURe7yk7GY086CZNFwz69wV1
aDgOkGgPbLRndH8DiESZokk2t40CjqH8+IjJTYPo2m7F7ys9VQdkEV68R44WZ++HQhIMhKNV9+/I
6ctCGWeFyCIowwWQdfgo1XaAVc7OOhZrQQg1X8ElNKOOvHyvsDpf/T4TN9+uKn40JcAg8Z5+pWlq
j8CcqLr1X0APcrmSXmByH30dv4o1MYdts+aBSgdkuQwTigwvdGkZRneP2wgjCbb82bltLHCs+emv
y9TIs0x7LK793sOhWmijSErA/sz1AOvobGoBsL73FL6FxNDkORk6nPFRtiLG3IDnZ32Bpa7nzPub
H06M2UGnEEyVQMk5E+R1A0lDim1sNPrE+YVCsp4GrZE8EF5VCICy790vFfVUNpf9nDqCkGt0aQtr
HU0u0ec/R47SwLYpIySmejUSYLjp3XHUGK0hb53NKSYzXMlp3RKLMVcFpeT3GsFp3PZrJv3I+GqV
fkVrC2MemnGI/S4q6SJ4VZ7DTj8gk0PK84SPGqoTWdzewCIIQZHnrcM8sv8/tZxuNXse+q94L3AK
YW+xjuo6jbQv4bk6twMc0wtK/HhXSlEGucOtXUtEsqYcoOAEQgjpD3cp94FFbRdIZGCHmyf7R6y3
muWptZvOP7Ter6LKGfkILkNZIGIL6p789K4DlNT+HH0dznaexRWeyzUoNMwzJwBs++u6riksNv0n
Sz1NIa8EMCMoy4b0cQ7VEjYsk4P8brVOC3FUkzNUH8i5jYNvkRz77N72dZOxZ8JKE1uTzdcngtse
g1Pf9O+knKjf2C1wQ0x4OKV74qPOlDSb+ZpjMYceeVy9LJim6RsYQfjbtnd1y8Vx15BhvpyKvt1+
wJiO+Eqx5XMHf5R1GXAaHtsW5EJsZ8mFAplKlaOMB+psPKH7Yu2qgQA2vCiW6Yfkm94MUdC3KBye
rTSmpwMy1wE+wjfuVMiLruQRofvhmm6qUkuaPxCJgV8/zj5EOpVMdez7c+18mwN33FGdKQkfFeCD
TZjZNcJ/EjYNdjl37oCj3WcWXhwXxGcLw80Ewi0qkvwGU4eqksfwLBVwhszzsscI1Z1z7OXjdmQ7
A+qTI+opHbGOvvexXi8l797TImsQUNt6l1h7VlK0TvhrQaBPHVlGSXrHYiIIcKYqP3tL/b9fLHKy
zMdGBo/3VdLqagA5jJEpeGGcNBxcF2CAuE9zBMuDgDhp/ruNYlNMVSJF51urCxJsmkLz+I4cf2zd
k5glh1a6zOnTxxYTp9/isG/e0Ux6u2RzFwd2P7vFToB3Ff4OwlnYUhLZL5AlturMVtdO90CjFlKX
/X+HGRB8d1N/NiwwtY3VWIaLJ1nTLPMlXee61M17mAYRBMHwsoynUh6iTlQ4Krilf5Kh4oTgP9W+
M/6qEvJzLPMn5vcSqXYVbyfm3fW9cgjZ6+Hf1iDVOCtAv5Q7UIMyFNk2SlplZd3Q2R9/Kg13+W2/
auZmFNe7dxA9242EIEpYDA+piOwIHDh3fFy+sjxh7GgIQ4DO8l/9H0ngSaxg0knYejspGePpa6CJ
m79cc25zCDqOD7WxyMBcDQi6SjKr42x3oDgd/biziQ7sH0WR5N8LlRqJpXmy5oqaV1QcI/Cli1mh
9zMtGTYB1T102/ZDoeV0hOf/UP3fYzhQavCk9IzHHF9wZzwB2OdPPdnjNIU/Qbt9kGRYBrfPFfuf
ZaJkbADIPXYP9XTzFaQtPDsPFzaIbqDmkB3tK7CV+jW9fJsALqa7PoZp3vFE50z99w7eyM2Ll3qy
ZnYYSCfCCaGyK80d//W+ILJfq5LaS7Wut0jDKTDUYd+NQM/V8lBFkEAJOFHe7Q7CK3lZjAccEUgT
mVYwtd5hz5TsMI8h7n8sLOX/cXe89RmOOjsXQmCtSEQwXjxcZGgdpK/MWddja96sSFJADwaBC17Q
Y1POodyTk9hCoF68/uYMDKq9FvitF5I+vmXvmpGKh6kdcvB80BCet6YXP/kzn54gptbB2X8xPHty
E3K3FHy7AzGOt+U+j02WEk2FLT42FxCkUWhQBm1BpzWqiqEBhNLzGL3oPCAOzbVpW0DNKIgRfTti
6+5bUmRNLe2E76wITuzsYWoILtvrkVV0eBgH/3kuXN4RtdWWqWRDyG5Z7NrU6QUQmxNAgtpToN2F
bE7k0ChyDRwsl1/Srohj9llIdzE6A5mlYaLp/dVuY+tzHZ3g1yWBZrcj2Mscpcw6nWpIqD7i9r19
0c95a9Ctv5NqnL4uoBzWTeW/517x8AHsp81GBC9EPA4u83hJEF3it0M81Bl2u18+BgSCRCEFMawR
hNUgjx3xfNjS2GRy66/8fTJD10BfzKa/aUSGodYsCPo2UNHUkvWHLoTHt1YkkKo6eK1Q+t7JC7pt
7UlePxJAGC7oD8Z8OYyqhbRix+PJpFEDBtW2rM76frRtUIgysBTigtaqK9KU/opJqCnbWPb6dHN1
s34HHPYiEoz9662a2TNXarm9GJ3PUjddPoKHgUSLdb/ynp/4Ld0AAm98cD038r/aubAY+6qMiGHw
CDtzqoehbZbQCPscKOM+VOgyHKXOcaxbDBCYe207cbJqw5Gy48PNmeX/SdK/bKcuMmdK0JK68wpI
nLvl9GUXs02I2uZQEae4HOl6Su+VA1gLgu4ODukoCn4d6VVuriHeDt0Sm+7bLowqTZilvQe3F0hj
Mlp4YXSYw2sOHdiW4X3AT3184NofMOaSPyTEcaRM722rrJF6w/tgPXN1TQjKgzAMsw6mRRBImhWQ
ksZPlB1cjtbBPkydznK5YDXQyXNxW9HGERSzBEgld3uf+BI7Y+ALSPAZi2etrCWnaNCSGkI+uhES
kyvP4CoSm0JcUrnvQIQsJqxRkOD6IRs7Cp28C2GkMqFuz6EYpH4h3T1xNl3kHuovMF24VFSyOAfw
+7WSyGA47YtqOru325Lt+5UXwYsdrulDpOM2w51Hrnl/dx70EDpNplGUJDvCasbUNUHS2cY4of/Q
Ndl6nZv9psRENFronn0pEQG55a9sg6LmdHZJGp+h8YtLzYdTxhMQR2OYSERowTJGCZPRd5I1FqY2
J1mY23e8kTkuJdGxuVkYM3iXBlVBcngNQEL97thowifF//8ovwiPeWv2MnVaqcM+bJjKPxUoPoD5
wwilnKx1b6SD2wfsQMionhYQgVXNalTCeHwoS9IZc9OsKtU3LkaSAZRwkuNoqKvVpoebygMkAtLA
JGrd0RGIA/qi1lEOvr41ddzdOOYMSIIig2dZOdRtVoxarObKO2Pixt2Z9UOaHb+eLmECCHYuTOa7
IZuN1G2qFjeefebo6mfKo02BFO+43wFZepISF3CY05WyLX1VSEUhFP9+c2D7SqB0sgAl8dP2sny6
uW/V5P6tovzDfhou9JzzIQ2i3Bnrtpxj0aRWnGImx5oU6ChQhcrXZyZQIPRRwXwvEAw7l46gxfV0
BwT+5yYNNRXVfOsJL/Snil4VFpKChkyiMrXW/oeTQS7g8/ghZjGy2N1yCiveYwLYq0ViIMhacF9l
0jPQfFz40xDZGzjMROE3dvX58sMYRWWDHOBqBBxGta0UqPbNt8MyeUiJXuM3TIZWouu516i0K/PC
hs9wRt/9HuPQxd8CbloGsUUdT/kUcAPtLpZmX3cmUGwFk87w/4CosaVO7K8QQh/ygfY6Ezd3bycM
LVFg/KWeZ4cU7uXBX/tt9fuR2m34Y8+8jvx3sBCC1LLFGWoYipoSLX0HiaSfIdj+uvW234Mg9n/p
XMoBee2asSP1TgALKHt2+jNinL9Mb+PElYRWcizZmdX/QViWjhbaWEZTQRPnfCz6krzrP4iUJQr7
vZnae7KF65OEkYbWnCtqEAYbHSVZptaRjdn0w0BKhxWvIORyoxacfvfi6spm62HATHFIgT4/EqNX
8hiClMAXT9HLqybsKPVm/7fc8QX2Xn3zLmpMCG2Q5Ncz+53LzPFtnwCtOqukdKQXvYrttNah9nnb
SAa8uYKpCsi78Piqjpw3C6PyMNwx1oM799NS9yTLdgNNXUuV0aYyr7tcUtxfXoNTunYDZuAdVjf+
h1HE8NTsOmA3Zdm1HLf+O4upoPHm/r5M8Ki8rgB6hdjM9kDAB4Myt27hgqk5RqyyKY4EssxRO4ru
sUjPX6Ts5WDx7wiAz/dth8v4q6laHrbt3No4uJAQSyiziBhfGXhh2KEt8kBaECj4MGWIQPaNKnXA
EwtKv/eqRuxJ+JWTNFsyV9KjxJrkOlAqqbVDpWShDzy8k9kKdbvVS4KW5a3EnXpIZ9zXJMp8nQVR
VgAEELL5YsB6z1fU3WN9bVMxDHqthA1SMvnaP8WRwksdDYwfJqmGssnY/D0gA+0GJHskwI6IeWda
zMmvDrFje5rQfFkkLPhe10sJf7OTTnlp/UIByZKEmYT1myahVZheToA4KXyBqfyPcmciX8uq64GL
13ywWWot/iI4HWdyQ67BQ4Y6vf/BjPBACtKxeHTyzgqJpuF3++yj1nTSU4VMB6BE0w5gha3ZEzo1
gJmQWA76/inWRpQGG44B9YbWbSUceI9XZ3/ryR2nTMcvO5221vKGSpdG4G1bFXOJ9Jwkz24INhh9
SfLlUJd1UgMWmH7hdcX96s4VDgEMsw20Me8u9oHwbmWPjo44BZnuFA5dH5zyz0mxItRxuoxd4epu
JIX/yf2wmqFf+UaoZitk3llytxcMk8VMMU3mGjDqgeJAEKCBPJTQQh6oxLEjuq4MUA9NlfkS/K4q
xQjq27UI/lElbYZFleBKXGMO5qJDK3W9tWGGvjwPiOgwM/nmniAOi2zZlrC0ucgzw5AYxB9y4BV/
2PAGVRQ4ugaOpLFZKJogEQarHq4zXuHBDyrnfKgCrTC/IC+4MBGYaCwQVepANsbp7VDFWhw55H6i
r5hq7P4Rb3Jtq778VVSSWb46dt8djiHub+Zh2MNIoue8eoHWwDlmxirCekPA/QX5Yotjip+nO15f
ye+Je1nPH0+iZjvZfXGS6Czf73F3wOtWIl3a0Inn2MHOHMeRxeSS5Q3tSvGVU/ksYCOz7v4tSwSK
gMEU1C6cTLiQUL5OOfzRLCK/k8UbuDZwGpYa/asACIQE+Yze44+i4BtUqBp9Rkl2PXHhR4dPT2Mu
j3Ns2qv/V/K2a5wrczECIIy4r6nWc9++iT9TnjVPE92kILCoaAXg1I9VT6fPGoBJO02PhThKkUdf
/aKligq6Glshzzb+520EMO39Ictg6lFBeJXUkaQojH401YY4rJOZBFnieEtScTtwwNsxYvSS4UVm
/XrmwvXV5Hqpr8xdXIPRHbMmf9BjzxF9ODJBx3Ngv+tuQHUDmqM9kmMRkWg44oJPRMtKSlh0qkFC
9aJ3Hu7BXvVY45BRHNzpIGfqRU5/Ws9TJPrz6wslhspXXaZBuiHS/kwt0Qu6+CTPv0z7vbn/3L9o
Og1zUVTY/dVgKIkPq2if2XIRH20rL/5aCJDntzyL0AkvzkXMOJJiILRRcORgbAOim/k6fBEYPQY1
mafqWMXqsAO88eo/d4bbeOv7LmcmW4YO1RUI+UcPy+RqN8/0mvYx3dTK+JAePChoK+Eqq8xNnGY+
UYBNZQwHQOPMtoG64IwYDZil3MNFu8sUb5pZ3haWSQyY83KkNPwK9+bnYI4LGfGuMPMVWO7qdMbo
+VOUh/2FTCpGynxtEeO0cwRJsBMar+7UcZ3Y6Jk7PVNf4CkajwuAtGA4DIaHqqEGI/DwQRwNDhox
qY8hCgUlB1A1qeTMKqCgijHSv8piPBNkJhZU2q+IjIIdBxDyo781p1OA7JbaX2nScGdIZEHFTcM5
orgTCJETMktLmJ4/XdGDQGmv28YvEvaOD2kKrChS97v30dRJciZQH82FNcnGjMSDQIJ5J/TCczO3
RQg9h5Oyyo5Kad7LjfNp7A1VXT/8alzAuumItAyWlj8/8bmfjnTG8Y/vxw3DglzPmByp2KgXMw+z
FnpNos6sPXxkNy0mqj4+JlEYZEyI/zoHgAwc9jbl9kgi9PhQOsaT4FLt1qB9lgSwcMTQnQCD0VAK
NMRM6ph10EagB9RTghww2KUC5MJQjPdogQKNdmqQ8cu70m0CFPcBd8j3cxXx8y+8FJvyjtpbV6DQ
T/alG0Q890+QDCc2X1ayg2lvDeYEPNURCqiN3YAsbv0GD1zqiCqq94bAZ1hjgKHjaQ6/1mNSJy4D
rJnqq/H9pcqnI10spj72FDBhaEJzWIbbmSrI7pzplLpfhXOy7pgv+3xYtKtms/hXg+cHlRMEVvng
oLUX0WqtkcdFcMD7qgJ4JtJOnwKszd15q8m9IkfXMps5LOpO2GVmDR23V0PLGKX61opMAh0YTlu/
WLkrahEs3nkPnmF+I4A4lTpPBI6vGVUwlRRqwvZVZJx8isJwlBE3XV2OXP1KXxhX8UUo0qVMKu1C
faHCWOJ1Uz6Q0fJLIdgLH4NsIuvAC1afquydUgBoPoTOvzi1qV7RhltORC01ycu6cC0wbl/0qtnu
G0HI4ZRt2fAML/m0plyRQkV+WDxQ1F3LKoXfi2RzeRf2g2r6VwcWuZJGaIChO5Q/re0Ejv/p/seR
Njgh52D0LrqaZmmb6AxEmrrgV0ajhTabLrL1GK74gvJinPgDst6V9kwtM6EBTSS4ImYQuG7dsLo+
4AvevxUnZZBK9ALNwVZvb1+qTDltC+5kLJzSsi7NWe9D7/JaeCnEmPcIq9I2dCttRsnA6GDfkng2
OixtRg/+kfTSGaN+jUOqh6g2Jz1v5NKpM93KooLKEjWqdjf9Ngd3iFkRpLAfR2OuNFofRzLSc+/A
KMOXS+ksmGC3S3FUIWlOLdpNUB0uz7NVYvHv9Kp5OYVKkBNWC3RonRwc7jQYePoGp0KewH4Cbsb3
F4VWyf2IGx9y5oIrWffg81QUluziHBcaXuATenEqI0XfSZFaMEcg+XwAuvv877smduyepKSFOKHw
Rj/OZuTQOqtbe/Tu1OWkrlOHMeaESK3dy6YfN+rbQ2QMwSyBE7Ia+dvIqN1yiY9td74npqkMAYCw
A9pwTJSvhvNEOhZvLAaupL3wjctV6Fke1Y7Ts1jzE1BXCFaYDFtIMAVfmL+uyET2oIPS6mzhYH2r
oOmQypoO/nrrPOmb+kkln+SI2EPHp6JXjt6JcUBoRxVI4T4/m4eskftDbV6Vvu8eWqvIg54TNoVk
y3L/DJVZd1RBKoBJwXEYK3sss0gkocINPFC7eajefMnb1IXy9ntDArM0hDoeRGByog/oyTfI9PCy
gtkyUgk9h3nbGx4FQDryVyZZ79TUncYwlAJvQJVEox54lAE3X8vlPFLRV4anCF2RBEpF6pKAlGr9
J0p6ci+VFPzwV59DPiCoghLL7s7tDR03GT16nygwb2nsG6KLaajvlR7208Wt+6lhBtsG0xL+Dkwo
/7MADxgGuStg7BOyTASuSTAFeyO0A/IuAa/tgg3XiGq42XnrVlGSr8RoDzklZI6U6ZG/5Bllor8G
gRwX6yt7chJBqEdAqF9YS18UKrvTBo6nIK3fF/1HcibhNUu9+D7WqRdnpzZPBVDw6eUMQq4PYT7X
f59LNErhwdTR7jiAV7YkqVJOvPCktOp56gz5+udFj4DpAjYclp8najbAWBGvsf4rjWTN0yZFxjoT
27lRvQDVTSG9CW/YG81m9FQgs4Otsybss11Aw3aSiLb2FxDjg+Fs7Hfp5OQQjwol+2fh0DEEQiWB
ikQ0I/64UGx+PYhDE2/yBzP75eJB2gb8/6CPW8bMcQNoUSa7PWRfL2KbsrTfl4XH3ZplwFWBTK4q
nJqJAK8Ur2JoQwU2mJivoHfBioJMuUaS0j2SnOWaw7BaVvFSbiX/9JyfQdW9dM4xdjWpznXmUof8
C9ImlIgNUSsgx2zEbQzgGSPMLv66uGQTGB3XvHoyVbRhjjY+v6a+NWssq/1tTUOsqBiNoPoQ0bS9
r+vAH6X28hoN9eCrsiNxOjz5lOYL6voUvzxT/30+PJoPbRgxAYyIAZXM/+BFiesBo0vVV6XHE9Vi
gLj1/XZEbpGHlVCgk3erELn2koU/7P+djFpZRhCAWtnTe3d+2D9j3lJyN+zo7Ee9V0aFEehch4wq
0iyD/EHCWRrNC7Q3ddDZwCFi0whub4EGP5QHiTUr0HNYVs+sYQTupiZUzqLVc9LArbfs1E6kE7Pa
EDUXz2GZ6usanS9uBCRzfNJmYss1bI99Cnvi8DxqwVcN5BVlRCPAf+2lc5EJhS/kaBNIQpOkunKc
hYYoFKRIXQ5gVRJDhIxOzyNHJq4xV3K72fsaqQND3uVfSkxJFtrpBVco6cflsQlqVgqrhPp24ZKD
dc5VEZ1uaNdDLwlj9pji6weQQbh7pN7DvU42hKWIJrNJhHNn6O+9B7Xp6MGhj8xG/nZuhjDb8M4e
cdOKeJDp8EUzGX59DBxFkCsuAwOxc9q/J2XNF2TuEjdV+hLYkbUNfIiUrCr8z+7VOXu1vHvRBKPi
/vRQKDCdh5K7GVvmUaMVTrzJUrTpoYRJxYH07Irw1ZVKc1D/BNgJqEgC/tu9j5vpCduFTUMHUrf3
bxxQ2eBUCbM02kLi4m5bbtaJ1lB68uYZ5rFLgHaiOyCUzQCBUI/3iczqw3nkAde6wJaJMFirrTaz
QgUKxdd3fal+vP2P4Kmg6JTJKIPWrvEx5uzsWaKAzvfu+Si0lFvx5DqgV04EqOIa9t1zLyhIx5kE
W0eXt55AiEb6UuSdYNaCF6KZrD9SJPmJLW5lQxFfQVWaFaX/58O3tHwkNOPI5nJwljXqQrXC4H7Q
KQVhUV6Ij6N09G1fFqQWv4duuHBzZfAHCc+dZjuBfl2qUqsVWfQrF0M/J51YpRpmwcP57sZTbi3r
eNSq9/l4hDNRjbIkx3U0acVqLhFog8YElQUl9lGXwvQ0wID+CJ0Fk962XIwMJ6CMr3b65fu2Khg4
DOvnGwji6KyuZ2fCYsP4mSaNjngaOGjLKtCUd9RkwH4W+3QaikZtiE6nQs9xVnkKDdjibBuuxqK0
s2vPch/5SJMA5CELne6JP3dsQRZNaFDxfVYvsJFQ988b2vVaQFuTs60uAMuitBzLv5P626duZMU5
Q3d/N+M7ZOsqcaene714vg8Jz/1lsMLvFZzq9ryMup4wMMotv6xVL/VD457QY+nLDvLPfR3D4ck2
I4DDSj+RCdkm8kqu/m9glUDOkO746Fao4rZ4RiOJbYOFZhWkIA8sLO+pHVcHILQEcJmzf3gvKffo
WHFS7Kg35mDvY+yJS0ZDkfdGlnj18xezfdaPdhFwQ1LOGjYF8grNH4AXLUnX73SOFrZmQJefa3qu
AatU0ws9QxTDL3oFyjfjbuLybcT98w0G8i02fgkMUmo+lkz8lw99JhP9evozKYFpqtwJTFvn1cT2
V85JuenjT248Hs3NpVmb+hX1+I/n6+P1EmuuDx5OmKp1dpmgSZUIy7vkqpY9K0J/EclHyX8XRxjA
2ntg6nSYXQZBy5ihd/qYhG2Mb28zVUKVQiPmSjrG5qTQ7wTZji93jVw2KdUITdI4ufOnBghDuSYW
dCuE30JUt0r3O6xp8297l1A2/Q73CkujTZJranfx3W2QwKurgpx4KKhEW9R+KwGzTLajIkSms2Iz
ejfeERZSuDjB/0SmRXwxy1rMAMN7Z69avAtwj0XjHSsUe2mJAON1OIQYtWoTOdFebfxF9sdBkkAV
yLN8fv21SfqL7Q9m6rkh1wkTRcj73I7lLtD15siWZ+GLhpFm0q+Vj1w/VLYhCYxQdOU3k6Hj5HBN
kHKQHhG43DKj8+63wKdcoTwvZgfjahNpO8pJYN1vGXu1fFQF7HgQUJpS6a2JkITmheb81wif0Jfl
RAQltMuLD2wUzhV/5eqOs335qqVXsln7ZijQabj8LUDpmsNlFyKBF8C4izMfRk9KdlhWcLDItFST
FPhW3Su3tSmNCm9jC/LBJv/rnswYrRmfgT6EviVTRsqhWbw08uAeJbMLTnlmzFz9I4m6TGN+xujy
DKgXZ4e+JEnNztIHXjBoJggQkYvG8DMn5sHFoIwbdC0NXXilUgmCFH23OWCx149Neh/9M9bHgQqe
vIYYc8bS22xom15m0R7kYIHWphVsFRRZ21wDvtBIsqM5sgif6l/N+quv0DRXQACSTkUDiIWwypBI
ojoD5ldIOlj+rRlqKVtYeOyBXk1odclDEMWA8IBUBHks/STbr48Xf7gokOfU9S0nIGmBeFF1nAnv
lq2kdLnps96wXAOP+e0fr5b9j/lIReh2Q9xt48a4NN9B2vvR7UOo0CxOXu+A/MHahOo7WzVPj7R7
sS/Ia2CaVyCb8uoJnB6zmWkoRw25MGbGI2rmpoCemr+Sv5/Pl+CkBUuUhs9VbWgz6XzMH7x/CqOT
9qSWGM8FmrZxwp09dh1PntDTOpJ/XsVSXdTz9EFOkfZnJqOIPBhimuil9cUTXsONiL4/PgsUE2UT
kjZYlf95atw9G/5Im4n7JEYdmQbeZQtRp29rB3c5YOq//CXPbbplS1TyALtuHkGcHLX89RSHE1b/
SL8CmwB8Po30zI7Dyu/fWTQyGdy2kATJh223bpkeGaQ/Qg9dW1GFLOlSD7IQ3LPkhfjvTzKDJFyQ
L2TEobKUf5nPxxgCNj7HvVLW1nIkQy+UamANvTtfbYKj5w6KymC6SS9YxMvLiAqF2XOct1QMICx4
yaxPsKD8F6y51wEXL4OFq/AorjOmSqJcCBlD1RlcEn3q5YktAHP0KF4RRO9Pb2GkO3AQS85HNLlW
+l8vYD2vmhfsMgecusTv7fwa3/uaD14WDvwWUg3sfePwtZDE/BD+3gEmV1EHB8pNFsAarU4wAWnO
hDgUUh/zulGzyDYvO+QnKmuL79zCj4prGlflyOfP3EpGtc0fWQgw5KUrwilziliwbMLOwfvsj8Mr
27rjEQGUhD9NfY25g0IIVE/1/NLmuLwHbr/eRV2j+3E03/LsDn9UMGljIXyTHnTtVmS5OQ4/Zg/v
KLjoYTrvx5SFwyzbMxxJHTsN9LBFhd4eURoDD51xuCvjFqYoD8mtPqFJtIY20qGRWPzR1LRcj+pn
yiJgjbuG1wuc2qMSXL7Z8KClO1kN8oBrC6Q83/6ndxiWxx9d4Kay3jISFLZieAoD/PwNxbfN7gr1
OqfKkJSVE0JXRwqN4sa33ng+ytU77QRhA1rgGrsROKOJHZNHfK+NdT2C5zc/PNCr8/3mPP82Y8Bm
4duKzFxB99XbWbW2aR9bKzwOBhRfNbrZpLfmHZSPUoe9zDEn6LEBJAFzMs68xPqA9Ra0qiVZ9E/5
698yUot7aq0ZXi127HY86zY0j1W3RF8MR7DOWARAEyJ5Ur4v6qyq5Cs2a18JJCE6OCxpZenQwPS1
xRHGbEBp4DjczgIHVqCyU6cKMxmTs7gdZGjEuvFvSY9R5hA8MMkobFToLvvJGxxqef69S33SEoD6
piFc6GoDf8Sy1oAQ4c2Lo0iA9G/+6HQuz4fC+2fREGW42phMfGL/ZT1zXBVQwDJcRKVyNt1YBsMv
bTNgAzqyB/ylaWIk/NWNkRVn4mqp8baE7wYwIxqgXW254s/HE+mu1rA09e04kKvF7XhgavDr17Ug
wD/6ePoO77AWvSVqK5ZvBTPnqu/OlCHvne0syhUwjCnN1y1Y40Ikl6j2WRj+6vJRDz5X0XZrh+JH
HCqqSX3jEx56LhpmqvlWtZGtM3ad6Mr5Zs0w5d4Zu9pYxGaVcRRsHPZqVHIE0JJwNc3TPWN76tKH
Ya82bz/NW3eCirVRAjbrLDBWEnrKYg52GyDCnNnoqCGDaFnxgFEwOyG2ShNKZ1QwZxi4aD0pYaUP
zQUuvfvOV7ipUAzztWC+l2YNjTncYAmcZrCndFMeqdYZpVPPBPkZHuB6QJcC4DcIXOjM0iGTXFda
ja/tkvUsgf1Z5tzgu5mfB33/eDHpXACAnWJNvY7h59faVmU1JHzvLW2bD7UfzEd1OYDwAVEMmS7d
L5NGWccsPsuWdXPnKB0VLoqyGlUWkqLMd+9GjB5qmqfU6j40zR/cu2ufiwSIM0EohTQkdEQlX9I8
TNL57wUsPzzLzIB3qV8AliYgP/3iUt+cAFwxDgbt5fQkYs9NR0HRuEvtXh5p8zUjRVEjSQD6cXY3
LOim+cXHj7RAzFixf/ys14Ii8Z35AMOJqhNOToNEI8nnbE16MnLeWtcrW2GXckbuxPmcDyEAFIYv
xqAvzl85ZmP5vJNkp0MAt6jIuuaRNptvBAUufcqpqq5Ekp+FQsTrX6h+SqKM8JTn7WNOh+O/yqxr
vJD9rTufJIHpaDxVnFhxpJIAC35s1/BaBVkI/k5QFtJpfCmO9YUJKkEigQAgf8oD+gQAJHzewqdK
TrVNWSLO5ReJZFmsEqRYsXmZKXY7GNXsF5HWCSJpLMV8AmcRWmFgUYGtfahnYZV23G1oCktzOM/m
KOSJFZCm9wYoBcwz3q38JZVt+7XheqNTnPbB9GxdYH+dHcDMW+FS3ssWPVl1egBLQwxk2lD2c8Ps
BDOwLL/PB1cCqfXiohXkMlzI6H+NOxjclqv3M+aSpVElhN/fEemzD1MKnNCahrtH3ha8FRXu2zbq
wYvIBOVf+hmtTtGpJLhyFKDrASrLF8bmU1wAWqfLfPIz9PwU2BotxCy6F1Eae9KshI3ECEm1PzTa
Rb61Ul2Bxc1FBXTY7nele5URRB2bey4V54quKbLDLzH5kQCTaiplc9eVhWMlRunTVx8BDzmekCUD
7dxg6AqyLc6GuqlG/QCt9eZEdw0ynVk9HPrDiomGIx87SvxLtPNT6i4XnQgnfw0ca6XW1SK6eCEX
2yzhyQ2UH8LpJ23mFO0A7qC9/cJIyljeFlcjIZvR5ZTWc6kAQn5S/Bz5m7rSsn5dz5l6hDKRGBE6
Kw9Sh2QUsDyMhOxm85HLx9S/ZC6vSchmkYjM7Ads0gHsJnqsrxeEoVNc9AYIe9B3Yq1SXFjoMmx7
HsBiO4GAKBndh3Brt/K4TEC/sKwqvDJnNXM3jiSHbU3oAMx9taHMbtcSmLQQuwcarbBq/1Vda4SN
Pusl7SrhF5ngMRf9fiwEMC360duFWqoZjWSwsmBNEgAZ9fPXmW1wlOAX416wFhGzjMmKcU416kMB
qJ5+17aiTobELXTP83oHSevYeqqiHGmWDuXXd4lhq6j5dtIiBgGLZV+nJNqYDHsnCak5nrfw2w1L
vI9avF7+gNb5ZJUWfHYHtAgtKoPN13dfX5SrkirXEh+bMG925pM5EfbQa1Ct62SSLksg1ZB8963D
ugR5iZXE5krFuykVWSDtrogK47mQqNLAOMPgtdHodAqLhk9yHFOVbf4+l/tLlQNsjWKqPNkPyU2x
Pbz2wpRB+BEQliXdPTcx+xDHqkWrEx95cKFT637DTvSuD//uUXuGGkpwYmV9P1LcqKK0FPp5AJUQ
SNa6KiLasOuuE38wrcOhdPZOMZPE8Ar//460qtRa0WSgbh9ybZa95dgifcVUPpW8kcNB0tr8+pIC
sGdw5LuENawK77atNee0V/A0lz+OJvPcWhnFBKouH4jSookoPDf0Bv0cFkcbFiPK52qkulnoG3Ew
OZx+b9T9evpF2zegor6IBE1s0WdZZdAG4WlTbJlhzYUGtkonhRFIyjcHRQn5rvCksRkZMl0kABZJ
KPPT5a9QmY0rb4VwvEF9EGcUE50bJt75U/+iuh1NSmDp11G/DjAuSGWhesjdUcQV4Onu11xwNHYe
T3oa7gq1vtq290+cnpRDca9P74HOThFlgKH5mmF8CYdgIT8Vc8juufrVmIm9/oo/ADDjImz4TTeO
0OOAdf3iRtwbPNu/KmWK5xuegqtA+pyNpZO8nQ50pqq4cfPwPKOrd8MS6RM02RG2cYoj7px7D1Zk
jjLjZ8M5tfA7NO08J2K5IFCtsbHxhN5TH3i6xJB2NFGn5HjD+Z8ndgTEqVPKMmgWS8vCGwtsqmNL
36u4aw5JaEUkWl/JE+NkYMpcT2VOZxMzvGECFKk1J/sscKvvv0CHYbkAAbQXPLKCqQZ9LTGCvls1
KbUrXxR57hle+zM+o2xvIPWaFuWvqBFAxwz21cBGrRiIzxCm8DUB7U/56EhQE1/aCCCuJoRfpOjJ
W6A2OgHlcS9/1dKPhOqpIiwjZorbR5sjDfMdANSFY7uNIuSc+xOdvrSCsP4a56YjzaAls/lkifBq
80kT7Pfn2dqKyctkU5XhqZEcaNrRyIt2Jb1+uuCx2mnAnxxI1aJA2OEC9wLsd8etSQw0CTCwbmro
w0W7mayX39z4S8VJzcSfiNE+Sd7vdHK34fLD60mRRfH4nU8CdoFyNNAmz4YeU0/kTsDi3dl3hHB0
YSuTY+ez+vj5wVREf3SUbRX1iRHfdvmz8mxKn+IKJuYai7kR5s+aMv9lw5DbEUD3/4nZAp86zC+G
JQCLa5LLp1/1HuRDnTSZVrTeHccnoYAKPd7p34JUnepBe6AP2EV8QyKYxB2jiyr3UDyqUqMS1XxM
RXITrv+mWUxhSQ3WPAJMIL8VHO9cqrlmtB4a+8M+HZXJlMgcNPlM37iG+/6U5KgKKDqAXuOI9D+r
TO0iCvECmE2l0ucxQfaQY2yUYg6L31rqqEfZ5qTZp+2kDWx1WWOU6I5nar0AEzGd0rlez55Wvp2H
SkVscFSa7pMYjEPYlhgsjbDE9N0sr8vj7gnZo1RYmc0HMHlJrz+5D8sTsWyN2vzXU9T95U+spwJ4
FdXGTPwmcdJozou/4bTUZ1IXAZt84vL+KOQT3bNmTxKYFUv+5YfSLI24p4jOmYQRzulYOYf2cSf5
ABI/FrFwM8fVPogHZ7rIPkKf/Ia0yA/5d+2DkFU2GOh653z63uDF4uJu4qAH3XisQHIyGW3MgEPu
zqVAMXsxV/9LrPzekuieFotHdOjkB0jChENKYftZv/1ZS+KBr3P1GYiu/KozhrSScsNJihbEGMKR
oOVCkQ/Rne+Lf+Ox6V8Tn/vt+a1eCSyEwlkKH70dLcl2Ty31/Nb2nPsLosAG/zE4yLDkdpIeks6d
I7gT3Y2DpW0TwzEzXFlAxF55vbzDbd36NOMqG5TnJ+DlBuJ3gu7F6CuOBTZZW03Yy2tvJtQfo0mg
RUoJgFwHwB4A2aFCFsmEe0k0FSM2nMmaGD9mHVRu4q8NqPALbaOzjuAhiEZFMobfAiKcLY1imjUC
4it45hKjtDJtFxmJtubPIKUArGpFUbrtco/NK1NWlxTSMPkEEaRhfruXFFzuwUmR/NUC+S3wcAfa
G9iID+4uqy2EU3DsgL9KVTL5np3ha6wFw4WcIfR0rvHHMHxwxOQEbWbdOoBW1OCx2bD8P/Ev1jjy
1uml5zcNcIpxHDMIFUvayesqrac4wpbczy2D32b1N+GEz/vwGXmQwJTH71hcWCpXGzdOiRDQn0y9
7tK1njA5uyr9xwdfNHw/zbcgTR72jetS7cB73xBza/dGEkU93YE0hcR7exh9ZX68TgwCHgmwdYP+
nT/tJC0tPyoBlgm1dCtWdKPO7jb2JdgNCUDWiYCfKdAKTWk61XmzlovAfMTXfiP8cLtnxmvSOOD5
8/REXstZT7+J3+7GziaI2/hyVmYn+slFuHW65VGRnCyeZEu62J2iVL0r9JuP+wsaMzRFPH0hESC1
IOp07w6dbHEEmh0KVmxRAOqv7vQYUjDJ1MZfO3TvuqgEHg+UPttHkLTUfthdX/rdHq0ih+d14JD3
Jc3IbYJ7P+eW4ePtsoa5sL9nIUJeGZJKoYUXwgQR0bAupG3kc0J5b+XKbBLuqwUmHbBZhhEWSYh2
KdAZT/x59Rg07RCjBX2/a9cwx5q4luIm4Xi3k4wLGMT6/ZEFNXajtSFgldTX/n4RbX6ehNkdv+uV
TkKBpNe/t48bmtCbSt+7dpR4FhNODRy1JWiiB9WwvEfuAT3eyqgNlk2rOxiGP1uHj6MxTMhgv+sy
ovjWOfWXUFWQPIUdKn8ssAyzxws8pl+GM1ol/k5DWVwTRTCoeDu2qmFfy9nnG9BsUulXD78VC5DF
88pq9p3ijeHNVXlk/oD+L1cg+Ig+70KYs1AjMWubW0SC29SaqL8VN+rzgTlzOgzSd0vVVVj3+Add
q/0MsUOu1gLIK6Ir1s6I9jNfkY0B8VTNb3FVRiOofB8E1RBdOYVJyEeh4Hjj1/QUwV8VsW9Yw3xP
JyfL74lHMg/QjAZgmEHEKDRWMfj7r1PmUnyXmkQCuAJ7lAlt4KeIs5Ri9lChiIr6+NdIwqKSRO/M
8lXOljgy6vRCMRVgPAef/vD6ZMPjx8SWafLoLEjD6AvrbZ7C2HqEIM2KuzusqX+zA4620TBbrsFN
qRfVhM9++fdTuLmoXOlhrm77UR+gzBhJkUj8ctuVPawwEENwYs5JYEHwyxDb2L96mwwCCRH3d+G0
5sMijWLNet+1swgeM6p9iKyyyvF2N19P0Mcx6fiKbmlpKojdnXJjZF9wzYhY4v4+8XksxZI9FBWn
U2ShCDJUlvknDoxxQr+QvI8I5gsSgLzmxVfwIIyV7i/ySiVvoZNtPZAlPYTFdJo4xsKAakYl3z+J
eWIMsTIkZoChY83scZrIa+WuQPKSzDY1kbMwOYP/3psQRvzVy3eW9boadm/PuxJXUtxvHtLzFRDT
NXAasQb/VmFLqUAJR6g0pdOuTRWcVMA0BCOEF0VHiw6QGsf3/02PhLlvMr0/IId2i6MGvpSmk97t
I5QqOKVJyTwF5hkH+PhP5lu/Fui6qLAcHxH65bAC00ZWqREmFrf4raHGo8UZWhl2vmOIaFaQheUt
PFk1fg1Z/NIcU7RkyR8swkOdVveRX/tNg1a7GAccd0iWx9rGGuFMgeviMa7xHv+vK1hZnTD2nKOb
zGdtE03ZoUH4sjlsGOHphKlkfi/f3nGRC//qW0qfRP2FLK/k2QKZQW+dEPe2zL5FTSU/eRKEj44I
Wi7Y8QNAkGgAwHx4tMkT0WUYgNIgvsxgA2ENWSQMFvclKIcNJChT+WrYlN763oft7jbTORFd15aY
fzRKTs4fazrSymI8Vz8nn2Bl/Lzr+rj/E3DBYH7fGq0XNF/OYJ2A9V+DkyngWKUmr+Uq97koyPpX
QRto9TY11gSIXc9vylrxlPBK1oqsey+rzg1m3nOdRIVPygwq77NLhh7t/vBo9WpRiJXskmNZ5HbE
G/nfMKLQdFnPQCQU5F1wEJf2c/O+PuV+F35US5NPCUSJ8pemBZUnjw1mGQwhuSw/ciyoh+fVIry8
LKE5qDgkvbOICa3x4HDOCJwtZYDIwAqp65mViBPyGy9UiIxt3Ch253JwsHg8w1zBVNdB0X6qxejH
jREXqMnZmFwAxRdRoJ4WfgyFkmHD5jA7RX9YBMygu6qg2PD2bk8QYoHlrJTZOG3OsFW8+27KOUEw
L3wWgCQGqXSLJXlzjoIjGCzS1OfX0gY5QSu8VgYACNFntGRbegw3Q37aTKvTAxO65GgzMnD3Lt7r
UAqoFDH5fRM/OLIurPd0nrTJcmyhLZfbni6jt3tiBsuz7AaLwTqXgL501kFvYhE9DbCcRHAATBdX
dfwm/K+s/zm4e1AW2McIsS//A4OyagwQNLwEBg3LLYfgFFXXJFgfgdKTYSvPn3QEEP4NwHnCqTt9
knVk3AKIKc0x+/fEAwSzM4U7dJfcBC+EE83TWw9fYRE2QKuXs2kRAmoVLP9himEDkaXOMgKr9wTJ
YW7R3rpHtl5JIBL5wCpYgkQM/QVGxgWgzxwBnNpOMSUBVqI3r4+FhUff79VzefN88c5i6kHYdtTz
Pzdbx91yYgXYpl7AYmR2epRP96s3mvTmRGSZzNzoVecjIzajGmfQF7v+QL3ko1MXCn4X8RWQwdiw
whGOo5K3hIAFTlh2FeDJL5b1fGQAw7UQC7aj63KzQPjXzywYl8SA3+tC/C6Mdu+6mgzro/VjlKbX
hr6jq0uzJ8z4ZIDIJS7/lAD3VrOXhihgjngqH2EwsdHs6fcKPrtYYl986Bax9LgqFbzgo1u/ZbNE
QKw/8rkIdFFQrMJtr4uIddiOYQKR7rL9RPoQRPBqFGCs0iHMU7L1GibG7w9GJEmT3c8zCw2iXupA
YrCB4bEZetE3VOb4/CLDqTL2PHB39/uzd5jBhsde1/ST1O9Lv9a8EiOO/B49UwAdImc+gIai9WUm
d/QUwLTyrMNMWRi8tpz8qp9GODvjQy78QYgEowDR/8N7aEnjdBB5p5KMClzoX9GXpYATnTUF+ojX
dZrCyJeZdVFHIRl7elw+tqEz8TYKkAcX5KU8dvMb9tkcrWR+JzYRTIDvyHwrSeyedTEpKEIPtIRK
2XNbnNCK/SefyImBkzS1CTVCmGyZj7cITO0FlifSYbtO88wfdiS2J5f5ONBxmPjySWTY9COU0pIh
Osc/gvzFEq4W/qcc/061z/jyEr4usJIiN3uO4hjZgj8X12DbGaM+OQyb6UrPB05paKb5N1M29ek7
veb+TTAtf8kIEcR3nl6go4z0/9FWoMv8LHilcdQ/hdFtPD7pME3eo8Ju5XbcLWppOWZUSbXxgvrP
cy53y6rZBONkiKdONsuj6aHQwls0dSILLTeFFEHPvNKPGFMbMfRSSif5MGII9AI+tghk21W7aOJ/
F5HIZ0FmofrUNc7XL7iIjJWr2d89f3ESFXiC64fCWyECyKpS3dsLsNkosR4tbyu9D0Yg+m8vFJHo
kxaTmV7hwwh+UBt7LKE3b0tK0h4JGZlPD8nszZSVptCrGFaQW8pnRJuAmVGAKrzxFL/ExAH2oS9v
Xpc58jZNb2FfXr6MyC5fUlEKzmU8UAfY0gfbQquBqb7JR9d3CGOLpN/Kuo+KW2imwqueQ3Wc9w71
zl9T5JJ+l6WbkdXLUuOY1yy7f7ndyzg7wmc6RgrvwxMNquGJE3Bksk9jUbYVSUYh6amrRpNTmyDc
IMyF07PfC9mcNp4IZkc2rHlcBulP2D/U1gBXU5dQqmyAA8DD1QBidwT9mtn6C5i/LPXI3vynvfmJ
LWLVfxHOiKBuel8Ewx519w0pA608RhJtWnEfmyDStqgUixGUUsdrZtmS/Ku6Iv34wUTZIjdc5mZi
yWX4IdXJaqTpOwjkt6fr9UNwqn4bRPyiWfgigC0Ot9xe2w6g5Sh6BLX2uiuVbJMjajh9b1s7df2M
CnvaP6tT5a6dGeycjR26bqpa6YNnJqC+iFV/AC0XzdaRWxenR6/rlV9iW3Wb1EveC7mG1CXakHvN
kLqPNSikOW4PTBWl8R/S3Gwo4MRwROspKCbJTe1aXDY10FVhAOrDdPcw8IQvFjxjPzgoNNpu9wk2
x2HStZrZVgcNz4/pfP//GjrxWSHYmQM0kaFcQhFEK/hMHHKcukEQsEOrBCxjqW2a7lV9bz6bI62s
QvBV3Wv38P++ybgWRB/w6z7Rdq6A2sZP/TgI13g66O7pM5cXGEZSZSZ4qJlPY5woAn0WfirERV4S
AxIMmTDyVgtu8XtQ3M4r9cBJHKh8q5s51ntMcg0ek5hH2ltJNfkIfW3kX1GBoq9kG7iXjDPhIRrw
2PqCSHCPzUqVR9saT5xQgHcna+iTuIlCLPQOjBDja6JIFk/dXT8eVgQesDZ9xLX2bUMHEs9H6Hw3
bI8CaNr8bNP1p9XvzZ6OptpAYX+D6NEpXlFfVO0HbCjTvWlYTnclbYBIBg4caK7PbJOkiTE8cRAq
zAS+6kxKvBs0Arw28bRkG/A2v72Dvm/pqdn8koYrW5lKORDny/FmRdZV+u8cxQi00EQkfIdoc2qC
y6e8yl06xWe7ARfhze2F5n4TzobmsVUKxIUiPJwJmS7/vSCMM+SFCcjcxFztOUnZ1Q8V485g1+nX
ugvG627Qay03T2SFpWoMM0bgXUoHc2hi6uIlwM1ZuB/XH6uAkLP5GLzGm2coZYr6a+zOfSPlgYXq
oPO8cPhQmPA5kG2yAyHJYmtJREo57PU/k4HdnRCiLeznVamOkQv9NFJJmZRqV+rPMiez5UpxfGF/
eZ7aZeBK1Cnm1Qm4MovjTcScogXZdrQkXLdQiqQwBXGzoSrJFev9yTId8znF88QNXwWR6RnmWjrA
MaqJp9t67IsCcRGIK/2wLUyuoLCLnMw6rupArMyVIh/WfCdpOE3/o1S41rPlAi7J5OFJlx3my94C
CoNTGOueBIXnUBc2uuYga9sRgrKpgGfsjam+FCOrVE7ZrQgT0cUhxtowfe2VDE0QlnO9JYuc7ZWZ
9LKs+GStUoA4ActtPF0X50EgOjOboaB48sjJGydkbikXnDdUEsSNN98/KFxXHnP5Aa1zPCrOrDRM
nrv+Cau3QFPsP9FBd4HLyGq7VgaXkF986VaORlIZ3ouvYWBs/STTyUc8aWScAse7M9gkeKbOnPPV
o8EBbnPYLg+EMcWdqYzTQeJkcJN53QYDs9proRDz+vPgvTy11/u7+XHeUUBBYdGyI0KWaBUgA2CM
HeW9Nhdtrjckv+9KiDJe15nBju/7w3q6FW1ypf2d+sZT3qlev/f/MJPsrCLs26wEX0ko/k+qXPrE
dve8JfK5WVSQeG6ATNjKC348NrYJ/5Txex0Xta3WNHv8g/rUYqixUaFbNU8OZVdljr6T+4ptVlF+
eCgdS9FAC/ON39FWWq/irDJAH08oItuYvCpSMUD5OdeHHQLKNBMlVmBSmLxvpXeqh7m6A26nycIO
l9wPoWqe6wgBD1F0FlYo0WXo2ZP9HW4euxK43ImGrZ5v8OwS6MJ+mUPXBctC+b+v7tOW+k/DQxq4
XOuW7Kk0DL2EDL40zKfUd92Dtg8GxQdGJd4jabMVFxdW7iQ40P9sjCr6glARaAlJqPCdIP+50h3o
DRKHHf/ByRmZE0efktE2skyjnFLArjy1YC/N/VeGBIX5udBVHKj5Fiu1R5dtW/9Wsz0ZHD+bPK9r
K1XgKCRx3nkzqEBUU9hzApU2reGYXjN8IDo5IuhwgUyLqmoAVAdNkdoluau8CidvTYWwjx5odA0H
brq+LwAoV6H3Zeg4f4/YVlDv+HXBG+cVWk6unePheJf5X9X0R27U/8Ay0cyrCdoSqSEumULDavQ2
wXppWwldYl0i06+KpF27nBxSkd9zzvVXjQ/lo4nCGb0p6DFEhZ/Lmg0lcPQWrSkElEhO982biMLk
IM3eoscTKgHSrq4NY9DUtAgA2S/880zQLht6OufB8S2E85sxQ+q6+dOwuSRhPz8Tb45GRM8TWOEb
iOpYIqvEN2KVRJpKi/YV+l+GRDmiJFKJ36tl3/41MQehtxunLF4uzlE6CUkS1JrdYwCd4YKISSYm
lSvosj39eooDWHNafFIQMZE1yS1rlVhbplK6A8DQEPJGrYpg3ZMzQp+psZfMfoIWannPzEHlXWIl
DLNWZ8WTh7UdpMAwkdG3+SCud0YN8JGV6yTgSyCqN/VNYfOnTkFQv1gc9pyzdGh5M+2PytKHZMWq
EGu3xivMOBdDQsitjGentm/t5T4xEl1SJEfYL7n5jFUrvEdCdAd2W5OCPd8JUZA/AEEAg/wDgJp2
o0d2hbeWfJWUF0dsfH0PWMyFNBpKUAWD6B6yfsAFSpkUCtd5npuslhBHNNCarcT2qOhc7iQAzf48
1a96QJUl6EH0iReEp10nzugAJPPzubqqt5gbtVFH2xs9mR9FZkZsY8EDJrLUyPp/9S6ugXTtRoMp
q3dx2L3Niq8vwMTV2RQt8cU3bIWJihAvYmc9xdxRaI/GEiSqp9tinGu/CSjyN3J6SBb6B4AtefCM
WD+foKEoOaeJ1z687m8H+nQphnL0AcBgErTSclZFz5HWD5n6d1NkAuI5pEAD+AHkZ6ZGp4VXbRbo
4IK8Vv9K6s75OK8cT4IIlgShTktpl2tjm3yzX/VHDXw8TH9420RId2u5toHmiLPmHvD5qkkkJNbu
KzDyq7LEBLFAGEmXjI5UkDg+F3BfiZh/10v1Bi2AUyV7hxBmjbM+CcNaiiskVZuyDmg9bOb8MQaM
Mwijx4bUCgQrPhbYgIYPpLTHeJb+EURoQoNrtRfCl6mn/fFAg8wDYIcSGb7Q9SJIVD7HXF48JEXT
iCnefbCyEvr0CiDrz5jK58YxNjjM3bmVWpnCnpVPSOia1MFjmjKRMAvabHJb9B8FrUsvqLiXLda4
5TfUw9IzGGHfyF+7qC7iboEq7H1CxYgFzvGKrAsFIgcARoaFc8WMZU+VsEVTRpKVpxzebSRFbclH
E0d8QMw5QouVSV/UIEOuWkKxCerFoIy6+6GojOQMwoeZDaKs0Z0IB9GV0HvzfSsQ923RhQApo8b7
qjgewCbyvq4cqBd5ABtRYgTb4HaVY0Bawdr+fl3aAp3eDUPM/sxNwDjSLhQ5bmlj6dgKAptRO3H4
ku0dzFT4BtSWPYdChrqnJ0RD952DB2hjjzzokxd8F2TjZxEOYA4mrxQ8ynJMIGyGTX1jjp1z4lDs
D5h7odCuFk5HcMVn2xDAnAWGlWBAlRZK3UXRJ9KKdNSu8+J1XID3EkI8AripdRtEAqgMr7dFTb+M
XDRK6lzb+R+qOyxGcqa55p1gCjs9b8OBp3eGkVXleO4ssDUKE5YuREO6SfjehSEH/gzgBJyWD85o
/xkbiHIsiTHEuc4L4EStkHthu4gm/eKKdXDnYs4hYZK0R/VoxkWKpaHlKPHMDr04x9H7SjZBBFeu
iC2d46JsOKL5CUe8wPyUC42yOUvSLhhehJiTJIKAw6/UKTmNKQsiFm5kI+nyZy4RUyK99idObdQ9
uExBa+n3Mzigao+mlKg2UrEahrPXUHfk208hXqYLu0XsR4Js39gQutGvbxsl+OffW+G2tYOr0zNF
7gvrTqhdWJ9IL/qxYvpV6feRa9X1QUwOPR2nMmj8Xpi1nawm5jkYAaaZeoTzGGgdnrGxtmoV4l6/
oystPOto9RndhZjrGIDbM/M7elYoiImOeSMsBXEJVNU+aTXhwQ4glVRbvTfMajun8r092MHMmukB
QVoHu/MR8RnzefGIXVdvjpsNpvJw1iKr04km5T0qn3sJ2QsYlB1o9oOm26lwyGYE5Y+D+kPV61dg
xqvqweiqxyppg6fph+uFJXyMI78RIxSoIzvNnV7shpqMTbPKBw8k0PtiSo+w27GziGbl4vaw7SEI
3Ny6QeF/xKzw+vA2cqJO/bpJzMMc+b7eakv59vKPO7wyif9aOdKaYl2+KApDmARByiEBNjoszohU
LjgD7aqf/09hQkRxywm/xxZ6B6ElvQLIGumZOgw+zKMq+FkDq5wQkyy0tHDlBNsDHlgR3AVk467p
hohC4zhcimulVYyml6LWNK1eUjLTsRuaeU9LdQaJEaykCh8SrQ/8r5ElfdEcduzWSImlY6al19vz
mNJ9ygxYh5t/Y55GcgVZJT2HIg2hLpVNBysCZkQW9zAmkgUAl73Mk3eCeQ37HRn94rtB+SMs9IDE
eqluEFvPuOwDUSblSFB4g4fJm60w+ZkZh9h7tYOWc4CcUbqas6k/a3pnOmirOGA3cTzxyPdjSRjV
QVvP3rw0wxFiBmLyUE8qXbv+GOd0Je2x4vs/3obGG846twPf3YU3f83P2WzsljEMPUHwZfz3YKjp
GLou8pihiu6ruYGAezuVKh4L1ax/5gPn+d44MdZE97YL7vJF0QLGqqe84X3Zxg8VMp2H3f2GgBRt
kOES7mRtexo765UOnvRlGMZrpdcI9UWEnyBiUPgHdPNlfLMHszkWmZlhgo8Qo/yBwljsHq/UMtXE
3ovpM/QUHG8UKoyNApSDpczMRxi/4MqDKpl4jGry0/OiGPaACX1rcMfDRztyMKvyLjomCLeAUusc
w2eSBbTS2Lg0gBqpGeK7rfU327AMGR0t4cRb6VFipu3oLa86XXZULoNlZxgEM4ZeCjPb3GEz3WJG
Px52lYUDsYIPpwjN5U1qiOG8MJocLAUyrfV2MRa6O94idmZokbw4EkPlBsyzeTdifVi9vWxtoVtA
NLYYgy4qW9olC39aNKvQRhO7ZZK+AV9ffSRRZVWWz1u8HCRvb1wxkDAXdAa7wotf989wHZX7JhG+
L6ubS6DJ3t7j6MVlMdM5pdvE9wSlXICcq8iXYPRtb/qvGgkcEGOa/gcpU8g8oWEVl3frUO1mAued
u86CRIYAgNtaxsUfN7txPKqnLw5gbSaoL8m2JdcqI7/SRrkBmOJeN0uXT5akNfSnxY18etXdbU2R
Bg8mmrJ5DszsDl3/85TgqKMVn5EvKZuNE8XmjTfrmQHtxwlW8WkEWe0Y3vvSGfBmdeQUX7KUaj/K
Mvb34JaiED6JK13QoG6LDCBrz0AJdY5f1mkVD4Ckp3NtcCsh+qADJjWG/oKoPIYqCDR0wwXDKWEg
SkSk0j5DiBYXeSuK0BydqAmS51z3X+zrXjSWHs82zcgNy/TkGL67S7TlkWcnk9tBSjdubYmzeHmV
oEDUhxTUZEuH1XJ7TFC11xDDAgNzyOJG4EkjnpIAZt0EExfVtxxA/X20rOvKM3/CpUU8xNDuj+FR
rNiKbKwFSkvZehaVGTG2HuQFFZFDSrfBOc/G2BcrxenJ02jOTW/6wqMvOz+pkG+IqLGWoBcJb1yA
cpi2DLlkir11mCjZAWRAFm52bf2J6oeUD3uhWLtRXGhKIP6zVlJX9WnkvqKorl2A2f/yUxN2/Yjg
vUAqCOxIGYw1jw/ueu4HErI1EXYSv5BHF+H3xAlWXUDwuYtuu/Au1HoSEZaD/LPwG5u5hiTkBVxk
UVhwpB3JNUe/ef7Bi588U66f1ed0SzxphDNmyNi34NOERCQwUPTU+CDo8Us9DhmacJjaSNmm9hrD
DEYMNrrZRXHwx6egiin6oE6BsSWZu3VdZs15L6SZqBBB1HWa3g4vLkL7CxK34etXVhStZx10vcs0
LfSePe+Qq/kKfTl2VHAj7Grt/0BnDYo3n3rzgOCvjrhX3E3JsX0l69YgmJL9bS+Y0dLjq5bA0i2I
/EUXbj6Iid+fGlrv/++B9UWhSligl2iNinC9h1/W9Y7pPtWlL6vXrYyiH/VHOJ9gNhdpWsx+wPfK
rsJVG73L6XiYuj5qOP+PVERvm16K4Z0/dPf0q2y/ZvKY+TYtBUbECyci37xvoZynrpC/utkmcsDJ
OYKrBLMJs5NoK2OBdakwC4OuFSd7GJOZqZY6Ixqs6wqrjm3gsAVmB6dBqAbJc9UkOyIeCCU7M4L+
+R2IcQuvY+TUsHG830WOObZXPIV33sOafsdN0hjhX3Xvvtx+04X3NXBOanjExBKk5ylXJMj00Wkq
59bo//FEp9ARKLhHZep4xw16obpg7CexhsuqV3BSdChXFnJf4/Xw/7GhKlp/kME3QZcpx+SdnhDf
82QXbzsx5STQgzt+NuKCa4yO8CFiEd99KPlov0IJwIYMVKtzW2TkQvs/qC/bPjC+JqAbgIC+pU/4
JwwiBzpQNm6IMPMx7NeTfjUb1dv78vU3pky4Cvi0UXKtCSLuBywYe6GAgfD5dqB2xkzjLnoOUe6W
xjHjjO2Zz5bqv6c7nULma+tZmk4E8cPcVA6aT1aggFY/P5DNnjygoM1dhbWe0627vcP2+P9NxRGy
BFST2qO5bKANDLOUfF8duPQ4Vm2JZIZqoDXcOR720Uo++tKMTaY5tATxDlzvRNS5keXT4r9nvg9r
oEOOIyBQOM7iWcJoc+f3GoDt2HHEedpsn/6HZ+KdWsOoWxxquVEPIRjYsWIdedjn/6eA3EO1b3rH
Kvt6jTFlCUJDMptOKI3Bgsfaqk9uBAWh+t3PGGpOxfaQJWHzSv3+OiPqP3V/9AJLEnDY+2D6Tx+2
QfdiaSst4u4kXmETDys5QlI1xhlHKQ7qPVtqrfGEMp5d+VfzAU9slS7KN03rHz3rVxs+DB8POLll
gLl95M6KKlMmfYemBMDdXFvCWWebiqtGMyEE2Ju5rmzKwRy2mARQ/TXFqdjWeElqtxhUq+A9wP6L
n52/mpzJ+ZxPm5B5BTd/PAMC0yZtYCVBiQdhaU/etgA3vkLkAVvY1lCTJqHJOdL0qingrTDztbdT
FKpdX1DDjmjic42pkMPzHTV1kg0DEz712XJjMtoGPyWpLw98+XgIlN1Dkl2kl7Hjs50eLayeUFL1
fznelb4VUnhcH+uWWK9enGXBd+s3O0UN8RTLLFd+k67Pt/4TsRPGubqb6Ef/3djLem5jTXAuujdA
9fzAgdeFibfjn1vUfpLicKxS8WG9hwdvWA5eWtfFlWuwZxfzWoF0Xtko6x5upV9tDF5NV9rZ8C88
7r7LEViDqm2HdWQ4L5cYYoctk+4C9E/BSAg43+erdeFy1l5fOw+5IkOgRmkXxCTfOZnAw3TSyOqa
T0cestx2uDS83kYoA/TjGMvPxPeIeXMbcpaWdxHMHfTnYtbfKo1Im1/1adTNJYkneoTjmyb+9zUo
ORuQ9ofaz1PLxvx81stqqGY3qD/aep9uZiDZr8ZXXBSbQf/j2AeSAJMbifuedi2w1haTtc7BpISX
1zXxdJ/xctL3W18KdYWa//cz9aWYTRjcoPrkX/4u+FVoOtLj6oL7/LtotX5JW6+A8gtg5nuDN7aZ
dlUyOXNm2O19SIRB7pzHEl4ISQ34MYgTu6dZ+D91E8EpUlbeQ7bNAck/h2a7s8Kpc56LNZPE8ImC
eFMStEV4kH5OZV3jvQbF5pbF+fkcKavaC5kiNFo0P8UETeUvrSHCSzUEXg6B0dbRRkkmhHOfUTTD
mhlktXAzeNQaEd7l5oI90WSAM6V31CYn0JT8LNKKFgfB4kFM4hTgQMH/R2ujzo4oMKIUh336Smhc
ZVPqtlQq4PvEaXRpEtA7lBQGDhr0mA6Si9TOCnG4xqzgTn21Y7N19PmCu/adH1Fcl9/SXpLuQPXU
RVMbTgei6j+AbY0WjrjIvQ3sbpGefiMOQTVhezWDdHx0+Dph2Aay96WoXm5OAbaxP0e8aBOUVn0i
OSNps5ekobMCcgGX2qY1qY9zJM4ptOZdGGU723mThi9GISpK7s99wQLCylrHCnuiDXxeIuwASoL+
GIG7CL8pDZlVk5B9x3Jeg5PvHRu71HlE4I7NM3cpHPZUzatQnqpspxYl8KZbE3b21t679HnAiIn5
/oHSh8UqHxS/wLaQlecNgG7mCwR4aq95tBmmBnNa2+vkqK48GugkUheVKPk5VFAinUOMTRL7pUM5
pSEqjiNJWsBg6sN+6OA1BDJ5uQZ66fCvh/AvAx2vHKQkbsFFlU7mEECHk6xDiJAbTyFXpMdxudv0
s8XhK91yYdocK4uS4gYoY++nZleql2DD3usEQf38Vv4A0Tj/BGWMNls9/ibDFYwOnLyxzkbC8cQV
EfgULL7xBHqAnZ32Qhbu0atP8NGs15YADRbVmxXAYA1LcfO3vqQmTNEaEoknJtCCLMg0ZrcBht0e
UuNqauDsJCMm7lLJRQAApfbL3YXR/knD4kQvg75PiaECFx6l3sZXPl3wv030aifpXJrVlJzwquE+
tzmvsdUQ8heTTmxs/f7wCstzUFSfdZGgifH8ti2h6bDn4Pwu6Iv/XBXFOOXKmIAgDGEox6g/iKj6
3HqA4DTbzRm2/2jbSKzzM+/52tTv3oxG4WYEmRhS6VyTcj18SaiJsMsreh2oUo//0sAUtucYx0i6
RhcCJqMJhjcyTbbzz9Q84AKJyGHpdGlahCU+5dDvo7BZ/32v+R2F2Wx8kgXMYGdIHPAud5h+qZ7u
1wCSUggQOYIhk+URNUo/NFGAt2a3dm3a6sE7IefrQK2GMrdIRNysDpkfJBqZ70t3OR/sc1/BwQWz
N5SeBB5wZ+a7jSIBmMgZdWskwJ0W/T6UAD+NnQto7Uy5Gzjbt2TfhktyAzt1AG0DU7IndpysESFJ
WKZra9wAIazGzUahp9FYd5FJtmJuQsYavD4QxPyzS4LJJxIhiVdbTSD8+OQMulw1gjdZ8ba3nz2R
JlvIwnMTiCKSsjQr5MdgKq6PNG+bZ3sfB+SnKYt0OwzGc+pxdvijZGlEe1oOZRYtPz+rO/ldVRaZ
aJj2YmLVZQQqor4I9Y4ZJGLINGAqz63uTHu3yje8EpmnI/UAZ7dPYuh5pkpWR/BmH+/crul+yQ2d
g/mAz+7wH0TdPG5Ws+zf9YZDuddFy20FhfADKrUjL+lncjeKzrIJNtRnco5T8VHwI8MfwqFITOLu
JuTj7U0a8VbIio4zks5EtFP/88qWpPaUUL7YXvitZMBp/Br3r4p7NJ/4kdWmVz/FG4nLldOtcIlG
+A7TEBcfhBFYQIsvhdGg7tT/dP/KF5nIRiqq693EI95JBnJocaa8F+AfDBZi3qid9AJi06+aVyGA
DAVjAXDs6Uj7AYIX/UqqRrodV4+uCPr/1J0NK3mRZ/pCCrb7NDfZZcZTaehq+WWTVWXOJrO5VSTw
1XGYYKFeBMpCsGH36HuxJDiFcQeu8R3FbP9g7YF76f6zCqerCTMVcd6YXJ2uWAQdueF0KJ3XdVBr
I/ET37bLCa3305PpK+4vYfZZBoy4OHfOkKG2rPylwp+sft8KF4fmwFe3XjhTsc8nYEQpXWJj6NjW
dfXiOvEjusjDtur/smDMuWvU21I28C7QQwvEMXpj8gPAwuEWxst7vEF0jelHqrGIdU+l6OBDxnd0
kXG81OxfxuKmZ7xZyiIINobT9CTCQRb9eCYEwFS8ApGaVNIDKoPiQmFh7x7lH1O5GTtBz2EqQZu+
wJOpSyqdjNTS0lfvxQuOa74YCw4PH71Z0nyVf6LCqg9gMgkPKvAU+pmI1hWQRzCtat45ALyb7/m0
0hsh6cFBxyXov1JjK6oSHuov1zXyXfXGPAz4hzKRh2/x0mDifeckIL0tD8XhwUcEGc2ZXOj1xV43
+nCdjS+LpUy2dkAwPmNcc9T9xNSOi7OkapKbAbN3rPIQ1UwQLZAZXmu7uOhL1qjKhiqoBOUEJ4yK
0ELr4MSAjNSjttQxzSBc50bAFhxH3hN5/zRqcwd43boenMA7THg0pHuFs7hZh1aqlUrNsc1msU56
dtuN8qFTyigmsOIhOlySeqDsipzD7Set2YV1ao4X4W4k9FuLAqZjtRsK1GngcG042+cP+pW3xAJi
eBVebFe3qijxWNdK2lCKeuXn9CcaAPu+xhweOPsf0yHDNaeTkgooLJDqPFF4PfZwXt9XNo9uUfaZ
W8tJx/fem0od6Iq//ILAA0dcdZUDIcpBZvNEkK2asMz/9u7TNmWNT8fP5RaZt1A1OmLF+ViqDFTu
kuOJmHLOV+OrCX6VDlC1HpGC9hRmoMXcdkej/49dyjaUqaue+nVOKSeSdG4GRImY+YY0yqM7CAKl
OUCwxgGfKhedxbK2cidHyf6QxUQOsXdu7Gef5KCTN3PGSDJ3ytvCT7eNGiNmMLnaybNQI3+cKnuu
1YVKGJ1dbOOnHGnwx+NraWYlZuV+7ejCC+DVZYWp6FuUn/pYnrjwOd6ic97nLVZq0h/aViMo81Cu
FsVz1m1x+CVHefY+SIeFk1zIPwLHfR4pMFXqqGhQII/fXYV53HOliComTDGbgTH2YsHr/YJND43C
Hc1UXAfesiTufKxng0nX/CbOR1kY0w9JgDfkqwRHHW/lp1dVHHtW3aUoW8F3khozj9pRVLTOvf8B
Ho6ZRGwxhNkCpHP/2Gbuv6tS+3qyxgHr6xIGXZauC6W6i8oPFG/R7ChraxRlpO0h0bF4aYgKJiJL
s0hT8inny8s5s1rdsof1qUEqtO0JtO7AWvlfnCfor/eutu4Fb5B0lv3QqO7eEcOLuTgnflkCXMFe
vDqxx+Z/sUYQiEC7Jh9Y21l4Kg9RMoz+Uk4fL3SdqlXcj1AaH28DMV1qDRMS2js5F+zRCe3xk4is
4Flqf6eh6NTq692crOcziTfOAMm5RM4sOnK8y00AGtoOM+G+nPAJcTmPnqbGD9MwGuw3y+kPHUDW
u06WYn5wyVXZg7oOyZcMfZ6v0hhbQFfbGqMKtKGHyAv+iYm65liPH07CMmEdnAkfuFPpIKCK4S6x
U2NrgQjyD29Orei43XfZqqyKiIuKP6MUGUofHHs6v3gS20Xqba2DbBzkUE7KPOM8qNKwd1dSgzHL
SLW1Q081fCok6uJLRZcdUhERhJ5XteN3NhFia5BWOf9MmLiG+aU2F6UQMxiSt/SLh+riRon/bjCh
WMv0hXF4M1way0L3xCBWwn7JDI/VfnRQ3f3PVSR/g+sqCUkIDBXBMfc8FhyeYS1TOx86nmxzJVLv
u3NVjPX9I6ptKAGGPQlNL15xsD/AACL3wQElDC2qAArp5tWzbnVAvHfPTx4uRUmX8vbOArOLoOA3
XVzH/QKZ/H+skD9R90Yvk5chIa3MmwPNwiM6Cw/XXP4gJDrrP6kb/QXqG5tgTehnkbEW7jruFt0Q
SzewdpkdZAVVwR/tqtj5+klyy0Ez2X2o7CNBzSSNqgxaNoNh/wMz4cf8sXlWG3ezrW4gNfSp/g7r
lrj8oIiAxjryFo29ZrHNiAblf8qs4lnO4mT/Op9i4vF1iIxSP+5zOeakAlegsI/59QwMDwyhxKy1
SNzYk6/sFfAghqnkkX2KDLNR9/jaPVFjh4UIDPQLP7c8Vv6fWKn2Sv+n3bJkENDztDgBDFQJ5VIk
XUKut9yDFqpZVgae9Sj3vfqHerYZHhK2gdOemh9ZiR7qnLtpu7ktkMQje06N7LgYkojz4Ovt07MC
+ErdPw5g9fUm83jdsUdpuIb+vehPMmn1R8QZdLOswUdNJs7p20FKBpHJEuf83H9k01lWKt/cWb5a
Z7TSYpybe/dSAQUeYfWm2TNCuSIDyjXb3GCZitKAr9cZVResXycZoArfbVhYv/LvFMZlScxxaBsr
iPlqaYs2UIfiK6IW1SOlJ2YyVRfiRh4z84t4QNZxY0g6P8bfc/rWm4j4a0zmvLRQ6Jb0NI8ekR7D
Sr8SptBWGo6pNP3EDoFV8aug+Moy4d/ZX0WPoy4pg7M/4yE3GGq19iWy1PARoS3H91FXz5LaFCTH
C5mYrUPjHlGJiE7CmGlVjqYyCvWnAmkhcTI3JeDr/cwMzUh5lQhvVzEdxN2vWLM2KkcT9k1dal/7
z0CDQw+717/92NNGKowKri4fu90PEYJ7jUi/EhBHUdPMPFFhP+QMBVKQtjWD2dkypwLB9LYZ+dcp
aLUUx0tf3R71GY0NJqFEg8i8ryx/ARhHfLYHWBl4DgYwV9oStubUIMmIQIbzrEnaNtlVWNQ8XnTh
hJGYiN8GOnAq/6+L9NeGL8iAfolEobxE59G+GNAhAOgftoujHjKZ6TDzLSMap7uHknm3ZpApf7Qc
+Yek+P06RWn6ZAh9UeeElMyg30jvsN5sdvl4MeZpuDcfb7RiZQ5QpIwJD1M8MRCwZzD/Bf35kkXU
PiflutzfSjhyLDy342MPRF78RwhKS+kuKSac1YQSZDsXVRfKZbaM7bJ7D3evx5vwTok033U7fmTS
Ybju67F4yCohm73qpj3GFPDI+kwoGPJF1ATvKMvQ5RSsTz/J3WpBDYJ3zflwEtU9uOb3rQDeEQMY
Bx5AtcccfBpob6mekC1IsRKYNJm/l1j4ianmUVpCDPfilNqJxc7/us0F73qA1LroMTX9en7Vdfwq
f1K/ZJowXnbNpfQK2Vilw4WX+eA9uq2vvW8IcGUbD7QNi34XagrZ+2NetPhIfG+BFyxkWSmK0qF8
jNbYlDcJ9Y9B6OokmnXXhDO6j6K0zpQ9X13XmndSVcVk+pRX7z6Ho5yCZJlQheM5UG//H2Ld6HW5
9aqWLiY/3ETa49c2Lt9Qb35yVkEGJJhdJSp41oa/YDByLh87A+PR9695EukCaXctFtrMLg/P0StS
eXv+U49lhjUdL0G4gVgsiskkyGlOtIxA7ytuGfnyxidcafHdXTwpG/kG1VzlEEdAT7Ty3QSUOOGe
Y0fhsj9n5QO3u5iBm4tHwtazQQZK6KXn8LODIQ+ixawR2xQ15fGF8Cz52Yf6rf7D6MJgAPPgyrK4
K+ZyeRYcosioRqCSjAG6cvXunEEwFgv2kTIdMzGa8xXoR0T84IuuJm4X8e7jOYWIuqFGT0Pa/rwf
k0TshSqXjctUbleZoZzZznPGu9MANEBJEvEQcscy+9oj+19XzS+BOhdO7M1qy3sk5aeheXSHdjM/
5PkNFcVCB0bUvXdz3D+Ed+a/t/gk11zqTAVZ+B7UlafGSVDODAVT0jQ+/kpx/Uh48z8Jp/0MTDhp
kruvGaYto+n4nGbK6YSPOKa2Vf0J6tb6clHuZ/0e1J3XUXGwD279zjlczukwixuJvQA+qLR9MCdI
diU2YNmwJeM/Shs0I7/Eij/oe1kg0lnMHTF9aCosJ6b2uNzrZ6H1n1adTXcg0Xv+N0aIEefLNyrr
hIhfbwWuAwpmWy8fZeQ6PKrqfLxi1Ce7PThD6qy7vs9b/0AAHAvqz2bLO7OhCylhkms8e+zlbCMD
Nq8x0TtZYiNaR6zqz9nDfANeWsy9d+8BqLXX4n3ScYb09tNr8VHKUUaJx2f303Bv8KRBlSO6KQ/o
HFDKUZrLES7T+OKTuFNW9kRKLDm3TJFSQkDNxvSfh6RqdExV2W/PAx0A0EPdqFKl1nOtNyEXlZeQ
bdA9WU28gynxHkA4AR2O+mDaBS8XqOp+kDBrWvYTS0PQLfwV5+wqofRcvsOCIQdp4AnMWAHaFEtX
3q2oDIuqWaLbFuz1Frx/cByVCgHQBRGMa44IuhpcJdgeJVri8objb2dmzYKoIquiXhOFOJWnOtrS
IVnpNgJrUniRzXE++OSIHnX30qlQ0tdWWqjwvzC66nU9ACmrekSqibCbvDqAYLtKVOkwH/eDWumi
xTGrWiXfArrpAw1PofQrdhrPzxuyXb0t7xpC4BSvYjcBCZr7mP2ECMFDqkoCRR6OJQGY3t2zv628
aNLkSji9dMxf/jjKpVSrNQQjPOtJMHcszsIFHAqIcu0xJKrkz5cJw8JgVjtkbG+33Fx2b9nkhTi0
DVQXMiTeuHYei0WfMYcsyZ2RUz6owzUTFEs+KWMPwdixWHk4n/mMj7jrjvweYkYx7/MfOsOUiCg4
LaeJrnhqzL7T3wcCW2+1JaevY5kNc0Yl6M6IrC6dymj9/8GEQJbBmTXp+BiuBCgnfHKBUNRs9m5E
RD3OEP6KlrQ3ixTzD7ki9KMeieECW0pOHzRPPwI5NsGaty5EcGQr7WlkAAyaKqoopa5jSpFwlIQb
Oi4Lgl4B+K3mmiWzBz+yeWxPJNwFI7UI6A+POuAnMazn59Rc0/t6F2CaKo63fnmsoMG49+yNoY9w
EaqBTcY49dFklfRMP1t/bh43J1jLYymbx3zCdCjed9N1E/9ZZG3MROu3hi5vnB7Ifj7hywpzuoUa
8scDMyDEYzzRyn2a6954AinudnoIFxb752VDM49NjXTcdhjjoRcGqkooDTbBQxJpOtOLoVFb8Atf
gqzhsVHCVLD60vGDsbp2vG21koHgP9V4dSsBJv16iHJBEoQIAsPd7gbXny7cIZRr7pbxgwDNtKyO
J3SAeUWm+HXJbZ/7TZ9Fcbp4yIxm2jTt1cCmvS7I1RqAE+TeMh/jnLVQz4OzLsxiWqjZX5acw/Y+
HxxiK5h82ExK0yisYODoWRVPNy+NlO9/eZqtpwoU5CWSWiQs+lv3l4bV5P/qS5Tg9E83asQS1O7z
80CyRs7RUu69Fihid4l9pM3jy9INrUHzO902CHvOV4I3E5n6IeY5AZ8evQR8A2Gys+iW7pljhzlg
GyAjecIeo7r5+B8XT2L9LF4gNMVQ4AqIDPHOrYXlxfBcdxCxmczTQSoYYR6snV7RTMXr36xT/FnN
KaphvD4kT6uF751xG/1a4+CHMstWbs+rozGdxAIyeVQyPFySVWd+hPD+jzPGxHPF0YS9Q5iO7keE
EKXiqDdxXqGEaTojWHx6JVFN9RfF8M+2R5YfgkJE8+p9Uv8A+9ko/pShaIPR+J078KqXGTpeORqL
m+Y2fWbx3KtneKERo1kOEkbvgJuCnCyqwG618g6p9lKi+7k0jqwXnG8G9WbtdkdFqjl8L+JRAOvg
U/WbmrPh6mT3rIP4NgSyv6CPGupugcTo4OXwk0Dblfh44qwlsDYARrn1kvhD4s6WPifp8Crlx4CH
aqQboirt0k7SaqsAoPwVX7sX/pOkKqmR4SJ8i+FnV5Mxmewz8J4NzLbmzlEUaTYznmOesPHKjvNy
d3sec4S0XTZqbheTDD0sW9Ly8bXT5q0qK273e0sFJSZLpQryD/RbF8CKJqKTvCsFwfa47icxG4y8
cKRfAp9WTmr2VPPKt/3z2yIfQ7yyU8d4nCBB5PkHx0yjqwrqz8wkwU6+DtwmyuS3aow+3qOYdSPx
+wSWnZDx+6C3QHb5DrwNTnpY4mRZlf8++DMGYiC+mZXeN5v4OIlG03EFibUA4vhXe5JPs7tIHwKN
DMu1j8mVZsXQ5h9emTVLsTkm64ffPi4oOWK7Ko+XG54BnHedxSN8lUDcfGBJm3D2F5U+fbTiSMuj
YSh7tBba7bh68eAeqfB+1LoTYuGxHSe9RZTfhg2at/fEKTAmb7YxRSVb8sOscR7OBdROTx1ssWO6
PfhYyS84FV+m+jNNF1SY8xv9CXt0oBreRX0SuJJpGPYFJkRs2sGVXCMCK3WtWXmrUyOjG5r//Dek
wOi/ZD6AdjLa+OJvtD+8NAdgQz2qN6oX9qYpSmzetnJmVhb7pLNZslw6K51eaREA8PP5HiLhYuvq
ESxz5YHzL4Ha1vzYqpJp6gfX8NsI4I2wZT2inJxsEpGqxLodAFKQudBhkeEX3XtIrvAxvO0cr7EI
LzvGEMDXwWbqf+4JDleuLjJxYQvSAKYG0VVoXVZSjRKFu7x2fm9zymfRBh4nrUlftXSQiyhzRCdQ
AzMmmevkDQvYdLoAtq4k+4upe7hTA+e1uP91s/vSNzeZEC6ucLFe+Z4qPk/ol7RYZUjn8xOFyDiN
KGqE5pNylycUNBPIdxq9H1FtQoyD/U8ZbBlTNbRruWax75c+WeN5krNDIw0i7a4w0AbNxpurYHGV
p7k/cp7Cub1KHnhy+1YRX5ajZUdlwJYd7nJzRkC7WPGojMexI8qyyQoK/Nlvir3HIMQwuzlfe3Vf
DSfEidt0wIQYBtjY98ElpiPszCaL75kBDYR4MbTNRklaS/AFf9Sx8G40OWF8jf3SIT8u4T6H8zhr
V+9nV66GZD63n5gKLEHd1a2eqH1ZQ2JPbTI9i5Fy5bNXSzIq06ezT9S2/1Jp99qSfbRdZD/7a7e3
ysSizP0yyDKDi3VIqrYKE56UNXakqO82dfWgfCkuoAExbV+fw0XdYkhvqsLcInQ72BlGJFwaO3p4
4w1zCtaqBT8xQ79N+VHd3GrmgbfmcJQHz0f4S6N4tsrIsfg5wpKoc5V5SLzhUt8hruAtX/YAOOBQ
gvTku1R9ukYNxgrjYLwq65rLaAbagK//oyRumPSlGkWsQnrredQPxEBrbJu+dLdpBQSS6rgQQkeS
iyCOd3ruk2h611eSesdTFRzb2Hy65O0Dnba3Cipdp7zYmCKOBHnTfracYrVhowErAP4NEK4EROu5
rq/4AaUUiLnJPySA2SHuLRVAAYL2A4KKGwHHNRdlxFrkpCVB/dH2naO4gE2g3/XHJeWV/M0Yjnbx
dqG84xOQIq5oEON1mc59GONWOjRQihjnVsFomfuViY7VX/wG/rakZ70E2uKwYIPNYeTedcdBb8m2
VRxitVKcPc6Jg6QaaxbhsGCw1nTl4pmcAPnRCjH8ki1mE3n8tYsqum+vYDE3v/Jk5+h7UxsQpxYs
6LTF60H5iutAOmJQ5xubB8RY6maBSCmexfoB1gRls+ietDHFUakDgF9sPb40USGS94RoT+mL7CKC
2TCV6ZNqIbF5F8DVcrCvM1c08EoK2ErgBDYuapZ2u70AxdBw2rpJlAlJXEaOB83xsZ4ozJRJUH2W
jU4SmQI7hzLJgXoO6N9EDwNQOfZl/9ZriBk1QXftJF6EZ1FGQFRAvPuN3lzdSNK2hhuKTNylx46t
x4Zj0oS/6JUwmN+ObJvzTOgDW2Ii5kRljcXC3JKRPy9cm/vDw/pM9X38QmWGaZ5NJ5y402jCwFSq
PF5meWXCBBh9pn+BEDQDJqmMKr0ifHyrroiotNEkTe24Ka2X0RJ15B9GX/tsDDIefs69ZzqXx52z
UKaFFohhCE5Hn6/EeoaR6eeXkciAqFe/uhbL9xMeKqWf7x9tocYar07JXIcQrS+XvLcHfVAHub6J
j7IEl8wdtbWErpJxo/aoVETapaI5egDHWFZJW8Y9g9L8IED+Yuyvcjd0HVGdtDaLzSld3DBXZ682
g947pwhBW1FhjkUQwjwIIQs4VGEJRhHTTHmxqIMhJnChSSt4rSOd1ZHraiGZu8KI6nTdRLwXLtZq
gcSTBFTjGjJJUqU5PpshxDrHo8ihV6a6afS+Sy4I7oSYD42EcwZT4IgcKADZaK2BIDzIyktsVxkT
TIA0IYXt15nUgrq3gAltwfB4K9/wCZPilk67ie5guIbldU1BMP+fDYjQgD2XRETzuwEWwyBPzZfU
xhPP7f2qnc0RK7zIKBbEmoxwRuuHlXM2WFCGT0DbHDwx3KqGxVNnL/0Jkd86ZK2d1Q5GuFeHCjfG
HhpXMZZkD75Ef5wDrxP3PyD2qDbX8K2328qnqhifbBN33I3/Vb4VFAp0q8KpTK3206ghT7kJ1MHf
IVHsaBuVF7HN72L65Mcs79Xr0OwrIvWXLaVYwxWSdIXSYYgDYtXdMDdwJJvCW08zh5EDgVOV/iTW
c3WVtG4c+A2Ovi2KpD2ottEjDq184VVavTviMBvXJA6SIMEQjhjs0qonINxa0+l6DbMhbVvU1IIP
a+yznyqS26MfocvwQI55YPxCgiPO1m9gMmvL0kvffklrsaW7GMFDUdxdDoVnKv3DICqRpEF69TNL
b0LN1kKuFClwXsV+QenrBea6k9WaDDgzsxdDJKXo1UwK+RzpV+TdTuMtU6fuoYT5br3tTkiM++Cb
1jTMimqsRT6x9LeQf6DpRfeyd2FjrJWTg5fUDjlDcP3D377MFwiiF0GGRtUDHW7fSkRfUYVYf6ng
FLr2oKmH8pnKLBZGMUjL7DdLn+Gri2AQo6oTt7dhHK3jODNhCXpcgS0BmEtSt+FwGztv6iwL72Db
J3C4Cm1jGQtZMkK42Zh5Wn4pzuxmyrk5YN1MedKsC+G0/OvumHt+Q7nNtuN3nOPpyxKSX/9xCVk2
coi8X7TZ7TWyZI+w7qqiDXqBoCZBmJ8zCcy/RlvJyclzzKiYGgTDjxSvUS5VfFXeVOKwhOXqZjvH
qozStBO3hjxHh4O54Xn8Wl/IBZsJJCV3wo2TmlOoAPwEBBhgRYmuEwPpT5aNYI8Gvwt0joVSaf3U
y+R8c8Rgy++Y4eeOYzuzrcB2lDM8GnRduP0Li+6qJsmp0jwTlZGh+7LXjOO1iieQSyUOaE2XCU7P
n4K3Ga4vt04lWZ/7lH1RkYAEM/p30LeOdbaNvk+WqizJd0v9EeJJ/pJ4cTg4DevJCuJRgkJ5THul
6GEZm62Np79okncrHbJsQyCkMy0Ucu6WIpt/ZERbGdbSrdKQXdvwnabGlVto+Eh0mayTJCLaOacR
+u9lyRRXRvpmgPlgLtD28O6w4Ig4xln95bWnm/pzYn+llRwaomqpO6P1N2AFQxjhiZlk3LT/+YJ7
6r+saAOYW4eOUn3UN6Q2KCYI0b4oYcvSZ21vMekARfwz9cmsYQgsC6Q4fDmRFF1PvaVE2OP8oxpH
Qtrrs0MC4I3NdqQw1RIQv12yIDMaYsCNnhtOR7CiLjj6hZAhniE0loEqKKduGvgYQfdpZm5UAxk5
23Vg5V6MwH2GEwOgwjc2VWJMSAMiSKyOcJAG+kt40rRei18Mrmz8TfRbh9gaOrpekYldznXB93Iu
cP76rXEHr0mkOjaG7G0P+cBq//etD6Tlg0S9RDl2VVc3clG6OCpVLQX0ELDc7nUU8ONFsCdxxbbZ
AjnEG1d+WIhrerO84P9mJtEmV+vy5s9AU5CNgQcdItmjzBShmZnZjrSlB0qiESFyyPPWB1HSaxuA
CX2j6YFP3IH/5jiK3isIln3iUgc+3bRWaRZEIrlvnMQm8OLULt1k2AYgx/kdawsCgkt6OrXRkbUf
kWVQeJzLxh6QoDxibGjfFKz1K/aKLp7muT8zxl2LMxupmXCsPP1Z9Qn7NuMD633DIwCsfBmwBGGQ
S3Opslk9T8l5x4SNc4Wrb8uBrJO57UKfegiFEjsIDgk7K8wczPye+zIWDf9EI7CcClmeG5HCMMdW
alhNRSPEURzEIfWvb+S43ITdfbzxfmCYSgKUD/7GhUJtO6vCoiFbN979a2U4lFBQWh9IrijbXh0y
EbmnzlgSutScT2sjqI2yDdHfOVpufejoeswKToHHpaXAgQbc/VDs3iC8p7/3NV88IvdsfPLFRke6
6IbFIFFEB9qDFPVAy0UbO/Qw6XbE8rzLKqM0/b5rxtNX0av39170SSMtVW7dpevWMpBPH9P00RrW
WXlTDFssg6jZwulmeuTqMHUMuMNlPxpO5qljGDpob+nojgx3UwloxceJB7JCYkE1Fre3gfsTxU8g
nDASV9+LKbD3iWV9xegdCAG6MVT5bJSdN4uwW9CPHPgK/7oCLa8K0gShBxvUJxVBoTKnfLKCJPU9
KaYhoT4u8pznzuKE8j+Dh/v66H9S/KijKyffHQi1D42JVGhZOtauda2cF5Dm/bnvrPSNiDqx1CBD
3HJ/qFZI3zXxHOHrIuGemfK3ZxaK0Tn51bmjDHI2qQFVFZHd3lcZptMcOIefFH68ss13a5h3X6+h
zwWKfTnI8PGcl68FLxB9vhSbSmM9hB2sNIZDJcuQI3iJFB/DoBLe1j7+bkv/jI/TOrtkg4QwXOW3
j1GrJ2GI7cGXNRKOuEnSWsV/vqoT9RyM1wtziJ3xs/z2GINGevStsKerIr5SgS4odCmS3/QZmhXM
gkcxqrtUvqWAQ1rLhHLkbT1b45MNxaSTduBx6ExrDjIml17eBDkaW7uy1ZEB6ByFQaOK7Idy4ALL
dZ8AKv2L262HNRhlsCeRLK5IyrCUTI/MxyvlXjP8zM0zOIH0ocLZoGi/zAicvEqHhtwyhQPIzULs
arUdC29FsKFSWzKcGRqneDeTDF0XoKfkJLNQ1v7AhXihZSHl5j4QEvHnCbgXWYWDVyunvCMvb7BT
2ItfHEUE+Fc+aWt8RGje0pvsrnvPbo9EtAIke9YTwe9tlmYI2RMkLKDzHS1swpq9sg67+nfgqC59
tdBeXzsm+J8VDVoiWX2XPR46Ke5OR/OV5iPwHI0GGudT5v9pWFD6HmKV0OiSlsAEhwrcTQG3xUCa
Z/8Rpz0gXECHV7Ecks8ElY/avl95PYTJ4i3FXH8ekhjG9RuF0G4YKK9qpAkSoRRMr61Q08iP4wCS
jtMh9WGKTrOsWeGK6Mq/hTwGPr1kWaYtTg/KNQn3VucyezGekKpClFl0yUu+JFJmeapt7XFmwYUS
FZzGRMCFXEcHOipO91rOJpHpyyhVjDNZBkD6gYMU9oKaBLP05Q96EyK/MQTw8LMLctsYKPHsZK2J
WWfpPOvSwp4qwRmO8aufICulonM+1zjIVvH3Rv8y0VT5MleA1y2Gfqh+/aUPTWpobu4GeAfbpVxY
1Tx4LiXrw/hkIKCtWml5odmqVbPaJXqJnyuwHDpuFwR814SYRDUZFRgNkJRR0lbUmr86RqYwf8RB
bT2S7d2QX5UFVzxrcIhKHrRkAFLQno+gHsv1gS+iY6Tnqwxndl3xuNoCm8MsjUOkXAe8yqdGbmHN
I428EobvmxOvX1mft3vxmZFu9usXRv4yxjrunjUdGv+8m4gD3bFBQyYLEVwrvghK2pB6MY2GxvYI
6wVwoKao6s3hc+R+YNcotio9b7ZktH3lwhlxoOi3dX0Mx2hnIBIvaIP3Sfjm/N3gQrBwnolLK+uw
V0xYhDJN5YvaNT/V6bfaMFlhHyOGU0wg6sHIg7hO9yd4k+BLUKTtv/Vm7U88B/egiK0Zdr9sdr05
w7jIPATjJCxBa/3kbXnSJuKt8KNUlKkMKI2287A3NEUD1s3slrGTUMYuJuffT+J4pTyKIMxoIsNr
oJxOniqALnkZmowXvlFJj7HR2IPl1G6fHlo3oLTH1rxniCQTp8eXQFcP2r1g7h+uUOoq+emaavD0
/LtxJWKOgxb06nFvxns2V0y8yaxcGiDCWWmCdrLAmhc9kNQgiXTtsfPkNmzq30V45k5QM0uzb7IR
SK7LdREc/TC50Iw1O79LrxEls+H8anY4TPnPXc0gVeGnK6YY0+bD35V8HHOdjDO1YdDAVfF7kjf6
l+Pz6wcnPnFwhbGv5sSD+pmaF+16b38Z7VX2KQ1OXf0uBmfUbNgEoYQTbgLMMbAchKpcp7IhmEcb
+XZd0F0UZRtMdyc01s2m2zjueWC8bpsnA5vVNGouCb8jKgtK33nD3GYKstwMvCt75eOA7o3cZu9L
FCd5K4jxADBL/g5sZXzyZZqq6dCnC53Q9rqxLukChEMO29hsWXpXRiZqjjM8kWOfln8KvJZauzEq
wbRfb9AzwVSbnOg+dPsJmq/kzSqC0+HdNYqOWEtYm8qHB27vXoHvhKL4XPVMzUsdYB2nfvOwQJGH
i2kVJVtQIxpCMJhC1LSpy+LSpi1iacXiyYkc0z1fWkCSHUapYCGa2gNY0Xm5KEQu31QA/xKdd/Ix
KRBp6eQ7PGcB5pla8GuCoSMMmiXsgupOKotcdIpOXvO725+kNTuuKlMSB3Ows5qJiOhUEcrm7O+V
BgN3PgFweI+mgUfwHAYACM3mtzDmWi1QVJrF2Hom6B/HCEuTQ/6Y+E/216YvO2eTt6Xw2WYUeshk
fhXLIA725oIn2jB0HDiO255xFlU51GXLdDnet0EzmNXlZZshwFlhB16BmMsR3G30pE+Bzk+4qQw3
2h4xJJEK6mywtHaJzGtmRNarJJ2nYKY7I03pXgQKGiBtek+00RmRdf53sh7Rb7uuFPg0ZEzhbkNP
hJ8AZAAe8Yp8hthcodP188GweovRLu3OgLGcNnqjfN2P6QOx+yg4EogoZpowhalBqOorR6pj0gkU
/DcBeLTSDLK+E5mMeKdb0oCFPuZgvVuu5tOhElHEoHY1tPCcFhDJ5Xa9nSJIm3/zd3ZoSR6FVDs/
xoOi2jGZ5fR8cp2qAn8ODylZeTmVIwuOyO1aDf8ulpZ+SzKW2SDsZJ9Z0OJmLtAJIPEeEu3oeqhd
w/o5v8R/7m/kqASDlpOOlJpe1DWDO8FzS+NtEW3+Dsw8U9pEdnqUzMLmjjPJvSN2Cts/qa8V8FgU
UFEiYKFNZ7DuccCQZssihxgsDsq+obBKbiPZDzMHei0YW0pO4H0THrxzGK6oR+TK1Hfk0o7WLm6/
guI3ZV5LEdMwxvFpcLE5YSiC9wybJGjOIPWZKSYFPMzpji1dq5bNuAARUzMAa3n4+j8BjYfjUymD
CKAa9hEnBxhRmc0nmQIfraiLyrGbz9p/wYKlIE7BGQtnEgAByvM3lxazlIAR2Ol/sd7y0lz9gb/c
qbjCZjqWeMXiFFpXqj9wnu23BbDnep/2Wk76MLWU6gXo2ifeJ70vXUEk62PbhH+1Kcus8L3p8Qf6
sOGxSaacJU9g4XdmGWBBQzqbxlJZFzC2Exk/Y1nhGWnDkW6ftpyd0pdUmG2suX9/zINGmirNLhTF
DF9Qc0lxQ4+DlDUwmv9DUMl6tvC8I4S+3EHRxFLNwl+yYpkP1gHpm+Z5D+Yas3ViEZr+TznTUaWn
8CAGt50gNpvA0ekTMsHUi6y5N7+/1AXejUNXogwgLj3Frgri5AwLtfFYw1La0SigZbaQ1AmCXCOr
nJ1RHc4HT5iHFTARbxek/KtsgA8XqM8+UshPSFOaFn/FBp5Ak+1gyg2c23WD57R7kIIMmKlYqVOp
o2nVES1m90PwduEK1dNbxMXiuigP2jo5QOXJXzR8jK/Uwi7ODa+dXT3v+1Tyi8n2+qkxO/H3wfpu
wRcg2WrcmHrbRH+HQROrwd0goiF+2NHQbHmbVCwCikKZ0IZ2iVhtNEUz70AN8RU/9Ea88fUxioOD
T+QaM6XLDl8uC3aqB0xPlNxCCYJMq6VsmV2+ZE8MlwHyRcnGD7TQdH5URoAk8j17i8412ZGV5JEC
77tlDmM+knEuisE7LchwW5x5eGaSgwZ5HMvGrCG9A0hi8MxXIMmuJ60gatIwfR5R2esVP0SMVuG9
MJDjnFalMDcAaKuAeMhDLr7XvKLM+8k0s5svET7nX+zIT4QDULCM1UvNVg6s9ZgwC5bUg7tq5Gmh
nB2MsQDCZAAFHLmWYjBTt3sIOUTH/AswDn5NVdq9NMeycAvSaR/EI/4GR837Ug8Al5vzagVid1K+
z0Nkvyx4NqnmkQ1C9Z+8U1zEqz6n54h1sTDEgcSKEkZWa5h54aTCu56p4bHGQ7gHldBem2KWdn6v
dMMVIb+ga716/8HnrV4Z+nwTXpNHk9sNomwbYA8OEWFyf2KIUn6GwlIMc4SaY65KDon6kXKxUiQl
3aUo8H0qtnRmfef4pd0y4V7zRQU05iyLAu8cU2nTMR/EQ4JLcF9jAA8tNvTKnhpSgzsz+KeodP5D
Am1+KzhMszESdEeY2189+bSGSYUBr6ggq1PQ9cFOx8af0lKPn9rQVudg8by9EsnjrYr5bcec3zva
ttyEWYVTz2Z7GB+UXtF7Xctn2uNoB1esPdaLN2npxzTSfBbNsp6hgxJmVnRAugCMyaL6ofTU1bXU
URx96qppgMHsFmTNNEYl9cmc/S//ZnliqR23jDcOxW+P30pJg0ROMW1jcW1wBZ9la75/vKCV4dqM
qu8jEvVvY5vVDgMSRbba2bniQ8Vp/GHdLHFhmt/naLtfjIgzc3wtrv7wg7CBSu9r315Z0eW/CNy4
RASYZOWJLiz1A2FDOfB+cTjNZwZ1/yp95tTfKFGEosv3jPxEkqeFZNzBNYFXkfw7/7o24xC5p8Yf
j6Xun+/0J+cZVG/PqpQpS+1dJQr+sAKnhxr/z0CrthMO8jmz/XL90fdValTvPre/2ueqhezI/TTd
YJuQgVK+xDEPTOgIn+tyM7O+CVd6B7V58oE+pca5Y8cO9bzourqH+mIm9fC6SoSOOvHBOUDBOJvB
NxHY3zyV7lKT/seX+HnYcKyVkbJhnjnVa6aDNEdd2xlku7HT1IR6r+mHJaSdOGXw3T2jRz7Cjx9i
pIXYuGmb0Sj7TPInX9Zm6yDvui3PvUpV2BujjvPopW8sVPguFjayX+XrSVOMJGWWQweQu3jU2V5I
keYkJ4heTiVahsFTQLANTlHY/b+vL2CQj5PMMFjRHTyIoSnDSfOfB9o/6vSvgmvt7+k8fYRusgoB
LQyB6WbuRKHV8sn9bNaKnIZsQf7tSfY0LL3kLLeRkdlfX6Nzi7edrKLIr4OlEeiLPaBgYCnSC216
f0m3FjmJmx1eQWKBxW5tcND5ULHFiOXzDHJwK3bAe93lq/PxOa1EkUVUko3Qjv3JPJLTVxl/GqQd
5z0L0fqekGq7URQrBF5nmAQMbvaGe9RcSP6VQwvMOAesO5K99hdveHCbGBLOguMXgbaYYJoXj8hW
qAa9GBEpDKTSI8m2iudI8iVlosYeeq83U64crSacBlA7iifHXT3OBuW7/Nbkkg+nN1Jcj34oZQa7
+jvN7aerDxClAnwfqaZU/8+Z5ZaK0d+khbhYFfsSUYaJEmFRMsjK3lugRu9oamXIUYzMSuQlYEZo
t2/zjHoVds4SoiYe8F3cVv2SIdndlA9syJbA/bvZifGCUJvhfeuO8CYwDsQHp5IqZY1rXvt4/kLK
vGdEU2u8yiPfiSZXEwzkqtOATnkHPLHYTcdrMj7hh7mop2t7H2Mk3+IrRGvuAAawky98kDAJFevs
WxhV8x/NEVSN5dKZSFOpB1PNGBrO+9m0vXOJMbfoHucu+ejdIaWdbaFH7jU6IFNRK6yU9HTZOEbU
3JQoftVkF7M3i+WdR8PqnDrMZ3pk/EJ2/duzp4AHPtefDq+Oyp0byOL81E+j4Xw8ngeMMRzwbqkg
9OqU/Q7Uj1+dm17Yu1/nh7lKfuGJvA3CFqzvOp1EfEXuhbkT2jHkpVoRq1RjPqkgrzh1tRAyC1Hp
bm70TZUVqraNzBofvG21/uT9jQSSQgI3aMubt6BA40M5PCDwRPIe2eP4grRCtXQvqGrwNbuHMtMO
esAwfcNBcRSrfFhAozbCA4nkD91i6TpuuuL7OXvogU6rr8km1ncs9NJx031OHvd5ZIUQT6qe3ieT
5354MQNfmSp28NUY6kuePnc8UMLiDCDTIacEMYhK38/gn2/6yv+Zw4HvDxWRGX0DGhTIqv3cndsF
M3wN29nGePs/kU0JFPNbkiSHx2qORS1oMUeyHNxWwUDej5nYOVGpeLREbsSxNYwCxFm02ekQSJPE
EL5F/vbtFZmvTzhJOIRntpEvHhdODDSrSGC6IgwX+aUZAwTfzxcneAaMQiG9bWz5Sbs6uS9hGjni
3ENRxLIHxR7/0nkafuZFh5/c4n0O9gRIM+w2q4XYX6N1K4guH/xAPslFy1qD2IhfBFTV8PQ8f+pr
EiAkVIaDeKHbt1hKWBa4toa7oEcUfWdp9N6x4AinRSRatVJ5H9+O3sQUhE9mg4aLFlYEYRTDrLtl
Xvu45qODpWJlGVYW+Z1ZI5zEV6iHyrcJ3sdcQXbs/NpDj+isG9D+3BnnKxkr6og4mv9O1CljO4MT
R4pdTtFd77WFgpKfi6CVUsLGy5EBFBBYZL3HFXuIYZ0U2Vr01A0/VCL49V7qwo0YCRQCKW5rfcdm
ma2c42Mydr2n8FqPllKo9wn63/+ex+DAhNsQBAn62TiQ8WK22C9Nu0l6psUG6UAUllJCuusWYHrS
i2RMNcBzCyrDjQQQ4N3HxFDtZiO5rCv5+/Gmt39pzdHxzKYVQFVPtklIczGYB/ZU9PK9nsdL/xf1
F18+6J6dWbiXLi5tCReshFUGhmyhfBB/HsH+hskXCA9Z/HUxgFasOOlci7y136Cm1PsIIdkyD9Cj
At00XSntmGviN+3fUioBojewkVwP6JElcrGCPXnvlfSxxh5fgO31xJrDPGquR7VFkhmdutPF5X2/
r/ou5xqiFsVCmTkJPJh/O+IPSwbL85czRoVD23Q+2FLIj5bMtn6755eQgVCsH5KwR2BFAGMYoJFR
KY9+qq2uxN+6ktIY657KyS6NTg4SpGMxXeNfrTwbO7rce1lh+ZNHyuQ83yBr6Me/iDZBzhoeY4m5
psDYfX0UFuhfEJ/Cxf8As/tvjARhX5K/ip1QegIW924qfFnto1jSA1ZUfywOhYKYjbmnMzQQfh1T
knp2uulD4SXqphPyVUFUcP6SwqQsbpg3Sb+Sw8I6Ow2UsylB7O390bfPeIKVzD8VGhKuFeGeLSv9
sjvj5oqqEkUeNAIY4Lqs+zaCzrCEMASwfIH6eTXZno1FHDDtuxN3rKMvgTqKjcMZU9BFAwXU2rq+
jCdCVTfb9zu7jA3w2i9GWLQju2oHNd8mqJ5xXFf1eF8p04i4gUnABwtdT7D96oupLjwr81D77GDL
j8QuhNqPImWG1XXWMZWi5L2kEIK/AFpyVLZJpZ8Y/aHiYTJPsRAsCVkf28uyiibJhTTpyhuADSXQ
YUBZU/qjORnMPAyblnjkmq4H/YfGOf5uZP4KQjvqpMTIuzni9Qs1YyxFt0TioP7De4hB0B4KdhJE
ir4Cq21L7hiElXU9++g0d4Xmia+NAvS6i2V0/gkERwKsNKhd+Tw/eziegjwf2SeFPfESaeRcB1xI
PG/XyLRKMLvlK7tK6QppsrtZx4JSGu/Gads1Mk1Z9WejivPJh+sesKT6IKM8TY3XWw8Z2yfDl1Mw
zhHx2+gO042J/TmceDVRPWyJi5J3MlaNLAxRe8UueLcktNCShVSO/DFpDESDtvbLpNt3oHYxt+i/
IPApXoNkZmbwFHi3PVOe1acwSVFokxKpqMJHiXuNSSFmYmX+E3NzukaN2WKZ5ToKuAE9CTMKkB2l
psfDQUs7c/eZTFJ7Oq/d57PsRi58r6p+HYnKBrXdg6fkne3dFl7yNY4+N72mwhQieTqen6fM2w4n
Oax8shluuVontRRjO1YF8qmKEHMEnHUC0Lr2IhPVuQoR6qmOar0TxOjbxousIfq1hY6paZGYs0Ke
WnirCBmZp7J1Cohgidtdu7gsVSKWBGCTtkpB7hfXoPadlTpH28Zc6aXKDmm9XP2TI37JNQ5on5H7
nQsH5HKLNE/C0ih8IPV/wHV9g3Zk0lGaMbBD8244RU0Dh8YMuyyhBRBrwIPYNIj09o7iYbTIDxCf
8VnNFuW/YpPqEx6L4fNzNwzhrYmwjK4MgraeFuKzeGw6jJwa2zPV+jHWAQqNrsqHxz1YfWnde/Sq
GeVnyoEIIAbY0b7jJ5fZLw/FZsw8kO/9thogZlGdoFnFxftYik5HnwnSxMDaAyGmz3gKDg/1wszS
WMjBYgJM35keufXWgYfrEB9xBuuSpgS4lfIEx6ASU1bmb2nfOrX5BYKQvniKqW6WsF0oFwJJ2Iv1
EXT8gVLNHdqTknscYupsR5i4VqYxCOISnTHeHmjjE7+6T8baLAOwvo78lRxzvpyrNTnp+KenOSlv
ieULZ9+oHa0WFO+qYSNRn5hW2lishp27r654QW0XrW3gEAOpR+UaJLM3T7PxxB6PyEp1+hsTScXi
bM7wgxs01Cc00ugmjnK/KKd83r9mQQZb/KGmtM4Of7i3rGNzQi/RoU1SzLSBbn43CFKZwgBo1TR0
lqBbcK2pMTlGJeznIqeWU61v+XzRrtd0zqMYhoQ2G6uNB9ltTrq2Vf0NELHd66T/eTz4j940HSVc
OPx/vsu8pRDnPOmXVjuf+3srJbdiZjHq8Feh9VQa67ACDqG0IRAwrKb4d5EdnBK3wmhJQr65UTki
6NyiHiP6zZHIJ4X6tW+A/DxhVQsApmwCLj9ftHHKksCmphESW4DCrXAvt5c7LySk1QNBbbIB2IkO
g/w+ZpsBGoFQULhvDORYvbDzOkb4wm5LUrMGuyoLBPDgEdoh542PF+ZqphHK1pb2HFL9xrIcjpMO
QxanaHmHs6e++Dx7EkEhQjg/Bd7Zo6bf4Ura7uYghY5UeolHlDU8RJExKBe6V89yod8zosCN1avk
xDSobPj/wqtAdjcPuU8dgXFeLecTkSLP3dtBytlL7kiYbF5jRwO8pg69jZYuQTxr2CfLS6B7Hpoy
W5xevOqOdcleJFhAcMa8XcQ3gpw0oixbYksHbJLpw8DIh/R8DgbS96xl7rgUL8hVL268ZSzlwKuM
0tiPaMRXOnbstk4hwPQCP+8fxfdKZsGnDsV6babTm2UmabsLsBKYCWxGNQ55fA6idcWokv5FEJhj
Tp43GGhqkUgobVtzz8gFdbWlcuhnZUtc2uXSdp+ylFGTaAye7CVaD5u+gUBuFeeUV//BhZey6bya
Mpwh/UUpyVL3O9uEbhNXti6Uo7XZb4to/flDcEWCC090RzGbIcDtCaihfegQSQNgVY531cLueJGT
Ux6BWRYaDDy9WUvgi8FCKTIhLH9wsJF3LrsydKmW8iO9WHld2rxAtGgfTN/u+lz+CWDK3SnS0zSl
ijnvXXiK7sXozGRSxjV7hAF/KPA3R3VcjOuRF6tcUdOjtDxePOtolpYQz2oRO4XLz59StBYwGZwU
EWIvmP4bTYwl5QKAUb0AHjv+5rtIc4UUUQTJPdddAjol4xs+2WM3IPPErgJcjrxo/4uzY7ymwgki
bH0/GXUndxytEo4om9oZxUhntuENYRlyLSb11qKv3dEEDiBcweGtYw3da0F9khpSuu8wMh9sddJQ
Nn5NC8nXP38bvxy0D1yvOgm4e63HIBXWLMk/8+Hxog1Nfvh0DhI5A/kCU3HdKAm4dgFLLw0HWqJm
PHUSuzRpnNBIgywaF2hDXHYnbDQL9QXNdJUSmd6KyzI0XIm6wRkoljMxYeK84WwrLGOCrnpi/0ht
hwg4zx8mRluRyRkGlIbMlKUX5/bM1MrTSQ1MgUZ7JUUD4851sBPvwGRdzA658S7qUVMz7EMCKL7w
2Pznx1B79Kak7cGqIuiqzHLFkV4cPlgQAqigfjV4sark0VBAobMJOi7V0k7w/WvaTbBh6nmZeQ1U
jwqnOp6dTgxPubQosAsrx3XUIc5ObmSXGs44AcdJOMlCx0E1UHzM8OY4pqFpTlDHZqyBOFunxHR5
9iwSZ2RYfmc3QmLOTjZ7mmlZCJnWOpQRFcn32aJG8LPHPOvXw5db8ceECGsbSdbf6sXkZGCcdxdH
oCdCU+PwDzSeGijHWvaO+WEFpGL6Y5lNz/RZtM8UgkJhCpphVLTEH3O/HY/EGQz3vh57DNbJCI3p
UQhmkyykzO6FhmpmGgvMLRSEftr4XimzhbxrhD961FSMxvfcqIzJn4EOblyex/s0/K75TjRCiusX
TXOGw+GIEAE560BmikAU+gyUcIHo8W/z+hi9VcysagIz2V+8bQNJRDq93AyykBt3qtgP9o59gO8+
RNhPv+APfIQftfD4QIzvcbC7OADQtNhC0l6UxixyLdkOJBMVQI4cO1pcdlb956it8L6zdSP1QfJY
H5sKKrgrlmkSau0paki/zzsst6foTdowO2qG64HHE5GJGFWdfgJBVoaE6dfiG2X9yz0rdQoNzgTY
Pzgo6HzROc/MQC+HtaAPZPeDAJUYkD5d9yANzgzWS66ig4P5dqiAuTN5FwrQ1qCDtFcWN8nmv03Z
KCtIc2ORTJmmeMGiRfpBWtPlxLIYt4RNDFSpHF2jPgzdZFOITUzu5qYyKye0NgHk6IeoCWE6bBls
O4J7gROdIaUzLYYMMhnUeTDT6IIBAMz0CBO2jWuIjJL9Ei68A7caETLwCT24vo2gEAmQ/91rjeZm
X6OO823vAac+vOt1zHsvOe8OLrczLHUZFzL3B6RcjIHtd8thK8XtXaxJx6if1y4dXoObKeUo9+ME
utdVUexE9C126WYY/dsc416I9uU6ZEnJ8OxFaRIrOonSwkkO2g0UGCk+XxLIWRs7KSZRdaOkaYw1
MkTZ2269JEpHE8KH2LdjP+IAzzCAA//FywgQvniJql0igItp/BcH6Q35Yji0derR8RY/8UKILDFh
X+JUYuBsqO+SllttHgJArgnyzvaEOc7RNGBCmhXkYqYJnE/h09+wPVgcCcUg8IiyAQ70Ey1FqcTm
R0gM8zMP/mORkZ7dYCJTJql+4YCfDZXHLslyl8p88VaWo5a2qIKCB23buxJcRx73+ItShYIAzPF4
qJiJ1l7yw2VJdhBsj8xUyZpnLg0PLpAoXbYPUybhhl7aqKbvMFlP5ZhFfJ4C6a2GEmYzCbOoLR/e
AJWU2l8seyHSvBuqCTbVne6B9bzhgu4kL6YsneGbpoMnct3Wprf2A9owhbeNC3yPx0vkZ1es0B7y
taEHAwjKtKe1WDB7B10co54xMmLBMuzuSC8vwvkX/D8KlPzHOtDwGURZTODEwpyB1mGdkqfm0nZm
rbQ4cKdrXENhETMDDu06LSymdFxKwcOsCZ+92G+X/YFCYeaYL95yVuIJq+VVViCHTP6i9TFP0T8M
WLu3oAuA89TChcEt1ahQ5d+qhj3FIQO6wmVFS0JKSfIXc1OUe9FtuROFE0d/3hLQnXO2yxB4TNSo
kQEVws4V/oq000P19ewVSN87iO2kZaPEBD8/A4uEyKcJBJw8uoUymZMiCl6fhXsG3weM2OyNJnzL
8NMirsJ/tyGLZzwKPiYMeGewwSaMm/keJ2KKRFdjlVxDGR6HthsxRHjD8iBnr6zKwn948UoSo4ib
6Iw5V+PnzuuoIMpzDi8ox2VOnn30Bg2QX53LYPNOvll0MQdFkgVrW2V2VpzBwY7VyEP8fnYgyGqn
7Qjv0yh5opXt0Y1a4rNMIndh4HSs4DQejJITBIMftDZf2r+jCWA63DF8X3FDVy+5sTd9wibOxtgo
IBwmMkJOCsI+FpQk+l1C4JrJKl776ZVfj7Dv3l0eDXWM9AaYKt3n0jzQZzXRzvcuyfrlEhuXtBe3
FZQNoUPFgVW5qQB6ZB1W9jRz5zz6Ch6a6V816BEQcsNyhv/bOvKHSVZmLH3N36UjJ78ZBAMwFaHH
1i3Ii5iMWsTK5vOBaJZxZG4ZsS2wtiv48yr52M3fkoKdXnjjmey4dJJupCXgdR/Ab4XP1Z3ZCSxq
Fb0WaoQtTs11QqDrDfq52AiriGzx0fgJax4hK5BVWe46g3x4GVsR1SL/I/oZubk64ygu9bFiuvLe
Cb21IVBk65A0AgeQo8q52csKvgaAEhGnXLy296EA1CN1abNAaG7GELhFfbWdgGbb0/7gpr1BobH0
hfW8/3RLa4XL5tTCeJnBbihhdtEzZucB58l7VesurDHGfb+ctiX5pijHMzNQkprZL2khStFfaP6V
XeJ0bdZynEkE6O9cwxN/+8u2F4Tu84BpIKebF6tTXUtq8+aV3fi7eVl16a0HYm8wSu/3eCswejNz
5ZIn8VHJK9VCDNoMY0L/etTe3D3quSJ56hNeAiflVNlhbzvHV4wAKgahJq2jmO2FeRvYNrSZ7DqG
SOt5vnfitOSu2h87aOrs3eJZOBoSj381i646Ki145PlIjpATK8S1SpT+jyIdGNz8BotnQcxBdMco
HkmozYl9FMiJnjhHZ/ZQnj6VEgjsHbqDF4o9NwEZbcsTfmk0hAJ3zxBnmU42NiMee9hsQxBMJA6H
OKfsNpV1rqgOSWy6PThbF4Uh3UgIHPWKyp3uWBFII3Q8+QsC2YH/dT4m/iJLtuYFaF1inNo2IUUg
lyCsHoFhrQNLhA4/SngpUhuuxovaQJhP7N3rakIwqJT9f5AdfhmfgDc3UcJOpAYtk+2DcTdXkxnF
ndepYova39SF9iCVVKdp5mzn8261mjF48POgeCtX6Vo9X+TIlY+GEWmW/A627HVJ03VyyMOgG2mj
eOJA5f/SF5MeqleYbtSc7QoLnJQTB9u1OJYzr6zcHaojy1gT5vpsnvnapnQhwBuZpnh+C9Ro67G+
jHoFUJLQP7DogDLxbUaF/wLpf6YK+Etz6oyKxqqJj1vhJzpcjdB3Tgm3fR02p9VyfrXvsnBjBVY2
LJyclRI2LUjDF68fGdDvrOie0Aa3y/iYADFnSv7rMEWFh/tPL49Esa8RClD+4Uy8u9eZP3030HUL
NJ2LxwqgKjT7e3a8AZ9RwsRHZUpjyvUqLahvt9HYTLwvix6i6nzNUzJRIpOX8R7ed7xLofLXmav0
mmOqGnFwKOWpy1sOFUUhDxQQBIdmKEndIv0i8s1QFlo8ifExUINeVQLUY70jJJZJud1vSumAyj5d
Hw4cWBZl6DdZfIvPv9rjvEgd+KDwBQw10WMDS5IEJXzzSY6ZfXXnTjQLq9fv8oDPWz3UuAwovdb3
s0s4xP0wg4aIQgyQCNvBNR9Q7dQ9Pzp33yG2XaVX9pkraLGiHFUkQ04MdDUdJbg8Kj3VeoM6TUbs
Pc1mFNh7MvBE/ZjfUOtprjPxNoEZvsxuCbg1/Op/rIw80Za3xsSjrMQR1iuQqIv0p3nUw0Rr5/dR
ZBnvoP5Ac3VLVvivQyIrcnPJ2Yge/uQXG5WCMlVH5i3WHNYPThYoH29qposyFpA/MdzAKYzYz5GL
YAHZqxR7uwHlwA1OPnbYDSNHQ5++h9rc3mBIX791BqgSxIwISufmvN9VdWrOpcK80Zf25Xftjx40
vvpLcIzpzbF7tv+7LZVYyt5uxffN12+NXsg1TiQb5UH9qHyJylRwfV0n7weE8UTMrTVJd2vZi77J
3wG3txGL1Y2dCp+hTfY+OaS8Sx8wEiS2GtVDfQU0zsy+NdiWFlwvDyrCU1FTiTkBsUTSyJVmHOmE
ApCVJ8t1DWixRJ15GYRPkRLwB6m27bI1tz9/TGT748Z9VmcZOHUeaw+0TKYW75S4SR6SInk7R96D
vSGpY4yT2ixKjboOGyHDqABluhbhob6KX7Ma/JBLcvAkgAuxBIGGAlBpsKDD9VXy2DB63brZ9x5k
IW73Urg2YPj5xnCXLUF0DnXS69jOAhC2mh7iYPOuqGrAkncnhxRg+6ifq1P7kWYAkZ2Asze05Kr4
QeZijQkiZR0Wtm0jnNCirq4Ew8LqXcWVzbee/9hZjD0e/P8o612ZgIMXuCbJnyzqP41g87pm3nAX
iKNmQ48qO2M8Pt0bWnkTRiR6zF/nDSoyLroRbwZ4XIuEzLTkDo1oQ0QrQmcwB4CLEaPgfs/a2UbI
8gcNoM0GsnaXQ3qaFyEUy7LAAhqAySovvX5wjfRevUxKDV2DlAcdM8hYPuIb2ZPpTWAWpp6Q79p1
0qcoaffVzwkEDvKbdFrAltsx6unjlC32Se3tA3n3jT4VMWR/fBm0Vc7YK+QzylUkwAp1wOIqSTGr
lW8v+BedN7ip++rvbJmoy19dVQGlcY0N9LwusayaYsZEZWW6lU63/70fmf/uu6sZXANyB6NCGFIO
i0Y++V47LA7nbfNs5MBO8dIdNsHcL/dmu2pQEyJbv9XX8FA7COKmlvLP8PJt0Ptlb0RMqxp7nRjj
dZsMqHo1fT8fyXpz3bKy90Gi9QcZiPfDd3hw1Yvchi1mtNde9nYlkWbnbEmaKULH6OIoGKQpdj3k
bBmsmtHLjv8Hh8TPSxT/NAs83AXuY3GE+DPrEY/3dHo4Xv61weNPcdROssAJWWEW4bJ6RR1MuRhF
qG6IdAsTHUYPvlNiIZtk1sE72ZNE17LX2oUMdw6xxCcMdJEItL/8NOiOomCjnDclwqIh1qQ22d9x
gEoQHO0E6/GQV+1hRiUaD+YZA7vKyb3Zth7NQ8PCcbo6Rtbr9qH7wZIbAVJe8EzrpPuBFg+oZLRj
YGyrN53AuCMSV5ZYfGPYnqXmvaHX65eaxVKLHMTHicORELkX+mojrteFqz8ovlMrslLqq+y78Yxg
e2SRB7BlckOwk1leZSUJP1ffqRHpYIncHy2dZfcFuIBs7clVoDgeE9WZ69x5lDe0utTEC41bJx0U
RdETVOjrTe9EmfvoS3ZICtidjFe1xl4U0Pes4kYM5ZKNjzhXE52Jv3w/qSxCadv5rGWAXOwr+KXH
nDYHCV50qC0KE7bNFnVJu/rAxGqKoJfZTJtciE/sYROz25ouNFu89EpPR7liC8CgxvFsHcJ1cwXe
BS8s5yeY+j0wmg+g1Q8ix2We5gy2fpOtvtO0MtJYGZDnU5mJpBaFsrIypVUWayjS+haKhqMzDXZh
1g/FzTPEY5x9xbGmC3H1ExgxE+QWN5VKhKB902ye3TUpISn9u8nalxcA23TP8bSEiXF67cmaVdQY
HobApzQJrIqsQ4KfxoJKwWacMol80dW78sK+N7XSTbVp2ePSiRZUtsv5Z95zbq0alAcwijah5N8o
juUUFBu/0E+qubHwGfYLmQlwepi+Acjo+8Qu3aPQXzGNJhAjJJb1Y+cjD2PsJ9hKQfhIDW0du26S
QAqZI5DM6yKPTs1RvFaDygNTSiWQnFIE4s38kEJsViVdh09LtyBek0IMlpdn+tAdSCVUzOS4IvHq
e1OyKSpenNSUPZpnYQSRl2gvLiyRnuRaWEUlj+Io3rSALTgTCkGzM3ottzH7th8jW4fSLebfxjpE
8I8Ic44H2k1f9awFqqtobKVKkMTQV7vpY+hBqLzXaTrMfcsON9wgUitoy9fkWkzJ03fouHHXN1ex
0yNqwBRXCBE6yMBjKsXwMmyzkQUsnqJajG6S4gUYODRs0qe9puXADbZ2AgY0ZTAlGg4JHErNthvj
5rrvHyoXBGY0cVUNlwNTobJmOeucvHrKmxR2X9KrfmoEpGOlqjZWeH5FwdysuReLD2XnvIUr7STw
AcAN/RiI0pd8xlSthby+QvM0BgPrGyVdCaS8bysHcGV4ulHXh5wuXKu4QVRjj6tL9DJtjZWRugFF
EoJgihBiyavt3nhwmqmOvB7rC2o69njgcYIC9HgBZu+w8wS5E++si6CRf7wVdbmfyitDnklSGpbe
ZJlJFck6BKkpbGCF/Fm2yOWGb6kHsGmkvzzuP+xwfA76X+qempdtsgKhTMwe2f2FdJr8AuXnzn0z
2TEfIP6/0gBMiPYjKOveAT9+beguRIMVyhSDNZw33qzNp6xSSQmACosUDKVKdXjLUcWFD5HkgbmW
ePsLwjeGCkqiPZv2riBr7+E33vBMv8ah5V28iacpKQOxlmukVi4LY+m3WlvHN2kMlQmJlN0eTbHt
HVwfeQd2o5faaQfxeKSVlI3hBj/kBbtzb05xD2I/cPeJVdH8UMaTsKwQqe5uE5wGRvVA+9gU4BYy
BGkqgVXW01uN1dB7SuJlOdqNuxUpe5dyB55u+KLed7YeKEMOe3PQtW5g7II6wE9bo8cPIukJ9Rv/
Ho7KhmOPN37sHalODvLfcrqwmaln0h4kUQqIXPWNxtwG8GHc8AVccFhpByUBwQXjG3Ln+BuWBeb3
TqIrRJwHRSvS50R9AGjyl4137hCL64aQP751aFaubjssfc/bVXkW6rA2Cl7nzh3osTHCB7ygOyA2
cMY3/LbQ8J8fspoxPCWoXjvyAnxkckOLOjQC3O8Mc4WRZXgGaKD3RFdKRflaGmLyMF78anl2UeH1
SlizN5GK3F9GV5uXsS6OC7dPubgZtQeUIbI5GF1KqvKz2tRo9cOsY7fXZKPOwDJuSHx/OFLt0ox4
Y5FmfYts1ZrD7Wr/pqksvnvRlww3pTI3jwibvynw8g7WOK6y9Ihj1ViYbDYfugWNbVYqguP3ve9H
CxUZ6tQu25DasbvdhhsmtW3IcEg4tnq3gJLzYKAyAI2XmbvXU7534shPNaSnrij+utInpmobMGI5
C+0VYHbghH2NPAFCBjdPwNb9J/j5bHo7llw+YjfX6fv5vHbd6vj7f93rPz7unYefjgU/4/U+LUGe
NcyqjX3KPo+E6OgFBb65rh+4VNLDhfO0GQR1/rv1eAkPg7bTTEBWGsg6iRGzUpSHTgP5PSXBfUlS
/unAH9LvhCWGHmGWlq9l4mi8uq6oQH1aE2+HOI5IWfRTewW8rxhVrNA36j6Y4H8MTZExQMRNmN3T
3FTARl377+EMNx0kpmeIuJYqUYVDaH/83OdX7yFI6YOi/sxT4XThoXtExNJbNh9Ch3m+RO9DDOCb
Xk+bmJYWTrAScsks4dEU7qXQbJ1qNZP2YtCT0D4zDB01Wr4wB/+MejHbAk0iQomjo+4LUQDUcWlL
WLmVQisT5PY7WmknPU+evktNqzBCQVTmrx9+Xcda7Bv1OaM9dQFIl3Wm37K8eDNN7pWNqhZmOLn4
ArQ4LsPEvL1TDeIPaUp3RjTUGlGeX/cpw2PuutR9A7hnnQJe+nuyBuijaInvpUOKSVcNC12RRaiS
yBFI3ugzzxaun32usj4MAXfdfA/pT7GeAKQkd2r1eZPP1WYDdCfSRZvRCxV2PMS2J5Zgzx00C+IG
x5fU2zPWG024v2+tLlN8HqpnOMMTq391Me0KlzYcXY/L3JbTIasG54RHO7FL8NkdH+zwYnfmlf2g
Yx9Nhunvg163eTYi+j8+TjonKOwh/fjMVtNGSjg+uizcQhGSGIP+WHAz4xZUNFCQrFJgHa8x+cEK
qNLUyBYVA/WE/YN2QEt1wMEWWmL2fco5Z+E8J8pKPu8Q/X/RsNztpbwDUy5iDsn0OZUmx4oyZMCL
OLTjdKe3lgY6VbjI3JVtif/rYvYSsjcHiPpOpOH4JZZ004totuLUSquqPzkLwF4fweTNOVhVLtVN
usdWRFkFym80HzLkY4fvHbbVAhkie7pOryxOvAvZJw5gSeKKH172VwX9BW70MZYr87Z5Du3IzFGg
WKZkeGfn022u39DHr+baj/xPR6Ttv6sbE2G1OgOtUvNJtQvhr9x1fqHxb5c3FDANHgWtdrrrR1hj
05doPq9f2/abVWlxyc1jcNKhFcOLGlXSBFMtWBGYDZPDf8q27CiG/POKOrYL/7H7hb8507sM7Gxm
b/FI6LzulJ7ZBGshdoRVRvKX9sT+hhk9xSd/9DK5HOkD6L2qH53umY6ET8ObtPprgzFBK+HjgYpu
AMGq/CQFLwtS8G5CSaITfwLWSn9Pz5WcsDg1EjpCwG0gsqenw5TAAPM9GzL5EBQPCH561bDYm9Ls
gYuLLY6XEkKTEddqLUZP1SM6B0Od5n6tSrlDMS53H0csHxclUoyyBS9XRoVcKqtkVsIO/UiaxJZb
qCmnAJMm8nP2z6jvWbpwDserM0NbM78cnWlLoHHFWdpjJmDxN7teRpE9BXaCNGjDY5oKrlWFrf+K
Ex/iw7GsvhkbQRzEQ0HC7cd6dAagTGKNhvvRf/WIialoPedYBVrcr9xLPYZ1suAd5h6fFnJvwnhD
iDDawajWY7tN/RnfK3rmHtvg0Pis4VXHSlg9AWosC5mX5OrMywMNRjHv24lcuWIKMkJdvJlRyUdZ
zELUr9bg8RF/W99kozb5UsL+ejSw+5zCbMw/1XuMVgGCLc96exluG0JrKAoLXIJ6Lr+DvkwlcHsy
IfsRkdppQnjKMTSmDxGFr7r9bGlJRzqvuOYBL/VMDyyeEZMD2QLk6cl4xyM9R207NLN1GKXItFq0
F4rqhPZp30HJ3SRSW6J/bzhVOl8EXaXKz3+oFumitOGwMXK1QY7zv5756XXL4J14ZoArRW2nXkhK
mT7ACohvNUTSX5yxCy1hfb6oyjpppYXk/20PEfkpMrxQkvA4Ujb90dK6zUHBGcW5SUI5bXYgqigS
0mVlvEqU+4zpY2aixafV+g5FKoI89LVYt8F+iV/gQwn2t8O+OvSL7HSauxkAvEQHkZrsr9tVTw0b
wAEQrrZ+nwMoaAP93pqDoeplcAuIE0Xj04dzgluEgtxR2fDqiQkiq3tJHK6us8Qattm0Z5f+XQgz
2cOWwV8JUtJY8l2C7lQDTScrndRkPRPycBR8D76WOP2SEjVB3frZUh0dNQQvf2KrGNl8jCzanOV9
ZQyZEsGAPPE3rpdro1KyZjs6w7KhlBXw+9aKHKmWKpOAP3Z0jMnZcnFG4TybVK79kP856kGvDTil
z6hVuAfYR3Ot68/uTVIe5pCc98opBtqMMWZKpizrpiqvQiY0e0i0x2faaigRmZsApJNfxhQgQlis
UUG+b6vY3Oll2JrGLahPUh8YM5cmRXVjoxZwJMAC0QkSJUxc3GXAfS8Qt35BGEFNFfO6poRVwaUY
ykA7+8RM0y8cLquZVBKmmjWCfOpoVGpqEM7WydUviSi8mg9Qmmtpt6znjkZHuHQZPJ6HFNH3cbB3
3weO9UcJ4XcDp/+4EDerjqtLe7JuSC2NvFuf24xawe4RFP5lllC1cxYPq+tlrIYRhvpcJ82hXyxi
VkB1qGKfyreNZQTDt2i/eMiqV4XI6r3IaPBbQ8tvGiWdCfna/yoMJUpRJvh9abyzuwr4q/oIVz0Q
6HmZ6B45tT7yM24YRF9TbIpFgtgxsH0KU407UPY2LF5/SBVMNAURORGRNo0c28odEUeYRTY1+BIr
J7XCKTkFA5Hyzxd5IcYJ99O16AfhmBO37tVP+SJ+R7S+4s8eqlZZGJTgWPeviTXYHhIPaCKn6Jqs
A4WwJNxBVDwXO8balotdLARmUP2Sb3+F5duc/CSD4JpA7PkJATsQSS3Pw1xXV1CFKVkYUk+9IeJF
4Atbdp0lKbzIsS5XQhZCwp9AEZb6oiJMygmS7nBIPl2pZeYSDNNOciDAXFJOs8oWlTaoywYzxZ+t
74rHKY7vfRQV+t0HuTjgyT/s6jbr/HbuKAkTQ6WxroIr/3nHzCRklK1sgDretlIocJawQ4Z+3wex
S+AyOm4ZmirxwYAVEFTlIK8uCKWHpaiEXXUKfSiQe0gv7RdsiPBRLwiAES+Fc9x80zUanj0J2NQc
RgHofSZUsxV7OylU9/kvXXtktYjM0bVBsXbOve5MTOMzUl3W42C9l+Xh3WdZTyKSZOX9e9rUHjAU
/ctS7aDVHssjbm6jB7yskdm101nPUU3kAqx+tcdNEG+zzh3MoCMMk9rkrb3/BPm4JKuRQNyC/P6C
FtkOtkKBLgw3L6PePxB+2kY9S6tz4qB0zdKOknu53JPjR5FPubwIvde4dIFHog1DdgRpG2WZGeBl
qUVnK6+oURxQ5xvY5Ux+0pUiDfjqoIYg8qr3EF6N+J89gVFz2gxs9g0pg1NUaXLjl8WG2jdi8Tjf
oC9Wn+xA0EkYhJyL6uzY0ywZ1nJP5y6SCSInXurarbB/JAZHPE3CzZ1M6ukzh/dtKkdK2e9D3kez
0R97D3wjQ6AY/VJM91rNXvCLvuL70AZCutM+5WLHU0t40N6KsaqEHqZu27qI0HgNpusx2O5pquqQ
xmJ4zV9GYLBhSV558IQGSDYIwP2md6+5ppEn238pi/k70Z+KcO8Sp1c3V1dq5nYS6bq+M+TGSxTY
GS3qj+47bq80TBtoIvamOB/oqcd3Hp38kBtcGzSPEC04lnYQjC2Z7dovansA0sBf5Js4L4tJHgni
S/B4l6RSz5yjaixYDWH7H/Ra0c+42m+xbfkSWpCk90u4N1mvN9z0KgsEdkqu5Z+VCpo0Hnyc+N4B
Rogutgn5Txxgh7Vxlje07jgcfqFPQzMTLn7AZhWzZw9kGWAMzPBPedc5mHo7NZYavfewjWgyyVcQ
wbXdh1pPp2L5ZKW2Udrw2ntBh66khD6Jkfli2C9FQLmuo5j5ddPrZNF4dhO6KRY+IblO5VEMykLQ
Ux92dtRejqke1XiI6OCMw8Us7Zles5kgc2uZyg1iQMQxZNHaytP5QrB9X9/FhZBrm9ROyGVywCJk
LWG3ysf7xSDmZO0uX9MJAH6g5ZMhUBGCq2ReDnbJ886XqfkpSpQnuZqxyL88aWc2pqesbQxaC2Ai
nC02M3cfHA3LZiGsQvbgYgQoADuslhCKHu2iwAjYlO/wtVQlrXyQeOCbowpntmSvP1vo8yK4PaQr
e/ImBeS5/bWKbbcdyIE+RLPB8Mo4NAN+SalQbF1o23k3ytLSIveAvcQUoAMUqgQPudRRN8mIsZiF
VSP/Rrf1v7zYk1TpiL09hi4O+ckwPIIuejCEyVz9sIBmaspZMnEi83m9yeWLPXguDb0yESHgXRlE
qXpGGJA7lwZ+bb+T6flpi7px26RgRYsZsHFsc0ocKr2jIJugjByMQ1FjB8blH5nWb7HTsFDaRDHx
UDZvJk0ByvmGX0GrASJoITGwP6MtMJu2+w7HUHp4nYd9NR5AAEW1/XI94LUSKY0kwD7az7cyugGO
5X3D8XezwqzhE70VYBYM7A1HArA+QKrCYZzaAgN254OyeikLtPnB9rzc/Y2HmKvhTcxfjRJecsko
N0X4g662WiwkLFldzM8ujj4i3prvxb5ARogv1MwzhlshdTEHr0SAWiLbk+oGFUS3t3QWss3mTkeH
1nCbfBtoBGa185YAZ59yyI++N7F3PsV57qwKSCriq/BZq+MfcmuhLhySvyXBJK4zSBo73PGhexW/
/q/uRgFWUVsfPiSdB0enviNR8i0ZMMCS1x4pFbhwzEwmEz6pyLb31RHlfE/FYp963sTc5kCyuLWM
CSq4L/UQ+yuciCnCptpFVCBc1vE7mrhnepwRsQ6NebUpJIe5dfQfp/no46uP4MZo7/7rMAKnGqsa
nvEwibFhBfJcMx7oATGk4CEBhbL7DpZF0/4Wniv4MzFUfZCgeujauVDwLCzrnWd/Rtmn/kGr2Jnj
X45TrtN0PstpistIgdNrgH0lQKgZeK7tWFKvnfHptttrREFHKlekZqskZg7oa+XlL1WrHMXUZ4Bs
LQhgegP3odZFmSulAkFNWUWjdRiOx68j271lewpgJYT++KOq74SMOdyZJxq+EAdyBn0GN6GZto2a
+1UqgRXYjh/uAzEC0XOvgs03H7nI+L6ZCJhGJDi+S7Rer+WSloxirnpHp83LbeQI88fKgdK8nZm8
rZSjhzFx1HJFBFtfHXK41L5dij8g5y5gIlBvcZxAUdemQWtq4NCtPq07L9KOtKdEwxgkBWExDhYk
diC76JFQ+9sDVDC4/E7Lsgr0xwpG1cxF+tRVoxIztiYcF+zvpJegbfgZLveGqkWfQ/nIeVEFwc9H
bSvsI3R+dOyQABD1Hgo6YUc0k/5Q5q7BK1H2slI2xu/r/qe8A74hkYC1p2uQv/WENx9Z/63pD0QE
zv4v28/j/OWMIrTZXr55n0UAB1Mm1fTgj6GzVR/8qL6n/3CuLFWeWes/HLO+ohPcJmmQr/vorRDL
ttZzHy6mGdryudUQif8PKhmBJiAacaqI3tg1nmd16mvAbmsyokyC3HBfe9Cz4tww0+b2N1ZfY1CC
3MbxhXrK2H3TNMpdzWyZzCoZM6nQmOO7VDd20JF9Ik+JU5ZrigZCHRtcQ3nXZyAUX2/n7s+BA0Au
q3IqonT2FE+10h2wdMVW7I+/dLJpXkTO5SJia2uytNKLPWu9Bk7teGHJcSeVnI1cef4Z7k9jlwz1
1D20rRe1nIjfobsdBI3vJ2tgzZWaBoAIdPTeGejKJoi84jXfl2zPgIAz9AcRxdcCb+2Mxpb6gpWt
UrjD2rNchasrxd7HnckQRn8xvNhTXqaXHtseUknMYmjnhak+lnitlrrnsHDXlN5lhm700cQLE3S0
c3cZRasWoinkd2zSTvpHYOr1lR3b6NEVs+I1IwEDtLs2UzroriyHRCgUcP5mNFu7ApSFWl0dzT/F
cumwDQMjj0xXFZEqirG6DNF55uip4M8lx56vIcpbkp1OenQNffJChz3qU9FCW2M2kCvIQPdkii92
3KrMfnm5x5arsH6vnZzJEIkbgGey/nyZl1geo7Y4SIIzjT4s5ISZdBFCJVvQ/doOivGuMfzRLtZi
2qlhwyn83lMTjrVNeVbVX/jHTK1ZqSJVT9NxsG2QAfLnmOmQrBBskivO+R5HDSfPN/vfKx5wouQc
5jzudVuJNG1faFmeOuVmKbimOx/0iVKy2KQj3pf1XgpX0c+dgOVmVNGP0Ss21fUhsSLLnx2PoaUk
uKw1SxWeK0zskGzElPdOYXKfQuhD+Nhg0YExNikXumbh7vmgv/+rPYghRuoZ/MhOUkD8gE6ADH+t
/zLYXbMj9IssaGcpwayfUpLZMiDzviRvAErPWJTdvCFJy7Bp4uzpxrPo+IC514JibTQRMGsZYy0V
I6Nj2EqiGXRUmFY9AlRaQhLOhXc5uK3nn5sqQZtpR5BkVzCVvberZ69qwGq/3li/dZhtjtKRJASK
o+GcjCkjmB69C15t6mW1ao1EOo+h2kFQsYzyFnwchVaI0lP++OTBKBICP50p1LjiyevFReawSiZR
0JHWuqdP0Y7WEsPIwGSnDTFsXlqtdy1St+CEnFPJgQ1lx3IF4Ql0vQP+WiuvjgIbMRf6/eK5nrzv
XHZLEgesHW2yaq3005Ha+1IfourB8Z9B+JAyH12M2V6Wi8X+A8kUVwUbkVLwHM3wNtEdDGOL2pLH
dqCRyFLvN1mAbHo3lLECIsQns0dEUlfi6h+Q+BgWNEdc+4jCYtGriht7u3yNpbH3g7SSzyOV1Z/K
t5rcp2F44JkscQYdYvZ0J9+9VsaFcc5gK2lrT7Be6lSbICpNkiWtxPeAr3w1Y2qrkcERJ+FmvBcR
yQ+urqU8G/T1ug8zo7dtPUxfrdd2SBgHZgUaPlM6ECtYKHTuhuPgrKbkvkJt3Agd6irpJ7Sy+Al3
hX5RLm3SfZVI8xyF/YJsmJ59HOBgq+Ol+bIcIc/iPpbUq8oGp2HpiOdRqaIxk2AqNib3FhppEVdJ
kl5GbtEzIH03tdB8SYASzY1NfXmzgmfzLtobTMybtAWx1t+bp8s+tigny6bAE+yUiilYVC/g1bKf
g6L1cYvHXswzGGTSv/vlcs83gR1I9JZOfEJPyZNKrFTSK2GUzFuAMgxRru4SftHqhOXxiesHHbRS
haB7Ndi+NrExdhlLxWygFGuee9yYdgoCMZwughxeTLDhOM+MbrZAGMf59dzYptOl5zApv879Ne6S
iAUxpqMzT2HeA1GqUdTycQmoIfqC8A+pKdsoD0tlQkhbyviCaRIg4QfQfjeZhyUe6Nwg8epH+IsB
UHS8xluv+MiDHd3v5eEg/QkK6997gvGOUyqP2h5S0Bur4ZXqd/yML4a4cOhTc/1JTNOHOblZsjvP
aFataYY6tFncCI1MOXxN5SYZ0kzM/F7E7ZB5oduhlXLt1+20PLcraLOrMs4p5y6AzgYB2Hak77aC
Wh/8U/qgTgX2jvDWV4P4lAjiS9IM72AN99wwBi5cbUvFBag1EZV3eHGAxl3ZWTbA4jz/FuXwsa1q
R+rfX5rtW3iV27wi9OXuAiSdSOhf27MITRp9ChL+r0GSP5jWjz/ls/GJlfUPPcQBeziD1DbBm2lj
i64ngGN1dOjsY+F5rXaRQVbNRIX1zCkb+Xxfe1MfKV4Jr0qSVl37Rtn/ybXrbAp9sIBJ22fCFCvw
MnmvcbSaeRXi5E1MoyQXuAB3Q7tJJvgzAwFWwqgXFWiYP2X9Cfj7XhWJiFcUEZLIOcm9AIfKLSo6
AQNnW+gfZcK7NWA0p6hEnwPnQK6Dj1lj8qGEGDi3BoTkT+KDrX+/JTqEJ+MBlb061huszel3CBET
7h6491O11jalO2/boY5/m/SnXAnBJitZue9diz+V5K7tl+IhxWtG3L1ruoyxNneAW+sU8FbdXPtc
TxxqqlIbCSmCr15mfLdbWs0O+ZUTrnOn+dGuJEqPJuPlBFFbAvlPcdHsHuc0xf05y5LIQXe+DF4f
Fa3eocrHVP5ah3Y2WlI9vOUslc3C9PrbncVgfAEDhqpf5r63d45EKXm5IdMYWQSh/Yaj9dsFc+qh
k5EVyMPZz7Mro5aGUIIhliV75iDRVbuR6Id/b92cMieHzoyYCyB2QwVqACFXwfTMgSBsCruWicY+
vQc3SHSEC+d7tofs3iH6bICMT8x4FBh5nLNf4a/SxXNF9Zc5w9KENG/XMfifXExLVlYz0W+rEOyW
Wg1mEGi1GOveUgONzQVNGovBon24goHoIyIwOyiKqTahA9bAqJjZkoAAQcAfrsiA4+1+cT08uEkz
lpfy5H59PnjsRQiL9xho0ExnXA44SWdiKyr7OHKc8YDd5qGKmoczfCXSisQQkELiYn405k/+01Tb
JZVkvMZ9pPOQxtfi42aadD3BORNuVBTj6vOFf8djkzoY/efM7gplSB7qsxghGZoovr+bcneTSKff
QphN/cSNW2ZnStITJ+yZHwOuPDq42g/jdPMJv5DKaebGb4pjCtfBRn8izcmBeCbChJafOfQNqyhq
g65qkmqZyE+VPrbzm7yw56DLGhosfR/qbBCZgBlqBst54Z3eWXSDAB81rO6ou/C4yuwmlBPd/rUC
HzGnc7qABs+A9pcxE0P9NpzwrzQ3LLKCcS94bU3DchDha9glcBMAuHnbU/bVvJIPJQ2s6ytG+e9q
gEQu0rL2Ujt2l1Cy+HYf5CBfM1STNf7/NT0NqgDb7vr4rubuvHdCOpbeWHGEnPsc47EnOo1r0FXf
FzAsjX3h5+zEs0MPi6s1XtXCC+VwgLTJF+j/mKB3Anv4Kp6g+jm+A7s9inSGNoxHDtY/e4e8iN9v
kwYYp0WOFLlrXMA762cYT6RLZlXnpisJZLgtr3yEMLK4lQkGxKrRIXeSUOx0UPSJtutmUUOUenZ4
OEnL3v0OX9KYZaGuVNuqoUkZZZTYl8lssMxN+8zpW43Y9KWxiC6Hu/jnOvZMv4/KGfiEn/5atZfZ
qDhj8qNh7aRt8AHJiM8Jg6Uvp9a41NIQ77GAUkXErSl3cFURAuoEIiIaQG7pAtmTe7PlP9PC7p9p
WOM9yRXVfRqd8ZUZhsqZA360Oa08rrr/D/IVZeJkS8ZYN4Zo2bPbTa5D0xe+93h9+SQ5iSDd8Cmo
lpxPsHYOGxqrTUlv4koMrFouSjmkTU0TiukJINsSZVwlTpWDMJs7HbJYwJBblURQ5wQV035jsfRa
UwCoo+9AjiP+IYipuKuOyjcekYk/n2+4tO7WapRHX4yDR2XvAec1mN43ovJvqR/yrT/r3011trjv
A2z5goC1Q8Rin9m7ny0fc3rpq342meBqvchbDDsp7MOwQJ1GX4/HMh0+vufE7KC+7CiWXIum/z3b
bJNtZB9pCpl56MTj/F5rUUMIeYhnJiYk9Y4tlW+ffq5EDjTYSZphysbIQVsXAtsk9DYSvna4varF
KWcRDXKwFs8MKTymAmuJT0o8YlJzfjGe2VuHCvFui5OiaQAydzNZ86TszAMVNi0q/7eTL9qkGv3F
MtvTQBIDdF/rkqgqc7gTeycKiIYarNTOT1j9Zzkvs8kSc5JfoS6pHV1DHstFkJp+wXXhmkxrTONc
ptNXHRAgT7aVgpWp8ydYwXJQcbXmovuA2kk093Fn14fpI3ZVHn9gRy3x8O2ILO7bu91mAxMtg33z
VzzNChN03jB0ISCCiwgtrJ85FKeIy0cmKWYtxGFeyHYD/ktuOqAFfPLXs6RfoY5UOfrC6wNC2qog
QZ166fU0v3iaTWPUmngk+Z0UB2gqbWbJF4zZ9lOA13vw0+PrMUa2MbEOGhKidlAseQQj+GDr3NZI
QXyLnBCqlJWpCaTZZkVYZQddnMcoEaVLqI7MuSztQ+KUFHFb0GbEzfsjkoq8mMJCcjhzEkziM0qD
wX5jcPBtE1I0Wj4kvCUIj7rbAVDTI71xiPDcwW38wEWmUwg6Nt+6Zyk+jz1wC7N9dQxBOHohde9P
uC99mms/eikc8KYXGl/6PllIt2jWkCRiRwYVIvmUprpB53OMzJD8pY62hxPPhobtbnrZiFfzy7sl
Q6vlEi1zRRNaoL+RumJGRe+vzqN0dOQBkd1HnH4CKygvUDDzcDlf3Xs95jfzPZUlkQUz73jzwEe1
LPxUPBncZiFJTeEegg28oLyoyX6GD3TukKKKNgoAWT8mFVKf44OZ82qzM5Sm8lpK8PGA7BEA7bQ5
ZavfAOmFHbb3nhNKcbEoHrzrzWDuVSxHAaHRfOjFZp9c/phiW38J5+yBYyD7xPmVRxUjQ72HcW1O
EqkxGOHSEZkgCNumaP96G/vPD44xraiNg7/uapR0GSWrE75f6WcS4HeTHlv+BMpBWc9+7QSjfvxt
mBUNTFOuKzFKdU1YNCPs/smJ56Bo8UovFRn3wTLbVaZx+cFBMtxAZ2dYE0rI4yx//vaH7Go22i4u
v9rOMjuWWnUUi3M93X6A9wtAxBEtiMDaJc2ARcOq3wZxSB83HqtqMO7axxFFzRKtCALYguHx5FVJ
8leKhoT/hoWZfJGHMgZIV5Z2aLKxUAzD7MoeRMFfsqgqviC85q6V9tOVE2mV68eOfxwc3uC4eB83
uDwbWULJIZUSKLkdj7sboUlFtSTOKQJCyJUZ4PsnILrdghTaO5+/StoQzzW/u0abr8y9extcAgjX
adMGkYjEifASdqslr4AQAcJvmrAnMxE1o2le8HnyPxuTB58+oWrGPEfVRtDRYYEe509HKCkf6lMc
HzXYFYHbN2V4YZZZx/qdAl9a3d08fNPgvzvoJbuy3/Q9ByWdEwjmK7eaX6YIbTFipRwf85OZneqk
LyBK64ssVQc/HVZ4CpCG1K/LL+hsDLL9Qf7xdwEimcamN6C98ZOUbNVIc87hmw1TEQkvC6T+2SRT
T4q0wubrw7/xEDSfY4Sfc9HPA96DE4ORfxNALHDEhrTDJDoCHB45vNqL9yLFA/QpR6EPOQtvlbdx
HVwrgmKp6H8kQa6trNcMzsLr1xuSs92N3M4X5gAlafqzFJdRKYI1HsnfzAVoE8BkrNBsWgdJN5Tw
FqGvPHviEobDJqfbFcPV4zbn4I0klCXqFBlrLqgLqq3bDoSeDEBTvxCEBj+SFbop9DUtR/bIv/KP
ORV4uIk3aSnv7s26UCNYVFvBVAUpofSheRUpGylkif0Ah4kX30e3952XcVsrrfcWUMtpdNd7F62K
VBEFAhq3IwYDabejgktC0jwdhqmjN+lPyB2iUO1Zt68TD58218w8/oXOpzmzlfCTWUpifJEor83o
k9IO2/1LSEP5+/8Bdmx2v1yMDgB3ABsejO08GfwNeNdDpDdL6NneSe6Z0m992hG7+OIH4ER27vLt
5vPVKAvaK0USE9ND3Tc1HDwKjQX3vRgxWVcPtU3mu2m+Sx8DT2UFhGqyny+a5NvnHG8UnaxBttEe
wOPZv1LaNSH8IRk85zw+m52VjXpjZrm5XfkMMwohdPz5uxlBJYgt2v/wTlAGnW/h2NtzH4XEwa5B
oIgKFCySmrgI5MA49B52Ccwh/8bB/hFymMPdR59EfUI7x2B3uNutaot45vJHbq0C14tZLN9hFeP7
jpo6A4pc3hkDXnaln+8wsHxqHJWLcrwaaBtEUUF9LArwwJJNA2H+yteaEVkMZdnoSpERJuMFphmH
bma1S7FEydxDIK0uGqT7FQy6MrIsAvL5w0/FlH7v0iIrtSKn/JE/8tE6lbVgbV6ojAaFyMj+hKrT
gj1mymaRnWKThul/vkgQbIwifaQr8M9wG4cZvruvK2lC94QD5OqX15U2oL6JlI3maQ5cBntJ/l5/
6yFkxJVJ1vHWirKbdus0zB2Uc0MhD4iPEI23Hf5eyfWweDDtG9ytnMu4y3NZEP28d1YdkVICiWMj
nDbh5g0Gu6mdnTqHO3HtULLyS6ytxcxcu4+FpwL9AIKxv0a+rbgi/rQRDemCfosBpkXO5+UoYuNG
IsYfcx3dAhxROlKcCxsOsIP9O7QNnGpWrs7JxbKZcjgBNeOAIyRG3b4dsTWSVDg2FI4nBu1lNcNs
84pR3zA+UeZvqlcCOZ1RLxyYZ1Y8fn0onFVGr5Gw2pU8QFe/3rIuhsw5ShtdBx7zdt64Bb5rdb3U
7pzEOGVeYia6cZgYTNQunSR/tN66bo0btfgt617XnRg3b8n3er4Jz5i6nCrNDYmJsWnBZXw5Hi6H
saKDIOiHEvbiBSw/6YKtsmPRks8YsF2SG20K76UK3hopWGAQHAr2oNNqLG86hZHqM4P0alBslDr8
S4wmyG2seCzrj64TsEY3uqNGKAL2Tuby4bnRpjAr0X+Tx/EQEE+tM3HutQm+FLADojf1SP/dkgby
xnLgcs55QHOlhGTjNW+IMVxpO2ZkWqQ5rdjNdqyafpSGF6cGshd8jz/hrOMFE5HExysMvwOSVbyX
xX0tvSvSHUYzLPLalMKyiPEsxgwAfKd/mUJlBF0H9VL+umtWGwH9kAUT3Rt5XhJOPElsC/S9m97s
3FNENwxFm8QRnR0IN8M/4TPYb0+3ixTI05TzHiOjdH/TOKCbnoNcQ3hgO3uoTzJ0T2i8FeQ5A6gT
YNQ8EJzEBsQWb/+0wMtE5p1q/+D/tOD8wFzu9O698PIM5Zbgrv/rHe6ac7cbGhZyl+bq4mHhVeHx
kO8+CddJE1WU3xt4dKrROf1rjspWsSEg/4EYy/hxzAgRW+jkCRYxWus/hlsIUM6uj3TbVf+OmPOp
rOOrPNjfvly2MyNmtfOiEKVNT7eGvF/KbJPp67qk8W4SmtHO7e0RoujL2KsgEblUxQPKW1ZfFvhK
AJyqh02dzy8TAvElgW5rwKOmxvI4q98bwoJzIanr2fpEIZECDO331c1SL0H1LvxNdQ/YVDIa9v1q
bFJ5yqwUnh45+Ao2p95/I/Nmy8Ifpyk2jiI6iehA/qj/5tSed87CCoErq4ZucRAna7rMHepFLZVq
7WmdXmETLzsuw1zrUNjT1YSO03+C/8hrUjaq6QE+me6Q/avoF2NZEZV9e9g8Tin9q9Ej4yFigtko
kZwom0B2ixL2vpknpABG9fNKtxfqMOwu5+9FpgL2mkUResEWwGxIlRNaaQJkxfy+MrBGQhA5cQz2
WexQWJzICcb1teWgYycQvjA89qk+E7kXqNaNKVul8YdljuEV2a4iSRShgNkHShsQo7v9mbRyGr3K
CB2cnsbmFw6AlQEX84URR7+BzUk18V+hrYJaG1crlwV+9iL0SPDENyki3zJkxlWsOZFAyzvzBxm1
rOw4o+k605gf2PS/hDnOSDOXFcusTB2Wcw8njxxvBO8/hyzeW/4Gol44xq1N+3yJO8vCPbuWwgIV
ADP8nAOfRoSvLvm2Dt7hOSqQisFio624oAiT9hldup6IKG1KF0yp+og1FF6l11jTRcqiJzGqeHXb
mpAA7XsBqf9UdvFEuLxE3aYVeUEa/mwMxMZsDhFoa4LIgodXID7UIzDHeI0yp5JBsAq6L+SeK4C5
bwWsf+m+GmvuSXvm9zY9+/UCkJ9dqmNrHiZnFO+zl/bx+LD3ZtcxpEFN7Es3TyYGY1cbLZ4hFUxc
HKLq6xrT0f26ymrFz34Vm2EljEuecH+djf99w8idSW8Iwrk/ASJTvzA3ER8hfdSPf3N/XFLFOkic
3Wp9/8eCtOw7LUdzrKLHHghFxTcWV33+wCLuncfvjrO2bIPNFSz9UA15d+m8P1bO6ax2jPdlIBTy
yjY//xP9tanvUR4SY5PgowJ61kz1kkqGzEa6IFE3pVZaKf8f3Z8Mt+tThqoW8UtqrLdOLN1EXHwd
wJtx7ea1erRiYGzeLb/4oML3ROSsPpyHEk1+2P7cCpExbQkKb4LyirhDqQCv9Cvjdx8nq2YK3T6k
kTK1cTni30cArB4QhuWw2c47jmZnrCNwcGuDNrIpj5+BkPuk47czacQzvCuYdlJhHn8g9ZkF0iNW
Jm5upuSD5JsTx1St5anPlhksjKGb43Vt1fhE0g8POIU26JMFsUbwspODddlptNnOdWZnjnvz5xb9
UnBSJpbUe+U/qrcTnCkxWeyLOVpXnWBBo8rDsRx0ud9Z/MJSWx1E5baYPiqh2FQI6T7QNm3g86G+
NqKt0ClS8yvfzV4v4enQjSmAo2GL6OzFjh1Gf3WQFORVKNfrU+6S6JmM4BpK6deplRkRkDf54Oit
dVkXup6cGMy8oSirDncjoraOFnckHJc6mJX16KpTEgL9kpX4k9JQnTXIwUe+HQBz+sVuzwecUXtM
rfbqgUTKUiABz2bIf4BTiJF097CAFZ6Dpuflai0DEav4kbcPzJb0UNMtbekcJABbMbtHxKGhyho2
Qi27PS7LmBs2Te2FZbrJCeM8laN5BuT/yOk9nTssAzlx8JLj3opiTH6Ztb3cTEfD1qk/JiJXF1sV
8ZVC/XyqvRP2inKPs6A9MRKOX1lFhD63mEZXDTia3VSPKu1ULow1w39JVhVOhbpQTOpkvbakltNt
FRJYLsnTQVJ/f/OvpT0QQDr/3ewLBYxdUDZJwQzNu0VysU0judcdiCKtJ8U7OPCaS372KKvu2Y6h
5VsQ23dIPHROhG3ewn+Yzf70/Xsc0fEmvE0bW6SXpnD8o27hx0pJqiNrdi2Xz7xMfpRArDJWVl1C
nUi5DCXa2P8baRr8BkYUHbcsoaGXpuwrVN7xxuv14NQ07yWLvuqALiplawisgIoF97eiUifE1mTe
9lS3X2S6fi/l3TPrMzIGIkmhGM75W1tYtVvkFZ7g/PjU/QIO+y+BrrPKfsawez8hvD5KINFmp6dI
bidX9EupKQdD40UI/r5HV4LX2CUWKnKP3gH7Yr2+i/mG60km3izD+nZMZwAZHJa6bhKW+vYtKTpY
/mEEsuN7i7APrQDagfujIURa/GPBMRIh2zGBd6LDLy5Gx/KSpyy529Tln0bUCg1WjcrBesBjY+sK
MocxX5ltTVvswKGeUIEyHPpL+sev7ClYzyq+1cMy1t/8VaInY+PVYgmpO/ld553mtCdCbZlRVUti
cpmiMXIhnOvAdteGUvwlxPNCPIe+zRCGm5Ob1yMdRESBr+8MvV2vRoVzl4z/bgk3gweL1gp0WjuI
2QtHCR/yuu0/Qj5641V4ffLzlJaLj0QybY8fa6Fw1uVcBuuehX+L+afpAS9t9+VgG1UDo//BrrPU
qGVld4Ek6WfTEN4g6k4zUq/VVTiXda+BPwW9ZqhOY6vJXZSQOqUMqWr46wZUyBHqmD8H8rPTwXUK
FOYRLaxiEy6bXYtELuCU4SZ3QPjk5PBkjrFewXGFs7fHXX1hL4suMAt/QofRW+Tu9Fw+02dgTVT3
z25s/Sg+rQB024A35qkBNxu++0W4DmweWGnPf/9qkTz9782wzC5YeQEvMpMkAobiWUia5i4xjCfj
MhLlGsVCvB6iLJQMZj+uO4l2PoA0FqpsFdJmg3lsikl7O4simBK3+SYbuQYIp9Q9dcc+sK/i5DJf
5C3qP0poE/bE8j2Lw4iSUCWtn2nB/oIlE7Ht/iK6PwGBLOr+nesS5OPROtqI0L+XfGfL0YqkP4v0
k4dAXA4jEEQ4CTbYCtPd1U+KokGJiNCY9vX3S1Kr0QEZYSMfnVBwGU4nzL3hKh89tslsuQLLciJC
BM73rZXbQfDJTdeOVz2k5PfUMH759XUy6oWAT1LSpDOQCQmmCkykGf1hTzRvuJChQUfRwytSV/yw
oFtcry6bdw6+70OEeNWwJYeIniROQWuv6yoiNPFv3gG+JlZVc0psro/v4cDcqMKULKAxwn/LHlKV
UnhdfjzC28Fo1sXlnMsZpLtT+cJvRaj7YuVImtn1TMQRGfwggDUNopYp0oVbOxr0Nxq69Sp0ILGV
UV6BiOfdrLUvn+2HCxSBWQ9Q2r9bIatXeEoh1hR32RvSVbzyXDFXFOhwwJBI6w1ihqnHoevfTGAJ
O4ivacjC5lwRkO/iXj5v/VzlqbRsvCpay9d4dIb5gZIqw0pgNqLzQa0KNnoxfaO7yCztE3JFzth2
89HhwRqi8YPbepfJTCeeVPQ5V6okg3wNKdLhbwE+E0AmKjYtK+sMIi3qargfBlR4plK2BPxyWhjZ
u6Qcjm7m3YAZWbHN7eKvb7NlnR4Ge4OOziIRAlBUrAOkrz2HT1q7JesxWI+uUiRPZLM780uympsb
6XSME6bUvJwF1wiJMS7/8RhxLw/R8HwdmwXr1wjn5NGP7RhaljLdcdANmYrT15UuI+MnLdIEU5WM
YADZd8Atve5vbccgGce7ZsAg6KainORFzmH3pic3egtuFn4Z0nm0Vppw9YvWlsq+iZ2UHslynwgO
+Brtw+hvzhAvgp6teaKh923HULjpzIdJvewBEJp83ZuCVkkzifsZxKFgNzPNpv1rbcPei0ekzxA3
6NvBmm7AAekUij5ElwD8Lych2jqqeg6I/Fag4l+i8LHyXdWG5vnqBRjaLbP18OmhMkZNxxFj0uUK
vag/9D0YT5eMgYNCESGUoD0dMEbDX/vsvEKkLu6QZ2hM2ie9VgYWOEB/Vkd77FTB/8d9YaZX/r7G
/0FNkahWersqmqnWBNSRH1yLCiwl0sNdgP2/wGq+zZZyAj1hQQYfv7kt0v3axSjruY3aY7lX6TXv
nJrLQ4TD0AIaky3daMBhLpSs1kIS/f7NB/3IMgVZV0OqJq/r34pa9GrNtwIt21yvesAikemfMoM8
2IKsIHlOHwjiJbKfwkOktDJHCORPafHlYv4I/oPiunDz1amVbIigepArl/EMxMAvNs2hyfE/V09z
uQVxMVo6IaWkzAUwpGEVLsQLrXYfXS+Erf31Typ4FN87fNWOSn2+uLlSN/21++G6cGNkbBN6O8oQ
h4et6Uy/1ECkBytY/DvcMcrCsuR509lJHDI/2bsb9BLYClL8T7zA7S8w26urZt4uk0eewfRk84ZD
8KXrUyCS4ePJ57yRNOSKJtTW29fBNTzySqWaB4aehnYAWowa+nLmovqWegfQcqD3FSR/JZGpDkgF
dIWrIvVYj82n+XzIqRAebaZglzCcifoQeVipzlIpLOlTcvpRQOxoGV2f2R3mrrpSc8S65TrERWxY
wXIo1XW7/rZwMaMEsl5P3wexY0BbBOMcP45n3yUJiOatwSeHjyIJV0g74Tj9kCW3DpEHeALIB+gw
mvFWymL7whTzseDjjIFFATn+KsIYvaSzZmIUs1u8DIg3jxT/YDL4qsI7/ioHAwgfXRW/F/ODqLmr
fTt2P7iTJ9UBFfP/T0ULCHisLXFsV5wc2WT335e13E8u25nliON8LSwDI6x2vlSCfV1hnwnMUGSL
Pon9GjO20Sx53Mky0nk3In8ZYVjlOj8AYLV868dHejwVLKZztSWx5D9ILARo9BE+uQ1O8aVUPSfS
EaHw7AAuhuOCLJ6ryJ1j+P5qJe4HHnWCQd/FI2aW+IrkVPahCFgk5hHzwHzpf7gOIAq+IaSmxGBn
bhvZGIPTIkvzNjCdgPMTc1+gRMxmwKowKNv6TPdK5k7xc13rIl+LUJnxwcABBs72tr78AmkGkwsi
OjbSd7U3iNYpCj47MsdF6Aqqk8YbZPEEI68gWNk/rwX6pC7irZhx4jDalFl3eT5RPB866cLDfF5i
nCEJM30iarEDc7rnMhwMzVHt+Gh3cPcdLiptTj+w8SBZ2weoeZQLhWU8qYZVHd6k2pz7S/AJ3MlZ
c/mgDLgr5u976tK0kvU0qGYAQYU+xO3kJVyrefdulx/Ui1sdblBfV+pS5qBj99B1QyLziXXKx9vm
yISJ54E0Yzby8BYKQWeapnh52OdXvWPt9GzctzeNPWyLursQ3gyX6sKJm7c+zFzyQSfTnN9ioyOf
538/4PGVZllxBWkiUIaSkiwBt91Me9Lj6OT/GpGv8UVmQujItKIX3l9bEyXjWrNp8FlF9MJV083x
ytzQT8SCuf+dY46kaifYHNRhK94wFI7+9ZgjexfaAw7ZkrpzCqllTN0rfhV5XTOFtxqkMES5xO2i
2gwbSN8d0JLZsQQJNeuvxKvnJnsry5vxqvYJkbh0QZfLsSXtPkJ3M7J9xwFuIYxskq+6pGhgroEZ
9Vzw5Kv+Rd9bDfaSewj1r/ayFiuAOn/QBLkZXqcno8PeIBue8EKdjPKqUyUvBKrBh1mTxpd2ZooM
UnGiG4Yhsa406yghl7AaOrulAhM9VHj7vFbj7OtpqAuzPHSmNkQGnFvvq+2xIJtBWnXyoVLCT3Dh
T41biFwD0zbxJAEzuuvFcYiR3wepDvNCvu9libqWcizFbWoClSAZjDjDrR+w+xdFnpCL4DDBUVb+
XaIzV8jHzOe8q+YINJ7RAb1DgCOLPEUAitmqYsihw4sxQgbj9uce1wsNJ+f5RZNvynxOeSy84VI0
GVPf2X3Qy2pJsWuEt6Vadb1Dl8fQCDAEGzEu8vqNEAW8TT6IZP3lqpm7mTRY27RkJrrsE4gph+AR
QgV4HGlJ2m68jFxJBUUCScG6xHzVtnER2HKx7XFi6YeIMd+UwvZ/epjvbWx9tP7AkfFPFZsICFC7
HDF8XTOhHgKJtbP3Ro3MJKvoY2HxWF4a2iHCZasr3D6qOu//7ezeglLpFhmf/WMGpbdlNGv6/u1S
db6k2TomU1F5MsenlDrNAB6aFtJF53IbcICQ5xu5GyLxlWdqz0T/GLEmr3d2YsQx4tmAc8fvSJUi
THeWnPwHDCy+1ZwASBIh9t5xLCH6HUWk/3jOyn/3ZFljUUM55bPtjq2INEJqGpoiIPjpGP5AVdQJ
yBD6MuF/KXd7nvqaFRpPE8lfWIihT9UqlhidSFn8FZJt78X9clM3eX4TSkQUKVMUGXZ9ieJph8lm
zovEhlzZRLNRQMQmXkgM72BLpFgy0F9xbkVcWP9i8fXvooABXc1zPlufjanlsNEGBMO6/tZdXDWy
6MKnBKy0VlG12lJzN+WwRw9cFD54p+qKo+KddukkwxWymo+9e5Vh3JDSfnUvjEJR9z0SQCkZ/xfX
nnal9JwHVALCHon1NqrOeiMorX5Is6kDYe+8GUMdGR+8mCMlh1N1qoPRoQlBeZASK2mp/RjR+I18
ZCJ4KdTG3Lmo5uXYRQLRJnWdkkGB0Lk7CCP+PotsDYqRsbbl72OFG4Kk0r9ZMg+twfDEh0Eafb8z
Z6s3d/P2mLX6tHus57J7peeG4TOKOd8NyZNpYpbj1W7NVTpYvNM9Si849cVCHbkSQWqLX5mcVV8E
FTP+xwDpjPElN/wAGMxi6oWB39NwDH7An82/saDSupiBjjDKHLKZIhJdQEMMsoZRlWxgXBXfsf1m
/Fsc8cdVEMGft9EPXfIeoVIgyhJVUt4ksrM44Ybb5UXB0snyNlXByq7NsTCFm7o0Lqd7Tn859/XK
tYTfipBPNhBnVI8lJiw0M3noO3smqh5gZXdmwe7U6Empc0t1MZtXu31xKhPEH8EWeAc8uex9XlCR
X3ARca57M1SEQhQNa4IMWkkTPHnQSpbuSscuSCqixT5fvlbn6E7CaFlFfPp52VtW7C+0IEBCgfY5
eOk744SRAHYk0fENhJ4Y9/l0nTfik9RGIus3jP4lB7/juvBH12KUf1BY++fpl/SqjPDT6ghycYqU
eVWQHriVWi1sfnQbEXu7Crv1tuSdLHO0u0sFg0RsqjqvWITiQxM7KuVCA8oE0IVGt3ynI97jZOQc
4I7iJwPh+nZPwVWkmYjefHYkwEFQ0P/GXWkj1hI6SXHQ6+k3ceRPzGotaRLVAD8vXWLGexfSdkUp
J9OiY2YCN4zGMhPs+BB7wvfwa076C1juJlXWQ3wxWLU5FM9RXDLGGeumtCyF7aPUMTC/LS+lf3dF
LClwk7IAPVInqcYfKqiqyGbZGHGNGGRpVoChtq2LxI4wbeYJvCET0uUAxwa2hyMoCR2PjblTgj0C
/KZxG0cRse9D0hJDolNFtiq3wSPwnl7Mc6nmN4uVDmNF8EfLGvtkN7xNySr+ZLB2h7RQXIgm0x4Z
Eah+2d+p3pAEnfji90dIcKVePvXHW4TNEtrnKSHvIKkmV373E6XD9VU4HWJWYdXbGJ3kDkB7IIhI
GJuK1e3ZodLlB/wXwDLiXXLCJVAwR7g/so5l96FOS0qRxyUCFD55Cu6YFlYPX7yMtHrA2MtxkCNp
gvSBUhGF05dtLakpo7mmufm8bkLdvoakr7IFjcPLR1WRFw5UdLspBeuAPQb71LXMaSj94WMbzDNX
jnyskiSnTuiVCr9hiTrBi9h1YWPnXPBk11cwBWJCyZnCN+CoJcOmuKh+TLDFB8s62B/9YGHwfm09
veErI/3FEAFev44SVsPDPn+QFNbcfp1/O9lqloRxkmRPDydHUtaSs2I8N3gvGLG5AnQ9PpDmQAul
BzgFuOxbboFebNHz110re2tTzqcVQP2xE8y2uoDVs1txkcwtV+KwKPkF3jbsvbOpkQ6bCgVpTHS6
vQc7TMCbj9YizYbJrvN4Jb346mHM5ae479tsIKH73dYxoiTNUdjbaPnnDi6eqVE+ectNlRfhF/LF
KxOuhC7yEqUX/7sKUXC8slvZdsoYg+rwSyH8O018dp15KC1LH3iK+ggx39VkdgCltKQp8H7EcaUy
SNmSffa5UsBWssD+2DCUvYmo8qNHUydyRPjtwICLSKpCfEMTKI4Zv9Un0kM2Z7g2lTEyk6pQYvoH
fJq0D8A+2VAdLlUNKUmIUAuHDscwdqp+o6W6H2B79XelVjoFb3QgLAKu6UOdLPODtSOh3yO18TK9
1Xv47uJp8+Jlnjkh/ToE2efzXnxIbO9uJY99HQmOHLWxVI4eqjMf2VKZmHeUmH5kfn3mbbAybHCZ
hwwSrlPTGVwCrV3bmvkVdMupbt4hP2QOFWlPcGXZmHGOBSOWE78GLHcm5KkC/f5QY3asg1iWXM1g
2mmyJDzyMHeljVQzZCZpMzRoP4WjpVv43ixILYK5mwfCiLIEVwInNzZZlzRWRh0W4cagO0idPw2y
8HjoTnsT3XJMDM1P8Zj7txNdsbro68cJqztFBC9IF7zxwROttOxKiFY63Lfm6g+xoBFxXJZe3W2B
QxzWMl6+6xntg/Ca8zMthWmM0sZyNf/NV2PNrSMTlFp6xBtCkpB+KpyMIM9jAZzQ9ADEJgp6hqGu
MNX/HSstGUQc2TGKqzVAjFDWhyAxCDlKGxx0/wuLY66MbYFloy1Ql1tKqKUmVY9urkh0wQPNCjDU
hp/LLCY4zhcyLaWOBdTSEkG3SZ23UNZjswjrAsHGc6UkM8MFyyPNOI1rRqgD5FLCDtbJo6Pk+jbW
Gp8We4ekE8SO1v+sYJatXSzKwgXP8rHWfIZxt/CC+As1Jts+5P9sdRxoVDeOEQfS5CejLCn7vo3x
5RXaMYllNxqzTm2JVg3+uHPxaEO7T0rgaj+4Lem03jo81pnIJcIi3bPzHvYs2TRkeRyVFmO0sjLA
VnVCni8dS78ACdnIoYZLyLj1yZeFDsXMuh40g7D8oiSdSmVxjzi41V+ednFDXoXMa0h/gC3o84mQ
jMiqC72JsVoFlEPETN4LPwa0Dabz3xu+gv2WGr8OhZk6Eaa1KyL5XVW3euoEW9gzhku6mbZMPQV0
WtW81BiasENbjq5yEfu17P2cqPWi+B6EHfl1LyWLErGCmgVVkBfRjHFl2IWUO71IUFiG48Jy2Z98
NDqCgl2ZsagwfyPGvV5msIMMl7m+/x2hjf12O1O+8AFU64o+bog612pZBfnw/ApLaQgQWyyM83E9
YxoAESE8KQaRO/sebgoxrW5TqE1/6ZImD59KyZJ488tqipjklHTswgMk2UL64B0tIs05P7OJ3/vJ
qGMskJgR1DwEtjHLeGb9waW5W8IbmxQBr28N5ZMd3UPkfRP0bisaBpGdSrisy7GO4f11rVXdWiKn
0wXzR0VFpMaGlrxKHTSkpMsZDjCXfo10KRVIQ54qmUMD1o1v3e8VM7GxmMz8Kfjca2mCU21YQXO6
aSyLyrKJi2exOnGIqwVkr0AyrsR8r8QwB6/VaopP+v/dzrbMVf96ifOurZY42VUh7IIDrT/Xd99/
5ChJ9MGrSO3wE/khDYHoFaWzx/qJlS5GhUR8EqyYiw5GMxKtW2h8ENx6mipYBht7/L1fN+WumWc0
XW0TiE1yHbOBSO63+f/9YlkuuLUVIIMEQr1O79eQdTuF/wurjxkgufSiDBeiIBr/Vi3V+Sp0nacV
HDEYrEzOnstNdJHjkcDGBiTvf0yq9jLM4XYq0vh0vKdrSs63lg/zkHW/1cFYLqGJZFi8CUEaVfBw
JCYoFsLUeD40Mu3NGJmmJ2YguHpkZBiVyIh6c1m+9XnvO4gfR1st+h+Sxt9yYZgzALtXDS4AOrlS
YqJUNN+3f4XSZ4Cf/HEHcgtMKqfmWU/IgLjd+f9t9iXMpb8kJyQuceqQuMUWFFSStCe3cb3+sxvr
feyv8WC27O0QnLjH36fXcQK6OUgHpcDvZvYU3pQVr0VUVhVAprJ+IgW67ZaOQaBOct8d7KJce+Ox
4Ryq7HNsS2GH8h1Yt9d1ZlrHfPnraTRy7jvI5a5ZY+3T5AVJsrwUusr9tNUb3oDSV8Nq1x5KinnZ
75MPX6h6xPtSp6LwXZ9LFvSLuyRc8hN9hjOGW7nirTm0luxKzke3G1vwBYbAlLv3U6kNA2y3d+Ig
Y3XvQO+Vn3lBACb6PPLrgd+H/n7MWTMkKmwi3NINvJEhbKsbg5O+JN3P/AtGFKVJ+59UajyRP/Zb
aSk/JJM7AMZqesqHDllVjmAkzLJUhYsPDOzTaySxxYRcJxGcx3aIzygaWcKGN1o3WBhqCBBRfEmr
Ue2+qgEDPtHMqlu6Dllw4QlyuSkIi9ieLG7GzYcE0PkQ8XhOw69j5SasY4XPo1K5KgZHzAAvGY//
aq1PLR2DMG+BrKPybX02c2I+0hWynEaJhOeW+8XlKnb0P9DvdhZ9MWBkngFIb+c9+Fa8Msi4Sat2
Cpd8EweREcvVPbhc/JVG3+LT+tdKTUAsEHBvDe3f89BBvWr5jzlZc+2nPKT9S24N7czagUHg6pxR
KRu/UAgZx4DcTZNRk6FwbbzMtTyh1wMkxN8eyLPJN07XdOgLsV54VQdmwaMzVVH5LCosFT2CCF2F
d57P215F5kxSPVdKHEPVZ382NaCvZumk349IWy7vb3ydAw8Ee7klakmSrtfXwRvVVfOHiVmlvcjw
EtG1KrADiuBo46NK7WZKoUIVSKHs6/nEYVtcQANqftoMtw2QzjLU34pnv5antALzvmpl5K7lwD3I
paWz8XS3gAO9XjL9YNLvmpYRCAZZlohHyNJ+lMuqMhVtrC6bosIKXwWGnqaWJvjsfSynP2Orj2ms
+nzVs9Ier8boRpSTdt2igaC1R3AB45Q2pRijQAcVZXPRVSL34kGuTzDh1rlpj0/uw24Y6uUp3CLT
6H9pvBKQM2gk2Rc5kgMieSTAVlKXIxSm8zEb9iy1KbQGjUkgojPPx7IUSxsXOcT/pNjGm6HHojyz
3cCLxnMlOVIdoiQVbaOG7OWkgUxcsP56xEgtCB3viDBUxALOBQzSdlKlPpU17PyPoUCSqh+Q5i6K
w+SeI6KUz0aeaXTwscGx3rUdZyAwGRi1owELZud25TXTGBgekt91d7RjK1MDiQxxjijWu3FoMjr8
Hm8JAtXzYIYyMfGfa1ej3xVdA/tATiI2KDd9NtGF9S1F9W6LgJD3E/TwbtF8dPPNXX/mJ5n2UXck
2lc4sZF8SvoJNrEr7nGb42UUg3uFX1uUvoR9ig0Hwa61haab8iYjieNiKSzJMg1GhCGBmiRcaBu6
Ds+Ho232pWqhGX9S4SpjIxCzPLURwM6Nx5WH4dJtgosIIaUqvGVNY/gIzltDCpicxkiazrw7sOep
vJSc++s2VvZ9oDe74K/ztpDW8TiIH/eW+L2VQO4iNLu0fpkiMIR9adCnJUioJZwvOCuQphf+VQ/T
ly82iE1mXfgOGCl5v2yDzqe6TIRVevRTBJL103uLTKc3z+9WKA2sBh7Z5FqO6mTjt7t/DXkTiGdG
0c5hAL1jxUs47w8DIVdJzr8xL/lT0KblIfOpWVHpPyNwLyIkCHMCsEpYOLd5EElh5/r9b60zy2Ri
erHBw6RtE0yHEZpU+VRTOsrBdM8yfBJ1TpO/YiJ+W1tznRhh0wU0Cj3dCVi2uByfCbWAPlRz3lz3
m4I9fTUDlnoBe/NWRIxBx1VtDVO/YXvaZgz7gJCzttAi3w1TJm4eAAwFrhgTtUz8EcQlEWI0JXP3
gUMTbA2Qq5Q46RQaJzfaF9Ifcc9ne6OjLVdSvaBnbGCSLF6aiOpUBWx/v7u4RrrQ6aGQCVK3CDoa
MW8IeEyFTOafTdnAXeDHwQ/1MGDXbmcNx5gknocceKu5JitrTgXL7AciO+zZi8EXj9YhbDM+Q8fK
uL40CEmu9s7/rOL6ApEnvWi+6Xi3ic4YH78fzbeOLLw2VuXBrI7Ly/ww7KMXK1aJRy3IqViuqS7l
0FQUlNCRk2CIV9i4KSr/9w+Z9v1Rh0dHrlSNBfScaZvcS97tXYgr3fN/wc+lcF9rgxn2zG2OAoAj
vdyVs+W4GN98s9a52uljBOybgEuoZ/I+CyjBpwPu9mrAR+K6yfUELbehemlPFj/XmNv3YUDRXfoy
v0BJ1QmPwhDyFcTLok0QCcA/LCBoMCC8J71EpNmO0q2NfsmyKfgOpMlqeqOqpgv23QDg0OPWb33I
V39ze60sbRwRHYF2h0KCl8ccq+UQQhF0CQbf5JSxo6JDpeV+AO9IwusdwjjqbC5pVCur3QMik8jC
riAGDSOTBS59hVht9v+AzvYK5nja3ZQ6gRcJtGlHYw+Z0SOTb0m1ek11pk4bBLqENnHacIph8eYr
hDmb/MesF56k83cw7cHBNFi8WxBxO34Zs8KXEnh2d6E7flLca5cmxj1V11z2dHeWNIM3C4ovUPnd
+0ELfy43RQb9UyBv/wgCxl3D/9Sjw+qJXok2Q8RK07+a4QTAP7+I+lUxyLyYvG/X9GMxke9JRVGf
POg1miuHWROjWOdwG6vwopcRyCI4aKM6T5Xv5aF1pqFsI/3bGuy3DxcMONxG/jXVWgRliZ8ZXdGP
LpkSUAn0yL1Knwe+1L6stnKQmjYw2qWhxH8BYkGE8NXLZ1THqjE4oJS4SzK363epjoenRXWkklCj
1d03u4+lbLGw8NHF3Pb0ZwFF/K96/lVYxUpCS+Kz/oszBZt3bHmrW87MZk54Oai/gN9NWWF6Mycx
Zpein+DdLZhCtUuVUuCp74HcMsqp/NkHQxXrc7x7WhXJrO3P19mzfhBz8nnQ82PIDEX23ZKDD/Ug
w+2LxNxcWh1T6uevH26bzQPK4Mk5iMDXf+vZzrBeL/Vnr9Kaw+RQ+emcYdoAMq1gfFOHH61rnXha
MW/KME9ysXwJNzvq5CM5je7vphcbJjLejg1rna9mCtst1hh4ZhnBRNTBf0hzj01kZwgxlx3T/H5u
SKJcCjMJtskK8eTYzQF3IxK4I6CmWFDwsj2SNaTwqVCUADKmvEBE0o2JGqDQT53tN7jp2OVbQX1x
ezYUN4+e2GJPDIEyPM7QX0Ubqyfm13zwKTNO0qSmsdg6kipENqBnct5M77/InAWTEW0l4w5f3SN+
+55ayP31yIIFvWBnlmHvgNkdDflw97MD9j5/63otCHEz3oe6YHF+NLMIzBFEs91vwPtUavLH40z4
x6hs+iKYJ/bVjWdANABx5agRjTtUmyf7KvxQguHY8NnulCof0thQBhh3VoT4cDCPjOj+gHp7qFGM
RRe+BmzGsGKJtRxykudKLPJDBbs85yOyL5hc7wNo+KpD4sxRVqbdDOTNyQBclOVMrvai6Mcic6x4
3jsmNxy2w/bQVLW4Ae8IDXHH1myl9bSxjI2BsGUB4p1yaRXWuQX1XP/ueaO34ugqK0hkomouqspJ
HPzqDfscnlFQMjkNVN6gmPc7fsTTomnJMhEmFzcqUc8GCjnjzGSuPmWjp+DCytOoa19x6FX2O0n3
0D73PDJxR+Ie5AadDQW9X/gQAwqFMafn5wTjwSndjiEhFKVP4erlEqv3WvCA+/ATwbuTTr3WjWaQ
+hKqcAApd1XqTswV2cQBpls0M70ipoA1ERjUtNaS66f0ELSUYFOxueLkQaq879fXDhbaL3JvSliI
ruxK4CQaeI551alLevx8TUnw36p0obnYUugdzQWtG5tbJXQDSo4KX0oDiy1DarxuYl+aHaG9s9Ei
5f0SR+8ljjHvoI1gx4+2LmFaODv3Edbr4eNrnl8vXdKt7VvTVK8Mm9ma9etogAx4MTa5OcM1/JhN
lZo61QRQoYNAD7tFLwKF9grxzpwmsbUYT55H7FydEosVERDAFyIOzAvR0GU32lPVo76KzCRR+8Oe
NeiEr2UNQbrWPg9oQvpucapGGWgHzsY9nsVAyEobKLWsW0pX5wu+51qQUW9tuQs25XD67b2ou9W1
w7pfWqFX8LrZTJSuUgZXPqm6FdMNilpO6qK6NpEyJ0LnPbYN74kwzneM7BRXenKMUZFNbco+GhLe
1nxnFCYFl5Xad3vPAcbTCnnyeydSV+J+VW92on9neARJn8NIqqtek/BtE6SAbGazUO7Gwo/fmS00
XKtz2RSXgvPHgSCKpo7XetNI4jmUqWaCmjf2B2/nd5Z2nPpKZz5V0zCxqD1SvdYV7v469SFSa6TB
/4EgSYP7/hx0wWqWm1Kq28dwF5vBRZX+wNhwGq0aH+fQvuoezASNnCqm0HBWLUCB1cx0Y7qJ5sRu
fmb0a8eS3GLlG7oMAG8ssYGM0Fu20rIV/XyqMEdsMDLFx/aBYdHIqH847MoD0JKa08tZhhy3WfYL
jl8Wy3/KbBefyLQUGInf+R0JtfLkOzIcI6nvmqj9qTML/bLeOJwQOBIugLXLzgP3VcLLug/VfPNT
JOLfWr7GLbw16KtoysQJszddgKcvMJZMvG8CIxeLNMVDxx5mSzxvwEZZWWlxeBWbyUs27oAk43nu
IpkQUJasv3hNfo49/cPEfWu76Kmjrbs5rNpbcGSVSDb99fXMbu/qVZrpm4wz7ki2h7KWHsTXTlEA
2k6nA9ZsdQCIRNY0qo+eOofI6WZS6AO3l4Uw2OIqzBmrSY/z1APL5jL2LMHNeR8UuzrosNSU9Mgx
MIF7vUYrLM++zgfsFvWxZlk5yERa85z/YOHK+0DnGljAJCVK1FDdVoikQAyI9o1A7gPa5pM87RVL
X2TpVvPRjUjY6LdBdIo7pRMpFFh+FO/DdJ5mceq1uSZ60dlKjj/ss18WZmMF1V+1z4cGU6IqlV4u
5Ufs3ggv5KgYQw7y3JjB3DIaWpYyhrsj84uOoTnfxZbn2mwwsjrveZEeXyoi1hZmzxw5ZF/qkSaj
S84wvdKP0iHSapWBkql8Vpod8QX/fHTD83ijFQVui2IEHDyn/kHtyVGtZNx/tEFQ1bLtrhoX+w8z
3RN4icrK7CUf8teXBe4jYCe40GxMDHhUMff6zCqmQT00/6fvmRHoQBZgNWdxguinAU8Ja2abCme6
+cxzatP+ZC1jYV1muJyUJLf7ilFFBGoBnUW8vRtEMEk9AosMMZkeG12CKKbhgpPxFmsMXzvIv8Wv
yvuyamH9k70fhCQOMdEYDHTFsZj5BWXMh+BHBXAhFHTWNiw37Mue9vllrgBtpatWjOtb4qkBVJ8R
T1ezxEPSk0L1e6ixChpnofMoVEjLxUoyyJEpg01p2ASDLNW0KanqXzQhuarLKfC60pGLqps8HYqs
YozHVsIkBi2v1USeCXCVogLa1pF7P32ntomvF0CgRX8bcBFa90Rs7O9HcgKBDU/oWUDXEEl1/Gir
tZy0wy8vNPYmQQQ++muGdZmwlOe0UjECu//J+mZiQ2LJwJAr1LSxn/b+iFM5YgUqsH2lKRLW0zF0
46/I/4xLvM2AtVZTUBruaoEsKdtQeVGwLAMKuosNul23Jr159zQiis2MS2g0AzNcNaOhnz3f3QMw
e+noYXoyaI/4E8EveSUtVeekSvJVohCQr8SFPEr2dO0YlHNjnri0wDHZ0JXLXqb0AL5LlOWBMFNL
usTb33phVZQcpw53C5YKXhMTTStFJrHrxHc23KKwvW1QtYukLci743T3D6DJ1Sw8PwNTiSTNWtpz
uh4oT6D1Hb14+EyW/tRvLszcwISQbUmQqY4Pi5GXoYH2TkbsBTcXFZ+8G6Khyu92LYt94Ya6KN55
X1Fe8DWQnx/lQswgiP1fl5KzPx+fG0o1+Uq/T25yL1kPeDcrIJd1p4Boy51lHacdGLCK2wh4X0IQ
d311MFpvt1y+BCHv8Fsren/ZuNwNtd8+HeBfnJ1tLTEVechVGys7HwnFRdbU1LG0kt5qzdqwUtHi
pX2wdegMSkln97fDj9zCr2KgpC0vsfqUcS1wf58/f+6L3lZzgxw9YLa6zsnkvArhmYuqF34Svcxt
ri9UMvxZahBcQ9P4XvVmptaM4bS9TD8qBOOt51j0dfOGxJigQx1WMNc6AAPqic6wvoE8v1SkWVA/
EnOryWmNFMWvkBp85yfyjRmJDGuadSCf6u4PjdvSJIgoeSo2zgA4feX/a4/W/c7DaeTSHUVkB7h2
6V+Ix5DElmP+OAbyziJv/sVuaFABnWTLyOO8RyY1530keyWqx/PeUyUCU57qcybhFm4f8I0+Mz7h
YcPRn2kE5aF0ISqpRZQz+yBrKmSytGXL9m5x/Kf8ZF0Ef/oOQI/b0P9GGXnMl0nkfES0AXRslmYo
pxJskXDXJheQGO2I1QfMVr8HATHY2XCyYHT5QTzpE0buXeR36P3K+zJUibXrxJ3S1AQhe9vwknLt
+Cf+oP4zDcw0llI/ZN0+m4A4D1jiv5+YckAM2Lq0xaSCbZX+mA4NnEEKTbr9t1SGbgeZYqzSPLiz
PiBqoRAIhM/FzcnkiNXeNHwCD2ueHFjAXoWqsqDukl4b4UvjMRWjV1E9X0r5NER+SpvtShAXViFh
3/TswD2CWpSOh05KZF0hYfgoD/LvuRaxb/kHQp8xQNJ1PvgH/Dc9rCWNDS5oD0lcWiuvxC1egpIk
A4asT9uoRWdqtFeJ5Vs1F5Cxy+13p8HyVr4OMGNt3MDvWeC28EH/DubXaZKFD7jDXDT2hfqx0iia
SVpsEG7b94v/R3n1VacpDl6/vTsWecuknqTCHZvXgxtNEZR2pVJfGHkifMCUTErbADhO3y8Nu3aK
pba2LihzY3U1ItUQSx8sh4Mqy9tPZp0fow53Z8GS1+On1OIPQXFS4Acz2H4/ABwYHO7K0KmCHB3B
Wgv3GSQa43QWcpJ0bubitApms/YD6crQW1mrly2TRUDqlghCpTNSzcXRNrFtXS5dSiIWkEPoBKWb
AFvXigic2LaWMYn8+3/NIZCmI2t19yqphQlKJ/8dpnAh9wcIWTrxwnxTBR+8agGQ0wAdP9DIIEl2
MGeCUc7PXoNZsAMbSs5FEx9hHxRXE0FPoRUc4emW5c6TA+DRYglI38T1oq3EXXZ5AL9sKHWG5roY
vjWwKCreNUfg3UaLefH7PQo0J/nOomKL4NbB18dbZA5xTdisBIyiczhazgE/P6UGxZIdr2NCO9ic
Wk4i+10qq9udR8bsIY9xdU4CfDH11Q63rU5ASprhVNNre3AfctgKy8tpb1iNl9fOSd6Nlk9VdugF
pntWb0xuKTYSzCtAksg9Kw+4Yt0WBz0UaFolzQW61VM9Ps+mEre9GLQb6i8kxNvTwv9oSIdBGEJa
J1fKA3Jk1ZRMt0TK1c1pMLDw8drQ/LHI1gPBm6oDLZKsnNZMPkKsvoQOFCx+GXam5d4AEBqcfT/3
CD1uXI70vnk+F+91rEaPY8e9w4bsOlD5p8I+hO/62EmPsqL7uGjAAHnpbzTYlNSp0Ni3FJuOrf6k
GjHm4HzMmwef33W4iiZa9JJYcA+EmDCD1TBEbCkF0YClJ12KRbqwtA/ZOsQhKNeNRcpPVGVFYStl
d5mFdVpcLaDg7v8uT667WT5Q7n95fqPF7PiTIXF7Y1EnsVTWcbtk6VXqrvUd1Br77O8RW5lIaxT7
4yN+PZsRCZoiULECd0xOf/a9e0CaAZYAsS0HCkH2bzRslD0a/fzzc2QbD8Uuxjn0s7wO7RGAH9JA
aOdtRnbmLVsFLN2nu0akDRQ0EJFw/1Vk8X28KeVfl4yo1JqWJYwKMJJNIiKN8ayN95NWpwa9AVir
/7pR+NE9mVzA/9lwsuENUSgZg5fPMBX0SXJ626n1J4mD6jDOdYM+u8jSFjUtuOehI0XBvNS/6E7P
Wd6fa/vOGpo2xU+VhrJAphVD5MFHoJjB59NpyxJU44T+oB0HGxDIxO9W5q3LchTnSGL8WlJvobDv
6jiXvRbN3bmRmD4pJ5bnv0OXlUMf46o8JeC+mZKADTh9zBOg11PDKfT2zeZRW+Jp1N9/F/dIwn7V
PoLRZOUSvbPhdHfApmvjxJBCQGNims9fo6RKddDCVFZhqRcvdqArX4p0ei1embzbvbz8zeaWzuI0
B3oMflsO5EW/XSktwq6bgbozNgfJc9cXogJhcccleyHGKeHe4rdLNSpZ4bnUqoSS44mEHvoM0Cye
qrzspUC7aG00FOT5HEHjkA+w016fdBXYycxLMkM0QMKLnFXr93iSNWDV/JYmwkd8iI1xS5p0SuRP
VmSAc+GgLoIcqmwPkC3gUV81Cw5DSGOG8A4ZexDjB/kz1VVq3h9+2oNEi7pK9VX0Y5yNeOT0x3WW
28dAKG/+ifCm9XvFBS8BaL9UoL/DIQm/oUFB2Q96ytA+zazAmTBYY57AMsx5Ho5xm7AiEOTtaj5B
+1YAxeG+kQUovsZvJFfo8sJDHn7UNG8DBzaDqoxerzTtkiDmHN5S3iPrJcp+OCXo3c2xVWMUakt6
ODrSkPDu3vKLVYdIRR1MfRXtRXrILtPjsYrkatxPiWaGucnReZjLGxflsz17hV5U/1CEueBVuaXn
oRQY7W4Yyz7dcquDYmN4Zx8Ql7TFfnKqezCY7/D1cdEUQ5J1SQeoHQnP/Q3XIMwDxqINp33JVJky
zHPnmvNDZTSuTNBqtJ0hok+uL7aqUqUTzF3kZphtXPvvhJ3kfTzKpg22cE2cBGu4oPtPtN6dAgG/
i7sf6EFY0wRFQVZ8lP2rBCuM86z6jrrn8bsbtHIFX0aBa0YNpg/PnyadoYizzj4XLUdVphm3vRvw
ZiQpqJUff7+fMgTawFjvPb7473KGM7X1ovNln2ChAnvwaeYiK2z0N38XGwcB37QGpDRVEaUxImEY
SXxK5bJewoIgGxPEkmKiGb8bBXiI8d86lUveK93VW7fo/ZDZMQwqXj8tS/7Tofyjwl3Jbs6ADfOD
uIsOZ4VtO7gSndN75Ssd3SbytsVNDJHr+WN0HJ+oOGsX1Fs1jPIjtSyeNb9D9Dr8n5HiSO5a2OX3
wz97+zT5+3LBa2GO9EKY0bBtGoxQUvOfVie918eo1lNB+p1vD5bFkCHZ5JUb5F9uAwk24BH6FWJo
U8tPpxQdmnMVhOVnIWMWGE8lvbOUQp60Tk2y7FLLsWeMZe69xmh1/ZXlYZRfIn0d4zi6A3CUyd4X
9tlsOSecbZMq9vly+lf+3nEOMA1WKFkAM7/7uCAgfk49cvW2ud2XYWmTB+SnjFbUaqHW7XJiwoQA
JXAIkQ+jrvXzlpfBYQCrTqWNjdPJWG4Y8a6W2Paa76Q2K1kX3j8iQqjcS0psm4Wh1Et2vT9L2vgM
AKJIfg3jYKCpCtmQrncjlQQNdiJyiFDpdg8vrq+ckdufu30L8IIVol4hvMbMpbfnSHLXHksHgHRB
M6WI0JG6AxxpdS0nCgtqkRYAs6WEyUnJM3FKh7IsnBV491ERHKbTbgBOCXLHWOG/CG3IhuCq96O7
LZbyoaZS5e/iTmnU2RPzK+uDMa/5tAfMpuUze2KVUWYPWwdbZK7HVIjt02xzSXfTsxMIN2qHiFiq
RLu7HY2X4bYl6ZK0Xv8940FcjJmYTyo3wXMxvd74+6pGrOWuz2BourwkVftfC6HK6H5Q4plgQMwx
Lcj/oDzfoveduuOqL5eQN8je5+mLlAEkSbzk0vF8Oqty95womUA5EYlVf2XdvyMfMJc9L2sztJCe
elYw/s4MBcpWMj9whM1YS5pVgS8Zd6CvWfVXxZp5ow6BWyXUir4QFKWoPK/6HxgovmOq+bA0jOY5
rsbIcRruYGNtrVRdCHCrLzth0y2/xZuvILqDNGHWA91hqAJ9rIIVfw+mp0qp43GLCzXRrID2yNgr
wPbKDnIAmgOYk47XDkEGENbILGZxpw8wDH9NxS/lU34eIyO8tIunQfVj6wB8XoaTG8ur68hblpnO
B18b1vSIpdeA4/OFeGEs+iqgx3AP3gCzdZOyBhWRqw1DL5VoF/YLrVdYMgIBooKWZTD+0zvE2FDl
STz7vuHXxtxkOUn/oDMmq1hr3swnt8SV7aNdS8gNxO15jk5tUPl80e3oemuRqSfzcBz9RLGc3fAl
tO2evYcdR4VmmDflY7C6SMWA8XB4AElSidCLoAJ/B8nlkZKTV4lQO8AxXCHmoZSsy7IErw7H+TYa
4IWxgDwMhRkNaFwOQeH4uiksLQna++Oc2y/24eMRoHYPzzyjT7en9l09hgrLv3qfweju1+wbbKSC
x4EOcBTCjHzWrivFjZWRB8LArmkGzF3woX7zoTQ3j3ZP8kDNuLq0fa5hirbswnmvJoArDPzZlrGp
2Nqt0LoS9JOkACkHKShvFaXAzoEzaEH4OyNCpeV+KqVY6a8olDmCsEvpXQAt+QYk4qP6Aom6ATo8
+dw3iVNXwHTmJA13Ahg5WHNLGeYnNoqh7F6KFyKvMIVs0c5fTu0K3wuUzt/nQuTycbrskOXDwIwi
lhzizmChREbbjuBWQDw26vHHlXN9zgPlEmeyzhq9XjVRpJHV0LMaBH3jkKOgqp0c/PmGaQdYo6RQ
YCeFo2qeaZah9C0PwRdojT24ENcETP/YkEV5YJkmzLkutwBmrkWp8Hz9ZgAtfcZXNICSWbGHgAjv
UeQqeH0IdQ9enbSDLF9w2RBiOCS3ey39ji+Al0uNvmJ+bA1j1Au0iy/CJn65RKqpn6xVhpuvfFsg
6RI8jn0xnP4tlTXQvtB9YNk6UW+N4/LACHzIXizJkBrT/2ULjb8LbnMEITZQtqZRUqKnO9nu9ncE
dLaE+IA6RjFdsfmaeSIlQGnkqtTEMhN3e+UhJ/smdRqkt8WyWXDdfmppYDosmROn0sPTfY1wz1zV
whY5dYvL//abMrEW6k5S06IgVon+y7Eumarw4NLCxZNcYrW1sJNOk4fDuVa7uRxa32LiXI0u8N3R
zfZ81KuouCWOGvaE1P2N0MCkw8XQRrJyynPBMb+o5PPZiHyuXBLMeX0e9LwMg4ZgneMpcbdLe54L
n7E0uJyA3G4fK+N6greDqFkOg+NB7AHJz0MbBGS9SEGDuMrOtbd8XrZMjzYFKqZCyqiCB+V4XAKq
CdOaQb6M07ory+jPyBJ5cSkV0US7IQeQXryZX3twi5R/+mb1Wowt2EEWGaI/ETNzRuq9K25zyZe3
bzAcUMWwjdYMVSvhS6SAk0BEjFzv2L/sPFUAoLluK0lxRgioyMOoPNZhIFRwdQa7UoU9EpL73AKL
IREqMP6mv2GDYHBbKZQXDFj/2XtODGwftIRzojNptHdJdIsPOYWt17FGAzwefcs2J6dc79VcOIr7
zEKEEzczpPflc0GtTAd9RGceSVzCqN4Bddm2x49c+cdSUOrBX4DG/i+cm0vYYDvo10mFnwr/NfYx
bJN914r8ZM13iSEHooW2IThewEMGDA0FC3hQH5uu277ValuXt+o6wIWRGWYkVGX1RJUYyNMRO6tR
hRtkUvt4tJwvVCkzwQu63qWhWn7R1EdlWuaX6299f447fKG1pNuBReZJuGYR9Av5obOzrMhUiyfj
3I5ADS2Sq9JHialZlQRrh36QJXcf/1AfaeE3nPJeF4sT2EsEHxVjRnIliCxC37x4Ze8mEy7JOUDy
uQeNjTPjtS0WZgyRTKMiaaHVPANEw6Zr4t9Rj1am97JLgBgU0GI+m+sv2/lYnEG7PgmJ9lopDhb9
XRsl9HiAqAonZYMrKftSunrL0UprGRrYGklKBI8CcsL9ijg6ZbS+K6fniHfkY7x5nkzokOEvUo/2
5Jc4iGyY+hrk6Vq4wUXdewcXm0ghOHePdR0knA9+TFxat7NQy48oy3E2xLAHoyUM5Z2G6MA3i59H
c1xn85MSYdDQS5c+oP7PoQN/Xz0Fz472mbJvDoumzgp0oyiF0ZPBoYBbAa15qVrGCgkN0jGo1qsL
1GFQay0Fsp1z26D8Ethtp3MR8MqoEuD316+wld4FHkhzlcipgd7YfV6DMEoWFQ/VfwdykmlsQuL1
zNL/69MuJfc2OzUAuUVZ/sf4W64r4TZUDuyASevbo8cUymYHjvTgWnfM1lvW6e1bSdirpGVF43NA
KDbxNlfN/RHSL2k4bXVaNokTlC8aZJ9YPNi2351GwZTAhTqtwbJxqRkAoXfoSRJlt43TeUsp+rSq
uI0P/brX49wIjnnHACfTrT5o/mTHavp1G0HTGVSAOcr4DLXhQaX4+RSNZG8pAwbSRtZDe0xK49vL
DyKlSUd3cExGt7eyuLD1fsVwHMAdjY15E7MLJD+DV1z4RrAal3tQp9MKBL37GYJNM7BstJZxk+1J
b6ruxjuD5rwd7eUQO6MFtDzZ5lhmclmpLX1L5ufgt9duy4fn9NEBysMWgQkUrZgJLPykina+dp7H
mRnoVYHF2qAKCnbnCRks8eMJEJr+ZUFvzeVez8UxcjRAu+zUZ038ChddBpGvIdUVqKdVMcVPou9Y
AmiivUt1JVLqmgu2w6lvIEczEirdwhZqIiwYXyeFKElEy39G3LcLvqg87NvI7fQ0L3QVwSjWuBWr
6ojrsNYgsob+FpG6sVCfiehztMOHHrREjwS6c3weNM5UaaJoMVNdieDikn+aTmjYP/704cF3pous
ekKq2dJxvO41N76P4ZoghwRVfZof1unyPaxDiOeDR/UvU7MlU/dUxB1vsTsAuikR2uX9yXiKGgkV
zGzjhwF0toMsoH+KtiE7sQ3zbgvC3beHNTuEkxsdXiVavuu29zD5SFJcnD7EGvZU408rbUUhbOx+
2ptflboP4N434rWCT0X/jH2IpofLPOyOVyqx9ZrdaqcjmBZhA7Coir71xcFykdD3YTa5AjrCt/2w
dR8ADNhb6DTd4GuWyMf2zzuOrN4tGXIttJDJ8EcGZ6ZOpntk9X/N61YYaCT2aUvjfdLmHpWXJtDz
da4OZM1ZicKdhSXsOrBCFhdU/Kc85HIcRzal0C5YfOvKS5EjWuckbCCrsAFTdolUDF/yqKDpooj/
w6yhiSw/8/ar0jq45dOD/o7fQyXjxDlrhGzvGf0f+WGOC519f+txkAttpsInF/z1xZ4Cyg4qtCb6
iXc/br7hSIPQgPBm1y/KAGPyHztZHqjZs6Vm4oLAZs185HrTRiOXz4HIkt4iwTGjm7RLRNS/1qd+
4cdS+f1EQWrJipiQRmBbOKKL1sMDv/cWq9OmW3mKl8R7vEyUGH9rddYI3eDoTUP0DMSBioxKR9A4
GLDnVsuxQPwCoaE9UKqRJELvzsfo2nCe5o7zkz7HTBJ0EqpxP8SnfwbVIzti/ajyCAkdtzUknrhi
oyFHNAqiUpbwA/fgwQ2hQzjf2xo4dGahoK8ykEerV2yvNq6jqZZM9i+SbWtN+E3GgcBewAFPG/oh
wxQOwrAUClH4mprETCl9aZgIzgQmdpB2fCvbEwLJ0aq26fgxPlk0LZJ36ibbw8rRq/UkYWj4ZCC7
SEUdyTnULQu9bEEWK/3niHutO6C/WPz7zTm8SgbagHKTWSOl/uGihI1oUjkQjw8ePHouAQBPLme4
QtjYMZdufC8Bi2mOiXw6OnofZA21076S3ekkTnjS6j2JxNdeKzZmHce/f5Y8xT/Pc813G7fVujlH
1gsm3H1LzkdpNA7FAApRm1bEtCNizBdMyX55VzR4sBlQmWTengws616oKfBq6B32UqDZPycUUMtp
kO2vJnHkra31WaVBAdb8pD1Z2MnBU/kYEoBtjGLsWRhNh7ZplH7W4E0IyjJPSVXbRBKrKd9VVdkt
4QnFbG37/VPIGpHhAAC/f3ijrGsXXMB+Z/A+JLpL3TiQqqCE/Ub0EK1ZZF0phWRhrQFo8zuiApOf
1cbBA6nk7/Ox6B5iQ0TdOiDfkFNea+V1WJT3qTcbdTyomenvd73eLgbNEmEuG3PoDc+9SD4pdGQq
3T3y9uz4wFV27GRiAZGeq8bzT0fzTRuKD0e2fFFjAFSfj+M/TbZRXhVZBhde868wz8p295Tcnf9o
NRwsQiKlXYAB8pT4GiE0w642fjXe3AeG+NzwFKcu0TE/KCgwPrG5iTKPxP4MyV+efIfdsfbnbeSQ
fVp4FU4pp7ME9Qh92KaudOXj0F2doLEGj/NwWpqQgureyagDcqUwtc6fO4hPyqIp2Mtlv6xeU5iN
Znpeu76wFZgUiYEGhZs2ySknzQpW1nWcDDJNqraqD4SjPlM8dhDPKByvE1FzalqQBh3ZeZT/p3XE
nwUtBq/KI8rp/GehTrtL3+r35H7eg42hJCcP/mdszmUChKS/LLgk4vr94akkgh1zvvvtR7PCBDRy
x7xBOcSaWsVuQTlAJMsyYGAnD/IXBaIhcy6u5gRwMSmdiIkipfs6gfYaMU/pTLfqU4UCqerMQtHQ
CZ9UmCOzW0Ya1X0H/4hvkLce+Fy6UGCeHMka0kLxwFR6rMd9huDJaMrLYe089VRmNaKr9REuEeLK
sSDayBzw5/Zgi7ks7xOtGB5ARR4f9+PrjwFQ5YqxjeANSOrI8BV7TsMC1ITxNTDlI8EI2EvhTzF4
b/cCYA7RAmIQJp+IwMobgnPKCeUbOdeIlEiCgZ19hKlXhJUR7BrX2va1X03+8hKQpCDZXx4HbQ6j
bLpT5hnoBJXc8a6t4OwADUGAoIWk+FJ+1ylmWcX2YOFEzWDFer+mvEEJOCVwLL9Ws4mdu58WH/Ja
pqDzYgiiupNVPYdDDx/Y9veF+k+m79+n1vqnhUcLorRQ8Y2m+za1u18g60+lPC3dasbkP1FKda6r
NljPBXFRtHakp30YMIEW8KJih1ml39QXE/M+lIl2Jc898bk2SccUxfS5mJNhmqhM7ZzI7OnhyHig
heIJZxv5zIpJtWGfCg6Yt1P7OC/IUJoy+LvpHRm26Qa7KAsV5u8/IUmmMApquPf7wyGQNdlRSIVK
QyopsIGOO1G1kwseTnKBQzw3yZINaCFahfxFAQiW+OeVGHRq/M1P08cCzXUuYAzAiEvl84Q84NWN
HClwm/fXYpHrIJZw5FsPKgQF6BdYRsbHFQjDIaobCab9cFiVmGbjd9+7EMsB4TFw4l3EISMcZZeR
aa9o3gaEBNGhfyZXvhb3Vx7Tc/vmOrMGC043Utgm8faFXQMuv3h31qG6W9x6RgCb60zf+jyaIOgz
okWd9yvyeAaEPl1vp5oNBVpKsooyJ44ZULAmqiBU/QBUX1d/ZhNmA91A68aoUaEG3c56aAMvWQjt
YK6X6sRkEt/43zPHcHEqqr3LWVbi7Tk3web3NBywnd4Y5b5VE2Tz1PjUClhTSfqaeC2r7mH2CgH+
n3JANk+vY/cqfLgkbwP5NlTf1BHYpKHZ0oJ0iHFTzEb+lXGZbtvjGAwLV0QqWgpbAL9O0hci6Z5V
oSUjaOxhoDeV2OggWs4/0LpQmtDyLT4MHa85OhhNQf+j6YMyxkZmO0GfF0kH2qUt6OXwbMwQnXAv
ZR0SGHSXrwCYAvmL9bVFuNBkLNibMDpjBEFuolhJazUg9LQGp+eqtTuUm8LjljUnn9VGr4feXjl+
AaiKpYoSt9bRbQXGcSaUG2sv3zOkw6ShSxXotPHZrvG0rPm/+0oxTAMMPoRE08hqY6MXK7vhHCS2
MNJEd7ZhevaRx4qpVRqQvO6JNrvZSiRF+Y+jjbaDol68PGkfoYRYQif98Fsmh4MZZwHHfvWPibn/
RD1ul0WXlb5HKryCT519eXEo17ReHNPt51inNzIfHnivoswdgLVuDz2XaHy7iZQyagsSfPhfYcPt
FzHbA4hkOS5wuEjktIwFUXI5/H0cGZDoNxXbH5+oU1onPaGmRFJIQ3aiftOrNkX8kykfGZxqF2i0
aqY8i9uEWqu4IAIuYOq3bz/9F98reOLErP+lsY1WuZ0Vz+h57YmBctzaC/x4/x6QqhztzAnmg2lI
zwcamHh69hJuFmJSK4hslVfHExFdHSAMymOpUeDVVsyXpEkHH2iZtsfJZLtbdBaBNUfy+ub8Lhji
yMAtKONDS/jFdWpHGXj0U6TtWMptVj9y8+Lizq5c1dVeAysnmGT6n59fp58KrrTz02rDX03l7zCS
ixi+DhtHHdibhe5ELtbnUuTPtykfOLs9OYjVZdq+xhWik9AI0/xY7++A1Df2cLxEa+LA4XIme8hB
SvrrK2E7XRSFL/WIYqsXqE1tVOsjf2mRGs/hR7/FQzRdo1suFNzKpItbVTWJ8gSabNlPeA6i6GOH
GHabL3Tkg6zCd89LGUX7tYPo2mo49Kh5TbA+UZw07GE9XnxKgJ4Pk5hpFfa1HiORNOipoYFDPX7s
So+I8Zqc6Y9Pb7V/U4ASqsytSwumjNRuUxq8Ve3WRFFqiqi/AdmxsJB294VneemMGyMrs2sxCmDI
wIY/0CV63A5d8dw6wO6GA0E9uX1pm+gFtVlVtKDFfegjMP5JLNJ3QxMuSqqlSPzSMLNvHJEFrbYT
Dj1m1PLDTk3did3oWduS4X+x832ylhS05FdJnRUyexGChi0izeBwMXtafsaaJdOdm1R55fzkjkuG
A5svp+a//Y+TvylJf1EPS84jWoj3qoOwI5eeFB5WlsfCl65JlvBjWyBFbfg8IF/WbtIW7jM6M493
OXL5l/LAeXfdVWk1laHc2KUiLZEp9P9UcHXC3/sYBf7K9z7zf8iFtiSwsf7082Z9aSF5bbkgjsMy
SThC97/Cb+xDQdL4eilJ9H73u9LDVj+HeMNfnoZI/qD/iPAUfYMPo8UkFYIJBRXC1UnCWVHdet7A
KeEgK3c0UMRzgajdLvfe05up8hqMoTMfQ1ZEFM9DOjWD3qL27IYr+6jkO6mbsskn1tBWJuA9Ji+g
S3gi+olg/y4wdn/2bMbiwxSYKkBrENOIcMc6ezWuobhbvLbpVrzdES1qks2w2uhqQvOXdg4XvRuG
cWUiY8uXV4a7mTmib/mzmYv425jklgubTXEJz1LXnJRGrNkMs5QUzlHmne7v0IqFni3eeDDCXQRZ
2AtvwHy/gPWzU8yXKB43C1B/htwMWKUhb3rCht3BSfKUOmjUtf5bS8gvsxksY9MdiBq9EvFDTm+U
SnYxMZTd+l4k65qMCO9+WHi/fLVM7dILZc8Ya2RT2xaSpdTBUm3xYYw0evIRySW3bLsXQPxPT6+b
t09MER+uJeY3N54QRe+WpSrDIqzA0eyJZ/ecUqj1rIQiBJlOsmjrruBBP+yRivPqrTO4HTzUHLuQ
rwFYuXWHA6uHIt9Tij3IQTnS1Qqm8j5SbgrcGCD3AvJIS3/Rfn7FUDEK0EAgdzOeJuMUwOl9KegE
BiCz8ZYHfilx/aUTJIcwH1D0IVrSGX8acS4RVlk+pW1nxduEpNqDwfGev+ybJQI4imFfdDn8Pcza
3ufsgM8ck9HzxfJjYGbSRxv/9kdoBfgRzBmYCMQqH19aJthG7hdkAhnYyEzIQc1lHvQgULyQaJ7Y
hTyhsHN5tn8qkW1C9vszRLBbWty41EJNySljcCRxF479jy11YDwGBaZRRWhiQ920r8bk1/RpuDKE
GDcADe058D5psXz+uEPVpJdmvh9X3dn4dDdvxp3pPf9vBaIfWl0XuLWftw3cmswvAirpHzptqAGz
gmDMa6GPbwKNqjhRwyYFfshMqWgIKke6lWCOVojHwkJX9kXf+ayS+wdWB7PCkilcJUHArrN1Neb2
0MHfIwSg7qfQSB/ThwXiSVf4P2pbVThfhT/uU+5HXedGXuGrhBqPNMGpT1Ws8RW38n0LzmaaVihm
pThu1UEHYTDVTfVorzi8GdT1JtwD3O8TrSqtbU1nyOFOdaln6mqbiaB6ZcfT3bPFx67NW+O4J/Vz
WWLlRQCYU0je5+zFD8BobDmtCE0roJCd49tL8EsR1kEv37AON6T3g5IzqCOPQl240/ozzejvG7cV
fkKfDxY7B4HkyU4uaixi+AQ++9+CpromW0irVCrycwUzQf3HwfcbqM9z4eWHMY76EN9KFlpf1wXi
wV+1TSwU7KqeGMvgVVIUd6NTQYsZ87ff7Df+3qICfWRoKR+lk5SfVt5uDpWBg0ock2mI7dTCj7tN
W8wmCZR8RQ/XuJdql5QjbwULOzie5aZxS8cOQfzuRR0xF9Cc22ATJAzQlHYxEecpv5Qlf+MZzUUP
DtM4z5MWFlm5J2eswowSUhTmB3JUEFQpIjb8QzQxjAGI3IycwTgJLNppjnZGqGMquiZXphEtPOcR
8xyng4GoBxWFhDZIE65+qtsnhohiS+kxNBo6kK2g8BMkS6zOhK69eXdKfpR1+WocZf68/fOy6Qcg
EMyXWypFJ5iEgYlqlzvGDocrfLIX/0cooz78GIe4LpXCxoufLyM/dhVrXsGJikptRj2BZBFsORc9
sJ4/59wlxaxfoavKKp1F3Lok2DKudsoo2Be6SUUv/UBjIozPAb45kc3I5Fl3cDt6mwLRX1r5+nTb
fhfyndz/LgIfg0o45eyzP6EoRO1P0B3oVgBHF4kAcFMPrjM3683tFQwm4v/0bowdKwsNTq9CnTSs
CfpY2Oe9IOLVijehfrjnPgia9hGiDeyb1McGjoRzf1t/3bvLf1FkYs6fLlJA+12dQAiVL77aQrQs
jm9UNocdYS+AmSr7EzMC8ApLZsQOZtnxtaoJWPyDe5gbD96A95ZpV8EkWoofK94tu3N3aXHGUxOa
yu/UVGTVLz7Ou8xRSn3fZ5WflrueZpA8vQ9Pmay7F3t3vEk/bjyC1+eVCKRPYA1y7WhqG8knwzh2
5ItOr0ntjDWvkArUH+BHum7DEHy8yMLAtjNXZY8eXoAoL6dPXx7uJNalV1xsPPRwZhb2Cc7iJIxp
s4e72o+4KM7i7chfuSdzUeR2lhcnzEtWaIQkD9d2KBudRv7R4LyXi79VrXJkJjeq/7pZAInRkCo9
VlikOzajlOiGbaVLRRBddkMmgjEnZ2TO3rTO7bEfvQu+1UBcn0WDiSagOZ+e4qhsKyNzpYxawgg5
K6mz7bfvfiMULI7t4WCIIC9QsL4LqxqEEVwPK5NwAzvPGNIL6/tf6FSEdlxu02kJeeRf9aC9DaOS
Yf3IKZxWEuGlQIR1GASQzuip3i4MXEU9/vYs8DbqaWoammENieH2qfauSHJ4GrXpBOMT1W/YvNFs
c/7FDywjyTspxCRlIuQ6EomDLFbrW/j+Ml3aExOzbW7p7lREEYxrSHv4zAj+xvPmWl6saE/IHxCt
0YEBbPMUun2W+2J445cl43knDLBlrlNHPfYf0Hp0zi7kHSimVDHnXOgr8DODBjPDiwlZE2yHnm7K
PkyiKgnN6VclwNc19FnB1+UM6vDvgsP00SpvS0mfu9QBm5tKJqPGXEWgNOSJeUMpHywKVx6l3Plq
XuLu8VJAo7iosG5esmmzbcasjyG0qs5oYc5iKP0dzEl4GSQ+bBU/H7EUPkQYGJBLrkmWJ0FCQ1l6
fO2U96Jd9kzKN4XL+ZqT1o9pyOaE+Tyigdhpiscqh83S2tv3sufMYrEzE8StUlDHgx/22EZHNBKm
ZJ6qqibQoItKAx/6/ge4saVeA/IlIC4aPSUr68o417IN3f3F15fDORI9ErWmhOgMQ1yCmglQ4sc3
iluhwRKWpS5+4CcWkuuFJ1trjkGINjHJyyGFJnlYRQVZkXakDHPov2n8WY9FwjfeXVKI78Bd+Hqs
RsFApT1acbXL1lntmB8l7YvhvNtxfHd2VkXT3VJTbn88XY4/YovwgDXela/WhIifJP0CzY2CQfIB
/fWDEWpXy03JpiMQ0YuqrHRozOSa4CyotpVS8wpIsFuA2fW6qfbgbL7jp+/jV9wDIoqGXlfigqFv
8htauke9P4+IZsyqVfBuqcg+qA4VJjw6yaTVRKRfLQ1/2f+8L50UrjSvm1KlaOe7ULCFKi4zROQE
IoCSrY7qVr6PQ4hQ5hh1h8y9uVQpP0fwlCMn6ZysQdEjrawg81Pwm1+XjQhMwmAawHcWxCMEKX4R
sLo5HzrUB6/p4dZzRx4Gp4+DiHEWHKw56poOCtAroOU6X1Pwv1mUTEkecx3Y027jt1IAfCj0Czlz
q7TzLeX1Gp/0U4UGg0X9DFohYMGgBOm0yQb06w77yTouvkb7OYGbgb6u2gOKWXqZADXiOBmMMLFS
4DnQ11jUO1U6gORFC2n7RV6PYVUix4i9Zfw/+UAsQYYL5qnP1YJld2fzXT6qbZLsTc0WHYiVBx6+
G0EQ/6RouP0XRwdqVXqa1ApZ1oK4DBYc2ZyCQJA3oMZrrMvCcRtDje4/vo9m4l5wQHORY/K91nQE
eEpOkX2OseRejZ6bA1GGnY/QI23YkA5C0WteG+CmPLmW5pxKrgZz+UEk2KMYMXjKeuJQAQRZ8+q8
FMXv39ZkKsKqdxI4gOXcp7tpDQCcQT/aEGKj0yzRZ4jfD+/j0pZ51dKtEBHBMvb/3GgOe++/W1Yr
f0tqx4WTS9wxv9cuqxPud+K2gciAJ6u8KYcZ2K8W0mW2fGHz6cZ7PKEEfG3G5AlBe3Ase7iZRHwE
echkoon05KUXqZcwnZutJg46GWjoeORuXOG9dboVOAIFq3RZLsP549rp2gjQx+ZrMDbnjk3WSkHA
SmjT1Db3YiPtnhP5rhqlp4Mn9UDyq5JGyWFLiGmIV4ZZ/ktfJiTix0ZVbu/Q7U647xOZMPiszJQm
SjDWop30eJD/8fhBIA1D0+sC5AIEF6KZdTbv8Gi5dNu4S7G2QjRRrmndkbSzGWeAD90pLFANS/CQ
w6cZQvdNnAJE+PugW36xMweKhYxPc60dOQMoM2acuhbGkpr/X37whZPoV1QytD43Fsw7kvR9PoiU
CCGJjK59/ixANIyIOVXye2efXd0y1Ho6XNh8pjrefAJUlsywxDSDj00CGUA9zswR6I/Xm8ynPqeo
b/H0/ugdXjDRP/q3DmhUZXAvxgMn+Nd9qb+MR9cektMzJ8PpbFAA1Fm2ZbVDZCGrR1Un0y6FlDPe
JsttMpRmESxmNf3pzSLCxvGRJ7LTNW5Xw8WjmlrVLAZifubXn3SXbG5lnoopGf7wShbmfYTgYPiv
BlE73UpU9kaQ0KHbLpxpF1yUfkzf9X4D7Ph69T/Gk1gCmlr3EzfT2xIjaChoLJnPCQQvLGSejMWh
Yd2MBqOjICuIfS6ZeArqgAAu8Tn5RzViMu6lQWsDXwK769jXs8TNTpYw9thi8wkNQPJbOqNH5mK9
SSt4Yxk7KbIlMZt8PQvHjY67H+z9XUMTttfUTnEpuz1OP/OKTGBWczosCIHhumvVj8+Gu1/HE/3q
zFiUwOKGD/AIsp7jbU5Vox93LrbsSiZ7V6IoVL5GiI5guvOZ/XpkAbhV8KLFAQiLTMrdRHTa+FTD
8moj0Zh0n7XZv9qbMe2uNUXaymuVVkKhe+SFpZduc1iH5PTeZ0lAOxQRNK/BMoJH8WIemmnfNKzZ
YGP/W6Soc8WDI4F/SLUyS8jn4Nzm8S+njisnfS/X55g3fwPkSHWDf4G6v3mdkxfqYfOBzIQDdN75
ln8Jbw9y7HakA0dab67vewE7i6uDQ/4BIpWKnMRnGyCUjM/DJx4QvA0yfNRYaagc1COZtraDZvhE
C3n+tpxPmxUwCY6ILmKvEs5sSU+ozVHbNlOE3NwWQ6tUsLz6h4rJqR/X2+XncceIIoNV/chQJ4PU
dCYQWYVhIszuKTY5Mq2smujXDm6G2PSNGcyVzN+VX9769dzaKD2u26HW/+Mngcn1aRyV5ESl2ISV
R1aEWP1aBEckH6Eyji9jcxttblzA4luiSFvN63xOMRMyfUmrK/HReORreoMq9Ii7ND7qviWWxjbS
ZYOYBWeC4oWWOYcAQfkFcEtkCpG9A8Ey1Qmi4lTaiPFs1L1QtOwrHKm4G2vPWXCBaW2+axcSdzW3
pm8wJ8dMCnyKGPhr448LQPFyHvzwNlNcvYDB5FZ18vIYB7gCaJydmzgBq5i7vjkQTO9zmO/20hV2
N1rVwhDDIdSHDYmt5PAZwpuGeVLbOPiTSeLJvN9z9Ir+YiVCwABs05glQOGYf/VtyLNLIUYi+hsk
ZQa8fj4eO+KndMQofOS8zUrjZqIpuwRh9dE4RMEsH3N7T8YG/N+U34w0f1t5qzkzpM78JvmJ7ZoM
+Cp5QdNAncybFw6hpm8acxUfcdGSIZsVtLJNfYFRD4NBb9n6pbveXWDt2fj4Xr2kWxzku2wEZ4ei
mlrf+lfqCvdZKbgnQ94wEtitf0ptMK988V3M66Fl0EX0TjZ8GfoMf9C9go6CrytoKIlWvSWedsYL
6E4RZT6VgvP43ogSSaN53D4cNh3P1Nd+Qx/poKqwkRLZlUM5w+5jYySKFB/UV80COdrrnGpQvBU/
Oj+9ki6+XJ/M/cGYMhQuuG4VCdJ5scJSfn33Vl1+bvQhGE/SaQvQNEe06IKV9uHpyhHq9tYaIjI1
v1ZFtOmzMcZk2LJ11tz8W94Vdm0WXoPx1tVdIZydbXS0FiH1dkY0F69uWC3mGXu1B2KWjXNyWMNo
7mqyPuA9TzTbbUfw5lhkmDv/iVLKd9NJ2XT0tWbgJKrHXT3VjjkmZp4NKLgERdM+LwfgF7+JmzCD
QLh9jOwr64unU7gGeOjzXUpohe6rVYd/gVTjt+v5Ip8uDYQgG/fsbGpcP1M1itq/RjNDuvP6K0+i
H0h4xQcXj4IcLltDpOV9DHPVdoKK6pjp3nhadhrUQpYYbj0P0zWzgjgTrVON+nDP/upfPP3a3pUZ
VkQxaFHBNdohhArVGvrMNGp9WJG3v3n7mvRLKNkYwjWRNYxKPlJBiMkYGFdtrkNkFf8uvzBYovTK
PEzqPTSfLojHV6SkEb5ob6TnOEe3dxtKmrfo64lFSUlgaFUJpL97Bvs+oxa0ifiKPE6v9jS3Xa+L
XpoAPLclFqooajuUI8SYYsCSxmy0y4cy4No5Wdc8yjJdMve0A5CV4s6sWeFq+3Hs00QyryMcyZ5f
gfvkwnYAfDA8GBOQsykiQk8wh+ENmC5d2KEuUrfu7bW49OGbtzMxf++jWUKNx6SaDdhrCepSmxMi
LCNBFh7G3BajKPnyOWoFAdaEBNcZhkIebwPeQ9LrAdvRMYBt69UY8pHXhUD9KBOHeI1p+zmmo7QM
HhoVWCGXg+hrl7VFlA+LvnA9ml8capwIj4qApqb674Yp0d5BX4kY9OQp4wiMm2Toe4LKDbZaDK0S
P3P4T/OHSFDyhz29uLERcV9/l/HMfffaG33Mngjhj0HWYNH0DXKONF7OurDcvLjgP0qM3WRU3gxb
SiZaJZrNVbhTd5W4d4/7qHy48kev9oJtuxrOOrP+TCz4SyVJ6bcs7or1M+IE6RnviP1S9YDnOvgA
Sh95qD8/hoDRtgsK1FvGVPce6N9X94k5JQWBcgimOtEWt1WvrRUa5aW+/xdNo9iF0p1KLzV3It1J
YBb/VHIILHN2YYMgk0RAvPrVcNY0iKrIYbadtPIEoQW9cKTk3QXMYKEnIq3LsAeK5flDbN3q0I63
4MVTNCGlReFlp4klb+ylEHOSpavA0sd/qSd6VyI9IVdQ8eYb5X+m3Ems7GBXYuMeGqmK17jaqFn6
WAmtgvcQwdKKq/ZXGcDdA0xnVGCgLFSIJdTD7/n14hIgKmfWlktME1FGL2/KNVx3jB9IXZPxsL4G
/E+/qGa9cAdP1eBuVSlSqRcISnJsr6LI/eWaFALEGS+d2819NPlBkSr8o/xZ3WzD79C/jXRVknA2
5OaDBi+gdM99aV3BJonsvmiLk6vRqLRaNi+Fj2BME0Wp48zCaENV0TVZUyk1RHaEZYlufzvQr+9a
1l32dArasQ4cv+evBwVnkiUTbQEEAQi/0Rpc9PeUUJ4T3eLbFOpNu+5dSbZkHipWXqKoRU/JrNJQ
aulXKxiZhkDMtA3y/HWhblPYDmC8TN0mHRmKI+9mBn0SjjAFUtsiFtr3geC1JwgZLxbBiSpvAZNh
3CY6Ym4tuEyqggHIM0P/CKzwnRNK8OlB0EPC4VctJ8EHYvDagjl8I2XAv0ziUeEQfmQS65a6hwcZ
h+8/dV2laodBsjsd81MHLJHmcskhm4IIz933IHbLjitCEeOF/KvoUc0QN/AA6WT9oURxAYBlWI0w
WKE45UZ2crF7xkZEx54A8hQfv81dqJN6Lr3scfb6n653+JFsctjL314BRQg/CmdeW+lMqdwXJXHA
KfkCkBo/0aE4Pa/JDxiJy28KNokxSeNngojF0KRW51ixh0IdWS1TUamLKtf3vK8H1ZkUsw8rHWet
j9DZEteu/Z2q0kTa10EcGoW7+AFzOI2rFZoIbX7hPkGh7iINEhmvVgDNZxi9nwXm+xTqoPD4wHE7
oRae60OCFY3KTOicHt9FZN1Mx237Nt1BUAgvqSztUt8ZP5IW5PClAJD+NwgApgjD32dt0smdS9I1
CW/+Ce65URVQap4ic4S8AyaExLLIVZwPYrENJHVtoKCj3SKzIRY40+MV6PGkSgXLuW6jaUPDGrZ2
ldUCxCf7ZNEcSpsehTLG1/UX6/O752tPnuze3IBYpoLCx3imNpHnKCl5WTYXzRP2Z/iL3brJvvj1
rVjjxjPzKqksP4bUlRTPHIziJJelI+iRF2DXBkFldjDhVemONbqK1uZwMNQ0n5pIPfy/L/QC25wa
Wdr3XewwBFz+/R0t2/Gcma0cpjti9c3PIxoYYNOGAhuDHPPLUWkwn4MZfF0zK03MFXE1KVi9qLyx
dTmZHzNcBI7M9310I9v8oAXXLc/1SlLnkBfnTFfBTJGosKN2bBPpU563eBaidRhwmkHKBTpd7eAD
nAAr7mlJnvPNNTEmswt2iZHSRTbQrGwfXjfvYoMNNHtXIclF5bWKqqHZwlx/sZUspIpdK+oR90R3
Qwy4QJxGz0wtXB/6XELpQ9Z/PNs5W5TxPqYDW7SnwqmOojdBsB54kiy+vy0FOom2LrjjMpdhjs5m
Dg4HQZm4r++JLWpZ9npG8HJ7Euar+BzsvnTMIeg08JdUQ76lTt8KngWtaQweePmOgNpz2j1km/p8
cHSXN8b5VWyDLPkVay+tf/zQcyaM8JVSSo/a1lcrV7DmxlcOyKS2vovzei7Y5ihSPOEAKpahzSHe
nQhuVhRoHialirz0G1nYQAVtGBQOx45nkoCxYvvXdb8Ritf9k0wZj0UHrQ4Zix0KAdM0B9OYrKyT
xHoTBK+NhcMBmJlUUX5nH2zX9SM9MmYjJeXQSdU1g4qaIyGoZDfVm1sbUdfuz3sksaguaA8pLBXv
Cx8BAlHiiU4MAUkQ/7Mqhg2frgsB4LAZixxeNEO+iNUNQ9tGHDW+veGUD2HCqV2KeKERTRznl3li
yXO/LLVeV5Fug3sNDRsgL+dtUam9iPy6RcvJA3wbRYRQzEMt18zq8Zn47hbldNOXMCjxy7PI7u7L
T9mvI/eORh6JvTDO0a4A63eTjqF0ThFNTMI92T2+pWYJhLdQYS1M6IEtQCShVAJceQegrWdFPgRD
XRN+yeBwZpL1U5Febtou7Ye0uN8MdqodZb8QY+HmqcGPQpiheaUz7I3i8xgnrQUne+GbkluCVhAf
vrHPCNT3OO375Gy+RuY8rnOGZMJqkUB0CU7ext2Xn59BwYzUE019IvR3tDdpYcunWA+5ieBjLbTV
LiozenkXyQV0Cwwskag4ch/exWMhUN4Wtfu5q7yIWyE8CZRfLg2Ox++LE3fj9gB6Q/KNSptS1ZDa
ecFmrlssLXzgpRyLQjvy1ng8ySQSpmm6Vc4MGCaXW+JYALH2Doip0bByN+qSIs/kO3UC4nU2pLGP
OtFt4xQjtcimjCq7LwVK0GCDW87DbDNajQhm9VVEiEb3c7OovwHg9zXrTDL2IbqA9Y96uGlRboCe
KrJSYQ7qJqhKdyjsq7GqH00fvhLM7/QJOPU2bB45fm7vevZ5auXv/Ns6XkEIzH90QbMJhOWHHujJ
r9b3bdntCuOYnoDS3W0phP/aNwqzSP8bXyvv/69oA2yqveAOpkQ2FzgRLymc9RMd5sRo4IpoRrxz
WI8TvNBhyiM87nZdIvbyvp16A7kgMEJME1lF2HEzCR4ZAWheTiALOlGEIRStd7np/Gc7jzYOfRFN
JPice/ecV3mz6ZJAutAAdd26DJzDuJ4VJeqWAMg69lJTPBqMMTmfFA/CGDJ7c1ldyN5XY04ngUPt
d3XQVLSUX1g0vXRFwRywgMqFH2yIBpK+XdfljSpLA7d57e4+q2diT7Zvtg0xLUrgI4Dsm3ygHUJ5
0YrXp++s18sZHZpGev4PNSeiUqk/Xrv1AGhyyNb7cczd/7vHycyQtSep7ukBoAp+7EM/eKIrU7ei
wDjnBowQqKA84VL8FSUbNsR3DCXz2u+4onwQcCfaEbj9VpTBVodO4NmuziJcPxczYYmMEt8WGbBS
ahHvJFS4Ou3uZEhOFGd2YBfnOCFw7fy/giEyuFHTo2xH+wH2Mf7Hg57dnWl2q8M1VAyMJpWPe5ad
YS41xZQEiG64X26JFHjW9C8iEiD+Jsx1vsCpOTlhw48LMpRAGTSYBJINMecQ5Uj6+qdlZIjCK0pl
di5rbSAsUIhtvwWDpaNAEMG0F0/EQim+HZtXQI/PedQOHnd84CZ17M7Eas0yQjXODKH9mltC8p06
Ia7dRwppd+b4HAB2flPmkz4glHrcgxIsqYboLIG2LDdTAqF3VBMQ8DM75X+wesDDj0i5euMU2DMA
pYWGQm5egQTMv2ySXw2dnfbFmtqlnCJuH9w03t1joYaEv1qFkBwiAwjRpDyd5hMQuXKcKdK4luDl
xFEPyGd180BhZj/IN0oOuF7ozTl3OCXOvJFpHzc/6ksa5hu05yYfADLNJis/Ynz/w3sNg+124rs5
Y90KTwjkul4ZuCYJGNiLAyxZI85Uneunxm21ysRjRLinCdvnZaVJnuLFhn1BOqCqoj9ShuzNw9jb
FsRXLaUCvZvUBp6FBmMoDVcywGOLuVuWKVMmzG0x1cN5soOkXDO8Hzg8wcRuZ95Bz5h5rYMnNb3I
JahoHg/2PZMYXbxZpVujl1grwlxq/lB6LtdfNr73j3C5wdlAB9R3qklqHx5VZAtlGJ0qcnMewf2J
VaTcFCt4SfJsBbqRvAOfRv8SHoAreTqxc3rZPVRkSUNaY42T/RpGTlHJXIwhG5Bo+FN1H4DAP+FA
vdbsNfAdacj95QAocWUbfSbJJJmPgctCqwRUvFjRZYGEUfnXVLZKxKz5RWkenlxaoeSk1C5UGMxJ
nhEp1ns6hBXsdsRb9CJtw3t3BzIjcBpiOPIVG3vPq9fMzzSczi/Akcd8DJDbtVXvHaObzC+1Ajjq
Ep6jBnH+aY7xKtGk4jBO/FQ5hl7DMygWzyw0Nebfgk3pQPemfXn/jgFoZkuwz8wONHyuBfI9CvBY
YoieOprQcENOrX7+PtJB7qR+MZppuZz/KZiRoIowLDlwyyCUPgj2qtHPgTUnxWMOgCoKJ1yQPwrx
dJFFGaG8AZv4ML5qb3KZj9ANKFoN7BPP1TIMQRFVPFQb2ODtebQRg54RahQFGH7+6SEsau9uHi9t
1SZiDiAJImilIHV1c+iZXeqJjB3ekdVn4jkpUSi8t5AO4TZ442LlKUevHi+bG7/xvCzn4FWfzLzk
9fBMgYC9pNlzVnVGW/yAFe4xkyAMGpaoN+kMx6A/3R79x0ph9ynloWqjN8bmYYtsJMHiBex5Tsmd
NhS1AiQkQviLL43SLanRAbrnCagJ/L2Yt1IP42depzijWRqvyNeDDJs8e/WXPJqOuVkho1v8fe3V
THNTFaTvleg9wDCe8AoS0yAH4L+8+lq9Ar5FL7VADVJ09o9EEygZ8vk69iCMahS8jslXwdsH1rlE
ltF2PlDYzTx8X8K8pDLvItZkPEZ5jM4S6pf3GjivGhQxD7rScVX5sXhMWkgXEDg/s8e1q46Ola18
alMT20C4hEp2gl6hXhSio7KmyHF2UWLmCUBQIPE4Tp0NznHZjuAEb7pKYeAPiEDaaUzc15BauKYd
aErZM65XsfkMsX1/QLxbR7kUCmUrd3AnYjahCsjpZwNIDGlEzIwyIM0r2N8H5q5czkJAc59FCzb8
mqJoPNHnc5EF0wTkstxqmtVMDw+0Zr3SRTsld7knz/LMH4c34SLKzLij/HpJJ5Z2jqaIV3lcLQJc
4vBciKkRb6JK0dfK+ePi7IAEvCL+QGC8DzS6Yn4O4qdTJULTfcgQzCwUjIOoRQVLXO/l8iALk2+A
UMswr8Nzxw+vDMIZT2dY0JzO2cTq8glSM7oBXFhgQ5L16t+7lv08cvobK0tQMh7KXcpjE5HumRx/
C+QUwPhwcRPVzhSGfNjvTOUANPnSCsqTaKv+JrpP1iuK6vKtpyDp7f+F/1dcnUoB7Y2zvCOLz/D0
VZ6Y3nRIaNi10/qyuTP8DTLybfPJk3l0+9cuyEwtPqQ1uCAr1nu3dLjYnnpCfmNq3l/hlSaeW/n7
m5bu/09JDURU/WtW3ziWHFNt5agwTuqPsNGDJ9itpkb1Pt3Uy3aSOeENYawzDmTzb1tiW8uehX/6
/bQZTaGAiHRscyqNpkUCd7AaZ7mHUvQkhikag+dXiKWWlRCzkXbteyDFiRI0GRkJU2PKz3Joi8Nn
tfm+wgC/Dc4hUxFBczJkvwMxD9uJUmPDsGVCmBfH84EDZNhb9w6ue2fKB1p3WX8ZcoMCLeVJYYRK
JAn8cThsLM/vfIr1iv5m49aPTZ43LssWJf6AQ3kz/uGBig/7kacWoNquwmWFWIvX06ZA/p6Kzrr8
quMy142VZHa5rLmterEFGhmBZKOrubDQf8BSdXrWllPVK21sd9uRPYRCIz4PrcLmRQ1fDz8QO7GT
6fvPPN93ih2eEa/ooAcZLScJLfPxb/52t6UJrwlJflc0IHWto1K9VcTCqDqE7/THISs3Bm3gaQ+H
4a5wjMK8r3adjUH9dLvTJYRJlF0CDTm/BmGxIbIImEOmFxeA8GWNvL01OUYlI6iJuZvEpNDvudbw
fQZ2J83hBtL3j3vBtv6WdXPglsfaCD+cdIqbsmaAPi+10BIZZ0UkxcRUDa9eZz1PhywSAIF7M3r1
oACDLgdOBbr9UvpNpDqeJnhylASTL92mN25Xf8xEFvSnlz/5rB1lJBLrhmQNvt42MvwRnhoyJaMQ
rEV9c+SZNwHEFvJQlsV2MUPQ+cP83OkkMm7zsNeTWXiztW959FvfFtYxcagcQTq+jn/UnvowmfX3
xGpJ2agWOPvCJ4Wi9mmMl94JSVv159OG/0XugS8AwmeXbaeYHkvGRxYhPdMBELxRq84msVgv422v
O1QRKinmeSFt78TKMs4sDrC5upGG4nrBfsV72AjZYE4y4TccVGnIlGrV9chKIl/T8ptVL7qCqKs8
WKDdNiwLubE34FhjGGWAnL0SKwVKVFJoVQFrl9dZzuv4wgwWSa6WPUsSaZu1sNdvdlRnuTD3QMev
bhSlWcnSiUcIJrZfNOLgo8JUhiXnH1UGZoy6ezEkCaygggw2FyJpWvwdhfA8xW2ePKnOptNEWJbB
1OWslLZbCTa6afLXVxhmH87XN54/LV+Ay+JTl7+MIA6mrkAIEYZFRtMUNty759fJGAsNKrlKMADW
JOjY/bhcHiAtN87JDFI71al4IiabN+a7mSHxQss0p/0SJS2DFHmLHLB/gwVF4eUZz3tEpnpA/PTs
UGymvUTOLPW9bdMPrrbOZ9emQZsVqwUEl18kwj+1zIvQcoKrWv5DHx71O/piuIDkwHW0P4CvufTV
3WL2os1yIFjY38b2RK7fmBz9NxEvYQBg9GvTBol5YqE2UEaqNbBY0dcBTwMxWPIiP8a3DF0NVIJR
fb/9VYm0z0NYTSPtSfaiKD9fydS0VsaA9E4P3xNHJhBoxO5dpQgghONuNyqrVph9gtkVpRQ+yRsP
r6pDZJJkpDPcrDNTkpZ4uDym1CPwj9/zOnpqfAkwWs6+LKX4mL8YSEdqgjcApXnORzqfwfP6kCZk
OXGs4VoAKVkyyytx09JJL0wwYA2WusmfPHLhFIiQaQalB0CIh0pO0hNEHuaMeHqBDJTsfUwKRZGr
f5NRvhjR3Fe3TQ6HMjH7VBNOkcqQ9w77FpX0ggCyPl2hTjkFXcWCQENJ5My4WJV6x/yhYz6wMIU1
Eqx/TyiLNxm6QcAyp/2vo7g/PvtoVFhkb1sv7kMATSWMZhJFyWxESPI9xR0BfLQpoV70ZCw2FyFM
ha8qoME+nKSXAlK0fvv3JB6DKH/jiE3N+jqJT8GCPbLU51XQZ6d7Mzzd8PiIUC1ZCIwS4uhS6dSd
NBLPWa+4oGdq1IjFm0tYYidhU7C6Ul+ygPZUGAf9hBqd8m4vgnAT7qLga/FecSHGBWlQ1qbGZl3x
PftdctahkeDpXqlccvrmuDmYpWXDd+wBN72EG4MnvQRuDMU3sUYUb5y+UkeEPoqzGyW8mBnSaA1s
QjsH+B4/s8oWTpDRm1inKc6/SsHkvtTigXNi8pAWbyZDvamr4rQm14K0R6ovkE/lQWEY6IE71bMw
k96zugvX9gEJaJL+z64zYjeSd/z532HsZRzQM2k2r5kHkMAMEsTRlAaOpbiFlSxcIZ0K2x1qhtHm
k0d06I//qfOggzvEvfPhiudi4tmhKfTHY+ND+JxkU8bu927kVSQ5zL5lTQt4j0m6vu35Ov7oJv2H
MoFgiUgXfGx+9wz/zkGccsXRbs1E76nGy49hMsCHr7FO/iTPG+VBIN0lFACoE64hWFSmHZrTdGc/
EdUsaVr7u0MT3jbX9oE//REgQ96hvZh3qmwiSmdYep2yyqmnaK3PHG1tPNFiy7X0FyTUR6UV80is
NLzEkKTkclqg7bUrhgJuqRj1ozk3POVid1KX7+oOY/Vtp73wT+9+8twwhJHt+VijlL+LqF+HI52o
nVt9GpqbkuiGgGAQPm/zk84SkHuRvksT/HByVr66t6MaW2BxP2UczzG58DBLPcaKposwALSx1BLV
GX6sI6XednUfDBsHHVOrawMYIhY8KopdGnoNAw0sDsn1sHK1lzjFiGatKK0U8rS8SBpcTuQiXeOe
JpzPTWo+ogKZVt0gS8zAM86Oj9zzSjehP+83zBug1qdIZpVlX+JuLm5Keq8t4AqJIEt37wUyKXpt
XAvA8fHWaCVP/wKykA+KJgOBYXSatvBBkWFasHYNCzENaeZgbUblBHJMKBHs0z3WQnARaBwqmR7Q
Yc4TJ05bAPNLD/7uMroobH+pPLVrWdzhIYJ09qLvzwBUvnayuepouYpoBsyD7RaDi39TNF6uPX5B
vpLI6tv884J1lHX9LFDjyhl9HZamz7Y+CsMbSIxSyw77VenRVL5Va4zcajQl7M67+v0G4GVn/GCM
5T9aeEQFZaKLVT7BJFi33mUbSdrSBahOeviUSPLbVGu1g3/O6Ns9peprHgqDMNhBtncUfAobgnxK
wmXQOFTbTeB2dT9d8uxz6hirRj32OGc+86vNhzqEFqOZ+cnR5mqtu9Vv5peq2vN8FaY0BJk4yhPO
mTCD14MlZL2sKw5xU7/4JtxINWsrE/nbuHHJpoP3YUuPxqapzobAqmhUeVEewO4tnOUMa0nQXRLE
TZL1uuUYgEXxwnKNfiEahylpNZxJdqYh9Rur1vBLapGs4oJNmqsPxT0FVVRDPFKA+weOv6PcN6Jr
bS5Ce/qeZ2R3xrrf7nlgkd7VOFDiONaaGLlPK6hljTkEyP2h1/dP0OSLvhXAOL5dS2oBTFnNQi8T
WguGgMEmLm6cY4LXWNWhi3spKDHkbZ+9sWcDMLSJryUGuBweKlF/RDz1p7rxHLqXvgCV6optO63+
2yz/lIRoDgqGGtn4Nrl1zjX6W3GZ4l7Ia0j4TJqb6Cxo2yvecIYbZyjfP2ZruyIO/xehs9s+JzxB
4OGl3PQw/gxeZ6T5p0Xa5RAzwE2WMzXFp+YFjyaDIcYgjSanulxe6xoTyCBFG36lov16QW8l6HaE
vT1nQ/30aReNipH72SQ/AByol2iLu8/beAYn7Wz5A/8iRsjlW6zCkuySaStxJiCLrA4UVvhkYL6m
15XL/z2iX7uFJ9MGJdseOclA3V22SkKnHCiMa8TOlAgIipNAEIIiitYl99H/fWug2N75KHgnaLpH
4OaNhmZIdQgiABQL6DF1zDAdeDn8puDFYDoKYrB5g524J5ldOZ1wUohRjcvb0BUpopNNl5bwVfux
PCzLMeybTmlVMnZO+tMolgyYYi/mMHsuc6fUAsO5y5dGlc3S5Wo1dVz2wwlwtXzoHz9Smem5epg5
ppdv9T499OR3OsiqqtlMwS76f5Ftz7n+SJ/YdFvG75Tyh6OWlti1wi7/rzJdo5doSG1JraQz3F8F
A6XRRqAVlhodUx5+k7m+mj59Q+FzmvviAHwCiqlM6O6Dg7He4z/Hz4rtWOU8yTQA3PICjoX+gLnc
U5AgBZ0xer4e33aJmyLI+3XiQ/Mad0V3wlRx/wFAPDNmfanHBtaH+WkzdI4IVnRPM02SCgZqqhPj
Ai0uxzn/yOgyY6SRX6rIT62flYgpGrTM4FoNtfe9PY7hPVWjj/sa9mhuMMa/5K6RsKI/Uzm4uLUT
3UrQA6V4pvTnJ+3bxvn3nMPfEuBFb2N+GQ3aztLBF+DGr42mYq+pjtIv4LqS8XOQ0tO/jfEfPAuF
FwRkn3bOBZkowlKdBdM40Z83dHmTE974j/rbSvo87bgOSKCHhkn6ui1lauwGXvZPZSKLh4DR2scQ
SwKTd21oRFZwUqvBddahEvlUcu7e52pG2W7OwpyICeM35xJyQyFE6QdyZsDjT7Cbu/yN2yMMOmf6
dVxZJRQDWi+trdngbXnPXf5gYtg76F/+WFMqYXUXW+0Wc6iV/m/wbhzcMMiWGq1V9pe5C2mTXwEJ
0VRfbosR5pa5409MhbbGtXNBQuh2I5k1NiytS9aiTH2Gboa1rFtTDOt6uaJgqW52bJ4EI/SfUnHf
dDnc2GSiuNOdALKa0HnuTzalDEwMHRb2FpzylV6m0I6EF2S59txsxNyEdAPreKCvKz9bbTFGcBbC
92A96+VqZzXirmENDcpvhXHFNiuKnhDPCcovgoPYX4y6l7x0KXBwLnnQ9cx3Sr+8Srz40GsMxqHu
NSzJw1Hkr7KcOrtwxptuVwPyxlTnCNdm2Z30AEQ/f3eHBPvovqdE2EYC7hRnyDzqJCEefTQ2XdsF
Z5ypnqn+/yntZrMaTNC5fiNIrzv0xSPRC25yDVaSxZXu6IE6shDBgnOqLSfnaEmu7fB1wA7imIoT
sKJXjbwrRFLYyQLGZmu5GytnbBIxSevLX7jKJM1rxrayRkcRXDmbAKc/b93AO09KsCW2eZhT0vp1
wUdNpRUsyCms6W3lAzp6TdVp4tMHT2sSNTrM5PAv6EEJcSjXM6jX2K48D081qb9R0ntj+zP/Ephd
qGMiTlXCEJwSlcd6d+9U0Xltc0CX9tjuVB42BXk6TU/ORT1un9i0fys6hYV8iTRGRLwk8FKuzZed
MYkkkoMZ4drgrwM4H+7GcCKlw3WpkVBvvfNio7S8jzVFOz54G/4LRSftgkOJ9469cYivFaHXK5Tp
uDe9uYcsHI/0rWoS06XrPUQ79TK4n1SGNBXKn5k5qju29IlZ5Ogt5gsklEZu2W2fUkGQXirAhgEm
FHcmgC86phSTZ1UzI6PfjOoQ0Q1N1mKbmQG8+tPrmYdY3tgCQ+wZKS7OK62aTh5M+ZdlBeQ8aL0k
HcIuHoCXY8HNfxpZu+aPkHvezaURCXB9+igpE5kdTOJkRSAabBH8KaERXGhGLejOK9GXVrk6N3wl
mpXTd4X/5GvS/4UC1Y41D0QSCoqTnUE2V6NFHk5Zpzt66LRphDIoTN0WhnUTINgTdwNoI9qRKzxf
g5Zo5NI05jo5Pcatwwc6Jtptg5xKVxEmapgWZwoYe15NJvjG3ooIa+Yaz6TRk/DkJddqe5nGOOcy
bOmjXBRqOZ5qmgVqO71ZC9pVAxx7qPrK0RSP7y13MLZ+VyEA/WsZmqhF1lHf1VW+M16SzmjRs+eC
qx8ChGBIe1rnQDoJ/MnSfb0yhcqb60Zo1TkHgYEF/emSbRjwdGHl2I24U6Dn2BkZYraaCe1jyAGH
LZG2o+eHzBFC2y36hzUaKNgEEwH3FzGKSX4T4WuDaVPQSTATkfsV9XicDcOhFJ570DReanjtJDDZ
X6Thr4bBTwda0D5jl5CfjDUJJzZoZ5m+HvD0nFNtZniJ06F65AYzIaq/T1LqUxRhfpdN9i1mSZ6D
/Ng6WkC6df8NvZF8nUEMNK+i0eeDIVIjXcUWJHLdaUb/QNRcK3JGPmvCZ/aca8l62e6rG6O2wUfX
DDciR+RsxKKA8FByFJPWwlCjmnF6KqDlhVyZ0PfrTVsBmn7vcOrhX1Qk/6Gg7HMhwYZdsCFCWuqo
P2/mGAi65Zywwd4eE+GMWE8OkHaWBoXYqS2+P9PSXzbklm5abBGNZ+8+IKaj04tPXRHHTVjWwpc9
JW6AzJ5GCIh7KauVhJhhOXgtxIrFU9Diq0VynOFRLQmHf7tnqEd5k7DgEkt552diNtJYub44MNrm
y6IfBPFbUDWG/o9MVwE27xV8rdCtDYOhMo13Xdl5ZU2En7gNA6v1WJunobVLxi7StNLCpOhFcJWT
tlJG4NQLJ+GiPdESP+N97H5UGWh5+0wTqKUvF2MkNVoSotcJDUJE+kFfL1WO09zhNA0M8a0fsGtT
feHccAiVtiNMdKrDUTGivQAVvxvPtU1rYUCUHLozwgM/zy3exba8ROSmJxMsM0BlTcjgp1FccNMw
3d3hvGrjDONXW5UCNuDF3dHHlbnf0431MRk9Q4AFgwTnYoNviOknrxJH0+JXC550xxN1ctnv/KZV
SBVZ5/4r8VBIt3y+pGFK09hJfoBhk5QUb5SDmd/8FtklCkfJ0AEYBDLamnSkCeEwmypnbOQdvUJF
CNnCzXBbmLOUDI+BQ863FyAr0toy8JO+99QSdUVe5l3r9QR5GUZLSP3fBQiG1DZ96OiBDK9btbdh
23M10keOxD4HX910eSEc6la6oqjcDOD3a7+AAD7KBbSZXC65uSjOy9c+a2RaYM+MnDK/qKm0bYMW
w7HB9aLHFMFDkpsK2cZk/WuVMWwzqXCEblux1Z8P4a/P4s5WijlmIhT11ofXmEmjL+5gmapcgj99
ljJ3WbJzoG8/KGR6KLrmiuYt6Lo7Z6lLVZizWy+A+5e1mpMP81EaYIkO/7WQyBg5PPfTp/njcgje
Q9AXzeZ00a+e3zKObHBDHxOZJjGPZxb2Pq7/NHEc22nvAb2a5EJXyyChVrU8aITnNmBp9CyW1JG6
0ZA2EaguqfCBlGt/boVKrBuhIJKogghp6+GxB7DRiev40EgFbgLrrCFV8V/gzazmV8ZwzNeTyI28
fJyPl52Jb9lD+S1Xiu3Oxc4i4b/qvPL7EPZD1yEoJ7jpxL4ZY8ddVmTvJFrNRxagngGtxInlQ0Cu
Bj7lcgxmIIZtFKcB8TzCubs3UvGmH+6TXQ9TTrrG+It9NKleAkXOnhyqe77LSL7dBlWxc768jWEg
xOnGeqlFzJtOAQVPAGDwWyWZhFiWZg7w03KgUPuBPQqBP5/nhnsriLdEfEIaEctSKcEXsE98fKOg
FY749Ev4rOz9ZIvUl/c8sWtqycny1+P9sbEnQzkYY6IBzw7oJrniGxcPcsstAXI0AN4GOcMCwK2P
bYeulOl7AUrtXQ9Zq7D/15ue87354RfRD38PqSqIYUApVuYn3MX+/KC82LX3cmQ7E+kemAKIWBE5
RxOOx2aOpdQ52lvO4uuE79JFPyQlmFweaiS9KgfXsCYunrsh+GAw2wbki2hfdjAqvj70tn3xO3vz
u75hh/eMkdXgy0pVx2unyCLqs9kMWDpyfX7XLZJu3eNfsUKKdXfD7uHPrsDBd8M1RGZHRjHFW/rs
whzTNRa+xpU1pp1th061jqvSzcOKSiIdRtpLtoXbzCblu6h6riFMuSry7/YlJ/5+ZIQxbWNG+PlT
5YhXadZ+gLOK+G5IhvGiBD+WPqkdKgVtBxmYhsxO9G1hvUIKCF8fRpqa3wB9r9MQTlvPexLaCm7f
GmHGtLqNXOeiBW/zUmEsZSblMMTCwsz4P7g5B6OFfiwCK2yxw0+MAgbQbFeCGglWVkwt9HqtwcT8
dSm6lpJcMelkDdMsxrbLiHg14hoIi4n5BvYhvFRpz8gF1SB5uLbcr8pHXkZyUhFwjK23eUoLk+71
QEk+r7XULAhvN+nbu4YRcecQzA1jZoGILukwkAESYmfWMTCn56w+p+zGSqWmRliniya6YODqZZH4
ZRrYJ2pfOeCsD5cOgFthgPWpbE1NyfxUomULRhfSFTDYB3KP/+PUe9RBQM23iMChvI0yObxlWBZz
ZiNur+Kng6nA9OsRbxT4t9G2JC3LvIpbqA0L6tMcb5mkVMid271dNQvmjXPTu3b2lu/YVN6EDSRR
aySsqiYPUBYU/fwOMnX7aEqpfjMtY+VGF6De/qThNzZpRF2Qa5q6SMCuuiod6fLHWaMQpFoNiO+x
a6jA2pmrLI3daDr19PGj3UZYsRK8U+r0mMTkm5CkYyi4o45F8Fv0EQe+bxiEAffI8Ih+tfQ0QHf+
n3bGrW+kaVX+27kEwC+CeXXp2ThEXISBzbiQLBc8u7q5hvUaIWSyiJ6LyBH++FP4F+0CreI15Sre
Z5nMfi3Tf0uoU26cs2647zMiDshtcVVwyv/5wBMyowuL1u6yXiihB/9vSxUy8+mmfPYutbdA3mRh
BbYU+BLUEcayDQV4aK8WOx+VzWYwnS5hJwDJbPt4SUX+/GOii0gfjShD7OWbcQyFomO0DpKlDPEr
IziorAT6Ld7T6rNwqEAqbk3wYEnFceq9hGkr8/sMqRyV/RbBK5CuoWyqt3wKYZaOQ0eESfT/502O
HPyRnYIFIK4+JjnXVEK3mfpi4gQimOk9K5xRhsl0hpnAcJWRBJrT4rcW9HeIhwKN1We04Inc+CG9
AccS9aTnVZQlc/ywjgzBmDZhrIZFLgigqzW0oMqWCsXBi4JWveX+Z/DoEU+5/hu0eGOt+pOZ31WT
Ls1GqveT2r4qBj8L5OHbf/UXPeY2NxMLrUD22xxsvwfppHqNAYK9mIh189bHr2vO1WpZNG4pQlvQ
hZLczF7cNQcSw+x6D4GzUoJlhXJMzw2Lji9d0L8obkcZK7d+gG/nEQ7nAAU6XLc/nDXy5+HLpjM6
Jh0Y5t/97oEnUJ08KhU/FkbY4g6hwgoZgx6gdLT7BgTymphXEFKVfSAJayexTQTElBUCFhCeFmDQ
k3DeGCvN7NHdVqNmt2AI+0Dw6UVAmS5ff20TTXmaBs+ZitouB/96aTCsqSSidTpUBhDXkp92F0Hp
NVKokB4liKkBLJqNg4YK5/U05/Bowxasv76JOFhOGRpYF9e7rX/d3bCl8MjT1EpYwKQm6QJkcSxF
SuBCBqm82fGqUVWkoze+9jxgFealjQB4B9O9evRvaOXJ/cWhoLL+GShEivvfh+IL+bTVtw7kl9yH
tcOIxIv09L6eacAA6Fot5aUU0Qo1KGbIB2VNClRCIwgJRTBgOBk3b4UyGnlRJnJN+c4c/yP7MnaT
ncOkU1s52FHm8P/ZWeW2kKgF7aELf2kn4G2rUtrWwJ4IpfHxNLVniiI5aWnYRHDA0f+b1FO6TuMP
xc4/UYkBK3A7TTrs8xIHpm/U+ypFec1MOe0aCC5pjd6cYfrRtPWvn3oOzVJoDBafH+WDsAniAeeL
q5HFTi9JbUN7lidjecy7zuGUJMSEQLuPdrSw/oa3I9LEqV5Y0sCjjlvvnWU8B5GZxf0kHT5XeGy0
+HQJ14+YxTqz2/IMaaRC9/O521LjzXqhuTNKHFAiz/ViT6KmdmR27ynzDBRQtTdRNCwzRDqkH6Bd
no+vpYPHj3OQS0CN7PnV3uqO5rREfnKRTywi5Af9se+OYdQXM7VckOQd0LP9BBuRBoVAPt9V5o65
5r8F2tTTblcozm72hA/i0QmKGeLhxpwriBasqAnsszgkio3EhVAG/w1vkAqIEfyCNRGGB0AJMVKU
rNxRLYVQAe4WDd9jqTlJw0fQpg4jycMA/Yt8lHHIn7vTAOnm2i/3Wrs+D3xGJxKb41KIRvMwkaLt
ZnR9OTWVltpn2YSuqTFOa4myx5xAUReRq79sAO21dccV8twEgYSUYgzV4E5MCXdR67hfSGaMGBzl
MPNTrAqmBkhHM5qCexsGqpgHQ8WqIa6FzEpqh4IBwaVuvBZpmoSHYR5mrtwDeKEPg/FuLm/9JSdJ
Tb7n9ef5VG9iZSTF5SrkUyjsjyCq+io/ZI5Nhb9UvZgYtOlWD1qf7DjX/rYtWdhAgAS7D8TekYsv
BliK4TC/+ewMJe+q8IUQybG4otFEgpUZuRTSvehv/1iFzfcwv9NQYkVaDjDdtJbqMckynKzyq4Ru
p7PcoKB2PEvc4SNoruxbKUu6mbXsZLRMOSBuGi/13PqRK2tON2uQGuu3zBRtdvWSm7beE3j85Fxy
3Nc9rX/26KzQDuipsTAOw0wC362Tk6khFvHHEJjatAy24XvDjKcQBv5AYBV1Y7Iayu9YNNz38KIg
l9RUWGIQz4CV7rPxsHgaplobH167n0L0vfFk4hZEIoZVlzdb6+qQXUVDfQHijLseVdbvAdxoMMm1
WbvYLyWS9vwC/b18x/SdjACeXbJNUM3ZM9QBV5qlhKYUOSowosaJSvBfpSHquzO69OOd9RA+OKNE
9oUWaMj/0EtT9WboD0Tkm2CGpugX4cZAe4OiCstoj0M+dlI6DZ5lPC6Nmm2GFKcBE2ngIUBg4Swq
SYKIiUx6YPDh6+2C7pGj7DOBU4JIrX4VVhZA1BTuR0kiXUbkWSnVcqZGjs0ME8NlMtibtClZdioL
dKxwfV5PVKICi2PrI9BL9pm+4ruDAveRStNz0uRBVDLFwGqvvPpmDGf3/atZAtpw5pjSTD7+RhqX
w01ytBiI9r0voJxr422UYxmmsCt7Y3EoSvAXaZMy969AtwaWjnk+q+uy5ut/y66SB/+Hj3IOLQG/
9h5NzQ+PWyEFSLGxoLXBrrqkzyD+Xx67GURI+MC995POH8KwQ/B7DfV0ztnscRByAHipAQ7g+hO/
C0HeiVG7Rw0ES+bLPgkGdJG1tP4qOD0CB0EHognOFfxXD95NixGO8Fm7Wvz5xe+HQ4ZX7nScAK8k
oHi3ZKr6QkGg1e6zUQ0IWiZTS4gXi3KFd1t4s2QdAnnIfW15mtxrGOR3QoK8D4Syx6htoqZLJl31
1XiE8xeFGWPMBL5oHMGHqNKS6Cjij1Bpk4qziejPk8sexniQy9U3qR8Dkgllj8w9boUZGz77aIH4
tc3S6JVnocKy2rhqXNmFlAVZ2mt+wQAuflwY/7K3Y3uyursyPxT5QzZSTej6lvYgiubVvuh3HuAy
q+9DIiwVoqXlcPkaw2gECfQ+Wf9fVA04HOaJFd2D2/QEDM0tsLHlJdstLwa5GXAdCFFHO38oI2ap
Prrg2BwO1xF3NyZg/3Ja0uOOemeO+hT7IBjU1IqvTLJt0GeLsLIgIInFgU4I24JCqXRJTRWq6c8f
i0mWzuhSiB+ZNZdi8AuR2qYcyJiC08IgCAmBnptA6/NB8fl3f0lteH/DiiPiIseYLWFv4pU8/czN
+rUNY3V4MWxUb3hapvNRWA1e00AX9ijeSOY1NJfmzqQ5D2aAwmdq/MKQ61H5gtRwn/0fVY5cmTMn
2tm7KYezHLwmMQ495qyXO40fw2P66ZkpycFa95bJ9wHhjmXYP/8Bzn9QvXbM1xb5rbmwhm9Tgk8h
TuOJMsve9vTkyWJRpMMRVkDXPP7sLkX1Bo8FP5zkgK7AM5YGDcf3299/4VnFIE6lD7kyA2et/eVQ
UnRrJFw9GRAxBHoEQxga+78QykWT6DE3z3H4FiAma+jxSoU/KNihoAdFDqlvALEFSGMEBxCRj1KH
Y4o57NMYPSU/qLD7y1/7bu7t7xxVqB78mXmeiV3y7M8CgGvD1/ZCMvoj+0ZIWZDmQMLb2aNSUrnJ
932EZybgsQRbHOBKnh+lSAlOAW42jzmbec25p8yhVz/OPqHPLIvmNAiyd+zzVhfAswMn7VlJ1WZ3
cnb3ccdppbV8TnXJiE5JQ5/Zuumqu93+jNvGkMo1OH893zoPx/FraciPwPIGP1s4wCv5jtaDokda
lAfdCcbnaeGD3lDNLA0Y6oG2pxgeZpSxQrMiWCegT/+bDFXA02VFXYlqcy1bf1C6Wje4apl0DRk/
8ziUhbYkYK9polZ7t/oPoCzs1e75UlJbeKUqVdT2LxOWckaX4E3VnDacGs4cF5PXgQniyvr3smfj
DEarJCq1hOkEMPx2Oh997O5juKyKDnCn6AKIo1Gd89O+gYCwxVfic6D1akv+ThtCGAGudQczMHrY
JM9AtpYFxO0YhPxzccWvtZPfcI4KVX1Ln9UdBwBbjJod5qC1Jy559wrpbtxzdKtgKwujpEsDR7BF
nIz5p6l8Ve1QDBFVps8LNyIcAX8hXq/+uM/4x0TtU3e+mWfUtS0ZXXT7sim4BikDBwcCQdcf3ugo
1Q8figAHl7P2tIvppACP/k4kb4D51bUohDMxNeGsc0Ta+HiouPDxnn94V788629KA0yz6W419SOv
E93pKAKaCIK4E9Z/HPilW0I77AhbdHnDBGykgb4e2wLtnXXFs07iiLA86h6C0L5ucRo14gYyPjDM
Y50BKzO70/sht6liYui+tUnv0ssPLl+qxeFGfGnp5YjzKakO/fr+VHlUoaTRIS1uhEuHYgxjJOoO
G17N/A9p+uIjSl7Nz+nxIBF08w5AdO++CgtDg1HHlYOGRX0aeMB722sijXrW+9MmWOEB+lrEpF75
q2Outl7scsfTky7AlMynOWwVuVVkRfEV4wQMS1HxA+ppsJtDxjX1ldpx3l/lHgvBNoEmUSmU48Vk
yd5WCfy8FwRccItLBzkDKvgi7BbwFcbmUnw/xA7NMwUWr7jqiqbXKqlhJSrMmX11MTmeKvamBFLX
TUE+TbFBQuSvsjITkwTuijsA2Kzdbju/81TFYkY1R7pGpsD4OjhcfjtQcDmaSPU/FP27zOJBJsDg
tzD+QSHp/b2HUHKMsR3UVMVlJq3mpcT/wbHKQFT26KP7TPcxQVbZRo+kqLexSvp4gnf3gIMn21aN
vLoNQgFHoiZwIkvKV35SLCnQBz51J3SsTBBH6JkLHgoSwkPJ1uWXtQVPzHC9NnGn6QuwvDcp2K+B
5RChROdr/Tn/QOGrrF4VTIHfx4Kf8Dcrtskcqz0988Osjno/5pMpJVd+5tNpHuFsSDGt1vKaxuja
MU1MfVxP5Bf775n6x+ADLygoHZC1Wi3Q+v60yWd9FNmMAp/Dvzxic0NWpxoC30EhzZHwxuEMbEj2
FMBRbmtsggO3+iTrK7jahJ/ax/drV5BJZvp4GJYoEoUWEUbLNiNOe1j8i1vGKGku4uL2KHwRWITg
5/rfTDd+hABSVGnKxBtF4aSkipYgOGSH+3n2HRoUNg3ws8AcsC9svbHb0r7rl3wL3Fd1BC7TpcsS
MIzzI7McBAnVVpADXmcAybTE4DZfWeij47qBQtQTjJo8VxUG18OXHJzxs/MvulaMpko8v9rYWROq
eJDdorwcxQ4p22w83rrYON9SYx64erSNuqrXSBTKC9oMPl+6GqiItjpZcR5etZ+nBVCEWkRLVnjp
voobW55chhatOF2mYivgLpz7xvDqV3FnOGdIKRkfVmn3n/LgeAxYOVT2S/M5OnXYE3Y8b/JtHgiY
uLL0ls9M/8HvSOokz/CYp3xJgEA8pIHAqfMOzHUzc6pYos7F5fSLN1R2P0SwjV8bIH7BB6gVWUeW
Q5GC/u+JZbJdOYaKwfno77aWPNj1wUsoeDkrpjcsTpDyFx+LQISM/KPBskxiQ64cSUuULDTqmDSA
oYGgdrsGTOXh8MDVKPq6UupSkyhwotnZiWsfqkSgw4vbbazK5+79HRNThwQKRsWKpOAXvc5iOTZO
l1n0G5bGTm4V97iED8nyiM213hbq/wl1E8DdwBHJsVTw8tHy+8jWjv0Px/Y8aZAGO2lNFLVJjKgA
uz5vXnmJwi4+bXvS7Q6y7Cs5PCddLuPLbp3uaGmoErOC/+OPwNqF6t0r6NYmpy//dzqH3pDr/rVk
0/nJpgSeRJZKldIequejoMDhVh8sY+tmsoxIoftTzERsDfCWuEh7M74vA4d3aO+aVFaye0yqHSeY
pi+n2zGtZLomAV46PSbObi67T/SAuhmYJNMOHjkY0JDbrEMXf5LRbv2nKMUit5m54fFHAI58M7QV
XBONvGuoa8YZ4pYRbKRjH2S+jAbxnn7eIHvQ+hXHRU39Yt4DiWFTwlPf0yqYwH1nU7RavirQHNBX
XXGyjJCWJHuvkSWEGcAPWP2dUOX1CVsByGB7K7Bk+ffO2GWJaiHJw6JJloVr4lYwOKHoP8om/Bbo
Q1rRgGE5sPLh3nYdt9bReIEHOGrruR5GFsMU7pI2vVhfJqLubH9qRNyYeaf5Ta5kMcrqdSuHSpXj
D8buoIFAYH+s4MpiEw/U168EDVpJcuvfB69a2fF1TGFT6qgkhvwHqAS3IFgbwraOrmKLLTURBRTJ
tbBibaOE0pwnhxjdKFs3UMMUuPWJ0HcTwC45v+kte0N2bLsdVr8KaEV09VLplSl8294q7rlkjOdb
Z1/aEZlu2KlB1HLtlKGu3oo/s9BkRLkGvEdiAcUc1u9Xi5V2ycNiIeF0IVDNnmCbN9OfbjikiA0p
3QTjhqaEFmDlHEPYDQiNgZ4rNQ+3dSAvWVeYc5z4/Z6YTX9QBo7jqRQXbCSRDbOU+00vy1ljObBa
5KiBwwv+IBZHFmfHA19Td3jiunOCl2yzpREQu7eiXfnYTUyWw8vsXXzFRbnsb7DOAtXaWu7TJyIc
C/bkGnh2QLeIAOyNdo8aKZiv0+HfrwbywTTF3j6fv1iiYSayFCo6jwCwffEEYeZooxLadqKV3WWG
yzdNMfkyA7ktuFOHoRRC3PUkqp2UJLLmewx6RyBv9/uKTBsiyrMjr/6RBMAsgvHCIDJcW3o1VJso
4vAeH1J+/i98uOtrSb6qdoWN62bCXpZ+FxjbycCK0a/Wjcjh3ar7uWxwMLNF6hLlbBPvkxQyOkey
R67zFZ3gGxTS+6nLzWg9JQypXWlYmSkrNQ1ZftuM+FukjopRg79Kaa1crwnxYhNYMB5baX4fPEQb
w0ourZfNx4TIsGMs7UPl87izYk5WR1UfWj/YxkRth2lDji7wwl/1zNUUWD9A/50G8ufEz4QX2Ysc
DKomcmmzNgznCzkNG/AidKC/3gjhb2WJCsAyEa5PDou0t11z53gcEgBhV4bw6k0ZhrtRQ1o7KBFF
IrUS6+nbWBKz4m+yAMOzS6X33LJRUABmfTiGhKLtaZgd9t10Oz+uP8fvgQBmyb2fbeRNdqC/CNWk
YW/BFWr3cPUNHCCpKuZWpSgldK4viwQUf5AgeolP+Nrb3tOhpwrt7sPU0sy3ob/YVX5GAbSaVhPa
ZmaBYrCWVrjCjMUf7BKbxLdEmGziSyg+FcN5v/3xoYRBiKWzdu/uQaQXfMyGOf0btUbpVQxIAAKF
1GkGRHgYMIQLqNTK+ufqXxjv7myLnZ08KVZf+YChGfneuV3rBtz18g9pnTVtd0l6bZgv52+Y2ppd
S7Z0IQtnN52+fbuDqnkOYw7pPNDKX8KLwswbIq5h3fDxIGHmVYARkTln5lYxKu0snMMC7pTip0ky
nk1D93yy4GYeGUiX3+gGufenD0S/P0l6zHVmUU4aMXKZVofp2jz/Z6esfggaBy04wsAcQIY04s8J
osV4k5ZI4Wh5F0IGDJC9MZRB2MHGQ7OlwrEFCiDoxq2fA8LujCLrlbviaTWT47bikSZFQUyFlW0i
KrQJa7aMmBW9/jgSfrFCC8tWSWpws4J00HtmaXl9W4kl51INBaqvcVkMGhPSWff1nLob8Sumc/Uv
01VG8wbmklAzZV0arVqGrnqGuALKKGtRy440m+OlXVjFOjKwUa1Atp8rb5EBq5vWfjySwDZ8wSWg
a+qGAOQGaEo+ezImmtMIkMciCEYeQE3q3egFbFPGnTx9rLiTxOFjjvrj/cmC91RsqgNr0z87GgiJ
58NWviiOspr31lz4+4OUDhhyKdXVfO/rhhiij5DzNMhWRqVDclbocftszpirbXEWCD7ORxaqS53m
9popG8ClIk86/BQPZErEf4UOtIMUz/yx2qfxUyD2gWsawj+qm3lHANUEV8gdmfJ4OMGUso050Xeq
GdY82bTmf77DJJhZT02YnQ36nipMpgCZiQNqj4cDOfB+uVPH3sZME9LMyBXsP6RJpcSK09BvGF8n
KeugvfOsyizCuxprgXksUJiSeC5weDNUlLnBvaz4eo9evyvahJgh5yNscmlR0TKYcHYtc3fNhVKW
75kWs27rfjkPl7ODEFol6+SzvNzYNZ8gcJ1hbQiNxqVdFYHiiBuWP2sU+cZHFofB6QwyH4nOc6SK
maSC2Q8l9/dwe4lpJGIwGxz/52QD4Sb1xiZ4oY0xH3xXRXgLI6SdNgGWm+MWWaqvgi4flDTgs8bP
JyJn4a2Nx7QYjnnH1UexksIWVwYVOcYambG6rXFfr/grpBV89qiy1XBQ1iydnhsz3srsq0XiPkjz
wbwijp1nq9F7yFpdbtjouL/xJRKOf2tpK4WEo8yv8/6IDg0f+aY3ATYDsrfscxrcRj/ZRphiHMBR
sUFtqNtUawo65uLE2bPAuArT9ZR1VnOeQCRunlmeObxZNNSJB3Rjj/A+Uq2KolLw05TIWNs46Ldm
M7tBPZldoeoHnzyYtp2ZgO/LvtrqvBNhUE3B3Ia1hpLoVA1H0yLwrNtfkXjUuVjuC9oNzYm66XDb
VNmELCtUwqfHXycuhM0E2Dsvv6II8fSOlknm0dcTzzkOwfZFKhWq2Vh3Ru8oOVnp8DLZVQatNbfP
Tvm7gm0FOXMoAzXUQ2tx3mrbTxX2c3EGIhEO+l+HEUyidkKvHXmzlql+LF6/1A/fO49N3a4ceunr
LLBhnFX15O31SfEAYSoxJNVYhLxgOVJcNY7+sWpurREc6NFzU2ELJ2Qex26Wbd6613/4fLHldLkt
mDJd1e9TyCda7c5BDqqh4pZgUNpnyVLrdA6h/h33Lq4bdXBLPWaoXn9ghbEOwkBo0OkU5IRAIdQE
CftkiEn5lN5Rpc/0gHLzB+SBHhYh18jkI9kc8djPvWkqeQ/j+DHRY2p7s7yBVGPImnuo9/W1PWjc
omlZKU9Xcg1mz1I6i7uJy/Tt5C7/f9/FLXBKIiTQHePK88+kOF/xt/xKqi3SM5iMGGTBHuOUAEP+
BmEPgsRUaucPZ/FfjdSpGP2YdI07x3LnRXDPrgHWfSTN0B4dqAuFU0xsFWsZnVIa3riW1Ml+2CkP
2bBBDHh3bGS3OgAQlAU5x5iKGKIIDTAWN632Wm3NWSol+ve9rxdJYpXeZUWFM9emqxc/dIMcgupD
rEyh3bNgkeTlmEvEeQH9f0g8KPtzNHkxSlKOVme1iEEa5d7TRL+Tz5ZtZRGo4urt4roeghrcOm6N
KgaqfpFK6pKQLqn0QFPgedPiyVZB8FN1fthZYPwKj5VwIrpyILnu+0QuAXwvXShA9K+R8XLfppxq
6ySTThSGBGhK+AodUxI03MLEx0HrOeJVf6n07S5eRZa3J/tgdE77wfmeJSaR76pR/BPI/cE1K99s
Y24lTDf5EmxP4nAhN4kcnuRBaxjNHxkL4r5OmW6W9I9mOESzwbSw8Ln1aMD2GyoamsXDxCLQh1X0
pa+Uytuo5pvIpWIFPCpq9bfjlnkb/sTnUfsBdX/IAct2OaYrpAlkn/XzMoL5YeANVXZkiZrF36tD
ZQRO+oYEHpCcVDyNqIH5yCMIIdqxW1uFcfRbw0LALUMgzeEEn3cTjVcOYndaOjuF11pv5tjRK7Xc
+YoaXadUfbIScRT/Hy7CbxnsAFQkrmy4bd/PDSh8iW5kYx5h3+pDGdxx2a1jltYJDefYLYgxed3c
uwkncDsUHfAiAIpgrR0RQfM0KxjUMKY+UgkxDZfnlQyUiyMV/DtUWXiG9ZcwXBaXmmxgMtnxzH6r
TzQtzQrikbjVKnpAos/tK8aOncPRhLJUnAR/9UDhXA65/AeFku4LlaClSIXCc8DRbwUPIkAp2qcz
SXnD5o8ZRSfY6DXUMwmWYMJm3O/Zw0mGG+eOqh7Kx+dKQ1t1yuttcDd36GwPdJ6/jRV4OXot+bwR
p2OC6mBIuFHkRAUWGN/7/FpSeIgpCCoClvURS+UpW0uKxvWKtCF6nAVs7pUBmbd/Z1N5EUWFuBQy
Fa3sfUA+Fk1BcfK+Hml8mNgPFbz/F+f8HKnmJP2I6Yjqe3/LLxFQJ+0C9YItP8mFCz0otprKYe1d
ufULghUM14L7pi17g4WVPT+qttOQspQLaDXbubWe6T2oVcRFYy3c/gZ1Z6FL/YWBmmAJ1+Qodnv4
lAgtJRzQScDpdKKGR0Pf1rDKU0jwPbCCW7QV/L708RInZppQZbV3XtX25qYYb4NVzs5+oa+OkfmP
prlTWT46wEIWH02DN2fsA4nh4kSzd1r4pjozsMFz90XhiZx8QwrsA3rMuS/1GGuj6F+NSEuO73XA
j7lx2pZmXkjpMyonl6Fl0gsbif6BFqtYZqOZNfteNI4XkWdadbfvjz3szbwvdtEeax5SgfelJXGi
1B8jhpJLn+seHbAaK/K33bJUIQevrDucsbcE5+mBugeByy9VjTwWmZltT4T0miPSyhhtcsUlPp8o
K6H0ZbE1G7v2llsifRjGAsmmf5BpjgKFJdiXOrirwI2L/EN76GLwymftahwZ3RRWcj+jQFeMezse
t3BcIK0mRcqsuEIlTqSZtjH86v9NXcNdcjC6qVeG+m4Cvck37LfwdZ1a7X7xwL9XyaIaLEYhEHIu
J7JlOGTesR+X63LFfMZA3JNJXBOzbYoxJIHSQxGMQEicEUEUzZmL75RbcCCFJ+Xf3mGwARrzENK7
/mHXHgALHp6ojyBv9KmbgJoP9oDYJMS8SIBmHuxU+YUljMFPSnGHeENfBucAssphGt6jrLmNKGaA
k0VoNuzhZ5FFtk8srBRcYATrd/wh92KDj2zbo7251KHJKjqKX01FpTrVrBRpKAVJH3/gM+JSVI3q
LpyIJXdLNtjsC5H+z+mKpex6ZMGbW9S82/tyTA9N85lZiFUHpUVZn5/PGxr9aaaUNASJobHbmhMD
0R9JxgIZlANP5BUEkq5pg5okTPR+RRFeMAIWqqPewKoo19y5Nx6cgv0T2APTWcO893r038fQe9lx
HZehmD6PiMqgLJ8av9RlOCtMQfDt5Fl3D/d02JNztIMcf4JD54US5zxKDRN46gLnTn+06bVMx35J
eXPLiqLLSBnd7web+ZbKN5t22wtZ5mt56ak8LWUN9h9zp8l89Z0vUcLI4b945/gU7BroKJGiMLL7
pypcFbGEc0g/5rPAD9aHaWAGRT7iZNJvSCwYFnkPdJ/WZEI9/5zsKGWFSU1GzUM3W/QHXlNgxq+O
AM+LPSBp26dbNlGYM87fv2uPULL1gp05+2kn73Z/maR86OwaXSp5FUOcnlW8xrJmcW8/33Gpvi3m
SJftLdt7o0edQn8dTQskk8gnPqcMl433FS4t3G0KuDZ1X1GK4vPqwWVEUM6dLAInDOVWdiAfnJw0
Ti+CQfI/7tVIc+x5MIi8CKhZNz81Uaq4AiivCk2asVUDLe8jJe9QG7XWbETs+81Qz8vvhBbDkd69
GUCCzWbdAXT3AdwG1FBPhAJpl1qK5F/Ia5tEeA1k4t39ZfWIwLDSTgcw/FCDw7Yv3QDp/c6k9zFh
nHiTVtmBo3V8ueQFdIap+RnkCJfQpqX3I+pQPy8ocoYD89i23hDEnsz9axfLAj+fPZ9C+lzyrqie
k2oHuzPvdfDQo8f3rgwr4mjzC47pCjaLS7MsxX/qD93p+FIQA87FYUfKvqtYP5ky8VFh5uqhmo5Y
3n/F/SufoY6Yf2cUmm9UNCSO+CiiTsmc1NNkMoVnA7+mVHmkyRZMAUUjZIf8U4DW0QKwVR2ZccG/
DG5DhYZyDSShHNO7BkuWcG1saD2kJQWcCHMmXwNXH+hSX/1eeoDj6ah+9Td/6Cn+fYEQ80KjL14Q
9Cbx+RJoK5E3/4BT70me8ZVNqLEOguqfHazDPrIYB4Hf/t63Iw5Ug4PMwEvchiuM49LZGFKJsTmx
U85clQ8O/yZ8LllBBisValaSxlQ3rTbJsLnilcylJDzhjpO1w+Vv1xQbhGHx/X239iaE4Zg6gm+O
wiwYdjlQp6O7RLVs7/4xyLv/qItcZ4Ui57ZRbnQ1lEcZCU1GXXp35ELV0QjcWE990/LsX1w5+pVE
QDvyoe8eeh2d/fk3yIeJVUo5JOWutLjvSuCuO/4ZKVfDY928vcmyNqw+t//U2cVzbBMU4d5jfucQ
34/5Kcp3emiXhVAg8XhuZxxrKUZh6ZHEXI9SzBOXymthYZfyEhh9H9TByK6WZvQEp3cFSsm6zd1a
ivbQKs9xwPQXDaVo6FmCFJFR4D2JPRt8ov0lkIrFQuQaeQzkrIRR7KWt0x75BjMKrI3weZRTi7M3
s5URYZAx8YJVqpbRzvDxXCs44xrDb8/cEfYj4+vI6iSPmfIX57z1I8VGw7SAeOGWgfOotXEhZANz
Sz3UOQcT68RWiZP5w/aJpvReKjB0O0jcyd17oTVdzNgEVgG7T3aE+7XbHr9wpEjL1cOp6oIQuOgR
vfnjAT9xA0H9KcWEjZt3gjYYrZh1bDIBprR1+YbRR/URW7EEJmysrsVHv9vZCoWewXLw0wegtDOk
359SSEbtGBD2YbAWBN12HAB7saO7uQiCH4V0LvobfQ4UIpuYwMVCw873joEqJgxOYjUFq55GYgJX
ShdaucB02Vj3IBI+W9Aal1PeiK87xOwG+ou16pG7vACmh4HX9MTk9+c9V4hGW2+MAOpuB31rSiyp
iY6TUZt/yRsH1aTsjHfkP1Sj+FxPRcc4TXfFMukEKq8z87I1dIdtM4Zg9X+R6gV61/lwa7IRStog
0aUFOsXLDLLy9nkZ1mLlfag1JWKr48vejDyWpbBsaE4AHmf0AIXpaQ7UAkitv2JzvB67/6oO5WEU
DhCc//iiqVQtMC258YNqueURh7hnY4eOLra+6mhzrw8Qz9X04fhGzQG+oUddHBeDxPTKFUgF+B0n
3/GfdaiW78redLiB2+r6yWgnKsDGhgQ9RX779xIDywOwCmrmyGcnotMBXsR5tESKuoz9nKWuci0B
wn/DtRq4oas9cKBhQy1//WCTrdmNX7LtM8ZxEyM50Cpjcwvj9DEtBSsBb7f7yR40xR8EMXmDMVkT
kU8AqdSrFBROGM/8s4iirw/IkXZ1zNOYj01U+7tCPC6p+eenQ4mRnBkkmwMvFlixy2XBnu2NmFR4
zIczAND8M5ZyqIeZ+l52g66kGr0E6XfjpQpkIrryW8qPYH4dHXTiM8DbvQEGH9wjg48NwmRafmby
dY7pH0mdjc1BpkG5vp2SIMUbWaiHksYEEqZbd0PQbXcSwyK1QOzwONsXGhLL7sPJ9gdN/tCKBH38
5RQFeaZNF4oCbap5Mlrj/wWh3KPvZuY5R8pRe6Em5Y2Xb7ekpQh9QIdzOvc3SDTccIUaavff7yZi
Xkzye3KQYRKdOb9ndbgXvUeApEx5K7e+wspSyPzT/Ft7eJNyM0oY0H1UKBs48abvFM2yoLmgmp/3
RAVqpZ3Mz4u7lu4gjvTPIw5b9cWJbq1DJGP0ZJl4yCcEPanRIbYxZYKpX5HSGCLwRgnRR/FIuAGA
Mj8q6mbxH8zr6/xXmczcyRs7PQxb6dluJv/MCDMUlweArD460zlz3Hk5L18O1X78CZwNjKIchVqc
reOzZarC1ge1LLFG+CEae+NI9qp2F+THuN2mYyBAmihtI/EW1MhNt7J4+rPMvgSsFGY0eeUkvyBc
a8qW97KaUGuYNCPjSVIACLZ46a6JJgkSJ+goI7DTUpeUKOZX+t2bcZzUa6qKPKcOUZmwlToANnga
+gAI0hsj4dEHZAeoyXzpNkgKZkaJv4I3n8hmksa3l/7a+kRHJTdpjRPUaEajUqhgnh57K9WUcBTx
aKf3vq+Qm/snMKobGbMKYkStQzjTToi3T+N4uRSGazsMTHRADANsmN0aTa5HRhi5BB2tqqWG8Il2
SQqxZtyXw3SXN/LreBhtP1cJrULfx/CBo+27f6ysP8SOULNAxgWb55Vee0WboU/sIGcqre1I4Bol
OmnKMIzy8rb8vCV+yQ5DY6xmlrgII5HYmoZsRkWnkXUH+dHfGCA/9Gay9OCNML+rhBCda+efRZg9
Wd5L2EglhUIrX0vKh+2vfKFITIGrYdPtIfy1uY+HLx+Q8UTCKK8xzf7qIOdzCDoAedEIVvWJ1VfB
ue74Kcor9QkMdfLwlsmeNAYw6E+03zb05pwA6ivFXg74u3xu9gxhzU2oDF5G3gjbbzutCKZZNzq/
kOFrcvC/2DR7KihTKLzkAFbLscdtSHMmDbUCgHrWfSA9z72g87Lvdtwt5z6ev8k07dRx6ZjG1UOQ
E5W8+93homQE6X6w1HUXmPzHsNfRZdk7GhVTedtOiwLBxg4geU9BpJtPlfHqawIzKnJxHBQAnlDa
u88g2WQTEhqRWjqU2QMWOx+vav5fPD6/9S2dhGbebLPgF2I7x0b6vqSyeKcRfOPtPz7gMhqFzyCM
iWfmu6m59B+RP25YNNMqdU1s3oxmhp6MnWIsVSgv98FehOabVSm1Fgp7DHcYH3Bw7RVPso1mB/jQ
aXVM+m0jejXFGKde+k79/pmFLq16aWZ/c2DQCcQKx5eB9mw9nhm3ClZvcIKoxWyJBwfTO8qqpRct
nsoKgzN2k5gSk0/pihzyOV2Qa+pL6omMtHUmNUFVOmTfdkZ8llF4/JrUWTfw6N36J1EOGQ89Gq77
hf3mC0a+O+l2YEWBW6pexB8UmBSSGMqMJbG1+JlbYQz55X9ndFrmmPLLpCoIUQYJdyX+4E3YS8iB
YLPW+NHwO00bff6JbdAyh85PDzVvktlJgyJ/+y5HD+4g1mfdygo/byjQ4atpJaYeZsBWxXzT0nB5
++OpcIv7TU2nmqX6WZdYCSv9ZJ6X0ENQEIljFWexUwW3kN82eO57WBI0W8ne8w74wETBR/jakVCO
rdde7EzaXRAujq2+iOPRI3MXNcj5jgbJI8FtlkuATjVaEtGAY+wPIvNH7Lzk5jAVzcpLK2873/ej
B4j4IEPQ8kc12eSnjDijCUdlND0Qr4fJ0l+Sttk4thwCg5PuWkTHHthYYHyrYp+lG9UGcHgNjE2M
Pr10bisK2YrZpy6+5CU0Z5NPr77DTOgtHM358LbooWbvpiztrETPoSMlgZ+8AgUCLepkfatMlrJ+
VkhDmF9F3wwZC7TjZuZ4mIpEZo6MELH8R8zPioVzV7hk1+8XckMxM9Mbu8/glfmnsHXD336uIMpR
yvRGSWn6G/TTZQFrPQoGCqBiHGtVlPl0hvo+29vudQEfrFf3sUvFBumPxdNKlGGz6/v3o/EipfQt
ENWBFiQXe2w5ejYOl6vrtRr4d6dvw7SZGVj43EpVievkweNFcWM8XfVa8LzmS4VGyEqIbEysrWMB
eBhwV5qHNN++eKWTlQ1Y7cC1rQBl6vNt6TNkVW4PWnqysyhATteYq9aO+neGYOJQ6PCH2JL6vaF+
5QXJFHVpKAjTijXC7RoDZWSj038QV0Y5qAfww7yWs8F+PHeR9KkttC2ZsblU4s6Ys/USnDWCl86V
6AEQCD6ivscMrETKU2a5hvf1XCgt02SHHY8MWF8BqVXPXuYaXiKrYsxLZLO1TzyaZjKinrXEPYIi
iLYYQCRvvnghAeRncD7Ug4ouO9h5k82KmcZaQUPs16PVGhCIiG8yBp8z8snMQdvxggJNg/KVp3D2
CCbuslB/m1rl2T66IUdI27ipA8y+hBAWAwKngcIB828QYBfyE2MfP8dkz2G1UrgWzLF8IGCzAHf+
jNoRBMzcFNRLqhgjqNaRTicQh/wPrTjSRWtnFezOtmmsiZlX1iGqtF3XIP21uvYplMFkT3GIWDuM
gSl+pLmoId45GkjMR2cnn27zgIX8mVU/6AwTO6nj1g7byQI+Br2sfshQZEZdjCTuMtG3YXk3ch0k
V1QpbK+qG1/K48z9ezlKuNR7sGcewherM5WuQJBs1o3lSy05FUVAVJBzk6g7x4qhNZVes2jF4UtH
8EHnyHAQc/nB/WBzOaYXKceyu1+hhbo3D96sXVeKJUKNmq4HdMYo3D6qCFXBsOTRyW3sAwj9RJ8K
ut/N7SwOVwhE5hDkK8IyfRAOiV/MkL50Tf/TRcRZ1wf/GuE5v2C73QDfVi6Vc1spigTdtE9hjA8F
YECBNIQbYPRnpxF4XKLPKqfsW2J/XLyoHHdcFeQ/s83LqUi83TPyKhRxW/YwyMq4N/9eMQTnso0u
1VwfOF5wrPj/OTg6hl9OXluxzGegByfv5miAtA9oyKUo4Dm7awKP810WZAg2UDbkicuBDw6bPwzz
tC2b3NbwZsuhCobKKKbk4VDXIenj2n9VrS90LCs4fnAZTLSIW8ptONy/fUysHbtpA/X8F5ydOmly
ZebkDDsdYDZZbTUV/RFn8/PnFU6V20sxYA82e0G4T17gl2xgBjksP0fI+CkpRIjJszMqej1kLE6L
CngXXYrnCgC9rPDhv7kDHMafdLR/68GK0HavOnqxXFFBfY/MvIUP1gybp44YaMPlBf63/L5mIpaG
xTGJZeoZr43pQwjIf2o7ionEEeH+MO7tdDfcKukJOUOizC8RhZ0ahmBS4FLMkrK0o1YKdIk+g9Vw
+e//A697g8WLLT/LdaifLHtOwM7ygb/b66nwsCdi+DinC03KCrt7P1G/VW6zTwKXJG5J6fMN3W7+
12Au5qtzWcpbRfMX6LUH9j6ttB3XwwAVHL8n8Lkt5rH4EBOTYUB+ABjbxwhf+KInQya3rtCS7/nz
ADQhuE5t/5Ah0LMDT5vbxOmK3gVme6xIwNLe5EEmFQYRZxzFTMbvuZ/YuEyoDynWYvcCDe+zrc4Q
8EKUPyCWIHS7EjgE0YPDKwqKjLTWQHXwmJWUycSDF7ck6VWNIXeeI3+NY2ORc8SOr5z9u8S3FY5X
c7pEzmMdTgLQXb4jCDyREQ41ewo1cs7M0E82Iv4qm85vBbkOSOd6cofLSuWbzFCQf0FYDaypmK82
ePFwgaafAUbi0QpRFyP9gkWqVb49altRrI7FajuAr6sJsPWjDp8HqK6855nX1IwNBrPu05CYNwLJ
SZUZPobS87qnawFg+H4+cHQOBRBoRjW63dqwHHmTzhravLaZ3SZWKJWX3hVgaD1/qQ0fJt4XY/4J
aocLH1hEnt+Vpu8kZhwpE7YqMlqWA8+mSBNUQdbhSgvB9v992vcPBJB9Ai6vRpW3PvxtGop1rOvr
RPLxgRrEU7W8lUq8OmUkzUQ0Foa/gcV17SkHF81QPQz2qX03C0mvM0A3qierzCozzXWK/80j1y9+
O1EDGswsmLZ3UTSRbIpRk5rS/9knWIvLEYla9YBvF9BDb82ZzvjpBUVOnWe0FGWvvGkUZ+vLffTR
DEuYVB094PXNuPdmvtujudvEaIpZmbUYzEVxc32jwC3ZC/WbuUKEWN77mgtXUNLn0A6R4tl/OSo9
SBluUdcjZk9e8Q3q6IaA91xo5DDQQaF3Rk2h75i9pFeCICOdxe0o4D+3FDWne8FDDQebPM09VGvf
9TnL5x8zXuubPgHnh16vwlUrIxlkbcnBN7rWhHTrV+/NNLFugL/QIa5z+uq/4W7p1eLlk5pQjyXf
/5eT/hU+gZgenSxqD/auGE6ttyTzyjdVY1zojjlEB4etr49MM1WblXD5MDmgTPqK5f1m+WK2PIAc
RhZ2LC89CG+Ddt9epV8ItirrNNEbm34hEbr6K41Sw05jsOaD4e7/i9hDApcW5CPmG6QWVX2QGHiD
pSqVHjtA+fcctfxEwonfpBLheK2Mg2PG8VbFb/ensKx3KhThbZnZXLmzBS0R7tgkJPKWuECzEYh0
SMSnbEsL8l1i9dPTLDDdC26LXFdJ9Jw+ji6Ij9aA2G3qQJ1I81MjTZGoNSKyucFuH1C0K7o9qMjN
90gPL+86o2cw7NiIxDfEI+3tEC9Ezx+gV8QfiHiX6nPMyVWqYxQd9y7mQrHZNGqup8Rk/IPmwIYJ
4N2S95WHuvXKnLbYyiS5WycybM5Ids+quw529r3hccj8bHdDA7mTQbfCaajDPCZoYaoDZu+cAa5y
/Ka8pacP2BeThIOaN1CWg5/mysfV75z9fhmVC3hV5sv2CJu7x2waZCJwsuajrAMOgfOisscceaov
hZX6d4TjeaIxvCw3wtpi8F/03j7CR2fkkSJ1yIp+gKQ1gqUty2kIrAo0IfHl2zgs+ZA147iJ2a9H
tTtnr8K2X9HbbHrgxfgMVsLMZ/UQ+2FBiryBgVGvUzT6Zdf4nw6xO2Cb5KFwgfhJrc4L0RFmYivU
YlQgchYRv1MFRc9XgepRCPmGGBA+a8kunNczucaqDeylj0Ol0Xl9trVJdOsT993NxKWwQ3kIfULZ
OZCWsHt1eIN3CM9gWz1ilFtZ3/4HPcQwe3ELJWk+c+qIieaGzWBWOJ0nyZQO6BuB5fRhqS5FGU3L
tNH54/BOg2UReI6WJpKLzrdekEjzrc8SRpgS3kErtJ75k1AJzfr0595zGKckzrYLSid83rtrchpx
d9umyu/3oa0MykLok//ynNWSm6vAZgRBfAhjcQkPrBCH1ovZnNM9DD8UlLhBXvMIMuiyI6xovzDr
gD3kzWAHmmJILgR0aIzKlQaQtHXCy2qEBYim7DUvtAy0fJppbGEWamcJiYMclcqHI9vCsrHXtBww
abJY9cClqWIz2xx5JnGjf7J9elgusUtX2B5YnyT9CNmJjE8kfx01wW2pxfkpYPIA2yPEsgyNoojv
NA91vkfQ3DpUlHwjRnBrr0yNiPUZ+7LOiHMj5IYy68iBH9PMy17ZI3IZrGhSEibXBR1Dc4aOugFr
lWBgInLkDbfmEneTmpoEWAZmMdPd9RfSriMFNmxNlCWvQMNmM/InUCAyith3LwU93xXAG5gKEtGq
3b94xUomtiXin8hzV6daFMLDMclHEyG4weiclGb/LYB+EHPg+q96ZLpK0L65IVzM9dwChi1Dx9CD
eAEM0CAZUfS+gP2/hjHUPCj6tEWhN9iNPQ3fMwaCecfJ22fd917NoCodbAJ8hZ5Yz7nxL15Nv+1G
iEqgOU3MK73NHHNG/iLDYbxw6zfa+o0J/L6V/4tD0r1YKfME6zJK5KkNwKd2ZI9K+6gW3N2+GJVX
YwHkmPLOwjxH9w4C6baHWh/hddiEUipvObQaGkOie6tfH2eiB8sNsvkFnWGIwTnWCqpVEZLKKsNd
LuQU1WNdaQtD5DvgtNfw2zGZO2hFWqcw7Ev0Za7eXekrMtIH42p4i2bYT9D3y0Sa7hnOWCRnVmOE
KEpa+wmcSzpO0J8wBiWisDsFL4mtIZx0TwwMs5PxShkeDTt/1VQjxxiLBi4OA6i+FtV23BmBBZCq
Fu0Is9BKDrhcaDWAkOnvpdYHQkxr5O4aSGagKQfmdsyvqkE1A1zX4q+GEKZOjC45sLPmkiA33IGS
6iNVoWqBawXh1oUdPRdHj8xizMODACL9Pr0Em4jkQ/81UCbeMlq0Lnj16ZgZ9P6mGWEBowpcxJmH
AAD6NNDJkvY8MM175y+xC1ex4IiUCWzJUTz3Vsn7tbuqC5ruSUZYUxIzVKOWzqyi8ucrCa6VDNBT
Y1xMb2mJweVqFb9/NwL3fwyDsHxuc2pwFNP9xp9bN23B4CmUFTLlWXrbq71L1ckR7OqZvnTl+NOZ
50sFcJoUuHMUad5RekBXhwrqAYUf7/gB+dUauonKVzHrBri7gWqqWbiDori7jhIehBBi9+3/iccK
Re6zHezswGTsECW8Wbgf+rTpFOwW0lJW0FjGpPx+e1HInpImCaNM4vCWbfScBU85Zb9+RxZF5O3/
ggKU+VlCsWLWm9LLtB3awM3UGGN3LiEX5X3vzDDGY2lGlKLED972hyn+oWvDkTXUxKfPXSTdz3mo
tXRamt18fRXoyfFzAreOve2DDrRoORunWtK3Jou7PB/x8pomr+cl9S0T3IHR+aTZtyRfuVCyZl9r
xwZn/QorQfkmHPZpyjTzxhcW+AocwVbVodeZjZDn2EKRAh1UwxzjuEPPlzF0lm1a+793rVqWsUFw
O5c4wGIrN2kl8B/KPrFZuj5Z2V4tY4rR9Le8t/mWqw0w9Y6T94Lk/s31WlActRV1qIbQbV4HybhM
CMaSs9tcVqTYOET5Rizx7/D2Q/7C7CK5Tp/kvTCAtHCjg2KFmeeoGFyGZ0/MVXpymhHf0Gj/PcnB
MDakAo4a2UrK8oHcVut6PdjlzL9FEntqSZC3PNeEvFGwGN2yL86BB/HafZVxIyc+5HysDzE2zTRe
tolDndpge4KvJHXdg6k7D61b1Pt5VIbwdpVbAl6mNYyd5mWsTkzPIZZQxx9xvX5eFEwQJaKI2BHo
EZs1Y3hFt8Sp02kjeYFjnoG9cUpVjwBUnimkUPAiwApuc9Q4HsLmKuwWcz/dQcTM4lgUeTVIbBlJ
spAwxEG7ea+o4EF0JWI5fLHFe4hGF52ZfvXhMkcSlpPPtGfOvE4qXfAshx5nLzlA6d7X3VbOE57J
EcTHyn4T6zr6rYO0wP6lgFsi6UB4Llq1jarQU+G5QAxucoxob4nywcE1ULFKzazckgoExXLJRgmZ
TWFoyC7Gmi037jwnlrD5mInp7/TzEc83B+X/aCRwVplzh6SbIv6zCh2GhEWbzUSmuotEM7X6X4JC
N9fgC0gIEgJYmUlZJLW6rz9yeobBlUjQYdJ6aky+9m+mb75oaAWU3sAsUwUEEvupUGCRTBut7AYE
+nF/FTcgnOQaC+j9B8gHHpub0MEf5BB6z0W7B4zqpOdZDNV6TL1YRt1N9rDA132VTOvbtp6w/iKt
ohdXYN2Y2mxomGygZ1DR0x90Nz1ZNBosJFtkNaL9TIE20Xj2ZRGcOaNhfxsFWHafdPALf/X27zKN
46dE2/MTADBAUhnSyHPaQQlOkIJnbnu5gdu+aw/gjDrCQ4EAF0ZJBCixOhkQr9QS8+gZbxWNVCqH
q91e0YSRsTO9LK+hAZrmUiJjMfiZWCVViZTz5bgF3YxM27TWFpDLkflOn/khDaCpFvFNbmBaWO0w
sv49xIhFzNr48uxAz19n56Hz1xADegEUkH+mgaQR2UVz/CJsY70mhLvyl2FZNt/U2DWozMZzyirQ
AzC4aUmvyMT22b910+bvaogUTRgv2J0FaY6Vp8yd2PU+uaXzvzMk3yKxx2wL6xuE5OtRzMmS/mIP
Ra76DOAS3PWkS7y6RrlBiiTRQf1Yet/d9XPaI4ikzcEoiZLPx8AU5Kbvv2IqdwLq41mFlYbHGrmN
agcp8Cn0M3l+ETxMkB0o77xihho6Bz2l8/zFOWizhqzj1su1iVR6Cab9v5sb6Yv8HedIdDsUYOQG
nyWDgC6gd0704YOE2euazPky3K5K2Zd6eprJBSHa2UVVEVqcOmMQ2tly5jwhg0B0iGcmF/VeaS3d
2uFDOmEXJlFoIOh2r93pM7EyAG8MARJkSHJARPqFtPExzppU1zmATYoZdqYaGGUrSIQf27kQUlJe
hDWFQzD6T2/t9W5TXMbiiGaygHA2ZYvxUgRGvsnnxkE5uX0a4G+w/B2ujyw7ZXhk2xz0MnPTGWmb
mAgLVcgoksj26JL+sbXY7vKmbwyt+Qc6gfohFwBUMkZa0AFQOIkOwnpt1Zxko/klSmg0IaMfhh1e
8blc1MCaCVfFXe1xtAwrswdkZFs3IYX14wNswCLTJ9rvm2BX8KCmzGHeeH0luWnno4HIJT1T+rJV
3DKSFDr1OKXYT6Qvj+mA+rfKYAeJpjvWtuTK5elBORdvx+YJDJGitCy47xCVlA5BzL+Zm0iaAnZy
qKSwQxMAYRfUuWl62raId45Svq3bn+/offlGFvLKxa6ESAB94YFFg/SIWDFY0jxisGoo//biAYr9
1IKrYwmCN6pMToe9iy+/moiL7wGZdAVJGD93JkYcHRjtgvl7EuFzwd8gn9U58hqdvibjAYxv6wrl
vE8n/s59lHPv+LeDz1FREwBrWbSB7SyhHoG3jfUE6l3x6vvZtKyrdNuGGWR6n4IX15wSei5LT+Ec
YUbgm8p4a3ONJ1lkHHmvUnr/qY4mDSzyEuhFcbLjqXrPoOe00AAH44Cnk5YvNRjgIYN3pFB6CvuG
RNdnDjKv8QI7liCCj0V2gk6wtabl1pba/FLBnliTlER+2E58VuOwVCgeLBT9ZprTNbPWF4sV6c19
NOwPYSEO7HNn72sXst2gZv67A9xU6PVf1XhM8fPLWWzNEJi46gyYnoE059CcE6AW3Ni4bYu/HBNm
JZee2zhawBoJsKB2SHbA6fek5JuS1/6rZ1eyvI4ePbAbfxmvbvYJP/mfUoJtBI5oz/wh8UUC64q0
TOBC74aOMbHHq/ybt0WHMVrYHpik6c3oO+2kVu7pIg1Z3CH5wz32RrvYkyb00JCWRHnx7702x0Dt
8azb3M7TEmU8NVpQHNjGp2RYkb21Suss2TDmU7VI8NLST01DF3WZVdzbuSUGDtovfQVx7lVpI3wU
yFNszawR4CCegxzm5XX4NUjChrz1Vvwf4rMY3B1VygQm2VDX67oLu5EBQVNLckMT3PCYtNvpxfi/
UWH3Ok37QIZ6/34zDOU5HPdgqcoKRhq9ZXCjDKAfJr3tpobGG6F7EhDuMPMiqNmw0SEImNtO5Lqa
zjti5dnYz4FZ2lhMJlYFoDxBHNTJZO0mpEGLSPAZ7rO3FoIeDvJ0JOmgm1jjeTa94MmbDGs4xFUw
+P3RcO9Uqtoo5qoH+5cpoJAMTJcBxBPyRge+FlJZP/F7OdWovhPpIvZy+56Lr0EVHHw8+vJzcloo
WYFdvDUyUP1SkNytQQeDtMaInindJEYMG9dGeub78T9N+dfjEkZGI6lX0sb4Uro2FlDG7fiqeXK/
EafA07Ht4VloFGbhwiZnLhQY3n8EHuiCUDYE3omp63IhnzE/zB9XnA9Vi2GbSFvzBEzAFLUl8gZj
JDr0w4atPHyzINwIrwjP5ghGPrIdRuQcK3aZcC22nElBfPhngXgWCeWjgS0JY/lVzvOlotjJU4/3
Q9OIiLEWL8UtdITYXifbryiDNu9Y3+Z3zhDmpZN4XKS537v2uhr18Hpf/nJHWyZ6R78+hIrzF1CQ
Xb1SvqeJW3NoaCZVUI3jDI7iBdytt8AnYotRQryryqQPydiAZbVY72tlp7Um7Rv26N6iW8qoKCKe
1S6AQo+qi+/g1ferRkzCVsFVq5Pq2FXx0EurW+nv/6B74nkLiqVuBy0Ae/Q9pIRfqxD2TT/KURlH
+cqC2f7hFPsv0RUeEreYuxHs0nBOyO/NIWgXEFJWBJOdOG4P/TdlyCyOs4rtRUSdv1VbUKkjw/jh
MXukDuFRiAysOrxXvwocnr4OQrDrcnQqd9x+hILchDo89hKClAdBu4cwHG4sQheQv+8Qil9rl+Bn
tMSxhhOVyBKhVCqFDhSsmjgjyGkwT3S8aYPgBQu6pQ9KvZjVpdE/f9msfp0T0NA7kkYeTN6galfU
Gd9hDtd5ivJ/xeUj4viMYjalY9a1OfdzU5LapXz/bxQ5uvdeZ8DGrRCZ6h/uv2UyNaALe4peasnC
tiVtMSFVij4dpYQWu8M5PynqQjHMPQOr/KqzXrA8qiSuXlpQjoEgTZB8hoUL6wV7dozm4rT9gV5O
V/ZjhjrJEZKv5U+WEyKvu2b123xcdnsxjrrxNor5xO5z5+7Gqk4CT/HIOkP8Rl41HAu2X0nmtGQ7
EkWnkPI6FDku3dpyetJuzmgGMKSzn00cD2LW/N32mGxk9dyEZqeXVBArSkcSKKvQmKYT53GUtkgw
vU1V/6xL46mtlPpEK+QjntYtJzJoHaqRKzqQPSyL1eQIrV10KY+olW3ApMHUybQnNfNjEoI565rB
iSjHWC4sqlpoajzPu86wbWo4IgtmC5YjQSGbeb96gFLu6pC1p3ofkZtFqQwUCsl/CiRoxMsJTxwG
DR4L7Rlg2FBs01dPzOrKSho5FRZBbDgBNmmQkg+dHjilXNdDHmqyUd72PH26VT2/Jzs07aBEwjLC
LjtBys40DVS/XpIPM5cUS3coKK8CgCBP+AyCb4UFNDcHjj3idbBb5UDKY0UmLumSPYu2Ipa6Pb1f
lwAhiPu1UgUenJuVF4oQ9Hcdmdei7x2feiUDlnBum3o5zFBCRY9qE9rJxfJzjRALBqpy+ZzAw8wm
I+8L3aTU81L0zG8YU7bjHArHas/b2TWNAiilDNs7UgLSUPCtTD8QM6JI04HFEowPNpVwehfVjYDO
a1uWKSsUi7zb/jniLTALud+0l4JrEDqG+WKeW+vtHwtinUfJIJok61bFpTQJG62tIQYxiPol7OX9
wIpEFwWamgPIShG8xanjUs3rVFOzB0XVtx/BxN7p3uxl5J36nNeFEAHZXLLO16DN7MXAxbzrQ5Xw
FLLTBge0K2P7fBngGDZzpvSi5sAAzOCdM25I1fhXdWHz0OMPDWa9+7xx4bFe3RwFWrBpzQjzb+G1
qeAbOt/TZlXQWmJCoBD+0vTIXXUWc1rqwc2lb4dnxtYQpRC0CJNxLLAEZSTUqwH7BTbgxIRY6m1M
h4aWQQIb/5XFZGk/gi7rRtCoQZcrMpL8BjZniHpBJ9TfX0M2U/RgKBFA9iWoWIieyV38BPEDuHIq
SS+lgEy15tPDthBTIG9Vu4cjSGAg1czZIuuMmbg5G4xLwogyq0dlyp54Q0FSWEZiGoyD53TlHm28
hoA/tapo0DCMUDVk5cPXP9qa4YGwaF7IQS4bA/LeO5mtZdoBPZXQ8jASr9ewIANALbmbxrtNz8Qh
WunIKgpV5JpvWstu+V9cLvMq1DpuwlwJT8si4yc4JOlzWTBu64qWRjTsrxYbZk2B6hT8RP+i0QbE
ZjDAEx6/Hq2stZPJbLZgTviqxkPOJ1aGsLiuKL+In3pRSpFbJyG1xAn8f5kSYxYo4PmdrsjBq4dN
2h47Y0vqG4+v6YnUhCIcaVIhTWRVn59dnGPwVy1qR99ZSm5ovK90xrMy/VqKo0XlGW4/7+gWL1++
ai1uPnoW1APhE/pE06cIb8r1iW+Gtqa0KKWVNAk0fdgW3HzqYn31yVXnS9MN8WyQuBgHm3Ynbf0i
rA0+Mc8XlvpuKK9CTwu8KvZryDtwtLYYI/Bmj0YnFXgNpPN2/Ht8w6PYkTqutdbQkt7sYnEwUQt5
ueRlxH/r4BjPYrJQw8UelrqHfMDNlbc33N0jWPNatLm9qViz55addkkqBFh9HNzApqL3OtDSQG/A
kdYVQW6TAmjBZ+oiJvJTTZrTecBXf+yXyCFl/nid/4HMg/j6CCB503aRQOwkOQ9e4PS7ulhkcLEY
7sRSTM7JJEheB10/ynFfkvKyo7X6mHLjg8n0b3cOOC3EsWzbKVa/+fLPmLjTMp+MeoY3NzONnjDW
A2ohV+LHqO8DKJ7jBw6nmpR9IcxMwj07E1oIQ6LGpUg9YQ4tLQ/l38rGuT7l0DCXhk2wPLMN21fW
6+JwsQKrxDrw9MWz/q0kfjqADSSfYIgbp9REu4NzchGjSgKl1FkZkFHgMqNyr5yHwPGocXI4a8q3
aRxNZD+26s2FDQ3FM+j89PbWT6NWr1AdB95Vfm+vqTb4K2hzMxFensZ8CS91Orru9fBBVNVfjmPq
iuxTKJNsaq+OhX8zXGQXZZVV+6ghcOBbHC57vvDuNtC+7DUWHXWWtmeT9WNEuXKEWB7dfOkpMVID
IsiF6nrbVOSkaK5qdnO3n6VwPcE05SIgw4CJniKumQQ95J6ORJNPMC0sgmaRnYKK6pS5rZK3tMOA
0/R0/BEFL8Sh9Cz3gqI68TerWxSsKtqXuGNkcwF4BamHFm9XTM4gOC0KM2hyOO4tkaZFf+Oxjg90
j97CQEfscYTcr/P4fDMfKn2LC7r0gyLLf1laxbrTDhSFHWk96QF2yBBhGlA1D2t5kMsBxmQCr26E
MCC+fWevBIENIWUqjwixlVnaQcjmoWjzgsRbd0qx1QAkrSz/5nwwOBkFNK6NWyeqyr+/aWhTRjyV
b0+W+rbyvntsq61+a4XLc67sBdTDdudla/34jPndzmUbaKPwsgqSOfzjpbq9LLk43MKPQIFGcBeB
AhUwnUjHnRSxN+fUgEzImtvazvQw39Dj/w3t7bVEFrszkD8xkxsA1cmm9e8GDfIpKuaEEWeM8SSx
zj01SeacQHECOHy5/NSemfIbkdJ9Qz4hGjwTJRkT4NTEk7QrCpXSLUVMc7/kNSpVReTsExW6QU4d
i9SRRysdKfvdknfwvT9nZlZ04uvt7WUZkkwRzGlmQLHCZ+fr8sjORlXFxHbHlTI3waSxb/F6kma0
R8W5zGWKnxeiImyTKVUQZrjEGkeujXYXIa1epkI7pAVn0E4vwKERoeZS9OGvT8Y4mllxqeBxMVeO
4xG6SnqA0daSAGGCeTcLD4gDvgpYfMlyFJn7juLX/weTtUSXCUG9d7IkdSO/t2hDvGsoSUqKomh4
QDAWlZhuuoJZ8FG00vIzOZcC7AUlMvfiQ/NMdgwgioPxRZJACnmU+AGD/rPUMOYWr/9jZm/NW7TZ
W7fNHD42H1ncqGMIhC9ansAV9ohmgT3iCV9Fmxe5gte6LFqFA3MdkXyJBYVzLey3yJpCCm4hxmZ2
yGcDwyt0SN/ua9PSON0vNFNzUEgjUtMyy3UjZuEAK139+cziTluWQRX+CQHNhp3fhLtTc/6v4kHa
iVnDnYi0xqQ/VWpEFIcqq2rLOrQvzn6QDxgSmrL4uQqDz+rwN7TzMN6pZPaysIoGAV3GqbGcFCHz
+tSfbQ7pE1w/4Lb2kNV/j0V6Z/vuXJ4E32yTsElLXkJj6rJQpY/wpxp+CzjuXzKnZ9sb1VX3JVC9
cxhHJpHJhQC1ZV1TJCXmdDGRzjMAbHt6I8eTWeJVAcZINKwqliPJqwttgXYtExInTVxVyY6zYUya
+5EEIczcj6W/x0qRTCjSPj5PVophy0O8xc9Ww8xoFrgdiiX0iIe8BW7ce10fdFX/y6mQYqR4ZJHv
eLGyrKnl0oNXI6cUYIkQBWZpN9HbVdfijguuDloMa3coMrsFQBzjXvNkia1k/+M6BegbcCdRWteP
EadRFWlQ8jBTwdwbJWOSJRznAGh9fVPeJw2wtb20qjJvH2WIf5thJ4DUt8PA9QGUAGnqJrDgUMMM
+Ihg6O9KV2jI9YublJ42zhNmAz2qHFTMrXlvCUrV60s/lWItv43r4AlHuB4siOupX/uLh8EvZe3R
/3dfrrltiJALVhZJx2z17HXI5X1bWJ3+B3bvuZtoz7ClCR9NO+zAFvhkdzN7p9/5zEhRxeCoiXJn
XrJMFpye9G4U+TAJZ3yPEY2s1AiJ1AKPPCSClh30MEY8KaeTKQXZKGEvOyu/cTOL8Lm4TPy+aTLh
ptPU8UHG2tXhVJmUEcZ9Xg0IVtfW3YaWAl5txqnUfZAY9pvaizDXXNwXTfB4+ZRzu9b+KQRPyknn
Ma+lCGxAOu8wiQh/zPjKe7SuPpjrLz2KlLogu1u/g/0E3XBw8c5ne2/CY00Iub3hj3x2lzqFhAaH
pRl3CptgZya3VpcoccxR4AmJG9NW9OMa5QF7ChmjuO3L/8QnjDGPrjGc5qZS7+/VSBojZxVqdWkC
cEIiXXY/+vkqcZHmpvByZuLIcfpBTLNQeYa04JeD0SolF4Tyrn9mdsH7bSPPv5yF0aEJI19fVdOe
dngnoPHwKhWDEkIOdI/45g27agxrYaHFtvZ8bcx4lXbW3XM420Goifhg7WBJnX9HSzM7VuVBVQkB
+TOkcju0wzEqv5SFrx22iFJ9dYKnfHp4VQWavcpKm0ISCQzw6MBA+bqKhNjL8IsJtFdpOYJ4Hjir
l3awaZlwn6F+E/Amjx3VbjOYajI0toF7m8Ck6ouvXi0OJXUayFMrEFhDMkj7QeEwaMPrSTmTSRBL
MBtZ6NFKoRpPRt5ascPVN4JAF7Z5a5mAQzC97qWh9AycivITNVzSt+P/MfqvwWgazAss/3lK8x/1
csY1GY3ahqs4EcOgsCG7mFXtK8c3NtaU6cYnHfbC/EXKnMqi/8Az9+p1U92mM3xC8v/4iuj9U18L
zBoivcxfqJgjOREx7M5qIC0JQjAxs3sqW95G7tPHzu2RxFItGl07Mq09af+MGrXvOOsSgL3AmXfg
9BNNYXmgLaI7WuRrfCTpMuW7YIEqtlR0O3lVLqKTZrxmFtB9yT1I9yRYqyaOXXZsHZoQNxXNt04t
1rjvQD4wFD44Nozt9o7KAhSWpTA3xtD5R5D1tcfEyNKEitC2Q9r3GzpIMhvisdJC1UL16AFgFLK9
vM8SPLAZ/pzltaUdATdG/RCYn2oob19pwBSmGepOrY1CFAzUmKCqGkplaCi3hAthC7T6hJx0QPaG
fIGSeqixtdnex/WA0qzzPNf9dy7Z6JJPGUpK64nCj0kgtGo3OL0F6ywfkwvEiSndzoc5yDwQUSp7
hpcgjIIe4Du6Gvo57xY/OKfCuwyhzqe7n9Oet37QyZVGYSAGzC5VS6AVwjFjSbdgp9JzYO2ExZxx
j8ncPo8xwVZxTE3NQWl1xivGnOszR6y55tEkOpA5TTA+/+BDa9xdpB7XiHBA5EPKk3ftQ55na9zr
LLN4mGk8FJBnLgH7c0vm1tnXkvm2oR5HoGRTGAq3U8elqcU0k0S+zWbfaPvY3tu2ta+G2eC6UFaP
k8h1jSwooVv7qr6SE9RxmzN42rp+GpXtm/HVgg8VTEDuDr9tLuLXF99QEiHqUsAeoLWLjPgBLD+S
zgrycWYXVQ8uOy5HDt6lvtD8ZVWsjmsSYm54/IkOWs0Y10WCgRusr71mOrU4uixfsANASFk4QgRF
LCLwyLNxKlqou6sk0RRENkIR9yjdRB5lQuuAP6sKd8MjDuASFd95d/3Y0TVUUFuvOZsj4H78R/Ns
OsLbLE/cwZdhNreMhxlMENhmq0iGN6bBwMSBTfcceLV1ptjXtvVqeAeAQWQIbCKmOph1QPQrw37H
0Fgp9uGGy2Hp4wOMFd7XYGgy6r6ty/dg1VLhF8FQKRxdW50vDVni5ZBIcPb4eHJOw2AFk1DYsRqW
ljjmhj4lQAoPvL5LQVmlqaN0nGn8PBQqAbiPCOleBdJb8X6zt6yR0TjqpRYG3GAO6NS5+CPfkL+t
uQXP2GBgWqpss1XxYTj2Xrt1X15wC9pEBSws1rPxoM2CbkiEbaa42bVPEjSmT+kOfuCYadfkXxWY
x/iCxYC/p4Yh2JKlb7pmLHDyiXG+rfsUR3XACSFPCxDnUInqPBwraI+BUtD8HXmJtDKOUbQ/leDv
6jvPy6xjeDBIznxvij+CQ5f/UBDKRJbdYTmK8NnuUQ2CoafsvGwhvDZ9DEV3kbigS6CqUgXL0CkP
YKdqAnZAb9lVtVwhL4l1hzou8gjVqhQ4i7cHeww2dQX8FHGCRKy+780L6ZrvZRvPBgFAmcWe2uuJ
GVV4Z2O6ZbStzeHNNMG/OYG08wQasMzhJYn/I5ireUQOHmfOy5V00wn9jXtKJNK2uVg+THAVx5aZ
5ybmkHsNiv+xqpv+XbtP/f3GpUkqbzv6JETz2WTMzs+UzUziUQe6PAXwqIyFk9TjaIqQuGDciSk2
7lnVh5g6C0FVco4xh7li/zb9r7ejGZykLzV+vQqsnitRCTg3VegZxrdKqGIO7LsCOvAE59qtLTXD
xyZoASz6Y/xJkjm6f3M4neDg8J98zMldyFJhLvfmfkbM3H0Di+LwDp2cvWpV4fk5IFfHVu19YljV
kLC409fVPzIn/6S6aR93VtAHnWQwCtRju7xlOcne1Ykl3wSDJ59Qvv6CAXKJA/9Pc3fnfUWT6tGx
/gI4JPYdJT9kXgpdoKQ4ohAqha4eJazfhmQJWLc6niR69f6oPZ/+C9OEZNYNbtxd4BKgW98vTNrd
WWM1HPf70OXJlp1rkA4mxT8zp27+WSietjW9ezrWpS4t7n6JpOYBWJDthN5CTSWEr5tz3MvGUSLc
8D7PO0Fnacs/6cnLw5Cb5/iDev/6jso2XoVB0Gt5SPuEiAgz5eDVTEGvU9dYxEd3fcoqmCfMPZmt
AtrGQ5Qg8QN1L7t8YXlkkCgGG5HeOT2te+HBVdoMUNGghivrtO9ylMyx9z96haNRyItMdMBcAq7/
NFtkz/IpFjEGednEkLBb6AlcZVjdPUjQdsZQhLZl7Z5mlTS8y4qLHR6zNirb8Jr56feoTSjuTztT
Q7Nsm/f2Nrw97mtz6eH1r+niQaW3xjUsnvQWCH2VNYiPz0MSBkj5ntsjE5rIveejWRjDMMLkwOU4
beZ7ZoWlrn0p+9Yd5Jv4x8qbfnfKFN7zOXoKf5js82aJFNPZlwP+LQk4WaFFQMqVLijKpc+3B04d
TIixndvJVfQWaS6lBZMq9FfXIFrJPFF4OwN7bwVmpECbbu2x7P5FT849eXBvwGYLL7sH2r6CuO3h
XrBJoEPdaoEOg1/0SrAyVOUKLjizDa/gg3eccyZR+lEyk164u6MFa+4fjiC8DZ2g7UgwVhOWGSqN
gGm/Gom1I5c7QtGMxzrNHHqAa20DUj73xEuzmQEL3ZjuGC0uJkVWoOKCsPB31dX8aP3dIcdTy07E
yj8mN9+9X+DQTZPWHmuHOr4JAgDdRgcd87N4VMVcw6gbZTZScQ5OU7TVzm6UdDbe+HlBP6Ueil7M
HmJOLfZDeeeMhnyekBJl5OLZ/QhzgjBYzsM6AqcDF9BNvsum7JrXiP+PXKax+YFK6EkVTI9KZrlM
RdPHH7y3OpfN5DjPKoQgUJdOmLE7ANE0u/OwH6msCvypl5Q0fvTnEGVqwxSvLnCQ561j8MO8/mov
r8JzU18qZUyY4IlEqB0usna5csG1QVsfaIb239j/YPxrkKo0mDSD0O1ucDNOT8GFEs4kqrQ9sOEK
3uFjSUhiizODEjur+ijbzTaqfopfa3x2d4SwzrZum++adLyWhdWreesKvM110Fg93wvtYkRlgAUD
IoK+NEkSZZLjExi50Rrs+br6+dwUJEn7y1yISTFUilYfPfNSm3LdLz/Io4elOMwRhd953V+rZz0+
ewJayqqcXRsqGyAwvZaXY2UZG+4YTxI7w64QgXnT6xcKseX/zOMLd2MfxWEJTRTPwSxJk+rsAPMo
fhW94gd/Jw4vk9S7pjdNWP+epcgRxoemFT29CSwDqE2fUw9gWY7shtEZslHVfb0rpE+fjRWqKTWa
ASukEGc4Yp94bamGfSXgKaL0xIVyKCX1cj+xlA8oZacZgasfQVT9pnF2fVFP530CfvFtZBxPEaSP
LTh6zVjs/+p7gkX4FjMsA/y19VPhVo2xgxvXAMOb/LLIz4YhuJWBi5u7bOwC5yaXXmoGSFcRHrU4
NH6Pu5zZ0Db4rFHmVB6nizvkftNJZqeB3+tZBRAtlXjtOrg7ZXX2vlD9BS/f0bBJKmx2eY+oTf+m
LM5sXlU6T7/CJhZHqK6hBUevvXKi0VTzjGVRLgV6r+R3GqgHT1ZUNouuhn1g/Uh8iNsjiYHsXnTO
7KQI/yG6bhPdU/Ak0k+8OL0yeu7ZnBQJE5UakYBqWerNDw7QDKln1yXBEKZpyzjkNokqBj4Cyp8u
vkvSyaYKkglaRnnkiz3glOeCgPWAOtunMuh9zXXzbiQFxUfYcAkzUtgEQHVKXqI0jT4HuVVD4DQg
/F2agtOmbnpmBP2tpg4drNwMz6lBWrZUwssrJbO5AY+5KSZ+tJq/0FQv+2BivjLbKBAhnETPdlf8
slG14eUEu6FlRTgAAW5Uu+iyT78gNEk+Y+0tDjwfhrgn4oqvCZ2CWbzaiyRkHtG6Px2Re9fqNcbY
wF7mc4R3++Lz6foZGWSN6os5afIfOA6mAyU8mOLKldocvLL/6z7doot36nPZMtDffQ/XMICfLiob
K4UYKJxsnwwTxvCtU2/hdxPhKiq4BVxy/IcmwwSUPzfZQ+9B3yvn7oJhzFJjeF/SA9MSdCiv7XEw
Bu1vaqHO8sM5q9z9ywTxN5z0zh19u0zT1d1kkNtAMlBJk1SV5vWtNl2ekeg07UczcaQKhLlQSLoj
Pq1Z0/nxw2B+CI9NzHL3gv2X7Io5lWMQSc6EnnmbX7XSpnir3bZKyRX7XNQHNJUQ3Qs+3tSJSE6E
KFTA/Hc6Hzl0y8R/Rb0NsJs0flwOyYe1XY2kLVroc9xK+3ZKwqH+/QkQN1G+WJ/5uL14iTMtEg+K
61GwlCZfgn+MLhGLf4avpmHznBwmm2kWio2eisqWSgquPdqZC29k2lG7qCkuT738s1IA+zHevO69
iTS7iw72RiOMhHpYxr6ktyN5eGVDw5N1c6llMVzXeoP85nU424F74nG0hvPshrexcWA9rzAavWE2
iODaBvdaOBzA+rX3ANjpy3iLkyfb9S7B53gOJRHv6PGXcrQLY08xyGluwowQH3cBoDDfgaUuAsg3
V8FS+8S01gqxuY+HokzVCLwGQrsKU8e3Imm0GH9TNWTY5x6w5p5wfhXotw+/8fyb0dW27rij1lJ5
r/vtm6+n4my3cIhw0AwTF4GvOZnSxIw67qD45G72qBGnekRlNlxcd93PK3JFF2izA3nBbSxBKdod
/zCNNw/iv5CLrZWl/LaSrA+8FbpBZNxqVT7gmgK+jCxuKVpq53yasBAXWlaYCoCq6wCobtM9a6Fg
LRBLFuog7VTB90W4JLSCY+UzW21CawJ5RzTU28T/fycERkq2jDAeQdkLB0YfEJIdSe7Mqls2HdNu
zt46BFOARute2zzgE/w46ZebIAFWqyWCMU9SEtBT5bEqk3HAs/mnkWZA5q5exm4nncspFR8+XcBY
cJiiRL5QZZ7HPZogR1EIxerbHeqRA7oJ3uhnBwQ2xmT9HJTEdiZrGolr4tWcp4EW4UteQ0dyRPyF
ioloxABz0WMNLhxqTE2nKxYsVqWcvhKExewJyiM1QEbNqMWhIQNX+a3FC5/nn73BrdYSzqHXkGk+
vJWigOqiwNT/Hrm3CpHCJmsuTcJLNavMTxk6Ts20QaL0fLvpoGMiHCvLzRW1FxA4Tt2bv0kUA3i5
pg58l0HBiXrdn3EkfyrickTL3P4CcEgbR/gEbE5yIRVOR78dGO2/6IbzLtnC3Sanjh0WGvhmC/RI
bBupfZ4nkgwh+YlrfUydujW/LwQXg+FOwsBARznJMoVXKzQpSYL1IsYPfc1y3fSHrjKEMWx7pUNx
yKtaoz6heA5mHd1qyQo3QTug1oRz0Xw5mlnfvlfgEs06DsYJe8A1pa7mOQqEJ5eE3SqIHty3/W9Y
7VuhFpef8XEUuO2QqoB++cmvKKl2fBuupbgajPQKraG8ScALZ6JmHUYlihLd8rF8lweGozT9nGj2
V6PENCWEzvqwrtCaUsLDo8q2gXD2hsP6+fbsyUYuQbRybIRHFc1+B1G8/s3KEHXJrE1dFm0j4olf
b9Qzys3s++BwHfsw+e32Bz9RUyXVoO5k6NrtMxIn0dyo0LbPaZNW5mCeBqGNz5wxQzgRH0O9vv3c
gCsCT4WjqXn/Re1SHfRRFcZ23FCfc6z/nNwPQggDp0EW0q14fIaDBBhpNRWGAEHp2XX3NBBJf1BQ
lAQenendN7oWZJ4TxYyAlS2C+xFfBlPS+sAQSsR3/+n3zhj54FjTo7q9ZFMF+sl9WzC7mxstD/z4
VFdnG4H7Y5bQjmHDfLaACj7ZvAMzBZmEEnULfSnwyfHxg7X5fdFfyVlhuu53mr6des2dcwwpLxec
sFPdSs5RqQXvkosj/V5ghodJpCITlJEd1/THtC6j0OLB1t8Pr+d405Ey/CQv0GON+7jHdYfsrIiJ
lWWQ0D2TtbY7dHnE7Xk/Dd/Qf2FnLehDIW8Va60uYX8tKzDs7YalG7HSqfXOR074906Gu862pKfv
hijrTdJ8Fwt+ObFV7ScQazM1X38IHXvN8h1Va1NBwj+qzeksGupDO842Tc7EPlgGJJU2y1CgqYEw
jPNV7+RyvhKOxD5yNtgONSeTdSp1HaIx7GWn07/R5On/k2XRaX6PApmO/57yhuJYhX1IUFa+cD8R
WINHyvJVgf+S9BkBNI8Z1RDhljj9jLbQ43Hmmj+PffatGxvEM+KXn2Or2bL86FI6t9HuuqwhLFRR
MJQbW3U8Wp0yccTGeTc8+U97hk3baxQTmlYwPrl7O6VgWCIbAf2cCmRtqwjD1L+WNexma9I33251
vc+lGEpXIOMXbjHiqrk2BLg7eTXjXI3EEhDOJZ+ehugKY/amCxYiRH+gUUZjiJGwvPlzBBYSe6KS
Kqgw1Bt651J6Vl5ldxILh9ijYzjypXgrHSDDMMUOcQmAA1K1T0iImbXuvK4TNOXVYOgPuFEw0RD2
Pns06X5PnAcXtFwOi+CKTP01E3IVkcnbJdQF3p/GuIx7qQU6rIOio1LtfBMxi2mMnPHeLaK7kaA/
VSjslqWmFi84h6lJDtn1/4PeIybBkVBtbcD4Tm71Hp8MH+MNNn7nz6DdEqe5noqPsz+54EoijObb
7ONxHdvBpp989urVkKuzxsx4wk/+kFgdZmFEb6YbsKrpLVrHsNhzVD3DxexkWGSCnpF+KYgqk+uV
LI5rkiASPamFH8cEyP8gsR5Y17pF9DAQrDWwQX5cHVgG8whPL2toPZI1lwBVw3fKpeuSpzJWTBEj
YV7K4Qp/ogFYje/TXuGtwwmbdqjkqLpm/3PiAakfgnrhqit5U0LAXjxgpGxGMP3pikdzwPdzB6Jx
el9o6hW56cOuyL2hZ7KMFZAqS3rD69KQtvCxIjnjUHz/0NpYepJeqnmI3lmy3dnJvoWdQmylVRJ2
VHHQU+xpCxgjp0hT2me84hvp93x+Mblbd9PU+2P8oOYpIXj2g10AgkKkgecM8Mu58e8Fs2FBHBYl
qTXlub/yIChwxFAYZVU7e5bqEGHso/xwOuxupEE3m5ZuAO5wkQIwQLKYDCrkx0EZhXQUeHe5CKt2
Lp00ScOBiHpMnWI+pUb0LNxbOziyg0PLFAlXehYcoeQm5Nwv3Y22hJfzhbmznKcFB9oKdLquwdV9
JmZN6FOs112oH5JqewH/xTYN/bBX7rTAQoAfLjlfeE+geIUtn13vbK05b6ktyDXmot2MCAcML3HF
Wa2Ay0lh2SRhsGhcVeqUpJC0Zah928Wv9Cw2BS3d7yZStQLSn67ifM7cTdbvss9nrMxwgx8H0OPM
LDGPii3SlnnMdNZG99faoEz3aAGaiO+azdpjSagoRhhUNgORqWt6sC49ipfs2P3deMH4kHtDeaXw
MmuWBU2yfhZt0R+jGw2EpO8ANaB7TDiBJ6o8qASv9Mq0HwSBsB6wUINC4dPJ/nCM7tflGRJ7XJ9P
uX52tPSf6QmdCyswqroJ3Arl3UzZtZykKTw4zTsL5XozKQ9LnDHJA+xN2azGmodVR+lUv3WZJ2yQ
lhL0SHAQ11kmC2WhxsraQlj5MV0jL2rXvyLO9TPzOaFxEybObEzTS4qNyYD6OfcsiSOIbCtwQNbI
tDrULMMqAD07sdW46TAcvE+bBNlB4ibKzzrOEL/LTg9Ti84OI2HpV6Vh6CCtueOlf9DagDRyDUwt
pheq4fnV+j8Te0iTbbjuPnycb3yJtrYpftGhnrBUTrICnY+z6HFSbSzeOMfavqb7tnDIcLe6pVU7
p4bw1CH/BMVsRavO8SfQNWE4K/TKBRP4Trp387Nc6fA/bjkD9cM+zmsgXg5RvuIyZ0R+stopex6B
VOPpN36n5dTMowjtB26MD3vVrRjhQNN+YfMoFeuGib7rIiHoVL2nlohKfdXHbQwNcSNZtnYLYUsX
FL4u9pQkN5y1rRpcXMeS5WG4B6xCWQvfhtUl5dv+7GiGzuH9JjZI7Ny2VX6g9dEQcUX1a5RTH4Cf
zjRv0J8ThlvF0Uwr4ghG8T/UhkfMHwg1RfXWY8Yvge63WCrpFqKPmpHT40LRXj0AmYCk9rtTUTS/
6HxDCFPBSR5O0CiEmDS2p/0FwBN/VtprDgugmYqp1TVcG2Qo92s+9nj3zdOEnM3ZNelzpNlX2e8A
vLVKweZYfsWJ4s2m7O5et5sPCtJXjYRnrx7TX9KjPNYLxjr+oiQAq9UgefEYUHBISOVSvjkg6ktq
DwZkrJAje2N+hsi8WVJF+A1l4qkC95D66Prrsn5BjmWDjGgTX04xs6pYPjLw+xvDvc8UDxtvkO2T
o7yFu1fuJpcOvafNa6JOJjDL/g76nQVIoMZ/v91LLQ2PlbchLL5g+s8+CgUn5HX6yvpxTaGumCIY
1aqwURLEhlQAICxxsIiBRCNVn19xLSROTVTuycwgVZgX/L3+yM96Js4OUqVVppdSC2IZ6xEQKzAP
ErJd7BLqzu9LX6eQhETxU1TTnk8PzFsP0tmhKYPD/nZUj4C/99gLB4rUTAWo7FzUPJCJYnqiHzt/
pGknDhvjFGT7QmOnfbulFo2awUiPFxa+4xp3cxyzwN+LTrLF+JB2ZYELW654Sf0hugE9q5fsJeSG
omfKIoIM8ihx9RssDmswBYhLvZe0tyEunzOfsBtwrwC0L703/twnU8SB1+Bf1aBJt0cBAFoBh0h0
7MhoWeze95ODlyTuIRmMqC3KwenkCy0AkANlMnCj3RqC52NysZgYX3v0WWd13QDpqsYIbEbQilsL
ffdkv6hKKTUzo/qDXad5mRMSBSww+nc5ZQdO4Sy6g0ebuHMFyNoGhAl7QCu3qNCXf/+S26vIsyIc
cNawGKywDFJNRaha+7ZjRp/gmnNJH00xht1BJUK/zq/2Y23mT0rJq9mS6z+smmj5ycXVF7BcEy45
z5V6OOwhO23aJG2esEl69uSu/k6oHY0B0XRDbKbFPzL2Al0I5KaSGvwYwMB/g6HMh/PyWm+pnueR
x07rhsQm1TICGVXE7I4tCGde0oOh1QCv0Ajrjk98uTdXIaNtq1CuEh9QXdlIzXY+6Bp2AnShbiYT
Zeu46KbBXs4OiAJ8d5Vf9gBqpZlB0PrpaGm8aaQX27stnP4g3SOmomuluQ9OMecUZM59Sc2UauWZ
0GfHFl/EBI9AisHlMu6QpUEEkN1rog+ZLFTqeac70YrrDZtfYrG1oPu7hvk9FTbOKeKSJcGSChl8
GkWdMydDBksgA4+YedG5yseNm7q7h9TYiHSN4Gn092iS3O+phOwUJR6ivOYUIlNA4U9mHygR3eDj
0vwQR/C0aSOm9CqTnLcL4URl58yHId2WyFpdDn+FHbEN+qIA82QMXDt39tRoVOA0wsEqVJfbq45k
uYeHVTNIhDSWvo2EuJp+s4hihOBKmC6Lbkn/g3CVRmGMLRiFX+skmHR/svOFv2Q975rXaBCBmAHC
4XwXLlKTtVm8LP62RayiF1V4YsbR1hcPh7DsQncySurpc1ZBu3hnc/HRC97t78g/3qsKDYgsdzpC
XjGKQdKu4m3qx521SKRvE/kWW3y3IHK1I+LddconOTpQocAOBbBkMH4NiE5xLZ1J8drJsb8UKxbk
4T4fpMMRj1xXzsaAiqSykqrur0hrZCDAw/mX25I6DhnSRTo6Tt9IAmofZapQgV+3995kc3hL+rPM
x8kiGmbJUm0a0osTflYqeHlzON4NXHctzFuFx0yGQbtGZ35vNnxFQmIvbAPzN2f/oTBnYuyviddo
MueHDgZP+v36W5RArkvK/2WDwnl7j1Nywc2FUdOg0vY1ewoW8p/lKXnwVH/Z2/cVgM4HBjCArKzC
EfOeyip20rHNWjh+CoNpJu3P7GoNqag7i9jIDv//U8HlKVofcZNfe3KuFvbjqXlNyDJEK+C1kg8e
57BDu6Kv2WycBVjxFRzMv/B5vfp0aUYm9KqaJ3QEneY658R1ACtE9jG14gz89ywhddWTyMDJy8HT
yNICrNdfYUyDNUNpjciSCEig+oM2vVkwzvXWHaiHaIxBftqejulq9zQtuz1nbzi6q63r0tDniS75
FypzYMjTo/QjTFmJ3MDbtrINT2ot7+4jrOvgkfsu/w5c8hynYWdcw4UvA+Yh6La4Shrgc7n0iRFE
qQFWWgcDPTaTDEqb6XRKhD3cV3gTIwHzsknJuivH8Qv6qMg7yqL0wKyuobZbhP80QCX6syptNRbY
sfizksswOXRuZbthhft24qw1snA4ItG8Esb+8AO4u8EOW34P834C+6i7sYQdsKskAtADuztuzE6P
zmmb2anLZ2vsNsAOQeKptqvUDkDCDGJFa0f329QzAbRBbNDtpQtXdpo+OWckfLCOmiT1RB8xTAEK
RSWRZYJsObhZHeG6pO/TC/41tCbygTEQ3xX0PPCZAyduWI5450YT7yTABIn4ZPHztmE+98TLNHBD
GrJVZ4m80UGATsLC5fGhEtbjByU+8t830GfhmhRfa9qSRXg56Zo/Uv42DVjeUbZ1YyrzfiWel3SY
RVaPEUBug/O1MDsNOzoON4BffiPKpRu4+QhV4b/uTyPsC3YnxyDzy5b8LxOHCe4lz1kbu9yIuyHW
gzw6nBAwO1gplp3Bs+CXY/IoZhSR++0BgqpGei7dbETMQ5qCR0D7G0bH7Wa3xhk1t8AgcyUJaaTD
vd3oyjgVGOqeWDpo/mKB5AOsbp5V+qe1phURGI+9ysOWMtunlSyX2j4idqvfIRMTKE9sWBwXJKka
YXa4t+YfVZrsTA7NV+OP7GWTag5PyzjbSz1FkZp2lISlEFE+jiYDZQipm1MmI5NwBi5r2l+A+X2R
aRwKE+pdskmb2zhvkyei878+6008yYoXfBB+xttw9NpUyTdYE2uy2sDnT2HuZAuFsEeAC6Zhxoej
/vRJjTCe/Jyq1mEYtBwmkCo3BNDrEATxeR6pDJinC2ZhmkrUX2+lFdUPwWKm29VxkQ/YhgCwA5UL
OKl/uwv4ml7/ZwNNIe551cjNDxG4s7KjJGfneY55eF3bjg7afZWJwgnKk8X8/ndp7UjhGgp9udPi
J6RKW0Iqq2vK2M1PhynKgv+juviOBBXFBwkiyiwmrNUS/9f4sbn99n8R8rkACxvrquj1/MxcBXiF
ewymJoxb2v4Dg/T0SCPzq3BdJaR50r+GQZ6s9PCLoBT26Ui/ifRU3sAewWNIQUEEKFUdZdMHwfX4
skcW6NPiD6VmwTWAbO8VYSwiehO8hxqTh8oEifAstz+muomw6oC9DYdSWAZYSYeBkOvmT0NZukt6
+FzPPNQ7bZmPwz1PLZ+5HQWp3YxjxunWLw1zSrC2Wt0+RqZqZEq2nP7wVrhl9lFdDVAREW6aIbs0
UKLDKg71YlXEuldxmNb/2+Ss9AO6+jwprVuM8K/an3kmZ5zSEcBMX1S1lz1sqo0uy2Xj8ISDC1kn
A7Xn3Gumnf156gfoITsvVk1k18OU84DOT9zOQLaZbOfBSQlhYOcYH7SabOE3GnEK/8IGyw1N03Wz
zIY2B0PCObLPgnnh8P6IFQGcpkaku9iDMazmLap+H/S4QO1+dz1iU0NqjQu8bRH/ERS5FVsiCWzv
G5+ZOtQccrNfWlzaIuu7tacbYNlU7WHjMDBwSM3YATN2i8IT4h4G7GaSs2oRwZX85ow9RsqJ1ShP
ROmyohZV7mOilrrRGipYf/mZdDdupb8Rmannc/RLYr2mE6SyyJ19aXs+yoYEaY1DFTWU9FM6Aq+w
cezAxFxQzTKU0iBVARcRTOgo32dWzSVV0BgfWsAJpnSOFHf3AelVMncjioYPoZF9rMGd/B3Qoael
IDMQlzKhJid3/frP18eGTSGFj/SIXm11iT2XWf/qQVg5CN1t+JytAqenErWfVJB6HgI7EFXmUDI3
NCcGVo2juUW4Ql+LKyB6ojVqTCcGIcLESlJo5gXDrzidnDBicZznBEqVqBeVyMdt/E1qeM5hY0Gf
4CubxKmmTsnaf8SWeFU74GKHEc3pKfm2GagIRYbtwGZRmRAgyrAPionQyKp6pm9te1QTnoe4JbB9
sHX4O6FJRXDVUMztVMf79pyz4eXTOplNp/Hj6yGsxhzIMLQ2rIBeQ0g46E7MXxBYnpd5ou8YBW93
UoakdskFwI+wxkyV9fR2BGQVgsUUhHCkfdSQRQuI9mdo10IWpurxoahPGENNhtZ9STQ+7Zq+j4oz
xZGDWMGW83cVqa5MAcGasfF9kgPkQ9Eis8YVIaMV+sSKaRXl7fTit2MhcssR78SODR2WAEY2kc0t
1b12RMQL+wXNt0di2iTdxGlVMpJ3r5lFDWOJEubIslAk/fcnL9TESWTdxNwhbSkjXx44AB/79IBY
j55siFxd0RKugzVpJ4pkwiNvZ8jhrocEB5X5wvhZ9a2BvJ8+fBHsBgjpSBu83pMP+XF9OnUn5VMj
/FH4blrw4a6Q/ZZ9MvQuZPtCIM+eg1b2nOQrpTIu2WDFWBs3U1ZOVwkEccb86276AYZAkv279/7E
lqF1kB2uc5omAxUsuzYSp4uazX1CjmuVeMvuWsT+Ycva1edQAwOrGDqOnt6RTKYnNbnQiGC66WAI
xBs++bOV6rnjKrgdgCyH9R3anTP673wwqwuNNcKUNxAjRfy+Eo9Zge7aOdubQxPDBimTTeBPMI90
+CevcV9CL1K0GXESj6Fg5PhYT2v2dmV86kZwoWzl5wbPS9D53ECt1B67yVIHPfpq/4fxzpEgBHBO
XIYMqjDzx2YAA0pzff7Tu3OhsYZh0uCsH+5d7Q8MlqkByj+iznylKglp8QtQfYZsuzDE0iDIk5Om
oxr010bw22UwvSJM3pGbZ/5e1gmztLukXkVDOV0g2Kabe7vA8Y44konc7amzHkeFYWEs/s2m8MB3
Cuf2oxmJNw77gDKao1qZcq4IYPI6Yvm1vZcG6yMZL6XKMKPf9hmJGiszl3IhBvEfDYt1qEmg6kq9
gmCxs4ZMfo2G1DhSR6YrNUB9KSs1ToOiQwQ0NdGySAJzM5zpPNX28pqoY8YtyqsNSxsVBg6muMDH
jomj+PrfEjfqbJ4kEXg7SmCtuy87HfA98SwQsBVgm/xwCQDTvuFCIJJlARIl4T6Yd4stEdNbBAcY
TIeJa3md2dJvLL/Wj0aflS5pPpFRo4ztFnXS4KcAEVm+VFqoqGdGMY5Nsy8/vr4A716yKdCuR0FI
sdZudTD0ASnP26qsww7xGcYiGpuxsGjIoSYzFX7E9hwjMkN4VreFg79FG6HvIfhDmFMS0vsGprl/
/ZpuxcAfRcjQWurSEj1NrITQ3jOSG3BrrVIug6j6xXMY6EX0f5B5MCzguDbtwbhNMgU8M67ddQmk
oFgPxdlA+yMaXmDWe4jDRxKwh3OHW2YBVLNRAr4s+J+2uXuBy4L4XAQ8KphNTaFYIiJn6FKmhaWz
j1+TB/ZY4jzkuGdDYF+UHry1KRDQCl5gGW2ias/TMFDkwLCHOo6POCnCLovof951c4HceOMJS2IU
5qV1+x9VrZvWe9wH1Vqu2Qm+ryN3K2f6Yv3fTb82qCJsTkiUdAiB73dldmBbcw6Wpu6czfLwrOPo
oyK3m14BEwX5CfbK1lyrDjU23PJbVSecHahl2voYw9DDYP9V69aTIN77/V9hmCQAUs34oEi8zVOc
VnnN1kL5MWrzW5gnIf5X9Lqr0km9k9pTyyBrfLUrjzgVeQUhAbyBAPFhAYKKpRSQAPdiTxzlHAb2
orwuw1zFVhXiMhgMenBMDNv8t7RSYATYY/ikSfOyyIUmmPzR4paD0xL67ymk04DW8xPXikrW9beQ
gNTnfleCBsUTasxTshU2l1p7n8nAF+iGq6pAzDkoz9rhRX93BMaePj9CeJTjY8MjXR3lFhklbV2O
YuCFKGjnUrGxISxTlobm8o9c/X3AAfgS8/OKtkNzgEgXxMoTHPcn7YfILXv76zd2rQylbbkSewWB
nPxeOejTs0g5GUknrKK0Vdg+Am+rshLXYZzLE9GNAnGJr7VQhj1f/lWToHPjVfMOqqKiRYEq+28f
RdSiGp1USk4JEFXi033mx33rOm+qpxNVMwRmdAmHMIV24KPGJ9+keyBw5oQPmk40c0DDxiqnTB5b
/L/+qq4gb8XynVcC/JNf8kPT4iFwDfIJeR6dPe6tMJ5aGmQu2+SUVLaJ59iT0KMeaCgcWv7VMKnp
H0dHo/l6e6agxdiyUsQ0LcRpWa/CKzbLxan+fVTSb8RBD4qyFaQuV++5EyIMPT7hJo/gLuatega9
ApoqiAuBIjJiyx/8CAMObrwacNUyDNo/tEvC7wF/JxKdtVfteq9phBmNzV1/Rw55RK4OmbesDp3M
Ia8+1b4N7EVeYJt9sBL5SW9Seoc3kcaGz1Q5JPCnK9ogDABpS3ZeYIzjgXS1qNNZp6UUB5JiJ7kf
Fi/YUjnUjLsuPfKCSwvisUj//syvUCh7FbkX0fm/lX/6aM+7YSG2kLqNqDD3xTN2gje2X5cjfBdo
yyx862vAQPUshGjy+P2pPA2/H1McZbAGv5GIHC830Pd9yQ4aJwKNyUVb1SxY3965kQyLRUJL37BB
/7OvP8r6j7h5XvfdHzmcVcXIJ8QloqwyajLS2/gm7q5ROj/VvT36+bSyVYxBpaMCyzfyHL0l9PGQ
jcPNyij4TAT/Vlu67P8ZRg4uyT7bBfWmCPmPkvgnP57WYULYgmgo3AtOfWd7CRQDThat/74cWA63
wUD/rFbsuT/9gN9hlD5s4rdI4Jz/C6FtZ2cFMOnI9aFiAuFv9NnUSIEOE32yk1OxdD2jHx+QG3N8
HGjVjEmgRN50rmoyIqh3pQIO9jdUpBqtUEfGHJE7YWGD1P2sMC63k6NxNvg2zW13J2AL9YPahK9K
4dK2XMNfJvQcdUEPwl4cYRS8o5Y9SKZ6PU7gFkzfoAmJZEi4oI8f0+O5lld7VNDoNue14OX5RXCH
JtOH//VKwpagSHBge8xtFl61pQlbBlACKElOBmVC2syKvFGN05fOCQHlxi5B8adAG/yokDsZTETL
GRVvz2sP5fXGOZ/mvY/VDdyQmFVRteDBEZwRL5yQVUoENsvY/S5rApuzCOPNhf7Nfpz80oMr3JGS
ROPDXsALWRteBbw9iAlmxM7+lbCJRAouHDZ+DN/6XHW2yc9gfjS9+ZYgvdWtsE26G2EKf5LAlNBK
aWV/IKicBfu+KSwyAET8IquUd0cLx3/w/yIeTWB9r8ZcTKD2GDtzDuc4rvpoN85ESW2Z4uXJWant
WN3fgcLO13Ur4chvHHMEF7vV0tVskQqPw3Q+O6J+KF9fN8mvglpOTuNI8KxIXcbQCKk0CTJpM8Yu
w/cF7WyxrtGQESGOQ+gvH/Oj+rP+1fJwWghpMC/56BKLKBE5XolE6OkqJJ85++UBoqjaYVwFlksC
r1OghB3NGKO1Fk0u0prw4rU8D3Ap9m7wpxrPbWxt0Irlac06d5pHu0IZxxOV6p5IwEaVVEpBuy7k
PNRsXurZwpb4Ez81qdm0FZOojfi9/sMW7Caq4FNH0OrWKYQB7j/gdgye47wKGrvJteBDvUEJ+GNN
6A0dZMdRI2FGXbZPoDKc3ZkbnOd2k0n+UQDm5pgxQTzVB6THLPHwSEn+ABo+0Ytzh7+7UOsAyU0k
I1LWJ9rwHyIPdpe6zw/NJIXaDlOFnzsUbgwvATNJG3zxxmCd+1twzAQ1ZbZXua1GW4hjBdY9XmGH
ug9K+GhTP4ACuiyPalCUgLSGaa7EH3GxxIUdV01ZEVphY+eusVL7urZPvPFrgrGSUaHYtPx9KaHd
Il9knwn1DoDRFuD1Or/1zicq0AhiiRR9x0Y9ELtKm9WDfTt/teLCSaa7sAnSrykIoufW2lS80hJ3
c+nw/JV+47vFaAxFJ69XOWBFHP4Eylo0tiqG8qEdvWLxbJ+j/pbqGJu1wMf4VtUEdZANeoWDVZS5
RE70HXHZ2Ek2oOJhfVftlo5pyMpcfSvLaH1jls8fGn+Zpe/GgJLSYdMQCk9PdaVcfAA8jcEgNCet
MoKj9RHP00QWpfGdur3JtIw9+Q3BMAswbSnbvvLdtCHiLAlM66hNz4d7t0mE4e/8uV3JnGugzeQC
/9lbWUdK56ZTaCFWRgsDx0HEO/9dLbonl6IM5AfpTXBpYpOLChNRwYb6e9+Jt/4qexfN6ajpsSdx
8gQIsP88cT4fVQHieQdvxaXStx3JWkzMF32AE7MUtQi/Q5LRVrA5OZVwThXtu4om8D5dbC7mHpag
760mUxMbPw9fNl7NNO/ltUHW7zxVkRde/n//b5ooIhOUyP9iIaYMAXmfpFtULyDMNBwmd8dp9mCY
bPCoCdaxEb7COfXmcZfLqV0+Ejs0dGeWhan0QfQhlngmVo1ATyk3CgX3gtutcI563OUEeTHsgGN7
t165G4eVREHvss4XkNWU71LoRMz9FXYaG07xxwVH5eYo0SPq9POqXobcwDzHymxxPb14b/Gc4cOy
eFNGVwz5BzrMP73b2KyMk5Iv5anymvVRBwkoAKJ3vaxLvLU66CVUDQZbRWvxQ2iARYgifsdlb+Ip
WA4hCbyRkaX16L6XYVdpv1Fgp6/J5JBv/mUmUeDuPf1WMDt53qOoLm4jfX8BE0f0xyYWvr5nOyd9
Q9uvIjYxBShTKIxuL/axItyhbcyZLHZSnf7a4Ih+ryb1YbKKHuz+5tf56dim7KlL+FTkJgkLcSd2
e2v8YHsEjpgnqCwE1Is+OskDZKpsJ59+yDKnf7gGMzFmPY1115f3fbhgM8YXUPI5zXRaPg+/cZSl
7QW+ulI/IgSXlV5x2bj79jSXQnbhLqTWKQYtLrqOnIOZNdIbDzn1nBTdeTNQ/vxI08PzJ0jxiiXX
d1XyngFfMbiigAYHmfvKUT3CkAtOzLXTNNU1W1UliddkBLfnZUxX8G1X3Y+iFpdnHabgHgMRC1bw
na5i6bJCYH/9lCok1t71Mb1D4Gu2k6zyRC0u/i0CoDzPLoVZDiY55x4N0ZQe02dIIcdXKaarQfy/
H2Cf+H36Tsgy6QRtllbXHcl9J0TBTRpJA5v/AZHVZHenurtQLBQ3NBkGnKFefIZz9g6ptrSw/2/u
hAC8U479HCegC0030+5rA/pspj4i+YcildaezwVyronBAAGkQu1BXBywOeabOV4kfCf+0IxoA0MT
f2mZMiie55uy52zkQoN0A2GbZ6sJ2EZvVHlm9Rw6MaWHROE9JdAcKopWPFPFt1U9k7PFKmdH+JSs
JDTMixZNetCkAPIXhKNaYiFLsaZf5+ugFpRn55nTsqtIWszZnmOvEpsp2dEpfscrAACNAPgibxce
wkjZE8SdtwMNNra3Lg76qq87dUvy2n4F77lu6CMXXA9nsrhx7mDoyJefAjpDxLIY+SCXkQRhSryG
7Z5d9aIhRdPaBCsJvuaG68Cngqnp29aMrY6hBqNSO5U2FB8+Ml7oCFShIaUZeK0BqLuwEeud0DaX
DQG4YxnJUFFHHKyqlirGt3wXXVo5MQ4stCcNq+CVdqw2F68IZQP9TFP5E6waBLrIp5/p9gxNJnqA
VcTwHpWNqrqkLn+bEF71QG8N0PodQif+G0E96h7y1TmYMbN1oy+nypljnDoj9jkL/zGozhRyj+3A
2J9BehSVfr1QEi0T/yjd7e2Z1EwRXWyFMhNylZ525d+Mcbros0sT5Lw2izFe//k/JG0ngWW5x1Lj
puTZefGh44osgkDlCRKzEEXPLTWbST8E7K0VMlhACwFWm2Dv/1oPA+L/THpuRKQff27EEANuIGAz
+0/PK4izJ/VSmGejk0BVoelspjoAckcU3k5guW/mt/7EKf0MIl43LZxR1QYw3JypPsN4Cj2NOC9X
2vp/jDFlcmLhUQtlgxjVaeD3yK2gu5fb3/b/Y9TGg2HS6Bo1gA+v4RzsB7biKmcDzHcKmppqRazt
zq5xqYqxGjhh9Qo4sKIXR3j6/k+thPCcAIa6G3NkhzkpQ9ZdxHiuVtsN3dlTEvVvMRqWSpdkFRJL
rUFYI0xoBvHew6sxczuREe1J9VVrj4A4DCQxI8Qapda9GRDYQoon581BRuMgboZmZ4rxiWzUdwLA
304s4HFnTsieoF6s5SW+xMGvQnnFadITfZdreES7zzvxmg5gVhQRE4hZbFp6wx3Vr15kFYWFLjmF
4SxvotaMzv2OTTOIiH+Nm4kttFZFqZvadBSgzZynAKim4p/DCgswI/xK8cyvLNjTybX0btfyWKXl
Et9aRNEs6dDWJd9C/KjTri6n4Zb654P02AG4nGn+m82m10gY64xq5vdDmv+gXA4rAmBKXV/bdL8Q
nfj1l8NzDprWvC+ihVjYT+JmjaJa97CX6dHeNYGIYkERDiK/JVtHLx32WqEa+3uMjeLrBRANpO7m
daKtzUnnAPkM445nAxm6crgTPYiy2dIbaA/FYWlWxYoeZ/Jq3DsJevcZSUlMnvFqkEPGA5pBqUMo
2XBgupwKF/MLKenu35p+62CrgY7LIhvAh1tA1Y/bkk8e6E8oYo4JkY03HdULXNjdNoptZA0VKhGs
ipaUt0AUtu3GVADscNb9drC3NMvvlk+D8yYY/p9hUxC7qe1gBKBNqtnyPtyNofIocoG+b2Z/B7oj
C9IVHeArQ3xMQ2EFTOAgZi3T8LJnpM/d8jLp7JIBcOnrw5QBMogO3ADTULBAsKqnYhash5Ms5Z1e
jtgi+wShodj1US0MNuJfbcFisXXtmcH16kRptK0T1tljvcKZZ0iNCptDkX38a73vQiezQevd1l4Y
17niyMPXjHg8M+G3yBSyP8U5qlR30nbDEAlts4KoJnN+vmltEdDm/zy+yUo4hse9vinIqRxmePqd
pd3HEF9GyXohga5unBbaFD6Ar6Hf09/M/kiEsVSuFCjpTDgsqH+z8z8yMamrQ1eOUFqTfDrrjN9t
sudD23FONYZMKHWb3J73K4MZu7coU7SlTqts83nQWu9yT5Wt4CGncM0PQ+Cn5kFdVfL+I78Ax4QY
m1gvXIBBbrbuWWj1Xtn61pJkQBzvsBVcbZ3/5vEUVIQ7s1C4UVPSCw/8uu/9OoRwnrusrFoeMhOa
RYjpGedYCZqqzEVhUGRz/gGxYfftJrtW3mghVX9oNBMv94zbQaVjQ6a9E7zSi6GVwgp1jP3Y0/9I
3oeKzYoWdjX/CNr2rIm1G6r6a+9uTg+/MbA0qS1Cs4DfyuYNS0B+na+kZctxVIRW1vVOQQSX8k+U
wDXpoJfpW5r5rAqPzJlgBZtqJHsAuRqkLHFAg2KI4iydTDjsFgoEPEJB+HcevHdGfRqSg/NBe9A+
i4l4A/0I7OgRhQiRfz8oKgDnfNb00S+gKN2ogKZTS48zeafwwbAj2tcIWDt+vOKSM5Wwk/HQHbWp
Z3heOZrKAKl3uMylLp/OqDC8YQJEAoBKUw3OEOrsgT/JRVkbcvDrnIrfLpi5kcADb+Wuq9OFSMSP
eCuirJJ5SiAkjV5A3UnvmurAqZJVvQPyLIDXVHS5Pttp34nHDYpcFPvKdXPn3T/aMWGXpaCfY37+
x+mZKpnEfG/tV/1yinAYC6zF0kM+CEzqCtx7CqJWaCu2i9FXHztq4BnUhmV8hgSXaaw/NMPJs6jc
itQZPifq5X5+EUyRmJeO1BoljMMM2B+k2hwPFsllKhhXG5EqEUwoKrbu93BXW3IQdErjiYPGGSCS
h1tHm8+NKgkvV/h9B+p7yU5xoujg9Xg+4O67ykt45mWpTjlUImw1RguOu/2lVlW+M80eB9OQZzz+
ATgbU4Fmuh+AvamCXVhVCVBuPvCczfa99Gok3VRQbXgT5UEsqfkOe2ibpt69Qq0wDjqOsM5Ks3Vk
R2ThX5DGsNp/n3Yc2swljljmkeZSeh9DBCIMf0uOyjED2DwnQAe1ucdkkdVw/u/XhbtAvdHIYoWu
gdOy4oAe7Q9g+UTqCNXp6kcUuzqgud01vxmvsQTdB18/u/KsjmRmg4yW+CTSJDQF6xQu+i0WalhF
IZgewG2ZYZ2jYgesqFHBH5V9X4ZlhFr06Z3w+vJI6bniUe/8ExQp5QE53o+lrda+GAx269FD6tua
+EMCqI+sJ6M1lxQfNCuP06u6bdvXIfvEF0usBKVqB6w+xHgIGJXdpan+mWHkZcNu7Mg9n6OYMK+s
UzHEi22Yyzq8jPMRryEaVyjdQ1tpi1OQQPPLxiW87dUb/1/sp8aLV9c0KAI6dHHKgIizU6MvTH3/
7s0GKEg0Ei5xzRMI6FtQabdC0YyuXKhcrJxikAGzDMZTLdlJjLIcDjZ9/GMDy3BskQ72JUZz5uCr
xPJu8/1QiZWxpavanD0BuQZ6Ru2gqAjYsZvlwyEDEBSvrAgLM4rQ1gbDYg/ANaXAqkuO1TeSFhyN
75kZabIJq58+C3gOVha4bGZymECAAXOHe1jepi8/C0Q7rl1/1Zswbd3izVtpYH7GQIW229ysorW5
kvhHTz6Met6+fekG8JiLPGIqh3Sr+f6f/3ITN+vhAiSBBZ0b3HrtQnpdytG1uvOJiMFWKnOupWHo
GNc3CC+g8ENVWTjiD4A4aa03MQTnJQIOuKk6Wo5raidLTKHLaOANbB1iziN6FXSzUf6FyfVZf4nA
d01XHYMeheS3qFlvsT3kXAfkWwUmw/vSkI/82v2WsquktbpoX0yX84Lj8iRStXgPrOhxAn/w6AIg
HSZCA/RjdBts4DshF3eU5jgsvxUXw7/WlgqNlCjMdaZr+YSfeetgLteYsbp5BgB0DAf1+4eKPWRB
tFcsuSiA+8kDe5rFsXRGpEm2ErEjgoqwiS6jJd5jjhyiNeC/VqkqcEkFHVRAJyMhiq7Es8b0azv7
YnOxQtcBZhaAlTNE86dUkCaZ6V77QhD6pxV7wjRs9eFNtY7sYAReLjofDK7favPg9pxLFZPpRw+Q
UhnmiC+cbEkbYK7RL6irJhr9lW62gcsNHcP9M4rapZhUBP/p1r4PsrxFq9dsv0Q8T91o6ZIyl7h3
vrIjO8CN5FRleOPKbfQHyoCFfK11zFtzh1TYt02/3sZIjsDbFn4TFUDs7oENhE36f9X2DJzeKJyT
8HxjP7LQQIgB+1YT6ArWdWjJ6PJhwYlZsq2XE6w6SRIu73r8uQ0EN3NEIwwUgDgdDmn5sSNmFLsj
4H6K92BI14qlbJ0t5VaI8fxUb59KkLHQxTLXlx72Cr8IrDgxVw+9UZ+8sUjsHO4iDnKtQfwlOBuf
e8p11cIhq2Pp3Do5zclMw1d53JPnSPyl6CXcNfj+Rfu3CUUCA/JI+OFiZg4yrtxvxpYNuTDl47TH
7DClVm5z32jlmo3FZiHarTpfwrARmj6lVzpuoSkwt8GDZagFaTYAFlkeKeDO/4zAjO8oSpU/pUaU
hr+ITUm881U4B9JDHFr2IhpB+o7xxvVMgOU2FkcrMprZKjmxb3bENrseg8ljSmOiGSxvjgDjd9Wd
aAHPdnD7xb3P3DQCi/sIW1s0azTVPhDgMOcfReGXs1KhpVceZhmZIcwZQXSa1nqvBKxlzyB7v2RF
PUe8HmJXV5GxDzASPoWXpXboKAfpbhJh08/5I/W7voVo6WXKOX4AIXtpiXLGmWwhzgy7YehyrPgJ
OYkWYt3h129npCJ3loWeeoG2r619gHrVLkh5kRjH+Ah/xyjIDvP3cAnPG22OVJgCJRUn2iQ4/p6Q
GfadQv2R+L1BIeu8ECstKBkt86Eluoe5dosN46Maj/jASLIHeSHSofu8r4rWKwFA8P9wkbxTj4VT
tR1cN9tDCok1m/XZPx9XpOI4ibICBEcwAiLzemfAFkCd1/VLA5mesR6FdAFDdzEljFjlKjviiNq8
xmaTMV+ladrKhcZx6x0xjSPStTSEw4lFWZMF7kd/foHJE+wPABV4o/fA5RtXKC/p4Xl7I7XGy/zu
Zmemh1hbYA/WSJ4CtcOMK16TCiiOduenUc7MU22jVbkNGDmvfiH7YV4bg+YOaevZTrW3GI/T0Mqq
3UDcNlB7U/j3ghIXWEr4vJ+W/lOsyIj9sFksNh4YV3iBA3Qo4iNKxAn6KKYgJ7e19uSvt54/Np+N
26bef14hfiSxESR0dDBXZzAv5rwgQGKV+Dt+f9OFUQa/I+gVxwRc1zaGKZhKGHKROdOVxnCJntDN
NXfMrEW1iqKeQ/ViacSn7wgZ8PDTXwWON06pQ9M8H9wQmH5IRdyrZfKIUNZtXccaxWeJ9K9mMsK8
XZbnyTU02hENXr3kH/czPQu9f8ia32K+maDCzyCPm9Lyku28jhla6T4wvYgyg00qEALp6ajyFeFt
6C188l/OnGNOhUDrQXdA56iqfvY5cKDfzLN7xcW0pbfvxpuYRIpYnsH08HWig74n6pipEiOKR3TD
qlfCqyYHPZRunBH9spf23lfVhCQUddc3TWxGwxVMkluS0qLb74NkjPKfatsLM5hZVnKIotr/ZqQj
eAxCVXGYwR9TcnZ08W0B6yEJEG1Yblm+5WJahzqT4kOadysaMPSJXDXZdNfC8HCy3E/SgQyo5FaE
dTXc+/h1W/gdlFQFjli9nQeFduVEImCi/oCjTJQefZxRLZyFgUdw6ECP9HjxcKTocOFxpXuDqYdx
rSRqKLQkD4JSyQj8fNQUUaG9HdqT5YMGMMU/dyQDpJmOydKPFq2aYzqoKM/mVrH6ZgzuFdcuBLSu
QHXI7seEy4baflqN4qNbHDyOgIhO5IbJEHUnCD16YNfzgvYqrXf32C52TKVijv3uZjbkr+lQcNrr
6+gNYU+goKlhHJCbSENMi713JBaERsSzBYREMbUhbS+GebC6oS0DqfP8qollYt/uTYPkZVtwNmm7
oJ9oB3wYv56NWq0uoBflfK+a6EQo6Kv9SQo80zojWn0g5Btoq+5dvghpw9zkn2uWLmAu8+oL+/oX
lj22oJkKnt0AX8ErbhZDyeD3npVaj7USc8euM3bPLDjL9Ox9ctjH6rTfPH1v2u5cPL/KRqipVoZa
cWsFtQ7ZV0gPtHmMOsbNPOa4jkrv7XqFwgLXjaxbXknavN4ERxCtC07xNIOCOIu51QTJJNQXnB21
WdsvCPWLM+wwmO5h8DF5aNdDVAKvHHNJY0aPumiM+YGsBu0j/WG8qxhL/Wcxn8DwvrMh5oflKQWO
SkTATo3y1+26beZ5UbrhcYitARUvQ+yi+bCqEC6driZZjTzqnmPP9K81lJd3xKKisFH0X7LOu1dy
oUovrUExz9W0FLZ7LN76laTNbpJCZX+aY0KTNvxSyU5/bOitzd/+HenlixzdvmOOIISR/8lqVje1
ubieJ3317sJWXh4S7vg9Mq4XauFY3IxmIoLCIQnMhc61DNIJGJ5gu2S3VdpNwOSZtcYeU/7xQA+/
FeZF6OcwVE21cWM+tYjuYJitNN2vK8oUdqY0dy0pjU7BuLbMgt1SxXGs3MCp1H/V3q3NgZq+7TED
7n4t7gZyXlCZLqfNoBTerXBCvy8NCzqFjYQ12nHXH0fvx+8aZnOOgcLrqLiKkFoBdYEJQvOWBgZ3
O07Wbe7NUPKS2NYjauMLsdC6eL5Q9m29LAq9AvzBNmXDLpLS+8rIVKeRv4FKxw3bhqru0bSxXG97
W3+8slwpLvjmvBZvdpK3bYNEtZBA1vTdnbZn3pPqSPDrr/sXqkGMDGNtBU7WmBUAlXPw9fR2GBXa
VDP2a0yb1/jZy6cjH/FNznhIAmu0lvUzODmYfuK69YSxJ/gqaWjIIY4VW4R8F+zUtfGS4BuwoYHO
42PFU2xVhuYyqDi9V0DJB/cVO/UZmmIbJ9qFoPBN7Sd0UTIGbhKXtMVqDyA5KkzjayEAxQ21KYOV
VgNIXSrAUEMX3cqi/sgzFffuWBAAnSfmDNn2bvkNLU/yZ/M29TIO20lVHkygzIe81yUJMOM6o7Lg
PKyzjal9bIB6wsJycbHzMgrsENm5MbppXkuTWeRyMc4ZoGCysd7PW1nqpD8u12VqAq8YqBbtzfkR
r911ZNb0A16xwBqsTfaYB6hdkt8BuCOcGoL5QUPu85Mp09ljTqlAeOI+8b65xeRb5IVkOiWBoXee
x08dUgNPdvb31A6NGHwT0YSeEq5Z9ABYTRMtojKUhjEzADBH+Tp4KBBxJLcpl9pTMGmCOKAAdgUU
lOLNUK6VvdbPGGJqosFzi6T7VIO7mQmAIOZMfoT+ShKchPc7ooZEbCnD1eZXDPtGjKp7tRagzsSE
vCZX30c9CpcNF5MpbVbiWux0jZVn6qCKeoDaJJpIuZDbsQUpN5MWJ3BBBzUKodzFmIR5ypUjRxnj
OWAaZ/rsdYW5bishCi/02bMF58uaqrdH/01EXRC8mw/SySXKOdUUgNCMGuVw/TNLwWjRGvC7KMQN
/knww+iDcY0Vz4y2V+9o9EQK7yxBjVqSKGIn+3IPmSSDRvgMVAOP+OpRAIaSlLGB6TxqrMjeS43Y
4zZpOnt1aQ+ErHk1cgmHW/r+gsGNCD3sUe3hzjy4llaJ+nE1xK7DhJALWma3G9adu1+h9UOHw8cZ
VGilMJPYI4U7UmHmar2mt3MW5NN+I5ZAXDEQpg7ag4pxEJWO5hcGxzwuIucCI60Jk8H2yDqmJiGp
FkUI4wPRG992wzfAGeMQasSo7T10j0ixMskvgKKNE3RqSFsCxfEm8l+A4/ValSF90TtFPuP5H9Vo
2RDNCUrHGKGuw2KIiXg56s0IY0WocHMmqsaRMM1eFWdhMANbCgBk+qMiB/n98kgmFvXYFtQCcd1Z
ewq6K6GJDqZKWjwAdhv/HoglTpJbYETXT8LRk22RE3s0BLBbJLjsMLt0IqdsHtxdOFIKFys2vm99
TdDgTTSKv0OLJVmzlQSTLPrw1pnuW6vp5UwGkqoTr7nADVCKbHVlIkTzW7T76IZUTd+byS+pN2WP
LgrJ4EZg+BjmI0O2a/DfgNzqWhFoR/CNQ/Yn1p25EvmCpOFMfO8wueNVicbSvmwenh2Pcwiix/3R
jRutcu6gosOdhZgj1pjHgbhePW712OGwF+Raim6jHLCwYkdCxLOTtXjosj0s2smtri1wtAjOAiFn
8npGq7QZ6QJt2J3aWmM7g3MWhpA/7XiCH++x5JAdzPQM5YQrKclaL8kgzn4fo1rDNodX7MPyyN90
lnQMQAHdkVBWjcrsckFjsHc83iZI6jTTiTpZDzeT8hBt7kEXic7OG3hXkToOdghgq9WjWFZZDrRl
J2PoeQK7de8MEe2r8lR4/sTcBh980Z4lDHKKyUn9clegYwX78NhNrlgfkxKPbo/QvQjf3GbYJMrR
vfejj9kQNK1yXZVamoXSByl+fdG7k9AOuJC+uMPORKBoUuVXEVdSAZUpl59fFeUliizbr6MMP6dc
+k8EZIyGwOy5fUVyyWMYapthl700Tf+BO7Lu/0NNPaGYJ/pkQsUhSU2bUko8PyPz0cVguAB2TZrN
Zm0ToEunVmMlhAPoxA//0fSo8V1EbVI0RnRog7xGA3oZxnXYl2k+VIi93GHgnoDWioEKjW8UCAl/
GB71yeujdAvLinkVDJqIYznijIb0dpczgpvkVpFagBKOjB4CrOt4Ew6KO+EzYNXrhsjZb7arRqjt
Ozy6LyVetwpTZX2eXEqHG5wnWz7t3Pmj8FBle12z9/ogFz2Yy/QjDTFpDmWmAsBzVYm4WwbUO5WM
BSIWFQLtQ7lxGO36cSNK+IlsDSIaH9JVY/kP1+bUv1R6Bji1No0+GuozCuN4YuAZ/RzF7M0aw5D5
2/e73evuHS6ZZnkywJIJAQjzGeFA3hSSN81Mek9iCIk1XOSAvv4yriPTV3QuYkzxzqrKz3Co1st+
p7Rwj1J7jT44MirQYIXuLUdSbensD/TT1Yo7qpJ3peCf/CI7EVOxI2K7REPgfm5rtKI1c6G9BGD4
h1VmO0fpqwRfhtE8KXP5mxdiID7WKW2TuR3wuXntLpjIRPEwj1aQ5dl7pzCp4Wsx35OLVEeQdZs9
Xuu78AlR3kNAActO32X+tAgt7l4Let3fbGfvbWGEukIl0dlBtGcRAt7fvM945Ih6vw+HyT4aAtBK
0uGJWhqiBl1hjrDBC3IyzZsnngzLNzecamVcKwwgNV4oLCZmV8AaCW2WVPEpwXqBQsxlv7EkQVR1
TACOdibr1GQHFAqxEQ+5ypxnjVG5dKBqq2/PKG5HB0bXnz2AerDMupO2/2qDK6yEf8302++BQX5B
dQbZ0aMgv0ND9w8OoSRanXIa8H8R9MGqCk+J5lsQFF3wv4EfDwx1Zfq+hu2gRtuco857C0BI0TwT
LUrG2viLLidO2goUQdw+1AXk1ItBrMtFPJltxbHTdU1HJeTIFufaTWcei7iYXXO2uYBNKLM2GbzY
yvDYV55twuKCzT8iQDaEEdKed28YxpMm8AYwAHy+tnY/7bN7r3d9CQKSDoLJus33d2bktyjfrWPh
Y/Iw5NVpAhrX3cgO2kSyWXW5p9UTMPZSAab6gBuKJZEQ0h3AUO3JJkdYotyesjYuFFva/lEme09+
nt3g7o1aRW5+Om5j54U6ELMJQxSK0u5vlQihvZvlYQCWOAhVR1YCQRDFmSNi+n3XHCaegAxSZC4h
3AEQG9xtEQaf+ysvLQl3hOwxPla8HYYQa/lJW+uAy1L1GQ6BiO1gqB/BZhYWCkSxacZUqcxP9bjE
V91gDmur+nu2ReZWvvgIDcxeE4/H7UvjG+/MHvOy4aI32diJggCx/2T5+5v+/g5Frtz9KZY7mJ/T
6tkVdFsaW+IWbVTgoZT1tp9VCkddwdnaQtGtf+qRuEcUWS5c7Ii49KnFMY4W9wDtypU4QYlb2IT9
17avRFADlJhr6rBQ46tqCTWNYt60sN61Y0bgbh6MxJuSIFTrLroODl/qJOrpv00XiKCqCVlGtRSW
MQRn2sKeeCCo26wFOMIg8W0Q/hCK9sjfjfnnsMQPej+DbJ/tfoVzXw2bWgqUW8lAbR0JmSTjuOiy
wpjnMf07VG/mz8K8ouE3Am6bWrOGTIhBf5h8saMBMu8qtVXTqIvIq1LLn/P0UD6JkhATb92MXoWW
3EQnBhdhWX5IXMJpTduQpJ1lr5piuqAUMUtj4EHnbG1XA4FPVZZHmVZb47tRBKMnd7ojljUPZEp3
RHIWh9XrK8Ix6AIzt2ddbi8DQRiSW1r8GSphFpR1ALNEvz1i0W4iJ0npKBo6TLRg0Doo8JMCaVvo
cMnuY97ByKMtMpFb1zpVLR3ukl+Tf0Hhl4myl1nsP8oEztvf/zcVMV0Q2FGLktQJOXt6+F8x6cjl
1NFdiYyWnnGZ3Fg7DeY+GbFOdOVTTc8TN8/ZXVZ6t6vtQxtiy8HPwcgH+EeHz9iz+qsI4QgNPsaW
hDR0WgrwL7uqLgPikaJkLvjt9RtoZI92h5tMZoF45gbsR4N9lh1POOkmdbMtjj7YpgVjKjj/dXBK
ggJg0n/bzgenyDbJUrgfSVtLg1Q/Fd8J4MpV4+j29rrfTjOBUPjRVuhFTFx4Kben44mGKTTTnXSm
r6KHmjj/5IuG0xEZODVasIkPtHdTEldHbjV2plueck2TmaCClLh1o5gAos4VvplpITrXMmlI8oy2
Gma7RxDSMMWmaMO4nranUaASnveBwP9hiCm8Mb1ce8rYV/EslWGOdGd7Go51+QiDnF05kSmTLDmZ
Nyj4qgdfJrjIOl3L+NdUgBiEup5sIaFn/Oqvs4kLuwB1YkJcLVcmLw6kLIjUEfZi9z6T9C5xm0Lm
FALyLe/0uUbcSx2WeszubIIOG07ju7q86NCohVqwgx9nEom5iRWWn9GISFzyqhVO3QoJKrwNyBwz
yy7i3EdNsWO7lPWaj3UQbeup3ScIw5wMalPNizsCJ4AkAwfoHDNK9oE1mgF95OJFCkNVuyQUYGdl
FEc1jNe17ePZGlb0tuk8Y1oUQ7nnPUuFpzvatWJzOmr/+igzsor/5bGFvsNf4lGmCIeFYs36+hzW
YGry+I3LbC6aJFVpf2DUU63Af3L2NMzXNrDo2Ywo2KIQbqRFyeTauV80g0kq2mABi7fmuuQR+sjK
9UZgbv4jK+hQNwGM0UlUDBq+WzgEjkmVZTEQ3l3hdYzGpEyTggRta32BAOMUAdM2/zLzaGrZom8X
M2vp7xOmPK5vOgbrs4WPC5ko/oBUJtmXu1pt2UODwAerh3GuuZBkn88/y9iWrXVR8gDjRoXdZcZX
b44Thdwqdw5/PLKpx/OrD/nuOzWy5XI1N6ixXG6YquY+q0w3yrSDXqXH3ZTxIgSsXBqlUUcFNoTd
WoXEBPfojw9ocphI6RTf9XlblXwQWiUwlznVXtAS6crm/xN2kI53udk8rYr3Inz81jBtS0E0zezW
0778nvr6kSo3wPLT5I+zSqIY+FGJ5+Fu1t92PoVt8B4m5eZQCdK0qeuw3ETmQCYp+G1Cp39A3PPP
m+uze9/UkJonu2wgzBgGSrQFOjEVdZyXq/amZzxn62Nu62NfNefpN64ETEhelVHbvaTqwRyt5AKb
2AOHQqo+0IjjNkWSLg+tvgRgoMUYXUfas528fEP10HHswyIDYG4q0n0iaeVlgOV94sXy5ghI+TrS
yD3d84TZ+tuLOsgQnGt0CFquqqTvZQgwD0PzN1LQB+r3kCGIzmV8wqoYSrz4S6ADXztVFS2yaRSM
1ycM8bOXb3e87Nsi39nR1FaAjJnksuN0VLxTro4S6R1jIfyaNkn+2oRzsz9RXQmaHtz/o78c7K/p
uuipIZVcRPAlIkEH6pSWcLi+5gizWZMxavwDmj+6+06RW6y768Hd5uK7CrRfS8pkQP8g4s1YyWQK
c4SSWtFs1EXEOYx5e5AuyQ21qTZVwc3oJ1P6xFhWtBwyMp5CibBWrEOBAmHA1/tVirA761ALKdAx
71Aeg0pOZDVDfUfQ9BpJBZ2pfB6BDJYLsrd72gwvNNYs1waETNrcYKLuGGLL51RHVD4nlhkJ0uV6
6YAy/ETtNToAdsMYD1v2E7l3gUQY2sYRRHYxlxTe5+70br3fWqh3zewanN/HEzJsW5/8szUouEIu
zXPbRXUGcEwGJShwGv+jaCGvsj/zAh1L3mgs6xspF0Lanl7EI3uZi4D6VahMot6+4K1RJbMtIH9T
ESHOuvBpHXd0msz2mBTD0C6lXH7uB1I4K7VycXAIru9XyBawkrcFBN6CTIP7JLN4zmrg0QI7YcuF
dvvkJfKJn5aIWWoSgOI4kt2AciMdzZsuRFYZR5z1VHP9bHM//wtNETsImV11Zv0CKzhZkTAqXQGm
o906hxQJAsNgB93DbovXrZMlxMoZSlKUZpgU912mnIVxzXG5XnXvijGuJfxPIIBi9w2yPg9Y/eqH
p7Wvbk5zymm9+DJk5JBr/6N8aZoJZZc3CeWOyU8rqU69GTrn5jx/nJHBCwxM1gx7OSNZ0uN9JnLr
wrvQK25yzxk4lfWX8Rrc8c1i46C1QQfJGnqf0ap0+C3LtHpI7s/0Mg4Rse6EeEPJ4J465xM35fOb
FTx9kaeug22DW6zqsjD6NBNK7xMcO+bxLWHdROYcLCnR2zhjW5Qb6CG0LBFQCnayOAtsWJodDiug
rRxo7PbpPCxItr64OYb0FMzsMB/TXALxdBsxW4NcoWvJxkisyp4x3WK+9Jf+oqeZsdWkpHoznvTc
v35tEKZ0XfdJD/5IcmMa/30sUPb2OlKkLFBWNztmC3zAs2dQLSIL5u2IQHk6vgl6qqnFl9aapK+I
AUGkXTynviqu5aueGR9xY8KvwsS63qdIsUF2gYju+nTW8ExLV5Be4vLkhddJkyPtt1XtJszUIZ8x
kzf1kY/SHJFrW6tqJYPFbD/mcWDzypDo02z0vEbCzzHyYiFPAiaVs3U1ASorA7a/2J8Hiagj7n2K
ktfDYQ3cn0Ly/K1myRjX/qfUCi5A7I6d7Ogp3/E+ND9eDlM7QB8lHVPlvqvGJ+KKl2Gc30vFgmaS
oHiPA+qSjz/ortFfL8KaucV3HoKN71jrsbt0sR95A3JCr79Xnkngxt7Ky41grqdtU+OO+jBK0JSO
qnTAdhvJUtQdpT6wAfD9QqfBvLLUuEKI7YL7P6GUeZ/WRn/MRY+Ukijds+4t8d7q18eQVc0I6Ryn
vwo8Mm8McQ337yCCDxnyK4svKgrK/kYP1tnrdc/fJhacoTsV0Mh0YqKCf1XwNnVRcb5PG3GnlCl3
1ko3vfwWQZOKuHTQ4IK87EB+YKQix/dEts+1UzJR2d4trb/Bv65r7KxFPMRTsUXsEOM6kMOsRv+n
+hRSCzGDjedkOiOpfEXPG3GXlQQGWTgWsMMYLlR6CrmS9D1VBoxPKWJBKm020aOuVvIdxWXn9oQM
jGUBuHsyFWUpxoH5yKohWSmMOpgGn5ehRTVpCC/09qImhKN0Cwp2Gd+TrPDajNh43n78U9FBaUWm
cZ21GpNiPFID5BUkhQKYVzIVgoBoxo7G02xFrZCtw2jNOgJSUf5MjulcK2uA7SBRiVLXAUSsd3BW
ObAk2pLXDHeXYFO6RyefG5cXrYYivyhcU5QrqAvO5JZihBbKuw3/iZUdImWDTKCLGpEYPVfri9GN
nNnIkT8R0fp7GhVv8apNsU9B5MPXUwPJ49GXwuAR7LYrLOc1LHQGcCWEWrngyWVoPXZYnyUbjyUU
nlkgJ1R9OhsUcJ+oox63JfOPkF3N7lTa7zQvKVXCwo14rUFxkE77tMmBqGDnmo/X/ZH5R+tpkO3X
9EoAjn5CLCbeMbdoxefMxJpNXm+iF+oWiewqZ4QHdAfDgPauHsDjwYTiABO5Ek1KxZdXOXnqemFB
wKwSqA7VCzABsWae113f9MkGh/iTn9ESJUR5rapLqr3kEeQthlMJ8Gngtk4dJatklalKLU0IhuqS
KYgbecErX/UeOHNfKJuUzOkktM7iKpaUbp9mAVrPXbuNJVeDr4Jkts9bKH9/YPJIf2riaPFIZBIv
7hzwjdKzftIWU1P32a7sMmN1bR/d4UKlHnY7Rw4JNZdyNj2BLD9cry51NeIS0vgcnbIAe8C++iDo
E09Ahud2iel/Zyo6JdIvmfgl+5CPodMRQUqeyAMB3wiF/yzCTCN/nGZ06ix5LJtW8lsd4f23pt2a
qDLwyjOYL3gc3KXBCmYhbev+6f/z1k3PGUB4JHd9qOfi9rMQdM4e3UqlKJyjCzRiR+Cs6bc9g0nI
eLTikNnpUkpeTfrh1gVIfGhw1NIuuqUm4c/f/JQwvMC5zF8ptlF8/FISTwOKCMcWUDfAjgQvMoHO
ikt6gFd4wC03d2OqdotxEOcY91hzZftT/nxxBKolV7lDBs6Mbix7x7e1SX6VCKrymxznpa/2Keil
7FYfgj48oRGY0kkhH3R4sGRGKOnJW/D938XS/K2yHYZvAbG7Q67BUCEHf0fd6L+pUxdacqyAW/wl
6nq/vVzlvoPHIbGDqI8DV6ihHbJdvZ+ChHF6z8OgHQQ2HfhhZunKs0gD8jAVvsPRUyAy7wk+S3sj
GuAs9d5iBoNimbj4YIKfQ4MA+29FQVkWdtqfinxvRp7EVUpBhSafqDreJl/WSbZ7G4ex28e7ULx7
dUZwK6VgyQyVCan7yxJGKZ6rr6+6/DEJmWHzvFnwhH1p+eCUSC8I6c5FVHJ6a7PtVfXKbLhY+HcH
9ifPinkQ+e7Ie51tJujOlzMuD6hhGbKEh6uVutWdOE6XOHM8Lp6aKugaoLDj4Nhhlg8ZYcevyDvM
PjXKh2qgCcJHlHg1AHRk/I4GW5/rkcc/NzH1f8DfBBL56AYdCNQHYjZ7hj1xAr8l/WAzWzc46vdw
WhkN3GmnDSbrqxZwtJ+a/VUg4g6ME6J6VZlXvDzqWeOhxxpfut4Vccr971FExHe9db62cvvRTV8T
ECz3LlHhb0ItibpwNMEZ46eh1YlUqh15GF5Q0p50vxDrdWdU05uB1Tmc73h7ifDB+eoKg4/0td1I
PaVUYLWfO1jhLAelsQ2L1ATdmGArEwOq1jvT9zweiGRwwX7935LkfiLrLWpgFgOBzvO6QyLNPZV3
DYGmy7N4zA/+cjzvakW2A+rT/GRXROlwuF5ANEilQb8m0vJGdJNyH3T4gdn/NIj+LH4B8UYuadFJ
J0hxRutxkTISS2S95YUlUbdInV/RNLbwj4i8QnmG3OOpeideVqRJdvwgeN/wWPxZQm/if/eAWsGM
k5f3076gSVgTJ/V51BLMPcRsbpcPTWcqMoWNj1WrZ3Quf+p+JFkEnqjYIkjai4CL7zJmGg8dZvMO
5wWC1idBuMx4G8y8uTRIYdK2VsJszZ0acvB2NSvDA1VA/1nRN2BMsdJHWhZe34pSz7MV61OL7LPx
b7CUiofGa6tT6oxUtKmS40GWeYNRhAmdmbHfc954OkWFBbhWBJVt/8gKsleH8khXrBDDqKsMWB3B
5Lcy7F0jehPg3r6kPQT1ER7szczkSMU+fKeHRlE3lVbKmDLbtolDHEgfxwVzuB1+1XJhTzY4eEKx
nXayu4K40mPwEAHEFH/JcA8xq5tSeRG8MYqAPi18QlVw5NvV8W005zqdRq7G89KWEBa3DDtqmlDb
32B3nzbGPfBV68s2t6ywq2Oa1kTWWNJ61NFgw3EajQi/TMdcoEc/wZl9z/MLLSxtpS9npiszX+ni
TepxeYmZocctN3XETSnBECwoITCo8VxJWkT2aCuAoM7U7W/rKgp5Aavy93l5znSNaVDbmlhpV8h3
0pM4NCxk7KysqAg5+R5dIh5nWxGlBKnaoOv9diAWeHumUwX0PrisMq3hzdJi8yBxP0+G0VDEUBIE
nmluzJi4S2k9NLop7S6Y1KToZSoHKDQwvumWSJpq0S7kdlhaAmTBuLXdohOfeFtkOtvCgxW79oFM
SPsdcRy3D0XA1o7PRIemiF4c+BgzkYBgW2gbr66+P43jtRL9v0LkEPlHATfyh/rjH8fvp8qR38L+
relNUFPtvMsiVlb0mZfw5CXVtDinII3zquEKAUIN1WR9TfkgQ5KRQhFXX97FtWSIi0nyRpjXYTTU
z/vCZKidDlcBhoYJf8r+YCPN+izpId3rcHwKGbJH0lnaZRYeMcAej+talaW57csIN01W0fxRpmzc
HT43o1Yvb233KXfT+OKkVFCkK8p+PBBydWOlAIfRXskVc3ijqh6KV5JXq22wlOxlNBl/XuBqWX6a
O9BCJJureOCuUVKqTGrwu6nNqfInGXNqJxYoJjSuBkuGprvOtu/MkjFKZ8lgVEE7N7/8t9ePDDe6
BdFT9fwVfFt73ZBNzdJwdm9Av4q4kamMe+ndYDKetbQd6ItRiogQUdDNJtJ3LhbKqbacSW9BMzuR
vckxLF1HJBlRbpOJgDpLT/f5q09kmdR8RwcIKwVqzy5I4mHoFSGRtVIM23GO8QR/XGF/pq99hwe5
xYQVhoeMMtn29tnTtpHuPSc1JyTMUKtiPv3a75Ufq4/SqEgGjQ/ihdT3O7neaqaj/1s7deUjO90M
j4oALcnWg83PlRGd2wWe+ATREseZIn9D5IxY7bfwhNZOModmGwzX0jFt5PmHS4leMlwNoA5rToLu
EUCNz8PCEBFd0ppRAYQY8qo1B4ccJF1mbVL2wEKBJMUk59adpcV866Qpkot1UWlbV4VCBPQAB9nk
h3TnXbF0Hrvhp2EqzcUKSZ7JdH1Z2zyIipKGpqwxHATcI8xkyuH67S2Imkesb/cKASsaGHFhc32g
GX5ooV4C7q7V1XJNgvd/d0iZuuxzpteWrFtGVLlMZ88nJnCwNHLd6ZWq48aqpl9p14LZY/KJ5ZBA
uGp3tFsZuhMziEauEW0BOmCApPABTa5ueQLhBQXps/Na3fRc9qU6iD/XURGYlemnxOpa20NA3EdS
e5s7iNIA6FH3+5G2NT34KLi7eBoqJCZyiRAj2DOBMLBLYGs6+2mZT32pDPLsXflRgL4Q40TH7x8Z
/5AUcCCGQe48ljWF/qB7MmXBFva4IwMWKW2+W6C+BHFOHJ+mzatBeN27N6jEdnRb8vbYAQIuoYFw
TgaXb0gKxVBom1M7DJJX5qV7KcfYtS4KlUnTc6EPq0hVt2fc3DHEJXgi2wemB+uAJKnDaUDxrVT5
efAh2cKtW7+JKD8aZ/AiKlNfKzl6prXyimoTmjrDjLTrkKJY0zmgdpZy21U2gTkNDQOvTnYR2x/a
9qH945Ox2GjiKQLUY8vVC3rJ2lVOGhltGefpDaQIyxRzrc+v1j/n38cv/WwZo8RkWNi3J7UlRfC4
d+PrTUrMPe5paAUm6sJBYxxGprEVXYH2/Hy6TVe96w7sArQ316wlehPH1Q/Dh/zEW1ewsXlcxwHU
W0s+3rpRQTe8zi/adyqiZFCGXLyCnAx2jeL7iwQYjD+FdZa2FXQsIz1jRo+rrrTaOOSv9iE1p7Sp
XDAUugpsaeFVc5zmD4LSSQX3lxa2FEERW7XuxdCiG+j78+3nSwx0vjFILltu2c7QfcoQVtbwz7ve
qYY31JBWcgD5mbkZrDcCrRlH7Z95JITKvQrhUJIePniWqvyLAljvL2hPVZpHsfgLPhPlN5ja9zBX
p6/ZPbwuQLaqg19pWj9Ym370tXJMCk8A/lPPaZIqLUVbtDwKDCB6Z+swbDhQ2hQrGiShCFro6LCp
8obhpOqStLgJFC6SaPmzLa8Xlz1mXSyJUhCs8II3Zw5jIy0l7oQtSM5KlNOOc8bUbgbP3+dCpguJ
BE0zb1r7DTyMV4MqQST3j90Xdjt7G/bvtV3a2fZF0CTZTqIKsrPuVnMyD6SPhad7+vEHpOqG4H3P
uUcOMzNyIkyuGjyQkMwdt/MBzEbs+7wqtE0rrVKwTtP/8EYjSzT4/nyUu+Az2hss2FaR7IWBOXSa
72XZXBncGAjxOtK4IbE54yJFPwI0omQVG+r4HEQKLgXwbEAfxNnm2G+TuCM/FZsNiT/IotU6eT5i
XPNiPTcKPqR1gxJsSqHCeASq5cGYSCwg5X+/oy+KD22ngTQO3OykwjLW4qwvX2yyPIINHonMIPDv
3eJsIvNB70AatkudkFo7i7WdmlhDuW50M2oVUM13Yy+98zyV7wp8QfxoFgJOZH616gke+/wRTyIJ
ZIjB4H097ezCQicSEhpnjrRDKD6MBKYhBkKtq0+zc+s9sDUqufQKtxt6dMC5nV/fAFXhZZxROZoO
jhOtsyRHERCvaN/ih2c1YBhs/5H9z8Nci0pALQ3dTD+xKrF1pGrm3g7k5t66d9KgJ0bsGC7RoeUZ
CbgOlZXWq7/uriiKld0SW1LVpWaDJzAnyfclzdoRFTRiSx+r/cCGvD01wNp+Hf49GcFdzWKKzFa7
eW+8WaeUGjXFyJNX0RLxoIIEp8fkRSB4Eut7PI7y2Trf9h7BvjlfMejLiTirAJLhmu76sKLgjt1M
0Pau/LeNZj0Z6CWw+RJSSHjh1KO60Y0/pffXdf4wq+GaycGQEKug0PnJonxrgm+j8v57uw4FEfbn
DLFUxkzQqqrbzhjBn1PMA05xflNU4qKTUimLXEKwHW0UWGCNMxHyrV3soe6lmIQEHzaVS825+jic
Fy1EKKEcEQVQGQshXo3M4T/tTHgDmUh4S/jSCuNyhhSDs3o50IdLEV4MusxYbvqEdJ0AOl9GQjpe
TnbOaIIZdBGxVqMWxhxHi4iNcV6Y4SQOlQl0wlK5h9AmCGrhcscAxOb5D7UIrlQML08yKCNKaMAk
OWf/JhY2sTA1WceaJRTWK0ck6R3Il7eDoglpDvR0EzmpbF0VJ882xKVDLuHyM18QdFFixTxNNJe8
zE/3Hm5dT2nl6CtXhMRr+1gTCe4wJd4r+oLDeurpOpDP7PL69jnahxkqpn6wZ8XP/cWfxzQaBqRX
QSRSoyLlHy9HWgJzazwmwM0oK8k7XAiW8F8tBOmUafmcGAHrQKV6MKd+tb8GR+6VTsQ/uiZSNVXb
UKZLgwi+cKr9Gz3KUjYrhRut65C5xN4P3xm/VHBOvM2JfNb9DL8wwyLHgjFT21uZGH28iqJ0BFKP
TlAkLgxhwSTt0wf9G23OdOuthkGc8NnRL31d+KeUDLioziGGOGtEg9KI5EyQNB6QbsrCEe+8QbL0
WaSqxhEriDqXFvPi4cytFfBcBtE5lPvEUOSOAZS+KzHMfHH40jn8J+gVis9gWc55/TwAr7tTOg0+
FHKzbzqvo/UZFCunQVouvqmPPiiRO9WJXthPRdX/1JszodZ2Cx13VWIsv1hzNzH97TdkBcywGyyz
ktiDsYmFPG/Rt5UJPoR0pABPWojHWavdNZMvy3yAVrr1Zm0pAHkVsW6eErsqCsGa1B3TIFQ6Su+Y
o8iYmZmDYVfggPmUk1p7oHbjN5DIwfaGV7WzZToxZjp312da9M/NDl15sRS0OxqIhzIfe6qF1zB+
cDTMsgUgOlIaLaHF/ffM8W8DlUruFRfLtL9XpYPFm2naaER58HwM+BETdFV39fM3AT0c75DQ6eeD
myjqR77zPXQyJCL2oYOC0czN4+6cplMnzneN699Rs6J2Z3MRickZxQQXcDx77FlIYSpOiMBWpVO1
py5LybGcw2miedSLMyzx1nJS4+qt/TZ3lGRlCgT8BfzAm8Et6n6R9L9EYv0EWsQBh9gT3xRT1g7h
k8ST4EuXCeH/bnA4kQv1oQE0Xj7ScBKk14sioe7QlcYFJ7IHpig5ht6/SoHN4hALp6EbMXrFcv31
tSYrLIWLSXyoOqjq3kxBjvSEZer4eUh5UX8eBzfIV5JgJIomEq39NimtxnxVG87/6w0lyQR+pzIx
jqMad2KCmP/719UnfV0dY3Q1u4uGHC2vlNiDF/mLpxKHiDGA2EfM5KeBKc3UG168m7gc5N3FyVPj
+2HEGfrxJm0k+rfWaOcMpjmNJXfJ6GousuFvcn78i8I3TwsWwSxRngJmA1Od0YyGgyQU65XXVuck
t2ACpa7Po2Y0fxGPGwkefXNxZLVIuoVAufEKD7rnPo+srWzuzvhdT0jp3jEjsrhRgFvwlsyTk07M
5b2FOLhdY4krQ6EPN7tzHSIJS+i0yK1VBjtKFE1srC5vIQqzdWdz+qH7YN526+C2O2iQIUx2atyy
QWdwS/GQSyNSYVIORFi7bIEE16tPe0rTclkMbY3sGvBF3pzI52HHtrHH3f3x5x/NSRUzb6mUtf1p
xUytjHkq5xgDM+x3om2UfWOvbSkl0KYn0to7TebqsvE0O5RQ+N0bm/1v8NPeLFGArgYGo9nBn0up
9FWjkyh3akbQBZhWyqMvuyMeGCfgqOpfgIFpq1Ipr3KVNvowy5ZnaeldvEh9H5qEI25uTDVoGa9T
yC2vHzPDvcBAz7kRWDTV4g9ZJEDk7XD2qtDRpp/Lwy3uePwi332Y/fwezlJR51MO2cYX88CoGB72
18mo8GjRVtQ1GF7vkMgq3p3crHtpg57T3L8E977rUk05dBQS6xCI/X5NF0lScBWLjOX+m5bIypsr
JS2Ps48FYaUPjhch8cdGUDvptDB/sMcO8bYc2p0+n80M9XBPqTlxTeSyeOpO8T9IKldGg8JNJwks
0TcQXf02sFSJOabE6aGKIuxnotjYSeyWmPGuZNbiWQpNdJJeNBZyTQMMUJt9abxbJ/F9QWSSHkbA
8ZZXD076JOp0i3poZdkgC/mQj/EURVp+qSb7pTmB6yZoZ/TIbfOyRkct1EKuXgHCfWt9dNt67C+z
DZdLr4ciP63vOG7jH2D7ZfW1mXynIHWQ5RTm4t7kTrW0nhAmmd2TU4nqr9N7TWbhZO5Rn5QZI3Jm
B7csY5tTcWlhWpM1bcIkd019AX81z2zR6N+O9QIQ3v1gh+2/QubMVkZFgm3PfzpTV67WrgNcHqeM
67Ha4TjA8opgVwe0CTITebVK9EdHOyoUUDLAwrbHYTaF4fhoJVXC8DiAXYX1n6hxxUqF6Q8KHh/P
A/6zUhx+rUSrMg4Bmj3EhhT09tTBYJL/2RtfBgE9Q7QnLYnhT51Gym5Up8b1hrdXKAWgSIeWIpm+
8t7ERYTTKF8gxbOXu028Ib0JlGX3R6jhxNuPLvnbm0rGm2yBJz/4FpD+iaIQtpHCQZwi75vl8vOP
by7B1/OcEZtnvQ9hzlwGPn8xA14whnbsvvTqiuu1LcbL0SRaEvOd0+wHjbVWm5ebhUyMYpdEmlag
2qfazKyALTBBJozRnNHGMg+nEq+jTvxDQxaC6vFPG1Pg4U3Bic/GA2PN/a3UV8CuzY3PboMBToMS
z1Zb6FWneb5rECxdIHiRNnEY/UMd2Mnc5EgBquaucefGAqNO5lskpYsOp/eppI33zzM19w5RwwVX
4T+kdC2e+PCGn+E2CPIy8TUikZ6qID0wvi0JCUA4wOBSZTvpgV+h8X+7D1RDROMH0n2TZCYl1X/+
d6hwU0FmLk06ckp24fCmnSKhSoM+EYomAOXh09D3OPnKSb1rHq6TwEujDwSg0Z8EDWpb51SdB+Cg
Jk4HVrSoMHH9aqzXis/vRyz5R+LBn5mb0d4cSZ3ZKeyG7paCzQW6qVParUgsGV0KAilY6187uUVo
ptMVWCVgdv9EQi06yFtCIRK60wLehkpQc6sYRP5H95XbAkozGVo+iVsM2sivgkAeLg5UsHrQOWHA
bwluFs/D0Lt2rqbHMe84rmBkkAx9jOhpP/kKX6HrtV8QI61jlqnsF7Ehkx+Is7FTFuEG9PatHFZq
Htn2Pfy7o/oyo5OLV4ephc5dUZ8O0G/pxtqM+itTN61IzEGsL9yc/SXq12k7Egpd/yGXcnNha16h
FHKThYTuqTZDZhSdxtV/fTck/5B+/j4keVcPDFLiPyH6Osa0USylS149h4mDHc5wplAzc3JiWyaX
AIucOhQsGnAUkMWAJJ/GAtmFLaSRrRLcFL3myZfBIta0LXrbVuoWjEIo6ox9B3j8aOaD5gqtkDlY
p3Nn6CcTBocRMlh61bgjs7x/SXNu9B+TU2Fb39Hg93MObY1xVg0v1BT36lS3e8hTAbi1TX+Z0qTW
ZskAnm9b4tjykDlgH79nxac15ozLwZiFCr383AXsg39mOfplKcg1vKaXda7e1NN8CDHnViRB0A4E
vmgn4VeeluN1HehPbzNTCVnV7jEcmF74Vn+Iz+/xE+xLKWRGS5asodC4TNIftB34oz3G1PG/a5bC
AYRtNUctXYzjUTdaFTXeb0+tx4c8maM/NPFi3D3bcR368vVAClXxmd2BLA/2gnwVXAcYXRcpyCZ2
UKCtUprpVdtRvMNcWggujNA/kZ4cG/kaPh4MbSz5TQUCxLyasRoMSh7DibZmZBIItJzxmvj/+p/n
hQ8SsssGZLJQzHEm6ow9uBo/N4c0sDOhm/viXD2PV4hWLbd6DRuREQWgkT0v6nxekQyAInVmnuFO
Nl6opFC/VBU9PuonjaksrEo5gEEjohX4UVV1vO0WboxrhbowR/3WdLQ56Jr/kH4xpmjn+MFC79CK
4m+0GtpMLEegLIUjWm1XdOKUz7WAjq9+HyRaTGKrh3CGMFat5njYVlrqoC3zPRpY02rgne/L7xBn
Nphb3JfLw3W+m+dMbakPNVKT/FjqzYx1ZHHTaATQUNcVUHf6VWhSXRS5a0iBo2MYwn6+N7YUTl+x
pBRPN5OIc133gwrslOaPGSi6QjB1gCQ2Rwn+Iul1cp5KD+pOpl7cRmejlNU+iD6JzjjERfPy8czX
2tvL+1RJgAegxtihm1oZF9hsOuD2PhW4yItbzAjojy3V6U6+OyJlVqwDwm3TGQG18U+qKPaHVvM+
PMfcWbj8V3RjiIe5/CsY+Bl54oBpqWrM286ejEmvk8zWuCdFdJokQSbe93Q079P9luFDXTLSCApZ
jB+/0fUGeOxUhLG5ZT3v00oxzA7xqg5bgwCC3oBolY9VhaqjW/EJyIdPqw1o4Ucp41bMIFigan5a
J52MBgdTl8ixtIfPh2KvS7FIiM1WzjzOLrtkBj7dF2AWTx3WkAz7hG2OWSRmkDUmnNb1I35qd/ye
TmfUWA0Lx2OsOwfvkmMs0vwDsksXwOgUJhQJkJd+QxP6QyaP7MerVs9Blmv/SW4ffXrGQ2/fdo7p
wC+KAR86Fdu7l4964/Yb8vhIrGtFYMId2JrphXBO1mUnSt2BbKzuE4pqJx1cdfkrLJezoFKIH7j2
znzG+JFJnyJNaXL7JwY4L4x6OjtVy3bJss007qowwq6qQlee4wevG2PTKARMP6JL4nP3E5ZnlJ9N
N0GkTmsmMA2zlu4WfvAFProR1mtcZQWLs9OWKVd5ZhYOkZZWyGgN+4BUvQJrF5BX02Q24qraQtBq
PA2vldzthr1R8JvqNpXyh7uglMRmz2aF7/b7IrTbvhW+zDRY02EaP/ZY72riB2hNl2eEM58eiAF2
iGqaPCY0R53BnIwStANTKNDGNo0VUvW8L83lmkNm5+An8P0WXkxRwS8EauczWIcFQBlbwmI3MrAq
cGRMa0mYgWDhMWA1vCZD+bTousgFv9tkMEc5fxmaFyIaWFunNnI/ZdmPs5wX/lPW9JaU9tvDEyuU
wYN4tKqBMRuOtBrAZwf3UUFdisUZrqED9UT8AndUkfhnSI10AAHRVApQ+1ShMH+e014O1W1PvQs1
8Ipnm1W7ES/uDnGHhhepdOifCXk0/fx70jJxvk2T/6XqxBaUWTmOTg2hopKYQC7W6fH9j5cpMDml
NNENTqViQTn/CQL4EvoGB37LiJB/BRvQuxNTaavsaQv2LzMKKXDizPCK5rUFfKB5xL9AbJmPPohF
xkYbZzRdHD/bLzGUW/c/K5s6o9Poezc7udhqdfFSdRP4r6JFVy+3rrb7R0ijydaUgBi9vV5Iy5MH
fjAs0jt1Is1ib9K0/iJtn15mM/iHLLEeyi6GMVdF4Lgt3COe/2zyHPAqYsgPkh0XkexyMm7wvFkC
vOZTbiDFyyJPLl41ll8V/3qdUilStvg3SsTF5RQtqYrQ8pb1HaNeBihGbzvcAFxQM1U7mvB6zAZK
RPVGCRbQPB1qitJLBatyMliPIdYDCLaTK5Uym667fSfUBrhGJrG7Lz+QRezhXuKQqmshKD4nUyv5
rOcWW2fK4rjpTtqfP4pUNDxEEqFkvr4LXIfE47I9vFCSrej7Wai6khwLDdN/WrDOp8/JxiNh1c9n
eoFX0qnKWCWtC+wHGJgH+XDnYVwFOWF5pjI33kCARMt1os85SpbxCcqpQkR8Pi5v3EsR7BXGZbfq
Yhdxb+7LVy347QFNf1oMrhTQSdybKXkcvWPEg4BKp+NhMjo2PTkCJL+/iee1wIVfXdnsv/s3bO5A
2+iQvg2WylBGDo/uR9fqvOCABZzKxUaA1a8gFTFAm7wBPpke9YMCrWGJNth1QgjySssAFSQWFBxt
rxM0DjbqzhH1QZoCNQdUkNn/yYGtnIxVXldyc1Dk02ix0PTsbefwRVHeXZkQzWKZprjz1RU1XDbw
GeGLc+kJgpPssSFW5LcZAlL8GW1dB2b4/4oLe8Xz3A9W6ck59RW5haKw4N9K5KOBqfpZsXmHi40U
a3s0qFKufZk6KVM+PNDB7InwvI4CHCbrXqgm/jXlwXaAqHKHJXJheYYqhUqYmfNJ4cHTjzzNL2YP
ZChxpGRDZkc1qxXJ5k1iMA6fsy3w88TlHpP2Ko0FEmmwiik2vsr4WWAFS5koztlUEcj/oBqzLusQ
C9gLdTyRJ6ZudoE/zbSPl3uzt+vL7jDJtSkr6MSK/zUqbzx4revyi0lmGX42Pbauc9TPxq3JIeI6
Q/QDl9dfTKia8uHKnilBj5odEzm5NRB8GeBIctIYspbtPgmc9KTcINlj8kScvzpCthT2fk+rh+X8
LgKz8nAZ+dLEXMoConuIpLEU82GKWUBTAz7iRMhVcNrJUFw9ZuvC/ws9ENusK+fu1b8TMdNsO//L
ZFYuiqJp6Sd+1smVa5t7VQW4MvFBowbDd8LMAL8frBcsJ9yBwONMLlEBZzng0Y9u1hJ32LJrPgDV
yiT8xfG00WST7QXSybrq7VBf/VmlkF0WSwuTT0HeiwdKUOCppXzig4q7Jh3E+y+TOSwnL3MxE3Cz
2R4Kvmy4svxKp4VhZflVxAD/htzFdNYngzMlrHFi7jAJcM67FHRi/s7we4c/IuiqqZWtgIo+RAbv
/t6hEWiROunZDoCIpDL2ZTsFwOA38iHWGbEngO585sw+GHsglQJUdVEB0Lug2ifBcAc6LtJmWsyi
z3h+nlhsUQvW8vlOG+XPIZjZE4qyOoGu2//tWevUesyNzU37XWN612y28kY+dz8s50PL26ukux7i
N4IyaDCIpfuI2hQY4WjWdgZZjwyAPQdCGOHuFk4tIxyKz5LDkf3QIJdKcUBepeDio0oSkpRwxaod
BTzcJMLlx9CLksGeuflxPRUAAHyas5tiB7ozVtWvumehkUjpUlEfpTnJQcXzltTJTxc2pwSNn/dX
plV8KeBYSe3N954e1wu8VKlTTZyLc5PBIdO0h9TpHD5lxOem1Wk56I6ITtKPYAzc3K+Xr0RV3/kN
8wROs3QN8wqFar9PrGjIZGC1CivvWK5gvtHHCSgvF87+N7tuT03aoggsnZZ+1aunOF0UdkzFDiyy
exOwPFPPPMEvWAKKdOajYDi4hCaCdYCWW3nMZ4425CYzAzumkGehggyS6E+dSLIyx1rQfLQKkwoM
kmWSrAPlDnD3pMUYEkybw2JdVT/MkqhKW/E11W6HSjwnDXqbfItwJMCscLIpvDZVKReWkFJHUEv/
tk+qkYTUfLcp6S4QmL4nWBGx3UmIrj5qK8G722bsOEDg+RIgwm/yx0jFTmuUWkggg5DAdE6VJtIY
kv+d8uAvyFop83FW4oo0kW6+3COu+h8O9yaFX+YDjaC9bEylrxpPWtcT9kA72r07krDP2FrsQJWB
n8v4qRkD62LDtjkN/dsHM/4fotuEooUo083J8UfrZkPeoCmpadV04Y/DhfRVuiPp7u+NXtoyE59J
91X0f9Jg8oCkGpIY7I2rPysiEBOSLHt1wPItcGT92Sf84zM8i/9c+YPlWMYFTrKF+CPlddDl4pPV
hejZv7JzxaH3VsU/Jxxrp0CX+px9ctI7WFnTvj9olMMyGVDsrBMftK5ZosyiLpXH3ij1rzXp1nh+
U0JHrnQ7+kcDBMnNYzasih2sv9/5K81lBqKOQkAmVMLIse/8yb8H9XYllFZLOyv13KdxsikTiP11
zSFT0PAu3RPOiFHqmxEmwLq3OnVVTX82Z0cNqZ2P12h9iZdr0fpP/LWaxis8VduCIQVZYyOZuohJ
mTTGRQlVqO5gHgySKokZ0uZWbMo0lDqMYLQ4Wn+KAfs5IEhxM7RooMKt+q0oFKtW/kJQWnVTe2XN
CYL3/visxxlO6JyW4S8QBBvKmhB/O5Jl57CPAVQmxS0tP8Sov4FVyAM2el4obOa1I6qk31cNvZZJ
QBXTNVod3O74gZ/31z53bH6jCCE7V53XXH8WDUdNm2qTBc3uOVmtppCCps805nrbUm9jh63V+o56
JKiGV+/r8jMK3LgQZ6VX/7gEv1NaZRVfq3O1SwB8wyFTH8Yj3B9c4PxBmt/ELay2iAozFluEDplq
rbJH7fWU9V9Nfdt4CkOnoCOA0fjJQgsssCDXtb4bIdopmdv+R5zNwlRQV5YxVchO/bUjxopyylYw
vOrffJ6wg6dwZkU2LG2EgtvQlXDFzU2lNnJbKDmRcIo6Zzn6wuP2V59Q2vTKv05hFviOv2AUYRJG
pPCF7/lD7CSLTJfSXOeGnXGp4lQOsV68SzI6ziKpx2pxXSc2VNvocvQRpdLYCJhwlmYKMwF0j6s3
Pokercm9sKZI3M/O6ngJN9hZfHDnDaNfn5cL0K6kWzUZcwPmgn0Y/nEV155ZwX0kxtPlMTrBA5sd
mlJZNUZcwq8L8dhtrgj52mvDtAfmyd/ieSX7AlzEP0s1sDhIdFbYlE7GXVSIzIedqoEkxhuxI3vP
LIUYXnVwmdaBPiKGSPxFrHDqL4FaD0D4a99jjz1QYSbyjw/bs9chN3Fuk8ZxUfXOtyxYpVLTmDpy
wdnyHvwgJQNXGh+UG301mp/uevystuIobQj7UehqNKU33D1pLNwnpD7By9apeJ7ucKCQTI1Z3hYP
eDeWo9bQiQgb+XxUmZ4IxUManowJbBTtEXOBF8Bt0P8m8jnel/6f9wTBsEUhhETv/1uxK0mqySX3
8DDrDa7BRWXAsGCteoBvtx2+L5nLFqssyAd1E/0vMBQCpNmdnk5KcI82BN2CWim6lCrMiTJFIPmU
nNnrW0Sz7npf/Nk6LJrfQjpGyRbmJZ4k1IN5aQx7zcsbXyraGkGcUSqLbnXjo2xTRIzPwJT7/5Wp
iAduGRno8VkyqJgIED18JDPR7gDrOb+6c2IBrWcQ85ExoYrtFRruACevsGF/Zv2IFEuot37WbSGc
G7gGG5IDhMAOrUdhGsxzqMwbS9qoObcW1bdvdbztroeqT3EjyLy8c62+d4B5/BlwmsAbjINh6ZpJ
N8O7ge6yY09xc1cxDBz/mZQzlzGKxfNN7A1nOX0fuK+o2CsGzzHR0qs7ONJAAA2486JEb+BPBhJM
N9KVc1SxXX55uvMOCJkFqorXnj7Fy8wYpeOZp4WrOqcc12xcaA7e0hUFf3Vlugrfl458VH00p+2D
DbGu6siAEPe415I+sxsfCM68uHtmaDVyN6kUCP4MXdNoLTO4vqaWE5C/+tQd2u4lK8PVKBYatqgq
EhaorFn1ocQUEBNLQ1/F6ej50IalBjLsMaQPsFwPykh4RgRgU0A9R9zRl/B0ztXvfDbhLsclVUyb
11OusaE11VJTqL6kRQlayOXh6Uid168cj25XmhFu+eadrtkPLhSM68RfwT3IE2r5SaidzOREviNP
w9JGAYYhnBMuLsd7ewG4lp/EXTjrWkS4D+YQjKC/qd3icE/FqpLzXeiERXjha/2c6PVQ3P4I2Bm1
xBLTOefmYpJY04m7/ZYE2CPIbY62BEbB97FUMC67sum3KWtdw3GguPaVqpO1A4q/Gkw6hrX/vIyK
Iiq7ZfIv6GzjHQSXuO8RGvgrk9zEmVITb1LRmt6887NupAjaWGlWO/BRwc5qlN/WY36E3Wzw+0ZZ
gJ1kZ9+eul2hEcZfR+BzkPxYln/gyLjfz6r7YJQsXPJ4HWDSgYXQuI32TmFOdlnL+etU+hvFquc4
LSIHVSvZfpNNoTraX75H1oO7kNGyNMFr+E/55tGOhAqmyYFbdyhnn5Kq1Himbqt1XkC2XBY9eusC
AUPqy0yJrVSrokQ7PcZz2CjqOWMklCcU+fMUEwo1csbOTrtKv6y3ko8jfwR44ph7YVyBlgcNwj4B
YiPHI60Mbsrip1ZwdISbipC3ERsRsf//LpgJJh139Pam+ywxcFyS06xmpivu13P3k136H5C+u63a
bZeoYNa2kQBNsgnydGQ/xbTFraFdDe/9cQs2PVbFMhtIt0OQ4hb39bggI7kWgEjM3JjJ9f4rGVTt
3qLeR8Y7aLqnHZ5Fw+5QnVzfCv4L8jTX+pu1cVB8PD5VeDKyLpByRCQ9lcT5PRkAFOpe3fll3BUG
RRupDOuZV1zZj4xqUvfwlQpZNZUc6dXtNeLmNvhEm0QNlLSdw+rZcQwKMAV0uhjopy8GkUhefgwB
VK6dboObhY7PfKbc42Zk/P0ZljCk8m9vGO0iCLeEkTFOe+ioo9/ojxVV+tDDE9MhGq9tonw2DiRV
A7aM1QBZL6IOGj0c4HIO673TlNJ7whgPQV9OoVaNF2y7NJPpqSeyYXlh/Y3Yv0ADPMRAtSEpZNfH
ADeQqaJ/t1Fboon3mGsRzBu875KpN4jqMnuX1DEZZjmyeMEZD/pnUKNBWsufQMJNkvlpZ0ySZj/w
3ulbxk4lZHxuzkdOG/1Ot4Q44hFPirCv/ljHr+b9YaYKZRDvPaeOl3OGhjyujSZqNvCz0u2yc84a
Lic4MHW2d0YBG6m64P2YUuD0qlrkTnhhsVZ3ooCZGUA6JqycyoT7lRiSHTj2+xii+8W5TBqJ0mOk
JhwvKPinoaUlIJWcNyCicZebwWnUPVaD3AETQMuFTgU0UXGtPUzUT2W8k/neTQ1R4gpSIORRHBIj
6ZMdf0FDbaY0+z3juKJyMydLCn6//BhjuRr/npjUpJLjIp+UpbxC8fE5r4+lGoteOMKR1omz+/bZ
Ag+rmjiKzYEO+rUg2mCbnnVa7dPhB/R5z2/mdwArhCGk407Hqex7ClXW2XvtNadLiczNYiCNs8xa
Ngsx5p8m6yDvOhFZZT/XIj8LwCKTcy4wv4wwEAJozzdGvJn2sbIKupJq53sHfmSdhbV660J5X1pz
Tw36aFh33yOkoz4ylif8yTAyohzGtqVdzpj50bg210cI1PEIftxIwC+lrCYPyeXVkvNo3cj+bW/3
Lm5trMdjtMR4zLexc8RF2ShmpZJlj+ybsu6WJ1XCNdvOp9k9S+zTwPaXe2od5kTo/oRUfqVJn8Rv
7K8+QzJIP82Ni04LaCnUALdSRoBbahS0uNelPViAQlob5guHO+G9Gyf+ucCYFlTlisyjp76C6l1g
Uv/X6R9rz93p51qXnCNU2B1Q9R1hRaiVgY3mFM1HHW676fymDAP/c1yQ4hQIYcc3dwD5qHPwyHph
VZRwUDSrLUijRgxxZAPaGUELezfPYh/GfB1j3kfIPZvxBer+WPKA/OJWBtgNmxxj1OKlPJJ1eCWR
o9I3lXCa2K2g9l+y4dUm/exXV1gVc+OoKLep1H8N6NGjXvDq7p2OdOyi/pnLo6FrE9uCAgGnILK7
eOoEGunIjDHEaV1Ddydxpezr9T+Be1R64sCHhoMXwXCjODPk1Xwss2hW8SFanlMix75yXh0ziQ9A
l1g6spjmZkaiIft/BvGRsOmrXY/C4Ib54GrMTx3oWnJ5y34m46oz8Ohc1dok4tt/8cHtAer1317Z
mE+DrxD68Bxa+hSPRwp8kvRmXAG8BOgRLbmxeiK9oe/sShiSGHFoX2heXnm3gMGEy0qSUSiyR9ew
RoFM18yvGjU5jmzCwhw9sYtfuW+mjUooxLDJB19xxufgaNYYiCe/mBLuXzMB9+ifG+xT05zC5eiO
YGzRMFgToDGc6e/A8KiTbO/qwS+j9G4dL1ZBKGhGAwSZ4d6QijgqoIql4E7MIWY+zYMXXyla2Un2
zmBj3hByM4t8P4kVuSp5kmO4vwE0RGga4m5OZqKU0CqZ19h1I3oANZJiDyw2Z7wllMbyCncQF+tW
tbUejUZZKcaoWXzmq7JF8iiJHMtot8zlSyTwoHUrNVIypZH2YSQlcr4U3m3IXZYzAFVYKkdhuZ9y
GHcN2XaEnivKoHeBCrnWbUxjXJ0a1FSqX4+b4Ol1LxVvM2jTtVZxKwEJSx4OPqCmn0l7W/tYyrZ6
mFgPlPj1QZqbcRtYWJU05rDZbjpQK78ieNgyBVQMne7KuXZB2MeOmT7XK3y8bXNp1t+BPoxX7pyn
iS0EEoej3kwip+zuoeqF0cDxZFobo5KyqTilwXAcmNdCwYEJjIcaKU8Mv/0dUrMHPAHoBN06S/nu
2W6cg48r8fI8CW54xlDJai6y8/mWUivLUaEn2oIkk5JVf0ZCyye8WlB5FrXHQAmGHW1UyQqPqPOp
A+cv+kDc0eQaMvdShBxEXW3caj2CRg0bhH9YN+PTHxBbIDClbeFhttFhwERxAtBVWW6OkhBQufy8
GIc81D7ERD6Ia0tTfs34n9KjJKYek5Vj9+N/SFV8A2j54+AWImZvKOj1A/BUrBFcienMkFnaQ0ZV
CgqW8GCXwUzfkAqinCEvzlCssJJH69zEtRb8eXq6LbOg/BkLPjxLIixSArrXSVikhafeau+GBuqa
Amg7fnQrNLVsEE04rgHZJ9W6c6qNqHZq14lRZRIbeVgXquz4Beyc1l5/JWZEa5cC5s/7e1xEYu+H
HfP/dp9hpBAZKRqnUWyA7ErYVgazp7vpUbvRwvr4cbOzuuieIIytsfOLXeUiKY/YUlg8TE0zl3NU
8mtWyEcKjvpWahp5I2dERxzRgDd6duC6dT7wPjbGsyML0somq8iog+ikIwB3ueljwqx7yaTmPkSz
bEOmuw/5NvbKaq7CIwhpch/+z3XaZAXkTIuUUcMzVXCnqjUqmj2TQCM/wbnTyfOIzTrfy0YukeSf
UJHSrFtbFW2zcr906jcp+OhM0dQN8oVzuocIBNEEuxJ5yaan0CnHBCsETe848QxZYZCUfYB2z4Yr
ySenuDmXE8VilwbuOhe08MZ/BuWFvMwN7SFIUto83O8h9visyuIdQyO01mY+9nE0Wl2V2S504dlW
ljpka9ceR2qQVEN45Pv6bbwUYBjHWh/M0PUl7YvDstPg+aP1XT812dx9sDpgSYA4lZZV6nrLi2mp
jONrcK4O2cpcmW4F7Lab4fn1hPUjhx3BlICM6fBfOIEazXAegf+OEzsK4EZ/fgGNpwpYWAAMrXX/
zFWzQMOpgU/PShsbi6gPWap7nUf/fI3r0q+6/UJUGAiBHoSJtKBzNmlFIoJW5SarnrJwRbry5KZB
d8gpkHZd8T3qlYBxj7uKLNd+JnSB1C7dE73mrLy3LNGXJM8CMhpTsTldyDvik/7J18n4ARmtaevN
hm1nXl9qGwDgGY0+delib7ZpefV+EnYCxUMjwW5642RPiP8DZfBuic79/fpowYbzgP8TW8G3GNKX
fjvRs1pRxnbBIBdx5PZACqhtXSyDmqiP/5xjX6Te6QzEx1tGAr+qfMO56jhmO8oCq110gB3EkVvK
eEsufiEiaXpsf4pXP5c3DF06uwhEQ+/MOWUKlPjAbAE/Svd0nZxjpMsw3MTiEXbb4FxL66EDZSLR
LYG9/pZIIIm0L618BqgivtW7eXCuLN7xMkH8VvWIb0SvejiFtd8hGOeS7sJGclAqsoblNK2USQad
jbxZ4AhsZ75zpKbS8H07nA9Xf8ss+3QNPxRSGCyCJ6nbCd720TIUHU3so0SR5zTgz0CW9h1YJV2H
f6vwKZr8ZzWG6vTZ1w0zgIHO8FTHAXybnftB6Tovp8AXYzoTA4WoMzoJkJkz6BLVP5yVIcJV/iju
av9nYsSxFX9QlZsazSbvmgwgxrPaHRKZHNprkrBUlD7eejzh/vRLQG3G+nOTfM1aMmMINgCtopLz
45uon7qPbEPBJBxFQx5jJRbof3apKrT/ixgziyDosM8s7TpDcW5RyWYqzJuIXSVUotLlj4W/MKQ/
OLyNe22d+PF/tTWGcLukHgsP+HKwLMnLcKMOrceEA9A70DV/9TThUgN5zI3H0bVT3p0X65mMfcSH
xFEqb1kvNMjwhVisTFeKk+0JBEipj6BkCqWyTfQvSAWPl3GHdMjTREY86r/Z+GanPT4GUHiBxtjp
S3GkJRn/vEBCo7VMsY1Z0SpoEhlIjOrlAft6aqfjRg6ECebXF5TRHzYNS89Irsy1ORmsNQ1oXOuw
0m4PwNiWL3O/xv0zDdmX/9Vc5NvTgYfa87Ei7hiBb8Kfsgy5shHovugRMzKJBXK3+uDpKA7/o7Lt
AXwb9yXLD4I8n9s0ppgX2HP8W3yjYUk6TurspRI0GM9F2uALyf2UnUVpFKxiXdi7VXnuvKwL77Bc
5tGdki2F35sEq+DwkJYD2oNGls0DbewCzPqFParO7I1hR5Xxt+c1jPilYlfxLH6jl6YBQbmE+vrl
Q+oDanBZhnirMgUtoJHBAv4IPB6yFji+4RfV+VS8zzm+w9sMTv95rpu+lf5oJg+gHMGhSzehu2kv
qGmAPcJo75B+1l5+3QQDYe9Te8e2BcENIJkZHVPSp77sPw4+LcxL4TxDqdAUod8d4NLl9+AMocSY
f0TeqBKn/OhWJwbYIIcYiulmped47X6nMZ1Ch/9kPS5fWk8zQk7/S6qzpKlcFZ6lRp4s+M8Zpwoy
uXmTY6KpILUx3cuMeP34h1ikeCD+CWpfnV4Sy1g+HBPKacAR4ZoBMACbwbijluJPypTVUOOR1Sr2
Y2AauVAbZXEBo8vsy+TrudXlIXdpHREQBliRgtpQGrHp9MXw+tY57l/Ivzj5rFosen9hmQNEUFOM
cycPnXhho9CmUrnzwAkbSW7icrwUD6F8dx4yceWuLAkuIL0VRyr4TeZS412u7GLu0rkpI1zZd6v8
i1SvF03LDv7qOPtwtKfHA1xA9PBlWX3dzW22+u7Hm7obFPLj1jg8dlTdHLNOmyhwKSulKOx9B5MR
le2cV4KiCQjx6KLPbrhkMJNNJt+13fuT8zHxFaH9HcTxMypykQttR+bkJ+UjsTdbHUgW+9fbsTeh
D8pHtXi71dIYV60AkQTvNgBxvPIvkYkDhdSbQf6VuLUwIjlP5nF3odqBgq0UxWetgDB4vjlgdIE/
y/HgYuiKJxVcJAn8JW9ezW4wr7nwy9LcoId2YSwU5BvmuIMls2l5iK7jF+FTT+C05ryfZ5WVhPZ5
nyiPP6Y4sRTsC18zbjSfu0k7XgUPWpRtqQAsVr2z1n2uDK9m7ZfKj4wUzV3wP9txG+TVnYYTFZZz
6t+XLX0mtqyJVGH7qnpMJIro30hZS3LRi1G8tS7hWzK5jBUiGE1JBot704dFQkEJ9iL97T73vM6s
9s9Xm6zOmxh9qohKOGnOqpBaNDMCXpJ9RopJQow4dVtMOTmeCmEzpgKBEoi4aqi1BTk3xUs8NOav
09eq3fvsZfRUeCwjTpzMStsKGpjy2JmLV4rLCR6UWg26HAI0nngnhrEh+mkZVfawMdbr9s5X4HDG
/Gt0ZTPdb7GM2httZ5iDj+OA36EW18Hc8uygEquLrBXQ1DotXcVGjVv6k15drlon/Fe3SEO/+ZFK
2o95FSPTeCmOEREQrJHozJkURU8sfZUu6u0b8am1eZjqRPLsT1nrq2teXVN2dbpcunqOUxzpS+Dj
acN6gkjPY40Wgi3E5eHokNtiLcT3B0cUULMSfkekz/Oolk2Pc7ky6MWbD2KavG6mKsC6WDmL1o0O
iXMi5FrimaccUDdwMZa1uRPgm+JSU98qf21okSYzOZ17c4XncXyQrycU0MAWcwfPApqk3y9Z0J3L
f2DhwqZN0re5ZzRDgiSWm1ZamOYBxNJP15PJI9UTxGdipDNBTRK38xUFFKRYNLJnJguFaG98Jtn6
kiEoQklPpTxbfGrBeS3vhE0Tb6cbELV/LonPzpV/6NgpSVeV6DUxxfej8xGCmUrz4euI8u8vv/Bx
7d2/pfx+ZgRl4p7elsq5WhQMrh6AUG2opIO4qRy5vha1JhfLofl0rrtZPVxz9kCUQm+8ZwsADUPC
I7CmCOI/pENQ6MppWi+VLfHJo4TpLwczLiycK4wTwUBp+s0r8yau45W3LRWi/SsVklZtWovVozX2
caWtK3LZaOjJjvLOiYgIAu687U3neEcDnkLZ5LA3o6DDJyyEcO4/4VJfDxwyRI4pu//oTQQvviBg
lGJdwDhMYzhy3WIa3slamuDTxT83RnI5S5oATtlI1ZpX4/58aANHM2yzBp3pNjjB7XyHDFV2tycR
qApQsj5DteIPvDgYNSV4pHfTtVDLFQ7ATMlYINbQeR2qtSIvvdDy80wimE98VsnN0LXboicx+vfo
+xoMrbbRrdMaEfgZqaSQddqvw7ROx4S/c2MTo7yV3ouzGbcruXcr2Ly19eJGJHsAQP6sZJEbKwkG
z0Xden6M3zKLHYEXcntVB6feRspX2R3rZJ9ZafXrEqkafo8sf6feVSvRggP5HRp8HUVjL2oVF4w+
Bk9xz64DJKLhdM96Zatob75MweEFE4m1bFUe/pPtIqFtGcTe/mrGiz7b4Da/3obXlRd/Qz0yte3o
njvH7sGn3Zi/AOMfU+NtoXn/lK5CMIOYDmG3+TWHg9W6+Il5CRF1HtO1DWrqps259nNTo0C/rfGW
Tclgd6NJS2JmksRC5rFFEhaE3PFepJ/8lQZ+824Q2yl3fwEjokZOve2I4lgCzSiZuX9YPFeMF5eE
msZEn9q1MTZBQCHJ7aeua02F5q3OzAnnGxv8t3k2pI4mh3FtWit3K2YeZFvLzp3nIhxRtOJristo
j4z9a52Xem4HXjriiL2AdGAkFv7Uw6ra6w7hxpPZMPngxm6VM6ZI1UxH+8msEywBG9qUcgod6VsX
ooEAAHm8MkUJKbsldGToEpcIwwgTE9vDbPmX9p7eZmX0a0Nihziyykrh0ljQMIXqVATAs5VsGoF1
LkEmkv2PVDEESlNmeVv4Dcrnrj1xEGKIyt98bL0ueFcvI0jdthXvb2KGO5JcL+687grplBcBoPIu
CzavcAZk3Rvy8EaOjCxBF9D4RYVhYXuuPFbsRHJaElk89kMVKuHqt0CeSgeXwWLS7YFPeqGnAMfm
t5zksDMEYMf7H3ctK8Acg1HDo/5PizffNwuM0IFJDUwQC1i2KX0rWJ+i9kW37QE2n5KIcp5KKD5y
SFwdYDAtusvcoXf+OsCyuz5kPFb6oY9KRpGmJe7rFoBmfkT5hb5wrumE73LUNndm6Gmqpq/p/Ta7
37W7X0XIPNfDqvH+G8Dzap4DreClCa+0If+xpNXB9t86QPEPWNkEvbRkOgMtItywtL/F1RPM3aOF
YMjixZyvFiFX8fL6ux/C/6B2N59ZqDOsDOREt/oVq7afcb6UKwRT4gAKWRJ9xnAXLcvKqKu5aEyG
mcXH2bBWIED/9OQHgB71VFdiv5+ONm6IEZymavKCZ1QukodWvX1u9Zp1/rhFbz8VTY471O8uluHu
v2ebsby7BG8ASxH7TYTHcQtZZCOHE06vNm5ejwWSOY3WK71ztKzk307NqYgXB4NpweECWTsKSjY7
eT7aN9OXN+1SCasSRbogsKrNm6v6uxeuzJ0rPRkHu4Q1Qw+pI4FuZdIokbCV6X3HMok139an8jXG
wtsJwRdfVo+oBW4PrCswRX2Cp1XnphMVCGxzDgzSAREaTj2YsY7Or6UJqO3jo2DOyEWnFTeppTHE
0DsLDfFxC89feOFHJbgcuiIgfY6KGkQQkDLUx+sG8U2WMlWYDTo7+X9UF6f9OmncT+wZeJ8ao1or
S9cnXr7bI6A5AduYEv09HpKF7FWGnvDjrPWLooKU5oYefIXGSYMEm6M9T5RiBuESvUr/0Meyv4y/
5K+CJu1f5MWRfuONjNZ/nMHtN7h/gBTknDLGxmhvPK1T7CRyhPqlF9EuSmH8R23Y2RQP9KCX02Df
VmUcShMgNm9XpQw+8XNA0aiJl0OEgcHdP2unUNHC2W4nxttaDG7o04PjjtzFGu6aQhzQFnlY128M
fdh4+ucY69VpZaUneMkC2dbeMtd4ozfB+4g+1nMjG7YY5MAKGc0M92Q6hP15kJHsoRW08NSivpyw
Kvd7xk+ait6NBkflsMZ5RLepLfwhLc5cCEOzLwUvM/248EAzYc6WZ4XgNlvdt7osR54WAMInEr9P
sB9o5SzwcIs3GMkVtA3OOvL+dt2X50OVSy5C1WVQH7fYYCV/ytKuzD4+J0NEFoKQNHrf5qHCQOhI
1F7HQtpwHiU0fHDVupSFC+qtrykxNDohrXPERigQ8sQKUIsMW5UZXofR2yjOh3HM+/fGly1fdsfv
azttpaFQ6ZEemQia0C+TyB8hezXeMzXwF7oIEX5t7bmVMD/0C0gmMCLzokOK4urHWlMOtGzP0fl0
RnRXyW/pBCOkXypWXY9KMIPuMWs9CHOOsRbIEp+82P+A1ZB9H5jTcKpD2EJx9VZrjYNUCFegyzk1
ibRD/wdlZGDS8xUXPeIRHNSeZPOJd4ESA5/5+1QD2Gnjqj7R5o+DCF9e+PBfne4XKgpyItxONgxF
oaKyoVlwN7rosNhoFJHmWWP1INs7MMXt+wFebrar1l8PKeFCA2VR5a/UzA5qAX6lZCIf/lcAgTSB
/fo1RVjVsPdZ9iIivQxses2wy/Q9aHKaOH6YAVEki+cNvRqEZIOHxr0PRuLIYW+m/LLgvGPvV9mh
gs2878Nng2uT9vM9hxZwrOiwQfZu7bizKGnzjlzjvswlD5tqn+JZQOXvFcsWEaeW89hOHhNgjGTC
pMCN3rw/O/1wmwYJanFV/6uvd79o6+uxTVe/YEA6olqpi4VWnyoI0WwmdBooCm9svcgOPjsXUNo0
y4emE4y1tJmzMBqcBhDe2AegXSQzjbn8T0POsC9+UBw/9li/P4HtDl9J/UMeO8Z4JwfuhItsKJ9a
qNzsRMehP7o3nznCzclSqtlfs3S2TK0HNrXji0OleooKJS+F1JSCaGLH9wrgxli8bcr1e42zwRMM
seofuZ0gIOxzChGABPCrj4zhedyVMKANfmlv4vt0o0znn1Br++szkL7wgOGXU5dfBlWfJsrOyXOM
Lq+ZNlhPfI8yWHBGnMliySQy+wATVb+UBXrTBppVn7zJ+RdBfB4WY9029sD5IA50GD5Cn/wOWznk
4jbtlbsobvZmuCfBBuJCkgI8Fie4fGD8WK01v+ygCKLFwrV+Qx29sGrxmxEG1BnTgWSE+aebeDnx
ITWHZQ0lPkuzU3FLAHJHJWCGQADH1a7Vs38TfLaNzH+MJrjTd6n67s7s5DbSClH8OTYywsylkP4u
FayfKIOn/gi7948Hcq5hV5Ws3MM9adNX+FR+jAvdjjyENbtZ/P0zQbMa9bED/BuGWWTCqUl9Ap/B
hJbq5k9KnzWWBCpvJ2w51V+zLdDBeBd+FOkpFNxaseABUq93akXJefgk+b+mc/bAQ40MxXWFZdJu
jtScRULfDXK9yyDwmripWV1sxE0Wv29PnSdzuKrYAEv+gjXLBbgq5QRgEnjcFjD5GctEiNC8ajkL
WcYGkL4S6rDSgPLifkKQQ8g7xeLbMhj433/6n8Y+i7dK035njMVTCUNCMWcTDJE6d+ckjGk5HAI9
m/12djcZsDZ1AgXsN+xoclGUY167Dzw4w3k+gil9kGGyEjjqfVLkP0hsWwukOX/hTzLT6GzUAP8V
8lXhxvIMYdg3jP3Mqc8OOeUu4D6KFFdEUQBWjWc2pnrrYWEJooTjm4qPvGMo1Vp03XIDvkxRarRI
F8YvbZ/LTWawWJCpRuklbrInXqTiJsDD3yVxtAbCxk52YeODqwoEYQfyyEfiWvpp1iuKpfsGoKCv
iuaIMyPRxREZuthdkely1vmKYOHClo+ohvxiYk/co5AaQM5yhioNYdtbtcY4uTBj+dIxQtrMvTeB
eX/JoziEhkLdeQTZPIWaocnVSDHwNNszQdFLYMiJ/V3SpKunlTP1iOK7A5fbn5cEsDrgeZ/3FSgU
ljAsx0VsYNhGMtu70vhpELAxrMRyGj60lnN7JJVMro/+6L0zGb2QAz7N85KBFb2olwb5IdS869qI
eTIZvR93ifXZltQSVd82hfjKVFVQ++m/tUp8HVCBrDZTrVWXtmG6Ly1DQxWkVhVlVjC+BLfGfHEj
6wNi6Sdvx1KKGau9gbrwPSMODZdm8+YatfxwKxCj1X3kcuEzYr/hZrbRkW7l0RNcp6+2QYjR4pzr
D7ou1s/cQVJV7QfzTKlsoS9oRhsGY0/anqCD0JzUPYb607kUUMkB/OwmBbGV6IdFbVRJzEL8P2Pt
0LqKRUw+xlXThbCPgoZHBIhbEDaHbVgOu7V2KtatldzNvMcj3INxiIo3m6MPaMqQywaR632keuCB
qil6pb5unFehP7QWA5nu71E27hBNXGYw6doKLjthKaxS8kIIFEI+D5waJVvleWL3Kuv9bz977lzm
xd6WidB70p/3z62hcPfeslvI9v1lyOAw0kdOOIgFW7N1947aFx/F8AgRLss2+ngAldZ0BzYRd3on
C304XAyGqfFM2g5dINud0lNBvxqfMEf+M64GDMX3iHLAFLJqDx3hZQiAEyDnhXMAaPh6NcrDHc3a
Rd6yZJgOBFw+WqdvRCtZ6p/MK3unzmkHcH3iPOQQo3Haebwd5gAmRz1p0zZNPQm1f/ZPVFwTPy/C
YPO4URPCcHH/hlDWW8rmSuQBH+cQup/hWW6a3/i3o45aDb6APXI6R0LkWDcaAEoGJl6dwLaqGV+K
2YzAZ8ftdZnMvtaUCQmTwCbk8LGmNOAT7T4pRH0OJFuDHj/eAGa8VzbAD3TXRJgom81C6glcFY7H
VozoZnXw/JqV4KMS4GPsWyYWQSifGv4TEp9RykYMuuGZt1Ng/DY2NCan7+l0EzltY6zmy4I3nWvo
cCM7Qt/fFRM81ke7UHf9ucTWKXGheAu+NwZG8NpGXi9HtQS/0qKnLOfv+jB16kZ+otJH1o4zWCMN
G8YlMvdy9gQ6xVwNXuoT/TIyZLX5Kbf9x58nKdLWAlnT9mjJ+IFYhrBowJibtls2N0i9+WDNpoqe
USrpIkyS8q0FiiUzq+rcUL+QB6q+i/eQAsZdKFKjBIUJ8AwhNFKtxxvmK4yYHHXGyzOc5ShtsY15
JwU1T9Hz+bWkCikdaMBbdZ1KgW/OBdP/sIeBQn+3weW2y0HpE2YLPob/z3K+TooRL5Y3Hqdo54F+
gqoJn5ip4swf8RkhiGXtvm5teS9XuuPCx2S/wyl/dP8jv2c+WKgEI8XvkCL3fS/bTamN25KkfRMl
+WboV2kUwUxsX9+rw4n8af3e5gCbA3xL257njMXOhltIaviMXsOKImUPmuewTJbCxpqkjqC07I3e
gcokEbgVzBSSD4ADpbkcTUo5zfKc16JCfhrX+MeBuAJ6CvOe/OHfZ4dE1FJiau9ytNNr6g91+1fr
mEq82TIbEcIBq9KOHlu007f2k1+QCPyQDk8T/aq3g65LRqY0WEEUktBGKpePOUsh6+wQ2ph66dDM
m2u0za8vza+ZW2PNd9Vhj7tKaiWDDI/7Dev+C1XbewDi57dAIaOKGMfKc8l7s0GDLEbUTFhHa2eq
LEtzo/VjXUhTzuaYMl9rrZ/8qNXkfb+e7XFgrSHWImQ6tnLufCfoGupGIJ0m5wHyZE6k4+UAS1dj
K5dzzp6HOlg6P2f9GdbnXv78fS9ZG4t1S81ZwaN0hVjnUaVdkFm6Af7BmYammiOoX2l6GArIAFFi
ziBxdyETg61RYOZSkgLYGCNsltbtV0t5HlKCbfWFEarQyXi09kExBnpcNhww5rRCMCffemgUxcIm
RG27ntPeNQyA0BQm9vzd7w1LG8bsUkZWf1OLwAXZihCpDY7+HUvzLPUlhNl91jQPGIjifOOD5tdr
4flUOQjMJ7S63SzSQ4tbhdSolL4StaYd5YPgOtBqdaOOdGm70p+IfVp86EKMdws7NNx9FFPLhX4t
Nr6oQg7Y1xxdicagqxY/QZODhafFryBC8v/tix9zBnzTXKmrbeE7KqEBNBF0mMtxb9fNm7QyHh0r
29L1wqsRUJU5w67Qoz2Zwi2JZ6RTlc5KSt/KNVvVVjPbH+RotKiBFdR6SzpvW/3sPAovSY4FYJxk
gc2aW0RNuU2ytp0tLs9lSpHtmXa+Ot5bj0csCrSWbT4CYlfeXdpuYKcxclr1/q+BKjOq4LolZnky
V+CNlyyXDvvQu1vgZq3tPmCULQ/o4NPtlFmEcHf+2ZXQROGZN1mnax5m0RUD1hjT/Y66abLplZsq
F9bVtZnxy7R7Z7O+ZyDk5YQgW7rjt9ByAb/5wbpvNoC9NBeBp1EQY1Bb5b8n53anxjUo59N/xTva
CSs1YdobLCBfTMH0nkQxPwYmN7fmaiBnxlT1L/ogOPMEQm+dxp9UgDuemXjow7CHylGKUAkvZ/I7
5Mac4ZHA2Kli6ktSHHk7YQUViUcZtc6gqqehgjoyYIYkddaTyEgDFDRJrPTSWCgGthqz36ddsvnf
lNuiCDCl2IHfyr4ocJHIVGUxe+s18d80AMKqbKkjHT3cEaHX+i1TbV1fO7/0IEZZsHh+y7BLhEyV
rafle5qdvQOHprY8Q7ag5A7PHx6IiohoSGgH+ErG1e/JCgFTxuQy77HbexOimz/Iv8MsU0K8WynU
Rcx44Kpu6itvOc808kCP2u4h44dBwrR6hDJJ6NI+g9Z/ic0JepyVzo0A5IMLpna26mb3DUqOenC2
wQlFHziKZFh9CGGQNI9b3kjKEuSojNwHFBHUWJOlCccGPYcZY2Y/qonXuJZPyG5OzXGEi/y2d8oA
S+yE5SXJ+Rwkqtu+0rGcTPVWOp5eIQs+ZYovZ73efjUoen825WTXfAdIxuXUaqD4SIZxp7VKF+xJ
2NvJVnNVxIGlcpKJfJkMXWWwLdX8vbSvVk3ehHVr2JhqBnaPM3ApnW7cj6zAtoUfpK9JyXh9eiKs
e5EPWGXvX1CVOpNYpvLqkh7wcfOQKbLyCRZBR25bh8+8GchuAIG/9mlmF1bZxYjCLjcfeQ93m5GM
hO8/SLHTF0Kg14unM+4jxPFRC2OYoAVf33ead9i7xrxx0GKSFWo2VYqDqOIw6FAYg/DtRQFOblPR
2IQEewwA+lSQJEhKh56UJGinyfFTOvuMWP6SLCiSZslfNv/SYJm69wAKixWsC5gctHc0NTwrMtLD
C6X/ZJ+AnInQKG9nd3nfAfOm47T6hh3+pHqWUI2IbCj4jeYPKkRA5gBE0Z6Lov6WhuTV9Ed8ZuAt
4QqG6xoKiaekSpvYnHcx+KlnOjCAHIHpmswMe2rSl0UlT1dzefWl9scpW8CrEgjL2EvMg33g2G3o
qCsOBx93llJfajRvFDFdP2J/203NL+lvBYRbYXy15nGHF0h9WxPFJE067wCCA1SS5EBDnJQqG6Ug
6fkZQK+KKug9hYUY4r80NxQprrabO07ZnmwralDOIwWfJ3P1tZlxfMrBG0tzarK52mf6fnmDnlCG
ERi1kIOo4WW8b69dKAI3bJil0Ofk75SKqrL7bi+kkLQ5eeVtAyogruwYJiRqa36lMHYaVwfeJqz0
GzJm7Q13ri3YDLq3oqsS/nQymxdv53jfZBHuQ3v2dFv+AAgGPneoFtD8Mr47u2pI6cimVj0TGZBA
OuQ/469twqdwdLhMLRI2USUUoWxVpQZcnOSLEExc/877Iae5q6a4s3q3lir2LOwF0HNzMVBmuwe9
nP/yEUBgBejH6DuTjo6iB2tMZoHAYvj5YPDPRss2TVW+oUYkJyiEazhSGPWn5BTFBR+wUCAqgvGt
ZUbXS1W7yWXa9nKbX7w1HKmm7KdUQmsWZKUBy6OK0qIqlAHtST3cBPIhCb4VrrcZTjD7fyqG1zzP
arFuu0ZSYkmsrbnPR53yzOgfrUnZyKeNyKKF9yAW0faI+qLrt5h7LusUIV7JyO85wSkW7OYEPp+K
PiA6WTkljUanW0Dshw+KM4sn9JLsqVbSzlTJnFqGvlAqggNyWzTB4PH6auS/sitTXHkL2UiI1j7h
R2+wvQz/A7Bn9u4w1MSguvsPrKj8esz31SPITONyntE6CUnXiGSUkzPhJX8M9am7SA8ZhSndGi21
2kqGAccjmyfCxnMVWiUON0RTQf0VJCENceGOhhQb/+73vGn5RzbbfJe0mb2N/P3f+Mqa9zVW877D
r1jRUVKrZr+fCiuZIBdEJPOjriur552c9jc9HHhXDWkv6hmobm6gxjPj0lckkU3wk3wwDe5SyRY0
fpYMSUog6sHMPfpDSTGVVgMV+v4mOHqoeSStxPzaErF1FJKey+f0LT31PN0rnWz1XN2okyL8FBx8
NbWcdw4ZchKHeGvP7wKPTkVeUceXbeK/9coaFVQX66ux6i1XjG9JF1BesDLeIQgt9xH5X2xO9DM3
Aw7jdmKGYBQSwxkt9R+r9PF/CYlGXS6pDr78G4e1j0W6Mff7ehcvKE+voN8bVpOGW/YyOGamR1r1
m/r2mfa0CAQNIeuLWIjQ4nLtpM0MOXbKJAA2YVk1lQvbNuKWF2O8ypsZwkOdhnkz3rxMndjYLZeU
ohZrBMB2oi/YhGpPY92JflCck2pZ5HYG+vyvokHgY/x53udm6lIxE+YLVLNcKrBVG1s2Nb1uQBKA
nGcV7E2sDBBXK/qxYLh3OiJ2+1/JCRa7mQc8ylyMtwLNCZBtX2K+lpiR3Qk72EfDnRWPlw4v8098
sXVoOyIXExqYhZGeILiX+QvjlR+0xSP2n+kVpPp0nSIiqK/HZsvCzMHrt4tJG1E2Q9hRa049LJRf
6rBFZ49SwCD9YOz1tWtHqMqai5NFcMwbseX5naTO7RKl+ZKtppKwtq/dtGcUcaCWeQOIQ9qePvWd
3MZUnfU3xmRX2poN8aRA5e8tX0brqeulmS2DZPzAzwzMBCGexrr26TAp86ZBL8S/5/ZZUttvNXjW
iOmHB/NBQ61uoScCd0DW0vxUiQXy9KULBFYrbloYSxsl3wRwfPRuax5U4Og0vrPSvKqKTnFjUq50
jIWBo9ZdKdZVApY/ycuQnId97PIHMs4VtjELqL6L6ueL+ZiDM2VIVbLaiQX2nwJ9/AH3GGFGYPjo
Tt8Z4IO1wXA06pXVSWXyOtIPPyzu9/F6bD5jAFCSIOC3TFFb6iuSkhAKSOOc9xx18j+dSMkN1R0Z
Y9A9jELOpozoRgTxZXV6xX9Sym4POnF3r7nXyAFCPgNmpyROtm7jU+/cuTk9hq1Ete0waGxADTY3
i1DM4swEC9NPLrQUJpmzuedh57AadR49FRqfjEPwfx5aaZyaZ6Xu/xRhSd3ecO2FbyrkO9VIxXtG
Yq5ZE0RQA6z57hocxDG9sOeY5j8yKzvPt8JJbdG/14UBbaOF6zO8RQFyjiONvKoJFfkhOF08Nv7R
teuxPwqnItYcck7LN6He9nHoaHPMDyg1o/kxmyEBx+VXucns9Ap5FEI0qZhrfX5p5PY5erXN1AZb
p0iNapqctL5OxgCZcRlivyTNw6NSTcJiRfD6TWqcr4nNOS/2jHyqoyYDX1Ta0pS5dwQWjIEXd60E
scsk9+TrC80Ka+F4vjmLx3LCkWqQWJSdsWkLyTnM+zFHHQSzXhU1MB3YfkMHropB3UyRRsfEc66O
dYv9JYHOzAvRrp5WlhasrSg2tdufADplVLSq8n/0pnGvIXXHbcUK1ezeZ5J0Q2gTpkFQIbSS4ZrM
/nWMKvofRinJVuGCXzz5OAWA/CLq1X3kw9QpEm+N3kPr88nsgOOlRvlfAu6BnPz9/gm6fhjZiz2x
fUxwoKD0+KAijfTi7Q5uzWw+hLlA6j+Tf5ShvFoNjVBHZ5+qWX8lA5eGzJ+Z67//lncfbLzTWZ+l
3yL+cJEussQFNsYLsPZ976gJpSAbl5+jMruz3LWLNA6Ej/CU+VbOZUFU9AlJfNZD1gUdjijFichs
pQlxLd1fPkXn0okd3IBEPvuuAXxQ6NWjmHsy4KgTIbvxrxhVVll0OFFmISEc2+9Dx1BwQN7DnTis
GYbNBcIsg/5/uXLi5sw/XWIcvF35kZTGQpWXkq3VTWQAY4Zwp4OPsUqNVGV+Xs7Qdg/XnuDTZ7V7
VvuiPG3hmEIrHCBAflTQIzWjp3cw8l4Ujw8qBALLYZU1YFE5bkWVsGL8QKYD4ugoKEfmAgLfK+GN
vGndbdU2TTf6u4Me+9ecs70g12IDvY0kvmg2t6wJUFxykp9y3lLX6MZTyGtJ873GgIqHHg7p//No
TZ/qWW40YjYvfegqxNDNTGATK3tmtmx9B9JjvLDISmopSEhUCwbk/E5NbasW0XAJiS7Ew/RLtetj
pHi5J+7/AIZsoJTRnbubHHhLFP/BDcpoHz8mGlGtOaVaOBAtmhXM7OT2C2RdYz5AIcMuof22E1Iu
BvYBQJc0xypYA3FEC/dKaH79N4u/OKfP2YhXb+uJaAXqQrtIVqfxc6Gt1voxhqcMpD8IL3Y7S6Rv
hMH1+tv1xAaYDAUf/l0hGkDFF+lHpTQNy8tD0QxXYAzVB9maDr0NyCSvc1u+s7N58NuhJGSKn/a7
uSf0iokVSPz+4UJJ+4s2YfByYNJ6SuqvlRrS57RZIJUkesw1jqrrI3poJTXio76nPoy5N0wP93XT
3jtzEgZ++2kHmmDCi8jDV+0B0A8bmC3xb9ezOp+XwY2pyOvafn5isMgwRs6J5W7I4La/dM3DLqye
d4mCYT1vYyjUUETAZ0r3IQowPPhe6kCYhpUsG7bEt28sg3NfWREeMzrBGIRQP/EDTb9fCU7vQMPv
2f35Fgk0KnX4OTuERC1nvY00Mq1zaoYxHiG9Uro0k+HT9+VureS2p/vIKBjy5j4h5nyCobn9frpM
ddQ6kKkKMue1VHpSWUQSDdmu5uz1MXfBsjUZCrm8UB4UBKQMhtW0gBuIlZwHNwpRhhIYm2mfBGoM
E/63P/kl8CdA64rjGaXjXxSYuBU8KaV7nESMIS+pX/+r3uWZCidT9WM855GFxcpNyqiklkC5MFV2
gfduT3s7gOQMkPJ8n0Rvtz7u7yT1AdrFxqCHEpIW4krINogd4Y5hfZe/r2WUAcxUEnbbqbWkZlEW
eUWLnCugeHl8Sm+dJ672ayKdqfcKcZz0Fi1xtznw+3cCc9DpUbcB+wEfiClW+JD3IghOxlaPmE2G
wWbqL9DMF4gRhFYDKGwf3asbQRxqtIj7RhMtpTtihsidBwyW0jUOX4GRksXqh9HrLL6CW15gC85k
fztk66SgLMY082G6LPR2wTQN7Xc38hjd6FeRPEz8u03gUe/XSGbCITSFa/1SORPd3YS8NpNbz+PF
fyvU1R1V6xPagUVsOL/JAORsf0IGqdqsgipu2MDLc0JCTVYV++5nHRTHxGQC/G5kvpS8c3iJ9ET3
TJHCFFMQPTU3nyDxIdoT8fnfmhrjw3tt1MuqlFpZGDx9lisAHQoXHiUYYD+FC/F1yhq7jVg+zn5o
Oem9PgoaSo8EvSQdCnyH6Bor30GoGLywAj63ks+3xbFbBfvC7FAKRfRNAaZ68sfGr8C8VHCD97jA
yb5hxuDsJx5iGQ2ddQx7o5bIa7tXF9I2fXyyIKqbGc8oLEMaEu1PA2o01BCzco5HMXMPy+tI6DFw
cG5EdSwBi8kY7BOgFYfypvrRJgfP566UGBg4f72ifwgt4wwnM4S+RZ/t5TkrJdbzo6rvzCNWQAAd
OQD/DU80TdDmSAoTp/1S1IIAcYfFd0cj/F6I06J89boUYpId9y5KCecDRO+JreYA0KOsfe1LPmCl
J6atzTnemr2ra2sq6OUAWrJ0VpOuMXM9HjKYCQd+npn2ObF7ArB1hq3CBUQ0GnXU60hTdKiQeLsX
iP/PDljmJgnSq0PQN23Nt31xmw2HYJPrA099yqq4HczoXDi+AW9tTM2ejedSks1fnMxN319Y6U1q
NCtwErZS457tZ+UEx3SFiA97B4o5EOKP8kn92p5SwV86zZRZwB1ANua1jnGvSXvA4QEVf3IZ7sip
VTvd+UJRptuth7qz+D2xkBdkk3pkr9jVOlO74df9c9BvYwDan5sipJf+6BMXYipN/Nv+Ttx2OhmG
GI2jya9VwXYYYkox0mCY25LoYNZMiOhqS9JVTvIiVQQucgKeKYVPUEJu7N8B7pbO5GTHihiMVIz7
YUlAsdqVbhyJbfM5K9yY4F8LP6JP50vS/6UsCH3O90cBoKRBH+0K5xVoXWgHipYZe/PJYm8ZscjV
nEJ2DNkUIUqotvxoJ3TyCGA4Bmvn5+bwrF05cl5+xMv/awxv7cWxN0fAtRnFbOarYvT880Q/Fbxo
dhXVGgy3G45zdPu74KJd8obEbiOpr8RxOLqypR9r8JG+E3T1rMIKtVXP+dWXqZ+7YPqn6G752SZR
YHOnUfhyqKMopDLSxKz9kYP2IhWwQxNVwYbRyI2ReT044FL0KIkt9HUX6AH13YD9EdEPUvdE9r2A
qOulAJ5sFvMfUqCqbjIgB/r+bUEzUyxu7rSr9wofvTfvihm0nHts3j8UuqfPUWac3XhO/rGjS7kd
ALQLhgayWDwSZGH86NlVkKPEcjUoA0HYpv54hKTVwS2raJ04BGtk/zfn031ImQKsM+IBH2M5pio1
2wz/l4juxXGNfu6TE7WACPyJPPGTT4uHnDTpGzJhLEnds0+v/xfjetBKZrbIrO8PEmgFW26rpMqk
NBIuUQehJtvMCa0BeYqlutJrjSHzBgr4NsLRuENaC7LYybhOmlMCx58RxUXjAEUhFvpyycA2S6Yh
AQt+l/7hR/VxIoaKJ0qTMMXhwi0T78BdGpUE//EmIdHlSW6C8PGs23z6LMnKBEgImTrHBKZe9zFs
BtsAQmn0ST6hVSmQKV+1liJjT1NTKTVyHDMz3E2k9DNql33JSLojiSqcCks74OTFlhV2L/b89rI9
jzc2qvYPfi1//Q9dZNisxb3OGZFzb53Y1sCiiZqRdptGLspGGegjaU/HhQnlvoj7ySDldFmx3Dsc
ApJOrm7q7ETkBPp/pW8aOTOT6dUaorhmkvA0jxRZBNql8AznyTvg37Xz9x7fGGoF/tal5xVGOX1u
FhWuKpBu5npuIV04CmfEHU2cA72QVy7rGxUKMBjSi7an+6b1hxJjZ6W4lUDX2ZuMfL/Mz4Ym4iyt
0mp2at8TrB9EGaHG1OfjMcV0LqyqI6vfrDQB/hXUbck6i0Gfbo/swROPGOolaThh3NcahU50Y9UH
pez/NTuBYP3Nk7spewwu+/uMLsVvyyvb5SsIIGL2gMWbN0IlXn4KJAAgZpKvtw2rnH5AKVJYphiz
04jiCEK4PEJHDa5TkyjR04xB+4lwaFRR3NKcPmgp/ubBT6hlKaSMUx1EOdLHUZeUnnHdNfPc+d9a
Hfd7MXyrxiDMe1DLQL/P/4CR1v8roMNeMB1OnG982IbQl2FMvkwC87GQU8yaqo8q6W+k5Sz1L+q4
+Xr1mqTqhZe/Mc8QqmXcZD6GO/8pqR0STM6Nq2+J4w0HvHnxOwNkiBmC8t4y5t5gePXWj50C2Hsk
LzYTzM3COfwkuq7B0cyCAhFAUGSlDPHN3LfBJXV9/gcVnMoK5ri8OtOgaX3hvEfFFpRkp7ZIr2yM
uqtb8LywHKnVlyn1ks1w0ZyxmjkJ4Yfe7u8jJhUFC2mE7hdTrY3RMzZe1O8XEbtQ3GP92BV6Z/eL
pEgxa6OfFEQ1QKUq45DVPvr5WvPwKP1572hlZGxjntHz4TB6EBvdfxRQhX6ejsaHJRNktvgNtVC+
ArRBP9DO9rjI5nAXb9YCT9r3gH8ZFlE2lVn47wzQSfiwwkveTzWTasz4Sz9vlX+34AaVQ0/MxiUt
1A6uya45Z8+TjnOWzZzoHd/nRWXTcqlaGVIhsj4RLR0yKqYdPiDo3+PjYMBqqHFZQQlkWZDuSHxf
wqxuzQyskMtrJzOVeKigdw0q/BITSjP66pEpSW09NJVPACgQ23nyp+IS+8WbMllzVOPqkKeHLp+L
h+wzg9rbzTq6jUSKdErw5jhxDM79yDBrYHGCVaAQyqtqydnQyJfalnXIKlJKsYx1Jbg4EMW2+ZnW
bTDGcbhzpIzjVUqWTMAIbOXobHZUznzKaC/eQitD5OZMMnpMQcEtooqu5JyUU5f1EmZtaC50MDkP
AGa6LeBvExmNaP1n/YB/g33xnYz9y4aBrcxuB99ILm+q4DkyqX42Ff1dQ9oseAD3FaccTvcA7uGg
US4KIcS4lB40XCszEyD4A/7OCg1ZVcfW3wpcSstuVzSHdV4HE2uBpJFBFVW9wg7K+fWKE7idHo+2
d7OgQnLyaJMlMqVl/BXNgbO0uO4/9nH83jH88Cwx/uO0CL5w66IbSYo6Dv9zv1Bj6exGLRSO6dMG
r00v91mGDYDjSiqC3IYZmA+koyDcQK1yDz+EtEny62CItyYTJ1EogPwwy8CEEicW3+pCUBj/xPsF
v9HCgRSsYFpozdZYtb8l67Vg+pTa05tGp7sfXYHWjLIeTmfwyX3zKVxYjIpU6XLLBKhSPosP+ana
NCgDSgmeYU7Ev6XQMEyYU7wXObJCI2dk8OkXmQ0bVAZH5KfD8GeNujktOhq2mB+P3uyNOudZLRCR
tKPfRPE0dVm73Tco9oJTdrl1Amw/nTCwWm+pqvAIUWB0JPpBHBtLHBacz4qciklEylZMCE2/569K
Zw3+j7sXuWbeuY9LAEzQAi2M/GS38p8hw2FWfYsvvFw5bTe8uSGNBeRoU0qP6dm1rWQDJvaY1T9K
xG+jdbuCQUCgbHPOl4Gl5uKSk/JEmwSU0yf2OWb5+Kzf2oHVbwJyfNIq5dTIP4+oh6vCGzq1Qdmk
079XnO8HLldBVfyGgqakttuk8tHcXQ+E7dqgOuMAK+C+Syo5Z72JjdrbM17IToeP248ZVeJ4nSRG
P0qjxbpbn0a1H+bN7h7WtJSGaf97qcbHQmED785SFCnhMHC+8hqzy96CMB+1LjDNdXUYenUnFqJk
etpDoWEIT19NGnX+2LjxReUYnibA3b8D8UKBxlHtZ5EDBsEmslHCrc6Y39B7RYbQyCXQ99O0QiqL
U2P+H0LWy5TYDpuKhUAw0riSQlCgInDMpSBrh8iszplXyQfjVouBSGowB11eZkZlAW0uhWiUbd9h
xlY598AuVDdsBrBx/exzYIwO5vJpQ2Rkhl3ZIlfiQAhwqmSObQunxQa+A1vpXBfNDkreZn74ki5H
bN3Em0o1ufwDI99lbAqQOHBl1OwdX93wX6O7dkcDunEAsMRk7qqwT4ScpxBbWTJNac+MThdmO4v8
f1julVYXum0QZAoUVS4SScued98BnbuSunXaJZQOVgvFwfymruZnn1v+Mnbn+Ji2zv7FeWUzBSaL
IC8+Lw/+YDL+6REvvvHPIDTGnrr7Kd1IV2arRNfQIHZqmrSRFuKzWnloSSugVqyGu80rnkramN7k
br9HyVejdLtjE/h+8/osFW2VoM/y+WbeYdue5ws2jGDXww06eyL2l3CUlRbnGInmHvNX5APlQ0y1
Umi3VrKoB+nVCW2tGS24x94/XOch15PvRDxRs+ieZvJIyOm4N2eWzdnhh3FPyifxg8Ba6vfNZugh
EXDwjTzcWRMmNgFFGaecGHujP2np4LQAfoUR+l3ZeFPqL+ATgJLMwp9e7rTcrrMdYgCzAGak0htm
5R0DDMBYMQ82YzCkDAxiSGZtksYBIjwmmudLiT64pxCCTqQp0gPaiw2OBu7w3p715LD4aF7xUhaj
ige3G0GKE+DbMz++MTB8Eihr0WGLSWQj9CvNX48Ae8yopM+vgiMvD2eFnS93YW4uuFF3OtnmMZ4U
U/LC7IPng5pmEqlApWLwJUT4gkC02jCC7jV1X6fAfW+sBGBhJfVTiiB/D/UvW3NQhaXMQSbh5gSx
CkemHftbKcPt+7PI+mGLIgOFzRQIH0FQ03aZzv05TSvGAI/PfdKv1zJPxQVluWPMaoUuGXc6L3mx
SULRW/O7B7K7qxPggR0dNWf5NV0kdaQqPpiV9m4K08w2NwODHY8/E5v0Jp4VO/nTf7MDddHRSHnq
LKP7GAmScHqw+Bv89O57spJqxxh9LscMbEb/UzOWZnH6Q+mmroFcQFlMRvaBlhqF7mtunLotT8FQ
B1D9s7DVf0t7a0XF74qM6G/ZJSKwoJBeytLNHdO+ifBLaUVWhDUHu9VyqE8M9jNBAwBGOMJy3WmY
L2BqVQO4kZYDVpn9yMqTpIMJ7ImPxZw/Mt2amtYDGwq+oVhopytAmRQKk1q8+oRjhyzDAxHj9/nO
8Ng78uiEDQdCgzEjH0WSPg+VUjTtUQmR9d2xy55C8+k0CZynC10DqzTLYqoHXxku1uR4kUN+4uIJ
yWuLM1uLt9b2f6byAIa3moyC6DWX42Z6pt00Dzu2LnZamh/DP0L/Dj7s+xEUkur54Av1x1hj3baz
2Kgsg5T6GaMPwkH4iEi2Zk5z61NTTQvsOxsAEzEFnEQwYA+W2ccIbP3JCHTnxd1hz5f9pd3zSPlV
7Woo5C5pAh+wxkCq5AXaf/mduA+PAiHVG0AvRs9FwrYERhB2R7RGUH57xoB+D6S+cPtjKMqZRZVf
veuup4mcieKv424+OUTyiPEaSSj0mxxAVfXl9L1N738lfZ2KIBsh8wf49t78D/USs6yif/vEl/4t
Ch0RmwY6Wldqj/nqE/ZTF5uKQ5mqT9msB8YBgf2UWMFCr81cPDPcUyrOyuNaM0c+3SR6UVnkrHjO
jCPXBd88dCbDqlZ0EvwXMutNMGP9Q4Qh2pQfHX9pm+sGtPyvJjYkP3x1u7MLlH+MhjlVzfjq6v2c
FRo+bvZ8GA6Imjjm95LCcYLMujFzQ6QbRqY1somUh9C/TB23+BR5FEr0UNQUByP1oGMtLDqRwB5B
66hrjq4b7WybgxW80mRFt3gK2qjuw3BuWieNOcoXQmqwWBIthXrg0jX0BsOhukOJW09+AhgFdhpe
IQv8xWmJ2ZAr0YhiZ8rxGAUSuuqZcWvo7rjuqo8l3BZwf3NK9CPr1ZRukTkDuwCQEiG5M3ENcD2Z
U/x335X5mbYvTd2Sk0wXhr64JYxertHCXcmejh6IunFNp49/1GrsvhUyvAhAeKQW+CZ91bJz+xdR
Hm0cbIC3g2wKTqL1c48Ni6EMABnmS0ENY3EsX3/L2IQS/8Sv5dIlr4lMWaRRzUPSQE7YXHsy8zJC
hnVjTXvC0zILqGMCjpd4KZL31pr6/lDOLNJQMn3g2K/aAXTcXCe00u8H3B+968YPOs44fi5n2Eog
n8XTS3ItiR6KC1IfRsOkYd53LNBESI6r76etOBudNjqExvL2Vxdc0Ji1WzxUnk6Yv6n4gHpkletN
/Y4BWSOl+AlNV44h5Nj8CQEu4jvEvxU0rih5k/RRy97dgsz244821MPDBFER4wRAyVZT0ftBT763
x9NL7R7WHVoNh+q4Opag57Sfd6TFvB+d8Bpp1SHCzjoSr98bT6nwrn6UkqoeUSOW1btP+Va5cH+8
+zc+lv19BPKQpwUzT+5mm8/e/AuBkJE2Hf6a+VdOUdY4xBgBQlz/C2q9+Mk7kGuH2SjQ/FKypImK
SLAuFDnlC4BMg3y4CJsQ3cTmLZKxGyfpbyDEvA05ouX5eK69TRvhOAFYU0p6Ej2fOlYTn4C1sj8i
X1aNojcX7uCnA40QxOmNi1GdGUCbfeaXjxCPu128JuktiI78w1zZF+tc8ejPrmOqT2GbDIS7heND
rg2kyca5UtBROkEttMIMVjVSQqdegiEkCpn4bgpqLerjfYS0eadLrZgWKT48glGhb9lOMOmBfG8Y
Tj5NKWA2VS559maxTSI9PgwbvRkO0Yo10ZeHTR0xLfGl9OMRAus1iN6JrYzw5XMxc7Z6bMrsGb+X
Z7ZyoRIzPJkSGVjbvK5vpDryRVq5PD44VBq89kGSDZ4eS/KPwEdY8gbXKvVY/lujsYKamwOaM4o4
6igrDgo7xotIC+ou5nGZpcJnpAsjTWSbcU1C5Bp1AT1TsnQEFjYovRYBS+gs+q+3hGBPf1QzUx1W
wwQj2dRKZnWy3AteTu9FcntprFro+mAy37KE5gGlQ6Bbn2W6CPkYco9UE7nkWF3cqEZx5rO5r97X
snozBLEe3mfX7ndGMGtcbhArF+YTPeFEliGzICJ1HhtKLtv+B3wxof/VndPZ/e/JURWECa5xt9ul
LdwJawL7FSVwJBHtAC3SKIaFiOt/09xy6LHYpFoGXzGAgQG2KHzQ+kdj6K/UCPMcicWKVeMwxGgX
+9JL4yUDHozkxuLHga3YgLQnu7BMTfdy53Sd2qWLEgQ7jhUNP1JljwW2I8MRnaQj/WvhHNoMQV1R
0dinlrETcQUOVYBC5zmfeqlEwxhtVhHZ+lfGjYEwyK0EG42wov93iSSd0wXbNuw+vEnnG1uUe3qR
tsj/CgRydl6RehL07LfPO+nlKhZ6ZONaE3Cv5obBZ8a/g/Uj0DPP9g7Lm5MWVH4IQlUoOhFHsyh1
DUTmVvmNsLwoXbbxBLgQKGcY4H0GYfdeA0oe0HW2ccL4QytqkBPvMxHnQ8SExyH+6Ah77WSnDWGU
4rYAtFPrakAc1NefLhFaCUUnfjjELhSTKmn9am3c/Yuy/AWcfYkAiXTCVynlRa6WUVpzJbGUWAIf
qbdn0/YCjOWNKSPOkdgaDTzMzcF1HtB5Q4oE6Wp6BFBchgpOIXO1csLGIvBh55aeg/43RxVSBZjY
9kQDZjFK0RfDtevm5WPT3qu0PvWAJqFLP8iDesKmvitw12AjA1k3jbwH+hj30iA2sVpQohghKE0d
deKbcLKg9mbEiFWel9zBgSW/7Vgl3XcujPZqMkIrihtxfLiRrpWr83eV/kEgj6Zp85UliYHPwwg3
2qoir5+ESQl5yz0qAci2F5Qonqj1172r7OM3Pr/DHfvnK494msnJExIfZXqghM2WeQ3I9rsekvrk
lYgajTqWCz4+9am5XodPd1xvNyvHxVYXop8Nph6XbPbbTu5L2shoOsIiRqLeZ3vVGddoWl16kTsC
lVh0ZrUc3pSOz5uwDqbuyaFS55wHEgWNyuKgmLxrEeT08++G3KOt4kduoW4basAh2DNb+z2vVXzS
SdAc/QhFGuyioIt4wmtQxIO91LnTpO80yW73tkNsEIp4uDmaXBo3OJlfAFQnnvUK66x9YOLRYV/i
HcZYgdRCS2azk0zoBri5IHCVUVHAmxXq+TAXtP4yEQnTTgRNMEFbm60tCR7XRq6BCMNQsTigEGX4
saH1505rCkZEnArpNWMApoW7v7I7dbUl/FSYrI1vpMEoCjW+sVjVSUBkgLDZ+tE25zLbLrz1D6QD
ZCU476KHiXzyJ87W3BJvWRb6kYP9CAYizlrPj3OS2kSp5i9YGif9eqllv4qbeG/62xoMoWyw67d2
y7sswLlXxry5eroYQjkpAXNWMDb1V13E4IgPpeuIAoyvVdZjsGsTfkHjPTq4YEn+8bQ6wDfY+EVM
x0SD+i2pjGME259b8nnMBmMozbQ6Jh/o4ZmREKJzbstA3ztSBYWxC0MEef7hj+BzsfM0JdAoV//r
3UrhLVwj+J9XISQ1Pl4YqzTDe7mTtgFbIyfk8JNDLwFKIV1TMqY4s9tTpLqQJnMsewX1EfbUsVpQ
rQAo2wxLADd0KhH4fvuzeddLvm2+hl/UWmN3f3K31OIgtlJC1LD/MaN9TEWJrMSLfC71h0QRikgf
Cwu3PNq3WW577wPuiOqOjzwn3cz2hjPcUetlcsp2VSI4z1vMTX45jBo4TUrznlikZozm/2dSh6cc
ut6SoxgwcHGQa857at39FLmEw6W9/fUoEN4mRrKWFB4XvJr8GuLX6ub7LIWm6lHPmkibBdMM5K0W
TcHZ9hRnrcrzvRBnHI6e9Ki4iN8WJ4C5eQbPO9Q1Gi5YWhAyzyPzNzuzyJtUOvXiICbLz1VuLXk9
tNc+eB5BfTpfhviZAQbMmYem7255F3lhRN5tN6OeioXI9BDAxA0IPJtgF48Q/OqkaAaPde1/t2iX
kSGQjdG1hn/I18o73t7zsmkQJ0u+P5kWkrU3twk4eWWUGmVC48UhmCwQuskr3Ztar5CoVDiyBNIB
pDKZre0zPohzOPLeTPJLKEkFz3hZVShJTKKJq9AAf7L+YAnq5u+r06xl8bZSo3dL7pd3AYO742Qc
8fvXqHHsKluwrcxkBiU/o/Bf1FY0TvIi/iupxHgkWIK+42n7YHChrwokQ+yR+ZPpOH09G2GEBhI3
qqZd31srR8lXea8LeX+GikgSF5KUWFG28WEtbSNNdtqSs6Fuv7vLwLslzC88mscxTtBs/GGR1KHg
PwOrH8yb8tcRTVTN+YEQKMEsK+QyoskMJzOi23JV+vsAeglUvVSz4HZwWDu/mn8aS+Qhtn+9raJx
ZSQ5Fn7CjOIFaFyo4yXg8c9NplGmvQ6nW5bbcoSat31QEBj8rX6sBdTRVbu501HwxjwPqpDWQs8B
ZS66lyTOGMTVo5dXGpphlEKJlsVxkA7vDMS/PpUrLJGRIp1fg/PzhomlpuEtmBQsxT9FEpIZVR0u
LKw7cs3uqs1anr8MOrYjqTu6tRoI4+wL+q5MINUYoEjOcTw0LudJpqvSs6KpWfj1AuFuO/+PwXVt
FPGHZ2Fxpd8phferZDUXgOOp8u0aEehM9FDbxa8EcEhGIPqPn7g7/furHonOXDR2YB1mzdYubXZW
73IVAGvB0gJw6+FuBjN2B7VucLEijvKkObcppLgxOLH5cmVuJFTJJqZ1hMIMq3o/FPVgq0A90lPD
3f06zHmslIerOnabJtml8f6u9k4hJaMpMlrMhWD5fI57I9vFL4upPs/w952OtAfJzi63ud2hK8gD
fGTLOQaljrDStdavnjGbY/kwr08UEiY4NL0Pcisrb8vhvhdvydtGekkNz05l69i6eUlA78hsJkuz
KDimwl20rQrxA0N+hkgNiHmtvCZNsMY4QNWeNynn/CxH+f/72ZhMHtVOh1u7gpLHIAkG7zkRxdMv
LXWtC8datOVtobQtxsih5AYKGe379Hpja8sG8lcp567Y+7Z8gG9TuSjPJEnkSJPYQSrm6rM51yAO
LcuDuKAQM2e6oXLPjruU+x0BF8w8RaX4tV29Pvz0G5TL3I7gYFgHD7Wg/N/sSDWGcXXHpsP7Q3ZF
Oy8af7P24TeGMSGwEZKZs4E52Km2ItzkBqa0TWjJZSzTc/s2RMBhcP93ggnnZ5w9UBOtgXb17+uv
Hfw+/e1nmIE6kj+4B9mmPPx89vrVz2xlJJYQwdt6GXcKd/ifd9P0nTQ2qYMGrJOVufb0+d3aQ3Nv
2F2oGvIVaxMY7LXja+5SVkMbMk+QPiAGDC/ZAfa/v/K56kuXU7DxR0KN0DKfDaMpfD9YBkVo86aN
9eqAF5ub/K6RigJ1LxmrAnkioA57BZPtE56RExjg6VJ4jujc1e0EecqlfdFj9+AdqW2jQuV4XMUx
F2y6apmtlgSRu3j3n//07aDDE58GOgXMqSDuVaYZ0+gcVNkIFp2SIOlrRr/Hf7LomPf2M+YHMWas
TAYTRj0ajdAOwr/V8DnCKO5SDy8yb4mosAtlVlkuBgss6VJfL9IsRQUbPMNYvGNh/OUoZJxDDkOf
R1aTr31bcYmLChufEu3nzOvZPu2rd0d79HqR8RPAmWmoYl+DqIxp5S8hyR0I6oLRoJpaD72o9KMv
kg4D6dtRhhlmOqu7DyifJomAUO5BCio9poOUaBQ5L3IaG50xHJpKnBX80rbNbOvyGQps4TaGisum
321hbRdKBfkobVLujxMDEezTcOL4es/05WlvaNGQ+jpKpSCw+kZjo7RMSw3r13MDMem3cUiaAzwk
fy/Cq59pE4u+rGOkbaCUK0MEJBa4aj1fsZ38ljfqqyQPXHjHXfpNhx1o/BASCFoqGLjWWcrVPdU4
shXUJ2UM9hK5o1Xz0Kpq1klCAPcihmgX0+W5Or7lShbXfYAYWYBCMim5ldBn5qCEHYa9Vws7CsUd
HK9XzsA98Zurf6F0BFxudUoZAKfnuyaavhpzXIDCTp3Kfws2Jp5JXgr+Zfui9DoHo9h0Sa4rySbM
o7CXbfF1VB6wCpGvK4Y98Alo6y5GxObzamNhNOZDt5G1uWjyJwtn+uDfcGN5s5aNeQhhCDCTfKtI
vr+Oxu7nITg06ve/DkQ2iGU6cCKdoNYmHc5/TZPJUd+LwHM3493JvSG0sLQ/aKREsiupzJpoejen
79vorFTRy6ole1+pdVsA2EjprXQRlRx+2Ud/hpn2RZx5gwwCtxbrXy30OWXr6eTosnNzedT08w9t
02LDAEykG0lThCxWsJrPEhfgEhah6uBbbR9ArqBpDHelTEudxe2vTD1OHZLmc7bRBsdZU3qzFXiu
291POuEqumFDx1gs9Ll8ITHPfTHzGDSGB/hAwyR/+NFnYLe+qQ0Wxk5CgcnOwVkFWq806BTYCy1m
o10fJZSeioUn0Ops8ZUaYO0zn0mx24VM8Pk2TsrF5i4Js/qQ/LYnGx6tLqdxAh0rntms3WypdMlB
PiNX/IsqyTTRvdqhsZoWOuP7udURaExrRErVRuLSP4tthgA2XQvou+rEam4AxJZB/I07seOlJDhL
+XXPsmfXvQxGAijQlksrwH8Ejtn0sUUsdGudaM58GzdjdT9haXghXYk43PWBDR0DaO/H1jRzNIR+
DdLiIXgZYGXx+tJ8Gsz6UDDxwMCfl4e006ahIgXK8/kmOJIsuenjqlE6dLxHYJprstgD9ImkgkTs
jpbsuRTBMOpNDb2MVB0L5JIAwwD2zOslc1l3tbr23DpdO6rdzNe6wRm7WEdZf01G6Q+ju6BONZSE
nnpEdp7I9/7BgUAWej8QESZIiBLg4qf2d0IkTNmvGJSDG7HWarvZyqz7UHse14K0uM4dmoq1MXJv
dURchCTUgvW5n9i52h5HTv4AA1RuCRlEUosxI449Sk9YoLNwxboLlLMWjVggNulvMQx3vufFephM
gl2/YbmwDGrKLgCImVDDKtaG2Eue/WQS+1yJ7992M8aTI+P6Exy1+J1N2hiN/SHbL6Gobgc+KJrp
k/y5tcZobXL1bTmpNSN9s2PB8Y2yIn3gFnjTgDJJ35UKXvUH8m4/xnPEm5t4ZvDZ7PK9+LCOHBmF
5tAKnk4SaL7xveK8Wp45o8xUYkcTX1f2XUPNFzn1OezeT59M88dPTUvoKwgHG59a7IcO3nKtVH9E
QaV3Tj8sea3jPJ0vHBHkUZ11uL2kNRm69CIgmQX2Tgpc8MeZgkYcjbTD/nP21OsnoWkZEdvJ+mFb
okXiBcegDoMDAVRfH1IwcOLmujJZXgXXoJVi+/+viZozD38uUy1h3iaAeGy7z/UwKxiHyczlDpDu
A6ZO/vUsfuuHgtE53xA/EtlbgMS7NkF53+nw52VSkvA5feErpIbCqrGZsWD3UCpN+OG3dzT6TNyP
idwk7GFTPTKWoVVo6l0XHXN4cKvuI1cXH7uvZfDsyeNDXC9zbqZfFzk/VpahQKS4qI5I/kTFPyG9
xTiCHLYKmkjOJlED7WvhbEBRhayz0fwPQZ67wJMv88r16+EigxVwmkH3OsRE55qRdR3rGuvL6M7q
hoVqmncd/H7sFBQmv/oU8ndakPfJRTWzfhPSss8r4XST5J2AtqSJyfFw8CHkITSPBAkrUfoyU7YT
r28+tfdFCUvkhtLx7Dwf1vpTR+6MtY890ERKbEdZbmS8muKPLWDNjeifzRAfnJSgD3riPEdZUdND
Fet7k1tDkklvX22Rc83J86St9NY3CvgSlu5zS6mRFuP07Tf9l1KiiECbkpYSWPFL0xUw9H7mJ1qJ
0bpXFlWFacB5jE4tfyiTjkdQ8EQGj+mUe5MQfvmEiJMw2FMmgppmc4yijiLgIWGDcg0e3BdrBZIH
pPz0x14ntW3gNaWQ1yM6eFnlUSRcX/GvfnUad59aO6VYGFWv05yqVhjJSmOZFAOdtxhfo57wkm2L
P+FMxgZ+tpsS7QUZbdtJRkdBPtB2eY6aa/Yg9yMxHuvqbGdqrjq+H7Vj11ztcBZRBhui2Crv4Wur
ekyM+3Ong2tomiuIGR0Ifupbi1D1L3570/gQW7WXH9hR8ldGBNCsr7gGp56QfgJiupoYSiYEj7w8
//9gUrhxfFwfm3KJ9MyUdMV/1wkdLv3mNl+A9XuxB5QpFI0fvnXU8tRYpiRe0UPspDI2Wqd5xfhw
FWK2xtO1lAbkoquBIJInf5WVIqMd3XXgq/cpqA5TiseoZKJ/0OTZda5ALq30nZiboGbk/zqdwlC4
YM/KijLDanCyvXtjZmJbYjGgEhodxvneeOU0OtdCjPY6LEjbpf0WRz9wjJJhNq8ILZ8tOT/d7rdw
9fEMk0GpFZ0MSVGnP/VXwpDPfmlzMokX4xuIS78WGszA38sJQt0IqvnZ/6ytz1kET4ZAN2cJIgZn
ARVhYX3pPcqjzlkPPmxciX4EgTJDiteEcTJhl1f0yY06qMleu8p16zIrQa+qJczTWb9QeT5kb0fZ
Dw6Qr25n3pOPQY3ue5f0md1ssgy7zfZyl88+7+L1Gx7Mfj7oVE00genbsKLs0AbEIQFp6h9zaiaX
AiigZHngZ6p5NGT9rexP1NdGLEB/LqN/VaGqv9Md3oiUyFoOa4GMwJFiHDqYMnnZOwMqYJH3bDwP
vFpMCMSoouucA0szZXdJxD5DZEkBLJgFWpYpIPoXhHdzgsU6tIHGdsOUVsgHcf2pv1l1QmyGV6fD
z5zk5+YIdq0KElQXbsfD7h9TrNJXB6fK9h2NtiNHRZ7weodxfZxWOHHDP75QgAPioAe4p0UH0bHd
pobGrI6moRi3Px8r35cKWyqweuLXPIXnMNk5/dEglX71T2tqiBnx8iM7GJQM7A1TumnNzlSVCa1g
fsgV2vBrfUdUAlMfqfNMal66mMk9V1rrFLL0I6shm49fCe0jXqmtv1fsA4oVFHlTSJSSK2HLfe95
458glHboubiurOMrpkVh8nkC1yZOnepy3k5kOdW5t9wk4Vam7hnkh+Ht+5I1H91hlnf6OV23c/rl
aqJzAfIxd8ivv4wFLRl25SdorpAnBK1UZu85usDC260mlHwPhzgKtCGv+zDsB9/qk/mW6gOCMZLG
WM7g5Tx0L5JhjPmOr0uKXCoFuICcwwtArigCc032a6sTBvbyFw1u01q+iDhUC3v42uiQRtE3LVtJ
3wuoP2ctaq6mlys6LxtOh8+qLgP7Zfj+JjpzlC9khkpeXfTlvoDR8MWyzovlXHOpYmztoxHy0vga
pLjQSrKyInZR+prOeHx8PRSaX5ORTW4MTpStkgdMQrkA4ciJ44oEMce/5snLuY/304iSKOTn+uUZ
xhL4AJHh5zgqiHgV0KFNSPAObNwuWmkeQGsdGc/UCpQLVwRATErniHpJrQVayRZ/Nsc1a3hUZOAP
dyqMeETR5W4Ni0nY5uXiRdHgNYH6Yt675suKvMyK1CuzQuuFICJUWbcn8DfyK+YQZ0UcSGmGHOeC
DF4TGnREcPJ5xxbe/SuWi2G0VP0uX/aQUxM0pztKrDjY8uxvbfH4S43BuRMCsTX35tJsDPBIbiKQ
sB8Tj5jw0ThVQf/JUh0hXs9nrMyTKkuv8r3GRJBbi7fZmmwYXu0kS7CXgZan+fDRnduoX27AJDuz
jKMrlJa/FIFxSVT/XZOh2zHobr05FP2ox7JRN0RevkF1CR9CnEToJll7gRCJz4hrz/0CVbak+kfk
dSqKdz3owvq34NNAdDH8ErYYoE+lsFGlKMoUW8XAYxHZFzWa14nP30jBURBDqYW+3fekUygvm72c
vylvoy9MKeexxC0ZCExwlDMIP1p1CjqiEGjLIQWYOuUikUjsAkZzLOVCpwnqaGY09HP7fX5hs+aL
mlmyZDZSy/kp+mUgTYHOtPy/QQ3I4Nkv02OlY1UTqYs8k7NCZHCPukHfQyJD6nNW/fO0mEu0TPA6
fiLumkJxjBCKKfEv4Uo4tfFd5ZAzhcJg5ESocAseymmiR2xiBGewLC9fLaauviF7rjP0jOxX1XtS
F3lLwsyr7KeYjajNA2n2rbet/PrBaKgEi8u/9MKqugNQjs2a2a2jz9n7UlWROFHo4EvdhE8G4J63
aHPPbAy8SCCJrh4shTAi6ljHWx769UR4EMxTHPCF2fdEerNwkvUuh2Nw1U0sJEdx4/I+GrDCHnf1
ZYFQ58Eb2d5FrTqNkQhynwpI3Dzj6UKjN90ZTlKAJvnTxLoFbiWGSxqEC0VbqHqcO2TWpfsRwEYM
ywBFf6T1CKcz05chyZ3z2MqEFJ/335hFsz4Wt8dq/V0YNk+nAWaekUpfw+vnvGF0OipJmi2kcUNf
XDY6FoUdkR2Krv0dWCx5l+hAYN6XnJzWVMC/XNMrLVwdhVOGBzMJ0NZGcCHbjy9WlH7B9qwGq99Q
pWW1lDaI/oob35FgbtID38A/UhGKsSfwk61W27wxf6zuNZDuzyLHCwgDlDmzF1ZDNPwSG4PmKYEh
OVZ5COR2+QFZ/M3dnxZuu/HhWLcStLzlo4Yi5EnYdPimlvpyI1VA5MhAp4Rgvn83q6abpsOVpaeO
N/QM7V16KtyXrAWEBAaOmQMUPCvlf1tLNpHZ6lXMifeBBatufpGD2vap5Hc8zFWidWMhfpxDyiIc
L6vFaXzOei2iLuTOF8cIFtJWsNEhS3HVj0BzR3v87oGEKPmIOeGnu9qgjPKn4i88UwJXugUuqC4b
VpIt6Sv1HkuSARWT4S3UgxVdxUW2PDLdoITZS7jNQ9M0qgWwWtYSzMq4T7ETjmd3/xubp+5L5ZRe
SOU9z4j4Zyr5PYPK2i/5YWuhBx9WW1do9cPbj7ed7Rh+LOIpdVNb/ThmMROmeC53tWaOz20zNa2u
rxZa2UAWtzO7fj5Yv6ENdfqRSM/MwX4RK7BnMIaLxSfLXb1MQw7v7MrpLXEtxltA3FbfE3n1ltb0
tyK1/gl1nNsVx/eiNNWre2dAl+ygPxPmuvux/vVM4zLFczDOt5HKLaR1MV7S5niK3si2hDhst9Hx
sV3nu7LHix3NflWwilG9RzzY9T33HlBcZPuRcZrJF8GvFMYI0keQs08Z7UWNa5OdULUTt6JE5srX
9tMmkTGBMBHvnNe8KUgdXXT7h/zbPFO5ql3UoB/6br90b5fexIPYbCPZ4HKeWrD0kV+C4ZdH9UL/
8Wj7KgKaYFbymFvQ4YIDWLdpjfr8iq3GTFF3hsP+FqU0AAb9f++EmOCLCy1qclNXOaTB60EbqCIa
KR/Av2SIeo+CvBjUiQGylJklM0yY9aSaWyuiM77ETmRuYNTLi1o9znHstPTzzPBbH9bX0Ndf2i4z
Fbpv/V1zuhoi+fozmgdOo8YsCt/92qv3Wf2r5Pbj/P+39o1minPVTfWnSl6cmqGFxwIxhBXri7SG
pER+1PtqXKMUqRS9mihit9vKWKJec/WKERKo6CryfTghZw/0Cbd0vbIufKFcp2KrYvA5ybj5tUzh
lEauTMKRRIg/1Ra/jBzchPT+gCpj5Waz0BuKSFoHe02yYxDGMQNP+e06jjRDKud6pzYzAzE1Wt2J
98fLUOsbMgqEPSzbtGODGmXDEsTAyWtwwN/n+njaIVOgkm0rSrMOYlJi0E1ouVLvq6aXmVpXluGB
k23y2z/u//hyiKwAj0i1TO6cBjjWQjXV1s+xRRKItN3Rx/CHfx6gHiNvQNW9YZdatji4OM1FPr6z
a9erQR5PG/qKkRQgyYdIRzaf2Sj9auFpCa8L2zIWb/i7OSiD3biufgxDCnhdnHmWi/6iDwaIqPWn
3lOkQeZezIRDoQ2CMaN9BYNaC0WPbArPp5BH6dHBvTYboy/pNJq/9HX/G0oHSUJhIIcobCUVrd3h
ILSEnkAT2Nrr+dGtvI0zxLCRIsThVvnlX8578xKmhFdsfmKoYRVPEoo468vyr8+FNl2QAKOTi4gD
kxH9Ux6DU8z2JmRwRxfr4i2KRU6I4Gm6WdRj4zmG5Tqrtl/9IF5LIQkql7eY65jS8YqV7qCZTlQq
Z+G6lIx1tw4jwvsLULDu6a0OzhnylhVWuD5YkASuhwQ2RiA8NpswTn+jJFFI5pGGMv4VLm43TNzu
VgWQCedBaz4M5CsGzW0rLyydGXUKDrALdqTk6rnkpnohSEwZDbUA4wUPmfZM+sERierFXw+E5hYw
zHtYyetYiUpNjA80QbYE0g3LatYFMym2RT1gGnHtT/tr6/+Txf72ibMm5DJ0nOXNI5rVv3x16L+z
zeb4rgKOoh/GJXdL63aq1XV/MkrWvVSuZUU9B871K/l4JVjp0fMk+2UErM+rtm0mBEuwSbqr6Dnp
jmEHTmtCbtenKpWzb72CRFnBjkYQlZGSTqlDjk3TO8bL14LqmwnqWTE3BVDzwLclI+pX2CgtODvY
xUKgu8uMTskuS1bdvLuw1q8RR/2LWbFTgeLOJcVGXFhh21UFfJ7zfumGfO5H8bbhY3oSWrgI5XbL
XRCKiCq2I/0ofEGXb4plXlTWinOrNaTPB145S8GiOh76Fcs1IJUAn+ZxulBoO0eSTGFaEZttwRhR
GxiXW1Qe1WJCmluneT5WXyw15ExDnP0u+1aJWUVcyVjiqln7IT7NbUB3FlVuPS8boaJZg+sVcxfp
ZCUrhgsAyfSDe6lfniA6VFxx0MDh+n5T+9JV0tAXMOHopMraZGRjwtvFAAS+Qun8+hhCvz1erXBK
gOvmuRWgl+IiN7dTRDaehCNAMcMRg3722a4U3kjaSPKvOMrx86rYiYJfKuScGEH41YXJR+0cVGvj
3p2y6/4j2Lo8LGhkIQUgEseDtSyowZPkyz8BR3LCB3creZiYKW8X/DpSG0pS1nE9y4qp3mIJH2to
Bkzs5X6ikozzYKvW5qBofnAb2UOOTk2vJ3WlJ8PSP8sN8C6suitw//V2E/b3rP2S6bmVeZp3fbdS
l++iFMc23jJrXCJ+E9BRqSSdCJYXMWSQLgDNH3+RCN23+DuqUpwmlbgjRbg2rw77PXw5KDzNJkZH
8igqtcDY9e173qYqdE86DytB4ghiXOXrMLF541ZE7ALyJbFRMyRLxRGa1t0cAg251kUQVwM202GK
uBO9NhRESPZi45OnDEgOTIk53xPSvN4LkaiX9DuBw3QdwJDBCrmHfMTm3k7TU9GAAQve4K80hija
MkkJJiJOFngVoxRYesRUd6CeO5QRab8ePoNQU0+pEqHhM6XtSZd+U8TFc2+/6RyN71a9G+PdPr3A
eqZ3ZQX2Nhv9pbaa0WAnSnnuiLSy8pHSSM5xweH48WOPi/Hgon9ru4OcGmijtg8WwxHXYH1MgQp1
nQJOgy72khAJTse/6Jtl6UbWuoycxgzqBNkOmnLSoddPxJ/Vctog3UIxu4Bl9sIYAnwevB2RfQiA
tU9v1tO74mAbO1ywJLsGNWKjA2ee6Gm9XZ8fVOrzsRoeixjZfaOJFL+pMP8Q3v2+GM3EsZSZaDyg
+3wy2crhoglImhwoHwccAWnAWcHkdSbzZGsBALDiLiFKUn3ntVJ7DnUwAGquxTzdFsbwDRxMWLxd
wUodIUBpW/Ox/l1a7pg5K7WkHXOFl9D2mF/v+dcaNxBt+XCENFnlBGT9xX8fi02myCM4em0HZgUE
vMvRgrt6Hshm1k8vY8OE00gPF8Caz9Mu6nwaJb3O1NJ/PnPctdKXgCLReIooRqOGojLUOQt1Rie1
0Pjo4rNECm32lAkrXlRv4tfYsTa9WI9UdB+VwTkmtvxHrk7Tr99tomo929u7IIrDS/7jN6BkNHzU
PuxS+8C4snBLYHAeBThTLs4D5doioPharNnXoEnxbWhw7DUGK7nOd45cG7HDk5jWK/LKfYO5W7jB
ArxQLak91x1btfvtDSClUXFRIm1V95dBD2RQy9PgOdItiQ+l6UVi7QHZVONaekEM/Vz8Qc+tC1oc
aaMkR1x0fO3512AfjE/qSOlv5JwRrjjXFtoIlNKUS7PL0fvsi8BMuTMVLzHzmXa8QB6GWsdMfmNs
Q9EDTUNsbSsCUFe6dde9UggaMsuNWfm51corzrYis5Hd5E2xqFWZAfU/yySl5aaU0mn6lurBgn5w
QxRu0SeGJExpqZPZTwIzjPU0RHRgR9xFmawT3UuJhJdOE3+TuGpcLG3IKoJ4RiZRXz+5plJ5uLEx
8PV/TejweG64z5GYJjekz37i7ZKikwCuXloCpD4/lWMFubFCFix4riR6FSkwAfzbCGYM4WJSOnF2
EnjDTqqi9IBaoTcWmeZKhtYPA9L9LCAdDeXyets8yy/NxP4SnkXhwOaS1qR2Iok0TIVIZNoX09Q4
1sbEZsBNEzztfasuD3mHyvWm/wmEDmj6smI8HGEi1dXP9szxk5AY2oImKluoX7SKwwOcGqsocAxV
qoH9GKL8nUVsyWKC5/8vG73V2325mvuf3EVRftHcIFQIPxSMTmEa5rUpwbG92YN6bNDiuKCP8wd+
f0yJeQ7QQBgRsVlAQE9aXxJm8A3qAzN9n/zDjEJyiyLvQaxSrRuU6nKXqLsIiRTrbvDRF4J+Vj3i
lzC2Cf9EZtFaE9Je9KrehgF65aWQNBWnfRspcGZBzFw/ii9UMiNaH6w2kgn+ZxqALbsNNt3oeTWJ
JNgIq5JhdhVaguZ/FZOnlXAvMGv5UT7K9/uNgqf4p97Ptw73SP+rs6RxCrMhfWx9qqfNYtctpnjJ
Y8L9TZJRrysLevLPMSxJWhFKEFYXA4lO1yyyT1kRSR/EWg+q5jXPfMCR/LUm0ghQPLPqKXF3gg2t
ELfZfrRS6DDAxXuBcmesS4XaY+HlX4XR+vOz6JCxrdUXqlbbzGefzmolU6FR1VQPWy1qoxzUdYaQ
uIzHQ+lFpjVVJW2JQt6/X2bBgCO/mmqTLufWNR+6u5cSg5Gr5xBhFcNSvw0QmTfNk9fF/rmoabSh
h98khcfdkw3MVZV34P/tKN4r7jgTPQrLZpr+AfZgwjnQP/MVRSLVQfBGEFYqz0rSjTmzm/lse/ni
xroT1aJ56XGMqUM1JMEvGQgxEwe82zI2tq3SL8K9GpjQIjgS6VBhIYdWx7oX2eoBOVGin72hbUt1
93+gSqmYa/TWGkGbgLiULnK3uz+9grUFQazqt8obw6lryzPey0M6YiVK/miHCUkpenzOiDffBTIv
5yKXr3tpV3X5ZP2Eui1ea8y+VJSVbORbThvBWQizt6IybjpCf2MCq1QXsjxeG7dfzBAw5lHAyMV7
WLV2k9fz35eXEMraGHZXs2b86Sl8kV4K5mvocUqNuobV3Qg3+T9lHk+0m2eh3FDmMKKBiAlpoMfG
uszMm+ekGbI91DChpSX/JL2mYTsMMtwXgaZ0uST6D8v6LBQGacbWlnHYV0IUeHA/b0hXQp1bhtXH
D9bF+/pamw8fbgdTIg2HsPQjpb9DNLFzICaH7modN4+EesMqD4w6QrPzOBidmkeZMFLLhcFCsC4x
rgdIJC8HUYvk16iMIe0WKTJkIPrP52Rh/Q6aiXhAx2ageGIv7xfwtHlonwVKszk0HOH0h52y/mB4
pS3vZS2sv/a+uFDLNYkUJeNP+RyZ2WfmzCzncBDJPfm82UmA6NqyUH0jhFmMiI+xLqNijZmz3jrZ
1B6zuC7CIlegjfVWUbyotEZPWnq2go5xSAzU77AiYObEkgK3Wp8tE8EdhN/u/jWUTeaA1f+Vpkeu
bC1x4kgrrx/rkjOumpo2CNTKqZnYOAqu70eiHBFEbEzrqlvSk4QymivihnlJfzkufnqKJRnSQRe1
OjG7yf0DLxpAd1oHxIx4ux8Epnja+ZHRYTQK1XKbaVyqCUd5qFqbAkaDDhCkkM4Lk8tOhA70P3FI
UPyX8IMHlgBvGKfn/X/nGjeaplm8Mk7Ib7xlvJxiRP1hN1ZYnOIq3G/Rnz6CVuMDJjcEQufyOD84
/84SFCrHO8MB+qkjUJHHPUuDWUYfxlmPuIZSLzMoZkzBt7kzBElsmqHmQzx/lnnTi4uSgplFGv7D
qOByh57hyPGhgnRax5qaca7D2SKdMv+kWWPo9MCRr3WkUF5+waTnCCbLMVpPNkc6tH00QwFosxzr
sP0MQRQVbeIPkJBNtv+5m7xIIWAcjKvI+6pMrE8SMIyO4RvfbYOYGis2j4YQ6Z5TJweAxI0ojdWG
IAloXHAVysLMF71y4Rt6hLd9r/+9lR5bRNqQ9F0L2GCGdXOA0lztnRR9xyZi5fxJeDnMkXv3P8lh
CDnzSALl9Gbb8uXt8hhzji+AOwoJkbAbwMpmMmxyoCh2qu+8Sdu5zTCEwMNc8x5p0dFqs4Mq/fsy
/GLJEm28iWZjIAlyI6QiTG8r+ZrYim7AVtcJochFZQBLihm8FXAKGhakRzKkM12PIa04rTQbLJf5
mFU5F59D/2Qtkb8ek2B8/8xB1HNaGy0YguWpXYMA9UFO4vx7IzVc+2WVzM0nV7Um3bCfvIviN89k
rv15N33cuK9Ztq8dX2aKVs5RoBP2/4hJ/KDWBNS2hda1TIUCIEbD6amHtUMCa/9dBt6MZ7LNFS2+
sRZLPzlfgkULVjeLPWQeoWJ+S2NdFCuedZC9+rk812Xn3hNSDWF9B8DBTiIKiL8pP/nLCbuFTnJn
LU05VnGDaXNe3touYhtURSLo5nuuy78E/upO4b+UvPq8n+H3rHQFAP3hOL0WoXE04c41H3fDwXKr
VQ5bkSZ4pp6iFwFzWFzj/FHK+mgclgfiHqOatqcKJ7qlBV6zCDzIlI+XEB8K1dm0+yP7XdJiF1/Z
y3aAAhQJeV51krtfkOsg5bC85XNV47Nh3FrcpRuEsRwNitjCcHf7fnmTZqcvkTL8Yeul130d9uSs
qbZYYCNfC1b5xIGtFwF2UaYciPOa+B6LkrVrlmjJRs3slfIEIAlpapRIa7XWQQJEymeQcsLLidSD
1KQCpHyECRvb6ZdZv1Pg3wRuiQi+s1X9W1v6uz8KKdTB3SRxsexjfK8MMbYJgAq4txbJElLEml8E
zh82JxZ69pJEmNHXhLgWkwadsSwkNUUxOCw92PPh8EA7X17JfkFFctSJ2XIuGrxdGl2HtdAmCpSf
10QN2J5SZUS+CUqOgdljz0LSA8mjTsrTE8MHlHk6pOwDHzk30BlS0l4yhyQSu3WkZsNS+UgyRsBQ
+OfvAoMobktT1+LdCINjudbJTFwe8Dlg37Pf/U3gWjaEVm7SRI/iJ6OkQMge5Ievg7skZqOS+xuy
Xr+1mB8Gh8SUTlEpPXO7jU3IsmcG7wVzvstLTP4s/oqOsmOJLBo0lqt9OeroymRMeYzXkKANvxty
MfQvzDbKPDFxl+GfjEImBveUyHxUjlH9mzXW3nIcSIdIky+28h7E/1wTtGA2WI4XhxKSOi22lz+b
/5zgPGnCysVlFqrxjEgQn/smpQOl6vJ6vejFYZH4l0aGF6FpKeDwg2UmYm5zY8UNSOk4xP8JFh7a
ozqGT2m2aAWCDS8yERRF96LPGukiZvMyR6T3omJWITfl30441L4s/CDh9bUfe4enbg6uXAL7bCVL
hZ+7c33Dm0d1I0IC2ulJaBJ2QHcz50APA7887LI0lJ/TWT881eoGIKbFJ5CYEUYQGGQIik14qKhL
5PkeQSmE7xFIAPASGSJBcHdKqkz80xMFagQNuQBuzHyUvMqlV4O1/6aQpZwRaeRz/J0zFFFwJYXz
AAiJ/YasXhuZkGr1Nem8Uj3IkiqwyBi2ynYEyCIorfvUn2BF7MyIekLqYDFv3+lMeiDWiecUuNXy
T/+KspzZR8xaWF0mbYmIKLL7C+e5sA8CeBL3TxcJV1sw30WDBe6x0SKCqld3LKh5q/SBxqzJBUbU
dWttvHV0u1gfeHjdvjCmLMLV6Oewo7nVSx7lrLpA4IcuzhIFKvtvN7/HyO0CLtSk2Z+LfoIlmvsB
y0VNkXU8cln0i3CaCKJzJCLtBV4EEiTXg8UmgtmZcpntIyeau5EyswSq3JpIvmB7hskG1NjEpgwz
njwtPDQj8KArYMvla7kwqO9IDXTz2CKbQRvS+uglTjPeQxT98q+0yTH8innIQGkoshNliyioBeeq
YYKkkiDd+T3syO6Fd/KHI+6qGC9T2ArcFPabpK/uS6UcHaBC2aevNHB/z+sfnRwsOpbyz0STzNAm
OyEGCO0TzXBZybEC/pgsHFeVb5b62yq2aPBtXYBJkeJEW5PCI+/edPE45DqBT2epSdoDXYPxUDc0
EhM0KlXuiBDvPa0fcV6gu+3YoNR3CkoCGPBV6sQzdgPyCurOVVVktSeTr2xrnUoN2laXk+bsjAuE
TtxW0G6QjIytyF3jFGzFaa3EjIpQVcMykUrUsTM0AcD5jIp2OENsmZJqCynW6sQQvprzXXLwxhb4
QUJPboWA8PnuNrrzkZFFto/0gsAyP+4gl1Rd/hztHHlpfDA0UmeLPgh/wAJ9xPtJeDvZB5GjQfkM
ObQidZDembQOzDC5tXpjbg+mXpEXbFL+lqq8Gfa6lkcS8oroPrB5hlasPpiLS3Lye174FStGjEzr
pe6lVTENuZ+SX2QUTlY2hjxJTJnXXU6DTc/s7ePwEdIQr9J53Wjm4qgrlhbOS3aFePWKhXgon/2g
6/mkhUsZH23e/pHDAdq9dHVUL9v/lNN5VYRX/V50C2OKjdRPTsQMY7dKPwp4Q7T0UWwaJrM8/CKz
C6dvKuHC4rwag3bLGidGsQql0yEdVJzgMqtB+XJyQtd4nlxazMnaCvJbtrNmNIgdw2Ii/+Gy/tFn
DjnqhS6SIPnKpubYOKRUci7sG+GCj3P0z984Pjj6j1Q2xBz1IHSmGqexCbQO7ySd1/y0V79UdFYD
U215halx3oN+41XCepZtfvGfaGs23VOKC4+uQcxs7l/BWueJm8EdPTG3LD86wSnLe1bOJ/w6HAtb
2Bt0yxc9o1PWXmqkrU1XjBuhPvW86NxRDAJV7rvDIOXuGfEWQoxvVrkQ2J73px050Fo9Ijh2mO5E
6Z5G3WbgiwMLyMxtstLAfPOIHidu3jeV05KwLeoulWjlUJg4ORxn/hgW0X9txDnn8m+Uq1WRS+ox
eE7BTemaIZyC2f8Ay8wvvDs4zSauz3iVgAGXI+gAjdR7YgvmMsou15J/RUp/yf8/szEefYBevfpu
VcZ9+dm2osUltbdk4Qm9dAi3m47MwZOBaXT+/pK4OCD8NGKbFj8u1JN2azLrGGJJ5OXn7SR5NWH7
5DewVGNCScUts62o/yrR3P6A6wW2+S0PMiSQcXbJxuoWmw8OqBVtE3qoEzLpiZFI+IkAueUyjtco
YGT4ngiVooKz5vpr4ILY8A9jdJPqMIGYuXLSzDn5AE+EisFCo2E05G1B0KRB+JPhijVLXSg/fwOt
zhn78hJh9yP0GPAdJSaELtMD6LxxJak8IQu3cN5/vkntamxBb1MWnHOCmqkXeoc5uWp4OQKnkYja
M45ZaD6PgR3WTdLChlz4upZy4TZSM0DZn+d8//3IX0peb3zz1png3UpiSWJlCypU3MyaHIHPfwC3
4lE8aZ18rOtSqi/TxLlpdysGKFc38lQ6k/KG/XoI7ijxcFZ7vlwbIHdaOKQfQhZJWMlpkdJzwEnm
W3MG+HjyG/iiXc989ScrfxSnaowKJifgxjjY88aHJdyrqeXUjmXpTG1ZPqypEsgQTDczrsCcbnFB
6/2XHDqMHRfuwZdgsE2HTj1R00FtEBfoLUmFfre5DJTf7zzYYLuI/QlHBaNGt0SGWtMLetHyLcFC
8lUr1Q7sXEWZ0Wv5hl0XOp3hMPwNyzwABagPBZ8vTFEG8x3ZSWj16oJjbSrgI8VT8ULD8pmZdgTq
UZc++Fp738BZb2xJDSExFd9Z86qi7WObPDycgqP9K6birlNEQpsmuJW+rRAaEUj1PfGcp4bmorOs
+OPvswkceD/X+we9d4hs0l5B3n0AVLBdXV5L6aN+AL3uk01QhqfppvWmjquFP1+LYhQzOZ+Ff0ju
YGOHnu8O/ENbmRzgLvuPoQbLg1sowTUqSLN2uhXV1qlKT0pwhEEvIqKM9ACNzV2rs5efFr1UFRo8
S3CyrawBgaIqAfZROF4QaOopzDiD9MBOOfnTv7fcXjq/amCxwb/yBeAAAiPGeQt5zSysI1PCLT3p
/kst4J4rkY4+c9x7XpVvoFHrn+PTAuZBr82X3egfrdJmwk5CwXkMYdHM2QFOWsBfkt0eU3WRgNwn
a6aRuWKOkNmcEpEcCH0s2UPU2QkoyJNoZEWZegHsMUYTpFjRMfA8aeqai5IAoCJodTcR2eE4dMcH
b2jVU+p7D6hp/V7lR+ziipibSb7ZaVAr6O57RwIEIRgcdwgkFnJV/FF/+eR69mUhfUPT+m54VgHq
rM1KifQHmEqkwTXViQ0uuBMaHjrWB4ABOZin+RlzPoNuOZtVREhUuAX3zP5clAbSCvHyv5i73OrO
Wye1ZGtYDb6DMEuHpa6cJc+YUjVS52ktvS4Jqpt2WcznG29v9600X1E7qrD2HyrDUjL4egjkfzws
DEMuWCtzlgWumHzuHNkBYJBD51oKFMYEAXYM9bAMyoW2+SZbfGCXCRKg0wWalGhg6PDMpVIT/rOg
Gs/rYeZn1/n1IB5KlYW0mY/MR4Os66xzfM5ydTT2OaBoKXa4AMXlWJ84LmY7bdvpWEww19e07wHE
J63wSdpPh7f+E7bkXxjVeHpmHt7WuIJ1jU+6tBKvMj2NBLdrWIDzX7lTmqHSjVG8CPNdTubwFkKC
6LeV3+jVxo8UWgpVbVVdJjnA09voqrjN+3QK6fmNshMeZsHO90RCaI0CeaXcvXZ2NEAS8Bu6OkbL
qAWY+wZyIfdTdkChRfYiNjqEE/7XpxkYuynbmbP0Lq9rPr7Uvfmvt44f8+W4Vdu3VZa3q64z+Kq3
te+4q0Gjibg2Hm1D52Mc6lmBrSpVpSik6YUnJryQEMgroxSutPauw8EWiJsarLOo/hxtjA08DKvn
MBXAnubuzQz7E6vZL9BMtRckE19XUeep2AFQ1A3T/FifmGZcPo5G2Aooo4AoCUZW4HS7WpLcgrgQ
FTlVQT4UaSw7hwP2sN/obOAu0X/ziywMghAy+AF04GBlAH9LxSbcrhLwDLrwPqMvTH5zoKPUttPn
5071OLvAmTBbPkGJ0/B06MEFk4C/e4yU9LNHv1lsyXG3SOBnoeaa3vjWoOb4ZLPfykP0T9ekM8Kd
OGKXJ9bOcT6bSKycuO9lsIUq8UJMOMtSOEXXRzIkSXiQKcohzvhDtIHodNy2Q0gjWfWDVJSlyA5e
wQDrtyWYUu/J/ImPgM3EYfGvy2PFj+jEm4MptiyeJpV5wuGqq+ZQyu+4i9t8vZrQWAc9molTREQj
9ZSIPP745DyTCn0NaR9fJ2bzm/dLkeYWZQyXoHu5LqTn8iN3sz9ssRtLKH8yNGSUmd46geklLFb5
o1W2Nxtxdx+/DRz1Ow8gA5biP77asqa7/vOgcZXfr9CNHBwjzDaHSlkabhwVHZENjywGNJkKsMCb
IbzfKfJ8bY0csqxWnZRcoF4D3SV5rSVljtJZTXbJrIgMp2EVMVVLcNveDw/k3Eca4VM5TfozEIHY
ia+sYM01pTDqIxeDp0FnTFErjAMbqWOyCMWUo7fogkkdwQukdK+QP3CtAS4KoIDNG97c2r8JCC8k
4W6MoX1Qo0m7r5cYLJiYP+mVVFugnvWDtAFA6mA193uDkyFxOd+4O4Phh/hOoNuKuBS9xkk/vej0
mumaJxQvWbIyLIoVg/zBIAJ6Vk3c4RJgGRpHsj0/NQ2Vj8CGTsfPn934x46F5zxNsrL9E9wugZdr
eZvu23nyEbVB5UyaPTzOm9p6v0sK1ldwxTorCLvNM9J6+YPpbyjvEYKJbV8nTzxy4veRRD5v3F0L
uDsIAJaSmA7bPEznZ6icT31f/hOxGJ2yNFjRDkOhBJb4Gxokwzzm0ssHiiE0jBVgMsyKxvRCMky4
Kn49+Ccm1MK6tSgyinZXzxSwOiSSkXAz82zb4CVm7+RPMNrFMcdp6nsdWT56uqIw3/IFX6qnEqek
zU03ma6zuR1TMUZ2aoQkd22x5TP6Mi+QRXpofsRwLvRWBIKJibY++vq4ypQBSE6rjwstSdNdinL1
tgJ9zAF9M9cOpvFpsdkB5imYIwAu3yQmmjk0OqZbeyhXuRD+yPi5Ke3+nHm/HJOY1bgQgqHzv7jn
8fFdTv5ESdLvDnTdUsOPylvXkzDc5xBzFVDZ4EQwBRtSYVqtnlju36TDsZqW0lKCxArMwnunUhFt
nRXVakiKInoPsM2hf8tg4pgweZrVKbbLNp4FV16R+l/Tmr0cTgzv1MSO3NbaTR+Fr5oBTpa/B0SF
RNyEbHQyDI3q/7w4L2Hn6pcxQN148DxoIADLcXTCS1ZLSn1KZicc7OYXv1wyraq/p7WXMFgBAZcf
QmYAIS2/psWATIGhK+cEbhn5wgKk5YatUdnWq528Me3j5HNt+j3s6vn89o/SwlJXwGml1TI9LevG
qWlITITB1x3egO/YxOUAg0RwlzZijhhmJcuCFNcZXCcaOzOfuobGpmj7QFxpXvpX4BmVDjHmfVSL
SAX0DAuAPn4ok+8EilLCOIUN+J3NvJzM3QHzpuMMr68Pa4gBxQGl6LSqAxT76Q3NMFRiU61hhRao
kKTwYDFe20+2hW9FNft5vYc1zxAofkkmgpGbMsxnTEeOVlGIoV2UjI0X782mZwbbQAZLPfT2THjp
zqu0iCezvHqQx8BNt/ZPYYzMLow/TGE410WFU0/7mRGmleV1kVRljnEpieAHRFeBv5ZUCUXSzdtg
sZ9wILveVnQBX9zpQmn4wl//fx/gC1+XkuOXbHxCPmWZsul+F0kdmtu1D7kRRU+HwBh5eaEsRWMG
6nqbfuNS7ZeMJceaxsjfPSXXkP9EppKljarf4yq35T5V3c9ngA21pp8a82GAfAS16n41TKeTwmgk
qtRysrWKe1riTEbxVZZgwwjjgYVqbvac8Vx1IEEB438mtz0YhVkQpFqdoQqq5rgBPnPCauK8sHly
xhKtbJ4W1TwXoc/Oobnr1wjB0bU9qC3XxO2LsV3FLRO+n7VeOvQNIyJYg8E0s7fFbA0DCyP9D8vq
PvwEyRfT1zx2ediP27fnSzquGR6TxNuCOV0Q1id1L9FWYUj5m/r0cZThZxrzFdKORinN4u40431R
xJtkv63LrJHJK25/ZZFMOEKSmNMJhc2uhdwOfeefXQUu09BWXdOu2Z/cmJuyXUgzrFjEn9zpfoIX
CzbOowGcBk0BWIDzLlPA5jCxvMmuhCShcGDWl1oSs9xq9hJmvd7a77gP/MrOIwvgjKW2N8A6aogf
8VT00EAKtz38ttmnzbmjXbsBwCKPKBACKEM/AY6Sq+TBv0NRwAl0DhjfbbkCG87mgrbDrRa/iHcn
2v9sVTMUUlhZtiRmwmUTdFhsVjZ4LIE2x9Sen6nA29s3kkv0FLnrk00Amyt2T1HKGH9Ve4O9b19Y
9PkpY9yyV+EzgnhruAMq5LT2+xohPi0NFCX6qusw8r5SvlmPLygsRwnCOSpmZnY9WU9xydYUYzxg
RFYrDyX/ld1v2Zv7g4tkBEsZFOqnuiUaa7nt7rrr2iQTq5sQbAeG2R0JE4fp2fC486AjHgvy0pbI
GfZ864r8yH2hz8f39w2+qojNiM0+y4XSdaT1SP0yGXDnTK8F6bJ9nfmRkyDn/IW6JXQgKmMvPBiL
ZG1rZYnZZw1tjBQMdgoZcgA3OFHVjhmE51S4U9zaA+o96unqHRE5n46BV7WZRPpi6Ytxop1oKfr2
gTgaUxgSrqlpj/Nj+9H7G5gBvMllK0TCzypXXQofx1sSzeHJgtqk7lWt1fBaXRReUpYwtKQz7XYa
r6pmN6pSv7sbPglKPvhyjp9i6Wo75BhIuUr+3m+Gcjs2IOtzuLakc6X2VkRpIr1nfj/OusFjyPuQ
BCBVfTffW7+FxeO1bDsYIHC1tRQYLYDXltmlxSID+vI8p1nHaD2TaOgfshf1l9aa+Nk9I12dvmc1
xpYtq6z8bqA3mgb3BmUTwD1ecH+iFuQODXp1IGPJV85mVNCL7BrfckgnoC6OL1Jrhe3JA8glCZwr
oXiNN/KOFKy+pV8fwJzGGuey3+ehIehEVcXa6ontB1bKtqBW3rU45sfa4wIvK41eHQ3GSs8tza5S
WmuZf4ZIZ90FWAW/L17nEi/Nie1JswzzPHlnxVemLgDe1ZaOu9cPmJxDTO2ycxSVhBAB5vIBNFcC
jIZ61LU42yJI/oFeDIHuOZLNb1+uZnMeflLc2fIPlNicgYrPxSP9knO2c1UbtlQ5s2ZLn5QRy/5k
eAK4N2KCHPVQY+xL1q37tqEIeQvezwD9kQjYXV1naAgWlYMo+bPVUN5dI4491eOUA5+ypZWCBq0m
AiYE/rAa1m0jksItWrvApx+LtM5DsAvojv6xf1CB65AW6eS5EZxsYbwcX8A1uKBggbOvpbDo7czE
My9xKBkB6u8u32RSjXtBQWbakO8azfMeg+rs1aqcJd/OOvM2HSYA6HJU8Agsq8wLr6wgYF49vQmC
7OUEVTBRTsz49t1+xIFxrw8tr9chDsRWWJVk+WoRhlYEzoZ9xDUEwfXDmAu0FePvof0VWRAvhgsU
1zV15d/InaRV9uv2r3IkLhKm9xkx/gVkJZHeqyUp6aiv8ooLRHir02AIMo+OuGdb1D5L/zJNrVqs
wGjQMlUxsR2xokaSVZ/sLbBgzJbMU+gQvi5hN4wU1oZ0MSGwfj6gwMb89vAS6BavUQLD9/8Qyc9g
37OBybuuwaXzepDsOQIyHPbcX1mA4HXpqWyIR48Q7YKqK715bPcOEL9Npx8rfUJ+o4b1fLAsywls
CUgjZzvUg1YTwQ6pXeYAPkUfGpVR28ErSl5Ada6s0I8nem7ri/6in8iJhExtriIhAWM74GSsnCmx
hV0KUL9wEcwWIF7ys+i+/vQVX5FBYMOuW5lhZ+5EcwQWP7f3EWOcPJWn2TwSJgOy6TFcgWr9X4iP
LeWvWagyxbFOvFiuZD2GJADP2nAcuuXktn/GmaR6b08ibhquUnYGOte7yO4H/Gm0g3K7v585MZ8K
TS+iotrTwiODYvwTcLe6Ur6l2ZLJRWF7cK7DZyuTaiEDMi8MsUmSY7RhIccg/dfq/5gCdCXaOXAI
h2sKcb0VmYZ/eBoETZE65knpikRuOqv+MwhqW8Egj3uHd1bt2SkhjqjVKojWRXNZOb0G3gyHRcit
HNoyKtBuS/AS7OM0CyrCWmprnhgqqr7DyQYWWgb3W4jp3ef4IJBobZcWPc3QZsNypbITnrVUOebL
YKnSKMe6tyhni6PzvzQh5cM7/ne8NAyW5MjY0n5AF+UydSRQMo4Ro+ZbHqXg4ZJuXdiDR67bolJ+
jrNyLlDy8tGkezaD8xIcETgmfKWCONas+7L0pfC7g6LyJoEHHLvCdeCPxNoz7MsHCcF7FFVJRhOL
Qqq+4L/viEflSZ9bo5zusbwYnRuK9KKQDP9yimMkxaN5ap9u3kK7PqE3XJpO7swzrKmefsvYEfwv
x+JQKVYMzwGxLF1l2gk6Q3E1UM8UXRMT5mFm0x6D/lKyCv9t1gzx7eFK2ewyRgNLUIKF45Szsiju
uw3QevY+UoBXcDtkvC58XJ97R4KrmWbInHD++gzDLf3k4klNij/q3xDe6HtVljWfZ/fgLBzrjOMe
yBlxgEtxwLT/g3sturyAeeJQupIxh/L14zSngDU3N/fhgabzH9dUAxyEhtt999rlUHkYYc/gglxC
HXKtLr+WpjLw4Bz6Gn1z2yC6qpbicqlByWLvbELuIrdpCDYt2ARnmN0Knp4ONKZhqGzqVG8GxlqV
rm13ovgs+PD7P/uMYMohA2xis0lX5kicKwPIG+LebodHCY7yohzwdCIiEAm8JtsozDRDvC2xHTj5
mpLAPHi2HPX7ssaMq9n/6FiokXQLdB7JaptgAN7Il9R7qPrm/FofZMo3z2QTb4JehkkQR36ehg1d
E3zW8yqQvtpNohY8CNyrbuVjerNjGTeNjN2tciKVIllqxbkLGhLCPENazgbNs8l4CGEYXZ1cgxGZ
zr8UuEfXucpGxDksuz9UT+H9BMii9OcoXNOGHLmqnHBR8O/9b1JqjKhkR1DhX94b1q75bnLdi17z
9Il2Exavzb93dd2b5zFmqMJY2u7hv5vaoYR3DCyQ7Mhk2MnB9r1AAvKeLxYFedsWXpsWGkhtSqJk
oEqrRNb9el4YNf6G+3G18FNMEUCtAvp/QkTL+gUMIJH0WO2SthekB/aErYThJYKBCLDuQQL2mN2m
JrABYGB4528aJ9fyZ9b9dL8vvvadC/UGk3urmVJg4cyjybj58bKUql1VK8+QLylLVqqpNGvPmAgf
wb4C6U0/tKK4OFil6UhcBYhUBxoNx5HBFGhpYZvzbYSsniMJFmCtonx1Fl70jQxqr9VCXTNSoh/y
AtBWZ7zGKrLUGwbTjaAj+qRQPi4ku6uv1e2vJSNO6Q8DKQ52sT09gVrzCtBm9u6LFS/bXgzmPaxA
RFgqj6hmC9hdUDRhY96JHV8rvoSpyQ02/y/JV+btqcllKj0GbMjbbimRC7Z8Cv26K7Zp7Mm8s9Zb
h+ODQtSK2LTAIBMM8p6lsX09LtyyViQl3hOW1Na1hIIl8fLnQ6IdrYZTzjqcC0rNf5n69ilz3omP
eQKzsJsFe0pzTyMigk/EEhXsmNHhB2UxHik5TvszL40BK1OImckHHETKmIBIfwze9N6iV8HXW5tQ
ZnK5G0M6w8H4WN375sKEbIFubf69F5pFT2I3Q28TnaUYv6EujuRNhUpNT+fKRpdu+V57QyV0zkq1
aEUbg9dd/YJoGZ/mZ2hWlxO4BiaJAIR4ijuQqbGR2+sR78mJMCqgxYYiOwdPlmT3Cpc+gECRUwP6
H5obqAJnKmHn+l1L4FX1VsdvTuqW++NeRC7EktW9fa+mP0k+w1Ofu70nAK7WOH1RfXDcGvOgSlJp
TAN1XRmyNFDlJ6+I+tFRMQ7sFWTn2MwUlj04uzeHZJv09HmRuNZOVDyOnUIp6n8LJkUM/8ml7LS/
4ZRcWnKvcTAVQk5HEFNnMDhPV0a6bGiqFyk5VyePA0PfEvQ3l4poClOJtfBUk0I1c1qNN84S89wH
VWeOvxvSKWDvHBphvre6p94FRgSnKEne9mSnUQHAQuOSLWwPHoWahSBcEjX8WnHK32PrGhKAFBvV
dxyn9dv6IK/tvVolvZjqTbicMubey8uBc0q3D3ljJVUwPpMBE5i8LaMXivmwirjEYtP+175BZMto
Rod2kUV8LPQN7wTFD+utv14NnRQO3nkj7pPjFTB4bJlPiUybpHtruP4LL9GWM7tevTxvyPd7kcgK
C8G+smbu2O8oyrKnOiABZLH/sGJT/m7OWQBBg5vOJdl3YI5Hnhhb1go15QNkWudW6H8AZEXsAbjW
Es4XDcoEc2qN3opOiT1bdubWoxuk0Njxw8Ikv/CJFYulj6yYJc9UU/t1ydOkZDVE9e3Wg6MoPvcI
V68Fy3yUDJxg1xNt9D2Rju9SiV8q2YKyKQhbZLmHBQs04OHM616dNnjFyTWYAXBfuMYrEuIuTihi
G72g7G6O+b5xjqRi2cHXnzY4RcB9flI2dj1jvoyeuV7aq/gX5QBPjv5EJojTMoPWl+43tv7Dk8nO
XKCrnI1S2uR0mUcGB5RQ2Kei5VYoakNhCPiBRXn1pRw1GLMgmy/9DSYoJvrrtGVGyB93+1qJ5tHz
APnJJzeBIHivVL12EApYEwFrOyHM+3oIfEvZ0BahaRiSsu6BEUaLevwbYpAlz9IhV7JsBtTIWNak
FXJqwTMjbia3BIBEu2E60LDjzVIsaBghlV7yt/H2hqtVTU+qdMdl06szWteIaoP/UsUZnNIYBO1r
ATXNAT9ddtLGjDhf0htPs3Adm3yGdVd1wqfyCajJSXRt1L6pAROKawU3dnnIyT0PwvC3CSJcopaQ
zM52DRyzwlUVuC44wkoBujVTjB/grd1m/2CgRvg59a0nSQ9fuoXXtXZcmLe8l3QyHN2Wxo0IH6st
JZAQHXrZ23jjUckBxA5mFDS8UBpKpTk57y7ojkgKtV7/IraLQ+RTG4nYcc2yl9l3L6INTc/cbyKT
Y7xutHXIQ9/yyIVBtz3wFYa46ZOvsq3UoOG7JyXjpzFyDTWQGnpJw88ZdtFQ4n/6+5eDvcks9Oz/
vlXeIVLsQvJp7ej+6BYzzSyVb74dDBLzkQgzwJ/UMRDnqpb6+M+iRVaY0x3jqycpJ7/m3/kfgl6Q
Lg3uKd4UKLr44W+r1BXR2lAv+YHvcSy3BGdsMvzCBlktq8hPZhmIfoecrZcbr8JxXXX+/cNex9he
l/ATo4/4+hE+0qsPRusZcPcNPxvw9xI6dagzycYnuFd1l3bbtcEE/b7FX6SUwrELgh0KtNZghLb4
zaOpY/0tT4GRlq2OraxemzA8uGpqiW70mXhDJStOpgSH392KoS08lN1EZGZ90SjBEUPHnCMPYKgu
bBom/52z+BGAABTpdUcoKCo3VXsP3Zj4lKiBkWLpY0mKYsin2meEXHVFfX/01om2fydlsw+CA22x
IFyePPBi1bW0ff6t8oz41d9rhUvhE/PR5RietffIiMS7xfjFJFgT3q9anqVcYitpNSfH3XVdnxZt
4savfV+CCNJBlhsXm5A28OpTTIttJGC6WzPoGWYvRtgTe+HAzf8u0maFQpdczYPVZXCrQqmx6BOS
vObcoL67ygGYQXmI+zwQtxDSBH5gFT7qm2O1T2LNb3r9iQH63NbYueycgTy3396r6lHnX0M8mh90
MOuvu/4/ci2CS4q9+mXOT9YD2YhUZCtq0Y0plUufxvCOLlCfMue0C4o+MWTJfmHkeHmAaSaVTv3e
H3ff9wBgs1n53MJCP+cJyzy+OZP8ChJeXmFJnci0ATfUN0ygawvy4saAOGA+MFxMSwtsVOJBSGaj
+XmL7sxNOCwA0rfx+wJWa1FNL5tJD9rVdx61RQsjmlEzfpS2LKyr9a70lesvPEuRWZhmzwGvfngw
REBbGLKoeQmvZq3N16q0UI71gaJN4vzcMDWdxXcTpknYvRA4eT+UbncQRJGfeS15PLKqwLHSE2yg
1sm36RbmKA75uB6P9dV8V+jskgKBouruWA+tnjYoWU/GJoTdwHMgwd2QPLycOg93v1h16KP4Xxyn
6MsuFyJqmty5yX157ByCgYekDxdtgTh2dTkKFE3CgSiDMSwaqZndaarjZ/YA6XHtS6ogdc537suE
3qhIPzG0lcbIzcvsZWtO6/+YcHylXSOP6UG6UNnmehOI8Q4cZA4INx00pb/93a9S0Hxx6aTdeKgs
RKKKqoxBJvuMLb4vREdEqDeW7VcwAaToUTQbv3d3bkIEWERI+YAC2ZRDpA3VELzdTwO3X0ZJttBw
s7715NLStlqrsqqDrG/4tkrB/JkdQcuCr+NqctT5ZlTFRhQIGfiFSLFIsSbWP4xuInZdF+1P0dRu
bgapEr1xoE4b0WCNjmakjfVn18KyAQjbneeKdZpaPlYqZk91vkxAXrEG8A2ZsFJ0KwaKupeEg1CL
C5vUACQ2JtS4kY/1kvuBz+jQ7l+w8xraFs9ix10CcHJsSS3bglc2ljPta5PqhYMEdqFJkjWSg2o2
oZcKpWogH/KQYR6KEi1tuWvYIjWyNGc89x0lSii/o/2ulVfiUM0hkuAlfuM0sqtypIDp1SzUSVe3
yo7HwuhE0mZePRa2FHAAIOtJAzG/l3TZZhe3kWugeEDxklWpLcrmfQlfmIwEYeA4XwuOfoywEXNV
d1M62znh6BFr3C1Llw+UjJGkn1/mfiMq5CzcoiSe3uSqiCBIQLR7tVgiudOcoRwOmjVMKnufe4yS
c+pihfjhdy4IhSVLYrcH8lDLt+IQvbZg4TwR09fGpuQtFbtZyU13YPgbq1DtVzTNBHaYjSYe2lkV
bbA7VhdiL5aTDTvL2C6jufKZkbbySrWFBXOTflOay6nJZVwFfqFCWXPIkw7ULHr9Bnf1s8e41l87
kh7oa5aJEC+mGxbcy7PNfXDnx6bx5YYhDuol8Z72Z1nfzyyeoCXiHN7eV8NGG+4jnLG/EHXU+iA2
so98bbi+7CGWR9kUw88wZqkqBJayhP/SBrTNyXk7B764IIwVB9rlhbsyCvxef4QF6ArSOTuoaPuM
GuAs7cQ0l+vtiD8zjUQiEZaMRm55Jgu0uYPXe1EktS+rUlm1Zps5m3MhJA4kEuPhkTM/PdGQF89M
TrBQPZAsCQo7m7s7nx94q7rsVb0jnGgOhvqiras1HUS3k9xBDovjYOSCWJ+LqYT1ek3vIhRQqpMD
F4f3xdt+95ORlHEbCOEQwKvLumNQegJYgDw8V8tfYDS0/pGqGE6M91JPwll7c3QLQQ6AITx/Bkcy
lEIXhMnkfYhMcX4dF9VTBY49ve7ub8Jk6NoaDkrzhUFB6Dai5Bc8SmAtzTjz73y7GPYmnol2qjl2
vxO56aSnA8EHMh4fS85C++zBkYBbTF6VIGEWd+vJFxvudi7RppkM31zD9C7/R84VXa+8vQE/Myiu
V/PTMJbpq9J2C0//Z7OPSXX84B6c93FXVhoTIWn/TX8GjadcgF7JlXG/1R3Wf4omhyCyCAtq6zPr
MOQRqkfTrrODdfB99EiPbZycg3y16kwWuYNwpY6pxtNXilEieetScoMb1b3Is6DT9eU5ANlD++St
+hlsv9547ddGI+OYK35K7BQMWVJWp1Wqv74mto8cBMPFaZXVXeMdeZlWFeMw/r6HTcjL3iirsZo1
5ZaSln+6zaW21fUENGE7uGGSYSegB3e9xp8TfdFhwAj7N5YkuQUoYHW3zFeOBMpH6JNTcdnOtCDc
2q+UViUmGbnl8Fi1d4XFBVaLWJbCDa/NWDe558clWxLhCZo0fx7a14h0iISpspzswIDA678Uzjd3
2nFB7I2ipL26Krl80C8sW4r/ML1fBH4ahOHgZhV8nnEwP2aPHAbS69k3GvJj8mSdprISSFF+fTHQ
daP0KPlKqLw/fIhI5ooxkK1X5p8oiQldT2Iompan1mUyIE5OylP+j+wTzq8S3GAU49z804YgitTy
gi2dr7vmGx9eEnqmS0O8KykXoTe1h036kor3X0LnN1uMxw/1Jm60LQIzppnChfN68nVinr7baDDd
X1tQ/nEyu+Pt17+Q+8TVCmL2Jjhm93Ryvp0XORxkQmbF1uhLTcoOAFtfTVefs/7MEy1LhMv5rBDk
2CrPFBK1S9i0zyY9DDACP7TWBkO1W5P/cNdIkW8DkaS1KVwa8K+TKaPFmCFjP9f1RhVtuq0zusrX
0VicT9JrB8qjJ2FIzadjjnRgq+/LqH1zLPXucmChINjo/nY4KpvOzcaW/WwWjxcDuYdI3GAogaSR
yShndw4sk+Bfi1aPxsSVtVtkOotlh4J7Z7O3GbE3g674C63/bH3obqBbH1ixH/DDtFbaSwRq5Yo+
+O6m3Ovb2458zex3STLeH3UqFXVS8AaYEcdM2UPef/qHyHMzHrgVJDWwtJre8BTTBS+8G4qzIcqz
eGRqXYbOitF/f9Znr6vNjTBSU7LVoH9elozaq8JT2Z7700J4fUiWDKu/Y7sd6Cey0o3lR7JWuG9V
A1ArW4Bb7d22Bf2Uw+wtstzZXgRBWLtxh1dEATe4Ty4AjVcsLVBvjsml/R8BFhYC7vEodygXiZhK
CxOIM3D6MhFOl40xq6KcBpKE6K4oxRQauRcWI+5dPZ/YGjGcbA6qSiRYkYWAZJvYcsKNEXjO7/wv
bloFMVzP4Q6JHQIP4M6cy2S1MgPqlKZh52DYB6d8fLBs9W+EyNfolPIhKYIXdZzzI44TnjG8BayF
WktCjd0FWdLo+QlynyLDO5ObIGhzdmxGaFl8Kc4OrJEW2in2s4vPaEELxy0Mom4qwXiUsHXneiYm
Cy8F9NWLvTLqYp5T3EOfMrOj7dsemDfeyFVfxGvnIrQ38M/5Zq95AsCUCRELEb4lIgMcnVL5cy9A
aMqCtVBZ+pr0O07vv7+9jG8cin3H8dII4J99T7zo7ue7lS3G7qI5iy5P5iSz9+Fx8Qoc6tinsAlk
9hH3VQIWrAHG+qgdC9aO32KshgT5fzZLs4AHHjLYStUcApnuqV2V+peIvhTO0pqA53WjD97SpjVQ
rtA7KtpJiLrs0pNuYJtCqfVKvbNEAEg60h1KGUAQ6OpO5oU4wSEQpFDIU9HcSn+xxvLE/v+RvkcS
3zeES2LlvOn3tu6/emkeAsbvngyR1y8qBoHS9T0DXPfF3SOgBm4rZGmj+It32dBTVEkdPHPOh/W4
H196trcdoke4a0LVky1FsPzlwIlwgyMOUD51B+UQaxYxmHWpI9Ba9XH3cjYx6aEkMtWB6w7ePMM5
jqHzm3L8r2xhCcxm83b7pnHJD6avQVdL78Y5NqmUE+qedf13X88sPgtNdEtsnv+G6joKFjGZdoLg
Lgm8cDTQjIahOYoG/wWe+vTpg59J+pd1mRTncJR/0t1m5L7SJLGFdpS1PflJCkbP8eJ1E7m6fhUw
Rl9TxChZ8ZFmHE5fpVqriGFIpdNBQu6uZLBn3c4cxGcjlgTP00vjYz4E5LkFf4ulHjgwY8jHR/Pj
t14Lz/B/3BMgNDCGDGFMJl79RJqHNGAInDpskIwW0JLRcg3lfc7QbnBI3NeIF45WOv++vC4CYAAp
swe6L7oIYEMy6ewU4Tx2fRKKjPskR8YfC89UmXL083hWIAevqyf0Y9mt7S+gAbI5oimNoC3Z95DW
8ctanX7C2pZkTjBnCl/bp4sZbT3K2lwo4KiwGFnRXFOZno8jVcBFksGm7+wpG0xDTQrTuZSxAZFC
wdtfRyhxHnoo1nxs41A1gauDI31QE9OyWMZ1XCVnGZG8b/COshcRnhTF6/OkmKnOHm/b8XngPfOa
KMb1vqxCSCbejuid1BSdtX5UCACbsLxSWSXz49JtzARJ1wefN8kaS/4IiOTEFovwPz5wRJAcF0u8
XyXf/+YZAXirBY8u2jEdupT3A9UgFzXImKTSvP1ivs7xSgUSAow60jhbibwZw9lra9oV4IxSG8mI
3gjtKf6CelsfeoGHLKNS8kfkzYLm4Kv3OLHQeDrxfCC5YGGQwz9BCohenOW5AavlGNVcLFhsFqly
NwYbhcV8VNdPThpZAxw8hTpFQ2weGJ5xO1SQqytfgBJngJ8eamZrD8eOw6eLyvywnwEpJS7/ce/V
DLmOVzzX5DmDVallhXCMEO2qyLu76EEzYiJKxY4DuGIL6rYj1eNSrByA8gZcXfWTQKj4EZE8BGO4
Iw8KThopqv8rz+Gi1Q1V6arZWYttOLqdDKNJKN/BYWYzJWd0nW2U2+ucupcyzWHGGl0N+QcYxsSL
VYlAihuG3n85CHy83yX4nJLPHfXyNzwgqyudMEV0FFcfyYaMPQp3cU5yDxlAJbxA9fq2kdZOfH8b
yKqx5LWiS/B2YpMv/e5oUsdi4B+kjzCsoMOgizktgRXxIaYABBcPUfNUYr6yPcO0wRljrqb7mop4
AzPX4SA2uXwf3sjR+0Jog0wJoP8V0sESPc66NGQBuf1sc5KSiSN52/lJGf36PT69ce0+C4XmGLxg
+iOMM3IpPfV6IgOPKgrgtNEf8euXUfn5lz4wxYy3DCJGk5szVfT8as4ooppoTgthX0VYwFMQiVkX
24+LiYJLxdPjV6HqecAu1v/C/qaH8xVqgtvMg4t70GAAH/WELSEWk0gHpAx5LPCrBiHADeGacNHI
/PL5ZsXt7ztPn4iWHS/pz4JxBoOwK9qw2LXikTZOy6SnLFC9bUaWDJjPrQpnxUsRdkq2ht7JDwzg
Fy9vLcP56e8jaIurEU/Ronh+rz4tGzvyDX7IYyg7q48E+IKSAYoUSqRUAZtRNZO0g9fx/S6uQ30S
gaEqnNg5hTkMNs1WVnAWrxfzq7KhOHy1p56H1JmP7Vx5rOb7EztvVsuXif4YHJW1ZURlcAd/L8TE
cGto4egnqjmVx2Um/WHR2vVpdeZC/vAVL/B2irGSvapwDhlTCf0lzZ99WO30cxZr1y5Gzrwodne6
pgEKvo3ELRnRvJYLaKNh78wIoL+uDlxPLGTcCQmpgGRT6ee78ucVan33j8YO4FD3ugv92tuvb3iG
sRErwm+mrwOEm8K6m+ibubVlQN+zkLAG9FBJHH45zmvNpEIWdKTCARcQlWYp72z0fRXxgO+glFSI
zJVxiDwqU6WC9Lh/szqqNA6kae5gFh6SvTgpxwvQn/dr2ObkZmhAeXyGJhOApuvCvhvSuQK7vYZi
6ugejh8DT5/lZg4pc1wu5GFR12kOtcPOe4K9RjoxnGWt9rhRBnEaQj3ZVLUP0/syFtD6EJeYatzW
LmdmgxwB3pxNNUs/MdGGkyHPddoEsf39wYRQahTxTg2nKd0BOjH9zvSuuV91DmnzaU6LWCi8t9Os
HoEW4vLxqz+lU7zRGwPKiRK0tIurO2OXxIbC+6j9ZVx+VU3liFkbaR6+3bVGpyJGYk+ZBKLTRdhi
g2x0ZLCSr5zC9URdYlHtDDfGmm870jmMow9OHBrNRstEZ1MTBOOlGWdUa21DvZBpZXyGYuZE4XF4
6/ROO3ZswVNdZyQjpFELhHLVpU+sbPx1dI5jZXAxdNrCZhug52JOw+nuHVFDq31zVMS9hezAFawC
mjgwn6WLlkKXGm+WAjfIfBlFrrVfY8laB6h3Lu7VDiQuFPO571fhBjdYf2AJ0DqBG2j73igJ5aL6
tdQdH6B2LOYMxvgRv9o15UoaowS3lDKQlUvYHm6Tq8M15TqKoSJr1TdsfbXdIhdAoe8sMrH50DFB
z7G+LvHW7hjdRBjKrhXBbeiZzEUKS5HXjpA7dFIZbfQPNFktKWQwvtyu4YOCQSnBtQok3TLlUo77
yFuSs057xVkS2X/sqfMT0c+VedRdkZSBJgSNXBrFIbKB615kYrpzgaXgfXUE6e70+wHqejPkls8w
+fzNhHsVkoOsCHJPREECeG4oMujGIb8zfe4QOXR5GLF9/j+3ggXhRh7+j0TYe21/514P5Hm2liVj
RP4W3c34QKplxlGnm2XotUxMomo3WK/8wVg3uuiryi/zOcPTC/Znv2XsZVitwmJ8By9HlqPnkhkd
mr0+I0ct2hxUYERzH/RYcLn4eQe1nHZbCJ7vptIhFFnT6KY/P11uVbCsLlovneA4ySv7eNDYd3MW
GzI3pSmmPOFPrt3SbalEkx5LzlQF1ynHBRXk7qdaR89hFj2xi8agQ9upFTFESvLSJA9fCQPJztlH
yYByLWkP6cl4C8c4cB8gNxz6BA+x0dCPqdXp3Nypoe3YgapYWgXya5ue184optnT34ahXT8a34mV
fSKK+pxhVU8457EE+RkWDYuq3c1CF6IOC6qt/btE2wtDXeJJTUzT6t0Rg5LbVYocJcF5AA7f4sB3
hz4ZqXBohWXS3WUxwJiBNZRfn/nP0cknJDV8yGcc8iVXGbVFA8b19F1zzNsy6RG2BTWBAjeKGrTm
rkPo315d5jpL6ajyczCmcvwzPGJb60MaMQcFz4WagIEnjzg/xnis4bulc6qULcsA8qHfK+BJBDK+
8l/8b+cuJnPX2a6lJmWPSN+DuUdYX6lAKEpY6SgRRrfIODdtU2rpIgMlDfVnBE1gvdklHkmqi3yR
Fsh29otKinSn1BxuBB4ne25mxnl5OqDkBQJK0w5L1bbYOaaNLWIaIHG6MTXfTGOwF5NduhSdwNdn
emVgaC+t9RllwOXgZzoJHa6U6Z+Qiwey43wM2YE+8VWIKoM0TABes2R+iWMmwtNXN4bprKo75iKF
jwGr4cVUCOCXPxKMfraqTyOm3XdzDhUHjkqyyz5FALErthDD86afkwIq7h354B3vz3bCgZDust6/
dAnTiCJbdt15+3qO00zPZNksGae+CjkDZ+2BgKy/M3LnhTsXFf7oeNVacbgmz9D3qWrjTRygNEDN
CyNxl/VVzoanEVnZTAsWrXt4EIkQKoZUpo5rQ4Q5ovwjCD8hCS+4gL8HpRbPC8nUbOyXxNBNkVfX
aPGTOLQR7WG6zTYsH69Nh9jvlw/SuQE6DGuKjVzWbrVqS0KtxukDUBSiQ5FhFK/0XwFQKQ6RgBBp
VKQbEA8MWLwcx+S+geTgg4sSw/+08y38dmmO8VBzZBqzguYJT5DrUdb4vyE/kvVAw5V44UXaylkL
IC/9hNif4OfqTEm3AEKZbnr+DtF1kPlQabqxglcQtGLNYeLjON3M23NKUoVu4zPSc73YYMSGt2ua
YtQIjV2oQQX9PhHRJ/q6FaTIkGesRnXUwCWinfPcUVM/jHr1+tKAMH6yPBYoF28tysk8wKCWQ0U0
J9QdEJdiVRHjoGANjn1TJ9kASI99HPnBoQtxmKFs8GEf+l/OHVGA3NBo3m4JX7gF2C5wjhu3FXlP
Ypt17dQXSaGJWLaTrDb1/FRmPrcKpvRRgRseFOYBiq0Uhp9zxrOKhX7GruFUHhalThPow7R42Edm
HaXYaz4GZ32w52ZH2j0Q2q5WEQ2F0SqZGcfTGXY4urZVK0cQifnCk0N0fIEKozOE6jspKG5QJ9o4
FJ0NDIR+3tmHqLNsFveB3FaJiQL7gqBVBg873Rq3WwgURzNSo1lOOTJlO0RX9lPKjIdBrJvpOi0S
9KgLbIw2pSGwP6yrMNQb4oqcIZkCS4ILpXmtsUF3o7GO8WiTDqPaq+7ui9Eihx5Y3r/BKn6a89ey
t08R7CevyKqpIGhVtwe5HWi8joJLJwGVBOROUVEHrOHNn4op5M6+4xTKUWcR1p3yJO5FLU22JkD6
NtLFscIWeCRYC+eEBpmN8o4q4A+JYvu/XpPTRdtsBhfBhehWschmVEwioT6PGX0c8W0ZMmH5N5Sg
65lKZ8QjEX9GE1zJiMN7fQ8PJoIsDpINnCSFwc++/EQJmzCLMb5J/Nqo611LEvjH/5bKiu+EKTIq
IQo/i+urc3VCCNWSjD9828CTWXFZekW5RRTz7wra2QaMdPF974WfRGZRtr4l+SN7COYLacYU3zRy
GnTlA/korXtymjmbqD0NrU/reLCs1Q9k9TVLEePscOjYeoyxzSBYUJ+sq+t0hgATnaCYW93M/BXT
yl7labyhGym55XA83bOa3Pe3CB3E6NG/MiRHpU8hmcQFQsxQqQr8pFvyd4+F7RaNaAVqS68dXyha
UDF8Jeuf/84NDwlY0KaWAfX3IY1wzKGfA7LXttdBebkM/SM+vmT2O0hXaITLrfUDNwytOk56Gx1K
8gHrgX6BeFMY53pah3RapGJnX9Uhc4SAcNHbJtIWXqviTQUpG5VAqozEiCrHooW4ppYe53hu/e4u
l4HzHWQkQYnu+LOqqOWhiYYGDsn19jSWQ19ImJZ+4Hmo7KVWwgTEXFEBUYKCjq9ttOl4bE5zhnI4
0WBHRJuosEle/AmA90j48lpl9UUpPsQ+Yc/3TxXZhoEEPJGRLH4fcINorefbFyHmXpiRa1A4AUxJ
BJ53p2GNcxcNvyjEpLLsf307ZiqRE7NHs3oNkM+9d8OqUqHLRlxwXHSs9dBVczbHuQYTBUCGo3W8
DTwAZN68wIg8OmUgcmvyMjhB7HHkrrj9TgQk/2FZWnVClzhG2UlseFQO8f+KxUfTeOBa3UID8WHH
gNnaiVDTPx4tZTg1Z7kO5IKwrI2mxjwZTA4yXYIgJht1b4C1F17jCATIFw6eMbom6VpGlvd6LK2a
v5GsXmTDAcU2NlEMGbaxYQguwaen+lPwoyC3EOOAjVUpekN4axSowbtvUkHShmDV/eS+5jAkwJ+B
MLZIK7n2VNSnKpkEJsTi2vgtCH7RcVsOjChF05vLk2Ml1LnWHFBgfLSUjIcgqofp7YBcUUxZlvGv
c2g0xKvyQXKmKWBkq7qPPLEOOxBSAxG/EHZ4CN9oaUOxM97KUFydPrSk9d0MKSWAqyls99UVt1+J
3AsVQYDPxqmnyy1jeAog5zIXLzrDoP+f+TB151wZ3VXQJaq/uCeG025wpSu82bCImYgshd9JDhKI
24SH/2jqb+RmJY1YW+tjDKezdTY2N2+tqXvamd0H8BqPJ04qcFnsnQfqDwxgGIzcjkC6OBNr0FRR
ysfeHnyPZcfzwlKOpUxpi5IX8AN1bwww99E+11dfNkIVx/5LJQpOiju5p+H/z9Y9+/pUUtqXXQ4W
/TnTtSpzU55P8exKRhsncd0EV5oUv8MNfkzpM7sVMO9+V0o34JJyR5iM0Sn9wTC4KipCU8pwFif6
iCsKrQdlzzSnNJA9lxyzflO46KHWREKuCclKulpswBQ7iL47hwUSSc2KLofpCas7hDchEjQF1OJ5
jR2JjX/zqgUpIH4NBaS1sYzu3kgF1xCclesSoaByMoi50y8wdp3RzZmgsG2acSeFuCf2hagh8PTm
lw432wFqDPDYdOeRdWnqkeY06X4R+kH9vnQAANNho2SxGY1SNdOTLZ4p/FwgsNYU1inatDClWBgD
f7XA+l7qojdUDqcGkp3PpvIgi7MLliANWcdigbVCHxMbdUTIauzNdojNIPEA4e7B9h7tf0fh2Hgj
9TSjpD8cdOULoga9KtrlphiS71guZl3TfjkzSemu9yx3JUIiK88wJ446P5VjjINO+oocPqaRx6AF
J4vthNV6QsgrFHs/7R4wtOLhd6s1/pzMJDrBj/kiLMu1rT5ZQ8USJ8I9yNcWNegzzGPj5oqer/hd
/NgbkYmHrEfpG1UsJS5Yf8mKZJv2JMoI3eV24Jw3awSIWBfu0IF+w93blysbKMRcBut5bFaF70iA
oRVRaCnPAzpx+J4a0OrtXfjM8ngd3g5dB84oKZlgubRAwMAs0ACC92ZM4pBtHaemG9AwMJo5JmMX
lNB4jxUC971dYBOpSFECyqZ6WKJuUGPDR18LQbPiCINDA1GA8gv1De8OdXlLa+NZeaSir3wh80ry
/o+znFNaa2XyxtjIixQxLaicE61k/6C27UL1XJpsY48Pz28y0ED4yGYhOHad3dNLh03ZJhEgSM0Y
O0QpJ+ao1gFMUO3l6bZsu9FvC3SETU1UQm64U+yGpqj70rlVBmjHrVBLQbR+hwRGqwrGn3zDLOzq
CqhQuT9pYXfxk3AUXudg5bxH1rHvu7KCVT1sDY3iHRFNPnBSK7nRRORt7pSEK3YzhWpsGN/ByNVN
Vv0c5otO4864CibIOEgQBu13Y5qBJ1Xm87tKwPtohMGXYyQHzgDpWFElt9ujUwrW8NxIbK9wCpkv
6ldh3rjylBCHta9C+28bG8w2OJL/pXwsserP5ssGqubMyMmsxo/IIX27KS4oXF4tvpQtH8krwX2n
ckEpDHfruwhNF0bg6oUVv3/wFS7o/p6DKCcu+uXU7PL4wPv429ZSEWTsGcwrbi4WOn97QyxglIzD
PWs0DvCfGvbAV+EhHfNpZ+Zd3jQcB0/JR2rrfxv/Rnzh8V72bnAfIdc29djovbntbZXOKZjkXoHk
h6iaMZGrzkn28Gst19xhPh86N4t6fvr4RmnOCKXDbJ01fW7G+YiGRb4UlYU+gvh3Dh1BSMs1CfMg
Q29f4FCKq5Vh3I5YmPEGXXakcNoJ6oNGkkRl59wHoMZv5O5E2I8pLE19p7fm3+QPhITYXpz2hltv
ZCv7JINiY8EXFuZ64ckz2goI5Yr7o3+1dfZ/2Klug6pNAzyfU1pN1cq0yAMc5XozkOsKy3HJprKT
oqdAg+QMJFT4XOh0Jmwql07JZgE4G9BbWGBlkxvzWihsA9po4DAUJmkZtBFszADZ6P8QRo+TMeYT
mPOwlKeqMZ2ae4ckA3WfeJt/AqIKveuCPvs2/ObYDuyRchU7scW03V2Qk2q0d6pffoz1jVN3a/8w
z5zYPiAykwHeToEW+QVTo2nvjkU3hgaPRCiV6GnCFgJkfqeiju3ppCEmehIipwbQsczmkAFYqvWa
xw015HQTXffkzRwc+1+13y47obMfwazo5eupnVViCbmBHw1zTMcfo6cG+YTBxWvqiU6Z6zDOlFPU
pIZ7KpPljfo/rCPhLu7Z7h1q9k/HfdPsdFDNjO9wsMGW8E/F1XOLwsn0OjhiN2rnOE1ewTgxRbak
U0VD+ZhJgGWIHrRCpdgs/qXlR1fZ+K1ALN7rZb+xO6LIcDY0RKmo575k856wNGks25oLEy86J8ZD
sdh0zyT+BeqacL1IY5SStEeVyalD67R17vTVXyAkCORhqHNee+k5+u1vNVJ1CNZnI1aoS12Zrdt0
K2gXg0d5xmaJuhjZoksoBgvgV/OyEohDtEuF08MlBpbBKDm8youvYYbcR5jc05YmJmgaR9xeS/oT
6dCb98wfhSN/osscGomnKp7+taOlsSHt3PIAfAUA1TUIZkm2GGhiqnEovDGIhcwVGmKd/ph/FMg0
lukQfFJHkSG+Du+HwQctFFMjteEbVvgFiBgVjW2sgzS9K6oYiP+7FznqGu0xNGPG1+3kQy3MMm+k
QoP5pH68JBMCg84MLHV26v9djWbOY62Abf9Mprpkwoh6+2+lOu3RNLwheLXyZ0nwQC5dD9nMA8RS
eeh5PySpXxIPROlqqNFXZhZ5gpLQWpBo75lr2gf11at8pwwgo5kuFkZwkE1npr3g20rLARgMBU7P
q80lK9pW3247m0q1+10wZtGBQkwDeEBMtlywnnoKSacN23GXB1hPUQ2jH3Vg7u5ZEzOGIueHMdDJ
wjVmDvwbR0PiTT9cf11NZ0KyyKqeF9KuD2r6svaIWQKlLL32lHbT9304Ihqden4LM4vvy7lzojWh
KDXdktqpx+Wxg5DyLCPjH+XmtuyleBH88f6dOiTe/RJRioiMet4IGYNwj0ZUbwLg3EqsAtEY3ECs
eOo0kJFe/kH9KPTTr2kaBUjmm5HdRau9J2ysI5bVy0ViAg0leXxEOZLPYRbzAsldsxv6bOvy8M/6
xIFiom/+YjQ3Yyioq0WiaC4aQLIWRyF3yMxwrxxQapWBsjCWlcNwOEfSqHebSH5EsWp3vnSfiXpG
9DS0WUhVwg4Ada8HH9Od966+vgA0dZH6RFrGgHjGYwPaBF4H7UbIEwevAHNqfniDitOJ5ktjNwME
SjrxCmffki5a8Hhahg1JtF6Blodd2HXq3kBshPISuCH67QhTO3FXdTQ1rqIU1HtCwOJTfx9YBfAf
69vXUMNwQCqyINVTe5ecXWky3Ayj8S+kTJNt9dqBD2M2xPl2Xz0iupcq364KcqoxzzwpVdYDCpcq
dzTcULJQcWBQsqeki2Vk2j7+MUHDTfAM0azZ2+YK2K8Xjti/fMKn8eZ3Susu+ay+hr77hR8UdQ5U
1bWnPIU+0icLzwHb6wokeXEeyHVSvuf6dYS0wMEToBHDJ8JNtzPVb5Yk9nFaoStqHTsgWPViT/BN
23gXE1//pxVVMI9kXjzCDS3LyC4FstY6WiRwp0/CuZpbp8SEBrDp+Z7O3A4fXAtmyR///Li04E+n
ZxSUxzyFY7ll2sRfLpCj953goO+c6LduKysJOv4zfskWmSyNYlv4eNeyZNqQ2ZLE8abnRjkSw63J
7AAtC0u8v+eFd/STsxg5XLUNdpauUyFwO12+mvfib55uvrdbCpRPduOtBkHYUhJWnd1qsUfLECKH
Jk2r7A8J69lM1rZZZNeoZbheOvVnasxonNEd9T4olCXlyGr2QchVkfLIm19bNfi8b5lg74cqiGEB
WCFVwGqaMd7EvFF1XNIXhdFviT8F0/ZNRcKU4of8JYUCrPP4tzKNVZRugiKQH0omuPJqUQ5fY2RF
ZPjRhopiZ99rAnMMcFGafKWdn47wXa7OrJf5xB49yNKgzst0H3DrmfpW0FejU8qiRNJ6YucjHXC2
llUEoGjTd2vLp91pFfxNfGSEDOWDFtfavZoppvjo9pfESxqwczLoMooVtVgH0BLGzpzHxlKc5ps0
zytqofGCdlKvOtkfYXf2HC+dFXpX8HjpeM2xDQT84eg6eUy0c9kM+EMYD/EvTIa6OwuAskcb7qhG
+aOYATm/ZkHd6tFl2HYtc5HbWH0uiP5cRNn/5uGN28MWngnRT9QsC6STo/QK5YdoohV9elSCPTvK
YQeLH22eUTQlOJldrQP/Z9iLQ4MwW3IQAOwzz7R9Up12br6Ixw7sEa9qDffO8yi6thP+GDe2j22K
Fo5r6pMGFPasSOg2PDq+xRzqS9ve7fST8UY/75kCi2oeret24HW7DqFuLAr+k0K2LzCBGepDnuwf
jzvpIDXBx5aC3vDNL+4Dn8z0QseLYWMluN3BQhX8eshSd4mo3AvgEmRWFUhlUpvPFUy1xR2xP5kA
gzQoFNvpyoOESWhN/yr/H40w/blmBcEm5FQW+ZEWhy5zUqj/Ix8hg+3mhDDuzNWs/rtjRLjJM3El
4t8K/2mxG0DFicmhoblbMCmvA/Afwi37DnT6dhw8bfb63SCfcc2mo+G3SedBgHy9X/fGldH9ETV9
xoIirl76kjS+YxL3P6qOueBBTbF02lrxDVLulkDhzfixlsWQECx4GJ1YTnNRZygEAd+vJF+AEKZQ
WzFMrMvasJ62dTDkxw1yRbBfTEDhM5u8W+GtWMkGdrinipkneNqKNJRhNuJeh2mV21UcnH8xK2O/
ROqOByf6pt1oGhcv0pFR+upDX64wNci30OPKaT+IGrcnrOTfQp+dI/7u6iVALZQZ2TpxpUWfOSy5
8B3YGSbFAZygACkLbF5c7ys+CJmIQnZeC8HOyS7GHiD82LNtWjdXYkjrxXEDw7I6+tLB6o/TApmz
B5ic8os9JTrgfMt8QCfB/0YeUc3rDfs5yCqApPRQfsZGPSOu8lONlDSn3MLTpvtedpbKwqkC1r0Y
LPEOlfCaW60yIOby60TH6+JBEoGtQ4ZSPoWQQZUMenjhnFWyafaHbfOyipKye+K8j2VkJc4xntbt
MnD0+D34W08tqdYluqLrbYUYX/OaD+rg/HKMMKz8Qw+Jw6ToBUZh2f1L6ZXaaJoirSk6ubah0o9N
JtZU1guLQ88gDlnwPVa70yiaY6cIuLrp1YSYYXLXv0IMgc4dkKaug6WAKY80Nog8DMSWOsPkXPBS
481Ca9AqB1Hk0Iw8mIJh4qOcQaEMz7CszvCVtlEhNOkdxCWV4UkOsoEUyjGf3/S1Aul8JFmWwb++
v61PP4wn/F2Al8rsiZxt523IuN90wY3MoFr5I9Zno/v5oycfTQpzYCpKIGvY2O8r/uyv/kPtsMHd
mJYOPaEXA6/20eg6yeuhrPzBamd825lacCBUbn3JFdFCJ1aiSSrMggBtH7EkBSrwqFZ72GShHOld
lzsBBeaGA+WP2mOCFQuUFIhJsNNkQU459Mcrn1Ezja2PiG18XYqa6tYETO5TuLV/p+w3HaTr9VlS
FY797t6ZR+E4zjviHDm7h/c2e4ms/lD3Qaq3MMzG8VoXeoBQ6rO/dK4nEHxulA9QMo70jm2SHllS
uEVF3do5lVjXeKSfvWVStHkNZryQ0eCbTIVxjF8ZsikktQVe8YR1gtRSvj85X1dFz8ai00exAJSb
qnFiiFfiDF7OA0RzfIQyuWQk3EhmypXwozhO0ba2uNai6qqCivPRnqFKf6bgUbPIsTOg/B5JoxuA
FSwaY3MOGJr7ZcMKNezO7ekV/UmF5FFheipLcVKraRENDvt8iGZTvIs2viTQ5fPmPPByHEjo9Xmc
tUSt/beWffEtYvqfgnedQ79BODvzRyTH/v+5IDjVibOlRG+PQWynTtrUsEDONm9RF9t0gAgRl0du
O01WsUQYsFiPsY16wIY4cNgzjVM5UypaJGQYGg3Jsj7XKH7pY4RinHfbi6PuWWKU402BbgKA6pW1
A95yJaizpacNtZ0Pz2kBnOjUiRVQFZaaDHvtdMs3GbivsuvSWFYXqhQM3GvCCerMNhww+pMyVCBx
rMW/cOMFe5JTsx3s3ZmZfVwBfUqow2Bup+rmqlvz1g1afFyrGzWL5jeKsYu061itqt/7NayS2/n7
9VKlfqWDL2K6CuEjlMcltD06kMay/FyYy8b8xom0IZFJxMbvFQEvVCnr+4N/5VnK1Juk5UjdHHNY
RBl/QnBCOZN+D48MdD6uFxH6GRkOoqU17zWfl/6I44liMWbRzGlxX+cqoNeYv+v0U8mwm2jpgZ7/
gQ4lnBdWT7suGB+D2phoDVp+4mxjf3w+BvjP8H7PuI7b2YdbXwbgsPn8m83USmKjEnBR9Lhi40gl
h3cbDamaDgfPh/NIvITSxlwv7lsHJaAGFNcyAi9oSifyjkfwQTAoksehVKWucy1VAqDYxrY29UR9
0H5iNfJM4aTW031fJ9+EMQ9T/4C+dNKMs5HdcPqZwtUa4qn3nW9uv4O7ft4yOa76zq4Dvi/X4QEH
i2rI38sNIDdIFc5oOKDx8y8QTyGad6KB3+CLzuohEQyWcLNxx+abDS6EIBeHscDyDH93/KxhG4IV
MDg1KCdHALijMwnwr7ukQXQo0PFnIGHl+djUnRf3pFj2OkeRc2+ZiRlLqfelDrg8C/WJ1n9F3lw2
tthXTXBV47xB0nQjmjcASmJD0wN8/vcmwr2LxsjJG8AfktaQJMx6K2Xe/AVb2ZftxFW138a3W+PH
pa3lrTIjs0HY71XYWQCrotm5KjEomSptd6d/sD1nHk1E/jzNNmXExCyZ9670GmeeK+z5tUCajKUC
m+gS5i9LJE54CQmZBd7zl/UNLuRpwg7mfvQYz7lNmFVnXyVxIkAbK3L5xcGhB9tEv934xZOkvC0R
nBOsIaSZIfnFogPckOCgSmw8bRRSF9DUHTuU9PWrgrOuG9Kx/9hn09xPwIpYnIK45TzktKhhRmqo
MWDFC3o2fj/3xkEMXnggD1zv+VbOp4mTWlB3AWaCO2rKcpfJ/8XBxA33wzsAyrc+VUjEAqX2CsEO
iJl3RmAp6HYggHxkiupHO/WPzex6kP+JBNohDG21jST5bEGEhuyhqkZOy+kYiYlkhDxuOvbhrMiq
cUAfrMI5S+7ruzKLrufwFXGzw7CuryMlWcxBXCeuDUr+vUsQq97zvz5XqXxaWTWvfHA2bt9c+Ivk
mFxcOQLQh/1fd17obqsVKhMBvmC23zfereDm19EC7TNh34Exv19je8IkEpnDg/aI9Z0vjgohfUIH
nt2Z9j4KQCERlUL6nSknkMwgX08rC7P482YP02pzedGYvbdd1ro+WMaGVSdxmwrQ2hZOhSQH9whd
4z6BLCk0+16hbYA0c5z12WMU8DOX3xb+NZvXH/8lJ+J7setWG8E6x3rF0Y8Yuo5ENUphkUBJrFl7
9s1Q1RlpyD3orWnEBfQ0newtAM+DFMAV66W/oHeu7jP0va3dwe9PH5QgaIQ/joiwZ1WHQe+OX5XV
NE9CLl21tY/8mYXSYVLGsbcQBdyKAeh8XQs1WQCSwRXsftIS2DYhSEwL9kw3L6puXXLhwLn/m/1i
ytC7HFcKY9+zVybrSPtR6JbgMN8dJ6q7wxm2EMXW9sNP+/NCIDi7+hgutb0FNyAFurWAQjtByjl9
Hks2Kt3Vhc21mGnr76pmPYF/oaAA/NZ6FB5nFwt3C6EYs2ASy1MWNLL+ehn2ZgNrmo2z7HGRwjR+
ygLgXrv/SNBZEvFqAdf6wE+UVED5pEMSD10wA4NnPHRAq2DddAtSPHjz18suZracdTxwxJh5B8CQ
AVBJ7Se3DLBF+WzR4CMa0abPvmxhzRSdKjUVMrSiwlNimD2I16I8p6D+2yb86Lb3BcNyEo5+RWbG
PsB056lOSBGOCSFdvvehkuqT4NqRitl/g2Ip7pO0opReY0YHYQy25bOT8TZ+MDFqnJmSDAAaRBpu
SyQwJa/CUNxIXtT1XYIBL0DSuia4z5Fae8CJ7vxNX4HPOLnCPUAIbvzc5Cjd8f2pBW5LfC098XLm
mCayATzZ0g1YF4oF0DMmDqj2zSfrNs2SfPy5kwZi9lg6POcLQ8x55OH7LDLU0+qSrjOR4/w2GKUU
uViLqvmjP2zbiWkSwYEkGDQ2zTEwnqpvEDZNEXqQSphfpqBfEUvkVIuYXxCUgtcWQ/dZPrr5iyMT
1J/6dOtJlFLyrqOI+v62eW1FVITkKLHrhMEl7KpG+ynvM20/8FPoCaBxOzGf13nUKfCLrhjiGxik
8E/FA3B9Ne+jAx/6HIcL70i4mS76sOiZQVOpIy7daHJcNFrEPNW4CtYmXXYzheRxdykXOZnB/4DX
k8rraWMM+lywu4wrrdFCyIu0YRLRCe18HAmc1sDc8nhB6f8GfjueVwKRa7z5OoEq0OBIDh5hDWSo
PoXcmjK7hJKlQskxRvKRLvcF4HVVv7xu9UiclT+aaAO1QKwta3yICljeCsS7zKMiHOJ45H7YW6yG
JBtgX9fzbjukzfmA4tOV5afyt1BPccXLUC03dTtHIPJOazccTkJ46zcKWF0tz6uQLByB0aj6NLUa
V9g7aqIb5qfNcIv6iOqE4Yt/sAwmwxWXzzBsA+LpJrROkN1IJjWTSVkw9hL42Z7Y3loHNRQdZ79n
tlOR7VFbtbdA/qC3UZs0aqQOnatrrBMpn7/AtdN5CNpJd+CCU1k7fv2dZyzXCfJ3oi/3klPGchhF
QEEddq3ST1/i42noZ9fxSiGmFGPiPeTSKIF/c+lTEc6KkCuV3F6E/fqa3yqjelzXgmsTQjZc8dhA
T9jrnLUWEHTcGLylAPJSqNH7yWlBDvxh6tEWuV1Fi3XU1nCtvC40leUgHX9L9MzoyFyfz09F3bhX
m/bHkU+FSWZ09ryFd3pyYT3YtiM71LNZrBg9DLVeutBnbcP/floIqj5Ei/kbO5r0LgDP+O/l+9JN
dEwiXujWXt3Pv4mXPltXTUTYfU5nRYVQW+x/Al9BY1VwxoglOibEbBYOiPhDt3VLm2lrFeUuK4D7
jT6SWgQXTAeO+RHqoV3pTcA6cuAOjhTrR1tFXCy2NZQAakDIDrssfvUeQ19RAsQ4BtyMiy8I9kG0
IfTLAHECYVywzgg2Cs59NW7+VcKJESqhtUZCt99S0tjWW8rTx29RGf/LTCTa/fVTnbxODDLciG3V
e2/ITUlwLAHFSLnn4r6q9yMLdFP9DXg3GtyKmOxRR0gB/aP0Wf0RVrxecRJ4URAxQi4vbClfs4sU
zcy7U2VcaYisfS+3la7IYQ4XzZJsV7s54ylD/knEmt854IZV6bTJDGuEL9oTkB3cgl+/n8PztYeT
fQLHijTYDmzok6lFe79LWmIzqWJGAVzQtP1TryzDdgY4NYUqtnrfrB4+61uKP3GgKKmOnGyO4fmL
rV5OuWQQnssMSSYVxbx0hkNzWy0ffq/F9wlJ5fivQfwlVVtudK7sVRmrDkSbXrW43sjLb1MSvAch
tXoo0kcdhxNGVRdRiwJgYzl4pGTafqA4LEkhI5sNyPH0C8rNMCERh3HoXsYZuz0olTSPrIfk/E6z
5GYI8z8rv0kxXOX7+Z/ssFAgFlzuEQ+2g0TSDfFDIaMe3o6Ing/UT0MBu5B9ClpzSJHBgsRMgsBn
/U8OXFBS7dcn7gx6JidWUIxbpKUMkP6S715URcOwwwG/prPH9RPgbHTrqXWIWIrZotridyN/vzAc
CLLHQTFOpfolieV+mmtREOLXmXjVsdXFtEl+4Va5EAN+0Mr8LIk2/gfIe2WrbI6m2BmFFkTe8Ntd
25bB2U0GhAPe0ue5/l5+mXfjCP7nJOmvbwWqz2VB7shUuhnBHY9m3Uq14kMRr2YYLa0BTEwf7Tya
bOtiOLTLqhAyQTgdtFZhN/Ty5qsudFRA9D1A5VzR8b/gD0S1kOVJdPlEA21fN0zzs04gY9KyX1hT
s+cGdQxHIEwgHuvHidv0RvqUi+vZzOTguCi5fd5d38qFOY6sPUoxSJoQC7R2D9O2BRA+WDfJRLxL
aFELEBdDCJdNvbhhy/9yumgQeASQKOjHNg35DSa0STjDMleKxy+jp9DbviEbTTqk+GolZua3Ze4N
yUPCd/fD+x2h2tSxXKv89Fdm3LATMKTlFwPFkahiQbI22ILlT8LBe6Qt9XiGZwSSjdScTRFczyJG
Pxs0HdGdIML2sWukoaE9N7Jis+j+sFGPnIohC0EDYMQakYvmfinZ8HaAIt4fVMquFvRiwW2T4hC9
n8rtxB38Ss51yTJ3ubWjr8MyoEuMBF97QUZ6pViMXZgPP4mhCi/7ZwXUNA0SthzRgYaNXYaIjYmM
5yBzuFe4ITy+rp79VTWml5vL8qNqQiSbHDIeABQnLbSP3d2P/r0DREvaZSVOUm2ig0DfNNIsA9+r
/fVwDiyqTPnbZEDfD+hWQqZlT5kZXiTGFTTJj37IXj75xOZCM9b5COiuabl3isaR4EjZZcctrtz0
df6E+HVPN45GW+oSzY6kExchvfghhfA9bc5Crvfjys7+cZ3irA+xbUwf7L9K2EbWULkuDRpDMG2I
xcjVf1+j9zUphyiicsm7iFyqhSaZocovO0Hi/WO3EM8OGWubgUTQ9Sr9qh80F8NIWZKrwQzETnXA
MAifPHmQh2x4bAoSvmo3rl/Eai3+1/7xY4VRDdiqOsMUylM3y06YbKQfwAMP0jR/B73DUWWFuFyl
4XvUku+KTjGkhomLyzOZa7xn9zFStZbB4+NsURKgYQhUWgsQC9htihNkqroqV1msmGHpV1o4a45+
vQCYbTjEnkMF1LI61SExfG7+Uvn+HlgPYvqGByt0zGsg9pe4b5kI6NpMQcLwJcnfTn2og1baf+9t
MyTUbDbdrLHU6KVhwl1gxyP3TmqSX642QQTuweftiDCjbqW5zFMFnbxdlxdxdZX7gE5nFIQ+5R6E
OwWeOftgWlxcaN8zNINfbJ+GL5JWBOEQLMUmd/EF2wfsMaSUVExLUP7z79zS0jxxldn1NV52p83x
ZqXl8aGFqnMRvSC1oc1prBXHt8mVIBN+JOIZQ/SkXMDCIDg/K9B73a6qbkB2Rawrq2FYCgaNTEg6
2k9W75iEIPLV6QROYDh5cj3vABUuvUYfICFT0Nxh4qMuGAYKqg4vVqxf5zqoNtoznj3odQVvhczk
j3I61Bcvy8MAQsKRQpjAWV6em15/MMEy+oP4qX5jKOJSnbaR741wVkzVS9zXa67S9bz84vtkvhSO
FzD0hjDSzK7LTBP2qcDpJhPpCJGizN+vvGKWhho7oaTL9XLdk9uufKIXhszHzM/sxEJyMNQcsL94
fmBcgfxD+uCfbKMnpO88XRR29/BNxDHfPwmak3VCrCpwIqglrBZORN/U7PgH3L/ftU7i3LfZ6tLi
5AdSZZSOZiYpMUU6zl3Ul7FpDHARNHRQo+YxAF/nJZlOm/aWBqOZzOPmaKqralkTil0GVYUFxIsD
Hnlql2gi5izrMOvkj/N12zBwP3H5Q0NBbbkrr/X2sKh5/mR+1oDa9ZSogCU7JeUU+VVxQcMuH++O
W4ByhHPm6gAhfp7h510FonUx33vBMjEJznVMUj9Xi8lZWOEs6hcpNgu6LKPaimWeW+ts+OvsKu+W
ALkXDECVfZFbyYHOSqFHbp4FsSlBdiAAnp+JQ6GDI/CxkiC2lGob3TaI93SF+Cj4bDSY44RDR7FB
5gUrWRuJPu431qxnzpWAiAlyL7HXQpBCh/vigRH69xzQkqqKHQivsT9C+1uJ1jQ5dXqCBMWMbb6y
H8MiPxNQmhDGaQDnnrj8Xxs1B+VRxz6wUscz/W4wFRhJkZFEfn9s2UzhvrwW5iTUwSyuiTxgioCt
s5c+JnFjEjLvLT/jPGR5mU+0t0U1PRTS7ZTn31Q9pCAouAAAtcubWzlGi/aiUna/JuQjMMkagqM1
Itiv4pIskNqlXJ/dzr3+SDqPP3AaU+JL0spq2ic5qjWJp3IEj+sNMl9mfeKL+IsCg7GT1ibaJzcr
CXFC/VJN0TndZJ0EujrbmtFhT6fv3MakhLXmRkw3vqJ2NvSFUJDNMyVe2u8m+Dcjfu0BTCBsu+KC
V6FbIu2QZzRCVNeRiToA4PHXhEsqHwgbIjEumlBh1QhBKmKygFbylUCi781HG6SRGlj2o0dYNBDc
IhqU4aWKKJsM6+Lsga7za86yKy27417tIThfiBKGo+h0R+a9RW+inLP3tvKBYORWQSVVDI0M11aY
U03PvvTXpL+vKBF0TLbDIFb2yt5UWy259NRr1nWXPD0IKgLDchkwxt+NV8foEB8fSViNCWXhpQ/V
7GdrrPvibAGpEkz9bj1BOH9hz6rsLYy2BjXMYfCflRhSytXGPXLqfvK2WLNLx0Ny0Iz0kVowZOKL
cg1FwP8Ln3fHBe4Pxp9Nd3kVyb8Z7OYthXvHvPAXU7fL79021tpXapxUUSdTx3atY18X8e2ts8zI
A1g6Px+gF+62UDg9StUWw5jzVoy89grUbqgAqXHCFnRtJQ8mb9yID+VV4tyygqnyRQg8ZJMqC20l
FuuXzkFrK337ksdHI+2st2TWgrRUnb5zXN5c+a5JHFZKImFIdpHg0qE4m/jGkOnoH0EO6l8LvD0P
K9YL9iFocNc4YFJWtccZGwgx9/652OLKGG4jA0rZQUJnUuUuI/hBToz1pjaDGIbtm1O9qL9Plb2W
2jYBN7PKmZzxq1vRvuvysLdLG1Rf5n2xKwIe8AfV2JSMw4TisXgjXeBijjytxFHOTU/Z4KOln2UC
Fx2rl+03DDv9Wkl1cOc2hl9ubDaRDP4rGrRavOlPOTx5Hd5QA4XNHxTJu6XAY6gtCtkvJSmLntIc
hbgtCkx25R5MrvEGn58vrm65g2Ods7DWq008+lU9K1y0C+rkSN1XHrTDWgRdm8Pc0AW+rQzgyqUO
YoJEHFOuJW0ysWQnMY2iwNKlXQW2f9gkbyPKASojxekC6lbKyTkGTyP9LEgey+yG/9rzs6ronwpF
rCpjOwOeq3P5+kvrVl4A8pdqiE+0xOce5C2SsAzZHolWZOok2Mv9dcDj4SAroEd5JwAIteuutUAX
I6BAb9AILPG9az9JPB0VvXTwdrD4VwHyACV099tlgrPxcmvB586AxR0TQWcU8xMEaC6IE3hovN/G
qRKHoSByt5nW0T3dV6FStjCPAinWH9kmK9GLb3OiQRTxRr5f3swGqaRZspMQ1PC1yB8JrzPJPDYh
hBYpAX5/U3nWgmbxKyIkDlAHgc9E/E0QmMC/bX6p5xSDB9nxAbhiEks0yfUTURqqMhg+DfC/3SzW
+L/uaNiNZwYTY3NNh3iBgG3DA9ZzOGZCTDpyPNBpQ3zvA6c81QSzTUXnt8gN7dG24sUMELxty99g
RLMcXE4vh+/RRlpWlz/YpExEbPesRxoGNazQpaxj1j8od+szfte3b6Ndc3d3zUxQzJTITdc6a0MP
X/ln8JDRTPVTRdBVn73F/hpiRSjs8MIjZh1SABKt3qJP8KmSLFaI+GyjfeyzfS0wPC6od8hhAtV+
Fr+8wI0eywKlRzNZUhTOEzKyCSOSW0R1UsOM28l1c7HiLOqoI+jKUiISMwUYzEAegAgjE/ZVIDKA
iKYVAX4xe+bsdKgyjk+/5AiZydwWe41Q6Txw9PLjsUuGBMdzhUkQPvREmYHMuVKnfHfI6kY3AlZ5
iqY97SZc5mB41LnCYTw3aFO6O+ujgLYIrcmOutMtbGB/dYtcd5zatQ3mrvMYEzP1UwLzfSa+jMKS
BzIBO0Z6D06ULbIQyX87gWQMMoNwycINDMGerJIrwxgyBPOLDqJg5FFKUheqXCSElndjB6qRVXRx
ou1uDbuPTuaihgQOT5V6dLYlrgiOPesrtTDvhHFv+MUD0k+JMcIJHNM2+XJOyGWiziRQryDvQ4cf
kcdtC4BFAn0kVZAXHwgPjG81UT18vZEPGXjHkpjtEZPVxzwZlxyNHMTsnW+u//IraRi+Lr5uJZ6Q
6P9lFwarNikp/Aioj9lSubXcns9zg2PQaryBmIUFZfp1fqHwITB4CatdHU5JHXWbyrX4RWwuBeUq
iQCIXFoLYOMIa+BzfFSWg2A3hDE7PAMQ5ydyMtVHHQZrhLMsXv2uxGSjWYh5/AQut/p3cKOBVU4k
7tYiEQ8QMyXV4I0mLwILNlYwb0t59CJ0XZrjmPZAtMKk86Bz4h/uL2rwIXW8aH0kfh8Pd7CaqITu
I8sbFp5t58YtvLasHt8fW9sh0IdzvM9Y1XlybnPjVhc7JVw/CoB5F32OzjME2vkwuE8mtKLoP9ji
nAEZHp8qOJjkKJCljY+mIzjtSiM1zthmD+tOUxCG+r7HA3cTHvdKW367AbMXSo20myAoUqb+r8Ij
Td8lCgWnVvrDJFk/mWD4v8Q4dhClU4Ir1t0qetY01Cmf2ht7sCC8UA9GtAMk2xyOk/DhPeie5vGY
glhES/0ixOJYpiOMWgGfI4lYw2GXZn+zxoKIAhhC9fXx/XSMfc3nII9tKRnJTYD+716hmb6HJNaW
Ff5HeRPBQB5iX0l1xzz/Hvn7QmrCBjpwAcZMHUBTgBqu32nGSS2nCaSihBsA4hkrhybXDhjQRMXX
zNnR0BOxkrunbQpD7hnj015792+yZJ3UlB4MJFW1u/BgU5v4BZeRTMunsUfst2u8AerKO4jHcqb5
FZ/Lalgel8lizM8T0/6UoiMPYcjew8brDu6Fdb9fM+AWr7fi0eFyiUeOpItWN5qbvJn5wZO92x47
6qURRCc2KWoRV8ppQLy5CIAuNTFITAILqOi1ArPjKaArJ6+nWa6xoJyUf2qX5swlXfFwzA9yjw1W
ir3KCKpp4c471MIpgygWOq9rDgsccOuwC0DoobwsR/m6sPn29cKtN/SXvu4RVIFboLwS5uOKS6K8
QC8UpCASjXDEUgrOoscm1VVMbJalsFI5M3xZqRpMZ0HvizlrRPOmbYJnCTi2DyQpvNmMU8h6wlaP
Q5+lSWLF3nYnA+pt5RRk3bO1/ixIvsTwUPaZ0ujlAAYcYDRBF3MggFpHDnAwcr+lkURjSd7G5M4C
CtjH1QvNhIrPKAi6G+0m+/ft4BUNV6hYF9ee2bYTF7dfu1rMvkl8Z9L4QlhZcC/iHlcE+698UMwZ
CetGVVshc17Ge7imuxzq/ad/eVRWTX74fjQS0tAp7WBQqa9shpTZUflGNgwOzsS7Tzmci7ebgQEr
4g0TjVcd4krxiDBWjfWUivCB1tdodrgiD6h/KDmsXJdTjRfDx098J9uC8LyNVd/HLZ9owDfkfCCk
A4k7Wk7ulyKtkqEBeQ8PH4/5FW6KXc/zv1x7etPoSKBr184Z/SQfLT9fU4kkuWOQfupVF3qKZXZl
A7J1JnXu7SX/dZG2lHFQyR6R2fqOnMcrgWikO23CjP5yjIl+NB3oNm1I5U0mx3DW1DFjyEC1+N5E
oDukjBIMR+fTjTveSczk713ZkakcXCLaCxNGcawmrbzarF5xiYH93ULk4vk9UCx+9LjN6FcgAW4f
Xs/gyJUWzzsEctj3vvNSRpmGiQrMrLefrFNthDKnr4bzKjE7BA6HfAUNhfU9cgM2feDyL26JDHCV
S7t8dlfn9CfJQdMr3Aq3fS5DB4WaGubt/3jqGNkz5sxk6jhALsHxKNTovU4i+wTMjTRdOUAFzLxf
ini5qOCkbVT5vm3g2pbmq8FsU3YFyMdAN9Gql1B7Qy2H4iq4TwMxMOpIaVGZipGlMB777GH5VKlY
IpyMaqvpDH0sZEzMuEbpLFCXsn3xv6Y7dDxk01W4GE9TwzDbjO+HbmILArbpJMaZX2ozZpEovTJp
8EOmjDUf2VvivTmtpe8RWm+efp8rKD/jKbjuaDpDT4e/BAqSCIxzzuKRJnCs1ZVZYTOgZr7BFMWZ
7ctCjUw/yGnZgJYuA6N/WDje7CpF6lT63Xw3v5I59hFwm+d/QbQnt8sRlvKgpywK7glKChgjWJwe
m+UfFLOHLlu3a9HwLT57hy9xEZmM8dJydYr9/rD59jp+5cIjFoO5A/fW/XGouOkpEDaiLk8fnebU
fMTgKwXgcALRZGygTQGBCtOSbsk+EQrkpJMRhbsMJHI2DSp9AO8RIZf9RwftjoYjkHu5XoTcPc2s
MJpQDLq/Www9NZwBQYrHJ+luqDnJzHjFgTzRe1TXEGWI5VBIbwDZhb+cWkzN4N9Ul77ZWU6nlYqJ
I+HRvYN9cJE82Q+1yXIsvTrLnEcHdYyoo8u+H6dl7v/nEz2TfLasw81C2QVMlegmkT9YxqNhMf7p
BIGQ9r5gpVDmzd2HSVBJZ3X0f4M882wmVYTJvGiEbokJmOyG5Ou0ALZy4kzBUg+JxLI2lZ6fOzP+
OtutHvYlKNiF4Nl6qOcq1CLqSC3gLJZEOMLtWvt8nhOum0jEqYpkZgYizaGTViPgNjRFQ85p21dC
cq7c4DRGz5SQNlbUxHvdQcdPyJGsTpIxinqfcawS+YEaGzUqkPe7OrzU8LTV0YG3+rmsF/6M3SZz
E7CCuGSbOP9guujZ2mBcWadnvCTYvYhcPntnDM4eYc+iwl015K3cQGMrepTrRhXRlQvqAKNLqg+/
EBm6DZETwO/CbOPfujq6g/hkTV6C1BB/BA/s2htFqUZl4ZrUGhn+zSORRaNfyoT2y7K+3qMW7fk/
rYkN/L5rI3sqUFH7S7Gohc5+yI84F5JCBoM08tGqbbi7E6iMhZD3JF6eDv1sKQ+mZaKcs2IH1jEr
c0Jt5YLHxFI9LZD3VG/lKVk/13eN9MluFSu+xvm/+h4ZETcqjlcsLM4lFkX+NhUej46FAX9mlaxK
gyoDp2//icvggXweJqd2jRbvsiJSXaHGTyAP3mucVQwtv3dXezX2blvh2j8DkGJ2Xe7rE4ndQH0l
8m7s16k2SeEYYUG4RxlAHxt6R88Auq7NpC9EBzyLjbBGOps4dxQc41yovym1zoFyIKDTFxO+JvC2
76g/WNGgxzwe7Cl1QQQ+MYy+PHBrS8jElw3gGpHuOaLMoaCT88nNSrDGv5C6hX4dlK0p0w1e+nKQ
VRTnLHh/X+68BAgTUpW1DVHfcbnI3ibvKsc8K+e4yQU5XVM3VZ7X5muhw/MGWxQbv/wV0vm6ji1C
kxhMvxqCwvU6KvPWEXlUYr/LyC55nxd1XMT8zqCrILdUulPVIgRsg4cFS1jaOLXBFLFnLTnM7TV1
DksFERomkS37KpNSxsz4QzfnIQxmHC6D77xXpa4e90ZaMu+iSkh4DPVVJabKsSi+GKneGWkggiag
ohKQzW4+LQ0x3q6rkGW9Nuoqe3626dWXLg4DCD/7wJpzIU8HdQnYZs2v3vnGbsxhVgkYetts8PRA
rHn1fts9UZsyIb5sN5CXznxDePLsI0Y1LV//AahX+Bby3uMKM3o0kyTwpctu3J5dCqc2nJtzu27a
BpD9iNeUOqdZfBW2vfVnDmLpPY5aesq9aqDKWbohTCkHAzIY9bP97ZfSnQXf64DqWYhUcQV/qJ5X
7XoEQ/rm2YJbLJWm0bAQRsh0YgBgjuRbwAkn66GfWsIwOKZ4iZD/krWLlJLc+CcvoIxLJavrNKlK
yrW6cJXY6MZ+Vn7BYkykyENHsdHGLOWwHmtoSvp/mXo6rgXXpqsA+q5ecJLXZ+5zaEVBc7mI8AkD
ygp1egz+sAaZXK5V5K3WqAVxvaVFNPKvnNEKKot6LER9GwNUsm6n3xVTwGMFLKXK6GfUE3DwL+FQ
IoGcJHsVd5jUA/HIoh31Ge3JAeoybbulRt0/WF0LQuJgs8t34g395+4VS/xbrgcse09TWUVCuQkx
aWmjrM5UgNB3bNCxrxcSZhmnmGS8YQvXCmdybkOEEk2XRcaRKRFbJ4MyCgDTOyXHveM22zkd735q
QA41gx6+lq3fDIU2ZGULKlbsn4yDw7zCe+GPE1fEcEjH9bpMOJ0egIBhV4xYXh0ev32aBJlBMe9v
ve20hyHVdNWXHD1ghHwsimc8jmAVBIXBx7LsxtCxf5e3CXeHRFYusOajh0lrzS6dZ1mOJBbY4JB5
OCTXObSN/sle19a9syAQ5Wed9QlTD/cRvyTXwdcfE32HHeNe20nlYpUJu4JPon5eR5DE51KBc4/w
vC5NdYVeRr9+jrPHdi92MWSpvNhVx0VlJuZHlYJdIcQteBThWgbHrhpaNcndRrZt4IlebXBacMMp
ZUt5yjs9eeXeTMfAs5xAL5KOAcBPpXMW3JcvaqAkASEBpVTqypLgwUBwrljDJSrZDqlsKzzu76K/
hbnLvY0S9rsu35e1QIm9FJmZcNFEBOaRpXbrDHeWggP44+ljbDf8xViW6o3KntafCOsvlNtUdOrY
p2mSwOCC9f/sO5b67GZfYbxJc2WvhkAgkV2nAoCqaa2wBYF/tKVmr3sN3oKtGOoe+SKjoK2nIH6p
8B0+HsyV6bHtH7Bw1hmwD9J+WI1ioLDq2UrRbnNuLtFdoYXp60RHpGzfZ9F7fYSVbCuE56UQO7R0
ZZEkGxWgKH6Q8h5sCKujEms6X8ufVgfUW6Dg8CL4Zu0bN53OTXQNIRtW6aEuC8lQaZDSuiiCftYi
9bcW5PTQ7AkCdAlu1B7xpmcUMlTW+MKlo9DpaQjTjizyFi5kBgbtoXRii2kTfk1Pd1963Yg67Kc0
33PhFMxWyn/rdvpBTBTBOHaTgynbKCvm1wmhoB6lxo9QKE0e3zH3qF0Fy88CcjsbvvMb7CyPD/SP
Iph4PsvMyPf8hZVRDS4TEYm+FKCQNzp9ThngJsPfHkJl2SwawHD5Mjs8uzLnoDIzV8O90goKnMc0
GQaCH8PTpuE2t3fuTsJFGsWcMpGmi+gnkSiDIarPgS3FBiSEDvIXtuYOAggxQ9MYcO9K7Xn/ruxX
HjVU5y7i9ety/z9e/DvO4pnYD9QKYt6FUFfMwzx3xIkNTZgW0zRIrz5JJJ01h3BawqayXVbJelue
pPkJxyg5TLtzGWli51vhRnAjK8ckwezLDxlCg/dGJaEN+HqCZxsFwnNkbOYh9AAs4uStzHu/MISb
F4TWOynq5TxkG9s2Muz1BaIgF8F60QZ11HtQQ79h8tUYRtKve2WM1/VirGwXaoK8iYp/LNWiaNnG
bQ+azwx+yBZ/fVXXah9E5ozzDhs2y3E0MkObTBj7fFYT6GfnmCKo2F4p6D/NAcOY/uB/Ii6bSlG7
ju/NtUqbPSC9gwrtKmaEIdllYttDMZzsldEmUbIUsOdaed8uq2gQ6geQjKPBSDYokdfkBH6yi4tk
chdjhHR0C6h/1S3w87zgcQ5ZR9NHnih/82NWnVn1ffA6tggSKNKkZPNfpzSCSkIQ5V9UibaT6BhP
jcP2QS8v1pYvq9TJGUKSTKTHlriyziWpGbYMNM45BOtx/CU2Ng+tMW4NzQzxmxmzfI7dt+9YDtyP
B4FBvgxMdLwjtGWhqZbtqWampKj6wt+NuBlhxoZeUz3UvkS5QuW5rgUGQ5s9T8SPcHuoP5sBoo6y
+gUc/wP9Y5/fuEioU/wmmpImGZtQEi4lyS89wTAlxhizpe3kxL8XEkUaXXYSFR1epOGUsPB+Cg0D
C+YfHflpHYFbCVRehGLGl+Od9PTqmeKGuXHnKrxaxHVO6mP1jjCwm/rLawaMbGDDKdi4aTt2VJ51
YLOBuCak0OYF7Qr3ldRPu1UImSaiPblZ/I+Xp2JANiW7x2ilr1I4LC3FEN4pjdbMLoXaBSBfUBk2
NpwNhTgTU7UJM2vLP/wlEMJN5DubqUBdHxjjlLnzZzdAi2ZWpJMFZTkdZXoVqTeYpaGRnSdtC/DD
/MmQF8SeO7OfwXnlZ3ue2HbCvI5zUd+Pag4g4wPop6TmAoKlqf067WMi4zv/75D/UA751jOmzrdr
fHltvPcB/4V1ddnNTaNdsx6fPMuwo3S1BxjJkLOMQqAHC94IR3Bvg+cQtNjtRo1Y9MFwc0ovKSbF
cJogYupcDmSmJ1RC2FDKAVw7MyzfxLIUQsWUD3gqbTLu5ChGz1XvZXkAbURyDjzfC4VAKrOhgwcA
dkGYq1ZDiNmhCFGpzGiRExoTpYz95HeRrqPr619vVSRjJ4bjduQoP9rKJSCpQ9tBzeI3nfjSYgva
eh4ekXN4FRvnkso/dTLbT8cpYPEu1wgwgrTzx8QJFqNB1/sKBCp7ZqublIEf+uUZwSoNHdU3tPaT
mee5NR7w+00CybKNIH7Ts38MdXtfYfkkrLuOjGDlpwODFUBEKWvMPQiJsuz1/o/F2d1M09T/dSye
2hucGsZYcJCxgeyS+1YeinFJtmfm9PlhaQuNGwP19QQhLEmnrJguPEdz7CjWqBpcYY6RqkR5t/fv
fUO7e/lxu8GLNok9zXg8JrZpEltcvdrxBg7Q7IBtW/5DN/wFglO5VXpW9VJk62KnG/Hq7Isfilvw
CFupq1e2gUUgfcAH90y9WfIsPBjt+IVDksddhLbs6yh6pX4cQGHgWfVmjw7dFI0a3Q/HG11fSoZr
y3DU5W0v4QWTOpzHd985nYzjiOvapT8OkRZnsVq/Yq2QdMal9hxh/Y7JH4L6sP2AgV8WgWTkbpTm
ElwRVc9c9DUFwShC3MQFHBenXJvbVcT7Dn3d2MN2iwRaZulJfvew1asU34EOrpEZV4jUy6Tc5vUZ
CAcgqUSwQ3p31oKm6OQJdyhGwiG3j1s1xEWVBTKKx6Mdd6SNAgTq5J4OmR11wHMGYtm9KgV4Vb21
NIyCwvf6JYww+srYhPZrOiZoZimUh6RJsxpOT1+OsIrCYVEHSSVc3aI63yqNGjLx/Zne8DeGWqFQ
pfFc35OmHw1rjCrD97J3aiO6rvitszGDbZobQfZSRpw/W5Bv4PGmg1F4J4P/WEQ0A730nZzK9e88
mqk3TRshnkJEP93ObAgB1zxhA9Y8llW29dNJl+OVzqHUpib5wd3gqISG7MYM2Kk3bpq0voPUwo6C
mxBSbSYllQQVKQQFkut/sTreJc9sX5eqvyj4i4OgdCEuWmdvdGmJ+JuMMaOn4AdMlRl/V+RMyqgG
PoTTyIiGuZGk/UQjloatd2vcoiy8cCCn1WgQ+NNdyzVlEgOchWWH/Bhq8iML0/20dwzyfhYnIb1/
EqChnk+IOZGqcXQkd2SFvSN2FUQjvUFFzfKy+59c6RUk5KafZFHQT0KGygBhoLkadXhaFO8NTNX/
WfpCb3A73j4qBsdqbtn9D97HPrzsbnjAc2WrqFQVLBNgtT5/NqpOhSFfB5YD+9zZAwzBahL7xWe/
8bqPjW1BBsz1zyorG5/n/O1T0AVlUon14BWw85AmdK262RWWWlay5FjW6MtivZCsB0zivu/JLBgm
eJgMUbgSAylsfBZohjX0UBpbc0QgLraOJ2Vs1xCV9yHsZPgbKD26Vi+DoxUw76Gjtsyk6NBMJddx
Kl+ABiBm1++TnISX4PIk095F7zn3FN4I4DBMExLI2uX0t84ZaymaGPve0zEdUmoJ1Jzacm+h5PBx
fwwm8fR0Pz4dp8wFWtJUmr6oSVWkR/fr3MEIZhOzRNLvBQCa+Sg3TefrSCNgFhtntvIojw6IR9By
CzKZ5p5l81THWRqawPH2c7lM670UE3ei+a58NiSNnNApgV2nGufPBAUAO2ls2twSSjFd2NgXMqU8
wyWMJGqtCLcFrqkvr6RbsBYFw5NgtwxCtE0wTx9MtObdA4VtayBjgWZikYgIg/+ouCbCfjak5L4n
b9YHyCoPlJR7MJdxehjDEqnQvVIJcgcnA2D9tuKg3svLcU2ry7YapuBtMsl31Rho0zDcCZhiUktp
cUfmqkHA8KjiWOI+hA+ayAlW5COuw8NesqR4tz4NLXlgf8kq09iuEYQ+e61T7ZbnSK+8jqTRAfUa
HeJr/WAZwRaQAW9ExuPIRs2fQGrEmppf5uygu166Jq63Y0bttMaIpwQX5tR9v8bmZq2PHbgMDhmx
dshtKyx+eT4l6M1LJ/umGJKEE3AReS37jFmmG1LVNIZcHCr6QZF8octXyUktUf3FlkbShu13b7hB
KHFxKmNZ6zK+6SVyR3V+UK3UCYnXzBqTq/iM0evICnOtD86362s3hE6ryWLbSqNElhpS/RKopphH
TdRJyLgtfYBzZL+EyloGUGODQAoyvl96YZUZCgrbx/0D7ouiqJomP8wC8r6/5kwqVPK6S36MGfoe
2eMikCIlHAf2H1QBseE6sQCtXhXVbcWUAMcLMUMHcOAYQbQc0+TUscK74qK0XDSbTvRR5uzp3sCn
xHp0WRnGGn3MwkfZ4EkSayuWlqOmEiweepWfePwhAZWKSA+iQW8FShGigY1EmugxMozgaqY6o+dl
V5W08vbI9vLBmLzi6z+DBDB78yvK+cvmZAL+P3gy+Er1FH77xG2R8+cImBKkLi15VjJxlmPXW0R7
Cy7ECP1+nC9ysEt0EAcZ4aab3t5wmHJA+gLchwIibZECJTcyJJVV//or+Jq0GCmT1lYnG72tr7xV
CoeFh0e1bCf/4uRscomptk7CGUL5DnX+faq9xqNyqyDeiofuNsIbNCrdwmUskqBwKt93mynU7GiX
U2LVe71OEq8GYvPSAQBsifXyJju3NWTg5znZ3RVtBqTFHacNyRkRp72ODtFuwkE9x5Ubv+6g3bzd
AF0sKHAMbLRhFh+PbQ6Y8Yq6EJiZd/jyQ06sORbd+QsZWaFazOQiHr9Bt9f9sa/VWIwKBVwLMhCd
yTk+ajHWXQZDmjbEfr3dGQhyXxTDFHXQYtyfgGuO/L13i2KSHQiPX4wVjGprDyQ252B4SdY/dMsa
1o8au/prV3DLziTz+1tcMSmymR1ZwA1MzdHduYVLxG8kqHDBBACCzHBmVLP80zObxd0QFI2yXA77
x+KkziPyiCtCS+32iVUQqrHhw2/W0bjeI6aKLa2ORysNfu6x6BLylICL96EC+b61TtPSpp/tSymJ
wME9HHOXwASRgttjf+o9O6k3b28yZ97OdCGhp+J+v3UjA9YkzDJLDhnAlQJzpDhIQIe+fZAML54x
a1T5xUNHLH+wdat/ZsWju3j3Cg0Q3quvsf8h4Wum+pUBxXehfADZVLZs+0zbW+vHOkDrhUjQy68i
1a9L95MUjCrKMxSStJjABy2EuYg1p6fXMiB3ckBDZmmNlK1WagbxFBWqnHEAgbPzcqQMu2p2kniI
OqfWi+FKnU+cYL9wRUzV7UGaMZZhWb9UYNy5+/64lvAAx0+VVV5BML6uqnmTR6+BvBYEbIyexkzZ
n6+LhXb2mAS1JX1NyaxV0TAK5TVv9xflNomEETEghTNL8XnOwUBKNThz0gpMW9GSzchzDfXWZCNW
QfD80DEE7j/zWrRA7115r05KPhibuxwRMDUWAdQ4A+878Z1460nH1B97eieUYoLIl/qtypZlZI1X
jLBjv3Olw2eFRnwvoJJI451IAxnRJn6dVJjoIMj7jsI6UYOl5aCmmE53QHnGwJ8xt1d0lRqU8XbG
kWzSkabBCucxBtm8BB0cpXtax/cJ/NmEboml+DyhkrwhNtcuFEWY2Aj1qMA08KiLSinZUJzRxWab
60/QrDJ8Im/szKTOC/VtHSSbXhRGQBNKuc2g5nDay06+5gX9kQin3mdulV2z/Xd57YeVYgfxAh2R
eBFTvXO5Y+JBl+mVUUTIjo+SSZ0bn0rWDlsuNhOuDYgjC5JsIWE5FERJbALesFgbSw01wQiTO8zf
tbUuHzYV6dt9Unx7aGfKq0IepDbXWpa9R7UhcPW5t1h0yoDfXbPnoFiqDIINSKxn4MtobvjdWAyH
tdYiz+3Zw50wHGenEk84u3GrPgFqWmdTH/svqgqYApczqwSKUom63g3lJekkZtU36I9/3O4zkybs
aGdgfOVdlhFxssx+HAcZy2jOYuJ13xLiYY1g+4I+ta/hjJdwlzCZh0RAKMrGAYH5GNf3GfRgatkQ
TO2Lq5aW75RuPxdDS/dXpe9Jc2daL6Lhi7IFqoOtOdMqa7uJ5OryIDhXW1AmMwb3JBeK9BOVrHgh
PsMUmywrsNVB6trc9jJuQSeqUbP/IPYZikfBCRFgTQykqaPAEPGHt8YmpMEzuZcl3RZPtMimKsT1
/JuHxBuV4JZU9LghW4p3UU20kA8RFb9EVG04uqXrnPyoCCguepZ1RGfzKoWRBcxRtDuTjZ66PbyC
OTaE2c1yb7qryjPdGA49UEAxOF4vfUnSTyA7fycZgW/QaYVeHCKe1y41mVj4RZ/zyy+bF1Rn0gQz
UbuOhocY6zNljI4+QI2D5oIZpExqEp6pUiyJle7zENPQ67uyqASC41EgXONKMo+leEex51yf1QjH
DC/sI4P7ylF9HyBoUGva9LLbbEw/9pL+qZHeazGPyYEMKjTbALujlUMpB9s8bKGuseq0b7tun2UB
br9Dr7EQvJkLKFJdNaiY+pQHwfRvENU8nvATGJ0+VfyOS2w5rAB5GClQ1uq/Swn9Y/vPmMyIe93C
aIOwCSIZwWOO9ZJl6gL3HUSm0++/NIzAUghRFiPSo3GpaITiKsCFiv63WyA8KFjbrDMC0DqS9Rhp
4kV7Zj6SjqQX53WMMA0nubxZASrMGXscm0hdjTVEaxqqi7lEckjOEbRlk2Cn6LwsF8+2ophbZ69A
KRCGdRD1zpY4W3dXd0AFY/yKxvmIdr4sv1TVHnzf0TSjWSK+x5WVa1QrTjq64kf9m/Iktll0F8VT
VZPaFFu6oVqT9pjY868KCaBxXJDXf5a5qZpPUkiosrNIX11etfvhOc987p5J7ybMujTWCI5tR7KD
P8aZ/cRoUvC6dcTxbVJrrtIqWl3rAU/7dkH9TrBnH8lvq/nO0R4sq0XoU1W0VBoRBnnU1luxvM4X
AbMHyVawJDh3V8zACygGJxLM6sYObaL6nsoE0BMw6ei1Qtd9Vk21Ui3Yb6MzcHhEjjUD20MrbIZW
QQRwP6omosI3vmc74OxzBPiuqsmodhCCduJD6wUyOATDKQR9XI5F+a8L+eAlFAEUHFgnOmbWBxRM
YzmAKUkfmyT6Ppd43FsXCWSr6WMxxmb7sHQIt1r9oaSthi/D6Uh2OJdews9GruYdqzkcJYJrYksG
ImgQ2GP+LUL0ac84yw6e7uZXwOxgNk65smbRCgRzB4n3NCdoM16G8EBVGHbvvom91fC7sKhbDcVI
heCAfLQc77nR9xuFuDptZ5P+tvGgydSk9LOzZEi+/kI2zH9cZri2GhMzA5Xn+cKNOOdfzMHjXeDQ
UogvXC7T/6EGjKGmii/lAIu+2ivkNayp8y1/0DAWlYyTn4meMtcNAhCFADOqLFzjlOv8Qo0hEtmY
+hrrtjcX864tWh8IblP7T0qt6CAN7TrAzXntwKRsDIFYVbSj2F4dhSUrYFZFXmMVnlExCAk8A21Q
iiaEI+nXyumx2DdS3pXi34K6Kq/TpCkxjT053aE4j0O7BOLnu7alTm6TJ1MmJH6L3pBfqPEmLmk5
3qVtJs3P5MpHuqJMTelbjKCqqPjHu2zaDVd5/QMrhes3bIsEhJcDfq66J6MdvsqJCkt+CcZ2lARY
eL4KyJzxBWb+8wjHeauvKvIUzVQmTrRb4G/oJDleitw8H0EIaVwGrxdaaOCGqIOP9d4eXsKZ7BBx
FFzWN+Ab7xBLcQDnBiUtilidB4qzkp27JnMigZmAxvUvQZz5Y1q+KTJto7tdHTmpSTMRPrlMIefB
3morDd1u6TpO2sp0/LInN7vXLopINGLlU8QLTMyHsXdHVgUrOGqinDC5u3+yNvY3jDHXduuI+ow1
RsAp34yJKP6v6ZR1+l/KdRFdWVAxwb9M366SA3OcNO7GGALqtNxulR2CQk84rDEpTWP2poRxgONU
d7Ub/FO1e0DjRutf68X7vEpnDVGLHt6Dq+ZZg2PaKeXEA9ImYNPKKdEhB8xwpnMCbLbEKKK1GfOy
66dMugxN7ABfio7co3r76ao6G9EvPMXg/CkpiS31SxhZVN3m8kMqBxtM3bCwTg+m/UYZZ7zRkZ24
4tF1444LF9QiPYafn74zK/dG6pMrftYXkEsn7jMXbD9fpl+WV9hhOx94NZPcJkrdOil5ZE0XW7LG
DemBQmRPVyN/T8EmbS1ILZYCG3Tuqdz9R4z5GWbiHmn9OqMWoqfgJFzeOIiNEL4u+ClvNXuRXuKU
idz44G3icuVzJkN3dqlnealu47vsFdbcqWk3/2SN8g83EaVgTY6DGGKX0Eio5GzTKg3/pEUJ23xA
FPduyU0bugYUIzUfU5/uFPFUHlY/zv4tRum6zAAlt5InuduMr8Iy4125wxSBeGf0VrGSXXsIuYGT
q2XagGk7V7EGLYwvx61BI4Wc9xRyO+ToSWXvLpeNG3EJF4oZ//hvPRiQelUeF/QTIpzQRCulrNQS
jfrZRv2bGsQWt7CEMtMdnhNGZdmWbxdyRk2VV1UIGsN1ftxhyyg/+AnP7Pxzv3g+hEsAWml8rUKU
IWSKpvInPWhCWX90QGnbF/96izzjkp9SQzCUKFDdYWzenJbrRqRoK5+B5B3f+pZJoIiP8Icvxg53
Hc1FDPmRxrAOzeYiczHw1iMsD86Hz6iCYkzQa9UMV9MjEwBLT23LH80GnZZEqkE3HVvr7nNi2Xrb
8N4VVq4iQ0V4mieaQj6CEooBIs+ArtOp7lAlfZMam0pNH7RtTqabHKZYmRa0g+642nZMxGx80zkb
k+tQqWen62r8OtUEtf3Z0HpGJlSiJcL/SxCsj2cDhSkVvt7DxCBRLPndMlOQ1kzTYFf2eT1p2GBV
Z7VgtcYG2D7CnPvIgB/WFzXO/P7hTNYv3NJgKymljMeJdpulmqlyy+Pk6tGVEkGUVxK2qfiHL8Es
qLsuF+qLELZ3vMwPK7TJzX4L/ZZHzwZrkCtwtW8YaRj3NyTKOlIAVNcuQKOGWc7bQHXtzcSJeOCK
vLkHFuODPfbqRynN/LPIbYved4jwyCRvR/m2VCMIK3w1mBvnYLBgkJK3+BGoH6d7eka7c+3Rd/FC
JH/rspHOF+jsqvNQ6SXc6PSHp1H0sAK63GYQVdtpD0mvr3VXRCDKCbdaoz5Oev7+Q8tdKFHANOoA
WrMgUKZoWXFHsYOS3vAqVvyNW+UNd4s9Sh/u3dLCDJv+pzLNUkElzy9NNxgX/6+eUbFeUoCvHMU5
2zJlF9FRBcR6g9KUaXg2a+iXID3QDvhpEfoWV6HIK4C8VmqhkmnKReDcGgpJnBbLFWLPrY12EWqp
JavW20qEOr5uzV5UP5xy0pPyOaQoSIZ91x3TH1J0nUcSkdNTUNvyJOQP/cPX5jApcBL/RVWgHOxv
jBkiEJhLXZAfD0e/W6RbTlVbMwVCzle+1P10E3NJ3KILcjpmJYd/ux7SKloZPe1yWZHtShEvDGUI
qWuftnR+3kZ1CWQXGZ1Bw9f0Y1W+0L3qV5yT1KOtHYs6IVZFNLn2YCnaLKVB4UK9Xbl5aCe1w5nX
nsmPT/9x60olfiJziD2H8N4k4U97EXYyPp8Z2NUVoIyOIgWOQWmrezzezTP0Jt2OnReTB4hS5K+G
cl35f15GTX3SPOfKlwuGp3W8UEIaNSWq5SXXDvWK+vJrpVasBV0fm22+XVG7YHIwAnwLW7LopyYa
xu+ZmeD5XYKl6Hq5kLHJCbkyZot1k5wVU4Rd9LikBoEhuSQpM82RRU2EeXq36BCdjDygyO/MSiPP
LjT1CWC8owJ6CKT+Y4CROUnVv2p65fEzdf2sZ3Lempe8eQNdOyCYzfRBMOlR698kPUAyedptQp0V
SuwA7mlJ3Ckq2qybUTRsxdresTClx5bl2BMj1i3Ur/1m+THwuXeMfgz13dfYF8OgrLFpGHfXD4ze
qNHgIWveuAmXZY9Dc2d1gYGgXxEl6NGnmWgvKW7/l7RBer9Qxvces+/HuQg2ZW922hepJcPLAJ2L
tkBy/P7FB7VDU/lkpu6FT6T4k3PYLCZy9xeL3z9SxaxFTz7rw96EV212INjDsXBii8OCRUWHSJAJ
ilQ7xVHsyDJTU17bTintJA+gePLWFhFnmres9LABEpctlMESD8kdm0qllp5mXLEqJwTQ1Sj4EF5g
bi/L/BZPzWec19rmJZhoVONW+1QfbhJtPWkcWMi+WMDcOfJsWzS9G4vqnyb9sCsjSOIMl4eBp5hV
zMp2LwP+/BuBPBHIZ5/ePu68+zEp7cclOBnJ5BwyOqRIBHsNR1c0QF8bn7pYWlMbQ/Jj8NuLujIC
yCz0YqEGt19UOSl/B3GmobBqYnkldXhmeBSUWNgIDVO6QNlF5YdMRqPMqELN7sWbCSpwhFA6Z83i
/JUvKmBiU0BaHKm7OlMV/1YtQx7Pc60koPvLxKYSqSmKtVqaguP4T8lzDhuI+yKhJqmni1wcSTHh
cZvjEexrX9DfznL8sk7tDqKhGz8VBJ54co17rkquCJUbvHAnZ+xpRReUrXCcbULPZhndRPkScogT
AR//Z5E6yHDc6MWxevg3clFOcx3ALuQo2FBYA1Hw2ZXpcXR7F5iU6/tLe0bPuHTEgya0aTVT8Se5
wki6YNU0defP/emaS9n15oXfHzbuRgujLhMD92QubXorBMURmUNmMbDLrDD4OQuD5WkJdBwvyEsX
knn6hoS5TYdPyfaI1lPD4GTFTMdR6hvwtitCpJmgzO69sospSFCHBbKJmG4Nsdc7pF/fcBXZOGuS
7RBFw/29l+EZse9fhzT1Kdugi2dYXw/I+ir3BuOk/MrfTUr8+5le15RxZZrbWUymq2KyVUhhEgUV
GAYZI4PjJ7WDEoa3EBbPQNFmGz5vdlCqdNwJrMEQF9BuuHIY9H5u/cGhja/VqAf4ggw7Ww1lsqr4
xChZhjDV2A4gJqQEa5wGnm7kfYcrug0i4zfsQdJPXMcdLXHjXLIzMoqZ9faFdJWkVjSt6FoeNTVi
gyP2bmlqCxtXWeKlQh1P1/ZgCwREBpAnlJEnfBR1/9I5LKr8Ek8tfbF4UM18xx6p9rRqSEPIXzLt
YBCIEsI0D1+qAX3EiWFFejbDP+KVLkytP+lijUUJbvN88OC85AdsZKqpZ9uM3lipwclE82Jl6y52
kF/MmV1J7FxW59C+4/X/Miwg76mWNeBrPhjQOKeGPZmOmrBEOD7b48Xf0+tmvCxIAwMThXMEggi3
nYrGqxR0AX3HrYQ3nfMqNSTtxwejO8omkdiwVa/T6ZK4hKoL3AF0D6+SxjZj6+ses4+EF4aIfA9J
QlmCV3iPJZgzAqfpsfy/2XMcFg3aX/BJXtN/ni0E70JjXDaaOTEt5IfeT00cG3pLlKppd4STnO3/
1gNeOfxLYvlQmw+9lRsn0TEedRPy4nyC8f5cOhqm/nSDIla1NHoCO8g4ob9GVlS0Xz+9DyJiAL0o
fU88EObqEwfeP883Kw4dlLPPM67FQ+mYJF+Q9oYNyTso1ZaHaTLuOY/+GzHTjmZuPll/weTFu3eL
D8F/zbMeRJ9NTsOVscmn1ORIxJ2ZtXgskTTp5n3iER9UFD9Mn8xd46oBesL2sJfByOE4boGS87iw
AGBw+0yL9oXU/KnoBit2EoZVydcMVyLMMi6Umy0cqQomnTZURYUGLyI+EkUx6scdW2ppwzgAoEpG
MCdVwMcHxEXmusIjr+/DJDeosdI14q3kMlWQlBl3TremwyR/Tp6XAoEgyPwgt+kWzrFfQ5mQHEeg
fGeaFIdRFHTs3axzpcal2gbmcGaf8B/OBS4ihDqTjH7YSccOFkEGMiQXU9JAujpxlkuPJS0PPCSp
uvHxLJd9RMQhOUAuAy7IWEHI4wG794mmVtOOOg+fJx10Yp2dp21F6o4KKuoaRYbpsqjRIanfKMgD
ikIrh+TEF0UwEwJPNk4k+QVLqVt5sngYACvCLLMEXB7ugaFEWR+82HoxyAsF+2TeYs8zW17FdS5N
oLxhSY/e5J2W0N+Z3Efr2wFjJwoElaGS73gU297GsViPhW3ASbTMNox5Gryb2PUmTACMOBumLXLW
3Nx66dQdVkhPLSL+pg+YIYkHWMXpT9Wr8wtfZCS4AjBr0zUP4RcfXz4jzlw4TVdb0weh6s5Hjf1e
Rn6Us5dLvBIMP06Om+iVU9NjALEvA6wmanOUfJ9YxsX3qoEHbpBzlezCKGT6+97WUy2GUagaYb8m
NUApWktBVZrwTLei2lczEdnMu5blGFY3BoOglCfz2hJZKKp/R9r71SljzzFc3A2rgj6Yv9Uc0iZ5
BKqXROOUoVBjr3MCS1Isd0gxSE34iSzJi+lHh9dMIOMluH5XutVwZHAVqlYLI2/2s4WOW9+6nynR
JbzDVlqu7oJspuZkhReJr6JbUwc1tcK5fNVuCZagpBl1utABNz2W0cECrZiByv/zoAeSL/eGQfHH
jE0kRKBGJ6F4vEq5rE5f7wqcLaEBRs9/a0yWZv+Hu6pZoVcKdqK/D8mAQjyqz6TfwS6I2dMDlrdg
xKGZiyTyXSVbXxj1JouE0VS5Ifw3cSd08wVDzc4KdxcvyOi8BsP5EsRNqbV3afNypPz5556Bq9XV
V36N8GvE2v5BYfFxnPiFoQYBHJo2jw56VoXX6Wwar6KhBB0XlOOmUUbqayKQhkGtxJvnVTeWO3+j
KfHatOYbGPSr1STrSCaYKgoeVlFlZPrFWcUwhc1YyMrs6vOhalyNh9LZLJ9Bfaqhcxjh4B/HMPxW
IDlxTeU04z3OHRXObTekIOpCB2MKkqEPGESxtDwGZACUyeVTDHh5CyFXHHF0pf4wFwxHn8+RzDwX
RdxJqFLISg3tx0QRBu2gD+olVJsHvOuaN/mw3iIpdoxYUBKyA1nIuvB5/++QANeTlJpCybiVbj+/
IEdEnUvJXpcc34LzvuvBvoIyYcF3mPRw8zg6bV5SiMfh5maE2K+RD+R3z+PTZDUyoRPCGQ8n0nea
K5kuz3+mRjLDC6RFuKc4f8L0PIIw0qI6bqKIt1U8sEkivgSYPTfUul1Sp/HgRDPXZWFEH1E1qQTn
oPJWnM1xsJ/oKIdAi2KR6Jr7fasaNt2IpgV4flDFqokOPqwLwssG26ZJXKyUqAQqyjni4JJm1Ipb
HVebFv2+Cw/+KsZQ/uCoLJO+sapkYM7KhLduU4bxR/zYHAlOFo1gxv/QWTX5Em5IvypqcMhluDmy
RwvvZopNgfAsShJZKogn2Nl+c8pYbq7rY+1bFfkfENLhtX2Ar6lgwHzvVvFxqMKkJXG7iE+lwcdy
xJ/+KYaiWsj06gbk6FVv2D0QSpscuBcU/3iKcXJa62AhL34Sd+QnpFm3EelTMqz0RDhcyIV7YAuy
IrVfwdgbjjI7rEgTq00fx1TnT2YJgHQpXTOr/+WmYLraTOTVumZHqEsTEVwTI7Oi4u/K6QKMqm7O
7OsLZEV0qIzFPmjkmPAy/oN5vpqtLL/RVtvQBgkEshTulr8F/EqXjY5vz69yOptD31NQcQsKFwgO
PwseLspynunVGH6jtlfPHCJQg8N4dPOTCDcdQoQnpq06S63a7mmMCUq0RSYdy1fgmHIY6rEXdtTI
U06wL1jNwXb/ZKftZZ0QoVpUl9Uw3d2x6bb8ddXdCsXJbSJrPwIcT47Agbgl6S2uR5gOalQtHv30
yv6yoZRPV0EpI1RBqeCoEW/mX+GnEpHe5AUoD7OWK4txMljtzyGGrisTjj5AZ9VzSPhoROCkCCV0
UquTN/zlva/P4DCBBCqoV3Yy3R7P7xxreJWDlJzRmKBHPgkM4XJ8Go4xcwXLtyHcZQBzzVMCJzZ3
M4m5UoaWmKKB+Ejhpz0U9SJ37ikGEfnAgQ5P2mJAaNOPAd+HqGYP31jxge+9rfPrl0CGx1F3FIF+
kxDGStJGOEccOuHORRKFWoHHyk+ED/OxXHJjLUMwUzF7zuAfN4aD2FC1srFom4HCrx+mptH2+741
i2SP4darxhLjuQEMqOpWzyIJFTUGldC4PpKiq1wvs2ix+GezYStnt89lFpPTAndnk3e1k+SJdtMr
W5VO1Hscd9SOAWg8DVdrMj1Q1us0PGnBDZ+Hf+0FCOLZUdvMM2KfqoK/Sr4iukWU0c1XPsSrp3tP
+0tUe06hlqv03kEzyl2dWD+tx0FQMI2c96azugiBz5YjoPCMeWbmmpVYN3BJDNjoRxHvXFANVyt2
aAh7PJvJt4b2cKwX7QXe1ieQ+kAomzHBduEzop3Ic9E683PLDWcy2CBX+Hd8xO/tVxqd0ApROICk
cE++LfH0KUCo7BhMPUQFEJ7z0cJ0U0JNwmSuV9jQHbP3UZC5bHW4TX5x2gtv+t4bAKxzNKfNaUj1
ZLGY/LZRt5Q2OSy29aj7dZUpvhChDBpiAQPQf4bUjAkIcDErPLX0Om7sNXDEWKfRX+iFdiAgeGE/
B2T4GBjZCH3ScQx22+iPW9AAbvKGh/zeQLO7dZ1yE5g4LctYobmednSIe5DLNWYANK4kLaoBnq+J
JNpW/O5Bq8P/u+IsTgvLS5R99EP9mvHE/f4pEuPV+0UNAYBBv54gEj7WhCnvW9V2eKRp1aiK5T1P
TJ2hAKPE4AUyZ/NjYhXgZSe7E+MdcmNhH4tRGmu2gUcWEFciGyivL6QoxgTdOV9tkbV4+FpTByQp
h+sNA874d7qdlxX2qWY1ksPLRTSKQdjFbTwYutVDba/bnuHZMIu9Xjta8Rdlbjp0RhRJaGGpYVSD
HyfwB1/ICn6sKvXE/GS7F9lBvw6xhng1fr4g81ZApfUckvMax5o+6DA1ydVc+N9cTySEjHytI4Sp
Pqjrk4zsPU3SpCa3md1f8nU3s3hM45Ftc42DN35IWg9y98G8rfFY/ZZQ20xFqLctoY8hn60oaPlp
ykTwpbCmMknXLFF96VzLsyNLA7c95DPLoe8UkQ3WTxte80cVBArYkx/pNSSyLF+XH7gWtviLgjkN
7EStx+muJkZeNFAoJRef93Ws8SKBvol8HlwKmPQjzUwhDDg5mEc62BYdfGYGmF3iefabiiKdfBhl
/LqP9sMmcmE+PL7X3jBBhf/FPvDjogbGgpBWTN9Ku88IgNfIDtFDMWR6N35YS4EnQD3vp57GkrRH
dCkcDl5eZI2A03HjTeEDekdsa4+ofWiEsuNwkpaky7VNnmiPJnXsyf3NCq/GsLx5YYP9z/e4slTh
sVVLlKu68YiiBSxLOKsW1+ND5EMH2jiDScfIQj+AYINboPjBaKP/HoRIr2HWzs97MMy21cgX9+zP
QYmYSxvMoIszOSDdcKN7hWB7/y9LWOLo/OBarG1v48UcYJ5OBrmcax5CVrOSl2Z1ExgAWTETBVd1
08x7LhXRjJOd3SHt8FknvBu6RroDPxtx3YCnzFuugf1ZXHhGog1YdHWpsScHFg5evZK6FOErWLjW
OWl3Uw0/9aSzgkVLm9GsrKmDfTW2Djr8qHD4Fg7q4/xsRb4IjWb6D8pIRNH17NWd7HszUfk7s9Gd
6zULA+9SXIsQmDsb1dEsa4oS6W92PO5Bg7Zo8Uvh2rk8YTy7DId6g+9dTILLwnRpWOHn1Svgi0fB
MalryI8VB6acEdWvoXu377+2YkSmwcmv1GR7fBRKMn1lOjV0kssGYI1sO8fRSZJQ903Y1w9z5e6H
QQP6PVKLK9Z8leEUP7poXd6SXHToPu1SDK4devvYR4uYQlaQRcE7sMvdDB21OtQSv/WDsXBGRTlZ
iAspi0Pzdyi8Ma2T/FUfSd18sE8tiCMb1s7iIFXKVn2lZkwA9DfcVvv+pKl7H65dwf4DeqNw8pyk
Gt2Xi3QE2mPJB/4b1suy2+eNeDC7QxBbpNlbcRUlH6WNHAESq22uZ9UTcnKCvDc5S82ATFU0DGDC
HVVELMQ+FcQIh+5JxPj5+TWR4TSIXqG8S6PwGO7t8ZjavBrQ9mpwp4HSUivgWBVB/y8l3ZA/R3x3
esSDb5xZOlIW2YoJSwK/5F3TmbgZKaMYm1O6l3CdffslUroR29GVIarFFZ/x58tCDOdmQrQNSPJu
Z1Kvzv43WHomkZrQj1yZ9mvsDe2zmzvyPPAAULMeul2kGyzrq9jb5aWxcEXhnsV7BiN7AnCrjlGT
s+CeyEPpvzao3zWsi9Jh63Q68iyQbsuPb5vHumLQBB16SmVnWaKH3DlR+HNAj/F+6RXEOTQc+7uZ
oi5UbOTjxNXhzEh47v4l+Pt71vLHiuooSHvFGJD+koQd2BS6ld+h68yoUAsAXvRgMPr3w+u8cwHc
/nqRZZA4Q1Etq5ly1CTuSnfIJeYtK9xuskRaKF2tpNWQHsybFEKD3Jr/gEQXKdewtvIuAILUnj5J
bvi3B9OPfPlKC+q2gPY8gMN2//wuX2kDS7vI0lT4vYhxhiBXCZopQRr4c5x2/NVKKAXg6Jaq8o6Q
/tMUoTHBRfm9mMdMdxqSfBU6TlglT6lLkbgD5mkDwdU/mLcUv4rtOo9EFL+pppBFuntLDOGOrP3Y
CYSDh7LhEVLmXybTbL6bQqDlJSlquq+bEW2DbAxZw7peQjViaHj6BT7SoPJC89rk+4ZmKPcLU46V
mtpjddqMisN/JpuTYm4AXzFYUNGupu+jSGTJ8fOnVEjw6/Fe9bxbM43EDWB3NHYPkidafmT8Dxpz
vAOFt1Bt7DNoM/ytZs/3kMaY6Wv3BzQSPgcU/FznqXElNiPLY181Q+CRZcKc5jv1oLNl5kI72L13
6D6WtTl8pCo7uuHiRFc4jy7K3uXRg/dLp8KgLfEKEAxHxIJOztzqfkxwW/sg9wetC8PgrzB2IcjC
nRpkPfGIc6ANGNmdFTTQimrmytUzn4jppy4+kVlYiKuzexhpTsL/9OrwKYi2edQf+ZOy6XK9q2pG
0NjldB0WOu4ZmFHjF2YVthdRVvTNu/fVNtOBaMqH2ogex5p+hrkUubshwUyo1E0PTfIF8RQNDm/X
9Wn690BZAjQ/iJrL33Ndf7+YSfqXOrbsnukal9T/HbYVmJCgTOUR0ceaT8cKSZu3sHKjCzJQBazx
fJLQt7bXxPorTNyvDZRuabQFlRGjALHNFX3oXuP1Eop9JcN4mOvaSMx+wmyPR9lFUirQx4Swel5t
Fz6AW/0XQ+yEqrEtyuY/3bDRGR0WYXP+1QYIAe4xT1yekvFGhfMfEmHfnzysCmX5QCwnO7dw7py6
XLD+7Lzzaph+oD2ms+yHoG7UwOOVnarFzg8B7ArBQXno6rhF7plrauHrzBxxYzJfVc7qlFWbZZO0
tcJLAx3xwCuX5fJEKJMZgEseBsFJuaF3tMRkPAEab0+M16gdezRBvEzwT+g+dARA64TAyLuZVSA8
PA6xG8M9YRXhlrUUthXvbLCBlfaZEOBLgx7w1Dl95Ruygc15G394fLykT1wWyOQzV5jFbr9xllKz
iwHCotx5h4FdtSIgtO4VBLY6+DfW8Xwzr8I9I8+o6MvBZTkiZV7yoy9RykiUGtVimFe2sZNT9BP7
g6pkbKYsmbM/rUHDIqD0a4VelRSIgvx9jLYw18qB2td6aFuPj4/fRrQmMj/yPPHwP02Jw5WXNDNs
9N9Rg9cdHVeJcuAjyK/9zW6GeJmf0/K7rEV4tKmineqYP57JIu/MOlEpR+Gr134fPRvPWaGI+I7Y
7ayhM1Xv3fnkh2mr2jE99D7c5iLR2x+Q9YVaKrR3ttWk5//8Y7w907yz30bn4FuQjOB1ZoxyPCr3
mjBxdr/f1ao+4rv7/qXJaXegJxXjn9Tn2A0/B41kJg1kx9DkVP8p1C+SwR4st5PJ1p6DEzn+UFMA
V0IH4jNDNLA8dMKgoOLBnttUeUNk3997CIbrVMVEEXcXBsXZYBpk+lVcojc9H72/1sS4o3pTe3ce
1IXO0LCdE+xLyKbVHCEK2FZfuhZstUs1eMszKRe6lh1UCnm+9eP6axc9xv9JC6EGH98lPAFa5mW8
U5xiU9KCGjUPKKpDFwMsQ2GuG4U/nXkTNbftj3hlGPf97I87jyeDoZ/g1rxTDhy7ve+TXWcWBfVQ
qufkpnYA+aCECfH/4MU64/KrorLb1iV8d0RiO8mJp+B89KoDM85F1M5Qhns0IiDlyvcEvrPI95N9
BAC3MzgjOCioDw+n9fh8EqRYdHwZPQyC+5zD/SgzOkXzrEB0nMVimnjXIkwzho75tr/rQdf92rHw
rk1WZ1ys8QYFNZ7UCOw9srehrbX4F3uHSVgVgcDptjcUlnDkWLUZEVCxXD3OiWdoZgYIZi5lJ7/I
BZSlE2pBrrAcxiTRkasSrKMqqgNXGkrR+KnM2HvLugCGvlCF9XIxyNB3DE3YmKAPfA5c/KIntBCx
uY3JYqWgmyPororfLs9IMrJDeBodhG328mgBeKsxLdHgvomz+tMv7clB7QXr1H20MiMJWQZMT5Wu
j61xcB4Nm/c1b3qtUoE+JaOby4Xbn0EuveEg3XVDBGdrb8tsnI1yxktEFsx/uYq8uby8ne6AE57A
LIyJEw9MSD4YFfkIe4XVETQWS0DopEzIXB2SrxT29wTyiZQnSkes1pHuVB4tFWux4NBAf63PbeL2
+kNYZ0VazfHaYd9clWgK+q/vows10kKkQNNYy/8nd1jz0ofkhxAWpPiv7xfeakXRA0U+0c5dRDcH
THP/GgRV9uzFOwF4LDg072Gvz+Y+LCenaTVZ20nrXa9ktE1+oAx/gnmb9yLeZe0hjjUpxe/MqMUX
/o72g94Mvn4AST/hi5Fnk0XQ6TQgIenBD8eFHEW2v4WNOpTPZbB1waUqwEuQxff17jEfBYUF0Kj+
F6lNf9dj8jVZmejZ9ikPp9iQDWVesVNh6TLQ+ZxTG3GEUOpq1qXOcWImGTLCFUtMiCLO5qeEl740
MiucZk0e40nYktP5JNPjIO4t5GKKg1UB4azH3/sPJ8j6h1B1J/gEw8BzKqfnjMsy4gVMSLHEDSlb
clXfnW17eeXrLdBN6VdqGqjeoTV3zEjiGjvPALBgtlTHnYH5LyDF2x4gAQXXxYruEqNZ6cwk6LGA
VNM0NhNbVIUNU1NVdJ3GmGhjtTcLDxRaqcZ396sXD6Z/UzUUkKNJ3iftyJpnUuc3J0bkNqTFV2uO
RY4/5kLDwgsisspjnVN5VtaU7FNQXwx3s0lqNkgK7vjS2++eS/Q7vkNm5RzzpC8fUXrASi6Yl+tS
KEwnAPIxUdgxyDPYvg3v6TwHnbuy7ubqN3PbHxgOiaDK9fRZLfB03/+BxGdUneZnwf7tSVh/T3jL
PutuZ6HN7PB7UU0QtyKWUTuuCU/mW0yGotPmZAnPor+4lwchklLznXhHKK0wdwFNYMaTUyy5ZWII
cEmnRe9CiaKBeeRoBDqm7SF2rKmBVD193nVJdbQaaCvnu9PCLnbL2J5haKBuBb/kD8V5R1UNhOzk
ooyDXuJpl+rtA+D0cST5RwaM1YVHpWNZXHpfJ7GdRFGGBLOX28UdVoTPSOXgHb6hL3aR06zHkPph
TyHV85TogS9UFfiyQgBVMCtHGKU8ufCb/7QCMqBbl/ZSbAcU6ELCjatz9R/eKKi8U8hA3h8xwFwX
aRjaMmVXpfERTMnG4aDzUUerieU3YiDj5ckNnDdTNcUQR1X1BZ5H5fENv0gO7/ccAzvyoEAPxwkR
wJJ6zx67w9ekZ3rAEx1ouHdSVObF6nPWYnstJqymog4l7IL4Bpn7IAWz8VrS49ZaWvGFaZQZLaTZ
BE7WOjh6ZDZ07+Jf5vV6+F7yAVhObC02zhnyA90Zm09NxzKvbMseGkOfVnWuBOuTP8eUNksSuJef
qmPg5SC/g/NcKDHzX+GuFYUV8B8Buxpn0E+E4Og9bGJZy4s5VK+8dm7BjnOBvQyOWy2VfY9vyzjb
rDVUJziXf46Kfuva+GIxsrRwoTLyQzbB0d/Mc96zISTWSUzLzINlgAjBtfL+G2lcGUEIo+eYmSfs
WOoZzas/+kS61WG1FBrc9aVfhsKO2VD9CKuzfeNut9FlUG6Mgpcv4Iar8ueydD59LPSReqODfsg4
ARhIfzX4vZtmdl9V8Bbvz13rVWLGUQHFa0BFZdM4Tf/4L6+ZHXstl13qlG+DECSNR4LcIPUGkHAT
rTwnI/M9QlYkVv1x+SJapqEFD3houx67NjbvoQKUrQRLahjiPgqH/2BBwE1hjbaMiMarieOweyP3
8X/bwWfrbbBrb0siHSLs0cpVXtfgQXgGeHquaf0MskgStefvRmgLQYBLOsKzpP4PpRbUDg5nvLnb
yVV/RK59NflPUAUDlxe63Yko8apGC0CseaKJkVq9jpQsh1v/bbIEQPZ69gfVXuYEzDBnucynqJ0O
SQbMNPSZ+NSVSk3ApfU4wiSHTtQ6QuYhEA4Of6bUhBUOPLXIyVmPgVaOo8z0U7KOjQmDotu80+in
//w2B0ALEXct0jOCKySrCaqeD0buDO39ueqNVrlv8wqY/2MJzda99cs4tHHMsljljPVxwnp78g4O
AXgqUzZcGwc1+gKBlJBT8NfOTpXmfRk/aLuX/ygQBn2AqV0hJ5mMIi99MDp5xQzXYDesB4X43Z1y
mNQJlbR15vtkWn8P/6OXucJXaRjdMYyuiUCHkOiHDwjSToUhNVVZFr4qZ//+dMfAJV2w52yEh/Rc
HkuimJ2dKBljVQ+jM/P+AAypNi+q+k1LRWhrOIjtshuKWGaYiMQqgFEubdPYCmPN02Y0D5NsJFPV
bJtNamK48iNuSZVqY1/1EkAqXNzWoynwUhs5sI4uhN6SiaDMjRS8Vk0/84LvC+XFPXgJh6Z8Vo43
P45DK/fnyzrEAXZzCsArxFVeDQ+DvTUnOm9jKh4A5O7owy0mSsCYziSO5UPFEaty66w8CS6+Rsz7
573fuleVHeyYhtBc9O21UsgoiFuFV1V/4T3Q8Tf4kOIYLZ91t5aUf9C7ptHXmz2ASzstIoRAogdl
BIfrojVFLYcCBanvVXh0NvRkwNJsGHvV+aV5QF6jcd4xSaNrQo9YDQofGs7sLIk+4/X2nkdXCHFU
LpEQFNSdk+6p+F+eZaORiN02tFk7BkBNmB7WacuLgqxFFJO2C4ApQsmWSifg+eGlT9VytS+GQFNN
evxT/v6L9Ur7RJrb/cjs0CS9+S1Uh1iW+LVhvGqWh4Ns5UZw6Ius+uzMQO7/EGxt3lFM+EX8eMvj
dczDZ5FL4+DchwJKfioK9IBqr3Gj4u8jMix+6QfQkNIvhTldZdpeeyH/pYVs2PgLd+B9PnWy8azq
ELBQy8oKOLdp2vmWFR4RazB/fpblumZ2VhzIdjQfyMgyf4IEAmBTRBQT4TzrW0SRGTf0hrwDdUwb
wN19yJM7MfiZ3wr4J0jzGsqinItR0xjo9d1FpJOybeYEl2syhfVIkw5QtQR+Nb33vJV4R5Mc73+S
TDJJQzxE73T9VbNzBK5GLsOZ7d6Na+dMGNshi0/rX+oec9aO2CrBsQFLACeR2pmy0+hA2Yzrg909
tEbhuZdLQo3GoLKL/T5yM0riNyDXAHHz5r6DGHg5h3NjxeaqxJNZORxbwAtS9cemJsI21rjD7fwA
K3PcB6cRB6jPTGyR87b38QZccFXBnejvTsxBxifT5qcc3RBBRPC0Gu4qt05vOtwEnj4UFmdlgriP
xwvBR82DNO38f5PJrXxTh0HfFK4f8P6t8lJ4SmX2kDjpcpgzQLHBQS9yKszY4+8QTtVxb2+ze7Jt
oQpVlmBrvwQQ060sYgNYjE4MrEx0vMe6iG0WueSohRaCu56WxCwC/u1JF5Ghl1HTLMwmSQQqUpjN
n1b9PRBuvlll/Ub471RWxg3x4vansGtGbYnBsMMJJPUxi11ClX+YZm+lCLvHIf94cbr9Ay4g7YMW
ypmAQinDi6vtsRMf3xPWgkI0O2xj50sHsG8r9cQ1zUGpYUqeR7pqktacrvkf/iqz236KORAf6Mdg
8eEVjU2luzsL+KB7Noqd3OTUOolOSXaEb6R5bJbS7+jgm0mF1OqjbQSVcqISthVsx29VwSvoCqOJ
rFLvVCoJ8WuQvTpznxdxw2tLC5TcMANjpifeQecwAA48AlMnDjtYVmRzNwJdsblhxhMV5N+hQ5/b
RMjdrKtBE5CZ79YxiMLRtyl9ngGPTjKwykxNsXyVdBgJu/zXZHNFoNyTRAaLgL9UOyaR4g5b5lQ5
ZfZ68hLrhdhCkayQRHgmhuxeGhrQb0i8M/pjGf+3uYA4mwtdamHkjgivRpxWL8e4vyVY7Gcq8czF
ore4eMkmjbz+oWh0a/naLb1zQboEbXVKy4TQaUj9tvP5M7EJ9mnul9w1g8woV51izZk9FQ1qn8dq
jmDQZGkLeT0ntZBbua2+tyFTVd9LyAczGOoqrhqVCYlK0TEhnCUt0hg7a1YdPvVugE60zQLqIBhd
SKwSbCQc4aO7E1KGCTP1IYK0fy/rNAy4Pfpjk+7AfD3zvw6a0tp957Y0k4nTGRZA5I7z4xO4n++x
cbqygcyQxSzLLeQD9Zjqeig9MZwUGuzKO0GiKdC8HUm/n9CRbjdKzgsrbP8Sk110wUtM9xERPsm0
BD9CCoApye5o8XALI1QmMmOqcHMwkAaAPhQNLgxJ11kKERviL1MxhmhRqZQ6iPoY3h0hs1Afi7be
AL7IdxxeS0BDiPAE1Os6TLV+r6QBZpzq1Ysyu+ElcfzCjozEz1hki+KzYXM9JcutODeRaBA7xLHi
k2F6BV5DdwbGReFN2X5Zn8V4U+evJ2hmYqk7MEMSO3U2QVxfTDrMSzUWn4SYEJqer49VuveaFk7K
E9siqX9QJzt1RWRT/Axb61RO2r4wyUkZg3t1bjV6a3BIw5ajPZihKb7qUbejTPK9UgJqIepnwtV6
+pbStQqVeQM28WIbyd3kRXpJIyaybBMFzrNoUihFwB540t3qtcsv3K1y8Z+SIM2lIR62FqMQ030X
xnwivTW0h9B+OsLmi04HbtRkzMMmIA086G6NiNZD4RYGiN6Ngv17p+b8Y8Ory8yRXUk0z8C24NXL
N0TR4+gjaCcAEqfP8dUvmFj828iCi/aAV0uA2J4AsnO0QhMkEu1KW8JPHwLS4B5HyW082daEO64A
6X+9EsrPrbIvi89eT89l3OJ/5vc1gId4O+IAzWOqGkweeDvsF+ZrNTnwAc+FdT9E7028DpKZVUN3
Ng5uKEKxO0QBglWy7PUlNjDowtWgysAPGstWpYxG5l61Wu4PG0ZThFPj2pbm67D1xc+/C9HVmA0h
62XSzCu9gxC07tvy/GwD0jpQG/haKRSKQKk1L5FR95BCr74mbLC/DVTzpZdjjlbd1PkEvCP77ezE
KPeAuNqPsSEWc+sG1kW2RrMCgmrGAPFtbYBWThSTY2kfj3QVM06HDzjqfVmWzfhieJ2rAfyz3WpQ
oGyqhMW1Be+QmpBPODljmlIQ0u51HDjoeXV1MMU1guyR9vM1VRs9pomadyIfqZ4xvZbnH35sk/C9
Y9bedHucyvVauGOHQAgIQ5ogoeX4NITkyQxnJ2bXtYB0oGm1Jz3efUSCgnEX5g7HyA/92SAkBDr0
UwqZTKiRFDi8auEgcIPttvGO8mGMSJsI17ZX8cNXT7V6KH8X09c5zVMTc+y7Y/xh4MynjzfQniC9
x4i2/fYx0winJGm9W9NLprv+wogP/h2eYmxRw38QA5VbWDGlgiaFUct8oS/eGEltUaIS4G1LxBCN
ZN6BCl6NZ/5Ltw4GXklSFgPLXCrrO52BW0HxDd9RVP638nAYf5Qk9TQGfwHdbe9LlXCBrMxIth8+
HlflOAOXA3DUv99AOHHf33q9dmN0lqIbJ7q/hxCuzFIn8Dw9emEbe7HbIcTZwKViEv5n7ozlSsnm
THjswiS9igQw8MMR71p32SJnmKxJJfC57PKyYetTscuSpQlqs8VuDCpsuHQWvqvOs6ivavEKUjpS
j+KIuKJFghSDILshvURUXF7T0QZLujqT6aHQrO6wsqL2tOGdEkz65ypA3F4FJpcXmE4FfLPueOXu
sd/Umbsr6uIBAppt92Cj8McwovkSSnqsyguc0hqMETY4sJqR/rv6tGcctdbEBzKA9xDKzLbNZADz
nQ/MoEPiXJ8KAdMRVswzvc++3A5qkBC++5/4snvkrtDFP8iXOK+9fHg5PzmZCEjOrZwB9Uo/zBMf
66mXx4777Fydwsr4a19yVfAKWd9nmeh/KGuTXxA9cM+yaY5ENiNeVN7tMWwdm4nURbpfeoYS3c4X
NVjK/ivPKp+Znez4d8NOEmYUTLsjq2aIMRn9gxfWBHDrNV33v9Tt+IwucFOUqR2ceuFyHU7ZWYS0
gfIg6q5uabDftMSr8gvYq6h0kdtgI3ILFDvGl+g5T1f7SBqVafBkik8aMetnb4v1byc5a4TlA4yZ
jmfIj8A3NDI1i9ScARgmAf1g76jeLnpX2vKFTRxGEWvHUCYRwATc88hlkLwIiB+eYaWFfl93cOlX
2frdZo14TV0bbKOUnt4mkhYcL+D1sCcCZnUx7klNfOX+MBZcXoPHtJWBpb55VwOJT0XBrEcY9V56
tDckSerGpXyHEkos2e/NnKRgaxHgB6rzSNXFufR/XcRoPl1NVnHal9iMjyMQN6iTR8vTVIpYOE7G
mCNBKTfHi4XTWDavk1sc7LBSZOKfQdxJBv0pjLh6pY3q4OCdSjBCt4ES3BrL0jNljncM0IY6o6f9
GNXkk+A5BzkOABGrKrAjfrM0tWlJEmt6+9zFBsetcuiBpZJxLrRvsa7Aw5KJ8A1F4eEUTIHAhFdE
bFTs/fGX7QlY71vk0GMFseOVPE3bIGAX2ybbDZyoSoVREXYSTQrivB7p2R6hIOteUqbulB0GDYPQ
AdhznD70Zzqz12p3GfwWHefksLIO9WgqGo8sx1gRhV4AgkCx8otpN7B2NCxS7pYdhSQfqQlQUoAZ
FIpEOyueDNUBV/E/haCTV3Zl8U/DtiEKhIcohhctmeD1XVZZvjT3fM0IgSQ6hLfNOPccjfuHrzmx
xWjZeI4+e13tfcTCt448CP69VUnciJ9sE5on6xRd4NDNy+YOVOMl1AGyTu4on30ggHswyS3cJpP6
noYPrCIzt0+xLblbVW75KFEFvs/W4xyTroH59vAx0zabSkb3+mjsFSSXyTWYgNZ2S0PUfVORDAnG
AlkIyFviKbKxhQYyWciCkl37ZedbTKzwEJRS6Y8UaX/QiE+y31XUe8t4Z5SB0WDXqyX/x6eZph/o
+giCOYsWmx4SESxOuYsB9K5aF1l94t9hsUBON9+cdCnVBmpjcE4ZDHn9pYEhplr8VxxknkbQc1+H
jp1FfxPIAy6RHZ0blbBZctDL7Pbq06y3bJOtmJQUthWjK8qYUBorOUmpcXo+1Fz0t7FiFhE0HyoB
UQbCehyRCakxBVeOMkXZ9viuGEcjkx2GK3HWMTxCitO1cES1yclYIxyZJXhqvZcuUG7uTI1mIEND
UonCk9XZG29vBVRL91c613zmGt0Yt81eJV0Eqe6Hck5fyW6CLmOdNHOGdXs8pJ92lokdjviRGx27
Wcu+5VO/QDcMclXQiqzJXyDD8xQBc6XTapLOsmp1HRKnGtwVRFFGSe0DQ0+uj/vvRhTVUVZd7lQ3
sOWxo7MapXwkcWBGRMxunuZwIEzhOeETQJglheoKmrm/tkMeqGmRJZV063DhuEeMyorcuh4MMwDq
QG9r0OtYeTBeXfOKeNz2cxo+FAl1AsrRtn2leR7FfivCmPY8XFkxQnu2LBCiwQLTPcyi4wOASDgO
Ncw5gdJmdk4etNCOgcw6L7/hFqvnYlbrFR5JO8RonXpM2NkMpCB1D95tgBGnv48tBubax/daFt7Z
7x1Ng5uF+SDCeNMfNPbXlaU0fN/vCRJfe4OSeKhFXSpfIVhTvfcEl/1yOpHgdDf832oMCu03OkPV
lJN95NRQX7pkZLOuHm8cfJ+HZ/WVIFZakU2ACikRlIWWBn118cz24lO+M462opXBcic05Knb1fWX
DVJuO7UU4fxK/jV5HE7JN53NSlSORvl5H+KFCtsdESmUYbbqejeKuXstAt+xl6E1m7mEXx+6/l7i
512yImyfiL3KbYWxrVi3ZCHB5K+yuOl8SBW3fiPG8dc6YNBcjSauP2UL70KDhbYBXPV25qPiN6nK
TSthIREMweznxtFrTOwPxU5T9znrwBPXP7UEqv0mRhP4ZwLtZDs5HzoyZiXiV97LyZDsYjSSkMfo
Fz2e1Os6OdaJ/hdbG9bfjvQIZM1+R7VMfvb7OH4PRby95Y/gBAd/JtO6/1uAcOA96Ex5Rg989IQG
pQzTW48re46BrF6f8kMGw5jV9STYO2iACphfY3Udg+I8iX/LbhdLz0QIwAtuPj6YuMT+PfsyZ0YP
1KfN83j9TL6R1jCVRkInjc6kFbSoGruE1v5tt8I7FT4q/9E9g/O9ASEkCgZS8Z/GJLUuMQUuazhI
w9hkHrz/o1MAdU/somykuhTQWlXQd6oo2WYhnyoZanR95/SeWADteQY8jL9eh112KDmnEkRfGxVh
o3N1qGkqrRRvRMTLN4cWC3QG6fOMWeV2C97+om2xhYQ8kubnzAm4t7bqhmjFrXeImOF6JOe7uPng
FVWnf3XrDB12conlL8GK068a7xdIMcf5hrJcNmWt5xyy5hiZdoeiI9HUyvs1X02/cLna4H78/37d
5LAPglZaXgRn4CELCvoTfmUPbnq24FjPOXBR86ev1OHkbySxaaRjJlPZRSZJhSxQnolR3rKgP47q
dxlL1oWv2Q6FO1dGCTYbG10bPylOCI4W2AaHyYd3z78kR6X7Obc5HTfHv0Kt4Um/IOGSoLMVhRcF
HjthH3BcFHR+k47uzQMvX0UhQknFMSdp4PeDQwioMqQgZV+4xpHumaw7K41Uqq6x3cBVEjKzHmLt
o72/puRmj9kRGSP04Ifacdcjz/9cLrxdrR6PWCHgls+O90TWlyfUoSJvMM7RlW1ffeYqoBW2Z3dx
mOxGk7sGjHjkx/F884nl58ykkntTqUnRnHuYiiDll0nHtt/naPEYaO7thPe+ukzHkJHgGMVddLl4
19utGBC1RdtEbOvmpin+GFGquffdJvJunKLa7jWuSltuCjaR0hjZIG52NLle7txOFrGC6FvJAPrN
QQwGDjBa8G5wFq7MKcmx0ZEPgXOn5FKY8pUjOMi99Q0/o+ElwYqcC55rI1blcf3SDE9ogScMiv7P
y5W+lA0BzxgpMTxazpwteWY7HGNdWRePl9zVH40G12KwtSrKJ0BIKxrItVqdUWzGRzCJYQ2HWnPY
q4eCew8nGz1AHoS/bPctkg5GjE/X0vjGn5dAlFcaSbgEB9HhceZSbuyaYFOnusM1nMgJ8/JRc6NG
H4zo+sND+mErjescIT1q+i2BVYDx2E8VQ5cHLJNWrj0tbzJfwqDE6bhxWz4dSedyzWbg8tzF0s2L
W10pvGrn+V3hsmXS0Q1KMhTDEFXyC3q4in1Z6Iz2hOSfHQ59baCqeIR7OIALgVRin/QaqZB1gXdz
v2fx6rTqxBA+CIDH4H8b1VZ3d66hkUeLLAUz0TYHFn3GntjLXEVYXGgbvSqvD7RRpS4TmigT50nT
/ETKAASfg9H5mKvTeJgWCueSXzr3Bu9EoAdrQXBxhzPoQZnRZDbCIud+mQDhYo1Vzg8MISXqIhdh
upldyY+UdzXf3Lqcvu8c0ySGnFoZTgXFqnjoGSCNaxHq15Fe10Hlfkyr9UPYqIrRr/vV0EGnfZnM
PblVXEIft7tg6Yav/7f+9vw9KDPFm04PilHWWTc+uUpykSR0LZ/pXeDICrcMMnxXyO0GEbKUJo1u
O2tM51VTt5xC2ZIp+JPYukLjIq7yfTsWvv0koy9kx4BO0a4QqM/6lusdSK+0AiWlZOunFnukok4I
EUEMj2N0+8ujaYxBoWRvCmCF/dvHFqpoSTReMKhEb6rpeKyGvQSHqRZa5oWKfhffv/QHlQVRDZXP
fmPj9IX8p11902MqPnCtr5RvUzgOqE6/PfmeTIF5tcIBObrv3YhvAtr+x1HfeZ6OPkPmpBv2AgF1
MosEsoEZHK4oqStGza/0ibwfNGFhfZmoTVCpGu6SVVth5/fTzidLFCIWplkxH2IBxFiMzI1c6MDa
JGVLoNud+/ydBzKE3883IHd8bTfEgKa8ZlqQyGJWevtdS0LXbArXEKkvqK4/TBvmD4SVoP+ivEDp
wa3bgy7MzHdKHBhbndJki2rS4n+bPTG5IiG849X4g8kqYoteHovRzpM2lgadMMmHqES+6OtCkreJ
+iYiF2Ew1nDX6QP7ggsgTx/TpqOKofPZwqvB1BJL0ItvpI0GXOp5VLaA0CU7VX2ohCx/OjqggKhM
qwezNnDaxPV6cOFZ1vC/sWZqy6jVBf2nEGBzoaPL8jm1pZAX4C5rZtMCdLdwvqvpBxUzJNIxqEs6
W6jGQ6UoNvPz+TnQf8DQ/5q5EdvTdTx3aQ/XewoVLdFCFUjV5gXmpF9SS/w+fXKzN8RRhYm/goei
FlkyFfzVUw3ADwb+2Xubx7kL+CgapIjWrjlUzlrsbAkPft8eV9pM4dkNHhQB3p9Hq1rH5bn9uSKI
Og6gfHUiG0kIOShGgyt/dIwNw9qIWPN+JGJBiW4nAXRhPzprdiDIlyu/Lp4Sjtzj7dkHdpvNP/WN
OGQ5SghiFJo089TlzTRrpPqZPpW89ym0IGSWxiZLhPZXL3bOE0nNXm6uKZjgomAXu2e1iUJPH+hJ
epVPI0yFnnggHbkp5ofOGDwLSm+to8jJfeBwpTD4lE/Vr+m4K5x8BKiXseZXzbua+IKoYRwr4Pd4
hnRd1hE0qZ9NAaMkhwc3g7vIzvAtet/jENUO/pB9HMgDYKU5xxqjxN1kfZ71kkiA5lfF3aFieatX
b3vPAhGUyCtqcrUKRQskZ7F848vPui7GWtBOAoWUJbFwPO7lIBwQxibubrSQkBDo7i8WmW7J1f7r
a8EBbIf0V2Wel4gvBFwLenyUZ2iQj63xcGk0SVdOpGCEUHMdo6lf7Vea6uCP4XI7e8cE/4bMdsxH
MYwovA9UIMBXUMf1Rg8Z2vzUZVFmCumWNkfWHfM/ttH22XAAY0W8yastfJsrt8p7cOcqNveHt9KI
olts/pJq5GkvmrAWvIgT3xIRN4o4kf15VFEpi2E+cYKqLXpIpXyhSKC8eB0GTVyF6hlj8VjEoWmF
W0QoWFp5BTszuUxXCxJxBvmHanHtuR8b9vl/+czAxvb1YWriBsRCjx93c2srLEgRm7LKR4xjlGo3
HRrBpGhM6+n2HbDeYIVgQwsrizi2C6GMbRKdbhkMl7uDyLa9ocUS+gb6yQ8mNRgW+ajKIBBNvuCi
4FtoOiOmk2crSHK91Exx6YykfVxIGOjzflzfam9YrEwmivnc8KOUzueT92soNe9418zRWi7/al+6
r5DRUsmXWtc9h6MIFdV1xDjCBZ0IibRJlO9iEJ+Si0hDwdjkHMVcSnnw+LVKRnzvx0HEz20tlOPO
vcbwj2Vp8u2sE4HCgvsyKkNId6HTFmPN8X55aFG5gHITkdj18BTkE+ZQmxO2x679ttyTjH+x5Vju
mZX9h8TrFQwCPl1jGJIzufjJ6CPlLvG361H1eIQy/95CqrKZW/MGrpzhWBqwGCcNii1DwiFUUkar
K5g01oDHXbnNSNFUZkecPoSPVuIM96P2Ob1SW4iq7+VIl6+uR3L8pZATQ01rJFf319Um++IBCEst
mWnfNZubaOJppcZblYtJoo8776qWPfqc0D58Qmnt0/jrigsffAJ6U2QbkjWXRhz735Y2yqdN8yQB
2lcw1ALm+Nw+bzI8gK82WqZck8Nn50/6+y4jvYeC65mw7cDt8x/ue2m6yShTRaLQnPFzxbQWWwfG
sNr6/h0MJ/Iw5PuBncwETj5Nf3BsV4Pq/wQyHCMyzjeIteFBduqmpPuXoBg0iuiozRoVFi8/lumw
wLVrZjWhctNkvTagBiz2drhNw6cKzXRWP5/r/xwWAc6xh41zPvYFXSg6vs8GAhiTGskCoB/cCNlp
H3z9mS5ALIAUrNLeoNvHQryDr8Wrp4xNRHPu2qDy4aGn4eC7po1S6D7BjGZs6jxg0w7/Nl4IS6fE
uQP1GFlioXq+f2V130xKqLNDOiTt14c9Xb+dkU1887Pl8x66Gw35czTKt/A5CUtwW/YF9Ma7zayx
3HPw01/SPtDzqxMkbHRxBbyx/QLaqejSwWcNEsLjmy1Tkojng4SpmVCQw0oepZAnxhbGNVoakla1
9ClvkWG3+Su0opU3SvxguSTTyaKCV7nOQPEeCTe65+7q4oYyv6gxqpABVuW3S3ZEIyKTSY3sDMIp
kAvakdryxfG3pQaLvC76QC7awy2sTrnm68/3XR6jacwPzUkeJlrRagZci2fQij7p20FwDesnCKDZ
Rnr7k9ilC/khWRsKwsJxwTGCZ+D5OZpEn7Iut9gihFDc/YhzI1UN1CZuYrWKKLbpHU12aN+f7O31
HrlqQVUj/rz1Yq/RktTaBehzrbAO6g7WXmMHX4XzIbq+24+Mwi6d9wCTH351afG1bgy/4m5iI3bs
rLpepvFUProijywJjYTaOUc9+l9uA+mCuheu/ijHJawEV6w7CNGcr+jFeLdg7JYMoN9L1xqgtok6
Uzz/8FMrJjDMND0QHaDBZv6otnpz4BEZQuj0359q0WX7B5Ut6lm/j1ygt4Su7hV8pA1LYRXZPhB7
r8Zcrk3tIw6OPTLBstKJAFweHwBIpr9uvZEmDjXhhnz03RwOMVMyGaRVb4C0gEoGbBhBcG8CqSFw
gIc7vPnTezdP9Q8q7Op2RWzPOJfp3cWi5o04n/Q2ahdcIT1RuWxWX077gyuMKFmdCOBuADcDdA4I
w8WMp2z0qO7aRnwkA9ovIFOeZPUKoWsOQeA1iLPsjBnBwV9bBKcXEysXIi07pGpVwCNsTNZhi8Ah
ZvnNHkXrMDrkmMohwmMjG5HOl7wkhzXJUoq0E56PnfB1SLscilWueZhMeewpqZ/sMlBRVMFa0sv3
xFytxUnrR3gPVMrO9l9ZLkhjyGT+DNnWq8q1+2Iv1bIbW9a+0Dbq4gVfaAxiGabwhO0xGB/NqMvh
kvEp6KOByEHb+JD2XTb/a2Vf1F6nfaP8JK8MzvAWfORjuibLaZT5MOpu+hcRrSE3aM3DaL5OLHzh
fylOWQjGfibfAUtXFyz4o12hrO/R5HG4ON51uLyD30jZsHGBeRlw/tbNMpgcAU2B61TYYuOFmjiT
RbKRGzN6xM3cIx1jbY257CIBuDtXEpJj8R9J6TL0nhmHC/oosC3UNOkhCNrf7E5RS1Bjm9ALWSkh
4cV39KnNSm0xuxikw1c6Rv9mc+brKEuJIT5J9NuAhYj3pZWb+VpTL6dA4TPHuNY4vd/8g2enxBmW
aOmTYDHVB68KBNezeaWfzC9xLi3L/OcSj/UgXaZzpErvHQTbayXLGOUvLNoziOakRkL9BHJHvz5Y
mrv5ktblPRbYrcISpJFTdclxCZuHAFjgCy4Ut4mtXB2pSkNrIH7JVyyRvGvE8WENzkcGu0nk3Lix
1J4SQ8GI17lay+7ZNq9JS4XkiT4qF10T03SvWHeD6Xv9nfit6AQDneLX2n0WslvCJR9TfZ0gvAEo
yNlVKy1lkaD6539ftRdPY8vCQi/B5zPPhnl2NVmU+sMzTgts5eyv9OnQNsnELcvuNH/cT2ofURGd
GgFBUcQaGlg7iOFcBif6ZvLTHqK8snuItXZv+xC4cud7GWwYsGaEwOYviuNU28Sfl9tCYLWkcm4K
UpYdGas/uVnZM8EwF/hv/CYF770KMe/ydu0Ci5/ztOQLWIu/tyY7280u3vvICuQKAUFpw+RCihCo
XCY9ww3GWR+tLMTydylJt18UtxRaazVqhJMW0SMC7SMiS3Q7rOYP/JhoqSUzDL8ORP9sl+k3x5WU
5iEhwdJ8BloEdV6ZIjEX3aZCa4DdD16IBTZVY6cubJ5HcSuA736moAbw28LhKqrMV0tArO2/BbNn
YWPTdiCekUN701ePW9h4odn1CEzUffyXdMqwZNc/zq/QSkudMW/65OBBBu/BbGEzG0wxwAqWv3AT
jAwD/aYrD6L/0rBGPMscwcpZhL/pj627Bm7W8emxw3rvaYm3qxB9euDK5Cp+YsjH4QtaS4VfkXhW
zi2hwIarqDWzyOydwFMj99myBAIO753CF1agMOEiSz4IC1iw6QoQb80RFtzdYp8HgfqBwAVFAlxy
mletk9DZNS4+vF2PS66rMukWh8vVu0yDOhvfmJR092a+9qu12zb2Gp53+8CiWonv+ZZj0fmGWUrZ
Ird5bUmyGZnIcScFRpsuXt6pUhxot0gil8L0MvM9pQ0/LiG65bWsnGHVESdVyyRpbfuqmUqS7w7C
vA64pVc7Z9EjDqzZwuZsJ6etk6sPV+tifZcC/tao9vrBflxyQ8xRcrVjq9sS+n5S0Z+XzcB+I/MQ
dtmDdcSrAFLivV7zJ5rQzviMEyZA6b8DThHyjNbeIvqpIjVhsrgfgyVWfqVhn4ZCTXqAdFUfbE7T
9hHTENR/7TjdRLR6Td99vepBuiKRiWDkyNpYwT02qy8EzwCDLGAp6PPsa877HTw5Kl61GYK513OW
dR47lfXKmR7fKPU7c/FlG3YuNyI6OhYFrciNd3NwVtpgEYHfUlw7rX1RJfKNQFjgWBQU6ZGXikVp
wJa6KoGokdHh4QURtI9Wrtw+3sRHzmP+Ei36L5KRxVaxr95fHG3E4Rm8ns/AuaUk0x3HFjVnlXC+
Wv1cIpwV4uGDxsE4v3IFuG4XDieIknMPBLGrn2DgbmUIlg8rnHc/wgAwvNkSrHe2oYIkA+mjWAad
QMHPvlbgTQz/mcP32GbN7M2RoeGgtasiRp85fFr4PECUKrNCacHFKB8HSvVmxr9J6Jl0qq8nWIGS
zCZiyJ/BxO6pk+RkDGN8fcVtwV5CXEHa1A62eqZj3O4R8rh9P1QuouadR7uw0ra4bW6Qn0WoLhVY
+AQN9kq7o+E8xPCXBaqNJbdc8aMfvgdnQ2FXcQdWSXryNdLSCHqIHlWxFKzQYty01HZbsWVIRYSj
CHaXTTtuEZHgpv8sbgMPKw+qxnTiAMMWCGV4MBQgkSB5qebg2uofLPEWXbKQhS7Ejz8/vpK1VtbX
uG7EZhPIPSajqVJTdU57Hdn2jMxKHIPw9Zaku/JzW56ygOCPdW6p4q5MOGDvzl/MwTEegGzDZm0O
3zam7HBf2TpKTTdzIkngGYGMJc0RYwtC8ibeM4ZcH5xlsrSjMI6/wAelDUfkgQ1UgZIdnJ7KLy6V
KR06tB8sUnaro2VAs48u+0WmYAY3o0qhTP2e9Ny5gQ2l0wZG1MtFH5dqnFeD2UtzfF4q8pdeX6E7
SqXazdJ6av4V+lWsG32M3f9z5iIY+QChp6YUCreJmPoO27x581jL5vfP/ha5liRC9qzHZoQLJO81
67Ic39Wcz+Ar3uAZdRlBmVToljo+Y8gRSRCLJ+ycPAuYl6WkO3rDTNQgVVoK6sPQuZcDyAlyo8pL
bUFuJzqhcj6rRpowRXzxQzUFVYiLEGT3HI2T1Mq1U9cJgZ68V0/OEuzhAdLiB2D2v/NFaWhZMiyU
pGuFyFcwQp4mfVCB/DftyebYl0/vsad/DSg8bd59hpdWnUkmuwI3p/49+abO5ySBWRw+TjeQoJiQ
IM+f2nCJAPVnwKk1idFNYtzOxdvrs2tqccCCIzjXJfLaJ1fMjzjh9oHcJ6tSja64sffIfzK5xF3i
iZsX2WNlrVD60eKaKhaqjNyqmQxpiN3ZWmH6Mmke0A8IHJl6VdWKu2zdkE/QFQyBfuvXijniObNU
H5T/xHSTnX5Ei1/uh/TiH0mwtgpSPoxeJFKoe4hD+YFyT/Hq3KENCQJvBbc/QC1lncbIf8oXm/L9
RGIMR7Dh0Xtp6RXlsQ4GxLtYLUUu5U6Un0qYiua+L/w9jZif9yRHLMnJmql1+AAUTyofP9EBlBt0
IZo2YbynPdfMHZHU/7maL7auIFUPE2Ro1awhKhYkxCIS7EL2lOpMKxZxzXgcX13R0aOR0B5Ls+Em
FaFIbrg9pg8fcjwwsj+tkxULcQjr9xqy/zo6mmPsJWrkak0quJ6MUYsEzuux+CEUus5Z6q7Y9pCv
xFfx+6fpPWUp/y9SXK13GMDsdvytCCWJfjir3SV2obPBdsbKbjCn4LvnIVuQkfGgVNE3NTwwGR2e
AZ/lQB6+o88101afon3eiePYJUdwkyg4y8utxqEYDkGfLSq49yeQxRcxFxhQiz2SPz/e+ReQyC+g
5e73981sRjDGcw9pYoTTliPLOhD8i/gAJr+xEkg/SpbIxm1r/LMTpMEC8Ru4FqllTUvZL3i4K9zD
6Qp9Ja4YDXRwiOmHljlyA3PyzAgXuZMNEaRbqSM8DTteZCJKKEFNxaTtVrPb4Szcs+spNIweCxfv
/Zd1QN6/U+L9Aj6vAaMiiU5JccrrDTkEf9KhDLvOJOMEHgMPla8Dgw1ZgW61Yp3z3TU3A3ud31yl
2dbb344/LAJu08nJ3vRtLeaOoeroqvP6SsbgGj5/Ek2zeEItsG5Ri9y3Y10xlJUG8x2cQ815mvQq
EJQCljWQ48+8ZuIgL/yq/KawdtxO7djG/jgLhnvCdX7J/uGvrBfKW4W7OgM0AP2Ch92pLvOwOYhd
GpwzEK48sVRifIp0kEKBHXoheU7Oi8Pjdvbfs0vYJbXLBlv8NHbXGqMXI2RKSqFxgbKsk+YYFN0q
W3dfuBv7tAyI8l3HiuEo0rzyBNeyLk72HwWPzbg4XOgTjVmrm8MAlwpdD0BN0o49MgXO0wvqUwKU
RktNHZ63aHMLfnUPOmBkQ9JELN+T/YvMT/+eCPxk2EAVlmaa2c1V2cz+58iwol/TTlI3Rqnq/NB6
0VHzIbRmWBbXxHwS8WajygCy7ALV9OLTTQenHLzox4EpX7pYxjmLN5r4dnmfvhfcba4Uei4annul
6w+42UPK9nqAXnVd8yRck1tFUVFMe/5hwadbSod087/tERIOMgCU58ad6i2Cqi3/BJA8F0vk7ouM
wBpyrsLv1OOuPyLN5FQHKtUqKTVjgR9b//FMijQx7nKLa2lBTtck7Lat/rJdfPOesTHJMOjwfr0O
UPjh5fMOeZK5s4l4LfP2bdnD5HIsxWmqO//i0WXByWY4du8sGJuMt87PoDScpjjMwzqoy/vouguE
rb4hVp/xdvm64zKgy+UeNPPPBgw1zPilfvY/AfW3BvYgg1D+TTxSlN4HHqNKPOl0/cY+EyMcR2Bv
RVqwWzqR67pr6Gjpwrq8iBNTIpIOPlvF9Mf+hnmV7+GVNlxdznks9iGa0IRA+A2iYRiOAYKCzFWp
+AxFSuZebGmSswuU2dMINLKaYv1eagi+4ZP0HtknD14LE3x77DLVk1UIe8oLD1NMY0VltHPbRRHi
5132f4tp5sf1o9ipkhQUgWj/bwghoedW6+GwJA4KOsjWQgxd6pzjQReOkTNFjO1kyhJTt0pQF8eU
4MQWleENbERcWARJX3mv9WYMvo0/Vd8kQhpFW0w2NwgT+bcVaisiWIYzay1jPlPefHiHJda4BLuV
08umyG8x+3ZLrUkNRde344XCSxhH96ALc0KkRC4mjZrQi5d6ktJzLOLW4lEkSl3qUBLTi6lPCMnU
lIBs9+Y815ZjATO5Ahg6Jro+7DRPlEp4F9KbP/2vHvOwjutYn4AbYDCr5GHA56A5KHlGix6DTNFq
SJL+janiFIJ+UC8oDvPgMKfpFx1kXqaP23W9hQ3Pia64dq8wgTr7/d5dX520EkMEfPxM6xhBcCXq
QNxeh3MAVu66ETzsg7f5XiCXFG6pR78DCTQMxQXArUVVIg98CEkrXA4xwHndcbf9EWkjHDDZ4dV5
VHCVkHzwOa2mPAQEF6VBBAmw3HYutW67kYYQ3U5acf75d15rblhX6CwJzHFCsl5emh+Q5VWr9uOd
t6/yg1wJbxMv26kBJf7wwnd1bZ2Ohdx4fOn/VswVA/PD4KysJVpNziDebLYyNHlesCJdXmC6oXz5
+/z8kU0FFgiUw3jFMGwI6qx5KmJoRxVUhGnxc8o+ZNZ7Dn9ycQFnjX6Ywx4di95f5k9VBBoRsW+9
OtECekbp8TcYO4jVSz/LvWqhEVU8A4qlmVMFX5zWC2qq2XRP8Tq6lvl8uF4Mf8vWFScEOUPJjMog
YR91JlhqvKNXjzf/QRRoGt8IID6JHiPp60j9Egw0GsTbejL5nv+bM/YkM5IboVuFr2xveIS5HtG2
a/2x9dFyiNHuLni+hYETr3iM3k1O/dWLFyye9eR2xqAsR6j8RvmjDUCpBCYHDiHVXYZz+IMmIwvF
bUXFj/u9K+zWgVkmuFRe82LdSrMzf4oj7aEo4acZhdTwZot5LKhz0A+mNGFaauW63L2rN8kVytWN
fCGkGB77GmF+hlG3O7175IZEW1LX3Vmi2jdtqs03YimbRBBtCx6dFu24EwWU+pHsECqkXcWGOXrm
YURNn7I33xQe/+Jp5zU5FN4Xi5m5v1zXj0iqmbVhZOvJNnWa4+7ijWaYWz6qg9ZjROPf6HnCrY5s
q9LYiOokcHVTiIhbx821wO0BimIHxMILVjGJCCkKTLKGGSZRlYqcIqTvXzauesoFeaKMZAxO2yn7
JPY6SRjBTfQE7ki4PKeXMAUJ/QQD7KMdqNwTkbVMOIiq3/LjvXtfqbRmBWfN3aw18PuDzkdVk3Ry
OdlzibT9xwoWBI+DP6lyfHwesHGnLPZgwN9QNTlgzyVjl8+aP4fyD3QUhfwS/g/OAP5n/cjlVU4p
NtYAkZCuv1+p5qTlRn3/8qH+YXGYgUQJz2sUkT//w6KAmhyBP86T0aPwFoSL5zqUn7Ucw39EasDs
HddzLzjqBvM+ar1gRJCgRgn/oxV+bdlFmQw9D/W40VAXzIAOBz0yTgvmVvcFZDb4ypWlxY5hB/l3
3xlPlU+0ocuxk/ccpStaDJG5pC1BvGPHPsZjbV9QZuxk0L0qLf7bMHecxgJKjyeUyx5VQ1dQWxfS
7i6U/Fynu8d+eHQN5WJClexxlYRFMEo7WEESdlZIyrwegcnCYgVXkVP1AxYfeyCLQR7++nH0CrCy
aEF9+AhcXd+ztS2VTsdulX1Q7Ip4Az/iJwj9VJ5Ybb8xkWU4h3mfixKdDxCBTqsdV2YHjmJomyXM
vtAAS8GnQnmbBJac24DqH92Xg+bHs24kxIhT0FLWsSunL3ZAttnq5+scO+ARuR29ZrU9klSV7iRq
KMLXfRh8wdzws/m1167HVKoX3ClYgPlC86/0hYm4VsfLtjDQnVK4E34wiBrHPpP1va3ku4kjEY5O
PKUkGYSah17w/B5EeaJo/GESCKM4SSYUnBS6wFPalfu9VSxAeTKqRbRk5lwbjIBZ5t21MAZ2ffsD
oEk3ggWAJH1pX0WFAbAU0xPS/qqZE94z4CxtTCXenkPyvaCvX5zpieUzL+gw/aBOcKLB+amGWK4b
sms6MRQ+Dk9Eb/oRciGhvA96wQgH/e5g2sOoAAMGMhaKZGh8e0sspG4QFE9XgqwIvJE6LeAxvoOJ
SobCdg8OfbOwN2PGIn8GsQO/HcsXNkmlkbGnPUtqyY+Ri5mGQ3bDDcGsSC7EMH94gu6wwijiZswx
9x0hBCAEgqyGLNfTbfhpXZ6gehoBQvNdyLN7oSoUYb1ugd+W2RkwWlv7CGkrYZqiXG4vKHC3KiMR
xPE5qVp7GrkxOUKFRlNZgWU3lEG/ubisouSn2u2qWzeQluq1AgNmEHOIOjgTfoCfJpaDWvWk5fI/
AVFKeLp0eOBnRwhNnmIE5bNDw/f//jiQgoydj+82qkvSnesMP5ie18Z3/m1oMfd2L1EOTormR6qm
ZLIxbAsYQI9GIxUrfP5mT/9sDuy9saFb999BNZd7PGOQC3lV72oiCYb8HjxVWx5kawerMFJ15AMa
ky7EMt+PVBGX/UeNcYQIahz/L3lL6EaokZYF2gSjcsQVUn3ijbNYIE9D/JKHS5y4tIBOg+JngFug
GF7CayYUzX2lKYXGsG9zQk5wtn2dIUVXPoGe2RcSdUfLAGP/cS0ZEMF2/4JRECoOQvhaPRShrUS8
LXFtV4lPpfBLXUMdu9JPdZQ6sLApHISdtJoTTWyR5Pn/ZQhyTUst9oOiPGx+urYCJNUzzjlzcWpH
wj3GfFISnHX+Az7U/dQHQa1h3QqAVnnH9RextzWXJ7wBOZyYUss5JKYslqdUm054h2EkSbRuaNq7
FKPhid0LrY/B1jttkzvwS020RND06E1JtSJkME4UIH+fO7MO4qmtp7qYKKQLUTb1vpqnN/1eIDR/
aE9L9slvbe5QP6ISyQF2iLWYUerXdcdc1sDO7bCrKdzVK3x6i+ydqVJTqzJLr9b7/Et95+hUSHVl
y235TW/E7TrqA9wMsKwq88DrbSUVh1Yxnaa3YkO2lODkmZnKVdZwWaFZD97o+Zv8eW9Z6pd+nt+I
SoQjUDft54LqnNcOo3yow4F0PovvOEEGK/rRQL6HhVRyY8L6xWrtsGsDtT3bMQFAVWWn7R3BvA0G
h4xoqe0viJasnknKnkSmbbvLi1mSCwC8yn7EGQRiC/6LHlAdId3tPcFbwHP2ytuheM8Q9qkkbeyg
sjRergiUsn1+ZT747sAQ9xopuYeQu0TutanPFsrJ0BC5kPTYAO8CbPwLnfZG+CbU8UPuvX8VUOXP
C9l7st1ZnrBF7oFYltVp5+4ruL84lulzhJI3nbpJ2yJYpkcurHGHAalN1Knde75FqlElHPAj2eWH
pwXP7b0ZWGeWsVfVCxo5egxBYHNUVyxmxM2c9CAylmsc427ojRKXuj3KImeAFqFxs5LNOMbohoJg
w+H/wcTgcFZc3rYr9QRwjhxn1JraJNgCYqCsBfSd2jx2HbWOSPByUejk8p4o9C4H/IMNwLVl0VN2
ye7RQpE+SHIBM91K7XFaDA2gfBQZ28gOyL+zb7xtzIkhvt8SlylpugnbsFfHdDakrFdUiIMY8BfC
QrRUpBDyAde7LHXBjFMNd5rYyDVKToxtJX9ih7J5pmxx5oB/11M1Mj81CnJmIwGfQEWzaobOWJ2r
LqBNav5FZdXEnzrbonkPA6jGLDbjkkv9mYEqQq9XlNnvoK4sy9BSjbGgSPIHxL/bTGkZS6phh9ld
wm9X8HWBLGPUdbRlSNmHwpaJyPTsjopz2xJCwRCRiIJn8Kgb4gTj1qw48wJnZkxlN60yn19G6EQP
EwY4XTOFbSbAkeK8VieOgHSSvFw4iwkCD1g3LR2eqOUovHw2ILeFK1rlh/SRY4/VwHlm0CTIkipy
CjwxpFdE8FVNQyoUkoiv1Y7R8yID+n8GIOSZctL8cWN0P2rDEkYx7E1QueZhaAL02e3L1ZCcaAlA
WD4biVpb9jdkzL7iWTfXvdAWRTFllHYDShM3OmFkwnQw6XrU+0/aNRCOUJZ2KgOAX4Yi66Mocjt/
8tDX1MDXIOn0mAlkPlxy0cE5ZTFTSHsBJhFY0u+KmTEOsD29egqNq642J7gAbzOwHKdKF/MzZmhr
c3njyobaBfnSdZGWEIC05/Zrx4dRDH84pY35TY3lqrq0EJwkPPQWHPz4GLU7pZ/ajgG1tHAfBqz1
x83HqfMod3O2KKKEgTYHL2fIPaC7YSElAyJiPRg6RrOuB+6UgBc7baMbIejCJjMUDXgi/puJ7y2E
1pYe3z5FZjl+3GFaSstRzJH6eHZa+PfQz+qyZJiAbRKIh3GbQiw6FMpr1Mi+vrckGmJufZhPJ0dJ
YlnyaIrEzu6KxIKwBM3kUKlnLupRRP9s/sb289DlXs4wh+In190t33ntoEt8MerkYhGxQUPxO4Hv
vHg8tdHb/VftPOuPz4QXOnWSHuAUaoo2j6ndXfyt1NILu3LrRkk9CZ0i043e3XvBtuW+Z/xqLb4g
XdAzZfYVokVWpkBbtcYEiymExvbKIMjWt5YnTxzqG4pvCVAqhPtnx56OD69q77iFb3I0JE2i+Cy5
J1crJP2RIScc8BmRYf5RkOUj6jydQvats4wL+5N7/cOSSsiu5mMFOmCypQYoPQDUo4H2NdNe4O/f
o+N+zW0gCqW8ZUluBagPsD4rw9uUjN38AX/HitafC9QET6ukGCglWKiiQ8JBnJPByRHTKgzvn300
24rM5MiAipCNSTIQip0m/7go7v6/YMseJZ0sC1SDvKFCGHl31GkUIVBfEHW6BeYs6T/cVyvej66t
IyXBo4Sp5vFze1p/b2GUrLEoOajVX9jkaDqsZFGMNc3U/qqlWE21K07/RbTMegSGRhMKzqz1en+d
OJWqxHKLWIg1UOSFqN0BiyXBOhFJkp0cUBCxkHZgpZhBKFaHvtXKQISfKOopeVpiNOVoB92FMvYY
eon5mJJxwIJnqAD/UvU3GtJ1rSoXGG8w+XyCScvJbXzK7t6DaqyHA7iLplad/MxKicRIHmtGElNU
65OEvA7Pwx5cNNVF4+AgR2htlwopYcIyNNLO+16y4W8GNkhj0K5w0CyZgwHpd44gg2oDvxBl3d1u
JpdKq6qBhSC7vipJM0/OudBGfb3wbpVt2aft64WT4i1VjIQFT6wAxVfzp8vrDP4DAyXZnWidxw+S
kqag7WO7g/hjyjCahnaWhdXSbxyzDa078xSET0IHfDax8tkkcVcKjH1cFiIRViYxton+thI0U7mJ
C8yUXF5qaZF9njlIgOIXfZIJAZb40No6pIuHdwOD8vT7Z6qurr7FLR1IU/w+2LJG2em4Wn4UTP7v
cJMaMaSI1cTHH6YlNquUKWbYlToQCPNmeU4aExp4tPHAkAn8gF4kJw6T3WZ903PO1792LgDDRKzm
px20hm7gDZaUbZ2g0grVu5LcrW1lcoif53b+g/jgwLAVFvK7B96Khn3eZ9ngHUUGn4DX2snqUM7n
mRf2x9dwqArzlunXhFOJpHiI/xMftySCUv1RrKORUb8dHOAZ5gMeCTtzEZYpGsrvx/bjUO7UDRbG
d/OCfRcSW81xOarcuxljI8x7XvzFsJP/DCS4kjc6RXe2WVe2aO3NkXp9W6aNxv2WCYPTE+PoJMLC
Set1J2dc3LtTFPJgs1YYFvGXvMOho7WVKvpwYP733GXkGMxD+JbDVrpNR9OuFLGYWlPdc85T9hSi
OwkACLo6NjePU+tppqZsPUnMay47LDVLsuPVqfnkKfRdU3x8xoOCYFE417JGQnZkmB7zNuQBNxdr
h4w7tBYZ5sc9ED1UgeiUzVBN62nCwkXhhzz2aCou8EUNsrHxbdD/RQ5PmZin/lNwQ02KYM6phYy7
kDrgwEzHibS2uLQjyIEcm5sAsn1EtJakR8ewyX7H3MWlJvtxHmP9tTYpHzXXWb8JH66QMZt8VD5z
WrJmE9QAVaiD709JHSmUQdL/j0SKwXLCHb53CLWPJabmPN6OJBx0W+6GUM2hjMHAL8dGfqay/z8T
jTtvhpuhshN6u26pIMT3gY9vgfLBaC62f+QP9Xe9wm/Rsg9ryWbdU8IcGD5RAHxcrCXyJQ/RW1R4
n/k1XeLsSms2A1rfftDlTyTZceOSE/PT10jyTV8yBzlrEyMH1QWECJCM7sWVK3cXIK6YbnKNj+Cx
INT8no/H68ts1iMIcEI4wZG9kPO7qlKDYsfOuUNKkqtAe7WE+J4amfXLE+R+Dm/rEUVjW4EzgxwH
aX+fHhpa38yAipZbFWZU5CrBXiYcqorAivjW0m2+Tpr04l8yl4bbmZfJ4xIt2wT/UnBPfXYvt/R5
T6RJpe8gRBUQ8IjDL4UgF8XfluGzcCS0QFvZUrdRFF9gAotjCfayf+Csm/H1crG98TNaw8xPseqV
nEYzaHO/7ksKfhS7noHk48e5DHaxZ47wz1NHcwUQFn8zOoiuZ5XQuflZNB3eGZtfdvoA9mTEDejy
d0yGUD4aOjQCPDOfafsEg0YaElHWBuo2OHdG4iVbMtjvPcTZXJF8cwCqLTT5Fcnv6WtLWLaF7/ak
LF4l4fypO6LEL6aNW3SWrjUQv/hODMrX0myDIzc6RA0syn/eyGz+UYWuUguRttXBgbzzSbF6b65g
nMuByAuFExqAU69/j7jCnspk6ayOA4o311WNeyC3iWxGvAm3AhTSoG3vDmS7e35952yrqUI8her5
DXJSi7WeCa0eGB1vc4y98NnnKKEfl7ZlyA87WS3/mVWCgIMBw00cgq8MUES+Eio5tWcb9tTA9Gfy
ZWhMLWTGiqJER1tqx3ELPN3LqqJIpSDDJtpZVfgjujCu2vOWesNeFzq+Hitj/9HU5MBXYhGEkTQC
kMFB6w/OqBl2KBkxHoHgQofFgmVGXmKWVb6u7nsGtfRndaZhSYzqU5GS6Zv+mF0qSkByMSAJKAlH
xbKsrfnJ3wgpsQD4+LVj9xw2tEaEO0B6z4cwpwU8wHm/tzzegszX+3ap2z5O1JFE6hpB3Rvh2Qe6
heuTJiObGwg9IV/UYo8Wsw719L9sfp7435f7LeUqf1zRpLHN0WhGfR/n9PM/6lBJENFNWvkAf8t1
GENpYtr/I8ByyV9vz01TO0BkjgIuk9zKcYqVizvvaglUt2qX9blUosu0qspAuhewKL+lUAJcanBy
uzR1X345MR6/PJitmGCShaXJR//OvAyDK7gAWWjzuSEbTPYFyjEWB/6/mViRh2Paw++dTEkk538j
R6DqnL9WStMC46WxX1YFEfjXIr/jlB/p+XKu0rVUf/oyJKS64y6r4C5o/tj+J9so2WYlfuPI4LPO
YsaKN2GP1QW9DU8ZuLLBAvOFMd9QMdcCE+7askWEo7qiZ3u3xCl6igBf6J7TBrYqGCbwlA1adpGg
G45H4O7Bw23WmOqMlzpRDEZ2up8LI9hHpuQvjUAjf3lnuiGBA35AvL831zCfnf9MmcQ3A+4UGcQJ
Q8AnB5VFD6Bz3CdlN1TlPOFPvKjxZL0wBFLuRkuz24KizlHJtUA8PY4S97uTmZQbMUoWypaVGAb3
nAtVlxESvdPKMV89HJIyuspTN2vaBYF1NASBlPg8GIaUVkGGHTy3IFf1X4QN4tXZB6YPl5ALMPdy
YYF2g2TIFsvuzzTPuN8LV1qY2QrNkzfYdGYO3KGzMDRtBLjqHCDaB7vLUy+k5qHSfnkNJDa9fxLn
ZwAn1+nBOIbLF2OUMS/1HbRCPRh7MnFZoP6ImbXXljf17SqNfIJS3tmzDeT+V8pF4I9PRZdiRFoT
sN3o+h5R0mM9u+9vuk6Hv+H4hnY00DfzwUWEGNb20KJ3gw7VxR0VRXlKJ3fsCtTBxmY5t0Lo/oaa
ZqmMBI11SZPJvDNCSV3O0ZixXa1zHRR4BGFLIJkNQxrWv0ak5713R5A5hmP14g79YRtTTvLsIcsU
1V2/dNnJPjduE/Q3aMVbLOZDwFU20bVW/6f7Nd1zT/cY32L8Fy2jXHNgUongZe4BefjbuBf2KBte
EMYMGq4gxFJF0UFg5OV4cmA0S8SNNV30u10cbiCWtvay9BL6xuvXefbMZi18AZS96bktRDCHsxJU
1F+EskutW9bBrZckqWg5D30EprEQvJX6hpJcSaNoC3nm0a3XaakU+/ut66kPnflWpde+SY1DkysV
TZ6lvANSmRBs+eUcNZDxMEwGJEeYSy+CFj4CYThXJ9bfmjBO5SAgVEFt7ydvDFRIKXxmnOzB9ViN
MB/WkSIi9PMJHWlyddC76pO0sSWFiqLBkrYjA0jkEGhXkV7dS8ug9PgxQa4BTFjzvoccErvFrhir
juDmLXrj6oOuXeYMArHk0DO3Rr8VtBpxyB0zr43YeHBNqou5avN/lMvZRkTaeMHJL1ygLVgmtm5n
xp8Q6CSkLgd6tQqMf7l4kbIHfJhBMqhJ2/6BadaIcNNnjCBvgijf6Rw6J0m9WMO/9IUd6FGtDTyO
RounbmIPNqRGWnxOhv0g0S+bsSkit3J8VxvmGz0s/N+gmpquAJPs/0SZx5CK3zj8Ux1Ht+cg20Hy
8tfrj02WTReSWxszazGsDmiyJ1V38eQVliqY908/hDveT3Z93790SUOk9qt77/tO5YctcIxquHxG
EvrWrI32iGYt/ByGuz6uBLh0lduC2rMvmhP86auB8LR31sNwl198YmMX6Gz1yclaBM9niGSxsnZ3
aXtHLarVhmU/DBU75I/ZsFq2fvVpiMkNCXBLLw6gUbYfwVMtuW0bwvWgbGfg+j0y9IBvNaZo/xa6
MssUOtD2TJPPlxE37PeFgRLbhU/EZ26br5AYZGoN2YN2YgnM/1F5yB0smGuXPkfzQLQXo13vZADM
jQ0wVfxugzr6UZfv0QW+9odhxOtSIExEenTCgnum4toWef39/kNY6KCGfOaWpRua/BGme5X65RDB
E67ps3nJzpWHLe0dyBPSKQQ069WZARHwYVsP/RxYtV5wvQmdLI/TkWUSp3qkgIS7lBHqGKWE25r4
IA/xwPsgQE0ZVGsuaAiN9MB7yZkxe/moDBZ4KVSvJ1huBDtzodbthqh3fxxPCiOuDSgp4zOMNd/i
nctTfSlhPCMCb09FgbNF2jT5sf4zSoeQL2hYKPPmp6XjNR7v0KnnrwoJWabNaPZ1TR3fEXwd3Ntp
tDgTmvDpbY4SZfRDDJjX3cHt1XeIGWF2uEyh7GhZ1SLMvpRlPbOzHRSFkQrgaq1d8xnOI+yt8zdi
aIB1z07T66WfVmFSrqd43K0ejtF7M7buHyvinwyuq7H30Z30HrkU7s7c3UaF1Dq4wUNkRLnZOmiF
GlC0DMwwfuldqg7nfL7qV3BkkU9bOtWCGU24JsCkaFftDGRX9u6atSwssTJe8A91ZcvBeG9FZldw
mTEI/CiWfFcFwjEkPWIZOYk/Pildvoe4AkdtiFbuJQbEw4rffGUpZQ7uOBlVsJSthapijMumoVOq
XV13EXpQJTJ4mH5puB0986eVBp+dIV1BO69S24WCfr0MYPGmBDsHl+PNrLvfdcKP/JfitXkT8Ndn
Q9BjnqeabNZyU+7WW4LZCRUE0ZLpNm6Ocv8blkk2yH0+tLZoe/TRTQIADb5XFX0ZhA49qO1mrcb+
By+5svGmo9KU1ewXsoHyQKIp9nwFJv16mgXSExvJB93nCCTfLMA5FJHiIVln/+YDB9OdvBSDWDxY
OPL97DC8ba6NXTj39BoW/HGy0PPm647X3lkghMbl3JaD/63RcXNFVZSWiX/Q++H1/grvoZDXfwk1
UVm8qT1QFNmPgNaxdli/uj+95FV85DeJTU5qcGl2t/41+Tm/1C2ybEh5THZiO7l3jMSnHt7DmBb3
fZantSQTA6n1XSb6t4qmf+Dyp6CMi2TylBl/BTQ6ROqnuk4SIKsEsZJY+/Co4xD7c4kgMU+DH6Cu
busvlij9uHsDn74Bsb5zsNqap1I0VcXEZ5oWPNAbAZb7wfqWzjyb2hlFnTF3mUxYTvx7pL1UpCZD
TdZRSJ5BHPWz4F2vNCCBCeoxq47i7Wy+c84W6CyrnXaHJTS9qAbdrHDtV0ErergqmB7OhQfjbvI5
v+pir7yDftu6KZcGGjvr1sCBwKDin3usa9Au9AUGbNCH68SWc4zddovbyDiSn8+Wz2+82Ki0wjPL
zudUp40XCDDPSbO0wNGBS8mjoQ+YXqb3f5PgkVrGnAbfCbwgVKoEaJcOSMeN1pbmYjqjHxESk8kk
8CU6h1EFIbc/wWdaHG5CZznZfmN9ZrepemzWKnGDnq4fRWYp3We3fPTnztbcZskKGEEMoYS3eojn
R2rChjl7jofH5BM0X9ISYehaI9nd3krJgxzGGRoZ6ismHC0DOdhWG0hxk677Z9NYPNcvQhq6E5Kv
hm/s4O1pOI52ahop/EXN6PkwbNFdRdxP290r3uSeBrk0EUo7LzU5iN59wBGGlAUd3xPXw3rOIE86
UZeXjrIW+6AZw21dwqgQM54CHiFdrSd7GvqhpWNqMUA0/L0hOzCVY78zjfQhlAJI81BMB8kNgdPv
3aRALq5yFoJ3vsdhxdTXj7t1DyLJfdyprEfPqdv2UtNDaRxDoOK3SLGXRf/WX8EEPDxuoViPoWts
fUNqYtl7aIWCLew5Sf1H/h23/+C4sUVjluDfsiVhCmRvshkD0WdlpluofJq2VPNYxP/Ny+P8VHIF
zVSzqKM5iJIoiHf9rvluiAmqBtK7lzxCRJPrzVsU6pqqup7aYCgnCp7cp7IqVe7niZLZpyr9egV+
gyj+31bom87trFZmT46ovtqdzh2fn1jJvG/suxtuY7L5zKfCylZQIXCDhtAPH4OpTDlTA8P3/BMo
qL7f6Mz/NeTs+QHU0HU+hzbr/fnglnOL6d84LySG7iZr5OXDIAo+CU+zAUeSPfwGSG52sPjmWJkJ
nnJggDk8MaPn+xbjHIpXuBynIxmQtodzjf65zi8bEAT9E3okit/lyr00xWP047dfc5MdDANfp0dK
JG54KBrCi5uN1fYHyJ0YY6L24rv/HVcxIzkcEP5m3CWoycP9FZ4i2GD+sznL9MlJOhJemMArHkvm
Jc7TA8u7OVJ3y8ZYGI8DKb9OzXDorkacemAyYKzb51KTFWq3b28HXzcoVrgE/cbY0OwLcfwsWVlA
EZY9/8KN23XsxtEn8/wnpqmOaWvBcri5vS4vppFOqA/nDhDdWcTt8HzKFzmAaMYE0zrpY0HKbeiJ
8fQ0ncRjYIr7f8YiGGw9IcnqhCuBqIsleLGTO9U60AuG72QEfm1fQ8NL8Z7bZ7XY22nE4+sYWhMb
r8YXYKvkwN1iS1ko6r0noLljmus9fW5mQXXbwLoGaukJWxCNXPU0hpjq82cxg7QCwEJvxaoeixpi
PV2VVt1rjpwDCSvhXCbTg6SShtsT2Wlc4Wr0e9/OYZ3DOrwA6QpGX+/yX3pPfLMlYOWlggqkonCj
VToiz1QHFU6/hMi/q/lMCo8eMH9dRxAD1yPmb+DbwDw6DMDU/8vCMfJDQJ4YkK0cuJGWliwEsqNE
aMNpX9ATTr7Yf3lYECmA9+TRvmMjF3qq4rW5bbsGV62SIP0XZ+DeDZ/PVsjkKtG0K7vZv8nwIIlg
oGndKIEyWeJ85k6Dag3HWTGqLCwtt/Pqwqe1hV6BCoWOBjcP1o6HbCIoOzZqO4w0VqkCZPH2XOvw
boSvrI1WEDvDr45D+qu+H+g58EKcGA4m/6Dlzidrc8KM6ONuXzR7Inb3GRWHNF4i81XXPWxATAWd
ABiUQz5EXD/WhtTULsk93oIdXL5G9WWpUGlC3QkYFgsmaMAaAesB4Mt0JidNIfjcb0Y1itU2tqbp
nCsNF4x56A6e3Fd+N0N4UmTX3ztCNFpgaKdqb2suTSNUOq68Vl7zjNEc+bQO+VEocLCQfWhV1lsL
IY/tWnwzr0HKly7/eFjllvTO5zpQHdwxx0UBMyxlpLQWenxcbwAv+aULTz7ACpNsm/J4/tDel3+W
KQBipfmfkV44Im1ERPwC/WOqkIB5sd2wW0rra8CEBvRgx4Bmb8UHQQAbGGFEkzBcHp9KdUTtYE0D
3Iwa1SgU5OGppq4/fia0+agJGPr/e687G9J5FP6S9hm1H37+BvKOIbXAuNO8H/M2VUXN12ppA51U
LzlHbmjuhI3PUq2zeO+6RkBhmtAQqVgyFmW99K9GgHBUTtGf7+/tiPe980DtRXZayDahctd99eKn
hDlRUc1dza8WmPvSOIL3SffS1qxNazUNUJtXxU06fbQdlH4s2qHFAXmzUSMnvCGUWIsnb5zdQlAR
JTwZf07+maUv3i7NaSHPApfWQDFpP45HkqOhRHVXHuZjtTmSfzsBxkwtgaChZ992chM3msS75/m/
KY33b+RefuUaiKWLhUx8UJdx8BRh71vmvUpj9Y6H5lVKODT38VtIBHazWa1VKlHjRQrb9brpq776
t7nR6jTZU7qRfQIp7dvIgV8zRuZ/1Qx1EUXdxfbayqHOJjZBWOYFK5AWGRKeJZ08nZWAXc1EHGM3
d6d9TLq8su84hE3E/2qwlNJ4frKf+IIQ9DCw4ExbPLagG8ilcqIRCwm+XB8fl28/u1xeqzlRzKgw
NkPVRVIWAEOHenWkCrFMxwtoQLZttm+nXe7KCOra4SkJ0UJistM6SXRBn0iUJcM5ogkSn4gzKtbF
+nHSdG1ODnmUOAAUDGuh/Q/N6QaB7DlwpALLuPkhp1unK+RZhDOQL+hk4jLEgMo/xM5eNAjHAp/x
+0GkslqqpF0HQiZSd8WXy3jdgcpqbMD+cUUhbsJDCBqKzhFDumB1x5+QONPnf1qAg8a5vDwyxmQf
O5tbBJnNHL/yG/VJzqdYbjE73cWiy/+vjSNbfepoeG1eXisi0virakkkSqXPWu8ggCYsSZJGSS7/
tqBjeVorrYi2uQCSphQAmUXmhKdUqOCNG+HNtQhor7iZzdopwGmZV/1ukaqNX5iXqntdVvJAOEeL
vGDp34tw5r9sJVpGAG9nUQQaGUkoaTcT9Gv+qkCMFK5+ziCDfkt/ju5bVWOZmNdE6mQd8BFny9nx
y/G4BsR8mIsT7HlFGvfNC7x+2ZLUbjvM5SR2mOnzsV3q0pYEsGTimugbcjh2DTqiR51VaWZWJZm1
CszwINsg8fACRqdsWPdvbJoIqQmaAoZT42HWMV4tYawjeEvwoqV6852zXC44ZAtM7epiZA+7l2xT
w/Ai1/Sqn02cGJnjxCNGn4T9jPIDsJOgZ2bMB1oPapa+RF8ij4LM4WkkVSARTMybFw7Pr8AQbT4O
kSCGZ5/a7FP3FAhi9joQWsC3cxB0A2VImwwJOGEUGoCy6Xv5VAYUAusdiElK9bu9cEn+OcqggRCT
lpl/7+n/zwX/kfmsftxv3ot1K3SeFGBo6C/jV3onuB3M3t+z7BQoKHXxG3wJkd+DPhkrSZJ9tG8n
JopU0uA9J3LQgpDhG5KpFb9Cz6GwFvyNIw9h7RZJ55/MCFYr71FGE6pZ7KBDfQMIrTb34vJ//lOd
lzFX/hAPCR9m0ugDhcd2S0xhSVknwODzBWkMM7/bH56kPHz3SeZQ913qlKi7P1qP9LLsScbuQkeZ
WrpkntbPhrlyS4qhdhRCuZRfl9drIMNG60A1fQ45PkKazaiHT3qzYgKZPd60BLv8ILJJsOBLD2rS
fIHtDvRlUbvueFyD36rVnw9KKc+nssXRSamlGRFzmQdLyi39BeQQRd1eoEa3A1BtNRwz2lLd4zIk
aMz142EH/zGXN0m4E7uu4+nJPUNdgQIOLhYn3H4RDUvR5wlpAlqdK+3+I7yQG9vjas2mS/kJsBLX
zALvYdZ9pHQ57DSkcs0aW9epLBytg1N3zptqKRG0BRq2QW1EAZQBc9t72Srp1K5pocQ5CQfsGeea
KaI7D+MD+9Nh4mUIROvvwp7jp9yI3q1gtIZbND4mpy/GgY06F4dpGnk6u+8BhPqn62U1MsP72Wcq
04uuqxuTlzPQ4pRdHhYEIcsm1ka8a5sh47nP+ndYc0aBpGTmaTuCccrzaK628Fxj4nG1mjs+Mgr6
U0uAHPg8JAnNggbtPUidKiBwsrIjm7mKsUueBflRzQJdCtltWQSDIaKru32OhEMxskVdKIX8H7yu
cPvT+eSSJkeelsG83iNLK1tF5AAApCQvIxzjM+QcHDEtrLVCKlAWFcIBt+AyJcWqz6M9fmTpbFqN
P/MDkg3UpTsw7lR8s5eMrXu1ebjVYELXSkXS0bhAP7mQMOOqgqED37VIC2UYFWJMDCB4dmA2CwQu
1hxXLsAFAlyULY4mcOrwo9nodOuKTYn1YU+Ho2SU8gy75KptSn8+rfEwfpOc5ZJhheZxp8gJ5ajc
mG+NOuDAYEEBLFLZV7hcv7DOpW6zVA6iN0tENcW40uVr/AOGy+vRGyuGRQvgj58gpN5B5O0dyUDf
a9unvnC/GrrAChkuv/I6dDvKhAV8/KH+IOhkqk+cItGWTj/7ZatrWhxQmEgV6MqPgSY9coBfeXlw
ZwdyMOH3i6GrRdPaiWa9NcfbccIPO9RwHXAwWnsYBI0+Pct3nbFhYslcrQJGLgE2oPyqMZe4kGSP
NUeAjsE9yER5ZHgUBPuN/ESfs3QpYjgIX+t4POwp9KfnINnNqe5UraHDnGIgWP6ca/SXIa3H2oXT
ilFxEVXfL+ZRiLRZ/+ILBQ3Q5shUuVI8xtnLTOmoNOP1W90Bb9idE7n/3m8tp0GdFUV1WGVqprWb
w+XdW2JgQUnLZC/+yWim8coq6I6c9n1cR9NseNaRFro8pCT2GAlmd3oNHbETHRtDK2dQ/RuiOX/H
sWOaTP1tyiHcMCBZoaeBO3gSJq9t8s5oNwF+yM5Mp5xILIq7ybjXlK6xriWt8UfH032uakHwziR2
T3tedROsQ7Gth9YauDWGoK8BUyADstz86CPnssGDk5MH8pvKRTIdUnCH1PX1vzCt/i7u/PTRE4Eo
pngSXQ+qYztehc3pmLJiTMt2iBaCssPyuGEdDljrbYS702X2sURPmdEdXkhadRLNdDquHByRvKiJ
ceVRGkqSsXyMtUEZ38h0qe63eGf8HBQNjP6h/iuKVGmZObLvJcWLN9kKFNhUFvFCRArR8xXIHk8O
eJM5mZuPWeVjjJ5H0Kc/2yvkeTmKpVl0l9L2ZgDWMqAZ5tY/T1suh+oqzzyf6oGScUSQGgMtgQ9u
17MW3N33GwcLXJsjTWzZ9jA16PUk4G6zsHe2ICJNeemPCPX20HUuHaIDehXPBlz81Strroz5RSYa
kY1KbrxBGKgLyh6stzM5ThBeG+c3MpGc/qK7Axj0JQWOq/iz8O/CM/og3uU4z5xZImv+xkuc4t/Z
kZbTMGIMmptDne9+EVSJU2xJDZa3gjpQP29+y8DEm87PFsWiHAzVti3mcOTw94eREe5RQxBcAx10
E3iZ2sko2Z1zE+nwln4GJKied5P5r2WPu7BjMa/BUnMSmIMWSR1nePxO1dqeAjA5CHPqn3nLZv9J
OHkO3w4L0WkTkEx3yaBo8OmEIRqsnu1MFKfICgu6poEEs2cm8uz35FvaW7EVMe858++BKYVqFnmV
EETZobjgCM6Ky64MdiJxHUbyYesmuZP+Vr5MIVa8ti0rZVT9RQ65n5l8j68TUmeGZK/n8UspS43S
bMw1ixTHtnXyn5VZKN1AMQ6KwzaewkKEegjU0tZeJ6D2TZiCOmdWRKHToqS88i6mBrnzbbl+LMch
BnREAAK2IzDgqUWrR1+D/wrl5rJeDdingec5OiqjU12jefvS1V6Y406OCrWRbM66SJWE7PrqmBSK
6fe2nPOM8Ll8wlO/JdXPiVwVvrNKyOO2K5IimCLEAlGhxMTvZvO+0HXv9ooFdznPeLhUyy1YHi3s
HQLB4UTXlB6g3elTzlW2uTwbYQzobBwIo1g7HVUg947KZ0CuJjMvgjFwyhxfxiEpja9j5n8yx+Cl
jgO+Vpr39Kij2RslvJtvBj6MoGJJwRJ0s7mlHvg/TuoTBQzLElm1+DXslAuW1MIVQHx8xfU3/SgZ
ndCHZRNaDf0lQ3eAMM7+Z9v4bAiF7KnfPVRTledGOhlCOmZdrkg2yrM36DPNpHiDj/U96ZZ/8nv9
zml5iez7Xpz8CGyPVxlMwHHdCpLsIj5tLMvvUAwoEo4pXFHbkV6mqpbvaAh7/vnBJj0LOndh5709
RwFX2ODj94anMB+TW9v4JxA5zx3QJTgVX2e7zKJw0yVLqCAIP6L7rq++8jx6QansvH7M3bSQpuPl
oP++x7zkdNpQYXOUn3JsfOMy0j5G1TxOenef7O+oAdidZUIoct2f0USZOagfVZslckDxF5Eibfrm
T5RFVi/8ASGN1vP8zkkDPYcplelnGiNTiAN/57ynKRDiU4era4QZELo8yOl/vyVrR2YgSxszrG1R
t9pbj4Hjhor8nxbsetrvoJ4SMKLl1/iRuhjmidfl4CH3eoKytEnANGxSYdXANoM1/t2Y2vNlYyxu
+v+/KpwDpRMsoPnrt7tqDrlSQ/pwDjbDWQMfNb409o/+pVQRar69fmV1Bos6Ux7sdCZV/JqgLa2w
TnkW1GLutjF+vNKvTiMLxz00pQXI1p07+XDYsYb9sOMuiIowDxA+lZmNLvh4/4FpihqnbzmWaPRi
ftfS/utCWKLXIZQs0w66C/NYAPBEXAeAtUxxLIm7P1T60HqGcLyyLUsL/XdUCa3S7FGbUAQrHZTc
W8+qKjQnaCQrkb19hZ+ZyLx5mKt9xNE92vsmXNE2uedXn4NslEJzCWH3kQAcmnjjqYIH9dh9PQMM
rMlDZFCu9ui+mdFOu5DRU1Wi4lLhrs6NEgan2YHWQjBHBCHQ7vZUo4WWbzFFEBUNJLE+WdrLAOaX
sY+PyybuXorFX1QJAd9S1LRX46TbVtOnv5T3h96sDEzoXfosmXAQPyg1inYmleqZVYQJFvHBt3L+
eb3yO9XMCDlRYxMtSRnRhP0E8bfMR2UI/LvfJenj96sTlWrK+raW2sLlzd3cJBcJ09nHRCMoYkYp
zj0xpOyFQELJVMxyHKSC5U+jWERp2Q2QWf911NSbpyKfsAZx3TlhiOiaBpmqumvzvhUirjGEmZs/
1of6eQhg36L8x0tmTQrKjSyX6DBTNhKa85/yui1ZSzfF/8wwRKvj+1qBRqZlJK5s0bmI33AbjA9Z
VNSamrsPLOZ54OF2anLl8qq1pZo12bYehZ1KxEXgop7yks2FTq/SrRj0dp2TcDAqZUxN2VtiJVbV
XMzdukShR7oxPP+DqiAXdLhQdLR940KAQYjc4RBAVE8FKlT8kIjjlSehVxQjiXdsnvkNb4l0KNMd
ydxxWyn0EvqaVfHw33tlvVDFYzbU4FElbyiXz0hW1DXRDs5bB9Ch2AgJ0H11H2PAqd2IDmikPlJJ
cnJS7awmsf0XDFGoG0HAp7/0/FECdvf2YEC9Ee0NdQgnjZnt/M2VvsQXXUdC+wPATPAf8EB5MpSf
AyJSlm0qUCOId8aiyal4nyf2+k22g9J6+G/tLdA33OadMquz5av3ozk6c0xBPSWPJEq6GyC+diY7
hSUFl5e4ykadkelI+si3Xyfa5orLw1181JnT4RHYB4liEzn+LZ+J5RAhl/3Sjwas4I6fXFuP+Rm4
Bo1flCgg9o6Ss+jQYsoiT6A5GWB0H+0JY5M70VYICirwAuTOWBHHBZk6tWqUyaLbtKV6yVcuPlF6
XSZZzfwRc2B7UxEqTLZdN2jt2qxCeI/t+aoj7N5mrOz1vcnwJwxowK14wvbwppF06z6IGql2iJfb
+4AQ6t33o4R4DMQMT76wviZhzls9R9cCw5LCipKD9x2KHFwsPPEBWblPi20MpLSyOTlaG3IDwWdp
4mA8GzvcCST9Zn6mw71IGztNWxfTGTIMZrrivBig+ahtqAhLcBkkzsE70WwgpL1+mlzN1eHca9LE
3gyukHw7GGQDo6lxQdNeDvQF981FUvQ15MVV7lwCtHN0ALGS8wWmeyZrA2pHsPpKdW93fs/tGI06
cYBN1Qmpb/3/Vmyo9k5Nb1yLDahmupL0cAF6QOpBewnQfZXpBTQ4LlhUYsWlLEHVeSNMcKqoofZs
709jPNJqVNewhO70NEAP6VtoG3Hx3HdEbzjZ/5nJ5VjYDDgf8HNGQ8sUxlRnc8E3r3gN8HFsZXxd
QMTArJ97r9KbeWMn+Bb3LfzLPtTJSQQhDKgYjh3CL5R1G5cbAjhOM9YdE1KaHr9BGtQcuO2cranA
t6mbM/zhQxn4aOX9y0wKPCDUT3alvAItqzohr5cmNXOstoOMG3UOtPTshOgy1sR6GHicUZmpXyAa
TxQL96vwpW7Yee9jolRDbcCMecyZ/AZZYAiIJlojrderEKoPraDsFagbdczGcwy2OMxk7vfh+KL6
HjbYYMnXpPOKpCfjZQXw0R1C+0MsOmzNP8wK9ZFK3srT8Oz6iPYOthZXsaqU5mW/S7AYS1vlXFaC
fM3+Snlbc7YApf1++SDmNTczIufBlkpQYnPRej2OfC94U3v5lFWl7lqNmcXHuz48YK0aAbPdn1MW
ihbnWReu6vkBsH+/pwK6w/Co/LZ5Kv928oj06P2l+TUjXuyGQ1GkijhXAcAUGQemtQ56KjKWxawj
xy9h1kLulLoqIrHxiKgs6nH7L/IftJk1drjIhJmHgpJdiLP7Ws1Zj0KBWTP7U/IyRHdvpIY8ihKu
891lzEG79H+NYZ+DFMGSqThMta7g6LX1UDKRR9uiDtDYZGVM1EpO3rgSDHULJHIRqmIg+0x49W3r
YP1C2nBAO21OzhshHPDE+6RwWw7Fm0UyWdKDtVwYTyfJhQDMNpSkQllV14StaBthw1urcQgn6I9K
FylOjZhxB/P2+5DHEtqGkudZwjjPgUiwEWipaPTKJ7wneECT8pDcKmJFn+jroxBXRbySZ8B4bk7k
DnNdyJzKyG/c9OiZbAWYQBQhO8ts6Har/2L35lMswRV4OEmJxzeeFxyDb+4R19yokYWTCpJd6auF
+wxZCpBEfc6Gbk5SVzN+UqVLV8yZqR5U9IJcdodCtGUIsieSThfpPDRsstfGM789k3YKav4Lgn1i
xn7gm57Qbv3L8YMHGVY9m56pFk8yTRnRssP1xeMDUMbarQYJIGvsC+NCCsk/V0LRGE7rGRMRaU9N
iswqSXyI7WmJNZkHX2cugE6jV4QeMtl/JEqGp98qZLVHPeb5n+azNZ7RaWrG9VUYuKkhPvihGC3q
OA2FsKLdNIqk2iR4D73pIjuEHmTCrkUN8wZvrLMUyyga7plSX5DVFB86bc5CXwa4Qh7StZUHZhM3
47GTO1m1IBB90+uz+UpDKJNr2npzaFDtc6iYjvM6JIDCiZ+fouxZsgxCDiXYK/YDTOfxeT5lxgRh
BFB9KEMYN/LNE9rqKEAuHZ60tvdh1VakvRe2h/Gyw0MD0IWPYrPy52RknQVL1Iw+kVxhO8zz+2sz
PnELSBMnyC+Kccc7nJOM2tJtbfyelI4dtCyRJfKNrmMlRIGqTQGCFcqUG9oWGSg7mQmST85LqTtb
7CUb7IbJLrYu4TFei29c3Yx6mghfz7wXNPlLKqI6itF8/iew02OluURaZ6g73bBLLZR6ID9kGgwj
sqc5hDTlyp1+yRNDqhLDGyEEg6Rx699x9UDw/27bKdlHedmrTPgUUr1LwyfgqqxOaEVXgE+6FLNu
Kg2Ugq+fbhBXWFprTU8q0mktEiH5FreJZanSgYBHmkMS9vYqSTJ/bblS7VuGMv+vu0qXr4hxZTFi
L3QcvPM75WVyDE9tJCtK82NGzR6Tie1mHHlnxCmnScja+ykNwmg6DiCpwLM2nqMkzsKpo/taV+/c
2IRRiJ+UK2JTSlCoKXL0R3io9AymEnLcHr4RU30zh6nEyNxj+IO67MEfy+pZ1CgHwYLwVVafpstE
QyWrjGdv7uukGiCd1UtX1nNP49e3aPCRMvZasnsZneSn7khoVjQYekk9dCX+7aMlAKCvkmU0ASFN
Xh2yDbjpUxNtjbaWorhKKqTYTKnLe7VYDGxR2HCn568PkcVigUejgRgoZDk9+zhT/KPwuWLe+nC9
B//8tYgotJamOImq7X+8Ji+gL14ka2S9xTo3S6QEphB4JUDUAXs5RBKhxeOd+Nn/HL+IpVKuVEVM
BAoHQNvTViHGj0VCMBSBsosJXmy03sghbloOAEfpt5s9juMpTS8PTJ7coP8DgJ1evwi91J3QouqR
4r5bBC4DY3AbVgak9V4bR9EB+EuIzmcC24LKGSRbRy6bY6L3C+cHeeqzoNcztlTBmdJ36JVENBuv
ogLlIUO/fdL5mlah0x8SZzB+FVe/D0aaoEGRYZEgY7iegf1pE+SKwM+V5CNSu/Z3PBRgHnM9dQlt
tYrhuKG4H4KVe1mkMIj+Uw48b14D/je/o/eOZcKbiySZX8B3Eum3oyhWH+kKcKeMrITpFyok6oTc
SPguOT/h4Wt7XHrWbjpfQhskfql5+V33fFfYUFHGAKDcvBRPuMP9J4KMPK2OFUoswDtGv0oA4xXB
8JQlqmedEnyjUvRuhC6QLkjF/knHYW0ccSuuXnCfQjwMHVXKIXbir6k9EGb7bqh8pmou33b8ZKW0
VLxvYpwYs65DVJwbX64x6PGAcHic9rDIY1DiI3kwXb13IJwc0+Wb+Ab+u6HOGYutJXIqzmptGXqV
/fXf+plU19LGTBAtAqk9ml7DJm3849d/J2Pdx44JC6tqRXdcWQYXBa8fM24Inh+B6X1ITwSXc/dE
PsgGS0JntJO6faiydzu9EQqDlmakqEzNKYrZuIHyOPpcVKfFyvqc+MjTBBbVUJkllM9He9G7OH0z
SzSCNSOP/NBhCqryTLFYomSqvHDjpGuF3ZhiervviqODxtbdJDFx622KHMgH6C/RixLQ0Ta9LM8A
sGkUVU+mmPUZ1U4ob6sVwUvfIMBVHPjL2PGHucH8K3EBO7xNDYs1mSzYMYezbKy8BB6GrGrk+U8w
akb+HQFRs5h2GvKKqWqXWucopXWcIHQhFjr8doLT4xLC6eVyMccoM42GevXZPJ7sADzDMs11bz4R
Dnmn+uebEeA/dqiRDmEpoEIaRXPtwv1WHJSTrYZ7D3QtNeiKIcpIdl2CuMm8dtjFeTXJSnFAOIs3
kCk0zKPduJUzvR78q3WgL+pQHrR2HdaIpUrUkFTrEkXoYucxE1VoBNQtTQVgrm2D6cnQ8AvxmzXu
xobPdsS2P6wJ60iBXoFBWx8n9mwcYChu+WTpztNHG5HXgJEJ8HUP5RjDIe9XAhZ8eLxiu6CX3mFG
DaEKAWld662s6JLDf1tr6JYVvoyKfmE7PktuZCjGqa8GEXLBvgihOvZYkTSeX9SFOZckbZ6pRzpF
V6ClyxdfemecNGJJg2vc+TpxLGAZUKJw99LSePy59qRqhER/u7ginAiNy3L+H1In612OvODHDfUs
fmyuaNu3OwSZC8hFNFQfseTKXmknHo2Aq5862h77PFJdJbIakdtaGCNJxaIiCyUZZLnXgmCXyfIU
/sQlxullOzqbe6pU8utxIewYO2STT+lHg2Fk6fZWIKs1bQjIENMBzfHhVHoIDTllABz0NqawsabG
tUDtieFqZfA2STsFODlZSWLpRIY8nOrTu25sVcuxoAuFxIK5/bhyk/K7QttEP0ec1YstRfRP4+Ek
b6gbQTa6OCredOvgCdkRYAu8myB8jgcSBhGrqoFijVMwsbnqMldFRGxXbqJynyvxawHh0g0RPuqk
eXO14it8yaPp2DmqyPq7jzMd1KvBpiZK/sZ4nRbR/1gevfapv7OW75/SjhJOmRwSfs1oKdHqHcrc
5BIU2tszdVXELbTp1LZ+Uv9BRKyQjgk0MVSPu3thsPLTMCUpXX2bGoEsHWVuWDzcGVIHaI+7CF/H
p9aEY7W7XtuZVKcb/6pE8AOc//ae1zmjxxUsmj+Cg4TVCLNiyiX7004/r+NPHfaPcTSZsWZHKgyv
jrd+gEYRT2qzOajwH5/tmixN1GXCUutgwS5F6edF35zTtENmzDZTOzCkz9+FmxMQA15ZVIp8RIO0
Le7N3i0Az3GcEcLofvLhWgLSWimA0dV1K30GZG/sEX93WRqYG/amCaF0vZimVmjnY0e1nXC0ZQKu
JzNZLnMuqq2Qzn23vBu5Zd/0oI9osv1x3syYDBzxiNYweTJ2jPjjVp5bXVPhcz7QF3SdpL8+r1Hc
1WuUKtG4xzvvBvB7ffpPO5sslFa/U1vmdlPq3iy2i7ngR8i7l4SvKPEPIJhQ1a8j89CpOY6fq8kj
xU7fo0Aq6nSHYHGx8IW8mszT8lXLsEnH/ip6kVlpFxpsRUVK1htIUotxzztlFqrI06mmh5I3PpVe
qPSWAZJULTHuU+H8GzyOHiwDxQJTkt8FL7p3VU0/aCpd8rsCTQUyL1/wqVPnpeX47mgh4pW9IAsg
bmGPZ+9VBnZPGicSUH+grVakGNLWY2YSsoxo5s+mBIKs84Bam1TQLpq4EttmCM9fCZfFUQ59pQY3
sdu73fFjDY67o/6wWNMS2L6j5mkVxJ0B/P3zCbZZ8D2rGNu0itNCVe1VebK/WnFCWwEqkDEcXOKh
W7EvMKtJ0CeXF5IJqEmjHCsZ3qeqp/hKACQ0fZ1WOJlPCLjD/30Nk7MXOiPcK/on43YwrYoqJPsH
caR+/KtP1ejj4GPR/ecLz6NPUuXS33uvfGPlBTc1KYowNFC7XD4267qoisa5oVPIXYIH3QsFcdFs
BTZWpO34YE+a5yrPVfsF8XFKC6ZYBPgftyMQ0t/Cp/5cg5ADL6Dkrv7GjI7/rXMvoEfgD0XCPYS4
fdap3foHByAy4YJH/D4nCDA0G2ekftbuzNXA6vs3CZS68K/jkMFJQZGZm3N6v8GVatTBxZZjY4FE
moMV9wIMTB90LVDuVFY9KK5mRC8jytIQZvoA0x0KnylFBcGmXEwvoAdRNQx4LuWfoC1Xc9c+d2rn
sI6SL+oh1LLyCTZzmbMeew8EJJmKwO5SXOAkwgQm3Xx7qCjOuP8ERfAbu7eTlCFPhFk0QU+n6Qzj
MVeOTXip5mLIQJL97RnIQs4B+p8/agy0PVyprZfd6BDXA2C8VZKcjgfg99bNxUXO/xuGD910HxST
JcceRWH/cL7WAtzmRS3nPLeEjPs0BWhJt399ahr7mIouDRH5qRgR0cT2eDbgTMPVhgW7F5Q79sNQ
TYaH12dnCtQ9D7Od9vKCaJH6iw2motaWKBsuJYunY+EI6UqpC8pTHT5Jr/V6SExSKZcnoyRiWc4K
06qYezhOgj/nMfNRDT5o3z+ymKF51/GNoIJXJjE1qg0Tn9KpDsRwvMHNFpZmrPyKaikDxXJX+l4b
KD/ZFsV3YnJGpqCBeIyuTKyWFhBmCU5ukfTvrTNoQJPBB2GG9ytPk8wXb1mVp2LuUPF7lspLS/1d
5uViFWj0++1Fh1pbTDQxhr6k6BwNAiGYvNZdjBCuIIrTHDzqbClPg+4N61Fft9IADs4N0iamBV2H
y/pS0ZH5FTx6QkLHGm5ldWp/Fqn6fA0+H+TBLbkhy+MWRIjJstq3qigj/Q5QZ4zlIXicoDUMOKeJ
9n5TC6JZrkU25l6o6itduq15X9nL1I882NsSrEdcVfYeZIiInYNMU2nI3oqv/93mGkhEtGri6IjG
rYEB8iKsA09+BgHEFC5txGug33ZjYHqAIymzIiqwD47V+yOvbozwwRcDvcPfdbMyK3tMMPCdPphq
0A9mgIIRMnFf4HzJ+mIxLoj6pcMmOxdmyWJL94sz5LLD6SHMwsyr7mNrLq3hoYDaBBJzH9RCDwx2
UJFxF8Bl8ZHv0ceVg9X/PAXo58CnQy0PHe4zHJVCVVnoeFZEQ2o+E/wSOoa+Q1eug9j2ZtFdjQTr
btMy1wgiNzsnPROdgHHx0q7AClJYf2g2AJQnM7ejqJGS+SEpKCvmdpyrtC4kwPDYozhqos2/mBNj
mGiHxhcmSmGYO1+Rko9FDc441cQl4+drsjVKBe0SL1oqt0IPL/koGzPfZGFtX2z+Vc4IKTAGyw+U
syVYTnWSLhQgy4RgncQiUlPzC7ZIzO0zU+hzvaO5OP9CzsN+0wr0J5QrtvQwTYoz4+g2X9QDlKpR
axkUQTpN4+0yaW5dBNjIWMlaole/4EN1vuuiAxg11ILmkytIhinPgx7zrNWs0eE+IobaLDQa4W96
XcW2ISI9kDph7a0GNFUcZ8WNG3S1UsAjzJmMzS9KuWAvbtMUvAqzLt2quQ6PtGBqyKfNvZLkh7WH
yJeIgQoqQBPE2VQcIso91KWmNg0q2RXGxzbDGuRJ5HJAPI5kSnbD4qhkLS1PRsvXlXnXetdOaub9
6mQ7tfvKcRkyzE017MuITSsT3zDVU4POczbXHpjQxatS2tuikcSnQKJ64F3od0GMLrNYnzekAY6m
rlXbP3Zlp+c8pN7B51NP8tyaHHOKZGPJ+Ie4EZblQSxRiTM6EXZLC7CKRNRNPj8DLaYOMvI/5oTk
d0VV8aCFbPIgcMjcyhcfs5Vp4s0+GpsZE8iZMkXBkK4U2A0eRbNHHlqDwJWmjXfWVJovZ8X1xVYu
xJaNyMAnye1bIiKxlDIfPu+nxczb0ErygnmvPYYsLX6dneLUW79w3i91ZonDDn45chU8CcLid+5W
rNef7DcSATVhde5luNCbv+tFBSE+Dt+/2k6CcgvQLQlZ8qXxkJg5HRfIM9Os8LlK/8gRwyQDFqE1
cMstYype8IgAs/AteHynZ3yZXaxVQFZ4ehj5/eqrzexh6PdYCBS8RYX8/KtpPgO+WcRKaLHRX3X6
W5sNqLnu9sVWM/oxbYuk1EboLV3NAYo5d0DOFw/0vdYMv4ooj9Eq4HNFk4WiQP+u8IYJwobkCI3o
6weIK0aClZu/VojijIf+gHKGgMVfWq2x3DzK7yJCfKrHSe2cZMprZxGkgHPC5Pt6liv1ag8ZbaQA
842M5U5wZfqmXH7CAGkW/nUyk5cQWDDFOP5QS4eIV+nx7c6sL3YjcEuR2qDuGxzeyiCe6iIgjYZ7
VNCxBJBVC8kvkEvtCzRyJ3G7YlfQ8jK/6zEnRlxWUG9IlxmC6zh0h+gnrLdwnznaRxKogXtM4LGU
hLjdCtrUAkzu62LFb91V7LYbQgGsSX7znnDtruyp0NYdmHr5FJv+wQeY20CSF6QjOMLmHnxn7/uT
cyBMTibjqpnKJHj3XVWSQmQCBse9t1ecpbas+3EVmyFHVEaxyVXbM4E3Iwjh2hR4gx+Oea2M5H3m
v84YSdF1DUoznxi+3VeU0OkxtTrOwwHEZ8iM5uHI7A/KN1uOzzjeFG3KfUq2awkjVpkusPuz9alv
HUEuwfuGnxDIHS5xec2TS5FQATCmwzNTXPHB2lNdxqY4+EaHx6aUnvbCHXJyZ1frIKCyO+9cng5K
7AfGC9MP0ullwkqcawIspjv7sxrcITDrocr/nb5vi8E267jnjWDwHkeFJZfUR2wWH2vMZj0tKQQ6
gB7ph+LjKs5VV1ewemPtzAlDyfgqTbJprpDukU/xcg0b+pPAAqF9kLY3wKOe6DM7jDPng0MSPIXQ
V2vc91Cu2O7llzyZwwo8j8BbWyowfFxVwCjBR/9U1sKrD9h/3ntlN095ehTGhxyjSPZiyhGfR2DJ
VI3IlIGV/iPf6xUEr1OXYwL7Zw4cY3SC/V22cPOrXebVGPRZNjQdzYOcAdM8fYYWKklyswLTM+tv
WFA70oCCkufty9SQ43TmNuV9rKWNAEm8C6B018y7P+hrRp3k/JPAd0mt1SOPKDtjjJMYMSA2XHYh
RZBPmZ4I/F+0yOLNCSJcRtoiq32ISNmX9tKMty+27DAY67ZsStlqci42ZzrGbtA1DjlKZgl8Ws1R
SnCRJ3fYDddwcb3f28RzUAYkxr2IogaweS5+UNMcilSUmg5eMr+dICkAdua+xFf3p7MlMdAocSB0
qBuuQ6w0dLm8YxzczwXPz1tjMjQlL0vWJAQnfWPe6YAOdfXthmV8XBnmIDXby1xSG6mOa2Znw59n
YoQ3iJ7NHD8ZgOUre13q7jdU7QKvbSGDA4HM1vMu7nR4KczQXRjhWK8lOlW9ZnHm3Y2yW7C9G6I2
HeHTUbsRQ1vpKWKTw3C77QJKq7ADzIv5qF3UdQjnCyDE5KkZQxET6+GK7sfjruW6TjYV0WsDiChM
lN7GR1HW+VWJXBl1donn931uWunEIp47oYDESP2N27QBpWsOUZON3kKvHR79zqRJiCKNvgBm5C9p
0ixetDSYNMz8ORlMkcWYadv1vUyEpxWlSAb+1d6WUhCiSIZSoNRiVCMI4n+hNGBBVLC1wIFPiLPV
jCvg7uL8JjEtsRsfLYNKevH2icwEoXYPdYDm6pjS+cTNhe5sj49wGUe/8uyNSxEdDm/wryFG9hRl
muIascsTziqi4rqIRb+abccPsNStwRee182xgSKF83xn7QiuKyKCYkYgs6NI72xNjmPpqIVZZVXu
h+FFUqVFluqaIFx3zymhdY83g01VugHUqrnpYe5YKGQqblwcdxOrslEXpDxG0hrXHqWtBlyd6vkn
kJjsU9kgBfbEeK5tVmFm6bH2U3enxQthrmghJb9LOqO+LMn74SUQYGT4Xf53M42Hkmd70Dq//NsH
buO4X7bfoeMDIbOcTFtd5bhmYsCiGDw3iXZEepa9ku8x4MQ8XAU8eHVT+wCTF2ooNkMAWH0DQtt5
xvgaDNobMwxgcf0dQ//iB9B41HqlminipApybFQrOF0sU/G0uCV1GzlYxqjNLJcToqncAZP5KqUt
K9sF/EJ3UPgupyHE+a6Q2gubLYTu2LPnD/NSAdp6oqWNIh3h6wVYDZTxdiwA90Er5tTNfh4OurYJ
ev6kHeeZM4xIdor5KbhaLQJbeh0UAMZv9h2Nj0PVOgvJpQSbJwgdA+dVcbKU/r5UjpdXDHV+Ccdq
y3zL2DCwcox0RJYFkbrkiJwqz8rm+aZsscHQa4Oix4ThwChBbFHaLRLiZovMkbrrSYe2+P+cw/fK
7oxlLMMLQMMYrRGu3vljLLS24/e+x/ocyGf1hkro5PpXJkZEZOyIjfIdBznkh1YbJGUd9MaobKkh
dNRc4EK3+8uEn+ot9HO2pY3p/uELtk7xAQGsFiVXzPDnyeBObp4hJjn6jFLx7QWwxOT5KnPEqRFQ
+8bB9h8cROorcLfwXPY+n5B8RdrouIpogws08cxo7gHvzSn0rGe0S2YJP5o5YwIGEV7tfkd4ZFae
74OwREb/pbljhq4a+08leqg6wdk6MK8i1olICC8fkOnHCksnaYCwIZup835n6TqbEPLPip9lPX60
6jdOeJDGp9RJ+h6i2rbbQUcqC19HNjNqoAEAYejqoS7olPnYN4jTTrOV7hluQLmMzCXVJu6we9BJ
9kleDiPu6szVgsv+jQD5hwt+9FYHA1XHcsK6Gkb6Uf7WUUYpLwd8kFsH/dcC9CdV85rRpyfdAH9j
RXMM1zgOXrh8F2gHvxon1JlrXNDtRuptpVvDJ8PXE0p8JuliX37/A4mMZa0gjxhxdrhBd4htsAcJ
BADf5qZCRp3ok08MLU1+qVP3OvUZy5qVbdmyjs+e7hRUcijB8hS6AAmXqEIW17cCBBX0vzY72Z7N
XknUxu7F8hfzmVQis/qD7NU6NzD+OUsjXxf0PJvEw3xP1eVysLYTRWXIlLuR98AHYBPJQXL694+M
vHLa5v+isTDTAPfTNZ9xaWX0XXxbUjimnCxnbDFjZ+ImYowDR61oLqephsazFP12Pj7NJEkM3z6r
K/YL2aas+kghYKQNgsCqvpfRm+bjFl3hbyTklcQppq8mq+4uPWgSkApc2IYl9CfkSamwgZzeVgKK
xJbXudVSGNkjnuyRo4gg5ubfAv8svnJKLPk24bWQ0kT1PG63sfcPImmmrP4lrMx4C+TddlucNVpz
rtfSJATwsy42NJGMJQpk4epl5GRGrdITPguOHi4R+c0qqIqtNR6a403UjEYiuYJy7zLe2SzEUCWc
8XllrBNEOkhftTM0bUR3xQG82+Fm5Ewdi4kv0F4IIrvSOgtfbKfQ0HncdpGMPqPsmdwwWrE+aPYw
rSf7tJ1Xb49Z4zzJ6//4FxsKRdDA9zXuxqAF183ITWIsx0lXHDIA/bQZ3qzTDHiRr+MUmfj3ThIf
0f39AULBSzd3SE5DT3oOYxOf97jQvgpJO24nBIStXld84Pno5To11NkCUSfGHmdkw4GaXhjDG4dG
r14AFZFqyiP9arSylwYHtexfYr1B8wF3cHZvGgetbHvgnbep+a7kUDLRLiBDgxqCQYt0CqO/kdZM
ME2l8oL39fCSJlILJAVZ3bVqUfgedk/r18Hhd/OaSR5sUpA9DTpl1So4wHhbITyRWs5i1RLvII8O
vk1kaTEIfaDgOWydRKBBm9T02NeGNo/hLpVBjExjEEHHjy0gTNRn8XS/i6Z/JN4P0Tp30dCs7ivW
UkW/Fm0nbr1Otgl8acW2eLJWkM8QzGhpMBulX0z8VJmbE20ELLWxztOKKFmeHJg+qfAx7AUlCouH
sE4ZPjznLl/dozLKx8FHWcdKRuwO+mwuylOcD+16TRltgRfyg2M8+qUJ3kuBfBPkYodwiYWvOXnx
znYQ7bgc8k+qlAifgKAmZhrHjMAvd3m/0lxse7lfTWCdsg0UhFjCgbMgNWJ3TsMYSTx08AvEJ5BO
ZkCNrukb3hJjp0w/eccj8SIfNTamV9QdDKP4AOGl/4H7LqXSDTLFQ9gEsxJwaukmj3AzsqkyE5Tv
eFDCmwswBhwdtEl8zGU4uwzzjaWa0WBQyZQfNFz2RRYSlVFcEmMQKnLuVGftuwFzSi+m1nwwF/Xg
jkFf9OsTelCEm7eJutB7x4w/QYmRgDAcbA5rqsgn4XCZANWo02A4omVp+n/ccXZjY4ipp3JeCRVj
WW17ponTZ3JFu7hykcPbQpdDB1wi3jxqLxLmdw2nlo7psByhGyMTS1R59bYtOK3SpyPFFTzh5u/o
oF5A0daqhHaYbXUNKilUkRov1+KmRSHPBl9MyW4sq8iTzd1wzrOkvjOmCwIXBjgPGbaym8hW8Sc/
i2dgO4MFrdMxTIltqDFrX3takPZGR+teYtvCDRMU+ZrF77B7OTcaf6HQuyHRO+SopaID/vl2G0Tp
RQWvDp7q+R3oFuD2npxNOcBYcMppmMKQ0BEDbXPaEjIOiGFQGBn5gk80DuTYX/mripeqaeuxzA2B
tX32eqiCp/+wke8Eb2VGGnP6D/Tzw3bI6CpGhA7pQp90+dkfyU3Z/RbwhXyYgcBY0oomBIkFPpo9
dyj/EVww4aT+6Oa/6jtteGkaOSJczf2WKavZgSQGGirANfhIEoEbKwhvYzvHEZMGr8AujDbPfuQJ
0/hAXtpGeZvD2oNuSRXtFc15ppyBwCVbQSsL0Hlh1l2UEgo/+uxRV2ageQ3A0vZvUMbPqy0df5sm
HWk0gQun02TeSHKkN9Tr4N3qH8+C82CqsaZn5Ns3wlS4PKQPCXNL8qP62tvIhUzT0lG/V8Qgav88
kRUDy8r5HHk3XvpuO1JKnLZ7O6uSHDGfJ4fOBb72aBVpGrTlGuf+ZkDZKnxSd2C0qozvFDvFMy1Z
QpSnSv1xW1XbxC1i64liikU8Xdww9cAAIGhHIc4e7PglxjCTKcVVkgvLeLA2MT3CeO//ykGsEqPF
xILEeyVscT/0H1IL4bAYiw83NmloJyH8rQnvmOsfHn10/JqfbbeMSoCCEouWaLy0VH4PYML29YqA
vkTmpygsanQmTq6Zfy//Sjb/xuRqL1pSVapkOXSu/G84CYeeIFEOJaU9s9g1c+KByArtZNOn/6NG
i5UsDNpg24dSX+s/6d2/82/YMaan0Zm3GTQXUCqnZqNvaKEPvD6z7DvgeWZWOjrUeKt3Ud5XSTeS
VIULl7JmDZJtpjCSKvcSNZlghUE3WZ6J+pktOWYIeN/H/enBmqjVeppAoR3FkQnyRCd2jzjCliWr
zKWhTrgzXSxN5mFOnp2sccP7a6BCgrlw6JR8muIDeNjOshHv5uxr+UigZ5Z8c/i7CCog5DbhJ+lz
MvZecDwnZbXvm9EyEqNoQljVaB9W2+UabuBcZQ5pHlg7SCeKma1NmTQl60OkcsKSvmGFDyP0JUR0
hjzQgc9apXgJ+PonfEw2pWoZwvhmgnHtw/PSKDpqHgxXM1XE5M2EC7AZb1TpHETMTqB80bSKJrzG
kLd5NUsCHNskfO+nmRfSsRejPCim0VQh0YuMFNxBGxGtIRnia6i3UI0mJhlIKj5Ott9UGtAVrgLc
sG1gdzrtNcPDkVRWPPK6iOHn2pCk8iDoB4J5KC/R2l6NtEUlrLRTVRuTcDcm+SfS/a+jMk5bKLFY
pJTB9dLeVn0fwmyMAJgiKNZ1lwMWpWxAl6ES+ib0F+Nu4aCNZ12xUGnkUVLgA19NjWd0n2CT7oJi
DVAv9kQLn07opTyJe5FM1H90oiapjbiOfvs9esO5sMXq44sOO4S1jhdIhWO7uqENLJS1NFgnySVq
8Zn5iz764feNFbVuYaqebNPV/Aex5qNsnB36iOhBAbvhDHAQ3/BGqU/owtIExTPG8b9KeQeBeLkg
YvcBjlemwHip+qLIyI9+t+Z/zKWp405oEuOgQyNo3qzd8Oq+eSXuwchpUh1B7JUQna39xpdyrEa2
VilWqdqMYhMuCkKHbYvchH+CFtFPw3wg3ZOnN3p3AYILsEIXU+CdQGkZmV7CnmjZRcdeaHB7bKyv
y9nGBcwd/l7C0ubzoHNrpjnrqlXZB0bmUvRqLGas5TSmbR9RG1P3ztNbxsxQ8KP+xPn5g+QCTco6
X4EUR9GSOHZWG6iij+dLfYEGf92ZiTcUDNGOUe9a/MnE+gV0+MQsImZopVy6rs0bNY3RhhBWGvPX
iiFvpwtWJ7SGaQSf6kuODVxs9Ej9Mpri1W4T/5Pduzo2toGk9bcfYIfsi2O9mj3Kx2OcNHNLu2O+
qB4Yfbm2O2ZvFPJqpkX4FDO1eVMOUt8vnXcTTbYbRWMDY8aa64AwCJTseGtPcf4hlHgZcNjeBhea
rybqVRVigVIJSt7aD4Z79PdKXOOSUUf5WxQcTwGlDbeK+ctgmtomUJzzVNz5EvbX8e7Wlaj90l/o
TKFZ8keksGMY2RwKVgXqll1H4mixmz5TpCHlEjH5jkRcn/knznPIHnAjsz55ETpDnBl6njhh6JPL
WnVhtSuTkyrwIWZs3aBngvzFTr3vs9Alaz4SHBPoFF+jgx+1ImSu64LqfK5seM8QWD3MoU+OfSca
XeQHf4msen7WPpBPMztsQsCR8+6S5ymRyYllcRKeoTUMtrhyluh0tjTrPpvqgzj/kcqPtxQQH5nV
fbfqh5SjaO+7oEteeKDcCyA/rVnwipfcmYLXS4MGSkFH+FY5jX5Q77KBr7BQ7FrAvmarTXr+auZG
kvOLGcAB6M0OlDhIJBZO1EaQBoPjRIexeQrJxHJlJ7NHaGgN8PeckMyirAODuS+NSaF6i6tb4IBJ
RZq73KeHC3sT86JtjV3NDjqATvH+XGaVn9WhzVGnrDxCy2mK/5I7aCjVqPB4uvAooW46qQpIfZil
JAdBSECHEyhfbGMudzrZQV4ugYUpGwlY0V1JEUUqYfPmYsqmEDE3cqH7GhVldgTRtMyLVJpz67q9
EXfLMtM1WUO8m5zAYonh8sRvomnFVU4LhH8l1gsyazq/b+rMlhBCL3p9KhmoF3T8kc1TIToVuSWy
sq3kcKFG4lvwwlh4kfw2hYo4hCaWNBwDvIKAs/yq/NeE3KVr62FVwdpxnv0VV8fykDb3rlpL2sU6
UpoNFTHnH4kRK++XVPejSeI2M2Ry74dEZyHC4946FnDOsdB1wPg8KPOUZDEnZ2Zco2DDvtMwYO39
/+7ZxEEyM537KOrPX9pPqGiJZKU+lP/YVig4RFRAOPuSKrDq6ebEiHXr4P1kheaui/au/+ziqJg0
MGwlcjty2rmFbbeeJa92/7Bt0MF44Kwi3sTd4nwIG01Cxh7e8bNrlBliVXicJdd9L9Eug98/4ObT
CaTg4aSeh7n09GLQ5MVVlkSAukd1F3n/GJYyTkrDquUlw5/miCL31M3abgfHsFL1w2P0Q1Bvq6dE
wmAYR4pgLXVg8KlgC5oiuu/O8p7ESjYkSRTaN+8J3/zrUkvjTOr3pE5+EB/xlA69NRpEyiWHUJec
axyhmf+rC03i+V9FA2q6PJOSn03EzNIyvUWBDenNHhUoBz14NQcUu9jbgrsBmwUtDxxwllsnJWfs
73ShEKxZqEZuuFRAvGf3yuJs0CLXGRQtbJCxsRjkmK4wmlUM9dQmXLVMZwllPJnjqxfLGC0HFqpb
nMvzUo4r2EiL+a4KKnVCMITQwg8SSsal+z4tc4JcqZcdw65BliTduoIMFjWefvKNeA98HiFLICcp
EX5Xj08fx8NFDigt25+hYT+OqsI/8mZ5iA8xUw5JVR0SkrA+FmoWdVZhwmuPoK79EkW2meQMPk+R
jp7hj9putkYyTSD/eT4N5eg05KG6dTeRtbl0Szwv+l6YNJw78ZVEKIWQpfyzhfbWPjVrwrRANKeV
vO1JrUjRPYrdfGD0Hojdh029wAEszZjrlXlNUnSIELY1CoRA17S26wJqd22vQCOW9i78jDzOcWcT
0TyWOCxjaWc63GMkkql/iLlSkuwMJwCzsFqRjNMKBY/NZNmYYPm5YCeM2Lwb2UQUO5tRGi4XXkzx
cay2fqa3t4m2IsCVzbl83FV2SBt5cz7GvbX+3agrxDjgXLR58tZC8d7Po7fOdtYJahiscQZIO35f
s8e0D/12OFb+H+LmHAA+heNtWFT7Dkew0ovOn3xkhFW6IWHFESgWgCigXP80MBHPcxhOUx5ED08+
xD5JWzUOWWLGKWC6T0IR33vXtKPV5hW9g/vpmk/EaFBe9V9rMYsSCQfAfUnVnq44leEli4eH+Lhh
j9jUDnw2Kr/lP5i8Pgf5FMfkKUSOZD1Gmw760PQoMAkpl+YN1Fh0neNyf1FO32oIYOpD2XpHBpRL
DYbMbdn0iqpgeA5mPRBGsS/7AwKIe/xdsl+c+AVOHroaOdb9ydyENXqOA3hFGQBL68QrbX403x4n
zcLDsY3Ma8BdLJN0ZPkeKpy83zNFBa3yPDH7kXOusLpRP56SvShu58ZfW8SPlXdOZ4wFOSO9LHE2
YLbym31kGC8ClUP8IECSEn6DE8ja4eQJ61sufeBIKpUCi78X+bzs3v2Arlb9zLTOc93EdSHj5Kbj
vriT94EZlwyel/Pp34rNpZl8xR9yLb1+JzDdFq/TmIgUnUekuh05hxB9A9AQ5jDSG6ZuwKKQcpUn
d3SsoERQ06oGDk+7UDBmEprR0+qycznOsHEsHGgQgwYfIvcnHs6FI8ta7QIBBOeQLcB9Iuvi3iRm
kAzFVKXJPq+7JmkS8SPry39DPmOcRVMva8N+VR9sk9/yY+JLFfTmz5YAlN4rKk5xuuxuI2T4AMy7
r4JgjXNZJH5E+DRRtEUbNLz+Vbjxv+xjtiGPyavuyotcgxzFDafZuG59uNWo4rdvrVBsDxRiYiN+
e4KYfgKOgTxeykKgA74dKvDznOkJd6U0Rsr8G874a+AKoITxD8+tWjpx04rwL6dlalgSt2js3dZT
NnDlJg2Ey6K3WTVAB0XO9OPVf1vx1sgyAJqd/TC3cK99YS/XH6BQdT3GNjHtgAYnUq0JxOiSG+J4
5zskXkBFmR419IVQB9QnuKLPZr/a5MH7JMBElwcH9w5EH940UQKYdxrelqtgiFlXhP/cZwK8uL1M
nHMEDj4Vd55Hx0g7kQKvH/MLL82DeWQdHD5Pp91VR79giHG3qL3NUacVok/PcqaaTwY9v5lXVfGQ
U3uDD19SfYgr/XbfxxG9pc6nsYIqYMY7DKGkMqstamyr73QrdASe81qbeFQvT47dT/tGCvyyeaR6
HNI4DXy/GBpyzOyM8/gsGsoQbDS8nqT7qXWRY1/TQVrmU8mvC0wk2yvbAVSBHJlsVQ98T+nxLIUm
9MqPciU02xSa/7vqrQzrMY1k4fSADetsib8ljID1L/kSgaMLm5X7DQ3DYDkc/TWR+jgZdoF5PqOW
mLfd/lKzOzAESR7V/0ha3Awlk096xR5O7iMsdiKpcgsKBmxDLWt0iL9XTTd6cbcSs0X3z0uYhtI7
FlikCPwedemH8kWDG89UPM3rfhNMFjWmuWsHBnrALVEyXEEK4UnMN2My/GrsFgILapBDcVsdBI94
L+C1oEkQq6DsI701TmQggvn22EtRYB2ntGTPJTZgiGPFYpNOzkh8x268tcDLlsmo1lR7Y/DSHkOB
SKQgEpGtmL5wK9UWY9/RljkC/k5NHCBHJxJ4bsU2kekMlnCvNr8oZxsLM6FyvNHCmn+1PYj88nVW
9D2+3yHjyPK3tNfKpVMicfCTDP9UxyfsLitpcOSa1ntYvH8kVhEzuHrXlmKDrqKXYVj/pWMgQpB5
jSQpOH8yoJMhMT6iW+Dh96Rwny26vN9ckfp5IL+WLkvbFb8OpAB/eH3BwK0U1VAnhHolmkFs9u61
6DAuqPREldMDRBVdxLTXmN9OXaWSHubtWkFcZ5ZdI6U4ZrJ9He3kSn4mMEBHQl8KwPJ74w7r4aHe
hZm0jivAu9g8/cptVp42KTPQ69D/x06ih9Oo0no26iucCbK7SmI1T8L7c1EcQBcudsS9x0ikCjPD
YTLAg3x4kispuZgiATJYbuVpnTleDvJiqTlnDTfXIOr7UBie/vQNHQs1D1pQIENU+KyaR/TMMrs0
R+EjwYIqXh4iRXOa12UcIooQwnCoePc0vZUg6BFZ6zAjKBKehHoK1awMl34ScC7Q1UwrQMdRf92L
SPzYlJa3MsmlJGVu+Ac1ZmwyizTnnYTAM9Zrs4e0nRK46lhcLryL91nefrRDQbzwJHfnZvW/9rNP
N2Vnx+5qoFeDkv3YDs37UqbjO87Ipfl7xoFgmZDhmUDoO/TI5ExE7ArPfoP72gVcTb7DqdHylNI1
8dQPuhuCbfwk/VBEpgnJG+rqe0H5XIE0/ACyuon5Frtzk9BWH4480KgLDmIhjX18FLA6WDFhkU4V
Tx2Y/Eqg3WbdmyPSYDczQ8oSffaXFD1Q+/4eY5JSp+rzA8ryXzUBF/FkJEs+46m1/lZv2uuFxtcw
6A0KFa4XV4yycyKnvHj7xj9PkU6d56bEbRcQNJe3pJQjuULnLSm3q5wzQej8CyE6zhhRXKy0VAHi
+TheLAOFmAGDs2jRNYPgvNzhccErjQanO6BIvUuGa+3lZPQktO2BQfuFGpboFv3MfBMfxzzMtCTk
58lPRmGh3NwpCLi7yQvxDcG3EfPwo96cGWUBluOOPiLh2pc26EBrjiMNgY2DuTwnTymWwavfaheQ
yGqyU++jVVN3L1EGEi317j/wL69cP3rbcKDS/Vvs3CV2u6J00G5MvDM8MBf5487sb8eU3Og8VsPP
SwbFX5liLGL0EYJ0dKQKdETptkZ4CxEQ2nigMgBPACC/1sN7uFDiGlR5e2UbEMyedmArezBU0t/s
UC9nA6ZnFeUEla9CZozCoY24N6PzRsqXYIleQGfaWs7Xw919ab8Vrpzj2N9N/bWaV+Xsq8BKIU82
YtvzsD5pB0gRP3DnO6wd4ztFF6DRxJaHbgadikSgORt0EFIMAjYo/Ha/s9cYzpevVHOkb0wk3TMc
F6bNKDtF9MA3n5AU1q+RxgVxd4M6hQ6Ob7SDy4sJ3C7Eva7tP3JqLP629mr9+0c4fTcwWuAoBWRq
Wmt0Q9HJMxVYkaRdnsUj+j4GJjfZPR39pOz14rqrNLUl1os0sbO2kE/9bc16A/7/WWay1tif2dHX
Qk2/tdDm3ELfsQCkbCWSs1Nmjt5wWmCkajzd9a1vU5SuX8v4Y8yX3nko+qk4C5fFKX7/y7M6NJfM
K1S2SSWElmYnWfmYXvIP53j2ZvvDJfk6I6el+idqzeiDcWru+YO0OdgXLUrSY/u32vKTA27KJaco
kG1YztpxwjPXYfCZUxWlMUYHr8DDCvRUgL7MO2gKnxwvnZD0PuiTRzkX70lLR3Yn1kqTgBp5tXYS
YEaqMsB98tNMyhzA1oJDA7g7VascmPxwrdmY7B36W8VUR5TzJgo+/Xy/Mt+0BkDgVSwGSZb2yK7Z
cIdkfsQMbj/SN2+Fw+TosQFc1GIYC5b+ouQxBthYXDvn0bRt6ezHuZF4++kS8VKeYl4hCkYvhiET
FxucfUvYq5BI5sc/BY1Jv82HszW1+EEAnzPERkBEIUAQdoyPFcjfG8HDGfmtv9f8NxAOvVlYeoCt
Ir4kZser5+dZr0krgcPD+AqA+7ugVlkLY35ffKMyyk69ALVDwZFPy8m1hgQwJj8B2R/FdO3MDazy
gxDvQCpdtuyPhk2FtgX4HPQIUvAX7SFVts7JV74MibdNRSLIZ3gXNNmY5LwHN19ah7Alt3S17Fns
iS5eoXqUQMOKhD6uw/EpOiUpC+0of57vJjH++UMkVRuDfShDtbCFsuJojMZu1qvloMaL+byaRCom
iNEjYKrALqDcr+rHkqWtaLsEoKBleoGgwZOp4TjbTaVJu4zpLU1OR/GSzoK+6kLeR7Uf/nfRgWrx
GX1/SxLjPsy+vlaWFjjUchXWgSiNTZzv7meFqxSUeiDdWjRc7yMUN+h/lpWO05lKDdmGhATICoL9
LvZvY+FB8HBRocmTm1tQkMf3TzQ6HnHm+/ewlnUdkYycjsVcC5E5ry9h79UlqtWOu1CNDomQbaxt
rGUVoAPD7PncZX1Uo6fb5Zd2xgShjYzGkazQYMOJtkgbieBJrKPHCyAQPVCeYjWaGGe8YA17OAZN
CBuvvkn+r0Twn6aKjSebVuOkf4xzroNedxhKBPHHaHaxhONfPmejrAi0f2N2Hyu+Ddqk6pnbOkLR
IkjUB2y+tiwTmWe1XM1Ja95UtdMWhLd8wpvk63Ih7mCNt0sANyjdzE7YGz4zZAqXMq5Z4a8/Sf9X
klDqme9Rh2LXA0lQaAW+qEo+zyS0quxIGTPXyxQaZZJvriE7NPsHcbT++ewixzob8fQednMSJL0f
kfKIYG4RaLQ1xCFn0x1ZDESAUMT1bNG7LH+4zaaOZ2jjCR4rjzoiynUmdz+0m8EF2ddzKZETj8Mu
KQGTZAf4vLWwUzI/6CEeEC5SKwW9kPsf8q4aiG64Mv3wFnn01dCUq7wat1HxB+9ZXldFoZn4TqQU
isORjsENJJHPBpfJ9/FiL4QdjMmwn4rGymuc/DdIfABBJAys0bfUNNJ3zJodGmYvu6sxuDIqMSJf
Oc9CYIIs6Wwjqff6qIOIlbQRKKmpLNWRQd4O9V+9FzXsk9WPLZOE/uhn/+gOQuIWhe5faETSHj6E
tmq2PvxdnHNtdtYgc077OoQLeHLmWxL/p1g28mW0Srja1/RQu5KoIzs9Gwyy+l3frzOtGGjot8AL
EIvrC9GAGdJDWTt8SVreOkqLulQVSq8T4Tk14n3I4z7yT/vh+Gp4eMPggdruRoAaOP4KpAYaWQ6b
6+Bzq0I6gfWfQYFVqviN1iu8KSeQDdmh28eVhQZNcjF6AlHGVKffb7zGrGx1ms4ytzVI1xvkmkwF
k6hU5SMAGFGRfKifCc/rWaa0YZYGr8wDx2FiTo04sVAPLll2VHJvvjPfhegt0xR6bVBZ8iF1Zp3t
HF+7dF1UKDhp4dWFtSq8jTqBHgWcdXk53ni62eo5qasaORB++Pdd1l3UIUOA4hZWQyPfsoNHjHOA
3bycKl2SqvH1EkwzWA+bmBOcPU4ekO9Xm5xwCaawr1wjhw+I8exZGt6zTqAG9qPNdh42u90eAVCZ
Df/8WOBtjhf7s1JrG/8vY1Ha3eec1wXTyieb6upXiSspf4bSTq5PvWAKmxWzP9BBbEOZbnsAHmgs
wulpMhAdjmpKF/DLPIMl1Nk8BoO5LWnwjaTrEaRggCP1zq88VsMga0aQ9ah01bpqDFeVz7B65heZ
JGzgI1ab/6UdGA4nYF/6HDKZLvWu5r2wuHTJAr5erUPK4u3kukOFzMwnW8vbCiP3jpchpZiAbdi8
Q3iZ2FuJEh58ZIrAWKIo7O4sT1wL61zWqOqdL7U535xvDbjya/KoJuAnkHtKZKYbip4iDV5pVS72
HbJEjKmiRXTyRJTTzfQ6txaQtqRpsSbZwFPsbTlgp1CxazCJYOh0mMr2XcwsqpULWzi7BxK1Agt+
F34WBT+8a1B9FtRYhvRYrPNMMFfCBwJDX6XSZBXmMu1dSm9JJZ0p8xkt4PI6sMSiArpJKhGD5v1Z
evpKENQkH8tVyh1qqBdamdUjitFoW7rFyX+jYYkcD4HML7YYEAedxiFIua0wD4Db/BuvJH7OxilH
+VEJQkU1HGAQRcWyUF3pGnKCA3SbbfJ8iRSX4GllTKLdtHXK2jAY3p/InsgT/19FOr6q41Rzu1Fm
7MEKCCvUeO3n85HQBgWVpY4t2nn8rZI7JZNWrpsOUxTM0sKfz+GwMmvTyTnpUwiavuAH4J7VA8MS
1UkZTrmtv3K2OwxN29bAXMlVuRphsnUkq9KrKeYgANqUuYgCb+qvwNgoo5ALe+yRshghX1T5oX6Q
SOyDZbWR0s5SjzP9OIlcOV7+I3tlGNmD5Kg9NN360St+sl0xc/gtADmRvjUB6U4XAo7EO0upf4Dk
gU3qqnEIipe2cNsZx9VRrVeLslmU/gKKV6z1y808rU9FoAdDiysysv0r6aWmA0DXWm6IutosLVy4
dwYohAv7vVdzZokhKDe9vsgyKW24jxU7/Tqee3QWvBHr42LY6FVRX9nOHJtO6IVa/G8xoESqISyd
PLLXnoy0gXUoF3hfojiPaKR+UKRHA1WLsRlVkLi/h2CrO1KQMOd+3UfPu+6Q58dF09p6hZFd6+iM
j2gETrRl4BN3X70XgDlum/zf8cNf9q2AiOmax5VRbFHuQB7VN64pETMohiqvihbcOkI5fjPpPZzz
O1b11vEQfi6cnsD+i5lLjGb17cVDkQP94LAsoT/imy2bjz3lF3hjDplNWuQlwMPTtN/zdDldugVZ
C9oCgq3QXJZII0o4aCVx4yM4l4pazvADMhV1R0tcAufOCvYXJ73w1yHouJ6QSso8CxzJ4ZuK8Lxu
ZetZ7pyJPU6E9u5gzhpSsr5zSkpU8YnzjHbwdidvBQZMEk1/ct+6n0v6Vb6ZGYRGWiKWnP69ui/t
bhEW1ipOPY5KIh6KsgeF1lOJR75yfXEOIvB3sLvxssj9YLnA3nN+a8zmyMCl7ZhzW2BSNuiACFBC
8eL9AjH4r3PRsfnt7InMUE2IZlTgTZu1/Upg/m+F7pJ/BykgPjbUwS8Eh7G+FcziClQe5fHKCiVQ
sl1oZaeB2WyEE57gjQfQ6W3NyNj+IC0ayorxQHcCHQlnfvgqOuMWrsRLr9WG8k0VGla3WqL2VlSo
BmxUflXYEpTVBEIz0AEkb2IGn3Q1TUnyem0bWv6l9tRvT4RrWAdCsRwoaovgenJwvVcEippVSqji
Lcy55qwP8qX39oM+4oleHJjXQx08XMOo2wNfNf6t2Ur9c9RiisEMfBPaE5PwKgqTZiLTJLhzMtn4
BDvOReFX1hocPJ6QwXTc38CWtPxCksB0UvURYMqJ6Ll+5Pt1fIENdEiYnm4Db/8xyWcAwhaNEgMQ
h+rOYke2mONEWX/Pxb+GWOIIdqO/jNcvKSB0eNyJvO48o7dFojLOjzeaHPLtY017l6vjaLrECCLb
OR7kKIYFwf+S2YSpJy5AVZ7oW14vRHR/8YCmiCHrLpufe/+W5LGiDx51RhYBnzlqB/XVMuzz2ofL
qShZjUF6Oj6j1soIpOfEZSwmHeQYWw0SHvrEaiF2Gr7FKxyvpn71SM+j09Ew0qtjxJuJiU6STfb9
NrNAP5CTjFPRjAiS3WkwFer3uX1Mk+TZfLYuxTHXVe1UeMJ7sGjeNji+1rAdmqMiZZR3BUO/Fv3r
+cm8HzxyiyGBc9D6PzfJcm0LdpOdVumXrcEVkuHTAP1QattUukZCP1LJsAzSsWhny8JOtdbB7Uv8
1rTuFGrKl38xWoNKkWHiXdhUP33NC4qswq4IjWROyyTphYPTd0WSsZ5tHd5ifP5O/LAVB1zQmJMD
wBKSvGEruPgX4jsSh3PyXQgQBC4XOx7mvOC0tYIB/aCD9D75IkQtpNxPrAh4T8mFm7qYjM+2wQ7t
7C6UU/L5ziIp3NR5CngjvKMbSm0AgYEXzuHUvdg8VD8zNo7voH6kOJAqr0OU7MwUG69NtUXGPbZQ
q+6Q+v0UqMQpHUJL7kHponSYF9WxssdfiM0X+YP3W+i9idqKLD/uByUiHMQIJpIu1OIAftA/Jw7f
1rIeRifnziTV5aH6isA+zDyOUzMFScOovCiLMYlM3zpHVfRBZqj1uWZM4IPLQbST6Et3iWPq9un9
yvYU99PRxKoOmUNEQo+7DUeN9kNbxo3YAp8hdZcM1Crr4SMbiuhA0H5ZJgEqMSHeDEktmDGJxxkw
PrFUiAa3ofUkJtNskk5DFFIcbGJ1pBvR7PKqg4Ix2kFBWRwnSaT12awsPZswv2TuTHkFdS27S6EV
HOzzsTV+D+JmCK2s53dbpGsbGvuuaQhOJKybQ/kBZ8FE7U/nw1E5ZTooPx/EMFPMC9rEyd/XKXht
U2KlXkJXNNn+WFCXhSg69xWQkyI3MgyaDg/QCII/vupDIk9JjBjkZqZN9s/+Be1TMctda3ghS27/
TcrtcsH5UK3JjQhidbBggeBxuPcNlrxzN/0YAWtEVstshsr7eqhgFnLB9TFUFpxmEbItTmZdWLT9
pGo7V/uzNHPq1NkmVb+jO5j5okH3ard+KztE1JK3ZKCLJcG8u1QGnD/jsJM5n+TwkVks5J6WJK98
XY3V+RGf+es0qDehDamJpFUESTQOUqtCP7QRUVgYcoROigUCgEpQ+7LOGh2XJFo+EuBSWhFcKJsX
zs7vG61LMnPOpNfySxv6FrAM416SvZ0TyEEt/0pWqq+NA7MI9IUMSAwETo+bJ/GUTdnBvum8X6nU
8gCmSqdeVVJl8zWLqiNlc0WrE9EnesBlN8ohUOAOLX9WLe7s6Htq5aAqRic9fwbhaxfw3fZsBew5
aIdYYK4cfdbXHZzdb9V8GLLpsxyXf3vvsblEbb35oGMqh2yQXOI+6mNNqMoyqBgg6/6JXTCy1z6v
51m8olCkGgD+Jg+0POX00/gaJmev2lZtGRRvWn903SW6FXdDU8j1Z/EYHFReNZ/JEY+eSHdwl8Lt
lbwJUt3rdC8bKOHKEQmpgKsqzwxwy2WMnG9hlSKqcUCC9g4wJZaGsfz7I2P5pHjsVz5yBmZBHeba
z+tiGk2vcngGG0ybpsWrORyDXFI9c1FiHOQqmhzKVi79SyHO8DVafv8zIJJYqPfBTnnlIHQTOQN4
M9ud+gYcHXDOQnUkIX5Z/DWiVSmQkAKDohV1XQcC9mFP7rK/xJieWWZbQ234LEOTvCtmuoKQGREY
5chW67w5Hul7DgVWjWSw75OZWL3yOFQjXYNFM0swarPZqCaRxEBrYHn6wBmptW4dll/dhko98C/D
3Gky80KJs1EcA4j3iU1mVRONFTCMLIJ5iqRBSdkHHYHWg+SJPqPMReZZEcq3oEk486y0dHC2jaHS
3I+pzvNgzzaG0LbDNXwyv5dw5ESD4Ky5gBoQWtqWtIwcPYiizjbuOOPREMvdyL34ZGs4jb4zmcvC
VGtCucMdU7OJezq6vh2FIpyVP92YSoBISY2RZMxT2Eo4IRqHnfEcceN3WuHkIJW70A3HqAFUyEMy
2y9sx1Zmzms7xJ8iE0GCnC+JAVn08pchmVrfZuN5Apu2ZfQuDFy8A98m1h4nuFAQfAyddTpc3ejb
pphfOaiDOcpJ+lxBKJXzKGxBGOT4t14gGiKA14vNJxdvGLA15UHje2gRtKm2MJLD3683RKDwWIK3
MkHcfV4ppiPkWp4+Ky23Ox6vu0r7DYILvqA+HYP+AYqvP7RctEHYHgR80Ji5jG7lBvtBaWFNeADJ
kG47x/7CtgGEd5HfHNsipifbTWlqkjXZ1tWitrn/7YPObXXLGkNryyYPkyb8sbtLWG7Q56vk7Qnq
n3gIKF4TUSUTmub0K3MHFys6fwaSvacPe40LNXMrKrgYt66is+ZfWzy1KHGK+LP8j7eE0tqk1LAJ
/W1qxkptRL9an4QBYKEqHS08L1ab5/0Gp5PNaHbvvn2J8Z6Vb5o7XazLIj1mqJVlSlawJz4ljVjQ
uAUsOAAfk7f/N/+ag15vPw0cOSjCmqVq7WwH7Wbe32Eymn9iHtFqFISQa10bGpPrJJwJsprOUVBv
X2qg8TXg75avN/PYxSw9KWu6OZ1pDyCKzn7ncDxRik71svmRO9FO2piH9DlSrSybRBM2YQ1Twn8p
4nykMFVmIuMINp+N4kJazI6eY9W6H8/g27TnA/LV7J+yZWpMMCwZ00Ng9Jy6zv4cadnzYPmWsIYH
a465jTxNm6g8T41W4HVWHkRw0O2CSzUoBpaOjr1KefF4ijM0CVU9ybeNXKGz3kOnp/Yq9AsUOqao
XoAakGEBnqDDAjUoxKoQ4Gr2s2XIFbGv09ZIxaAN0v3JlO9kNWJRgb7HWl0pcWEcwv4PTp9nXsUo
2IUwwDhBooO+GgxlWQiQMjicf6KO2nywljx21hUwNMvY1RSqXMhO6W3sLxvZcZq6oP1QP/Vuveb7
o6RIWYYmP0490bXdM1RrBRBCMF4/7f4WWnNPjarmLgYWCQDUlHVPVuIvfzrKyPr06jlHKui6o0I5
oVZsSSOLm4TlUKJHkQnvJ7L+LD8FM6cmyLpxjbS92bOrmQ6QqMCU9pKLAR/IxOV+LTHgBfihBp4Q
7zrguLMcGiQl2yVC5wh3khly9b72OZUenQGz/JMdOqrpKUXi16mrECUvSgNdBDBr2afrTsinZg9X
L8qIbS1wuhw5uecKK9HVpRSsKmfqUoaMO2UOrdB0TVAEvEt4U055pJ6ojjPn+Y9LN9ZoC0I2GSWn
EtD1AoQs8Lk2jp4DBitqYRTclFCaSJ1lcICiTzjbQgRZ7IWWhZZ7LXm4cvQthiq1tmWylKl8Ke0Q
qzEYNI48iJp6AzGBYrTFdB5Jh1ccwsA7sWMIOSb4WumiNQrEEYrDkqH4Tyt5ov86wa0i5Na2+E2o
MmhAtoB/v3juC7uGBC2Cr6sHCpVQn8HLHid5CS8CBrk+q82sHfNvBQlKXTnlhcV2OqvLh6fq2w58
8krMl7UyhoS69cgSnfCG6t4Su8Irx1LCRlM5HKKn2vfrFq7h3XvmrpGw7bJGcsePV/7tsSSoHY8l
nKpBY4AyioJYOycwONA1JpVA0VQFzE6ZrajpheGfuf/SUXcyWky9ocS7+vQmz4pZZLyQ98DfjwRS
5mkJKMSdVm8jV2PyRe/EbVafiuLwy/F+MffADoUa6oThFxScwUm5Q5J5SQbwkY09gb2Bgl7Ryni/
mXmOrtH03WVG6Gx8eIj4GyclBNvOs/ba6Ee4i1lCb0Pe1cYXuV3Dw4xcd0/qO9LNc9OMXk9ozSIE
XBwDmhrSMAOXy5If6LZQh48oOrY9N1bRPRTxrlZq9n2YLGa9XOicXnzRSOnQv4aq956YzzE7XkHV
QrBm6oaflmM1+1OMD7a+rZ5i0RonKf2bWdH9jjO6TArNKfJ9hggQYIB1DfwZ2GnkUH4Du4a/Yi4C
VRwy/UPMywM8lRGWclNXWfEvFxVYWad2onLTFShzuQG64N9EerKBNAOLehpfNgSoiULCp/wEIsa5
ris8u5IBStNP/pGqxH0g16grcIgjD0PrqKvcuGJmnLvjWMp9athJwTgw/quTbBFzdXY4Xs1XIM/m
Qqo74ZXA+C0RFxN9tVlJ3z1qY5eSqDUcOz+fdMOxG/IFaSObJ7KDkQ+I5YmyL0Sd/BjMtj9FabGo
7pTbEm3JOF/itpTF6TSqcZuzrBD2enr5KPH15rJ64FYf1WnhVJMInfEzLBIXmLRu5q9n7aWFF9Uf
q831eutH2k1B+MxDSmewvIGPkmSeNXTxRbOmVgQSZtYeq4fGCh8VMskR/pELgxRHisLCOw41hjEW
OnoeGwPZwTbvHHRKimBXrgN3u7kmzDBZHcyaAegpzRzZPmM/Spk6fsWPl2vQuhziYPGIzYPobQD0
Rfnze936HM2L3Wt+HMvU/C1GhdEiAm5A9LJGpXl/04qCteTpFjK4H1Q4bQvVsxYctKiMRTZwQsGH
yTnHY4Zq3Shva+V9evn9Pl6ENedtDv9tYkBd/rnAmfHY2j09AkI03W9LjtyplmhUSun7KwCdNeIe
AuLdd9w5Z7AYHVxzos/kvilJ6kN6eqWTKBL2Caz3RS0T3Wdbw3C0fw4I3uBHMJDIR1zs0uPy06Nh
u7TZr5JNuEXLbkl4yb8pc3mAQF0ZC8JKw3LSjZnTUE25eHDsQeQvRK2EUMTrJI4tAqoZs5RmtdqQ
aBuem3u2kWNm8Muszr1greIlNC3muJfnzG0gw+vhGxlSOsJ8RDr8fglUNcbtaWxHWOYIbILWN3FN
xff9B3ODoCwKg5ba05ckLFIpmA1UMg0qaFTpZGWRHDfXH6ABfSKRbVR7yX+tN2oRMOxneaMApF9E
algFBGJNed6YP4HumHgv02g3DUIVddql2vtFLL5ksD3zLLeyzcRNm5EmyIZjlNY/bKb1+nq/BaqO
V8qzVi3lDmBsEBXOip9UlmmIftp9N078KDZcGh4y9XbPpeWvwJneiBUJ+Fffyzb93mEZH5Rv4/F1
WJpX4U/kmzqzYLQ+hmXxf0q7bwf4SnqQ2spTAlpLm6CzA+gGEtO+Y87LcJp2AK/k8EDo7c5g8m1S
5ScqtzW9zNLkF+4PS7clTshmssQC1UjvQWg/nQ59EAt0JnK4Ce0lu/eif5QpAhWOXAuYoB53UUgY
AuLmzlDSkzJmYIt1JLBt4XKsQy41P2X4YGLp0rLJqfQqvLjoHMI28LSu6O5T1Ntuw1z6zNmBNf2p
LDtYAc61oDVBbAluwfrHuosFEDUEz/iJVMBIuzoahuNJYnvh+u93Vv9ij6/WFsovoE+AdszxuQqu
g87sWTMBX2rwQdYDk432s2ZQl1jWiq0KzgkOZOFUjKy7ugHUIUKvm6TrzmVOMg9Sao2IhBZKKQFa
fOfyWBrhzeOai/hgzIuhbqAJPJxzSJaET7dhoMGX4TmIWghz3tNo+jId+2O7EK4OJw56+SFSmTiK
A+bvTL50w57cQYGw7DKtwWqNWJ38dmKuANHawSdR1EBygz1eVDQ1nrH2YFok8JQkAviPFOubws5K
ViuwlBWzy5TbU5lStDFRcikeppHOWSgQNwuFt1icyKgW55HIc4BN8V6y0ykF6YQE+td1cVlXt+vq
MuNKbeA8GjGKYgQywnTvyLLatv5zUEyAXxFj1Va6gy5xjHK6cdC+vPoqOibFGl/a4VwrZwc1/Yec
CPJlmedZYJjFF1IxwJqITauesNtY43dmyCaDFer51QFskJNo0ErwZLkwEGdgBLHI4/acwBmWr4sw
aQjqO9PWuH79rX2KXrDSfHMB3rZyEANe+rYl0vai22c3jBTiPE1JfrTmcbVFXm7awZBCuCCgUipv
AE9wQBSk9Rw0lhxlhXHzsOCiMhGg70PIy0ll1WcWNV+fiRK65tGoWQ3sSRezI+RlxQ15WG1jpPYy
Y2y2cHuUhCqrCwS38Uh0eMHQdNSqxQVhUSFUDDhWq63+WMnWhswyRc8IqnaaINQwfiWENRpIVsVY
w35zNL732zxxi9cmH793MxRKMQMWRtF2ON/9QRLG+jdCuZhvWuhbdwW1F2XzlH2rNahwY9Etu89Y
aGLzR7JCGWG0PveK1HPuJASqktKtT7SfBNro6M63d4A1gK1/+tTMHW55/th6fcuPDZjGSRdmGg/H
EicT6uCz8F3Kxlo425NrHlCECY7A2aETfS7mBjb/KJA4LcuyYr5fkbKDsw5qB6/OP3od/LZ4JoE1
koPUKgJxAa4kTeWkcS305tRMc7FKsrHe5XFoKtq6/gWIBxoZ4v/lmNZjgY32UsH6/6b+zPC6Qzfy
UoXPGcqYqMDwxJ0R776GUqVPD6K9Z2JLE9wUsF9zF5UvYS9nZHMoIXopElNnftp1JCswbGQoXQkz
yIQVeMHRXL78nTyJtsSinNF2kOxcHTz78N2EVQqC1veaUslp4Ocsw/Dh2F96UUtxyr8zqEzmAVfd
mE/4fnYOnYSgtP5tlsKMZ3uHNymXhnLUzz1ql4M+7Pr1z9RlNjSlBFon5BbU1OAikTcyTZsHt8+4
Xkz6HG7aUKMQEAbO1z5HZ4STCIeTxSdH8Q6rsZ7wBAp4cfHg2DD2cUIYk2e3zmzTrKuZCzssQXha
qZSu7XtSeuGhp0WDLxmEhfyjionccDjES3Cl0bVJErUidXTts/YgzO0fvH0tcFCQ4YWSO5tLCfyU
NofvqVxIBfUA7JVJT2w16RSR0FNLUvQqRMbdt4fjKEY9tDKFDHoiF5006h6y5KZxpgVzQ7JRvvEo
YVFrcBNRb2YkSULkBDa0EzCQd+VxzlIDGLdSRpDvi1FK4DT3Bn+qr0wOiNsrsofuskBeLC2yVRTj
/l0SDANYCxNUd4Rol6Y8A/1tn3oVo7KaGyHh0l0iLeFq//7zidfS9i4TtHBsG5LulHvUqt4AL4Ec
54ioNnJ/MMglkkFM7MoGn9BCj5ShcfBt4RAafOCM1xc4iEGdRXEqcp8rkQnDTf1Aks+rVUnyyAr7
Z9EFb3aFkEmH5sUcSg2iiqNt8wjgNLg/Z6CtXS5aDVVL41ciWEOTAj4jB36bf4eYrosWKeDXiftn
zLAglmuDRzCVjoo2FTaE0eHmck93zSB74h9Yvrz60EzHKrAuP8uywoZVCKasjxa6VmjJKeNbrOEV
pL9y8HBCH1Iwydo67Hd6DvyKMlIIG+q95hsgfvEBcooO3D0fawZuNFAPcXWuyCdB4LVMW6mPAxQk
Qdv95+pZgWm/Y60wjZiAUH9aOaRTdcsUOsIp+cv7MECDGnQBcJxFcxJuicO18DAjvjoSPGVRVTh2
h3+ST3Y5BUFTz5NfoM1J2b4+ep0E/jCc0ogeOrApPwJjFRZ1wViNLbXyNastqPoiH2FO+PRJfu1H
Z6pEF0olA1e8kwhXMYjosIeR/Q3gkTUZsAfzgt/i5qG7HcV/u/FUKE3PrbfgfaOgMGY0YcyhGRdJ
Cd+9xEN6LUgzKgTLDg/ti++Je0Gkslpr3jK4S2CaVoKO5MlQe4pabIqkYgSmT+8a3UfIBpEk1z3b
esullubdIV30LvHxo8X35zOf/XBmwTTJIFd3XiKfpbd5yAb1SfN1dfdLBDoA9fnHyhw8DgSMDVC8
9by1JEVt7YGCRNtf27jC4/kLmGaXYzb9HF2s9vwk4vuohix3HNbNNU1iTP9WmW7SHGJekr9ZECee
abZ+YiQZ1eYy/NpbB2ADcB2O9okFGOC6cXcCfbZxgmH2BEjqBmOe3+IMLzQUKrM3oliQ3Y9gIDDO
XFHjdvNsIxlhWXg8GdO0xlambGAxb25rS076GkOMYgY4XjMfUoslWn6aRiyZBwaKvs5iF7k/r13D
dCFQI/6hg0LTEIRXTZavFE8gV3Nwa866b8/caWhtWS/lFE/KoK7M6ckVDKdQjtlg2KxWzGWUHRMP
cpOVCMiUpUXTkKwMmTMTva/O0K2j0jjCNRuryjyWkj/TUZuHTcuFpZwiYgJaKg11Bzl4Cg7q9eqp
Lf4bgwiki9og47XDUDYHunTtOnjeWj6OvljcWeT3QjAcXPiTl8dE4Ku0pYqZvRHp2CL3IPWWAM7v
vaCVAtTp6xsZFKntpha0P6FFBjbrBfXEzjnSTiFhsJu5JqEv27z1GIwzwWehFFjd68nVNnHzfjVS
llY5yHHOwMaTu8eWZOvMXhz9dTPca0Hh3mtJDcNzV5hVPlrcaOfaFsR/NiQkaZ/IFF69a3RMpNv3
B1YLFs/wf4Q2GzrT7vIWjD5FoO7ki22X5339zm7/9Xq3SgarZM8CicZIxON0nE0kv9jBM5WzatBd
SMeqhVaU8vGVrPDlMSI3LCCH2MN8f4Y0cG8DK6Qa3eI98i21yxqcPn/v07XxWDDaZaxpyewJ6PH1
jBsiTTzhbgvCypmUkQHKdzpTvhtNnhymWtSs29NDlMavWGh2FhcLXQ1c5hW2CaEj34/nfPEEfpjQ
ggLasB+MGVOfzxoWnSjQuN8v4lUNc/S8qN2dvf65Vnz4S/0XVoCuGgopnYkxm+aVoCTY/+r2vtRI
Ou/GlNUJPR5zWyWA6y3GnJ3su9pu/NF2RsbeT/aTrz6qXXC2rP31gQj+1FHL4ehCzY8JfhfZUkjt
R8qWNathdAR7cXU/FVt6f7+FWzpoytRSO4glKOpkocqaspUt3ufkW5U4IjLQN9RAkhAEEeUj6PD7
EmoPStiwFR/TTyl13okSZnnGjbU2jXKk+brbMES8NZws0fgQoJtQLYgGJsKiLKxNU2uOVMlsJPOU
0I7t4ssijaOk+UI9oIiZ71SIqglSziNmyp6s2k6NXWx43vF2e5Q6RBqB9KNkaFarODTAb4iDs4cm
H+qPlC2YDpKDYrao/rld9rv8ZAMhDVs0cG+AlY7P5kmqptffdBLEbq0rT9MF8Ax619KGxDKEx82W
z2qCujL3zElVml9vTVlM3UwgQbYVujm/abIZNG+HN1PMF9PE3J0Toex7f3ml81wTp4IzF5qA/HOe
O9VSZzx8sQ7DNlxdwbU+DYWyMqt59U0U1pxQBdNvqjd2IM0KAA8fAxYBNWc3/9o6hF7d+2gypkEI
AuWZfbmSc2EunQB9QCvXwTa7CY5X3+IAsJt4p6CfCgNtrfzRCyqiYU1KAGV2h1y0qAch1B+yUpCN
Fao3i4riigFIcMtpOEhlfxLeIQm4aOtdSKQNkAd33eplMz3QZAzadmHK7GbmBusKPJyrAZbSdw/Q
TanlfM2tK+K0B8BWtnZbVM0bmn6HDBKh0UEJFQUyL3oQAxKpqI945cQWlQCmJ+WQK031WzQq/aaY
GYulgKYPyh9YdXdlIxXFNk3Wh4fyRPqFJFe5TUuylSBq3q8NJ9w6AkjcVDqDQ4rk8+TBpnXlH247
Mpbf00H5D22m0o+wcw7xxO2XN5jWACkJXwiK40g3oEYLKLcA+tZqqd6wFNiwO1Is0qCXhz3YhG4g
1Qk/vOPiR++3X55o2kczsPEOQqwVKuoS9dQjjOVysBxx1KBkhVIoiuuP6td83yLmzOLYYCA1RRaE
/YcXW7YRK3rF8ZuN8JmPh60eC9Ga2V+8b2LXSo7ZegF2MXvu1kF9VQ84ONQ4JH+zqfCg42H0PqMp
XoUEr8z09ZTd5SzzHI5Da/cgCXWxFul4rYm0SMabfB9NMI8xINAtYBIP1HxXhYo3j4YlQxwSy8Kl
cmARIL66vIRcaAclJQAavoCpXxmY4r99uN9SoBCIeQSWty+J9ncJRZwM+6JN/fKY+YFN/1vl6qi9
FaEpnrBS23NdEznYJngQ4lBqbWYs7rEAR6e52hubGyCzDW8wEOc1lAGN3CA2SdJHmUXwu3NgCEgF
MHceaHkW/6vkpd5/XdwUr7eDIUgfo+N/PYFODtuqyIfcnryvjcanNa9w76Y1B7bwFoNBH4rjJIS+
C6BGxGH7oJ1hruU9YPBg/Tny0uxzeqe9OSysqgwk1i2EaobYxnGOfaZq/VGixCPpr3ZT+D1RC5yD
SmKKmT4QYYdq5pCbgp3X03pFN/KGvxGq4FHTIfO1tGAG9IuSlOvQDtFRFelgh6eOT+VZR7dO+npo
0KRv54iPErivs+vKvHdLIJFTI448nMND5rJRKyngcbwZMBifP5NqXS2avrX1nwVs+xFIbShyLrkO
nfJc+TVoeD8ym6xMJRnXB63KlpbNgNJPeBTcTHSYx8XnEAv6M+BloXJ0T2SzcibkN92e0l5MQBmR
1D/frzJSokqox5fc8U+VI1XnclC62FK2JDNqNWe5RM2WPymLNGp9T3Tm4XlJxDpLaTgThtKr1wyv
3lDPjpSPw6kEBq3I25JHqMtZqxxEdo1QW+V7zoX9BzuoMIVF8EiiDO69kWxCQMIVhcq+Li7sebFW
CLGRoT78k4HhUeZnXWd3HUr4SP+oCgg3FQ08ixTq72f8PJnwavBTnsk2t+qPYjUL1jBBE6xx5HGV
Wq2kOh/a+/uYnrDUnRAXr6EjDOOHHz1o9n4b+O6C3Y2uSuwC08c9WTO+NpyvVgRobg8e6he6qYPa
gXkAi103iOQSHJ8GAP02h7YGCuzB8MBI4oW1SUhK3GOKBYt3UtdtlEic0SVi00P18W4MPB26IYho
r820SVS99oP6mbE6eA6Ub2Cow0xwEu7sOSKDiKuShw71NoSFz/VbQtmTdfb759HF7As0q0an4C6B
HNERrMKgjl1NVpdVxvapUN1NU+FmSGqbylGo7XWAnjoR+c+hOLiURhQwvMGtKuEe1/o3wgFV+IhY
RRT3vCvkyhy1EnOYRWNA9QCYmsAjhmNe6z4twNa1nHKw9NsiMXVwnv/7lEH5Zb2pXPYMp6kkmTzb
qaDVm4CyHhPc7rhzpDxdWJ/ZPT+MZzdiT4LgqBU0TIr7tFpgBsH4Xe7fZMBX0SBM0qSmmt9fw1bL
XQg1bCJczFnONw/E/rHCjKGxVrssDLzwKlD9gFXs70PsH1q27wtNFPWFJ14ISw+4aGnueFSpIzSM
Qgn5DuFBPF1e6Cr4r4foRoksYKB9olPOs797WFMI1V3AH7Fol+3kN7vV6l3Lbde7hpFzK/7YvlZK
U9ajAyNbgR9hwZIIagu3K0/B4HRckBReg2/Z8jAnCXam4A96fnHkKe4vpatH5B93o8ZucNLoCRYZ
NuGedBq8wnlADOpAAQEmgkVwIMJmQaVnqZlPZ8AuwtozMNdVQMuFHf44acWuCw1yzRD4qCO/h3Yn
nzKeUx3n5GrLY77iT2Y1lLLx1JYvnklBbysfpd2dfrrl8I58HqRgz8RRey49ahbq555A/TmX/VsY
TqfErWVIDgLt6AG/KAoxEqIjtOH3qqKqU+1v+ygZXTEzF276IL4iW7W905ExCByXA4uFK6wP7YS7
JzWSX0MypLtskR9h8os+4TO+iTIDI28H5yKi/f9KnJkAtE/6S5w1ttGxe8VwuPRxSRf1xVhLiJT2
91AqMsUACjCS0HunM0PMjb0ZGJ1eiqhpJwvfmsPhXZjWLPCl9thdAJEJQWDPSrj11IaicrM2ekqc
jPBkQxYnJkXlIRrOMyrZbW6l3bw6QfxxaUcmz0BZZFfHa5mY16njVKqoBvKJXPesnK2pk4ERyt88
xOTQ8wWUfl2tNP9w06Hq7BpSJ7WRxqucLQTsFP/h3Nvo9Uo0B3bknBc9XSoDasZsMBOa+IqejGdA
NS7Y6jWCVDkSXZ7wOSUY3XVeTHIulxq+CErVMUCptN20SIojBhN51UCfUJkVudmixAvL2UkCuv5S
eNjQqLyIWXzNjetQ4BD6JP2p5hRt3vNpzGWEfdv4UXyH+1LjFPKX1ShY7g/ZEsg8HU1PsyBndTnh
z+rgwEH59+qP3v7EDHTqsL90lTJVA6EbjkKOo9isJWKBkCsZ1dk9bZd9Fsy+8inLOTQ9BGWAK5Eg
PeRUYWTPBk3tiAvq1ZVRn9RazE8DQohM+hzfjgQywPzlls3PeGejY2fR3eMOipuUoUogdtekUVU2
c0G3JNGITNt8Mdwh8vjcjz0RkBFCYRWpAqdsD/d+ZNqpmWlKWppReItfFM2Uu2LzI2j4ebbIxrJx
bXw0R9pbwa40vW16fAiGwv9LCSHGN5a1gRRum/B3UsfsB5GCjYE8yPdaq7h98Y9mO7TBufsnTRHr
hRmnV+uR5uhpzcCN6BG1xttg/4GgLdv2H7qMR72KvCHmjMSBIb5SVxpF8iTMbs4NW9nVvuVAu6mR
I72cwtjXgBB6YLWmsAHoMgGC3fQMAPjYUv4fFSwHZRF0+nvGkAriBmjqz+caMQ8vGSxt/RB0NdVK
NECpJCh0eGBVAFTWxPmH2ZQ8RJXZ5163HFZRhIxyZh7JN8tYLrtI5qdwf0XWmL+buD2gGMnPmP8X
bil9h4peWsJY6T+o4WOBitr15e0DdePoCrcRvTk1zUZjgLVH8l7557fjl1CsFixFsgMqot6zyr/k
0NGEX6VXZdnHqw4oS9OQL8QTePIVLeFxpBtHehiUywLqtV0sG+OuYZoRbowqnGez2hrdFnxgOud4
U4TESrkQqIqgFNyzmGeoPdKkuNZU+S/bD02iQl9Nc1wTU0OyIv0Uhokv0BZCq7b/jmd2ot8Ha98s
T1YEx+eEuU3ogmXZso2PkJrKXH94gp83dIUREE8ZR7EpK7jgGDO5h/65IPFFF26m3Zzx+IwPdssX
swhWr0Cya9B7GFhjGjAscyxZaqtifK5D0MnPOVRyuzZnIlFCqjkXMRvmhv25k4EZNgCxlP1R6jdB
YdcSoNke6hdEHTPTCi0FI/d1co/sYavgHrrBZeFldcWUZFqchkVR/Q5kxX32GLxReSJxSdiIhhqW
vRX0lZGGP7LOPjzNzdWSX489YF5PJY0qh6jgaJ8bRBYm5ztibz+5Z2c+r4EL01aIgH/pfEXHVc0h
3jI2iz9SqUL6dMU4T0h7npYhfHW0soNf8llp6Zt8qOfhWgKG/AgOaZ6TExemknJPpaNg8MRqHt+d
FIy7fL7l6EYUdPYoqeYdaHGsy+ER+zgUIvG0I8JtHaDXQQMba78kIvq5DJ7o4C73IkQjqCQ7s6Jf
K9iCMdVUm1yt0y4j3Iodp8S2M6thvln6qfGuedJNFWwqm9+6YxgfNXbbHGOjPd2ZTUYfKadClf/m
v+UToUYGnQL+TTFjD5Ki8Zip4GSpqJ29EAiY8UVtAYxM7aCoU4JknvHGyNPiDR0IUaL/M8YoPdfQ
snf6MuIXGN0DItu17su+202T8/QwOgIFlZjM4NwrK2U21SbuVvaC0F/TyH42s8MT0gswSXJJhiKc
jiF5kUjpEYpQAkWXTyKaxx7tx7bxaTuwyhK2f/n2EFN1Sx/o1D3J5bc0wX1mNgYZg1ZYKTCQQ4vE
3FJeghfmE75GECH0e5eCPDBM9nxzsWv+FFiSclfzgBCg2lcLqj4CAWY/ocoTklIeuhIOYu44lIEj
5+Ewzcf5WTHb8RLzQXQ6skoBhpcMn9PNlUCFIZVi39+y2ha552QN+iVzW8a+qziBw7AYbD6/kXai
0K1FDo6NVSly0JnO675Sq4G6h5dQN9NVnl/0wA3BhYseYkIyrifTVAESuP/mJbHDp84+/i45/mOh
gmAiI6n2CPid3R+hqPSgmAE6LQLR00vC5rMiDcj6ySZvWwl+6DX0tvwYajdTgXZcRnzWOMX3gbEb
HRMMdQX8VVpeXWiCSKNlLRNbx0tBL9tx3TiRHsFUHC3B15VkG2XbFKCJ8qVJLjuCBnP7OJQHVZt2
K57a1lX/As0nS1W7asDSeJaecRlZKp3IYA9buqlqACD49rpiOrOmw7LV68eF+b+pY9918UEUdV1A
1bGDWU3CskqwXokfJ2F/dG+X8TVWmGNvCXu4LhJYYqmie8djNlcwYTNjZ+a7Vb4unLGbj8OFdR8T
ArPddvvxkCrX8meM5RsfKiU9XHbc9vmML0bnzn1foq+O96atsXojwku9uRVTrjRjA2EU1E0+CtLq
1yHwRwle+IoDzkRbk6dYxvCtyzQafdK1U/77imAJP3HUuqq7/Nn4CObzk2qo7iAHsAdtiD+GgMDn
47vNdeZMBGGuM6L5nfH0r7wTkNwNfcS0fb68eiTQoXX9zDMMdG8axnS4kXxY7oadQNwcgh0Nv/CE
tMGTL/Qrl0mlhwitXEMtQqUag8qgElL8Jsko1oadFpU1N/jxvBcpKz2/MEXqpJsxbVoDW/NdfDSL
FniNxEzsFYhgCf8b5oMkrfc+hGM52eC1xU4arsHkcuXtJ5ODGN4aNyCx5Y0MqMHdFxsm4t7C7zIs
ieY6TWImZL5634o5w1sygJa9Rqe0/c4BHRYSvosgo3A8+cRPb76nevCZJVFi7pm0JgHqMX9sHY5l
pgxRo8m88Fvisrje84g/Am5v6oDWCFBNO0RjWiFcLCNrVZHNdTpG/ONSA0MDa6LxjZXNFbAmGAyS
FYUWuh4+0he8ctdC1vymHa09f0BM+P/eXrhUS2u4oh0kOz4/dM6+i87Rzrwfvkzvf2D2EjmMCX8a
wChpDNwMHwV7OK06XDhDG5neMp3xPf6Q0WfrGLPrKIA7DV+bFoC0/kZVuWLo6TDumJJSTkDCZ7gB
s35hoFxYA9/2gsCkIV6V5nlJYZlYfnwpqnw3T5so6p/7X+KdIZDhHzIsUSR3YE+2uOCk7DaIjEHE
CQB5Z6LdTl/kWeB2XcXD7ia2Q54YFI0mBDte4nLiHR1ykb355K8nr2kbqKQVLD7P8Yga62BjeESL
GSBtV5J2kg8iCyDZo4UZMpcNMs5k0MlYqtHvNWWZgMyoMemDMXE2wcfcLAvj8g+w27kYm1Bf8MAn
lir5miEIQlkBHu2PTmdT7yozEv0pVPO+obnfeZQHhKKYd8MiimOcMfGYGqV/XyjRpeqGm/7cwrmR
CuikQKOnlAARCJoY0/gpr2SBBo/SM3HwE/kwXn4D5nUpqOXreGoKVV3jnh7WLs3BB0A4HOe8gHaD
ssvR46HixIRTtikCEJjG65UqKhZx99a4yXwqdSjIqk4lk7cvVwXNYMQswAn/orzqmM9qX79OIOSi
p+LFLYdZC5x8eUURa066EME3xd6Uq1TZdsdpJIj5xM/a/D0mwHR5J5xJjj2sy9U0GMsymqflKJLp
jaA8Muf2jVbHZrKE5m6gVJY4ymcqAQ1m95hJZcV1HNdcI0ZwitMij2QS/5GAGJAK/BLNMtaawNJq
a5M+9hZyl0+QSqaahl5TWBrVhHTUtNx2KJs4tgMSPzu7r/xPQLSz/QgQStCdzDbvirUMgpaa2Lwn
AnYN2m1KUmdKXG2rKt2Ln0mRV8H9IUUAO9gT5oY1dvzBZDdBFJBUqQxs02BCevsfwhe4w+xwSGbN
jVRynb9eb45e40BtUPJVNyJmNlwMcb5Rlu9K43ZZrMrTAHaXEYXmJuEZzTTjK10SYk/cDyY/wugO
LRi+EV05mTNkB1BVvO31Tv0v7cmy4vHAwrU5n9u25Lk1rUqOqqAspepKl7YAacla/wp8kuzuJbaR
JY4t54sEYzZWwv+thBW5XAMRjY8P6GJv0Ru0AZtDBBP4tBG2VynyewYhl4zVYKpbvM1Q4/Op3iEo
7ZwRtvMYgrFldT67S0iDmDl8FJT9O1P21eCBfxxb1r+Up5tC57ZPalxQooaB5gcHBCirMQHMlxp7
38SZzs/D24lzbO102XU7fib4uB1+EsyrkGpMaHbXn8zmooxMmX4/k6FeJ5GcccuvOZYvkf/d/Quw
U/r3j5fPXMVU7UmLCg0gR7IwKSR2R/HRtPQmSer7IqeJfbirx92esgeA91xlds8eESZpBBpZFOPc
KJlbxqUlVxrjE0HxCiLdogabLG+Z64HPoHWEe+iEuQHQm3Ur2pooKpzh3jECn73R0V3r8+5exjBu
tP2AccCBNX88yaUT5Sk429JALaHr+Y55D39N8Pjqibv0ymrjZqlGBDPm6GFmR7xEeFYCXAh+F/r5
sNmYBTh5PYvVI3XLZXMF5fBypR+3/H+oUgrgZDIYuEuLf/8MEpfDRQFAITUvKdwN9/tTeehDMeFh
WrgtKr41edpNBJANNnMmFMPKVHzte/cpOqZ03UV723ffKKPFCQgtZldxPKtVtc6RFxaaSVs+jCji
RZxiO6nkKzyhrpgZKSziUjYVE7Ib9QMdDV9v6inDHGzHjWXDBXzf9cPJPhqqeO2Gfge6bd04cRgV
vlwwWR30plERwq7ozD5ivRa2CRMVWa61xAuJm4+xlWy0l14FU/KOgBUxUp6uLJnS8nnew/m1Xl2B
Kf1ZZ6rSjxPTUL5OVn9hLu7n+u03BIQToLakziOSNRgkPW+iTza8ZExqi8hi/k+mPwczVZ5HeiL3
x9ZZBSgdoEdlacz3pfqIpzY1YmOzboA6kB6P0VnVMSs3vqXvq7b2lCiSesPf4ieDYT9TEDfnfUD2
Y72bDnK35FHGIcfy4P3/MTgwm1lDufEAZosgcNYRV7lyG7sXEPDvdCxHj6xGrvoOcG5LFMwliXL1
tIQmit+ERpzjH7jygIcvc0aW0eMd6lMDnfipxTIEoCnw+wHZw2QuDXUDqECKoM2fW8bXd8eIWNMt
5VWbDwh/UfTeqnSdftkcG7kM+lShkGns0BQDZ+wMYI0npxTdHmJPf4nknjhJjpq9wEoLFvvH/vcO
5BLoEnOHG9rxvWdRL+ksSlxLRhxPXIeG0Y0JHGsso8/lrFCxusZer++Z66fExPy4GVnXovx3KhXi
0K5FjXnRdUSJoQVPFPkniIr6m2U3Dmkd8bJ8JMYv9FhNt9a4V9KnYr3SetHV1k7mV4UJQA/P+uwa
sM4KezViXUxDI8DGqAJDGQ43XIgwCAZMcqR098DsaF1/CT6eKoF4R7XfI3JOAaTqKsDSkWZTYmix
ZX/zOxuUafgSihUZXjev1htHITLDPmjuAFT1NKn0mwZxxwSvnEYnjh0ALa1mmu4a5NVJF++objdR
HGouxUPxBsuKjpBQIgVg/LblA7NVAW5tnBT/z4EekCl7LusSuFAzotL/qjZA+Eh5Lgsn+d5kDwgw
mbMPW4wFkqME3hk66bowFE9U+2l7+EfCedBxSvHuhJ77tHYF9Wbotq2aRT9y5TC0zsPCJ4SBedsw
VjwHiHmQhChLslp2DmtI5/DQbVl3ecNDVpe19X5naTsP3sqartMl5V3nBxA/4Pb5m66SSuq/oPik
MobaGH/DWGQjyySm2iDCCQ5moggYcnzSyhFJ7wmaqw2vBYtp0+6QyNDcRUjWUbu6pTr4tqPl4aH+
Mwx5yal5KrVn2Njos3jr8Ys5oIyhXKM7uLK6cOn6aHwuFGMDTS6wgEwOxHDOGWySbEF6OKMbyfxP
nxXyTPONAbQIIzA7RIwy/XUBdsa0RDQS4lCj5zjpvATFZxA4bSJyuRVKWMfp0BoScZLcQZhup4oN
18xuNRc/e9EsT4Dm7SDTwqukG/Xe0qDVuj//lcU1RmIXI4Hr4QX8HP4ZKWrag3ca8p07OhkfIg6k
norpMljt9cfAzFEqmH/5ozlws+cjhNtZr3a/XrfxbgSStisYuJYkXNm9owGq7NF4/N5GOgzR5md6
DFODnJQmq3+ND6spJCTPxraGjGYU9QtHHO8nJqhEdWbZo/J0ijnmxDk84O6zGsCWLiIAxx5vMO/U
+HQCmz3OfIasfrdtv+n8xXvqE2wKa7WzcIC58rhQRQMznzzjzMCeuMqXD4/rRsk/F0gyPUQPdfEB
zYjNooawlnidfPJHoNTtCtbvCW9B7GDdwDG1bA+1blfHGQnXATPJj/rNjzzZIxIY81oCO17GkrCz
9gzeJTtsw0v+2ObXM91GWmoarwUbVW2zlqcb/AO7jHxwI2VXb7DWyDC+SK3CapMJgVT7OX5gvZp9
3kpXYzL3Jt+D5jySN2vt5m1k50bON8S5YQXVJQDA5qXD2z9gF/RnHkHwEc28N/MpKcveQk7WVZ+2
1JUATr5W1+qKUt90lD4laKcIrMGMP0QqX20wc9ILMX81RvG2gio6faZKwU3wK3084nvdmLASNWiV
DeP5l2pHzKRZEwPlNgUCjJWunguFFGIr58FtbWOMwbKMXP/vpUVbiZdm8DxJq37egrdhnYMW9QQ5
kh3WTI6YtkaNfd9GvS59LaHOn2hiZ1oaRw3P9qQFl2TbzWlatIyE3BC+AEmF6I2dcxsnxnFAsFjQ
eI8bvDO+iWJ9EmoAkCMr0HOH3kCok8V3R4lD93BmeFZ7We8Pwqn589Uou76HCoRxhF9t1Zu8FdxY
QD49bAUpwwYY12t4wPly4zwFRoCSvyu6TXOlGJNh8CBFky/XwKwasgbMEJr6aNeWm18rpXxcvxut
UETwgo499hEN7KrUDTLopZMVYjlfLCYZ6baz/g+or3rGkmbQypoqq/6rTUV1+pSjMbvpSoJTq7i3
GdDok3df5LggUKYCt92QPm+RWFIfyczJ3EhzaW5wQCZnEZkzju7rw7HXFRLBuhu2OxwCDaLEY5Co
QTX3qhZG3FKdLu6UO9aZ4+tdiXyMKmMAwjrCN87ChhwR2XKVoAr7xX1j7abxivrNtT1hnNPwNleg
sVqvWgsuQLcPjmOcncdWPJ28n29XH001weIw2Mehi4ak/ck5nFiEjLIH2N/80y7pjlvahgBKb1uN
7OxvdLM91or7r/4+zC+JqvDh8JG1N/70o8cjtZWel9Ie0oSgJTjEZ5GT+/dXrCt0IyHMjlgjrA6C
FOFZCfxzGlYv1hWhc0JnbbUspl+/+B2IjwDPlhPLfCHfH5fA1uKw2akpH1urR0ZZB5RKJEBQnNuG
OgVIdN7wyn2St3a1J9tqKWaPhsJMvYU+so83Kebixf46cGu88d2sd7Nd1I20OZneGyAly8cDWWKx
jzzRS5ZApTEt0VFfdEaf1mjxexJsU9a9tCiAFAtUuDB6REL0QOFsHZahlC6fHB5hXxjrFEtW9BvU
yJho6ZHoGOaKgXOWdw7R8g9S3PiNdIrtQW9ygxvaWTjg1A1eB+7fRZ+OhhxqW/QuKlJ9T9hwoSbj
vRtjU9dAgE1adaNXexeY0beMqvggD/6OWLGoF126cXJsQRzb9SwPEDm0qo9J/3qi0PKTisx2nfXX
I4gu/MsN+cNFQptIUhiJkSLEggr0UKzGnkKWTpmsUoigPsU0S28mkkmK8hpdfspKFs7NnexpdxCK
n8IV/RiCH5hDZS0fidw/Bag4xIF/mIJYNJLndUqKYF9sSzPm58Mh38en8NVeETzj+Bu/6NrzePKT
Q1PdBH7iV8otWskwBGa8bu/Bnp18jCJLKIAvmzjEB3u3zG7P72xdlXgg/bmS3M4JNLX6zY5mPLUj
ktTTGPJ18ZqhBb7sAiFsqBhqQgczSb1XqMcOd1CWW24EkfzkwtlVmY/xtOkO5bicM7VARa/KL8ga
9n5tpzhNb95jvdpwTXNW+RSoDNQacYEcSpiOTsGkjg2rP9bh7ytnDzlIPyKlag0CGd1IfGiiCyds
9YMZRhqyNAl96NJ7CPrWMNxHm6BtFJPl52wmt4WpzSZA/44Ui8XQU6P5jBbMw3WZVkkml/Z1YlkV
SQcRlqAm96RZGsczmhW9j2InaQRK5+ROn9xteln40zRGqwnqsxsChDsOG1w65IgpfDpGtWKFeONk
L8QgyL2w3U/SR6+LMwxKeOS0qbCuZYvdFImSlf1HbU4Vlm3nqTkFKfH5wjpIBUAzw8IPD6CbpxV9
KY2FQRWy/YYIxpWfpjaKrciN8HdaES3kN7ue/5Yvevxc3HCU6/wmJCE7TTnCGu2TnzhPaUksMgiF
xKqMpbuEl8/hBy5YQPdwu8fN2ReCOu/AHfimiVP0wYiRIN84iIfeZeuL80d25jeiCVkdsKNHmswQ
f7U0NuaFllFeg/kzMO4Bh8qiY7oChtEwl6oVL32pPE57w1Vudr6UEWPNshP8YyRrrco0iJxSR9tw
/3O9KNE35UXzB6//wH+SB+CW21vnDZSjIuxAe5aV4Jd0CeCycM2GDye26vCnKFpVJs8wiqpG4426
P+N+UIAlWhDDMoe99HBJQXgqRpeedbTQh+nwJSb/rKsu+Sx9jXDXIho3bmGyriGLRzuce+nnFJpA
YNJMTDGOzet/Bc9duHVNeil3qv4NPA2ui/5vTltDz8LvQXRWRS+BfndpCH75sX9+QmBBCo/yYFWb
LyjedXq7F72hsjwoYfKwFXcj3nuFK4JrWVHFCghutch2bsLLJxVHIfM7nc2mT3e8wY34w9wLxO9j
qdd5HoiOEom5dEIcbYZHXUVcTIRX6m25paC6GoddbTbkWNWKrq0OxB9vPTSG6LI8rN9oH+C6Uecm
tQF9jmIVN1e92ju//NR4Fec5jm35seTIdo/eF+ckn82ItIJd5fQhhaPkd1aso1iQEVfUT8x8t8W0
jO3pNohv3oV5s5eWbcQKb8NOy9Uv7sJXqL3K2aU28qXxqacS8xH4IHQS2oZdUXZW3czGFuK2Ix4H
ZP+aQDPiHtJ3JmOHO8wM/F+FSdJnEuDesAtJv1o6+SvDhwklGa4dtxnYG9ziF9r8jL9I/lMiUwzh
NlzidGQLUAPGOk3co0UaVPga2DRM07647gjV7m2tCgJ/V+bq1NGfwgNNFa3haiQkJtNVxYzbA/mZ
Lv79RLB8BpVfmv/7iGFHjE5qfCqo3+bgNJZIo1bD+YSsWQU9Bmy7PzlIJEz2HBTpPHjliuZN7gxk
GwA1YGkEPL4LJTFdk38iUJJarJvtiVFXBkY1ZU9kO24S1fAO9uY4s4ytwdsJvN5pd1kvwTab1VFU
PEFJCNl4JkOukUFucoJWaC9h2B+WF9CW1JqmGuCumRcAVXhOOkeFmWWtaNMuFe6RDRme7bOOyKKF
WlXj1mT4TMbccfawIUeMhzgwxtA5VyP6yjtlCTNTLMPidPRrORUMgCUVVh/bBCpnDNQ11IzYsjsk
Bg9lUuwV+tQYDdnuTq+FwS/j/rw4kj9wajXpe2S20JNQGxnlINa/e82K2YTokU/I2wex2XrjpIv7
k4ofpCIVIqc1KF9kTX2SLG0q+T0Niiv4Oot5ZmMmRgBU/tL3V98r0gN9guMF357AEnsiwPCn56Z4
5teZDwELr0W3ba+UiO5TDq76jakyiSWYNw7bEWfnsXax879LbJ8HGVaPNFIdPBEDTS++bYRX0jrs
lsvm+YKCXW4z8+YwwQOq7d93ZLXZ5WswtZwFPTUrGnbdv/MdI90lJrQkCvCl1dd9qnL73KLGWQrv
7eBtEZjYZGuvOb3qwBLHO9P+577M55yTlrrIt3fktSfT1h73etzqcGCfn487FkTtLOrJYS+GKZH5
sUg7q3WWMS5l1iV+9QY8q+x9VOUNcMcG7xwi/oxSt8V3+3P/y0vLYlinbRdy3P2+sc1UCyZxYwCS
Zw0udbwt8+W28qlEk/QjMW+DI/E0K7I1Ipi+D8V0sKIXbUqecAaKXnvMLiRTouS+gUEFE/20Bnls
pg2dFaAjA52ODPD+1bgJiZkOUEb/b/cwTQTGSJR3Y9eY80qkU9iWVrXXRZXGeybsR/8s6Zcvv3Kh
9MTP0Z314gbwv0WP7wrQP8wb6Z03v1FGwWNk+1E/g7Ley5eTZ9xNc40bw7L8KmXotUKEnVZIAtwa
D0huBmcpCwujK4+AzmHfTlrK50FN53SQfcToStwAqlC5rhglxVACyQNzcLQkqsoLHYDDGJLVuDSr
tY3B1+BspM2hSPTS/Fxd7+jEIqJXsbitQpycMbXO+MFm9Ys6OGe7BtVT7PaD7Aek4K5/rFVqSBrS
1RgkzlTu1rP20i+5imJoRNl7wwWHIxVdoBZiN36KFSS+RZtrMY0CX4wYPxBqk9d+nS/X6NDHJZJD
tvIwnNazjaL0fS1RhAUk6+oYTHuYukrjFcZ9IuFp3GQ5zznT0QJ8M1sUhQfKl661nDeZMsrce84g
RVgFJmBhSwvCHBzfcMiQ4+Y+M4wHVd30N/KWlBm77w4mVNPIctLX/3KQyITABK9SsdhpyWBmqQ8v
P7R2mbsL2FgdSGF1fxk1h2qtOSIJkToB+pZ6yoOs0nOS86LpnvunfPk1G+MahaJ12bkIc4k2L/Qy
B0AESyOXkdHewKS7mDOoMF1oJyI3ADSTJrpCKrru6Se+6QIbkBjkWlre0OjSLMGq/DBYyGWjcTt2
v7JkzNF28QD0HUITeWsFB8wJTvQN9oe8KDoUwgHrSlDpGtDM4ydM2WE9PSRZYuRdrbDl/gdkGCOf
anKF8BAp1G8coschx+W6B4q40VDmN70czBBaG8n5S2QwMmtvqvCLhNKOQI6JywveJa9WNVAqhFC1
JTpjG6dEOcrk4igedk/bOUYnfJso4ZypIxTB5PDFoRAx+AzH8e5y+a+nBdAUCYoM+ifRUkQVwaLi
hGjxGZkqWq2KK6uDWtfQLYI9W1S+qQJOlDYy7HKbaNgOP0QbyFCzfwJ3DBr8aJlBwdPFxNAzIYCM
FjmzVqkWl7NdwDlRw5VTyR9PQk8WGBvkyX3B2lGd3+6/AIrS1PsN/qTfe4VV8OvhXzDklAocpysc
D4UHAZcLCk+UqkVqUqYQ1ojWXo/Xa6U1YrgWhqLRQPif4QZlny06E9UF/xdASoZoyJRv+ymlBlmz
hGld6ibrA+wX9m1HQej6CM8JdG0Gj20/M2/f/qCvh+Ttjh0BAssuQx3YkYLG55CKkjeDXj9e+CTP
IfAifhQQajbGHQD+zIR0lY4xKs4fOr6QS5KpC45upQc7TWNkIAmwD54HZTzrD6yzwPyFDUeAKPqL
rVDKJlbfwBv39AXsqAksDvNviCXTsgfONdoEQAXHIXzwrdZv1zzaUqkD7WDv0ccqQdiDCDjWMPFH
9LIpr34yIutbhWX6tVDs5N2o8DSWJ1KL8XPgmVOtNxymcUUtmFzFNwb78tJuXkS+JU7VISDNFaUY
/+HktVbr73Js9lCqR6I4ip95Yc480vTXJSTmtO4kri+oOcgG2Wr//9LMr/U/YgCeml7f9PJ4QWnn
/YVEAK551OXA9FllU/7Gof79ZC2O0wwa+XuPW5Uy2mrh89LTRYGuMimikXP60/wBggAN+flXNIWN
3LowtC+5gh5SpwQRBsIsqOGz1BD0/B1Vep3CpIXB6ga1uX6TcZr1naSMz15zwqrU8iZeX4rlP5vA
HYKP1inP1i+jU0nF7LcQDYdxQjdA5gFLYcjOV8lWbV499ieimMaUn4JJ9yfHwnH7SKWaFSheqrnr
JZQrohEwjZezueXAS21haf2/ttowo+tmpylm1nGeXVTSIoxHr8GZEcu7+jHXUD0NmhVQtSKm9SYR
YCjrI3m0Xpb0dryrdUVeNWe3/xT0EajnRvKl/k73ioH738xvrGg3UvtXO7ErhiqIUzdOm5JAtfHq
491sF94w8Ub3UjfGqCgqFMx1w1vyLr9Um5iqrDMHcsdm5p8WMIxMHtp/XLmjYm1xciPe5oNDkSPh
CJIFg3AA/nvqLcvzgEH2iHf2XVhqjzqYu9pN1wzBFv8k3W1iZkVM5KmLkmjL9oD6nhoPXt8xeYsM
YfsG3Khjp6k9hTrivVNW/SdZYNKJF/yFAXozWagyw8c58NN3OwtNKtIH+/H/R+z6XaINC6tZzjeF
QbYI5MpX2fl5NNtSgCQlsMDNeNkFuAws1TtvQ91ritqZMdK1xTOnrcd1pmeT3vPxZQSqCQZykegv
KR597A5If7pKkdENmM5kQdFabJK0517goJ0PrIlO7rO6hClZce7TjzQjRIXNcFf2aB+eAGLznCIK
3Wb8Bkv//rzGmrt9QI14wTNtJNyiBcHPvjaPUtIRj+skTn+b1nWzi/lUWA07JZegf6ivV+bRbi3V
3CqzA22XN88e7E6gZWGU9DD9XoUEw62sIPKN+LP46Sce5BevEHNOUKGs2ppa2EgZwvDdTNuvkFIa
BdmOPrmZi/aFE2aprmMykrkM+dCXn3BviKVxLD7TH/uUzlT3YobUXVzQ8LQqMG7bOLlZHy77D9Xa
lqx5/Eie0EurImgsAJHJQwU6fC6/L/cq4McV4G3mC+RcVucPOzJlkoyoIC745wKK4YQkCO6NqhQH
1NkiVToPB3zAY+XPrOeb8kB/6U19M26/hjWAKAinb0EfcvnrJ77CxSdLHlOrweJH2evCumEInOG9
JJC7cTv5D7zmtfunvW4BSqjkQ1I3p5jlQT9MjCqdTomaebzQhVbNRbVR4SQkpuh7WIYubFwaIFRT
WKm/TtySu7ZlMWN04zcJMLkKCcrPcYKvE1F+jmvZODwe2OCYsLsK6X42khrPpPB6MW/1Nzk8x4QP
F+Y6VpHXta7TU6APC9MPtFlge/5JJgCC57xUWq670Bt3gXwg4/joQ9TImIjTeAX3XWgw/Nh1QbKD
1cUhtFdA8uMjH50MCdIfK0xMinpf4L3op/7a5Od8Az0IXVnpMsLBMMw3KPp/wwx80OOzn3QwMmvq
4HXsFoNpySDcX1XxmAyCTdMoRvmM5wS3qFRSdLqN6AmaldWkYuKhkkxoNyQYTxXB8CNpTcZZEKPT
xUjmemxFyihvel0Oldck3dGZgOieRyh84zRNG7ezbCa0/83wwnLShLguaticzJwU911LSp0YA63m
VyFHEyXCULKSnwKthEb1grTuptS0nbEXxxCZo4HHfubaQ3pvtWdIrAjpfgK9chOW1A9lKkQJCXBl
/DaA1XSz9OKwOed7nD2WDuZ8wAY4Ou39Pn0h3PT/Qa4Nl+NzJD4H/VV6x7dUh6RNb/o8wrI4nj5A
BBGtl68ZTOmNM1U+xpYNqBVouOLdFWINaxGEf32jHAXfXBvDzCoH0VQaQcTJfmD32RNk6Kcd2EMu
oGaqG2jzwrrSSIfcq+eQ17yQdyCAX5Mo1cfaMR6ElZs7tKaLZs/khbr4DYkA0kxIPipDLgKkkZen
aM8Rj9OF4FHXlolTm+H0CgdoasKCWru/aYUQ891Jn02O6ePtMraHh/pMISQDclBVeVEdQ6kwOnAT
TdSCjP4GayxvWHLcWAU11sW+0KARoN0XpJm/l7KMcHhtcNfm2mzAPTN2AbXagz7N6t8F2asv8cj0
wXh5GT6hCAnubW4QoIFEMR4VHlnbP+4g1OdFLcUxM2TfxJAs7w/ded8KdbWh8zovshtnFVuXAzGZ
jPmzZm1dCDkmVUp7qRhO/WYT1mJF6GYtRPKfo2+YLJOiclbjODsWzTxOLe+qJKaqXDWJhSkoONSk
2Yx7xgDQfhwRJ86UIzqZ7Xoz3McKYxRj2kTQh8K+fWmaFkk2Tn9LRkbmQCwsSGyU8/GrM/FW1qT3
XLHsKAGi2Zy/XmbriAZ1m/gyP2353PUUOz7tJkOpXgaLMHvirmLd4lYFC2ZXDuuTJy1/+ah4xJ2z
WkuOCi2jfTuIkx3mfn9VZfvBQFPxui1KGq8zUKDvrae1oMNBpw2/FdTtYURHW4/U/dbcFqtrlHRb
ZkXQPbGlRJkuHsisXbGU1MfV+nqxMdAj8nb688gGLQm9zXNEvWqeJ18Ru7dNd/3yxVet0nCUu1gw
hOeEO8noeqUCT4UNRKDY7mgRK3M8zQ7jJEgw4PoVK0cOwqDHff9ehATF0uZov8yDdZv7tNA3SH3K
8rooKmzPRIVuClJ9H5z+7Qn70ccixoDmBr9PDT/A1sDpzcxW6wrr7EOrVY1m+bss4FnDHys/rNfr
FEb+DbYW6fjMHH2E810IUyZDFN2q6rDcNaLkN7iSPoKjjuHnk9pmy815XpBTzhFjjJI+np8MFEi5
qquzYrVGHndUOnyZJ84WvqYAl9/sJlwi9onrTkSoKjzQaV79Ub6VzvomQeSUHcIiaDZvrTh5wdnA
s14mO7xN05VQy0Guw7KovJna3p1BHaah/B3f9YW3WqyPOR/eAYh0wp17URDJWe3habmbAksVWfk2
GY2Db/njXFnVG+CfLchpQAbgKONyV1M7908gxjFCvYYC6uvCyEhbbCkNWUP/zE8PjhY6IEcwYKPJ
Qr2V6x4IuphlSoipoYKrJT6E7sF+UWGQZIOenrfXeqor31t+RWA65l/GAEKbXBuddgcAbR1QfldJ
cO1gXzFFaAbLjOFO7RO2DyUc51NjItNeZfhr3CsPYsT0GK/Ml5xV6pr1BsLcjRWKrBXnjmzsDCMX
TvCzGoGI8z9yh/zX1F9DMeWXT5sAmKEj9ru3ATT3u17ydmUsmYer2Gag2j6hKFy/BkR9Pl3R+9X/
lDA2QIT3b2sxsAPfc/dc1ON7E8wh+rBNV6N+/nYmMI9/ipTZCc3hZKkr9S+9ly31F+l99NSWT2Oy
vpYSWZpkDolsaGMWyo5DAVBYXEERsssYWLQ6RBAlIST5hEp7QpX3wS6zPH21XL0l/i5ZnMJGBWoZ
HrYMM4cW8Zai+he6a/sknQjMRrXo/JGbD67r5FJJtgPxs8ZZrCcEX9Hi6snBLT9vP+RWllR0b0Iq
gkd3GWTsz2qr0OcKrGDesJvj2dq0JL6Bdpsro8U1FRib1a+CuXQYCeQLqG8fiTPbPgtWhSWnNlg8
Q+hDroXfj0AznfBj5mDxc70d65I4grl8TzCQVVrJu28LpFhlhMJSsjpd8h8SQ3Xmd5GWEDaPE2VE
IQGLEGBSKTRhqAfY+NKxJJtdZzPYEKRoJ3krjZac3qW1HieAvEm+067XWn/V+oGLmOv/VvC4izSm
OuK/kfDDVsRHkwiey2BOsL1X1f3NgLktPpfBMuhQ1y7TFb9vx0cVev+ig1Kerd7u4kzkfwY8LLX2
L/izosk7qRyPModZmqC51nmbl1esZD3TfnqGZL7Z2hhJiiUy3jytR6AgT7kLyBxKVqeiuWUnADQS
OZyoYsLw1O6y02YIJxFo3ciAuYRQTIHob9vxdGFYH38Ej4ObJsyyGl8bhlYlk+ba3qBCI7HvrYzT
cOTpZ4qC+POYPim142ZDozHfqdRNAWav/mqbUpc85o87zwvQYimkMMaaC3V9M2KWkGw8iunotAyM
FgBP7ljO5Apdg3pvm932H6dEm0qf+C0XXyUG4f+0jpsusAh3tECjONdNKp5Ufj+wC7MztgI9Re5i
54NS0maA/Qzivv6Ny+UPO5bZuRAU9sFoAGx+kt80XPXSbWjF35FAwhuc6ozfAqn2J9/ZcY1ww+KK
NT235E7wGOriwuNSXOtN/wJhoZXC0rHuaQtjd3d+LnQS/JeWBfKOICVbM3W4s1jLuY4Yzlqn2DRA
q6PKJCue50HMpsxR8H8uV9i3W/HhNDI+Z2QUVKgxhKlfJzmWrNGyNNBRWUd+KPyUClTKZt3KO3AQ
T+gXT2vLP53Nfv1otPe7WX3pRsZ4W5otDSvesIITJn1HE8NzKdzOEx2XbaCLs0IwV/1L+3nwvMox
8twZTyjxT9BiQPsi2/7K6P9QEGfGZLOR0oOVqc4sj09sB5MT4yxE84fJlZMHtfbA9F8REdMmNzYR
0vuMGNa3Yhx1Zxe+OyW5w+QOTjE3AWovJxu3WSaD870jHIeo/CMWlVNIPhkhF9BjdTUjn3k6I9C+
xTcE5Q7gDgcfKa+oE7NiQ4r6gJzHf43ZeCtCklX81LGy6CN3xudZiGw9p/wSRFDhBJ6TFLXAKr8x
gOrzoscXAzWM5VmhdpKJly9sN6gshKfwwbNAslv8mElA8QRiFQP+ZNh+eXMAkZse5lMci69mT7kd
X+c7Hvue4CWywYzyGmmAhrA/LdVrG5wuBCgoNeoHRDSWHHAo4tAyyoveFE1XGPzd0zL2bLeWg4sI
URO1x8mWbaH0C9mrsrwWXumXnYgPTlncdkHQ6sGsGnJtIL1iZZTL6F0CGCWar2y50va8QDMVkp18
lH7/9/TeBwmIHK5GSJvIp1EMCslJR6SjXPAaJyWk4egYBLCTCj3Wic7QaXOVdibdsSQs2w3B90XU
izKGZTc+CcwhI4E4CEnYPBxOhXvLTCPtNf6sTh/dHCn0NwBndePYOXQwudWdxm7iy4RGbI86GRc7
Z+jWNMONU1DiHWW0GH/3kSsXJNg5ROeCqTkBWGw3j68BIh+9GNfnbhTYlgeGIaPrI++3CqPSmnwD
+TKnxwRolzRXrQMEJezq5CJvYT6TJFTNMizMK88pBMsbZ6G/dowhHfV66d4lfRh1ClfG5YIlKJDE
X4PCM72OsnKbfbIPytIibriV4Csa3/LcBnJ7iZiKtBcJse82l7OetqF6qkKNWZO3xTP8J0IX4/4z
iCBlzWGnhfkk1A9fDF3X24MIZxzYujm/CEpRE3HESJJAvst3lmqqXq4d3vpxIkatY7JW2YTzL2xh
/ovwXUEh4+2bsTPnCwDyhCOzUikPOyP4itSZuw+rfaQbkohrcqktUKegWGIgQLBzoX5xTwI+Gl1S
A0veJgG0fO+nG2976yw+yx7kHVx+nnU41rSaEIUqkaJ5LAsjtYWl37YL0FcVBjpbJfLBk06Yy9NF
GhMzDBwRaEuCmiBvrO1CEVgu161keM6cj7y6n32PuZZ5pQcnKieY2CzLZtGkdx696m8JeBw+QANX
oYJLrwxSKJRTKfQfcj6Olz+Ne4IWdbSVwOy7axyr08YckumgH/6xZjQmfOgoZuw/DXitTYhdxOWr
CLTvzdbGA1RZTvODksnkxmo+IxGK6UrTYQgJHV3zyBHPZJUVRdbiJii/G75DQW8B/qgCnA6doiEo
WguCAVPZa3exl64h4eLdPylfR4+GckHcpZgFYjjS9JsGeOXmT7pYnR9dSOxzLz4LyOMhE3GPSc/b
n7wIHii+wE6hJnnjiGyp+oKqSA0XWJ4Cgn7VHGtLE8cbEInCYIVYVscMu7Cc5wLH0JkXhW7PYc/u
aIUwN9/UPjvzrSML953zVmGGmIuXV8fnQ+kT7HS2/KX/gDmZPnqIcqrP46PnnVBn1obfOAHXtc7X
/c9upn0Inp/bRklXt82eAo33V6oYorNvsrNWx35C5Ia6RHbtYqFMl2bPiSzHm3ZlsH0RrxXH0742
7GS2Ks2nwfZvShGLq5mJFass9s/hqkvTfP2O9UaHZRqlfD+DBjwaCVGErMhUtjtWmfdcB0RA2vZD
wrVWOfRJcz4Z9yMvtUOdRxTiIqP4P4zH6tvQDBYEUQTWXQiSIWO87+JFGavhxspfYc6YfNKKPykB
hm7A/sewz7TXGQCmnWybI93vIjCA6PHCneZakioZr75xf5wgjCZ1pGVS4Wk71/grlMzkHObOJ4M8
KEoT4yidYJz6xrex8RPkc6z/lsoVKUDu5Ae7ALoOQbNg8zrObNvlLOImtyne/N5k5MzK9GJaiuHJ
O+ETnRKyJBF0TZtkVJEBhqG7a3eUSdqPITVdl/6Kj/pzVczwl3pR76rdOpz0luceApZ00She+uFY
sDckXPg9MNxiLPFKKe666n8F2oZj0ZCwtQ7f12NFWvUsAhZP3BOryIyoyPiwfkO44KETXQ1DFMK6
888/2qMDq3XtjGBZC1lwd6mMCGTKJ3h/nNdAa71btM+9z6wjnpr8zgTEfXcS8MZi/Ys1SfyeKWJA
J6O/nTc6MZ8JenCZ5S+80S++VMuIZiZL1hTguBBz3dwI5L+quvrJE7cMT3LSgaMyHTLksG1Lsrq/
KqESJ9EE5BJ6H/ZK49gAQ3r2tSeBrtRW5h+0eTqO9oeXKPWlI7unKQmwpE8cJ3LHkRiCVhngLeZ6
/yxr2Ia7E9FhFmVR+53SzOP4rIGzsQfW9zkr5WaAGiAq1GtzRy9LQfT++spe1WaX1moka0bMo6Zy
qquM9Fyc6QQLL7g0jdb9Yw94lX+uH7UKGbuQbd8SdIWfL7KoM6H/EuC/DlAK+QDMMxIHwHySYDRm
4aHNqY+TFHXDkAbuSubQmWz8iMBZOuehsehb2YkOYqAWc/OcqdniXqEqB8KvEhcaAkKslQBvcAgd
8QHpSsCw36iONE6udbI0FW3KlZEGqC6kc5jt31eOu3WYm9eqDtQnAPLBHjnsgs2Y4n6fk42qf95R
D8a6aVd1bPQsvh1q7XCLxHz+hD3IKRrC77xnJERdpPLrHI0aQUq+xsAf5MyFkZFqvuTcPIe2qIdi
qqczNH92gcTaaDGdJITAkJYbDlvTgFHlXjxreXn6vb7u+jkQWPiMO2iHViFHlP0kJ6DhMTj+0tBC
s8ZGEXVVHDB9znYMTdN3nSeCrSv1T5MB85hnOrj5YBfV89Rz0P9d4i4r4jiDoFhUVq8ENLff2qPJ
2vF3liayfi1UphI6kmhnyNgDyPlJMoWos7zefgNRHHdQvdsTjfkoM5aHwtB0YwN/SIRcfWPQJwHG
7UNNTtEzMdeCJJsXAEV0QAJpCTRZQ9jZUP1QtelaTx7iDkgQviFs3//uU82uEGecFigl+pJskwtV
2gO7R+j3gEd7l/GDYksqeFn14Xc4/VjmVbK2og0ncY4W3EbYxY6yfNIBONw0dfz1zTCJR3jpPbsA
zi8l9udc7tV0nOTOPpedxf/yX8DbNJ8ClCFTCMFHopjqkwza6T5Bw3Lgtxo3WJnigGnWLjV+s2rk
IN6+Ac4Bl+f6ZqibaL7ztokdY+NUB7pnstRt28lA6/PZSMG6sobZhBMC82YOOPUboOnSZcfDpt4s
7PJdzy8pK39huQv6V8D/lIUN1BSE6b82qnMakeOVzaJx/eM5vZ7YXrZ4yflT6iwP82e2yOaVMKLz
YUyrmZFhsLF4xJ8AtwgB0CpJuIEGyg8tJZSvzLE5qFmNQODF8Mvy5zJk3yCIqJqfSjKFulM+5Ziu
Q4wHKuFW8ccEdADOhnu8pNCsPnbvHar56vgud9auUNCjv244TEsAS/KC4+yqQYjyJG3vmd8Vv5EK
y6mawmFvtiBJtxaevl7ZHBWUmP7eVhbzTze4CrAP5SLQ1HxQnMZDgLsI0JfE2eqxJdH+j7RxuamF
1w2H5MtnekulfI/lt71rt645V9l9IigykpByUeOX7DnDE1huaKQp8Gg98muh+Gtn40O3meIXM855
va08+2szAbJe61mAAK0SwklEI6kQO8A3V8ltuU+V/uU3+RtA5ah9Tpyxw/w6LaVaIEJvLlTcQFjZ
zM57ilB9PXbQ+60Qj/jPQdpPiCL4TFbFPPLEjB7VUh51EERU68dsz8ifaczSVUA0izdSxqsx3wFh
B4qKb25VML9Io4qUdcxp7AhPtwcEW0kVV7bL6D02fP24wP3FW/mp81QMbXYYTXZMJao6RfWsmYfJ
a7m+v4KWM+0je9LSGwtir+Uoil8XebUALxeYa1lbBOZwSeaKMdn3ivno0tBiDlX3H/EW+le6AYs1
teyTqiimROanNbQSOt0evdEEAVIvO3WhUaHz4+dt9wgjJvDgqm1msH014OkdWav4l8k7p5zb2cG8
2N1p0/YKcGrO1y973cTyB0ASL4/dnh5oygHBCnOQBMW9h60HbQMhwTRecRtCWk4KZOqlbq6HaOPg
w5rxmfU/kojKWXqWP38LfifyWqTEByl5nflP/SEEn/+XLhezIZkcPpbQ8XprRiU1wlmSWULiuYAo
s8So8utVFX0FjfR1iBy4zUd/AsH6/KnZqGZO4E/rkPUj/UMlccMWQbt+MCFMu51+LDFqqZhg78DB
A/OFpPK3vXA0rZzEbm8+36o95qnt1rM/m/qxakovsSHbF0c09JoxCKZl8tGj1auTTImvWkXPPWuJ
hCuP4uEIaqbX+rFljf8I9byRdIuuJRReXO0itQvPzkwq4NfUvTYecXo0pUR8OmzTmaQTsYm0GIKG
zYpFE4bHG8TASLzNn4L2KyDohGsLFwN8On3PST/34R4eako637GkT7AsCAWLE8X068jqja9DhxSk
epkjtYe7KPtakR3BeLZ4nmx1TQGqCbjt8d4EeNGz5eqYaENLL67cLTl9rNFYzTPRAbEgsv4qAdjf
pJ0gPJwu07dOU0Y+CFJXS5k98mzXKmwO4rcsoSLHIttxuWO+1ieH/phdJf9ClDjsaKDCvVKI3o2K
dN8rturD1lmuSKUdUIEhJINTFn1EA9YW06H14ZQyq/Q+eBcpIbtHxhIu4cLTrPmvQi9sepKEIDXZ
m8OnunQ16myo8Gooh11D5uwB/4Cw5/utDiCS66dsFcIAhaqTfICA5YTkI8gAYNs3hj+hpKEF15mF
oky9dnGQuBOiC5Rd9WWjxau7bS0H60WxgT7ob4yZHP9BY32JbJ9OHkmiAklY5xN6/iDbPF5RgVBO
8VCOGgFLzAtSRv5LoQx/zRunO6cCjlT8PmgSGMp8/QTdmsTw2alUyXzwJ8OOqQ+E2IBKouJQ7rgi
xfNTkH8ckVIXVUEZrTXv5sVnda7hWUU6ioK5qxx0kxqBNO5+qOZc+bH/9OzRP8pdeT5KOcrwsF23
R+ibyB4U+Z3uUhjGlVHMr0ZqfCL3FnTIyUNvP3kcgyouDr4exQ+xT/SHbHBaNc3TLr3Fa3QB8Qcm
mnl3eQV5hOIsgIRPeXcCqhsZ/Hz0fqLPK36SZH7vO23iinf8DDAaVjgQQRfNSprhUovD8dq9Xy1V
qOsrQvHcjDYgI6J2aNImDPr2VhIoWMVHrgo6tDE+Z9FZHYVBpC9qVp8qsA+4lD6UpixYqUvXwQqf
5rGd9YxhJmnCqB/xCjy0W1FOBgioxnFGqxkkMX8+KtbizAGjeEBtA342XKw/zaIrOSV5H2t37P9c
uI7RL/Gi1Lu+1i1ZCmR2pCXgAYry1ekXALe9fn6/klml6vHjbffoN6enhlwFAjU3Y9+xRLK0RzR/
uVommNX53d7RsTTcf5pcBno85uUEkkUJxV4O2iQ0morI8IS0sMmPYY9YelS0YYyOT0rZVnkymhNH
T5kzfWDDD8/tG6ChWWQHbI5XZsFhqfq6bFEViFxJd7RHINtG+54HcXJYkGXDw3Q/vi1Im/ObwUIJ
PTyVSwTEPOYjGYxaXeG1ZFRJaSJjnzmZjgDw/PDeHRApYdyrLlfZowtkfGDcz8bT+5O5DQJ8P+1I
b5WLa4bQgnuDVZ2MfCruCr41OJGBgzoSs0J2OdLjKRgJ6qXtJlBhaDjbwlogyovsW0yHTfo/iIdP
sCRslh2OnghBiRikCEBMqIw2kpCJ112KVeJ1yA8CIV9DXT+Uz1jfjGcn0ZbUcYNNYhxMeFbAgX86
nTmRMbN7MQZ3Z/Of0q0MjzPLtV9isKqakoKYKgQwRl0GRi9YnAsW/2KEnuBSzEirMda8hUzH50TC
iUOSXSpBbpbRNFEbGOBRiyXCdIvx7p4RSNzIUBX9wpZlPjc+Xs0YF1rzgAfpuQdf5Ez0L3W1pWbL
ACPiUt4fljUDSoO86gun8JENVbCDB/SPycAfeuBlxXEMdruyDiZURgU20TzLtB+gVguIn/kXoQnD
KjbD0x+6GdZKFRjUizHygEWcTJQgmuAzJMPUZxsiTR0MB0ZB4vRpfKvGLyJOTyXJQKNhqcdW+ijA
VtoiqyMS9LPinkFL9AzTwBYV5FiwXLD/48bkHhvPZlrsi8J5bSAas8SJ/XoHccxXtEuNXBvE72+y
U9j36C2wIn57j1i6gbgBCz5tvv0FPQNbnd02alh4k+BVZ1w/m9R495Fj2EO/8lAxUEcyTXm0oMVd
q8pgLlgWWGEnDZNFRbD2dFxDrY/n7FvJEJM6czyUWrHUYk/kFuiHS/6X9Wvr1P6m2f+wHO8yNOAR
Uw/v4KqBfmlebPoJVehBlsglyMSjtzmKNopPV+/PNrrZHzYDZXZK743eAIguaADgCTn47stI6h3k
BFF0BrnOEuDHvGximSj8lJ3P6sstBqeKMrJdBYPGfA5BqR+szxPx80yox3sJE2aHbpsxLhe/zPB0
wrPoHVW5nVrN/hYy+f2ZyofWQ8W4P2kupNCUTehFuXcyXn62K2ekFkxc7nldtsLo2WGUg/ZjFuJd
zlZQ08t3U3BeIuVZuJA1/1s6Zrbu8ftQxbrrO7TA37Dix10UJhZES1NOS8uo1cJtW3MB7EqnvJlE
7DFWK3ota/TOFcRs10gt/JusYa/8FV0SRYEO9yRm0VCKdzo8eVKjIyZ1fknAoBbgyVTt6WW1lr6r
alikhbxN8+HWwu1UcMwX2vyig16j7h8LGF6OBY1TYyk1YrXnEEYkkyho82SXGfBKyIxLyJ6qDJ49
PZQ8/zE50wwrEQNkMKOAIilIEER+4cqFOnsa0pLoZ/4dhVjsMuMlCkb+kWKTVabcan3cLb7oGegv
F6LbjsfWdhh/XVK8hi9boVx1WNmHL9wLsDeAl8aGn+8spUbEmN1b6WPaGY3Y+U1p9kQ5Hie5Zeur
aHawK+0d7s+4Ksmzr5Asqj7K7PeYbLoHNp0DcLjeuU+d9Vg5w3KlXL+hIH2IS4z6oaZQAP1RQoB3
nb9L1QO3EZTevN4T3G6uP2MUA2zU3q/YbzEO0IyMUgpe0x9+qu/8J2tMg6E7wmSW9+gQ3rDancSA
EZ+oRD9lVC8XnaMSmxwOinswcCWwpo/Y5xne6ZIs3S/rQKvm87U3zmhPxxCgsoHKWp50xlL1/QyC
vXlQDwjr2wg5C49jHva1isYN72unTrCTVE2L2if70qC71iVSqSXW3z0uXvRNgLfHX6AJdxzJ2jmo
LeaBNysAM7hG1bVTTC66h0X3MiHkondDR6EyWK2K+nwOF9Vmbq9gfbM3G7sSQiLykxF9kTiszW08
Msm4UEy0oL5guKI/SMkSOayU+KA7B3dwT9f7AWHNV15N8+p+MbjmQB1wsP7Awfg4UnsEnyqobOKb
aS/SFsYV2oluZ28M0Wway2ni/j9SHjEAWXCA8r271YpB+S5HHPKXBA72X1sgbbN/FvdwKkBvb0g0
J5S2zGf8Z4h1VypOGVbFy4Tk5DrM5wU8m+CbXdJiTR1SS+6hk9EU/BczJdFXQRgBSR77lhk58qYp
O4GxEaLUTQ1mlGKbcu51CkXSQF5gtoZIDtFN+nfs95TGhcehND+DD63sot9hSFnl6igYxQoB0HO7
+eg4+swuCVsOOwZgg0YGKnJRZFZPCSsALwb0BnLHn0qWudWn8QMZI38iPA6p5115B5Hr2X5gT2uT
2DYPJka5Oj6bTTmmIMfE1nqooGL/sBG6y7xKdRN49sdDxLWtxdc2LMqpas/3g3lyh+/KwYEAfUi+
CJGH3bO99Y7XTAZbJ6/2QitAw1jdnnwDZyG10vuQ/1PXYQmaMsIjtmw1/3qMPZwDyXFGugqTvSER
BBcSMqVY0M6dzd+Fky7R6ADTHJxHfIAgrfcy1FrxF+dRrScCRQL38bhCLVLVHQgCJpBeKk1ajBqo
3VBQtj8P/PR7SbNVOyPYHbN+g94JFdX9jGhNf3+1odvAH8DwqD1FrLWhFuVgcmTXhE6L4BKDb1LH
hkzgVhKz3Epv6TPaSnAkUqZVIzZLCBtC03p2H8iqpJhCgXIkhObOAj6+QqljMXqM6lhMJ7L31cMr
1uP0O0IhAWt4beAAZiMP7dTC5DyjBX9GYa2nqYFgCKCCm+wuLZrYNeAGpQ2192Gemr1K2h9KvW6m
tjReh8TIFt8oiCLhO/tox+YACRPL4IMkWw5GbkLudgp8YphqXqq4pv8awwl6iuXHs3WD6N3BzRTc
VLNqnb+9sL2msIYJHanM1kooUX2ddz1vy9SWbBR/VE3dpBBW4Hwe8htnqr9qLJ4cxT9401bSDcju
AmgqOqumgpLOt785C+6wEgoC4uKmDrbjyzsRIJdEA/9N3kNewJUmNrU9KZBToNvWnQNjnMTk5p6b
p4xBDl7Iqh6gaVvoMf+iHC1ExUvDBDTbswrQJeqpvzp9EbhH63AY17qEUgmbMZTHKiM+a1PHh8qP
/JrXYCPF+yLBcN0QTOQOmArjpL5coXnD0jL9/qRYV1abqMvkt6sX5KJQ85uhCvJD8XKWlJrtGspJ
b6cv+WbW22VMiJs7PG/y8Ov7BJseptUVD1zggOvQbqEMLEqs4ZTOYxL+jX56UrNo1yKOSGe1Nud5
QdK6Z5eCpXsmgboz0AfEP4eh3BqwaGMrfHI1NLhcvTn0otXialYvsK3Xufft8q91YOULGSBG6HAz
OVfYQ8d/ev+59o0d9tdvsVqbTXlmHK0gpOIMHDoBpLbBmnf2l3N8WmHwO3E09Mjb57QixLNVTzvv
SDMBvI8AZe7noX7tMPSacWSyLfEKiHZuMV5SmXgWr5hAtSaT52TP9nfK3/S/sQkYhBYa1Ijz1pMj
qOKsTXNkvIdPQJ5kU7mt5+0xz0rIUP/2MAbT0VYW0y7a2tjuitsVfilBOCsy/vqChARp8IzXQQ0U
scOlvrFk5DPRKeiwltgqD0ttquf1DQYFbumewp5KdNXWjqu+gATnL4Nspb9TGJCF19zCm2Xw6LaB
0lE1LTENrcGMOyaM5R1jBzKaDptUUyy0oFrc+seIzLJ2wD4fi0MgUn7ghJhRSpUTcrIJWswrfQxs
af1Yu106tcsKORigdU99DR9sRR0xv3xJu24DEqsnuAat4dCOZ9arsUOZf/DkWvx44357VkqN0nhC
XnCdyMwFn2p+sPHNVKVZGK5g3G3mJogs629ZNKXRfZnis8xYk+FzEuyZoZUh3I6SyuycxILojjvL
ZBNUrF6i16T0ObJGh/bQKWc6R55TRl0Se3Hl+6ClFFJQ/Hwpd5hl0n9KtB0C3O9D+TtCgxLkVFUy
7EQJTsfo66Wb0kOsoRQGtsLMg7QLFKH6HiwairVIMxVEkCZFuJcpOPzZoEsZEneuehHUD1wuZGwm
NK2ix8fGpWMeOdF6tp4s98P7xCPN67q2fHH0SOhcnW5NEIQIxF496FJwAHzpXGWtlCsMAo33R1q6
KhfrKkz2j3m1LS4rJ8255LE40Rwc9jUyrHX+/XHGp0/Tzj1GBZvYUoIFws17+AxI6Ew5fxKE2Lmz
pnozM5OaLiXSC4pDvyrMQPoKdLKsaqYgFxgBdZybRCy0IiByXtJCMsOgrNDAeF0SLLBxxjX8wEU6
7+00iWscxJt1/ujrwV/Jm1/C45r3oM4LWvqaI9iZQxmKYkMS0jecjE45EzZdePzORWdNybgztj0Y
myGC6W+75z/OsFJmEZ6lyU58N/x88Dviq7akXXDBHoiu2UocL0+vx1gc+KsVyNoJVVXtsaJIR3iu
09ZVz2Ht281OEN2kzL2t2irRK09rWzNABz68ECEMknHMF4ABfDqO1YzwZBYuTQmiP0uDvFErnqGv
GlYn/izIV+rvtKljpuXUwedmwEE/0B6w8VzzKdWbItOfteQQ6txEE564dPpneJZ9X/28GxvshBMV
XyVGbgSKIdUyCyj2w5DNW+Q3Lv0lb922zCYGDsJ/oex8S80WajMucJTAc3eTBDgOSLz2dsxC1J5A
yVohTr6EV4wTRHPIJE8shsOwATfSiFbNRV+ruTPveIb4FgwIw+TPDyCILRDt4YVW4E4bWVehKTVR
/bEqTnuWvwnrNkd4tIMFM9DfjDUe/WCEnYi6ou2dBuyc/8fW/q/agfE8vQNaq/XS/mpArU5LVRoV
agjtpfEDTqrMRMUOK7D5sW5JXPDhiUk11zK09ORQVUtgv+M3Zzmcj8esp1uQ5N/b6QhoA59RSxLU
rqZNhsbT2vSgvam7NuzuCLkEt6XODQ0TwC4GBibSGoLw/qGp1T+pKo5cw6erwFIC0MwQBozkcq7R
BM1AAf1BbRAJhiodcX3R2vRC7sM8oOxwU0v7k4/t5H5+dnTxOBysUfVhgfA/RXBemo5QMHGBGdBL
giNI9D9m//csZMm0MJskEQR+SAUipEkJndTkXUdl7X2mCPciwW7JDy70tplGDTlvryjcTliQ8BZg
yhQQazWBqNmyYYf6Djn7dCBIaP1vkRoGl1Y1mkdnb4zD8Tnt5x+2wUCjIUOosZiI8PY+8SK3Qe0u
xyqxFd6O+pp3K9eVAWnz7K/gQO2zscqeUsOh1/tKAzWIUI9u/3Pmq8zkoUJhi+kYoykK81EtJJTL
nbREBr9zPVYlYwINWyvbLLVcbXJj6JluGk9X7dV/h9W6IP2BE7FW/HHs6qAANXadunB8V/rzBiow
rvwxDc3YlQjf44PO8UmWI7QX7Fryncs4mbZTDAP749+lGyTXrDnuZS4KJxnkADfqRowaU9mfLVpF
tZpCdm2bhiDDyQlEm8rnUbEn8vxHrSh+vEM1EruERqloZ7094/7ZVnZygLqwSMnczioxv3CYns0T
p2jNPr+W2jgdtgRNrniFTJdrp3BcBRb4j1kEI2Knkcir5xNReJjhEszBA0AY4TzTj7V4qliwSsec
grioz8jbXTVtj9r/jDnXL31i7dXTAGd793KJxNyrxHbL4j9PNWremOaXfVDN+CmI54/k2+kLPMQo
3IS9SVz7BLz78hMPBpPx13YOpvREbmPkv8bHlngdc/Ux3qwaYLdtH6DfEnrD2xocZwYotUGUvOcU
9tU/vPWD9Z7L1Tt8c1aAGoVhi0wvovSecvaYOOv75C6ExqXt00OPqwtiCMsRSTP27gHS4X0ejg4y
4PXT825BsigqJrHsA8lhzQKO/d/+GrjU9vKtJ/1NuP7I2En5W1IBeuwoc9qpbko3z9c/lFHroTGy
Btgfb4fzNgBD/31N7KcMbG+fHUHiV6f8Y1SC3tjXwbMo3OP2s10rDq8r+ahbGNHXWkhPqnDC/Me8
0Zeu+ni3RMg6GTlBEs+HszD+Cdr2ietyuPDQCLxSFDuXAYZ+41k5ZGSW5d9xpFxPZOXdc3+Xh3Am
2Zrcx0mG9sCmeXWva5jT2gtoRl38ZHt6TakTaCN6d5CXP5Xs+w4m6DRpbUVTAc3bn035O8S2Kpr6
p0bXpGztTkx7C9ThKPmraO0lC1TgEzzaIYvGogl5ImINPBgV+VkPBXi03prDhAu7ZbBu7o+qN5v+
i0TJrwUyEGuOJC8xh6b0L20dNdaGkHPUOTZpxAj4Ybg0OztpbxAhifv9MwOQ3ueyDJ7+7R7jK/aO
110PpwL0DKTAvp0a0O/dEVdFvENT6Y6pqM0pCKV4FE9ZN3ViCbdNQNa5njvQKOUGOJAMbJ8ZMktT
uyQ0ZQ4DDge7Ve0/BwWB9ZlWyHQle6L4+L/uFnDYnHPCNu4BDBrEQJ1v2jwbQG5O47GCdkGNJq/q
6yK8kcVhqiDesre3C4YdgGhR5XY6e+C+y6/A+o/QxTIFqFc5yvU2XuRVuWibNPgnJrc+Guga4wQ2
wtQSR3H0hVC74rco3nHHzPtC9cCQyR9o5Z6I/obG9OLv5LUbA4jwS6hw9I9Wy/xSbSdmkVBn0csl
yHDPWycstIUIhC5+fh60akKSUkMU80W66bKm177zy21BwpU0j9JTmqRZCyCWGoaA63Zq/fT7KIjL
ecpZon6FOIb2hpk/HAgPaXZhZtw33PWCOd/HxwNttCTkylMCSnMlYCQ4BIxi41Kzwfu1QGUI1EVS
lTx6EP9i8gf2zc1sVX1Aj3+AOKayGUI+M8LEt4jlvevIbOvVKbm4Byo6V9pheRVjAHdvsne37rbc
9Top4lacU+LFJJTBnyLXY0v/EH2LS1RMqOhgKxyQLNPGes6L2FsBA2wumKqiTJZknG26npp9SIG/
vAy7Z0GcewBiXZ5LFZ2A5CN+M0xihbS8QBrvv1Q/TETKouqIJ1QALq6k+By9m9Xn7+PU4t+1eMn6
yMv2MNHW0eQcXdg1a8sY61onDxG7SLebIjr05A54lEPeVFaip/Dz+xgry/qfdlHT0I/mbRyXTXde
Fnq/3UgW+UeMw9Nts14fCcHjQSIBh51t+Rwt62LJmHndm0F0rjoieIWHp9CEP4bBwZlDrXx7DdoE
c1JiOUW0E2AZgn/s/lBArQP2SHAc8xOw58yZPfldiCNAxQEFdE4mwP8QWXY3nH7Fsa5sD/IxYlmh
1zu2rzCwkwzM2H538m4bqyRKvwr4cWBPZlzMpHomHv6rf1zby6x1FBYzvam0vSIZLM2ABPOQJ4fy
x79Uwqo1ZTrFPwFmvfanX6pO3TngfAp/YjB3SQ08q7e7OPZ+X/DBiruED2ntLrPU7xk/yMz8OcBJ
hEuT9Esr2J34ZEmpfz4bQ+GN5c9TRQTDcEsLrMCvp/GrOyc8tz8hno4C7mpkRAaxQcqclwDpKVRK
l+sgSRxyoyQBdaKOx2FU70J3fjsi8oLks7U3Q3+xzNgR2AA9ogPPXw7DMVDiMSb1eFyrZFFpxLig
r0rCz4vueIb9rk7QioFCfCnqbYRLEl3rrx9xTWFUyUG7P/ocszIn8FQO7wdqsDzzjxETnBXIteFE
rskweDUQ1e8j3bBr5LNphNjT+s+CW845KEgmsElPkMdUHol/INCpZSx+B4K6YowhHQkwHE98fgwO
aYcPl+7A6H+YKWqJYuCYidiwfbxsJm4VNZEEuPdN1n73l3dOIGtXsfLNtmK32cPVcq6AIiAHTU0J
21dwiciCtE6AtJENNdeNwqNNENRA7/BJ0wPQgffGkrCDiC/uV2zXogFreOiOyewy50vABnAuzRgG
qEp4OoI5wYfP5h1CXlt2f4r+Rm7/tc+yuCS5TMGUTdMtDgo0oUMEXz6N83onmCmtZSjfi+JOfC0S
WudTEWMai7HIrDCaaBU2b5YqF136U4p8nFR5AsUZquQHzIsJUpsOMfAtuD7t/FQX7+cG7RPnwtc8
slqBsSk8qqelCuPOz1TmafnOY91abAeMpjXjdAFzr0WIAq7nO4XLa4aX/k5gtr4YiQAiX7O3buP/
Wexw5TamwaOmSB5NBfSvdLbaPIzO/QqkH+ey2ZryklzS5QafBiKNamx/wi/dM5/szHF6J5IRVcOB
GZszYKeJ3ejgXVfx3AAukweZLQdsVIM3szekl2z1N6VYxqUudPyKdG8QWM28ZJ22+eF6Y9bLqT+j
oziOJcD53sY1dsyb+2PKvmKGmmBhncITkWompQ9ebG805sti0rF4VW8ELRGCpUGZrX2LRac4bWg7
SuizqEXw7q/McBAMme6Xz3/seCYU3+IKCe0d1w7UccOPDjGT28g35xMRvnk6rx8Kl6BTcoLF4zTk
JyB/8ZWg89F4mIYpjHAQVSQjouc3rE0jM0/xTulq4YCrlR1UYg5Pja7zgnm9zSCkGkwR2+fgXwo2
hZJp0fvrFsg2I4z7VxfSkx7WAb3fYmSbSABL7YF3jZfhH72+sCunpTsFk6+mOcMJSbl8TI8iuUAj
6NR5oQcn+fD88yH+XoCaf901toUITqCJwkZqww32IZ3zVtsk/r2XzD+3IAhz6cIlKCAFWqdBL1oQ
ZIOIKZdsHZ+IDnJO3XWIN4uFwP5YOt85PwjdK9GokR1lF6B4EQO0EF29CbhH4nNQJ4BNeTf0HRvT
ppg0A6PQT6saUTJch/D+IVvXQxFzNCe+ZOdSEN/zJi2JXy4/35ZesjPA/yBjxrHSMZWXzdoAa53f
yxDpXY296xc5W2tKN92AC0aXC0SXYy8QPrQq2+euwBn7AsQ0oKbjiKFDEmFsj5VdQEuJgxiD93QD
gXNu367sByjGCbiWZe3htFF/J1SegsHkqJI5KIaCcFcxr76s3AKnuz4KJ9W4q807b7GvHkP3aiwt
Y4u2g7LTpLn5TU+9CtT9D+F3whGzXkAdOF/p/+QQG47Kl1Wyw5eF29yPj7xL3yaeDDwI1rq4SoRh
jNG5y72HX/B7Q7u0z+LdQNQkT2IkDiZ9DwBS3O18PFWteZSGDH3cWXi1ul+fcjXEKu08XCn58EX4
C0z/qJET02i6fq2ywN9vIYnQ61d2/3eQrTApuNmcukASVvn1bqJi6kWd2QjlE7VUYdCmYBNiZLtS
yTVQKNggGzaGXYs/9xNKKbHP77sfbn5q4TMbTaAzcxMnguMdb7BBQ6uaYsbF+T0L03EOlqbVIRN8
kMicaIuXHRddureSiV/WmISC4uVueCruHJVm2G5DohKssz0pm5CWsLvm8PSahrKJMVOu3yZR5I/i
gEbbdicQE3kU2Gq3Ao0Vfz0zYSMMz4YY/bbFeYNcUW+jj9m70DXe4RvD+qVSbf5Cd0P2aQ2v8Acf
UJJSPyB26qCXN22Xd4zKGl6TwyTqhTUcaE81AoLwNKpo+GPw9K2BGybg98WucdTeE5smsMlYRRjz
SxL4ZiPK3M9unPTTJuifacMSxymIsfCidFFAE7BibEk46kt7i0rFVfLNrfTXnCFvAs53FR290uur
5D83bhmGJO68Qq4kpIYrGW7xHJ8c3BgXlkoEtelyC4/AXp76fVydg99D5yVPoxNiZC53kfuIfbU4
vYMuxV8oLOx+OQUbCSSz0EeBfy2krK0na84DJojfFBB2Jp0VN14JELbuPkHWf5AP2sNDDuEjhUhQ
24HA/g0cHv9pXz7Sl5A8ZRZsbbtCn3L3ontSCbQcaioqzX2hGUrXeimcxj//TtCSvBxW6/OA79NP
cn/ZnMn4/QLnSG70LWewvR/1Ro/q34/a8rC8j5vBrK/9QwU9qkDAto0mn2/yTIDaYkWenNlE1Uce
Y912qoY3YttARdBcjfXtdAlmcEf5JMqz0TPL7BAxyaCJZ+mY+ZrCOTWCfXtH/tH8mfB2gp+62Tds
wy9wJMzmmRIZbadfCwZUiNUv6ioRqu2Dfw+bHnkGn8UJQU4m6ipaDBOD7yBQQpeQiUZ7krXKdrMt
yIEz2YHKnxXK36+yov7dktK6NWItFqQ3SwllMfGYXHl6AKvaw2jh0pXA23Ormejr5Ei8MmYVbA4R
oyqGBtjSarmHIFvTfDmgfhR9OzaX11LzZGc/N3Gw3wfANgyKQvskLyBBajwa2pR7OPhsvJdgT1l4
fmlxvMwOgitiGx/vJM3NvDtPTa5OlN4Gg2fM/0IpB5jbu/qTm1ftBtNtbxvy4oZUMnjIA6B6gdor
nMBnjjvhrYynhhDt4YCxhy+sI7KIpg4PtmnzFZqaZyElTzx13WXOOP7s7Rucp4t5dVRdLEV8rpqy
ND99SOxEGEQp2HG5g2rTPa+qeboonRoWpCsPXMqrPKszvkHOa2Zoy3gh1i503Ej/d2KyWTyINqCa
cPWgsR4Zr830bbGokb2cKMuVJIvWCYuNtwXTcjx1Lm21MxWoo4v8lzw44FlRbhZtryGILklS/4GI
7wQDr9GYr3fFxZNg7DhjQVzGNy6ZqGkY6YyTvoie//wy019JYx2pEYSBdmuOlRPr9rL2JyvwJaI7
niPN7ANevxWTSV/zz8t8ybzetQ0wnkogYOuIowXJWNhiYSKB7h6iTHF23vPKNCHPelBuwYdY50mf
DgC3UkeWLTo4YxXAvxBweZG/bYhfUp0QypVpFzCO7RVtxNyg8Xy9cKIlrWDUky3xL/l0Cjv3bEce
2NbZGmcQ3qNE1p7lKCTjXzX5X2i4WPeclkUBH/yxJ8mOGsEXDb6D4C1P9/CpX3/0yc2hmzKp4Zm0
p5g8Yrd9IhOcSS/136Y/uU1jk4q2wvKSA1SHTuEiUP0PWG3MNQ3C9L+8B8jrDjXArnMw011TXpAv
hrGWMtYIPn2eJig9NpAkK7lmJht08oQNrFwV2POfQCvlLqOBoHncb66mceZaI5E/E3rfIoJdvw8J
ZLfyJzoo+ZWGLxBfZruV4ABTmYxJYFqJ5jZ3CS8u0cM0fBbCmpQvwB9Ezxru5AAvtjS5NjOQMFcp
Nvh9yiuFbsLdNNBIabk4VSNYDmPO7XdeDMgB1S7qR1W6mqaf5Lw8oMASNsUxH+bE4qhcK38wGke8
CZtc2XansI5vA0ykitR/SBUik9XtjKaIgeDNk0LN8Gf/N8JbHGgLWm32zH1YlSeizSTuy3RtOIBO
479P0ATViymcKHc7IX5uPI1li4BLzogSkS0YakF1ji23L14qIplxNUY1Zl6CVJkr52zToaniwe9D
0tKYqkCjTwEMfBdPaJnr8VfRzVzK2lzrNzYu8I6f0oarm8J22PJHnf0S3uQCYJsAVry8iaCjMSE0
zfCv1K+VVUEEtkFuH7a50u0hKgQWPHYWK+iyxRL4UAw52G0pq0lo7HqxMjCKxfwxJjhEWTYi0ht6
7/A+mfLytY3ClmFmIWHaG2ANZol4T8qRG7vglT5ViWk71N0W90f1ieLgnDhYPBM5HZQY4uqYAFRO
0wkfMfNaD1Eo8J2EV9oJ1LJZ3r+x+HTpbWESVEcV7WFgQDMjcdJ7sqeXsKk1KyUjrWcFUJtVut9a
BrfDbdRlqCIfME3LFOphVd9lSYJDJlMbBAQ65/G5cbNI+97OqAoHS32W0YX6ar+mNF4m60whNaxu
+OXWbZ2R783TTOruUBRYm1Fyz3MM13aqQxPHW3ObXfudAhl7HPbhuNXbcuSDHRbcLZxNslsj7RMb
Ss1ZiEBShrkzKNACYo1eSQ/XQArMH7hzcBAE6WhEWoGwFYx+Bw06lj40hbTeff3vc8aqlRcjw3vL
LywzPavwSiWz8PKZ1rRTPdBAEZsx+XSIVlhlRYdW67SkP+LXFB02ylKfpH/999Xj1yiY/rBaIwJj
qlp5SvFUyQSCZMh938JC/Df9DIGIyiezZxBk1rLFpYSlBBASetsHFRFOdssExFDCtyRqe0WzLWfu
gjuUBYcmp0ecQtcyf1banmDJtxI2hpw2SdqE+j/607LXtowtYjX7l7WYVODN40+pAA96AIUGUZub
0/TYEyaYysZP+3ZeybHK4z3hOCVfnqHfiFaZWO+NLkPxJ8XVedydvTtTUPBKg0IPBrQKYN0FipIG
8E5kvBHMNpHuZSvr8krq89D++LsbaZSIpHOsaBsTxm2XVYorNHf+bmD3ccLRk8GmT09++Jt4WEcl
G0uBXzWvTI35gjw1icWPzF24rSL9+vMqOBOP+s8OeX9qG+tRAsotGiTg6Y/cS0b1cFAiBYUi+g+0
ubuCj5/WwyphmP3ap8O62eNjdAjct8FW5/nc8lNWO00OLVzYsRHJ9UFkxDkPJYxwC3AKoZE7VNyV
0nYcKo9iMH9P6Ir115clHkWFxgh0ZDVxiaGe8t7R3Ls+PzW0RD9B6TXDm41F19dJAeiWlVJI7p0e
Zu57p81/uOm+i8xm5MJtv7V1DeQMTPfh2xs5J6bAqISixttdKd/9//ho958W4O6Y7iIp9jOGVOEG
HtRje1+6Lt5SrwVfHgsMnZsu6dS1+NqCKRc/7sFTPu8/gYemMyD9lHapr3mewMWYFq6WwW597CXJ
c41ilhejoM5uNFO8Kx/WZlLPAKfdGvVceBSSByBDL4n1txy1BgWa5xk1se4npMcNgINmLFxt3U62
Y9AFduP6aI8lkCo3z++MDy2R6IQEmECmvT4nNIuzcYGGnmAIQAYPiCwM2zMOYfpJdF7MTvrRyW1p
d1z4jE9Rhf2hCVMyqzgh3ApR7W5jmOTU1WHm1v0tS9P6t+TqEJcDm2c60dQ+IbSmxhrcEO3cmLLn
LbipEgtl/9YR8WU8UksLpRdpHuKRxy9RLUmGLFFInjatQHe7O5VGncmXHHD/shVefKLH8NaS3JLr
DvKrJjFRjiLpXQNbpth3tITxbAkzSfQoMOtB95YtMxsQOj6xkhPRaom11QOE0ryjHORBAN7VOlgY
7RCtThtl2dBClu470UQBt70fwA6bDm2XEP4T6li9N1NcNN7gMHEhrLIfwNBqCC4bVJcUQ/14O5Po
4S2hj+7BUJiA94SYPHzQDBU4eLkyVhwQRWx+XAtR0j3kHylBDBQBGejK+enwu3dGzehRMO7scSux
2t9Z638iuxj5VOvaQfDDfx2Yi01U9ZgfO5V0bqsQnb2sV/QUX9fsI5c16rfRCPZ7nqygqk/hbsOe
v/uXbbUAp5ixtg7yXP9oZVUIbRMdFPzaN67qJ80eCeVWdX6qoaIAGc9uWluUh9rUkqkrHdqjPka4
0Ue/OfZ2J5CT+nij2+dcJWZAOBxFe183H4T95nIJNvGYgB/wwnycfUiPPbMVeGg0fyrH6RoFiOM/
OrPGEKgFC/14GgCrp1HTGO6VsFTzrr4CYMCbpwFrU3VvKfd1diLlYQ502hDbPQcxWlpIxtyMGBrd
DCOQUfhIYkpZfioTWurDf7Ssk2mB0w7RTjamzzgQ8Dq1eDPt3QSfdrUz9I74vnV/6gFegA/OVwpo
7+Zhk/K2wAbH1rlEO8PWERSIYu8QT5C+zpnR3cTE/YYhKgHmPVq7ISgUPR1E9FGg0GZZ+wwjnqYB
/hx5eXqrtg6CLA2jRiaEv/iUcUmrKpOlk6eZXFvq7URjxYq2W33ZluymOzbfQvnwivwoL/wy5RBc
AxkUgHAhODwh/NhPGnmKr+0yy3zSTWqISm0Uc1hT/UdK/RfW3QLu3I0chxz04OZJAPoMo3A9JwN5
Cold2TU7y6kAhHIuB80alw3pM5k0IthDCRqzfkjk4SaVr4sOUVtkeRLZ7x030A18+XznH1GDI+0M
bw7l5IZDZPgvoJvkjmdy0+MW9cASdu/xWhPirb1Sh7x90lpAMGvDMtsmIaU6Q/VuZnxZyycxx16A
fdLB2QZSl1JS+eKaajMz0k3yHytYYlmTj/t7r3aUKNZQD9/Z2SVQMh/iHjvu0o3oDD/J2XtzUhDy
mgIUwx9+l4fL2otri3+sw9gZTpBrZ7U8qdPk/zZSFRer9l8IqrGIwK9brhbZgyTN68uxoLryoltr
YZ8VAR2wWofSomrK8dj6kOsW2wI2p4QbWNT2zqwRNYsZZsa883360iRTJCFXM9ukCtqv82Vv9iLa
3LIulla8wxnoO1V65p9kq70yxvqpyJzdun1wIkYs/GqUyN1L59wO2qYFy79130aslKSqtSxQT/lI
S+oa0r/oIeaHqa0NSLk2eSh1gNViFEqtNgEIkm00NzH6ER2/a1ELIJN0ZLR5ebzC4Bq5U0vjPjNv
usFj535WKoxCG1ZihiVLNQOoy3UqDuoHbihBGhTAnGM2et6KnJ/yiAOyIlIda7s3mtc67/hepYLs
ZVWAbtxYGeNODDzvEDqkho2d12HZadE9fiYxJNBWLgOMnjNh31Wo/i0TGGVhkugHfvooM3fue6zI
p3OVsogYrwqEq+hYPliBXzFxgrdusEVPAj7VAASu6eiGTM+YJbDrw+jvuL9DRsdFD+oBvGHscPYM
REJKZg7anldaszn4gqionW+bAC9HL3//Y9drawTn1g/wiOlCqc3pR5fS8b+jaPeg2MZtlNUmPSl7
r+ZHgSHcvm7s72wc3yJR78ycZ5CVeNWKRM4EzQG8SHnADfxfxQKnsxwPmWzVHFhGlxO0K17sOhEW
WX0OkbyoJPkdLzjemj+y/eYMgpWOA5XLWKpO0TdyTgmSzqc8Y/aJZ8CLmfgpgHYX1RIEd9zlZ4jw
yrHPDHoKFiX4cn8xp2qk3zaVYfJLfFrIAnQTvptCQYSRrUxnduBm3O900rXVGEJTAzzypHkFXUcS
tuRKnEIVt95ZidoW3N00A5z8mnSFHGpbxkbZFlUFnLu9od8KKVUaLBqcgPdsT8U2wBi6YJRxkF1k
CG3l71r9BmvGpKV57kWX8LgErxOsd2oxW61YNw6vuzTh5J0FM9TqwRwaZQqjyZPYnbV9H6dP2jwg
/L80tAlBc3xBJgHaePjv+ACKWkKOkuhyMq6NNnU+nbGtSsqKcyjr+m1YUKeVbnYRh+eW68J/j2Jc
uqPbD33KlNdamdoZYRymzq7rw9B8SCXioG4co8fUGKTbv66cvZqV8ppFskR042y/Dc23ZNRJ/eDV
UdT8UhJyDhgVG9FwBJeN4H0OPmfc24Kzgg5ejj2McV5LafMsj9eSLHb/YWb4jQpjPKV7YsV/m+6c
QNkiHvCrsfx9pDbgYfE07bxY24fX+yAJ/GzMyCjc7TtC+o9sGI5i5SkUesiPfWUZew4bcKWubzzn
sG9x8QHlYEUKOtMQVIjq1uGhcB68zM0Oizbh02BES5JgX81KlwEy2ndBsMo6Jmf4KxkwD2HM/pYJ
udC2LID/cB8geJwq9+ZibEU6/jK4x2T5ksOanBKRcLRZVfRIeYN5E3WiON2gJCD+pXLzvWW5HzeB
tyfmjOMlWwaFfUgcV9LbwPbLNQkSQTvobGk/t93fYUXalcgqlUJVirsw/v/DCaRI1M/LtukRtWUN
4rpzzYO4tZQZo5utLTKEuI7sDLncLbfwVoPDxvjyQkdulzTWm7xhxefJ6wmRoHuytO9Ef8W3kCsq
5dhej1TQeSp6nfR9QbyuaPtzAOEiHyBvAyGapInwsOjr4uE29fBY7K9ZV74bvoK83kuWndV6j/V8
q+ynBhzRgZKyyMgXmKLvV/D1zgciq13uKuu1zWH5OXcyKzpR8Bg5J72T5FYYZMkGKKAMFgE1PqBe
mC7YYMHgoYRVgIs+JDqnF6EhoAEi5YMAm9VftxMdlb34lJ6PCG53wlgC97ztUPq5ogOWJJ/xYiOv
JhQxF6rJztwVX6j/Lhq9q5PZsB945HVahFzU+cYAwjRaDG87bBI0c+1DLw7Vixn0yNMAC/0Gi5DL
lYMLQPzSfwwm6W2hQjDTpHEAijg2krRbe2kYwSiaplhYPze9BwmrJVGKtH1s+BSHdAfFKJzrvoeP
Plvorje3RjphX54w7vreDvO7PLNLRCc4IqDsYIZ3ueFBrHAxkS3FiSaqcQUe4lS2MPTVnyAdo9PB
B5H73O726lXzeVcAQiCoprzjKfpI/xLv/wac5VmiGFoOCeywv7IQGfLrMkKfr/h1N9uSWWKxNhXj
JGIOhh/G2uuzT+R6C8U8uCAf1eGrPbLIQAD6hZETnHcGpkZGR4u88oAnyi3CYWzaL2/VCfZvekrN
tNO3GVO3DS91y96hVCFfzmR7jvVpbLdFEta7rgq9G59racWkNBjxLDG0I4KEftmEkPc9f9ZjXDbQ
R+H/qhERejZwBH8IDbnpfING41myZ4A7hQyeeQ23PpuQUzl7ra6XFOWjcBz4bqZnNpnG1W/7CtU3
/cxGwQj8rZpMivYzvrhpxUltL599udcwE9hN5YTyLTqt3h82oSfYzlGQ8WTeOn+sG55JGHqdJTmT
4+wfFHVakDaU5b/EuYV+n62m9v8LkMBhNZr769Uys8UoRZkLMfAICxzOFY289W2Z2e+9J0T9iTmY
wRb5mqpFcHhqjjqMkSwTyqC6MbCbCTfPclacdKNeXgy3bj3YibEGPcNInJTWPGRinOeHcf27mcOu
kgjh9NWXxZfwU5OUwMtYdkrZs6k/cGN9AJJebrR3dI4kYMlMiA5RD0tiICvVkCmwTUHhQVaMHMwp
6F4bU2ljL34sNTuEoUR3nmhiLt+yNBFZn6EBEte1dcn+cKJfAI1Z9pfG4fLHKEZs2E1JLc3LaHvB
hf7rR2VTneeTF5JOLe6D6MBgdfesko1KImdlfyoKULB4/KJR3jq2fS5pfbnzLXGrN3bybZXi3it2
iOjnepcjxsk7fyYa+3h+6HpkbjlkmtWs76wkJt2DrPwe2IZUTzyYWTivwYp9gbEyr5EeKGa3xAea
ICeqrYoCXc/V/vghvfGvGedAlYz+wsc6nXLfWIg6IQNQ6lqL/L6s+hnWEu0T0kyt9+fq+nUmIJRu
qPBxp6MzKTKeCpnxyFNQihow1sWm+x+XFsjQEkoTOA/eiWgwDIBQw3VWdOMJ733KiQmiQs+mbAwu
ibmANo7MkZRGgJnazg/5igXnIlSthvWiA+0SXR/VtaP+0OmGCEm5EdSkg6VFnPgp6vHsxBYnnic/
9PGfiPyRsCZM1rj8a7vXZe0khYmr/aRKL6ynsDYD624LeWQxNWcYicE2HtRZKNDGpuZQLgwt4nWi
Z78tEx9f4Nl6qP4UOW28zWXaI+v4UlDceXWSEIzbDqHrNxUhpIv/1usWVqtHyvPzid2T6feI7U0O
zYR39zkTCsOk2VQyYu/AhVGLoYH3w2eiZz5h32GyekC1SJU5Huff6TloeOJSSTVTjzXFIIMfGQQ6
Ih61XzKD970cvXQ4C19y+5Pl4BjwUEbUxkJtk5zA4/WZsesI/l21V47CS0eHjsQi1pfsqev1tyye
u631IdP0hvPCGQBEOx3xPyAORK0u8eSioScq6WxUeBPC/jn7JQvRawmfPZO8h7Lg6fKRKCOf1GnG
V71gTNztB96AsMoTASb2n9VqTsQCq+FBmOmVxVbV6UfSY1PVmK0oFi4xoVzQrVe+vVdrpEG7z42C
IXRA22eST4rqczg8rhfso5gm9LfOF/35+S3poFNQl95EOTBmzymd+KgxnkS2xh59JTvrFxW87eF2
2zVFLiK0mpbf2WtWZGrN7SXgPsIQqLNQYAYRGF7i6LCogagD7dSgzsXwoDZMxUZR0L/iRV0Ro8wa
UWGwywMv/aEfqVUdr0n/Lv02/JeZUbWVA8FWG2LLTDbmCUa0fYJJla7HzBRUd+q9VEXd/ASJtYzg
kRzN/d2hwXM8nWI4o31eRdlvyqFVmXyuSAWxaKPm/0PhADf+hA0jHCrmUoFvi6AzAbCe6yfbA1KQ
INJ8BKUsp+JYefDVHajHH3lW2EhvcWqbzFJBee2JRGV5T/hRMEKkgnC/Xb19CPtAy06Q7mjTpKQf
6RxfPyK7bHRJ7hzDFokF7Hk6NLPffsJKLREagjfY2mZW6dn/buB+bl2YN22lfeMdj7T46lYcjJtA
SjAtvhC6kTYkC8pOV3W8EtgJAeIhGINWIm9D1ZoQkwvuWbIVYAmsp4Q2o4k0vQ+oJ05GLNdOh/8M
Hm+b1YIRQWyHI90XA+/+5Cm1Awj7l0b+cUabaQ3jFZSfbrIYbaJQE7k7ymx2bs51iiThpTa9COfz
qXD/00ODMQWOYgmYgR0XR3Qh/q3UbJDdYUWgl6PtA6tfo69si+OJ9zTPKCuxxJcck1NT94t4w5qu
v1oMgsrRc9vvYuyR7enMlbOBrvafCJ8xo0VO5UGNOVFPwE0WaG6LUehC7wDMujnjm1YqZS4fPK8n
ZXdjVWtUHLMKERij1b8cHi2PBmi2A1LE8chQW2pygLqFsho/KX5nji3iKoUZOU8KudLVHnN19vkN
8p8tUdXKU6/g/BML5YIJz1gEGJfX6MbZxLXtwCwrkuoHdTf8muXY/vGzr50i9hji53GQNynwg0NB
DcpWLGBD5dYAQrldyP0NZr9lI2VW3PKsWvFYJaeJ/RS/qWaemKOvXnmXAiaYQNlL9hLkL0lczm2C
cB/HL58DKSQrOWol2kLbsrm//25YTBcG7UEeGQdaDA6olH0k3WBgFfntuY5wXJQbDV+iKqF3EuA1
Hw2UA91wDc3dAg0lygSmPq/NFOjtiUFM7Nz7yUWqWeFcCk5HxjCYT84FgQ2Oa1j64EaAcz/umS1f
PJhq7vPpZJuXx64liFrLgJ52CUUP4ZfDwXHUOPG6ZepZ9Jlii5rDRT+0CDxhICdIqZHTfTB49e19
CwI7HT3/yPUXde3/m5wjt55mlN2DDhnWAEEbcaPLEarKF+ZTMns6OfjQy3BIP3dYsRNIMPpoVPyR
jHJhEK7o2DHMz1W6OyZY8BPSJT+ou38XbU23R/kdi/FVko65xvXkV2WB9DsMmGVvUP1YXYySLE4I
W41lghkCeG1sCRYfT3Mi3SQYNrumTUeZB5uDj2qFcBbwWhPs8GEcRMaAncckfX2uLBnoWSsVVOw8
WbzwjGCVx8dS2wysDcn4EAFf08ihffxnLEJnzXoQbpEKTJC5cVhU9gyonu2KOlDF++5gc272n9xt
e/2F7iz9hQp3+8VSau6Bjq3sYUq2ZhnGhM0ve5VyROkp72NEFIv9apJiDFf7T3gAQr5+k28oa9Ge
XYUu0HVwqfkVeQ7sIBdLk5bNb/fZQEO11+lGMj2lKzOoG5ZemLN8bb1/zUdObptI14GgzooV0cTb
bDS+6V33jNgH/OQF9UstVdvdI8IBy3SmiHX/AupEY12uMiOkOb10w4hgmXPXRCzW58AH+sY1fZHK
7Ykv9Jxj0jDBjiZQF5n5rOvqAaX8JFayO2xIwIhMI/nMy4rl+C9/XqzG11oRZgZ0xdVtEqBwWl9n
0bj9bN/orDWEbxagIk6lBSqAAkJlXsr6w4xr+khwkD3HNZoM/TQXq/BaePCXN11qid/ym7iwlH5G
C2UvEvAr7NO0poYLm9u6vqaUzRFVfKVTFC1XFFz+TNqHeA5lftqVz0vWKV7HYhSxRltSn8Zmkpuy
qcSn4MM87+yDeZCDKnOYVvmOsymD+M3fIYbiuGqPYgPwvAk0wIxF7WPTwzbFaSRfp0fcjucN0kPG
dyqmfpaHwxsP2OHcntefKewyiyuiRYuKSU3MZFRd8+XEHiwcNfM2dAGjatFP3xME0Ji3Hgv/31Nh
J6qWVfky16DuHhrtnlwuSmCpWkbhf5VPkovZ1diQbuAi9/1fLXDl/7rVtam7OLpXSYeNJwh6rZU+
ax9kJ2xhgp1b+BAmfXZto5E3KWXOx/0U9L3gl1FH7RnaVUvzmYP/6hVBfx8+KpTaNypidSMa4z4n
WtTA+ptWovZGPjCEHhVZ0UmaIHyqiYIoK5vqMCAXnGMzT+pNO/ypA9nE2XgSPMU5+kAXC3Cjd4Ef
7B/UEXXGxcLvPK/WJxkeCE1uBkxUTyhoH7eHxzNqbZl/cnii14VK9kmCMyRWlIKkK8kb34PhrE7v
yZsGaDTXqi/klcdnsbja2ckZKmU/obiJT7ERuvntjX9LFWwEMjh/BAjUVNcdH7eBQ66Qpmw8hAgn
0jxMdMmGIA3CPWJ7CUDIijqa1IpPiH63TU7dRFMyjRvp8ivA48QJMHeyUyvM9icsnVCiFJ4o4HK5
N+27/LvZGD5YZyrxEZVTR6oGoGUV8PNb5weRga1hARpFNuX3KQXjMgq80K+7kh+pSvs9NzLd8GpO
uHy86+ne002gQ8RH/eV1omeo1yDTJDNLdrTluOmeekF4P7gX1HjU7TP0ETtbrwuMaMEukE/GPU7O
aHRCJkRYnpXtuwYtGANyztM0AGwc+sFPnPKLlcXq/SxlQIBlJ9auX+/ZAhhwKo/Nev206hOhwgfZ
Io4x7karn8reVN2fCQWAQpZBK6o1eqFYRzwZnpa+OkET1yEwxUuG9hq4ZlQd9QDn3qFS2S00Si9b
qmX6EcLqtreZ9N3lcrrxoxYa7maFM0sWFxRmn4yGT9ClklmfjWqtn0OCjcOOqfaMoEa/E7MEWQiH
Di6h1fGfvbPTbN+haJ3s6YLd/11KiFS+Vn3jgMk1PN1h7+M06JiqRYBNklatFNa2pNdGfRFR2Ii9
EHFR7q1kCvWEjMLYDWextYeF6pohLUAr9Kw65/gDS1XECTOH06rfBkDISc9m5xij1Fz4Dw/nrbwg
VDo3eps48wbqA1sznFGC1itvvwnb6ARicC0ioeoW20mezCLQ8yiUE54ZAvyNPJe46Vk8d4BFJpcY
7XsmbO7/ctBg77fVJWvfJS4wHYoWbBBBMsgf26aDAeve9ZWGg4UiVy6HrOz+30Csz2wHlFINutXd
HKWjKcKE+1ARUMaltqHXNzIYgkNdcJZf1hbWO8ahvnW2TKE/XHByNlm3td62dGb9f5h3hCHMFqG9
h3zx38BwLQ4pwqqNaZHmOclYMnZ7UXOa8Criy4S5HtfgafbdogMIAprxJo34pySxNVGTgGl0Hj6z
RmngrOLIExG+sV3LVj6X4Vp3tpmz0Iid+ozfwpePc9Hw0GtJXdkPoL+77RlFZuU8Ec//226EufuI
19FZc7gVnRZ4ZeRJY4QXIoO1VNoff6fQ+tTbqGe63Q7VV29KhafWnOJ+sIP2fDJlkaRXWI5tqxNK
byg29kTgrlV3/8tDzBLOGBJg0W3T2acOE+JJR0PWjyGMyQqi7rvIBUI47OLpB1KQkg6ZgM1kfkTV
j34SAnbZovUGIFBVJ/QTgJ5PJGuqB8nL+FIpWaW72fQ7bSgY4mK0DVodOl761INFxbjhLmDn+7Au
CUMh24OKX4+WXXGtvSe00b2QTJEPYXvzqVnwzDFDo4s0BdmDIHoAbVNcpl/CnSIBBphqM7b7T/Xe
1b6Er1tPHfA3mQdOI4XZYPFUHs8+FNlP7T/Ov8nzE3XdZJBbHCVDsc9Jz+ycQgDIb5kW1nJL7WPa
bj8i1dg3KYVEom7DSF+0m5sv+UYNuVyeAIXBm7KAotHeMlT9TkwjyRlQVeI8wu1al7XRUG7oRgsa
YpoNQHAO96io3FBlPMLBffNlzF5uB/9lkvWjxYp5n7cAM/jT3vO1m5ANZmbqCZ+IG57yJzJL/pE4
ce6IZL0N53l6hEIUIqBsdrjYtXSUKownbYM5kbB+B6XSfY1Ts79unBKYFc6NVsSZyEz7WUeg2399
h6WOGbkO2gPD8I7cLfq68iplrzKRD53x9TOzfZWuSrnQSfpVdwOUHMvKj3C6C1VygLjG+uIRRHLh
KcQhAPm9KtHECLi/Gn4gtxnNRRsEpHLoaCHODFESnnEH1xMOlEtsVdjiSV2Wmaje9b0WM1C/y8Ov
6NXaosyJ7FXGs9b5BfC/noa+FJwjLmLLzT0g/kWpaxfcHhTY/IKEq5Rd4qscYtfWcPdUfYoRvjVy
e9dWoSgQ7lTa+Ol0fpqIk6Qgm2VEmfRhfVaEB+3XqafjczqojmxK/nhZDBsV85QjU9eIGZ/qFUIk
qC8fe72C1EVS2KMzZW1uYy7Cmasw9RzCYndHHI7oStI3OOufFfOYq2KoQMjClyYR25Qx23rBKDzM
QUiYdv/xoE0nqtFeCdQDuFCYn79f5Cxq5uKR9Ub7/7k2BAUoNJGrt8Xnm1DIx4czO+3hsw8GVVQU
cC3fTOvFUFhgp/XDZaweLMshEb3db8qTIbiUJV8c8PoWItITGfHJEmgiq60CzEHNo8DbJCOulhya
a4iGDmbaNPyeWEz4MVGVI6Rq9+gHj80rz5WQlu9QzM74yC6xXmafNMTVvj1KUpWgxsRdafrqLFoA
nxsBDVPM5pPkI5r7UorK4wNBrpLb5t+9We3WJV2pz5nt6QCriLjIlMMVE3D/kRWxmiDSUT3BCgvU
WTVx/5l106oSU9DnbWM+RUgHDfJQQBZtglnVBK0LDPDGPDpu9LsY/jcgWEw6Uq9xNbCe4T/3Wf7v
/PJqJ54aNCN3qzvLV+c5qwpM6rdxbFs4IV00uDox7vy2sVcpt0kms1/2tB0BSj5kzGgoNU7vtOvX
q68GYrlcgrMZGUQTDA4sAhm+Xjw0Ds1yDaPjUrVevMXnRNS+q3xIpHFpiA4AskAdMhuXuoLGfOn0
lZb2U4nL345oh4i14fhkD0K+8gV6wRp8gSZsj1QEHF8BMmjCzPA9NPezrJVyTEpJSvVWpROOZlWX
RZV/L0kP5FgKkI6NETqV0z/tqZet4v7t/P7wnfs/iSostgjJK/FnlgIgByrC9OI2EwNbS6sHEO6l
ADaDI9XInvOXuEM9MCziqHK3LcmwU0uI/m2rWrCSrVoScPOv3m8/zlQvO48QSjk1OdaLt4AYqiff
3wcVN8XT2KTbfXPWVVyor4IHyxB11XX3D1cx3s7Ig/rWLoDYKPZXkkktgAkQlsADZT4fyl1rA48d
OQNH0nRwyTPXIGuP+WPhhu8A/O0WTJbU40Sis+eUtOInet78+Q8d3yM35LP8+LquED7D6976ztmo
/G/IHVIiIVl2ZYzoRCQjjllafHSpblfeIKo7VdOYipbdz2uH04CbtVQwCv4Y/O6stFVY/lUYu4kU
vSpSVL/bmxkfJ/JPG857uWxImUqu1lYpR8wb8h/6di29E/Ehq8F6XE7HIZCDY2cyzlZoJnVLOISH
25GBwO6HDuIcLNIOYMi5Z9KrpN9roeWguE93mkYc/dYkNL0l7gjdv5beGy4cvKquO+los6lskPAe
bnJQGIELPWi+KAaOD/RctstEsf6HKwRdBAzVSP+6ip1qXkro3llpG3iaIxdM7Vf6yWPgZQRpdVWy
SOBjHAxEIP3jQyNkz91wssaNvmsGHjj9HWF820oaMlaYAjYNET1aJj6RfewnDIZi3b3lr4Hk+4IH
g1HXCQN04Jit+IpxbKAtfYYwXgfnhPvOgPiLeFdaL+GAIQGzlwLfG3oXIsejeD5IEo3WmOngcIjL
an+Xesw7Nh0t2YXy/rV0QCYsgp4sbCstX6wL9sGS2Rqd4Cv8UCIQwFLXHeQaKEbMauxybAyx8SrB
prfEHo2HiJcyW5Hp9dLko1EtGo8//J4rxKhuEwg+/q4yl8hPKkd5WK9Yg6SmlMdoFm1+5Bh1WZB+
iKmBGGrCqQNUsqhMmAGcO4pwq9QvkejHAmi5a9xHT0FAEepjWHVKY9vEhhDqG/JggcvImWWR+yfB
95GASiGyq/2PuO5TTqutk9tr7aO2rR/ZMleiyzwVczI4i+56MtInIHiuviE/L8nx+HgVzduoa71d
d5J68NIGFOyJ4AUezka59ZfL9XCrJDWYRKKGoYneZksOpq97jqUIkFLB3y9kxDn2Urqz75uDvqLc
sIZcw1MhcUWBOllWSjdUMjJxODe9jrzBfSWYXkhd0lotGVG6KZgXcGdzx+XQY2KdE9aRuxxDDzwB
NXujBbD7vw+ReF1kemrpebeGKl/k26bo/JMDVQEAx4jt1ewdmXS+2oUu8lUSnCoV3wViA4dt3w3j
LZ9AxJ/Izzk5UBxLHjvLGDZNeQDuXA0m1MZJMHZK3gyow+6HsD5lQQYoLcaO12pbAzD1qFvgKWix
JoZ1JfOhoahJwitP1OFbo3Cr747NEIKk/L8wx79fG1jRRfiYeM4dncUCGK4jNCXqMNf2qOoHMTM9
boZHYSfvb7Da4VJ5YOu3J4y6VAkQf8cwxfXVbS4LxijFUzw/rFQO9GvRnUww6ud3SNsbI7azhzS+
cPE4kc7n7USx/TIv3/Fb8ehmnJyjctmi5zME54O1qXcwRRxBjZnu8RZV7uc7GBuvBw6Wvm8WnUw5
IMdv8cK2246D+jfKzfyLb9Ki/S8rUjVs0lNgf7u9BGgLTDHXpWr5tNj7sjERzBhuuJz1F7fzxQR5
hU4d2HD1pzK76C9CRTGt3nQqJKzOkSY3p0CtNuKEhcnNVlT/tpvLOsg28LLXHm7W7eoRgvDNyFef
a4pl7M1xUJ4eruFOMaMWgBpllC5M+WJ1s0AtPF3TrQVvXft02wUwUF3AC3hChWBpCJ0GU6A5/WAl
POzcrZhapEfkjWu94h/UfiPEysV5G5m29mw4JjCe5ITgvQFEh89NC3stdl+gpYljbBlVF4tqBhMw
/os+i3kYgngJ2Yyld2SEjgdKriN1SzSnOeoe/cIMCBov05kuA3gtSNdr+keNbHXr+deT6eGot+9J
yvaJN30hH22sC8O8YmEbML2WBHU3T9VTBu460QupJUywocX8b59V65/x3tbz7hJbAwvczeyA4M0G
6Pg6F9hm21DUCmGx+0V3SyF26SMVw7TIM+GYW3IUODZF1Oi4SalucZ7dMX7xtrmr54Qwnq3+guCc
TolXiygoWgUbYe3MumC9STNcEclvh6FmyMNgWM4tWSWfh1f0mj/bIdrBLTG5+uDHzs/szKSAEqPY
Ej7kncr2AUmgC0TTMpQI6PmKp4KeP4/FI9MHjPvcpytwSNi1WQ2E+zArspgazHZ2K6ylu5Qk3j8k
sn2vqI8IIVZQY5CI4xWYYSXFXEhWSmqO4UqopJYW0jSb0up8YxrMJVMSi7802oIySV0cEZVbQ2ee
/bb8AU4uOeGcXE2HOROrGyktj98PqhlmifEGZP+cPWmpeAU8iw51l/MQbVfAh5+pq8hmvZC6eM6r
N57pueIZw7wWpzMwB5sGUzc6brZm/DMLTzcbIznzNpAj4SxSFMd/37SqVrx43Nfs+u1gf92LQVy+
Txz4rLJ5HEukdLN/KzIMgEPiV04lHwbmFKp/WZdNlMsoxxGqlamqeHPT4Y78rrRo/ShmZ8i600i4
Fz+Y01qd5xwZlYQanF9dGGiK7HprpdsJoZKEeKv9VPToIc0iap0JF20ALZKcah1KVhlaCdP4S8LG
V3JQrVhHzqLOnUlTqFMCLmq6qIDgDBpp9WA0ljAJQ8D6C9kFfNey8rOLTr/aPxNVeNjLNB4Udc88
CXZ6VKpmlhkfcCbNwdD3oPUHfZtkfOyp14bEmP8vKs3yiTGoxD5xA9hCfl80zJ4fdFU46zQRhf/I
JHRktRQuBrl4BoNBO3hXYaDD47kq0pGIeG1BKhlYVrNFMqs+oPs5t183iUI6iPAJ5pkbh1NUJU9G
tJMoMxOJWXy6F1kjfumDn9MJhVXP92O7jhkx1q4aHBX17PKUst4TotJcLIOHAqJPXyLlJlyGBMC5
n96FbaksXB3b9Vh/PgkBaCCHWYeOPp2L+FHMJ571Nk5kV/njh2u6PJ8kNu2E4z22FPr9iUedfsuz
a3yHw62HPmfaY9IiBbsmIlt/8LqWrEBjKNh9DpaM/rwHT136BRb8s4el/5gSJITEKFlfM+iFoAy+
3J+RmCiwR0BOqY5B1qzBkIaeOmPnG++GvxFi0QYEj5NPkvXj8loVbqjvnJSzKSVO4qGHBuXW+dg6
UPj7t/RgmKQHC2h325+uQ2bu+mjHLI40cRwroj0OEd5XJbhspzMzhjipnutXWxD3Lss7tJ7rH24x
uhao7I564z8mW5bF8o9D6GUUJwEywDs0h7iA2hXI6Ua2EfH7uaLDmfzA3UX21bS5RDUjJs5cI+f5
0fe9FsC8UXnCVbZjWLB0sgv398LbfzAexX7cX3g5VHOFS9omcp+i7H604LCaAvtuwfwPGlJRw6TC
6exJy1olZOuAcuN9xsdOqRKoNc8e+JmUA0goEns/raD9ZtcaB+JpwrqfR9ATQ6qbqqYnakc4xHly
D4ECywlHYOhUWnGk/euQ357RVRVAjss8ykx77ZPg/oUw4NuXtZEV2JF0qlfjj55JABK2qDBpS/qL
FUTnU9Eri6fC7qgwRO7PS8DRYz/KWuLUfF9iMpgH7dED0RF70F1yojP2nYfnDMS562GAwm5hGG2I
bGlrQBFja9aNY5vGNsj2SKPFbMZqiAxVwlC36TteJ9zHJMfwKOoODuGZ5SqWO1uUu2NV0QRmDmBj
sqs9Li0h5lq77JR12Fo93Zb9HHFZEvQccGvaAKgeyuyMgk8weD0HdOVP5gdAtElAAQC1BEQ1rc1g
VNAMl72Okr9PoRcQeSZKvhQhGIUg4sYLC/rUG6fj2DaEr4WWXgc11Mrv/UtAUn+wPhDBjb/mu7o9
va8xn31mozWdkDuXTvOI5brf8ARLc2tE88Iordgkcte12XVWzmy/Iss7GteiJ/jNPChCNoIe0HGZ
TumPF2cnXJTteTq/qNp9faf44V5rQI5zCSKUYEm1kE/0goiozwjamNWahsxVjYF+ZRMNk0EZwe6f
kkYG1f3NHUbhBIBOUa5gmcjMmh36tMD07z8EIrWQBcsRUjqAW8nSbvi418T4tYL7a+cQ7RA+kd1K
Yp4iI1XsqVB7MnNjwXYy57ZZuHKyReNnnYUQeC/4keBkg4GOylNmAGuIEQCGujOX2QxxovhRBj5E
dbGw/bAz4oUHBvoyuLYeIEA+rSEMSBtQftB7tHhVimkksuiCO2B232jDGuFibRhM6CdoT/P1KBPc
vd3olg+UnYNBQTmOfXh0LC+8Q+fE82kKbb6p8R2Bu0GXgh/rUMJ2B0rucMHVTaL9Bsf2RhBdd+Tx
sC5mY2Xbl6SnVz7tfbnqKuoCF4DCCT76MF8QpEOqytY95d95WjTJQ2Oz/vnekpa+2AzJllU/fxMN
4p5zHORTejWeUdI+jxQFknNoVbRBaCbK0eOY+KSYVP8dI6kjZOuPGGFQ1pBoyq6kMWdnqTd4Y21f
55zYF1niJg6AbHuBcU5J7FBt9XfnQrxzJ33cIdhZZwmpY7wFHM3t9DCN08W90xPv8cQFzIz5ivjV
25+sDw/l2SbitlFx88gK6gwO1/uH6dP4wIeLqJgdGxkxX93yIp6nVE14StZqxw/V9hCj5YdNsxYe
s1kPc4HiYQDQwiUYGgBx4mc4NjUa4KlzaegJzQd+x7kE449qFqwMWQMBGMfmHqlX/7BGYSQN2KIN
p7I/1Jnr1kAG5E53K9km14tPOQGTVNXnfl0W9FltQu/9vC/vzSVujucdLKs5h9AAT0HzwPDSg1uE
rHN/Ljpmf9NbUDUnQKmnVETaRuJzVqUjiD8uKszEWEm8baz7OqlEbjY9PYGEVECeOVy45+B8GS+g
2Xuhz5t8eiF81urApdY/a7YD9lUlsVNfGSIjqebEFd899UBOH0lhQkuwTh/rA621dZYSdKKZlFQM
1KMm5hIJGi9LkZ4Ld/jj9Au/H3jX+uBupZI1CfC3XWv/nvEcw1xyuGaN/wr6BQws58aR5nuAOynk
+gF6HBS1PZCg5pNTAcr35rXOCTct/rtCI3lR9YtEOBk+jp6UZNjDT4hgmaCuWMXpP/ldE+dX/Lx1
+/TjMgEqLZ6V4wvUxTqGQc23N7nK2/znlHb6rhLy84Gbo9EfXC+dAw0CbXYPtZUMdGGvoBNDb4vp
pqZ6X1efoPyEUgVn3677aF/Ej9X6Qw64L8wXVYENZUB/S+ahh02DlBOL62KbNfWpJ7tl2aBceMqB
CJqz2qJFo6NWEqpTnNyn46IUBYkuT5q4vnKR91wDbm2L1hfKcjfED5uhlnrgbxm2sF7lJQuJT/nI
2rivMDHNjV+a8OjGgpbdLUovHMIbXOrk7IXx2iWCnH/nW4rKrigZ69Duyj8XSICtuGB5ezQjhfcu
31pknVsQpP4foM4vty70wagxzEDUbZsjTbEGPNe2Br2F+5TPOKJivuNz+MCdgjHhE5LKYCR6fnwk
x6U7+vUL5ioopS483wINwrG1IzmSR+BJtM+72xlrQCgWm+ip3BXop9V6ZTwxoG/3EAffMqXWKPDx
O6BwiryyNdIRuc2GqgpSj3ZHqDp9ppcVtI1kpXqBOv4qzpNgx5WA5+bifHwky1eAnKVvJGMkriUr
XCdM65EJqJJBUeFBmu5SKJ86ZxCPvX035DqyFvB9mTXlgAr2ZfxVBZQ5h3ja7gyf/O54Tq+X45QJ
Y920wI1WNTQqbW6REPxytFWATfDBXRjEop42M96bbWxmCONY8xTbAvp21dbqL5fSNCrY468hYj+d
US0643u3glbG+Q4+9rw7AXrp1z3Mb3qTB6yidg6O/vbrN9hGXBiU807hcjt5C7hEze76vYzyuUgL
JWjPZUzZm+xGq6k+b+5zqFkcKoh49efRZVwfo89Mb9a70huLeatyGAXY9AJ+NREltZrA8Ik2jZ0H
oqFg15fTBGViWYLhMp4ldGr83cz6jimVVSviWicvzg+UgUsvlJ/T+MrOhtGc7ZSx0IBzExL2s7a9
8cu2BKnciA9tEA6+habGUJCs8mYmVqZA/6z/Oks+uGwmGsrbbrKbI9kFmL3AVKAoXyPs1mdb6FSw
YvdIwQfbiDu/vZonifF2miLzF9DvNH52LFJJBoYcfVGXKLgQUljMjyb8C7t3mRHiEzqMJSTBGc5A
DqrQSXA5mFRbOsfiJkV9WrniXuDK3pbE7z+dz0eRb1Z/Xz1ASHQV2iyd9LzAA0GWX221nxrpwnC8
uvgkMhzVCVFsi9awZ3aeIocApjDQU6eYZs/vVyKi6C6+W1z3MYHhFa1kgWSnSJTbRmepmyYEXWPn
rGEI4a9EQUG5V6IA5NHfVuKlbSlxKZPW2tVCwA8u4yvcAK3icM0mSv2gqzGXx4buHtqXrox6K1np
xYv11odevDaNOo5a5oJYJc+Uk0+fBAA32k9ysLYBGLErDtNCZLCNx4PJI3wMffp7+Ld2U3dh35Hk
3WVGg9a7nIPk3bXDaeXPYbJAY+fbfz5Oy6Vt81tO9URpSXkhwx/Rv2s8iIoUsuBmib+ywve+K19T
hByZJuXNykUCPC5+80JRYRUVWULNtr9iHWX9mjhq3Nfe99q6RadB6Wb3AnKoj8yI3Jhvh/iCGlL5
csusW0k3+GzFlVzKIqHh4VINNpersHNi0e5bJWCGdqGhWPEQ8e/UufjzNAJ01j1PUGn7BbQf137P
+KdURLm4Lw9178boO3p2+4gbCHW2pMQxhBY/fDUNRjbIJwsopafZwizraY4OXvfwbnGx5/lKcVV1
eEZLwbtFH/nLeGMR52prqoKF6ym85RRMx8XHyJ6fcbae/fmIANhl7UcghNcaXDAMQRMcHd7dpIAK
h8Iz25JWL89IS92iAivCesAyxi+F4y0TxwIHBKcZubG6V2gHTGTQ7QruzA8zOb4zPf9buuRgnaGt
if23QfsGP+LJ6jlgKq5sX8FaZVFgjEsoFc50AD8m5sfHIM3VTx/eBM9c2ovhW0RTGxLg2o6nBnx7
jfSmcjY6cDuNAVhX1msF2qAWuhLdMUJ8r8NOTtzoK7HJVFQ7uW6xMM/wgnUawKur8TOQ4Q2V5sns
gbBYpEdj4RkzPPjimwA5fmU/bQgOp6CKE7pxI/gfMar8FE5xxZwjGgDhIQXb3hvNEUnCK8qtZ860
xh0hvsFpHlHZDP3/vzlYsOjjHLX+1PdOax20Y8t3ha2lxP8oxg3MfVb8dG0NINuRArMwNwvjNwdy
obWxujiQUlDp0ZDhWpmSzm7e+Z64HOPO7gQCHMgsgaMEby3qp8BOFKEa865btOReJwakeG5gczS5
sTvvBh02F05JzJ13WLnhp678INfv9+0jrjaVqMyZq4DEeBJoaPIPDPBr9tK1q0QCcfuL/0pxh+4E
YPVPB88DNV0XczKQPYzmfY3VUHPuUgMPqNh5xZrc/0JwYZhovCdxN3hLkcurzVJecwE9EEZHlA7D
fQtS4lNerb+LWBMY1qmOKtsaKlGxnoRyYpmhFZunyd5UD+jEqyFdx5vbVekOOtzk40pKZQrv62dm
4r34ZA0/l7aVBJ70vMSg5YlzUNZRGlHBWzpka4b7mJFCoLbus32IkmQogLvRsEV+ZxUFJUuCoJiQ
BRBYw2cr6aEJ0HAvNvcJDf2SfWMUShUCKdBRhcN6CV24lpr99rTpQ8Y8ihYwjohbnxM66kCSNgTu
rk86v8VzDZuEtw01Guhc6qujAqM2738gc41YE1TcITM3W92qG/AnA4iKtV2aXygcBPfzePUVikXv
KYtTfFECBDdkmeUB80+U+LUTP+09qvdqOWXp/u5yCcXtxLTBp+aZp78zuBM/8f9ui50ahWL4PQGY
xSAcC3elmgEhovzCmDta7fCN0VcouLtTYQ4rlZ1CYUaTW3+MbaOcsn2ZSHBcs70zbsG+zJTYwB0e
2fie7aowJS4mRbqf7tUc0xJlMpG6/VJSkyn0/LzmNMUCRuM+JylDOd1ZhFMELTpdFgBtCEJ3u1GV
c3ksusf0ToXudJbuU1FC/GQtMrhduoBdNIr12JuNvg6QS/JW9VlyEnVFIt8oJj/It9fnqbwNnRJf
PO2zdUjHU6s3g6WiA29MVUiIgeQX0C5KHv4ocHU2CvK/VB8HYbmiLUxg6Vs8/lqi8c66KULwXhSZ
uxTw2/sA7kfuOztRPxy8oztRBB9bDXpN8fsCJIouSR6mhBx2SuB9+FxEclgI2EKANX7erj8b+BH/
z5xCR0FYgbs4lYgPbdNjIU2t7BuTVdn29JcR6aMYYvKvONU1zl4NlO1WCMdjaehYMX59hVPbMu0A
JCb4F9WFMY55rrK9UuwALtE/MvNsu5NQTJyozzTgssVm3S+PTFKyTidFO2kXX26dLB0DJ84Ynr+y
nqQzUzSWO1X65131UXlxpKu3rJtn8OzcEnWLQlYyqkXzRd+NvBTpMZM+T+inSJLWUqsg/xKdaf1b
gh8dxqwkbc7b66Wu8YiA282x0hkSCOf9hHVcX+kZim9T/UsFnOnYtoogW7Ya3JhAvo64SSlH05WF
sNNW7gQ8Xr7cjWSP4iHP2+hyuK8ymbgTI3Z3nBKnVnleB1p8SAJ7SqdFoLzD+X1e/34jiaA98YRF
ckPJf2F/laIiJ4zZvKotHMvhIpWSNY+8aVlUv15/iw4El1XxvAJnTkRpNo77MrP4vmm/UF3wt7oX
Ji7zXlHHDRoAM8f6o+EOl9NcRhYapMAM5hGAV9E+phy42oBhSZa9LyMNlpXKy++Ksy5VQIFNkfty
4FONZGhYAd7/AvJKrIjcebtXwpT+DnXX6b/icQqe8zY7jJB0oezV3ZluKXUZNwIgc7aJZ9mZnRyf
UXkbws/WnULV2OinT0V189qUVJeoAAS1GJH4cTiTRmxwE/NaK8muMhoyyNOOE37RnsCXpX6fLbDf
6PanFGSDbJRPqH2UwELdE2SiQ8U/k9iibOm6veISdEpd0AE33nr1VKbisj+CEKcNNKuqikoExdzb
IfONPjlp7XBHZ1ESVG/ro5UUlgAuo9rbdFJZGFYouBK/lbQMe0xuP1WTdVyQlcjxOIWiZc5zUrhQ
icygSW1szktB4c+NF3EDZZA7D+Pqj7MVnkeuEX0w9iBwk0yapWqJmmCLIr3IM3Gdo1fEbIUfdlif
E5hVBmcLzNLJn5vcACCOzDQRiYgeIP+ecsNIDsH7jrz2JZv3jS3H/AzB6iv/X5DPYn7ju1weeAfE
bPNFayGocuJnKTwrVESJmqwwxWDveZY9YaU+BRRlMQramSKT4QujEvIaFoATrBPZShhIh8fY783S
AV0JV0zwmoJ3QT4u0EaKHACDvmNLTCxqu5n6sPIxh5N7PPt5yhD6a8AgxhkyszD2QzRIpO9z+5iJ
5uvOfTeGI2Yvnka2QhjELtZzL+rsJeeSIGx01oz6vbN3K38QYUM/FXxd2w58T+lkGWg/B6qyktVZ
Hg7rl1+3RejFjVQnPfr2EALiOkFBgLZNtFbmqpeKwYWDOcUfkMzibfoqzxmHzW8TCoe1z+nBtvRB
pXXi0O+QE/Olm4STiHfUTjIMhDOVriKDWVdA3LJdQip+//tUlUSre643fcoZjveStYzjUk4g7AEn
vxLLQW9L5hJzo+xAJiX0Lab+qGQVwINE9bmY/aqGNUqZe4d5H5lCAUlrJ1WIYgkv8RvO+z/rCXuS
XJORwddYOUyaXg2Y/a2Prl8bMRMstMwsKcKcgYEVMn+bTUgsM/JhazUYaJube9Ci50MjOnEixwRW
aJ9Hdxy0qXKepp5mh+2XGgkJXUTK4lPDt+6mdmNE/gliHAJX3/BfGxi2L9GnWLUKHzIf8lGFOXhl
D17th0d5kas+uSe0fYEPHAuVJJ0BvhFkUcU1DqVgQLciwfm1ZvNdJ8aSVNuRejR7DKtn6TyMzvZA
PYNJJWNtdGlhLduFbLF1Sp2CNaTl0p6SBUCOYzhz/9d/y2JXR7ZP41Eb06Z3G53YJdOvmXIOnEhW
+fRVeNIAfnc9T9thm0Zp//Jw/7rgKkzODyuALjJxnTxROwwLptddks4MavG1CCTwBZ6bZxj1z3ja
lY6e90da0WU9Gj+A4YmJ7B04StzZ7BmUZO2ZGCE5ASQ9saM5zzrv8eyb7Q9YDBiKpu3uwECekZ/q
YByWt81QJYLno0Lg+glsh7XRBIP5PyxnW6TRR0PHF8nVrAlka4myHqOVhws6kEFJtSIjhAY+ONfP
hJC58qP3I41H0HvlmAM6eL6ktJ0fhlQuoBh7NFiWZXIkyQSyqCmpI2S7UD+FuHcF/o2a+IS2/EAw
h5j4Cf7KTOZEt6rxhUrZ2oMDSy05/R2F/aCmHV5X4JDNCpdFq10jhr44YhwHspCh++kPsx0RY7ss
WYtACTN/FMIymoeQ/aAdR7YBo1brcLtGIXG9chO7cH/qsfoUBprE0eCVts8QL6i6rZ24oV0q7BZq
nxSv0/YlO9sEwa3ul/f4e4yvRqu14YuM0TutOJE1xCYKkFevYgGrwznmZU71hsMw14rRQb2V9580
IXm1ByMz96D8XyRe07Ccsx1c+IdW0aFCGon7D0cPo3UNf9szrg7JYajOy4r8pZafIo0DzFRVsQyZ
z8BywxIYwfxv0V7ALmpbHI++SvNyQhUQ/irXUYpY3oG1jFWfsE/Akp85mNlDYwXXBOvpPfV2Ezl5
S0XTwuvVb8UsJh+I6/BhbkUn6pTt5XtMUDxad0mkOj7HR9WRAfXFbLuBVkNylBxopl1PL/kMS2KT
13+7gbx8Oj6/WCgyXW3oiBHdT210hg7ncVCnjbGUWxdPzM2NLTPdeu19JbDqr1mb+akpp2D538B6
ptTiHiS0xwz7fmtANqDh63H2h4NkW43NEmtGRfSKxLY6bQWfyNf+uA2sbWdmo1PJ6qrhbi/Nxp7N
HIUAKDLLRKrOyzbLZAMWgCCmuhRmCKqi2xhqdY0dtWT8V623rpv7KMyZtE701LX88EIvIkeFPWvc
QZGcVg7+HUlUcFf87Ecea9k5TBp9JWBfcIkvBIFmwZRQzL6SZmV2ALnDhy9XYgCRw6jmPWRcxKBw
vub1MrxZSGn7MgQsNgFFqEgwfKef4q9SUMRV5q4sPWwRef/j52A1KYkW/wrnAqlQhV6XyDT2dXTq
p5JkZZWPvsVqrTEcj5hag0OaydED0/OEIE2HjFDYdHuCRkgyte2P6sXgOLdjwxxIMcFal5Hdf0N1
txQek9In5YWWtGSwc4ajHT/bkcqxnMwwhT7l+TDYgemolrKrVzot+6jPkPpfrpAPwM74gxY10AQY
8HsKpMb4niK3piQ0aE8+JlQy33KeiE9+GJvrm+wVTDAOxcrR+lhGqSvxIGO6g9lxjHiotHy8Ksn3
VFHkYd2riR79XN5xRA70lIM1LEWMihzIbg1dkFJyCdezZ/xd4pLb2ojaJEX4HCki0zuEuaJsrQ7K
9f5IGc7ct3ev2+eGzz8es8OOdDnW+xFkTgNbtzxd74Ctih3zaZL5hIQ3vr36QvGssrPkAI3pUYtZ
plPTOlCH2GxAkOMNXt85aHfeocqR05j0ygOR6g1koWTPz7tDFXcWZv/2AV0dRSQbjpgJhpeQvT4F
SDCKu7c3mrSRHNiJY4IXm5ipVvGsm5hO214n4iRkBIVRGQaji/QfOHvQvnZAzG4lnV2oFKId7loi
56VKRz+CjX9lFp6X/75n5pNxb3AUkpaF4a3oqS5O30zuDZt52hmczxLHmJtMqHtF6ZDvC88Z57OI
YtWluFmswREZoMkV7NxpHW6CpKxnQWU3evQvJ52onunt8gpItgvXcOUBGdJJy//qfl8HU0jLhS13
Y0a2giCQtynpm/+LkltJo+zByXizRWdACvLf7lb6bbMrr+Om0HRy/hm/HPH+z2vv4yn9YtGSxhIW
s2VUaJPNKlF8ktplHHAl7oXXsF2WoS/v0/Q1APYSw1Ynl9VmDTGHVbHw1IeJCY0B+84d39kAKmGz
3Fo7vhAs4QVbDvVXks8B3PcXm/HENYXU4gjE22m/771EVXzblFY813s2lVAGFYPYTjk93eN5BkeX
HkkX1hvq0NtUFRql13sscCTi3WoONryk30oCWSw8vy07Cwx2RAnt/vixqC7a1wJsTrRG8NG6Wbsn
nJ9ZnfF57vqbns11+hhXwPVTxZkL7am4wHcps756VwBO18YWlA7NCeFXQozpDXv/piY/1gIRoGSv
m09Knbz5pwzYmSsK3gZyeK5eD1NPxWQIN5YlQ5Xf7M2GzZUhEVSec+XqnfWGARYqrc+n8G9tZM7A
2Brfuiwn7QiE47VJlZunzBcTCzuKQ27OTkQk/+GY4NHCxt3BX8va0s6+eJ4B1cy9ox+NyabB1TDe
gH2xlNISvEAkNZD5ksTQivIPi5iyqHoBPuIrQUX6ivqXmPCPZ+dZzQNyKSRY4kJNAbS0P3cXKN0J
sEZh2QIzqMZMkQaZP9pQozr48lcQgHLJ74e1J33HRG8HW5frNBie7wwHJDqdO/DbnXda9hQ7AfsT
a59j+CjUcOoSd0RxGYnBA4bn/MnbplED+s4T6mHdLzNdYZDB5Ye6ENK9vc/z4MmuhYjeATzVgdZb
TJ8cjx/MYuMsTjCoK6Jad15tTournUenDW0FlGiarn0R6E2Sf2SJ893QRouOITAY87oad7H0ot6v
VbNjQAd9mBHXUeN0Eq6drs153TpjMR5pPToXFtyFzI3xfGMFW1TQTyopDugBoA8nNHxXdBuCTqRK
hLfwhQejDWk87s08ZGiD2ZwYVIydqAz8m6vbnnqqoznCxP2e3SXLXpfRZRsk7Vq7drvJ8iWA8uuE
VAmm8dNVUO8TBKCJWUYmu7yeW7LgtNO+71ZAXbkNKr7IqELikTfpnSdEzda/QidxetGj/12BzKvz
C3SLziiS0umXY/Ggb2PBXMxOkVO6elr1i+CAM4+eKrJbNW3UIwOfrgj5qN0XF1qUXEGg522ljh/x
NC8qYBM/QUEIOcTKtMsUzJ0rYF3g+dko08uB+gO6Xvob2Ei69iyz3ztVUnoFliA39cN1GGXWZhhg
kYIXyu4U6AB6FSUEcUo31MET3ZreuvkDveO8RZzDr787DQ5dUX7V9CAhSILrUvT8FTefyNotChxQ
HzpJ0Q6uBksagAwcODTMIVIsuHVieZ+N4RsNMCTpVu1U+n2rDhy8P8be3gheDtl7q1Q4SorEXdVm
kpFOt53/yndl8KXv/HWRYot+sN5x6o/yYrDuiyxeI/IXW0TnIxWURlabkYfErvRCw9uUC6y6Kob3
dH6BerMG7xGLYMCXmtTDtv/Cq8FN9IByh149VWh3XHmAxlTRtDpsVH97O7NSArUo3BgowgAJshJa
iZ+CkZ5Xjr9+bS3IurnOmbhyeD6r0oVJBSCvjm1g7lkrvppVjfc8/gkiypfpAg1E0H42+R/p1x2Z
6ruJYo9OrD8jcaaca+ZClh2CjD0oE1Rp+tnKKmXITZg0SJXb7IsYqSOhiv5yu5oTp6bSamPCLyqr
Q9CDu/60lKP34oaiwonZJIRSl2jGTfz7ALXMVnN+8SoSuGy0V+2d5KiV0nXCQRTVm+o6XOOHkG1N
9BI1hdEeyN3t+81KTiw5wneUwDLys22V2/wIDqGsiQWaW7dGheUX2kHX98/1o9TCeSrDrIKG3v5d
BaxMZwqE9YME5BBuULzyKa8Cusux/Jo+FVrvlfNzCIES4sWvCknkAPFwxeDrudw02R1tVCCoYSnb
IudAV36qtPFAMsMxW+pQQsbfa/mdfbd41sIdLXua0/09pZjRulZuEy4IqLHQK+JXf2W424GVvVa4
zHJijv6FMQ8AMd9QpfXr/ztODeYfUp9qUSDjCHfVut4mXrioCapRc9diJ/6aaAYlfx0fpSAvbIYr
2R6GmqoZttSWWfiIHSsSjjsa3lC/qmjwE16+wZSXmffkK2tLdpEyavWKganHyyCrsE4otcbEmmtK
jMTJYriapzL3GXtTi26fn7YKCTvLMQIycBMp2K5BuXecWSxqKhbmjsjIVdlc1/NfcRCcLT5rqoFB
EE6aCDDRlIxvP/mxMYRZuqwA925My2NXj3Svp/qQVEwII/sg6mO1emqBghTM4+rc6uSE6Yjoz0Qw
bwOFWy/45GEg0eDIuUbTK7qoNhKpNfRLZB5UHQxLGV82ZhIIOPEM6kErJ5gVff3cGAvWDEFR03f1
eX8o8dQr6b8mhgj6psCsPT68LkffJTDjdTjpcrMqPKPulGnVlpA4Zii/bQAxCrECGeISoxejChvq
1xyuWRHXuFaLnyej9ysiIVwtZQCowWPQVIT0Gg5UIC+/LJOWC1ktdhRfVh7XSIs4PJK7lyVmxyFW
4erCOZwgErhTZ6qm8HmbxMsegitcnW7MHmi+GILhxUBnl6ygEGyzK1AphRvNDuK2YKdUdjIbiX+e
sL/vlgmlAImkdPlIlkIESc0HPNdVl9zARqlxlGqUhz/3n4iZkxxJZtX+AF39g81OXYM/ZLRTxmWF
q4TkpOvqT1ZDUxnMOMC6gOwqsYFwl4XZKlBQagq10ChuopsLI4t/KsVlv4vL+Y7vX9r6pT3NrG85
oPoLnnF2wZaPefR5l1v4DjOwI5qsPofsQ58keb4GytwOKJYhc8pqnoRxhxctA25wbAYcvWh9t0N/
5tmSzPbGALElfLD26PZpStfXQ0fR+7k3dIvlIjrWl3sZQEAksSKduF20pNvj+rf1cF9Yz9s9l5TH
8zXgU1oERgFbFce1f1EmDE6TbkqLHr575boAJOVLgbrHhyHn2gxP+orfmI9P1dVRVdKdsLNsNKK5
e/JY0BVokf2cp3y4wX/NBuf3Qnfx2l0C94pRzoX102f9Y9eEFQj4ZaI/cE67cnU49WJ9i0vYN+zT
Kj0fxSU2ZM8q/6VYQyVOJ/CtA4Wt3Z+X4FvMTukEW+tMiIds762jmDofgyjzyZ6kQlcoa38sQiGl
UxuK6Vjcy0QT9urJCnRa/qB4c6npJrcFcqKRP/1XRSM5bm5kE/vm3hbL7MHIxlleCTN4Td/sijLw
k4yrYEQR+PMTeCQMBkoApRa9PUc8AMBvPZKHn7niEruS53Hk8/xiIvesbFbfm+T1J9gYLjJ9w2QP
fXPZmQEeWeau/GFWOhpsui1rD2xChsN98JJHWgSCtxTfmuL6CysW1/Dnq8L8pV0ESlxypfRaukmM
sFV2adHyvRS2eUu00Ft9bt1Tl7+nVkGYu71F1yDs5piV8gGHkvQPY3TKgQDAWztXC9Owpg8IgtT9
tp+c2rvcjRZ4u7QoKoqnOpX9Q3xmrx0tPLwt/0EV7+7b7vNA4Wtjl3yfM2FA7f5DZf4mhYCspTF2
GQwjs7ZJmoxFJftqqS7KhJHXPXZhenyHlrfR0TM3gqrttjXfoq9m/QQSdlLRL2VzfMcwOjPYF+e5
d5MEOn3Cg0pbu+6eDnJzMnChSCvupu2ht4ua3+hisYB4pVfIMABLbrSjw5qgxVyVN6jnGKBHy2bu
fChJ7Y+oJsq+JZDd0p3blE8ifE0hTeMQIxfz3j9v3zAvMRPJ/R0ar8qc5fO+aovPaIP0mfUb8gdz
Ono+V+GFdFEWwcA+GNdjR+cQhtb8YvdgzDMp757Sf+OKT1gQhH+Rx9d5jmqat3mu5g8/57slfsq2
m98EdjOkO8lSdV+4Q9DhdPdgNcBjpUL9HiI04c/JDJFlGJD9FEX0R0XClUxKhJYP9vE2PgtfTe36
FKwg4bBDtbf9J2rn1EJnUKzk+ABZ4FI0HEesEfG7dZh5XmGZHPEgvCvZr9vfmK07Gk577v8kD0XP
x7ds2ctfkrV1k/+Ya5hYR26pcjpu8tXOAnvpQJxxYM6Co84YclfqpS/yEBBABePiWhQAXsvpz0JU
cZHPa2oYlzxmrh45435Mle6WaCoQJN6wzBGmubneuu6TGajltax72JL4aTecUsC43QfZwPd56k4t
kNSv80HsAWLcG+x3ROXSZdUFC3pZ8H01o5amkJmQXcdWMbftGQDafpU717geAkB5Ml7XrVNqFvWl
ff/qgxNa6sBds3U5Z80p5fntdWMrUXUCXvvqgr6194uPPFKnmK32nLvJB8xDIO64lrUQOKDa6rm4
q0feW2a+pZvcxGOI0nHWV8xV+aTgcT34AbevwHSmdZoWHIwg7KFbjVO3Wbe+XaNogLE6K0TcKbqX
J5I1L7RANIh46Qd4oPs4zUzrvBp1ykeSJXGZbh9OUOG1cYxsxOgbWhMGbxpwOpXHYJNJT+XEATLZ
5WBcxfPYjQkoNktqVgQbGXlx9Rzn2zOTecFM+wiWBdfCNoVNSQAvpo1uoBYNy8+splXYp99WVEHZ
93RVcUz5Jsu+Orlj9/jGxInY9+Br8ApRVkCgoE/NFVad+rE1qfnpR/Pcu/BkhqnCmdTNI9RD+1cB
v+D8T21EWAMY+x3Gq8AQHFXQDbnDTHkuzvUGRfktWBeu9Z8h76a9I1CJzBjvqjnTMTvj9Rla3yJ4
9nXHx+42wopNqLtKI90HF85HyPmlq2ZJwMEhdLfeDShnAFGrqX1P9cQeChRYgVeh9EcXQWJUWB+5
8bksyUxDrx7JF+AgFq3tQ9DPACk5sBAwKIgq5iNm59QCV6eF3/zjRwCuhOKjWpHHtv5btjLLmfzP
aHF0pves69Wg1XJ0mAxMzAgcmKTSh4leTY6buKG9KUMm7QFSD+EpsdeH1pp0oyrPpfq2soSYS0AI
F2x6r4FfsVNRQphT8tJMrNyHoWciUSnfbD/FUUtxoOrq/a/6S+Ir2QKBMFZQkBt3Ppz799r4fKcw
1KZh7G1lWY3UaQiSFJgeWA6SfiRUGbaPc902OGotL1Ef5ULNZTD2EHCBAXbrmGzMXTvExTR/NveQ
K41hSnetiMt5kMvZnpzR8dQMViNfehoPfWc8TfJ/1uBC3ZFRIfqCSe5HFkM7+EKrIcH+9Ze+Lpou
QpY2op5Akt4LQJSv9bpVW6O2ZlZ9u39nSr945J/UcuNmOJ5kp+DJ3NbsAPFnqcssNgpBNUFhqDs5
tjz+Q0PerfDkV4lIoIUsZmaiNkDV9iV9QbCg+1ZW7xE0lqq8GBNjYc3lo47EkY5QC1hFcGs5uHiD
E/Erl8GaSOWHclkmLdyyjpZ2CHjtXpBWr54Pkh/AjYIjY45CNB+FxdMvXkYvrl+xklfvT6KnrMK0
PK8KesaQprgcoaRMqyQxXL++WZdRFIoYscyvAUSWSsb5VVcblk+qqmeUNjVamyfW0xvTA/bqPFZ3
53rW9U+8vUfIKzdNvl2tbmvXYUmI6envZd//IOMlZca3LxNy7SLseki5/gm5Jd77oJ+puXj81+3w
VsHKMRiVk8vweWWyb4avxaGG1zp7237sjNDKCu/Vrdw59Mq8j0kd0S4tAjk8QhupqdpPY9y4iQBG
J91efaLQXiYCegUUBrH8oZw52XwwOF59VfQ8RNlDgJdlwH1EnDpdG3JrDYvBx838AQbgf4w3Zzfz
8U5wEV+J6afXC8SJI8UGB0VN/+be6+YqldY5n3CY8umhhG/FgPSbMNkHUxz8uzxiZNnvkXCA0tdZ
loAwAip5AZQ9IkPFDou9neH4Ji0iN8Xn7FuSNF5zMqFtwAvteWqBKNH0H8u/8Z3VK7xENI8Ekq5d
n38UUxdSrl1kksTLrvimbE1Jq+Z7ET9OgFLDa8tKNfsBDxZYVUKzp/ifBrSQFQgYLNFE+OxxjjHt
Nv4glA55oKFszI5ufYaltkbwffS+9vrMPdH0PtQUZLZmE1FOZI7vGWsIvA78UTS/yanG5Zbd1Dhw
tC5N3FPYIkuJdmpQOk8XtQkX26Hq1+ucenDFwVxG3ai9w4yB4wrKjzrpCvbK91HgHkabUXlq68F7
v+GBoNgRT2v6fpLUDh+5c7Qvm1U832vQ2dxN/BAupiudZ1QqdJ9977U7wD+KCS6o1HWloaFsVCs/
1Pz+VAkDPXU8rke6/SYrXZhPFUYYYr4zbE86LgVgoz2iD0CkT4XLmzc+aFtVtyklgOVho87d2EDF
vOqiKAZVp/It2pmOJXD+2NF7SW0SxlTZeb3sWFG57n7L22aV7doxWC03DW7uAWGGDfnxgKL2Ql8g
YjwSWuHfO+8mUC9hUvhjzG0liaampRf8Qumc/w4xlOo+yGaLRp5iWheLC8C3uLyko7EHuc1qOoqa
zGqFRx8jrEKL4AA/ybtnK2kt7C3o4FCM8RTLRxmDbg0og7vSCtb/HhQdZ3r1BqAN6as2WCTP+8Sa
6/WuZAjOIRFc59jdLLAZb9ap8yJGNPup2aL0sLjViNBtnbzRJzN4/PROoEpvETpqZRqqZE6U0qIe
UwU70VtdrvUXNHMvaCe5cDpC20gdQGXNMlS4mCE0ttWKjvYhVWVgO3cdBQoJVT+LCzqOlssIz8z3
/yMoK+jucrNYioNp5SSjoGyhFAwUvZxUMQ+SxNF8meVdj7QH3zkh1XSF4/ajiCgg5elG4A5ttmBA
zuoPP33Jiqt/4I/Y5wycJ68l1eCF9ZfZ+ENHvsl3uRyfImwNvXhR6fvsBqY/gf6DWqdDVmrPDkPY
KDfGbvzJrBc5LSuoL71quepZWiHnORbyr7NJ2Ey6aO+aCdm4lfuk0n7NQ4jg/H//WXg9xP63FVJj
NiczQFSX+tADz0IgV5zWDxHft+uz3gxvnOuOVh9cqZIpC7SZnBAmJOp+hbnAA57FXm0O8oJUyA84
spMBAR2wScVFMloxUyg4SvGt8EK8xtWtdsXyvaS4dPizEISvSakNjDnjPEv0WKiPbjUbajHpqQ6C
ct+kWW+hWhOgOE8Z/JWrAhR3fyzNROkMA/U/1t/lrv+TYwqmMlx9pm+RmxloGfSMa/kI+/Zb6mr4
AJVs4CzKIGNnP7lqTOGofiTqYUgfuKmfYN9maym+2JJbB53x/p7QwQ6r/wHpvElhvZeXcxfn4FQX
9jCZzhS44Ufx1GlsNWHteXX+N0bYuf9mZ8WkIr0jtf5kK8De0Z4Ac0G39KFp4hiYTruaVTnlTHie
f2XmsHVF/p0xxJi6qbTuzRoiA5IHZAWQYAxeAg6xMYZ1lggT+N2sDRcMfknsF/U7VBBbVqTJktfO
dFke3Q6rYKznaWsB9fYtfFtjpAkab/MmQ+V8F3VmysDXmDRDdFgkVuGbOWUKPEGAv6zpvdPeJnVh
dXoWkEzkvSf7Ag3ZS1Qqx/lyFeowNeG7JcPzrLAJlYMSAiLbKEOdPYCq1b0DUCiBa9dLhMmpP/Z+
HKj6ZM/WcINzA6f+jFNj91fR4Hq0es8Tj+9dOD1A+a634pjPG86jY32ojeQr3wKBT8lHToZVriXn
YG0QnoAVE00TFSvNGd3GYhJ1vcX7kharcL5Z2WQJcnCJR0wyeglbH1MZV/QiWCzth9NfdxwCuj3n
5I0GmLkhTEl5TQswjfXO9tnM+htrO9ol7hljtRIMOSk2vEvNrmDmZk7xIs1Z4RGMCTcBwr00Qa7E
/ZmJQU0oQHGrPgP1U/AE4j6waUGaw/W36z0Z39hbcU1qrRe1jC+Di3bd0F0U124XrP2L/cdW6hXg
ijjPbB/zRX74OUZ9WuiX0wrX+fmhlQb72ddzsA5UmSLO3hQ+RCplUnvL5WQZlUtFIt8hEIHQvE5W
GYe6UD2G9fiZJGAKM7BQP3FSKEJ65boVs6fqqBRcERyDujP5P0Fm9qv9lq2CwEN369rGKdwrPhfq
C2/TGZuED2zBc7jcdsPG35I/LwkDvJSNiCmQNsaiteDs0O/rXAqIBwrKd1SgVIokJRsIZN/e3PkZ
H2Dyzz76FM6OEOPf07A9Zx+30PaFVCtKuaNAFz548lLmpdZ6GJyqCYn4YEg5DDUQ5108y4BYBs5P
KM4Ii10k8n7i0uENITxiH+fGY20JT/BqjD18+LPTJAKiw9V7eFsbIm+n8ploInfVICePwmusbBqU
o3qDhfzdQyVCSGa3knZEDAJhlaWu+lz+DknvRi4ocWshplr2j5dR+Y9QnDbsaMEUz7xOhRiVI5ja
iiN2a6hdorKrJd5vdbR2vOsL0lhmItcMnXuM2TzbjsqWprpiIQS2h80SLVqPKfGALgMnXQ8tuZtY
BU6CUDSxUQIRnDHK+AzcQUUy9K2p1BMXv1vAFWiuZgC/uY+9udERjr8g9bbu7s0RZSibgetgpWZg
HnMMhjZV1vrNKPzQmSiFmVbWzXdfFXDe54QYJhsWGpQ+SsyGw7ujLaz/GoPMeM3JArkpqTwRo5+D
s/T33K46q68pSbAzIjCCZGnMzreU5lqy8gF+qutcESBONWkm9Stj2ZAWLhsjQWYHbEM67y7lO1+K
Bvf3unckjFb+Cw3837Hj+47AdAg+OeWBpuOCTU4zmMv5RO030zeXXPwBg9L990d/62QoZiu1R4HR
fkVn5zfGHN5oPciAnEe4+qBvm5mlfyP/wUALyCDJ4TGbVQHSnqKkI/UR6nXT4Bcp6p/9rF5h7yPs
fzZl9Doxa8iGfgUQpYwgXg2CTn4svyC36i9CWQ+Jo7mEj+5Lza0Duuyqsl2JnDusqxSmVYjb2Jta
IN0YIp1dXF0Opj9Slk6DoaySo2gjkMkwtHzxZ1Gn32YaivsiaZK/YB9RixgBY093Ga5TxnPM9jJw
LBYrB7xrUJnrscil6zuyOXvFrRnnrfYdntYQSwY2wmI1DMxNxGu4/CO1meJnNesc+3ZLDhNU391u
I5NyMfUUeSz7Gkgh6DFQCkcntNEgOO4NQGok8PPn9WOtp9mVbD3BPEkQBPzFbFrpiImVZ4TmF77l
lD64vFLrAMo+ERqg6eHvLQqHmZvAKKFgZ8jdWFR0bxvRd+ewSKIUqBi8+/kzF5a6FEM55WB1mAuI
phOlrfxZ3vD3jSmCzOW7FGgWzZoZsVrS6x78hxmzis0OvBMDDW3tcT0lKMyX4ov+9+66Br1AMkv0
3EV60w7pwqRATjMXHl9Y6TmaqALZlCWPhwMDTJYe/0bEsCOYiy+MSL9nG52ebQlNxIEy9VhG0Npi
9YNVjP5IydjzBJDUuWEsGxFfMxot0y8xoGRLMeyFFpP/0bRSWZZpg2a92lwe+U3vNVkSQxUH2yrW
8jqw3r3OebykgSLtVUy+F+DeLk7JiboSzPIEJqnVpQDwM03Qa0wwyd4Rs3Y7mjAkzPdL78aB+tg8
x2vDpLlDX7dJ/bXLl3wQk0q+UThLfu018yJUR4MgWDe+0p209gGeWyrrqoWe3Jz+iaJQbJzPEV6S
YfgykMNiEAsl3elt6PnOq1v5zeEThXbWfqrygP6Tadq7t8m5IsfCzvZ42DGlWX7kk+H7KuImD8Pz
GJrHKtq143Bzxe/oBWJagu39miHNo4qQzLW6ERBC7ok1OAezyBl5QyI09X/gU4Vdl8CcyEVfK6z9
vCnOLg7u2euNV9V21xvKic5EmH7zF1KhSOlhY1wD1nddqviEAkMBYEmDNPe6y3Tr90/An9Jo2EDQ
v+CrrlJbozydoWjaZqZ96/H7YonN6Be9JDBPDS/UMGW27vgp+L0rFfvkS4gRF81jkHW6WwfIIUtm
R8MlnPwEqqomAy3oL5mH0XMuo+UITYtFpP/NZRmAL4nwWgLcSpIF7QjvrnHBOmNJj5KQfweoPVGS
uRsHSNXNWQiagB97XCjBKyamRmxWEnsZPiQSkpnkRFouQF8UuSaCeApMon2wtk3nWhHsKjF17BO0
uxWtOia82098ricCK0h0Dk+dsXeUYGh423SF1FxMGWKh2A2LGzBECChNTn5cOoFxWSoKGKgOxvXE
E+ulWWRzSAQgsYvAg3vsebgJP24Ie6CTMEzbGCSfcX64w2njwXLu7ItdmOqZMCYcIiiOrKTfl1yz
hxBMYSu3nFCRtLD+Lvnip3bqhWMoBBGxtDGeRFswJLNjqxXWxRB9e1aePBeKQJO4Cq6Em0qiM54/
5NcMmiEmJAdm68A3Vo9/UTZsKqG0/tWE2zWXrh9L8mIuthP1ZZqPb8segKrK7iHmB8PSuyO0p/sc
/EmzezhCbQ3G2pY8uBlrtud0xuRvJsyl3LZ4dMhirf0+pm71duBkK8ltcowKMtQ6DF0GBPQVluYt
4GYNcgp2jfR+bl6or75CYV66jxtgpMpbfMKUimzB2Eoe9G1vl+xkLordny0cTqzgsjeSHgr9PS/q
hhhWZdPmWOhklyfHKOLLqf45kFgwn0c65xtkYlWh7076Q3eWNRtBDwnExbwT7qVXG6GJstL+UFPs
P5CWck8NtxL4UDdhy2Y8Xbo6CD6Bmfz2kHMYnMF95ikpAVIjYBNCb5FwvqB4Z4RD+T7zG5Z7PY4W
l5PG/jV2qs7QYRJVhlC8fg7Cif65WOYOk3feCJ9+NoJnItc/SteNhhAEFoYgkEU0mroqBKzVehsJ
kd8G9tDjncGrxF+70IL3soALBMXsg0G5iR2gXZ2yPQ9ji4B9wXOWsvy5kAw2TUBD8cjMuB6ViFQY
t0rJbioDaY2sBHGj6vsHKBFAoLNNBx3qORtjspjOANs7rBCozMDXYdR/RCfvRWdBIoSiycfc9JRR
/JwYt7duIrcxypPWP04vtXOcOWV4/TuyO6s32G97bunzg+/jYiqQmaxHahV6/wvVZmesgLDCAzq4
eGMtX7BJ37/4Br8R17hvRoH96Jz/GRyoW2VTW3lMJAaqiFHZeJTGEb4lJ+YTH8PJHW05bo0xDqtk
pA2G9idFVmGQI3WkaRCT8GU8QX3f0IcnpYsHZHPZQHQ4tSkfacwcwvThSe+tFHgzAUdykegcxFIt
8rBH8eNj63x1ZixkIADisn4fV6UtghQc2DkBuZv9OiD3E8RfRitTrDXhfxtCBmBGm1eMoXfWhU5b
EBfSS3lpzntqqIjnBlJqOi3saFpQmTKxYXg7rsBzz4nw0TLzr6oQOaoFVFgZGEFOSkywvYsGt/v/
iq3pyZneoIE7s7MYzMWXfF9mRrQrB+ZpyZ73erToCHGBq6/A7Qmi/MD3DEalzfDP5cuznNkb+Nyb
pHThJfcnOyfi9NYhtSB4wmvQ2p/iA1tFM+QeO2OcFtU2Vq9/b9PmCBzIqz8JSyAlRu6qvWUl1/4l
vVa7+wwauawnX34QloCoBpW4+/pENxQkv0VwIf6zmOihkkfdKXtPUGfJ3JiQlADS2X7xYFZtlBzF
4DVKI6xkaz/gmOR/1KBlpKUvG0WVVAzw5OqnXk4SLfXHR8JmZuFFM8ludrYllRWOj6XJrSWRysbQ
txL0yTpgurEXrMNOXZz5vF5Z3RPVwAuXJXNS23PZujr5E8Pa0gQTgiGbd6QJp5JbNbdMuuHcoL2i
DF2ujKqtZGHP8AaEV1mVv8c2EMQioeg2bGGzMVKn5JYYTXG/Mz02LIJ1tFQWFuZn0iVpi8fNxVRm
xiduyve5hEI5xaMOcT9GHCx26n6/lHk2y21oEHl3n4Hw4jJWpkaRBIGSRN05I8tZtlxO2qozGfbq
GLFvSkmXfNs3gu7RRrxrOVEzhG1WMxajQFo1w5b+xX0SPG6s5JEFl3bwS1YTGMtfwz2hZNF5LIQf
+ymqVPkz1AVUpXH3BqHsIS3B68l6L1CVQjjCDX9wJeJbir+2Ae8AiaFE2wmnuZESXUwv1+WC9NBC
OrZSAKXkJEoGq6JPlzSz0wQs2uDnGJZ94SPcYNxR12P9gZWONmQf/8Fys8MrwyjO52PFTvlaggfz
zCl98CZL9Tb/BWlYZlt7gnpsboQ2jiElCs63mf+rfGsxKDBbA+5pmQswCAF1hRou9y24e95+TMpn
6yhmIou7APEeoeW3ZPZpq6YIWFgEInnsRv8Eg7s637p1HV7cnJRsULSIhDAN+XO3ZPlYnThNaq60
uKp/W3ruO3zqB9ISEhD2XZt2WNZ13AB9rBnBN4ueEq4JmD8SxRw5xEnFiygiCvDJCv0dSGyilNtm
qcsR5yZFiBr+bSXplRYMMBF6Zxb/sviqca/e4r8OXYQON8EBHcmby/NhKV/bHNbHBtZuwdxB9P/k
xjPx+5c2zwN2y4gbox0xKkrkBIjiXlcaMH9k3EYjxaiWfz9z1wBed8/AuIP50RQRLRpV7PBP2quf
ZZdQ2EkVD7iliRC83qMfkxpn0HOA1glYU/s9E7c4Wt+ZyJpq4RxqlUqJKMjpVKWHh2EgiEQT8e74
9cibsOXZL+dVIloMrEOIfsNGWZl/mcP9ZKqdoDGjwruXqRUcNo/b69Gwk4yAXgyvxhXJ0phNcTDe
o74JO4IgilK3Beg8796vtrd3qqyyqZXs67X/jVS3iMRxVzw6hG+xt5SjJq17T70JJmIXccXGDf5s
gl7pIeIPSYe70YFL+qlts+4TYZxUeGiPnUo3SFSkeQI1yfrjdm/UoK4zygSq8jbTMHcUJIPWGLh6
cyY7RKcxFsECB0jYL9NBLiquCkOZK7iJR2a7Pyt7bLqTt81+rAbww+zmMmrFP1Dawxd+6mwjEl8k
6s3KcX0oO4V+YKv4kpcX/BPXLhz0Awdg00s8+rB64AgYfDBDlYep1iOQjJgjhgMpDo6n++n1qt1O
UF9ZcqjjQGQ8/7JhcSfugRQVIW1koGprMvb9qhZ+ULY5PXdvIfhnj1JstLU4UZJaTEfECqNmJcwV
zA8HfvwoqIXlcFtADvrTbc1bnDKh2yfHbvQt+z6Llk93kmEKvKHao65JzMoCTlFy+YOL9J2oeReu
cpff6K5TV99oucCCdHA/hCkvJpHKzvAELYV1rr7FC2oH+N0KzJj/MBeaOPPnmka7q9ylVoF2Ue61
b7vu2A5Gn7Txey0gBhRyjVvh6weZHcW78Ktzo/Fj6azf6TeIS3XrpnSzyqUdEOBhX99uMF2I5AuS
wCD6Mia/JHpfaXdm102YXQmIOKHMpiI+SF38s+1zAPsFhCkS3SG3Xb7cIGO6vLbZ9xffpmotSJut
b6S1L+1R8g+HKf6asm8jMoxo6GNJfSx6F6Tg5x9rPfW1t8nopeLCnLy532HSCQGCFONuRtSY9ihk
HGyhaxsFvcMyyZzk36wkgbq519LgojvTfdoMC0Rxv68NdCV7E1PkIHrZqlTyH31W4ydKCSmetUbL
RMnx442jy28+DtntdLtcDbUQSeBPp/7R6QNMgymc7zeV0ADZ/IjSU4E5B57hSlMNPprijCprSh3I
8PHapdOWWbFfMapzL/Bn2t/0JoKePpUEDrWei3PciWrc5TOP7LdnGdmkt1vdfn+k1Wernk1uqIDv
4aZZMgGdoA/Tn4lfX8nUVRFioaKbb88WvGu0BBp6iwdnXFIGbwI0VCqdXhC24BDXCHwVe0vP65r7
31bKMYy7xdb2QWz3188eW2qhmh+kKGKLH69XVYLWer9/c4K2oGjRa8Rx8NinjxLvPZqDVS6Cz7VT
I31f7St0IbjDC7YVKhngtrt7g2oNPplJMmpYTRZ/X4l0bdImKSC5EiAlzWDZJEcwaKtuHsJqGSt4
Yxx2z3kF9DXWAs94m26dPKQTtHY4xBO7QVpkFJn1sVFY3uUIHArfUQdysU/3WFBkIVFBFXjb9z5n
FZyiKvb7OBTQyBDM8U+auDsKzLpB+ghEdS+XfEL53fCazmhA6sK5idX0l0pKZFoOxQ1LHZlMIaWv
zzKIaeWU4T0vn0GjD4QLdFFdhKSsIG1eaID+sATEdZ7tiKcirp9UShQQfJ01u4cUNyVvB6MQGM+h
ISl48JehJFeoW88b/mZXb+owtBNfZkapoTlJ+/k8o88r4yNcoh4ONdkm3zV6xKI3Hl7xkwGkA6K0
pBENJjZBImq8/0NsYAPkJzr/xDi5gE0X54hdPyiNiRQFkcsugHxG6o4egxFAfEBy3VxToMthXPPY
/YQkpcItQS4W5wqDSn2lpNH64ElOPc4ac6T4K4+vfb9j/LC/X/JQ7k0Rhsr4DBoNGllxMBbt+jDb
HthCFzvjkTtoAzwBXk+y07dZmKBBVi7pUwi+5luLgtGutbzCKANmCSt/G6GXbCcSXfTb3hfLT+/E
5NUJcIFUZJelbscC2ayjv/dL3LNBkJEuMEgqYHI0i45FnX4hJcDr3YUhVzb/p5XXRmypysIem3CN
IEBq2+rKCgQuXokqSU0IUGYkc8Rd5+MilsQZ+IRElg1gWZXN3RYaOaS4Il6695Df5ESddWg5xiNV
P0C9Dqm9ve7HiFPcPiKLpJh4FJP3cGg9zXuqp5s8uQV9Z3otFRxbbkKXsfEMeWcTVZoFWYCtJdZW
4e8oxU0ZstNFY8aU0SOPXYBKz/fuOu5DEU1ODZaDI9COZHdi5R6dfv3t9AAnjrBZ/gHSMkJ1u+AS
X3wHCJpTSJ/PVM7ZmkqODtIPPdNh4eStnYDy7onvmXKTFuTNz5Yk8hB14vydRpb2NwvxMcXH+YfN
fY/QN3uBiE3+z/gY3riemXJeyijHtU9nUyPGxyh01M6iRPcdJ5Grg5+hTPSUP0FZjMv0tPUjQywq
MupHXXjCUjhw1MoDwihnvK89jz4cGySUUhYSJKnYasO14MsSYmiFBCbMnKhvrKuLbSHVesaeuyQV
SpQIoDaTpZxQ5FASwCW20FeVUNqiDtdb3QjHK6IEYwGneZPpsaTcN55QeAMDoyxuvYi0i/soRvcD
B9xxZeCU77cUzlnJogpVj0XPy/RW15djz0GC1VhqW3xz+JC3qaM4Fs0tBCpUqyFvtn6ptqlamg3M
m5e5obH2qKAP5SfJFOynNAHdmde3KayacXVfHX6PIaAy/TeXi8tLfewN4gCd9LfB1GpE0Y5zSaey
6laE24TpbTNjzkF+Ix/K/JWF0TnrG+sSYW6zsMpvv20LSLAQ84TNk0sS4AHZahN8NCyzMIPpS7fN
SBT+K0sylo5ygnrwtL5fPD9JFEf/yR0f5WZiwDJFovqfeNV0Y4DpGCZLDGBlT9b6mbFlpYxz8vta
xms9M8++RUh74a5Gh7OcXBhYHNWuWA8H8fUTVQ2WjMqA81HshZm1VpyHZ3qGriGCCFS5PYchJyNo
kHnFo6D6oEJWPh/7GFAbMWfYXAs1tqxHtyw5xRtheNVS0YdHE5z3sM6fO0tu+XywTwhW57K6n+2Y
NdFr0IWaI5LhYPcOEZdeQcaly65z1kcr3ZT3jotB8pD0wHZoar8CYbBQWcwnIxGpgCBIqAfAZe1O
N/9C6nxIzCTMxQFM2wYuAzq16WVn6//lRUGKG9Elf5VCh6CCLuuJrf+dwmKCuD/itJuOGBv/PC3M
kuSrD3ro8HAHmMFpwfc6zRNOYso6eU+9USmg42gJr89iFI+UCBiFu6C8OjZWgjBWlL+6IsTLqZM/
/T0PxdGWxfpSj9t1Bo/+O8F0m9IeCNTF8G2mDJnCJBrkf9JvIF4ZVBhxT5BSRTOPnx7GPBslWeb8
nCYW1klwwlTwMv45d4D6/T8T3dqlDF9UWyWRUF7fKMhbtvuaohdDuTAIYv9u7XzCkitcURrUsp3v
PEyvm8PNnuET/jxnA0R1gXGylXbkrjIkjpCjUATevo/1MjSJTimjr5uobKN/8nU/iW9NH/AJG6Is
Yhu/CoCa1YORf5fjNMMdHzu0QuuVL7xbiqc+i90GIP4Ch/uexckRa8YgFfMbdayGDi/2P94pkRik
f3gALIV8s6mytrzGwoZnSq8C5HOqt3iPR90R8v/GSUu+NitwsKYIFoVofQjbKFWZKk1niV6WRirl
FSJH1+Kvj6IGyd3vnUKrkC2rjIynIeHUEIMMcCLuOTl2bxVvce7w+/t9Oky6cLKTzEWmSf+kEU+F
ad/hJGVwMDNyUPFJwzwUcGj80qXBRdDTZOaPtUsEU35wiGjvA8lRw3UTwbcJBGPx+oymeOK+c5nU
ByA+0ahw1Tk4YRwIi9XNonDT0ExHBMCNSHJhofL7vxR1hjEPo1ONNyprPCUwLdIf3psCmvxK4yrn
wQdIXluUMNDHEqZZOBfrXLLXCtGp1TEtj+K+epNCyr632TEHOjez4TGx45VotsR64ojDhmo9MTWV
D4gqjMBN3/ibawVuPGgzdNTyXU64TNdMUeA84JnMxbAE3Ami3bsen6tVfIVfMYHFkmTZ3+N3cKTF
ahYIw5PuT3syGCkn/mLkZ+8yHHEx06xgcUPdgzlh5ERR2GTH3S8xMXw+PGwXJGlfU4qd8by4Dkja
dJu63tGl+6f2smfsuInCNxY7yy7y5EWtXtjg3OUBdQ6KzNbnTU/LI4X9vovQtB/u5ZQYbsbLpZoe
IDVf5zQJOuOzn666pQ9G1cvqgLIEXMGIMkjffbX18hQoNAgEnBcwN0opXZkYeMmgL3ZsiUpeQjlV
gWnIwklgMsiYCO3/qCOJUMAjlm7N9TAArzmk43s+jxBDWjtJGGllngqAza3A46fnGS03V601J1/x
DXDcAAc67DD7dUTmWOLgszjOgHRMP++r4fh8ytZWETN7Ohlq6VY+3aFAU2VMsIZq4ZMkIQiLipZo
YVyOIhM7qTF38jlmEnsPlXCZYC5MOudN7Wd+FuhF6szmSn0DW+WKQKcZcVInNSltXA9D3Wmusb+A
Sd4Bcb+tKOK83Qrq42GSvFXtPERl57aQH1Q5CCWEX0mmUswps/M7Zs8M7d5tMq67c9+iaxRJNwDB
SRYxNSvEx2cB9hJTZfhpNZeBNIsUOuivSDrALzk74CxGz6Tsog6j61vhxGjzaiHf4KL590C+UBdw
ctK9FNrl7If2RUw01rbsN/OnB8sLpGYYDIyoT0Kn4SAEObOPhKH5XNriCOiDSHzdRo33OQOimQbq
X7F0twcTuswajeZPSIF0wKrGNin+EswQYbk+QbSbwReZ8uoMKMLb7Fnws0FT4mpZ6JKC3HUBekYc
wrbL965GoSE1pJjhlYRQtrEB7o9TKrt85KiAxgjWnEl712S2PKo1ovLv0anRxyvCicn/ggretNnm
X9ZxZU7ONeswW1RA7i6HPDAHdRsTP1sxubCUgCDCZKud2zwP6PiQJCaBtsQZa27kLN76k2NLlsci
P5gHCVnIyo4tl5Hwr6Yb3qRfEZR8i2XMNfxZZj5qrAFznNPN3CG+42CpYRclYAiVp0AcEbS+TCU5
si8CbwuWBYWrrE3c1IN8oEGmdGWPU9X8tZ8blqHCyXa9CQ12TMzLnciYydT8yn69QlSowHTyfPq6
96oxmEUtEmqAfs4NVmz/F3PnaQBs/+4WNlfRQwv1KYiBruU5KQtnUu0y1iJNs8J3F3UFm/4vtbKM
UqEbJFnSDBwMyEvhlV4tPUy0OtK0N4aK08ncos6b1XhM0I0tGGawxYZRNikfLviaxYlKpWa2lz1J
c4KZHazmXDf24qgm/DM29WoOVt1O8QAZxu0XzwvNb+6qAnwEoyZryp7SGlC84Gj+l/U+I+/b+/1J
tgR8a9aDeX4C59Fp62Yryz0bIldj7ECnjrfI/a/FaC7DYWn1D/bPDyByJybYjEXzruu5RvnGanV9
J4kdpFlQLmcMwPI1+h7GhfSely7/r2Ho6q9C8Nxj7WGTKh9Ut8JrqHU9TV9yHHEcs7+i1Vz3BzvT
5gnMJIp2GjBCTUq60ilO+kx0zZamUbPBJI3HJzXh3l7sodfVEIXhp29SjZXaq2ZA84HDsL7hwr5z
tBISzRzoVjQSi4USANtmCZYwxjBH0SNSnw6LMGn1HIn3b/jn4MvKCEzsqxySNalvFQoFZ4BGmZBs
FIcjQMZaNiXGm1kLcMBCoqT6iiK6fR23bvR28ftWK9ilFiJhW3bnnh5mlYfvnQMJuNJxkHuVSx4h
x37hg0arqCW9sOHQPapuUWSgp4vbS7NVsY9u1ghVtQX90NlfiTEWZf82xBPhoxJ1iRsyBjB4S1v+
QwP0SmVuN3gBLFjr9O2ivE1Pn2esnHnkVxcv41kyxTjBRPwStcaN23xoCI/ZWjsa39SrtByB16ub
LSPUriX7k22hkwJdBXZfWC67i4mId9AH+7aA5LCivLTpoEF/IFpr3s8o796mVlV/6daeKPutGaS5
kU0a59SWXQ3Rdv/tWuMQypOFy7NBRC5rPdLj+jq2vMUApyBQk69tgrKyMOLnyDkWZoDobYPi9J1m
CPM8CObaI+PxU8PANnxxVJG7GCgCUm9MyCfrO3avvwj4PYeVXpCNi9fBZ8/h6Ku17lAn9ASmV2Z4
qsLdVl11Sy8T0vT4LqHVK0nClGDGQaRb8DCCXGFmYERmfRuG5Uv4TqJhAAuRvVFgWijL1sihPWAB
gOSDVykz5ErNVc2qrK3MDx5CmSFGYoCwGSQu1bejXrjDUZsIBhe7B6FE4u6XRj0Y65YDz/OgK9fz
0GqXI+8cgJzlBjr4/SE4BGZcYRxXaoJ/B6e6JrYWCmoGNCKZeb+0gHgQ+qXpug3GgZSDcO4fhbWZ
S7zjWZN+8S7n0q+tHUsHy1kp0CbmPR7WKBnX/zWe5+BpHKFmYh92pafZqlLRM/ZmxUve1vTOB8MZ
Spnpw2thYm4USRFylq4Drjre1ev6GmyzTMcNwvbUQCCrL21uLswlXIRT/mFFDHxLw5+NswI/2HQh
3x2ng7CFTuSYUcRPgV0ATw4vzf/vyl7Lrjbyhyff+Hl3OIpbRExiCQV+mlbXYAhKY3P0yOUoYG/9
wcjLivKrnkJlcUbTdK3XHfbRdQKdNBJSKHfTWO9woW/qaR/vPjaapdxKMRr5NOL00RNZfv2tcqxd
DLDrZgn2BDXaaCXK4wLQrdbKE+RuJek4I5Ta3NyizZRXOv2hYfT5FR3QdugruDIvkHVTrWvr1hDx
sUFklv/+CPoGpc989JoK2rzteksSRGDYx+j5IUKJK2qG7RijD2aWM32RutVqdoB/KLbtnBE+V9PM
22xhFqYNiKL47CdlfY+/ugVcWn/15OgTuIpdtI/lTFTNGeswahEwZq7shHkZteidrBYB0wN1HxN9
KqMZoVXvdC4DGIsNKL5dlSu8zqCvlNodapQgo7oINjnxoAqjXEjmJeY53e6CPvuFwP70NMJXKtE3
RcaYqpN7yf6NKWDOZpQhjdSUy9tUXnSvLOJGb1bUc5e4Pz6fJ6Luelhd4kJ2+AlcXLfAUvm9IjhC
ydeNBhVpPrvOHnVsjkGud1ZT4uVN0Rqj9eJ7o9yuYDPnP/gKrzjgFXdUPTFgk6sBQty/RcJ1vyFX
9Kv1JQKnYUv/JaVmxADVnN1GH9Pm1R5tOofQqBLlGkYW5gU8hqOZ8a0tGW7M7sgu9t0zKYw69UvA
nMEhUS5M8XAO+V0bnYuiPBbomf49JJaon9d4YtgvLVwlON37ygXsZlgcl3q4VDW5W1s3c+S+3EFK
SME5IWCQUGMmfFBGJtRFw7agP15yZrIs242NTdNIb0d4BAhpmeCfgfRvo0ooFm18XL5b5bVfBhf3
7tbD3NIVQYqATh4sf+Dp2PW2UCIEZtyb3RQQo8Ps9vVT1eN5/6UvbKdiKV5hfPGQAqJjQNMb247U
cNZXywKkKTpeLQNKipwA/RpXr3Yo5F8wY4eo5sx2h9qZKNgp6U0oIGYP6b7Vs4I+6L70NovcyWho
VML4UeKNlqNVMHbjkC7YxwMn50DntMDsUH+CvBZfq8nSYaBnL/bMn8kmBg3fRErkH/PfkS+pmPZ4
Tt/KrsjjLyGCm0LiIUd2UH+rloWnTffTZcxrRUrisE0ZsmQpuV6XS9A8A+lQZdAKFGZZozzsjsu8
6MHuUBTIn/0yGyRNnbcSIPDlwD34u2YPjne4QnV9i3GQm5Wl/L53fO6A9igjzc+Y1OzOs7X8Tiql
5XISO11LFUWyOsibsJUTfoIra8aPRQ+dB8IQkfWSFyahq3+X4ZbHdPtR7Zk6cToplMkiPbwVlvlo
22rJRmzIWcx+lfNXWxVzoRMFDOK3n76WnsfAYNs/GpbUn8NSTR4q5eOTgoztMwl35BoxD9/y2X6W
L4BdUHdWNm5WDmuiwM5YX2WoQHARrNfkqD6DES7XfdXPIYZ3IfZTYKZTHB1f3DRvYYHiC4IKMszg
yaHJNGT2ugdOGwOu75X3cp8O40iwrRY7jQHmWnDTILmtNnPuUg0M4AQSEFwJcbMb8XjhG6UBXgnR
7njenCPtIQOA/heM58CYMEizA6aNrc2VUih0QIehNRZR5xWHTuBOimKEZaQ184NkNvjv815E+mGN
Ah1jMhkqe21hQO6x8SU9UxqWRNYaTfGeaDARiQLTMEg2NpW3c7JarqnZiqvi/IYDjPzyXMZdY/mO
+JvtVwXVBSqH0k+hCX7+dQntOWHidYsHPGio1aNrIuwwXwvU2W3mkCB5fIVkSrGDBVd5041AcRiO
Gw6+FRNi9YgWKokXQB/RfXkWjE1Uaf7gfNaUYg/n41EaQikvb/5kFovyyFHM+l3cfjCAmV0YCznJ
tFR6WWgCCfz/dg6krbUdvPT763tclnI949S1wTkmI2FPe4h5kf3l1BlxJBZGEP/IaxQc+x0FT/8Z
Zh43D3UrR/bq5seyWtAbagjS0l47Kr+199dFHNzVAULVQfNXN4x8saWu04LBJVNAy9/RA1ei/IYT
aABZnZevvI8MSLHiEQXQZgjChXboNtO4GHkvjAUGPdWJh/pjw48DvzAVZ19JXiaA8fJc+w+y2oAv
YZ++aNYQTtclDP1Js6RwWmsM15v3q7RrCYXSr9mlylWAh0WtWFjLpHayOi5/cmyV1lMDDnmgoKjT
NsJYkOihpeO2IayEs7alY1saH1HTgs+ly9vflB0pXXynJ3tHflSjTKwLlhBxJTuxJ6NDsG7/E4tV
/GCW3ON8yj306pBOYcph5dqTqDjjd+r/W9i5BLNKSbhe6QYzjByB6pbAX5A2kms3H3SedZnz+LT+
0v73KuBE7MWVeDs4lVjEa5DnZczsx3c4vhTI4zh+zlGTw9xRaAs1OtqWiZVGSHd/UaLQ3Md6yQqR
vnJ32RRA0zs4qz9qPxqROEitCrhQnqUzkqG2tmfTW64h+uQqmPIvY00k3LlKbOwy9ON/4qYoNLGG
F2wUi24k10Fpzuh+l768pQReQsmRK7e8rtq5MXOY65I4MJyFxXmzq1NOy7cfwt3E5w0Syi4V0zEh
110oVD0ZW9a+6zFswtuUmxd7R9WTG8RcIveqC7DiM+KY2SCC2a4JWrOfCiXzRyvwbQ2eiFtCw4u3
RsTFuhK5T6f1R0EaDEkFw7DnMwbHM6rXgq5qJG4JXyWsQi8Iz8hr3wdcS1Jy7un11HvYlEzo/FiY
pl1eBGT8Ku3fPe3s3OqmpMW6rUUqlMnmCrLfdT4EZexNqLuCPgEoWxgvtvr1LVQVteTCkeS1dvXi
BkSJM++z/FARa09+iShRUwjYmYUGyQlN4z9VuX91N0tl/oK2ImajSrXXdWyGozJg6/mPyASy5tY4
wIxvKSVt9MDx1mWa+L/oYDiHOlc8WeusPGMo3mb3GxdTN5MPhuSgmFwGULk6NKf2CHsvGYsThs6m
KLLpatoh9EIWjBBBrAlVHAwNrbIonE/OoEsXh71Ar5XvBuQb3B6NDkLYoFtrC8wm5PsL/JXZuZE+
eJIFVtj4548B9/qYzmD4G+swF+Xi1yhjBsRG63OSRd+ttwF5pMT5H1zfQUgVCrhfbx7lEuJeO5/9
Fblfl7iKI4ZYN48dsmDwjwr6pVPo07kyC2sAnCfkEkPoLon+C67u2neCnaNps4OKbYIQFL2RQeNZ
5Zq6iWgEut4xxM7Iy0tuVcY5fhi14WSocOO3mzpY5owtlIJiZG3cGCC/32ayeRU4rgtjspLbbHMc
MRKTJXye/q3ommMwVi5Mli1G/R8dDW4Zd2K4SscGxhUNCijRClGa2//LlkOlQgP1Gb0+u683LkiY
n0MWaawDCEr1zr/93NkLQTaMsIOydg8VLhqCcOvHdPuT03R3Xu+KWx7jwiXxK98KcVAjzDqhKPPK
0OXi1F97MrzgFENCJWXDJ8fPHoYuhNcklBMTYyfWKuPXpNiE3xGhxzeRENzj3xQnXzS8egwyf+94
cPZ2f21xtvXjvJd6ai0qaDkMj0p3w5a+VLbDtaQcT1yj66dBc+ioPQvqwC7fDskVrdEaOnlEmlmV
M7kz3xWTh3bhdsJHemVCedZkkVGp9VoS734YI1hunZximN0d7orJmPYow98mSswvB29iQwxOAU4R
HiXn8s7hpWsF61kWd1A4YIFoAkKhgHiNHGOPet+sgGc7DWS4TUJTbGNy3svcFL7E0RnmLjQWA8mu
/1B2xLadwqL4weqzL1MNmT+44ngPnFSgJ7Z5UAhmZBgo91ll2ShfRRknLUmturDOU7SvRbyulWzg
LZ8pkNIr4MTCyDk8IHDMmprqi91+O7wWaLrE8ygu2RkkvosSNA3mm6TfM5mU7bXG5OM/zeeU13KO
vFlSfLX+KPKFc0NvuNCccym7KPfEynqx5CuKlgYeS7I3hzO+ALgvf1gQJ/sprY/v03BIaJzs/YuE
hSXeeBk2kenJszQipt0Vdh7qnfSroTGNuPSWnf35yNZ30Iaw0ApnmvNRa1WcVm1o2rnalVdpSqm+
F5hUSKGc0kSJd3e71WfzSodb8RyJe6NzZ1GmMLs5Fj8UShJgCzJCnX9xhunc1v4Y9gfA/PBoaMcP
zc3KS/wIDdy3vplMWPnUQc8h3gpgKfUrDHej9vQ5CcbuqtG/eX6V5NmcVgnlSmuVG4oe/Xf5I+St
MQmbsACi0qswXbGJn4+JT1IvQXAM3el/xvbF7uMTJ+MUjUNJSkJuqbrRmvQutw4NhOeoC8YuwPa7
ouG8Otde/hl6Qv4Yrlt/1BrI3rk6wOcA4/bAalNdRDRxiN3hSws6VT9HqEqhlcGcrc494mXAr33I
szviBl22jYUQFd1olY9JM/DPAw+YsyBGW5SRc2pf8nI67EidKAdAoXT2TyRfdgiVJeyBFyRBy+9L
X1xkyPQ8oE9R8nNWB1YP9I2xWhZrz2fPVNTSqqZxJZAqIVF5koq+KssnuSNbPPXgH3zB9UPpTBSC
Jneven7JhVTIgGE1d1Am5ogmk+9yHbMqlAW9e5NbRh2GoaXDJQGicdSkJRJbKXyLlmiMG9kDU9Bg
EadlRpNL32Iutmx/7bMs9i6F0g5DSYVyWZejAU0DrtxnR6ol/4u8CEfU5ZqJ4VEEdiKGoPrg+UiM
dlq5jIR42OBWvfg7sZzKf67wFpR4Ea+IsPhFcX2cnrUt4UyZr1gbSaIPdADleeiWiVP8kjTG8pel
UMSkG4TVzq/5Z9T1aBwoOlFx5NLRUG2EWTV/dHO2RJx/8Jyz8sxVWnL3mHVJdDeoqb1zLMasY88s
QP8AVyOEnENQQbma+2oGeHWAupL9Qdi+MxZ46ICddeqHffgJ0ZYjPlzo15e3Sx5t/A/3pWsCCEXo
TizJbsatWoZYMlZRgKStehm0lkYCJ2w2NnewhnJDEjGR6pCNvL6j+R2V6GyF99zRPXF75YAQDQLg
QlXd8C5bjR4te/0RQOs+xmeAERzAnK6Uat9PsRkYd4/xGwzvUaAPd76h5o+uCTzvoefvn+DnI17c
WnPTKJ+6NrmOEGsBDktlrYSx2qOGf17L701f1+KWvJZSSe9raXzR9OcfssU++/FVoSz4GtTJarBQ
9J93U4DGftXGLhNQ8hGxNS4Y1tcQ27jVyaq0aPFZhQ1THrv6/uD3wCP91R2+2QiY6NEnmBTeuy7g
c2nP++C/SXa7gcDnvkz72Vf4xvXQWyyx83vNfEvxT5mt3r1JM2qV6r6ElTVZrw5wKUut72tkixvU
mjnUNdWXJm+Tj0NOEhJt3ER3SXOhnxiyoJXYFf+eqTSFc9h0LTQvDXPhbILP6OFgMVSGV1ZftkUe
AtrkdETP5h/szWvS0QAKsUxrM2oS+tphKn2dqWdtDR/qpXcoa3d3MWoGNEczT6cuEYvoUHfLUSIg
pIqykLqHAuhAURtskaXVxOBMg4R9cXu7G4/Ce7khGCgvn0QmvAepaul6DsDR6WdNksZA/2FYCr1K
sw1tOiMeWnPSIIpn07WBGkd6UKODzQtjMbd7Bj9QvNFrKuoXj1rKdTLs9+6VwUi/iZOjLH5pywnh
t+zL/XKfj23twt383Gi9/otKmOrNqCCGZYX8tAEqF6LFFLY4p6oUuYZdrNzUMIxpRYe1aC272Kp5
tFU1HWlpGgOpupbfo5Luwdn/BrH5AkASkmkhuOEAag7XmZr+OxT3mglBmvt2VANSk2MPJ5JNNK/B
78Wglv/pzd24P6YK28vPVY03GGCgkzPCtGRUcp3RJrheKV3i2hIHjIqn2KZrC6hUQZbX2F/ixdTD
tZVsQ9RP1XSVbo2yFJhxYHGAZvTB+l0rOBm8H49wk8eQ4UJ20CGH9+rIg8tA7ZMyeMLeGHpBm4Qv
K3+qVtIh+wFxJoF0dhC/7Upo7mjArjmZtoL9loOouvrqRD4C47uXHVWxT3Mfo4Aq3Cn6/bq94Kgx
ZL6pAH5kbmrhu9R/3W6Hs6p9xHwj8jZpSeErMdF2o4eTvINcD5haJ6TzziNzuyn/hRHn0xRerwlP
H47HvXqY5Ewc/CbmCgCUG2Tusf+OXXigxB9pnG6C0DBnrwsxRU3XT8jG3WuERWV4qpOWyd5AiH6Q
W6tyTJiL7sElN7bSwX+ZijpAoppllcrwWJG25FfPfLBUdF0okzsffoEYZqwRt0pYeNIa+twj6ty2
v0orsaeXM0Q/T1zlBcJ96TiltZw7yGLVqlCWaQmKdrqzh+0/leGO7L1WCWXenCGpsjngHdxCc1ti
Ob/TkyACcvbAAKkQD9QuSlElwkcarPlhwXFVROYEMid4maTrFR5sAOU4a8JgD7jAf01tdKfehigu
Kq0TTkZd+p4Zfoffw+nPS77rdD3rewCRhFxLsbC2Clu2DKkk/eiOjPS8blKPmQrNiLgXOBLgPgZJ
nQjedohJBI+Gx9v1IZjxZLCiAcNI+c9ZkLV1+ebHGAsd05+ddy3tBob0fZS9MobcZpNKkZFzVKyI
wDfl1hSY+XAGIwQ/KIGG8TeCVegrHLIevrz5Ga7NUOXjM999ecRyHs61n8OGaRytLkYqzlb/0WFQ
KUpfkbUVPurQWTNRmIaPF3V5EBc5c5K9NKgJirQRSqowI4zvIP1UCl6bWjMlRsCX3IwhYGk4y9FN
/lbwIixH+CJ6D/RsvuNHInbQxaubMZTlAKsoi3VENum4WeGKBEpH9Ac3cuvmtZidQsYm7tYII4NN
nPTHI+j/nIRfoZOi2UuIRPHcbVdDJmHj6hC9pAHHaroPaonUXOy4+pUBt09++Wr90Jb875u7XDw7
RO5/7x4Lj4/9cm138cWBW22aP9eGQLrTvJJvWcwuYaZg87RUNLUxes6HjMTq3rv4NikI12FabgWB
ESnarYcklSh4zURDqRyJXe5ateQTnaHPgT90TgdgoTg9cdCi1G1k5XY4v+vxzXulzsIXTczIPBaV
nb/Fp16qVfPWc1UkiXwecRV+RSAl5JF2z6x7JoSsT0M8krrzVjN6GJTmFqGuyLGJw8ob+XnUxP0I
OJI07lH3iW40iPCPydA7Kgy9H3lNQuQP8XzPxc5CEfTJaQQ95Ty/4HDBipFjI1hYEGEX5HI2lFdh
ZpNo6Bu1ehHwNW9LtK98eu87BG2oaPIhvNvYxyY1gxKjYY+LdRHgIRHWgZ36Nhhvm8MHIM6khMpq
2f9cVMbfmqALhgDkGNDNfGANGau+zqa491/i0GXvFFG7LqV2HdRHu9leqCR/mKX+cmvlXqIQGIVm
EIAvG+SYEgFy5GDo9hayli/Tiadrp1VJMh2IaYeb31Uw3ZM53wCIn503AhXN4m575Jh2lZCJ5kDe
gw0kQ3oeZWm2kMNEvxJoBGTYLPlLmYOE6UELbiCOciVY64irlG93F57PK9LS0STxMGTSvOy19vNU
6L7zqEc+5hunM5h2LbNnty4YHHhJvZWDMFAHKyZZkuFBM10dYQbbG0CGfnLzFksRGiWrsUy0gBqt
R84yqj3dkuEXWVk3w1JI0AyZ1EeLGH7DoIs24qdONd2e7vpzBn58LqLOXg4nYGHYK0hwB/SFylD6
bD09TvyVW0lARxIbzdYpK4+2DP0Mp3YzCHmeteBCaz+CpiHYr5cqzXZ+AM525qS/j8nxXxubGvml
AUBC70CPl9ofJdKt17fBIJazbMMTUPDz97OzX99vXTlxctpepQ2/swYH9RYg3O6sfxZtniUH3tz+
CosCZJS9oBI+wyqUwqNs5xh6adJZjk4e++dPK7l2jcz9ylSvgZt2QzC5HAoClSiKNSsLv9r07142
Bn5ak4HUjnwqcnQJh7XAB1mlZSBCO1jvuw4X7V3qj5pVci2SHpyniBbWA+oNFOKBtiTcOHV2M736
x9e2Q+JLWan/WVEP9vKtDKj4evB2SGV6ub+KzRRQnrK1VJ88xJvOsNcamde5dOAohv3pkYptq98j
Tfe4zQzND1F/5UGqfSe2FfA4nzQkb68zmZBpvuNDruLoLp9bosx4lGVnkdblKA5vt/haSO+G4vrq
QDafu+tGcPZc/z24Q8nxPr///0R9K72R+w2tS8SvU/HemJ872l9DTwpMrlviu4aQxz3UKbMofbKL
LkC0U0m5skNhI7rFacJUBCdn0smoxGtWlaUllL0mo4KIOeq62OGYzvaxtIU/Kw4jGOUnJbAr5Fvl
J7aLY1/W39ll3S0DPO6M7794+1/KRE038eyxQFO2BJWGBryceRR5LBjrtz5wPAuSNC5QWeaEYB1s
CepvuSgdkLAmBztW5L7cQwBQNpyZ4oH3RxZoOVdTIy7evX0HJ4yAJttrFbuMzAtNQIYJuDfdNTU3
U8zJmXxIRtctc0vMH6bhRNFSkByGue7Wc5MgX7NUU1Q1jf62DrEBG2XLV5BFn82cU//MB5f7RYaS
zCLj138OmN6ej0mTsyJWh5udVCG2xMeWxzfKsubPYuYX+qxSLz3uXTAEHP2cEfhBwJ26NZs0xlX3
vI89bjgeunDL7b6Y2/BdMhOe4gnapeo3CSigKRD2Xp4/1Ye1cCvtZCIv1v2Hq69apq6/BL53WsTH
I324yZ8sTiWlTRHhY2aeWN7yLQqDaK2+nsNZRm3G/Z2OMzW0o3Vj0n5+UizQnZsFUHhSocVzHOEA
8cgZrO+l6FG6upBx9t9HV4YfqQ14tOyKl4RlFkNYj4+9bALw12VqriKGmdlsj3mw5V6eZ/lba8GG
HQOUB4GX/Mf3zRSz4kL/dmp6m2s7JZxMrDFUOus7LT/mfaPPrtxfT5wmpIM0dKfzb0PTlFS2HxDb
hJGmz6cnYtgrOQIS7GA2fv7wcNXg7YnPNJM3gdYF0j8FqQ9rMsA7FRPYLxsCOu7h2CQlKSYiHBlh
iXKvHbCMEodxhmrsktsvKGvUy6W6DJfLUlLl9vpE5sWRLT07aAyqJalyz2l0bhj6JwZw93FG1haM
Ipsu8VfiX2wI/Akx7rWOpwK6I6Uc9s/VM8n9ht7pVjrcePwq883oTy2OKiuffhJQB0wCyZvX7E4e
9iwpl3C+wB/nXgRvNfV4AkTbJ+M5kvwzkdmnnlSkDwqIxuybqaHATQKFRcbhb+gVtdFFx5UZWKar
tmOv9mQtuKREce/P2xxWYmS1yMnQ5F8xX16k+bNEkFdWtH35yq2NzJ11/dENx7fND5JIyj/Dx/DR
R8TefPqcyHF1GAID1VmOpwhpc4gAheA6NmXAstqVU7FN4OV87HtEHGlvcRCyJ0mfcoH8ajhcp9ta
00kXq3sCP9ndiLjbpEwQbbNemXyB01mWa4h7FAVWmlpnJ6DeA0zgbX6Yk6nBSzB01DlT7iNlPuif
ioI7BEZ0/NpFO7/bJ5he+fI11dXnWQxCVlHSvkeFl4tw7jKltUe24WzRzdltRCHdZ8gZ7QPCk005
TSdIRBe7G3Ycv19F75JEza0HyGkHLwR4YnJ2NoD3cnspemK9ktHQzNvlvj/UO7J9lFAgoyN5F+ts
SQ0pTQpA5iBwYYPxOJaSd9q8IShuTEdfDFIG+NkkB7uqIZh9H1gg77W6VrZEpBG7BwbFt63RfIPb
bjkKpncCW1Nqd6GPmjQKpcfkA2z0QzCQR8CNiZxaMCM1Y06NOvlBmS7D8ydSfLsImVWdF6zvGUDC
UWAk+0DS7+d9An0YdxG292urKRINnqa6iq3qqePPLgina9jRD84JpaWq9Z1IhnLRFunXnQzfVMct
TDOCZeZW/4KPbSGBEc4C8C+NZa4H47WyBT8RMxqwDCMitC42UWpDFFr2PfM0G6bxXlbp1mZ00DD2
jsmsrpb6HCr4kvdKkFGbUhi2zV6KSljrAkzv7vFzFxeerR18aZLn+FChG6IbXfLiFLSkKi/txlX8
V8s8jsxxBEiDJpezs6RdJDvo54/XUUxXacrixPbbCVAUFxZNOfiIZZ5ymASGNKeCUNT0EauPKccZ
vF8tFlXLcCr8YIv9FezBRZw5lBdHje93yi7SAhkhMiWa6a+9NY8mmlu+WLOxlJtG2zWtkJ5kEZiq
p/VKCuy6mf3G1bdnvupzVmji5uSIOwoYveeSnv1VxOeE5yrKEN+k/GfwMutWBYQj6a7LPr2A409v
N8d+pHgtOCEI9YgV2j9QnEfPursuc3HRzsQbSu2qB4F9Qe9/G9liz6j43M+6yMWxZsnK1uOvB4T5
NuKXTcvtI9mD0sHMQWJEyFbJTziYkjpFV2UrtFZtQRjNzmf3pYjC0slsxwndmPh81YPHYhZkay2k
QTPBR1njbcNCbOWuHZkSNZHVBr1wUZ5ttDmIn4vppZHbeNjZyCOQG8x1K7gXK+EeTmgZnnDtKD2m
3uEnal+CHcsiubDkFwbEm01Z42sA0+Vdtbfu+C5N9IW0EpKrI6VjH/6X97Rx/a6gDrs3/bO8KSgU
lr+1sJTcW35/dmhkromoReizgxV0CVKd+lRszPUSEb8v6CWHQZx1+oXEHdLkWCN89fyJq6CTznpt
W3lISAIEhVGAbkD3oTrWN0gJJmKrVFip67XMPKFMe2FjBOWpFiJQg0yG7RBf3lqZhMK2hVCCirYF
QStj2U0wFdQb7zlaX0/f1yHw1E0W0foolcoW9BZ0zy8wEQnZu1pZx2wwBd7PsdzMo6nJvq9l/EOj
NzUD/nLnYqa2FLJC86bwX/f81vb5ITabh43uxawzXPicLITF47f5r8q6IliRhUTI6ae5apH/Ew0X
5DsvStXk0tUx1RWB4tYqcA2O3boU1QAHk1+X9/wohBrdTdZKVWNQXINAAdhjSg03fGKuqUrsi/ph
3hpv6yvkF8hjx/LzWFiNmn1ZhEogrwEbIpNBlxe5HQD86MXrISvcRILc8Tx+k5s2mkFsKkVeLauA
vZwbmt+/W9jIrY2ma9aVAdZjYaMg3w7ttL/VZJ8OZ+XwSge7db1ohcGXSdU9XabLuS6UTIuGsjXI
jJwMdcOqAUSpavbXTAfaLtkpkkRotZ7oDM4Er5abK6cvpVyOCs6vmw+/tX5vtPmwwJdh3iztGCIt
SdTD3wCRYbV6LIScoIcqTWjBo5trcD6ERjVNRH5TS8saeEEfimfhqyZJ0jkXsNdJW/+IdRpDwMJ7
DAGIQIhnQCRsVCgcQ+FRTHRvSCkX45aglb30rxP0D1LAU5OdPrHYVmFceortyhb7+R/6ZpCx9D9H
Sn891/tGj93We7CF55lS6mxy77HcUXNdOjp+RiAl6oEVH0GDxMfDRvvaq022QqyQ6iD++31ij0Wu
V87+Be8QT6tW8tJ9aRleBaE85s/yJYLHHxwt3CxN9vOrC7tdwqqyWwBcDMFM6jM7qnjOMcN20zpR
WQZZLqJIhSW5265NFhqjSUKolHnDzlfi/IWSBWTgPy4Wdjf5mv2YFdC84Ct4MPd/dSRFdfZX5fAM
OJJCVb12TTRFn1UhMOCLeRmxcAm5uY37AMcGRZvEiNn0ezZ60VGjpCRBf879FmFo38FPrlnS4DCH
bf2M8fvPxJXdXD++nJN9lZL3fFLxbsPOyGTiUFvGw5HX+TzGzs99fLT8tSekeMgsfKgtcOiX9vD3
sPeFRojc0C8vYel41KayV068rxaECbOrfMXsKoLLNcsxBDSflnab4k5n/0XoZbRhihImLQEDY7u8
N4Y13O85hk5nSZNYYkhrYVIifSQlHw+fw4C+aiRI4/y7d6domu62bozL8CGlD5UG75L/G93/uLQG
h1pHymfn5Qc9YkhT44H74FCRkwLRDtGVfL8CmEq+4P5ioJkQT1tVaLtajWltFzW7gTMr/IL7MzV9
/1eUOLrOnpPaTb9fhPhA6eSmNuRuXY8mBK4+Asx36sWzO9/gHZzQIrAlnl83zkLCT3tRY925XHEe
KvkGfzSBWUBxZxelVvSzoiTE5R58FoSpabYqMa2N5JG5WAiou3EYQnuy2rWWmFt7tiEJd7PR5Qfo
V5IFaE18zqy8Cmat3KTrrdrTz46HKIs9QkVbvQRSCZPdj+s1G3BY07zhNYIhJ/AARN56161D82Gs
+e+kmmZMxVfs2TOUN1t8lL82Sm9LDHsQw6oNG6VPHZHEKA8iQLO3k1E7MsNOTzvJcauwl+6zrw3W
zADHkrmC8NGo3NfFDFxHMPb7aEafR5kYsVYAaMqptuGCG2mi/lUj8MNtwfbBfiMWv3bycsNCaZ2T
asl5MsN5DQa48ipTs+RsDFUYbBhiU1KYL9Vbab9hLc4qcEOuZwXZCy4/UZ8Om0TXIN/ycU47LIcP
L8motHxWXmf+bjfhsf1/vo9p4icjw5D+FD9jEMa6UGb8+M4cjUdmmnN4qI/miJDfwlzGOq5FWmxq
MNxWWnUQoBo6b7NPE9Bbwhi4sdiFvJztWTlrIVMzDZ5mk1ZygIH8eHzr8qPJ0yKEmdYkCCwkGFwH
zaJNspa2iL/0uEe8tAV3P15B/+Tb9dgc4vrGlrdw4EOcWnakwXVwVMjekK9Mgi5NZIVxSJ6WauPn
fWdN+Jfiyj3xOLh1qEIqEwbBCbZG25mR4ahyYeSjNFBADLJrU/aQBJT5pMuxV4u8SCDY4t5pYRbb
AvAzfAnDTgiuPagdIML00FebiiqpuAkSWN0hIGrmuRHdCPssowBwHORUh/ZYsbG1D3kkfu9YdpkN
BhciwUO1HEw+vulghfBU9f8Zw83toe9LJQkOJn5PZNDbHBTaB7PXPbdl1FerjK+Li/bxNVxkUSuT
7hLiBNXmYpI6ZDlieIaYPQD6nZ4wS9zO3rTaWnsYR7l1U2FCyH4oBSRlY773+Ba/w5fMkYQiP28f
Yu1iPhS7dYCPplpeM6A5sy0BS6w5rW+N06pDQsQeTl79l9LmHE774CqwJCixaDTJ3QIvWBgDeFj8
XZtH8nELxJvJlIHiAg8ZgufoetnLOZNq+gbbGNue6zHIWjhoCbTu38oahpOfAIAT8/fhKXjkTLTh
TuGEcL7JdmyhIj1qplIell8MylhURjuJRnftc+GusP66wRULrfMq6K5VcqZvLabzJXS4or/WUEIr
hGkZPbdh2fJ+/Pj40znjzurFLsYKhpLFhr3zqlOR+R3fbm+IL7g6mAQudP56XecadMh2d7xP69ic
BVPP8uX0bk0iowBzOH+YmC34pfdBjOCzvzgXxexDbSxtuVuYxJ6owm28XLsD7nnU7YLI1gNZ2lfP
VUdXR4Ysa+T8FIy1M2h4eZmlh+2PYQUKiV+IjyGgXp7ep6hCZUvYmNLESDgd1pJd+Dk8jBjCU9t3
L6d1bfGiBv2hvd0nbNljPLbaiwzEMeqGB/qFO57wohOhDp98eCXz0ncaUbC+EBA2MN1QZtU/HzlL
QuGgy4Z/CHsW11YMkl6wZVdQ4BMwUMzotfYRswF+BFwG6hV2FuDuWpaeLDcFisH1P3QFn4Mqdvj0
HvJxA+K2F2XrkHl5rsnt21K+MhYpIGtfUJn88pjn1IeH+5oK1paQJEaFxUga3P+wAyxWmLdYjJJA
qFlXGP0WzXTs/xgLneTLJbI3phTz6BLk79GJBBYauV1KA7SZ2lAphPLUC5BJz7JOPZCUwPOwXeDF
FrEMzA4rTkVs2zWuuJB0Zb8LJs5ug5WOtswqONpvlkwxZCbNqfpxCYcyJBphYMv0cGwHVbKDpbQK
fkCt3AFuJrutNNIpDe54XEZB8g7YTkxnlp5BJPBDKgvEnPGIozFT+BOvl4e/Q/msqq3AyaWYQapD
e2lnXgNlSF2PKgfBRzTTy79CUz4lGi6xnH141KeLd+CKvDYMnfwFfXA8hFz4elGa79RiGBX0leZo
i1xdpByJKfPVymA9RVrOkFWqqDrs0m4qRciKT3EqEGgxuHWHlXWyBSjGEFax/cGUjF/POUxSL2y1
VRjCXhxi/KxXJdsqBeMhYM2IxCPN3t5te3Xlgrpcglzduq+gtMUXNcz8xzAstiQY/I0MPkfRJ75U
IH6i3elY4TTt9uaa5GKaorlfRe1A9jhmPmWxKbvn+809hujlkG5e+i/zbeYKWhjYbitb5mdzIN1M
nwkgdONM8UfJxfpeHaDimpQ8qbq1AFp1caPa8CZ3Fg+cc0yRA2ki/p7sjTKnWabqcz9Lstm7L8Uh
BwnkheY+1+ofjzfDEJMpjodkJCFYRxxncvtx0TMIMP55mGr+NskeT1tqwkoerWtuqedjtNB2QC19
LnO5ncLpOajKyrbM8q7QNAEk6FbMy3qlTASfEOz91VfykNFPZBBqQ/LE80tozx7Hi7P7+mbl5jUb
tQALRj4mZYvt6lq/+S/ELWGny+shiUOmIuWBGRDLfrQh78It+kMgP9WhpHRPiCAWbRomZ6mir5ga
qpu23x3EzRozIA3tDv0nDhHhC88tmVdh/7VD8+um+ZcJs9zMc676TxmxvzQ2/jGIdxd+Pf8JUYW1
rITpBMYMUKPuENVcc8oqlT8X07X4x2oBHGDJ6mfcD2L86ABd5ayBM4qitn8+bsQ6s/DckR7QF44b
A2iweKvYsHM6oNQ/lE4jitk452VKDFcsNgj0aX1ONNIU3KpZMLH7e1JUmHwh9fwuw4JobpxJSpaV
Dg7xb015zzWNediZyLN3+lgN5UBXyGCTUhFYXs1PoUZdycqQrlOBUotrqmBhyXFtld68/gRv3KOH
5FBsLvnutvub7T11ZZDmpVK7sg77n32hpWruQm8dz9L5CGwTa3Aqcg4m0b0kE9a2GVODQB7GPl5/
6VlTm3ftlGp9y2nAydWt12o2Umzay2NzbH+hly8+0ATg2aftxnDd6GtLGnmMxWr+f5k17xC+SI5c
AI8kg3cGD0eAL0VvvV0Ftk+8oUJAieNI4Us/4L4YVys1n/hRFksP6iCF6o9pox4TZtPkkbexh3rV
tGIl6wZejPQIMre3m4TZaNu/cr3vKUi1gbNkoMfgts5+TqtfJnNy+7ESkU7Ck+fgEI0tk9VaQqv/
8scEtRGy1PD3kNKwKsdVqlM+X3yn/w4odkQS3Wdtt6nX92WHGNpu4dm9dqVxa8wCU8gq/z/mZdWP
/DovEQDXRIrUUBV6TvqLFKVvbb6rXdSMwo6DKqh8e5b4IHQppdjMeJSnhyCaHMGwN0qUEKBylIpk
k7kxnliF5KTVr5RkUEWi8TprQDLvkVJgM7DI9EzsAJDhfR0zelXGKMtZTgQ1psT6JquYM0OW1exU
ojWFTF490h3QuGoAKqD0rvZ1fMtQrBR/GEdSzZ3vOJPcqu9TjG5IJijQbkJr/IzY6ScjHpyZZAq5
iTPS6891dGCLOXTCji1sY1j0xP2XBW95NFUqHiSbv/IZ9oyJYDMigBxOrimMCQ9p4Y6fJgmlRiXg
mX1OBcg3XmC7i9GJHky4ig8Ca1xrb/UbMkU7PQZiit8VmHdAjaQtpG7P/DYIS8YVd2pHLC+vdECO
TbdgObotVotDbtKPJwk11PBcvZJJGrbKrjw6dJ3R2DCb8bdEywlHOwypjL4d5EFUvzXmLzmDyi2W
31hdZHjr2COKjPxd3Zdrr/qIkmbuFOGJXNajpK2dUYPnMahmecFhCEjRisriZHzez5Wyzcbcnrxh
pcJY9Cju0Odlh46CXXF3La4gPSDzGF2esgIBGxqGrBOUK3aDC9N6IsWb54g5lm8hNdZaLIPvz3kn
ZvoyVz7BhPAusck4hibOgRu6sEJ2Grp5gQvPgRIiNJd80THGnT+r/GXVHyEMKjFZHRSMrdxco+mL
kFWFu6GTx5FuD1f7Rfa+M40AnGLIgjhh0crA93hxVGw6jZhBzLQcYOd2NyzIBK741l7kYqchKP2a
avFAGTd35OzF+uadS7B2UVsQgtyo9QTNzpbZ/5Le3i9sNsOrad1YtkPgVo8F90lCZcmktp7nfRpk
gVzmBYhgu1qbSr3v6IgyZgEm8t5psvm2Lp8l/N6/hvQyFpVl0l/WzuL45P6ux9AkMk9s/D/wbTU3
6hlL29LE7xH48WwbHq0rXQhxs7D0MXL0njk6QCVoi1eXmuiNphoy++w+bGKCc062Ul4tpdaX3v5T
/PT/wRcq/lCa6vTruvhMJDXRphKh8E5zLnbqPs3qK5cqFeUrVAupn8dW6tnaDuwNlKMFeJbGx1IH
meMpEiuVdYh0E1gNHBzlCzChSJ7rnBFw+C0L4Vb82LPjgLlzAMTlA8owppMaWH4B8WLMmYpSTKYB
zCcBikELJ3WG0mc+9iYMVfpIqXCfxKB3RKs/xDSpPWDfHpR7Gcr0TCCFh40xEcIOy4hElog2TzNJ
ACgwGORkunXQDOLmkj4zjgW4A/TRZbIMrYEi6djcEB8MFo0ec+iqtyhaltw20AIUifLVsMQkJnkY
yp/yPl11uxMEDDO+OAozUF5YZ75nh0b8/B5bxJMgelscw9rFL/+kNYPAGPszrN3vdp7SsZhmggyG
1BanteBHMeXNkLYZlH52VD71wxWq+I7TcuK9d8e/yrwxZ+gIReCPvcqVLe/Wg2kkQzYP0RZbNm/v
qtOTYn0ngDvt5MZ0hK9HzY6L6gScXxAj0g4faXJ/vUf+FVyynTdhMisuuxFYl/PyMPGB9jcrMj0r
oQQhBikuHxdnlxCbZLUp1l1p4YK+81Jj32gCBojFErLBK+MMjAyZFxC3EAsEaLwouIZFKgD1rYjZ
aya/XTNb3J/sVYUSknx09TaAKV5+kDfcqUcf9dpSlbqW2gQc/UA523sjjBC0ECLpaEtYmhNwohaU
C3B7ze1DZEji6t367K0qp5uT3lNE89pLvu/On7J5jMrmjvy+CLGRUq9HMjVNJx/Vn5tX4cka/IYT
wLDvwYbk4GVzy/ZBpGGaHM6m5qT9V/hbdW9J9NC6cqxbEDm4hubWpY/+wdo3t3jjHYucEasQGLVn
lMDVXLL16VQ0L6869TQByrRASqX1DSBV0bDFErw8kYSYWWG+6/b55J10sTzdTCgQnFA+kyj9g6gf
bO8fG21xWbkI2bd2d35sK7iQJ6j0vvAr1ccJHq1xjKR6Rz6ZofNJBCWopYLoOg0JJ7drGn6UdSEx
E6hVHgWqwJ2IA79QlRV6StuMIwtsq57KBtKoNJvmPAdC/o453w3iRP9Y1Aw9Xl2vaZCXXbcutEp3
wJ+9IZaahD0TbhdvZ5ScM3wm8+v7u5r4hdLiGzPn1AGfq7cPBur7KEdLUVv2lCf0aa/GZBMcHLYu
V1lV9Le/Nvjd6Fth3223kSEb26mLScAV8KRjeKWGfMNyf5Y298FO6AWGs2qI+9Cp29Lhu4TX/T9l
ToDkeN2rVQrYWHmnw6Xbis6TCw5rpj6GP1wQsiVVYwPM8iJCs3N9+e2B3XHb0PCxobGppl88JSUP
+Vq9O9d9lQd+Oae1yp3IQCGYxxaGcqGnFyLeyBD/P9dm/HCMroN8fREDae8P+fAoh1uKNRLjh53B
AOYot0OXoaP/JpSwN0Q7CT0QW6u4Fk6BDCAnQDxDuDFYYVaZ2R2rtUffsidpHvTvsJx/a1Md58o5
rePngjIHnfeqoAkfAhGMlpcDe/CktStI+V9sbIcuaysal7T77n3+FXt0Nn/0KYPmD6H0vmUpkDXU
tmmjigzF4z8qq70oIkU8LqGrXCu4kCzzzIdDYwfwAeCiS84HGm2e8e9c0Zy4OIvTayw9UEGn8obI
ev7Bdd1v54EKA8ihg+JOxTbLfmDJ17y3uJhGQpAGz4YeG4o+JWw8PunpoebYts15fxGzl0sdnbE8
pxggRvG6ulYYVeC71bajEYPQ79YGauXAJcXI6AIifS5O4oq9aQZvSKd2mVfjqdjYLbRKo9pUCXI0
v+oGIGh6lFLGTc03PMmKb04Gfz1UW27fcTfXLm/ixeF1Bs4XxRahXPso467p9IH9OznVb4wZ7hxi
LJ3Frxe60y3DMcYdrouxFB1KpeWBn79GCBFOjoC+Uigb/StrKyRvbX44Gb+196cuvMFHHjdAsD77
cxU6rN9wyeFCRYEm9EkCRYAByVfVJG3OchcR0c+j0ZX3LrAGUwhc+GMT6fnjFEFaqyWyVtfMv0QW
npvwhS/UNmCdmc9BKOVP7RLYeIUR/IQBBjnEAts/hVD+q1DsH7mQFC9+HTa6YztKxqyWIuzRXD17
CcIzwFMhz2IFycb5A3s+Hfwid7tOTttiPSlWc0ZqWz7FdzWD31t/5/E9vQB1fk4l3PfQ9Qgs9cVv
HAKNsXJRhMy43USe20/cmx6VRtCf6DcSX1OdF9LIcJYJ2vuDr5vjcKSi9FkfDVtECJD7IMLZ0k3R
Tce/9qNf+LWJj4gpbMatInWERP34u+jg2yrYJmECYBaAydrc/KWDxi6Hc0aQubrRnY6tt/f7ORWV
AqiK135ke2bK2r+ltfERvoMfwdUky04Zwa+VESDpQZklO9Jm7Gi0aM9JDgF3xLxKQULKN4V+BMf+
asu7CQ8NU0fJY//zA8SkIWOd0ZEPMhwiXhBy2lJS9T90K3Qyh9v0687w7t/Epc6s0AhnDzgkS8u5
Uk3TS/a4b+j9DoRZsxoSe2GRk61l7a/9ixYz1/M0QeFqv0Zj0HKXNc7NijP0NY/my2R4zJu2i0Dc
TH5Q2KtEvln1aNkEpTqBA8PmhM1Nvl7sK5L8t2pDks+FYSaYMZXiGGS/1ipyMt+8iXKx4yEv2bsI
EljZRA0WCfoQWY9Wgi/wXCQ+4C4d7M7HOyf7smkmLBjf+XT+qKaT6kkKRwKBIXHsXxRCZE4tQBBr
HoAYBwPJMwGLJQfI/8kC7KE3Lc6YjxKU8OIHVUH0qAC0KGd0ZVAEWBHrZz61LP8u+9f4Dw+WLU/D
WiE4p/JuHLwzOKqCoJaJFB45K3EAi/XO3tIXiLaRMBS9Vz5WngNp3D6+2WNLRjvl0v83honnjUAZ
+amtmB2iI9SJbiQ8tyB1ulZYlMkDH6Rf4xMM49TrRMVY9Lauu5LmmB7dyx4r4wbkSf3/g7MTza02
AvaW4fxh3I+/onG2bysv96dZFAg2x/eMbrNNy3weyNbIWtLQ1d9T5U8hF8uXQeRQrFXzIq0bLCPd
4HhnMQkYADryS8Wu2v+4tOoFTDQQ355iUthna4ToJLR19uRIzNbLmyuG8hs1brcy2oVulEJIh22n
sGcACiOlpXE/IzlWM0tfs7Enpk/8GMD3fisAhxPCeWTm8Ddw4iSnEb2xkj5SVPHNeZRs/Kmch+/X
EINld3V1q9u2i4ndxE9gh8MutuFSmGQK2yzl5A1TuiQNBdg94LsMchTavr/3OU7XnrOLpRw+7rvN
WaPru/SpnMimgFHxSih11oApwo9iYdXAqJYt29HZmQ2NHZWZWMCtJhTyE1KUj/p4NzszkdYm5j8v
xL9/lVEuCBciNLOrAYI7xuQ+UAk01rX3grv1esJ482CGfwt7kn9/jkGrMOEr2xQV9Jg/GUu3c/P7
bN/IsbmyoWOE3jN2GcF65l4W6MR3dDpzntN8gFX0zK4hp2C0Mb3X1vZgrWBk+O/DtSHAwfRxAXgu
sXV8tKmeZTKuVmfhLzJL+CnlWIO/gTTLeQ1/ORuVU+2NnYW8ikMl7TTZrqnrMncKTUxsvNlpXfHC
Cod0xUjMR2X+F7HOhgG7WTscK6VDJZZCTPtuX13RypX+z5T6uS1wffsIlIZRVIf6GhSnQVCFQJvh
Nrrn6CXj1EIxYxBj4sjVFcWrzHjoausTLctmUKv/dqghUJqshlJFM/t/5JGMeib0uoaUA1SD3TKI
Fqmwn5ybuvMkEFSIHAaSCfOhcBQMgXwkthu8R+Dw3y4IdUo4s+EfeabI9F2XVYXZz/vyQ9ARf6+v
CIBotDW+rcJUAwYiuQePhrybyiHcqA8ktjHib45vse0XJq2LStoPgYIBIBTYPmUDFIf+QsSjDSBr
cOtUX2c940NOaXYrrwLxDQ9BU05OQs2xcDHBBd1I9A5kzolfyoWPZWIV5EhwSu+X768Q37DlmG7a
cn/GC3jwGSH83XdIrUixJlKN+WdC4O6NC890tg16gEeQDBYlKgzh9+oTMpPcU8yKMU2F1lA01CHe
Q/vaOlcU2CV2fAF4zzx1S48nH07mdXOrqA95jO/iHzqN4pZQlc+PZbZb80XfmKhDVF1uLUqhVt1x
iqxt9Pnh75sJcBDmqSdEEn8NfRador+oTgCmGXx1GzMyWDUln+yAq5zXX5mXBH0a2hCAJhWHxqCT
5Jl5UPq3WAzafWACfncxjpRmB4gMoq5wtHlq4sr9Jw57234pbyGjCEa26eg00K4fnMpdA5G22kql
cJ/uqIEmgWzLwblq9vF+OYLrn7EVMdTkVNjB3bZ0aRqN9i3iuJ6CA+6ONaAl/mWADLDXbIcxC9ob
ZChnfRyEiavs+cJxdNznoKkA+vcae8nP9UeZip3mOjX7PH1R+2UQks/bP9Gwr1zpWYNbFLL1ruYR
BvlOp+aUPAelaWBuc3PH4Fun5HmD7rWomp+hYfgEU0AsqpxgDPfGn/SmgnNBzuAs3P6FvLDKU32H
2umbawdLlsrp1gUoW1NpYNx9xEG2KXweKpd/H4OmILqp9agSmJXGtG+ZzPCHQ8gf1aqOT+8Vm4o8
K8or/kCbE306BsRlDRXWlVg0nnvLd9qyTRC/AX8lQTHhxP2MUGCwCNN0S14vVRhR+VIa6uUyFmQR
BhWZS8kRoGSQBihch4VcaAvpWZlf0JHY4iKdtRmUhk7PglekwceTxebHR8R24yGij7WxFdG2Usxu
V39qvY+yk+9klI+VNdp84qZnSz/cnSHiBWe2fvl9cxPdIzslL4zOKdPZWrdWspGrQvftGnB9qWl1
sjH/CoqgUzvDp3A/bwxJHpO2wKpzYhDU9gcHTBcm8t6zuh+jwR6xHMyIxkGk2Vc5kRt9Ro+5tKRS
IhxbqhRCBYR1ksH48NE+FXxMEydbU6cI5uAF+Iek2uFTEwQh2eIAwLADs8235OfksGReoabvtego
eTaQ+dC4LeJSUI9rNfrnUQzX2KWWhI6ZNFPGWkOvjIMEKzuJGbVKXUjrgsuLvZJE32Jm7wW2T0Yt
ZY+hg+WhC1qDXph7rw/8TNix5Sn8K05rcNv4AIyEksS82Oaq972/iIQneJEvSXQKe/vHA2k7YM3D
ME+QaXWJHY3DhZPD/KNz1DBGt8FgPM076Ai1bQJIm6AmbxgigcnrvrKYYOJbHOPV+QRpRVpxVHLH
49CgYJGk7G2Laanw9oEkeUCOuEuUcdGvuK869InXmctWHC7XW7fI1Lb6IAD+yVyXdEZrQkDapDQ5
Wm8Woja0Pda4J2/jYo5y0UY7/WFNtt3U0PZPIKggwxqZu8gZjBJZkJiTnvcZ1CIm2a3UQs3FeUqp
rc7aGJOPyIzr2zmYOjaW6zIaxIqnLIsKFCcTmE0nTy46hm2fli6e0R6uzUHnKEwELxekkCOgq3fY
Oytt3vfjTSmUmEsyJuSgi7Z0UzFpiiqlU6xqkuuUGpJUuwW9UoSWcVxFo6UVjNxANgu204knbuI2
SAczVIT+4/39vmT9zVUxO74IFgba0hLXbPwnAJx6qonaDL85RUA+kkEhAAZh3ToOHr+PgNB6RaB1
wbKia63hz5b9OJo4NRtKz7kQW7z80bWm7iI2AVKQna0uKI6OGZqjdM462fbf5HqeBT46nDHwu+m/
yOXnd8oR/rMW7le1PsFtwTkCFZ0VPEe/LCSom5oMeE1yxwHgls6vTE1E7WfXCnevWd2yM1Trc9ua
bI4Dm3oFb/YFmk50s4ifrEX0UGGlx3ZYAXz1I1WPZmXOCqo9UKda42gp02+sxapkeZRhuC1YH0xy
Z+6xtsiUhBb9+D/5MQlwglgccT89UP70/ZZK3wl/OzZsuoPfPYeOK8nBhbvzGbDM8uQaFLwoVln5
AoKSC+Srs/u8X4jxwiSlVpEjZGFM0OfXgBLodEDWacnhxUvQuwl3mYU/XmRgOjGm/xWceYAnq73s
Makn5OWF/tTXYIElseirp6d8+C2Dlzbe9JOESByXInAvzTmVr84Vvt7H5FAYJ62YLxXHcWHL2i/a
Fk8/9Ih09QWy8Yvm0IvqRbr5d6Da3dGaDIEasXsZYRAZv41brmC6RqEoEJtz78ocdeYKrSyqqOM0
XM4jIr5Cxw0EVOOOGkDare3gb2NX6UGReHah2esN43wft4v8ZU8iLF2PO6QZzde/Kb02dVk9t+U2
o24yvJqOphWVJv6GVVW2EfJ6zw5VG8s3NaV+R0JiibQeinhnOct5q+3txYL7hA1wL7TXiv5P63Xh
/G9rbPG14/Am4T8k39Ve3794q+4g6FhOQAyEBluUgN8IAHmt/ljgRPw5ebO/E1+08t5V0n0kdIjz
osl6/il6rkPlbAMyjFWU8/PDe2ODhcE1Omh9P1m0A5kbjpY1kMrzFfb1BpsI8+yvx0FiGM3LFa5m
/7gxecVg3vXhqozap6pFPadGGNPjzFplMfIS4RBWVp6Dwi3iyPRiU8CItf8FS04i9b6qhqub+ZLD
PyNAxokngqK9pY17M+jCGoHt7yo0TrLSFTmTd3XWoW+R0khIbpI1oLu6zqdMLhP+rHBhDlHO9yNW
MACPhmIfpVRCElY/UhPRvmxJ7o+hZSNsPqEm0LivtL6ADQVaLHT8Z69InvFBdq35e/HVEyH8efVR
HYiCHXiT/m030xMxmEzPtiFqfBu8nASby2tCKuJump9nXitq1AvgYS3MlSRNvfj4nWamtAMBjwUN
ZtyQ4oOGSzgO3UuvUubvfWeptvOHcLpZIxcFJ67K1TN0IGxTjngzA/MMUj7AV7Q53uWTFur2YpQ5
BOgl04iPV0Dnq8Q811/ilQ3FQcj0IZrCxrh+zm2GF7d2LFrRusmZbyFWZHUU6x1j2h5Mda8CRahs
vEx5J+xNpyjqNgmY09j04djzlZ8ksWdrQyvx5S69Z7ymp3dUQQPCpVUC+c+Lr5E9yc9X9dKfCKIp
k5BBL9IJSkeOe4ju8aA46s3rXanJphZecIfQWZD7a6X3IVXHu1M/s33lUW9BVEbYdcqOZ5fIiBVN
3hvwGwRVvtwc5Pm2X+AhqSZq5pxb6s+m+U3+Fo4YNyX3KkmSDxsnvVEIDZ3ib/p9omXz6SDPwCEo
0MjyVzUvfcHdnaQKiv4J02mgajx4frS96pxJfVDBLY+NgyH2eDBGr2KXXX6aYibffmblTaCI0ytg
xjI/z55dqPx1hPHTEcvx9EUw56tVGeLqRX1ruElP1ir0FeERWJayN7iEsf/X49+vMpc4zRssY9Gl
cXWwoiNPj07miJtW+Gvk7LmgpcE7zNyJ6SKmKBSdgVsRhhAiu0JCDqiqa1m95+KTGNIssiPieB2D
sTgkhARRrxDFyczug/L98XftNgM24tpD7Juszij1RhY/75NDPAhjxIV/cwAkk5iNQV/d132rZdPJ
sKwnb9rRv6cXazlJruVm9D8bhh88oaYapMkKuc7WIeK6luWdSYO4wtH87CDXYx4Tr9ef5X4IODjK
CCY+w5tgg08cLxX4u88rM/g+HZyMebTpAoArVcNju+IqlJSV3r+K2Om2/a6qqfCj09qKLWlUnLKl
VUb3Ov8EHSYakj2CPUzth7zfD9gfoVVrX2k2i1cLlTPHHCxZGnFKJ1juJzdh7fGPbAZ/rUin1R+J
MxCEm3USkvTLoyvJJce+UhIfZBPLbY+hti9zPNpKJMqwBhBNYs6xwa689JEvsF896hbGdY/jyCnq
pkgqyn8rkmYrjcGuqpHyW2L3CTltVSHFNfOTU0ZHKzRBf4AZ74xbAazp0pcJC7jxlU0UbBWOSf+l
zbmws5exP6y4qJ11z6CPt78RcUiVlqJXHCBdOzy4JROKA1NJCQ5IEec4B3h2zz1WNvjX2mLq/McI
dcs7bfOFoCUrn+cRV69y3TZodgkMUB144hqqsQqIebxHZn85r187BN+8vSJwDZBsX4RwePIVel0v
7ktnd5M8U6EzWDEaX3rZleEqfvSECiW49Vkz4jJF9w5SkBldJrgJGgV2VSds1xVqOEg5Ia8ZwlMV
rWJgEZbplBPvlabTtmdQOJ7KQKa8Dw+SXyLdAH4t++dXPLQPJh5MRRbVL4Axpdkr1hchCDC1E8xM
97r7Tgu6+JOuOd8PMgfApBdo/IDxDhQnpNtAFuxM+wrsjRT2DtNUlX9lu97n8xlC+UebTy8Ay5at
tlbowe00qanJeMrVK4dVM8IoODh4zQOdocorPz1oRBcias1usjSOliHRDYwC4cyL0CgQD1QrpEpt
tUWQL+biX4tZuPheVlHNp7WVdfylIurBUtm9Ao0Qc97rFLWOfwi4c4zQlznvwhB7WQYJsI7v1fP3
ofjz/e7Oy3LExTf5CSnHLIeLSyiiE9Us5TO/h/w2SzbhFAqN9R9N/jJ2MMFdqXIT3bL++ptnW8MR
5xJ9TeyKdWx3EzydP7HzbZP/ZLXJx2x2SeduEhW14LYRGwGV8/bD0G61/JqNP9fD8InzM7wgMmdo
rWIcfe4U/td3aZf3PbatXS+r9XEkpaD+xfLZxCgVh5PS5Fneq2kheyyJESlPjdgA6sbmNqy8uwRo
vnX3oLQ52CRhND9KwWN501hbLyiMki5/9Sfq3bBTqFAC8v2dcqH5x9/PFpe/PLia8N2YrEt0DvYX
jFa4oZVG57n1Z/11TNzRRhIp6+6jtr3p3eNiPJro9QyxUypYkM3EqxfdsXELxijQbwFYriNvlomb
VzE8lJUvpevoSwSTOrUl/e+rTzi2TXVq8PG0vUXZZPe7Xn99tJPEGso6q5E312YPhby3y6epnKU/
s/nFb5Wy3hv2wv6Afdv9E18o3RbjkjBXsRvpaq7aI92NKQS16v7Nmay+6DAld6Ie+DrKZgjIfoT3
e7mporo9oQcVizDbCRIfehFbkLS0iychsFSl3waOi+AG1H4NxukCVqvUKbmwYWjg1pf0VCp3tqhP
cTL6nYOgtJ1pWNCfXxK6SlGSiEWFKF63VpFy7f2NRcFDjYhguNyX8fbJOKyP/xLeeyM2kN/SmYjc
iVC228/9k2n+zG2N0E1ODTchymthEZlQC+fqA/BGokneqp7dsE/WdkhJ12R5zRFuE2Rc2fnVWtBZ
LU6Q2AtYvr3D1xl1KwXnBfz73jRIToPTBrxXNPu4DvVWbePs8Y6mokPlpCy6zp4YH0eVj07y5r4z
kxMHgLKCPYUzqHjYEzdOpRd/NM4sWeg8SKpBhb5JaS+AYt1uliD6LRnFu4KoIhrCqPQIav5LEh5E
A5thZgUjQWJzGl2r3G03H7NgOel81UACTkYMyy+I7GtaiHOrTMcv1ymjtqqKXi40VRfC3FQ0EFCT
LjNprm0p8Z5DG2Pw7UgxntHwTC6hsqpH5QjYYgTmK+U/sgkA0fuYyLQUR324ePdZDDd3NT/dT8qb
tx/tduwoaTV1AWiRWWz168NSRqCVxgFFdrins50aVeeC7dzqK22JoJbTrKykGnH/HEokD81pwNVk
ClWEPn8p1zIcP+mmiPsbWsK1g6nkLAVV85a4nwbYNmiR9uXSgZEPEP/KJugEZazx1ddFEF7+8Pwy
O+ipuE9QfrD+kB4aDnPEtv8las8/6u+Ps6o9e9xFPQ2qac0e87rsxXzlsf1ViNQztewmGEawuEOl
9z37v+GsBGpwFTs2sDzjVYYOW6WezLghwPEsTUu82IYPGyjCz/GfbHolFbLrz3Xz0AgXowSsUWZO
4ISG0LKXVP4uL3Ql/LyHdzNuxJZoCBaJ+c2aBn1JNqJh7e2cgZNSODsFV8Q+8Uw9NuME1buqiWiz
iMeOOJ8wFlriMGiYk71MEZDO+4kfJfJkBxmt00ZTKUHOQ8i7E7T85glWOveV+dEPAkcEiZrmkvLx
YXkqN0Z/LiO/aMuA6VMcp5MRZhDqL52FkZMQ2Qhxffg9GE5IL7y9K+0TwfaL/yqJR+4arrQVHlO6
gSHZ/ygsLvLw8hL0/+cSY1SjhjfJJ7THgtuS000AA04UCKA87fSlkwyhsZ06BxTkGjoIUuOnbes6
wRzGP8bSeGCCB6JIHeadcc9gLIz/EYfRyWm+G92XoaXg+xia0U439z+Szx9AaoCCR6OOtcpDFPbC
YKDwiNs97V2E6HK5jLqEOIeGLfsrQPMOM9cZtF9sF6hW9survmwk+Ji3ryQ2Nq3gRauVdrkOyq+w
iVnDAjZGxgmzBpzOcpcDlnLhJtbYR3T8BBi1Z4LOO8oT3akYqNHGZPgmW/QwQmjVprObQ8rxyxk+
H8oUDAWDFQctXwatFU4fv062t29hZhQkX+1WucI47biAvw0oE3OQhdQlfBF1cRjBLZbgGcbylmnV
ME2a1YqaJFmJpV4bHh7pGGk9LO09YUwOUJpKkZ/7zY9o0mL8fHKdAyXw7nIYwL4Rij9TMRf3kp0C
awi4+yEtfWs9R6MQ3aOFqrhAOkFxYywFY/WnsU/MGRCqkNnKauKsatrnIcc/7LJp3a9O0uqggUdS
atkdxXHsRnWPVwNbRpWLcUaosGiWbcGlzgUUhVdIVjfe1tDgpQelI7s2fBw2DoBILx+zxwHTHphN
pLyn5L0Nsj3yhEYWEhPsva7/4jR0Ja5dy+kdzeyav7mBHEPMi9Feucn+AbqRo8F0gKA6mUgr9+TM
6yT0rFVQI1Juf4g4Cfhot+nTKQC0BoIsYFLut5x2arLIPckM1PlGxYFnJYRXQLOeM6X6xgKDs9Li
ysaj+qoeO7+4u139vfybcRl61+GALhn0uQmmSQ37izVSa2SioEXkiXeLGJYhuamabBdMlRXx27K8
o5vDtfj5vjC2UqkmWShp7D1weHiPCzK2yx3T4YBzxgvYr/Nkh+pBSuDT254Kz93DJeCtitjKF1aC
HSYGAeMB+NMHwamf7+Xs6lVU2neMGWzcj6bySLqh14RKUE8TW725AMooeJSXw99LuB+HgdZ/0zOc
8nax9OVW6QWhFVOCLV5l2NLnp1qrwzv5fSoJBuom+4zJbAzV33SGUA2jZVF1P8TsyFOZZTlQ1gJH
gBN+2PaG9PB6Pju/uH/RywxjGcBB/tvd3b5G/Ge7aJNs4E5IX/iKeEmgKItRnAS2FQ5Vs2Q48w2O
uab6r6VhurWAgmu++FmHo+JQVcWL06mG6yGIAGJlenwhRX9ISsszP2aacOrSx8gq7tUFibPxK/tA
hQrY1eom0tUZhUlki4w/QEZ2SA7GegLPWKhlNGng5GsXPcnKip/wS3JWUI9oXnf9ST/pTZQJXCkZ
DvtAxg8OUHg2UA+s1/3SGKUrTWQCxN1wBpPYonlwY83ybPrKGOuJVYR+de+BHoWS5SVs2dj/J3QC
TEyg3grdOaF00DYz8UmyFBwr9Sv4JDdcbblDpuZo/+RuHLsYC3u5ZrvKSe0agrFVnqKhw2bR3/X0
o1p7ordF32gS5wPrIKXBpknNa+M+h8A9WhmjnZIzsIlpHSQhmn3Ajl3PMqMLSlNvfZvNoeyI3P0Q
BkFx3mA8mM0EDgJ8gyhbuPdRp9xNXCZbR5eHjB64RIB/E7cvEqJ2/vrvYSA6ZR12AdqUE9Fc8R/L
mAO3PEG3OlB17MezCD+G4Ah7BUIvxHZfle9KbjKoQPnbRcSKDtEah7IpjFj1qFYAmzR2o2C2+PWB
iP9XKQJy45IU/i5q4c3QmewZsnkoLaF+yCcZ4BlyxSkIsYNW3UAlZmUkVjbLu1huOHjpFSHNv1OB
IAPKhPHnGDD5qafFxVnZPhnh5RpYvVwQfTPShawbnHwQOCVUcIKXsn4bu0HzpIioJ+oOZVOxHxXY
0D9SokyuG32/VHLp8PvRkanwrKVkhCOuWkSCvfuwRJzcMhqFHJbreXbbVbIvwp6/j52hzfAUqRe3
rhV6uj1lSjBHLDYmN2inaUM9phwbmGkRQ9fHEAK9vPtpDgqkuvFWWHLBjzRj0rldXfcOIKaYo+NM
i2RQZLdmSS8hYD3woKqWd8+ajoyYnOSzt/QPHhSFV1da1bu8hiPuqmPlfZ9KXdacJCTw8ixuvZmj
0kw1C870kfn9YFHPlH3E0FVRoNDlMMgsVoqbEcdGNuuGfaGSxSg3pR22XoDhsaXzWmhsczf72lSD
QIANRPxKOqDGsxoFeCnETUerr4WdG3aBLvbcOM50gtflZMgcN4AcuAJOmu0Dc1VnKQpaqqGl8r6m
aQIybQtza9VsUqSc2jnBWNXklfw1vCkbONvyxFw9yiGtiPFjr/cGRSeWJoMnm/segVP46MAbA9Df
U2LXxEOeeW3m0j4cCbC1PBN48YEd7Q49pTt61W5aFfdi1AxTTJra7KVCfOCO+79wcpbbiXjM/Waw
Y0kO1RHws9Tq3w/UOKHEckSl1tfIFNbJGmhDw8kQLWIgKlWj1KyDCez0jTzL7ap/FWjjEXWyD8ra
qVrAZ3E8NYu6YTC+C56zoKWH71fm6pROU2jxx6pDRDsAwTz/nXButxWxSFnS0nXQhwbrVhzakwf6
+UgmC07G+UlzbhO3PZVWpEZq45UPYayaFPtVjN2B9XFdzWS/VMiJxL9YEmCi9CBHoZq7P5Kz6+xp
gleQAtEN4zYFtqC49cTClhfKAY4GeJ7eerhdbZ3miMPZzc1z9Bo+Ua2pkzGWeH8DMnn4n8sd5cgZ
AI/MdvdLbeBa09getG1k+1hJB5+/EZJq2FgCTAbYsOSVjSczhRvLEMVR4vpfrNCX27j0JqkpRWFw
4YryJIZiWf/jGmE9O7aj5n1Qs/pbYmDI3CaS+aZ3PTGsiGI1Lk6E/nH+CanrXKhqNunxt3R6gbNn
biMqUY+RPzilEk7hOp314KLuZW6YvuXKZvaMPoAMihMfmOfpeNZAxIRvPoAfx1VLq3sl7+Puo3nu
qZ74efAUzSqghtxjbAQR1nvKks96e8UWk5T+9VzG/nXXte+JY5rTxxtK0yrIMwqpZGQCuSE9iTcQ
RVVZeXbgfbW7nL30CdfC0nF0RUAswFh/KwACzgMm5caQCqO7tNCdTxwHJSM51+IjXPMLRjTEBL2A
mW0Bgb6piugjETF8B03regE/9TAmMBDQ3Ze7pQZQE6gPZlhdHeYjmZnxALEOQ4mrXlzDfpJrv3xL
4amisZgA1bryjd1i/tGoT+sgp+XeINOzN3gNUVtiNmdqqE2s6NwLbRpkQMbN5srkxe1QtcbLfoK+
+AhJi4CWKyB+dWUMcYhXAriyIGDVTiK6bkoGYEo9LisAqKG+EI8Bx404lShMTXgU3ZYWHBfoUliJ
StxEQdusx4OSnlKNyNLC+dc26lUB7Biq0LCJzZ3zeUkP3vTmIQc3dsfUs+UMpMNWdtvUHiS6VoMI
iDMGggUE3gMn8qZNlIE8cy+nAAlO3WxbMR79LVc0hnPmS3QD5rlSc2Ae966yGmaDQOjkKtLOUZ7r
J0cU4DDTF73Of1Lef76//hJsFiOa3JC+G/WRu4RpKjrGo01H59/Qc9bY65/yGJNrv4YNYpZryCuv
QTfLsL2+bjERaJxVDVmsVs1ppL9zSyLykPQ++/dPnQlFP2AkNgKQXR/GJcD9msX/7uOP/1SpFNOy
uKzaeU/ac6cGcjxeaOviDGziNHKdAmAxZ9OJZ/5bmLKH8un3R43kwMkpr+6k9COzoXW4z038iN0j
vgk02IPm6e/uxyISW4jJy0VM5ZbPQ1wx4+1rxZUqe+9geshCcXnoh9NkZhvj8BdR4YQa4nJf3X71
h3AKjt0EAkZttK1Mw8LNgIz/Vss4ABd+yNvlzSH/ru5ZXWagGernS+x54B5mMDP7y56nRgU0UjZk
ojlmCHtU2AJd8AH11i4n6z26AVjskjcdfSv43nN7nmvrHIimGPoyTOGSv/RU/YYbtdhqf5CkW0ac
dBcyiEyxIJlJ5OLqAqZKTIKN4xqlnNIF2zTEc8uyrELwHt6+wzFyrDKE0TI/AM4N2uYsHaUCW4SG
D3QIaRi7+R9QxVCFBNC4RdlOzYtzrUShU8r46AN2WYefbS6JqJ1MyJAajK3Jt1TqDdphH9BUhHWd
w47iNtx7t5ae3buVbqQHcv48sNrQ9vR27AQCQl8iOCb1zZ+/g5l9EXFq4K4XsRkulApZLLQwAeNV
pphMsW5UscmbBzYfNHonxAthcx9hSfvUNckgPXnU67+Zjgy5yMvEZl7BCiEbFTcM6yyJFE/397VG
qnkY5DsZPpTtuoxy7auZNHlXh60K2i4eQJlk3Engw7RfIiyjxW+WuxuNRuIEwJfZSiyVtLkXEYJH
PIOE7Mc6USqyWdXNkfxL9Tjy+KFXl1Zcpo1g0QFSJ7V96wXjVLopOIeVoy/rO4wQoW2tq5dS1wq1
OOzgx9HyKQo3FA6KONCd9pVzpe/6oSktDdkfPiCh7KLcj0orW62vhIeekHgeb9xJhxu1lk8jNTPT
kQoKTM4ZdwMQkz0sJMUfiAzhd6EjLMPc5CaYAcTbqyRH3b2bBS3u9ELeUsA9u/TWsbbaJOH4xpN/
CBRQY5I1CFJEOq67WookQ23kZ3PbqMXzvKoewxQQkLZXeNbA0mnstARXX7D3kZmUdMrrt6BkwilB
E0m0UG4kgrkkj40MrD/K19rFR9P93hCj7OXlPIWLziXvmRmygoaQ28ayano9Y9mVYiRhPwZlSSoH
ibSvHh5B7+gizxhcjKXAKFOAtDXVQ4LdsaTqYRArJ5cFwqXem4V1thL+N0ZMtgY+2XBupLQIzrN/
FRA544HENnquhQ/2NrbUls/wG7B12nO/FLjQYuQJXfhqp/IXpboqBfTHSIipAl9PAwM51XPkSJq9
cl/tUY9kl/Owe7wZ1NLdKbv4jfGJJ89IS3G5L6oergexJhaWD0dKUCr+Ot7de6rS9/J+icPl32LR
nk9lwcQT9WXLx4IymoCplzOkef8tcfQd7cTWmlrgk0ONd71q/mmEy6BuzAkj04QVPxBgqE2NKpEC
4KI5nhREz1KAL/IeeIlXqSmUYa5SM86bIVUA1BRcNTy2pmKbNHDFU1SZh/jgkFTd1/gSEnkOdW7E
bkFaAu7HGqgTnZMKAUu4LEpGGTrL6M/F8byc68BvBfyEtuRrMq2gszHsHDLuHGel931ya/psbRJO
DxF45XJHWbQoKb/+wVnFvl6ZQIFdMtEiu1KinKZbDGbZf5Rt0D6h4+nqUCcaLDgZepwXd0yNcl88
XEuWe3CeqBiU0lznme/YIxIV9xg0hKqPwuQXC2DcszuULF3+m0cuTxe3DKteEyxdfbS8MM/QAPDh
QcXvkevLsgGjhuBwAI/RfCH3AUq2IKJEmP7j0Hfxml4k8afCYwCq1q4F6/N6H6FCmfd+22b+kqUO
tEbtsvHAkPn1Y7wC/HhL6lV6nBii83m5HPFDKg6tsn5cQ35yI9PXnjQx0O2x86sySelutB7qDww8
6pU9185wuxhSQEp+QUOPpdbRi3+9a5+b3HS6ltEI1Q1JnfBP2wDJZ0J4QqNHIIRxUohkHu6TAx8Z
sPjIeDA00vnqjtyx/H/zXn6t6Q0bMnQVxd87FdiOnaQ25k5QJEZ9O8NojxQiiF44l2eMCHm+DhYN
cX1PkGA/ynFpChPu1hxc/lNvFxrgb6L8wqhGOqrhVsD7UYj6LvHAmjHad11ATPiJPWgZ7Ezg8xYp
5Ybh1nKBp7oohdAveuBZFWuBBoP+cvOauPbFC6H7FNQUrdhLaX4qjQ4/Op2ac8+VUDkTc3CLNgjf
n/Fohkp509cBCSqVSf8gp1yzQ+lpQ13RNSVGzjP2qOvOLmbyk0RyA0yK/eRROI6hQem9NnLsVK0V
anVx9TalAKr+91Bk3DYnscNf8e5M6exPu4fuOXZbvw9amQJ3EY5KQI8CplR5Lvn9WFuvNIV8cpzJ
M61XgRNRxz+zM91tcouUTvuOBlOfV6Fs01gzEEvAie98/CG7DFXxueHPJ5YBs4iSYDzRDGIcITTO
XAo68+jZbdH12jnWuDBEWz+GoSSO5o9oqVC9ZLTS1P+FS5DKL5WCNqSBRpvivmvETy8Yn3PLtICM
Ea4+cW5D+DitLvPiyTgmW84yyGbck+kBv3/FcaegYBTYLO1fEHVHgG826gCHUmP6l4xzFFgiVSFo
/5VtydbwKKTvc/04yWb6Gzfx84oIgJqRidUyfO2f0chLY+R5alWjcL2iYJA0lTa+QFInrUVnHnvN
9QKVZEhRjeB2IiVKhHLTn5sHx6C+CwhFr2s+bjs3X/LWGEcBaQSVShl3BTZtaI6omKILuWAOuTq8
/GPI4PQfS7cF5UtUMaxx8id8+oSFuGblmuNDEZuTPkMfE+KMFnvPH3lA1Y7UiiLu1cfC8ol3cYrN
EpqhlTRjK3oqu3B6H3qD9yuPJNDqwuxQAhjJjr9BNx6KL9DUW11TwyIpU/9/7vbNekrrCMjBvlA6
ewkjYqugsfX9pwunSHT3CWtydSY5pA1GLEhWUGpUEyWyVk2FoS973okBr1I5MtNz4ButAPXAd9hE
rn/yeeVyDP/lw2dUlvQCVjM7Lx7/qDAoTd0OsbE9AjA2J9Tey7QJv4JsiN/It/soJG5gCkdFOxtF
N7Tm+rz59DjCVZx9xpNkX27t6V1ZLPx8EoQB7m9qd7sdsnlqHoysRQLZYV0GKLiXPDOcTKSOACr6
SzeR2mas2vFhFCTvRYWPz7lZYH1BM+pNyeDvkuYIQeI7HOYnXD6ECCYILuI84XVPLljdZrnGp9Y2
BYWv7OGhobJF2V+SZOTjMedI9VtTDHzDLqHgcxfdbPkDbXD2r3x3EbSbcl3+n+vbaGVX5Kj97otX
fYE9csZpj7vuLOfyDCWB7mzbw5Z7xZpd/npFB3w51Ab8F0hpQMIC/9aAGDg50ddz7Si7OJwjRJfQ
gmKkYqD1mSFWoWkSWIbZ0msKqd3tpgkKqdp8rFGUHXHFi6ft5LDdrpLoIy7LBlqonjPEp123dVr/
ewGfdk9gT0ml3j6Yxxs0vtbl67OwKpKsln2BSOxS7gFkHz0ndPRaDgnJoR4ohchAKkYe/Zy0VzNc
bw34G9tKUDegRGgcdkyz1MIylkHXaKrp3FWIOKSI6o2ymPB+/Bb6dUTQsM9vgTRPV5as2a6IeTZN
4v/YGVY7pwx1zL8DVJaeowpcyiUObJxtjWBtfswMrZKu7Iodqhief3q8/HiZX1ov5tP0WrkS7SWA
jD+u2La44/Wjq1URjk205A9ai951a6Qb2jQOS5BfZRmHlXcnG+QMJOz2bjk5VHN8EGefDwbQKZWt
CK3FdlY7luZre4qn4KYsCLfiHjEmJKAHl1tQhySpU6oGb10tOC8a1oERxQGGDSI5577N2Xmcx6Dq
3ccLka/ng4PeYIH8z8Z275FIRnW9Tkk2aXEWSD9kQef2ELYL68SWns0b4sRp6hRhlfFBptKw3Pnf
L823R9e16BFqPhIetnkgonjM7dCRDu/T93NEtFm/mzufNvyE15n/zNmoSJkjzY0B7eGVno+dlgbJ
xLFHU0eWXi7p/O1AGLAfXDJGiVq6ErcBzHlRToMMZbM9GntskQV3I/ucxm1ORZn82FTUsVwQHVwq
ZK6MjOmUxGK36f19sQ/suthrcobB5JjzNjgJAEru+DR9gXCQSS9DjnfswG1gMeWn4zi58BESj6yP
9CK/cjxPvhfs2vW0Z3xKf3wooKnTooRUJJNUpVU5EstWBLjUk3UAalzE3NxAYgdC8lyRFmRpy3ZO
KUMM8RZzKClGMKWnpNqGSBuyn7BYCu74gvIIprd0xgqDqzT53iIQa4EOKx9CL9wIpr0ivJUyapY+
e4lUNx/hHJKX4Nwoa+0mvp5WaW4oJatu5SRAZsuuwFns38i7sDyrHHoMM0FIbWqHNhEWjHe9SP/8
2arm674/2UVXMwwHPUsGWWc/vEycrRyaRUevmKY14RpWPXcL8zDkjh9sxlofJFMJe1mId1MDvaDe
Qh8PSCqk802wrK+Td8vqGWOEVc1bt1uLhKUpbDlyAP3YM0wtYiVDDpA0HVd0cq4tdVR7MjeKyrwO
DJZ8TNYaRqijEP8CABni4AD6fRsYsXJr4RnNq7hdUr5vB230k0yDV978kN+8u4tqhdKTpjl8WCzs
9eE0V3/w2onptDxU2fUN7KcavXG7KObpq75LSRVFGZgTOPAVy0loc7CPN3tgHE73dEkb4tWx1MKl
GZCxPyj5JArxEtI23LLZewj5iVgvJj1Oyazorw5miqCnht1ew4olThfsOHr+CiX+yOkGzVAzFVGl
lOQrrS3HZKOq+vpNIH8piSueU1SzcK0IpDnsc2ejkTfpvCrQok4nqy6+47KGJ1oQAphACvqqyhqm
Kk1nRHsqx07kNHXPDRue8GIdkJityb673teCDAA7Dx69zsdLKeTC6LfLNLTV5EKfEz/R3iVVBQh9
vI4Td1TaVGia+FQB+w1Bu3nBHgAfIcpK1lke1DCTwALdRXsO9wpgqgTFMT1G1jYWbfEk4b7onkcI
6v6a6fruDG2FuX9ABXWgQKuUL9wx9D0HhPyaas3MwBZl9m2HCM2IyZlLab2+n6wm4G3Q8NrPaxu+
Z3oezP+6gSF0f2lF+zEQNVKGmVqzDYeRjta2kIy0qZe2fKChqnb56h+kqyR8QhM6NCfLYoHGn0aP
H9E9SlRBhHJWZq+zOXfvRxpT5T8drhZBwItfDwLiam6wnpCOo3R7M85xmcBCxSNQF5Xfs03Fqsy9
rl4hvSqVMvxi8jP6nVP+5MOHcu+ohAhEzNVaDsOI554petXVXtGl//4ZRlvf6vusB2d/R6pFXYcf
43j+QacburLAsIZ01EW1m7Xu/YZswFCJadPwT8OfunZn5ogaZYCt9qcN4XvImEhF5OGyvoNPomNN
pZPLs3YQ9sTg2Es0aaZXZVCj2qxqLv3SSS+sVU07rQSaggkR3+jeFyfOhp4f5q10Te/cJ283aK2t
god4HTFI5QjanIeEhcfw2+5u7B4rNHgozkAD5XQAX62TB5JTgNMRMTcDDFqjdYs/aVQmtvUiVHfi
err9ESbvx2URRTINen4HGzTsE6cHZjt0s83P/rH0L5l6BESZ6PM59j6QAtqQez9WtVq+JTb6yzhP
aFh9ku1HRn4eWXI3MHWlMLgGO0qwTH/6v51be5nyBgPw8s4ja5Ip7NiHyOLnMT48jgZ2S2r1WFzW
LM1RjHhRYj/dLF/53frl/yIbBPhGm+yjKcZ+sHS+X49kyfrNmLaRv4erfnokqJubjDl6ktyC0S6m
WEzJGJZgKcP/CrBicLFwdOgGUG20+nlLG8k47FuHVSbcmFVKnVMXZkFjklH8Ihhh7MAXC+ysHHGz
12SkoBcM1+m5fToJdJRIADAIwXOdF1LJl8DC/+x1+6tl5uiZKdO4J7Lbkvx8pxxUqtzBnx3B7vlF
3qq/L7t8uqmqvSXOBthyZJMQDE4BwAah3QFiigolcUIZO40psk7QGgepKYXuRKYEZcOe29y6Bmaq
Z5NV0Y3UQqbm3qmDq6/xYQuRA3ZrpaDndcUDOyOOyvPkvm7V+jSytyH7qSRAObjr0gyYF4K7bpVd
UCei/OOR4Z5uQ1VgGYuXqy1S2k4WFsTB7HVLkZUYmIjXuSah6ELrOWp60KZjE4ydAclApct8rkRw
ySLjSZ9lP6C4ceKJn6P9k8UwTZMCpJ3zuaP9i6yML+Uf8DWJfPNsR1Qm6uSSwVR7E60zyERdE+yi
bks+VxMQmFJxG3imMPpVpou3SUzduFh0WOFjCH+cif1d6jbIyskiJWhBQjfGhpRx2L5DnBg+9vqQ
DedpH9Ux8aT5rd4NOSj3aaM2xCA6y2EmWiQBhk324cgqgVwVJiR8TXCKphIkmNSHpyO6Q9WQsQ1O
qE1aEQAaQBxtfNTbc/cptWFftkt4gFMmc8A9/nofrkzzKDQGaFWDS8ZyIRrmmXNvNHmGPNt4x7VL
crzG+KT7y+PCzrhD0RawaCaMfgtQCxHH0Yhq6ilZSn8QhTaoSpN8nLfcVmk0ZpsYJ4plyYOap9lQ
mFcu9Uvh19JBmY2VesoVZL+TaKvOS9Nl6NiHOi7jdVhKjrUXZDfY25/ixIOf5hob/gdRdggWktFJ
ZUw/CUmgFG6lru69mlJhaKT2j+M2L/Aiu7kmcLscfr6BTpooI7bJlJuP3BUe7k1xO17oETAjQK77
hUB7Il0Y4Vi1Kaui5a+m/oIMLB1/+O/DjA5orcdYqxp5MHTHh/4R7glegBGB4QjdoNH2i379dsil
JUOmKnWryLJ/HXvUbfDgeUTZwLm4cHVYK6ewvGcq/Ti8ZhIxjB4f6rvE1XSKQvTKNEgosblr+6sm
YCoD4aH6S0gDkgfUjPFuY6mb950THrpvNrkglWjJlCgFWIYQhovJpS4uoOXQCxFkM7zaWHQDnzWI
mZc9B/7BsieS3ANoF9amEpGYSGnguUy3+sXQT4Djt7k9yHiqXAZaoAMbeNzWNsxSN7GXYX+Jvm3l
nIShWFbnVSxKByN4hGXivFniDU9a0ZdAaA0cMKLJyYPhcshHVM98+M3d9O7ZfcCOBri2VIkwIDQ4
htOlPpE+rqm53YTXw06Omp+0p6BLab62QQrecb604UVhojQCNhQ26oj98cwrqODSXE8c+auXHxHk
gWsJLdHgu0QwddQO54Wsg4z0azE5n4Dee2223Gj0v7e4RZkiq/NF6tSHYLzWvplYp4hslmcfW+HX
7SO5RiZ+4stKbKoSksSPoGjoAQQkq8w2bvwBuJ/mcM+KuPLQdCIScXxlz62ekQ+6X4FuZf9nsHBK
N7yvZSvYTSkPsplXRu/e0Vi1WvaAedzPw5cr8848eW9WpGXpq+3HJnmPnK0Jn4Fay0WQJjvaD2Ng
Ou3MgdgRiP7GwklVRZAhqZDrAndhuisGG7h5ucqSQeUtfD6xoqPiBkmIvdr7awRbP6N/vr+cGTqi
zNJ0GmxPLM65d2LBxBwyZhjaytGp5O3Cqep87kJagnPT8hG0IOPiIzCDKODr0tBveiNdc+qhR6HQ
Vc2oN2p8l5zjA/l3PjXT0vidxZktIlnJmgr8CyGSR8TAKcWIiduet04pvP2RFjSDcLOtZy79A0dS
ajeBFJwujVSkR9mtS1P2nSgJZ0LaYERnz2vluwTrQ59JQqJa0I1jFFsOJcbi+alvG2OI4L8h2ZiP
Ne1cuJIh5Yt9OHalZoqad2ZKBSok70FJ/OsH+m26zmo4Hns3d6XSvvo+5fumb/RNpAQW5KjIq5/B
uZjPnsxZWmUortvV89Hhj6cBALhOqiRDmbiLPStrzgGktyKK3RmXVpQwLKulUSWnjts09nGTyDPg
o1uX/35G4cDxYDb3AVKbPor7ywUeN/GDoF2MJRxEiZj5Pf0/5RcG4w6MV2sgSXAhssJ9jajvq++X
WP3NWsXO1z/LweR/N/mfA5zLKsGFXlArbBKmC2A8KWVndO595lPHrUt/zkFlQqNZraQgiOQeGuN2
lOu5VfQQWvCS3hHLHFZKmYyg8y99dvnvspkVPC8reOoa4+4JFXgUdoyNXrEy9LwHZuReYyw2iGOB
+lpZQidaySq0jrIE64uNmg6eQuTT7+hRZuHI1vfqRth/QhRLl0Xr9AhfmZfiTNBZzgU3BdDG8G2m
xmMSkVWl5rTtZ2ztrTQBCwyOBoKCL94tI3brK8SbwBv5hLG4a220VDzSnBCDRQXkiGd+E75ICvWZ
7q0dcksAbYr5bbUHNahI9gfCcQ0ZepNjh/l8KA6YMVoZIAD40IlgAZQUDZ8q6yHyv8f/7ebjqZh1
04wC7GeqtuKZAgWtMNeKEiU94GEQD5uRwDR9u9Rv0i+zBIVs787XLp3VbP+yP8ETp7hl3S+gTTFG
TyNl5YtQAh33ub/hXeoIXD7uYUl+eATudKonp2pxxfhYFn+STyRa7jpsra/gq51Y+oAam8LCbKjr
wTSmJ3buk4ZAUB5lfIb7lPWjLlHfFq+BsTR9JiSr0gPG+gAeV2fp/+QBhlq8R1A8JPwMEB8poSfa
gw7z/oljbaH2DmYSrFm6YhdJVI6KOkfwd8ZD+wSneKmfVJiAqmvaJrJEIU0U6UAUlYUjJrF5h7+H
B4OpLUOSdOSbffhPR5DLam8+Kj8EsSpTJHborSkknYZPxPHNyyvA0EjpYZGFwPqxpCQ/QEsBFeDU
ayPPbAmGADTCPOtTK/MTL3bX084f0BTvv9m794sby+/tI2/uQBtfHMRCsWx+asm3k6Dpk1DhZqgZ
u3KpHanNApBaCMEKdrWyk0mD+jy2bvXtuzMPnyttj4U9E+0M2NOdS/+SvqKEgCnmmZ26i5H5PGj3
HsoNA52yV6BU6FvvisarzfUP/2/ODg+OGVrPF1CxtO0Bn6INsGX+gq+Iz8ukAZJbyw3wm6xIhyS7
krysYkQpF1RELNdx/P5N8fyWQaP7Vl6yYqKKBTE1lWJ1Ym/tGi7qLIiuGK4p7qCJQQ/cIeoXR1Y5
ZjZcTuGOF6tHPS/cb/nulp2HqQ9LuCq6uViDmBRBb5Gr45zUa2BikixzZney81W6mXNGR+pykkwu
qyiGNle+54o/NyNsMf0ArP3BVIJATdVUkPATOLpPtJLs1SH3qK+5wOJx1R1cWt9gF1QR8yy8frtn
dNcLbTY2EcwXHkjLi3VRsbvucoJeDRKEJduBCe1b9WU0DDxQkFH31EqHKhs7gc4Z9z74pDSoTbpl
vYm7/C8naNgBGBVKXWGIPFM8AA2//GhSgth7JsLLW7/gnqlFbRiq0evUGms1RFu5iC118C0+uQzI
MUb4YbS6KdPXrgIsqHAfNRga5EvNrow5xWfPNaJiCxpOhi+SO9k3og4CD+T5Gw8nwUJoPLeLnAak
AmydcBCGfARgVcvvI/cQDc6zrH9DkFYG2c+msmUuO99dDJ/SON/5Ss5V/HUuvBZVd+amf6ZcQlf2
Vxai8UfUEzvcdQV9+shFZuQVWN34lt5NAx7afTxY+Fgk3pDzz1ycK9Xp5XyNlfH3CvvyBV/vZ8DW
FmbdTJt4f7Q+lupoGVnZAVphEffki7bRMFSJKlubtHJ23pSAX4DXn3qg89w0Bxr5gQo0XT+d0Cdn
KSwPw3HC/vE/ttK+WRnwbdtBf3QEyz+Ig2h5lOFNzMIwj0qro6jskmwnp6reR9yUh4S41LDY8A/A
DcSpF9i0px6VIb7UnT9mtvfNCNFGR4oS/qKRGMcecIrJtIC5nEAqFVjQta2mhvc1mmjDeJuJu/bk
TTixgpw15/7giBpZywLZw4MyJXdvMTvIYNPNmwFXTyS+pSFiWdlxnfa5un/iLeRLa94ssyW9Aiyi
HXmTJ9WJEaPV1opmurGz6UG7wVd/sQH8cGtZFub8NoL5FwSlfxejjluavXnlmgJ8luC5IGChP0ur
cz7KZdBJDyncNjr9MGbhEbOWQPhxbzuxm2Ucn0fQZWNP30hpdYjU93R4SrNnRPzAkRkW5H951iQ3
L2JWfu59q0IFgD4Xu1XHhlujiwEKfruQ9pgEyRq0wFOnt5Ze1ZCaeciMWFobmSS0X2wQVoVOy3Ha
spImuNVioxR2vfYyffW8gSmEL9fiEfAw+he+jihfQ8/6xSkOAEJhutGVFkagXn85AmJqlXvNj2FW
+SlpeV/kvjypWOfrUKZYJk5iaYE7x8aJ9Xpfiwxmg/Gl6hfbmoKalSAMjN4iw/BPvhdeGR5EzGeb
PWqtRO+8IX8OPx3EuIODyo1w4Wb/WqaoKo8cy7wImzRjgXN/FFVwp+0/4OTDb8r/bfYUcIO0z5De
A8lq+AjATC+1f7UXTi89jEEUOxe102Q/bbhfocYAdz2B+0bHH4iaDEPkbR1kNzn8AF6yt+GHV6Tk
ZbJJa8e/IaJNflTzkddQeL2GtNLV5LcrySaKaf76JHjMc+fWO4h+SBnTlN77HygP1NVD5RcfEWJH
u/1dhX3opO3OZeORx8aNHR1qCTsEjEsO68m+0OrHgXV9w/b4/DL0g61c9y4c3kpCRKovOW2AARUt
G/3yoQ0yQ38VEpexc3o8lJCvHJODrshnPIvJMTVeeV8ldKY/kAtpUNjZR80NOI3d1zMB/C/JS/UU
MHuT/jqQBDe4DagbUqRJA0um/setRIvO/GZMbiRvmrKvbRhRvKwxMfqZhSDaw1dULPz3fnXO0O+q
NqPs5Snz+Gt8RtSz5asjdlUSW5O0ZqHvRaJqZVCK28Yz2LNf1o/gp+0JQLkfqDrKuLZzTWDr9Q5Y
KcwdHPKmI9QGS5TH95xFJ4DUufxUjAf86X95DXWxvQbKsvmuk9MhNqOQaHjNTe3g8c5zNw2LoRIW
XAcpa1VpoFn3qC2QX+Ag57bBCYLVhksbe4WJPTdDaF7ZFa4FBK62T2oI30dQiNW6E8/sOQ2LI5k6
9iskNHkWhBugmJczkxszmBVljnY4Ivqs1dYmMNdsYPTr7XmlgyEkPtK95CTbsT67oW5KJnhwxxRy
WLUJt9I39NxaKXrDGcnqgg/qAa4fjCZ2wOgibaBcdb3yhenInNbT/r29FMFnOTB1nqIFx0gsO201
tU+VjCiern9zRcD+bG1dZNGWrW1DpOCVa7xX2Vo1iju2oVbmdR6vaBiPfJ3TFnNF8g2nQF/cSV5i
fx0lqrYX4IyGUPW/JZJIlHo8rr4tseilLZze6XqBnfYe/RMQKydLGf2owO0DiEUL0182SaHtOwni
+qmi8BzGZpSiwW8T93knA3lOJn2DyI3+iwo7RaZzBO181+xgjZea3mZRsPB59BzpsVeCdGvcafwy
i/cPRXIPYYRqsawE24O8Q79rcrwRrXOxeJe84Um3H8rnLyPvQOElcXR+q+yocHYPc1ahXMbfsB8y
GLdBD+CnQQcIFAQanXGvkba2swWcIWAllV1VYCEuOYDaXipauSMJxr2ySR3bkHMzs9uJO3/Icvor
fdO6StA54ERBnZ1W90TvQ2vxXpZpMJ7dfBGCpO7r5CL1jPUYneWyoLF/XBkWnYZBsB//Fdp93A66
ncIZDq6idGk3Yg67NLsBa51k009RNF90UPVGst49Kgxg7oA5AQVyJNgwrkf3xbNar/8V3ja+gHHA
an7A/L7T4/hdSQY2IASUZfZUx5Wb6g8W2bI53f893R7b4nfLX3KnjmPNCJChczbo8qMD5taEUHIa
PLq5x+OfMNYwGMytA4uC2eyfVUQpZj0zE3uGD6fiyr3XO18i2a8G3IFV55gy730P0s1YjvTvRNhI
fYEWN0XSvePZuWrKkoV/89foby6gxBm7/dxTuqHEPXtSSdx0nUSy2CnMCc410oKDlzv+u2hvtOVk
TJOoGi7z9HIFqBZsMlF8tmIw9DLWgrg3bc5YdKU6R0sRC+JyYy0KOZEgre4F4LSi/6fqStdwyPLl
dpREO9yaS7piJd+lWuqIMWCFKn1Q4somdLA3dOeX1B6ZBZuDFCqH2FZ5AXezJfmUyO62DFfXjCg/
WZJhoP3P7rq7Zs3iNncby0vM6J3HyyhYxuuNXiyxmpaj5M2UnagUjrwuwh4G+oooyZIVOv8FT2j1
eq/K3KQ4ZQ9bvy8OOifxCEXIinGgC7L26N99UeomKr0lF8DXm677vYm6M+94SJ2Q7bBdSUACS1KF
EVoMhxnmhEuZICOTPPnrjbM3/28nrWmMmhBJkHWNzGL4CdfcZigE4GHLn+NhuRg4hHUdA/HGurGX
Xr6Kbnd08agb5IWWmQUc3HoNTRgwnMq1f0TFFNKAg/xlwbWMUO0TUBRCHWojt5BiJs5FaaJrapBc
TukZ2RnORfYen5VVve2P4mxFwwu8TaxwpbIO/Afl0kRjnjL55v1FGjE/p1Zo/mt8HlynUyzp+Ls2
4mbG1CFkgp2INCaFZX9OOi7341Z4T2UHQE6RqfwS1potIMmUIkePuYvgzlNi5PiTFWYfjcrwDblq
fPIdxH+fA1984lLLZwONTRi3fnWm5GbuL+B+qknG6OUTWPUNcRdm5mOH6+jEkoC6dcOykBFLaJIf
XowfKO2mylKGOWdhHjwh/owjIsrm1vLHTjOBBv6A3kQIt9Xdhd0QVcMZJy/QrM+mhh5nu08LS9G6
QH4PzOdEDZwH8tbUARxxxXfAYS+0dtzEVpJrBi2TDBcxnzRosZG6BLefeV1JiM1oN5/8/Z5nmQNa
L9ZlqXlC80AsamxNTSKnkTt/11AZlUj1HIdPgKN50F74Z8ZA7FD/7q3Ex3j4J9hKAmtL4+98KChS
lZfsMCTcD1HivkVOBs8uI9OSfHs4rjchU0W5+jLH3j7vv5/tagQssAGQ7EsYc4FDiB/z5z5oHEH3
iDPjoJ6U8ruagPD3GyUTsSndJGQgq1X5m4UO4TIG8fYZfMZJ3tHEL9n/3ppfLexIXAWToCZ41QEI
A06UppWGYy838MfxM21S3S4VYFNcx9B1pDAMNbXdW4nimOSilw9EKLBR24oazywC8yR1fNbkv0F6
uuRG7RL5bM8+AFf6ti7bJD6pmNdPGjGNhrMeQjJgMxiWgtPi8t0KPLXAgczJQZHyEbkxUuqFF4tv
k2rXMatYqSik8LZtABRzQqxLOwuli7T7jW/PGhanSKa6AF5UsU0xGMNTwB2lL0tsw9/v869pZLYY
SW8P9CNAqmhOAlmGL3Y5DvXt2yIjmS9TniF1884LrxB3LiJDn+PD2vjRRdp32/7sE39hi7bP+emb
+8skFMeRjY92UZxzHZDAhLTo1SL0iDet+16EvY4tjFg7L25jo4sSN3DW36HlN6orexXEvHK36Ody
B1tLj827QMxlMDY7uAOnBlXRAXUZicYk7ybeU5oH2rqPhWED9Lsz4jduQYHmPEkxdIYcsxfIlCnQ
qTAecwUWbICpvzosLN11buXIg801iYn31OCUIVYI+IAuksNyRP78nOjUzsKm3FIpsf1f2GbW7Zmi
dV/UcH9xYdO343UyrVf0B1ypVvC0O2Uzg07+Aq/Q02Bc9KnQN1XkwN54TFhh1QA+Bxbn5Li7yHtz
A1CUNeFz8lzGXqZeOmWLPZhsYfD2Z4mBhNQLAynXNIxl5SHLwDUruGqmvozfwwMcbDGjcD986aHo
KBIERhBW6DjCbTnG19XAE+55LbVIH6+BGTML0iSr4IwWwifpRUUkNsELQMTKz5s3tjJubdKamIVA
U9wH3ry9+WyDRs+2gcNrDsARn+XWhA4Kf7GIb78sQjzjyrFa2zbJVwsv3iHsIhpGKPqXsuDGy1mc
wXoTPlhxxU8JDyfDXa+60wKqHZyUERybwBEWLfiTt2gWcfaDHIGRhXm/CyJmEvwob/tag6oG/RrY
4M/FDvfhxa3e6LLujufvXscs72UoY8ALJB9L6/ti0MHNQjSQNIwEk5nUKwUbyG1j8bvTwgms8ZSV
OryvVq+kp0RY+9Z04fca3ngRPQQw9marKBI6aEtMKIqyiZGuQy9S9Qg6dUMF4zxfy7r5i+0+bASD
t32zmGbHwnqwi7+ytY9G1gsiqw8XhFqiCL2wgH+z6AQkF6+RBKUH+J74IpzykG3oLL5WYJm6me3u
xtPcCYpkpzHyvEKSq5z3yUwOXzV6qgTXsgTxTn5RLsW8Dce7oy//bGkOAY9iV8E+yGgbTjKXnVqL
iFivIJ9YuZytxOpsR/cxabIyMlnkbEQEkMt67QqFJFKKTqJpIfO9+vCyXdPzy09hC4rYOKe+8rDY
pxteGde1fxF5hG62OQ6TalkMCKhwcKNgWzxjd8tALecAQ5TbMX9CMbm3oAxoFXpJmfeTQi9px53s
qCd5oNt1pZKVoHp1OjDPcdBtOtSUyECHSEURutMTLBkgXqwyYq/h29IUD9hSfp9UjCrPVu8h3yon
pBMyAVmQHognGHPWsn2A0vqt0966itmT4staqrpcr3DaG7TBRkBDN1nL+t0gmE1h+GLJxAVXRM8N
kNWo0P5oyCik4K0osVo9+9gpHrPRisx3u1s0+mYKuzJ/8AFqdJyGfA6Gb/pMdOtYBpqye3vHNf3w
IH5OrNMSHSEgd87qDK8Z7n4wjSAa1glHBQoqxLMHpqIkQSiirPxcNx48gcIwup6CmY0ktvTixVwf
pE1FCI3BOMJ3bhyZBPddqYN8bgL3DOIvY6Y0sxfFA9TbU4u7H6ttuK8z7HGWHFD3E0xvhpKEtLXr
7m3VUkeHLftMkqn8eL5WJq1KUqcFUN48uuxADcEvVsTJ4WTZGsfdzy5b0m///SccZGJj2XSzBlx2
Vb+uMuzmSiv3nLc3JJrBokD2hT5bTBDUzP+ZAxKAkwSAJ19NBZhFiXJUN3D6xmhCzDuv+i7KKqTw
BUCIs816SYkrxHicaJ3nB3794Ugwj5UsSPiY/YeVMMq+j1IichLqs8mbHhnzCrWarTJ3B1HmWT16
MIubCrunpa3OONYfISLdarYA/TGNbn4VVBFAWtPazK+pwN8f7OHJ/iA1XqGtO14UB6vVAc5DafkX
vFng8jM02ObAEsvHM16+mdHutCrWCQqwQnHzfTtzlhw9HpkTdmcouE9xi4kiehkgfbZL1P5Ku1Ot
NByc8mXA05uml0Dhqyt7aoecz5ER4urkYrUuHbWMuNTBZRhwLn2Mu6Jqc8apdBJlD+rYyC9FF4hL
ScHrdvLDDXm7svu4si7PGNpSYJVtU2japRs649lj4DgLiJk0x/K3Ipj7ufpkHrQMXf2PyKXgTrCx
gTLYDBY9KjVETigciAIHzPNKZcfMfst1P4nMzVRZ/ocYr0InbR8MVtMGhLbN0eUTjMYTgtjl5fq3
BJUUtMd9b/1Xf6kADz5RgRo+PxieidMTU8TYGcOTrhNl9Xj6LFWtZTZVdhDhu7YsRSH9jFmZu6Kk
vLoZR7mUutLURHygFbFTaSlo1OaBYydCwo+kho0+idk9ZotJq8vToNEGxL6Pf1z57Hs2URSDliZc
N6vaWO0XqqIHaPHX4QShGr6WHiRY1fXhKmFGAFVGIN00lFBgasOFJ/Zj6vWK+fev71kK5AMbffvL
DdjebxG3oiYIONQUA4DiVaP4ye9e659LkrYJ9v2OsCpO4QUBde5wOv2zcu55o5LMD1l2H880+yQ7
XGz8v7dPTg3BMKf1EfY77TK188+PjNUed/Y9DlfzFY2crZyxPeXFm1HuNg7JV2FZk85A8NT6yeG/
S1ZrCvysOngFzxvWlsk6VLEHgoAzoPsRnMwG4mzJl0mpL8JgV3f1a8owVYhQL5tKDcvwkljXK0mJ
5L8QNXeUeQbGMvsmIVyQPKYZT9n2vujWD0pTupuofaf4+3KQtvlfIyH3T+gWwUTBQ4U/y5kQW4Jl
t5y8oPqgKOsFDGBneSvdQBjw7s07zke0Pd8VKOJ7XOe9SaDsa/0YEURewbrgJlsHEo5n80qBVbae
NYINarftaeI1RABrJwQTI0q0VKNfZQx3Iz0FjS6xs9vIzOvHuj9Yp8hI2/WAwN1MmxWgy/Hbs6N9
ki4IERuDPKs7l6vX+Znx4AwCOYQaT3bMeN3ve1x7riEA/oWAzPaZbG125qVkPmo4997ZksekGbe6
iTfFYm2rKjfrchhPxzHCTP4ai28l2XSfV4/R+WJ1xs/R/0WfZso2qaLvbmqd4gHQyVxhfSun6+aW
ah3e+nHGGis+1KTtGaE+ZQo2w+CIu5rfuK+2cnNRhrRcFm2AG1XADbxkXBKdn3ahLyTxxUQioskG
lRhO4+bKFoAXEUYVvOQmlq8BytXMe6Jk9IkISeiWCjsj8JomvMN5BBsWn6tUGtnwHFrkW4bmhNjD
E00fC+zcJMpSAg0HrdkkRYEbxAlgmHwduZ/DFOBdiVV2zvlDAxPJ99rukFsnUcryAL3LBJq2hxmO
g/jTR8sF+6/1Fcuh3ISPNoqEe3K563MxD5oM+ZUfCWQIYNWL9DhyS2ni6ZYloJvHBMmSZOJ91V88
S2V5iLqTeUoaH8nqGFkJ7n8mqIgQpETABVQPxNQ+T2dRjzHnW8xBniGi5yf8y/An8pBeJgJRNbyJ
fRZQ1HlWQcC17ljJEOKp4x2esgiceoQFe/vVK5GGRP1+yVez+NeDxnp6B09MQavwdknwqmnsm4IG
DEYGH5YEsbR9wuXZ+mr5InS/knW3aDfC+jmcRTZKl+7wr9fiBK9BzTOllsdbCXFtQ3zJbnVQVpOg
Rs/3cymWgqCADVOLa+YwVNmQCSoeyJt/EAaC5lE64qPuG5DCrH7dtHZkeDy3yjBx6DrOUhDGwkjf
NIoMffBpIIgj9b4kDVSgsIPpMbnjXtdv2iHsMHkvSUCPXLARA58wOX/MYV/MP57WQX+bR1cLtyMK
/gvZW/eYhEfO9g5SNjABH+91eJy3RMSh7R7adNrZgVZxXKtaCuhXSWXsEFAEhdoeV5/PbkxePOSt
JZTGqsrC5kM/0kAUJYyKcvyEJJAC1eeDAexU9xMHr0qXVl14NCBug/fYLQGSrvT4FF0ZMjjoCFlF
t5NITaWcXTXDOnx3kOciAQElnPywQn5yMQltGioYXZuUKzxULK4C+ad8LB0Ih6lYfxD/OpkPny3i
fs3JteiCBKmjA/cfqJ7rSgzr97uBKD0aKKBmYFMHdoBrPKSuyjRF9vEP+XlsdkKqaItRdN94kJ1P
8mVO9XyB3oz2QwSTxbzj5+KXrjomxXO5SB0tIJ2D314DoMDamm1xmZyCFPAnYghwxH+VamdUS2Nf
Lq1sZQD+5p3D5I9/vbsw+nU7yUM2GkRMrGTLPuoI9z+xu6znrZe9HTgIFeiCGVXiH0q4i8NK0wwX
CxdPqGumz1jVZVcpIOXWEgQRKaM79megSXWMDzDU7g6KmOIxIO0H8wBWmDBtG/9zos8dgOg3ZgFU
woGmsn3ZPh26TZkRXM8c2S2sTGnskvAXqnEvp0nHFbRoZbDedPv/R3yUXdbc5TOMtDcCwLqnKq5F
KjfbLK4cXtI4mx1+/8WsTtugCTK2IJEouLIQK+gSfWzH3t7XgIxsZgOS2WjIQh4FUt+W/du6F+ey
zHOSAGpciRxUucGtmnBVwoNgLd89VH8nUgk3epWpgxZtBwxBGnx0McrtzSmS4h8/bWaAvvXWFnti
sOl5ud7OGvlUKKt2RguXRZV3vWGAvQKPwfcYtIHzNbOvLNvoFKhN5CNf9Eqmmaro9U6VPFUicHEb
Z9BeVK0SFcPY8ZO5kgd8OD72cIvgKTYz39TMgVEI45R79IjoTZD+GPy75zPi+pZ0+VwpVQrEkXi9
g4BE77/3sXjdU37qjqMEkcxrjJH6EX/oFqX/R204ARLN47whHcLt45bkFSmn4Hv3F7LaWi8U2DLt
jfGX+I0D+hNT682hEFadOpc4Ntr+tN1Z10twSEcmni5c1wPqF+5fMK5qwRsKI0igconLwQsuvqf3
IpEXOun/1UKOPQyXWHs1AwaIz955iA56cNYpXk8+LFd5Du2DVEDFhnAR1ZB6VtlLYP8SYjUX02OG
YJJXFFVIHxcg6RWoBxkZk3TbmA9gdkMYEUR92sv4NPHwtifaEG+sIA+5FwrCPCp5UO8EkO83Mrfa
9uyg7n2RJ95Jj860WrFn+lLpir6S/2rjhhidzVAqJQb+6WtSIDXUE0HVceYdtITp+eKTOaXJLcos
O1BTKA/+xZbEndqIOEyp4cjqTH9XmMhGv5DfntN+mUb6f540G+r3FBQM94fXqN3sGBIt+91MzXUi
hm8+3HCbv8ENR0EmIr9DwkJydEILSYGSj52GXhA3x4EpBeb7WlUN9as7MejbX2QvoLrr0wvfz3xl
smUPShiSeJ2Q77ZJbLllGtHoagE5egH0avJBsRb+opmHMYGGqEijfFwUUzkiKG2Nw1l2AkAEPdTO
eaAvnpvkJRZiy33uVgfgtwNiL/8zoCqgY30qWbtgZsVPGWH9kd4rkB1a8nKY90vTciJ6k01mzEHI
DpQ4brF3gd/9zzrVYqYRt2SudbVUPOpN+ej75lLB5zywj9w68IkB2uaFeKtw5Le34omDCw0cAOi6
PUqn7peZSEVB0RTonO/F/qg5nMxC+FD+YutZo9D07gbRKlHfXKsiBtQDranzYkLbEDFc7R9fdDZT
bG00dVpM/HF5pqXQRpE+8XJ+dZ3T7N4IllPgCAtP7okomVwpbPKFNQyXTbcAMKlm2dOw3jrr+Jud
u4jFjxYgqMXLRkn9MYNR2R3vgKZBlE1BaIbMre3VWLarLOpxgiTosU641Tizon+v7LgT49iDQkZH
lQdjxqVo4yqvvhKk2yiahka6Du3ih4vo4dZWunSUilm/0XoX2iHAKzvyI2lvEHnVO3CYRtnK2P93
oA+RRI8I4s4sjP3OCjwTZr/uUzBes47TLZYDAY0l1cBgLn22ZYJCy7dbi7Yc+Nh+Q5BksD0dBMYB
bsVsOQyb4ciKSmegcZ0/tNweXnkwdqYdTCtXsbN0uRXXHO6sUQBUhOfVy1ZQ6d4IfmP7gYxRE7Ro
noN4qDAsN85myegHonyadj+FbczyQLdfsLIOc5rG5WEGBT9ZOPRFRTbd/SrjczofJVQ5D52gR+WL
UVaFtEhPzLtOgnApxRyjtSy4KdVOYu89RWqIW/gciivoGX+T+hL9MJrZi8U6immYIqeOkUj3V+Ja
1CZrVgpiqgZEPf+gLNWsWJjL2XMkZkhfl5o8rKvbBl5FsgCV6qvLn4pIsje9V9fMWSaLM31neiju
vN6k+9+Bui5vZG3t3micypEujHBeEV2Ln5uLxKsaZQOJFvkRlZiCkVoUpKm08tzOUsfd14sVoKT6
BlT3FQqo6yZsV6AtVFqdm0JDS/WN5Pe9ToHVWLFilDERxbbVserj30FUcUhuugJME/hloNyFYukx
63ZJIP3l+bBGXZ0WYf7RiXl3yOT6Gee33E8RDToja4eRuR4y5HX3GurHy+BY6dDxneOkEm/s+iYC
dhRxN7u7YAN+kWKH55sgQUCpSKVI3gpVQyEFfl3rboIYwymuQVtN69E3K2jh0WJZ6Cko+qdFDlyX
G1p2AKWo0NUbKlw4HFibzEKrvG6FgfS+Ir3Vpmd87HjDfYmPnVBsJs1q2A61slQu6MminOXyXXjj
Sk70RH4cth0TyA4IFweDRLZd0sJx2XTE8kkqfLz2plwkIOLtjx3lgLQJjRoQ+JNQVfIw2RTyxiKx
Qa5Mce7auaDRCmhcbOkF+uqTW9IQkAtY/N9Q62jG1wuTX5c4SjliQfSsTPkhK/OYyuZsBlefs8xn
8CXIkv0DMtPX9dbH033CQjhy1KXKKP8y41WwYelvuNxw4CR+zmNXWY0tKLL/jyG1o3Y++jSaCawS
q1ThduOu5ogG4xFnTJKV1xiIhZd6NGY+VOCSQea7AwcbTNJ3+6VimMNEQPkvjhq60zMemkSfxBmp
8pkyf91rgotX9BZ5sPiD0LHQrSOAbZ8+m3Q9jGC3GyW9YT7Yus2e9hUXkKUu9eHcUY5xVBkrKYMr
JzjF9VJuKdOIb4IIG8YxL4UNb6IKZhlXRH83+whAqWwQeV8gDJjDheketkcWnjq7c7MEbANzEFPM
brAjhjPKOcaqwLfFsy98cFJEIV4NOXgzHFymitFtbc+mNQMxuxo4vc+LLe7Tf6UiiSyQaZth1TlW
3nTe1nacXWtioXu3DAzDVWrzID5x7LczLv3vqzq0isqsk/k15VmeaSSQbupp6j2GCEdv0ZfLr1Yk
tO0LjXUMk0fY3AXy+V+nJs+7/J0ZTk00glGHzw8ET1FTtb6jKrr14Ar7uWwus6dxgjZwG5ytS3T9
vL8RDt63K9cF2Yj3y+onQkFc3ANelXte5HtYWnG8YA0CECnDffu1JjggFYHTyJXg5iFPA0OjpNn7
GaFGZeSMbSmHpQbAvdvJA5d5snhyj9/liRDYlIYws6SAcYk1lrFq5BSB4PmSO8K668ubmjQkf8ff
KapOJ/3Ye8kz/QARf12Pw9qxfSW53WRLnfJ7/jwc2wWUcRWsPU3ME2D+9+dGdx9dzPU9iwMTPTYz
/oYcqNaBoWgOSy9YbQbvMrmbI7bWgYzk4jzeTUkOgEOrK8Xg3/JUbBrqmWdmycoW6nysTh4aUGuo
1dc8aZ10TzPeRougDtLFQVMeziKXXNXWg3CJxGStctPjvbn875NGneMcSQy6LZStoz3TiWDFHc46
Z/5XukjVr0a5EOthHnYVKtEdK8X+iuSM57Hu0vKg7JcMMDeCik15S+p5BQnLfVhfo3qWXrpK/6LY
Q25VxaAgMMMeZMqOshjv3Q32Dw3S51uUXPkUpsfRXiCCpPsX1s2XrIzWF8G2qE47b+5GU9e6MZAk
ZtdwygGhSp1EPhNp1jdklN1W6baCBaJy+5GWTYc41LMmZGb9YXoR+Em/gxZzRdVgNBj3WMGKsE8G
g5uQ4/Wrow9KmZJ7Wr1m2hUIagihe0duZpuJfaooR1Qr1GanPSqisOZNDsZEaWw1LSyk1QEdsyDd
HckYfJcfR8sNcEnYFNKc7RjlGAAd5Mr7znRqxpP9bxo/HyBWM/QbYJxsNGspZQONeGsZ6AYGLc+Z
YDW8CLMILmt8T4ibo2m2TnnBENVtyMseUHDYHH+ixkHyfmJcx2PSTAOBHvjWgXbf+7dZhgZalT91
LZkA9e7OVaPAz3w9/lOMG5LZACzxJRr+Gp8qBS2db1brtXF5KCqxknvi54H3Af94Tj2FNJRvp5uk
cohOGQw7CacMQleABD1lVw0tR2EKckbYHV7ycluAF52zdEW0foifJvEYsUpIlQ69hpGD/DmcL9aO
6Hx2cQWDX/Q1WDEY62/rBoRrFaeFf4RheobtqH0gzu0gpDMnCHQxwHyuOYslYIiFpd0s53Z60kn1
rh8F1eDlimQtaUpW5dN+oPen6Qjr0X50D00eUGY5FKazDOdNeqSU3T77PhGwdgvWCvpTwst1RYzu
B7/PQ70+N5rP5ydN1+0Ug0Vmm+h6lMwOAVXm6EPyWcYKxM9urfP1ivtwacMswG/Eo8P6llBR1SdY
jEMl5PvJWJqS+LEfa57sHMujZU2/HhWKAfQGYnWWx6bIRGGto/vgy0f21huemv9mxQjVlDfVtQoR
Zxb54E45E37SSs/dBiN5jyVts53ycuLWCthuRZKYLR9eoO+gn/Vh7Rnaf7b/t6gkCT5oJrg3lut5
LvaLVo6W3wvxzRv0CQ7cmyzfLSbdH4t62l8zCDu+HSiUtFjhdwagki2FvhQrbvwV2ABscKqCgQnn
r7Z0gYGrAmRx32gItLDBUw0yx5ijflXrEAK0OK0ohHFEqYg+WzF3rz86PoTXcNPkg6A9iA6IsVWr
aqv0pOTP4oV4YSUkXvL+rdqRoaZMlCaNK/chAsoFJ9UischJ43imPugxTSIoDJQzA+ZPjB76LJJ7
KtE/Zl27ZWCLeSlDm03AKKuTst2CK/1PvP6XdHlJZs1nvAZmxqQcF5caHXXMB6CMFmqRXotVNcOC
kXa/Btv08K28IP31OhSTUTLPjQ2T5YFpLQysOi6daghXU6vSGXtPbJy1xQ/OY+N9FZKam0YRRqb0
expD/wCiAH+cuPhzSYZ2l+P4YBe1L0VtZ7OyxZVB2C9AXdrkc4qAXJtEfRZN8Mjj3gzcTDVMXI2/
zviqQxK7A8K8btHmX7ex45JIMfe+47jWvP9QCvP/kcbph9ESCIpKloRGXy1jIItA4j3vo0c7LLsw
nEAbyBHWoGGgEsM0dzVc+1ZUC0oizxE4PShJU215Qs25RwY8XRyJPXYi7R4PJkt/lAhlutKAj2nP
n3D/SHinttNEBGdfw7ioTXXqE0WN1MM8a2U7eK4Xp3gxxxmpss1CgWXlsdwaYGBkjDeqBJQMYGjA
xD9z/0op2JX88OVZRSZFwGrY+SOR4KYAuVxTwAedjeve/y4x5RSBMqdyyH5PKKdvgp+8MMLquxz8
q1MBe/lO0V++57ESL5d6C/Ce+LBl1rekG4mVYZOs+9sg0S+Xr2+BqdO2FvgdDx5mF65yHqlHMMEE
MBTb/fZotJUROWCyA51J5hPCPlq2prHAYB71Shi8QbyUCgIjSjC5nzlkFh2IrZjGtTh60INAru+9
BdwwW+Cw2AAbQt90lZLC5P5xJbPdULS6MwsubMvPatWQXXR9082QLI5SptkoCsA1EcxxpDsUzk0+
WrVN2k7BI/Z/BTu/vziBO0nSMcWq3C1MH4NCmw8Ip7dttz0GFCEi9vVFj8onh1UEA4KQ8qCDThvN
kUBarPdHrd6EUXJJzyQYjZESLIiM4moVLlMaimTREY2xtWxa2X+XXrQKTPesQBds2Pfolxb41jab
mD9HpIanoaI/dhoGbBMeNYi5v4erG7oiNktB4CT1T4kPWVSb4/1E7ijkZLqB9Je3b16Pxx1ttGLa
z/s8OstUH/2nl/gJrgSd+wjrdISFMZCGre1OHm6uwTVMeYgRJNsUwZo2YFx7zBEW2Th+kpMqZI63
82F83J7zztq4clplAH7WEq8TxoP32T2/EUOurObGopE7fPueKM6V72XwEF6lt1YxMRFGhahITzi4
IEge15orI/lLmMCebFkQ6ahu266BKHBK/blTf0AlrMVsNxQFUEmymSEGO6bygWzpSyd/rVfsEAvc
PP26kjcjuThWFG3vOuSpcHC2iE5Uq1dFSfpD+ojOO+SmcwKi8xdJ6Yvr5g4xGsV30TI9G8acxS5x
rg+cbfdU7Lpa3Lsoex6uh88LYL+EwiFOWwRxoM6g5GQ5ioBLFxDbILlF9jzhhHbbMkwCGzAdspNc
unrrdX8sYvUd3dJhbqE4S01Z7A7A+mSaFgbfZmiA7/cmELnC1IMhhonVJ6A+xFeclkaXjfhpyHoq
rfTeF9/vR7DGB6R8EVkxFFwebL8wJ+s2/AhnKzaUFb5kDYOTdjnYAqL4b3wrDLe4KW6t24LOFcrh
hSU/I02ZmR5ex8EChxcvjEBQx0hmrVQl/Wk5LLEOj7u5RBy1wlJKNxANCfTDsGp/r5nWoMqhSZpc
97ew2Q0vHNpNrSCmRrFSxMAp5KqS2ohUOOewox9qlJcpZnIJqIe+enc8qVqZwGeT5DmTjM613iUq
jxFVGtGgppM74DBACdqFWd5nt2RwGJhvUop4NtXg3NullrItCs6vk7+UyD9RFDodFebptV6ALaUr
HoD4IWvkJTnL2Ogx3jCCZU6TT06kB6cmCJKCSuX4mRRinLHZtB9ofapAw9Yj4uPu1W1CLZoqHQVt
0AOAux77pT8mfNPNsRRO/QCBFVM/1bo/rbwFo6biwWUpiSwPk0o1ud81UXqvQFOWSn3bJX+fzU6s
jCR97T9KAGSvWLjFoHRha5CSnzVDJ9qjh5jiln4V8LbPnrG7BNTt+GlTiCyN9x5XXzi3uhNf3arm
VBe4OS1T/Nux/SJN/d2ICTT6QAbGm1/bqoRRyfScad0Ud6APdLzcJlhwo/9W4geClPBMERxxEu0E
xePRLCCEBvUIggqmhKPLaQJulXqnG3SuFGfbOLkkBImKBmhCrUwOB0/dT7Z/UxPbLS3OJ3yIgqUA
jsDjXY1/KHgVLicHi4Ngfz+v3fQo8oy0NzWNRYxVk5hiQBanF6tn2KoG2a994RFh6QwO2YKwpUtW
W8y3qv+ezVg5wmfBmr/4v5h9eShkNV+MDJKZt0yi05/vFdehkGx/MKbr39CWuwJLuWUmoaHjYTwn
yZJoh19Hk0/65KUTM7wdOgyEAVg0UDQdrZCWLNwmrJbsX+jd5h9derPvE0XtFQ7J1F4cXfnZtJTR
aCykHpklIlgvZfQY9CML47wdNs821XJ+phsWNF71Dozt764CAIvRoyAWucdNftivnOQ5zLXgIxC7
+5L1JuC5s/pTN45VP8p/EibiK7RQ+UKh16nRaOtY8Tokn1CTRO502aohwV11eX4cpu4HVYMdLiks
KbDjpt2t1ftf1AmS5+Z3UscbA17Ij3OCwfclfZqJXD9XMphnLovG6/eV/67kMHRok1khPLRZV9uy
IRTFVMZW2XdreR5gT0zlv+ZCrOVyYgEGEE+OoGBcfRex7qx1E5UfUIyDSNqFlMq8trnwEp+IR+Y3
yH9HPpIh5BPOuiH36VzzGsIAF1pJBgf7vvvr/1TphVXzYaVLLlj6A/HkjZt7qAsj5Nrd8XtGqvGw
0v97YXL3MdGi+LBJhB4d7FE5c5740Wvj16H4L8tZcZAMZ6QdVgqnDNruqJzRfV3kIH8eC967rDyX
ywJAqt+4v4ZB4fOiMW2I4SEYasNX6pOKX+l/vhDqnSeyMor456V1pGsCJpAnBdqY26FGGwg1XBeY
Utefc0lRu3XaRLZ2zXGUmaBKX8ksub/u1QUhi1fE4cg0RxNmGeHezXv8ZgWgbCayz78/4fBe9L7x
MQfY40XRTL6TRFlpgf1yGrGaenjR8j0UrjPQoz3YOq/eY9bs3wqXLXn69crLCU8YsHEjGx8oKbhK
EYFKzKnQ1OGqfa0QKy2U+WcYF48X1aY42vHV44aiL99jZ8kO6vo2gTzxs8e3s0ELdq5n/IzuMSAM
meBlYsV+jy2Kz1vKnhQyXa+qleopAXvxXpISRVGcLayCaAmIgs2NNLWnaqh40/G2g1FMlPoUZkUf
edgOX5I2fQvVXCXofIEl9eSHThEzuIg5G/qurnF6ST8kxU+gD79FDW0FRIkpf5bG/6GoVF20gAoZ
pfp47YO/S3rJl4omE8DUpJza7eEysim3thINI2unnJEW8W+qd5rD2tfJdKJ55uK+5PXH06AjxEpK
ELwZlr9R2ugBOSie23ic5x2gEAgtLC5NBuwUJndCZf6Ej6hcx85iQFA91Cn3pYH4W43AjqGx9Bw2
fKle7gI89P9DPrbIzdCs75TJIMaeatoV5HTIY2fbrl0T7GTjLrVRaQluE1QUM9e+6QVzPNVh63ps
cJKEDtuq2Ar84nDAYKQrwoAF2AkNwIoUA/S+nBZn2oNemOHSg8ETXXjImR9i3kAtN67pCFWUSPoF
SMNO4m0pn5iitZz2zB2+VAb2YbmB0oGHFniCZ6CL/w+/c/Ugqo58gCJF8G5AcpXL9sDqlOx7ebPL
ZOTQHfkDva2o9gqthsnIbAOFG0H1JEHiIz+p+2io72j6RO2bQpEwLwokTcrsV1QhMxpwTIvnOX/t
H+5YlgXttKbHpa1XzF1xwlDB6lWq6SgfUPyszq3KcxAjrQYoqGB9snPJdR8WVrMWRch9OxYORPPa
oJ3/krTZr9WRuNqvcHjVWQxm/yZFM+Nqn21plFQU6InOr3DjQS6d0WyZhnXmcPJDqkv8vwEmUzKI
rfr5xhnzXPzRKLqj14MXUu50aSTMU4Lz7egk90Z2gzQBClT51BqW468WnKV4RkSGfIFLSZrisr3d
CCxJInPom9sTW9rKHufhpsxxnzFLeZR9XGsYkVPrNK26TO7xLIXipgOhNOqbih6gGmCyhPowoylc
vJzsRQ+2YQClhUQ/lOOVfKu+0qEYhXQbf8fh5scom3QMC1B0qhvs1vrN/VKRI7JvTgZDNPBde1TR
3Swws+lpnwz6BxL6s+sBAVNFqVZHFChh+8ojbf41CEgGmm2Qj+fmRp7HLK7yKp6hZlkuibxWK2bY
wpuwNTwLvtNPtnaG7fFgofnOpU+Q13I05FaU/j1aquzHWIVqRrsgnbXirtP4KnzRJAP05951pMtv
v0P0kMtuEy0kzrxSrPn4sAXBKBZhvflNhgrNY6IKgKoYhgQXyc2kd7tr/1xwC4nP4OhzlvSXS0Me
MrOAF6116112diXnqHooDrVXcnf9G7sdZCU4xxtbK2+9Sdx4XXdKt3uD4moeCww4hQNVuNCMCtsS
jXgpEa5x/fe8SWPMpTPHTZ/kkhDvmNLsWLHqlOaBpqS0aLpbAPPj7FDgwS0UArq9Sw5hRAv3xr/G
dqhr+Sbo/jk6n1ZAGca/d4nq0HsC1htsiB9QoFOCU9FHOM57WqWsFZwJKd83JN6RKwYH3jKOzSTn
RZS+lNKNJQhyL5OCGEUeBDbqpXv3zXpGFlIVAp0eE6NBN0OUoia4OIpe7Hdjl5NbtG8uvpEKdgdT
MBCnIL08cFRYlgnmjBnmX2knRtpn4/QACdGckcVCAznVkHvd8UBzlkcaCKqJOuvTisPRoaJVpvAc
nL0TXbY6nEhxO8ewObXUzCV84E+XWE2bZULLW+ziCY6wTsyOegDJwDSpKlQuEZyo95LHbHbPBcuh
dhIZUP6wawFZPaXd+NhSBlGXgEdwBAgGX+Z9OoWbf+cHGjt1yxGHNMFsE0Bkb+T2+j1+MJy0yZJl
fXYf7RtAyZW8IgMiNhegPWXIaKTo2fdPnPnzg3y0LVdTPLR0VQvboB4i5oIUo+gNTVwAzPvx9HMg
IUWrzKVLKtABSbHRV5ond4X4VoCjdLn6D8jOzYBKom/ZJyz+pJoE8FEZFJBWtFaEfBdcCr/TN68T
1KRdxYjfBS6wdMte+/a310I1gCxuhTtmtL+bfrtf3CiSTiHywtQVxNNjWO+b22Kh1K5ZuW8R0jbu
YHa/IjL8BzQ8ziCwSIQFvK3EtbO/zG8g33WfuDnw9lOcRnjEC/FQUO6JXcUpluIEzSEPT33BExek
eZxyc3NyzVMQlxBVKN0J4Pt425MDQ6wrlqrUlLJayR/cysYMPpEIQfw9XWk4cCRAkpU3ybcVjhgr
qrj4hLRH/bM0qW4qjwSj26pwkbllPajRF61Y+1prW3hc1SfFYIwT47HxHO+kkPU+QqZw4vg/geuY
6DjgS4h4HUrROcYzjMJo/F4eWCsuBY01hU0cUzB+LOb1YFJf1VDx4eiTcQD8kgyzxTmxVI2m01Co
Bqfjw4I82IzS+UTY7qF4Pt+J3KpLPQyWA+0l5OFBZZTW8JcunZ2MrMli3VLdlCDYle/ut5wHYV0F
UFdUnFoKe+wFP98YYO6Qv7UXhNYvpp6wO3M50gs6xDXvK8tUD0kHnahrLUuwTcuazaW2W6FWf5Y4
KohnX5ng+iRH0GuCF2ZESKoTYu8z3o8dfwgkhCP0G3T3uu7dMjAijmwjc3feNg9sY3JtOSEVz0/V
uLQA1z6Q/KG0CxOKYr8Rm2MDiU0LjB4EdXrehKXqV1lhtvTik/jTESotVqk7vIG+KbkUn426vvfN
vWfJJu6wbSF5Z1Jw1A66/ItvHWDx/qG+eykVFOYCoKnctmWSJ8jidhPIol6kNLGnnpeamyWB5Aon
kyc2iVKgtcmssIOrLBVpJHB5JGQsMPxKOELiH9/EPCN0+h3FrrSihbQuz7JcX/U413rEQXk08TKv
9a+Jbt+QwSriGf4NfnoBahKvph8LgDr/b6X0NQ4RkrgPf8l5nkU7r1HdNORyTpEy0FtEpUpAknCP
Pr/PR5q1LY4h1TGOhixKieUqjbj550r/xc22NpAkGYpZJ744hbJ/xfAMzHit8TIj7rPuwIY3VU4p
MnPEUZdmAQ13OgC1XQoeSNBTKd6RDop/WuGl7V3VVUnFdx5Hed6DdTx3ir9NzgOWMHYxoNBxUCfu
P6fe1Zuld3mT3R8bzu4DuMohofq3fTHrQPykuJjw+EY2NpKypmRyPeU9AafrPQ6aI7gfnzkVT0v0
YlwoQ2Qw5ZKlCo8djcr5sgfivVVFASKkk9e4Cno9oQ5TvrrLRksAdgtCkVVWob/mHuDQjgokWr5T
VQ5s04jQ03YB2AT1LrNb7Zvm+NasRKI73y6yyo41rfrEWX5WRjkoSeG+CPR5VQI+R4N9U83ugWpF
Xnb9GbyzmHEwfOqrNelLiTPX2PuCmRrCZjZkpqcDqMjy3WRyDlxM/9Q8/+e02z/sIjLMjwbUP06T
5/rc41xX7xBMBE4dsGucomMblsnlOkA65n233/2ItYJPcKhKU8oJd9mKzM4Rw1XmTsJbxXrXtQ2X
dJGUf6EBlFzsHXY92KWpihQGrogjwDDCO/afL77JPlpOEuYd5OqwgS3poYbp3r2d395zwRtAwcw9
0gti4xesFO6KYYnmJlS/Q41PBTXe/MPnlWW4lnesjbxYfHim5hDlcqOUTBhIbfJRsHeA0i/F/5pF
ifyZFNuCdNVSlWDv8azG1mf7Fd7kl0GRqKN2uM+5I+jXB1TWDlXP9WcmoKn0nlcZp+/XKp1EKShc
YW5sGjuSWneXvQGf2r82ydi8kRG0SqsQ4uKl+FvUaq0We4w5VRO17qWGbi3k8vokt+JB4dih7XD9
Z2mzyGAYk4wE8Et96ySGkN0ddo3F7sOuJWpqmPoJJiAjsf8albDYREinVB2s0ta4hwBlKkLcgjzQ
zdq8DUr0j2iuX1fe6Qn9unqGWmw0xSMWcCztzpUSU2JpsBNlAwA5bB9JBNtys9DqgHXOg03r0Nx/
guOmt/K2AHWTqWNP3ifdScKLjsed738rL87fIbKsXH/fz7tI5vCr6S9JLaZNxhqU+CsA3aFqJbjZ
bzsP5oJN6YzMVRVlEP7hk1m63fa5YVuMnEgl4MoOh8pHBWiEShpH3ePcFmHkvuV+q6jn0ipO+Ijb
gxofb9VMN2vNz5lm3eOgHd3sBW7Co6/CP2lK77zHvPU/NqNzfkOCEcy2ZtLa/PHLPZ30p6abJmqS
fwiw/nJrQqNCkopjjxFLj45FsYN9bf6g/oecyK9pI4WPVznxqtE0gq2ySYlkoHV3E5zFW+xXn4RN
urtJOYckwheZmdlupXCyZw4sw7yALKHkzyWcGnZBnea91cw25JweUh5wXVsu2gqQTBMDZK8Y4lwR
0QRNPMZYzkp1zt+R1pdrYIXX14LjCoAdbgs9rzBCSxdqKeh7lP2DRp6XUaJuCamiN3wQzE4G7zUS
ZbCmt6agjTzkCsjvy0FL5tP7xkOXH0jLQKwjlTYnwINC6JXNyIFt1ZoM5AtbREw4m9p9BOgrLQBC
Vd0ukC94wj4HzCsRqE14gogyLSAMP2qVVLlYe+mp8PYa1W07ihc4F7KVQNU1j9YvDfBHcjB2Sa8N
V5DCAlLQt8cZP3/f6IxJTegeL16jXY+7lQUkFiWWJxeUxHJFi2eWLbrUP5M2MrJK99WJ/omfyjAW
McA6zUemECoqTUbP/hiuI/q+8SmrdgPgOU/YJBG3jgteYsnCmdtyzHprPhTg3AE8B1uTD8jwDg7P
uAdDaSgvepk2Znvi3I/jIiSjUxGCqwyTBXzgmVHtEfPMuIe9zuArKQw8WOcp27wU8h2dvKHSbF/f
WaT01Ga+zKc37GsWqiMlL0ZnTB97XHc8LJQp3bM5yYxd+r4pELUE4b5C91nXK3IzY9BDTe9r01IT
CyVrN6jfhWL8J0W/VU6TYdoKoMTQQ4EOpOS4zFGG0/YNqhd/TBzxnxsXubwVuRLr3BbB9upuW4oJ
pDUJrt3V1KIUNNL3hGLCWnuYXaJH+LpHBfKDvXjBo5IleeSYMRuToweE4VdhBJJU2YeGxm0hxyjS
AwAyOdiUGPLaVX3JLNCj2CzctZz2Bj63rDib4ab4allyXuG2Sgp66mFo69zCdp7SH3880wToOwYY
SE/YIV3lWIdN7PL9HUCN0MewKTS3dUVHBabqp4D/AhkkUr6FMNE/CiQ80a/YQrxVVZpQGBUyOEDX
fKH9FMoEb1eU5GlBo/He+aMF0VOdLZFbCTcHx9Jlk4Aq3r9rwvCr19xWEm9eghkSOLHKmDdLF9Yu
SBxlv7YQ6/TA1KiLuuDjbIZp001H2SYh1qu9Ag702wqgPNHwvSJ1vq7k7tAQC+JlCfznwiwaG2S9
O1b4vL3+/ppUGYLhZtqMrIm2gBjNSqDusElEE9CdoU42KeJGU2DOXje4xIZotLHLvC+rS7xvUU4O
3Dbv+H0I/uENnkbCi4kxqEm35kPP79X95EXixRrLKcSmuDK5MsqB6JuF98+eGAWTUqEuvRFch8e3
fDTcseuus6fAAra+E7kP5smDH2AvcLD8OSMxnwlu6qZdjd5tdh2SUwY2TAlC5+TbyDeq0/a5DDY1
2T37cXcYrkabJOocjrc0rj0OyA6UVvp3v3JguWBmz3aT9A9Svtk3ggQflUcRG2aVsB98+/h7h5Ih
UE7k8dyitwys1vxdJe/hGuBXcAV8SHqqyjt7/aVAsd1G4j3LSD4AGq07wfJYxXP+QRglbQTiCmtA
Nelb5bOd0vHrmirEVd3+qh3ujwKfMTijEao7MVcFUVSXxYP/rMJeFhGyEOuWd/Hvm93O5Fgjwlv9
ohnO81cXOA4+1a7VdAa0XCs6ZtslptIjEYRL2UQoRKItyYz62HSxsrMVcEhsrg8gshrlgK27WqX1
61C5nX3mwDBEAF63hdS9PzWJT8Tgeq4ao3BbCEW6WmcIHP+dlZD7smam1SXKpGFptwOJyaJ1LdrI
3iUFTxFfTrSEkA2x9BbdHyewPeKQ+5OY4L0gGZ1oGZ9O9aYzWZfpePknvqgdeMu1Eh8OJnk/LMy9
VlEosOOVAz6iCn0k7GbC6/G7MR/QTdUpitvXdYW9fSxrg77qtVcEEiNC8os2vMK41NgkN+tUjLRG
MnoEZud+ShTdo/TXYLB4yRZA8aV/KvuQmR+VKT0AumKZ5gOJQx8+QytmK4tvx19OaSlcNqn7XiGM
4kgZlPlUR54Hv4ZiD0f3C4BfPVw4NjFhU9hw47uAHhOCwrRh/4VI6x1HbaW4Df9J8iNk3TKPNNaL
ZGsRdBGqo+M6fmFUCbvoAMuHO4PI1UiOLqyuboUtr2+Yz58BKQRusf988KG3Z1Lh986PrU+tNnxD
CDN+zM++31e4cVnMl9/6plILKAfglioZj/lDqE3NAwgLbsaRRAnZtpt2ph4nGCZXw7iY2vLdXJKx
4HAUQLc8xStNi5iiYyL/fHISxGCaJqTgClNX1q+A8KyW5ruAz/Ln/grk3qJa739HICXqpD+gz49i
W3l90mN4wEmRhyK1yF5NQuvRySOTYLYiHDtO/suGVbOK/5oN7VD5PI3gYRWtbrqLw1KTxtYDFvlm
cMxVC+cVFkSCFwbFdpjK4O0OrA58F+mmdKxnNBr4pdp/9tlLnD+ZsEFuUo+bQTf6e/EMjt9EGxk2
bmhGTpKQwmiJhq1956H+qNsYadeSzBoCR4y6WAzaOyRQa2bMshOAuG9hbwE18Pg6JwtlrF68zjU4
72mOQ/WiU2KvXvjwems7uUmBQ+ADCozYc3lH5C9TFwe7HfETgB79ytI1Kehu7r1tgiu6Fr+bn3w+
3a4ZM5h9E7G2N1v+R68a7X2cLWxwX5IVIJVmX5EaYtATzhNqbuf/zI01vwsBycW2+3gmSZ3ui5g5
fwB7eSk71NQVTrkohn2wR1iPL4phW4LpBLReHHMlyMHLQp+bhtlLltite6X53dXF2n5v6Hqt+D0F
n9i/pcaqqWsy1f+/kFEyWmBJ9GetYCM8VS5fNvBg+2N2VqsfkD5OT9vQLpv2lFDKz3DAQypty1w7
NJWrXxx/Y8haGtYQMdpIwFr+Fcgtj1sPP02MDOE7+aTxYyjer1UXTDlC4wjocQo5gRoWA6Juokbu
33iGpnrKrPjuikiXZq8dNEbRf0k4gppChaHoxF43rRtRBizdGw9QGzEHmhrBJm7Tt4cQjNVm9RZy
i1JRLbbbNvWKMKbOpM0/wBuBHoIBY8AsyHUndyIqAWPq5JI6m1rQy3Wf9E8kGM0KN/SikTGwtpkX
+f92koxBEuzZMKhfXAAvuMZkMxBXwPsIL1ezKTcZsR4ZM1jk183VtvD14ir+YEZJTF5j2bU3x0We
fNQqO5rMccX1STgoh7GkpLlDFb/P2wK672a9rwwKmuXMOj+od875FPuvy72XF8GgPrTU+hWsy/Q4
xpxLNfQ0cK3spdVECOe0aW7IHrMx98ENYBlNAU8b6+u92W0zqaS5ZgAEpokHuiQlf2ap1Hqy8mfR
jrz670Xn/ukEyBe6k2OLaucVF37uatRUmS8NSe4nyshbAij1r0VieoIFEwllQuGJYZqab2FMFG63
tG4q6vZyVhDtgMLIILnCRGIgdd6DbkepAkQX6u46qcBw/60iVSUe/YkfFbYF38gHaJ4HsqSF00WD
kTO/PpIOM1lKYZEZ3cZ5MBJIMZ8yQ75LAKKVopAT1YdSbQrNOzuoLmBgzseGT8PZv6tEshF41Iey
k0nlGjpmpAjQ45FjZLKofT0u/gfYlPqxs45Pjz1q4f6CSrLLfXxa0uKbxRo0KHwi7IpfWaGJyJ+j
n1A+1/i2ug7MXP+lX/FRbCS8n3xtRK8rSvum6xTB11Khj7+I7c14O0OJcLkwZIE8r+U+ad+xOyP9
EhYSvNs5n9K0/0AHS7txk3GXc/hmMcSNfrY+vKCRt0cMKE1epNHT36ulydjPJ4Fa4RA7oQ2eoH3N
q2xniMRVyImy8y4x0IePs/Mp0eC5kKktaLUOrSWasgU1J5dgR3Qx44G421I+oZNDNRmNFJNFW34g
fhkg+umrR6J+uoSUt0jE39RACH2xnWv7y5J8ylHgYrbSW3d58UiBhZnUJz6Fb8yDplgK6QbMWhdf
O5yWDcIQgQBIL43QToTQUDqi+VDIDJ/XnIfRwrOPu+yJ2NjgulcXesItvbNx2DXn3Hf1uDpxFyRp
UipT5rxTfiGTRTwJdo+Qz4AXrLlbk2aOG1v1XlE87C/+hGoCI+r9InU0MRJqR4D6V4OG5SkaytF9
njEJ9NmQdSqKbmayJVjDokVSOchvegbKsrz2rPAZkKfRY2FMHu05QpEA42/1GbZ7vZImFMuyEyAx
e8KQuXN9ZPwZySXci2g8tO5zvDYfyvxw944Drl8sgWpjCr7Ms/EWx84lES5dxmKqVQexTrvhSor3
snQogqUrSvKY7mI1Id/lCiySF2aNCKSxFapmiMzgsMj13+xYa+3Ys9TXI3XOdo9qSoC3GcvXsGl0
fjMoRvxa76oJMlGZs0ZLaRZFAD7lY4Mjqds9gYcT2EMkiD2ZeottymZtKZcmRA3EnDob4+AT1618
z0mRcqemkW+W/GM3IFR1AGwkCIhdDA0N3uqj3Mq4JAAJoZJWyHKK4eKAYQYuBf0yfEf16x9gblqr
ASSluDoq2B/LVaRd8JQvITdfGAdu9rfLgP2am/XA3IsZXLoGGI5LNtSu/kZ7LYPzJZkz8Ua0XimZ
v7qZ1Me5MEwRADlBK4HkuZm18pXDRC2YtrhIxinysdqjIIX17TyOqljAHGKjAVHMXoqWQx9e0p0k
J5Bf9AvPvoi5F+LrkJDKES2VVJh0HtVdAJt3ynX8Kf/81PKTqIhxXMri4TJXAukRhSP4P8Yjmliq
KpjwSw/tvTqi8ZJ3HNSRTOqe1y+UKO/+U3PjFmn4xPQBjvGqyS6WRgl/Yahg4+s3KuCyS842R9qu
5PTyL6ATd/SqVsPHv8eO0cVJEVQUGO9b94RVA7RKNj9nn4thAD7pWY4fq27ra/T0smVWNnfa2Idl
v1nM95NnB/5AAw6gtQDEhiJ4GQSOFKJwe1t1oBINqRrubb3Jglq1bxCK0a1zdpLxa+8Co88nLZMT
1oR8F9/ufk2SlsddfcFGMlE9BA3ZCPtpI7NUX2GgpFOQYfRDPYtKJMDCG77MIKlH3xvi0By3KI1u
5T74vdznbcZFVfXXi0wK9ZD3koQz7WbtjhDqxKhXCLkM+fy0XHPtQq8vhFooTnLzsj1+mwVjGUar
r7DUNRDFPo70tDbPXRtyT+mN3p0yAX/cbJ4PBLj4G9hCGnF1dV27p1xJbQBFEhHSisCWzy7s12L5
OvXW9QNWSPaGz840EXmjkRyAuOXZhJqIn1Lqak87nAlekHeAA58vEBdX5sKWdxxX670HJ45YPKqr
li1F1SB2ptmpJGBQtFeG47+TsMAxG8wu7BFeYsf0Ej1Bm86qRi3QenVtFhIwFM/LezanYDl5ZdPN
7EVaZJ3ezy1659DO995W9doB1HoZvec74/Dfq8HjXCUKzHOP+vbqSyuK85bKXZQv0YkvfNMT6cU0
55B6okXqEPX7xh2V7MhAE5EP55bY2ITdN3cpCy01+sVFrni3R4kq5KjxtXnSnDM9W053RXZBrgsM
XaSEJlzkbaSooe37z4CjgNgDqwzsec9eHSOYGhkvPMdMnfzXgHAEJZ7aS6SICscPfXedyJphlamn
MYRyHVX0Yy1f0dapKYh8jbKe7/gIhOOG06VuWGxJx2pSlljuhaCBxBO9AmjnuOpbNLUlHoSME3q1
LXME1Z2q0AC8Cm+Etq6++1LOlAFaveAMsii8u8Ba02kiR6YXYk64gxs7wqyl0Tlw6SxxI3jKaCu+
mdIZaSt1HudEZZJ78nWGT2Vx9AK9zji4twrMXOYfwYFJdyAjyz3cvgjgfndLBk8Id0hH0HW/RZGE
55lJ+TN0wcNGXhatmqnsBGIftcFAYFUM8VDyPJQSPXWXu5xPt3Qxt6IHXZWjIhkDsGt3OAEuZidH
YturyxzP1khap4HyjzfbeSP/NkSczN/gVvZFGJXjUlcYigSjROXkEN675lokRAa5d6v846gvPl4T
8stqbIg9H1aqeLiQwkag5RV94K4w3MuIJ3fK9x2PI41jaR4swG6h1QoCHF+hTHKyASyVr3C2m/rQ
PtrLpsUKk0q9q3TCAYOkgNmWmWl0c57HQIBe48rYhbeCp4KHp6vCEpUUggtq+6bTWBNgIB1U3wiE
QnBc5qs0jR+W7qyBXSvd+20q3c2mVudtDGzXoZjlzwYmqfrwDmboOYAebB7FmzUSrw007VP/PtrC
ClrQUVKorb9z0Vm5gnFfR9e3FlccZJu4t5ExuWEnps4H1dx/JzdWQ0Zqg1O7In7k+TV8p8ez+Sfe
L+8zrvDB2wB+uJ97k+xnvPqePU1tbKf4AEBiodxQIzVBLqDqlJ8dMKe4TuUC+JzfMpIpWVBVza48
ty9H1aQ2TCyE1hHAhuOovaXtmuXa0lTEsBRh8TJXVpIRVBptkdf47qw3jYumJD1hnXYDup4lD01q
Rz3EZ3fRKofVFBhn1xK41xBCbzZoePKghP3OQzttR6rCwdbi9P0eCNex5m9g8PCv4JyOyvRj2bTQ
81QbeRiRpI9KqUcP5o8Yprbv+n8HMVupaLQQZYsBg4ZkomhMbWL9AGp+lPSi/suGt+pofji/MUph
bYzdpKjaHagnQO1Jenfms7bEpsmIRDUF0m2nLL7Btbp4LoaDU1xzG+s/uwsfPjTB93lCwDFkUWqB
1n3BUCV/4U27BqEKI8amIqp8yJVhQs/E1lHOuE/Ek1iDBY81sCIAYy3euYv9zi8nsHhdChSo6ZMG
Dg9vKpUYLbMO/P6OQISQ/Vhm0g8nA4aRmH3hmSqkLUJz+Fcd43vTfBaE41Le7fxqtVaN4EAMN7zB
aEbFvpdQJE/8sdHGUi+/ask4bSYqSHU/v/abc2oLCnWFKJSug8JlGMKhm7Y3GMyb8Nw4eJudDQUr
1BH94SLrgi751/n4kxsTw94D6Z9der+c1TzgvquQf7Xw39vq6lBjQxWnxl+M/cNGvcbIqnDTnMW3
kfYWeNIQi4a/XKEBz6dxEyL6sD1jtJqpfxLLhvI6oKsd3DyoDcg7K53Xdr1PV7vJqXOlz4S9r0Un
A4dPp5AUUv5PJjqWPRUC4GY2+YHHz6lbPVSsKWBNzfl4XzqVcWkGoP631ssSIWrFLeJYszcIlKOM
qGGOTQpnmbrej8EbqkMdxLcQyrX/Ca1n8lOu+usQIJYax9y9KPDLTgYCaHeLioHEekObmD7sHiE9
cFCXRkrvgOXIZe85dNfX5LrTpxnYEm2zYw/YIiXbZDmUW0PkyGJYs2HZRbXrwGE8vK1D5uX5+ysX
A91SEtFaSwQqDjuwDTcyA52ViHkrurdVUu6/k8RxiUmDvY4o4q9726q+Y7/n+mJL12GnBv4s2Ng0
sDQKl+I8qdSIAyZTOR6dvfrTzyeZPQDoA89M78RKH2lw2G1jpBa5I+Gl2i0DgBUxOxRA2wWJTjWl
syTCHfJBIj5xWS4Hbzbd6nNjehsRDC2aFwEj086+GF2TrNIapgEAQgUt2U6i1NEWX1wC8TmZn2up
1Panl6ckEaYusVGSfRo3hbrJ1+r7sd44sVI33YjHm7OhHzAvuruOzxcMu8ASWM1T6Sb/1Rj/49N+
RYYd8FfHDm/NSe7M8a/FOSin5CG+CBmdxHiwTJocvD06O4yMXtoVxmrE1PzL8Ve/n4oaYJY349J2
eiyrV3L2O1DYkjVrv4Dn4/DSGfR9f2/tEJBVeMPiZby7/zLN1eNm64udd9TglTZPx6IZlzThryGA
yGAYSbqs3lxJ8VJT7Em/MJTO87MkXN0fnyR0hl2AeL/an099dC13TbpmDXK97TBSJa2V1zB1r7jr
/FP8q4P8FDXcgHcF2lpbBbFvKXXpkPDLmbbnaWidFlrCcOuBt6N0+xME/ZXlGCZF8mqm7AuaF8aG
1KvwXO7CjsfIKqc5HilEtuNLDXcKm/5ehVZLSWQdl0wMW+l+QPCnlCSK6NkqUm4Sv1wzfWK++wCN
mB+r8E3S06nDSErKWXsQn13WBxIHI0ZLybveHmbTJGknCqwLl74WY1bWX9iWxmiLEPgDNq8p8GO1
kAXSEHDhr4zNI6VNGGZCnJQ6AOHgUFAoWHThVcmKKcoibNvEoAdELQtJ7vS9bBnSP14mkUOJf014
h2zMlFRXeX2ByFt4F2NWAQECsqeKjXVmotRMKSAguqy7yLkTaN/YskH3JGOR4VWuh2XvwXGLQLIE
eC+ybFj2Ip4XdJ+b3CnYPyP0WQo52aP+kkqTCPz4p8EjttPqQ/UH358wFL6AxQWrJw40xuzc7oNm
Ob7Cc2ZeOFcbnMxUu3u8nBXWm4rO+aaLulB1uTiJRhmX9UJJ4XAbQ+exD7U+/CvNQUdfyNfnWZgF
SmWyaS0DciCKCrkBJXHk3Ia7b557slxYdodX9jwINsyZU10OOOwma3mgG8nj8TH5X1hCzVbdeW9W
Kg4JwsY255Wnox7y4wSeBKomFiErw4Qk7e2/GauTmG2cg2NjwjgHkQd2N8D0XzFIp0/OaQrK7cH+
MLCQ8eG4u6vdQzG0wcto7H7D66y5SQkNZa9LJARqnHjsVZ9/jwk1+97bWPz9znazvsneQxq0Ex94
2Uyx38UKFpYGV/mcTm8Bokk9MLO4VlPhTaSsBL3c1xSaX/9tySYpzqVu1yb/xFnh44MbWHE0bqwB
osNvB5eAV+J4jHHBEQCZwPcmmkCcD8EmGdWU2pZ2oHGsXPUro++DNEPyuazHyJnOjjf1P5jBHwly
mpa3zDzd9Lb1mp0W2pGyeLYzpRZAm5rpYUkZ4kiLpxTA5k09YBDAW5b4cpVTP/e9wUp7b937rFkE
Q7Pago/KSRf1aaBpGMkHjh7tXjmCwcu3GyGD5i8JjNXTyLJSc6Nlt81bi5jBLGqkNGu/O0fSUrJu
Vv4aN63XXazjzmR5qfxDizWcO0BQ696fNFYx83OhnXvy4fuQlH2SFgVjLmoGtaSC0bGyTVGjUJgL
HBNwBsVEBNTZCIgTTvOJoRhnEzDS0Pn9UNeUDi67Q/1jH7gpnYcZXM9s1PGKY/KSUJd3CTKWN4Z6
dCpIqneqTbR/vzz3/FaBWby1dVDoxvTMQ2jks43CrsHDCXCtebkP8zZ3ffGaudRWrqZ4l5S0ggxB
CNexjNWMFPlpU7v63ih1Jq7uOo1xhnc2v0JHu8Bl3uCMbteUghIBX4Kepq3tTDNHq9vajtzha0c9
queOfF3UHYo2CC6HYKXcSy7UjEPBGtEoBU7wVMYjuTL9IIdpqvlFPm2RMfOmxz978JJdU+JpxQGQ
XWRFZW62oh+W78XRy4LEM9OCt3NeuE6nEsqJaMuGT3cI1uCo0BDFvqpFukvai6XTGPLdD+UUn/Of
BR9sdwUcnmdMPwgmha6aann89YOfd2oAdMihDxCFX8JY4REdrqDvCZoAj4VpQeKmarlz86dUjL9w
CZl/BiJ0lX5qprvDHDYjafg6m/iGpmQoHXz5uTp2PA1bh56BvMthuEShXurJ6J420HuO0ZZ+W6Uh
UVvmxhhlbzLMyLqXK5Wo7jgzjFytjGlfA+g5H7vEQAtS435St8QbIwMJoyJEQNpnoiGSZi/x8YdO
SBt5KHauX5cAlPfBruIepGBDqitHZW/+nXoT9z26v9ssEY+dNpCABqj4QoVtHX5BuiTj6/gH6SiC
rBMZ2FU+fk9pTZvD6wVxrv/Slorijkzd96VkuARtLyZrKz7MnlVn61QkbEbHJmx3NJQaTC460fJV
xGaRu1kRuEluUTE+PDZHtxqgXk8qZK3hFYfaWACg1Cl+GGQRgOaymCgvdE5ldAz5y/kdK6JaH8TY
F2s3kY5fHBOSMdaw0y5i+m9YUWa1PeUHxeiNjkLOTbDfUxyYGKoYwYYD6YR2rhJYo+NRGZ0gLGBl
C5m+vgBxOcIXosg2wuAjWA/JqjZ42cOoYVO2S/bIC7bkG2n6fmArdfhn26a4roae0EQmBlUYqYf7
XBl/QBwdMUI9RDqzMAdd0gLrX9BomXzc2+VhEhDWmI1Kg5v0952sjTCgcU0d3THym8qAza1RM5cp
0U9KIEwvDLZ74Ypv3rFwPtPGi6CTSGpCR7Xa8HvwG5HLTiAuVoKLRyVMB90o62IBoyATwJgW2gPW
Wr4vUGeBAQ9Uw5W7a5Jhnn4e4N6DH6VnR92BEt3+8FJI+/0KgVgRUBipK87oJMDZ1aaVCv44RQkq
9CzUK4fOSU8o92uur9PmlD+HB/iRkHV4ZB5AGPv36e0St3KKVIbVVrOM7HQAF/kpmmGw/EjxPyW/
c3dERwQPBJaKLJMFAd0AqVsF3dshRbi32H1roAmpw/8HdqEjyyxNpKPJM3cGpfH+otXSATOKTSy5
q4b9UawbmA5asD0DfBQptvBPaUTeORk+O2CHMpXMg/XBrGT7CCZt0efKNDnp5GeZAMHy8SUji7l6
oO/TAIQhSTOAFxpBoMqPgW/YFREzug0UnuDzYEgE64F4p/Z+sAZjt2ckRmxhhNQPJ77Pl941JNT3
lQ1YyCvme+9FTMTNNm3cwD3htMxaXCnc5T210iPewVBnyB80Ous5scW4vjigoXaf1nm12xviDC8C
+IcdFIlsBhEHaY4LmksiOlUCgEdtPh1s77PM9YDx4GzhZWKd/9lN1rB4ivNOnCm/nHVmhyk/ypmM
PYaOQL9eltWAdTbTrJ/GpdAYzhDz06CTEQFH7vpgg/1ubGIyc8K4zcBj89HiCISdXB86lPm+g8pl
7CiJk8MvG6QK4xLap7p5VVXOr35LDgwwGT3e+Vqme2IZmaT72wB5KEcYx4UmtF2Dvhbfiy7ykZIB
/IzZyGRwKqfxUTCqFtCBRb+7jp6wUC7QQo5VhofyEWTsYVbUDDQrfN7wvSltwYs05ANqt6JVuDsn
5JvJTlvgR/DSOpLtjxEB+apMcY3T4mBF6L49s3eVMehjFu4EMmuSPXQ2rBAkWg3jNiYQQ2K5Emb7
Z6lQaY3fdpUwRd6DKmsnoan8smwksdXRYXbQkAyEhZwyCBEh1043q+ED1FhUvdQkWAFLjNtG2zWh
qqv5TWytzE/lf2tQX/34EJhH6j2mGx35SbdLH6lvYjnphKBiYLafgUrgfx3EBZZ3gCEd/G2NOzqG
E/I/2D+rtjVfv3xhBcamrykY6lSA0t1WYX5xPZtOr4KjGwW1L8lk4d5IbreZpUM33czJrc5qCAjr
z4l8a+3K75iXXvYhdUDc2gh4foCE6N4T9Gyy5/6dbGo6FGdajR3Q9SxhwPGxNC2PlkC0YTDG8VNz
uh1D/7z3FONT6/gWnyqDo/W+bnx1fVNV1/CJr8ns2e3anVI9bu7B+sCeCyJZizytQ7LHhZvEMJek
WdWEPmHKju56Evp53BqV8qVSC8oY7LMG11iOgS6Wqz/VfcqyEL+RqB3Spaf/wOqss/Squ7vndJmP
wM2wkocAi/tLXHefRG6TzkotarCmv0V83cInE1qUqFc4UqqdE8ufLmxhp6aVr8bpCxO3CdEDX853
cCKz32HiFZ0lAB/YC3o/bAjTds9ygDgYb0RGGjF6agftCBZqce8Rd4AszxccTWmuo5VLv+kiF4n9
R/aZU3J63+w8KVNBcc+Iy8DeeAO+XQHD1uvj4zVGVhT8ER2Sl86zOJq5ofpEvzY+vBuHCUoN2yMc
siRWYHhl/ArnTYhUfyLmiCbtjDxnaHZOi/Iv3F+ATtIz4aZsMvGVS6jGvSsp6q9esjC3iVKLRvYO
28XbJBFdx3yNHVQKJwW6y5UxfCEmMTWdN5TiCDDWOVyYveYSUAVtKeCcORSHvp+FVQC3UYytSqqX
T7HHQ17TF25NzVvVafz6QPEf16n/DT1hQ06BNFgNVBZwEGvWVUPIoDmmBP6ZlUtlCtH/emzDHq02
vVRWiqfxmUbDIYcGZemMFCgdHAcXCniBC5JVD64xXHy2iCu2NjPuevWGZNM5h94a6zCLu2IW8TFU
dSFOtw0Bun/QR0rpKJM/ZUG2Zi/2wa8tng+j+8z/6BwJmLt/LbwOsmEnaRC21ymBcbOlHfYFU6jR
VJktXWouCFmntKy4eh9WmHYL1hYZHSzwgre8AR8RMotF/4+NAzxkXGgJ0r4EE8NH0BEljadpZ2VI
gncNORmz58nst8x5VuNjrzT3guqHORkaFjpKxXdEB1tAnqe+wpB9vNxvp5+GS0CyU3EkfgwFIvI3
iLvJE3OmXfKHCbbfaJFCMTgeM5AJWsWnkClZf3hhlyzG7UHT4EJpfLJg02qlOv8K5AImmO74ZyFx
md2ry/1KrDkxvgYlKH3BUnXRmvXKiSndlnUCgGxTHPqbpfpjZMA1F5zn1CdLAMZbQ6pxbiXOkabP
EL1lqbHkuAp0Gk55eHw9vnsud7pEVkPivM5tzZbPEaNPl17KllovENTILUINV0JmovVqhV3Apm1U
lBSeZp/e+ZIwMAuco6qDmAHRhHzQqM8bm0JzwMrbsxUNLFyjDsg+/PjiS/G3mGDjhg888rCX5+XX
LkF04lVB0TfdqlwNvg/INVdT14zDLuN69OFq9UIMDGguhtmf3sBjxtJZGYDvPj1U2I1xcQwAWUeJ
6Xa95R9QCb5WMoizA1GbtvaeVbrxEzk1AuBAMIsVkg5eqttAy+MuemxSLmo5XiQxTWaF+544ut93
KWZ9vlxuoCD0SE/OzPhVPVga48JiGlmAoN/3Ul9RUEYa+2kL+D4gnAAnTPmvq1T6yPVWofRP1jJE
F4CZHmo46diG3txGfdqYrH1LNFeasQ2iIusNDdd9ss5DxRg2QO64kuIvqvn17Q+AkwtDikKf1sxv
x+z0GZCpiwQV0dZ42QDQS29yPe0VDG7Cr07kjv1/46yhwxBlrKj1dOwcA6JAclMGmBgRrFc5qMRV
0ZtSnFKWvJMqIGqUz4gh8fuDqYw6MJBcaQpFdK76V7fuvlS5U+Qr/SX/HYVjUrXC1gz4U8wukvYf
BS3JH1jblY+PGYio6bztFeB1RYIeOMpc274IAD7tI38f+b3ae5onp1mBlh9FmOynvVic3k/DNpTY
QrqFylR91ivvUfImgEMrLblsQmbbF3Fb9bC8DJU8lLmz/qeRhNgRpg99IZHf8K+mUjFkqfeOgyxw
FJS/HNshyiRFvgsv9Ef8qnYJBIrp/FfGMzuG+aQkFebq/GpAUJxRHpgU6PO7avCpMyBWyPq6d8Io
Uu0wtWc7fOKhi0AD6+FbIOp4VcBRwni93P5yCRdyxzl4aixZzZ1rvHgbpZh5Y8sGZuGG3kt0U/Wn
28LgjaKHcnN8ZaNg0b9cPMj3xPvtdRWfU8DDeR5veJmc6qqzmAiEiqBo2E70f45n1ObX+zD6q/P4
a4om8OOQEQEYvWVVCE7Rb1VS/AZY2j80x65JMceeNkaTCZhv2xYku60rMP2d9V99HRRJzXb1M5MV
7nc85bpe2IXGldo1sfRUJVJbkD/+djVBIYxHoeh0X1iTpd4U9G7qNpaluxQL0WRWkuQk2MKctzLj
xn9toxJHSstySnA8PGkrKQ6PjxWrLnjDb+KfM8ttC7aMg2tx3IyPPbGqSfvc6tGOG6ybhttdV7eO
plkr76/Z/U91Xnil2hYRssbELmNsNlqrg1CUd7pI5lA0BpUwmvD7dPcDo5KnTClI6Gsxad7L+xxa
07/D+eAnRS6egSLV0kQyAWJbh8UCbmTtFIsLnonsfe/BNIFxAiAKz5qiH2Y7CH33mmJjMzQLSsrX
+KdlFx+k7VMfmosZo+0Ye9YAxyP3bq0YKmIYGBv0tYW6eTiKlXXbCOIY/sDhvjOPpN3U/MmKzHnl
4mrur4h50iTPwpcSe9mZXNQbed1OIpovgQjNhmqgmEJWVENoJSR/AD+Spqzhel4NPQHHNdaX7+cy
lN+jdxapSmKTcbLXtbbzDjiaTmCKrP+HKnpnGTPBPysU39+vMtdinZTMlW4YbHVDh16nSlZzhcg7
eJEApQ22yPi4DK3H74lZkiLs1VDFzsutkIVs7FZTB3wem2qwitwoHK/KbTnfnOmXOK3WOriQgGr+
r/wChyPo9fMGANBXITsd6eQ42g+Y/3PQbUq8ZN7ZZzz61bTTvBMTerUyTSBE27IuH3kGvMbkXjoU
P8xk28IMZ+otJDjCvJwSV2mdiZhZZpTn2Ez5xCusWply/9bZXdU6MWZUzHsWVr2M23fqEgOZAnCZ
tfDHc0+Xq9A4fgs28CWqzq+HbNaY4+EcxxQb6hKYrDC72cz3WEq/FKiL7h8d9jMFyttz39l6GiU3
fFhlb5Mw3nJ5OR2NRD/sVi3l32JxgsUDknrWsmJZHUar5WVu+SU3YIWpy6L65z4ondAGeixe41P8
Zv5yohUf9C/xrKXEddycu+prdDLv5UZLejrPCx8nZ6FzdfvksHrFA0nAH/lOLAwgsz2UYBm4rDBh
oT9TnPk+FPydVqUjqRnzmTSvgFc8mEorKr0Dfzy0CYLGslTjXseAUuNJspMWUeSrat72LRkeUFm7
acP460r+eE4wxDPS4KcI2PB9uNCizz++KBj5sJqgTYcmQ4mNrxWyGjm7kmmnGIfrirnVlerwQxPb
Pd5NkJZ+iAH0a8jxF6Z7Dk1AnR+Im1bZIYpFO8d32ruhr7eNigry2NaL/DI/j2i14Sx3ieUaCyiG
stcp6D2+pKM+f4PKgeDzB2DL1CTlSX/x6nuUMhMxymFbSBQXlVwus7peRxYN5ih7GwDDIlnoAdck
Hxq9IrQtUQEoJw1bldqdhwRyVlKv5yLWmUjuTNWInkv+/c5w8aJ35b4xyBBvDz2gpP0PxPgwxgj8
2abhDrYvfe3xx3CbQ1U8n9FUpEsAn0LiKZG+SlHidmlLA8xwvDUjzod0d2NSGi7AE4iHoidx95aj
8VbGX80ZVwDsJGM6Br3rSrYnE5e/3BQ3wnlrYK1AvkFAlN5qgSWuGm/Q95RAxpNpAkENwUkgwBQN
5RgIWnbgRj3J/B1Eq/7cpqjns5stUs7SMw2ZhWLGgBGiNIwv3A+AeB0+Sn+kd3P5SFp0XtL5te2+
kjqe87dAOLBs9T1K7P5l5ne0ghhUSLldhDxIeLPbmjd+RirhqQRiNVV43vxdUoPWgfBxWkhIp0WB
iORqDnB8AGWj3KcHjvVbbqCYq/Y5YL+4yearfmT482vYtM1oeKS6JTWuliZjBAiTbiVdYpZhjr+P
zqWd83R8L3ylr3WaCxDIGpi8kLwYa3V//MdxPj//Xf7ixLXUtzh1X6kIVxGaog/E86YFnkYZEMxr
T1/djJxIRe466ILiex0qwb2xLsV8HTk1OQ6D6cLuWdcGCQBijV7RZR8O4OQDz8MH9mBdVYKfWL/t
tq6XrLxaaZ9uPN8AI8dpkl3pGxayqWBJfAOQLfYFjEmUuAJtOTO11kTNjuUMVWpK71Zk9Fg0xlXM
nNBdTK9kRXNznvVNfYNc3R1uw+6AgtMPMslCqOh2fDTEInWoqfsU3FkvSPjfEGC908YaPtXNGTg5
IK3Cj6zn/PTUd3CLx+A/nn1a3ik5D2oD/vbiqHjyY8Q6KmCTG//zt+o7NVExxzrVntsQpsWo7Xq2
wEhEnuHs+dnfaHG2pHgBh6UqLLTCx7WFj6DZTeMrRBbOfZrGsvFiXMc/keY7DaJVG86nlujT1ySP
vIxvxuJXXVvCpSFbAU3Zl/xYz3HKwwexMCxq0oK9OCYoJgPdDnAy59rhC3vOBv2wZ+nwYITDqGWA
JJddEbbf7w/T+TyZwt9YhaIQqOY3V7fjbOphKbGwOIDOjK/D5zJGb7tOrxMpEjhElanqVFwx5JXF
Cpfet3q+GTQtPnN0ImTc1/1qPU+QvONlfny+5/ZeP6xbJ0bR8IU+hP24yMH42VMoMOq6bWtAw5si
30D+0katcsxU3OONs9ax5Dtzf2nYmmenCk1yuX/2TLOef9P35skvYk0cpMuXnLSkLcuc6uZO99j/
H687qQ4N8T3G7mL6ZhVdYu4AYb48k1MiqNlJsshJUiNVDY60C5MkU+AEEKJJrLaz2BuG9bw98RDK
2EUN4mBZWARMw/12OulcbBGTtcR5CrSyp85vN2POc3ENPyxIhCoWpL2/9QxnT0h5bpX5mSA+FXnv
7Vc7MAAvTmf/Sr5LD7PbZRQViDh6nclMSihDk/fo3nehk8bu4C+ErxYGbh+Dr2X3DW3IopF9OMK6
2GiWaT3uj4zKv+79xUbDNJ1/m6Nl5ZEY0P8CAoxJY2DuFWl9je5bKxstgMSdU/rZO65EGIs3bc0t
uOg1j0sdJJzdihGJiOPjiiICc7z6sOG8LTxNwRXSJoVagy2MLvlLaHCW7QLPNoBSIaxGBuKMItKR
JFwefpaDNNm16sltkc6y2TMkxJv15lnwSeqJyAslfMY06Pluis1RQGwosq6fD4m6qS/kK439igeh
dwqwxnOTuMRWZgWnSbJeKGhPxx4Z5xnvGiCzekRR9DrxL1mucWme9BU0bhRQjYnGpCOX35e/9CCO
UEVsYy6VLhW847s/QAEMwGPMGQTaDg9ijNakFY6lkmqBxhfA2x7z2ZFhKSNpVqmizcmcG7DBaK79
nvgtMimMpS8S9kfcNJUy7CH6oX0nqJYjVQbFjHb4T67LkUOAbj7DX9ZjhiCYHgT0WjM1rCvPyEhY
bxXx7vvwhrihM6oi+nseicnSNnZp2U/5z8/AwWWeM7uiIklkX/qQRekHuuphEyc7Uabg1Z0PMIHG
X/E+zhe+jpurzygGDZRCMJyqMrvc2sieQxVqQXQsb0Jbpr2dfb/EbYJ5cwrff33ntp02qGvy/M2o
A5V5NWAPQggc91lMLj8+WZY6mYoYTFV3yQB06ccXK5zHcyW8mXeU4NblAGnT8lY7fQ0+POC2ANWO
77qk1hYMVaUqGHbPZSv8CuTfv1Ty8TgxBNm07xV0h3cmVl5b9RApbx0Vl0CpVnLSQwXgBtgZEPGn
aSzBOgTy35XNBiEJq2TWxmDb1CJtR+Uss92gAMOkXE1CR0zMjOSUq639BaHWYD7kB72o8MqMchqI
Kzf31gkFnJrZ32lM5w3j7bhdn7OAUlDoJ+M71LNnSHllZFmzaLBrtvX3GwxkEkdOeBaWbbcSCIWj
zgucYfPxIZMIQPxfjc1OL8rvsqn7M5MSDZ+AsBVe751dZu1/33qFp3hI3viSMNdH5XjGhAj5Zvcz
CCDU3BWWX03ihgEWMs+S+EKR0NNjH/PRidB6amM/sdK8/3ptxwFHNquRXtA7g6YwSPUVzH6RfPYB
/9V4UDnEi4jKEiOm7XpU77z9iccdJrvyqOGyZ2ZS+bYG1vi3g0s9KIwf5jSC8kXP+UT/220FlJ1f
dZlC4M5//uCo+PO4zksA238x3BRLhwFt65Uxx5xU4764UWTEX7OYqQNQcruzHtU85P1xGYvlizbU
x13MGf+T7ewTWvunhpnC0xKuVeT2yjlCZidu8dKRzIR1LGkqaiA2tiWnL8Hzr2L4nFHRRYdmS4j0
9/NijOoRtGHLeUdMdQOpd6gmCH4vevwhhF9Wr/v76J15tUk1Y+wEKQx8pBoS+VvQzz108XhKzrNj
qJOhPOKGRMZ8QexJ0UoZ4GDVtPimrGSRuHr2Dlk7fdXy+vJSW8iLpEzqoHlVqRUUMfEs7GbT2IlC
Z1pNs4QWzYxuhxf2S0zNlZ7aVosWMfgjPQAtgQW1K1liCnF+VQWGiXJkWcV4FAVi5Xx8anI/eaff
+tRqKU8etlplKTsLwqyy3Qqewe4aZ7lKNcFyjXoN186xZrjuaBFtSaMqdyvLLi72ehg6gx2aFqXg
jjUcbPeMN6nIX7KaSR6W/SipGjUlMt7EDAMiwOMz64DsXHLe3y8hEAjS2bewIt2EeYZdRsyBW3v5
fXgrQIbU1tq3m7KH/aZpnLHelR6dnsyA4sKECVxACSrWbf+zoo2vU0aNgars5X2NIWWDqzm6fGJk
38rDysHkrjnafe5rsSPLNI4KHp+On0GB+lqvJNqCCDnISQBp0XCOtTaFQl6KABUjvs/C/5SpGpFo
IwoMzIzAshPN5cyjtdXnfyMPppjHubDWsLbU5Eqss57OP0MRC8i4amklT6sdI3wxpS1qi1AGKK8A
aoJAOPZS5p/RBTeKbIdGdvxy6Mf6Vo1rxHLt8NfvxBSnHn9aSU3wWAEU22b48l+GdAp0YkqFkN7e
Kb0z6LawzKQd3c9jDJqzW7uCQCDgPEAQv1Tvz8QpiWScaNdnHcm5yaKlGoIJy06ZmicdYbegXTDw
P9oiCcYH5+/xohMWsgXo1vdtC3HuNm+zG7VOoIR+vQcKWT6GWTftQogfAuRuvnwKA2zCXSGufD7m
+U8yRi5oycRDFhZHQbvYfi+elj+++8DmwLOYjPMSXWwrxtgzRO5llFVGWaEtV2tXjRg+3kfZdXr+
HKe91es906epgGKR4gCmhXnNkn6dysY9QNDgbjj/QdVdg2sqUPzX+rYl1jOwna7fUiXc42m2H2RE
tAYYUquSykgzxgUSxnW0mLMgFU+qw1bExRylHyA0RlMDVQchyRgXJARKgf3zulwP0RQ8IxMG7ZPD
dMUO0+SqaK/sAz75/Xqe53rn2EMj7Rj88nPQIKQbofT3UXhKS2NmQbXiM4fP5cYqzTG/unyx2Eze
hYreDsaHWdQvDdO3Yb3xIv5fYDp4poYosuO8OzHO9GMiymakSCZWqhYf1VMz7DF/+gyBPmlakIAj
UL91w5dcqJF0HfEcZyyPc376Pm0rMQzPyjbmKsswCSrVTLVkc9TyqIKTpLa5OBIX5vtgmlwfb9Pg
bfUFCj2fLPuzM/Yqzrm+gvmHM/w99lp2C+7RKNf81o36d5oo3K9vYNhzCfUfG+u4w46fhdNlPnq4
0+eJwz7Z+H31et1LtmD+GBm04NlwH2p0zAHGpKsqeFRwhiBlyTystEIfybLwlHsDgK5/FACYj9Re
oOXztFUwtZJQqqF3aLW8QM8OSTmPK8ktwLm1eaRaJ/olK7DqfSlrX3W8ZPWxVKUlYl4EAPD3/G6U
Z3s4sHYGydKFYtAwwywcf47yLjD0YcO6bSrhnfnCXu3Je6MdrI/H3ObwFoovQIg3hziZDDSETPsp
3Wy1LAGf4U1cskssNHiSvx+MphqHeyX2/LtsPB7h83tVAS9TjCp0oAPLB/vtouL2qDKBQKBygtiC
QqsUKnXehELd9cnui0P1Byk8guIi3RVsM3+n+4Iznkh+pJ5ohmjBSLXhO0G2XoY/w1tp8w2pEfDD
vFk1cVyFUL/FceuorNDDKgUGY/ZUcAyOHEBDPiIZ4FnBI73UpSGpe+8mwC25bWz0wVBFU4DFB9Od
4cMkrvmR165jRY2weOH0l90mnmsltSSM74ux5ULOCPG0GR99t160LbZQBKOTcGaabnv1lkwfvjlC
QLs5B28CK9m9uCRIajfQBsacjEBGbcjvTfLdKzJ7VwOEacQbNIqfjRbbeE8uk3GcO4/dzAX5T7KD
pO/ishoo+Sp7LAMCzftzHwq6HT4Pdd/QDDs5A9FgpOm1rO+Wm9DAaegsHsFJSb5A508cR9PuMNrJ
ZRDai8GyOiJyVSuUat10tfaealqUFDT4k9PHrvjGhUobKzCmgPfTI+gEmd2Zk/yAQ4WKZb1Tn/2Y
nO0YPqToOI6iS9P09fmx/Ydp0ZKV2H7Qdxga6u7UjITc5sH9tSdyXvDul+KyKH8xp078p67S9dRE
pnIv+G0wIQzNnbExCEjBsI078B9xC8RveYJ8VsopizOY/lZHuSsDv9nDdv4p1HtDjaLMD53uEUqS
zUaW7mSEUfMvijxGqxjurW2INKhuBDjFRGLlzEgydmJo1O0/tocTGNssg9z16eP2UGN+yeYaYQA1
gH29MuxnOqiCdeiwCsYY62FXWXS8M09/I51ioNGh4PEPH8qahoGPTrC7o3Eq5iUo8joerDvPeNSh
yaKXziZ7N3V12UteTLMX+Drw+u6MRD1wb3Y8chBZqRvYeJVRa3S7kV/0zPPd4C9uW3J4SS21kEjf
WUODy4WNOWEfptPWH+uuJ2t8Ig+lwPXK0zDr3Htba0PT8TaVmyblcKQuaSc3G544Qfj6tIWF2E6E
8FMZIfxYSe/f9p/YuIDKz/nTLghDVyPYO5TShccf/8IMi+LbrcdP/b1Lib5w7ceF1DUItr12nZyA
DValvCxepPa7HnTFhiKexKg9cHZ44Jxg490JMkIq3yVmwa8Nf6BrdajhQ0+rPW3UyTbiG207vhfG
MTVRhmd/QHtnP/rehQwoFmnJbNvM+v7PBzBo1CSiJlnYwqBJwUNSDxk5ojVxd0kfznnALP6QMYUn
vL4besSHqgwEmtcmtnzMEI/azMzMsAd3SQP8uOoIgHyp4vaHM5NZaVxu9FbED/6ITNUHeig8rN/A
oODJKf9E6L3thn0mrIG/QxV5WK7kpro0f5Nt6rTbIcJilpFGfeACV26/Z9GicI8edaDxegWK7tTK
bbQeATlr64vHNJcxFzRAFegEJ+idk9mgnei8U4QpMk2toh+dmzH8nKhAC7mPlBdJLo0hGP9bSy06
JbjbczWEdN6JL/wwHnkph/RaC7XqQuvBDPn4tUHuYYpG/ku1SzQ0iVnIMNhgIHkzSdS+D8RnMcar
pYhA+5kNwfXwWEBbDrpAdZypsGVY2hr0PucgtFRzhwKl6cXXlvs58sT1g6LedCyzYpuYcoJvZmY8
ISpxPYR8dautTxGG23U3bbxCt96aV3h3j92iPeBBAUc52NuvjYbmqwQfbTcbgh3oJRDhGOe5f24l
s60CsyZvPWQCjIDUJRklN+O8RBfXrxqQdpe1oz61vVUOF4bHq13Dxd/qJ+gS2XOovU71b04fDou4
1DWwRpzu3ZZmylD/6U9+3fc7g+XO8XcszKC8wNgMbiY5QiN2Tp3efrVNNVnZ1AP1YPYN+www+ikR
gIOUlR7DCyu/JKB6AYkxPS76ccjI57ROVQWGIAHyQLQWK/TM8PYEVu5hvUao/slMEmtfQw4qE6ME
eslGRG2si2ewWl2/pfKjijUZTIJnU6IKhbORuYtvHf9GUoSzAl5IrJv7QPMyPpJNYdgl9E5xXUqB
6EraIwyFLEakX5YZkC2FTp/E5JiOjpZ6i28FeGu/6K1kGNVhPRJBdQhKLi0qEkebzWFGaMibAj9b
u5X0SAZ7uUjNv53UtkSR8ZanKnmXQIDZNmLB9OCmvNPuC2tGTnI89qkRbjQrSAdxgzjIWVeOGLE1
r0yGFjqbdV2UgCDlX31kZN4Vz/RaGCeNhc+pYriS/4Ri+W8fJMEosmOOlLHCuVfCZ4fW0tfCU/0e
oYp9CnL0q+COXcQ5S5R7Fip7t5gwAO0jxiylofIneGJtV46LLj88yqB59E/SfCXb1GMbfhpT0UCN
8TwB1SWml7zy1uGGtnk5M4HnkuZfSC1EGHlAv03r7luBNysPWXFy+4ueWFCmXL2BjKoy/MwqH1cP
84v5JF1GsriI+lH16WoSbf0OhSO872cUnEh+rPRVPGngOXWNKVXKbfZRXQeIB0XfC4jAH/tcGnW8
/x1oIHZWhJ02LAmHPd5sg3J9kIZE5A8c4lu8OqaedgeN9HavJ1dz9vhOsVg9KuVzU3LHWKEwNe/l
vS0smHJUVgXIgL0vFth3h2auuX2MgtTGUwakh+jrMmD/a6zQhxXK5PeU98/JJ2TxuuuVL8vXHk5f
NJ01U/MacqLAzE5NzGscJu5n0MtYumX9ATG8b+vXt4gM9LXhl59Jub2Pylpd6VL7/Miuedy1z1Bj
dY4sFsvcnrDE3LTXbdwtl7zgKNet0/SFJpYOrT7QmHZ3/pwexTSDOiG3VIfq92/k8kfLhZW2DB0s
Q7MXNasjIkdW6bFPMOiw86ZSDQwUnkr1K3g5fpW+d3KmwYD0cZCtMFkPIS+dHg3B6LU378+x3Kdc
1RenbSf9LCkn9FlhE68APhuaBGcY6UUge76mSIjZEPcee8xBk33t9lH/UUrMH2f2MzYI+ljptyeE
x1lPLM/oe3hgUw3xC6zxzUauTtN83pGiX/qp1CMF4mMdTCulnzz6F3hxTj2pJKJ1309sD1+fg8fh
wCHNzwl9cwqwcQqxKfU3wh5YxEVWiB6QMSz3nre84cic1ZpDkIbkHAnKS553A95eI/bWq9NVIzwX
Jm0spuzzuY2tT2h3eKcgua0EuvxjvjOEvzMGTtEG6DqUCBxsg+RdW97V9XwPzPWO04mE2m8Synor
6H9/ZWSgdRp7Ee4Mha3JWVdOUlOIYTTKWUIgQzmbi3nMYcN91CgkPIjWyClCxHUc/Bn7KRLMgg7o
Y1PxntqDHnrRZiFrIGsfxZNSbj7uiQXQURh4KMBwtvSc4qFUEJdfxdFIBEvtL3M2xhDA/99OWBe2
aALi7rdsV+VttcKcyRz6BPku74p9JlEM3SQATHh+QyCdDK6oiNqr6SJjyF9k6rlvv+NiNcHQZcyG
hzNjFSdc+qgvoA9B/eAb1imE5BEhD83F/lF5W6X+XWQ64SlW0K4J7V1HYYeCCqpnTMpuEh4ddl26
qwrS1Pb13TVr3pPbY7n+zeS4F/0XmVH5afqc3M6FuizUWsmsYpfzbhm3Zl8c9sj/KruuJNNkGnc/
DU5EpCTxbZ+lYFyU+aVQGbsAxf2qsFPmQLqAoF0SiUBTsCOtVuw7O9fZGfBXK6eXDOT4dlb1F99y
I0OTp/PQMrTDcXppE3R2zUFSMNvXoXzVGHx0TjjsJ02JnlAtkBzIGXlDqHpsJpV/F8C5KcP3curJ
EAX8YDul0U1d3gS6Nda2oLHt7YdBg91ls/wExGL5U/SC92CtkPGKP5gKwotaZ7Gy+0lIdpWGGrfn
+m9DffhUNEXoLwj+sKmo5UIlGfbMF52Uu9GHF0Bkrrlyk8dRdUqWkfbmcravecOdaI/u69AcmlI7
wBrLA8p4eZwWDHUgk96l5ciJCR6xcRwugQjsMzn1SlAa1TnjwLD6PWXR8EhLOgKoEMalRzgWInSO
54ezCU+9ZaIAQUCEJOAyNipAzC+KEv8NQgiSuXOSQmTt8iQh3C2tYKGlaSdLdciF3ZGp4f/1t0tF
MYUuh3q75ciJ2dWc3j6mu2c3Ow2aS5bP8Rc74H+2R6GgF+BnTcyqLwFrakUgLozetDODlIR3SRlD
dbXU8fT8ikIYRudz4AgbLwwvLH+TaNvSU66sDHesOZOTvKresn1x0QHrT6uOaTWw6lzWkzBLLTOL
oVVJQswCd/kB8adF71wfmztGsUD0iLqzGz9rTrAmWjmPlbehxjZty4Kdm5BRlNBLusAuyYDE0Pp0
+XQKRX9menW0ct6BF8egYo81B5teFszqS5igOqzh1zUWE+I3aBKbE3Jy5S+quLbi1PCVEuZqBf5d
FPzrHlfBtKcRl1Zj7dtC4bjmkXIRCfeCPHERDz4sEZVv+8wHyLun9Sy9TtvTQXjXEr3p+qz/xsnw
Daed++4VevwDoQO2zFxNFtIfH9F2vFf7uPlQwNvSeOiAlZ82azuokoIOn6vXwr1MVdS/hgq4bbPo
2ACrauZ5vRTahD7d6Mjyu+loHttr0FHnzr4UPzob9j9nczOIpxy84ssCFuM/GH+sX6af7/YYUJVp
apsoIXRfYGpdy4rCu6xEkMbwFP9guLA8CqYnpD7LonKyexVtQH9AWu07A+p689DGOTWcMvdho90S
oFJOTFxcv8c97OBRRtMprk8biYtA5MzUxyhy+j4dmDoBMJlT02q4wUsFZFe4vyKIN9qsz3xEDsSP
NbHvpsca5yNPDALn4FdXOIGtCMGj8lpGqI3Q26sz0UoLSPXoy97ojGDBNb1WfmJmepNq7r/o3lIP
/m7GIIo+/eyrt609u8XCew00GQY/yb66T6Yx8X6xeLawmrxlxLOEx8WjXeV8fHM9QXyLIKxXDK9z
rOEXMSzoWlFxho1Wt/otw8WkFOWXHKE3MF222HO6KIeitzJV4rS9Fvz0E6nsKLhlvOwX3PEvJTwU
jBinsxs3ZUofvfAUo/ugYI/pr917KghLbKxLeHhtSGOwh+6TztYmynNlX6ASmsot9Y/kZyLFyVA6
IP3AHJisCcrVqWOoysuq/DcLASTEaindaKX7jHAbj1KDKINWL5vWpXoc/ViBlX/iJVArE2gE/iXs
eCf0fTtRZtbBJSMbTWn9zhKJWgj8F6tnzk76p6aD+WcSGh3MqkESmev5mXz+AjC9EgyJ1AQO+sJh
3T8RvJcGKugC448B42SoxUhoFylx6hTeMo+oWhq30lkTspDtx6kqQ8/Hlil0mvPNu1OmhBLU+AfM
SRM1/VS/+Rd/xRoKuK1Ueq6EMZFT1v0HAH8W6OLG6h4YanftyLQKIyemD48qqI1ZYi+c1T4FOBN6
Ui4CPk3ryvcWMeb6UIXfZtYNKfYVoH2pA0+sDsEOU0AWHumUgmvoov9hEKcrRvO2yYeLYXv0gHw6
rf9IBiHQPmb8vvEp6ErtGmfEFow0ozPqpK1tSpBTMMZaEmDrYDgivUHocXk6ebe7W9DImmXAd7a3
Qh07YbHxJm39zPVDfc/fGzDkoWC+LR6VGJyYLuG3c3B52lCKqfLFMjPSqauImdlg7b7WU7qsMnVf
QLV7H8o8cD8aNl2xa0LGKDeYN1DH+2xl/t4rzou+zYlPrHLrp5lg6egpqnxp7hY7CXl/9VtHZ8rI
RmLqZd8qLV94RJF24hNT4F9ALNqXBLpzzFeN7Sxt32Qnn9ecJS9hiXaiLUV45jXa4V4Ti6tnSi9j
6L2+BHienJ35FikzsUlj3PCSCLNATT6SCvRJwky60ugVaOQJNRogViSvX8vz47wIFmDgis8g/A2p
4GsbOd9H5Fb3XXKd86Gqu4X+qe1ys7nPRq+N7HnDa1IrejGdHF7x13NRXrKUOHfJGeXGQdJV1kes
CDvW2aPXDaMETkWmPlJgbZemWobnELYKT9tAT24KZfzmY6p3JPhjN4A9PAVIUQ+Ml1UlC4I1xHfN
7nKS5UkrTcmSn+DK1Q3nQYREhv2jJ5MczYYfLlR6Vna5sGC7dR0G0D9Ub7YO88rDSwR8s4JpKyFb
xa/+9kIRYp1SjTHH/RPe6t52FabYciosH7N735kiMjSeRIzRTEyXLznr/grJ6cUhUFvLKx2V6vNz
jrl1YaPtwFxIX5crEGjKQfSTFeBAtgpPL7VdSqEWwN6OmHiQIzdfYgouHRrMyYmzCCSHynKdC9aN
88aCspAhYBCcYfuRpSeNudAte9Jt7+zUsz7GnZ+S6NAT6jxbHOXCPxOKM8byXVpnJ5vGDzeSNNUB
asNx3Vixiw9KOB/l7OaFiY2vBu8PQZsZmlv4r3T6lvoixhBRgnp6hVM9SLzLK6ML0nzVOcpPNtXo
xPtP/eNYD7kdf4+YRK0SmwEwAkobBl51cIpk/pWzT0E0ZfrmcVPvZ3+woU37UqO+mt7UL5ldu/K9
b4UXAVoSKh4+AfNmSbE9n3AkzgT7ZaZQmzYZeVIm7+eMT0jxT2FUYptLz3VsgQ3PhmqnJmRD7dMp
abDllpJ9gVU9DHYDxjpjdW/Qbb2b/ainksIDc/OOpjXefGrRF27kG5R93tYAxxUFUga2uDye7aCE
zrnuPUuboowcTm3fZaWDhaAYW0QiIXa+lNlcrCodCJoW8BgkCl7YNdFLpIXz+ixjHWElbU0wlxj/
IgcvSH421NfrlO9kyhOjl0RgLilpwqN+TR0oRqHs8JgrVvkLEfIujCV1KAxn2f1Vhyz3fq+fN2Bm
LSD8nWF8JNmWqcRK0S7VoMFEZES2pUEE6y6t2CakzBFrjRZ/vXWqxSgY3tVb6TZlrlHSWKjKbHqD
SQjSJH0Em3uCqY4llxlMXU2WEjRgSOIMocDHkNML1Mu/qxLRG4UtcVHibDes8mIH/cYuSPThaJlW
9W+4LFARkBPhPTlPf+AwwFo/9I+/TOMHYqGN86NTDs6teCDYl+pGqAdTKCbaWkMfCVFYO1V/L3Vg
BTlVPQtzlx8vqrZwlKtWHvaULwXU9GaFi9KxiHLvRxqRHkzPdd1zVRfcd6zX0j+lennB0fDrGSV8
DKfIV+qB8V2/1BkDnN3jEueQoPBLHioQMut20NB63+E0rMEOBgcRrYX4IZ2O1vTaRltyq/7cEfCS
CwhxKis0KUqTy3F9Jm/cwjsvJE5o2hnSXToODlLzj8L6cI6kaU3Ub7OFYCUAsflTtNqJ87ocXgPA
FC4eLw3Pq7YW9lx5SK5v7aY0h5mqltLkgcc6N7ZmsTcBsnKbFoyG+FAgof9OuZIP/jh/DU93oNED
DOi3kDIgf1m8TpBynD7zvXA3CtKzoFEZDq96CunZ+vegvEjF9BeyCDxFFbyWu+iaQP0gYLOchwVS
6xztxJ1NbC0hF/GZcPnMdj/sWXN90JhOpo0cUUp+xhTl8Sw7ufx0tm2XtXxzjDoiYvjqU+hI5Oo9
QpWsLSTY2+VTDV+VL4fgmTK/2TfCbllzk2+rSHmgW+9xhaa1j4KVBvg1sThZjmFLAAV3V4z+sKQ5
QJOSkLuxmwnnIch64XWuMkKci8WMub3HQtfj2OPdQTnOhcsaBNw5IYlLq8W6aTFMA1990TvSgCTA
PlKqqqnjd7KpZcHauN4gPMPguAipqWZ02vqAUi/IddqApOvf31GBhn/MDgcTZrDcfk5Hlu7AU5Af
z6tJXEXAKnlJAP+jwt0S5/l04FpRJKc4YNxFiUetbOzU6VYgJlwxO+r+L1hyN6j25euJt0K5x82w
ugETBNjpTZs7bAyi7LmUaeVUbzRDELT628zdV8+B4YEPwv3y0HKFGRHlhZbQFZRs6drliOVUwrtA
ZKAgUtcdg3FqnZC0ET2eEW/X4I9z+REv+aLwsf/tFTC+3qaa0bkB9wAdS3vQSX2QaBrBqaupJh10
l36DGg774RBjcOfXsPFriVzBA9rX1wBHw9crO7R5Rx1FqB1DERgPZkRjye65oM1WmDrDEhyooCx5
k2IptKZrmBfE8tui9VwwI6XUMGi42L2KiIpBYUG0nVeURM/cmBP0wswxckMWCQEPrZCtRxxM9IwU
LG73WbGh2wYzBO6H0AYxWujsYdemtkvOweaCHmLsVU6djHVrETY3CmL5XDPPHk8CH9n34YHE13kt
Lrhzqvih6Cst5ibuKDlg4iaSjAVqpVNlhG5jziN39KWdaCnlM6UOx63smOk0vTIfyJWUbJVwXE8k
b8sTWp6unP9m+88FaMPoSjjFBPjWIClHZm+daXgEemkjccQFTwK4oaVqgaIpGhbZLLMU6cuCbqN0
/kBgFVzyahIxKtd7myzplojUBvgYELQJGKrwl56FZn/SfZVfMs/sM7SVPPHH0wn5gz2Dc0V5EAUp
p8P8+oQuE4ECk7Mm30WAM0gBcXoVd5H9ZMcZ4ll1n3XwUV1ZIzR9uZ1cmKxIZPSkk8y+5/FKGhjy
BNVlRP5PWKlunw/qxq8pbElXoVqilEFkZ5hZxehhS+dL9aM+OilDMnA+2vPPEZyTN1H4/1yLxRKR
JWw+izif95CQhGPqnIKGR1IDub/7kiPYXkzV8sVRHv/fOdV1aJimt3LhzPN0FOXtVE/iZL8HU1WZ
B78G9klUwCt+05wvFz1PVzOkMz2JO9+SPhOrAJ0P0EggeQH9QBUlhp4z2t4piMO5YqkW/4/KAKwc
oYj5ob7c1aUqKUvxc5dF2Uu+ZHOhobXmSetlfKike+DBsInX3RUlbosS8lhAzXyWPlTiNvAFPKK8
C6B2hTOK8SqJHKHF4ArxBwi4rPX2kOFSTAg2yUaEAhbSoG0Tm8bCs8SiwWA3c8Vj9KZ8WzBV4vv7
Wkbj8x5HZZV1z9a+v0wJSguPMbAFodq5alSxQLK5SCmmWXuKcmpVTS2GR6t7Sf6MfvRtJ3fosEWu
kPjozUQm3o1YI2v/OqKwJmGiBvzVg2gEkTcL/nv0aa/vDTwBnB6uhkmya7n2l+YXWB+xvogUgi7B
v2R/35NS1Rud2ipLVYXS6KlIhIpUM78U8P+n7dsBbAqEN347DMXFvNrlstE0yGv0NxzWAXddC/df
3whLz7i8701mnDXOW3V5GCfJvDNXPlu0vc1GEYQailU1v6BxCWg98YlpNiljpstpFiXaroF0N3mD
3eFr5BOJtQ9Ub+q4Iyl6rgniKCP+lAyG7AVCOH6Lw843bkSuvzrwIkNGMasZRQaPtfXLb9r6KD0J
PrtjH95p3lcTk/ymBxTm6txzlCEOPddRwnFeAWL4nLNVYm9Lj9ABEYidFZMLLLobnae0DMeIB9UG
lUfX2a8Gv2kGw6qnUCaSlMgnpFygxgOPcwcrmx+3bHiciSwZA7eAv5EQRyIFSPLKzDG8gQbkqWUE
onkx5OaqkiFEuvOAw8HyagjU/T5cCYHYuA8i++5XjA3CVNG+J78OLH0qNMrkRH0XKrZCkb9R7alA
GyTl/dcxq7uRzLpo3CWPNepYTE635YPQJUUTlt4KpL65MeCgQj3zeOumXde4RHYfTdi54cZ4vwYu
yFryksY3iVIjR++MDhyGW/8O/f4Rx31PufKU4HO4aMl5Www4rSAZRZqysOChlXtj7InRwJ6TWoSr
zQ0vN9qAe1rxz1UHykMHrwJPDSOoWP5w2bxaqBfEt/JoKjuWGSW1ObdNTvUn5keJl9iZ8ZD2JomY
ErMcbLZTAeNF9jcyPxc+0lrgipUSxzGy9D9Xi41dsbhKhm2Uz5OFvODQ+GnQlvtCrXxoiV1k6yWL
l0SWyWb9P9orM0WyyAADGbWSZajKLgDxwssF7mb5hw9JB6oXDhbhXbFPqk7txb0CS7N74Z3obYRb
tbWqG2wT/SM5h6Jo7qiCDvxIWznYmG7iCgrDmSkaC/lnyr9fqWnnclE3V3SeZs1/3GnAPrzTau5n
6OF0QTu6WwujLwDPzM9IpZajd0kq57Xk8eFQ6GFGGPQa2Tp9DR7rLeIPb6YbIKLk/uvE1L17+rww
ovOoSETIO9yVgyd1sbRzpkSnB/r8UrNDfUpdrWgzVelq6P1cUBPi5V/IBlo/GZa+7nStfFAJkU4D
Ja6kV430LJIM9EEC/KMJmNQ+y8qfSGfA2XSye3tCwYzuBsEMu6eMhLPoop25AjX8BLJ5AFw4uMc8
c/U6xu8WnyYxwb/gFOWLcHd2ih37gE3/2ByIg9ZXCMcR8d4yty1bfKGlXQgu8kvPrGQ9NBd+dyZb
VAfhSVIrM3tesGXp06A/ucmcQBWVO3UiiiKbBAMFHLbfDpD/P5km/Yb4EhQ3AzJQ+13yS57g+1IV
h5/YHUKVmH030jGpwfrwqiWqOVqjdTNeabzN/xCiQ88eljiKXuMtH1sl0RDBWxOwgaagiEW2I96W
/Qzk+nISUhDSqD+lA9BDfX86oCNDetyEd9ywnjIsoeupwRmYgIy5nfhIU1RCi6x4+uIeJWC5Ys2P
SOnxt1o0rrlgcYjyRw0bNRtUEx92rUW/flOWMLj/676kq2kOJLefIkehfmZLmPfqis19vdaaPPua
Pcm5vm1q4NLonxxg/GBdDTdQbJ2ZP8fED4w4Bt6AhvWagMJQg0nAGpknJgIxvj3/hJsieB/UcV7p
+Wos8LSjB6mU6AXWJoQLC2txzFMeoJf4PsTBV2qUqhDsGe9SHZMlAlWtYeAdiAeULxhUfkmCOvTK
k/IAvPLrePviTOgEkR4gBUMnq4scZ6VMAGad0A7moAaiwg4uMi3YnZLDdrdCX7R0+38V4yXilzin
zyps04HSAAfGLVRaflu5+ixNaI4Rz+QxaFm3ZiLL2iDGRODUUKzGg6zQdHqq517n0sD4k184gzn+
Q69KYDs0K4OXnlV0kvihQoH0aYTE4lrpBkXCQaWsnZ3MHvHTmv3D0qVITzxAZw2zJGkopButtHN2
tp333uMNmQtlHCTlSMX9sse/QO9ZpOflT7H1vMBc9qJgdq3ZPeu+j0J3VdqgHNiOxMvZWYllxSKN
aPtgvAeF83nAqDmuiulCXUp8LyY6ki+uBPkYiVQGhJMwYsEg9Rlb8dVVooQPyZX8B04GTD57Rj44
Et6Svo2gywtTsSHMu1MTxkra1gL9Ll565+CtvMFVTD7tIE1E7RHkSxz41cAznckZfeDq/STKj8w3
aOVIjJM7tHXQkXL6iEBJyIqX3rx2DdQSGMSXBnUlbi9FyzyonUcHOdc4KTC+iXELlHkLlKagVdPN
yWrhJWAlczR3tEwqpwkGskwLq4OgpQ+FwaLPXQjnq2upv5qO6H7NkK72uLKjDKeoYeHQZZQB9OmD
JImoafEO9lFhVtiUgm1pb9zzzMQWbGWazO2R/kDG+8HwrVQ6GEuJXhHf1llciwQ4wxVxGXC55Ouc
8LJnwq8jTc71JbeFVGvBr14MAoNZFjfKunlwGmHdVPS90mv03rReESCEoEnRI5H51NCqBtIsqnFX
ERWcVMt9fhE71dLywfX1KqVEm0YbUJsfA+iCAs+IGz0oMRj6JDsVbLZ5S2+RTsdDXoXYlDNvj4mQ
lMCWzgY1A9uyipMhNX3UoiTDaB09Wt/j5n2df43VjyzF7vbtG0kVZXMDvj2pnYmSU6asapS4dJp3
ZY46ug1ET4prS/fFWMuiFyJJ4u/F49URMXXg1z6BqrUIFLu4AOC7qv1EAdcSBl7EZgHCOL83Q6J2
I0TipbBQ+Oa8KhSCwnWFUpPj5SsZ33427FsoL11uSzR39kxj2H7/BUHspQ10zrYrdaUC13RzYhqw
5R6cqkuHAidFCbMVl727UoGOXfjNJ0KqpDN4nFipUm+eKLKBE0Q4/xTGnQnd9xfl2tURetO2b9Tj
n2bJAAH/7SZxktPNClzXLnktgWZ72bWljR9hZOzgyRX7eY+HboLoT/GU+APemiZg2/cZuKrZ++Is
nEz6InMkHi+tHWgjcOQo3hBDWDDl5bRlK8Vglj41+wNNLV9xEBD9lr26UOi02TM9Aqp+5DjIJd1U
atA5a6oF0nC4HF8Nb0qwIDsgQrkChkY4JyKeYshSph4Q6bgPPS252oA4Hhl9XjyW7f+fG8yEfKg6
0SAE5nYP6NTCL+CIThAsdS4urTvX+PQyF07EwKNOsJ8DRaGupwLqR4Xm92eIt9VnYGeEqdDllLAU
8JOqjlxG2Zd7guiYnMirhpw2E5baBeQCCTesn0bQ5HHOFAtgrIluz2UiaWg0vTzlGeXt6Qm2yiZK
SKdX4n1/R9wLQwIWxrtjB866+9wg0xv16ucDM9jKwDGQbh+mswRBx6+hpBfl/LiGvSTZnnOyqeXA
AqYtqfEXliWzUmlRLNN5AuoGypyiIgMaXFKx1vp+/c/cB0eJuOgPU5o6IfUKevnMKBREFIKZkwDj
t44M2/XJdkN3PF4MVZ5RYE6sWslTjFgXs5quGAUAn4+8fXW9Xh0VRZVQSKb94f7zXf0/HGweEa+q
a3gRNPoKGd1wtUagCOa9chUYdr9g0ri/L1bak7h//uWYgsDNUdyt7ajgReUuHqTG9zqua/jav1Kg
1IDgUtMf77NOSjkuW/WpHrCA/KqTqZv7NMyMGKlwPLcyfQegZRAv6eTKbX+XSEvqmKfcK/IXlMze
u0K3szf/CVeAS/d081HI15fpE1OJ0to1dEGZevwHtloFzMBIanNVXVinRHfTQiPw+q7zTXgnnmrI
Z87rQz5JyE7v8Xylk+r63S0bCkps5zqayv2js1gCGFOeU9ikNCDY3sP6LV3B+HEo4wbxrtMdHF4K
1K/RenzLMId/3okJqfJwUDtIxAaGLzgurCPDw4GNqcD1LqaBR3q2ofSFyIvvNFmPrDxuUedi8mNk
cuzT8+l1a5kegTHPHmmoIRh5ZsLjxugyVqhO9VNjSS0Ulb7ZqZY9uIEE7oTIBmNwH3GjUHslQIUJ
Kci69X8wGxJO9fJnTGxpAVAdVQmELovS6ZD5HK1n7mpX+Z5Nl9TwLgxlKey6iRR9t2MTWihIj01p
0fHxsXW/nBnMOag4DBz3L/K9yu1TSgnwqsKUp7KOsZqzgsj9rS5n5SK8zhFRrnaURoqX+jomaKzo
hd8dynGZENtdz/GkF/Zz98QA42Ed8YQf4NG/SisnzDj7GpOxj2bBvYFVImFVF7UltQW7qFTaQRUX
PpAOcTusPzT97xCKR2CbP+3WHbVj+BtBgYbvJxAytUz9Yfz5xB26QcyJUgn0ua9eqlZu3Ygj8r+h
+og5/txTBdGontk3qaMB17FN0s/5uwwxrRN6PWummRiSVguhFkBekFF0YU9cmKDQMbcJsnCO/lqM
H+yskjEmufv8smu7nqeQ6wMmGnRybOoLWkwuxvP8/sFLX7bBUWYkVGl71ROVgEdYDWFW44rGdtbg
9lCyPtW3va5KMXSXEh8Uq0SDdvVCQ8qrpP0beoR1LhDl5vY9dbrhZyUGE2JlfG6bT4KKp42OKnrq
9KgzZdhKzi5sltjk2NmDlXqB9VbJDqyDvNm5q5RxsWjqZO1dgoQDFDSg9+2Dx1ao3FZPdA7M46Zp
oNK3p9GNT6Acv5a3ZJs5dosSQUzHsydlB5H2cdIBY3v71uWfcx3KrW5wp78f/g97ADpPBTSyW6A9
wLG2fIjnAHGpq6EGAnI7a+1gx1M5ESK0Nk9wOFAzxD06aDhrOepsgc0B/7Uk4wp7MTMzPL8DH/Hh
VY24/7/RmwQW8E5GIuSeHmXFx8PvDQ4wiqFUTtbRtP8ZohS6Q2qftbEZIY3qjt1yj0+6aw0I6KWb
25K0boUcGISoBVsBvIux2meyua3E6MCo4pqXhoGnAQKcxq/+EBFqUo6mYI8RG/3daeAX5Ku80LLx
qEEPYkSmLPfXxLIPMH0x+Kd/vnqRYnZ7gEo/pCc0BmzY16t0cpuNEVjNR6t4ACUTq3DItU9GFlMP
bdY5/blyvqxBl2vLW2jZvNG71DTq7jBDhNq1fZhcABb3L5Gw+m9+b5y7LzQcomrZctZjukgsZ4IL
+3mO5Q34wagjtCff+mk0XZqm6ridM6KcU3TAoLGGRxLPjh8UWkU+54yZ3WRgqbhXmpZ+3NBD6afG
J0WI4EtoTrbi0Ll/9uLROdyTnuUT1U0Sxp/WBgnOENfqI1n0bp8Ag0znof+A89+p0YD8IBFfJPFd
lQ1CWy/P8O3zKb+T0KtlwtXJk2lWOV5JEG+7HcRQdlcE3SvdJPshR5sEYSC5l6/LNk3dKvYvgXoY
2YKpp5OG8S1sB7WIXUgrMr+yLfCli21y0biUXL1u6h35gwcEpRzsTlqV3iImPm0swtdHV3E0BQ1Z
KO1q0FtUV8gA88Ae4XsUf8PvyPVtdMdLCJIqeDKaqIAW7tk/o+U7V1ttEk701esD/LpJLxUT0VxB
MoB6kizE1SmJ6m7e7zhEYzLwwMkqiJCrb2ffcs+LgOMyWkcIYMHuimhq1ZBi/rArvSeBx9YxYBdo
rKo0a362z1V2dSufZWqX+Ev7pO6xWNRz76yuHB0ZyAqDIsE3+WjhZtxyKUxRc0wmiR3sdeKoHNrg
S9rUWrNMG6VUol0am99JJMslUy8CP96LcyF2M7o5YlsJwRt6afq7O9svDge7G9hjAiMGo932SVqz
sYbzDeqaEjHGKYKDkgMISlVAKUSRM/J3S8NWAa7woEgokH6jGOezPVTXhT3sQDJoP4Hl5qlF1SQ6
5geQGbVtY7C3uP+kL7bLOZCpqq7tONDAwtydln89N1WI5qm2DHUiLA+CRTzxfM6KLAHxGOYSi8io
R3eRvkBxyMxYOOTk8efUOUyRGoHRu8qbuB/elCYr9806YfBiCTff+cczyfTGzUIVjbGL0AOIPg1C
cXDZq4i+urYbfYAN1lab4kErNu4uwrodDy73Xps6IOCyIMRPqBhpGuOux3dxQKH926c0yc7s45S7
7oIYdJKr2u29cbRenzHPAlaOFrT6dfrF7M2XOLzSRWIQROOpAMqJdKWytZ6XmFqSLGkQ7xgKj7mV
SDVxHPs/U/5oBeccOU27bqWKy/wXXDxxdfL7E9pTEQ1FOsWS112tFNbd5/imrf/SGMKkf674rc1x
qDPcz5MDDUKZoK10Ah1gUyeTnKIlWpkwkNaVNy1JXXCdFVKE7LbNTDBcT0oFPVFcLjrfRQkDSeeR
Csae2ErWTIP4ykRoPyBfZYNiIDd/GS1FfNNem/hktLO6Qr2Sjq69w1SuTFRtkpKHj68lva9bdrU+
HZJ/wxAxHV66sLmlT5Wk1NaapJgWxnzgM84G/XDQf1dWjpWH5zHHL5+2rX56Z30Dng+VkP1bV7Ls
glWOnqa/28GrifDgMM9S4wtIeVypBR+c4ZA2vaWOqW2wDlSMkwSuJa/BwK0zEYTvHzVXw33pGvg2
+Z40LHqjPd8JtUyAeHLM2kaNLiRiXrh7BwOuPQSH4hoO4W5qa74h2RhrcnS+r5z5/pKFX0JVNE42
CKD3go2R3Yc+5nwxTA0vm9zxBnFNim2ChuLLZ7Br7cJX0iOe0mEBAJEsaWRsAxfBjvagGNOfMapT
bYlOyL5kKjbJ+IdmbecNu/QpQOx6xPiQ7fYUktOaZg9s4NQ7oCjtvihGxakZBDbNdP4C1YtHH8EG
uGW6u6wRX5RDgcAzisQeZWrR75pg6xtiEHs1XPvcn3j65Fe0LhS79/RqdxJD2AtbhDEyen6EDZmO
odJi2gS0Zsg1E9WeIR2wfkWqRREA9zcbVs39hPZ7BB2+N0/JOr9RYHA9XXQT1R3Mwg3SIA1Ej8Ul
lxZY+nDXWPA8pvmI5KywLxZn6M7TmrlEVJPrQf97LlOJmvdu+woCVPMvORFdsf8Xy3EiNs70uQRz
0kYBMjm35E+Mur9sy3RpdqKJVmMqlR1dQT6armmmF04HwoSvHWYssA2qTZ6sBXFPquKj2rHnuv0G
YnUv/jQw+auFeAvpC09O5SlcRCPQWKUH6zEgGOFkm7AoijyWwMx4+7p9FnJGbN/9l6nGNr5eQ3y1
xF5XIhY772z9kPsH17zm15JU9a6KdzhI9VkrpMIkE7a4Ko1IeU3kvz4DnWPCd+NWwUwAn5f//zcL
OicM9AjeMHt5e4NCL9t0ROfMMhg7pOSLfC1Kj6njrt9DyossnHB2O7u4F1rSJPUkPYxqElqIY1zX
+RNlTmQ2Eb2FCqVCx+MHOK8M5TuqWzoOTUgGaDhf5t3oRqAIc5QwLG+RhoBolqOlxZaNtQJS7KqD
JJRs39CLszluC0qSY5pZ5H2QoOVxXSJcHs1zKo13ppAz5rzy0S/gyvl/Uqqi3BhElNHqA3INjS8R
p9+C3bICEQrGhK51uHo28LQD23pBpPm+LQPUyHQol/E/REU076Yr356e+FMPCSx2o+RYm/h6UbzO
TuUIy07Vhkrla9XHRM3jBVK+OwsvMg5HtDFVseZt93xwhB2QTvZ8cgCjg3/mdKT5ktueqLf2a7rm
kpJ0Oys4GKkOxKg4WcKuWlYTCaptFmOLfyFXvulIiZoJh15fE8mufQd9dqCL9E0WrvRXF+8QImaP
RICr+D12ae3oHc0U+WV4RIGDyXTISHCc2/gT37PYIb48mymw61XpM/za2B8tLWO2tXWaXas+BWxV
wel47oqL6Oa+M7O4JsLzGiZ/y49JWkhjGMeFtKdcLX51JM/GMTbJbxVl8HB2Uso6AnwxV0d9R5WA
3rCuv8OoagVIODU3iU+1h6wAXETi+MqWWnh64gkTkK3iTHCfn8Ha5b5TiS0ieo1NXI8s6gI7Rmjo
JgxqROYsLB6KgWSzJKVF99jbiWQcWtP68K+8SxemCX0oKbaof7SI9/fV3HU0HwjkJOpLmtOKuIsf
fth3ybUCcsHU0CcwvkrvaKixMQgd2AYSUaiv07EhF/LUXd9+AD7z46+0QtL76xq3f3cxEd79PFP/
3GUe8tq2O+Ej7YveQvKW58P7HiucUtbNLs7rj2XK4l7AfknV/nPVOXlpgw1xbSMBQulMrrmix2Vq
AQOiepucQoe+9nfZyPQeQQ3cYgQL/I1Omg15/ZHZKQH2vvY33/IOfdoZXTrzRg7VpY9v0Q1XX3M6
kiiVN6/Dyd3DufKFTuNC8eKgwC6LVDKP7W7JPKTLv/no/okMblGqeTEj2rJW9n651bxPh/UioPxv
ZA22fGuHd6SEHO00UDzeUBFTwk/q3A5JjQuFkSXxewMw8kDKIKPiy3JPmuh4Y1nl+3/ixQqY43Pt
3D8WjFSJ808LXH1bagKhv7sAAHRcecw+feKjy7FzvQGih54RS+3iz4uw8QoiM/XyqO/TsTap3POj
G+XTSiBsxy1xAeQE/2yuaJ98ewM0LOv/mEO0frguCpFQFNfuqShsZ0QSL6F7ppvS327nh3tfGkMA
3sUpteuGuS6JLUzNiiJaOYgIIspb+AQgrzTI4ibvhI3w2Akola9HYBrNJ/p1ytg2sqsb6lT4hcHh
/0nomZgMYys/l4r+RuQ72K/eZDadLneIJ/AvNFoGvU8R2WhsNH459oXviH5v8wPunPqrNZLOYPwl
fslKbbq2wurFL6VN+ev8xlizgxBjyyDTLSOl6cQV0HODceRDE3xzz5QVhhsTxcYx7JWg7hT3VIfF
1zWRFkhY8O/Ogg7z7kDoAvit9ywUeWhPjYKLNs8BYrUfJQfIE+Hi4476qzDKIO/C/p/53rLMvpW9
XjBASbS+L2HitcbQWGqQsUof2aMj1gXivymh4RsHxO6BJam93ftgiZUeNxcKQSy1CoOw2yMcYqSQ
ByiBwDZ/FvqIfzaZCNL6MIPvCqngmceBgEPcVHeqaJcifaFGsyG/skm6Hmv8nrS2g7pkBeflWoDZ
ZxoXkDBTughqi+ttd0mKICAXxRLlolUBbyIEsNz5PYk2R+bomqB1qQ28abUv0v1PWOuLSAt73ysk
RY6FQUkllAXWj4PKlLIV0BTwBaQslSqbSZHidxIu+kqS1YzgM6QP9dakEpMo0gWbWHT0MsZDR0Em
wYw3hBXw7cVcNSSwir8Xb6aKbdtPxWIoOEUQboUBifPn4mq7vtvx8fh6YkpKisWdk5D0+nHQcnP1
W+sE4cnPktmTEYP2C783JFKhcM862V/m4m/TBbk4S7jIBq3dml6JPy0Gi9uim5qa2EKQ51NSPTad
08mK6pvBQwg+QVKXApkukJhfIh5LYB1TIXZ2upqb/xjr6NL/cG2KRhHJUZApgE1Qf3Ee+JJjo/7n
BaJBMXrbdo/Z+HK4YLGflsrkgz/3Nyr8ntBaku8wr4bll/rozbOhWrhyOaMvdq/fH6Ib0veRRJck
mLsl1Hf/6Gq/v1/fMqxxvBlHEU1PbbXWmzJRw7Yw4YD0W5okZ0TW/FNmXqhWAsql2VifvaY2N7uM
b1FfHLxrxfp9CQeJQu4u2zJSE0+qqPFMq8iPtoRwBs9nWp5isRmjJwQpVBTwLej7/D3vMsTJiR3Y
7OIXIkX9q8YqpYqYnLgiETW1fIi5YphRqnm2Zst6ITHbuoHnf3yXXB+XGYynOdUCvkQjWNnHWIpA
riETP2S4DgcxPRexjNb24SWxI6M9n619wsaxmnq6xIN3s4HLcfozcK3SnSrzzlNh8HAzYOotyUX/
y6TpElyAubGYVetKjihE0qUz9jQpPTbfC3drKNZoM+YNNqHY55PAejAjSBuV8eIueJOVrtP6Vrbp
vlnWknL8wdsiss7kU2/FEKqh8xp1b/xZtOa2HpQcoQMecOaOx1E0U6f+9gfau2CpZMA9MfoLQIb3
H8Rd8CsOHcMKZ5QXHkTSV5QgyALFYxBdBfbQsc7fbUb1KUnJpnxOG8D95luD28N9xD7dcUkKObEq
eRoY70NzDYaYD2Cgpa1fWxHOomj8CxC0GBtzVSwVOIQfBeEDDdhCQPiAmctWFboxykuPvjQ0ruyE
eXwnD1X6/xlr00znu71kONntLqcDTKkUcxWgWBirGo8KhNRbHYebS+snuXqd0vLy8qlp6m3JMBB6
MSxEWCrZOIUbREI6YJiHWiE7nQUdcDl3TqGfLU1qv/0018UND/2qR7OpUAqHVzyQ//GKvQqhBcWy
xg20b6BQAs9ZB/VSIbuoPsr6mDMg+GdEd+NCW42wt1/UiKnppABzOlCIvZ1tNV6BDmk9gDtBXQSL
H9yJ5p9WSMoBxmy+ViUs6conW1/1f+XWmpdE9Erdi0/61K5d2ul4ikxuIfnQMnj/j6Fs1q+s55uP
C/SVbOc5T1sD3YuKvxhcqyAqcYHCwHT+znJBu+ZR1semSkbopavjwcGBAfGv2XGmh5W86NbLiFuJ
C7yVLLtjIFSnP8ZZ7WhON0UAqipTWuZb9lzwo+J/2PYMXLEVgN4ctz5ecxjO3tY/UlwUD9DFyUxN
YPnKBibsVsOap6CEnKhIbtGAns4gbHUBQp/U5W6c6MufSH/IPeNaxalhrWwmsQywqYPCFuHM2ogh
OWBbLue52zloPUQHyfoBKHOnGesaS5VrGcyuYdYc/oRc2MsxmLFbSfCP8cf/SHeApsglknSETTJB
iBn2z5Dj+DMNEWkHV3TLL+kqiSHtTs61jclHUoqAgslFLne/1r4HhBT7OgNIp+n1ywZWFDxpaMgQ
B8RYVP9lBt0HsuUbZDJW5E1oZl0gQYN3yYEV9YU0cCnYQD8GDX7YM6ekwxAuzQNxGvfiNDyQq+9v
/rZuVbYT6nfSwwLrSejtQNKXrKkh7oryk7IeDXWTV84jY7rig7unBtMJ0jhMJpzrNa/M0HAegkT8
nTZIvg6Jo1XqKxJJETySgMN6xx6kkty78fB5rsPsGUM5bVAG0ysuTbiKaEOvu5u9WmDncdnETW58
Ngh6BusojJ48J+R9sg7Dsaecet9M17UevUetUTWHlTX9cMo57TdIf6HkZskHs8qdtDdmGcG0SjdD
LHExAm1HwroZpWKcpYAgelgWHMQqJbjCy8fErGbzOVt78pCarYCKM/UEnoEMCES23AXKClmYOdqp
BKxWJwwtygxhI8L0262VFWGCKrginnmjSNBJxlwcob5EKueM+TWzrG+EjbcQe/yPBB/RsyUl9ssi
WFVKCaAUichmivI2OWVQ77enr1z6qUmJA0ngOK5ljWxhaurgOW4Ua4nx9B/MBHuD3+WW+1FIdwET
jn2c4/E5YI4O28bX70+ssvY/fXWe8q/3HdpKvFjZbcDxUhX4Zpm3tGqiHYBJ2A0Qe68ExiEtZnCR
OC1eMlqoY4FtxmPhHXa05gBCJcVhFFHkv0NMh6ZBgPA8jDJmI8+5eSZxfXkRiAEvq+enMU/uSxd8
cKLyVE6eF3WnPpB4SiiA5UIbEhHyBK69uODB1Mg6PCtmSPzuXsgW75qAToXhuw7z9KeAde1NQ6iy
q991hpCgDuwXyTv3XYlp3ps8n41qLFqJHa1C+3ZxjnU5g/D0jEa1a1EWhF3AngV5lclOhpJ7Db2u
Eo3mXo17CzsORJvF+60KdF/kp2r2ybruTWJ8+oTESo20og1tRZPiJKsR6ReBuh/K5fH2+9iDSMkF
pDJm2G2+UW/g4cpjcVo3yMpbdiefh0oWsktHA9r2amZVPDNh19Ea+tJY51HyWmu6bLdF5QyvoDCr
vanw/c+XpZuhzaxyokDIDHWW80/xpsw0qIZte49CXEKWRpQCQtwbJZ/+MRPN6fx7mfv54D5rydRw
K3msJJ00FZlnYugDisubxoFakmaMHLO76D3NXJ16aK40P9KTvmY7LV7oXWwB3bwfT/lAoElrqgvP
55tWq2DQ1RaZgiUsN5mqnfasivEFZYXZUQTAhPF2zmDcpFcxe8ik8QI5Q1X/1+V9091zHOeaH6Ux
BEnvXTGYg6/eadmYNIrIMjEJkf7auucsJzvcyrVdSJ4pbo+QHOi9XHUJll3icbT9+oFa7XtuFDxT
VxoK+PWeLkuLt5DFtIDGXEoMTaO7JIKjAzzp38+jaeIoYmMpQ0VUutFGKnPksv+Sa2tpwbGcROCr
Pa/AXGQC6Fe0dHT9+oVAm2g/TODGGUHDf0Rb1oSBy2HP1G/EEZ4m8Tr3+WG0vpqqXHk8UAqFAI3r
qoJnYl/7fblYxMTQzGBrNsintryfrVeDOk1NXuqh7T2SgIKHhPIrjdOdvRLtOMgD2Ka/KWKs7dYw
PePyD2zlJN7jS4XrTxu8+fM23PmsPfWbl8MaDT/YJ0D3dKpkXy7ZobeHSOsbR8uFAOlE1TPaZzvo
ZaiZgOzN2/vnox7kp//MO4R26EGWj24dwUQm+l6dU8p8ppYqIsYWtpY6z3w3Fn8TCpjt0BqektAS
Zs/saxZwXD7QzYO0DmYIet4dWlG9/X+hWfjx0lbUROcZSO17Dtxtw6QblPh7Ns4i6j75/6tWqiQY
NN2WKt8HQGvAg5W0bL/E6iYR5yPvlib2A+bjEgpNlLin2K4fc6q1bWvZDR7I2KI0rs85C3GnXbQT
4fWC0N0ZibdK7xveDynahLmKOPgKtxN3UZA5LxQh7fLK2TrR9hQ2aHoqykkDz/uZv7CgPGCMTvsv
lerpH8IcjX6utpKdgBV1B6guN4zJ82B530Qu2YOYSypzU2YbwQl4mwjjFyG/4YRl+tnYEjdJs/Dy
LwvyeV0n4DUaorQBha87NwG3y2dyqw3eUvpwGvnouuRQ0DD/Lvj3J7kmMiPUIFy9cq7jp8v3sw4/
QWlvX0oX3NmUIhlheLsEqCNEw4nh128Y9PtaDgmHE906+FKuSWl++dVpEqEaC/WzbAaTj1sbJT3G
j1NvOltau/kf1ivNpNc4bmP1RnNy1KPQsYOuWV6idryQiUj91g3n7mE5F9+AZ5yn54DbEczEHa1h
/SikaGl4hjIJXSDOVWvkoR+pj4cnHwuTXqTYeXFEPW9W9u+CBQMTenXjW5IWmqgzX+NCQTRhsvyG
J6tMIEjtK54PdhbBsv0zzgC1RSMSBR0aURWU8U5ZB2nWlF9drT97iL1Q170/9e1kpowERl8H7mKo
rsI9FnTWr2CFuMC8YxXHpeJQ83waoJ19XsYN4cFjRZjEYfmDkt7fClylVihqnmk5kYzD31GMN3ab
1jz8oXKyl2GRs1E1hZ3cJdUFf/8kb0O+LlUsk0KhIW+maOa+kY8wFc7fZIJXJvBJcr2ym+IyVNVU
5P2w7Kxc4JafchDCgjAUaniIE6n9yYY/PyM2XAgQPt5ZuotkbPFpgriQnMNSZl7Pc9aiP4lDcgF1
gKHYQv324cWaqY9AtayeqTZhNHhp4K7EY4MeLiCh07EJ98hq0MrjY4OJkp0jPOlYk5nEUFBXpduR
P/YU/S5MIhWLftPs5gSXEaU28d5yvT+YKSPaBQooukj0srmMZOqNVx968okxN55UP4uDKYQ2AGBk
654kpk/wcwNN3ZWOInBw115l++nLiZLIPrtYAhkt9TlKtDQdCQhSe+9GgNNEF9Sud4f9HLVBvzMP
yskpIZHe+OkilEXWDdI/nUfXhRlJ6ARRoaB+bdqJLtGiDgitFsZTonNNew+dKuzoJgMnnv8EMAvQ
iar1h4+R+ma9Xlodgj2y4i3k3+y8OEt4bb7U1D5E1qYzWaFB6Nqw5BNEp8CUKHMCluKkfmcfp+1s
+T/s2s40rPNmtkbltqQ0LQHl6MvfXkQLIbnTuv59JYibVV1wV8WgUz9MTEMmXsN14GhLYaL3wwIr
mSFNiXJnPnE/eXUsILOa9VTab31hLdX8JkmQunlCv+zwxnHBImow7GAVsfpPu66ihW+mJO4POxli
VH1j2C6WtdtY8fxmc5/foa83hDyczBmT65Iimkv+JSBksTXmwr16fGbWww1vYG9wkQYqNqTdY6Wk
cNks1wAfODHzdb8pjDaen2Ql19xnWVi1tqlr50NhpD/ufzGMBGXvU5wiON5JnElJ2PnEM0D1mESS
Fe2XpyBTE2EXWxT5laV0nRLfjgeIZyVRzSnja+D0wlcoxfEIuZRe+T8gqpjfqXX660tRlpbfrvIk
JLu5koGCBQfdEwu7TQrsQ5PChvgijit20exNzbXZIHdAvFWOY8F1X/cg/g367acXsKWoMvyvPfGJ
tpaVW/NiR4eSTA+W2gJnqqfnBrmYrDQRlQ87OZQLd9VZEGN+Nld0H4EUIXjivcM/WvW7GqJk0gvD
BPiyTYlFhtRN+RlAT+lkhO3lfqoZatTFQq6Arz4NvG2Q8XgH5YfD3yL/kbTaVbPOyTFe6KLWD7ga
nZNfZXhnme2YRS7QQnOzlRJNqKfM1d5XHSXLIqtRsUU4BRtswNpsnndS+UxN/Bgyqrs3XqUM/g+5
IYdYKsDGjh0z3c16uD5JOUXLV+kiCFFhgmgX2S+PwVq/qy/1mmTxVNII4DX2uHZWXxTppqzq4aoo
N9mo1lp5U/AHwrz9luC4p8YsSHY4on/vMltiLsQzpCeqB6BRT5GQQ8G1kOLq5u6VfTYTdanI02j3
az5und8HW+12o1C4+wAa6rdIc4kORRR7M6O6ffNvCVqmtH+fcR+cxw+pdR5Fan5USUPKuSpLeWJL
xX/bMOrkRoZdvMbhDx2tqpA1yCN6HqSH8jQC6uadJl/CZPMGZ0tNNlb4ffQldRoFHHFXWvDWbKfT
M4MnY1g8tVXuBE8v6VWwJ5SxuBfoUeQB2BW+OHY5jCqYngsELhGcKoSj9SZrnbbhgUYCzBJOFNjl
cYJ826AUbuAkMQ+y/r3yRz2ctnAJrkV5CTnQIhzxNTQMDrzK1TEPE65PbVlZ4MHwpnBkQh+rx388
PytnO5f9vVgnSJZ7Xpwe9gRILa379WpJSeP8ekFMQ6fTvgJuW5xMqfqvsD/fbHW2ilgFdSak4EwH
2NsIvG27Zsf9YXlSTQRhFQgHSkstNVPp7qLFS/B8Vop/wmzpGjELzqoAjov3wtWgF50XnrlLrevW
iI9zQ4PRhXXELT+qJ5+xnGXIsVAPZAtN/1TEv9Ny9/PwGEW52ozk3M6DjBSifFsdUFlbFui6LgYR
QIrNbxDCT0WEQwKZiJWIRAfCuyM2JacL8EQEe+NRpQSiv3u9aR8P+osvOUEv648m6LyhYGOPfsI/
eMc8g3yWF8r8u5cYcvqyEsQM/Lv/hkUa+ZpHm0g1oZC6WQjGSlAUrYFoRksKMDmbzGO4p1/VHp3I
ukAhVy1uUChvA4WNgzHKSYZ2eqjnbR2Zq6dUrknsN52CqZkJE16/g31kJgwTNPRcss4SuF5DQvLv
43t7P9xKjTFjH1bNTMmPJSLj6zDrnMOeNvFGIdLBMxopJg5xUiXUTeSM2l3NDOFUQ9+sycTo6/bw
+CK1PY1NW30NP2bGqcgHJi/tS05QojllCySpxwcTNC4Azh8/yUtVkm4clRQy/p1RwBK1/46V4maJ
HMyo2KQSXd1i7kL1St9X8KzNZ6SRjilHBiePxzIVlhsSEcnmOHIer1/B+ZkXPSt45zi3dYD3aici
ISlaajdDlzdTX5XO2hBa+0CVvSuuzDkOZRxwhboNpm2kKvXoGE3PgclrkZv43l8ZZ4qKhn+7n4Gm
DWyPAYIFKxVz5XgFvj0PSXVG7t7jiPRY1j0PLmmf43t/6G+Jicfe9rdgwt6WCBezMWy94E9Kxyyx
BubdzsgM1R2nTlLwdOx0dT9u/5FA4dXVyzKgSer7/NTc1eZhcIuLGDYkb1WQWwBoY1ia9KaSSp07
8raXAaB+zwJ81W3CgPwIVnX/hlBCHRcXLFO9CBGUsmxmS8s7uNsPwZAT2pTKqCb2glSUZ29ZqscZ
khl9uo/kb1I4x3oXjESNr+urkx4XMU7Sy91+3ohQg3a7SK3JLRjv8BSpvQ/vxIhuH5L0ewUOHPLY
e/4d/HAdyGrBvr9OniVS19YGvzJOjtCzrnfyMOZnhUHsp6/8sg5vwsBIBnXQHYMH5fw+vGEM25JI
vCRXhd5ggYS2WycPbEq/H5/Vhu4yISjwzzwk4Zsrj6b3qGBXiRn+erJeRs0OBUjnZnFIpEaB+1gx
59UFOhe5YTIMfHZ48WU7cA+/z+6IrLJch7yxvwW9M8f86q0XMYXeHVGu6Oa3TCpGCxR4avAW4O4U
3KZZnId0werFA6/jdscdx2R+H3XuP5Gk+WEaLMDlK4CJjLsiL1qIj7y6dfGaZ8Hr1Tkn7x96tfZq
PeqfLhSgwv5ukDbGDhHwvJusgyvMts2jqlXRmSIz/dzAJR6mwFJMu1r4DQcS2Ew1QPy/gLJVNNS5
ZsipovbauoHGf8T6f7jmyrNkBsoR/+SKn8mOsqgndtvDp3qBLoeACTSBPiU/3WUb5oa1ggWP65GN
8N/xIeMCNk8dn4apVReU6KL7DFq2alM+qKTa1tw8Kfs2mqAtAeUMC9XsAaaJTo6LmXmjutX2HLO5
l4YR4y72ckcahPG4VSYLdNuWS/cl/FP4J+HJfUTRZxqttXUQjIcmxV+ufpSPXTYIjxvWeBOFV+m3
g0ptJzcEXGpbr6Naj06WdKsh4X8L5WdKKNexAsnoM7tgmz99gaEZrU6ACPP28P6/c/5GQysldWg4
GwZGnvKpT31cUIjmVuUCARnaew1ArdvOIaVUejdQJXPiYqvMaUAXRhldR7I/oBm149L0Ocr30n7S
f5lMctAHM9SWpQjfFoDaUluhJ8J9P0hF+GXpLk0nT4Vk9T8ZWJSC4P1/PvfG89shAgKfw8dSwjnW
XfvAVdYokH6mW97KlweplBBuMIRFKiSzZ6eMsNT1laW13aCF/zwO1E/h0Nn8WO2oJ7aOSjMFYkL9
bdcKBp3Tjeo+aBQsOe4wxbuW32nEZdGh1UYbrG02ecCkvI9nJk4pC5gg3MMcG3IipVxnbYFelEew
01HdmElUNg7AHKBsNoff/zx1PkyoIvEYP03Q92qvB5BYMw60inAroHLzYzEWtZOeVm8YQuLfhGUC
hzXDATPQXzPz9QNJJAhAXYm19Oh8qzYWfe/vomTx2jiOrfshsrEvRwsj4wzk20kqbWl69afR7M7M
CY0iUuEM3K5/dMnJc1Bh0KTxGX2/qu4V3q2XaFRfbpSrFBLPr0l5ANLj6GcDioG+tHzTQPTyHXuV
ZgxZ253dv5Bnmm0QQkLPFCn2XmqfZPprmdBSU/DvL9svoO2UXzGAEslo586tEeNh3owm37h8XART
YKrs2X5jVxMP15MnhIjN3jPGYk41UFZZu2CL+urN0Apgzzch0j+QnaSf9XIrTc93DdTMAVEzC6CO
k1iA6tdB0z/ypLnmRnEEDB20jf3uklKDxFgu7/VuewUlo7Dor63p2BfdLD4xUSUuVSYabcAUMmrJ
MMiJS5XGr13JtEeGGkM82eRSNLfGco04hA2XQHNa1bPU6SHRdiFypnl8LA1ja5TQFGipMwyrK/s9
GALi4Z5j1hq5+k9ms01Ax/w9cxqe4pJZDx6PJ7USiaJ3MX0dAYBwkDj4MZ4eBMMzFYKfAVpySX5L
xYO4lhylAtQsm4d/CzwqjuOk2iIBTg01hieaBkG2Ffq7ezBEIdL/8jZOJVMTRLEbTFoLC+4Jzpcc
YZg7rpKxJtS5vrsWkmtN6+R+CVfrSLOK2akPCk+PZ4Zt73ZYAmX7qHmw2oCNSvcqq0xv1NwYG5NB
J38q0B7zpmaWIaU+b4XYbDADKf0xuiMIDLheVtyRiskeIjnxV7yS9A+pi4pzDmJn+2PwWLKQiVN7
HjfUR/kdOX+XPO5DfIVg476MPCMgRCq+q3+0irqbMqc9Q56WNHhizUOGtaLapKnKibPfT7ocACAp
6NwUaZGF6loAMYCDbnQ9Yn3gjwHZrUtJJUVTV9WFAPYGrRVGE3BjYt6gZE0Hhmpg0yQSRNPfWFiS
PtpsYbzC3n4PkwrGnGU+q55Ce1NwCH3NbjXfawGxPAabmxuKwJ3VaN0TBPIOmj+oeLJzg/J8zfhC
Dt3s+8J9F1lxzqtH2nhYyYbW89oFr3kuBLDHUq0BEk9X3VT7hE3Ui1e5M9lRCfLptZSPEasGt55c
u80TdwNVo3jKkuEx60cu1eDHHewZkRB8rpR2PhwVUjbphYzjOSfCDZUjgwKr03Wq0LK/Dd4k4B0D
xhz0vijHpogPY1xsf1QJBMIG4ABuQmcAkndRXitRJkQwzzOJG6lRq1zfNzW0nsgMis+NQtuV2knM
4IdtKGNrALhmBMU/S99sCfyb9lBCvuw5omX8+aVDsiP8IXYPVXKTrH7jC78uaqn4dmv5Q2cfMCmu
YzGaoBvmFnBGR6WZ7MdJn1cPVT5lr3yefvtbKOVqsnv0PDSY641SNCfSFDdnjWZd2Ub3mVMQT37I
e4eIMorhpGsgY1qVhdFIA+7PlCL429vtqV0vw25lN27CgqazqmDvJC7ChByJ9s8jvw+ueL9udlo3
wr1fWStK9TlOs/tepSZmftEv99DL/AvVrzJ8modiaEUdBkYm7m390TmyL2iAncSRlEyeviUN9SEh
NrQ4OTE9Bs1y3teeHKphranAOt5j/eMz60kg1s9dYp9ReeVfxleM3UlBz6T227L8XWHemwhLW+5o
NrpP4nBi0whHSG7vRmzZqTeb4fd+nJm0W8kbsji7/5MQ63yO7if2YoDBJ3Q0SO3zeJYcxf238pDG
eWVf0zLVZmit1i3pCcnH3GRfhjIg4UkPEMw1A+ZpyCu1A8t6T6k+5Xeow5SXYQpatptJAz9fu655
/XBFBzTkGsE477CZzli3WSpRxMtjnwZlOTZ6c2vVBqhbLXxIftgA/2pmmTIX3W1usXKvfjMxIdCB
tsOYwh1BrynW/gKX5ratXHgts5qXyZHndzVtm0YM8HQY/6OU5whwXJLldGtqV0ENdfyxQhypBowt
X+Mlx8ekF7t1F+sFRhLl1ZlFNhltasKkoxZgoBGJfQJ9GaIBixpC/BOY5mc6SWSU13rhTOn7E/aE
tSZkseoIFGxInYDvyoiYvJ/aKoGFvW7gNHFRaRwnEhIREWEcHFY/+iDtYex0FdzBUKGK6PpZkqVO
+uLjCMH5J8suiR+awGUm4tj5JVfSOcodzxFjnIzIkEeTEjTbBQwYm20rvaSqjSagvgd9lDEleHF3
ZaW7UeucVvbIG5LtMuWDwOnizE1EQWzWFMFzEVElMlEBnMkEHy4FoWKjS/pFXPmJ2pOEeT3SIrd1
A8qFIXok3Kf/y3INkhWytUPBPCukb0S3f3LD95oq3Gp+6/fYz9Zm1wLmkoLJzcgBZ2RTJBT613QU
xhWZvYz11WOELAp2/R3lnFpQS02DJELeoNZH4qBS235+c/XwRg2V8vw3BAcu2IKRbxReGyK5pggH
KJapWNEa0qH5nsP8YwkvzCZzvBGh8tgDPucbsFb9Zv35ey16qRbCSyWPnfAm+douqB3xlI5QROAt
3aOKpdubQLVauCgtsfDhdAZg97n7wrabEtDxPmioUmcJ63e955cGgTrSzI9oGyb8rjViZbzT9Zs+
dSrOsMS03vRzWqQwLNP2mazPaCKoYgRmUWBlifO8Mmuz/Cf2oasMPLyOjtvuGJ17gQpq5wEWpB4k
eOve7MMiuQHpmNJy+O6E4tPl8IVAI3VZk2wB1tRTfccRlIHQ9dHySt6w4Dw3fKrQFHqQPE1Vi6ZK
t2FRwEQqH3Ltn6DeRhWNqpOfL5HSjYz7tnf8XlX2qIGF2RTMdB6T7bqtkGz03lRze1dDriE/4zVm
5XqolLvIuNpXUgBAYN7ASfCK7Mgoa0xCv8E58M8mIr5N9lT5aROd5dbvS2jdU3kolz8M8OPNM65s
w//EZQro1FxrVYYdW1SRTGrdrjmDT6FlcZObzHHl/yNtCALy4i0g6yTWW1/zuLS4Nfyk0/nDmyft
E8TLW7nsk3KS2iHZsqW0isAMFUI/jq7XA/9qrwwf3owMjBIIMI60c7DukGBzDUP+k6uY6ZE5jgK2
kJIvT92rMdYm5zRm5la5S5L3ZYxT/szL+67Lq1UaLjVDUU9vAhDpGySg0PyqjHy5gZ5r19RqaN8m
0DCXCddUQzjxu9x8QtAUVkApxjyAxA9O47exOehcQSo6hKlrv18/N/ggtwpLSkg4ssYxaBPkbR6/
CuqyMoK5W2KklcVtgMY8FJC3MXZlJWje808KhBJ7Cm78gG13vB1+hdNtgWNeTusHgv1UJzr5lzCw
1XNkvBUrH8LBftA055/f9CfWKdW7mtGocM+JydDSXy1iHPFMm2k7JvS8mR+XE75It+970lHPa9Sk
3rldilD3+85zHZ6zHsVdjFWDfJwGzdSn1XlgiDlUPIyA0N59v9/eYOzIAfEmW7BZwWhtMacoi/vX
m1agJG7FxALF0SX+t140nK8g03dJgrDorBRWB0KrCu05TXJk729jxEM8NmeFek1J5mRqoNKl2GWB
brq+ErrWyjv6BUTZWqej/nkeqVg3kHlJXvdNJ5pe2CnSrURehpztZLYS6IRyLld3OgTe54wj15Go
cdWNsct++CI32FA75VCLg+BJD0fIKmbVzyrlynC9LBzbXlVdQr+DC0zSNsELf9JkOkUHavxNwXYq
DlVrZ9x2VUT9uMpi8FPSy1XtN3ymlmvPzkANeKinxl+6IPTUi6c0ywScukwQBoHaoCzLxw/VVcWh
kqF52B47MI0ifkR5FeoLUaPlcPUIm79BSeA/C78DhI+d0w1/ko0rJ215NFd1M2vqMWWqa8Xfe1f5
38WhAelsIXjGEQnNWO2g9eWqDSAvqyMSjO47yMrRXjipneG6wprwzYtO4iYLAcXxk6Wf2S9fxnuz
FMqTuWabU4PzewbHQ94joWyXYjLqvvZBFyc9YNnXbsJSCckqtupOlwo7iipK+chZi3CH6Bdo/CFd
TCEZk0jrwzoQ++9IZR3x17xODuY9Qp8hpBXNfEma+uMUELnv2+GAPK4Z1mFeA9Q2EhOHNoJ94s4d
juIS3tGG5d+3yH5ewtXnEKi5mFKt7RgEbsB9RW01nE1Uls/PbmZVVoiRGvULGAjk1fPpKlzbipJt
xg2RX9howkeS4s4J/n3ujGu66JTAuI2KOOEbaj9CdK0T4tr4PlbrLmwsg+K/thA8vJcu1SJG7JVD
PrrpG1+G4obKkd5LpPifcUJZIyczmKeqCW40aAxEIo/6XB9QNpEyu3m7TAVUBBnB4G1gpC9Kvwau
jeHH7AQ43meAPxQN+B0cJtaIYMA71wYGWnarjxLNyg5WJDIVJOEXcrpColc7sFIMqkfza8PrrXEJ
T8UconYoSY6p/kuCG/g16rQPIi2zZoeForgWSRXO10cOvlsyU+YrnSxJdxLgrlf3GRkfmGf32NsJ
lWUMLcd21GdtnCrdPrhIdV7M3PLRB/QLpac/vijWGsTAVTqyRPi0veYPrnLqHNiogFpbuF3v5Yk3
yQpnibVTB/2qbAa/pdEQOUw3wFR8mk2uYDutUOnJkRRkE1Aa8I7Mh/82AvnsL1StIIDeFU/CxRSO
jPUV8fpR1QRqKxrqWzArvN62yCWbwOQwHmGgJSBIa/W0OVJsr8VUmoAmVklWaErRhxMv7mmtmhKm
aDov02dfUnFUqoc4TlBGyz+6dPNU5mneEOZHK5UQ4KQzQe1oon16YHoQn/Fd6JKRfNuYIc2gOQVi
zqHr/E7dzy78K93EyzMJmfgul4sL93JiBtCDh9vnVFhg19CU0nBz3setUgAUcXsBjoGWjBPDh2WG
AUZUxPhETDQmdqCa85HA5MxZ2yvZIkDpvMW9Si470BwbtFw+fwS9nuCbteaDC4QSqVq1Jg/Nngss
nnwnzRpHGovAQvOvPmhRTpg4LpslR+HuuSL7OpAEqaprjELfZGN7bHlAYy/9sCsSTw5kEREtHWHf
m401YbLlz14M61jbKEgEErWGLsCrOEcuyZuo/89+oY0YnVhTagdFAf4S51SqB3b4dQOPZ6KGawnA
iP8zvqzab1C9xlUbUVljuGj6/iNfNsoIoOGM2HXja1WLbyNW3RG8jCRrNtarT78+ykuZhuCSEEjr
0UtWhJTO4pnrEvhaZgnZm8hzYUbFiWGr3BlSWxK4wCg7uhv++5/W4IHaow6E8C7Ape46gG3oxoR5
Zr9k0nOFHQOsqruaSxAByVx7LkL6z9Kajo8XmfQZ6om384q7rb0V+aeX5wD0U4iuZjmtK5IZmKri
p6VQugYnUONtJP1+5HZ3QEPU3Phz6y74KfVridsf72DFyH+HLYbdWy6XZTO1EAVHkYR7Kx9XRZu2
kJsnaROnBGWdWNHyCY4171vYdUFQwy2V/FUgvlLr9d9aMLpSq4Ae2tyAojIdK5aPajsYzLO6SQKt
aDvG3jnVvgoIaUoaM2m8JTR2b8d7vJIBiySznhauIt/S+xzbFqC85qnVY7mprWrfGum8cojg51dU
KpDIIsIC6ec49UMdFpY3wPhFuvlO+YTwFb6J6minA2fvdhnhFBiZsdnUiTk3mhZ7w8n/g59aLgwy
AhIdj2UT3ecGi8WlblKE1NIMbtJFxMaGhARoj3THkWeGYABsHW8tbYRgk+v2qCtZKwkDpQGn4/gV
fBiY6xyNPTruKmMMQ6EnMm1lyICc5rGL3floVH8sAkU0ygD+U1At25rI4QuWTuUmQ7WPj2jhDoGA
xKuq2Q/20sXUnyAwOZLREOXOj2CuIpUCADvexxSWK6XsGSSjxahvfMd9FksE16xJRk7VXAgZmuI1
kH3Qc9B6ZoaeC/LlzMaH0pvvE/CRv04Opk652kymGkXBQxhdC+3GI0OKrmdEwXEl9URAcuHbNmJc
BS2/sxWX6PL+1aAZWy+74pGq5x4t/xEokIqzDdM/uv5JWvwc4b0FRowGwG+n5NPAsh4qMQonf6xV
kq2njGzJGK7QxM+pim+7ShLwk0pfpFyuDtzsuM8QiCNVIIk+4+UzO45ZQd+yYzG+IoqiFPoo6RmE
IlmpPDGgu2luV24s8/4LKWDX8w+brJDgrbhwsHk+IZeD4TedV1NbM3BSNPUUVkjyZgQn4Y/un0T6
sdzk9l2/JgQkflRDuAI4h0a4JPG1ODTLvU4egQh5TdebuCT0xmKSn1ZwRr9RwMl1vuxU1y9M4oR4
LPfpSICK617SZf0/Ri9hPdHyCzwo1Rf9w0p+5bHCnKKK+RQr5IJKnW4weY7Sbd6+7Fv5A+DAw2ZA
924wNnpHihYL7rJo4uLo+DiQam5Alpam3vhWHU6QLVn5jJjZZgfMbDvMMXmmvk5d2Kf976vNuaM9
cl0Y/Y7NiwAnH8DuXgrOxltoipoXqhctkOu74ngwBXbtL2dZQhct7LZJErBd8E3td3KzrmO4yUjI
NCv5d6TEq8WIx7P7+rs+BHyWbwSX4cGQykPWNHwGqxZQ6xgeKdmkUXjyKEDRdIpNI7L//wUEb3Vj
+XVU68E6Akz85Fr2ADSR4TpDDFFtyKBBYBjqHL41W+omg0zykVKsY9czJBuJigI0nzHcBRUtyXI6
KSo6rDC5xTHy2+IlYFay/02p03EqgSsPLr7CfsqfKIKwgnqeecQ6wmlWEeqYvsR1Id8dHQdxLuPC
GegSqXSvUINpSEjX9I8LzSqETsEKuQX67HxjFj37jb+ONjvjLAubhVov+fMJr+rDBhmn0n0PGr2h
h0E0YnPnIr+4dAhldK/uX/UkDIAx/iGE79aWQNqhjdIpICfiz3Hueku6HFSkmAU7oHRz/RuYxgqv
g/1FqzGoNCVa2+wJODN7ItLHugTdLx6B2a9e/5nruuWJcRRTVtaXYSpmmTS5Su874629gXMdHRS9
aFTLby9PwZk88HhrOc9rBI9L6eCy3CqHKqcPjvwWl2MSo8+3k5ZeQH7X9q4vMMFR3qqsXFcxBFT+
MW6yFX2UuLeTHhS1kBNxlAX17MgczkRh3cOEHqoEvu9QcJ5+MmrFaF5BQqi1hzzHfRvrKjo4anMz
RUm8CDVke9jYbDuTuKeG0gbsPM+R/LpzwZEqY5pVGkZR3xc+7CvX0F73HD0T32ePW6/k3912O5x5
vMazEZP2n1NO9QIPrbHNd20QNE0GSZT21NhRU0B3GB3yRVR9WG0NtraEX/eKBZUUyLbS07Cui9uw
i0xLcwqPrM1XGGvt4M5hFHFOOBc+qxerQm8/XyiKi5jRYicP67NA7H7pi9MlfTdgaeOWIxO/V+Wz
SN6RYEg0gERbpEVmUtmq3tLRr0ELo4lawBEC0542bPCihC6O2vW575J9dBWuf51mIEFpKuhAbKS5
jU+1SkTKYUpNtiBeY4EuL4VI5VMkn043T6fYDlE93u4O+QY+y59cWPXfx5sA60AkjWBvrFeW2X7T
4G4jyTshK1gUz5auvQ5JnvRzvjrr5xa1R/ORsYI3oLeulxjXfWSdmc5+3o5FA7Dc/5ULIn2c9Js9
Yusa2vDjBuraQZr0nMjfpJ31VLFgQ2B1KhKx/8MOvcTxHB2DtmtJ1iPCnnqzJPDGfQipmFWLUs8V
kE1uDSMIASs4nsN+6KXBlSqQRcme+gv7WxnXNI+KBSUVXGZLFq7fxU8NkEJeUIYDDcERRrZGGvj/
UQ5NHmocOvHrvbJKiA6YLcREoA0e+9o1R71BMitzAqwWELIWQEHPeiyPEUs40OE2gmTHhxvlTjkT
qEv48NIbyjWKWb/uqkIxJD5Et2qQJpy+zopxcHTjfbjfrF3wLChwq1SuYklg2qRySoELAfSw4nlT
hnV2kaV4bSOMnBh/CKfZJDSL06nnv8O7egNn/3FvuOI4H0j0DZhK08cf4djVIq6t0/3uB1bl0L41
iHGLueEzRw/n2pkjH9V0Ec/EXqvtVTrBQ7T5k36xLZPv1iqBQyzNakV2EigR2LF/Nk+qx/lBvZz6
OJ6Ew6kmlj4AMPnboyC2JUyg8Fj2suO4iaBjlay0KnNutDUsrTPmjyvL7qRxfX1jgF4cdiUS0bc1
zjlE7yWK9M7ef3Lc3g27mVD0fdnIIqgS+J+i9MHNYOPJ3tl7HbDTqNHWUx1ISV1KC+s1qFJSe2Bl
9wZov9IZl3kw5yCBRvMU6zaCPwRcO+ddpLc+Y3MpjlHhDrS6Zv5ufbVaDWZHJ+iyh/kBLZ9+Kun4
HBYXn9K+pAi7o/+/htYYjjGFpPvIdjxOEO8/FOrEAk8f0in71n2lStwT4ERjdIWTOOcb8rLHUa2B
AJ2My8YGbMzy7eatiq2ksiptlpBeV407snEfoic0Yn1akdd8y/W0DyiXHinvGM7KaRw0f2wJ3+30
G36/yGq9ldhjGH5n5hAI3T79T5RF+ICbv3v7HzoDTpKPpwMFr7ckct6+g30YH3L2aAUsUJG9eAyE
6cFlO7V36cc2PtozTtKtFZdhq0g6KfoRTVKZnr2Q9fsXU6u0K9BiDwL5xq/Kn3J7Ais1bXTrdxJB
0ITS/PbVeGeZKNg+y5dN6W6pTpnBXDhV/L7IzF/jCSr0lAYPgGO1TlVaKHFikR8h3jNosNJ2yLA/
07am48R5lNsZHLkMdoQ5ZDRwnJJAFOJI3w+xDTrkveYt5lDZgYK5tF5mhIF0QBaZRItQ8Mw9rI5a
8JqkGUAUvn1Slt2eQCPjqXU3uOkt0ANNZtfOhwfErdBx/mMvRzdUj3tbsmxoPcPBlT9AGzHe9T2g
GWIEjcLi/5Kbb8itaXxjxrlo4SNIDN7hpZwDF6IpkD82aQbMzlM6EPCk7cqiCiF4hTddQKmH7zH8
pMqVXsoG35bnzyPz4WMpteRR7Vod1BRr+9crRTTYN2P3s3Hsp+hkwH9RaFPswmiPvS60zFugHjuG
VbJKjq44XFWZf/LyjeNK/C/FgrU68UMi0LOg9rkjOecETfs2dCXmbI60cWUig45YZ/Q/rOCM6nCU
AS9ethjehB1yGsq2P9by/D1D0iownYSfyQgBalB7I4IJ8rEwAaRGUMQUaENaEN4NNUokK9sxra7+
psqm2lP9o7Rmv+S4JH1y6UXfI+vFr9VenDwKaPnLDooONRQn5p+KKOEm0e99XM/B+kkbJkek3RFN
yyopt8LRaxTerl+alr1fo/+MwFyBti3LBs+ICVfF4JUhaQ1WsmUCT2P5D379yWoOww1sTaeffHyf
y2ZQKwspZd9aO9r8WOngMvFjIp59ihBYv0H7t5a2PufAU6pD/hQXlx9QrXNxkvpAGg9Zs9HhcY86
QcHaTddOag3/zxAfGFAjNhScm5VVWiFFiIBg98c8PoWIY3X0QIMbF7/1gAi++njSW5pIQjTv0zS1
hiXG0MSTOWeRS8ZcB8lWVDIvES669NcnMEd9Wa0GBPc1HWeUf2LI2pBPCHvTZJB/WtROWyQpZqHW
PQtPwDvLbiEYA0Eh04cp0RyttlLXMa+HSz08V+e9aSh1/FM6nao0IRaFpREKNcXEUDcws63LtgmY
Y2UphBQMOVdG0JtyYWVhHax7fmibXDaCWJP2HwmHUnp2NrGefyu6gmQSwZX+c8N6HR2H174PneBr
4vH1eqRZblSRYlHUt9LDYEuIXhzM5sgwA7xa/KFMGqVXcqaT9/Fiqje3nVnyg5YFQIeWkmhBcXct
xsVb5Go2zKS0p73XYGrBAinxIKQRv0u2V1g8ig1nX1/5TpxkLoM3qBzQkSxqjBLeI7hgKT2NB+GR
zEOESLsx3MnwLYa9z0wh+t+eduvydiICTNm/kTnyoAAJQeX+VQwNcktZJuVHJE1/chfgmEnTXgxo
PLIWnKLHWiq5Jz295NBSAOl0AFnD81p/QWQpwFO5PdTNoJ84uXnvHgO+FlMxyX9J4fv3NTIbWvgu
A1hjY5lIepJuNOp9LHeIfIbehqDci1JZX1+SKZgcL9EqM16KUz7XOGr7WSkkarSgaIT0pi8m6kxH
VrO6EudeQED/k4Li0nQpzxxMVvjF/5Vn20gYxWdgVj468rBzNtZAeK1IyPDwqB/iawFG74jA55L7
8/RK+ebhYGMA0Q34MS2AFyIS1t1n7lPR4koZYQEBZiouf8fNo3elmpxbFFWMP/5aWtsR3kooM29k
CORKdUakjjoPX3Hwn1u2HTKLCCFeTPiC7HCFYOe+FRKcOaHRr6kJOLKehExGNjjJjLyarG3YcpxE
cpde+4/I8VU3UjubfIKcDjPhjQNCZzGpQkS+1zuqujufk81cAmZYcrFJ+YTQTDxUYFzDldEoXqxi
TQsmNPmgMgs+j8mE5st7fnKciUMCmX1E2AY5zYNbTtOb7kvw6uh7osc5NhegtLh/Z3BJKOHbat6F
waEq1z68DBinJbCxrACxhvWIEolAS2f5LEsZ0kSdTmSkAsENHL4h9+M19VppMUGAeAFUClikkUpl
jtfS9WOh9N8huRfqI+v3EEIjHBptlsRulHf1Jv5RbEbSNJnrI+PbsQz/K5v4HS1O/Ps+73PIPBSc
AaVrDqD/2QHt4UOqehDfaZHT88LSlQ02MiyiA6dDiTbCs38y2zt3asbEVu13bEFjryYmVyj6es5e
xbr4YbYfpmYkvptWbgozlK7kOolYUvst9wJ3tclsHFKXguBBywKItP0KPn2Y4TCqzYznpiRPrSCk
yu8URK3OGPhz2AalAJs3+IwqHz0HpYfYVd007RxXcLp9ejjopssF/LagrdUR229XBuXUvJwtT3+u
NIivx1xAENkCCjO8L6by7Lfn0YwZyvUtHqgIPYSkBP8uSdiVuPBu+tKGds4CefUbdOvgBkm155C6
jJBEQv1PeXSy+qwjUsoaVoYOfHHxUbKOOw1RG+raFZxAtu/JuIup5YjVyNW8LcTXR0JP+qsKtzHv
d+SR9qipVqowAVJxYM7A1F04DoukLPfjkHkwg+aoM/ruhZZ7i5DDbMr1N8yX6CXjzB6lMmqJpYSD
K/l7kjtliCRFyTjDwmn5UH1hP3/6UCiz5H35Mv337c9QMO790SJJG7qbR5qwbkW3Q7UPujtKGZd0
Tr74WAK4moZYGnXAY0WBu1qAKkXtxhb6Gc5+BIoRYh+URBoKhkrliy35us82sGYfwjgt6nG7Btvm
Qk5DTXbVDyzg6i4w+ZDz93L8XP3A4LztrzmVtYOqcRltmXQcN5qAp5cWYXhc3ZxHutwIKhYBnGx2
qDgEHeDBiSauuDBZbBfYi/wwP/5UwPKf6L9OjMoTCyP+Kj3tCm6sWLRahLOWKGAsLsw3tth6alpK
wwNpuReFaOrTIe9qWV+RLupymxpijHYfqzAZA7JnlzjeHvvCOPnc/ZErhndQegyZ/3Ixs+BQMk7V
V9VK8QYBEK4b49VyR3Q2dSNP84qrfi0hQH+m516FmEQ+EnqPVqfne0x+tnD/Yw/gyop1wqMP1CIW
LcJv3QUNSGgPWOQF18nkSYh9AmaCzQmFon/pJuQ+pCJub3L1SCTKLzlRbxmDX+MbRQHdOKrD2ato
Sk33IW+LmgQy6ebiqvbbgBQxDeH3uAXmNhlP2j3tIvYI3fZvGuzNIOdb6JJRALkVycTJDdO6VXPo
W/MTKnuld/exzydyCJQ+1Q8dVPoKASnGpeBr6B6Ez9s2L4bqs4lBPBJgMmq+PcTkVY+3iusjrTgY
fU3lO1Re8LiDFYikgOvqPitTG+omBZwKCQM4sb/AKVRSq/plCsDN3EFemRYniDWGUWC6zW+mKj+g
X4sK05OB82TnyWztfDev0z8s2TM22xWqI03GC9oMwp7jMLx1kRHxu4UmlJeyfT74WkbmQZ+Spwk/
oh/weg3e2Pgax66+q8uZSRepYkCwkWRpg2m/vcsobB2sQxvR+FzExry4IartcX9/kTTVXCYHuixm
YyfyUJJzN05uQCoe1bzdQUFE6NcMC/03qFogWxMyB35x9URUYvp+DgLM3jqOl/10BbUe1GZtNpNV
IaZRD3ZKXBxnjOSXjtwf/LkRQvb8xyaTedML+uE7wufFWx6b7BG5xzAF4ncZquz5He4+js4/5KKE
1e7i4sevGVUbjz2Zb3EIB+dmZ2no9OFi4o4Kt4EBbTisM0HnxNQJXJbyADw1DuJeI6bz2kThePha
XS3b8ROAaMjbPcZn+E6G4M7V3xGr7Z0eBvYoBuOJ8Ch8ZWfQOEJBXnwzRaUJKWs5I+PpcaDca/Ei
O+qXCTMwv1HwGtmxCirjVcGBcfLxlKDOJw1q0a8vWpiRUbCLJqtkBGU4FZQ//1hZx5px51JgkHR6
WFK/xxXTAicqGsBBoFAFbRvS7Won8Te8zv63xhhvgbrBoFs+/vdkp20sHUwNk4rNhtmSxs6mfsJA
n49rR8/yCVNAOmArEs4u5JEbB9ty/pzyPslyuKNEJp6w1oYTZ0nZs65iJXUByhFf8PQQM5XarJbj
X0o57yHozs1SLnAcwia9WjXt1n9E+OEDkRQavaXm6TbmukxcjwXG9KaTaKi7zJBmbEFf1xtKqyJe
rb6u1qrDxgJPGY61J+A7qXbnHXog+Bd1JQjzUkh9SNcOFCthZzAJucq1/Dh4KwpErVY51iL4FOfI
DI7q6/3RuDq/eyKwL+RAN2KzswfmvYbwaL5cQrI3iFhBht0nilVm6jbuKIPG8R4LGyx1vUE6Cht0
JzTexY9dtjZZ5QUgGNr67VC8y7DYgJKA5B9WZ2pY84lQbrgmDCbvlsGvmNfh56qtZgoo4pjdwC60
CiyBVDQNPC0YFyYgq7kVDoYkdAshUIxoDWAldhj7nDY6OT6kHog9XhlMZ17TTYWE43fr9q9aSioZ
NRMDn5BrvAJJfijB5JqOfcSLFnnWUKOZS7BoDDBqeouM3JhoGkzHaNxeYen79eh2S4aJg3tz8L11
o5Ade5PfR5ARwgibRELpoatYWPby5aho46FQsVRULRk6b2U5ejph9ygdoAruQtwz5B5tRhIVSEfn
Q6XBMn9BpaoZtt1B+zfwl6SgcfhxmTkjvD2HoOpivG1jOE2KGiymaQiBBS4iQkhKp52k0M/TlDCv
FMr24TajyGgcwrKDJv2GhbOICBWLK+TnW2RYu2CNv5J+bRZAH4kyKiMSTu1W3SLQdO3BZp3FhNNW
K2276WGQDt0+o99s3ZJRIT96xixfbNRMPubbZMWU095ywafMJq+0bOTmYR0/XDuG7eHz3OuYHwTS
OqGmiOwMmZMErRhp1j80qfPwFeW+MNw332cYiO6/Ef8z4fM1vMa0Qsd6vMOs7S7tpMVjf9ysFfvl
qZSy0zDYo/4WVk9fthvk/8/Bw/WSFkz+1GUwrS5dtwg29v2+RUjIp4bXrmIswoW6hAy6d0d6T7qC
2/SlwRREWvEecdmONiq4OMcAhqR5g51tXj1Trq0I4HyMW0E3xhOWj0Ug1qbbmhJy9OgwqniFXxty
MqHBqgVtaotYtg8+OaN7ibEzvAO4yV3XIl5G0s7/3VaLR/cwSCn0ScHgYJpFNfqv+gT4spAJ2N6Z
1+FokouIWpVVjFl1Mud67VOOjPsQwtHCbdo5gvdKNpfOqQBj/plh5pq/JR2Vy7YxIs9bL6qsEKyD
Fl0/br7pTvCsQnmJwDxwtRlmdOGDMYqg6Xsbp/HeD7IUCMAmIqhhLRl4z4lmWnA9ii1Nf3Q5Eqn8
/p+1z5jhHQmPXxFTll2T7bAkRmXaCSQNCV7wW7/BeqMyTMKZS7XkaxmM45EfVlC0xnvILUWAcc7b
FJznOXUhp1bFzC+3oTIWkZz013zUJww1o7NaZd+M8qjrz9igwoa9yQE+qHkT+JQYmnDwnuD66FaK
9PDAW+lQv4ieXYiYizX1xdjiNbcD3pBN0VmW0otRtC/eafiWd0j/EekTDrDhNlgISDxjoiuEL6fR
7WF3uMNCoFmFNNr6nwVWup75hcd+Sa8v56JuCLn6+9xwEAXgfEcxAYYgJ6YtTE5YHozW/MQkM+Z8
7tW0WbZoyl/l3xyOAItjmnZTW6Mx0kQQJoRQ99nL3DXrbKqPlQn2PWCYRRG0b7uqSw14ULaD63tc
mPpgNWgP01Hf6vWFfD+HVaBYyAUK3U1bbYJ77bS0FuRkPbi9Lf0w7ArfbrnQtVfH7G6SMvxf0DSY
jH/L6r0enet4RnKsO+/3ji84sbHCw/9isdGjxU3/S9nknmh/dPA+2R9U7sLtQX2GsOQb/FjOC0RC
9ZFK92JlCAylUgm1ptcZ07HVqSyd88eqNefoJf7aFh7McGU3dpEQts/kLPJAUAynHJ7xr1hh6Rn+
EdNNBPvlok+U/rCvz7sdmlEo+Zq3/+kEfMYwRu6efgOO5mRTeasZSdMgxyIAkQUd1b/c8LXncevp
3+TsFkLfMdp3D4GfjTwZjR45ZSVP/O9e8htfsdliPu7W5T2+XBHjd/Y0CXLLMZFpVoLwvMTmMPP+
zHRv7ICiO04506Ojjt/HCliSJhjtpyTXp41Na68+qrJKJvmjVdYBvQGiUm62X8QvYsUr9RcMNeRC
ChSMILNTS7Ir6XcFPAwk3XobXrdsnmXwOCcZpKPi1AdH2gzhcB3Fl5x9pvlqeekkbK8LBQHLSSAj
1Kq8umZtcArCMNph4w3PPFcxIsYI6GZtJOvg7Z9IUK535OF/U75Mb9VHUrgqSC0+5l52gmulsda3
wU34FzajDSRahAjLF9BNb27Y6SJKsNPWbW/2QlmBg3xj/MzsCUmbkdSo9lAAp2yv4xgJcpEiSMUM
xZGxOfi6Og7RqrknvBoSMzkagP++fm3qDmYuGJaV0NYuJ/M+nrfuXWCzbvcWp2RqjgfGJPjFnMeM
jZWzJTe8oEwAYPZ9+x2veud/fc2HLcdPVEF/qcO7LGusUgk81LJLS6Wq9yAtOkGAgA0j1v7n/cGN
xB6wh/G/yW5ctwwOPUEE2Hxbglv7eASzYI2alNxzFZU7gZxgIDkx8jUmN5zCLld9flV+2kdl4EYv
+WFqV+A4KQKt+lbAvk+gonrUKqjvHFUfoiiGP+L1WT3WHyq0vvXAHO9kZwJMfkHMnU7xyAXVOOea
w9Du8hAsxdACOOjl5Api8IM2sIEpGjK+HktoJnWeJymwpqs1RryDz/7ObVaxhyZXVY8ooWLRoKdX
P/apabRX6bDiSkgBtPpBELMYmf6cvnzzI95tTSf7o0aJmsngp51Sr38CcKGgXylCpcmAa2RvIwF5
NBshna2AmZTZP7EZBsf7ah1pEhAO0G58AVv7ibrCTjBj8hGNlEMTOwzhKFgNX+lmacA82rwLWQ0N
7sk9aVaaJXJ1QQqFHZz6Q+MaUUBj97XbaovfG/QqY29K5Tofkw6VHKhIramMsRykBkGZLjcBcQ1+
JChOFvyRdc5CfzUBe34QDHy1hnYesrdA084vy9nz0P39VQYaLLt1C0AsmurBkOc75BV7TTL8IfTv
tZ2RwMfkOsWGtCUmJXQr8wD7+MVa2acmnk3AnCEAMSfyTJyJnoBI0s0R1wqtfCYgIWRDOc4H8b34
dMMNfjygY33R4j9DNCgB0FBX98N/025qEO4B4KL6QDo0wk8rECl7vWj/WfsmknUF/qCwR7k0QeuF
wba6D0+nqp4ODiI6jJffaG0o+yega015lgSkS5kZ3yIMrT4ftABD2+jtKdNDOsBBaQ4hQioPpthV
D/OiWDJrVvAlIRZcF9JEGz7OcF+H74JETWELUtgykyPHs56RFBPQ+0z2hYhBsc0CYEOGFzWc9JnD
jnSnuankTo+jDscJRLbSSHX9Ri2QNZOmPrrDsQ8SghI9qSnKpHbSxDCFGPWSSJkAvuarYCCWRQ2+
T4Jk+vZcrx8ykk4qoRppIpBZ6vPdIOiurWz/j5TVc3WO2rmTkdPvNP4cdxiQ+o14Vj0lnhV62fSI
z/QF2cFpTpB8QlyLADegyNo1UArH6cFyQE3HJaLbxgV4QzWSWkrz5UQ74QfXxzXoPb7maLl9tCTU
oy9crA3kBw6NrNiCYwxyJZzMg0mihQcd0ipB8sHuGCISWJeU6CgKBuB0bvhCOqf4wlCMHCQsNHUp
NiNhVG8io7Oqhiq+6ZeBOunUVARtQTgTNKWfXAryutqRKgq2BCpF/o9isTZCs28gvzxTV6S0cRod
Mcu9oQwtVs743orblXPSPktE74r9qpHgB2kMQqPhnSBecGbBpK0qHXwP2rp2cMITlNb/kY3QDXDo
4+1LfqDUTT1BCs3kkzvidusiXl/xfql7P+BU8aW2co5meN+XJtxZhns7rokeqVY6Q83U1PWqpL26
drwwIGeZfgrPol4Gi9aG8ni5c9EuGmZ+5NwvIp6mKvOUfA1lJdiktwEYx4/kdwcEMMNw7saCGb8i
Qc1GsS5z7DeUHfxhLF7JfGbkJcGVZyGwSf3ryKDcFi1Wps5BAAcTRtIWZY5IQkH/5KibFpiVcSr3
+sIytwCRf5nt6/N5mY31K9hS51KAvdgVAUVEqa9ZQXbDamGV1mcSJoNxckmSmYj5lyJszOdiiU5A
mSREk5IIJSR/fIN+3NOJoas2KP0pX4VBwF9WbyHzuNJl4zbnZAnusciRJ4wc5Dhe882KssFWfkGH
cTNYL+/jE/Jj5Z1/4T81iX6tH+yl5AqFoGccmeYgYufKOUrui5ykrCrqwzr077xnhEYGkGIwa9Yc
MvbRqMjq8p7V/9EG9+f4BWvjyzM1Tsj0QE/XnLoWpd+sPUw7ZKITdPn/gxboenF+VgQsCLMFvU7L
/vSrm3vLnGiQpxfxty7MMnL8tEJg2urMq53tHaG6wDT8RXBdzxDJHlLWF5165AYfPIqnLSbra4UU
ePxu/pVIjhVG28wxn87OKIAMwKrMoHm+XO9l54inM/oZShoAhoWurfsAi4RZXEbdutCk/cy3FbxM
4dqWI11UM1GXBr8tk8Dz+hAlisq63im2WdZYCDQdiMyOeg8U12zjiwo08LKLFLGdPBY8+p/jgpWe
RomyrAXZEVsfPHgXiDeXBMv6JzwnITGPDBuA6b8G8tDvvaDelbKf0+4L7qxwb/5duy8WZaaCGJC7
F8U9VUjwO4E9TZRXooIMkj9f0RM4EP4bghrqR88le5FIPRRlOjXODY7Ot1zgb0cOcuQLvIAcs3ws
2SI13QhtDmOlbyrO04HYNpqpLVEuGlY47XAp99e2Z7Lo11cE4HADuOvDpxF5fj5rHFbhI9D5C1MU
4e6evJBG/OCT2ZZiuMLc9L5Nowjhw/12M7ExXzkr/BAV5x5kyQhF8pSu1R1sDQV5ZE62NIm361+q
/xEytYw5XW+hDVww1lfdnDKt2giBTpq4Dsn068IQ09mctjQRH1nC6h/cB0bDww0LZaWVkUgmbrgh
R5o0KWUPCJQ0FCOQwNOseNEnDSxDk+4qWttWTRMHN/2j++y1ZatNzDVzjNS+zyB4StoeD4FBH/RU
sjb+wZEpXmP9IzmE4+ZNwivfmr/vCZzI6eRL5lH2o2/U0azccrO49sEX7EIh126G8DGrvX2lZsJF
e/xQ7lgwKXOmcuH3xqcI0gHJz+frYBaG7sTyhJE3xZBGl66t5bVy5NnSDPvRnK5r9iMoQt/4B01R
2zSa2RWSNZ27zqNy2GOGty0V3CB8VTXRpOz9BO0zWeZapMiqN5/6CiT2ciCtpRZshyRwWRHgaQbo
yNe6x8qWyaHRkC0qLlcxHGML5b73vchP8adfsLQQAVOBPLyJCBaqgeZyUxuMQ2EjN2bDp2hffzGX
px9v9kPH3yrlS5x2Tb+ZzMUYdv/WsGBeCJloNWNaufY0DvzH7cPmn4C9J2QvF40fUAzQeB7fQ1id
542BtHsRQLebC8eSgLL5koWOO73tABk225+0YUXytnoQbSKSXCslRfVWXkMVGoZgZ0LFtYIpDJdo
YZ325l4fN3sln4jYBf/FLiOTyNK95gNkfv3KirrXtvUZP8T9qgYDmQDoMpjyRp8/AqsQGKwmzXU+
ZaLU1YWWDxyGqrlhvo7EY3ztNZILk6w36MdiKvkNHvD45MRsTJfdkWJGgw0tcQqawRIIeN65puvC
6nyOtp8H5/u5Rz8Z0nM2IVYpGU0HnZ3nt1GWKiDYIDpCfLSYW5q0HsOEx78PulGm5tiPrcpAZrFm
MCKWCgrFIpcZJQiQ8BYGsxUAGt/lIZ1TXAe+QMurlbGZc9580MFgz/vq1zNGpk7ey1zCs0qDfqa7
w+mlKOL9k4u2DmhCQsNdXO55Z7DPewDeLoINhVGBOJ4N8vwVx95k9Z7i7AoIvXeJCljqQcRsjWGL
Z1CKCHxSNLGeBXO8f6KKD0zcWwCLr5bpJtDZ5ppvGPITgbFwc2SW7/YAp/RAHeOeSwHtdxtAeU1w
gsd8uAR8yCHx4r03P6jnbWEV7xFF+mR6Enfu/BZoMDn5G01Oj22hB7t21dY1qpZgMbRkgX7Ke3ue
8y1kzW+xg8o6eCFNhsZQemujMLH23O8t38xheX8QnxvbtpyNegl3YvrB7n2IGQjMBJ3f81dIT2lD
eOilr3Qs2ghnA00brwpgRHMAqzTlEn9M/VGVEEd0T8/WUdkeK4izGzJrEjj5UcAdDHWEVPPDjZWc
dGQBNcyHOesGaBnubB8lZagj1zT4geNVEenOBqJy3I/ZB/qEhlxApo55NU1TYES+pyMSsNv5e9g7
3Ca4kpHIDevXU25zl9TJNRmEfkoSOTb7mI3cGcn2hjy6TVR1v0hYB1fbJcssxwxx6OKQKBjLHE3E
mKeBySU+KTkzIFSlZTalRXaHudHr8Bewh1YZmnI3r2+xRnvULu4kZv9PxONdjW8Cjgl/BFd18/Nh
l4hoy09VTw7wgIgi5EGICm7q/Ruc1saYQCUvYo0jhN5PpApAfcTf/10tCBec+SMWeOKTZhwI4T4W
PZBymTeaoq4L7pliZYjtYjD8V+JHkG/1NUoD4zH3sWFYUG/fMFOM12UmXl9P9LHAo7HTC7EZ6kt6
2oxLF7Z7S0KCG+Fgy6Ndj5qhSLVcUb0ZAT+V15gaspTmUfypTD4Te04HqWKV7xTF3ke6QrjqrrL8
YBr9u0JF9o4DO9lhFY5TtcxmmtYlXKENXvPy1MTxF+lBNQ5P6vPDUtO3K8DDYm+NgxFhb0Dh3L7a
ImFN2IVGoTS7LkngqTEmPhxDck+UQyoeJasnwAds2rr2G3lapQAC9JNsZSXTAw3EJmWE6HuHcOE3
FzBRWTS6UCbr0ZV9db9s/6q0K8XV05QqfRz+/MSeMZQ/hiszt3vyQf6/3WJq5NKKn9ZX2kcaQTbS
cLrsf589VFqqux31Sn/i6d9r7SBOFWkw8Uk0dn8XG6jtRNmMEA3kiuFBaM6aQ0gU3ugzsiBKJCCs
tcjKZNpuiyIcRO1GjSv5GZ83ELZtX9Ecs8dxTvzZ6CuaRn192ug90vZF8CV1fAJLxl97cKxmosOz
TbW/QWtNFcMC6sLbQtYYRSTyKIsVIFAFPAV/Rfs6nYyHX0/CViNwR0FdPMBYCnJl8GUZmGmb/1Pc
+V33+ou4YR7tKsYTJ+ka71++6taKkiqVmDXOVx0DPR8dxiE+xsANTwVyka2W4+BySNd4aTfM3bor
Lys0N6isngVSDJgPCReAaZjJ2tNUCC/wYn5/f5/lXkZ4UiIhROvLzAPpk7lrTptUPNj7j5GhU660
pgRh6Dy4d9ltV41jW7pDgdxFZKUDL2UADRSgrLkLBVbuJK4tqaUh0ALqc6G+w2YEQFcMAhomOxtm
9WkwNdlJ5Kd29vR4yyuklKdvXtsYsAXMK2xowLAQ9CBQSLljeL/7EqC/E5A4Od2SAA4RP9kO0lWC
Xc9p1u5wIohUd+0Z+sB3M9KJr0F4hGmsShZLIFd/tN3M0iKWel02tSg+cPQEQoS5ImO6kZi0ggme
z11x8mhg/yGIRj28CdKXlHQvf2fKoEPijR/Td6ugEvgm867FD/eNJkj69JzesiRgcCAFZpPfoszK
AZpxJLSLY2kdUUe1hZYGVhHEOkg/cSHyU2l63xA7MHp6dld7k0vl5cTYHqbx0uNhlLCH3sFgkMGQ
+n6wEdEbinKLoNKHzJ5RaI1oAkxcWbgTKvdr6HbBuAo7UZp54f3xXLLpKka42y++EKwUT5g9tGM8
cVwkkEFPKlf7YZlZCtvaTpi4kEOP0T9VzmDnULDPfaRJg42zPJbeyGVcro4sASFjSH+P6z9x70UM
MnIHn8R/Pdh+lGxNDiMseJPceuehLHgXoHrieCic2eLpp6cZ0ttVrRaRclKHjW0wJz0Y/36zl6zp
q7iI8f5S39UJPjtm1pdOEgR7M7S5TDTg3OCGiO5R9Xo+L183+DwR1VAHPVjtOQKSFkcdYgDGQcLz
VQz/7dRKDRxqATklYOUGgR0D/oUrWec9eArXo3EmMfYp8iwIKDTql29m8/oq0pHZltjb5o6pmTBP
JdMj8u25vYj9kOiwSGLOOb6ovEvGRXVd5JNPxquhaANH8WqpxaMpiANTABJSlbmxQe95cSv3CZXG
Nbzas6Tq2wiwLyPT6lvzz/fl7B1sozHQTgmrrnYSiq3h3MKoiHAe+2zt+Ct8knFu5IxTGUkv+MRi
waO5nTuCj7fihRYRBmUqPqXprttX8h+M6Snpe4xwhnbDR5Bn9g9rXGh9eq9BGs81Ez7QO5mEhNqi
/OmUfX3kGFb5RA/Rj+3+/iegDn8KjedJFAWII0cZHF0aaLdPxK+PvzMQ0Dj4wW5jWXgoRqKR8W9M
Lnf07wnAuEGS03PQOYj9/U0ZhWGGi9wMpb+Qxu9RunLgX/ctSAgPEk9SGwQAKP/4VptaF9G7zx+l
257qXoK2slyyF6bLY7qW9J/Q8m5RO/q1QZfY0Fib43rgrJ1imQD5SClyxkk5ayAAmgmfVWBfW/Kf
n5fvjpW+fORgk5cPkWXLTzXtgtrQaxBSu5U1wJe9LxcVXqdrNNUQd4TeUj7y0LBp66OWEA+gjXag
wyAtqGY9AkhSR6NBL+aNFiIZKXanWosa/QxdEj8jZYN8f8sLEPv1CQ7Dk8mNh9L2Lr5AuiIHGce/
fDIpqTNQWtqNBty1hqry/7cswd0fS4ezEYhJANjVf4wsDrAO8C0mO5ih2L8t9Aq8iHi5j0UiFwze
qVbTKc7FZn/utNywsoEyVygpbGGPEFot/PiGKfyY92UZ1aVjWHim17aiqvUiHuToWH3Om07KsGNM
MP/OAOVCO9GlDHaf35WHnCXxsrSsVnewoGHUaXjGN9FAvntBZH0oLn6jl8eXPKZ/2Ym+kekSACGG
O2FWN6iXfIbvfzzhD6Hjji+LVDItNjhWj/BryQWQRrTAdeh9n31xkP1gB4Uke5CHFncdgvLTbvrf
K+WeRTb4cSKUDq0qXlqt2lufdiyFz3X+e2D9A7kE+SjgI84JffkvFwH//EfRj3WzsEa6dFqmt4bx
jetLYypZPZNBXVuax8IVBie6gW+wUxxhq+046Lt0JxPOIvipbT4vaj0CtYrniEHAmFwRt2fQrXBe
e8CveJFQj0SXtaGTuRE31VV6qpIzN8268avBEA6Y1b3Sq7FLXGkcECAbEgck50MMyZ1DRmI+w/ZX
1pd/DCeg94SAdpuSTyJDpsLGkFrw7iZQ/XL3GNf8Hka+WVi5h+QQsmrRGVZo2W8ZLwUfRMiyoZnO
bdyDXKAvSWbqHwfpUuXQWzZU7VwY/C74QS4+eCW5vq4tq2jCjd3Dj+ayv38g+N6D/iX3ak2ZtCEH
LuAzRVUlYEBjgkxK9uub0KaFFGi+WVIA0ZRj62106ABdp0X+Cau5si8dKYhKQPUWkpmhKTb2aZJ3
lq20yutaiVv/UT3Wg5fp8NcLjfopyPF/uHR102du8ZuVbmZ1OB70Faw0N3Vv/Xk8hH/pwgPrUsRX
ld+tam3wTrkiQxDhZTGydx8Aj0CPbGg9RKiHWsN5WPHtfpU+DHDGSIZg38/+xhANC5irzPIU0Ztf
UfkrMjGXJ5CFNxNC5GCT8RkbNZLMXyLPBF3MMasnE+UA7NI6TKL6jjGMR9/yH3RzdjjJiEuBBgmL
0w+cSk2YoMMGX55cbp5+lBw3COARg1HifwbbC6i3+PCT7/bD4KxXe5z+zmryKSQQNiBD/h0AUhbf
i5PQcmx1kKbZ7mQoKOtRr7VlFsdmZMtgrSo82gQ4UQkZYMYFp92bU3xWagYCES/tzojMJu9DeI8q
Qwjjh3/ke9Cwk3kgxApa1o6mzs++fq1oPrKjXW4/BOnoP+Mas4obePbDPetio7gMkv+PL2dY4B/K
Y4ZlavaUQQcIH8wv7mytY4jq6YQEQV9qosEBY2MJpxgsSSiUaemkFJedgTTluAkVbb6osWjCzlEl
+JPadaWGgVyCQMRziBNRrcd2z+bX4BK169FPyY2TcCH/7wvNUsFt7Y6gp8Z09VgMy3WfT48qltkQ
JkXxi4st9dxBljOrrX9kVRxNSUO5b78uKO3F4ih34wOkAG9/D1z2kPS0qLOcdfy/dm33k9P/MwjM
Y4H82AdcCnrIsdGN7adK607Ij9wgTbfzpLIFh3u88R86DN3HY0VLRR6PHhXSmZ2Tkk4LNN7eOTxi
Csj62HpuSQpX1ocztOwJbFZyK96TNUgRpiWiznEbGIhZ9Ky3AtpZ6Py95EfOWAxU0SILTEsDUXxP
78687i3vnGCCgWayfp62BtzuQbpqCsKjqI/ZhYj7Hudc+hJ08gVJyj7QU4f+kANR1q4JzOgsP4Q0
8o4aw7AqHnc4BUcBrWkFbD/Ovn3siU7aiNFzOJCzgMDndMRux7aYbzAqF0fMEfVvJrL2HAipSai0
66F1lxhAZ0ZM9Sj7hGXPsNa33dwK00iUY2huH+FKorotRGqW6LMWqdZgvcPZc3+c7LgZdYKxCd6+
zcfzj8PDJJ4pXaOf9ggqekP1MNVGuQcQ/9asp6uBKhWRZmgD2Z5CySIVt+WIGhxIvkXwNDg5Mfai
t7qsHal9YJrxbesayXghAaP5Gerg6IRK9ds3v+bpmKB9toNGbsAdA3DVcXg2K5PSBXPgDcOolGHa
NKI3SY8Ud/yw/0BlmK22sIjHs2DkWeOjI2mMi/UV2QvFzPBdPe1BarTBiydB9vy0MD6IkDv+QG6n
0u0x0a2qNXVk4QN1B6HE9gtkaS5DFiUOqIe13KuFOAqI3f1lCDi+RCW6xED3UXRZhVGwec42Y0f0
KTZp1cRgayYMciptQZYyzYNhZ43iJiDWzI4Jnb2Vk9pxtlSo82b+EgEVFxpAkYmNNMQDLzAT4K0o
pH6v/VzbFIVRsU1XuGdzFy9C/JwmvR3sNSSXEInPAShYL1ENr+G2ZR9M+c5ZsqOUKr27WBzw1qaq
+3kmpl1xwZZoMUG7q+dvr152NGGlENYEbuALWYj+4mWo8tMQIKpWtFH3Fp+5ul2XdMVd2fha7fl8
YauBQifHdxA1+XRDEgJYoQEzUmfuQ/sCZ89Qk2PX8ZnKwvWTU3DSH48LRqbzY0kuOegb9WOLnbw8
DUdOyjn22sy5CepNQJMzCHOwX3Caa+11zpQIbZIKiVfLKprENn7HLJK6sJZI6GWGUPIUBbGVeF+Y
M+h+/k3vt/tbtxYb/cdOpfVeW3EdevZsX+TYuwEUrwOLnlUhyWU7loFNN7fGmlX1nAGk0n+pTx50
cXx/is9kFk8Qc5K4ZxHItjBBFUmK/gWIA99K2zxFK7SCMIa9k0pTFKrjhm5j7O5V7m47JC5TD9kH
G7IUyroM8SIOGIFo0TMo7BXlRMGXzuwi9sl5+z21fCZlFQ7Bp9AtllbzLvEfuRvm6/kD/iv53ePq
RGHyhIIsXieSc5jjAuZOfJktCZMflDEps5tF2FPyEwDXCs5txVCvMEVh/KKQyZsoNiHfdG7mPj0Z
+QI6TJDra5DhZbjvUX+tgVydDzdXjplRRy00P+/zwocJR9pN6LvxwuU71bgKoZ+H/8AUFJYvqnuK
kAlvRRh91UOKqBrBEJZF/bdDBoOjb+eL6Gq4EHdyDXu4T1O2yEvfCUKbIW5uHLQVD7/WXmpE8dWx
0obT/hhsifZKWFwoUzRN/r8v7TuhRJiHqxbWLbv4kzi4PoQqpF2i1QM+72/Ium3JNhFTxQShezwA
sKcjl/0FtFAgB5XY5lwQinwyKW61jQSLYnlA8AA5/9HjqDjW3XClEdkLkwsSgWHGmiJueObp/hWp
Nujbku03ZoNbe1XHuOGe1KVBZviAJYWbn2o9GugSn/DSjZd6jYEXX3/UuX00EsXoLkaaUQj5C9Sz
nk9Nn5MfawYqFNrKogfGwFSF0hYGgmGaGuPmcXPdpWbWjmr0U2P4G7Lsz9LXv3fx+IIgEQ5Lpm16
c9B1nq2TubBOlk+wj7d6fB47AK9D5cKu7cCzRCfQH4p/9thteyZb+rEYNq3u4N4Cu0ugBgMqKeae
M23hMFg1a24ADNi5LHEoPcbcozoQGrBAvT/9Y8r1arIketXzy1TOqVcKiZgR4IosAwcusQI6UA+O
Ql4aCs3a9mGwfjLK89xCNx65tqhV7nae2m2MJYNHJXCWs8C0aLq9C7a/xCVnIs7agyQ0tnItLImN
G8TYtlz33+2k+3c04EEWF4MmeHVMzuZH5FRV7okL3dRG+hSRGhUIyenL2d0TOQbwurqlWWXtSWJq
Yh9H42KYC9IfWyEgZiQvtu3C+j1eRpN1vPv5eVYlMWBZmE0JFDIVDeb1x9d9J5OGmWsX9vBhMHAR
OK2xK6pYh/V4BRRNgf0b1yO4wgI0toGHX1+4LLTl3SMkaWuGu3OOFq4BZrkW6LOX+2NU4TcRyn6C
uWSsGOnxnAmvk/GObL0SJzkbkMWUYa3Zg+yvSbt7IOeDaxwmRyAxur5vA3DnDcFRUcTAwL/ZxRiL
wbvBy5KIcGCQ1ZiYEPvcor0FLkl0U8vMBKVlT3pNoFEXfIe7cToTUCj+4VeqZi/CuJyxpzFiCWDB
EGkfENLwNECSWwpRMdf3Aj4eI/IdMzMA+uBKkb5kA55B9rGjAO1m7w5+ryrMwoaYIde385VH/ujs
7LPRTakfCeF6VHLyqhr9L+kLc25/d/uHOtnhkQy1HuLeM60zfA6WO5Yi2nyje6YdFBnbojrpIVLf
cMSmZsgmMh3wAwThMYRlswPiW8PkY2q+riSY3V7JnxTwol2XbbCU42aJ/fGJI4wAIFzW4JYqWAdO
EkLQeDV/VHFEh5eMT53s2gHybcZGWU6QrmKtZVzaRaxxWUnvp3DUA4mkIh+iXNwNHmBGIwtO4MQP
EGsK9hZYC7b8eLVr1YwQUeFS/6n2rSymxQyXIhbqRMTa6xdzhT/H0v8y77uP+4PEsSmZXtgLee51
PiF4HITQRIf1LdGFwDwdbW8q1RlZOkNYSF2T+mi8H+hT4ZCGqjFE0i3RVp0cRRD0ZW2/Ppq/ZCRm
PfB//hsP4QAN80RyvEy1C/wP3OhPqg/7YGpYvfG8fZ7iMMzJCxvdcE3FWNSCimg3KcPRaXkKKfPe
Nz5ab/ead04wzYFmKiqVTVbCUyxMrig1ZndmMF3DTnUhSVH9yaNeQMopV79Mhh60iaCG9iEV+qCY
wm94mwzRG2dnTwKUloBETpAtJ2QYh4IA3YRBW5KgdQCMCbkByrwzltLdam+Mq8xlaM5E9kocJuvR
pgbEKRGk/Xb2a2LcfKDDfB1t+Bg6/+suiwbo9V7RPgt71EkvKX6TFWVD44/yQYbiiKRYZ47DrkJK
hA+Rqf4ZkeNmTq6YWLHwuKHy8kyqco9B214mRbt8258IGHFCJDVEJODtRIr7aFE+FmUjDScRaBur
RQTmncNEQhPi5GeiiexEZrfpouAolfBOF4nuRBNG8lj3ICETDxxyv2FZ9QcZ91BzWo/F4Pnzu3+D
YcR7FHefNM0M4pjBEhTFzgoB6+eX0sjCno4lDzc+5KvZc0ikTlHIqQIhb7nlk7oTONELg0IPjPBr
gl0pZqrc1SrqzU59jaO/spAVOXd7A2xVQsniUkDbzuMoUsxdtEj9SFZCpeYIkY+QshVSmEnLVCK0
F9JPdWUEMNiKlTwbQnh0J0RZY+WqBTvL7AMxYO55VjZ5zyV14WO8z7efngSTBnOxgok9304bUp6X
frk25FtRW+cDau00Eu3FaogAd3FNuyGRKe4ihvVnp8615M+DuxJAi68dDL6jZp5NfNpwcT1ntD3b
S1qeoeH//C7mNzL6zdaIHCFvBbW7j28tdHZU1iG1lnhNDTwyvauI5+2c9l/8/jrMNiEAzernOpFA
eH9L/FQPvf1On/VzjU/Pak1yvCbv++v6wAdPPEJ27LWXobBkxuiv9TuYiNzdVTzIIObHjmzg5ywq
xNBbdN9qK1glGBeY5HgiGDylxN5kYeyjxARqYyMc5lAfUpc8EYxEK/2czpvRIZG0PNnGjsIK84Sa
3a4ww8BsLYAnnsITl2QpkrsxC2d1ApZcW5iFpJyVKpenm8hWjTTqp/rOn0yplLrHWjmu/wXBVN/J
9Vh6dpesESdVDfSHa1NIFLxp89i3k5tnbrlwSqnKIGPlPYh8mbue/ij6LshUJbwPNTS9NoG5uCwt
Lx2m59teFvL9x65u5abeqGMuX7jxWUjN4PeqPPojdyjjbXwwoUsL9yvF3MlH7hkgxET0q86Bdfn8
NmW+yMbaKZE9uplqqYHk+1cEV4jsZWMoM8ZjkgmlH7fKdmwwzXiZC+uZ54QC1WzeE1Oyp7tyS0io
kgw2pLfOE0w/2UiSYuz1rwzq0HFr4fi+29+GcPDfzKN3HN4r3SsG9eV27bga4lcX+G8v2fmOHEjq
Cf5CTKZAS/ICQS61jwjpz4xBo6VzwDD1jCVIxWncIGZ3q0SbiZFxuA4kmA4CYfFbN5f+o/xb5Kct
unE90+tjCE44j3AkAj0PzAzUsFhqdMM2lcxfVLfPWbX9EiPHGEo+70t8MLc5zjJx0HgkeqElX6Pv
f+s906vHGGq2bcS08d7S5gFnnXmQrKiVwa+n9pBRExBTWK4R67Hip/cvIDbdAc2XtjBiJM9NY66M
3XAnCsGBB0zCS6V2diZ/rrwt8vC/rXc7fYVVXitJB97AG8Bk1U3x7EW5/rabP3IAt3QT0CryODTG
VdvJI+1iZrcu4m1tykTWAxkkQfpr35H4pD3XWvqyyTNXbuuGwnbj4s/XJPtMB6Pps4/nXTI+QWNA
jn7tJtnvMDueXkFMkNnCTxr4IiF9lX+Q9HvywQ2FAKhsKWIS4YHjRMtY/pYlD579dXmq3ulhu2Lq
zgVBMSwk/ftNpt76nAUHA5f+CuflkUrS7ZgxGgb3HQNms3FeO14u55TCV2//Wx9ypnWKpzJ+oAe5
pSWtaUaGMACQ4sLr2/ft10k9wWceTvo/gJCxn24JorKiym6/Of6r6ebIEfsBqkY5COVaRfCaqnD0
nh5JmSZ2jhB96IVsofL1i51xp1KERJ61k8+HQGrWlp5dxwdcCghVPYrj+R9aZ/QCsVZnYHSdHdCv
xiseIOQRI0FprtOF4rFz6G7As49xWsFfFFCQqM/L10vHf2QtYCRbaA85aSrjEGLprnb/tW70v96E
vSOo3yei25piSSG0c9ZmjvM4lVbz45UM7RecGAzo5HK7jpk9HtlBG8JEYwucWSpd6xshzlIhFMIM
kFji8PJ7UMSYvyDG41xGFQgjYZC4LbbzAxArNyf8Adt3hKLG6QDYy3cCSY6ks0XJnPW6mIBg29kp
quMv/5PAxjiqi0CMTg979PoV5h8FUWajretxmbQ2GDF5Ee0srrUeH/A7ih7sjupibTqHEH3NBDg4
o9R71visopjK4LJCkDXnAyQCLTDYO36e75Su79Z+lwBwXrSH1YZh07dVM0IDIe2TBMLcX0ghLnDV
ZUpbwqfDNkqOR3FE6Lg0smeUDQCfY/FdX7ukaZNW0SWAzc4+lL37P+5B4UuRPYpNYO+vf95ZRFT4
rLlkThYXhNLxaWKs2dMYi2XATh1r85INHjcC09bz1ESxxU7Udx3Kzp5/Zda7fAbtkb0aMlkOFCmd
9LpJ9M0j3Cl6+Ee5RpDpssgy6OWe97B4YLzHyhx381jysSHUSnmsiC6SH4wAr9I2UpSlCyUZF0w/
mOKWrpW0HUcd3S+ylSKL71ruABNpN/EPHcBwMPvSC3e5g+dUsqgd18Mte4v5lHilSEaFpc8oRUHK
CJmE5DL+pgqhcmSkfOR3NhiHU9Df8Ka/nPMvaXxv6IjTeXBNDu+1qF7HnqruTX7eljUclkyZvuSH
K6smsyl6SvTxAnauq5qVVpG/4L74/raGlpDP8rAmArbQMln/CkXwxOHg8xNnw3AAJE0PRHy0RL1f
j+E/AJcCXkoDqbTAdkHbaur2z2tGPKr78WsXn2nTtAIA/owsVnGyt8+DhSkX7z+s+VFtme3QKCzz
KtdLf0rRarBotiWAgZr80B8pMW7ZHS6YN3AhATl7iI9xwjqdNteqoTcbg/gxAh7eJPcobj++4yr/
56EAbSjoSWFHpzsUGLj3vn7EBzah0f7clRP6OHNRByGLyHV8/Wk5W1vX/S3MQOzKYIH8j9N8I4+O
L49eH3sBy3COXOyV1jiT6OsoXjSBcBAR4S++iZA87TuHTxQ2mualriGHHe02yotdmuJH21zODb3E
Rngr5u512U/S03ZzVQaHQ6vqwIGyoMqmtNx9drWwyeJ5HA44U6RkzTc8nEOPFW0fxTfsjB2TMYAz
voZQMnMj3uTgE1UHmAtIfFuEvvBr9DQC53Uf200lVgOAW0OIUSRrrbGSmIdrfW4s7/3T+mhjTM/G
PPValug9SHltID4FZ/s5VED1IusCpBq7YpRSoWZ4UldO4OZ7tlyB0AsrBpXMpTacjWdecakV6IcO
a/5Tvjd57PY4DBibO8fURYEXncxqJlz2QBl/z5z9NlLuF7JK54KabHHroyknaILfIBKAcLSPo6fV
VqpPTW63jcA/YtZNSpsKPvYmpY8Cwf4+/KT747XJBsFhC6pz0B02ueSFc8cCQz9LpE+QSMjPFY+0
znMeIaE8w/r60rsuCUqotop96ClbVQyM55LQ1I9c1aufoNjHuc9vpBzqvPHTUFI2IHx0hXNRjjzs
X/mNttKoPq7FFzxk7bvujgparJ/yszyQH3+hS/qqcT/uC3kQEYcGEHRCIPmutAhQsvKlER1znkyG
a827Vwhvd3fIJSwpD/eN4oDrT/Alqtdydvs3wqjyk13mbAZb6xL2j3xYLE3Fi+/vUAbN/fy0TwMB
QqUQNLJ5UhymWko3U+bmyxkphN8w/e5t3uokIghT0lXwgZN6b2yhLC2aoD0oGt8zHnadultXhTTF
MfUe6EzQHAPx2nb75sdX8QOy+9t8O6Nb6HNVaRxAEDheu6HsAF/VbjPIFty0h+XnQwBCDlCGTAJL
ECZK5ObFS5ADD/9U8bDiLYwJ/Me75XKMbmKBqgtLDcgK+CBRr0HJt5hX98+8Fn3EOJb60ap+XZFz
vyTd/5UAQ2FJNXHPaFZrOKck1skNqb5Yvn/ExFBO8jFg1HmERvSdCHeKZ8/6yHvqDUBpxwWsF1e7
3sOcxe8cfzAZ9V9dBpcyqyB2SGel+UbUnOWqfUsVQgETkdIU1UEtW7+k8uzvOZQIk0I+exgCR2w3
CYHERV272QCmcDL4cpymrd6xOQmy4WVydQ0D8LUoh8ajUEjkKHupxyTNldBd24EOb5TJ+Zv3td7F
oVNoh8REcw8S5eo4ZNKsagO7T34NDItQBnrEP44AV7F4N2xhvf1MkhJL6t2ZLpYjkg8eO26+pS6i
KSC3fYQFWZuxoPJW6xNglp9R80TQgeEadowqwhYoGXb5GvRFh/REzzKgjut6Xq+udkOdQHAUXyjO
zhxtbEjqpsZKSqPk+E3rt3ZaeuuLakcmJFwjZYWGq6Dc6MD1MpeMjdbHxY/N71SYVaTx/V2N0eCU
THAlu5YmeIKc0Siq4BP7IsCb9aZNhYY1sg3DZYFgRLJgEbm64S+zZddEj5GQ+Tbv/pDkf3lcnnKb
Nfxc1jVS2hMCqo3vjsD9A/AQ0MKEHbmGgsTxiJXGQxlTeWZNiY2PAiCSfQneKr7dWFkwWBxwJzXQ
5nISL6IO72oqvSPSODebNV59JfSuFH1HoWHN/voIQpSYTT7NHjiv5a/CKgj2Z92DcItqttFXgcbA
mOCKZGD0h0IcSw3+vDHQK/rkSBDvmEGxQOkHFHOD0SL0siNUit4xdsAQabE82AqS9NfWiN/UbY9B
YNvbtXHoqiRgKZlvgBkZT6Kqo4Dr4C2/WIzPwKblejc/70LSyIhokecty3mPhu68P4EPKhEQKK39
UU8iDQtr0P0d/GaZHWKWFrMpsY0vIE6MSuwkvn9jJaRJlH5qliA4a2FfS20OrEIm/r+wGo8woPGF
Vh3GQPb6bHzS+0xk3EH4CB6/72WItXSYd1NNky6kGUvIScq/L32L24KqAb5kfaWQfsB0BbNayOPk
YsHOkMolv4H8Sx0SipfOTXVyeb+7kvncvDaSewtX2xg5CJpqHhboEnltt3D9MfF9Cndj1lcs1yhz
5YGPtdqTaMCYHz+4kTl+t0v8btdPGx+sO5nqU9C0xfsq4djJVR/1hK4T9y7pLlWAs+ISYwDlbnX+
UNHdIJcCcV4nNYhFuQsfTkw/u3bpMnBH2KZxri8W9Y1nkyndVkSsnm7fiqPeAh86Vn3ExsF3ZEWK
dqLiVLsYBqwZQrWZS9ssxLIpRG0g87vuzrZx+KlwQjmMU9S1n5/NRBpdkE7obqnPNZ+cwH9O+55n
hERb+vOEpjMwNXx7Hsm+Dp96uYLqrTesYAGn2CQgAR1cstHzE3XQGpFezHhpjgJkxbu47IRNI/7r
vJIWj5QesKVavKhJL/6BpLQI+uhdFQYQ/0YK+m0OrXnAMkOqmyNGrzcCCStPW6AiLPxQSlnwlKWX
hsGAc+ML/tE/9toxGSMXGg+NNBSQzTNw+0E9VwfC+ejAUVuWUGGfs5eao/btL+Jwnr2bHqhSHusI
Ld/foJ5fOnEuxzK9m4MaFIfxbgXjrp5E9tHMKfG8kd6Y6EjIaBK89FdlRpHKK1h4wJCenRwTyz47
yZ/fA5CnbA3SjHm1GwvXBavzkc2J7Yt8UaE7RgUP4nK9sdhKnZ5ydsxyLqik5yl7/e9oIY+qBRd0
Gqt2snd+MwW0lFxz6shayeGakJhVxH3R1yOIPbxTmflJpKkxxCxcZd0JQI/cxjUKQSRzkeeedcBR
UD3fAsnG9tzSMTiF+98ntylPxzlCRyvRJ/TGm7aoO6yFplvd+4IxEKQhHRJcgnKInpncIcgxRXFG
7N1VE7i6Dnn/bvTmgYyUqJlRpvBMOF/Rn27+L+DTvZIa0vBVEqJBeTxMfgUkR/WJb0Vnc6xNrBda
Pflmne3UtcDwH2RAyGEHYLcyvYqAPOFb8+ieLGng3prV6c4RSROFfU+dR5HIwR4V9GP54GynlqKl
KWTh07u7W4oqZbQoQM97zbwRpICVT0ClMuxuakaAU7LDHmQe9hGFzZGRDV6scG/jpky5Q2R6Jwsj
vugi1pW6DXaeqk4kyTfv5OdWcAL/C+P1XxuGoR8zp2SvUUPRZG0l8cmpAj8PDwN2QdEnQCxHDr2R
ore+v7r3PiQMDWD/RCTMUEwCJHWd+2aPa6xpcwf1OtZDLiq7yeCDnfzpGcrHtH4bGdnasp1slL9o
verosZPoPtKRbkDCQODuvIRJkZwledBGtmBjDfife/9dWJR8GDUhbhKeCOt7Kf62bURe10ylZ/bt
ipusRRc1TbQnv4bdOtPWok8ylz7s3ZBpapQ/tPk1sbggybNU582U4X2WG+4Ve/Rj36prXd0AH9QT
GjCFfoy/Bxr1xbQb5LQlCpsuQzjrhydHTvVs1J8vfAPivEwoWXvLnuzIIqFOfrTN1RG6LXdBb8ZL
XkdCAleqtg/BdYegBCWSyGplspvMvA68ucCbE3okRUPbUjJTQiVeNMl9dBn1ahKoZd+8zRqxFl67
3lNbIEOSvhSwSqUpcK3igivjTBP101fhuEgstLMtW2qYw7+QTYdssqCsHMuceCV3Wwd3zXE6EzM+
YYZnz53l59BS8tjwYMRXRLWCv1kVgQZW5zgiZeDJZSg4aqWiWnUCnubpVoEP++guvXPPs90m4jXd
oDKuh28HBOG0ps5c0IduXR4XC2L8f6y5wCMfdrw3JLlumTc6WQIqc44azOu1kJ10iRSFCDjqpG0O
rII7kPAMihgoIwtJVLGqchFQQDloMJFmgXzLL62ZMzhcyZ+06qhKEatYJ1wlpZJf0w0D7kbNp1Bp
J6VWhl1HTCTkwJO5Dw1F0I10l5khbMGMFGNFpe4AfaNrVBWKiLSNJtH9+LS8/2N9FrNVW1njPLZT
bSIv8rsw9A41Y5acUwkFwui5RWHlc3X60mwNd1In7rXtpAZN3id+mWqds5k07MpyaHygp155TDdq
K+x2jilE2Va0D7FJOZpGsY4uuxrafopGmDJhZqpOmw7/na4c+cF/xIiyvdiDZgd1XW76r6BMTlqP
TSBOP036IlRYHCCYSK+7kG2GgLgz0HlP7Ig+Ey/Ffjh2wsiBJwVVM5ydYTedVwNLkBkNPy0LxDG0
fOJJWxyMcvOOw6S+L8kkukwx2SMpFNhiHUZnnsaxeZvlHAph0NhXDqrQNl8r7DFKg5vQVzukXZkT
oYwlI7MexrwLbI9x6gBdzUWBDSdQ42n0Nkh1v/R+GUpwVUu2I1UXfl/uD6yM4a8DE8QgiU5lWKYq
MZ7PHPaRxLgbxH8YfdYFTYd3kSD7v8eYOfCMsWHQH2+Hz0Lh0InNC0cyv1zb487VaIlCD47fnITa
w0TENXPwXfxe8VYfD1/KzIXrdj9OyaXeNg6gUqlpVN1RfXc63f/dVNFYnQXuLEVZcS0vQL92VTfZ
VmZtYLkmnj99s3Dafx9R1tglEYfPdXF2MAr0cNcvfc316q/Vmvez0fkdBADUDmMl2+ueLomCd+gQ
VxDAOH4njFk5zCttuW6rhhCx9rtMraq9CWQsPJ2xrUpe1I16p76vylQ2UHd40ZFE20QE0N3/XAPf
f/C1xUZKhLieb8dZCTLBHlhjo3i4XUvyJiZh7qk1B5j3+uuVQp6WO7Yw2SlKDxrTXkcLb2wNoDJr
83g8FxG9PQ/BmwTarRrn0xUBpvjUfqgVkdess7IjLTk/bL0bIIYkuhcCWIxRd1KtkoDRy7b2i/QE
yjkveyT5xoy8Css+JGf3mdPryQyrIrprCMEl1W73/9U9hp9Acfef+5jpGxja6rDvyvYTMeOK0l59
DU+ayYMrte/HtlTC5lp6gGV4RaNm2Arj9xggjLcw+5DIoX5Rs+ILC/pe0et4xNoppMLoSOdtRRNu
jE5gPEyJMFyl0EZqZGt8YZW6WyfWPu45bYU2gPi80nYg7JR2Azf+szIwHan/e1EoISlTTw5wCsaP
Vbu6mv4R4m0nr3Mu/WIx3T+AzwgyWRl6qvlWTsCqr4bnLM/8PjFL0fe/d8fNYBwiyo4M9tGZQQT2
L54GYI6/uGWrm1pR2rJjNT/E0I2f+dd4I9mH4iDQ2bkBX8VKOCj2evmB0dAAfQ8xmTDB2WrH2WcA
LOm+Sq+EG7G4yLAoo033zHQwcaQ0vG+pMP9AcN+YW439SFaSTcv/yfsjxeb84LxD8yuUoBYwd1q0
po9+O0t4vCVwo8nBKEuVrN5S8LBfwfzkWCx1YfLmt1NZMEdkKl01IfbMh+0LXT8/Au4Bgi2Rwwvc
YWScn3flFC8tdX74OctzoZyKvIycVb8zLiKM3/mwJUXxgbx7lis4/THQ0VV2NzSeyz/EShhLoDrj
nDPyPO06MVsUFpUmrN3jUnTjkusuAXzLYsI2zs5VgLQHWS+CVMFkwud5GAY6Hioocq3vlgT3WD5P
G+dHvnFBzRRA6lyTbC1/yHbx4gfQrjmM+9CIyRrPvAy7Ivoykv8HEz0tR8kdejm497qgpBsILHM+
NYWvaA0rLx7Z4eZoabEY0HOG4WN+xXTJz+gr8xK44HJHvcn84izAOkLI5/Fu6nNbEWkDLRmdwhz0
EDluoPslhgt+0AD+Y6AQjX21W/ToSbLd/pfSXWUJeg0M3f05om7GAt6z1YWDzkSUNTTmu6+oeD3C
IlsCTs0TdikkDwdMQ6UfBlCq8omYCjSp1BUh0a/mmL3ifAPPJaUTCFVkxwBFbewa85ZVQq7XnByW
MXKfISKWoJpRD6YOAs6ilhgnR+n/zVYHCeTsR4w8zaqIkP8pZoMGZe2kO10lINo2A1SqF0ISmXvW
V+iONx4q4ETrmV2jqxITO4P8cadcz7OmUWuAlTEUxB5ypP2RRTrdGSPU3eDeLDwcI48FYkB+IpnN
sm3PSwMacnICgz/w5VqWcQDVsq4P9GsUgBIYQCLToQ4zDARvFDaf73OQVOo5OUCK+EB+wZmGUWEE
kOoHsH/sXFkaQpSznay8U9jDKwTCU7o24Z8ygmAM0kPVDfMB9J0Cy05OmEBGKQDJYCbhnYI1JzAa
EKYxB2XL7PF8XvRwjsNe6upkNuNUPNaaoz9SYGOPwaSY75xBaC8LDw4BRvcNOPgH3p99ZhJCPMVN
y1WI8AxFZ0dO142qHOElnO0QipBiMcRyJj4CX53R7UFd3wl+XdSeNhQceTZ1YPSQ4simzHZ36j4q
KDlhTb+h0zPigUPTMfENK238FaqAj2GCZ1xtG5BxU/CVwhxJpvQ09rLt84G3KoUcYRt5jH9Fv2Ok
bSVMp6vRuYwVcLWuTxvp4h1+4cCPZkMM3DiMXffWQ1Csq+50CHCSfy9Kbzg9CLoTgxlriw27U92s
EF34PuJX5fWCt0I5EwZemoC+aY5f/A30ihlUZ7sTYWSkHSGRzNJND2zdPcTIR0w+BokTzFD9Flp4
WoP07+q00EAxqEZs4FmyWehfw34xYKa/gyzlYErw5qaP5e/O24CMYDe090Lq17uOW4vQRMPiByVU
YVb8qVRbGNcEh22Re+P6h4E2LExVYvn2EX0VzacVEC+S6ZkcVwbhEtdC7uLJdPYZqOMVtaFYcqZr
munD+yp2+17lCkO1KIVtal7+yXTitFMruwHBxR4s8+027ZdXzuJO/7bTuChDjFdpy3Ol5AixA+Yc
oJNl5Rog0gaBCLTPY8CbvBJh4MRaQL7fGuV9qVaTkocq2/HCH0bu47sd9h77FjSZT1okLs29r0OK
hHh49B722eMLrw5hoMnCVuR+XCPulK4OE1y6I2BuUK6flU/TXXF8XTMmMXozpCAhhefmSlMd2uIV
3eqT/x8YUln6F8mCIbQ7Dorz7V0VcD+64Si2OdCL/V1QdjOCBSpTVY4vNfr8g5631UXTik6J9FE+
EZunYgR7dMYLNWZw5qdRsAKI9OBjE8unKiAk04TQ7l89D+rMpUgM+4EI93Pgqmpl9kqwaPanUMAB
LhNHinO8IYP23Ocq2q4i6scCHegX5y2uKZ8FWPiVaZscsx25CC0CDszZYZUG/TUk/L+xwhe4sHeA
BJ+8u6z8wwGEIgVwSY7MY1n5tTeMM5ViaYGctbUp7kr8FRESx3biLS12FDA4W6CrQ9iTdKMcH3be
80kZT2vZmw9s8wlAFk6YQH4sCYckMNBN9yX7008qqFY0AsaLgQuXHviYL6AsmR5b+nn3yxZJo78+
GH+reNsvlwAYyie1C9/LRKsouOQZcWAaVnTj5XyuD2fZa4/SFvESGW2F1mz9GL2XpI/OvrZjFrnn
TCI9sOL9A/ac9XvZY4t+fGR3O6kRbxd9+1Gv8ik/4dTi2iP/lBoToIclcVVarSPzZ7Hg6VQrb6Pr
Oxr+bPX1iZrXlTtHD/IZCybstXdxGFqmjO9nxnTJZfkjmcRUrLSRpMI+TqP76NKA6uhKiVN3cgbM
nHVE4gaK+8qkRajIOwIBeKWIlD2v3dA39n4a6SaB/7o0MJbRVkkMnkqzByQGJhPsPxidbIFQXCPY
q1ymoJi4OyIHmD3/li3JRbxbr305BUfBWtmckyWLKCND6WE4a3Q/bxM2lQz8N6Kvizctjum4ExZh
17qmKcUkItkVJCKwluPtmrNsPUnqB0LXtBfoypr3bxKPH1NNjhUrPs6mYH/7EsXcv8pQS4b9Zw68
k5mSDgay5GypG6sQ/jJumkz3e0dSvFDoJVbvDTpMaExZ66bkBkx8yMdl8gh9bDjOWWp6rSAT1yQ1
6j4Ya5fFWLWFnsOcfFlbjxIil46Em2OTSRAE8APdhL68Vohkv3udFrXxTmHEXmBKckW5Mth1P0Y9
sa0N5q+ibVMqkqGWH0Pm8jthxARKgQ5sSNmoR1WDL1/WndKVcBk4GNWDFB7TtLlL23wenXGfpACx
Kku/O3mZHSHt0LG4TswMESmHU1KKcfhdkkGYVDocYdBInXfzkiUX75qyegf7pW9TRgxgObQuwi36
+B6iDqGV3g2dNHNtGtLnLq7n+bfDYIWWoXoZr713daCzCrbsRSRQT4Ik+2/tnWYr57Z3NhhK0XFP
usraoU9X37ARY+qPC7HS66GpN+ylPKof1WVjwdrmNe78S90CIk5qs8KRK3li29TRK+x5uP0a9axP
6FidrDMuFuv3UG7Q4DQrh9H6o2qIAy2EwqILCwm1g3nmJ2yqV3yk9kKcgbuAWkiDCfjuZQl7xRj4
Ul0AaycF2BxTug63ucy8OyZq+NqBlmLjFAzpMtf7yhM05cFAHl5Al+KUYP0d2fmJqfm791ZTtZ+2
9t9sso9V+2ySwYlOgv65tFYe4ZLu5UUKSiIXZSb02ApQYIUXKV3GdO/KA5WYRQ+2TEoUXbK0iv4C
VGIoa0bO4EAscHAyKGTfDWjagG31lFfQetDk2HREZv34Ri3dHlpRKJMm3qT2a4c7QKBhvZSp/6mt
RVOUr01/eT9vjv5BIF7ZVZ5q+13CX2VSxlxUEaX8JIWIuft1fO6UHKsHQ1dSjTac7zX7GzSiWUEe
Jbh4H1zcx2TvZzENGP/Oh5Hx4+wq9zRwNQ+8Bavebar27uf40jf00HycEsXtr08cciEr31LnoBxn
uxGrEpn+KuytS+yY40pN5/dNiALFjPNnUdlVRYZRqMx6d1oKSmf+qqwZI858xFcjzMK1/Sm4282N
NTERhh2rgQui8TivicX2VM4ETcAy4UbXbaiEf1RRdeZAD9bxDfanLaFixEii9TDsX/bqouJ+7wPS
PclIh0qBR89xIxKUcAm54M1rDmGhVzlWp9wTsO3ZjY21BFFl9mfdV06IlbI/GyZo3gQ/oZe6R5Dh
KWe7Ir0xbSnTK9WvZ2Maa0TtEOe9dvBCC1IgYsDIqQR5gR4dOMNGbnIrUD6ycwGdPHsEpagpY8SL
5kqMG16Zb0cFaQFsMYQ16dIttfLtH4L5sVkTP3y28ueEYHkaSM2hhABGFqoIuPqRxeYgNB8GAZfr
LiDeez6b7tElrnF9C4EJfuH93aJtvW/C+nea9rNtqGAH41uj+wafX+myxjfhHaCr7Wgp/hKv7Gbh
JPUcxzvhPEC3JdCZ1i1zrcL1zvJkTqIiMCjEn5od+BhnZf637rIdHxAKOa2+geMuT4w16MYCYJb5
5DBIGux42RFQZGwi2RLv6FK3eXbAEIZ8MWiiAzre/TiTgwU9+UxRiHJZtMbN3E4tBBphgEIo2ZXO
VFuFIQgmlIkDzqmqBuAaeRCOxVQyH/YFIOFksD0FIcWobGl73A2FdmGacqu4uRp3ORx3DSolKmoB
JHU6F6FXwfiaG4QS6xDAzWyrsfoLuPEfbzj8i0Viibgf7bq/9zmbj58HEbhbMUU2cZ83WWG6w7CJ
plcgwEdr9i5lDgnmShuSrq/0+I9Z+V2pOj/amlkmjuTvcqWAJUSUh0HiAu60kWATshpG1B3XBMaa
WTqZS8NWnz3G783cW8IXQoVkX+RKFbjToeRWsmrf00bIM+GxxmlDWN/uYOIvZKDKG08QjqG5zOZS
o9uVATsnxYh1ZuxEphrWEIN8DTjJEP+HLR2kKITSeCyLXW5Pg5Y8eYyDANJGXyDts/QzMOKDlzHN
dN2d1nsAavqgDGzRwYa88FyXrnHqBNHBLGPwSXVVVNLQa52AgV5DYBo/FAi0OXfqnSmWvUuwpH53
cfrUifkOjdqxAsEj1RhwjuyOnK/3fdtbA2puuXav6Hm/ZKmMDLJHaKSZRScCgLurZMNeiaPrZ1qK
bd86MMpAtwifR2Ef/6Uww6BxPHVE/dvOm3Ep1sip+dLypbj+tWMfAir/GL3knrIuRtiviKfdiyfx
AO0xbKwWp2sweFN7lHpP//EbPLwjzpSga+/WW7bX0kuEYoybnbHr5BdW+QWx2iqSTf1DEI448aaP
law0YifDI5KM/knnFhQJAEuioIhhQJk9RVtvJwBfeSiZ+VxpF8e9BHTj6+Vz3FC8nzm3aH07fLT/
hfyZtY54kHQ6ubHg6elPzhFAc3W/IfP6u3aUgwTtCvs6S03bjBj5uiyO/96Fqw8bgwXa9axVVn+4
Q6o1uPMtGkIajGtgUJXudEhpZn/IDjd4n8wvm3Wh6NMXQpy0zvqoCuK0hBen9aFrCFdomPC/pWdd
JaBvlM5wVi2qKE9PNrCrRBZrcH2XyhsDFudS+vr9N6yzLv3i80Znc6X9dfCeW5tL9oSmH+W5E7BU
FADKouV7NjNNjP4r/6qoTJKZJpCUYi2AzYE+vXxp02d39+a4uOxamzLCEivEqD9GvXBfRvJ1/84b
mE5as4tnVK4BS/BpH1dMnRFxe88BD83VtBN5PNr5eu4r0RMsmdzLUxx0YrXIQujLPNyVerQedHJC
dUxcN7vuZVvPemGeLejUz8dLGXbCJSI+WV1IYUfB7BimvWAfTUcEZjYolZ8jnUXog3OZBHJ2nToF
dq11MSjNHlLwJV5xlxajVSTT4y2sbiSicq3/7lZmla1gPkPFiA4yV643qY4oYnT2SZGLf7kuLaXw
EDSGf/AvRYzaMoDfMSjm4oXufnQAH9YP3hmWXiTtFDj2KDFDIhao2bbi2XWmybEWGBBJvclgqSd1
w1FwulvaS2ScM0dMU8wEc4vr5/A0Xlo0OH+e5JBZktboU+3D4o0gJiKRbNZt3/M0cPtgDWHfaUvI
0r0YwRnvI3fpI/rG6kykKNDGg0SHqrAEI4s/Wp0v9ztvf/NL2U+pEJxZdjqtcmvUpfqmJ9RM23Rl
Fd+krUaaKt7HfnBJnqHm89GZBA4mHkJ9o6DvlSlgFFkcZfJBmAITdms0tc9BNR6fX5DW031+o9fX
PvkBkGsFZtNhWEdXnv9zndoG5axAFdCIkkcX2MM5EJSlkvNvGHwfVpvlXQw6rGLTcvXR78FJOrPz
JQV1nDQJ800qwvhnUmA/kn/B55s+MyyzYUiRbIP3JzFwCuSPb0kw2Axn9NlVBH1LJImhhExoU+cw
ootAoaqEGJTwqbHVTMv1T9+JLLLmYL4UYThZn5T5uCsuKV8lyJgqarD0sGL/kE4x3GIQV9abOvae
XdyDUVA6tAQPxok/Td6ycXXwQxWKbd1vsQGiObWkVIS3diB4E0h2gvtrX6SCa6AFdKmAeLPTJ6ys
pw0HF8PcYQSvZWT/NiAEQbdtInNAC/hV30Rpe2xsas8/G0l9QyfnOdscrdKpUk68AMZ/Yf4yQK21
sVbaJ5x+56/Nzdz39zUIHs8cWbxPZT0nLWJhPnZEb6RQW+EHdYHuv5UXvuMN6rOzMZWzFCkPLxLE
6Gb/rlju3pDQi602/cI5K/mhTOMrH6u/nBQ3qEjJ9MnaPW+JNL5L1RRjxr/8sYNXRJaPEc+KhaFY
BTR9RHMlFIaUf6M7aIveHim7NuR8XgTx4RPXdxZIrfjX6T64yRiT4EoKUKZRR1DlpdGDzJWun88/
87qMvCNk0v16kN3Ks61pzX2Yf+b4vLlaV9w2AdgLVANbbB108pYXX07CT3PcenJSZnwqWQtQeur0
XoP4ZzhgT6nwTIMhuMQUngiaJV5BCNXXHV5/xxaB05zz4MHPqyIqhVskN5WxltjKaU+eU/qlSMt4
xsjU3xrNWEoWxuM48e4hcMIuWe9J3kxwN62+HKnBRvFc/OXy3e437vPPkay1w51M6LH65YLbGhTE
Kt40sYr2Z71kHZYuEYU4MZ+zvKGDUD9ul3I/RZsDm7/VWmCUsV91+qm4IVS2dxTLbItGzBTl2Gnu
Jy/3kxA+iXk3tAbJTkMBqaM0zhcPO2wpVVaKuK3mINHW9ZmrRDtR6wwEksirZvZlcg4zpFYTLbzO
56IYfTqYA/aRh3oRYpS2V8+pZw55RJuuTyvx80OllK0aClzIwlHu/ClaQBak44E3d5gIdp1BcL1z
bem1inuUJM8BV+BaOMNTrIcoFvmHhG/DYFQaC04Vljn21jtMkH+W19Cb1MSu4a8MTb2u6lMVh7+5
Ldro1hLW3APDchMCU0Ud8H9bnL9TyhI41uhdnfaQxQSznrBU69C2uel45kwIP/My7WsNMzxgPbQ6
dVt40j3PtG1Mq+FVbfaWhiRX3GJ9J5cKj0SlA3cpYXdVHtcwWDHDhezK3fOHmThiQ02E1hr81kuA
ALzA02sRSWnT3RAm8swRpAPdKWKLjQAhgGnraqqU6DquSCg0qD086ymvvNq5Mj8YENV/Z8yMiWgL
IekbaCmLkDb6ei6vpyvlbZEu0El36wv7CuIEqU7MI6SFuavhf80oH6rSGznCVHPzJyiX3g9WQM0K
zMhgQ/rQjZvSEYqUUxoZ6jihEiIHqpjRy6yYxq5L0XbNYBrHoRog6xd+DGHvR4uPPec4rHaPFCJT
vWcK329bATjLRThKyuqrx8RQiYbCM4XmEgcCZQGP+/B8jEPAE+96Ms8GQ2SLoT99CZaQ9/LaQIUr
NhKU9x1LfIzzJzs4gsZIY0TX8OY/4SG0Nef4BGsd2TxSD4zmws4GBIbirhqoEhxMD54GCZzn1TJu
opfx9VK6YRulMnj/va30aWH3WQrhNgQkM0i5a0ruivYFDpqYZze26HQTcYGsW6v4B30/Us5t/lp2
y8kRvTruqPEttlQbMD/SiT4xXut8Lc7TorN7hzyBH11+TkPT27J+7pXnQxU5KfEiIJ9YwdwnaLJJ
+a2vFW83iWS+m7IrVAGJazeveg8jwhVY/usTVxEHVo22JVlyVxCqOWzwYz6q7NAxwvWy1HYyLjaC
/X7fAjakXtjNRyXdwozC0XkOYqDln/D0AHRDPnXHRKComONw0S2rqJVoa/TfEDvNHTw5MKiRLZfd
2SQMB5h7n7pAwlTOArHtPK28LORAnMUxFRHM5N+E/SS+3v3MVFBXD28oMDfIA1Ed6PTRJHEM6N3r
qvyp/m/UO/41GBUfhkIG5T6rkBUOnWeSQdK0H3ilaCUU7ODpN5iDw/WrFguFLBYQk8UHHdTpFYFf
PYxlG231pFIFTunSInhrMClLo4LdScaZUqTbMNZx39VvdbcmeCf81qjy1lqQKFO8VTbAx/tmtn74
FIR5LRL0VKYozKjXj6YTP9p28dSTTZjYUFj4iApzvyw4rcUhKiiR1ha1RwTljYequQyqm+yQAghc
9ElO8r4ZY97gyliQOpvwMdUy+0r7WbjCua4kIfSW0L3nIwi9YblZlGsVklNBq1JLGsEjnbwTgJ+/
RsDkpUxZEmjScgB4uBhJPPYS3nfHxb20y+AoGnYMsDgQ4IkjZLSgES9RyKrEull8ju67UNM5ZJtu
WKpk57XQXRJY1C9QAhOfGmEyeXbZappECguLJG1rH0TpU4ourcSqlGWhk72Tz1otnVxp3SqeHNN8
xqhDtg0FcchTvNfKNtA7AbUQvLHMSp5cMLU+8gB0PULE9OYFQ6BBRRk7FlWiycg/YwBN7mU/AMaG
fYhPgLiv5fUBwzOOl9r37jnb5lLbXy6FXdRcgm3HHexcJysazyAOw9xWRwcmK/jxv5sGrDrc3G6B
aCNbA4LOVWDhMy7usHLc2pA0tBlrPjasDUfDNnthNE1WvhKks0vKiUGGa7znnadWMk4aVf7r3U2U
Yn1sAloX7R3Qb/eLq1Ie35QDcYiurE0us1r9Hz/MDqBWUVjoyuwH1LACNcebUmOYTPYs3+B8VjPT
GHO3hGrweL5L+vsGPRX5Zr5n3fbiUm/dOfseD8+c0wOWOi5IZBPnBLIb1yeCI1Qh4bkP3S+dvkn6
CEr1kWy6IGAs9OQI2vEZAXfmezHINlXpllYEPw5vDPdwI9XXSV7QmO3rMpxeWWssoHyD6V19tQkb
94/itSbZPHVM6V+8WkXkwQqe2/Z3x9wFAwMS5+2IqDT4kDqZXdE7+RF5vC5p1ppTLup6BpxJ7hBP
y/qXe99U/Aj4XRfjkhCMB+fj1FC39NY+3ESf44LwcMgx2U6m6z60PaSUppYgulQe5NN7IhxTOdnZ
e+zTeqyqdP1mkd40dahUWXOtPYXb+hDf1MnTxg4vB3cst5okCHnVr32IwJDMG8cRNdlYdP1eisSf
0pa59oc38j3FAjGVIJTdwkJwl4fkXQshU5CAy9EjNiXXuZY+prmwoGnzfKQutuFqkaS0Evrik2H9
uQVdnq7PwB2mfJw80HGa6S0lSqwdVlF2cirM/D8v/lolTLkb8x3QS/F9LRxUvHmbsgcjmvGLou6U
ikBVfhnfh43mCh7b/DHuiO0E+qIlIKpauEhW+dZAdAWSQZnFx6bDf4OuH9TN2rFdpkCXBhxZC8Of
q+jNpRp3Sgn/ljKX+T3Sx3YUXo1ws7rysuHBb3ort+aWuZ2bqLr2+QUOkk4iyKy7+WSau1ZVogwD
EvxdjEKfEzZ9gH4ZtvnH3s/CosZsk7+ROE2NhH65mkOp0KN/Eyn/2yzWJCJw1oO5Gxm6Qbfa99xX
nMmLQBx7sCosM97VYjhuwEvph0+my2pRdi0KVuNCj+HDjH/JJS75BtfPeglDnld+l4MZJPsvNEze
ecu9iWhipN63eb1ciwJ5D7Q2UFudnX7jPuEBvQCumPpKxYZJXUwyogjWkNRmPQWVdDAWgqUJumrh
uIyAQFD5+Ji0FTUAWhovSuin86RCEAcZPi72+0nb2iFwSDeFShE9EfQGRZ7MhuTdUNhvc3RNof8y
7NrWyPklogXn/xeZs1WpNM6pNv9dNB2NSWP82FYSuwrfsc34jLDZtHlEazeUopz7NoTWZsvh42fH
iHcdz8nvHwaz9/xmgWXTpvGcA5gvUaNwAZtha6lITynpoJQN5CPs77W3xT8g1sHlcgGffw0a+KCB
G3+JRm4Wo3T+1mPvbX/L6SxC00PjBfMVQFWnF1DHLL/DYWeObOVvO4Y/gB7R+yBK0peJ3kXcbqTu
zWNudsojZULAeDpmG//aofCZkGUDXxgYxyXuVRjGOIzrfgZqhSuzUlfd8jXmozh3CoSuGANOYH2/
Ml5Jx2mfRTN4msBj1rTN29BVLu+YYHeYdd77dY408cbxlQ+/BWO+4Sq902WFAcMiFIEX6wcZgFir
S1NideKY154P/ojjp3Xq4wb99rujVEyXuB51FcXFqNwo5VaoSJw0SMpqQarHhDSJEiGfAgulSCfM
SJaYWo35UpbGpiSsUQT/G2AgRTxfYh7nE/BlHW9rQ8H0GWJvYV45nO6L2C6sFFbwdJ/KWpGS/mxq
Kz7/zW97rxBEkDJpTWbABpGlTs6TivKx97T+fcTlJA+99G6m/KUBZtfXaob5p1gCOWl3UYSoB2+e
6KxJiG5Ym733UUA8b19+f4JOImafUzlEabet6O8oSrgyvcQAkQznRLVuH/fPcFfx0JDJNj7dA6D3
oPpCDpFv5+GAdFh7CjEYGU9nxvfI14b7FkfbyIU87Uf/FbBYY5PMWr/HY6YUl0B9ZF2BGcpXlu32
OXp9wE7mH6Xb8WwibaR2W7bFfTQw8CDdYkYS2Wj5T65URy1bnw9dmF1kl+hf1PeBKQH8dyUSZ2VI
+M3ue3YpSPUNMf8g1HdLuGmDDKVqYWeT4lbeJL7Pe1yqMkY313JB5axq4hpApQ/yupsnfxFl7yVi
85ErUeZuzIa/psoWvOo9CARQIb8/6B00Ga1tsD+PLVjatxHMxDYF55I0QgmZcqOBDYNcl6nmoDCX
71GtO94Yip4Bat0a2jnK7jvHNfk0W5JN1u+DmoPLCvhB/KugsOjXSGvPwRfiiAaHo/S80jCFhnLR
Ge5dQLyrt9X4SAWesKh6CrU0AzmBq7zp2WQzpqd1rH3WwNbwLFkyRjKhjdq6j2DM453JNVd2IcKU
8xuSwXdrE++/lBjXcq5sqczigyNoFlYpL/WyPF9BZisHUzqKVzkm+XBdmv8WulVq+9A8LuxuKubA
oHzv4MkK/Qc2wPtQfzAvEzdqRHcpz3UXrVbC0JDMJh7oHz7qJ9QPxNPT53tzB1uFha9ncrVLKDJN
UBDZVTBIFLEMvVc/avfmUc6u4PjxEL5WR64Qgnvg3JQY2K5U3x43heORdTtuXCMlSho1w3XXMrzQ
qeFRD3gpkL3iix9x0XXWLwh4qHLg1jhbHQKiX/GikbFPwgCJ2xJnkXmhQ2zMeqUBSAZ6cpMBW+/P
jnrz/n+ij7jnOqPz/vEpnwhGGjP1+/+oM/MF/JcmgU49TKpNVCBq1WyoPSK02OCxU1UdidSdWlB4
A4A5kT81fG9obgYglPr0nieePVduR3XYSA6lGA4i6jC78M9RFa31375eOy48R6UdfX0my7gwZbY8
V+9PaYy7irIHh7hnqe4xPh3oxSeo1/RtLTlefvxMUFILtgnMjHm+tCQNrpl92AKgEcgGo9cD1NmF
ddE+FebVWBGJrf/3c7QvFcWDtV5X7AY3Ct8WeH5PyYLC5jskuS2vtZ6t0Rmdu73G9sF7en7NH4ma
bYME2TQVrJCUAb9hOzInQBo8P5Mp4yqsWi1OSo4ZISYnwuKGQCVmUdBRcgjbbFhKTIIo2ei0hwva
HADrXd+RQELiwW1Es7ozM72glcXzxWxJvZgp30/P34uC7WYWu9Fx0OLqxeNorsNHr/7Y+qEpdTfT
PqO/YaWbl4CjxvGIewg2xwr4r+9v3QQHjjN/d9olvlNZ8z7HPZuWFLeaI7sNrBFcDh14XcGg6eVB
7TZFClNn/QWWpBI9Ew6dlWrwXqa1bwmRR4SmmlZHJYkLdun0f3ugsAm4QH9hmjsqCn5yrJHTplEL
cvOYWSmux2WSPiPvRGcJNexzS+o7d3KR9BJbLohb/a4KGkjCrmIzd/ZrF5aDvdzcRNdDSJln1bjH
LH6K8+FQ0VxG3Lbqj4cGEjwbfUL4YU5biAGleZJrYk43gSOzIFSZA35RhPRyNNTk9XkttNDmVf9u
k0qg8fKJ600BLOThSmO+OKw1ImRMOgVK/jiwqauPt2/+K1vhI5R+msDElUNwMir4n/IyTYe2epS/
MMs95vXUVpfGSJDl7EzF3m2VHghSJzjDS7baiBjm4hWjderM+bJbozH/pasej8oQ7F+FA3mnQwUX
ubdEQ0+xccaEDcR9/ry1dRkicr9TYOr85u5AfKLyKhZ8oeODxY7zrXXmI2m6+v7zKoAoeu3EHHT1
xZMw0qPsGlHIVCpeyy6LQ0ZA8ymXSXM42/DUk7ChkOyExXMbD5PS47AwDcmSHAoYry2HCvyObMPD
ByCnZmJkOQHKNyHiLG0XVSLt32r4nooX9HoGnE2BGkFoYUrKaML6UTVAle1ObbtABu8iPlBk8opZ
WqT1lrjFHIXlIYJrLqusBUlIVkkzow1pY/fXxX0LceaMin6hH7wvLWUzAjZd/pqVqOZZzkLxEG3L
9v7zNVoDQf4AaLTtRBjFNhFk9H288AGd9djVfT+WXMz3M/+FXHN2BDjM2wGQ+0zis/fEkO5XBLOd
tf4k8unJnU2ZJVDD2v7bJw+20S1pFnLtsHHCrfmyfwpLULm1rGzStUC4T3jvLpV64Yld+XKZAJeo
nuYhCUyRz/4TX/arPRUBms0+A30abOsXP7DAOhqyaFXJpoAOljGeARq80FjP83qdpjecEzgghJBJ
UuuAZl8MiJTjReJlk4A66PeyvK2xu3hMmClWsLGANN0M2G/5d8QV3LkwCqzInZqHIbOpRsiLkDrl
6ZhsyX3LU8/+yXnKzZhzgVWXhxha5vvPCGcFC9jVoUPCQkxZokFWO/JSsnvDirxTeQPxXO7gcsrt
o1pKhZVAlNsBIv06c3ajOo+HlKsUMvLJcDieXv5yWCY3eT/e8BLgzgVp7iiIfmAqj4SS4QTLvbbv
DKHIm6ib1sw4zWV5A1ag3VVZEisBl5wm6TuE3zdxWRfJxERrCJYVfXlFOvqi1dRJwzU0x8nDRx73
A50id/xLgH5Wq5Xowrpbi/3FDWWjlhhKBZEsuzeway+eJy7KZS+vIosIPj1HXRSuyRGS59/3hSbV
0Qkt23hQehj8KNNVPQGjUG0k31Tf1HNDIoA6NdYfHKiDeoLkNm25gVqNjF+sBbBifybzRpP7GaAU
kCEJ1JGy7XdQNO0X784AtasyZFttsHXXhizMUsgy3l8caLaYRA0A85dvoyFPfqMOzczi2hg3I3bf
6Th2NKvXUcSVRlpXx1daQMSvFpQNpZfM6haZJPNahTGK1iwOpGZ5b5WDUECQ6S+zqHHr2qnneYIe
8L2u3IXH+1Qv5uQcFCXowcoeEE51ikpEW9Ps2uM5kvQh3ZaHxy/y/YQPtcaV/9AuRV1MpCgX0CJC
IRLIW+ZBspA1B7CWqrm0UADg9EH6VcSCBpvZagqRUwSwSLPrJhy4ONngWcPa1ZBL7wbPBuJ12r2K
fdZNTw4xC1yNCXYV8igOZpOQRS7sJeTUFTPCpBaLPozDQpqzxKNgMDd6BaomoB4K+1pP9PeAxJQC
fssZwBnkw2Qshdxubjjs6HMs/WHR2XmbkHrYusQGd2PId9hfONmL46mppZCmJMNLbN+O9tZQtubJ
CRL33pZzy7dlExMLtyg8ASCLb7CIN/TqyMlOjXuxWJ7cNktoq0yOPlygOrxWXDv/6+awgbgVOxhK
YCq6iDyRQR3oA+/STOmyxF53CmY8wiXc2otvV35poCM6+gzejUUgU4lZGj/mHFncz/oOeikIumFJ
jx9p+NbP7ZZezXdf+uZ/svTtDQRqdceSjVXeEBIXopUhFRde7nk36CL71OvAa1q43xmTIPFmoT7C
mfeSpmM6pUt3ikXHHdJLyHJ6QMenxvnvpg1aqKi//UC2hHgw5gp+wXRkO3ygK0lxcgq5J50P7v2a
VLEUSpBHP5Om7NgIhB0q3Uw1uCI2aVg2ef932cYzRH8N04x8F6+wHWseJpYgYclhvWQRKvB5Yxvd
vlds119TMLSm6FUkXEK5GcxS3ma3qJdEeeg5fWDwaGpv2GKymG9Su0OtfrNU1POUhe7k7lXh0as1
41Zn+OU6Jwkrs4kLRKh1m/z/BojxV2gX6wZLDT+7wKV3ObmHPugakzaExTdL1qO001Bp+AcLIncZ
QT6rhLCUT2WDKDTer6uI5Lu+ZervWtbxfue/yUsjM4qY9G9SWCvONzBV9qtgPxYq8NLQOlJxq0Tf
7a9PV5bKUoNfsbiXgxQ+a370EPgXREXRch0ZKb23467Em2R3/z+9k1MWp89ULDbYNwEtqxxSGgf+
IM5cN87ALqjDxnkaiVOUXIfgqz11FbmiWVFBBl+b29zfO6jRC83KhVWLu1sFOffL/BEMKx+8S0Yi
ziLL2IU3eq05H5xcMroBjpH17uYq842+W5n0FMle/MDDqAH9AHsVzZP3/trD/xyvMpCMQ/b90PNT
19QBpUbLtUuCPeDmtzvsYMYilmaoxhZl5URgRd+jLuBZULraihIBB9dH43eDDhyw7hemb8Daomu1
onsbTMhT92pf08LmhzxwMUInSiOyRnCSd+nnDs/qF9lLlDZc5xomeBb1JcpSTBE5XgB15clrKgNT
DVa/RjX3XIRUdnFBR2SEE/3rZrSmUrQFEbwpZshEe9NePQwdDgctUSztpXAEffr8lN94Rxx4eRCW
3bwyRpyAi5caswvRvHt36n9UwrN0vsE+R+UZ3Tt5F+1c71kTU/qRKj94e9F7tjix/2I693nNT5c0
O/Ii7FvXPRmrPWZaCue2FgPiKS+ZUD6r84CFwPqtz5WZ9dW8slZxdiD0QxuVf0lFgVQjFpKvA8Nh
BIq6hj9M/4BQ+5JueewmC4en2FBFLANRBKPGgNoB/T+1Wup/nbcEbX/KK9kxH48Owcz2JPSqD5xG
bDTLtsAaFf/SOx3d1IIfSxAkyEx7teumoBEbr+EQ6aHbjl8D5nyNhs93fctM3+6EBLdBR6UbYT5V
QIPYLNaQgiMfmTLQkepXVc6Wa5sEiu4H3gbmg6BKzmHt6J83kpOt2DCaJbapQPZHAxbSi3crGmrC
zcG6NmBe+p1C+V4MbBAqcIohLzS5lj63h+kQ9bmH7SpLJs+K8+xwZn92gNIr4YsLx+ka6QUmy7/s
Le91prMe1UGgpas2HjmilYVjoXDah+PJvT2Y5HlSvF8YCIxLxvsuBoTnAhKIup9/enQm6JgMxmZt
p27Nyub97029DELkSmz+EaoAxV/Q0QYksVlZL3vpfWvzeI5ELKwmA9didDhTNUkd+kC6PlGVfkAk
GvGNck9c0ZbBPWnLmLRoxnuZfrQualXIgyiW3uZqBcbfzwaanNSSwzNIxNkIpzbE6Si32xeQT3DJ
7rtjzWz88MJUAP5EYj/wPonayN9h5yuFWdh/FjSGxepg3PPN3HZgDMzQuw0ZYVXWoLXI35eKVwYa
DmPs+8zyRrJJdefn2YRhYgV1iq/fzg4WU9+ISkDGpgBj7SVIfDmjlyqDjTDraijz8JDhtArknrZU
abW1mWWEhoFi1SyswauKrbKN54EwsqMHfxdGraNCMMmeXuSHWeNN4luWi3gIWZsgk/1hTQq7C6uC
GUgegk3x0sGCf666rijK1kq6L839ei+26p7pqoakqj8xNNcT9dZ4vcbd0jmzD7Rl/Y59TNNM3NJW
hwiKxO0nhRPsD4qy0szhF7Nq3qs2wupVq3f/yi2YxcVRqbkNmtWRe9jyUtKQF0W9vifih0i3XLkE
sIFba5RqCKvQaCFp+5coaGDUpz2Yz2zAK8zGb+3JP1mZTdkCKHEN/6rafQwRAhig0W0Fzr60y8Sm
oSkwumYzc7ysSthBFrodz3q0R6DvJyOjdnFeF0S6v+O9h1jKXVfIg8652rFtUkIUje+1+IBX2R8I
ZJYG62RrR0RdaaoVKLO/esr6r37bxME4CzwJbVpGggE2rc2aLGSnRbkxoiCnnDnVpfID1xJnHhu6
k08p+XsENTazoDvQrYSvNe9R9rIslTo7cLMUyLl3FTnjgF30QBuKsD31jVKwuq7ab74Syf/fXLZ+
RE4v5Gnj2dKrE1gZJLZ/JS6hcQeW7yszNGuUsMHzAbE5qCHV+5czYIdCS6DhVUo8PtTR/XrkqkZc
iDx46HQdjdUe3EWgasPgYJJs/8x48Qa4roJ0+WFO5uNSt8Za2a4qOjh665r5P/nyWXKgtjEJwslr
hpwH9N3bitbEqhmNK91uSmAyIzixhVoGtaeDjIq63kZdaDjSm5NsROg7/cbIH+HGc9LoyN2XwgGZ
9wGjaTcUzaa3VahkxODAKfklsdlvVn76fmTcAqTOM1uoI/mfLuFgyF4auSCK4cQaNK/gi3HdVLx8
cbKLgjpz/3euBmWm8XW6ItVhD7RlqzM6dM4Qz8mm4X8ecBw81p1ii5cVJJD0z2BR1GP14B5YqDGw
UPgnN/37VMh8imCZdi8zcUI9TTp+/TTDeaWHRPV4rou9tlL7vXNikc31dwzJeLZlH3pO3ZDK8Wxg
lRLCRhEOqcnjVxKM/BX5vqFIMH0BPiPiPPSJOeYH6VLlnjQxegVYITLe09Cx9OMO26h0SmR9pc4o
9Xdvp0zj+gFVtPBItLX5bCA202KqzW3Nr77sQsmDymIvIyAEndYlTx0s/yQ0/LToCJKagotZdBgm
lsFs9w6tapAfn5jPWGOkGe/p+wQ8nGFYTjFFRVAurSHihlOn0IKRKPNTjO70Co9w5xLHmF+PfO/n
Wvz0itmneqUxWCz2GJoAXZBzoSF0nCyjfiIzpF9ojYOcJXHCZRhvnLKNzI+WkgvMt81VhDXn1d/W
d30RQ1wDv46E8wL6INwF86uzhbf0elU5V2V4XTGiE2qMc4sEdWchn53zaIg0bsDbZ9Ckf5OB0p4S
H1Op9DQCsQiTce/134zG6eC+saN9hnFBdcpvqOghZp/TbmoW6krvzk+oEh7Qo1gYU/tzWL9vFadC
2QI/t/MwFPbSRlgtMrZAv7Qx9afcoTNcv1hfiLY8ufteY6Aa8gNdQwygJILAzu3RWTlQEke2Udh7
53vFWnmgIpM3l0/a3an5ON5Ek96rgmZvqqDubwiZxLPWz1u3uKadgcfVuwZBcvt1FsU6JZYNqbcn
BAKB2Tu7yHsqnKXVi42p7zm3Z+lhRyajG1TSfN2df5v0RCbbDUgSqXasnLh1Z+JKJQD1dClTKcZS
FUNGPBAypPOWQ1kFl6LXGxAy3o8pxHjilPi0MQjUIQFlnsY3bAHcrLRbMcZFBqSpNYMhqgjRGuSK
dLbAf9qZfAN2IHEts3zGqxczzunmEql570R/F6R8UXKcXuRNXEKB1n9qEuUxqjpo2L/NQtwoPjwW
uvGLtdGJEocsg6WngnAK4FVR0LoogU7okPZFusLpH/x6yBhml+bgYE3GIG5GFiKtTUFWDE2P9i0O
WSLmn7B1oEknLd4XcFplum7JBcQf7ALPYiL83SDE/EPidQaLy0NYiQOdZB3iV6oi/TPr48fSKOhK
f4KKRqE2t617u8Yl4AR606XCOZX/vMuvNn8hZ39Oqfdp1MDI6mTBN1qq26VLMApsyPqxnk1Afxc/
MJJuvgc/oie+NGJPflDtjSsBk/jm02QtHkG7SUM2RzRR/jzxLZeGQkSopMiZ3M3iMvHmp+Y2dUdR
wC+IQZGHh74atAmYr4+pyS/bH36vLYGlnROFjycdxOoqyL3S72KXt07tufotPSDfMa+G1AU4+F1D
Az7CFlzijTPM91iRQZdQvhams9a0x1PMHg92oQI9rETH0036VL2qnojeyIK5HQ//vU0KXOPWnt4E
wrFWdOCVuRlNHn5kEOSgaBCJVAYTTzGXcoRuQgFlcJrx+tT56dW8knMnbptiehUTzlCc0Y7QhCaR
67fwLh8gj7hJsFBwMA8H4fUIgYYQf7w3st9S+lTIOjaoiFHaey7W3jbiesYpWsaPL7hWDnVSnKe0
eUwBC3HOvM3QrEUK0G71PIjYyH3+mIpd4BFeyJQmxg7eqrvPZSrVhKgnU/Aza/3nmgt1LC0q0vEu
zTaRdxvpXnqagjSL6B5E+DHErokvB0ZdqjaIBm4Ihu074EmfgeF5j456aqbiMkZHElRL4N/CudGY
M3i0K/FE4KMBxz3QSVHw49Q8es37rFsN8gDG9hTjOVjN2QF5s6SKrHIa9eut9OMwBiBdepwMKS5J
RIHnXPAdtMn99SSEFnags1V7i2fgKmHh4h+WSRMJ3A63bRf7mN/0eJdvN0F1KAbG3STYPxVt+o/z
eVByjZoqrxmbyjUiGDhUdgWQC5IoRl0LScCutK5cTOCOebMThtQEUFR9+wWFzgtVfEfQIhOrKGW7
Cwa4Ng5LcNUFiw8Lxh5NkyKAbFstBhu0GiS6BCw95EK3WwuOLkpVaCnx5xl0FAopLokLSGO0jgFD
eAeIZUj6J63ReW6+LshPTYeA5VejwtD+1Vn0Km1jWejkV9aKjT3XPlLexbs6igQCrXFnc4mhBCEJ
sXgJm41gU5mLj5okki6Y3LHMUlBmIBSX32tycuTau9usRHbreaEbNQnqvtLSlJ2Ns0Z0mRk71n5u
K8RrNU2a1e1ljlurw/IGvZ2tZbdl4Libd7D37+pF6k3RH6cnQMO05KQU5Uv6j1Vbm/fi626IQ+Ud
92fR+4YHDLOhyTkIGCOZkWtrVO5uQm0tGmDaC2yq13Brbz8ifPSNUJZZ+qhstZrHXT2D7DwPL+1q
hOILfo5APAOHFteSnwwO3Pq58Y0n7jh3LQqiXvEsJ6KKyLWYVWzcgRRvt0WjFfq6qmXMlG3hz38F
NpSSVHoldSDRTU5v0UjUmnLttbsyyy20oxXP8CkUsBPDy0mjbJHTtFl9lZX5hztYGbbNKxbMDR72
xLSAzeaQ3rDPuEUgNG4R/pLQN8Sh7kMyBnTwy+gWQDPTjyg+yIp3wILopxTITHsesdv1a55JS7od
42aXqwyvOzj5UGTLXpwcGo7H0K6FDEwPv4fOdwIz5xSHJIgYZ0uzJTTSzrtkNQM34e234S8a4hcc
6nPDMHzZsCD2EHo26epmePKsQ2E7JmhvGl5J0ldb22z3kLlQdEtE72i/5i16q2FCggRbdGYTf8C6
/EHOk6rx3i3WwxmzpGt6DshXlks8KpwjuVvS0W95dkY5RhzsKW23YyNSvtWdeabNRJWW7SdqyKL6
LxHo9cJR33RStqzfhKVSgfEwnlu5V3IaNL2S0DVg+bFz8238gmm1t7wJd/iQ8q1s+gALp4qaS534
DgibhIN4PPteLncEtgsMvRCHHS96nHYcl+bw9ZLoNAScawmQuY7vYD+1oBnaFjngQKAfW+dOWWyv
jCxLwV47fMan4iD6V+lNEN/9n+O9fhjkmjyxvscGWYUzPuU+CPaKwWJNoBnfm4osk5pGowy8hD9l
d4GbfcCXmNx8YkSKIRRY6Acv1RZFJq+6k1TNTz0+RYsMBdjJWDcbtge87hG1fcSrHqwLommtiD9v
4/gXqjK/YBRUhfjgqGH5EMiSqzhyUpODSypW7jxBY/6WXRtyRbQ5fa2xf7Xg/XLmiF43KINmZrtB
v9GgmKtpD219UEeNV7/X8pZfOHipk0a2sNWtGQSoX3C7t1sojS7wlbrL2EsQRSQwjZ5lm3dDcv0b
G7JwsL3K5s9MY143S46/dUB7WI8SlzbK4PH8T8OCXaSvpLr5mvzHzyU/MOd8N/0NAWdwRo+Jd2o7
8x+Rm3ufv9SqEf3Oiwxmntk1XL0TnurnqY1pklfK5FOyABjAnnJU4J8XNTIpWS/o8wqRc+Fc27wq
gJiK9ebKQtGqzjJ3V6yham7dje/AihbMGcnWjRQT7hnlD4IkSWSbSnEr6IX5C4Jaskz4e8Z2AF4Y
xD5pXoHVmvuYSMpggkAJ6FlCW1TAOjZdDqVH8cl63iaZmm/gP3KhU4JQpfURpcqHOJqlJa/NFum9
rgaQQ/Pi1RO2kKHUoXaoo7OpAssU37iVz3NRm2BIti6yo/7EOw/B5i72xJEg4erAijgXzl+Y6KHC
EOc8y8N7va1vNnE4HXCZtSyPk+1k0Y1HeF0AhSbCEn5c31pRoYSO02E0fpIuxWP8KDMzGzyF2R0c
uDYlh8p6ME7HupjA7cCbS3e6O5O+zwAcVXucbsW2Y9YR7zEgA/m84EQsBvjC3ygISUfli+d0jSHO
Ds9897C/cfeY4F9YGo8ydVNYS9bV4AfVBYt9OZJv16kE0Im1qh+IpSTfvxD/jjSqsfY4PyqcOjd5
gtpwHBi9O34+n2eV267ssZEqtpFJKgI+2qgkHZwMHH5JSvlLD7QYX5jsmKy6v+Pb94KK2HjHak/c
5Hb62u7PS5G3XWZ4GfcklL26zZH8PHg9Tdy75verTO1t7SlAMkArOWMXKpGwqBoqzMMwbTYXOLQZ
E4KEunZRQcOAxw1UkAgedxZjGnYP01O2C180mxk9O3J/itEfLvfKWmRON5wuUUf5O7zMkyugSXeF
AiZCehUK6m0c1JFTHUQykpOrUolmmzXnRBV+Y3+cB8u2pUnCJw9I7DKrgnPo4JHA+N4dvsO+Uofz
sWI7AlJZcGov/S4KO8nwv8XzF1nW+wYtpAdcnJkr1EC46rRrDV1yUGlJ1FulN+KF5X2Luka7cA0X
cS9Q3bCbE6MnuLXEtOjuxcAiBOPg3m5OU+WPweHrLPz/LhZgrp661/SmI/fhCxB7NvtRGnnHx63G
q48Xrt+EnPi+LO32ZXmerwhoYpXx/lnYACUlTlcJ3e/p57Fb6PBJWREUNJwxeLV4W3Ms3/c4Frr6
WGcrb1lswXTIWYVqyDx0i7RrxHG2dLSQUbASA6TnJBChT+GIZ1d5vTu/PzSgLTMkmmhA7gCGIlgX
nqaB0+yNi5t4zLGQzQJG9kkXaPvCAtwLoNgjBog7TlJ+UM1ehkdZQCIajg4wuN27JzSaeRwCjcnA
pkbC84N1WvI50v+HiRk24zLonfu9PVZ7EYVhJtKbKVUBc/tSKfdGLHDPvZPp2feWCRkpkk16HmmR
N5po4DpPddV4SIhyBjwCC/RPQ3MpwvoBAsbIArAxhs4G+F8D+IkBgUOQbWWFNPNJl6fNKv/hViJU
TuNEOvu+g8hoeEFRxya4hRdgRFnDrjjqeoOFu21phAcrwnH/P1iW3QaTPcRP1fim4EcSubYQfUse
2Mb1qq23CWsKccXdNyRQwA1IwWM0matF0aoQnEOpWnBmgdIjlKSMQkGSuvrOTd85W6DqVPbH9XW2
nOLs4YC0wnc1hbi8JxmWZk0TPOHpEl+TizHBbtalOTZWjhnYiLmHatQUQvXV936KZA76u8vCMfm7
CI61RamIQSpz7K25nxTFNDAWrZdic9TmjL1kcjyQvlcwyW2kDAG8I7eJWYLA01yk5oZ/bD1hM2du
OTNYBMhLQ2IfOvSLTEbTiTS2RtQAhlTU3spPJX2QVQzqZlkPueIWVwRtmMbG/bdvvinMNQ+UUc7s
UmKGR70qEud2G4kERPM3cFWKDeu7u9Yl634DqKWJY5s2T940yCZqaMa0G1LStwnAqZ8fUmoLv1af
fXE/jU6ihT2O6JdreSOghizxFl7G0yOzIJb78IuO/SAK8rRr04hpUqGLD6OrNuArBIyqQp453uPg
6fTou6FJqkHAPo05cF2KWNh5xg21xEVrowMPDAZlV+YJZPlf61AhfO6LXgalMw6TyT/2wS275CGL
DRtT0/VRzef8HG/9Sb2d1/o5yd7OTVAhF2umX9x13aTtvM6TcR1MeIrLHFFAyI/Mjn1/cNqcIFhU
10xR/iPtHxdRprQ1ZviCqJs45fVJRlCNtbcHf//tCx1veMtAjQ++Zz3F+SLeCLR1wc81k7wb9Yj1
CYMCCINUpnwGFaLgBetzAa0wcDslz28DByg2GUnn0TaV38+Z9BZU0wSek/+zP/wA8EoXSNMO40vw
Y17fQSq0yVmSot/RCQL2O1nZ9EXUmiZJ0zLsr3iQsJkCL2TV1lF+hJ0w4NGiTwsamVHuryE7YKEd
Et4SsuxdAm3nIHnFiR0Z4Lo7TbXnk6D8+eHsUXh+2AXgb62wFZ6U7GshRD39PZ38TErrFPnY4XO2
fnrvCnJ83jKWDXGd5xczB4veBgJ5WQJvhxKtP592BDykndIo7h3FKa91Wui+rsJeI0/Kh0svOhCw
luURablHquC2Hpjnd3uPczs03vU+Xcpq8dd+lCwA6YZzPQyybePFBo5eUQmmeuhHzbF2wr+hMmDx
NAN6I74ZfrCu/vxH9z5GRR1PNjlaTvtFkj/KiyFVFanMKvxoztmBEcl1z63+lDTTsPk/lLLCSy/V
chKWYqW+5uWc4A8KlXRmeEes9tLmmBz19IA5e5/idMTUwKOPeOqKxPaRb34knBohavAiMxuPCHMa
CW+F2dTNpGKEDjbhyDnPSf4uSwwQoFdd22xUExUTK4rJLGsmymvFlRWKghNEP2SaXzezdyl3yO7n
wBjxjuim1+fLFS4KIJKJeAYY41uaGI0pqpUkzMlL5d4vKiTcz65vA6Dhirmnv38RLjbuaqeQuSZR
CgCB08Tn2nIJ0oR9s1inMMzlNeLo0IxuLj1YfRZwZwJ9ZzXfIo8nnoAFXYYZK+KWiumBm4f9/dGr
RaYb5lDgNfJyJ+u2KQuq0FTeYhqTgDWX8j7JfE2ildPIlZy77yqNhsxMPS81021nZkBUSGkwBCGN
RAShCUjC6dN5ChKsOwNRFYiwh5eB5cSgzSIDvrogoeq3ANomunE5uz9dWK99X94l/COngGvlrKvT
eUADR+yCXCKV0JyDebrtWoHxYScNdnve2/ebHCqyRYxXKZJ9ZXJZEETpa8LkoPqxsYiPIuNp+/vD
n1CkJxAVypqjThA8QBOKdfl9AWtiyMoW7DL6qh7KTAgNiaqDSWevDjKd3PdrlR1JQq9XqTFhAPQZ
z92InIgqkQV2k5RfWEbX77uL92j80Co3nqUTLpZ2LpuLXjrfdhtcEYBcKvjfYJuuETHar3riwhaT
0snA59t5mrgbGX97/iSLM4Ls+o35uItfGZJ15WWeW6i1gAtdeaMzYs+8yMw6ASlCv3t6QIjWwry0
e7g9tqHEoZeZ0cNGkj+yRMEk0pDlPe1VNBEpSpIj8TPuOyQfUcwoaoeHNCxqpn32Vs7aHPU4Z1GX
R7gzQjEpmm3y4xJJ8ZaPhsqRNYzBL7VnDTluDwzAR0b+S3k4mHa29bCqiFRCV1IC7NZStjfkAd4d
8B3+VFb0WD19seTjPzMrzEWFCQj7Iorvf+oRstu8yCQqER1aepAriCwVTXdaoa/BCizw8Ev+midV
boS4c1ebUXl6tCtRoBdk5EMpKCGM9f93n1dM7/mgBn1/F3TDUb1WmF7rkmZdaT3jOpZgKRuKOPv6
dDQdknlW4+UxjyiB1sFhkkbHesXAUnpKV1SvhLTwXfDzQdd9GekAkoryWcJA8jp6Zk1PXVNyTwwP
oeEnEcibmqPUmFF5rvTrSCx72z2ShIqWfVV5m/TaHus+eOXL+gjEU5Uv8BDejeUHA96oUUnnUFEM
NE00+rqBbYUIParE2dcDiX/vdRx2MO5AoR8ClAhO+zXCIznf1jx/Cwj+GYQb8y83kEJ7lJyMt97h
WbyH8+fDg2Rd0jhyGkyBjLljhYUsnt1Wp4Xp/wt2cprEVbZyEs7Dco5BLduOInhr8vPeQtoXow1F
dFRDmRPKNnMW781mnkMp6U3CZ2W4VUjDyeLaTcdDlrSwSGqxYvOVcvDtNj/P9LvOkEOio05ak36r
geGfZKFJ+8iwTfAMAQkvFZ/dpZ8bDKWcKxMY7IkQb31fNmhco7/ZMutnsZgkuhC+hr2ICG5BFXWO
BYgvnEpAADEy8LSMI4vmOH8frMRaIHPyQx2x3vqUKssvL1on9tOkG1Xte+yAYls+k4WHKQuadfxR
07mHJ86NcsH9xQXGzd1GunZi2OyPmYiekTaaAvmhlWejRstFcYsVN33xo/M45Lt0ZfgOD4p6egRK
+5xWq3OJWtiP23Hq1pou9uOjfvXnsU7ilmhPALp52zHy1qVLb6kDjLN+mq4HA10m9wxX1QYChSrV
Rypo4KhWXogRk39Wim5/NP9d4hBYA9WSSwzcDtngOjKlneIcM1mMbFC+E2EnGd40yucK0eq6EqDZ
tXwpdh3lY1MvQ4SOPiqjYrytfxQEy+noLnHYc5+baQEIpHS9J1Lh0hMBKZCzDaxpQ5giVdNZLHXs
MANETwF2ZwkEfdSd1Qhc+/oRh12bbNXnKCwp4bCxIlmvAKddlWtzGDFQnrlPPiZ5xliYvGpFtybf
Bm9uM2k56OLlzlPO+EUXo2sCGZ6w+LIIPpJ94FTwpDzqKM9eqxIIrrJZxZznz7xrrTJ7c1dGc+4p
ND8p2eWcRY3ccs8FIXBkQk8Kpjt8sNiS8ItbR6USk6TrgPmFXxOeD3jWKQxZYzdwn/wj7pMzQX39
U55F55X6KS4yLMwLWRvORWgzZBXtiKV1jXyhbq0lhqgPFttj6izVpdUYHms77tLKy6UgYDN/5PEm
W3sWLcdo9GjQv+9Twqxz/qGQnWHE+lKQFbWB6U2hAYxY/gjeHJfwwxMVTVc6C3ETgV1YFpre+xv0
OBVnVAlJpSDQVOTnvCzS8GRYjYkmuBr1SGnkSP0+DGAybaH23Mnwhj/HMMu+uk1C40UzRaAB1E9q
vemnyS9qWFrYVNMLYgZNDAD8i0a7nyouotWXQojdREt+Ud9137/Z92Iajio3sU04NdlX5ZJqLQnf
ApPGsZuYIPiLob1oFNXeXRGq1xLYloTSutZVGJGidCqMFr2AFU+6mGbL/iCimTkeySbunxvT0UoS
JVFguhM3uxi6V1jb19unbg0rrQPERLIrTcEyOT3ehLSH8qO4iryDsPqlJAEM+DNAqK6idua9Fs4b
MqLgFTMZo9FF19b6654lZtxzIQ8YvPWWyaChMklJ6TPtzKzz1PO2CAdt54A3pGXkaXreMiP+ih+H
hiuqf4lw/sUrvqlcnFMvcK//IP3G5F32d2i0RR7t4ICoy0pmfSbhYD15D2VLIVP1aNfFL5qneXzZ
4o3hIcA6CQb28oYVyB73345+IYIxawm9TI2EVG4DC0ejDkZOuVp6xx3MYK9FPULKlPssnAVZtOy9
xTwgAd/DJyTo89kRkiWIXSHuHFMzGNTiSGrdLzoA2ttiqNnHqV3NowkpksCEJQRZzKAEjU5KunvI
yPBoMLTJtRH8aiAzUipF+qU1eMPvUmL1HEsECudrKSslXGBGUqA8pCKB6enQLF5aiBuuj9b1VOaF
ntwbXJStUZUCrdI4a23nMM7SOsGnLtUKZjWV9dlMl4RojHSnXXZQpL2fqu7+tXFKMwmg/nRn1Yfe
IifXJzmMifTsyEwxWHFuoJktshh1pLlJzunf52L4vd2Ofo63GHLo2qba56iigUF5IILS1HzKg0T6
GPNfq6h8v2Ig18N0KTSsyIRYV2rrAgkXOH4O2CKpAIldbSPjl5QOo5Rf2cXhT7W+bB00kHTxLBUv
aVW1yv3XRm2EnQqFR/HI/0m6JfakcMrp+8Rms2tJQzfSIXD+m4Z5CI6TgZ116BN2BISc77MmyZu/
dS3jdnxrkpSAmLn/g1eUECd2JQmZ9F+7wLIpTIB7cPtB4hNmOLSivLJgpQFpWppDQ1OD7kiB2Kwz
sgjLGIUxzqpmOfp9vuurmSt6BKX3L88ZVKyv5fmpmy5qNhWpXqrBlQ0oCk0aONaq4MIFvpK+C1uD
1Ksbum7ja53MIK2Huff+wna8HkPIwvEmDdYhKk01kBY44nYUbUBF+nEyMnpVjUbi9hjcR1WGP3OV
Lq0zROHXD0oZFx2c89zBWrl8xxtdMNajbYR1Lcm87DNqI8keNTSjw1CW8iP3nF7Ih4adlGmZgx9c
CJOd4DRaUHCtPuMkA6lDSOE7L+nhtAzg3449ude1n3qd2MM9PJ8rZMgwb+FoTKsJaPRDZkA5Oryf
3l7d85cPYYB81XhVsSP13zKNhv4s7QxMBNVThC1ftgd06YD5DM/vbZDgrV0MMA3QD20s+MSo8GYr
iZsECJqzt7np7YpnYS2VvubKJOFnYcb4u1WExPzVishG3s+0012x9dzAvvKmCItjewqH2El1iw4j
8MjLplcr0Xl1idygQDZ82CAeGprlRgOCkCuHRFd9UhdSaZ15HLyhIkhqXFjAXgdG0sp9N9XN7iaX
sm8eg5uGLFNgmhsVnBpzIsq0+Ov6iiX4vMPSvm2nu30LmhOGsTrV2P/KZSh4It3ywTRNmrUvcBOy
hdpd9IwbBEBdZ5VwKhf+y5dPS5N0EMSNlikl0WKXqW+lXhiVjxgDWQKg8RSnFW8QabI0ms/Weq7D
aGOObWNk+Fc6gfPo2DCA/umN/Wz7hSywfyE4ABxebjcg+EWEI78L4DwE+gvZx7Pd/xNkKB0tlDaM
bC+4PdchAXKj98zZWRJCy+aloUN/XVHaipXT9tM3uCBm/SGAX38pAF4RrhjZpLJPj+25ovOoQtyv
dMfnre1cxFbdnVRBlt332bhN1FR7QjD+zpgUgKwZ2jHaMWXt+GJx9vlsQOiMqypzKeyS4OBPHQGJ
VNQRanwK9FUZibAJkBQXUzlatCl4dg0pQa3PL1Nzss/43Zd8s05RU3Bjn85Bd6hCIseji5AVn4H1
k/OlcjGpDQjb2PFxePpt0cNfZJFs3lyI9/h54qqWD/lD/cx52zPM00ozYCOVOeUuyZp/ZTHD2nTt
ChKB4CibRHHCCFQh073Wr3kaTUMPgxFrptLB2kkRmCEp8yDhm2HkAUWdocS0h+BbUFD1aMHHZzVJ
lwfynt63N3f+6i9Eg2nuoSN0SiP3GWdp6GH7WSHBgb88DyLX9BaXT6uulCvShze0yHkHJbPQN3er
idm6bGnS0uZnwOIgHR8Uol+u1XGtO2c17lDNL1pegdQZ2YU6b0Sts0ueEu+zCHMBMr0TEIJLpkFy
TyHpIfMbJYSGMaS3gris7NmAn5xB+kkXAtMMLBx6b7h+WwY+hfMvb5K1/FesXkI1m9M4VMO8r54u
bmuUszA2w1m96pMzg0rAK8IsZtUwvj7Ad+ns74ghKbz3ENGiYkXwqfNVIZ4E3+1Yx/cLn9casK9G
9IHrRa1JMtS/zyVT1ut3MOU2+8fbkcu19Q/T/nIZzCzkyHGakMBc2KaS9byUK0xqX/UdN+Rqg6KU
uQo/tjdH4mhlirYDVa9oEjZkRP4zXw5TYiJw7poxTb8DPut1aPz7v7My+LWVYxO8A8yACXMEwZGU
kd7UQ2mUJCvlfIdzqK787LrRvmaAdhGuOYopJWIWDN9LAalT1a7xWk/H5for19DUNzUxtykq1bJK
1h89L47zOA0x8sEMhyQaPfs0GljpASjBe/3X9h24Bqd7tQeasG+0UwUYuCUsvmP1liZhoYw3Phkj
po/GqFdSKf6cCgvnJ/O4OPCPiHh/EjnTRD98d9xoNYBIQxlOWvKqgQEC6ma7qJ9xkLmhKW+ZblNK
wphIZlQfbVypAQYzNElyOfn6H45wBvGO+jXGkpiCpmYbg0cC6dVUzUu6WHK3MGP8j/8jdewBeiHv
3oa9nu8AcT7wSeaOAPx3FDKx7j8L/1yvaIrfNuNF6Ba8/Q0JbPpnOus4V0Y2Lh9j69GlebjTqpFE
RW7K6JmHDLFah5DDVrfDHnAYlc1e1GIt+U4JGkA/KNAmstVuqfymWjGiXdXzE/3sb/ux6ld5EAXv
SIvG4i8BlXqOh1VRLZBVRKkigVvYvbH6Mwf9RqPKo+r1ujtI4+chNU/zj1z1JAhe8GezPp7SWsX3
EDtrTZ9UBFpYfkPXxXVJJtVDZ/SttSYbKoOIj7kesCw5Mdy79GdQ+200l5hWnNW+7+6fAKtPPkiD
jQL/h0K6qtV0/MQ7zZmbp4L6d0fAylhPAoTvPLZ31+Z9/TynMA5M5xE4frDDruBgDuZX/sM81Vip
+AgH6wMkJVTEB3BJbt90LraUYI4V75T/J4CKf+KMUzBzJL3Em4s339zOKkzVDAIZmVGyuVh3t/Ji
Mr39hmqZgNGlEYBMFIsY/9tv6IK4oiBR7vSlz4iHVTPFzwbqzeTJz+4l6F1BFW9+qtzzrDEWWU9u
RniUSZPzYdp2jXTPPFb4B2cunHojG+ziORVBx77yRSkcz1ESfnwxjbsAhvfagM+9YOD+tDkODACa
4E14NekXOKAkaZ5YplS7kDbscGlsKxz/ePaqYDZGyBvL4/jjkmvvz5Trh8vEBht5Qa5w1LLQnlwB
dJ+2CnJ4j1Og6Sdcf2qKZ9SM5VHsjLKcI2PB5AI4zQl31K/OUY3hjvvCsIPt6OWV+O+pwH4+zusb
wdtDL5WVyEcw+1bOVjSY1Omw1R4TUZM0HimoJ2oava9y4pQxuZQ1OOeoGafGUk9WJyN45dckabBd
uFWcCnWZmRgQMEc/8lr+DqR6J3Dj8Ma8PJQ/pycz5ze/fXvOwPVnYmjaUQ2HMaPqaIXDvYDnZWNe
8wDDKznSMTrX2lC1QhIx8c7MmwRb0IcVDjVmZI8exQofMHI0ja3WdENTWPHIw+lwYUzNn3dnOc31
1lZqZjZwu9ld5GLXamFizIHylZthPKdvd86+3JtNdNgnz0llUQUXPja9m/pQV3KKgCZR4rK4OOCH
2w5oC5OtIm5Q4omSmNzvpizf00Fcu73PZMp+rNt4GImu1cmjioyCP9EuCk3pidB9+Dd3XfGRMQVR
l38+i37sQqBSRVqulB7z7p/POz1w3SOiQVJ23I8S/ISGjQdU9V3vwlJUSzwA1zD2c0pegijQ8sU4
P5TnxgyVfCnDJiHjM3bjrpP1Lspg1QH86wSe7vuwCXNq9fddEbdGQDFFWSe76r8i647k1RYXg3ib
PqRGhzI74Pp11NQo10Kb44MCsKb6h86TcvYg/3rc/Nl4gUaNddKP1VM44RF0oIN2IntCxkV1jIF9
jp3PuMIn2GZSXnnKQ6izB2feeqDNJFvOivjjT+XSczbbcUJBLt/PaUNYvDt0VTme+yzNLUat4VhU
NeTPtRltkfbvhy3MyFw8M6zBV1oXtKTc3ZARv/YCW6n5R0XeiB1NgbG6h16Qw7pleKICgpKRhUuD
/i0Bs5aBaQt8ZSEJmVaYz9Lz5JO9spctMocKJQ4Nz6D+Qwh4wumtUkv8ShZYHHWyMViOuU+UKYkV
2ShYDI7hrDjXYBqgsQN/QJdjurHuhKzxkfEHGFdAvwu4WPbSHTjv90Dhk2yYjj8TdFLPQ2tUHrO/
XCZo5L/MjV+iGNx7GHb4tq2whuxEWZ7Wsqmfl2KRYTAe0zsHklzerSi/F+yNF/Ig/og98leeR/gA
/JKI26sZpHERon12YehIfMLkeGTjQffiyQORCJ0ztdT0pKSLBM+cGaFEjPra+QGP557N+qK27O5X
lylf8O9z1pZT6Luq7ZSY2v1QPtFus76VtnVbQwJXkngFA4M13AcoR2E2GgmDp/jlu1+NqDgN5oPo
wDOUVi3ObXhjCyVQzUPK+8SM6Y+zw+3HHDL+htHlJkUzWFWvncSV8mw9x17Q/3NEg3JZaLgQZBi+
ZET4kxzgnqIix6LnMlw9VHxGcYUfiH6WEgrsby7rYWqt0Yp+XFt4uA6QRGzpq36hGS31QC6NUDuL
zz5QxnogJuAZrOwRFxYmYAaZoRCsJ8q4qPUNJBLDaTSbdqDzxTyaZ3WInEYoeGlyHyeTrU+mQrYY
xi6Eiz2DkyPeyoD0NOPwoPEoTVPgAmgIj48QKkQcaeuxCd3j7dEjO0LBXc0px0B9/PoxX8s7xs2G
UIKsp1IGs+zNOixQg0v2n8Dln8JgU4cpJj9TIAZqU/rd36xkH7GPVbjl7kOvTYonBIf9fsvzgltA
BI8OQXdFI/sMiB9RTHojgb710AXTwTbvnHd/U50Uxrb8LSA3R4nPXVXvagRr73MvAYJ5d/NPrIZJ
sKA+i22sbHdqDpjiXRJW86iKeZRqkhdzWVb5eCrI36W4VMPEJRyyFnrnMJxxMOIQu0a8EWVGl64x
C1781yzM9p5/8SVOaifWzRO/gxJRgvzalezRjEnmkcn6HTQnjdNRMP72nhMGChxd1ICSMiedgE5q
weggWb8+AQ81V0KfxrFsbSrtS6/iT9hCJFZ6o+eA/XELrhR22dI/QInNllTB1atRQT9zL9VpkQ+e
gm6I9OB0tr8FkMAi2e+GnQpV/f2THhkDEDYK/jnPaXQVteE8GD6KENJ74XDcnt3HD0cw5wjpg37O
LfhL4W5lWVQ9LgzUJ7LvX9Kwocrfa+TdozkMRts8HK2NKqeuSKnYO+XvgF6yRa8zIIlfW0Mj0Zvz
bdMotC4UqbSy4+W9N8dENbWGSlusc+FXrYkxBZIsA6/Q+6Wcpa8DXK7zWUjsPLfasbwrTpm45SNW
/U0ydQ7/hw8lzx+a5ZLbKJWjmPjBtdJN5djlKYuRmMVNxJVC9KzO7P4YdGoTY/GDd/fqMxitIc5x
4QudFLUjTnsk6S2ObuiAz8RKqKXX7vdlhAB8LhpS1swXfM7CP1aOovScxBbbF+W4gYOSHAkuEcI1
F161z6e/l76/BEIm9QJ8qCNSpUuFN21jFVB+KsOFhPsARAxszfE5HSmxGmBBNDoIgpiLm24M6VvY
sJD6GMViuG4YZc0kuXUVvQYZFFGGM8IHMXVv946AkN9IqOMRgdjCX7KVMdmohqpSJM1iTCYwD6n7
X57mY31E1tl57IN1Eo6STKr/NmhcSbnXvSXBd7dUwgfASKj5XhagWoLbG/9aeyeOVxYz5T1VO0AR
czyRPoq39H4aLE0oMr/kx9KkfEfXmN/pdWqwHXmePCK85jaJA/9KWWyIUpt9+H+RqGkdCXAwWH9T
Vef0o5cLXnVKaO09ITTmb/IeMI2jc5UzZ3WOT+P5igTLlQcp/Pk4mSiil7hHiHsixORYRAfrsMj/
7P3b+6Qm1/99dKUYgzY1gU8WPoeAnzGfOfIh00pxhjPtwXQTvPa5ERVLPhL/lOZdoKtgdCQtWwTE
PaVh6IuRxsyiJnHHDdHC8fP01uIQykhLxSto/lipk3pvPh9FBaYKzAFukGwLhkWs1pF7y+RYUn0j
6QiOAeCWNInG4m2p9HKvdZoluSiUmLIZpG2cRXlaF3oZqD3jo+ip6/QracY5bua1cV0FrTSwgshB
VaUKB0L1pRz7mSaGKUKUESxDtnFosWFdGeLgvSaapTmpKjjslb5mNsdCHJoYoSzjS6z9ZHcBiBlP
ZbAnex6/5/tEslb7rBtL4XR8CitZFfLUUftCt+32V//M95CyI9WRSgYlJVlGLR7jMIZlB1laacw4
ufqmYIOSGP1aWuYHPENOxb3jydctUzkgCloPt11bZvcsKYiZRNBDOdsQHdXazaCDXVj/TteQVHPo
LDzDN8DbXOph3wvSDA3C2rR7ublRFUic1nYdXZlVKAm7ob+pIj1UZ+S2pLlN8qEMIJeHxN4V3soM
YeWuRL2RW8qOSvGGzpB2ybPNXSIQuJoK7MzWWoe6iC6bTQwUB/Q2xrjo3xKNzCB2Emr67c7kb7KM
tvS91nX5PZzR9xhMH98KZLe7Ikc1qepg1ZKKD4e2iqzbIBvpH3MSq7BmmTY94q346Wof+s9p2ZfP
3hInTK7ejtIXsDbX05XHjrdpAhZGJ6veCPKVBV55eS+d5peh0adomoFuBbJ0bTfuNag1E/tWbk4c
znSrSWcwYNQqNATA3s+F9c2enTrkRzsRCNDtjyAiPSYgoOk+R8KxHVvd4jiHwAvH7oN1tgC62LEH
0APyG5ige2I5W2nwHn/QpXXmku3I6ia1xF5T6jZb58Jmmmdryzv18vwV5Lh++hP2QetT8XMCbCru
YZF7C7BmR5WX7KywZnrMG/+7r9TWyZLOiSphpIRpUPFDRxI6QNJJIXxnAXoBRbP8oeXpQXH8yiRv
5fP/M+aFNVG2x4lXe3w+3/Uw3gfmEMeMxUrDY48GqiVTyWGBieDhhXyVPcLwulfWMbc0oBajXKum
AWVPJT55ruTnlVXNuU3jkqweMcoyaJMZ85rbyBrxWR22ZHWCXFK7qkovEImlNOS6IuSSJKdE95A3
13eXtzqEYFG7XgVLnNlOyr/lhOUflbd/KXE+4fzz4TrQwejCPT34qjFlPm3r2Pe3qQMQhZngbUTz
Br2uaSbooK/k/fGmF8R8ou25Xk3+XLx33BzuY6b/MApIypM5xdwtd3rxiSlvE2zn3c1a2eNOuZBm
XXqAtW6qkvmlv/MdfjFUqQuz1CO6XhK3bZ7E0t8AW+U/OGyJ0yjGyQaG+P+qUki9tdZ/eNCKDit4
JFDrppfz+0HNSiEWZAujliTM54yyDypkairDC/D0EqHKfk+2F6wbvyYdUm06Z/qTld14+rqG5Vyj
b251U41eC9xbLW+hk/GWq+NUUEvpvvOMJ1etbOWAA5Z0z0Zl5KRIkJLoR5UVywKQx2/gqNQojWqQ
ODLPQaj1hA9yKhLjSB78T2qahWpQG6xNcV3vwTkMhXYhU6f++cWJaeDM4egD0fhPnMngJUZqFEiP
itcNwjwUATX5elVREhjkFCPQbgo4pgk7TAm33zS5U1VW5kDGFtcK3EktY4jnpzD9Yip0gOGo3gWI
BXdQ8jGR4NgoBnJhIoYxPBQ795u/+6LO/P4VW2eByeQTea0MHo+pWML445rGXKXzQXp+e0Py4QMO
az/NBehD1idtfaPpAsEaucs10AOdN8JDvb6TQgNPQFwfx3IwXce1k/aZF2aA8CDXunf6ss02T4HC
NsRjsY5YTNfk9WLagZ8GqQAEe7mYaF46IoI1HPFqjJ1Ncs/uw7IATT3QEMEXJajwItmDbLZlnrbR
et5xeX9ztc1Oo7YzbnodGt7omw7eidozZFS2GRostQSecP8i5IPzQvljN8ChGMYbv3en19hDfO7Y
HOGJ5WsMYheWypR8Rfl/8xUbzYRSl+wWKPXbTVgWCbXrBPr8FRkwxJwfvMkTINt0Sd3WRw83LkE8
uK0BY7HvyfIsArv5JQC98mR0ozkB40iyEvg/y0oQBTqB+ZofZ1pyceYAJ1bSzqEkM0aYPxlkCYVU
KjE4ghoWqTlCHGQbl5IQ6s8TTLP14Z4kRRSV6bwjKiBBB+JLEKrQ8LLUNnfk2zYsyQjXq/sME4i2
whNiCdmJw5z5V12np/iNM7fNzreB0/KEoGOTvy/QDj80JMbj7gdNIS/r90Tn4L//ORLF8EVGLbTa
/uiHP68lhLPy3jU9QSNiiXs9ssMaWxVBhNF805I+gxEcP0OWXD+p1LwlG5vVJuUmM5+rgEOkjwdW
ek8lAipiYubtxAygnERWNPvkD22R+FRZZAsBRQ41mL0J8KR8uFpEgFT/7folvuTpaRqf3DHm9RYI
wreMo8gGM1PwPNsy2O7ubOIdgxF+9BeTxS4cgb4G66c9drpJYtNkpTRePYPbi2QncVv0jUyirtY/
xGHOKH2h79lcyzWmIG75Ags91BLxyFTb0WQnXfroQHCGP3ZJDSamzRDuRc4g1Q3212p39+QecmE1
V4MjgqIt55FaS4hu5QMltEUxMl7w1LoE1WpaA0PuzOuo6aQY3053Nr+MEOpjBHjA6h9SrB2LFI0L
VD8rLq4hV89VxgqpKy4S1nzyVhBe0L3ZNy+hHZVeDB6/Wv2u0Byda/IzhD4W7GsopbcPb75xX+pM
/ZFPlYsYyiuMPgEwmJCVeyKz+zylbgjRF3MvmwuzCpUE2C2xvzhfVFr1Jn7/DjTL6ZXo93okNt4R
VjsdJfmlE/jutU9LnZ7DX87Jy6XiAFgvyLOReE2esZAIC4nxIGAs5wF+/+/ueuvv196NASFlcXVg
BMBLKVM1w5NnkW9C6ibYpSEham+qrZjvCaTs9zILXKoAl7NKSM623+3pBFIlAMz9gBNNiwejakMf
lMgFvmIMVxdgCCzgokfQ19ORpxCK2ms6egQV/v/IUI8R+J99zATKovWOqLuk8a3TSQIfKAXvZTD3
TilkRXHsU+EnU99DtCVks3Re7dxPvVQpcECKrr9ghZtZpGeElVtTgQxCHo2q9othkwnVguOFXWCM
S6Gu1qiGmEX+Ty+I2+imT2k1O3WNCFf3fiEMxkQ13zziwyD3BO1PkgXucqJigzmHi5bEVaU02Ar7
JTbZP9FoYKCK3QnFAzcsGkVsBjHKI21ZxdtLIfFpxxBxVe38nAxQ+rmNvJjIVk9dea+3rrOMHVOc
BKy2+dVIqa9s/ybMFbofvN+058z3M7kgpaLjJWDtuHZ1rjpXcJsquT8Ai/Zf2xmJ+rsKhT6N5mxF
Zbin/tFO9dwGuOeeCsMAXjPd7f8bYXfvh0QkvO3bTllvVf0tVDr28rnaH2s15YP3UEqSEGwfMyEF
Ggcf9T2rRxNMLyrGgMQYJJV09if+/ZXvLy9fpilJCCW6HmuBTNEUrorMK11b1Ft8Dy0MBJvGKXPC
Pra9agq4A+BHRJoaB7D5LW7QP1Tol1QipBjJQjd0CCOK8IX3lSc0TC1gLqd4L55Jp/u6hqNiSFe8
mOIurTV+m6f3Nx98H3cYPXPc6onYNmOsl69iFeU/1WebFYT15Cwaz2tYcpqbcSB6J+fe5xdABkbi
M3RNgb1luQXVl//uz5RGjorZ6TJ84R5rjN1DL1Ojf8YWV0txGk8um702tO6csCZG+ktJsfDgnGgl
kOXsEh73PbkFIWPjpjFjoLu2K1iBMBrfx2ZGCKIYv5CI42vc+dOYw2qn5JHkciWFG++YIyWiV/vn
Ru8d+VxSAbT0fq3jj9nDJ/c9lDSf82J9UwuKYDIrISvgFoiol3GKxAfGDnXzpAZl8OWVULSp5q25
df4fu22D6qF7fYICUkvnvkgd0H04xlOC99bzcCafooRvELrEWQfmmXp963Way23yiOJJ+FaI4pSa
I8/sM3OgdUYGiURZHlb0pGiN2A0jeQrSrbe7qbsqN703qSPcjk6jDc1SuxNasdK16fZx4oEf9cgF
YLK34LtGGgePtX4HI2Ho3s6gmka9iQO3MKZ8ZTQH5XDKORLHmaBMhbR+X2NtHC9PejI/Y2Haitr1
LHaszwTxxaogeN82nPfJ/eKUu6jW0Qo6Ltsx1VlIcOmssrF+tCiXVmSQBmegw2dUMoiHN+nYCk0q
4NAJnFrzzmMKW1ofhkDUoWtUOrD+uL77gF73omqkP3LuH7mDf+Lw50fZ/C2sdPUEYq9rxaT4qvQZ
pyY79KrFXO6aAXObwu5wJ1vrqXEeMPTvDUFI87gIwJJh5oNVNp0AoVVb/hsbM7IokfZnHoip0x77
RMVJG01sfpol6ZaH3cr+y0GmcWfqpLp9M/mjDvrE4htb1griRvf63EMMtsKfKtTcL1lTqU3GawXF
PbikvqSum2xFpC4BO2H2+p287JfWQCWytTsMc/GI0nY3KAlQjwLIfw+fvLrvtt6gGshsqhBPPFal
UQH67/bMq1bs1G7BK09j5Eee7VY0AnLm7gE7mFyjzs1q03XZ22hweqyR+D7SENyw4hQQdY7TO/QL
w+mkvTTE/8sNNjiMlFitJ5vkvifh5hF3Mw/EEUdZgAB82mF2eG2daShYnmnmLVSCbSOUD32HCsbl
lxBXhyngPzyEYG8aBIR4AbierBwXQjQClP7FbrY7ZqnHJDdBYij2/wkkI5obtUNHChUoFVvevLxp
vLAhBzKwgZNc/wTLE8eWAPGjp4xqqgS2r7ATTdiN1B75KCpau5XDE2anuU+3mOevy+iSzxaKC6kY
ZQ7ZZ+WU+0VIqUnq7aboI59RIBAgjVckVdp67iSNuRrlOE3QobGmiv60J2/t0yctBZfiP0GduKrH
mwozDI66VQLtFM2cgYz8QmayxB90VE3WAD5XoIPcCuKlFsFNQqNKWne3R+SW5ZdIkD/dxRvhDWw7
T/AEv+ORl4JNDk7VLuWPKIG95iCdDFjyb2YszZoC0MHWAAXX3rv3Sg7QsT+MrPxUaLpnh+4uhXVo
zh/Y3RLRg47FF7z314JtwXH8iDwQ5mp24cbbZEj7Z2FUg7au17mi8NfE/l81Ma6HHWbqVBnNqeOf
2BQT4NmBzXYXaYxFy9lyWOpwYa6vvB8dxuyJbQtpNQV+SGPxJwDMsy1DLHH95SSWPrTUipT1Ur8M
GorQjSMiniDw1S9rkRIRXpHUATls35HAUZhVDem4k3g/IsahS6TfYlkS/RxTaT0VYpoaH8Oifi1/
49DIDpvkZ9ZxTv+NqDf1KapSMWwWfe8y4pEtDvS2IfJ84ZTVFwcjHNcf/Asb8bX2WmGRK5YQYpwI
3ObM6SbnOLLRGfSErrfQh8c9Dm2oeoZ4PjxolgSgWJWQaA0qL+JWdQnCi0gFzHlmpPx6ArtLpByy
AROl2qTGXuZG3b3szP1ou8OkWARUEZbl7sjlEwbZWJ2X2KhyjmgmrWtLxtMgnrGRaINs8eudOd5f
xMmyZuiMA0i2kSSExcg71aw9iFq7AYzrlC/5BJ0W/lnBKTC6R2G2oRm323g6Fw2r6hAXJ8hF5sXp
fS7O/af3dCagWjXY9qDMoXtoC6D1/qny5qPcoeCY9pS2BDAsBqYcO2zqB7uz3bkeFpoREfvTJstc
Tx+UpPZVRVFkpdg8sZXpe8rYOBIqqj7znM79WkUdC+VqoPZMQmLH7DuqRye4AJf9h386Wa1LYDav
/5m1Vf6g05CmAtod1GjlR/iNOfFWv30N++hnTi89XMLeW+SxpKBygOIU8Mx4mfKBFaMIizPs36oL
+sSVBewAAKcdPHpa+qkUUuZN6gqCfLp2eDEDfGwdGxHTKg44ETWxEzSobowLKQpuszrM+65zjx05
H7CFzfB5ClDyFiBe4Qyajc7HZF18+ZAsKhygxwJzx5KiWBkNBgLf5s654igaLz3kSyngeXWxbHm9
qRDKuM0CAicdrF53rt9MK3Rf5vO/tCBUOfNlULbnlHxFYpGIVFldgefHC+tfGqYohoKaGTcv8A0K
NnzaHk7cST+M9ocne8LqflPD9U7Ki5TT0wG6n+xn1/eY++0OvLjzhZHPjry5m1izH6wBIkAhEmlQ
NH+VKbtelpUdtBxrPAalqjCoMD3lOYiFdSXZ1r3UJGJTFxsejQeJpCBt7V1HFjs9wrqddFJWndAt
XtxGwBOzIQpbe9JvWEODGT3UYZFCEcf7qzKCAcs6ZuDfEGgIb7Z84db67h9FMFMHGnvsAE/69KVK
tKuqSlkcuhapwDo18YrdVcYDVL1dK3DAy2BC+nuRjw1reLPWU3ScuMxq/UaFB1TpV+KrQKE/L3Hs
fq4Ak0LXWfoykoCjQMMejVfKR66xJUcpwn2YrFCh0yfRIF+LpbavLSIKSsdX/WeQCANp3AZ+PB9s
uIPkyj6hn2aK/2xdBVyS3/+KO2fMFCe7EhVA9pBsqLaQPVgeNeUiMs2Lzpi0cO69p11KKqNNMohp
aoTa3aw5kta7szINKmfyTcF7Px8p7VXvX6Rq2lFZ1WddtaL5ebfz1H91ov7tLUqL16Wa3ecnbGS8
xB319br3WqzJ1JRfJ8xqLIEpa3q7WOI4jFLHliYvltMroJw9USUEoz+6BiVoW5JPD0HxQKHK82eT
a3vDhV3e5bdDVkQWjbjBdAB8hNlHrcgi4eblujnr4qPABf0A4XuJbY9DrmIw3sWYy4xmtSdttzuk
kJIDe1nwbUNlY6yxcZW88v6uqybJ+q2Wkxq1VinU+CKPs+SoorshI0NXNy1GNWmvHRHiqDaoSnSR
YDd0DGZn1j0zo2FGAFcS+JcviwiHjaNithkeJ01ZhQJLuRAWzIH60vrquxr3uTmJbU8lvPgP/XhV
y4W6PoQYBoW+gMjhetI+RvYAkTM75oaxcupJjAwKUeFVSLGFbqunQG6RMG8v5pXYQE3BcdxPFPne
IR2igf3zNf/8KprbaWevn5wus47UjPdoNbfElxqsv6l+M4u8BfwC+ZcdE1hUspLOJyasYmg/fbU2
phhLdrpYNuG+p/HxgM8rn49dvKV5+KdZ34s+uPp84GhgHU2yhCIkgNbW5QbbOCwtYOm8JQv8MKnL
I9BBUXRa4J6xAWP4Px/0amka15wuoSXMvPkMHeCNtg0lfG8KoiY6rs26mWB7n3KvYLvcIK5LW10f
Cuu/Wjol6JEDKQguILWXGNj9uJNJvsIoZiMU+WSOPC3/Oc1L4IYzYDMDZwSVc2QUMzNIpicDZTsP
eGvuDwYX8kJqH91Q4jP0PohCQifVztXjrmZ3DwEmVytqe3dl0NYW2GLMHyv7eP50AwmXYjhtQR4s
qwm1nKbyuKJ5FttQNnwS1tuNwrLMAwhJLCEtEw4ZNnLFhKgUg0bv/CPKM+WQaUYkgrOpvtjvipVX
SMfh0XG2LX8Kiw8Q6uAWg+K2k8FXWOISoEkpl1bjiL0ufDuzzRMlnZ33MUV1e+mQ0DnT+4DA3sv2
0p6XJvTQ0+PyETa8hN7IbRU+x1wdP3djrbZSWLp6K7zmBSapDZleHqt7XVP0jmDzt99aEgG5hcbq
CroM/kt4lhu/7/NNlmRdPy9BtRrsylgtpXuAT+/BaKbUjwwcwi1r2fYUnzNeJlq4fWnLm1cTy+pS
/v0ObLfmSFTrrXtFtst60J0C5dRMnHCfIqTtGxkWJLZJFmwSXUV3GUW6AtX2C/SNQBhVv289hcvr
4/aGqHNyfnvJDau9EE7t9/G5N3pFCZVXcYaD8RywKqshv7zsExx8TIXCE9TfIzxACNZvz2hK63VL
lxr+EbfgYizVAjK9wAE234UO/0UgyOeEt0Ka9S5Uj7d2Wp0XTI+aTzoLtRfzJsxWLxCNlOf5p4fZ
cFX2j1NSW6JMZM1BlEewWwUt4rjwpSMqOPI+5bbElDx+Nyvw20FG5mBQZjXzsSBENK7Ok+UgkEwi
0Seg2AB5kBdonmj5sChCpNK3FrPkT4MYxf8Ctrv8CtJMgTgwiCrhRKCt7O3iXp5T1/WxAOcK6w7L
VVoIEIUGF3TAfhhvEDpKHLCY7uB9GDE3iVcMVI7SN4skErAO1YRiVKKGsM9zOL2szT8dF16pf9oW
RAF+rHlUDk9dlSJ/aCz6iCqY6iM7x6OeE7l/nrgh+CBzMoeXo8uaEpkmQpovmM5UIe4c0GOk1z3+
jKb632+RxgN/SU3M+k3IhngY4CMKs2+sfuRwYOr5/La7wFslxg0gI+i4N1SlHwMlsJSdXOZSEJ60
8y2A2bASwo/03Jcq+tBodNs56k4ZSrTVwDChbUB2LWi2KUB9SFVTOgYQMSXstsnmhD57Zx/mQ/29
NukiLUnGQfEU4/eg9VjcvRZiMGNeOGTdzA28aUzP//K3tddZDbZraPaylckMTH7Vc5dsYsfZ7cmC
a041B3G/JaCIDP/DWiPEBZZoZnRct9o9o1ZSrL8pE8i4azsTgOBAURnOAB0Jqvc0p83tCgct2E0q
VM+MPtvHTUUxiAYCD1ODaRe5VEWmshsHt905Qk2vDsEn7aOPrLFZorKXk/sGAhpyjZvXufTINzzL
G6Lw1kuxkcc76y3ChSUNRoh2yyuGO+/4nQwc6K6H1TFPTs3vg+sAtyiDCtp/Qh5kYkuqPlta0tFe
/9L2XoauXggWAmNAEiUUJqS+qfqZg6+RH5j5WAKuJ4HAYdP6QVNL/7jz+v1EWjCDm97Ps4MxFQ5i
ydx4LXjB1dc4ChbyDjo19Y6cy0KXjvlzzFfU1VlDMQMysWqcgsPlzMccjH3bRiI/qtyYDBNnkhUj
5SzgbtKulQvu/qdp+t8vGIKvakhVWAjH16MAYaeOyWL0ooBM1qfcFLkzHfLmwExd+CTeSXhCYOTV
Y7qdQOpyVywTdCG5VsfZHEdx83xf3ZklHMmcKR84ryvqcsq14/26MeGKN1QoabRR4vSlTCWG24TE
hq2HkVyxaQ6oPNGaOhGiQHVu36tLEe97B1PjawkTN18gnXr9kLWdy6/ft/YcXhAWGn12GeGAEdEY
CRSyGyVxkptMeqqzanbCqOU/vrcx53WyF2MUcqAYsqWMhW5aoN2EOBPl15Mm2vIA8Rsxx5I42Gyj
du6ecnuLrFZpM/oT5b6uuyOEgGCMqDct/BbGeUYqz2H3QbmoQF2X2uA3Pj6r7+HbjQRG7TNvovAx
mqYSqyWtFfhM57d6zsGYqw6VQ2X4rurJiJuRnv8mOd6YzWCcONtvadg4n0W8IVu6sLIU27XVY4gi
dIDcLUeLJON3AeAwhdTPkMHpOkBGCUfNEzYcFTjGSQwBGSODahJTuD+/Ih2NufyCyv+JXfUYAKQv
VR1FOibh88jZn51f6qMOr3Q440K1tSnh3t7PzLL7VCPOxWXDvVLR6euSS0ux2DKXY1GyHeFMTKfE
o32u/4f6Jc1am3nhdIbLli0XRHkA6xm3y897x63mTVBlb7Efkb5gIlYnLLUXdCnWguP9/YG5Y7gA
I299t0tomnpL1T4q/ksQNFkH3XvN7vH1K96nRnmwUd8EWwyzNeLe/tPm9xjgLeXkuzqjA6P0rlPq
V//ZZ3dhFCDj8at3hoXV4ov2pAH6UcMNEWJyhV0Va8+08Sw79Ew+AmVenQjS/Jzp5R+Y4+5sONq9
CA/9NE9IhxJWlYy5dHXJhMBSke194fFvJYCqqILODo9BJCH+CMUTWNbzjtqdL42dG9h/wSgnR1yo
E2XyPv13vRGu5iBhOLDuOOJsMR/tDocMiOLy3b2k/qE4+l2Sd1IWSKpsrM2WAxxbOY/hO5Bs1rFU
MBRauuFIq8z2UzvlMzikSLF5kKQC7rbxe8FExvukFNCdbvS3deD9jwrZY2LCmBymAFQEyr2JmP4+
nr/6joFfryUwAHaNrIzWZfYK4sVKO1PdAxMllWvORQ59phYDjJFBKC1HrhwOoLuaDbxZfCueSpG4
0R3hZW6QH+Y6ycHqM/BuqosD/cCVVhge/69X2Cz9TU5EuNpKy/tLNCpyVCF21mPQgDeNPjhnqW00
6MlcFH4sqFWZ3d1cQu4XUVYB3/VcUQsadFpnlhHIiZ6kO/nLFaUwz10H1uyBwpZG2TtEusw1ohgt
swIhk3bH5faHD51DeUvXUPvSZaQUUfv9/Un88rdE3X9Bxst2ArI65jhELbq41lRONWDJ/iXYsvtT
FqEQrmT+r/lv5eOirbxVzJsGr9J1K2jTDnc7ac5TNztP/+1IPEawTIktxPwLfoX7NwvYF/UBnTl/
12I0s7x9w4EGPRx1xkYsifMneCHukqP06KoHRIPNZEtS2aKazTB3kw1rivF+pvhzgWrOMh4/TzRl
SbwRCpQDj4daqswoNootrbkMDDg1gVltNWqhTNgaPYcj97fIRaZvXjLstW9XKo4zyAIWhNafKICh
8fznFDPoSB0YluX9Q2M5x4ysAIV6S1w8/RznCDjgrY/SW8hFr/tMqCxfEatSU6y05lAQfbasROro
nFcosORj7iYBH93ooMXHr+fq3Ww8D7g5Dn++Nt3MlLqrJM/QknWXjnHQM+3WoxGuO6rbclgC5D+T
1zLGKGIrK0V3ZplDS4XXdrUWrDO7zH/6xrkfz8tTCriaV49LgIGDCLVD9o8nO5caYRZPDLYmPE73
4pXQXTyoijnawKE6GOBgjzKGKAqVfFfPUy3euqrJG5dSyunW3N2vrDJSF8k+N5eSBRMsYSEGyVxY
mZTVoj0KChqq6FMak68KVzCO/uDA+7l8smJl1Ab9SB0KP7yHODZJODnGrj/bW1Gq03wu0YoXz75x
ptjh0ONCMgcCXNGoQ5HkisnalPthfnhHppUBvMa/1TAyaC8Bd/4akkOm1iw5SyE0mPPa6eOhCVRg
wREj/t4LUsepM2Oc/CO5FErsJNFG782pZFa9V7hmDJIY6oROY25K9+MtOX9tvPNM4TpBx0C4KZ5d
NgRv1qUQSkPOe9LK84799Wxyvoqj21duKlWqj0/NRALQbTyxbdkSEy1qqthqLD8u3KAKER+XwKfq
3g87Oae7F1JdXh+kr2d1LD8Jn/IId8mXuQ15u/qC2iA0j1o0ug0MO5n8bjMcE+fFJLCZ8GW6S8ii
iZSaQA719grjceTSchlOcT1dObmTkUMuqtQz3zNOlud9LM5cXdGlgSXKtvUQzJi+uREMMF3lfr4I
7UfsmDRFAnMKWzUSxbl6oMlFZeLWqODBjQDgl0RS8C6KHeUp2KhRpwsMPvT4moTgIqUYseP+eE42
NjZ3dgbECZK+fPMNNiXVtU7urUUPh5IhizMHsFAEHHnNMLKUJKLoBletHWNh7XRDrWRH9oof626+
NsTom/gpE8MncZfHTtolmJxE6EBOlNLG97iW1f5s7ySno4CKjC9/vVyq4tw6/+CT63WLDxQCMw4q
q+FIZ10ifqAqAYi7Cl9Qp6Coo3pXlJj9vI7Gxnb15ILPswqprwX5qvpIx1dl7S/IVW7tXJzSqXKk
hLKWlWBrMoOrhFv/iIkcf/9j9yONsO9SBr5x1IXfOoB4d1fWZGfvG9dOkTiHeKzNYFhNhJdyMP4W
xRXk5GUH876RKOvqeWOLTtDNMoY2kZvXmqhaJul0ZsPr50kvK78q4Go52AiXnDiAKyLy8ylj+o8T
ygx0z/TNcPUbTCDeSKX1VmmUGvpPIC3+I2w1iUHQX2k2rY0N+QknHLbdMYfNoQEsdxEIrcjDHWG4
F4PbUARz2Zn3o4d6xaH2qHP4H6npg5D7bs8ffBYSYbJLKuw2XQ79iFoL28OVAe30wE3XeccTutjj
SXaz+Redb5/bruMAGhSZot/QTN8kldZdCTGtPJ8ZDctJawVH0Vtwlut+drV9AMnnQh379QhVtGle
Z4v4USs/eNoqGdRmrouR4+A2NBOQgTBrG1Rt8NxnHviGlQ8vwXX/YybUjsblZQKn3rg3icHHlgTP
T8JfcWFFdeZl1yW1ha2W/yf2KMGN7asoIhq8MxT0L0TaSOMsySNzEf/D6SbdtjePPKqDuCcmcZdo
IwuLQVhRIV5O/qT8kb1eSZ30hV0nRA2MOGWsgjMBFeEpcElSMC0vsebLOHi9dYfO80CTZTvjPTY+
JC09Gax5LVLk2q6kYTB208oQBrZipXkD8SLZm7wBz79tDYpSKA3CDDHnAAmeiubeY4W5Gtg/ACLi
y6r3OJm1QxJsWf2ijCq7uLBbRFxUyor4hSu9zXUl1BaUnD7IUpyvw8UMhYsnq/dEZFKuVrTGCnRJ
vjqmbBKkrQC9bSckJxjgPBThzjrHa17ko4A/yrdyIP/FB9z3e/1xYToVpYeDcB75p7tUb/e9mgru
Kgc0IK47WqVe+RA4nS67wS+gVVXhatGydXfueCpHgeScSsawJgZFqwtKYLEunufqR9vyKSIZt6+F
AFa/vf69TF61/eNUWQHWdra+gS/2fJ4t50wOtiXvqBouu4GAkyQEiFIoLDdiQvruFzS7P666OiEG
fGO7OoEHKJnUQSTL+/a0q7zjRHfMUJ4Ba7fUwLBnDajwbBsMpf1txCfw6nsNpUgVKcKlxHId8e/R
Tpz8Rd2DxY1tRgkX8je2TYr3lJ8cddxeXhbLik1Wobki3/SbJ5FNSWB85nK2KyVtKZQ//YQxKHoq
d3FG5zxONrDwJzIe7WxzicNwu5QbEX3Fdshk4QjZVtMAEEzoc+9OTyrUD6K8VDqqYpOKBgEMtZbm
cAOLC7XdjaEsz2moj+PlNlAt7M0bxDrOPc6JoC/Buzee2ykS4bAy/NrXLiUI0EPtGKYdDR/IhuBp
1KFCl3dCLQLejuDOkG6764qsaooq7FFqbCA1fV3SFCfEz4VXo1DTWL1nX6obupfE/SUzJCb4YaaK
KdabcspXNZWfIMD5s9XgAsJg2PNbFUwpR3w+4CK9Rie84FHMml05rWE6EpVtPJAzOxpfuOqYpAwX
mGB9jYz33dR3hbvv4Y0fPcjLwTpeoZC9W91q/GgdGlzO95pd94JMizGIvAQEIBdoJCeWESvEk92s
ufjDazepIvh8akCsS2zJqAb/cJnOwlPGENbZIJ5NIuAQBVHgGxu7KRM0C9FyUFqxHNsnw/0e6Jk6
9puDRG5lR3P1l1HHfBoQ+NObE9Nps+gPfPw27yiZsGE93fCnzHOe0jrP44HL9Ov7fv5lR0JSa8b3
bDU3c/a2vgcJOE/AOex9ADf3Jq9A+hIGesmnylKnVnnHU0338dVilDvMCFHk4uBaWAHLrrrQg5rC
LUz61jWsh9fUiokPkq59efndCkG37ilS06zRLDgSh+wjTwpRCV7+7/pzBVESdPfT0PJi/T/+PJ0K
PXCRibKRo9Sr+yPWEbTJfmlfv8H+LU2BMKcUzT93X7rEXJo5OYilQ8xFgdWq37g6+bn0if7Eh3/0
s8txABrrqpOt2M1rEIexCy7J4jMgznh0VfrjhrQrg6FQYQ6L2NKJeC/WIy4TVPbqbIicKVZ2RKat
QpqU8JgFZjsHa4jbiiKaa/KiX5aHBfiZCbqBIBpVNp89Cu0e7zdoGWXsUDHANn97FHbjSd68SItv
I0KxFjBGS/diy6wirb0LHtAEPlQ+w68a3k0qRajIVS8eC48xpFI5rNbXiH784sW5dkpqd03W99XK
cU/bLPjHNtv7edmM4/4wJokcFcAbJNIixnLWRrRBR0by/GOEFwyuFvgE28lzP9Ybr/GvQR1ekiL+
qeW/ucl8W2cAyyi9/1zeHBi/ynU9cSqpM0M4qLb+zo06HgA2pSGZW4S74B4p98Z88JVc/MvCsba/
AW/lBQS/LXuf1ihyxHAoZnSCYSDwwAjqXRbtxA7WFpNp+69ldgWwMlESmMvarJvaNmz569zBJxQ4
VBPg+vSPaM0MsyNbBwlg65Sg1qJVYkPBL6XZJu7R8jPbnvDJKcwF+PFTHX16xHog153VOWcCV/Pc
g2ao44Lf/3MzaWzrrOSKhI6vFVI7fyyJHv4RoR+0MKRza2sWWhk6XGeNofCTkMzdmDFSnXK38I4k
HBWIepb5nQ51kFqWg7iE/SRTgW8lNY2nInkr2H8qM0yoZUU3KVWaqoDHt3WKWxf21MzvaIj36xQt
R7doE1hIXTX+C81EFBivKio9r16i5yKDIDSbun5v97N5rvZytbJ8sG6wNv0xijbQTJ0WVwKb/i9Y
lGSmbgi74qJzd8BPXx/ZSmcl4tggqMKUX49LSnjbtTxs20DdaGhhMpOefgkcUKK7Wm/SVBZu6jtX
cMD05IOPn9FmjK4XKWBot5naitUpEz4i9grkH9U0MfX//16ZVQBuLrVacG4THDQpAH0YzmtUXlOQ
pB3ssElZYiyJJF6uSQ6462W9/MvhvgjU4ZJTUnj2VCe8DhPa3Qku0UOXloPoT2xW/q8sL67DAtxR
OQhCG2Le+KXBZcedcT7m0fUVnbmRF7O6G5+2Fu1LCSZYBTFOnoD4jgqNFy0wan2DoF1Zb+yVDJ1p
uYfcHbtmbeaM5j5KtFoVg8UVc8OrAg1ah78z5wglybnF1jayaH9QUrwqE/50D2UWjPsFVmb0K6RG
gCdV16P8lw3T1iXYZKrOxO5PhdrztAUDxvthgopBxbnonV7licCRM1mu+5TZwMvx/Gvc0gF76nMM
5cO11jl1T4SNbzkiFJo3FIi6/CvrSavIpvdFNeHQg6c+VnCa+rKi+zwJ/lbWL5ytxER81uwQdxyk
B10jtY6GkaBPFuHHnCyxV+rQL5c1tO5P7Kkxb3RK5w7EHoiMoPf3rSyrss1g6zNcrspFRZWsKo5p
4brRJ80qOGk6y9HoOOhrGkUn0FjxIwYepplfHg1adB3QmglmdjOKlWhpiBX2yd5xkBTqs7UEc+kW
XtDvOw/XhSVWQW2B7uvTCWjBRzExUPGuoyL9TDeSpk/Q/tHFKuoDwWvw2NICqFPUJITL0EjWE+/8
xcNNvXEkYwX6Ph32TqSvVF+alDdJ92hN5NZ2YSDm97aJcNj8XUYA3t4AL8ziuoS6uE7ydWpo3uPA
YAwRl9SDRkzw1lgPOKm/iKNVZg1fi7L/vvPgvJi2T1zN0dMb0G/Rm9xrsGl6Fta7JwhzCjLTEwXf
q0YB8tW0GMLAVUa4cMc+jwkYHgMS7kG8AkQwt7swpSXeTRblosN4HRCWjg4LC2Qrv4IogpFv3Snm
dnjGa4Mqx+l2/ttdMNwxBSile5lWfKbFNDrXM8TywyNObywBuZsU2defEd1PQEZY1nn3r22HB7f0
bbpMdWHtnbau1PWOWm+3b6LPMMfGV8M/+UwnWm3cr5xRzgTwoHuHKhMO0Jm0cmxw2dcn0ecreq0X
vcmvur0PqcV8fXwDTozwt7sPR68g6oQQqRKogq540xOaqAUvUX6BCIi5vm1/YP/mLWIsza8unZfY
pKvNwQtVeOpSvc553c/V8oEqUmg2+ZrNPBZJerccgNT5N/R3kCs928ZHlK6tmPV3I+6trD7B8aXv
rFVa6i1/dbst1XiHKailea+GTqMEjWsKmvfYMc+0FbVs15em2JTVQZ+UfJ74shKoGgz1lDY/bN4B
YTw20Ef+S6NVoOqjE8YtxtP8Z3zM/iZHFsOVW0GEc3CpNd6qZjg3A6evQZTYFNR+EAtuwcYiu3+7
Q//1XXm+hcEBLq38c4MZCJN2cbdV6l/S7EuF7QGpvlKJ+ZNcfYeUmCG3UkyscWhkdLUcF4abmGPQ
dVlV/urrEc1qBL/eiVMaudy1qqTzwFm/c6UXW8Tdnh1TURldToBqnLNRzK9cGmKpwrX4y1Sm835F
k1W7+/QGB1kpnU60ltMZ/XJ29Jmh8GTD/Hf14K3x0bI4wUnzNIS8UgAS43o6OcXEP9TIICd1nxx4
vG4xk161SSysFzjKnRHynYDDwizaGU5kdi+BA/vqve58Hj4/9bwtPaARgEOSS4a8FMCyDuSXJNmt
YQfAUnWcejZVNbhCyNOiwBPve3V5xekpkq8yEuhnqUWWQx+5R7skXhPELct6QdRYAbmpAaSfn4Vk
gtZmaw2yNpVgzpQay6TzOwEe7029NTrjbfX/wK6h9vvRcp9dJ8ykC+ku0Wm8khullS4WAwgtIsyV
wG5S3FrnHr0uuYLWgCu9ebPTQ7YfgKRbMPbmUHS6BdmTXUa8VBj6PvCK+fqMWXvQUV+/f4xW1PIk
MS9EHr2fGdrQFNh5TGDFMETqTcQYky50UmUfz9Cui1+KK0RhSJQGyAH2ypPfZl1wVSR39dF46Qnf
kYDyde7obCEkaAOBq8aRaE12nd3mWTkzIOQt8WyCNQy+9BPSCHqJY2+GLCvcYXzE0MmnSksTu4xC
wumgvTKYI1GNXA7unQgj/gnHQ1YvSWcpiaH1wpmWLLgfHrP+kE+RcHahh3Ji7IHST1EAhXtNpQGf
1X48Ce8Oc5qjlyYTcFvWeDQ6DlWfiGD7ltmUKMy1/nYJQd50mtLNgfZy0TAvBblaJRgyj7VI9G6i
Ne+y5sPmrJ9F1QEfTFFYB8IhvEaFGLVcsOQsCuQpg5PfyUCTv+gAdx9SdMAWNjwk5q9ST9vyDYTT
XbZmMnoQwaMZZEmIkSqa4TRzGuokv+Y9o3ztv+NoFKBc99g6ErKHl0x5pMl5mtjmksa9a2w/+2Im
rFglkJ4Ie2/o4xiHPixMmxT5YTB89ZCMRWKxyTBTzPJFK7HtBh/Iaa0g78E4rKbUS7BnR0HSZxOT
ipoN8ONkXZoeIJdQzVYOlo8Dn9ZYS9wWnKnS5blGYjoID275tty1CrnpOxJrRCM5eGWcTHgnK1hP
042eE3ut6ALSMRs4alEWn4PpqAOdlQkkPQekdK0mMUfWGHclh6mopdIIxt093AKGIPqv6SvS1Wkp
qiiHvaIcg8ggwgwCDe3HeX72weoe/mIFoUuvDQ1o6qOI+kpZ3o+NMCwTjz+kofcqJaAGrriSaL6q
DiwHxgemo42F6ftqsTnt6VB2zd4c6foB7kQXQKMyLYWahkODxl4/V8I6L5XA3/cdJtiH82AH3iFP
8bexeXcIuEGkBxknRZcUWS8BUvBGh2EpRx3Ekwdgxb32PkXHuYG6yPoeUUxchns6j48V0Ewv2db5
tiTF+RnAtdzX4QXwYUO19debYb+czR9jeeOufTTlGCp2/W7/p/LMLhtr0ViE63LKTZ3ZJVXOtHu/
6LlagUF+K4d2VyqJlo8KWmVlqBMlgLJw00QWmFuRb2fSCgaOd4CIEy2E/jSYxjDzstOxu0CVVcJq
FdDlXWHMricgD+CoeRInyK7DdCVoVvumVx0EBwb4z7RcBxRYXu2mJY2je+72iEcFzV/g9avkcTuz
X9iPHuZOQbQkJcM2+hDaSRQtA7MypFxX4nHPYOISfya/DwMV2ljPUpz7C0rAqgNFqcJegM48iZ29
3MDhz9WTjsKoEBYShFavbEag7owrMQnSNnR8j/YT2ZMwkg3Gvo1B1g2tPrjLGTFIKIixVtPLqOmG
EDU4IlUZpnbHvZW7BEkeIAw6WWv/C6ZBnlQ1+TKp9jnva4EcBl0PbI3lf6O9OSyXPJLUa9EFqrkl
jbvKNY9cZpbW6e2dz7JOSykpOaFMZAGfiRMHseyqvE1vDGEQvx8zKjXUOW8QjtwAMLhHAsa23aay
yAI3IL4Rr4HCTbhoAm4XzUA7BG0qAvEgevmh/UkaS0x6UvI6mllRv+OEVl4OQ2UXM6GGrjBs5LM+
WTVm1YHBVdEN+xaRZ58JA5Z6ySCCN81/TxMVOHREDsxgZcw08Rkuijhcu66EWhK3eaKeki48TI2T
iO6RsEVfm91XoPC11l1WoWQhUq5aHWWTc43Q/4ybMbazXcUla2L1wyxZ78/aCNpKz2U3zGYfYL7J
qvGKJb2YPZLxJF44WrqfJoB8HZyLQ3XoCqrrceCjGRG9gYrUkJMhIWVQ3ZTMPkv59qguTNOX+oiP
6VEsO4uLNrTmQkB+ZHatM2bErX8EJHMkDSliTGxzpb3OBl0FBBJbQCdraFyzbzNH+Lw6PXoYhVII
V8cDKStaPLVoEGDPf1YossQe5lFJdo1YXvKRrCbi5VGqIklwtNftqjjZW5CChXgGxHKghn5g4W00
MDZrmBqpZC22rFuVrAK9Gfei9orr3Lfrn74zXG9awzslJXFZyJ6L2Nzp8N/cq62DbyzFsapW9A3P
57jnTszLzQw5bjJTCidRnZxevsqEeu7mD0ICrodLpRZy7TKF/dnDoQuwpcXhoNwdZaI7hI/aqTfb
hlKk7uPETkG+ABWqWHm5G0HJoG/7ovCnCrZ8OhT/VDJKviYXqrNNPBMzeOI47sYuHkjzx2cx7Hox
HTZA2XhsNrOP9SBboYsLJuiHIGB38Hkk9zSAtKOSZ1Sy0pVAlDnW2J+hfReqTvsEmLdB07iG+Dk4
wav/+CUNy1H7I5oyWFZ2b9taubkPUiER6eyH8mTZiQNXuNc5X24Hrv/mSkPf3uoWY6RLl1WQT3JF
ZVaIAxoJWqrSf0Y6Ps6Q0A9NAvfni9EJcVdU+3Z8eO9Vv/n6MfehsfwRdMBQL5Va4Xzo4wzG/AWf
Y0ndI0Ja6M+8sL0tKDxB0aVKECndBgs09FYUca3NY4wwaw2CBORpE0p3QIGC/yBe+m85usNfT9Pg
j7EpruQ5s3E/b3fH2hETmywfQWEIPgNDFxKWCzBjXHhwjDniBEWj4rwDZR+Yj2tThqE+vSy0d5dd
seyjO6cKJK1OwORrnkIhyzKjrebzAccgTS6eFDGBuGONAN7BX/9eeW2kfhRF6exGFv7BQxNagzNl
NIwCQ7z7NxgOBm/veBwnoh1AsMgN8z8OpkWLARotXrlCK4xhlQIj5VdOLSBfJ86RSeVeHo988zsa
k2gwAqe4J3jAxscPZVWk3pEbYJRtTjSrWYUDDwbaAOiwuOsTg6JRcU4Dk/O6f6/+rEfkh4Ozxec+
yVJ/LstsMJIfZ9xQKjfUoIn8mFKvlOdfBK208ZCLuKW92F1H3gyxeSwcAUzD+NXn3zSj1643v34j
Nuji7oZdjajQn7GVxPNAHMCoLnW9jTaOQGY3ngmjQEA3fSPNE3D03SRlRg8MpyfqP+nQiwLDkhaj
vMjOzGDvQnWLVNOmUSuTAltLIgP0SPvNqCWXmwP5csdGrxPw/bdPINU0cZEksb8MgHy1n2+/dBTz
Vx5Vb80zLe7eUud+5VPoGK8JDdJZmLNW97pFmj9rl5m6K8VCgABgdYKFMNc4c29IxPn4JN/JyfzG
fbzoBIJSkvsVnfo3xSz7fQ9qYK6bG36KkdnEzTzFIGlj4O+U6Yxbl/g7mGS8XzdRYTxpySSdI7W7
hG6F1EIRv3LNKEscZf2LchmyQIAVlSqrYy9IiSW+c0S33DJ1o/ZNY4zaBmaON3iGo+EtJ0VNlNw9
SyuNH7e7v6cD0y2vEFwognWe6gTuzOXi0uU+wbo594IdUn/1wHk54S1D2ezCoCO8gY2vNh1s74Y9
FymEnkGfAaX7zm6EDAha2ab6jyFDX1dkGbyKnkpDOkquKeIiT4u31OfPgGNKROQc6hfJyKora6gl
TZOM3cFaXG/O0a5trw4IxjtCeSDTMkgmXHltwG3t2cOE5wI9Bu+uadJ7cwRxp2HanRe3UABP51kQ
FdaZwQTyzqedPNwwlWd6XkFZj0OyMeqFPIupRBDyH1kRQqu2PB+zYLNdKU0i+bGPfmnT9Cb9Hb3m
BEVnqIxxz2uYe5SIsy1+h+ZWGSnptote6rLF/hCtdZqJmGJ0LIGlAq4XhjgKjFDIAfBBuKRKJezO
ZDe8cQlnCE06qO6rwL9g/Iy3uKrrMddKoFkFyDbPLrKLkEqiaIzebmHSf0IUKZ5CzQoy9V878ahQ
scshaVp7+ywEAIzA242HVaiYZtSL92dO99GDJxKgiE6dfXm/xn8PynpWAqavTQSYs8Xh3uUfdT3Y
2NVfX7L3ldIut4J2ZLT47Is6SDsUSVcWAhUGx3FOZjQCM3Xn/4oKQbWOAA1oNhXW8hUj31XCKvs8
ivb2/y3VIen/tMLUPmTTAIPbT79bTqQABC8WfTCg+yMY9uJ1hP8Q2i2M9zx7D9A3B0rtw6H4uThC
KXtSoJQ3XN9TLUMvbpVT6CVOTVbM/8Ch1u+OFAprabvj6vz5VmIsRAryZw3o2W88rHi5izhtTQbk
EDZLfHFlNOWbiOlIxJDcNWiLVzlaJcoo/jeLwNADYx3qIEvBSA26+M1cFUhy0ieWRWVftSk00iTX
2lCttYrwK8KQ573VIcXUCWLKkSWuHavZjB7kZkyxQnha1FeLHYUE/N5aoSyH/inkC6xPMGsea7PI
PfUDu3YOH3aJLQQ1lccEQKo8vj3vkz5kUEqJ1cOzNXQbvi5k1kWe1y9+JstHTTeNtP94uhFZaL0j
cm6fE+tiWLHxX8Gcpdk2pVLON0lTchjJ62eqEfmlmxqjLnv8vzBeBhTvxBIG33A7Izfc3+3+rbLz
hhG/4J8qYAv/u08kuaKJiR3eqI0UqtvPl7DV6xKjfnnB1rLHNFh8NJC2ABgTLOh3oYz2B2GMjtLl
lHaO5rVLovqCh4UGXlRhuDVenZsg6urf+VUBPkE5uPrC3CiJOy7LVc1RuPxoCMBCC1WXjJkGy0jP
N3sJDPpsuCo5GsONoI7hLiE2/WHmToEGNhuku5agzHvad+JGZx7De2MXVfrQKCa0KX/Pq6ZgAwXo
4Y9Cd0o8zz7HtcfQ05C9+uF156JVbxjtIQSYEZmH9ablitf9s+kEcuoPIIa2hOHlpg4JTk/TX1ZN
0Wroyv8Zf8+eniuBjweMe6w41b2vuWkYEjmazfn3BlSWyaep39cRbBls488KJ17399x8dyN5NWu8
GgGdlKYbOP48ubWL6PEpxaKh99fA1qmbewmiojr8ujz+dHgxCs7OB4Xkgqily8S0m0hUDj8CtQLI
v0Zx9JK/f6uKWqINfCTD8nHFovxIKupwddMZvFCba96RSC0etg6mOcbNcMj5d3yJg66/nIuqEKbH
iOPG2w8JJV6SnvnbEYcXCcwmW5qUZOycvkVMhh+Y8v9aOpYjFvHUcmNJpWKBYYvJ4/reRgcxLbvz
CZbYSSX2yTKXZjZ0XJ0IOARvzNnT/DYNwR3tygrvODxzWl8mCUHE0m6hycYFgzLp+NUmE+0qGRhl
xYdll4ti33GJGjYcIC7FtDTT19oLhrWDttWNL+CvroWxurkbCmnEbwudBA/gYQctRcp3QZqD50WF
nhNfF3Opr6H30R5olwW/pdkdu/X0htbGre2GYAmVxtc88ui0Ricv3YL2F1TlLSI9lcNmLDlRsPhw
CIr2W1KXdLQTFDFmlLt/dNMjRBY19Gir8uCNVkaCXBkzrPZnVqH96etMN82dMKZjiOsunwjdQuMO
QwziDwrgiBc4YJah4z1U05+/Yy+P6u4USGlorRjwHkpwu9OheTOxBXleAbODFgV9KU+lY5YPJmgx
eYosggjhRl8HjxaU36wt6gkSCi1b0Z3cgw7H6r/Jb47vRcB4ClbpDhQiHlqGYubT5jyyBPrGtr1C
inX4NNu2j+7G0PI1hoR7+vxcJUJ7lWzetVXxMJqJMnq18KsHfAVvBH4ZPz60fBGZ8Ib/us81ePwT
IOb6hxbiQlwLjOz1fZjUVXKUxhoK09PRSyyuPihUYidXJBr+hzouZZaSp9KACaRJ8OAoEWDGxb9o
jxOQHwRPNZ1ustJJD9PDSuUupTG9s2lNs6QI0gQRjB0uJo6u5gOlArWujE7ZcOgb4aU+vMdnQUKb
ToB+zepqPRy3Lv+ZveNtDK6Plx7oWCRq8pBeyUqsa3v5G0veocqM6xIyzvXxIB8l4CfEaoZpHjmQ
/fY8JCnG0+MnmSM4ffv559zjRLoWHmO7Blh3aUFV+OIaqu9Q+hq8bNosos9/noxkGHBmJZMG22AY
l5uTOh7jpZPgZ5x11mYTzobqW+ypzghgQIddH/jD9X+rTq9HlMF5QjGoipP9HjLY/hBnAHH/aYSu
mIjE8br0quul9kIpVK6gVATmBwrlBJKb79VV8TY7Y20hAPnmcym9Gy9hwroSVzDQ2CuwSIT1Bddg
6QjITsrBdchFM7nr2U9izWGnMj7ucEL6BtMJfvv1B5OWr+U/Y0gi+vsEVPfu0coTMRwWIDPC+Tt8
v3JDkqz3jEjg/yMwqt5jXsTgHm6nFSO6FPxJZlpQxresvAugqA8pAj39mR8ta609otz2ad+SS4qs
o9tE0TlpHyTaca721vZP/KtditPs1MksOBNjyz12AgyiV/lMTrsRaob2cLCw5J9DxXMwA2bAAy7+
rsuEuEG+jIyEnqMd+k1TC1TkZw+myXAonnOd+VMgQBFzfToZjoxY3ONX8z22ZBy/JHHdoRqSK2Ee
OKUpCMP+NR4QLfSERiuQCOt5P6agVyieiaSLW1a44hspSbjD4T+F9rP8SiQwrMfYSEu6FzlOxtUo
2Vtd7V0kSl+qxS9EjnWWe1QcuSUaeLk6V5iJabIdp6Zlw+1DRxcA8HmzWuVg0pLGGaeaYbqgazjz
XyedCI9YPQcDanwPpMa6snKvgGoE4zRuPm85PZNCtke4WAlPROljxmfLS1UjIlB8RNXx23uutJA3
GKethAQHrFv3OEMEJpMtT3tKVjSDtZT+foakCAbBAbjbJ3Tsj+HraFpc6wOI7t73nrk7H2Q9sLek
54HE2MxSH6AdHIVz1sKPGFLUMmu3TFwcbot2PxheCCL0nJP4qbOl9rPsIqQlA1t9vc0chXmwyctJ
OnSx0dbD8NDIZVP/6orF3VUN1zaCEiLDU9tmlIjck3Ik6EBTxIx3kDl8jeykLMTMchFpxhrG2Ozz
iGhzYpSWBH9v672x1ZTYO7gT/3GkuXmUcg2C5nei14H7RoKbddrZcZtpQZoqidLjxY3jME2GCBB4
l2dJUHpaVYEMwjAsFtseDm9sc3fbkyl5/uy7PakftSg8ZOdiiIvV6V4n5iNpU5wTIigRaKp5rAsd
NEU8s2/JHQYxEi5Y512IjACXiDetiBOdzrXvBoDFpk52OfdR0NbWilHNiO0qrD/YDKw937GLq84+
7/MYRASoklvdb3NgXfqju3rZ7i3e67BYzGeV+n9eqQ5pFYggn2U43CEcVFiLPSNgz0PSgZIOBSuN
RqlaAseodjJkB/1OmzsH1MV+mih6iKWV0BlXNjYB4gbauc6mlxoiA2CVlIEojs7sJFrZEGOb8asM
m6K6iiWferx2UlPnFMDQgBwkreD11LCyZ+6EesJB1pBTbz1EAD76ns1UqYXdXLrXMwU6+mEVO9FO
X74F2Y2g0aqva2ua3BY8uyaGadhmzI6xMOk3j63shOZ5Hj5YwwedR/wUnJ4foWirZGcuBnh/X7Ty
PcvOvzPben1EiDDRqolsF1+7Y5YzXgaapuj/CYbdNxEhRmkii4jGXyMGaubQVcWbf3s+Acr3QY44
uVl0XoabD3vlsKAeG6IfwmRbRyVYfYIyeAhAJhfczZ5Dv/NArs9IujTiRPkf8LAewcXTddqbnwro
ycqqptNQm0vEaV3Us1xutcTiViUfNXY1mhkpznEKL2f/f+GqleTGSiTu+52WUh7n5mfy+6j9yobR
otKSktVLYdDFCV2hAdjI0pEyjxPcH+/Y3+etOFAWs29wnepnAQb0On1QLw5dfN+PFdHTBUFKx7Xp
TZYek5KpvIf0McfTQbQ95cfNB7UrMnzgZCQyepTnxR8+hNqICw2g+jhrUQtuzK7Zb1JGboj3/YMB
v+rfKam9rIqTPbJYNIm1e9g4NhGBfU5S/P2JNbhY3U2Bor8gQ84MaYf/ZimOb8KLuV6D6DjBpUcM
F4hMeiJcpz+2XfTKdIPK4K8uxSinjT8iuRVVj+29+3Cgx+ZLI2GdpkOFwG4W7gUDvhrdyq433bzv
af1dBcd/Xx1mIlOKkiNAm0yOryvnE3vP+XZWJuWxh5BOGOcqnwITky03NAcvHrwtUIS9t5ya0Jqa
iQ9icVxuL8GceN1RlROnllB3QIsPCSpQjloCUxEpNrcsOod1dDSeds+epYMd1eRpsqgkiefYJS2u
m2ezdscJGr336eOhRxgHtyNKCv2blP930pWgMmp3YZvdm6LMp7LQHBIpxKd1rZmD0Hxw47tXclgv
MAtCV54XSgJ0XluOU43zNjgsx42pOQxzbw4LJn0tctZsCl5DDPZYaTvYajh1G/eAMvEGdnVrSrKG
iSEL7/Ir3IJbvnaNnY03QE3fvEfFTDoF0nRiGZK4vYhnZuYxRduCLNPa8QtnTYqkTOhMT0JwMBUH
iViDcHQ644aKq9gK9/bztT9e2XSiV6nmlZBGMhAZqLcwQ8eR0d4MOwVHfhUFzFdS+unteB/tg4Eg
3nu+V18Vf1Npl3B3wjUHkAuAi1fcLZrPO986OCDX9vth4msf8wq0DTJ+IdbBy0ANgVZMXdM/lzpZ
DciA8u1NtGRiWkXZzj7c6ocieAbZqqkBlqf0Z0misNghA/8xvhIMLqbpzatTb6bIP82w20APh2tL
nPcZLA6UT/No+WYBb6YC/9AdTKK91KiBwbrWDqgsnHpofVLFQmVjKEuzVq9bpFoQVqovJ3CeYPTD
CZTzs5LRDS39lyJBa06/OUuNy1oBvoY9Ow2gkpFuQkgfgbhmsh3UwY4oTpJBCPoMpIQxFz93uNFV
8P3Weon6uiMrR+DMLfU2QNbxno0hJS5LMpigbhWeaVSFK1TIbhwZ+McvLrXaPuQWHzF47iFts8gG
gAwOnD27jABG7HyCcuqAnXaPwcao6j/707GJcHjVPJHSJrrzzwla7tIgiuzhTcK/zs88z68xivXz
26oCSAlXEYFDMvPXYjmlR8zYS87tuUur5Vl2IeoRJol8Va2uRPsK7XM0S8h9FsQmz/xFyxRG3VSE
Ea8YEjVSxMQxjHgXd/QarxBic2gQ620QLpDoX2O635Le4i7fhTB86cqK5O5sFWp+f82VMrPzDbzd
nt61jzJhSF2gKDh9gpgNHeaJwpBxLLQkpEU0XiqBggDQ7leb2aw+giIWAZ0zs7qEyaTwTcilyIOj
AfGnZj1PKG4n6H8QEYuF8zMpN6vBE6NqhUZwRm3OS8ljOBmHLPMi7iXAC7UAtj7YPeQ+UKlJG6lM
3zg+Z1K7iDV3CxxeU+sPxkAsfV6pjQqjVppVmF742NYVsBrqqs2zKFk3RZu9UlHYjEVkMQOuSvNT
K9RNBWqtb/Pt1QT9G+iaTXnqjgNDi0rZhmyX2bs6umh6VUwCnKpkcu/89wFFFaTo2dFVt3KFGbMr
IZo+rJ9mG4Kn5nkskQpfRiIEAjGJdJZhQnuqrE0gj/yOdQr55lSx6Bo/55MyyIz1omQyN7vMiNM4
Zj0pwYWAanccpOAgfmkiY0+c87oDd4tXHpaPRkGw34pnABSjaP9JygmsabZ3I0es4+nUKHMEtLgV
/xlmlF8S0KkQCQtQsBIJXoqOrFyhlUZw9ie/8ni8P205zo2WsX1SMrNsv0NFnduMttWKzli7wrcN
ngqjXT7rx78r0W47yuAlIt5v6bzzWOegvu4gRUw7PXJoAJ1JaLn2dX4HclIOnvkQ7PDULUes+7UK
HYnj92cde9CzAUnkaWD+nTexkrh5Ol2ojEXeXMZDTbDC4FRa80sGReKdUV7oa6cbxwJbO4UOikKf
Uv+jsFCgMoqwwtEboEBvu3OaL9dJg+gX6vuC7C74aX3wCVgGDFuzGmpvPVypnxnXzpw6zuOJRvAB
I9/J660+Fs+Cb+wPqIiDv82CfznoT02yUkEocHx8s8fQUCN44O4REc960/S46JZnhvt71lnrzHzK
B1SqVToRO8uTH0nV4i6gNq/i168LeBWIx07P20Ep9DOF+rr7eMzl0EuW6zRsxXLqkEeh5LxoxJjv
26LQsXhlT/lP0iPf/9S3+JYxYNx5hR1+wYybsnlnSMj1fvp0Dq9dzuSNExrplyHIlBbaenEwWLJb
E9ZFmIo48BnSn0ag1Y0IUPc8xyl8zba7Kno8R2RLA0Y8VbwRiqTRQYt58VorIiQUhLMbyHPmjzWo
4pL9L2QATd6quBQMpbxzlGWeaLMoK+Fw+ukZPQhwMonpWcxW4EycNGlCp2rhzgzxGf/esMG3Cc0C
PrAO46EBAcPNQ5cq1GL2I1A96P4Gn+aXWGCJlH6/PhBWns10p1Kq5tBd2LPz4aPQbeVZgeZDfLnt
L905wnAnsPoNYir9ZKg7cNKLjOWit84jSSfJJMsVNwLyC3lPEtchBV4+llOzKg+ToisrbyKVIdmh
oJw3u9uUcHmyaK0usg4q7KDqB9DXi6RwHJ9p85HwL8aIXg7RgajP5VofNiaMNreWLplmy/ijxqBt
sSnVT4C0mGnqMJ0KFskP8u9mitrP4HwEGavKDXHS2tCZpkg8v1REqjjTR+F9a969XaHEkEkVDtMB
+XhKr4QfFLMY19HKfXN+/LrtilSmgm3g3HyUdipFw9E7alze8GlbGsS72E1cfDlV3usyL1sh49yU
SXfulWn7c+MjS8tft6DnMQ0jUwADvglyOMPOkjUck5LQem7gwlAOs6NiQ0VQx4q2c1/+LPElLvQR
BwAm2uVxNbE8YilIaiLJ8+HbmdbCJM3GZlAMtQgl/qaKSQgMHYYKZ6ydOhJmtVL4UZT/n3JuC76A
LMd0IvUJ+AuUruoaTfXovW1hfKY32uI4G93BNZNyyvevKXqYUcB5KIysPRMZsh5j6mE+g0ztYc8d
QeNGT5Tlb22fxxnKfajfQ+KGDRKpchWeKYpBAx6SOxvGn8EjyZQxUU6RoWG3mDngufAllTEhOx5N
aor6owb+FOjLqEwazgNd4ykychaO2vLkwnPsEHlyZWzkgLQiwE1L54B74LvWKZEBfgoibg0KMqqh
1DsFLPjPxsoSvdpqetIj0umUEQ4KR/6vOdjiw91+1wU/FPsjCarEPUp+kUVWgMok2YBAm59R90AG
z33K06w/rOjbaaHxgqT+/2QhuS2F9iQoNb6RNb+DyGgo7czrHB13khQCtr92ozu6syFRB8IPp1Jm
EQ4PNChx7406p+o0l/r3627ct1/Ca68yXbmf/Cbkr+nSThPc4HH0U4hO5OAmNHxHiVYfQsmB8AwK
28TFIhZTivZztzBS430uAXAhMHDtshb9I9FP7QeY1xbfOoRGcakIdfV+7oUe2mP7QZBl3FXCVKHG
STTjGDb1IUBjEYHQTCQtRNXs8MOiUPynvQs/7G+8MNJpZR/dwkDV8oqrj7mlHAJaLNwwv8jJQR3p
tKqzf3rwflUOddOcZw4kKfkEEZFLulA+IjLdC5MDtdsK2dgtwVNXsz5beesMBZYcAwSfOeHCSs55
XLuTdK0st9dYH50hv7L9LChCc7vauYCi3LttTIgWStJRrTDKeu7JP2WHAfSXjq0X+pJyEZs2W93s
CXYRooDMDiIC9T5zbTW76RNRZIZarDSsJr6cl3XH+Lo4sUYXyLvLSV6ynfUqaCInh9c9D/WN8oUK
WFnV9eZSSyHVkVu90bGWFPoNTScEHgFp49VUMaft+LLDyBctDUgArIWqgCgO/sUXiSiFs2iuG/jY
/E17YYCfWqJwq97L2aWyxhfaZQJ9pj9n4/VJdAvO4KfKw7WHD28WZ2u/A7EnBRKt8mJVTGauwerM
dmKUFmh5fXM4D8D2nY/b3QdZgEm/AN+hwJH5C0fwFqKBY8NMJIFqICmIIMxaXzaDNP2bhChenAH6
IJp+q5MG6XVO7jeSwssC4htakEAJ2XIVraE3nNuzyLaFPNAe/FPCJU/BQ+AUFbGO2MAy66l8HQoJ
Ml4GTChn4e3yf6L6s49yFUzYudgeO+JCGVyJZhDGHY+X06OqzP82v6o5z62rkbr8Pq3K81V7MdGD
KRF7svnYeW4URqt7h+HOAQJgAhKrAAOdHowIlqLXThwnV68E6nlVe27l9so4puxH6pL7y1VywnEE
6PkqX9B3oosscl4wGiuaKs6HcKR4gUAUp3lhltguN5IhV/F5Wd+PH2noor12ggOHnUHLPNnOHZca
Jvw+KDu7b2mRSZYR7btmKW6+YI1mMn1stYvFcD6O3A2ZVPjBaU97ba2E2vNmOfKiFTSr+Y08mIlu
o7+pURzoB3SUKBtT9QKmBSZoBsccnmqX7JVam3owAxq1X22ViQeA5HBi34sOiQ4zS6npFv92ZNwM
XNQjszi9bZPmBi88Dmxw46oJvixsMwhEmTLNLG+Z3BHGdsvH4mcccVfSh7k791LHSFyFyCZityy6
rDoNYBw3w9BlV++4cc17PGOGYcuiWjJ69WV2F6KziUbGreOz21A5EivVOSwZypPQG5rhaUe0WJ5s
Q2UqcjBgaEVaIceio1v1N0nsQnHaa954tyMxNw1M5FHvZMPrUku/8DEQq8tBJilFTdBuJwzDVZOT
AXx6uW+DuXCDeVN76hgnpn2HjHPfO4iHMAQukzPbJwwWnDLQHQt73dgxi7dDqmzZsITj6sYWhgSD
ttavJJ0aXsxBt5mlL+nQKgLM6mawBREfhiADfMKVFzZRvIgGaBlPPUiYCDE852TtFAI/a/Bq3PBL
0qm4Wq6M4wHrwvzOldTyMHHhrpH5p+VxOFoY54luU2qlMneVNra423Rn3r1AkpWObL3nqQB9L54h
nRXYA5EM1RywyYY/IPSp2X8c/dBfSHpQFO1eXu2uuMMiMo/4CiM27VMAVjFG+QFaboUbr0psaCnu
68yhVcFI1JzKYcv0lLm1HCAPkCBdOBZJyt2deGkNCnkHKmCdInKUlaUfXYgDpTxMknkzD9fBzMVa
RzEuN2mLmMrPrbgnGrx9I0JT6Cr/h+us5G88Sa13Wp2+k9qgGyw4MouLMORV6pWB/lgRI6I4TFvR
sdZWJRtV69qWJhwpjurSemjYx6DTnng/hQHDCaqjfdZkAtMVvVLybsccqZLYEgASIeIaXLiUXL9l
b8cPJu2sb1TWci+pR+46xRDofhdybvO185Y6StKPW3J1dtyX6aNT83od02H/imv7poUfdwF/DFJ6
jVwfxi++/f6E7Kktvz1i1rxBQrqPdiBQj7+bFG7Oaqa3uRlizwHRKAISU4U7KQJ3WO3whvE8/6ic
ag7NwN+QZjyHenDwa0CNanOW7M9tWHBOiN6MSXWkIWxlS8kriHZ0+iRl8vSD0uxOY588aZ5Quzh3
kkrafXB7UIMo6+DQ6upKt/8tPZUaBjdcEHwbEoJ9qKwn5XVCppg+pDgbiYb1lFhmb73JMRSyRVz/
gfr1XNKX5XklTghbHQXE6N+TGeLq26DfFOEWaDR3p8jes1MW25rxicZc7V7+zDU4Dzd6a/WyqwKd
tSWp0xnv1RwbQDvqozlg0wt7q6Eq5HWc7T65EIQLuFZouPA1AM4FGsz710OoIcUb1/w69F8DWlM4
bihuBOP8flsBxAf9J7dPr8AY0CeFxehBMN9pvct/AGOnrWkgLiroSRGg6IPJncLX+NxIcVafY8wD
8mTaUUBeq7hEkjjiYEl9IVeh2/oExynQnuGXoLLttW1qyapmKa0x7bmdxgEgbMpqiYWrd9JQZpUr
SKR60K//eNxGaRg0JCNr3mav62bd428zIMauqYDoTGzcf0dS5pk+tQeo5EvtqDY3P7xgKNqQY6ni
mr0trfD4RQGUasCMS+K6jSkZwnFknXCRjSfnR59eCb747O+duMcpfrQA6eMpMe7hiqUog3Jo+iXx
vIWy/37yP3yUe9AGTTx0u2vs3R5GOyymlF0qwxL+jJL4m3Gj+mSVzUv7DpYH6Fwl3hOIHSyoqP7q
96B9irMBztHeXltd6U/ak9XzjpGVTZC7iX6ftAHJde5Wo/j6LrMr+pA+84nVahj9jdNHIcEAi1OO
soASsgaooYzFqFC6j+QoBfKEv85PKymKmG7TPCMyc/+WdpG5B65YCwMLpZjPCCpWgcR/5Vrezjqc
DCTw76auuJKMEAE3W5e87IF5hsE2x3ziJjyZEZ6Mpm1OHmGC6qp5VxOoWcMzEpHs7GRkCqwgvsm3
BFsmlxfGmqTD+3uYkd9ZL3/Rrk8bR13Bxc5uUvyjxpWP2LI6fa+U0wJVQx+5nULtUXB+sC/XjmNG
0L2EPep8FehwRFZk90IYz3gDTPH1zrlXCHjwZQJWNUxR2wp72qzYiBR6z07vr0PvVkz/B/9ECZYa
LJXV6kpGOurrtrG1C0AWYECEin4zDjFl2ZraTKL+j2x92t5X4JNSa5KdI1OOGS/CpjcXWrQNOzqW
k31s8fpjT4CifGKyhCuBemCWl5PUIrYDQcQsMenooHN2gUnGPiDdct6Vxw0dz5aXrLahTK/UfXJ5
UT1rkTSdKXYKZDf938Uqcrw7s9eyuqLWkhHoDoFe9L6iOdcX5X2r+SHvsrulsWRRtkBD524gw/8I
QeAW0IniSzPUdIuQWXCj2t324efae/07YBzTIrYM9F/cL8Zrz040hDvFHARFOMeQnhQ9r4wFnjFI
zn3axLroiqP3JnC1oA+aBZYf951LUmTXS2xr2p5ikgLKTpI+TzdmpTBEjRVfBUWYGjB7qTud1HCl
MEfMjzqx7wXqeNb9VhtZP74B25/cDKSqWZsUDQ/msBTsYFspit8q1cLODUW9IaT1KwiJ0XI9T3tz
+l8jgf5kAFAR7pHInAnUcHzfStUWj8jvi/LYmQd5yZIH7Bri6EeWCJRy6v7W7X1x5pniot1AGT0L
wLcfTFaDO6dHEfAKtJtp1QHFJX/pgLyruoxX5PHT/RMmKqarap6VeUSjeC8dFF+jO7xgQKuFv8Bv
WNC6TWZZmrmYXlE7KfPiA/1Cn01WmlyAV3lApeKSNNOmHyu/ka95sWDzr8+f5+TBYvLWVqAcLSqj
Rx3BA1ETRGNs08bIvB5o/WdKgVSH8UwZz6Ey5SCTzK+QgbIcJOu77t+Ia7KpI8jnRQYZu64ZpAf9
hQl1Qrs2sJhcfgAzv62+/mY5K1gXx1LRBj/Nrl0OVd1gkhamb9MQAts3klAy3qCLav+SFnNopLXb
rmQL15HlR0nScrL74Fup4crGU4zfY9Ff8NGBD6f1xSPKdXb/wb9RZBmc9l8oDbvxtGt8HIbvhVII
pM4+CBBmzxp5PpyVCJ1JGwCUZRymBddsigun14fPqGXAJuU/K/6vNz47BjK5PZteaK+QASB7ldUY
uxADyNAU8NjFsV20fGRRmK1MxRRpNHI3IOVMDlw0W4eOdHX/Xyt/qZCxSvuB+KSOXTkqWcKVlgFv
HqvsgDex8rIXCNgr1jfdkbvsvKOzTAKk+SO4dXemsLtCXtJO+wMq7qBeJ6/gbWx4kfY9KBiJDtHF
VcwPiabZ7YTSM0d56v5SQkAmU0YbkCS5+gRmSi7ieDdAxPWkG2jMLWCL3BsIfMQAUP6MccIJCqCa
tDfYUubfDNkx6brJ07clqs1u4D9kmY0LuaKJt1oG+4g2BLBiMbRE5jg6dy5KOV1kHRCcIDfOoyc5
TJEJv21L+sHKcON/EyS/g9tjuekkxl+YiiTyklQ3CqSGg5klZ9AOvXc19UX0H/dfG6cnsqOZGW74
IbsyveavF9ljNaS0HlU9umrMdQetaCNBM7dwahnhOvfdlT7Ohkbj/RHuKbmXv3slCb6CIMJdiKMK
b6vr6HIjc0W15/fX4tW57nkcgO0t5z9+a+AvsLC8EQn2zoSkT7HafBrHUTALmOlP5zXQoIgdKaTe
dpoCelG3UV5KP/oRiz2stcEIlauzaNql2+3GebXfC99Ru4Y9n5Y25ynWVHuH7h7Ms9y1GMujn8Mk
cs4xAnHrGXwWdkNivzjYCMN6xgF9aV6Css7gCWpE1ivvrx3Y9v+1udDIbsDoGxD7P4XhJY3FITES
gs3XR6R4PQ35W0LzMpBnsIluQCm2mD7QfCubGezVYdGzYGaKJqaaNIwWr3ttLVEJ/HVyjdXYuAoF
H5x7smb6yWBxjyow6tPZIx8Ues+Am6mn6oidOT9LIEGbcFC29IwJg4TFvhB/9Win6HFiTTAWYqBd
4PUrlkf61TTMt6UV2fp6j8VsPuDETtkWB1jvnpooBoslpSyQlTVzFsS364g1bps8KCWmsLMoXZ9n
Stx7sTs8klxQMORz0eUq5WY7+HDogpr9DRW/xK96zoEN4KdAOQWQZuLwPCTIq161W+sn3+50clJH
HFNMz8UTuPx1065cIaDZMrkTjha/R5+O+dYHIcNL3EjBaF+EAGbji6GrNporA67rVw3fyrJUsiGV
B5W/TpCDYGI6Nq60do+IweLdJrtAsBEViqkkypjXEMH+Q1Dlw+8tIl3Kkt5lRZSUb6fzJrmh68HH
4khKAcyy+oID63h+9xDMr6VIKxqIXo3p616vPgY8BKVPTP85P7wu0t/BpnP7hkvKP62OeqRc5FiH
ZSxMMqKZkaa6k1kxk53WUY/skGBzZQzyPc/5x2e9l1Vqww0vy2uOG+K3ySh6i0KVET8hZjGLgKxt
wubRf44LF7rJdj+FDluF2guEAsRxVcHM2LkBSbRTovXOIiMg+F/1X9LzqW16eDe86XLnaRitHSij
gMQ9VDqrIT98CQXTc/MeFU/rQy/MkZVNxMg0fhFhVeHZfjBEQYeipx5Y4K8s0/qxIXTkgOWU21z/
j88zAw2kYuQXDGcd9gXz3LhlQ65FR28AZTNpLCw1aF92U7ux8BNwmkQlQ2KLqpVdhml+H87HcLz9
NFhZ01fPk5GEn8WHw2eHaML0NoxPg26HHao39rTV22g5RqDBPMivq1w0O6kRtcQaxRrnZWRmEI7C
k7ooc3VfcF4ZnY5JlWmmUe53lj7x6W23M09A96p5QpM+6KKXw5yv+M+nP3a4p0sWIbhpXTyfrmje
LbLNStS0cfk+jTnuPSAaPj5mf0jgnMlf8Vs4d+3Z9RiVLBshorbYqKHnfEmVhCYIBo69DT3/0iga
AQQ1rxY25uQRs7PGKheYvmC93z1RJlqSkPRw9GX+MLuQ4YSYuPMMFgz2IEABecz5FgeF5vxDN2nZ
5dEFCTy5B8XkoEI5KChNvLgYDaV4dfn69S0KuAAe2rMMkLquatHUvdP3t5YjYEtYMK4Z7jH+4ChG
TqEW8B7MMkjLji5aSjuQlcmXoh/iEvhQ4X7f6j6SAuPjLLoIgznyl45A96QxewAzfjdbsYlYUF07
8Yyc6KNKk7hqse1o/2SGnH/rawZXEiEWyxg0FQUxnFlrrYWCG5viuUVW3yCnC/l/ODLgMbWdkoKu
1DYn5/xzzsuTHrigLaZEfj6nlVjejU1Dda0i48UnVP+gBKn2fHOpK9pv7ZNrp2PGz1WiXDK2ksO9
oljzswOhJJQeLY9UqQ6WYnBIKNZOc+FjIJOXNECxcxCVy+s9j12ZkX4qLT3f5LrskB5El4MWmPbs
VLSUDMp4d1En0xj1J7gywuk7cG0bGvvR7+XMeL5VoyAgVTKpK6jbT+VynryFrpYw+PbE81rcyz7I
mGfCHc9pTTQ4lsBHCYFYMPGF6OJq7+vvgoYdUmuiwfHVXvPJ36q5W0+cUChohGoCkpE5hEi0Wyu4
V89AjwlnccYth9V5u4UurAT4rtondzpkIR8ji7qKXpor2DhDXHrrgHBH+trnHUWysHhtSvsU2ahP
QQEQnEjGpOhZdUPRJ3Kz9lSYb6+rOqukxWUcYCJbC37txG1VVaJBaYhoO+Rye3JOXlCbb8kJspx/
xz8VgUY8RIiGQi0MtEPYZyUKdL3mUZTt/WK7cRMUwFlZmHQgWgXkVTGB69V40g+kUO8usMhpvtfQ
+lghUnTa3+cN3cQJwvw3r9dmvCiHpq8o/Yus376bVMUaC3DUa4BbKkQ6JsN9CMxA8vdL6kfgxUnH
oEwLCaIDwprOYFnyAGWVl0++6hAY56k4MFkG6QDhBmhmrnUQ3jVUAtWyPs6ynKfTKIUAcsUGI7L/
yhHmbPAZA+ejGjYbSsVIi6DMugKpru5ZNo705TzdzeNIlSuWRj1MJGOWCMoC9YRY7OPKUPCmQDBX
o9ElQFHEYgdNZsvFm+bXMXUyic9LX+pzMEEu/M7sAo+mIj4ZhmRfpVpp7CrDeI96ZR/AfZRvVQy6
IqscNtWf3sC97u/5CZMwedLIdLQtZYvPXH6REOipsZZiZWa2O7cmaIzBrTIJxOLZxyhTDrOgMWEb
YTMhxuf7YZ1FNEHK21ej5Z1R+wQQxeB6Bad4p22OM3qUk1s2dyMy8iwgrTW17bJY9RqefCOJ7pd7
cmVnSDO+GT1FNpvSV1y6xteVt7g1S+0Af8FBj4DaDDydY0Jez/3bE2+Eu/msU6WyCxu8St2F2Jho
j2xc8ToRM6C++xLJ/jKoqeVCGaIU/yjzhEoTekkW82z57Nr4j3pzHSdtXzjFN0XK9lvLRb71RU3e
1QFFSQQ4yqZVvB9avTukCKZl+tjnjD411aijgZr6mtGye6ZNAk7+v/VFKV7TaZm7Yc452CcmAU+H
55AC6JFyA2wlZaMolZ9zQMWE8lkcow5zsH25IGaT/Eiz53+Le17xHTm4isa+yuac8ItHS7IwfRso
Mlfb/NIV8uZc2qpUtuNR6oWjmIu0xaQn0UpPX8OzhkIYRXfnq5f1lGEje6NwhtZOmcxp4SEU3glZ
mOyG5AY+0ZWOVbyxlu03pYiMEQXUjB0Y+AFVwID4knp1umHzmcpfMuiChfC+cYi9qoLGf2Xcb/1Q
ShYqzJr7mTRU5EpWrr9BwcIz2vu4TD3RmcYasbO2eVeiXe8Xh19v7q7AqAGkKT7zj77cwcoU9gU0
wWvwpjRcdnZ79q+hsmpLoWg6AC+ZpPsB6SbbD4kpXdfIPOfHLXyLm6hNc+I4pXuUtEa5XTEaFr7O
0fILosB2Q4EP7QYFRED54i22gr4k/W8iEDW20/KdhdEvi7Pft6KPazjx7/NONNI1DdTrTPHvxxPY
7x6ZUybvO5mZFTIxi8ABdyM4dcR5m3CCtgXRv+z0/OZxn/jU/0b3L8DiVN4oPHHWzi+jdRimZoXP
oFPEdTelcAnZdYtCP+JdE9h3u9NFf232bzBysZ64LTRI9GhPcMNSrlnQeJivAkJm0bOKb4moiSEz
Lm5y9E2L2zT1OyW/0oIzEpwSIq+vWaeSHavCvSi1Bf2RabNuxOzGKItLY4sUzwRTltoouttpsQ+h
FPChMO894cTyZZDMts4rHvJ24tKOlrLbAaiMVRmFeEBzFIo+zwW8RYT17BWR3pXmO9n8aXXeb0aC
IPHJlFIxNnMwmjUpNnwOgN9x4fP5rayR4GWx+d/MJsUaC8Q9Ih/YAOeydzLHUyKbCZtlovPODPY6
2jMIJ5MbMC6fuymveSFioDorLcOQAAutucJLvvrXcsX1nIHNfQJpEChy90/DsOySK5GmCTGe91S5
P2HJogxIwEDhDnhtW3iQd2qlZrEOS1aW5M0FUBPXv9KhEbVhwwBd8EXHFWSYbsH5PsbXkbBFPcgr
V429tTlqCmLPgfjKcjW1v1+mXZakYznGTat7VOOJOWD97C7VDt3TXsZ0L5NAFrj5Kvnp48lgRzpu
QMoquaj9lMHAoL3PM6FOBp3gqcqtCm9obnbBpUOAIJDvjd9tKSUoxSNNePRSNXfA6gQPS2YS+Q0+
Os0ecUcXXOJ5MiywVCC+HfYw2rgKzZ85Zy7Ub6tsaADUEtA905wMPayb9CQpm0Ir/OJD1Ljr+CEh
/ghGtH81FKqGYJBF87ruif79untIng+i+NbwcoQ1XAv4pSzws1ZGBvwaaDR8ByzrV7oHvSyYslDS
5KBO6/lK29+YYNtyQsxY6fvT8WUs1WxLV1iKWcTEwjAM/+UWq4l3u7DIzS2VeK7gmVzAuzdSHxJ0
CEqtlytZ25hI1mV/YhEAu07dszi6ETse6Bf7BTW0MuiyprfPFIfe19QQsUy4x8As0fXOTsCkfuXA
meNSCQUSnbQLa1MBGUFq2/SIQrU90ECLBmewZ1vSTiM6LIYuvdE/jHPLYPRvt6l+oxS9KWGWfeGW
JO/45rnhWBcJp8haDMplQwdNETcJSmuzTQMXRQTcvQrkNckIfbzmJkTm6zhhrPRPqc1WfQa76fri
noS4VwXL5efBGgrMpN3UvCBrZaA0nxH5yi6xNhSWmepQxjqY0zuUgAlXqgm/1+E5dA7JL+oMFQSs
DV1GvDpEHSY6x3TE3h0V/oHP6bMbKTZ9lw9a1BKi/X3B527WkfYY9u7saz+lDyckNWmThcwt+VFf
osI9F3LntB6dw0HghuwhWBDoAos0z5tDjyBd88Di7qTXxeMNwHTDw9V3/R0r3kXARrrSvgF8lvNa
A1fjcwUUJjlIxI6WiNmMUpg/a2H65IHAoVFihjnrblzmprUhEAEMR+8v34gRKZ0+EuPQEJP7gcFE
CamhHOOjZnbFmUjWf7/X/Hz0gCHGYv0cFvjzqLFsDu/nmZ/22n8bYhZ4+N/v4ehIRVlFbb5CqMwe
sXnOLTyl7HA9YW5WysTrT4fnUUMgJwPe+1juGzgunSRcrQVshnnH/EJ2gUO2jRosngJnJY5bXKqC
cWrBAs2FzAxd3umN1OjdsVfOfzy+8GY5e5vZzXXi62cLxorHzt8mG2cEm6LpSns7jXF750YCN5pd
WgQtuUv3oA2AIth/DOVTIcJBe5fLeFiad9IU8FG1ASxzaS5zq4PDOW+8uzGAT7FCLDqZQRWLHcsY
Gq+yN8JPyBZ8ZWNPfNHmYtHcaTdYcTyoxw5HcCYacq77dKmiZ6IYcxEEvbr8PvGSILJlPEFMT9k5
JoGAskDwTB4FikyVXMSVwQLsqmEvHIV3psw3zrGEKSF+w3SVfvvMwXXMq3PndG8r8JfittBkz1LK
YDKB7nrC5gJ6dRod8ZfYhYTzQ6eC1AJG1eM+gNjF8FNFEyVfvnkm0Fssdr/rFNsF44zuDlcL1WeV
3x6lPZiVwv4zIDvUJQz4TdXCTQwrk/3A87u+9JBy3YDredOFuFICZ7kx82D9/K/QjAIA6JBhb6eQ
U+mLgL3+6VrWTNEcffo9cFkxOWkv/J3Uox2spkP5WE/Rp1YyV/M1stAlYzVBwep262mBLGdPlDYQ
ChKneqUSedXNu8KuCrJgpOJ3epctpPKusaysDXZWjr7lPDrFv/8RoWB28EmjBmcvM2MjhLGLMj5l
9BpVh9gCsckyAaHH4XFl8EZyuULtc1S1UgChl+TLuiMjtnMqT1CpL3scYQtx7/PGzBme3uhFfyHb
binqVWobiNepE4QOG6nW/EQ0xZ4x/qvG2fvf1F0qAQYbyKl44qEs2bhq7/zsbr+RiN0MRldb7evS
bGML/+d0RdyRcwtCZSh0Sr70f4V4RhPXkOYpf2YGepDVZyVfp8kKXxQrcEzi+fcvD+huGsNxnrOa
FpFkuRqHT7co8Gkj58Y+Zw4wd1s4ygvvAGRr9nwjQ95i7RtxVRJM/n6YYc8kWhfSO2waBtNAv0XR
9larj9o3VHeJBObtbt5yAxY62CkeRVTBUR5FblPsCKToJMr8Am+VdtMH4RKGB1xEgsCeSujKSBFR
WOXoUXI3jTtc/m7tbWFmQqAxbWxq4oDUBg8oaKK+srCchH7dsupsuyNRFQ39YUnFkK8JqXI/y4Mr
k+iUJY5sgLi7uzWhWQeAD2E08kPh4ZEFIxLzD+hTCcXlc6EpruCvD8aiBK7dS7OSjVLbUKipZxPl
lCWus/u2KHTqPsZ5y9RQEhMm8v4MZbEVWPLW7Ebo9p2LznS+2EGVwhMp6zg6SHvh/Iah04wUlG2i
WA8BMnuf18uWILNRZnSzIavjqJ4fuD5OfstL3GZuYM8JjHXZlxt/LmkVbpFQkUHJp7WAhiAr3KuD
t/YSXu1Vb+ae4COgklXF6PPJvVa1q80wiWa4fyszHG+jJG5JCEmS+LlTcByJAjunb7k9CxDadTI0
ywUf2FnAMbl+6ErI7PHwA1WkYpTkcBEWuIuEPd5OQW8+QcxoWlxhm5zk/MaQJw3Gd5e+GU1d/eba
Lwira2Ie9byEbnZbvEsjsiWUqv4x9ajNPBPa9EN4virIGb+G8DI31qg3oVIaOWC12XKkmre9CROP
muX22colHWwgzaWYQaRSJfRpqibJQVKUF5LmVRRcXP0navinfeD0YIkiO7SRhXCW7HhvNVokoMfG
TFX0W852B4UDiBDsdpOzpprgqiTpmcvmWBOkyEqzw9K1UwSq26Ubp9dvBdRHAnchMw7UtEAD4nrh
9EpS/qTFAQDUq0gf7+j1x9F6yTE1xnxeZSfDy7pKwanJBDWQrK71c2eNzisc1SXeMxu3cGjPlZvJ
RlkA8EOZDzVT1v6f9MvABVDGIIivWVZqZv1xacXaHPXBEyzc/SbuKdZM9RN+fcX/Kqd867yHjfVl
ws/TZDIwa/sv7TH2kJWhOF0dO0RLpp0V8eRvlJUoCMa3SwlkYHrL5oA37+x1mvmkCKAXncfhWsht
Iwa7b6aLaCWXTwekvjNAd+xFyiIMuCs2WhDbeqkA4BduyWlZ5J2s/DvPhHrJN7UGrWMrZz2v6jY3
l5vi2LWtkAmz1OwmNMAwe35eELxETkHJtdD2WviVc/DUKttYFNmA7h1907CyZkqZxY/kDxqQRL0d
+JgIrwOoUFsHJljFz4LqywwkgZYLpNcDjPYG3vQieJHinjXTJdG7I+A7Kx2ZqLzjGlY2akaxUIfJ
SVaJE0DLzwpTXX2x/5NNSPN5wDZnhiWupg6t+xQNtts0mWvQCnq6fVdWDqyAXSQHT+OG24zNi5bx
uHYhm4Ftl1vOD/gniAr/KpEFLqjvjDeCAl9B4d6CpJjDq7k5eDH0V8HIzccWvAwWULQa7dxvKC2c
Lb5AxMLiP2n7KzC1FZTpCfMSUUyWH0jtloHeu4TV7jWu5G2Cl8K3DcEnWtnLf3zTsIJD3VIocahh
kn6ZXIbd4do/nrPteaWkbxNY/O27viZMukJoqmqlC4g3NPoLZ6Q2C6LCQn9IJ6VzfGn2qKEvn+FA
tVyC30++7o1c3c4ZANgS6PFsrp/qMdCGRR1eGMiyE0yX7PJoT7/zVzvtSLVzfUbGnBHKbP7f8ybs
R9/gsWl8sE+WnBbY+qCPEncF6LJVE7jpQp5ML2xUmx1+7Fm89I5/lee5DxcHtx009BNUtsrHVHjy
aw/rcokYCPBXvKSITrC65R74QpLWaiDVkUxjl0ofzlAa+gM9ofUikeMZcIK+//0PZ8RHdzrD2Vm+
JSsMx9gOZ4Gc+gCI6pRUx5QWLrXN4fozVMh1jsOzfUiG+VPFELMutT0OKA/bQ+i764P4DURnFZ55
I2Rfuw3au15yG5+U4wjLE6r8A320dCbMPhr2Vo8AE3FiBwDm+lqr4FayxoWe6vQZcKYqjBDUNFIk
L4XGGpwkWJF3RlatZNMh8opBRdufZTRtXwm7T3hM4CHmstTkGqklH7+vX7F282kAIxawhoG4/9/f
ABBoNyn7ODg60CNPqkYlT5FdK+32o5R5IBBQE2qqEbJcyYieDLzjkA5bftKJRnAbEtYmdT6I76KN
biaD+CboJ8QevDN3p9pwr5O3BvmWAstAWAV6sPeRBkBzyjFW8azyXwVFgOCxB2l966Ir9Ppw4MfS
U6CnfpK5Vp/6s8/tvqeNqXhyhP1NjvAzQJMb6mWr7k0QHYjGtzj562u0LxYDwPbMdzi24EdG21Qt
0IGkfktp7s7g8honpLaJKEvIzVfpkX7NSfoa/0h1d7hvdS3EzO2oMFY/7mZfEXo6Egq8Gf3o3G1p
hnuB9jn1VRyZ6eci3RNgjKe9I+KvclCY00rdVESj8QWwWJPzBlyOmXNm6KaElzN8H1kuahgVhmZL
JSWs5qgiZo5bxbRlFG4TuTy6qUxuCdMf7BCRFFaiHa8GT4aSN4C33oexczmnXWU0mojYnoilyUMN
wXldpO9cX207+n1YZbjIaOF9oNLR2HnxYEDsyC+R/YIAqpKtCKaE6/yGBI6him7oqJJp51sTT5iu
/stusl6QvPTJ7LPtN30P9KqfDHcSGkxAJjjETYP69cjF1AvMaRrra2FX5uSsojcug1kmBw7XEo4q
IcDuNDlXr3s5aMwTaQ5evNk3G+eWeiD2CANlMSkuHzuKI3z2/wwqgjwP3A7CI1MTIMzBWSdJ6doz
uMb2bxj9zzyJmO0pZ1dMR35R+PWaCTfTQmYA5uj3hXA7bKZqS3JcmdqAU2g3UuEHCj/iSVA32dM6
NYQPLksy+o2KDNMbsI1aAOHOD/DElMmVCbXn+NyTq6xQuuKQ2840jhnexU+r4KVIOAYe74EVBZEP
pO5jwwaef7T/WAuytmodDQstkkR6CqHtjZUeT49k06GAy4yMmuEXYkbYWNHrjKCvRp/nE8Zy8YZ0
KJFswaTJz88Kjw0i/tlQbmBTzN5ULcB3v9cWa6gfmB33SPajKrkwLOHYa/vsSgjdR7rsmYQcan8e
LsJ0dNRwx5WrUroxlaXpo0F0kGs0XR77KXB6hPF417nvr7Dc9xEhpZ8BcpnoMj/cOiieORRRshto
EU1scsT6/bctZBRqOaqtobo8bEH1YVXikaWYsrkrr4EYOEGcchvLdt4hYQpTTpVnDZ6KyqUkP9TB
7a3+LWa7o9ITff63HeCaZQq5vyLLTL9tSoiTN28EHrko/wkDj8RPNqAU4cevEaxgGLQfo+KbqBEm
41H4HF1IBEtnwKeOVatuotXTYZ6yTb/6TqrePg9GktHBhFBsQLmKnuRvRRnlDMnO01vZeDOk+WNE
j57O0xPsloaUV7S4Ogoo6vOpBEak9Laz2mZWMr6Vk7jP5jn+INR9C7GWaPEfP8HAEAUbjlwsPXS6
PmnXEtGEkCzVztFkieUEsnY28hO8yzoENbsUMDhmkCpn/xEA2ouNp3dc4xanqqf5kjBZ0gwy2EjN
VOS/9Y6cVkuP9MUTLuq5ib+xIlADR/LBQN+f5UosC6JNiBvMDDBnlUGPcNlMTeaI8gp5SqP36UBp
9hfMk1fvLK3KZHxu4aK4g1MZCGvF080ASdm4+wtsMutVBxDRq9p/EiSFg0UrQ07XeumlSJyXoLob
XmiFzLSInE7zHNAtDZtnhn9Gu6bnY/JY22NN+Wd44VgmSk0COlmmMpQ0lRS07WFyJUAChtEs0KGq
rZIQ6pzJRr5GVgaVGsE4uXWOiHal+GzcKVSPfoRcOFbOOGYktR/sZuQ2Qcsgv60BkZmRh6IQ6R1r
7Bw8JClZ/AevlMkuzjDCtmbcfbKFDa0pyI1RFx1N1sWNSvglleyazO2JN/vxYVbZfhYQYJFJD/5C
0j5IiuXsBrZhB4xeJhWvz38SMqunpgmxcoW9J4dXt8g2uTUCQjFp/aPqtuonzStg7xqVWlnFmlD9
Be0uo0f8JRG6fNgPh3U24QJdKuvGIIrIaUbDe+moGXGRSyNX8jFaZ8M3Of3yWUqzFQhxAu5Xq8nY
VQoKeB2m7I/exS3akYroSx2lPOubB0VwwnInE5aolbbKJ5J+yvINzQgzUPnoX5/2OxcGJDp24ZfO
tYt2mUGhxTiLGcCzSBbVPmbhfjeMK0ep4zu0+wSQa9qOsSDgntjB2Bx5Y9pEdbJWyKY7lbgDQAGv
2M+Wil6wPeaetzunTI3gGnPuHFWR/MP4eh9NP5vRZFESqW74L0hy6lcH2QtXXYnaJcoq6+sDyZJ3
Tpe+py59pEh7WofAz6CHqmAEXJwN/ObBNO7Kxt8L+EFXbESATFNLNi/uqGwAb9I0OuyHQUCFqgjh
NSCvUypLWoZjWBzxpaUVBcE8gsKQQCp3SsHQluI0rz9nJzpV8CzhDQXIG4CWQBEwbKKWVXLesTor
npRbGl+fnAEmyElhtK2VDVdqb+QRjQ6npPDnxkJmCKKyRyNNWRHP5Us1LFTYXMRiMCNSmouDfGEf
0Jdjo3i+RWD2PxbZ+DERsPRjNpNWw9qK9mgMjgtj5tfTDWW1LTMeU8BYLyBOTT5VxHDF4Iy43lRS
uimshBjpeAX/Fn1k4RxAdxmJVJHXKOOpy8g3WmQw4Zl09IZI7dO3KXV5gsn7Ja15AXSvbJIIs5ca
sTxD6+TJ2/fGCtFCY0kwJW0gLN3CPwmgW1oQbskqbYORfQ2zvuTgpWf8Fl3BKDXDQoLoidoTwuRL
TiFQ8nrx0g5Oe2JQGfmpk5M9yCPjmkbYyZojzSPpSG8u7Ij3xtO4CB2ARqyIm7+UdxtmjVe7qBqv
JiYk7LCNupg7KYlAiqhxxMvp/gSLsIcJVT0rW4vwsR64YvAzOZi/UAlvlS2EnGORKf5gRhOZtQq+
rFds7/8HYOmLQSYX8b9I/r5I/LCvXRs+yXBGWhceSFrLUXCc6i3rFr6Gu63To9p7ofCLxGCP7RFU
PshD9O7OCt6hDN63IvWxHBRdO6DTKBEL5esMXrjxo2ZwEvoo8uJxUpzD1w0ZYhYeEJBHwZcubkpO
7VH40N0LUz8Tzn9pSkmJKXzqaxipcdztCrDG0rGJGxz2mpybOAxLfEdBabyPpBlaX7AaOB3pHFsF
cm86zitG9cQGPvqAzV73LvpH+62vM8PCqS8pp+VMsu1nmZSjTdapAzN7cChM4GYyHGWDA/vmdgw5
7Ucf3PdxPSqmxpURm4TSGQpacM1few0IfgA9A0i74gk4w6c+eQAjLJv/+gnBi0Yhmd1P8GXSdtFK
pMQgqzu6jrUwTS4h8yuMXtHbQFLIBFLsX3Az2GVc86aUdzGRsCq2To261tpKqO4c0/k9sqvZ2qMF
LaDg5LNWfjPtt3oTpdQ4mX4bXIM2NblRTl0mLfv6+KZvCeoK7ic4HS5S3gSTFbgxTBlwaZI3Zb3T
NnFl0ij8rmdElL10icCYlxsBO+NS4M1ia4s1L4TITpn/Gm1vOzIbzYqx/ilphwgHu8KHqMR/2kRh
JDo3SO7q6m7Yp6NxMjThsKDcUWzQqXvOrOc2ZqhMq3isJMrkNVP16i6B0owSmQ/uA2aXFWcXp0SR
XjBUxxo0iSvzHFsTnfy0Pc4zFt5nBbIsns3kUzHoXEn4ptzBSJTRt2B8ME6d0JsLf+Lt8oYBV4CS
GG4EYT/Gw6Eo3ZAQYqVSBKVPLtmCxj2kcCeYPQ+XcwkN/QNADGwZUxKmnglqStYRkmZSaZ8WafPm
qPB/SKr0kxTDVhvm3eGUFHO3WzYwPmmw9EkMiUobXOfcSZlSSmACWmYBdXOkiIL9P030UmzjKnvL
3rTz5i3ma6vu3OSQ5tYDlnoQIbHMNo5gEJ1FNwHLXnarqg4/cbksxA9BpHpyWKzj2Ekl2g7C7WdP
TH5SpcwYDG3W0PDm4FrxSAleBTUBMB0inX2E9b7jny92JDAOz/kAPhOpqmHlNT0KruUm4Y3JZzdg
+eDkr5UASKD7oIPqfRx8UUMDJYLNvbkbwktR8ei7TFCxPGxlB65woNT5wziOqtr70CegPGRSUmb8
+jerpFneh2f4BG6O/Fi9mVQ1NkHPRjMkVxgDICgcUQeLXRZozzdMm6OADe+9wFyy4W2fnFeZl3m5
TDA96sjAun8JexqpLzXu2jSmcxnS/TSzYro//fSUBOpbFsqG+kxwAkp702mnbeorD/uoFPbeHbSx
g6rWVLfZZ55khXSvxFSaDuQERpI2YrP2SFr0QZHPporRzt9eYtdaWYcoAtVREdfTHMg3HoDXW8Jm
rcvvofbnSyZp0olj2e2ta2+1kH5O9YiJ/q/7GFv3YCP+dcDbJwkjCd0neULZQW6rUhxg8dcDiHag
thQuLqSGAji/n2aCPd4Myjx6zzn1zHDClXnGEoORo1/hR+kKzKlV5/sXDVSYrk5qPIlfU0lqpKeP
p9nNCva8V6dAO1tvEFadKz1tprcjJtGGG0prNCeAq1Zr/7NpfYhnUusdjkiOp1DmLjGRo3prHJ3g
PjccBjR/x9yf/yToQfc6vA21NBnEQtxx8auT6DKT6opMRayzum4sB8QmYbbXGyrbFa3OnB7Kmll/
nl+NyljGKCtxDKOoiEi32/4IcUmc/p/B8QHeyPMxhlRRQA8gAjuk1ES4RY04/gSs+DVlY9zMns6u
k6KL/VpORAu463dz7iSB2u4tZfD0tGmAanToslGV7ld09bDqDR1314Gct71xGMypMnxdG0FZPdwN
jLeEgwVqr+LJvIokQ7HBy9xl+j4Hfhz3nY7qJvyWdZdSOD3MgLtOdD3iAKiYAUIU5BcaozsgceRw
MeZdDvKGoT8HIHihrCKW+mOxokumDJG3U7f8Q+bkp+c0Gj6fhkkrx6LPjANdEFL1okh6AgTA/WE6
CUHZJBISXVLbosBwFfeXnZQ2C98xw3XkfDESRgNVGdADuOA5bM9GHS2NxNQH0dRVD+gnw+Dl1fSh
btlro1hcfqQuLRDxGJ6jX3VawxTIAgnSjjd6pj+TCtqS80KWQAVpexqaIq63CvVUDCXf4KIB2Qzq
WBqUuMpc2XxrVDeTrrIL1wBGko3eCBBqWCWq9X8CJ3sxVtJkcnmWlv3lRAzMybykj0jltoGMNJZ4
1AJh6YhQWrm3NLGPSoUxhEui1QKqEobL3L1Qg4/vNaj5WA/hNaf/Urek2rUKHJ4IY/9CS4pnSgyO
PuG5NrfkNlguMhqr7ToHVn3BmMjI2UACj1jbVYfSE1YHvqsYG/cqG+03FdSuT2Hr2cHhjcpDmzJf
oZIFXnsRA4YtrFnV6bafcd4yLexw2J2pM88sir/tRV8MdMTNInLz9Xg3BDKe3xtOfmzIf2/mGsYr
yppVWwz5aGVMDk86MaGKGCaQKVf7q8f81Z3BkxicnQPpX2cMvd7Mg/5mwu+DkF4HIKQgNWDq/qZT
ij0dJzSxPtiRnfNEpgkyVZc8MduIq0v8qGykcLxihXynBT/2dGQrCnQH7b5Q297qzIPseZv3jluS
Mhott8g3NkrKXihKJSmB4PHWWbnXzMIKC18yypezkR565e0w+zs43RJLSNWx91GpDPczdX4L2r/L
msIGV6ffm4WoxBqu1lcCKXusKJuE9TzEZm2ERFbml4c4xI8LFSz0+ltvniWvC8knmMQjUH1JSH3I
nUC5Rn0F3rO2S+M2CFlfqlka4VNltwPR8P3L3Lfx0o+8+5OGnMsHRujOGTG/gSyb9oyFmqSQBndS
lZ2yx1SyEGZvhnEqrCSXRFyck5rOQTnTjggaV901kL8BAMUPuh7k9olljh/e6wOfPxh+K5/gDSfw
/1ZAtUUhulS8/5eLiftxCrFSNmPi1vpV8jAG8rp8x3WjwLFMc6J2UzSpZue8EV6R0HE0LLML8OBB
gPaEjic/hB6eR3T248aqMPHUov00189cjji3SFODrVelJ3cT0tzFneT0oHHPPiSnZYD4wYI5D7kg
t/SgCCH+V+YETp6hDEpgGyZI8CC7orF53lyWaiWz2JRGXB3b9iwyxqdr6SBqrKRLZBpqZkBAOSrk
I1nCrOAmmRvbFsZIbK7R52fDdguk9+HlP2mMPZtdWoBkPjj2DLziRNupF0Bp1Dr3Q50A10aha1fG
rJbNCGyccWKOvtkUMPUnTsy7YxW3W2xfv5Xq0vUEZt+/yOWmv+rRMNslkWYPGts5At6aj0BVqcNa
uH89hEr6iOsIpCZp//J58FmFA0LaN5EQGMtsTbpcbtUGnRjmio/X2nqaGD/OuGJgXRYV3GZ1379e
PnhOWz+Q+hk5FnoytUm5fisRD5qNcjJDEx4dpmNojjlvdz1U4TN8Xkz/ZIqiOg+3yCYb3CyCE1cc
Jpd4Yze7ohMbSdAPqhXiYX++WNMidJ2aTtPaBCp/cUF/gR0DIxynG1XrbsVKNYnGqYRO+TlnNQy5
kvrK+ifUa3vkHxasHGGK4igUDf8111vXdDi27bcmqhra0r4m9HQS/Xn/y7sepzN40agVPUzbEccT
l9mLPQt8oI/YtJ7BZnHJ5BqS11wJ+Wx+RFeNZ3xkpzn+PcHS0YrCkOb0SzztdJ0yJx3MGQwoPdFG
JWTu6QT+aju3wvnC4vkIFD9uB0JpBVE2PzV31kyUBSXI3XCZwvvlzLph6favIOL3OklO6U8FmVVl
AI0SvIyxYY3KwoOwXRnNEi6uJwU/gd2r+O8nOmCWYTiPBtiDk4I/8YLTn6wZGh6fTGRDobhZoF4i
Vh9h9SFLwJPxIeFqXmz07JRa7BF7mc6rqZJERpCiSDLmCfEIs6JpuO+bzZPWA9MctOeqQMCQ0lW5
V/gVniw9eixg6ro3dIOzz5ewEeZlFAVcRisFvo4pDiNeO+w9Kb2/ajCX2FJSVzOXrrNGYYl2FLAN
+nY5qNsE1+Bk0Vo963WSJWXuCEpz/xvQrOroqJu/6pwjHmZ6gWQAS+GxAEx8Su0w2d4lpmkO+gO/
4wo50WpgPObTO4uxVq3NBnsAqJ3hu7j765ZImTOexSdj5VKgdOu0DZ+7LOsyG9MbjTM5+DFe/8BU
5vaL3HoHtneqdjzlWU8OwagiwCfp8B/mLXlJ7YEP/YZs90M/Y0h+3zPyOltZ/ujFg/4vqzWhiC7O
wS40W/6H7EvcFjw+mWBxxVmGCYIcNNPSb7eCl4vrSerTARsBOX/ADMNgnAmjKU1ptWmTQsscwVNW
96J88w33XE+Drfwm/WljdLkoiEPKP6b6lA6RZPCggweTH5tkBeZWNVwK6bB/WFfS/GAk68vNImp9
5eSmKWEZbB3fDEbPyQxxkyG/4x+7PXgVUn5tKDma53zW18AqpfLgaJGoxy4LC4h6YfxN2af9XQpX
R8qNL+pR29WpSY1cbQSykcMJOqeQFe3MnRfAQJRmjV2GzW+EBaHrLX/rjsr9rHkB9Jy2t2UQEB07
lBbHxPuqboPrypel8Pi4rq3zlHzUN9XYW6V8EmoTwQrj8U/1NK5LBdPwOBcQVW7fjYS6RGg9X9ZZ
0uzq/nIim2XHhqeN5/+975ifGwFwijZIPsDK5A167fQhCb1GLsQ2mmYoHwOnosO8w4dlQ+FCAXsy
AnY39TKJN7nE9BL7lTFOnCCRGyotJ3bxF0rJZTR3GOKTuJsSaqrub7MD6hUu4Jo/XDYLTa2uqeGD
pTCx14qKYHEBYlJeBMcfJKsR9j8c2tf1NfQ7yC8DNXa/AT2m4Ou/oR6g/CfwfI2JYBriQFZOf7Un
/cSoHQ1iWTGAhtfplEJbLjrBAmoqG8UbRDvjn+Mw8MBWTgn2jZiv9QbA9QWf7pa9wJpziFt2COzC
2eTE5PomJ8euALvhwWRuwqVFE4HqgWl5MMX+GM9pvnxjJjwSIKJUlo+g17lwHi+7tKOEVZrvAl2g
q4A4rK9U/I1y8CfQ4ahNVNA0jtVOw71JxlXLarE6OaIz+k09ywccHn7IPcCkRDJPrcKe7Lt7Bt9k
5jQeeu8BWhwyUVi2ERatnaLdOcqSVZk7NZZq/qgD+NcM9d6qEkwFWdK2POtfk8IYB8RNwv/cToIX
aS71gdnpR3qfoba+MXh/NXi2C3exRDw27CFQhwfgpk6tUNZrs9IgOEByJJqbn47Svm9RBLxDuafv
d8epOYS7xp9s1n/cmPLt//A3tbNg9RAQ7FbhqgTgli8aAuxUz8oTkvOQSDZeeoXPgS4uN7Vpm7DC
PPGaC9izxbYHS6nQbiT/HUqnkGK8XDt6jRA7kDB3XDlSnGp0e3+DRD1EJNOM7votslEHOk6kVEyc
vjf8nK6P2xkLzw4iOB6AsmgdAO/Kl8VjJinQjhYkDOi3rXFMMBF2rsGKzrfM5VfLBDbjouz2j9Fm
08F8Q3/DfHFDjv5esq7g90xpcqDbXu3rsrmgW62LXMsK6mCE+Khm4xO+7d21sIhgF0V/wTnpDGtK
Dc1WCZuz0N+7i6iXi47lNbjdkN0fo29b6zh/Dl8CnihWPIuDBBBWbot/kNKhYd8ufXre9++YewT2
62DXMh8dDCyLW1I4jqEV+h1fx/IsOXMdpXP7L89+tTblA9w+yVlOePmNOo7z6zZaJaKC4FyaCfmC
yrIbyPlerw/G+UK9e0zi4D+EFNpDpOYgM46QmECNlyhFmDMQiaqBegN7JagupdM/V4ExTOXdoA6I
gWQEgNkMhnLEezRBGE135KwknV43uXOQZq1UnNgOakzeF74oBXaLkpwZjeGVp9pUU8RWkLKTTsIv
DpsmtUqGPeSO8oyZ8HEQ1BxGT7iyCVlYgPDIozQVGqSzipoxlOjoN2YX1lpCJArwBGdQdxuKCCnK
/sKu0PWhFolgNI8W2qm0W7C5USRkKv/awP8kGsj2qsRQPx66aAFLGlUY5G8apWLK3K4an505amTh
mcg2epFQOTh6E42LXqWqguEG+BDZ3PsTahWmuDdO4RE6xl3V7hlAmXh9/tsa1SZ3dGlcrFo6bsRG
zUdH8yg6SHjzUEFKyekyhQHWBz7ed2zDdFhyzx0JZUVdsM94vgTB0jG8UCSx3U6+aViSXOShx0dV
bwxBVhBsgPYGwPkrBe2qnFLR22CG92JBSKmFOW8LXukWz09g39u4f3Ar3+djAKVXIb0sytn5g1pr
Zy5E3v1qYMBzPK/B0SQJxenTHJfqyT2iXg0VQKw+a+COGkCm7+g9Ns3c2yXBXlUxcewvXyMey62X
Xr49/2y4q2Lz2PLBEaiafEdL9mWP9E6GxoG5n6b/hSEo316wApS2E2n+yBrTTuPWgBYXdUmCYUMY
7V4QWP3htbId8YGlZr0KJP+EayG54/ePjT2svXk5NLkU/kiUtHsv20mLCwnpYyjkMp/6opTctDhV
B+EU/e35BGSGMTEDW0U1uW2lpHJzN7T4Zl1FmHpNvDIUR3DhvXD/RfmCUTj5bYz8nFzBd3VdE63k
u62er+LYqewziCmVMou/NFqMwrej1q9mw+/m5Vd0fCw8f65tAHDh4woZTFblPaqIcG+KtcRz/i9p
jcK1ACAIqR9gxcwCtxtzm4jrySyRS/wdG7ysd6tILqBsQjFSLHwwzcnr2vzMcZA2BlsA+B6TwDlQ
LhmOmWWb9yBvdA3J+g1fgau+v/q4Gt+aOs+vSGTiiccYJeAzWkd1Bf+gkpGwWNwTswlow/l1EigF
tLYEO6udurmTIbDf9HgWWClC6+8n2wpynLfep/459IiqwE1P3TShdroc8mW9akJkb7A6ocraEIDF
xYwC3sQh7fEj61kmjPh9rN/u74efijAsZ+zK58JaoaKkcErMOCcfEgWWE01Lodvk7qQshw33I1nl
g8etTzzEmSEzp/c53xTyuaAzh6wPbgeHHj3dpN85rjWOpkZRhn5VvyH9QV9AKJJi+VA8tNjzG5mE
RqbeOcCNaGMHbSBliC/TYll1L+pquiZpamHAxr5B0/DfduZRVGLloD4M6k0dvJ4bZro2qh4MhxJO
cDAvUr8oMqdqePw+NaeeiZPi473nOppLpI2HMxs/EDVnrB0f2vLh7ry8ofIOwdZprmhsCKWNfFAA
ohTo1fvAX4u9GajMZhl6KoQPePdYMxkaXW7raFRrS+3QGOc8jbh2KS5nZFmQ9nd21Z6T9gU0qsfv
LfiBpcWlDPZ/JMFdwIPBFTtgLoozLX2bbozhBfojUmS3c+8aalx7oU7Xf4gReZP89VlKBvo7mV0u
X7gYTnuAyTgsZyLPlkzaF5unsi35kt4Y5d8x5pHgJaHWNZbd2vM9+OFUwlw3zwl2/chLWU0V2rlo
xaXRTvaw64FhLCpMrIvowhy96v1LimpNjOas0qdPHHlKJHjdaGM3qI6YhZP2lVeCtRoVD6S2m6iA
sKkmZAayGZxfml8c91ZLP5+K7z5bbC19OLCAvZOostYGSgH+Ng47Q7nipB+JDHc1B3H06oowTesV
WPd0shJRES/eRJS9z5ihKOSPpco/wxL3r/F1KPlVr1HTHn2BNYWkVTKY+479OE3ufjiqul8Qc6Oh
PrnVhHPyBfZME1fBM/pY8/dfBEOAMHnPGgNVgW0XtXQy4PVLA7oRrufAFSf8nc4Z2Yt4592V8eU5
qaeGtKEVirzephsk//rfi60yuaBpR10bFrxbyQ5DIg/mI/8FtzsUr4amqjTnhO3lf1g7hM1Gql1C
lS5y6+KlIsrGRCGZ4WqqI2ynXoHbOgXes7IN/qZXxY5DKwhWjepVuLKblqO/3GIM1uDdLDhVLIVU
3EZ4YrwNzV3otHe6OG6C7FokOJ97Pj0G03/e5RIKFQfG1rB3m7F6BCSllucg2uyPhX26fAsTBptg
kUQpBWL5qM7rugTBH8y32x3Kh45BgEggjtm2NFk3L20mvf0iOhJM7TaYu7fMc1Ds+ft+qmmLuKh7
F1KfpIcBH5t/gpU2p+qPcfwgnjDMMHVYmIu6hJ8lfvvBoELg5tkBsdSC5wZSeC5BZJcn12p0R5KG
VglT2tPNWPPHP8CWfa7Q7zNu0BjThSupKVR+ZIj4R6tGKvn0qehnljZSKp7LmPu2Sf6VFfYc4ig6
8MfMh1pIt1t/fK2ZNhR8ITeYsHix0TR5DiNtmopEbD0Ze4suGHGeSuGlaqwvpWVWvsmEBE2U7xde
LG1arimugHcQy/BzkPSz8+f1MdEXbOPlkYQVFsBsRJy0z0SSfAroxMMol1XP1i1MdWv6Y0y6NLXj
FFLWtbx05YFw1hQhQkWwoeve1zjMNc17Rhxc721oS2l4FRe6Jtvo0kl77FgEyaOyghxMiTnzEBHg
awikyJEPk/nqufd+dpZGdE8rWWU4DHh7dCRzp+KzFfaKLv22Di96HQQRttVeoWZGRVES/7TXQ6A+
+CFpVUVrmQeTS7/JnOJh+X/YcbzscBc3zGF+s9/5gwpjYtoC5i5mezoPD6v8ez/AAbMp6fVjRX9u
15mIJf+kH1OghHKK1St0IkFOGpT5pn6fUW9RFI1KybXGHDq1rn6PABT8+AVLekeM23rrqwnp2Rxf
ifRksWuwbVeszfYndVbzJzT01YwsGsy1SfiGZY+i6QRJ1DEdgKMPIb18qR9piZd5ttf1FLCIoTho
tCq8UKHIP6GAjykUD1QVXGXwTeub9cC6DApgmgLuloj0gZlRMJ3DP2euDR2gf1IhYyKEB1M9dh/0
RDCRFz1gC7u1RuMRnxETXK0qM0vvAieZ44g+ZzULKAuTI5T7Qf++Nb7QYttgJvKAl/izoOXxm6Xl
VVuz1/sM2nLVcBBiM16LFnUoAcL2idHy45sc6h1Hi6xdFoT3i9v/oo1ZTqzbPXi6O8/E0onBJutJ
nnlm0lnkfy7hy/kibpjItC6QD5fS7J/LeUgGqbqYM2fFqdfwT92/EO18cJyotquVTX+s5lGmO9LL
NDeZaMFI4RDcpV/LTqACLqsSjxOU4d+DZCmhbicl8gZeuQclK7aAFCRvmo6v/Kb2GASVcGI3joCt
8r9SFvkbSVi8CdNDQ12smarw35OKCbsn0M2HG8Bsy9LvU2oivmA35PHr/3CPvyWyZdunazp+C71X
GEPu3FQ/vlzJt/Z3t6ihZNTZzAUKSz/zccJ9neONvyrHEkh3VY/a4D8E0WGNYk3XSvTXJlY3fMji
7PdHpslMFB6jPlWRf8BnT5QW0G03HozgOXfQLVCnfq3AL8QWZCEfbZFV4cndKw1ipQCn/uU3A2PX
fIubA65Gc89WAL4/RJgcfkK/jrRSo1tKWv9KJJtKKDxWGtJuvQ18qKRBdpBv00ZngSzWk8EIwDHN
cGd+22gQ/Xr3lTiY0YWjC9veRWplOVOcmFBVA2l/UwLd+9Oj9K3F+PMIlyoRJu0AV8iPcPLFZfNk
SwSa++h9VesAmXYZERzEhV98zgqLQrRt2Hn6sUd7ViBvbmpDq5/x6Ug8Kpa647q57782jd92vrHG
YuMwRnSsypKeSka+hUp2f8aw6Bcgvm0dk1Igy2ovqRnkOBVqU07dUMoOVCidbT1wSblXxx99PynX
WRqk2iMqfxunIPDugjilIrUvxn0oIw04UgQRBFU7L3uxUtPGgQPb64TtoReiqzwitxDSIQECsYNw
uxhsxzXIDH8Tq5pDOfxrqWTKUVdoV/7tO3YxCgkRjzwJbpku8by9UTHtKeYNYQ0w77wCsvVWvEuz
iH9nB1X6lAP6nSI0q2HJ7/9UthdSNja/P+RROQpZ1tIInw7MXMRBOTbB5bnInHm1Of1sJxQDvo23
wcgvKjJeAE98/Fph0FDfIOxQfk0FqCRLJL2d/kgXfkak4MaCjhqGCGCKwh3Xf1kiUJTB1I4l1GAN
BJh9My+m3O4KRmaXTxAoUg1vp2dNBgFG1pSGGJ3hkz/0asXkKYg8HH/mB6/esgUeHBHbeYlaLv0I
W3Kcy8EGGXHqXayQBbAcmiVKphB0Up7ZOl6zfqbty4D49tW4imr04Nzx9EFgYmrBSXPKBDadACkN
0XwGFiKjjybUG9Ki1TVIp4dE61NT+8THJb2Zjj05qHlvSedBjn6YJYdyTrO0Vn22Rv1dP9j2w/Ql
buTBwFosSMClBEn3evzSSQKi4utVUVwK08Q5aZoQmh3wyaarcLA8BVMPOgUOoh0p76VnOXOZVQKa
iRdYxbswN/rSdPFP4t2SA66uYXJkPpClIidplXg7wC7K/upMH5gg18ttXJcS0mFUYmaWpjDCiX/n
wMA1V5fLEjxkc1y7BlES3/WvWsMKuZdwD4Xcej+iu1gt9AjWvA3PT9GHKhdEL9VGTFnR0K++1BRL
yZ6wxnLmo+YgusrwUr0Tf/T5BjhFE+Nj5Csh4gMURvctlSyLHaz+QesoGInphoat74LuMVUJe8sZ
eu+Fw/z9CSBwnjxrwDH9EK9hnyGzrSJI6M79h5iZSUE5d197LeNhEdmfAgJph9CQNONx9kkjRz1P
WOh9SDCNzsgonDF7jlmZC0eb2+yAVG48n5XwVJkJDO/a1tYC1SPiN91detTC1gHULgm5DPl21U9I
93YZBn3bHgp4UKhC90H53DU5kKzAyR5Zb0rqCTP8SY4kxrlvtiyc3xqB2l+1AiWI/Kk9ijpJkJV0
1BVXZuNp/bC//iY6EfgJR3UG9v45keZgC4odaIMphm18eORfvl6iTxDlaM4on+b2KXa2X+8mj23D
+35haOEJWBVOpkRTRzmho36yFObA11OaEeqsJXLHj3dVHLoDPcaibe9geDCG8ZX4kn+FOddYqmqZ
t5uFX+CgDG9q7HMsCc40RV6vDNOC8qEHjKOOsLil77GQWdnsRsKWHJ3LbrbJp+V70voB1l1Ax873
7pubkOTZ+UeMNV+k9nUEN/DngHc+55BfUYUKGVmPTbvnFIh1hwhCHDPxGLle9DdUWaWUMwbWDbi2
rhZuuykEfDeIDKpJ5gRWaEPPaTbwN8EpqBdVXQ+GKV8w6SQo0hO+w6NYEMOX52+GsejYX1EDJwvL
VwHWvoUR5560xgSTsrdUiAhMxnpFnNsAM/DooTXpDBETh6XxEzkP/J7/0kFQU+OH3kQ42mVdHaiw
XoUSAXpyQZoBhEJOV7Oa4hhWAJtGcKTck/APXUcjIbo1mfLPJ+RmtS4VN2Af6sAV8wQIBeKsLSgp
/ELynyHbsoDH9n30t0HoFfK1FD37wDcqnZjSE1Om4qH12xV34fIfDIFNDa4WjVCJeupJJvG+8tTT
Panbo8kPEgFyfdqhQf0OwkLFDiGe90sznU0XgtGsCyf7UcCJV7EvzHTqILtZhMc94JAM9prvtEJO
wKkpbQPLEX6bZbVG/XUeI9UF8pQb7Qr2IrQU3MsK488Po7sEb4GN52c6qwnBxyuQE3WC8jrzutWI
csB//8TgRog+LGrLiiaSZjoV1no72aFEdA6zjPihX+Occnk+S+lk0RWlxNWx3SqGrgrqrkPhV8Mn
UGQzI1vIu37RIFT3IZrT95CL7Rz+NH/3CuW+xJnrw6fFZhSA6ReBwugHE9TimtUQyyHMHMom5tXm
OgaVXMtrNviz2uK06Gz+tvP+jAs3XHS3v1EpsqqzSKhR1utBn8ZiHoOT6Gk3gDBYUvHdHokPipn4
DwkTEjuMgMI11SwHl8YUQWu0HnKmwKZBVu4wdnUMRzb2o+aIAS++TxFTaBlhA4Xf6nqde+AXqWDo
trIk6ZfaN3wWSMXW7WJFC3+auw0oSPXdWarMisRlQbPN7zJ5XSYRqCPNI3sFs3gnnAN1sVplcXnh
qhk5tCjv34H4Fp5J2gGAJsdu1s9w2RdryInZjBCDweVU7xG/2Mz+QvZdSO13ZOmOP2+Tyz5cT1g+
96HAIALRoGSB8u7Z13XXM6VNWDGVd94z3FKIJVaWMHJOSEZBmZLS2zU9MNgnZMTJbAl4TgJ1Sv55
sKvUO/NV8YYNeYk/0CUdfPQuIos/E3jOtmlyfDountqbE5iERleVXzQAcOjJ8nGc4tW3stD2iQDg
l26q+57AzpDDOYppCYfi3G8k9D1Z3sr+bZfqs/jxLVcOuj0NeXDsVfGS6aklXWElqqfLSCmTHcv6
xxeCvErkaUf+w+1vDmBCmCb5epQwsQDOxbFIQ39Y3zs2/0SAQQW+vzvqw5mqQg54OdbL2mOAtFtt
uS8ZMIK19NkDLGYai2jzefrFkt8mKV/8GxZI6UsfEtRpfsi7UcGgfBfspLS/oz8rFZHmNd/Dcjr3
kUK5frhuD7s0o4M5Fu7JCdWzx8y03puYYWlpqd7DNH86uVsFLYItN35yfU2tCDXn89RSK68qp4jO
PNfqWlZ5XnjNWJbwYn5cTonbH397rl6X/BVG+7kOt1MjC+nKEsEe3yjl8wdeckZ01+MS5a5vhd9A
MJh9QS97uyZAj+CTfIFgwfO+6WH5bugEAM23uJ2XiMmQf3ydVdpNu+7T+qpELPsvuRLVLUx/4POC
z1RDU+BgPCDxZrSBQUngmZKu6IkFq8dNygpAn9vFGDkILhet5fzoY1QUhTy2eZvfRR0mBVs2+ie5
YdD4F3WAG+HFrzDJaFFGK+VnyDYQqczIaJNNCbB+bj6L7g7SSNyw59ocN5bde2R3JTNEXCknL18D
27eU3KjHAgKAbpPQm1T8AQP4MAjySUFOVjWeZ2sDQ7oCxQLAFoA4t0i1A/nIKdGhG49eLTb4LKY8
/U1XT3T/4IB8gWbIVmiMaugyxdKjUeqLmmppnNgXONwBRw6Rp9NNdpzxPwwHLtNuycL6C386d1L2
F+IRP3dv9Sd5sCVfAfr4doheMNWvIrh9jjnIAf1QqpkpekC0f8RilpMvbOWtNfz5t9B7Hajeh661
Q0usMlrSgJkE+iKGquJERmN7jC8Qo8ywCMvsfcb1seguVjV/AKybIc4d4IxsoqR4i2yzCPJ4l4zJ
mVpxfejIdeBmkTyU5IrUAUegn4tbymImV3fojPF0fwSqnCDWaGy6A4WLI7cbLVlN573GtZsj93Ib
+1nIQnMKkllDyVBDrAagIdp3++FKc73KLQa0BDInWTXy+rycGjo1xSgyzF9Hwpz2pM+6O2mrh0KC
hxoLGcdtqfyO8i1RXV4zfbdwV21VRXEUZZMO1asjdxQ1dCbJtfHqLf/Pq6Ii92e8Gl6PhnMgsvXo
u1gaKe4XcyUdc9c+GoGe1Jh06NtcdB+H16Wg/E6xFrXpuGYh3ky/PUgHTr1JpQx9D8zAFPmNq+gp
9hqwS7gsuGqSRtrvV4MoqYhP0K9Fa3FyI6MxDE7V0fxVSgAtUCYbY62fBfIt73ECYumFd0UQTvgd
WaZxjfd7247c0bHbJOPOL2hEpWMUDB2sk74Y4Tu4e0+O66MJdMopENgMHFuami63TE3ot1hHuJV+
puAwtgPQq7oBVtBlf9JO5vedhSHPR3TRn5GkP7023DajtZBKZhTc5b5BnnBoGFAVTkStbYRsxDRk
AdkEBHx+NTnSqclFLj6VmJPuo0dBcXX/AuX+CxP7Vgua64vdoXj+4esmGLkwzHnNABgX2i8F9PYQ
wjJe11SIyGeNKvxVz0XfrOjH08ctp86r6yOgr5Rgv751MynqA1g2ewNeH9QmNXHnqXeF/fpNA15K
Av/98X11Luea3YLQoCNBqU4F56PTvSxJjWObot7SvkLjAK2bPiXfVUsrP6JqvS2Q6sZ1SkMGvcd2
Gu8gvOMZLIAj4OuspHYlObdIEzHglwbiJTTt6Azuy2WrwFCQ8r2WlOncam5f+g/EtpAgBEiA2zQr
hGeR0phXu/Ah8wB/9+5GuUXgeA8NhroAgDw6VRIsNtcMPLp7Xx39IroPpjTOp7lWIs1COisP5UPC
j2qAybo/IGSQVv/YuuwDEikyGLUObJ84JkCB4Ai9d1bPnBBN5ef/w87bzRmlZc709admEWAdBTZM
GcP9fGrULONTaWtzWZdntEn5qiqxhOQJIGJ7o7bndm4VNn1ESu/cYFglaMaYdsOgVbJGKZ9w4r4q
VZutjpZ2tl9Ruur2kGpVSiCHDxNH0+5y5wmCC9stAqJ6ma0Z/+cOoHYDbfWc9rvvVQupOL76dXbb
+9xRWbMxfJgYQdOl9IXhQH6SqvJtBjSpzn/OGbhKuoYZrk6htCp1CD7V8JxiNUPlJZuZIXZ9bsDS
Xp7BLyF4Q2WkkP1yi0E4USzQ3zliSRbwUOibNFMG3W16+279i4K8mpywEk0U8UZwIEChxo6gRwkN
Zzaz/AZliRauccnUEls9Ei8eAp+lrsIpGaLp0agkHFkqjTD7PFEBo3FmJYuCnIsr8wL4OARq8Mca
yEFoDbsYVIfg9INpQi11yw4HIWTvF8RjC3alnCrOdt4Gd4mVZmRvME5oeqpGBkL8n3gAVK9tIFxc
cdpxihqJtTKYc09Mey3juFPv2KWPLqdZKdDr3julOnvGAEHqTXADZuKbwsbeOFI/OnEDQbTWLs3v
dA9MuLREsboTzUmbI2U6aeLobGEzOreauWIw3B4s13rLHtPjXF4yEoILJZRKSLJqnvMxEEbvhVRB
l2qysMo+8GHaYwr3IqAx655Oiey9xBApeQhX+n6aUfm6WpejDc2bLsD3QRb3SQeaedOswGmjL2kP
RARbD5odM/DQxtrkNBVN3rfYm40GxTmMzVw7cAPUDn8+1yLA7H14+s1yYW3vfKllE+rPJZaaMRXC
FyZoP7kACwV/tA5Je8R8wv43tqA0xUJDeCNLzU4JYirPIbczeQe4RTi1kLaewa02xQeyVybJgZjo
Wb+fizDFOH+o1zGrnN/Z96HDERNgIeYbrAAvX55F179TPGVYPtjT2ZeV/CKn9Rjm/DqpQOjGXPFb
DcvkHU7+HaU+87EUIW/3j/MCupLavsmwlLV8rKX2EOPXnOZqjsveMc0iBj9hLd8AQy/RaMOaAM4F
zGtYtIolSyDezIhGyRJh/zjQgWtSNAEBV4lKRyDxPEAklL5CW0PF57DPj/41Y0INTySdyAjMAxYw
BrA+g3r9b7wuI6kLOYRdE2dpr2hinWAUmJn4A/1FAXJysIH7zdv6xCRTRZLDu6yNUhT+ki+cJiBs
KwdFr+CtDZReYoFJHTJnpefbpxzn6JyVu77hI/O/Y7rOMOdcvZJRon20rh0GvZr/ELTNwLQDVcJF
DqKGx6KnXIVk0nLTsNM6u4cTlV2b16K9XbxaPvchnHd7PIvKNIaNv+wUDI+ta4cLt6dEzM35JgfI
HweoReI199JL3jv+m+oGpdWE68etdDhtjSspY16TH9q6rIZhXKC9R+V9M1S8avHuvDn9zBhMxn1k
5g/bfGZqK69UlrkxyM4TbN2O53X8Zj3PU/GGiZ5tlLVPuWHw1y417yEDwKn3pW+LAdmIMqQ6+TQL
rOmzw3U2Tq+MYFHszDBmsz42rgEzBYrSF1jv/V+dY4SUgV9yZ/xCTO5nKYYVnNvT3yYgv0AynQ/v
bmLMI8JXvnmEzJfE/Tql3s8DAgnfVtGVJqXujoBwTBC+pTOVxlQOStKaGPEjzq6YaCZkUTwJoYkp
KI1QqlchRlad8csIR0tVxBrc3PdECmmuZkC/JTDxufId45NfKSvrnNfXOBKQ+sYuTvPxlQu9YW5i
uCoXlflIty4mqIGdVwDzfZi2izNt4FP09lmSEWhcsG8HUYPc+5AXVARfNn4yFzFwXYx7bD8eLzS6
bHApmzCAKFRtnn45jyb4amzqplq0fls9nNFFyk64yX61EvzX4MVhvG7zBQjghOBMVRTWdk9V9AA1
ddC+BpybaPS1vYx2X99jzggEo2UgZBRtFde10z51SSMfUj5D9W+vl1KjEod1mVkoy+B8+s7KN1My
yvyMV8fDvP43uj11SS69TqVPno7B6ydrb3k8qfSAUnuJNOLJX6a5L0FJ2V8GfsbPyfcu+m9/CDRg
HkLBZXjCMGN2bUjjXxbcEKMf9XNi8hX9cUmSrh9ursm9dIf+6XX0npgEXMmOR4m4JwdrhqTWHnzx
lVWvwOvf7/bgk5pBDuMz1Q86gVaY0DHDuUxOeujdw1ClQhxy/+ritDwuVnC9yEHr3GAwYTwXBYzS
5ijdvhJLSMBjzjXJVIyMgY8urPnm6KrEQj8xrB7vHwy4i8uDjzMkMiJUWdkBsJgT1CQCGqsLoWPX
OHUNLM7XdrnbsT21LWdt1iXmXnwP8ccIEKJEi7JtBXftL+P2D6I6hPLsrOmbfqcKe69kS/nIxLPe
iC/boENf1lwiiJlLo2hmqxMEolLhRUG63e3XLy4RbNgrjYZ8exaBSM2vTLRELyp+lvpfc648JNkg
6nWjnd064Cy2/3mkD79puepZn+z8ShP2JnDToRWyOZryss3dbibjPDPcC+hE6+23cGXIVqz2okj4
WyT32fS7FIKZ+jxPu3SMcnj6VqC5TCxOS+UTm0wsCSEA7pcWeH9Ht4n+iYCvVUi1me5ZjhxctBEr
v8N4xq8MeUWxLlBk3UQ9AUDdmGfxkX7dRPeUlCx+/yKm4BmMEWD9Jw95FF2dk/AbY7J/BG4GP3T5
P2/3ttEGtiovT2RXnIAPNEjxgFZfqY7sNW7BZxApBcXAsqPolfJghVswjzr8xoXfXk1roOWKBoqd
149PY90ksxY8OxDiiafQnATG1SHCuCtI9vKkZ4P61hbwcFuOMAfkhMhCjEtfu1BC73YfvQ4/FJqy
vVxuAgCLAQARNGrY4QWH45EXMNKwyo6iNJxFH5MP0SE+ZWEIoINb8DrwaXGc0Rgj+4PpKa9DrtSA
9rhwLPRDch17nyutO5m5gGwhVGIf4cjiXWSrPDAjwDVFzQMvZJiLYzJYbIOChkYLrSEK4vPRGGb5
QLW9J2ZlQ8zIyKjjL8GmM4KRLh/MGUnJuWnvZMzTwu+2Dxdg83ABA35/ZdZLcamsJvGrcJFCnZoQ
gxcw2zYdeNg/LxhLDZXkR5BXd6L+dhwT04rUQm3UEcU2BgqwUtC46Yc+UR1PtG0mBBFl9sqArE6a
4yDYevICX7UUXjXEqnfQ27ayQVIjI3pKICBwDlMN3ammu5R5BKuucd+wdpvQAeMF8qgmwOjpXNUz
9hi0sgLGlHGuZPcpzOpZMrUz8SG336bi2zs0gIxXG4hb61ncoJ/y5IlnJuvIMlvRbxm1CjW9MFOZ
g1WKg2XRWQOTJjcakeDeT/ARTll810VqLYG2QoNDcT0wCweNlpeiCzdGWejmmXSA1NKzFucppxVh
H1n/IZMXjbT3ptJzQwRjlRlaL26GjK4OHCF/EheOwFMI3MLvDAnNRz7y5NH/QjXfM4eJo82MyA0K
kgeIAMs65dfjWn0YXzRs5Gs4wuC0BQUoqdQV9IBfQj7kLEnabJD4HInrTQkcXzt/Uv5zQe9ZGFl/
dYu48QQAXLpZs8aIc18Ar3Mu0stIFWFMNyzUcMI2lGF1postH0vZYmIQHGHucDlU62SkI+xjRkzK
wq6RACCMOesIglZ2b32V2CnbmSjKBG39AOvRo9v1DVl7cIXXJshtOT2hqcwMjj8ssYn9yiPvTVR2
qR1QoDvEVXOKf626367tjTQMcF6yd/w4jbV8RZYW/W5njTosAhpLrBgaUWiYlBm4BwFs4FF0XD5V
idlHzNHJJ4/4FI1diC6mkz7V1Vp1XVrOSkov8POC+N2obuv+ren8FFl9scwoF6tThCGiqtV+Zyid
bxLwCJgitLQS47ZQLkHi3oehE04X8O2cDXCee8SJxKyrbsVIJdzbSpZsBU3pRzMRhzJjFx8qLvXz
a8xRkHzyl9Ot9sYEWuOrmtlRQO1QMNrTJif2bfVDXYCMJ4FFHkTZIv4svzU9SPQqdwZDTRAsi7t+
dtfD8QIrZjVHb43VIl9RBCZOJ+msuw5OZaLqRwOVHlgZa4ej9ESGugS3H/T3/yKD0cJ437SoGZ3m
TIzAUt/GE3VZJ34QncYEpQ/hvG7R4/gqRa7Ek8JUzv249zSOp2WLbgmQJo2ul3v1MCC6MIDv4/Ul
i0jwxFUohBgCtV4nv5PFscIWHH5Q3TcQprLx/ABJ9EGZKYeePTYxheAQsEyi436zNgEOQ2ZDdFd4
krFnYOGGpVKx4yYTAJzIAPVazOyCFu5k7op8MpK9Lci6oexJydZOcKmu+wwfBIvyavlXkrT6czMQ
czlgi60fj1+B4RQCIabrtIHlFcyec4GbydvsAbNMNopx48PR1e7uu7uatrVhrX8j1vU+JEIUR0q6
FRZ2sA4jIBDRnQoDj35jXlv/I1Ae4j9J6wbaGkTLV6JpKr/iAbkmUrBICF6qso1F/3b/N0islKtH
jLIxU0dCVUsntuXwKguXiqBQRgNPuGj0S33NSfO/l10LWCB2qEjoWc+x5OgDeBHmDD51HbMjephA
cDjMHYKpJHOlLVjQinHOeTMR7cDUysNk51p7Y4GoziRhtgkEpHkft+GePUM9mceGkAtyW0+zZQhP
TzD75yr9AvmSJEpBw2WIlqW1LYwkf0OtFRfNjHr1kMvfTo5fYwpl2VXSyCjxjT+AxHKJu/PbIU/C
l54Y2OLA0HeP7PeuoLE0xwTKd/PkQfKYQmtRzEokhQdiAJvIcbNmsNQWRZj/Vc8LEaaX0ZHPcRI3
5xg9Q3fEUsVQrtYo9sMZfyyPNOpdZM+QZxlOxqdfoJFjLE2hS4uwRkoioB1NEotrrEc0TKpHJQnG
0QKQ3lR8odK+45vZyq9/Nvm3pfDBGHXQyIhQT3SmVPqsoRP8yRf7WmzZsh7YPCp4ptCbSzgcqoqy
nwILqVeuwAwhkdB8X6zUGxEJgfQ7j8Os8ad/4qV680JIhVP75jZerM86ubhy/BBK39XwtGONkmJa
TJd0D0upLMdg9Vf++FqmtQITnpGqQT8hoCXyWUMiKxC3xSesephI9tpdOLwEKbXLy9SVBLlY8bb9
OzYJ8h1txEJUtqbtABsX6jd0Zh5bEq3Z6aur2Uw4IL54zm32+ZWYknkmH1i6eTE7Vhj/DwZ8ZRzP
Zcym08uQ+FLmjENPspavSLC5z/bUueegPpkkKIzN8oFDogp9ZshKRtP1ulOLap52ExNQBvUOQEjc
Go7kh/7EyNJr5GVz1x8Xd262S2KfR6VOI8mUBAhIvLLAq65GSaMZKcNGVARvIE0LCzTEAmISNI3n
3N6hgZ5ujqE9aW26NcvuBrwKA84jSZ0JrFwZ3taEkavxT08xZibc37aAv/4CatjLyF6nX6RF9IGg
JVFIBT8hj4IQ5QMuqJqikAShJpZiU+cBK5Ge7RqInvb1N/gKZ1cLC/q0QnErARUOJfe4xw1QXXTA
EImKW8oK5aeGLXJs6eVWpuH3BEeOOL7Fw1hITfqjrtlG+N8FhdAlNSNm+F9STTE2b0ach7VyBo+T
BuLBOoby8kubsDY/O42ULs71iH0ijknk1ZA0E6viKzWeRkkD9ypgUbbTUiGrTKFQrE9RIKibO/kP
0o+5kLgyB0tA2mode9bLGBMKdjig6s2w33WCiMKB76jVIYHvYV7a5yWkBgUZmmujncrUDqtMRzeT
ybzvfyXcQMvYf6A6ecEaRb1OUrNDocvLZ+eqJ/jC341+pjfoOpZwDQ/5wWPkUBoYcYcczrw6/keb
zgd67ef/0LKeeGCQ4oCcHZShIilAWpDRldw0eTWkKVXfr38yZJhFBnZud55IBw81S7+yTk6A4e19
ffqMh8aJ2lxK32dhzkp23byKclbVnF72z1LnXWWLUUVfloM3I5Q1G2IZxyiG/T4hCghr6zdvluvC
Spjntq1dTUTJqvi1yPwDdKHgdLYJpbhg2jfAem+8xymd2ZlNbtl2IkGOLBSoQRTy/F+6LZ1GMPjF
u5FqEVHldR/IM1dLJ9lZzpqwm82FXHZk1ViTLQSQZF9V9Cc/Gu6lcSydGgKct+LNTYLeQDI4gkfX
C/Z5DdtELZSKFC0oTngpAWHXlj7lVE2f9evLgUc0RXYBvPt7kSb+o1xttLrCVf+NGLe3e0cS/Uko
NtOZ0o5XVA6xjP1j9pLvY1xRtIPbdg66/5e8RYnIM3CxCcwc+knyIRnuCrF/zW5vIhlzt70YYiK7
wuoR7kTWDDTwgGEwuJokBQAPqCo404EaODXCUxlAIaw41I0SJ2b0ZIOq6X/HXASy+xic633Kv4fo
OwNDgQgmFOQob9MokH6qGSE5vNIMiVp6tsIlyBdBxAnZFCoUysMxyztnHI6n2Zn8vFe3Ko6HCEUV
bbYxbs1T/zmo3bBPpuVSZ1FHk/p8biTZCypQLNK6tmq9LEPmk4UKNq+5q0InrlOq+XYbzr7ia992
vPCwFOy0RCn7VSFWY3mgLg1ySuU2tl6NWU1CZUD0K9e1m856VnYKJanqVlpwh0bcCKhpEKSeB+Tz
d3joQHOe7zp8iwxgab2M0Ltg7EWQCqB1F9usRUY2a7428fpj97rKn1wOlwCjw6HD6xrIli13m2gg
qSZBuTXbM9RLs8nTtULVY1CVttO2Dyh6r+CegpNkcVIcY6iq2TR/1G+M5z2eZK7IlWDFfcXChCEO
oz2J0gdK3Er4QrTEaTXm0hPyIQUB6QIQXCzm85P4kBbIbpsWOvKg3jyeXA2bB173FqnCWTByXAUI
hEHdRhBL06gQ9PA1UOrc6zX5CQsDcF4S7B9RVKuu8Cc+u366vhs8nbVLwMT5/7BGsz6bPmTLXNRj
oRA5bBNA7aMsFLs2uxFHBFVTxCzHYB885eCJyV/23jLi/3e5GeHpdrdxjE6ThUNZrD/W8151fe/w
Vj9ZrfTNi2+1K8k5n/5hqcslyNx98qoSdOViZKDjSLnMFrOJ0zDWEPb8HAy4Y6AMe0Kuf4WLaDLT
C0T1f01aDPgT4JflsETs+vT0cS+b5+7rPDju2vRAK4/GM+xxzXnFkAOxXvk3ilAvUoFmJAphkYMP
9G6DYJJ6Focca18LM+e18/tZO2G8QT08TASrT0aOkyRgn1MKKXhr1I5EaPRoiCw9hFC3BUCje8hI
dCAF4fPmCU8+lD99rDbVtK4kAmTFxpzN1MY48LzaSv+wa3Y/1OZcbJ0hG4M9WyIn0/bDCdEKtDMj
0aTadY9urKgqIWQsKAmxhRy/zs2q7Ysi0GitbgI1UH6pzuVVDudBuyaAPNHmohoUWMVmBW5+eRI8
b4mUqoXjuuru/j7wTsPBJ9yvYnZjVljtd/d7qmY2vli1pZuVGCTfqXQ7N/RljFJ6/pZFwoFQOhlY
1x9ZVKDu6b06dFpa1xUQJH5eEf+yFW1fbx3otfGtNaaBA8RaPTMySQdNqjTJccJYO74+s6Q9aW8b
us8e2KwwS10j9yR28U+STHY2XcVJitDHcirCuB6cXhwlhFwhIQq+fonILY0V6mr02iHijcRZ/5zT
9cSED2hTgp9VyLSTjduYzgYAElYEGI5BSqxPpdUQiwbPp7eR6sObX0MfGnMZcUpVUlGQv4M4dAxp
psQTEpLQo63bzP//euBsj0IhTutV6bKo7nUaFVdV7kGlKbtzqLItl81QGq8FqjOjo7aDGG72NbAq
SRRGQxyaFjimo0Tx/d6v8LgkNfdtnqbM5c5xqP5R2GB43IEwQmUsAxlXm0ECwfVyzyhg+KCImyMf
LvEqr2/uwBYDarZ0NlZcJGQW5girtwr49U1NX7Sux3og4ruBVdFDfoVq6jJfYb/uhtIGCw7h3PIN
vpyNiVGV2gkwEfRJg6wX3qFuoGXo9OJzwiE5DHlHLj7XeyjG1bFfWXT/RAQolSOnOz9mMqz9184v
ssbMZD0oJlWhIvKcWmXMWZ7ZM/VpuXlqU5xFhB5nXdHaAtiOuSSC6kg3jsCttbz8IRLkhNQh82nj
O817SaSFDc33z2Y6WHMgMr9bZjndAy+0YTPX9dw7ekgkC5w5f6GE0OvW/H6qWYTFhC+mu7RTttr1
TJIVUWJIAaC7//6/Xc5AUQYkGUoPsrWgF56wNxDBTj7qrzZMVHT3fvJiqIg/11Cl5zKeRCyzTJQC
hUFdW/FpcHCSV1jYI41uTKMhsGie9e88XSFN6OFkwGCAgu54z+6l7nrxLf1pKaApP0tv8uk5cu6A
Z+KEtDD6pnn6cHy3sMJ8VP5EuC0CWVKGvrSdetkxX1WFm6LMXg6E+vG31IFxjfTGkaI+igiEtk8h
JrSQQ3+ajIs2T4pJlb3NC7wCWzQVBtfPuRYhs/flxT2Kj1MM/lOjO2IkkNm0lCZRzHMHHxOUqgL/
EdKtYr8N7lSi6NoeRCTsYbdd9IhD9qHKTvsOoD5pT0oKgq8aoycxBnadBtUBDwlOMcje9pmAdMYj
8vL2r0tPwuv4PkuleqxfzojqgArI/MaM1T+cBAe0NuaacRsS5l8YzUzTk/LfW0fpfH233Xn1yVHB
Q6pIRVryxCsNpwj6IizIG9CQpUtza7F5vwsMB+LDfPhBWpXDX74BRqY5fNWEvepkkeA0la3KWAiY
evhk7DzRZn6d3Id8YrsRPYH5PgWywWcU6jf00TF7L1cRykHotBQopTqmzOlWF25bc4l3UFez2N/T
xhRcruUD04aH8D0sVnOJlTFDI7QKRAsUpUDnjzXDthkFze8nUT3ceAhZZI+GsOli11hW3kQcWB88
IEhb4UriwP8EHWD2E6olwA4nB9B3lShE/wJsx57rU6lARHOvEwvH8RzwKc2AFvrS46Igce1YXNzu
e9HLxVF7hahBn4bmbI9K8ZsNeM2wxDB3sDpYoH9eyNISR1xDjHZYMI6yekEq1RrVRqhWhgjRtoxL
VlKpzvORPUurnvNI9s+EqtcN6hZXQlKbg99gwNFgZk8JA5A0KBK2jdzXtikrLryA7pX6ql4+ayiA
G/fO3tfXOma2tp/Fcm1anca5ny4TpT71EHTpoviOUOE6mQfL9NEOP91nC91d6s23QpNrmrIQPdbn
vXO6GveLSCsyCyZaquxUIguOnTr8LT+oRJOICTDfOkqJ/PSShUEN2isHj/Rant6RpomsmRMD487R
dojPVOm+WftfTeZw4FLK5Sx6BYRw6aisBlRFnNt72RpeHhQ6DEnOdfZ8HNB5DCeI9GYuQRkBZ+Of
gPZjS8Y3mI5V1Y6KaDKjdBEyqcW8SoiChetZ1qRt3mANZPr2eS5aNAtjYgFqkYhoMMXTNKInqMJj
wvVCzgdsQYTsKQ2O97SBqVuo5ZoL+RDeGtdwWRaaLjPlxIZO9zBGmby+0YhmTw6T9mzyGCih4s4k
dQYXLIzZLjjhT+css5uxQ3CbX03nJifVbMqWE5vMN+4+G+n9B9J7X40GgIYQZ7wvOjf3Kz7sq4FT
qOU8IMJN8P3bTJPUojDHcpnCFW+A5/LbALo+ctk6SzaddbBKEXgy17O+hFOBEe8osGvics3kj7Eo
rOyYJRPx/ySPX3Teccr9XVjj56Y/2ps23WHxrBaUPIEgnKzNt2LIqdg0Q14BBuzdAuQjAcITL95Y
B2G4f37CfZ28wEqjzNgmGl5GxX3ho3V62nwus0Hh7l9Cqqj8OSHMKPyjNBh2c+h/ytRZzM3Gy+hG
CnOPsZF2NEnsxL4GKdQjs+S16fKxbKy9CCfJXRSeOHX2MJeeXWwOVHpmS8TjxDD+m0bweFCPWk2v
hSWOR1OI2lDxm0tQDY4xBapzyxwUU+mpHFEPm8JSrmP+lfvfxD85jIkTQVMpOUAI27DWMIY0Mlz3
O256Gl3RocTCV0uZkV0JTJBbPc6HnVBI8qa/vZgvQl85CWHTX++bGYEfxteeCRQwUEbi1ZMeRBhg
G57QWctdYR9zuVPdzpTuHWhbjnLFP5bGktWSAQ+9+6gSDuKizyQF9TTrB5vLqGLVS8q1q2o7ALCg
5IuZ5pfwaAB5UvWZKBRtXhU3KY04dYRghAp/UZ0NOQqQaOPkOK2WPgPaNN0V8smF7yMrfmVhg3ZZ
NEEmrZd4wRSHtb0pu22a5C4/Vokcl6rG/qTf4r6AaKmMjklbEZrs4VnJhUiH9PueFXz8iLvMShwu
KfL9s8e1p/XTDRnhjc8QpUImFoAh2NYPNrHgthcf6JTIP5/tZtALhPHVEJTv9UZLRL8HTWRbGj+p
RPsTlqrQOve9pGPcXQMwohkAdxc/yAwloCiaxHbc01Q8eIrfBRKL2V9RhU6D7CE3JdioGfzZGz8Q
kjS7YFFGbQ1gWBWfteSCm1AFIMH4rkgzms2unbax6Fmc3o2b42MXVkWZmBStiUOimb8sLE3Xm6gL
i1AUPdUjeXZBKcHrT4sMsYwvfApRckk0JwNRrvzPQH4sR3MftRRw0Guoph9N4NS0OM1aU6AIFAks
q6w4Wk7H8EmXfKC3Fox/OErpt0W7F1E4spBzyFroluc/9cznCF7SLIuNBu8ckqALQm2RhEL5rI9X
bmb469RqkPCAaqz7uEb3ztg2jQcfCxqKCY4gZy0/TI8tL0QBuca9/Q/S3XsK0W93GO1lTGnCOahj
QQSFAg2KcWMNK4ET7SpmTtWBIIA6p0xRuOsm+v/P734nuHplxgKaHqUDnGUsOXKzc1C4rmiQLemI
6maV9eJ3dvlnK54Vn9ZOzsy5+PVnZBXdGoqng5emo1NHUf+lV9x1FLRgzjs4lQcXnn6He9v7oGIs
I9ING8SgSAv6B5R/fJow7XJWzdWzMoAEhwuh/Vx37XQZUwNZjUC0hlSRdxkSeoe0WjDDKZhTzHRn
rTqaJWcZswrRwAHICGjdEYumK/WxlLTI9VVohASBjhMYv3DEvwSWPXFMmV8I/wJaOGB2GRgW8GMR
h1QEUqsbyinDZj2kBkv6KOXk0a2+rsPuc3DIZlcOdm+Ns82eN7Bjh3pU5Cw2ogrcWH/CRG2fHlub
WO0+sz0fiIm9qpEWx3JFtoWGEjANJx1no9HAC30jb2KrCD3Lw5bUP00P4nR3DaYZp+8L2KcbJYxc
VzX4oxd+KjYyL8/zh5OAxxn2p6bzg4oHgs+ei6bUhpZaUj7uWcD/26Lk3AH44dVRlxXQTjcCQWf6
1ymho3p5yiHOEGJl2GXoPDYgv8WJBvZ3nBOWUAknUuxFaZGYXCZYKGE8M5CntO6uxKupaz9Mpjf1
o0gjmckk59SmpxvMEeN3oU6k7zGREkijvSXr0mEVlXx2p+lAaiCNHcRgvdfmMjyoUH/B46frnDrs
DylmLHegosTToTArRKy/f6hAkf9jzjrmr4uEBcatvUmMOnfthQs4jlw6xBEKPQ9ibXMLJIz9IZFx
hQLuQU+roKEHHAbScujq7OhIjXJZQyKL0XPt56aqEjb1A7hh7eESRq/nFaiWxFOVSA8TQn9BxtWI
gdV6oE41GYs5Gk8AQLbk6nBnIQMiG+kmGh6rDz8OjyqFwtqwhy3LXl9OjNTfi+quFmY7sE037dKo
p05OA6ksnaRTEXuUiODTOUepeIe3x1+WAHN94TQatkLjcpHF7vyDVQKA35xTKQjQx3YODVSPejS/
InTZLzTqM5uxGz8CfDxrucr4lAGhrJzdjphxpW9re2XPsMj0+/tdP+rRyVXMRlPBJh4rdpdvTJWl
F6CCkrKwIMCnNO02P7/rQCuHYD7qG5nRZu0A9dz8kWGtcZwO9NUbu1ZJBswJXyniNWPyu2GJwXk/
DrK2kYXxMv1n9cC8olpDF9Qw5namwD5Sc3/v8kK/LUBaAKQHPdpEFWdw8UL7PCrxO2itxVLjXwfE
50ZC8McG3nAD9IYSPW2YuiuEy2lvGKgd0IHrtyBtqGzCRh/C7kjYiJ4oKDoLN1QXSQYsSr9aEgxW
1BnZ7BZE8GdET8KWQtKE8v9LSREKijFC51PTUjNfAa/eP/eOq5V56HbBcpuvhlY0DMJIyuMikXiM
2sOucmriKmMGA1dYn+JnYA5jyLG6MdYX/oO+l4awwT32pBgGxJsnZcIXJ5eBZgETf6pvTGuDaIU+
jIv0nAE0y70SGa94XfcK7ndnhRMT3KZT3cgMJtaD/x7HLlgQthFY6FbZnp7z725IXbUbDBktQCZn
AsDuIUmk/QpSFF5niCV+KMdm/Ct+7/thdqsWn0gDoS+eRfgffiqTgjzrA5t30ve1+AY92YbAfQAR
giNdx2YrJHkXHpT3SWhHW1/dbhmlSE9/q8auK/0u7ZZHrPHJc0MvnJKAFebYnJApus/WiwSelosn
w+UF5PQeA6Ky+KoUGxcWeOpvX3nYEBMo8K+ule9uUEOgM2U/VDhlVqtIGyge0VJ16gb270pXfQ61
F3cw/Kg/2yEmbPSMicSUk3FCMKfhJiucnyzTF6lLmgmtUduG0gp4NwRPD1mvfNRxqE5Uamk8Au5P
xGqwEfZFP+3THzZDEq28tXEYiB66GTA9DYnX4EZ82GcR9au1jxD8fza442VCgpQ5/OL//mefbsKZ
ZFpZekUO8XVCpNsPHpzIlqjD4oZ3nQq5oFXH2fo7CpJePtv+Mxi5a10+4/R+qghfbKhx5efxK/e/
xh8mW3BTnENUSuuUwpi2yYA+5yWxUENhcJpOzD5pVGORP83/X6rWQTkJwkMo7q9C/uIQEr38gO3K
zmE25ovexNDw5p1FDwK6JcI+htRSiXleLgrm6bdEJk/B4mEkf4OGw5t0PBxciAWQi6Ag/ecLUrLP
t+qbeOIL2rDxTk+Ga1KPsYjUjKGpTC0Ig5co260QZsT5AgMs9LR8b0cMPeoFObMQT00MNiEQiUxN
8Y0D8HTYCXqYpDnRaUGme/uv3M4xJULsnKqutiDA5T7JoDTft0qz3F+llLYKdAFk2fDpWZTgGA8q
52R6bi6jkJERos8k3JGW4jf80JtWAsE7xyZ/EyRma2U4LWuj1fPwZD1lAPNBTw10Jd3I+e55IhS8
RlUCQmUcJAkkok2qkK2WKejsVpV+xFCrFFeT05z2K0/RkcZKnCGeHTpUjlnetQbG7R3viA5jLIGy
LPgw+fgAf2HvvBKz3gQax8doj4DgWbT4T2obQ+j4WoBkqOW+LIBBPzWoI+inTGuzfZdOOg1/oNyl
3BANV1abE2WUBPCMjrDfXWHQfeI/6a5EZUBlP5A4JKy9XhQmbZxo9d52KZCq5yC6xI4Smq/H4fqZ
KxpDzRkKvxZTn0aQgpx2o33PXiqc7o/1545GoTEPS2GdjM809diBrcjP63tp6Eex/Zu00VSgnNOc
lIEO8aJnFUegAb2MJIXYOrxnYFVFTd7BsdITMQ1ttbb/vRohBNyRczDBtyc0X7VuQhp5NzNXTtlz
WKVmP0JxkDewUzI3A0y3lqJiaCNFDTRA9T1/9tVuTrYN5Tv5vnTmvAfcMR7GVM1VINDN2O6I1ozo
XqfsjYd2m0IOlZ8ChGHf/pvgYapDUtP7TAmLHzTxenQdRMDEViA5tLSkTYNRpiV+fbZ7Szy5ecJD
BnGfcgC6B9XvazG6jJEsq9xBn0UbLOBhFi87zLo9IeyzhyN6rbx3wabtXBK1991DhTbmHDAx4o95
ZEOhz6oJxVT4dKXhwmEXTik9BnvfmbT/xtERSpOLLY8XozQ/mkEjlV9ciIZ14fKv9VQG/7L2YMMy
1+ja2hBXVzDsdaC1XxX3m2tNFmcEGurzXq8yRA0sTqFzBGp4AIu8KrYBIvRjtNlETG+evKyb2cSw
ZMfKQ63+yiFRRm574RvF/YOjIkvb01Te6/P8vYxpmydyV7taKRzLHfc9668/f0WF+cYDMsEyuX1T
NNHkiLQMoeWTHFdcPsHdxX9I2EN17tkIz3WshP4yVrlndP4sfFFpHF395kgf6/PmMrDwRc0DF38t
llaDDx9mh4e005Lm5HZgJWnR9EUWgfOtQ9FCpOd8/PJlx8AHtXllMPGYVfp85K3zWRgf1udenq3V
MJ7qbTnlyndYYlOg1heMSEcwxR4Iyn9kfYclSRCIAoNre1XRlsK847/sOG++khWTMPzlb1hffPfR
lzAuTOVmV0wJfM99TCq0FwjUTohZu4vuaIQMheXaW74c0v1eyuqUvm9bpoxlIYxhZCbS6x5PQ+He
asnMyNjhodHVTS9y1nwIPpOA0Jj/mLta9G3u0XtBQ3KtYJ15Hn8gJ8ZDuKrKqkaUC2uSiAKxiYZf
CRpL3q9IAL3jUsH+MEtHr/LT8LxS1uoSopDidiEVkAwI4QDCOF1aDXS6vsk8KGzCo1Uj50F+WHV5
DI5DmDLou1jFaeUtGs53zk0pvsjWt+gp2Q2T2fzaqDp0PLeB6L+QtPlhpLaU7KbBWxJxet6BFbnV
NHED9zEYl1Vz1OhYxZ/8vpI6KEtE6S5QaX1BDE70tS9+FyiAoI3lgz1I4GLsy8nyavw5skb+4mHr
QTalsE/PmD2z3RoRsvlNgKLFdwfyG7Cdn36ksT4zKcmFN1G99dGu4LTzH972vWmtVSGKx09ah0q+
XKPbFQWTC/IcDSkom4m//5DQuEjwpDwvVhuou+pvJvsV88xr16u2Xc/rx5BxiYjRyOGaSUmojcsr
FQ+0wR6QbTsxxue/Kl9MzXgI9eTVWXQ4YgOZk2XGt2HbFNDeFLZfhqsypVyy/vwsGRetag54DSFp
qaTnf4IXbi5A4vpKi3bRKasYGeFqhOB6SjfsXmISEMX3c7x8ECP09URNHsYNkYRuvRVc6OWHKn9U
gqpuP8uNPp9VR4UcUuFLRuuiS3OhAmXcPfraEq6jjXm2VblQm9ndVPLkqiMVXlKXu59q8Ih/Eckt
dA+lANq8WBI6PpETmA/Nvjh9Am0FPqGkZpeJ39C17mATT71jSDgGPaio1Kj0esBcs19EH4lnEx1n
6kVATZ33KKGlPgEb0XtI7yhtn2lYd7/AY4uNRop6FPNcwFfGrEbSkUkOOuJE9GYEeFiLCFtayBXu
Nsnz9PvViSxPI45Yl3gX5Muacxl+f/95eUXF8l3W7vrjkgpbDCugMesl2eSHtjqjmAaeXhKY2PfP
HmJMRFPVRyz7hMf08tN8nooR9tpn1FnjA5cl4eP8A+ptkXuXW2iBViP8xNHQEPNOZnvvs9M3CY9J
oTOOJQIjVlOAq4U94UBRV+oInzxlaSIuDFhOTt4oCCggbJoKkl0TLb/ZP2HBr5DRG7YcQpVf9saM
Pd3Lpvc9Jnx4QDuxNPZDrACUcDXoeulziCggk/VH6gETvPpa9m1UeVjNL+0EmbfaYGD+LhVmWo1F
YREpslSsxz/1pjvHKv2H0BoxYS+HES83mZPII/t4324Wh+cw/OvmuQMUUocSZp3+DeNmPlfx9JUX
91QNQxsZIWTfc0WXGKADWMofR6p1eyyfD+Ixja6dI28LcvATVyfusJcA6B4alnA6HNKssxc1zKEZ
tyg7Ce6FFlrn6ngOqi+yCp20MP3HOWAbTDO/XpwXMK2DzCkYGU0/Vyqf+WdLKL5zrI9IM9zjJ6z7
f0TN9hmroCYAiDudRMg3y+pU8KNoCnIPn1x1JSDUMXGbnXjZQEvMaTJAokI0vf+k9/b6L1vi+SdC
LAhXyVoO8zfJ2aT3PSpUsrluFj2VUy13S/Yj8uvaj2YgGbc5e2PpHwdtb1zVbqOHj+lnpyzj/YX5
3da+mpy6ChU2zKIg53loyfV6MCzNLjOAAUlKidwAVRgGH0zMb4GY4TR9oJ0VfIWtM5MuTONjaCPC
J02ksI5EUYILqLTLtEwLOZVs6FsTnFoPVVPlzCsKZSlBx16zcyg7aoqckmGzwFf5+jJCz9RUYyQv
xV8BMwGDXWwKNoXqadMsk8hOkjPwxBvhrEPVVeYol9DMeLMCoNCyopTWIdLuWnQmx4I9yOPTemxL
nu+/Bwo7LlpYSVksYT9GUyPeEPrEkcfcgYND4owKZBXwZ3loZYIwP/GVSf0l51ZifQdfXJj1WIzd
t3GDJrEMFghoNqya/58PjIy5Bat3uX9zfZ7r/GrNtjLSgN514g7tsKaMzH0eiVbv6bvZh6rMl4Im
sEds6nA+Magbj4FnBTlcg+EQW2eOV4zJXitc9jygMFOzNTC3Z6/+nmmMdFXCclowQEZjRb/2zyk6
qIqbgPWfj8tR4MtFDJmCqz8PPb0SG+kF9N1YmtGB71nHhn+ovyUuq8StBaJa+T2RUX5rd8q8+its
ItZVJWr4OBnK1qclIaOMdPWaQdBtfB/6K9KNeRKNXlWEPmN4fwT7boFmWkLO7ZPR7DOOVhPzPPld
0Rd7AtbUY/MV1KQx8PzQxuw8ctkSYDwyktDVEMmWNAiXqw1g02ns1BZE525r7s6T/BNhnlCXoi47
fxA5QKsxqAtQTCI4ByudDZe6yhmyIzWhOAc+yI2j7sEqvxo6tfRU/NxDLZuNyD2UOf4f6VYwCClH
1kcr285vMFVaYcee/stcFZp+Dh6LTu6evYwciKpmLDIpgZJYOuPvFT/j4DLzu1NdcDNSap9rm666
JkKo6769Ggz52DZei44O4V3GrmQaJS485KSwmu+NuQ7WdU91CjEJAHbM/NEpYpOU2Tni+OjeHtvz
YZUlImEJZBhHonU5UuH0d9yveV1urxVg91PiaV+UxIOk1nfk4baqseYyei8uxTOKUFi0+wMvcKel
f0F5wrUMNrGfJa1CistCnH/Evw6i3DlGWeRI8lkxcw6OyskUMvquRN3+sHVASZ8+64+QIL4GzqZP
+TaHiLahOCKNQC//qiJZ3+6kdcFNXM5SZvkL9DPYw/Lg/rscCzWTUAnHPZi/jOY01UJP88O3eWXo
EWgz2VWbkKo6cML+bXViAEcREr8i3sGm9Mw7NFItkKzmZKjkJWPmfgiU7RTIdHP19VgBiNTu3O34
sbHibt+VI1p1uzo1jlZoTGayb2zT8hsGHiRkI9RDw0fiUvxGuY531L8dGaQ3WjJyd8sViUedxisW
dR74mIAZuc/I8NLyTw9jXQw1awMJ00yFpCgqa0XiIySITycsM7n4wBluoMMqZjuiQaHLwxDXo/eb
JS6848rzg/fEX80BkCvaPWm4cGb3vzlGcjYh6iC0jrcUE8z8znmhUjq4Od8LifV4uTP19A3C0p59
56bTRj7HYCg0dVkB2lZHzV63/lAx49H7bs3DCsQCkrhB8+w30unX2BCmg47KBny5IVBfGkwQm7wE
nEzIaatw/WE2To+0ueQCcbk6/uPNrP7lUp/QDvf2B+hCtRlOeQeXdVhqj9fQzzGBg31B0f//o5yR
7hB2ojrppcEIH/wKP5RPPrV+Hl3HzkAoYJGT6HvZF0HICr0IqvWejzVjZSSIV6WWfaRQ3w1Lenws
QMP3UXhN+DOiPFNHTebIWxUae7wa6d/tlrKTu2s4PhUHXni9SBROGTYBzkvLWcDxLLGovv5XpKi8
FWHQt+/00UYkcN0MRrDsEAYLyURsa/qWmfo4aszQzoYGEaI9Hpmk5e0FzMRqfr2O5lybQyu5E6JP
TGz8WaGWzA8UOSBzD2rHUVZfbAB3vqApqofuFaIKqhKRzgrCxMyEZycZjL7hSrX7iBOw25Rw2ctC
EMT5Mi2SEaPBVspFkikinRN0y9sNYGL2SyBmcIx7i1NRpxJTZKacEPagrOJTYurxAPwKbJvTvCqA
hnI2FF9oTxXWsZcXuHFwD1PMj+uYtb7BvLHgUDg9u6pp0sGhgRwBCAsR6wVaEfIP2IRw+5vqw91S
lt2w6k03nGAVUbF4W6+Ki9hLrHzPPSAz2nJ+DkeBp+fpwo6/GoedX2kaVkscJQTO3kBjWX0BKqsY
iGbXiZQayBjPPFhYg9lxytHpua3h14PCGn3V5dAJrPBEb2bEQ0QQKiCNHF+a9E+SxLaB8EtAr2Ih
uJ40N6yOYu3YjKJe/pQYFWW3APsVwzWYbAhXF2GsQ+QZky2RMYb3wI+hF2NlpgeEnSxVOgkOGNO9
xm1ARIFsjReP45iSmcYhAPtfAnkzdu/jqckHcINSAO7Vv9Lo4Y+3lUpkM0FS+PVlfo0zVg4xXx2a
DlmF+11oQGOcb4FOUAVaNOVLCI7A9qUbxDgBDK4C8ZxC/HgZKP+/8cQEXjX8xoNnSSEI0KP9nVk0
+9hdbMInKlJk/MVtugZIC6aGGWpDq+eLS/oRMuoOCz/wRKuQOlNZI48xUeaf9NsENkD9gFyU/dXW
OCyRR1b8/gQ5Cstb8tofLG7dhubSSdHMj2uzswcYyMYThBWfOvEzzoAO7iK4anuaB2aY3NF1SSwJ
cGhqREuf5fG9TPQQeFjMeKhqpaIXuJxhLUcj1I+VN4KXGt2TX3g4/bJD2HEbIYT5ehkQjBsWiKvl
Swg/eYrZ1JcB0KfLL5AZnxSTPF3GxhuPNRnSe3XzV6e5QLxMB3cpuO/sGwiPOXBzEEBsThylQFxP
muu5GCS0Lacfp73YdEURfbS9AMx+Lf6m/7PIiWFWFkL+tvW+jLP3533+lPfnKJhRoSRaWVmHRB/k
fm2bkYkviZ4q8EFDkXznNeRFJtvpQfal7VoykPJWeXxQZUjZLwxYWPo48hmELxX2v5lc049EwGUb
4JbtdozHMWRSDbdgOesibKv7DK+wlHHItAC8pnoJprjSJ1xVTn0sr/KDhXglgsyKWrAhP7a+qNo8
ijNUhrpX9jbNitqnAzp21rJJrm8sLD9M+rpgYOIwaDsTsc9VGO8pPpYBlXBi/xG56n63DPJ0/VAn
UWxjQK97/wifNibonaAb37mhToqSGaygXhD8ETIxezuAnGAzITEKZorwQi/3hUMYcW13uKsWljDn
J0Y8qNng6S655x1YXufjbyZEmQrGlfWJHdo0cStaLO63qz+F2Sg2GC/k418dqzl7kStVq1JL8xEu
ZGAsC0lDTdet4FnC1ne+oz9zL6SHzQXR0N0ZwAo2pGwquCyJdcnYHXTla6wCMhqcYXYYEWTItaeL
C1xgjivc+2+5ZJ6CUW98okUKNoZDlmpYLgrc84CEpCx16iDbHCiEpA/IMwh5vSTC/Z0mkwxkI8ex
LG4CkYKbDRZoABa+KOZ+Workmztf69MVoHeTrsCqOJera/oW4ZVYJWSIX6n7YvDqXPgA28i8Gxqi
/4rYJqICQj3rWkAn9ueV0eNCRuTXKgLkhodqK29Hjksvla3l6C03tRnQDrqFN0EHBKvwomjIfCRx
3uKVbCGf25j3RFReBZB/PkOwhYiBmCiwhRfdqr7Ma9NYFyaNDaXxjhPD96sTEPj0RdeBC7/7kxHf
PZgxt4lNQz9sdoeUc4rXCbW8W7iF6KAweOfexFKFF/71U7/MNs6vVQgQJPWyW8gijBE6nW34jRgM
UeSShiULCfh3O+f8uJYsBacNOPomrFbD019VlqNzLZ89vJnwDTcLiysSzUnBWIsbXbDc/EIAWCrm
Zbp5pNZs2QOM8jS05KPcY/iPmsT0SR7BQFNPCtT09KvlrnNS7J5ImTBgsaKzc12P7iSZiLDrpUxu
DT2t1JPIwkKTISS8xo8j55MZZsPZ5v8t3G/VIxDGXe9I3Yx4NaJuVfDaixHZrDrQKIcEzRHYl/Ts
zAsIRwEv8nQPlHJdtt68ijlwSxBpQejlzbiSdRN+eI2zd4ioezC5d9kT+liv77CmmktQV7Gl0T79
Gal9lnT7lGhcBP14k4HZVa/q6UHn5GUvP9Q6ftWyAUd5Kg2JXqICvBWKvt9MCpopgBBgTRq/Cwjr
0XdVLVeIKoPkj8Cc8rwUxcjrMY0irZOuSnTGwaUM3BSfdyGpCgWV6LjkJDs96iZkrkCGHob3ylMu
c91QMGQbkO58J7QxzNB6XhW8eBDHiH81q26JxgpfOeYs2qdqv87ApGS3FKWrObf6BYQp/3K3HypL
nZs4vPuuSBlHt6gKxqeUXnvXXsIFfEalZjtYVOdssClgSMkD0WX1779ywYktw4saY04b3+gUJbdF
HGSY/dAYjdb93twjTkZSI2X/EEWwP1FtlUZ/X1HXTcb7KlywA90XTsKn8eF9/6ZSDfux+MZ7Vsuv
CSJ+CfEHRabC4HkSNgPiujVTjzMVZ7a7pR8Yx6RHPWnsvRXgpmiS30j/hYoobHdza11cYbPkv3GR
tqBxS9BiPh5k7bzkPbXvM8c2F1LUusjAQU3qsjZ9Ly911CcpHxk3drxzO+bW//3C56+f4YTQFxQw
Tr7mnYSSssDu+7JZPuYKv93q6R8EMB8NxvxplxCxnEM/yZ1tuVcbnL+hvtvoq9wZUSgjsGDWExUZ
CuDhW17257pgeAPO1TSRY1KQK79riOEEmo19c/FsllHenIXNJNm7urHJCZNtpDziWi0blo5ywcRg
7WUbZzCjYYU7McRDabFDzA+pPZXaJn3HLEUbCc+vY6DEZnZGofwE51apifNePS2KkuwrdcwrarL8
TD3rKcRTgpuW16bU5AMefPQUWS9xqk2UxRIkWJMKJFeG0qE+fdZpnSe84/drWyaS6zo0GKfl4lvJ
nt4X6tFbOkRJVvR7qc7WTBJZt9H4KwwUC2fyuRTfAfNOcMHdVmgn7LMSEjqoL29Cx/F2TsEOk4Jm
JsGk3OWf+lAxuLJXK/tjAhbHabVX4UPYyPHNm3RI8yKSpMiI8wrtQ7t72gtvejKYBPIM4rrOSgTu
rh/9bGHz1RVuLSDo7sSG0/XLFoE0t/NcrNqzAOFfZ/hd/z9kKcK3eRzdkw8WwLt+8/RA7Uw7NlXm
Ag6FqQpvsGnx1EfZU0eUHU3U+TE/SqHkySmPeqli2h+93yaHhLLKVJNIKkRXAd9rAap5wNYP+/vC
0WUmwLQUGRfC2m8pc5sIKiS89zrvsAsAQoArTHBGMNb8s2VbRKGaDWnejbtfE5djO0bFOFsGxGeE
6OH6eF0p1ZtrNQKcyBw6i5rqUosxTwn8SDtnfG4e4e5XuyTJgP+SK0V2AweEBePlEK+qjOpLqco0
BX91apXL+P70LWIhbPCoPL8gj8lOgG0eEU1RAWPfXxY9uE1M3h1hCnGsyg0hmQjnZFXGjjM1d1Cr
Bh0zLDNb9DeetXxr92gjKeLDxFYS5TfpgR9JIS2nEmZ5hTnEvf6ceUG27aQACS2HRYwDoGc+crld
9ZADiPc4lKJIJzlsGiUDB0C90sw6FU6nRfd5TPFNq+QQ5H6ZYlZKFs8rF6wumat3Zv7AVEmhHRHl
E9YzWx5sD58ljb7FnSJQYfzqKrcX4/vRyMDqLKSFhDuFXV2wuBL4xc7zuBm1neyu011gmYeoP1PQ
YIbOTjGlD0QeSJPnfyN80No2j85oNQTrNVus7OTIz2eKe3aY3I3KyrU9gKUFgFWgrUDpl7kmhTjj
dmGszZVe8Eol7qqg7LdLrNIqCH6vhuqk7SbT+L3wgwrZxPHfaNMLrrMotLlT7+nwAuHVaxhAVAwc
UENPnCk/4QzgqTwtFQlghoqGJMzBSFckpkR1TQfGMR/12yoSeNSkuduv+crKJVf94UESdSzmy4/+
yFeS9IpM86YJirhwQPXTL45oLWoGlOEweAfmgqQJneJCwf3f/6rLeXr91Jmu6ee6bQCt6LqUNGNx
A/FpIVnwQWzF+AZudZGfPmrMD22xrVfufHJgGonD6gGnN/bvqy+5LN84HNnZyc8i3Yc3E8DoYTYf
hWPkXZiTdHJLjgV/SL2Q0fdoUjyvmOfu0Zewwlc5RvAqKW4Y3ApUlhmbVIRFEhWEOMTthj90zH2+
in/VArObGtpsNbFNhfkmffkIsXudbwaKVa0GZHeZh8VTMlsYg8GKTwAuW+TKVdQHwBgplY6w+VhC
SYllxa2iNSJw1TZOGPCXo+8bnfpinLLTWcLgd7SNNXrCX40myQKJJf8Mn7Sjk27KVnkAq+PFaouS
V1h82x/o9IqNvleXpb7nafSLl8rE2sE9EPDqImHVI9lP0b3OJd+7qCbGX1tUFSqOxddaC+jqwZof
/P0+kATWCZ0OUlFCCBnCNC+TfRI6NTsrpz5mlFk+WJsLZPTs+lNB9yWazzIYyxNos2zpjFq7fRpo
lhIzTYR2noOZ9Tiu1Wa3yhp1YanmbL61QeIUt5R5+JBqTTEHd2vyqSFD/yMBe4I3asziTKa5RgYT
ayZwR1X71K8GYfTF2xiSVG8LM+jzyTgzwoQ0kyU8HFBtToHFu3ioSJLwuCHPWLCWjPjzLGYNACrV
i7SSTbgA9YCtfsn7oue6HH4hVRrVAbQi5MjvqkTUQgfo1Vg/xZa6Ylixe5YKXSvcTHNy4d4+oWea
C2RwZkjR/FG+NEZ2jvN1iWMri3ReONjvPo06L8a1rMg+AjlwLJ3rS+JpqVZTfZrbH1nlEzJxsMTm
PVQ7ZuYE9J90JDkV31iK1e1iD0MkLbwfzrsfcGn+ZCM4OudC8qQ9BLWhmmQEiBeAuSCKmbWk1n3+
ITenjp4X/IkHDmdFdmBBeN9xFPVyUhtNTskrSUBhptkc4xvdVdzIUIE6pTBolp0+jst2BS8GmW40
+hQKLEyxemogjWl1Zwe2ydP+X2e8SaqClgEypOWm+2b1BvLYcaCZWzteSJxPxs9bZn0bN0we7nYY
42cRKTaW/e7wUrDck9Eyge8z9zlTsrv1Memet1TYwvKsIF9ejeavnuAAMEf0eEMHRlslTskK36HT
k9eA6EKagnxxvt4FIwMBrHh69Y8ZGzLpyadlWr3kO+Ufpmcm2Dtcdv+92RP9bwxo+Y2yV16amtmE
eXS9qYLCytv5fae7mMIsY/20/GXt4L9sdfJ1m/6/nEJIj5zLzqD3a0KqCfmEdU1aIZQZi5rAg7RQ
FjbCc4pnroDgx6xR4jaLxfro+AVjtDA3h9DCNxDO9pU9S807w7iWrHc7/1kxESDU8zTpJ2U0Hyhs
xbHPi4VvaLvprjPkwbdOt4R2bz86LTwrECse3xYAdkMJT5L1gcV/1dfDfwHHGF7E3rdBkT6UHg5q
5TtGWRQtdpcExZA8E2DS8mmzO+UGwVXkDDbMUhe3fPMsPcm7NrzPJA1GCYDz+if+CpAFzAZAS8YJ
sJpYfQjg3N3nxy2qpBxi5Fzdh3EZPG6y6qtUs5pSUoIGgQ8IAEsGB1Kj5NI/97QwFWdCoWUjZZON
fvXwYy+PD2pX+3gVf/72xkHJZX+4QhL9eG/D2m/B4IvPKSPhgRSTJA/w1m6C1kyhToGFLW+MpEnz
ohyYLL87flQGqbAyxq0huqqK0Ti0ylL9ng1FRZAUPgBhn9fA7LTAJ8MgJ36RV2z1KjCnbPLcD8CD
Lmlica0DpKjtlf1DALvFgaTK20h3E6DzRMfwKKG0dSheqJbmd/3PQzSx5HwH0eqcYj+E3q7TF8r0
eFhjpvxcS3pTijvTN0X+ZeyDHdQMNJOi6Yt+sCPpT0mrFqv+/PFjIfmeT4HcMapEDkgIjM4lNA2j
SrNOaqCATzqHWvM2k2nEVDNVpn28GBpuH9PRWwuDziDu0zMbQcLJBhbsONMbLukWhNHW8InAcRZW
xrvvQBtq7z1CrKiL/T0GzNG6aBnH3+PRreKDP4lZngRF816u8cIWf65a0gpDGvbQS7ZclZAToRXy
uPUGQzg25pikAaTCnFIDgkMNEzR6E192xidE+hJzrKncdjAizOQglIcdaWKzhKShyrDXMRzmTZ+t
ARWf8sBzxPspKygHY6NZBWUZY8sCiJ+ItZmoTJcMlm+vdmMsLKI7m8QBhNOTf9V8Mglk12+TPYi0
qUxaSUcbNNvoUXqwkppk6EvVxnSeICuMKaZFXtHuJ3R8qxc3lyrmk7Taeh1uTFtsYlW6x0M5zRa3
5Bi2VyHFYnPSkxtQC+XMoa7Ml7ZvMln1e4dGiwQflQz8mP8dmQqxeroN2W9WejxrY5gXrnTkGbUI
Hc3pDDqifHhQMwJlSNaIuTK9qJdG+hnRYUW8TjKWwSLW2OlBGDuXzColL3IHFZ/OsFWxPjkLucln
2VZbVCgrq8jYnqhH90NAZMDCYSB49d24+4BdGTM0Hv4cMGodgegbTSMdKwq6/pufHoIIDUAo8OJU
QTeG61PCC6H2VfNSICETYURL7dEArOt4ohzVmP97834mrIicNgcgVwODIeR3f90OxBUUw4eC2hHz
hwdcNmjRNqYKIU7N1vKl8msGU1va4uqTDTZ17WOz9wUO6Vuccv9ll3Lf7wXkAwQM/774Qp1Ul5ca
IoZ5LGAP/F4L4X2LA9pvYnryDQYz5CncjTYH7nvs0tBB4JkPM7792p02wFGR8SlG/ieKlBl6+Wsw
AstT1Wf4xbSEdYunVw6iI9y6CzB919EYrcn035ZvS/B0Ry37ZwIS3N/Z9O1CI23BVezwW1URMBr7
eRjoWkApCLoIXg68bMAojWnhHcF3qAltyPpMToYF0F+iW3x0UmYAJZ4W+E/xxuVGBwHmSWTHEuZd
yjloHm4odzTkiFA9VVHUjJVMxuQxpPHAl0grve1L0AYZPz1U7UCYXNpwj8mIVvIKTDHsint4TB/i
pYgc+47hs8ZVhxjS4OWFRftQmrFrdD6/OGWfZofeNdxjLwflLu2OskS0V4fQ3OECknpUSgo7ZnIH
Gla4GbdNElHC2xjNlFe3A/qmtOnvqTJFA/Opq8exc+QcckHX5ZBzJw4c/GhdI2ZfSeLqlAye/NbI
MRNuTsD6d8DmOGLtorVR2mkNC/vCW2leBq2cLE+kPwh7h9KU1C0Xfut44tV06fLPgSPlBBdEAe+f
Ncwbpyx0vk5R6rzoVKTpqeL1oG5oWl7ZLB6RWdMCkd7npXxgNiQ1pw1yobaVKbQY8NF4KfZrzLlT
EzveEcUVpbavErKw2GL9lXOEihew1O19JrN25uh6Ot+CZOwVjiu3sa2DpVUleC1rOIqa6WLD9XpE
TvJwF6d87zCpaEdrzzEfSejWCdwSKRXF07saRBuaqZ/D0xJvr943qI/wC9vft5UagV5ZK3w08mVg
NOfW+gW+XOy950ZhXNeex4yak4HlGvUBStbgf5BE0HQMoZESzKWcGD6E1q9BDQWNg98QJ9S6yh31
lwMURm9GsMccsL7qkixPNlTtDGVhYYnmJ+5YxY+moS2izY4SHE+Ae7vQSVRCg2QAPN/reKDm3qNT
PhCu8XwwEj0hPTvy6treh33f3ggso0kSBvdMTnQuRKe8c5JoYfDjtVVyZklYB2PphaCegOn+OCNl
8WB9nCcpDW3n12gascebeenSSB9KNbL0cb0Q1zncwVejRhyjwM8t4tXXmRanQvGEG03dIIexiZ0p
gBwF4/XlRQJmHK+To1+lVeXq/H4TOWOJ5MFDzXRVqj5nx4thmq4g1x5oFCMYyb9bIeKGUz5u8h+O
Its2iqolkmFNWrjtniMz7JX+juhpxcSD1RI/dMWysfUzPh6ZpCm/2Ayw43lydkEazSXHht7U/KH3
B1FquqsD4L8w4D3J76gOCVeHgp72fLe35zEDS+lfft6KV3D5z04buWCm7RmIKDeAdw9jQAvE95Pv
dhNZHPrZ0rBbLwbAS6mnhT4jFPn2QNstbV6CT5qwwA6FTpJjwo/3k87mPXmQCXTqjN7SVvt1NSGK
p6rsS84Z7yVm+jr0IiJOfrvo/7EyhgxC7zXMJVADA1d2jOwUP1Q/FUwBByXSLPk8rcQfit3bDVe1
y77tX3KOxTc1vVWx/oWIwdSZvfCaNLGvwTeY3FcYm3tNJoYtwsSZthHEnWst2U5+g98vudv7f9hW
f1EYHI6XjZOkHHNMKzjbtoKnS54BbeiRomrveNGLgH49pPZ1t9jSANblj87VoWRDG5zqOmwaMcmV
3u5nur//36wge6jp6yKdKoTDhdkcjG2lD7JmR+A7yY5k73bihJrYnrYU+6lx9kFlTy7c71b1+D/h
imfD6LB943rngSVz3LmkhEm/6N47jeUmenkEVklPHhzlkpBEVJz+QLLrMOFf0FXmPUrLHPEEV0BU
8l0EKR5jR/dos4a67nBInZfYdWNa7H30auIFM7+njtbQRHNf4h3YSNCvLz/QfmGcDvK2Dj6AwXBT
HFpZ6xU0Wz9Jc0/YwIC8hOsfaX9s04ZCLt1ZQ6mzdpHJVsl8Ibq6Ktj7PZRVhrwM4QE5eM8Vndov
BJPQ4kzVZ+OnKD5+srN6OaS9C7jEHUukPkziwjSmoYNv+BgxpKwjQY7bt1HsVF6ilH3Ud8+ZJRwY
P/50UotW/rweR1sJ85flx0bgPJywDVPPdO2GButezDC+0gUoeqdy6YpmCvIJ2K6GuY5YHrJaEH/S
7NPaNH4WmRwFvOOgts8+dZmnQjBM+mj/o7hSvU0o4K2YbJ+XPcS1zW3bDoalfEDJl2J/ac8jafwF
IUZJ+bYIbfSL27MozJPZm484xQ+hS5wfVLr3cK6M7dtLaxHR+MHq3iOItK+ptC6DejfkjEsezdlI
fY4gnaAd1N1JjemtGHZJamQzvEIpCpVlWmOtEAJZHuVdqKS/avsulN7PBmVW9/7/c7ehy7Y2UAdk
GsWQaEjNtJk+tjWvBTwudmaNt9fj//WgIghA3BA4TiTN1ZhhUKYA4QksVJSBV3uHrHIDjISlXzUT
QJNQ/bvITTlrDJK10Ox5cGeYBna3G12i4hx6gAX/o6d+PmCSodDXInRZf9YAaKd12Bm+h82j/99n
5fl+MvKhzNYZUbRBPFZR7TXAGQWcVnru9EnIsD7LYSMrkwvpUyXPSyVJwKVXzqv5nb/Lz+LlwZU8
q1wfL+eVIM5JGNFm8NIdXdEFzq2Gz4y4F00gDLayq+Rx4ps1uloBwEsSuh897LAU4fj/XHhRMg3n
wpP0vHWsxDbp4S9bETchQwHvC8NsxyxXtWBRaJZLUOu6yarhVJpP66hLa5zmiluEV3fySp8mO9xm
zx72qQon7eekpOmbGCNh8vx8U9U+Yq6p8dR2NKl/xIiyTPsnYFygOErZwzRNS5P55v7NYmRs4Q0H
03DQJhK27jnAQaWT8C+M9rtKc44cbIFVuMOYbuiXjnsbxWXWmO57djFIPoXPAH407fMWvIth6iu/
JKKRxqFXefVron1JSecBYGIOAOHoUZKlsO5MElo3cCJIZNNwATyLMvMf0AagTC30ufRnpWS/vNhd
fbkDSKUboGulLok2rseRQlzQ/tqA1fLlzx5otYk5AL5rXrG0pb3TmvDG+sJoFmQNHS0pp8pQOAPI
ZfyD50wdztijvm1ZDr3heV2LfN80TVwZTCGJleF2mVhMwU4QGPQwssmdeSFe4cqJ1Ktjrq6nRv7m
RGo6iL+QwnW7qwb44NPBTOJ7fABhLGRDJsha1q5sgY8LFmk9KFqRg3FcrpkX+TqLz0IVCHMEAxKb
zr9FnyJO5ZCJoTXhjWZro77p16dHP6Kd1YEKB0YexeZp21l2tS0N3NGeF8aooKlrDS+ccnKXKMHd
m1Rl7ATjsaWxT/oud6Ixd23mwQN8kMf1zhiHVHnO3l//0UVmmnECy/hZyJj0Vf8j4X4Re7e9l9UX
6EutSEZfoIffVEDDrMwbg2WoptLzo6mxoSMV91nX1VQH/n6jj6iMgZ7yOihHGXpPiuvryS1+dgWU
5dFqYGOXU3fRT5zodjqdUlGLl7hCNgDOE37CZg/WljfIKFvvc6INHawwmcN224uFJ3ZR0O/PtKN7
JQpw62iiicRvL02K5tJfOp2E2K50xe+JG9v35CGQ9NI2zKoAQWZC8vcHqu5PMt/vR7W8VyosxhY6
qgsnpQlKO14gZivC1hQSwsFxDbTgEsEPzuGDm5kJYNC3sCz57DqwMglvSoERssW7fUdATnJdysHJ
VbxBFYe2f+aAaYBVIHDvlPactVZB+LRyBS5Lb0Rc2gsJfNkVEhcuRP+kC88c3SQaO5s95CSde/UL
MMWvsLWROz849vnv+XNrTGPc3dfVFC60BSfz8S2YGOMkvA+P5juQC/LFeIORDb9TAwE5C2fhM3nm
ag79Lj7tqFsZeaSp8RG9hiEvaUQa5z5nOGMbC+3OU3CNQVIzwLIhuAi0j8SDwvRi9Or3sglEawdT
8swJ77THdifR5llu/aoepV4BjI/nmlNpLHSu7yhMwakyanzdslIenUyxng0inzM4U6dAiMuL8bXX
hmKPhWGdD5IS+6eErF0b/bq7K/qQTVuwgJcB1HF5e0gCC0rzLGoFupqmb68NaPmsxCVzME03Rztk
SmfPLm4lEz5pp2LGdcPyr33WndeA7PrVYubVYmEvgR7W5UamW9wmtmOHzovAlpkFgHz+lPTsJL2P
ZOVi1wcwb+IAGD8BmEIRdesbMK/0LlDjrquXcw5RQZtnFauharlUV9bUsizJJDQd/6q2iSIstPcK
JVmekaz8a4Qqt31JPZ39Lh7GCqrcYXtLaElUTw1OSye02beDL00qhNE1tYO4J3CVNuABSazvECDu
8ovQ8Pd6baHcL+qBvLeVY6oIwq5M9G6yK8Hnfd+g2pLe8MEdZl2pR0iNuO6358tFHvmJkePw5O8W
AhLAR1sk8P0No9k7qIJio1bQqw1ncyKJrf9iFOnO4+BvlivivNSiWGWyLcFShGlgl63KHTrvhHoH
olVwXxPg+0b8iAuprioAVAvftebQ+AMRFRAZdcvwJZLVJDwgaIAwyzbPLvtgOsajFslnNafp5oYc
rMnBUPtG7ciBCMye21/M8QmB24doUyeT4Bpw1aximwSGK0QMTjqJc04Bo07PZ+qZyMIGYRKZhYtK
tSYpCpGNPQQ0ohnL4XqJWFRnrGzSxO2yU9rs3eoiS+TLuDDHmldoH81GQFNchsNcxxTFnDRUxNjt
DouHmVMpEx8cCkWr/QRHMnznHd16nPgCwGEufFUf9mrZ1BaapqPc/67jk1aoSMRyK3CQIlRMXap4
1Sae6WJ5CoS++hU+ijCnH6AKg3r1QynVU9GqiCWiCSH57Ve7Vaz1kSgj7DmOXra0qe4DSHXi3fV4
8SPRw+PMpe5wFis6c3ntmvgqRaqsZZCqTT1+DudOIv3SeToYPQh7dAnrXy0Xw9ShOsunUWEkgksC
MLRh+J8CSEY/2J+ZaeZFWalhHekeFNDoDxDMw4HDZ3NGPu0XmoJTF13XwecdCMWiAGkvIEPISrFF
sCCQD8tNXzFK3XHvwcIO3ehiHzSFhChn08vx0OpCcsef3nzUPW7ARE9TgoiCl2wTOSYJ5YQRDXXp
IBSH8dfSoIZ4LWeVNQXbOrS2adoZ6xCsLj5XppNfyf76PZ/vswIrmpDvWD33PPHA9IDY/DK+vuix
GWVpr2j7LY9Snu2WvQxABKx7EXSztxUGxotJmAbMBZrb+Su9w6lBOMUzY6SlfldPOHDraKoCmams
4rpUq/j/sPSpMX/f208DdMGf+oDPqt7bGR4qlZhDlVaay+Vgw1sj5s4OqpsuYOBXpjA8Y3JlVA4Q
RSZFFXAygRJCKMtr9eP3qLKbh2IHO9AnpNuamVS28nlBiLVonDNIF+pWbHokrJGGzvCDPiRYfxFI
Cp1don8pZsN5XSZg68cop2eOTYYzScLqwDxHHp58o63ak80h4B8XHY0jxqXYYONhTPxbJ7xT94cR
dMgBH1OOM0czMeS+vOmxwKDogRVW76iqPAdKo/2kyFrcmvCLAH55DWxx0WvB8dyILLWzN9YI/jA1
LCUH2tHm9STro1iZ3MRi5QmH1yuL4SU/vaa5+Ri3+sQCwlRUZ2Ke98zXVOt8EtP1KfAuszhG0X4w
5/z4zz1IK5DhaxsP1yQIGXhWl25kJhjRJ8Q+TIqNc5DrXQY8s8o/pT55CFh4lx5aySOhKoL+M5d9
UbAFmV4yju5z9o20vNyFvXF5xOlj3vBd7qCIXoh4dDrMzQoPrpIMd8l/7lr0O0FPvwGvZfBfrMBP
25P23OfxOyMDI0vdULWcBn7TgIWEN5MXkOc1EuGP3/3XfUMCfHfERfg183Zh8aa8jLZeBo0eTSLD
kX54ghMAs+AHKphEXnvp+ZVSHiXxhYiLCmFD+VtDjretS05Gmlnn9fzbv9/NPu4mP/Z8LlYtZTF7
gWgQ0z683T8pyhOWgFpwt6Ud74JwEYj7OFXM05Vy06my3H6pQmlI7he+nYKvMPHA3mkzsx+62BhZ
RtdyNvvT+7nmElzhqkPqHQoHLWwfy9SXjBOO9ul4LwJf4RHqpaGaU2CZr679vh36IjC2prwz4F/8
njUZxoBz1BqohKrTCZ2RL/AXejmj3/uY+BM73MJRqRTYf38G4Gdh8OGEFVft9lIO0AcaTOnHRoXU
z0L+7wTK8ZTZTl3/RocfAQ6clLdSwgJxY5hEaTKn/t+2rOCpfx6qfuaqnt5HC8XXu49UtYdluTQx
iOG57viNKH0usrnMXUDkEHT8X3ZoIAsLiQyFduiyHK9IxdhA85Yv9JpkjA40bnq3G4nKdU+1bVmy
z0PwbHgbE3u0M8BYAN0wNGiSTfc4zEiAwv8tx+Z7M2B3pnHurkxVjAUAbPy4L2A26+XNPiH1lID/
pf5E3qfnERxJf1PqwQ2Ki1ryo1UoXEXBzIqSOfybDgg9hP5IidAkllqdvRYzOIPFymbad1h4FX7y
c0AswOJVmnHkOE54HCPjilnqdNq23Br1UUZH9/bqTT1h0HijZKpzrA4J5jvywGS2LKquTW0FQmPO
ABcpfVlcCIoqUBuzRt8GmrGOVLp+z8OpNIjGQS+xVVEYAmYTFcymGBnwGleq/ZJoIwoKDeD23so3
eqXpPX9Ig6SFBSxDkOALjoe7YqhaJKWhglMOBUbArlgueOGJim4x6xPZa/AR2/ZAPs8ePPIkH8Z3
qJhjop1dezeTcUwkZoNHhIGj6kNICpUcEvyCw3KIetcijKgHrrl8mJ+QeYEY8zWFSSQwbLjrWbuI
O980bBlwDCcEDNNNg7ibVEvPevq5KpVarbFeCBallA2vRRIwBSl3dtHoC2jm2EkiT1/OHIi0IieZ
/mcG7ABHuugUTJNzpB0T2e57dl7+dNfh6te0ggKFKEfp/9thkfm8hho008fmWz38SBH7tZuI/akN
/K6hyLUXLA4NIg3XTkYURo8G4qseEdabUyu/pooHpE8pe1BnSa0LBD9HrzvyOG6gjrGy9nwB8fpM
4u3ee90KSOYVOfagm6bD1XEvnawrHofZ4oTh4VX0ueoWpREZrqiEKElrzgX4CiLj7yJaPg2BNMb/
86i4RzjPwRTihAUvf6nSxOfNIoPgLall43cHHuGIaBSxV3NRUl3Ziz0dE5NBm/zJOUDtd2ucS5JX
ZXfoVi2qwDLZw/AO++/q0AGtGEVB0Cg9qe5JRMSqW2Y99p1G4y0J0DTnYmLK7vTtG5Nv2wFtagqh
1Rg2k4QjbB+CKHJyDdVHsJ/hS42bpUV/axGWEzIt4KDjICe/+NVlrT12Tbn0jMCcOdaDlkFaaZYi
IL22ONGM3tqd5D1JNAD+F36NVCzSAMNfTf/lnOfWqxur2NnI4Xo5BYAc9fyix5KwcYlGz6fDLcX1
/MpDaFnt75k/bAMvIn6DxYvwp8hNkC6fRLo2MO+wGp2MWZu3f88uwg2tuwo93Vy9XzhwJoZT2siG
4aEXGuLre+K5TxAnojnoq+U1wiaswa9z95LUgRtzIo7SFrV9hV4c5Vm7Epg7ITuDmMvoIRaMCmpJ
4uH4zxDWJDvz3/yTokSzRisQV9XzST3lkqVydOyzQUmaGIp/GD2lWy8h3CPXEYZy+ORcIvcnAmUq
8M2GEKyymPkLHknnWR3GxOyvAzJDmPTno9MPnK1SgD86dCU81dgQ1AHmYvhlB/pTLXRbpBTzRb9J
sETfJPjp8ye3oW0iKDtUTZTcEhN/94n4Ufx6Tvkx9gTS2dsRjO4ovFYZLE51WpnsVuBk5JmFlLvX
qRcp6DpySPrLSRNO56xht1hPSTTeV6DhTOdOnfWCAC/3GlxDRmHX/2e0jwZom7DLuAHRTxo6lPbv
y73Te/vxCHvI4/sqvxKzJCvgGvtp/fyZUL59dg1dlZPBKQg6LYy/gnCutEpJ1MiBaTQ2B26niNld
ihqK2tTOXD03zxH6bTnDbkmefWDemfottyqkF+HsOgnrfBC9JWJFdUcQ3ewAt5anP+P2W+E1Fd14
CsZ7MJSxrIHX9xgpghAK5AEemFT4u5qAG9bKMhFl3x24oixHF2Wf0rdL18uP/gDgiaXpd7BXHvbO
VMSYhfmDFcGd/LPoiGTaoGjV2cJtsafXjaHcA/4bEf9En22jkuC/WkUWoJDQ7zNOrDr51nEmUKT8
FQvNGPyyZiinAw4IKSyhMwyhIh6XYZ6gBKm+XlgeVew7iuSHerU2avaO5g1osznFexaOQ4LcBtKj
v5EhwKbbssOlq5wITOrQ1ycv+R8KLAzlcaRpnWMChJhapV0cvvJ0V4C8QXn8WSBpjMQRpy0SOd2p
Jr11bKNhElgQLcvmSuBwG867+TewyrEb2jaPQ1VH9qsd9zbSCX7W/HtuvTfwxacevsNWrUszhqSS
PthAD4Pq5N12zbXWK74+YjZ/w17uUwySFCxnSFNYaNVYXrlTVCYVsNpA3TzEznRsOiZ+Zn/pVpnk
jXxpitaRfPyFzqGC1xFrBoJpsaeqt9Ulqes0o/i0fbFqn6sodAW/C9Xbj/HsSiejwGa6vgSiV3ZU
DmN27eYfe+qZKAmT3sxBXsLUkWON26O3PuI/j8o07kC/VZawm4kUOJktKEztAfABJHcLPQQ80HOQ
ZJSqTcfkmVqH4jbYhg3CW/iBcvgeCKbJ7KJZB9tZmIt2DdyZACi/p/ozwGzt/IifXxeg78fC5+vz
/0WTeg5zU9EcBS3VmlDUeLDZIfjkBXEDvGMJV9a1+XvZthh4laqX0lFdMntDwuTyua8n3Ej7liuN
3aISjFmCuri43u36LABgXPqTkKXfIuUB+5VC9OaDB9CkiRCNclBDRB1IAfpW8qLANaa/O30JkXNr
7KgONp+wzAQLfwPEmLpSMvcWB03VzHC+xZiBIkR+1jhEJT5uq3JufZCbARfu3XbBdFgNY7zgX9jc
penUhnzJ0m25jyx9ZP/nGZamne1mr8rRtCmhTTvRx2tHfedXJwRgv4hO7oiDU5hDHGdozWufaNYq
efQNAH3YYRzPLH7YwPPIFDTbpsivXuIrLWQMKjN0QTuBZfVdYm1bKpqCRAMq6J/OLb1KckITXR5f
ydIHuRqMCUAK013k+kQKMYPxL1noa+pJZELu6ZjtkIx2kPcuNSyn1MIcMlhmTHZf4rAlxDuUopNB
FooLRpJQLBdn3CWMkRPbeqf6tF60o9cCMQ4w6LV9GrSR6uL/lbs6mT/3L+7u0B2Fz0kgMAGuRM7H
PI+ntiilQ/udFqTFC6PSuka+c9fX/3PenBInZe1+1a/QVAwXDWnD8vT9azIpi8GNzLJjQq3Psfhh
7lSehPVpR+kn5J6Q9FXpSQ/JtDw0wmlYhRo8RO1LyxJbOpLY1ysqll2ZjVaFJxaZdt8xGyjVWOr+
FpsVvQg+AXTde2WVjS7KU+TFeWBjlHEmbyROqKcCMDn2e0PuKd6f6V9n+USbwXlOKAvWgae8dsc2
TygOoimUVqvxOIQCnIGE+UOBqq8EhhrO/yE9Y48B67lnSL+jQyNpUWq7IlGKF5sasNBlIsITBAdl
oPeg1NvhEDdPY2LULTqvPQuo/8USQD95Ji1Bh4K9qJtdrSBQMa8EsvPgSgqxJlvOV6ycGfMj6LVa
yRad91Blqh8dz3nbJPM69mAlK/JIWz1I7Alz/Eou3ILHP9l8beIBcXZY4FhjJhEGnrA7MbdSqFK3
2jQO/+HjXjEZNYelU/IGuLbGRV25rCqRzOKfc1FiG4ZfWfsEP1dYPZP62EogxAZgMgFAjwe9ZgoW
mhU/D4QAYKRmAR7Q3vyXKJY2hSwriV6npoROpharl59TnNo2atol4pX0bEFyFJyBMxBNonxNLAku
HR/B912DYNWKovenHPzNqKwJjNXvyNjqrmFxzzCbPPxE40C2lxLx2NexkWLbAJL7vSC2SdaQXk/8
Rp9ReImXxLNWcp68mfIojtD+ZzzemJoVXG4KBD5Te8vQEyvww9De5MVJkWKsMiwD+1JTdnnmOfuJ
3bBJvChM/nJuB6sBC7p+LA6Tm7Nc6xYVyfwKsfmB1T2G0bOSd2prJP1Cdml95lkrdVGJrWlmkowH
Ni25cDpKpHdB7ziCk1a1ue5/C821mChnuGset4OIG+R+Joqjetn9aVYNgMV9HNTucLGo2UPSPshE
Cijwu7lMpnsIdI11eVmwm/EfCAY3oSA6E22NcDx/XTQRaZz9dxekBIRe+JcIH012Vrb8UPgIYLgq
RfylEOIH6cdpmwfIFLWKV+2NHZT1LsXOj1T/JfV+Lbvio2MPV+yRUNUubDT5tUenm1o6gyaiXUvS
HeVUyq0rHAuGX8nRde0yv3IWALTbLB0FquKiv8MXnGtmF1Ppqp016GK+R2p+rXRAJmOgvyr0TEAv
iUgTRHR8WCgF3RTcZGomFF7c7mWVO6FY46YNWHGNCdz6TSkIANWSM01ckHls3VUID9FG8r3g4Y+k
BUlh8HlafZ0XH9a1v5/eTCGO2q7/aYdtN59jM9tyhADlAY5xtPdCNRvnvwBzrCggmYdlEvMsrdsU
TUuOCIXDB7sbKTEx5qjSLekVlZHg80fd/l2Rt2bjeKue9ywqb3Of85eF5Pknv1s6tKNemSuAa33A
yLfNhQbVFzGPWVIzOtoDFpOSR9u8Oto687UZt9krJOIREh/Kw8XK+YJNXRkpqVlAz9Is5rRQfMdq
v4NF//CubPsUV2RlzXlB4JqNMQsZLdQUUh+npkGJ63ajmcdfuE9ed/L+am54nx25MVLZPZX8sdIv
MLMgiK9D+a3q467eSs+JS9JwUERD8OzmPNZH0O4/1mIPqbGuH5amfhv3INznE5z9SHrPEeeLmsGP
5EkNMhWj8kZXT903ry3TON+HeMM1jKo0IO+/7kaFUX7VRVp5fLu8n02fedgAcCg47k1obBXuVfQM
g8CzLwMbYq3GQMVFWLI66PDXDpAQ6ErToEKlFdSO2j+fhezKyEBeHuBQpey9Ro3QBGo7hZYypiXk
d6jv7CvpHP9aXfx7byk7C81R1WF0VqlQTgIDv5awhx2RhKkeg5Xq6Q9QuvEOydAEA0GaQA/TzEB2
dcbYP8VfIsf7QM3pCeJwlN1RLPg/uOl94py1YlNPLxSVzZ8ChXYpWqfm1OwgKj1fLvZ0PF33WCgw
ZbOtElz4Xv4cfClPii4o6vGdn/fBf+9ctYEZfXXXh2HLXYMzQkiQp5fOGHbHUiYxVUQLXgdaPEcz
qdx2YYNi+seEFRIqDDGj6v/EZcQbhT72g3BSS8Sj/kYhM7Fzx9h17h1cx+blQdrgXlcOnbchZ+9h
omob2K6ANSO4e+FHauMIm/TvzIroVZ35r5Y1nz5nL3QXHk2Id858nsnIsIxDFsjNkmRfXr2CDmir
qjaCIDISeLK8OqVEvPvoKZVDetTp/BvUqfTna7JjvmeFfDStSoO7EeOf/ztij+pAJ3WdObWSDeFS
8TCUDJGfGVCYZUyLv5UFaJJboOk2CVFX4yJBuQqVzxVIt7eJvhyyKVepkztxU5NHW2kEu80W8TB+
hlcgBRM8ce2uBmZ2xxNGEmuw85pFW/DGY7KH+7GgGdgtpPq5rA1977gQQN+HrVUU3bRU59ot83Vv
Ib6Odm1RtVeqnuTUMzTTGUFkpf0DIlvkdLV37fzEhfbuFFh6UIcK7rpKwret3h+o1alqhpkvnB/y
BNUhCrPz7XObRpF5frobbS89C5yEHMrOk9XYI1B3UYhqafudDtGKX7xHnoJ/goPaadMU6PkxR+Gq
Z8VH28ZFg51G7kwJdNQHkVXhmZ7Xbx9iRzI1tEAzlFw0t3GUs/UjRpvYQnyfybeUs40rQcoc/7kO
XNd4CBA8gh7ImsAesPFt+njJJkdTNVjzD1XNe/ex+RO6wp90CAYJ+rbRpSDZ1ncg6sRV16tC1O8I
xmWV7GnyguMLixn6/3b0phfItVSQBNvQUvWR5zqEQGplCMPd7SBIXSXYj8ptmDnVEnqPpfKlSLl6
ATOqlrglhraYS3cruhb9fGS8VmmxLsVdA9siwr0jMFAC7gpUryE4cnxtyqFNoGTd3IR4shoIRQXN
dtFwEJBGPWgCu3FiyDUmt8AHGQCv28TVUyjPzoGmMpTHJUwNtsehudaUTTACJaEvooHTfvVrdOPx
p9wPWgKS+lc+2hd92Xqw87WhrHQXlUTEOo3sbh1zjVjlmx8Zs7Cx0CtUvihb/CP7SDxUBVEhfURA
Q045Q6XbWa+gpkTk8QDjZCR1gbiEvJa9YWmec0KW/TolMGBb1tzIQz5TcEi43h49TS3Akc7Qjn0k
e/uy/3uge+d/tJyFtZOnt9yf6m90a884Ow1risM9+3yG/nd7onJ1IftT6DU2jlyk+Ig4qyizOKlr
F8fwemwsKmrAotBeiouSeaRFFX5XmWFuFX5uvOj5wmHfm0fSLUrYcIPEc1PC7l60Zu8pY0WU/oG/
fzWATWFleqZnmYsBGXZjJ48PPpuMqJT8Mzheh+y/r7mXVkSieqR7kcpRNm+z5w4mEllvRMcHpXdR
S92ssl5yFrZyRVcwwD7zFYAbQaj9OY5gQ0Apos+PXjlUBcxdT3peyMyyl69SPmvXj+IKrPkLrkoq
MtHQFfbxr9Wtz9VqugXDKdG2MOV4OglQTBF/m6G3mmEvplrHm9CuAQ7nKpYXIjbcYORtbFhJdYy3
IyBvaKMPY9GQO9iyHI3BNEAi9T7GECYsCdRftqcaPcyz9f5Pq5/RvcOQtFuSLY0sYNgxqwC4JiZZ
jXLB06GtZzoTDc3pVpkyGRPK/rwuWyzlpOq+PdpiAf6bEGpGohkFrTmT+Rol8fuHcriacFXz5aO2
SHasEoCjfcgR8hAWiaibwT6HCC24a4bF/I7q6iCMdqS0zPQq5ePVEpQn+nnLVYD6iH5rvpqS9Dga
Qn2E1IhBgXS4Du2tyP+Ko+rOUauJ70L/pRGpfnwBXxPLZU5EJTdGYxg1yrQCEGaqmnd0JjP+G4FK
0zqsHypYaaLTkQMzZuAI2jNYpONtltpadryGeJ1UroXBdukU6VZ8dGguJCMfRe4Ggidpcaxg94I2
unPZhjRSOrXiK1vhUT9whwxYFEZRnpXP3FIptXBr/PGHwwrwTZynN9sCXGtj1LQe4WypE/vAeHDd
kC/VNZMzVsVSmGonyZLIZckV0FQVKgQIMwm+6+Vut7ESGCuXjsg4jUWDUP3DYNfLTeS4c2E58STD
SyiC0VRnYXVChhJYKWnyiuVJc/0PaIozIbPk3JZer0nJVBU9qVDLTB8uHdnrzmFhtGv85wK0f1hL
rvicVarkqQYNbjRrkMsDGYTf6G3oeMbN6yOD6MwnRgP2gK+glHx6Xg+5FU+vT8TsG6tv7QvfWa5C
rJwdwetcweXNCrnFuT3pE1JEtHyDfly+a3gPLzKTPswUGZYSey+8GnTdZLQ3HeVNf/Gdd7oYBQ5Z
7/Vb52tGLJp7fwoHY1kPlqxPWLVulnd9Kow4lWUBbpXAU5iT1/SBKR6bXTpsNQOwqvDsQpZh2iB3
FhPvtM6mmWEhQnxiqz/wNvU7K0QZIL8cQfNSUEtHRnFtGsF/zMWJkVsZEN9v6gB82ptLxm1HRdq/
J2rQ5ezasIGwYX7TN5yGF4Z8uWI7A41Wv38ddZuMulDc0fsRlttSklS0/P/+q7qXOtFQPv0E+s8j
4/Y6zY0bemFjXuOiO5W+rDsGLfT0ZdZm8RDbmYtbJ7wXGGiRHTbRh+0uGIhnw7DyTonnYe/iHG/O
QX8GoM7NB/T3P7Q2LTq3ELhS2HHRtvWpCZ529pXjiHx7Odg1eV60vukdOgk7/JBkokbG4Oc4pIBP
LRSu50JrOFwcuLoMm84ADYV7eh4mKFCJxV36Ac7iSGh5g1nExwJJccxhN0ngCvvsyM7msITnPNrm
Y9pz9uKfwofDPg+JBh4SEkLroq/1tqiMfdXjmrx5zjZA5O7D6fDRkRWs4r2HBV7IcSt7bZ4aFdHS
M9ThdLrYj8TRR1U/TQ6ojoiOlvvX6m3dMUXf2r4sUOZUcV+HConjvUImfAV2l+za4yOxHIY2/9Ep
UiX2Fuyoqd7ccT0UxhJJ9enspv3W2RL/WS1EwslbPDSuW4Ro2HRZsaaYKJ1kINPDczrK2yax46n0
dElzrS+4BDZoVlVf5kHeolDEJCW31tvE5lVXItFdcfR2f3Dwn290ZdnpKSCyRZ00dl6n6+UAdpTL
HMOTdaYULul7NxEmfXInj3rS46zOxnQu4WY0U7gTDeHRn4PHKwZo/17UcNnGMnGA/I1oiHWVtBO+
RyZuvKP39+RmNZ5ZWBFqBzUaFttPZ8O0BylzC2Zl57ryOkWMCU/se+jBb0VgoJ0XDTBYRDvtcrnM
iv6mLX9AGgEtt0jcU7SKA9bETpItOkMoneSyYA+AIlYlV0216G2w9isyf6CFIBgWjk0KAcweZHAR
R0+PO0TOYyPq6YSXZYa1edW+pQfJxTzxUFiifq3Y6itzIvph998S4kTsGOHKKbxsKkUH07oyzhHh
+lI1ylaDrHScjqCmmnBFd2/NH2Q1/yVgnutGrOTckoDsOGKGHxWDKBJxiw2iHFuMJCm55jRc9bn2
P1JpuMMU5R5pDCldjjeG8ccIAYzhzhVBALroXeoew9T1KaXhPaoGNL/BvTuweYr4BiplPweSmRV3
F9HM242qHso6OUwgi/d9ZyNujOLOq9m1lT4nZagleysES6CkZpfE0a2Mg+uCGXFRjIGbVvFs/DTl
fQRwJG/bnXYYffcpGpoT9eDGOlCsMZvOv3BL2pKzIPfPLMckjsokCSb9MWV96BtVtoWok+VxcINh
TpexqRu3e4f3C/5yTxClHZJ9rcv8ThZ5oMgczRhvMwMq2buT4fM6Z9KJpWurHI3mZd60wPZjZjf9
fgfJdSSG1mgavCib3PwUGX5WZVWikKR8s+rn83d1jbGlRL4xzhovJu9JF/FLcc6TNaUt2q58tI2K
9WsfTv27QqEks6FKcM+MUBLmBuVoCsFwsIrNtWg9J/YjmqsT761mkDg6VFay+3ZvAeoDWV81XLf0
gPTV5ZWxrxe8gvLBSGai5CJA9bhg7XGucYyaUke8cDR/dnQf38jV1o9oiUeHgachel/abp/3g2bL
BScWrzeE9z3/YXudp5zTMDrirTv8nErpGcxhZ/n9hUqlkS94wZbCtKBzuURhdcc3McyAEFOCI15N
P4RfaYxtK7mM6nf3ILB4j4h+pTXsPRYOuWcKP3R3l1gi1JP5sqHvAYum64KciyHIkOxtYLtpIwOg
/iSqIaOrFVbnV1nK6lVgxTYDEfw5Vbk4IWFb5bsqGx638XSamQ0Ek7AbOdnNAmqEVSmxpZF+dWog
raNZi8bSQMrGDm+RCpCOUA6wpI/Bgzl1oj04G40HbRhT6YPndObWLjC1f2xtkv9qpxmuggpgIbJc
PTHrWxO4Dhnr2X81B6FHVmWPtGUnGnEpQANwF3Ftz4mOijjiYsBItOE7N1nTL0USm49jVhoQPx+t
IQaoiGmL7tz3Cb8hujsWkCGfYvEXn+lGQqjN5uS9Jw/uiQiLWPq2o72VjIeOxAH3jPMqoiHxUOVs
3RanVycopdhpDya8Kmz3OGnJnZjrSkfaiKHkQ+NpYpbqE+cRlc6AcaO95Iv7mWmC2FQBHEr23ixP
oWQ89ErUDchelUIbCyH5wV/Q+hEkXYyVka9HD5Qm8zchiUsmOvDY+ko0A9KxjHrg5u84m7kmu5e3
p6w4C+3VKfV2Sn3bRy33YBS0UW39VFVYwYu5woH3C31rpPmvHMogEmfyf8rcEAtBQNcO/ZApg2Mg
iFN1HPEwAapszO04R1zG1tuC116O7BFcSJ4ynwNtkDTCKarPU2FAljms+tNYz+faHalQSQf7bKz7
Sltv3Va7zXFK6OQpfz5HSDj6PwSL1uPS0Odwr2Qf6MrAwT7CGa1HcqX7/P05Njuvhc9ZG8rnAMDe
sXwuQNCAfcuqelTy/o+h1h+YHN3WLNqHh+aom2aS4njStNt4uuSJCPK5w+OIHqKqbXt7LWSpZMNM
TTYDdRbM7zVJo70753k4EtZyZsJ/Rb7IU4PfaLzZpfHqgtzln8IOy/pAsy1ujSAcuISoIu0DylEi
OLJlbi0HkxpsIsjjV5WlLFiUBWAMMKkAyVVQOomImXSlKx8pMZ5e7aN0PmWeORIi/f+5/Gy8kozp
UzBQ4cOlpjp5NCvjkZ67M2x83A1GneLtug+7RSy5khGH45qG3BC7PlU8kroyhNaX7ZIoSn4xjzYC
2XEDPmSvrTbQcuD4B9Rv/DUOQX+wNp2Emuqfu1nwqf/COft1m7FfPBTCM6IGgt6u/6c+7xEyC9Md
QTKYBjYyIzdlI5AaX1ProANpNC0nfyAaiXuzeZayyp7C1/2IGpfUrCOjASoyZ8XAnzXK1v180yu4
y7ajrhCrFW/IeoXN4DGgSQupBdDO7dxSl5+waxk+6C67dXk+xKqXIJLxWraqjGCuSCP3c7+86hD3
x8QrYEPMiOt0fcWJmJz7wwsW5g8O3OkA+QMFtYs/ltyKhvYAQObojH4+wDio8CguZhZB9uUwG7Vr
yyxRTURLrEXYeFR4d/WTp/bdANFJ5y3yu7/McAs3b88a3w1PXerv2buTzn0BkCVFfC4z8exh6Vae
iSA3z347i7pVXzKcVVUPc2FRBXEMGxqaJ86xoaO7iguAIbkWlf5DH+7Te8rxW3mlzn6R6FjGkus4
h6ur+G2Mex5FiBQ470+ZsJZPmtyt6GNDJNbytMxm4iVxNRxPBU2YlMC2uwGciG7NdVGjErKV9XX2
jmKJEYV6jCJwKUsmPWViVoOD532RvnBxor53uyE4OD4+Zi9zESgqr36FNHfKSlfte0Ai/heFfqLn
ZRE4enC36i857f1EP9kelL9WVo2KYdKdl5VNStH1J6958No8WDor1NrhL5FWbcFsq0vLEDT38qs+
u9m7iM0AkW9ONhxmDR9vUPML/P7mIFBUYdSLSGS2ojsoH6dMXoMEZE+FVR/Zpcm0qjUktUDyuZfJ
sM7C4Vs9ZZxmczq3XjUYGGSDirjjSBbK6hfeFxh+emXuCEsGV5Nv0pJy1Nb68x0bZqOP6qGLunIZ
0SpW7HbvTpf3t5+mFxmSxn1XvgOLaa0IUFPPumkDo+Ro5HK7M9zBrC44+LwurwMHWMujtpJpCEWj
Ubv4ADFESrre2McdOXFdlq9lh9onRu6ZUWKBHCdpRAd6XoP40unYMMHkrdwdzgrVuHv3A/eulP8k
jgbqaz4oTiqRVSm6eP7gSlRnXeLmWPCzltGsWJMQyVhRi6lkc16JF26N1nGWe4ml6zSlkSp3Z/TM
YBUQf2qRxwLjpH3mdpsrdnvWWvXvof0D41huO5x7PS30LvlvL76Wg4BPuVQ5KkJegwuHKXVNtc/l
dSIF32YeQAYmYsmHSiXwEh+yBB5r5srbTNNCRjNZnKTvopu354BphoLk1mARdRd/ZfnTzmBtXnOh
brexBKCCVgVwhA2E7/NhG9+sRaMFs41/kw3GLw2vG0BeM6vyhg2SkA7dLXJ14gTF0agSG/UaI3AF
jcyNA0ymqisvPKay0HFOoywMH19BIYseNNxwARYaqqsnAbmy0Fz7e8f9x/hZlumA0ZIcDg5vLVMh
tPr01pqAauKVVVkbHSeGPu75GKh+HWqPWDD3AoILhhtr0+E8/qsBe71ovXPapBHzvKu1Tpedwu3o
muUcjrTXTjlDnhNVcTtVkHKYkDl8nc7UtoKLBF3EI60lJ0GWbr4NkVb3VtBzdY7voMayJ9qDBISh
pyR4H0qq7cMtb4ySM1BDd82hAChoSrN45vnlRKgEurcPOwIa6/G+HL8xfqF2TkL8FGOsVXHQXvFu
EKpJY62txqZbyucBUEw/qYuDhfgyW3JZ6Yl8/jCLEEu0AjdpgZmVvX6WGPw18S3L+EbqIJfS25FH
lAmr5F3atUMgQ6xwU6SzCMz+uqs2mmmOmefv0Lkz6hPPsUKh++Jd8Cu1RbXv7TCK3fspBXJK3T4m
xQpyucUA524YCMzQVbg0OdPE1btxKl9uBDEeIKDsG5cOJQwREMTqnCLQI9kkO0MGNIQqNNmDRetw
NeHJ9OkuD5ateL1G/6ZY+ShyeCgegj2inr2QIQdv0VyyLLyA+wIgPV3ywvj3MOZd87Nh/KfdJ3dS
v2ooFA+jaCDJX1ugUBT29EkWSKoNBnae5edcAfyOqK0Ls+Kd0ca+a+TYS9ABMNuLjAPcez+NR9FT
RwAm14h1bfaf9UKqH8k2bz4wCmOkbyYTYIrkdUJmn/nSMSAh7ABPgQ2aAhqNrNMnG/cf2m7IkUw8
uVngjCXpCdnLrN4L/WTYOvwxZeGTY/5+hsTHsfLi8ZLfk0cIpqdSDwpmA63uFb6mj6hw4LNmnUtq
OO+a8VKFIc0DfWbu1cjcfo7lKbJOwiaXREzFogXPzOeld0QMLGzwn3e8PqF513fmdzPN2RCP/77l
7WgfRz9pQvSr0DnfpWCvF28pYCUgL3jaYe2vtVeUaQbOPMuZG+jFHt+NYjKlrNYEFw5B44ahz87c
5M5fQTuHKpCRjAUIpRPeSL3SQMrDq9a5MwQDedANiMbaGBe5B6cu8lX7otbDvWFaN1Ue+bVByey6
5FCqehz7NW8YeC1FO2f2ajXBvnRCjqqcSf12NFOD/ndogU6woGOshaXW+GYy1s9W/Dj8SGrKXkY1
T5we02MSXwFpFtF4EdWhMn9LDGpEgZH39evG/K0DULpiBbhUEdHwKAKOgMLrd/3WcLty5br3qPWv
OQ/8OULcVQy5WhCtvt4kN3llWT1SHG/6qYxTLhL19ny9kSGWHo3Z81+IZD+SDc3sQ4ozLkqfu2Mq
zRgRn6FGxqYMj9MNprjLERpeyUMRiNjFti9aV1cQnUSk078JUG1CmPvrh2pWuAgCekWRtCQI0lkZ
OGFlO1S2Pf1N5Wem46f9z8dNJ4kOn0UNngjLKBaQ14ImLgjfq6HClz1lhXRbs0oPmQsdFmnc/IE7
M86g7CrQK4g3P2g+/FZso/0kx7TpWV4A3M49cKGXBE/but7r9I6TSFpbLEU6qYciVLwZrJWZWS1Y
FXX9FuOyJsWGTeV9N/RrpncGgpEFN1kE1SkKyGZOHTgFFVyDOs5s/RInpc05zHFPaRGN1BucWGpN
4ASuzXGhes/2psfWoFZhg6KxfR75hpWMZzTc8vtDljhZWkFiBYF+j33Zn3tkpa6ZRhCIvQut+ARR
+ECfRRSnnrlLzYrTEr+Im57JspFazX5IJt7umDKcaqtGvshhGbpLCQLf3BqX380+luD6WqHnXT/j
tjILjGnWfz3DsNz1IT4ffarriD2oecas+1UgmmQMQxf2sX8DTHU83UqcvPsPYUxEJV1q3qG4jjKr
CDjdi/MkC3EgSs3QdqZ6wc497nzY6ReSXztfPUThG4/bK0nklXcV5j90nhmoXkO10kg8Chjx9BCL
f4QKK2zfoNO1y/ZdKasdfNHodxmCuT9mkteaeUd2UzsOnkHC3rz8L3t6706t/a3LTzDuitq6UKsY
9rNKwIU9jI/3Tc+YxbjvZudNWLLQn4ypfB7+WvH7SJLmINjnawH5aOtZGq7fweNaAFuE1+PSHRTN
V+MRchP69UrMDG8pQZVvXJD/VC+l81qmDvdIDd1GChWEqD0oUTC7NFamIxWV1QVPH02mGHI//v1o
Jzf+1EpOY5JaQ81veU0qvIGp+7ICaFBx7qqB2uCVyz/051TJFrpu9bHB/I7O90qwzK2DjymQtJH0
RrzQyjiaRzdlopBxQYVKwHobDioOP8/MT7fjgvXxAVaxR70RjwXtBkt6V/7H7/Bs1OT4f/DBVs7p
la/pCBV/yA8YSif8PEKPBYUqmMcIvdrici5aNeUfPHCB32sUp+lCpum9oOT4B56d8k+g8Ua4AhOD
a4RxBLYhgRo0zAMujRKjXNxOYd3Ds/C68ANH+UcblmScKA/Is71p+6d8VyusUwpQBoWM0yKuOkkt
wSlxwU8HcTuEg1qU7a9nRDy3kzzgzfoydzuSjEbP2vPD6qCbxdvhhGgW6EGCIMhHmlmekSU0DO1X
TgOzK4t+fkJetu0anhVLtaN55506YpporLqSf8Je/6tHiNndAtIgJGR16dTiQF9d7kLEpV+QAp6q
yKwE5FvsJkpOeZ7dtHUvC7Chl+JyMVk3+4/GviyilNMl73iDgs+Fg9rSe0DA1jFsGbfQAB1mQ1gb
y6qul/s7NPT5IDu311PU6ADg4S4PzUY3PsRdgOfDMCKyCrwF8mll8iU/rnzKivnCsgto87C7Ft9Z
zeLB6hW8TA0egmKFfN27c6lGtHSJq1gyEmO2S3btDRh8OksjoRtOeHQl3nJlxI1ltsiw0sPPMbZV
85YXWYEHTCepos3gFEnfRoKF/QIhVqrQPAsGYGw42meqbGrmpKJhHoqUkpWXY/rIpxO/WGiK9K1R
vGiL9bY01RTEVqx/oYdkZlUctL7cT10d+T0KgBTyxWcutFixSnG0/54azlWdMhMVOZ4fuZNXUIGq
TETmt3OBncQibCe/k51Y3+Ec88D0II0V9e+ouyI4JNb5c1oTxzW/e2nBYY1F3P+FUysKvHDCy3di
cQXsijDQxqJyLG3GJ/pw+X6P6i0jWZNs5GfmZYQyEGlCvGe8C09kbgY602rPW0EJzzx/vHorMoOm
Fq93y0KZ/jBC4jXDJ1NhpP/S6tgXW3MCWKLni2ZeaR42SU1NBtna77RFm4Zey+R34oRK3mgcYYes
Spg4U6JJdu8uliXy0FDk9Pd7VzVIF4heATaxWUvRExqB33pm5O6fZyTNBQ0hQJsdtRInFiUfxvKy
bfPZaZkWIUMZ1+Xyk3ciPOBW4Ha+pfIZ3vneoVZvoH/GIqKT7hXTCFk1sQQSrezs9z7Kc2xs+h9w
bgMiLyEMvxLPtHwxRmzsoaEz6hh0yAyGZ8hiiiM3kmF0Ph23LAN9uYiSOeyHkX+crrk4roVL3bk1
gp4hLDQRRnDOB75U6brU/Mb3sRmKRiJmUAdxQBavPdhlPkzbDiI+JXG3KzkQ79T9V1o1CRxJ4G3f
vzpMtP+GwMhak9KL5AkkuXI8ViNcvw9EIfLez4p9fJpMxsa3kZbrbwYU5/9kvPapWllWky8b25EC
r7zUHWSfiv6aJQuFBQmjSKsOj9JmA7KVKmiVPGjwyXLJr3w7Kb7JkiEUBY+ehCue3oULirz6Bn1C
2H+Bf8eiQUgEX8DMbkQRJ67qIZiAtwNjb+1oFTlQ1tZJuIDTwKWsdqStb0Srwiz/I3vjsKVpQKyt
FPeU3iePmDOMBFst8a1+utGPhQtjzs5r97bnq0+6pASqgZ4tC8XWxq5kEKKH7gmXWF09/al4yuz8
5AN+Qv7W7KSVstw47MkwTjispHkfyPQEb91RmnGnwhoEFB6ubOGVmiDRUxj9M38FlKzDf/L6s5tn
UT6uG52ZMXQFt3AunkchXWN6PdgpPkTfcyU0YkxwEKhG64BervqQr1D6rpyKzr01bYpuH3xd4sio
FdBzBE6o0zdqMWPDQG9CEpS9NuxiZcAcHDKD8G/JgE2OmPJfpVdubyZwsaUiay3hFEfnl29KtoVu
RMxR0wgOzsYH4pWJOZV5JC3xkyuml6YOnMaltezf3mdmlpUgjvBAqCbct5U6H6XOHFDD1bQipOmq
VXbKmdCuNiKx1Wo0zOGmf/sNvoktsKexeQ3KQjdGngrayC809CBZ0o/+PJRBlMBU8ASYeidjXMum
rtI8XxCqIURlIp1AIOj3G1iGsnySHOztOHBaiIFXIbdEu2tcqaNB1sUNGBFRXZRn2Ktyw12WpXoj
iuU2jL0eWmKClLUv2wApW9lvJS88Q00WR6ustu95sv7Hx8DBrABP+xR6cl2WzM44FHt6jL4ET62F
yt5gv+i+jgHEztytv/2yW17J4qtWddMvjEBaHW43nGbqu4o+9g2XTBUeHuobyXl6Te+r/uWNEvwQ
YE6z13Zi1jNH9BePs8WNBkDPu9qlXS6WYyr/yhp3XXd9VWcMIh3r2e3tr+uvYGeIQ+6OtOBjDs/Y
VTeqt9Qxd4GcWp3VfuvYzaslqTfDRyeAOFgq+AtOz14EZLj6T46iTZfDopQOp0SMc5szDfomZ/6q
HS9NFcfg18sd/ar/gSBCYRL9UYz+dhXG45CWnMk89YbEt6dNGlQ9FBqcQBaF5O6INkgi3lhwHKSS
lqaqm1RDzMLLZ3Qu0Sur1ZSHz+sSJW2ucV1vHJxbdkiPrDeirdF7J5IIflKakEpfdODnk5KM/Umb
S8p8i4+vYmmYMwBDYGM+1hLfC3cYVSVadHzNhr+Mc7wXhDyP5FPQO2F8Zv34/rc8bGt4mv/lXKmy
QgUrkUFKSUnwZxda2LuOUZnSJpVk33zqlRJzL3+BFfx60zpzsBMhFfKPY8WoeUvzjeVgIFVuZxqN
K9sK6ZB0nYK1vflZ+NCbmMUdeNsrd6MfuiytQ4tbPsw++s/ODPfTF1GIlbyR6FAr9XJbdaB6jado
KQUZn/OnRY9jJ414BqbV8JJPRe7GKh1AvQ6ksR7lQ4jR036b5zFKfArkrO2/+yEPpztYt0Yt5TE0
kkrYZwhZ9T7lNGCa1AJAJF+UYUndAX23XG4UXm7omhdSDnH0JhJeUbO4wlQC8vZmLYx+ps7aSe97
mRHis+ueZ8HgN5/S5Ov88H+xIaTschmk7bkv0oP+bWQAjTLblIxBsd+lqTqNo1dXrSTx1fWvhukr
SLn/ycFaBUUTz4ilRLIYiaee2GzstnbNccBlNj9pWW4DUFoezNFvMP9TXHJnT5Xf1ulp4kFuodwk
m0wF7IhyMU7ROYNfOKygJWABM2XotMdaY5zpbUqhtFqBxk9s874WThvtYJI4K2AMVx50mt1xAeB/
1WekH9nf9aECmM7oNP3pArwULZfh+xyOwzm7mqCN8Cgt87W45G9FMywjYxHpCoKB+7MBfbkgYdRX
QcSrI3klPZzxcANRCEOrMTQztHR9PAocr61TPlJMVqD296Rp7w3d0SKFqZWKSqSakvlWNcUhNVJA
sPJmHJkEKGFJRsYFN1Fkwi8hdZkRDNuD2KIavV8YIcE3PknoR3UQu93UaldqWiwD44DCb/KxaoWb
TBcHhYMRh4rb5Dwi7pWpQSKw7B03yx34K16X7dKxu5M3bp7PeXMUu96AXtk+XtslxzH49TY/n/tL
37GmksEaWBeNwg4MCi0KVejwapC1oeD7mW5UYzmh9cDCdYVE4aYrbR1b5GtCttxYEWw0+zJcpSEW
0w/mJGKDLHrXKu0VgpPPpw73OS7QIt52pMkFEVpa/ediKo06nU1ftwgc79+2HbPCIp51Ef0pYbjt
4Ntv51J7hhpNnATVHoCPvx72qeFqqzkdcxyV8YDAfjGSUNBkO0NuVtzhIGC1PxYlnQs9rsCYNquO
K8Au9etbUQMnxOAERKiCdTvN4c6suHA38Aq25IKnQveRslzgilIhmoqoI3jUjPJHvCpG3EA/KkB2
CFtohA4ReHYzECHr8PL4DT0WB3g/mClLGvvokes2PapvtDNdl+mO7VyrWWTF1awHlh5i0CfBQ2oV
ICjR0Yo9rX8LTbV70FPIV7FpQlhcON7GF3nIoK+/7JZ0/KzMBX8k9O0p8d5uZgWzEpUkgn1pRl6R
y5LwDkwQJJqZhntsooVe34hLodGQHYxZbNdf6kCZZGSwfv3AtlNWrlsSW1jEH0jHYc0LrV305vnw
XbTYb1N3JBft4w9nGSZhG8UIn6hOLYvLfJVQ7LfXEpq0szYshDmDx9woNqvsoIrV9PmGBZ83P//y
bvcmJ+fnpCWYoS+CWm0iyfREtPGaSTjVmsy4u0Jk6XrlQJflZCfeDfp2XxlAWvgCshu89RN/KSN1
uuFBpwoUq8TuLwF7UthztP1pCuu072n68nlk19RXo11V+afsftTDb0Ya/hsS/GKlm7wplJdZnzxn
fGW4cwA0xWi1tXgTQhiml2zQhutDtOwDSjRvgaliHwaXu87mnbjX7jgX2PA11Jv7QLBBC22ALcNa
O8/cfxH9nA0QPL6bh5o75frLpEy+besicSKz2OAG4OMEpm2zfFVZGt447DiFJZGs4O05DnpOqhz6
sukGEZ4BKaHKUOIVRsyKcUKhvb1lWh44rnPugbyJ3WG/yesM68he3xMuCv40HJeUWpCniCyxH9GM
GCIirqs+dKUT+i14uRe0v2WhECCEkcwgSgvd/Fc4YoVV69DddlsRgE6GmYtTdifeIzbSxi3N1cx5
pWMzK/HG/PFkjzP4b2h6izq2dC4frSxySbguMfRqN0ZvOJrJC5eVNu+XpE7RBwmPp0QDZ9RnGlMr
8LsGSNOVO8KT/0QULBhbqIcEov8W5c83c28d4CUDb7iLy1pCH9RTcbItTjIBLXv7uh+dUsUX5WgM
A1N/l9OVV4rEkBSFT/slnTn75lcmBn0GpQUvcCQlWL3R5sEKZ64QKv/YhO7McDVUh7LpuZ96BbEP
DO7roPRAyOxYRWGwj1BaNyOFdNZZwjdfUg1cWL6oDLwzPALSSvXrOIs2d6ssyE3BfVf7xpH0im7m
m3QHxnPkk/8jTF8XQPFHru56PatrRuR175E0nfIF1fYUS59gsW1rTlwWXOGl83b7f/h1BCxWcn+Q
WAV5clbu5iHEFtxq3YGjsU0FVhWmkW3TF1c357TkwO1nqhzlDDPJfF+93kTuirbtZmfuhUCU54uT
c3QbB2fQR5gXcrtU5puzNqx9XxYrhVJ56JTuV6MlvMR/TUTYFvOKFrQI6JUQZA2mtdNzPJCUtoig
ckviEl3Q7nyDXGcWbTpWpgz2H8tqeksWqupOpsvunVq5qziEdH3PS61FIw2JCb9k41oR5zFMcd46
NUAoSrAoSX8Y/yEJC2b1okqGvOlXgZEQ9yqDqPOpNgK6Gu4DdGX8b5HXWg6XtQg7E6aR8Ouk/fbV
RBtLD1uPPg7IU/dwI82wnIvuevpU2/KZGl0S2nsSb33fFuZZICPA1lvVsXldBc58D9GlCBdNshTw
wGAHsOqyPzUn1xOqyV8rVKcrR6GelFi2ToohE3Io1qX/V0rZq8kLwu51VaQmwkCMx539dT9fHjL3
IFk7SMXoTxtMMtt6etf4dKaPOvmNBmGo3ucVu5clE5DtJ4xMKoc7LEx2Ih0esZX53owKpw2qtq3A
uRDJd3WloQvXOwkHSLjL0mNMjX149woc8D20ufJW1aNhT2ZrmH+P4gQBfi9FEVGQJUX2M5MwNkLB
tljKt3XSBdrVrFRTvVR0RWpjzfbZ42UJZuRCgUeSZuEzUgnySJ3eB6Ejai6MoH3tGxuAoqKoImqN
qQc4eKy3EYPkxBrgZroBLMe+vMxXNRXbfGYucp86h7d3Sjvxpo4av6K8ZpUkJwmg4RHNfs9avK9G
h+oUpm0MYouuMHwvzouhPHdEiLiCiU3FUAWL4dYhE1CdBJNQowhTxQm9ADMQmBiWgnEqh+/Ln5jK
jNH0x3BEujyVoJ9hClLFwEdBIidZNR5X6a0czGcqE7zbgCbDLa9M990+jIycIV+qNfZqisrYfV84
M+RKU4f09iVckJEyNjgx4+EeQRG52zM0i3QRG13hDl0kfWAN2/gw4l8Oi3xkBRvLikQhNrqluVXW
ns5LyL2P1VMEeVH3b7/YkmnYnGIG0MUtRX1D5E03RkNUmGskEGSK4p9uylQ1ai88wFzPADsogbqg
VpBrd9N1t+Z7whZSj8jshx9S0e2dPpXujV/kxQzMge1oe7jPuEVZAFTrwoHBHH2XRHftkUl4pSWH
/YtEfkcswUIjmHHqA6wbpzBMhcZLygNiw0wzWO/luouI9xluT1ESJvpv1R7J4/OnWlLEQCXdoCqL
VzmXO8pwjkHqmdWtTotJo8k3G1L82R78MzOTTEstYVnHmF0kTUKF/ttypTypozdMmAhc7UneouEk
UX1BtFG5m3n1gcmT4dA5IEGjb9QINt2zoMuQ2QUEiUYK83Sgb9o4//aQ4rupzwt2fPA612i1H2tE
avjbPL08CfB/s3rKng4ox4MpJP8CuhxuRVNJHfvhjmubLjclll65u1dMiHAoHezCPScswTmZJmLX
2D74VQWTGgCEg5Ase2xLj4RHPI46hc2H+K1mvYXdN7Zjl/nyFSPp1+Swg29H+dzNVTsO9nPSnlck
EHBg4QoTvmDmfr2zliGYDTzutDsPuqZGfEXlVl1wUtxdPNuiDUDr7lGtpdyHcWht7+AJgkyA65R0
9wjSH+uoxGOxasQiuW3ATgtR4Gs89jCvBPfZyOdAbgQRJjVo1PtYXEuwx3TnuHM0oW5gLk77b0J3
GmC95M/ArwZ0xw+s7pUtndYmPlc4MoPBpOfTBMY62ZcRiesrSdWFFl44J0TfKAodhONn1s9cXp7A
6ZpPLCT0fGnfN1vOf2zEBExcpq+2trLatWwbdJ2GyV7RB/EXghYQfOO1VIyrio7d/m1Qs8qMB4uP
7QuRcg5KhnQ6K/3znzrWDm/86HYHHr5fuzdtZSPaHaBFmBHVaWjreXFSAHVx+YNXwaqIU1hd05Ax
nCJsUpAI8c+gVj/1Z6386ctutnmWk0OFveXMzfMmniz7JOXXT78/gSi752gcM20UQxgfbCAmKIBy
lYL/SCHXivngi8+ef4xfhPLP17bHGzVZXKrwqzJ7anCg9vTUpdyhEJUczKDIXxpMk5gbDh/7vx1n
Czmm8G5HY/xQbDlj3orwWqvX/T2qCg+F90GzGeQBIuzzStR7pxQONQ8q4WlBQnsdJ0LeUcLUmkFF
8UsjqMfV0veZqtjFPiefGISc8QoNT4jvwRnubO9XihWJyCLANikRwnd/93Op6V50SMFupRLXIZA4
U5pDfeQ6jsATz1zpwpxcYD1ki1YSTZI9tIUaZuwFvU34BseZbOhiyx1lWjBr/CPFgzq2s44XrcrT
1XiZDwkUy3cClpSrhjkCXy0QoFAshwB2855dW6SWGPHWpuVta8nPgr9qjSk+w6E8qjdIpIqIioWH
kGOrssX2LE/f2y0/oypT4txVBlglMkVeBHs6GY602fUh62uxnF2aR5on3BNhYzviuS/ypw5mvkcN
wtv2nU2duF3lYPV6idrAxY3cz7O+NX3oBphZ//qypMyM461NFcPz4WqvY1tSMUqsjGyf2U3f4i8x
VvQKUZMIv+xuug3YzdloTkhYgdyvqYekr7tN4hu6ZM91Fwvj9cnrkwipv+5lGEasysWLLbmao9SZ
zYFxvg6rRtub/Rdok8oZ4wuZ1mO7gmQhlVRKOPp6Ck5tcaWPYpceuBxorOPVkUo1oZmW9gRML5XF
s1qUDZN07cW60wOYXi/vVZSRKd+3F01s0LcCoKKuK2mRESm/uGKpfV9lOrn4c/v1MgeoQe3D7EcW
NOsHNynXvwPGtDgvuFDzsMzaZYQxu/PDoHR6CJbla9CekqWEUiaFGGWktFxVVBFPAnGjUyvYAFMv
qhmLFL/r/lUl2IP1xu0IzLbCMQVIvOIvXMDhglI1OaGoUgGCWVwy/u1oSRNLV0n2K3WQSwpovx2u
TqXBI5kn+9Bot0kDjQYWU9gFBqzonldzIqGkyGTQYUd2Y0tC6yKBOixHALgqKw13B7cjW12sEt0L
RQB2FIFC1G2NzSNc2VxXRzX4sZHO5Rx4/gKrggKtkvLI3QKopCh5YFV26HeM90QvmHSf6tIXzI5T
Druda0WhdiEzqXIwNJdVJ9A3sQC04p2SJcoNMnyY3xH9cTo6JSxVgRt/RSzYnnThk2xwN3aq1MDN
pieaPQiuUlUTiVftorWyTKl5VNPi9JU4SDTaAqZsV/qLwU0x4ycHokIiKJN9lcApsQdePL87krZe
DCqz75ODoExJ1NO32katuaXodgyyf/mG/Q5ew4MsnSYuqUYKzu7GTZNQVa0N+2f/CQHC8kQsOPyD
cZdTiNgeahUbkeg8vhbKfL2XF8yvJKforKXQP8g2/UqvrdfuM6LxbcdfF2ZuChhrnXRr0jgWnpj6
M67JDT1VQ2gy4tad+L0Q6q6IVtUa67plig0sWnM8JsJypChyiHI941GKpJ+CdDH2hhQ5XGNb0niq
4SiOffFsUX6m8tj+SRSKHPVHQImJzbFawbeuhrZyhleI94CGQO7tBFqYhRmz4YIYwdZB4qWfdWNU
cfYAwdDWinlxM8HNsC6EJTl18ip95sybRP5eCxurX9iQwRqXpoQPOBUASGR9j/iRmNkOluwDPBUZ
EdmF2v/HGnRhKE8zIJIdE8CHxL0juAY8wYgkm7Bs9bU8/Dzc+c1BhGZzIYpUQBNDy9PHLIjgME7E
J8AHR+BK+M4VaaPvMmYNYFOEjujruZw+WC0b4r6DugCkdRxwoMOGwrTq2WYBHtzzin+bKDc/dXhc
N1EHphmgrdJthTQYoWxZ1G4Pn9ar3+r3z9ElM1hUAMI5STU30oQbvgRM/jyDxNS/XwrWVbU127Qy
QKKj75I3lAZdeXDpV9X1pvGEzv24l8txxWysvCZZDBLEJJZgHrGBrwce1D7Vv4z+qqHx83Yp/R9I
TrIMwS0mC0QdH5risaIvIbIjkhDJYmb1jKqZG7VAN9hsWArWgP8PP26/+Fur0VtPGTgBy+kkYc6S
dQv+Qkj5aRgT8HSlUP9RUOiYE1z6jVTw4OPArCL+046qt97mT0eYHy/Sw/w8Jf6huwhigZhAoI4T
cv+G8Wo1346SAU1m11zaRszjFZlg6xOWEcvOo4PFN1pDzZgLFEoGdmONB4Zw5PS4a3tUDNgbSKEK
qAz9jf0d0e/ldJUDveP1iVUM9f+wwb18VTb8EcYv2bsdrvl0ww51dUyn94x3/g/9vW1HI9ZafsW+
mWMebNbWyfT0UTwzLSJuJjVMgt8I0ThtZmXUKwVZPuBn7ot3ZGWz84Wttl3kagQLLG8qezXCcAVb
pBjk1dXbZvnVWmIUOKzCTBD2LwyxJeO3dcv3b77gs7tH/AUimsFxZ48zNT9pAdCyo8wTj+idL0Rz
X7n+FMTvcl6mVax0nOnnk2Rek6kem/v1d1RIN2/zHmj2btl15QthTXBRPO2jlfvQpFrBb1pMWyMj
005nGI8XZn/+tP06tdEGmAbIGwfXMY43Zw6ZazS2/0tX/WicVQpmV7iFzjk/s7Epj5TO9Bvw7O12
nEPxA90RKugPUf/ezu3zkr/ZoszHFSckxJPfXx1x/vjxNW1GsDTm+vjoDj8GLX43xP5UHnKgbReJ
EWhc1xYYyHsvDSiOg6y6MXMkbDX77uA5IAPq/vLzxM7v2dz9/+ymuDgtp7eu2Sjivy33mwjDcXZ4
DA6dp90j4jKLVzAochi6WIDMeM2uQLC1EXv7jd6MSZ5yvX870+ey8O+rSKx/gDOErsD0F4c6RkNa
XZbRqgMY9QY6vOW3Zs/vkbTTkBpyIqnSYQ0o66v45PLF+bBWLWo2iN6PZXlhQ22eCHdUY8pGAs+S
kch18YWvkDnq/dnFw1ClFk/EIxMlJUa7UFcQZhsQ25cvIHc0tA3o2CALAZD3spvwVgEdl8y7++8I
kFDZwb21fCcqIEg3Suqm7SKZ5otystQENcxusdpCv2IFTWs5CDh5MI4J1VyibDDxnCbho9f+Dhy9
D1WoB5uYTCDNs8KvHibplmXLpS+1kmWY7NP19BV9yyekwQp/XpRUGbnI0UEkk2Ryrgb/psxztjRA
62NkXhtiSofgA8FEubE4UlVJPfUZYUls/R8E4S4yTyiq085aLfaGiypt12cQ9+5IkbtArYyzvCWr
djEhq7PKyy7yNjgcRdrXuiy4Yh1UsygqXSiZV7kG9Y4LBBZxads8lK3nV+b6CFIjpUvkJcja8b8u
dWM5fQyynAkCP3tMyZcvJtJ6DHsOoZMALMWQ8TWmIbQpT/gT46CT5kThDDSUNW/1In0S6QhkqDKv
xMLYKK6g/hkgnmrLjHjkLqkqGcYet4ejTTB1ku5yzVETZc7fYJmZO+ICu6YlEzlO4sfsQ+1CI4Uf
39brwDcFYrSc1tUoHsD9AgKZF52AwkwlHtMdP5sRGSF8gCc1pO4LDIVRRmTlD7Y9ydmbGpqdaMRh
fA1talGGK+AhH49Reb2BklJnm1MfHIMBUrKw6z07KnreeTTSnzUEJpucwYTjjr1QhmOiuU8LPOoi
pznqf3ZGrnyS9ue70sCAjEOYjyVwi2wmA82wb1aqNMnMGY3ludDntvBW48S4RM5etC3gsF70kAvo
NYoJ+6WWRKocuyXRlN181NzpvLJqnhX8hRTM8uJft5Tv0OeHE2xW6LTilP8XXFnScb0dHjaOO8hg
lu/RyVETnRHjXn1uygl2F/5Klyx65+EDfeM2nV4xQs58bpQzYf/bqatSSqofi1qhPVJ5RSo9FMDZ
X+wu6Vm3ke7wR7SArSocyTj46w/VmfkndegncpAZ74YMqIQw+XVkmi4yd+3xn9EOEt/fbTkb7lHq
c/kpxQTzoy5Pb5EJrK8k0bZ9xC5vMAdZ9VpnLNzu61YT/qE0EoZnQts1eJ374SQBowJPUyURLAB9
KqS6NsZAGhthAPs3fQzfcuMcYESqF4Tq7t40oJtJSdrvV2Rd9T/7x6bOjm6Ts00mFn67S1jfDLyM
PCyiKnDvxNfjtRlWhfbRv65D581XT0irFreIjdys6gbmWEjJoBgv/QEuyP/e44us0CqJcBRjzHhA
aouoNhzAu9QIra1tfCF0sr/KWEEv8n7KL9g2RWY/aQ1n6GSH3ITqcePvTW5s6yr6x0zVfyvS4qWy
InR7n/ruhtPNxVlbOti6b3Om8o0/7TMNDItfBDO6szOjGUaMOavk5IwEceAuyZNPKJm3YgOcv8H6
hNU8uEdY86jtTDYBTKAQX5KJAM4Jf43o/IR8JOUXhqnxcClMhdkTRX86ZLYeVRiGePkPJQb234Qx
1xXAT16NPokb0pB6F4yUjgYx0MMZVwxohxASScGeYdr2CcAXDjeIOM5Kg5iEPXEKR8t8JYyeXgIi
83wNOmb/Ss+J8j1vyEknHSi3rZkZf8s+d9OX9qjt/iSDxs2fi+18Zpja14fB1W83w/F9tFasRDnY
6GINTNY3GnEcw1StjeVb2+HOlulIjFVRGa6ibByYJb8MzTR+bsN+XDFg8uNNBYmbGRu0CKeLBwSK
rbcXzwdjz7wZbAFQNQWnQxpoQk5qO8Cq6XLb1Vk60LyPcp3ANRq948Z2Ce0fllw+VxVgc2hffwVm
OUE9cXl5RZvEzvmRGnAUzJWWLuZXWV7WtJyD5i6dkNLxlhLQgBACdrwffQVgD7GuDULFVvDnBXF2
wi6HY2c1S4mfbdE6fytO+8QKkad7p2RBVz/i1R/gg+YsOsKNR2fWCWxGxxNadYjsOuxAHwgUlrlA
OZ9XH+96lZeHZT7h+s1Q0gf3sO0iMYARfzr2AvMUUy/G1ujXyVRXp+qc58ED6duvaIepYqtFgfSP
nTF9ua4PvFPsnyd91o6k2JDgdMp/aw31Q+b9XuYMlZmYttpW7WbCEUgfJLt4TAKQCtmAm/FtGpED
ZrzO75j/dBMoYMJif9SdybseiIhHHQsQs+tQrt3gP4GTxgDFoCOhLvfrW/vEbZ3ZFCUIX7MjdLuZ
snCyWbOA/mVhavDAH7mUaaU2BcRji2TuzHazfjma99uEm3NuvWy/eAHHPet3b/BYgnV90e42E5Xi
0Teyt2hgdCUgAAtKnpNdVYaViFGVjqAiB2JfpEflstkhnMLHxVcBFe9HQgpfufrxzc0cLjBnZaUN
BPBcbzYe0hRq7NdTbOhMjoQ7kAPH4wxLtzVuhj/bYYTg4s0/mQb3NvAXnT0zLkqPTIygi56xCGNj
zwvyA50+RRgPRdb8q15OqvvmLD+dbBZpjlGiS08BeFbWxqMW8MpdeNlVq8+FFh1br6HLvVrUbmCS
U8iH0v+BO9HbW7wvZhsdXdUR8Qlla4NPhEdcNm4xOXFVoYZsP6eNPC3ST2BYVn2STyDLZYRnM5gM
RW4p3CA0M55/IS+8xgLvo+76/ktQc128/oCCStOGeEq/tdD/9J+F8cHVmaa68iWsS6fTKfFlSzV0
ptonCuK5EdtcxsBLEoF+Uc4Txu7WJMUevcI/SIHA+z/nb2XUTRKkgaCsA6JEUNdazg4UkxAavgib
Dp3OpQhDyDTOi3jkGWtUYlLb8eix7ULQRVdfAL3uYIftRczvQq/xQ8godUhZGJl/jvpLH9PYRNsD
15LcuUg9Zr+5YvO/+q+PfJpKiduHVgFnQsLUu0ZxessCVZ6ky8i4Iq7HtG6LC7as+rJYbcBR8nWz
UNvkpWyug0Eg+8dc0jJc51jojH85iubETQyOQDoeA7ZoYTIV49vBPCOU4mUEpvHs4j91WpTXiIh4
FVtsLaOgqIYp7ti2jPudh5yUJjNl/LUmLZBEccaMVUptHxTK44e7GpaiqU7huio4qbJJNaLH6tGA
Yttj0b3App/cIvQ5XmDyW2T1P/x6ZZI3empi6mwqUwidKnysksGb8VIw96f5i92B9ptiIJ4Kj843
qUBqQNXFe0hoCl8/WdhA7/UZ2tM1El1wWbrevHIj9+5rwqTWdllouIrUj0exlC/ewMgHzGxuGYFE
oN+U4rgbForpqfpyZGtKxPV456wqG3fgKyp9nuTKgSqWeoT80zKDOayzZ8cdkXOf9iszZOzBBioj
USdUxYzEnXhlIjJtJMTKdXvsZKg6l/w0C4ryt6Ze0G1XDpQSxm6wbPHGxD7mUK0P+4akPJeHEr5U
y/3avMRHRPtNsMdAUiCF8f3hQbTlUykHNdxRMZBfNRNEU3+ozYi7rF8MKOas7kwFtePsymAdcryE
j4joGpZvc1GJ+TRLV7ZBG4W0A8I1fRUa0RHIAf9/mawzOd7K7yHoGFRXRCN3AXjqGIlH3VPulR9L
BjYRgZHuzJRZ8dWl6424KSP1Zg6eS20u9SAQIA8qtkYKdkaq9j37eiYYai13HcSwASL+AmBcnLWI
n1CYoILNksjBMvGbc6s32KQ1Jz9YlbKFOBoS3sEkf3b2c2QayRU0p6cxyF14QM4jIr10z2wwZ3To
wIqCRvzqQOjD38fcutRLMH1R3lA5PudEINI3g9rZDGWYWKNdldyQDK6sWa/TxjaFUTJTgxB8PHiO
5rfiMyUlOrWcrJUp1PIeE4E2ODFK0SXNsD4gt8IA2T527IG/4Nki688i3IgQpCEOTF0FhtWJTaG5
5QY7qiCoNt47Q9qyIW4yhLoBhPDzDYWblGyxJVjiy4MSdEZ0qkI5OvCe792JqL292BzUZKviD75A
qzEZJ3UXBejJN+RvyC/pXWyDjP4lGDzQJweRRRyixNUmVQTk4pv/CFYt+QTlFF3vLHL1dSPrIX9O
n8/qpGz5HleIjT4XmBHIBQcvfuTpzvJ2FDTk5ZrN3zBRK0by3BTfTaxkbTkEDJJyMgECwpLqXOvD
dyvzuZo6rwreWU7yKemaJ3tCYaWEq14No1VHvK0itrJ1Wo51SuXZQJ+nu/uWbhyCOTqOzp4jZKsU
cIAF33OBJiEhXUm8gsmmU6+Gt6O8meNFTLP0zMC4pkdMLrkaJhgpacTOK2YlrbeU9zspQuhDC2XG
6JXJaE7T6vPgiIipvrX/Xqiip4WLtKVBrJdp/LlINIpa2NTOztzyjhhtgXuuMML/UJrJMXG+xlBP
q6Thocq5V0u/kO1pWulkI50xbFgW9JfB4KoAwkmW+Qtt8T3+/4NE81lWrkeqtrBIuE6LjhJdp9wA
7bms49kYHfAPX6+JciD1vy0yqctMsWlzVwy/lCtGrMysNPRRmOvHxuLHHqaqGvkOW/qpfXdYyf2N
D89FVvrNkVtdHave/Bdp/8Bpa9E/jRHJcEOZbIhjlIV2DfdulG5bDrofWe3ec6VlCmSJYeGU+izp
ge+wAIAzioIoiH9LWEisiJrg/3EvrpZ4s8vtNJ4vJuTgFXPj3yznrDQ0VdbjQkrznYyELJUoSf7f
Uc9vVHpScv9vKSfCrE1shUZFT4yHbDLLf7Z0c+o+VryAVw1C5CKQDo+x7u903EbvIhQiQya0yM58
xQ/AEdvOJMLmdGEHjb7d+bAqdOCnCCYG/hqR9Bvm1VzcVEMiZGo0J1+beJyKYDWpl78VznT9JVX1
BxeuVZc+nEt8hvbHPilX5RBfT0Gg6VrUHaKTZ826tt44DbUHoKRnMUu2xKaWz4wI6VHB3449xtyD
WyFDbrtTTYOlPkjptU5qI32mRLJHDZcGBQVxmRcmtiO8rtavT3Zm6M8uYNfozRBNmu7oiy8SeeDR
058tUc8yX1ucMF1xxB4FvmZlRDbqodZmaUbfZeEmDoVeaVvuxXyYCmMOsp5h9dCRMTGgZnqR8UpE
4tVaCtPTkQuKfAqd1uUqtBCZ4mJwPXivVlIs8ZS/fT2ZlxBJLdn25PEcjML5GKx8pfFVEWQ53bwz
5B6JfNTinQd0NWDrquen0+uI1HF1OZGg9WflWduCEElY27zkzpJ/zYHzVO5eYTXEUseoXNzRe5+1
c7zZ8dVVYMkSizqD1ItoyQ7Zhw/sPWK9mhXwvcOhxWG1/0gYrq6yBrc6C8wQvxruonaUenSYfhyV
xqOGSL5Cb1ICFRQAyNxrC5GVRiV7dE4Gg4W+/yuZ1W3RCuDbRpOtilIZvGergg+AAf/A5QrqvnXx
3DFpsZuWLzG1IUkqzkLibQ2Hz976XmTVn/FraXNLfI4UCiswFQzO/RbzrTw2ntvitg3IWlCcu3ml
9pzlij8JaktSxrEeeqqs+HtYg0qZrDBzxI5A2HNTFwpPmkG5DSd/GNzL7Elu3RkeiiOttA86l1dJ
OlGXlD+qLGvI7YQywDTMCjpRpBUx8hGMVnMKWm5YV1PTEcXJxR0J/xPbUD9OJ1U6ceBgKKcVoBDM
4JGCTJkqmsEGRGNCb+vqGyHjZ7v/rVF44CPIynRGuRrQZe7XBILpPFKpIiWnK95DNL5hpqWiunCe
JypCQBBUOL3uBQ114Wuj3Y/Thb0MY3lbM7eKASQr+lH/2fXtLrhurMd9I3TkkesJTJpBAld9hXg6
nG64Ct5b3cXU35SBchQfUw+csys5Vg5hsuvmJKOzkWGIae8nwmrO5lLrxyUaxxcGyH877WJ8lbNI
fI75uqcpH5HWfKWpSkcx5dW2k1IdME3tSMfqbvhMLDIF2ZcX7rK9xNE1rjR1XRMRXfQaGkm3jkQR
PuKoDtGkbReAMPcpvEXy8UyIdK4dFmdFIvsWsxu4U4f2CObY5OfMRH2+ffGo8TKw7aq8xFyzljRf
Zu+epmJRQuIgwtsAh/u+Yo1hk13EobwaLrg6Kso8t9rMV4HHaPQT2i1UH71Q6UzhYny+lxh8P/w6
tVKMhaIjVge9ciNTtBgif65kEqN+VoNFcqEN10jrYp9lxtjWsjuBPjzwU7DnQ5xmpnjSPJkDM6t3
wLgupS4rhmulfcZ80KEuomtuDnWOc/x7CNdl+18HUVz77zrrCOSwgq+4CDUnnt5X0R+xaAOJKfKS
iA8kUEZAmIcdTMlidlBUFQx2cBxbElRUbPLb2lG1l7EV7iGDpx8CrDdAB4HEeBS2xcgp0d94cbgx
dJQjebl8OLezop0gzoquWv9KeFLWKRWSXj44XzFAuIU/zfvD0oRP+/78vxhA5LLziNquejlFGUlD
fWvf+j6Lp7b60q29cXiBncnOC534U88s7rlDL+blZ620uQM6vOs0qyZdaK0CZ/u9KpzQZCf0m8ky
iG55qk0HmfY+NtlCwk9qcMhD9gtYFP7FW1+AMfHYxyaIpqwqd1W1uP1W3xVZTBbwtbatuNPAlJzB
37VfL9tw7dwA4evgeRBj9W2HSIQN0C1JXsh8Fjbd/4LljyWGc6XxfMdZj6JD7N5xDDyoLqgXvSCr
cABxWouEEtbP3JUlblDS3BdaLcfEYoho4z5VHiJUqge8pGrbOaSWW7C/f5vMt9IGhKaRdraUkQX1
472T9geTdKTrSHGtxJjfLSb5yHSLKpIahtianQieDwvhdS3vdq6M1leKykS7F+fbD2qvgoWQ9jGR
5ZN5TW2UKi/6/9vdzgzAgFrDEPy7db54+KsC73DbU6+uLL9t5b9l52FtsOPhW1ujWHy4p/wiGcDm
5OitN8KmJTI2TzQY++O2UnA0Pg6wEg1bnT9ANDImB8s4yTtUZ6P1Nwj+KtHD7SPdI3Zb3YH1VxhW
tOZ7aqcHrhG4VOopAT95cYwL8ajX0Apf6fvjiHLUu/rbUTlFpNYIbJ5BTpKKyLvjkQ9rxK+KO+aq
ygoA6mX9XRNAKuytDRZhAjQ8Lu/MOVxUzsH1tmmGpV0k6RDmkDPQiwe78JD6sbFyu4H/fvaqsdoi
O02RgntBZ7w5gqBuiq8faQc2OCjSsKesbe88QJ8jmgH70iCyprLOzg4zFsKZxy9OP7xn21z0Jsdr
uG77jsn6iFRmiDnvnvo3oW3mEAPM5dRt+DLsj3VTKE4uCkKXQ9LWhZeFBbxXAShsXXLYf8q6+AyJ
DBfYgMnI9ubYI+CyrKFjvslznbBOeNKP1j5Y/xOXBL62+nzhskUAmtROCU0UOR2AmJ55PR9GUgeV
XPLegVz/qFw0XgmmV+zD5UT1l24H7kNdICJ0d3/BwqJBE0d61r3m58aAHi6JDWQBrFdkha5HTzpR
JOlD8rqM2W/v7dLUb8vt40BMXcsiDKGrcVt7bkC4SvgzHz1NMxhQc0a2u8EN0K87tSXAwOTXahHh
LzWui1y2LnxpSmRUH10sLiwYgaSweshnfZu11YJch/biw4eDpnhj/UMWs1Pl+6qqMwgyQAuLEY57
3YReTFy2ZgDz8z6foG11Hs8aHjJUEBWQzkxMx/KToV9aWCywK2JuagEwTOktyGX+YvQX1Po7bybd
2rVYIgnVd/HsFFTJ++5CrFyw7L28hXJ/FltbqMUslOcEFXM29/hWq5AhDa0ekCc/yD+/Z0H5fKg4
nWpMRwAyNEK7L0Xow0VOTixqxBhf5LLEu+Mimp8WrDxHuBkeMgtYHFuve8Ryv5hkw64454kESEe7
3bEs7oITktc1Us/64mK2KzjodsHHu0cKC13zuVS4J78TTVLQIZ6zkBfh2fk0GZJ23Hl2daYKtXAP
RgQu17dNUqTo30VQNkpOAouSdTMxDjLkVAPEFIOcLhOgajZy++rMGV+GxaOtOjaAhgLpRdtTnPvR
m0i4HY2v+WtA/WWRfvJBsQIWiyo5I1C91mBZyx9LiRaEg9L6YHmfKIR3j0d6aXlaIb3zVReYspZI
3wgbRyJiVRME6CqBNZCArj4iuI7crM1mzkOn/sCP5Rie0KS4BIHTA/kuPZR9TzjQvxxM2ffrV90+
TkWSmzloWNRUIvT+pmSky3C/z1YQ7B3VE06kq/v930uDTWn4+hS4OwJFT8rVlnXP2DFbKTdtA1bQ
MghQ+CZjparrry6gzwJJRJAi6HNmTlBx1ly0PgJkQZQhaMdTSbTVLu5XTctAlggwgvN0PKaT+2CY
dgHVZ0qKqENbtAbX+aG3IhCc8BuaMuFDCyJ7v0nhtO3cCPJDj1Yvvf+MlpWjERXGHFLN2472fRIU
8dJiTxOhJlF4RUDDFy61unSA5IPTajB9i5pXe/l7nPDc++5W8xNUMW7yOyEdMdXrHQ4c9aR1sk/3
k91PUCY49fz1GWYy3EL6/7WGwg7fm66eh/Q7Qa67L/gAv6k8AHShYdb/t1bYRjdfxW4eES1b0nIl
fkVF5tN5C5Ol5nfdtRd6BaFK5WbNOSoAh13xragmww5wcF/ut+NIKa7GipJIeUVe8I71Hv+8kaEN
XRzsI1QewsUnS9DT/GKvM+Bh/88awm2IMqBxcnqWvHvc6HTlyn9yecUZY41MKX9VSLeaMYAzRdHD
lvdFcJ3qVz4keQrb4i8/tbQb9mi2xz1kIDLIHxl3CmSx9SnuRqT2bWQBTWgN0tQZX6KBDmBJ1mJu
dUOg+LPOyKmudfQfxS2wIQL14KhWkZBGX5HqO3/HPfDSodoFW2EXKW3IIaQ3J4ic1tnl1XVGSAxf
EbpMsUTMhLvpmi10xMq18xvAScybVNbyioAcZMiKmiCUCBT3eSNVnH0PzKGBqKsMrQWTA6npdKFs
RSYUa6fic1Tz/11DxPOKfO0oloCaAbxS2kpMAW9TS84kuJ9+oPkgefcEwTPKqLqcRFH7fIMLbMCL
d6cy8hfd1vxCFLhfBT9b+DCqPE0vW2YUIjcBGLrAOHleon/A0l3iDeXA5fAReRuLjjjNuu6c2De1
d55KvlCHtEwnzQUn5uzH8LGtBAgyxd1vkUQl9lKF8yawqQAfxUdDKuv/0n6QARP2kG99va32euME
rekdShcug2Q4dWWXnYxkcwsdzUrGXNxM2gfC3XNLxmS8OuFrgjR0pMqBCjNDI+Et7ZwR9/aq2O2V
XVXbRNQv1NPwitHArQ/ilFP2+1OopBSRUJk2F+pMNRXfeGO3t9NL/cTzI8HthQwk/+OaxY568add
AB08Jiy4/k9IDdpZU8LYDg2+dCNCyYvJgKw6XSAjN33HFSl0wOkOi0RS+d36f2VyZfwjbpzheGkN
k0ndu0zk7qarTzWAoSND3n3RtSaCGx5HDYrx0jLPRgWhgUvd21TFS6Ndauc86Ve9bv0Lo0573OWc
4EaGtpnRjgXF1QjuWgf8rmc4tdpW7bq3jeZ/AC5ficWTelAHDYKXn2IUtR/ttmtQ4YQUUu5rIUr6
NoAQvdKAn51v2nIi3jyL7ryRlCvU9FcWHJnGLtVhjOxaFgrFvr26K+FfMRQWTdUflNegT/VgKzmc
Qf65Q+Fm5jCAZK66NnPSE3VQ+0iITl/edd84HNjBYHByRIBWczRIX9Bi5KEjgKRbDOlpe6Pal05t
jKjfUvp7pDjeuCwoV2p+dLXuq6Fm7iFNBGLYQL1onPOo6oYW7fwTYe8A7mpapkrO1sGe2GV4Zpim
OFnGX/kbHw0/HBVbvVK7Ze6qORGO82VIbFMKxM/9FloSyn087vr+4neFHwvbjyQaqEK5bTHmjeiX
WkhY9nx1rcYvhW1QMjRlihVKQuswCRU9SGfNku7CTgy0pl/9Ml7GL/BDR+59XCM/LSLSn3jvpr/X
qa1cVVviqjStWecj/ifKu7mGqDLN8/22lkK6RW/98yO/XkmlkxnqRbLW5pOoD2jhCskuveL0FWXY
hZyQ27QlhZy6wtbPBuuF+1JUNN/r2+mTGKlPYYiYS5xYofCVU8N8J0UtusLVtff1AvIXE9xJMEen
W+N4zlkaP1T8BxQ3hCp+uRUtBaN+WsM5EwSA3sSR9UYC3PjTuieKA/S13cj/OANn3bzJ7U6wnfkS
jdjmad1I+FNq40Rnr/wIvApntTXoyADr2z8k404J1UlaFAZmb9EQ48NfYE4FrWu44RGDQPB9z1+N
90/sAAhChahG+oC8fvKuw5rh6rLF6eqYq9EIshqNeIyawTFWWDvQVdX1FiAfxWxuBrd0uZXVJa8f
o78JvLfXw3o+PNMExnI+OaNncsyftK926aQQY7WNybk6GdPj8B1fLWCcUOc4daoa8hWYKNhsn3WB
UcOJ2c1otuXmqQFv6vEkQ7Sbrc7Ly0/r4CGg7pj2xAvaPJL4AuoWiKh+e/5Tx0ZrKmSLeAYGyiwt
07dFsmM5jHq2JGrN/I4dtueaPQF/5JwG90HeUiuPBiubllkM6KkCrtIRoDOKodbVHQ0iDRKeBkeF
tZvUmh+cGcuJCLjx3Agkl+Rj7phHJltfzDsXTTw8znQi+3ShPNpVrVhBMT/AF1kgSyK3iskYEmYM
S2Q5MDLmC1JYSvViwQXZK5oh+gxTMk/qLQlSfvuCwhp2lIHUL1G3j6QWoX497W8CpHUU7c60PSg4
rdGL5E1RuPlAEfawTFrLYhH0uHzai/1pnXH5T6nrME9ufDB/4mfli8qpsCi+aZYIMNLo3Ta2VHxJ
tikYbU0xg7slBMhBSekuDjur9jCN7wr0UoIhz7oskswkP0uT9WiQoiHaB7RQgkb/4gYQgHA+LmD8
zSkIZVvzwRwIM/LwssXf6pLdThf7XG7aBC9IXQDL8rcJHb9mE4t2tHQ0BgKmYhInezkK6qWnNZx+
H+jnTljhN2DF4hMb/aN4tcZP0fVYLnYdlu+C5h2M6K5lyVI7U76H1C/1QQEhPANEiXCo9vPl+t+H
CHPAYMj8hXVjIJN94O+jVWw+kvG3wzzJBtnLLj8Ld/4wyWMPHOvBP9rMcgBRxWCcZwJtvD46lnVi
tEgKuh3phMSDpuhKhW9FLrrPZaRgCrZKcTxD8pe6HOsAvAeq/6ZdEqIW8nHVHMaKAETC/h36ya4j
DPRC1VRksSGDMKF6x729rmWBTVghUfq3WeF5dEwTrGvtRHnIQlQzI0Gb3ts5mdr0ce1S+WYtpxZ7
GpWGUY8NIOwcKVkeZEQJL43cQSA/KMKDLajSo0BdatF+StnOpVtDMAse74BoBy04RCNU1tOjjGg5
QF2XIcm50mlXfr3SKKDkAozgM6IVE6wJsBBzNkrTRhuD00ie0MZjH7xxPPRbmuYUtrquD2y6i6OP
pZ5V8nSxiEPK2oMXvfblxJVET3r5eX+KQ7Tjk37gctFYeHc/5xBNPyPS2ujU0806PE8vXBOIX3w3
+/PhQPsoaCgp9SmHt28DkfYC8mzfsdHlB8ywIde8sZljohgRrarbHN0VyAOYCqq1jDrk6/Kw8eRd
hWk7gPOocAdPHhpbJgzC7bgGxO62w+/biCnCmkcoDNO7//t8AQlUQQEUg/HtPryw5F+ulkJ/xRiF
KoE/YJ3oQ2jvaCq0c0BnsPH1Khfdywf+nKsf6RK2BVwVK31U7ytnIrgBEAJ2ygaQVp4Ey4/lFpBs
auOeYz2leWoppRU/XULSoTr/DubpyFkl3DG7gKUQwJYysOMXsni8K8Opy/ZbMd5Pvlx4A086eMnE
aUpdFEIjZUr1U3XgmTbGKBtmvvJsgokAWCnG1XsHpw2H4ptjmvpgk+uaeHNZucpK7DUYNhggq15g
GbY7UheH+2d6f+LWVWOy1nZTBNIzhB53Q0tZUSYy2MFPj/12sCUP3dBgDt3PfpJhAU8eHumuO3Rj
mRrWvrmfgqGgumBsYjfYab+6biWFlPu8+lTSXMKyAn0jyTGxcZX6GAMm2y5uNELNUHXvarCgWMDb
nzCKGKXYVpzRlNPP5WT/lwOG7Y5t99EuIZAEIp7HF5Ng4pLAHuYgvxK0A6XSggIRqiGHJum6k1NO
ILVi7d7aW7iA/cgMuvE+Eh1ce2YRTpz/seH6YINU/5PH63WwsWgltJu8xLx8zX35dx36SageEhVB
9M5PECQpcbUdvTzSd1f1yXZP/Y7AIPkUu1Z13xxAOTtuEVxM4CY6813JMwioNKGNtDsXhhablTnO
ngIxn6hM7pZXL+UbceJF/9EpT2i8c86hx6PVEeApMCtityoW94MRAZlF6eNx8SsgrGgfxowS4iah
SWyJRvyKRVOwwhZV4oZCZD+cEzQDtBIS8La+xnwhexewZZFpmV96Z0W+CM5qYsJL07pML3jAYOfU
dUoIK/d+Zy3bQ6BP+fZ4s7jp7TkGBRkMUoRaCaK7Sf2szKQD4Wm+1sJPrGzoMUwwwhTDL5t6rId+
+5mKcr/piYlUw8KmpICGJkV5WfvSMr/nZFByXuAmCnGsI3gM99A/jUp6UZJnVP4RhuNry5tYp4iE
ShKSzXDe7INaGgfbmRzzfG9DQoXj00merz+i0i6WVX12TTzuGVzeyT/qnMgBvTGpRkLDIoe/pYt0
hB3V/ZAvBbJgCylYzw3uvobfMydXGxF95AYR3dSWawxAo3uVrfcn4QL3Vn37pRIAlD/K7Z0SWlbd
tccgGQssMn3kOmr2qWMZgPRM2goSFjDzKuvhUbl1/sVqj6KVBL6BJR0RByFMWeZtPVUVyCbLOr/n
Mc+ZlhoSUJQz5ZiGNJEeGavZLFtYT8XQRpSNGa2ZhReDxaEbHEMYJzka3j3VOpwXpQ9wxl43twpL
FTT8hre78aEtVvS8JEsduKR28gHlvOV8TTSxTPT1kKpTMuTJcI9BuSgsczs3hicXtGvwBKgIsnCd
tcK4tj8o0GdBlMj4Du+wksWzXM036X4ZegF5k1JKIACEy36kMDkDQzfYx1TB41Xhf3TjLIGpcUEm
XgZmiRIdf0uabFH+eVFzkjs5A3ogSDvzQJLiWXmiHYbj3Ezl6vlSiSGTQnRopOgNkEhJCdie9GG5
60rNpfWn02FLiaLxLYocj+NgYXG11ME4RY8AeeG/r2lE/h2/RaCCbQbtu3Jvirawao5WyBh/EwWy
MbibykiOPPna5gqUKv4fXZN4q8/PuNf6djAzfNGiv/Sd380wUu19tAzEI+ek8xMA2buw26Mdjgnb
GdyRePBDdlv0Q+kah47H08X1ZvHWtb9EtyqcuZeQJKdlzytbOchO6bb49aOeHT10aYhyD71K4M0C
eltAR/qUrsDrAPuFb9E1+rA44ruO9gRasAwywxo6DGbXQeoda91FbFtMoSNdxu0tCaYf5D8hk6CK
cC/NfMJKPLgBKJFbZyGLyRv+uUz1wbNXixqvMBym6cV+6j6K0tGNaJ0t/xuhl0oRM/Kbsc4m0rd/
Gci4/K0pEc3O/tDHSvpvSqHxRAVKtBC4cmo96j7ZR4UgkeskFTCSmX4mkCjl2Mi7IQPWBGw9O00i
CTdJLjdKDhKvaUeeygtjs+Fba8+VKTtQRW+FcJ2omLFSnv5HtfyczijBRGKqdz/xQPLS+laLmTJB
CBjUGe0IvZ58fmVpHzEckk4uYcoqXJYl+dsXdadILl7QwzttphYpph0+Nrkbffv0q9zDBpo3TIS8
ohB5hFD6ECgUHpHMpT7lFCWGpaKxU55AlZ8UYeug4kvgkzIhdH5dGDJpDvPw5TFEssZBbBxxF+th
WIHMwmPWdkw8SMUMqugzxoXsEvhgEvxanbVd+9LVu3atSWaA7ZGfGPRNGJiOZlChDWvWCBPmfYk5
H5DteK6OFOefYQ1IXOWG8YQtCtXJSalU9Z5gMfs0rwulr8Nq+jCRHhFNK2JO9lUpJzwqAv/Wh9ZV
apNcfxp/Txff4c9iglW8BM2hCW1Dgw74Xmutp2NNCkZaduYqO4oOtG95SK/s5vqOFkoQCfsz8qP+
xVdomhYmhW6z4laWaH6xI27axUcI9TOH564X9PSr8BEjIOm2ygFlXmAYE9e4X2b0RkhBfYSt2XqT
MVg6ENJZAo+FAJFyoOhJAdebdlUpQFLQN4ZFlt8YPNmTHy8ljldt2GxD7xuyOSnS40f0hj4ZbKKh
0FJU7I72iS4KiBfI7byzAHFoWm9fVFOWMn/UgTcVO4NnVtl0y0iH5DDSzJHSrIR21pi6NUaaq0sj
7YbAVeysgJND22XT3/Cp+9PYQt+I/ebcwOFr4T2r9enIht+u6fzPGEiRKGINJ2h1q+f9DpqTmpZA
wKM+7EfMm39uiIkEForuCgrVJKLQkcTnI+hG1CMMyS13fq3pqVVqNNZaP/uXrh2v04PibRub1aN3
LUGsN6C0GlF9hElR5M7PJarhCb8A/7OinUsl8Ak3aYbSVLMDaLmpj3tiUDN2R2cge9zR0/36GTLj
yFXn9Ow63AQZK+VpkLysYQqqhKt3ycSUh9HXCBFEEqf7oIkg/wOxDHufjN78EfiLNuskGvfiVpjW
uf5om4beo2f9WZ8aqNM20kYPH4CLqIYmmEdTZz6rlU5SQVZQEvqRpDHUgjf8PE+2HFKOZ4XB0dot
GiiKJo+NEzHBx71IUp9NXmQij2m1Ao7YXY78C8z61+bkI1Zpw4d2D1I8/wJCFp7e6pAvBns+6gDL
Si78HyuWXbO8NV9PnlcZQjejSadDVfzZPs1StT1JCVtu2aviPoEKhSJDHPV47M43lmEY7mfbVYIb
OtCdJhbGw6ZmFmi1Iu6v3f35qQ1xIWyDeHvvgRyQXOSBFIZoS46Vpfl6wbRpQd2bs8Kl4roeoKxq
obX0vdPqdBcJEitl07K+4ib5x0vSy0PctbsrDzitThVE7oChmSXUH4TCCgAFW6yT1aPvhBAgu/HK
NyppbLMybFkxAInLWHrBrumU7M7cIgT0oxhUzxUG2Iru8xtt6dbtqAx4j90iVgXaG01wktmMZBG6
WDiromQzYdE/NQ6qlmSu7Rs8Txp91old7Yob/j5uKWUadI3UWHbxo8AfKYNo20efj/81z3ZLdlFa
KnN97WYBiFBSS8vsNsP53QUbGpn0028hv7R3/VGMzb0JhyLAzy1/Rw5l0NURyKmcQSUxvb7Ry8Gb
UqyONovrLUadS5lmTnMeMWKDV2Yltf6FxCuh9Ob8SZh8LfMs/YdHKIwKGLOJprYctyktxY3NK45c
ToBOSU+7fje46LutehtDlPeA/oOeNzcdvqFuSlhN0ssCcZTDreaYihISgaJ8uBoukSj4jywoiIbI
gQrEqWGilonlVPZ/3iylWoZkbDJ8aXTGmx4CpzDBZp9UHcSzy4UbME6OJ2On0zfQc1fq9+5Jffcm
YOFc5Cc0dk0tMTczrLp7bklQHC09L1rQ/zo3vLTjwplhzk8cSPyougOVNB0qBU+C3By2fxrWpcQP
PbgDDYEBir/aTSkypAwg66UT5cxj49ApNz0Bdciqf9mZSldlSYll7cNR2XMBzJyAIzElavKfZfsh
BfVxPPm/9+ZUVFXLoXxfT9lkxii1rIXM9g8jmWnOoM8nOVL6oFQlwliQK++JpJRYm55fEAfYVF5j
Eb+T1+Rf6AaKIQJ3Jq2lT6mjkYAEyo873+e3CPIzfKqmlzTjyx1woe2JRGdp02KEynCvd0WhaIpI
3XXXnFhtvBLArX2KQT3C8U+rBiPkhus1nqumhA6LixH7Ht/sNXQLrrpsiC+COct6hOUaEZtiLnW4
Lm7R7qzqR/P/S15JVE16zgi8uKTnyYHTgW9Ialp6wYbPHrOpI3SgO7sRYqIAA+XWbtACnjleP1fs
v6GZoHZOPHXeeM6vi/au3ebNmccBa4D45piQJRh11tSMPiU7RYvVwYKU+b26coB3vGLVRQV0O/IQ
0untgTcO79GC6WbKU5hsxhnRPq0ovquZOenx2f3zzGRECfCe31uD6bi6ua1maMznE6jAlBmfv+cF
ASxPWHQZ1aTB9bVx1NjC5ux7ePMPS3OfKBqRTLPlGDkPVPFI3X3wunobQ3T/phSR2YRXMmyobJ4c
ZajuTTcphfb4Bfj23THa+2hYmrZZbOviSNRdXPpPoWUoHrhM+oDDnX7czOudQpLKjv4knPpEpN1J
3rSOfXDDaBrWbSR6l3AOQvUQ+clHJMi8gc+sszWdykFqsckfMAnlmZ4i2VI+NO6HaBouwlHwsEI/
5P8bCKJkudzTSw9KXyrHkmtYEjYsLyQzLyUWC5X/cwngBSZ9hWS/O2kqLA8U2OSHjb5UAK7LDygx
YQTcwXqyLRVrUkNTpsrS6iQSas5t5QK4cXFuekNaT3/uJ2xtq3llT2ftgYbeT/LlcaSHc4/LAtPc
fKqgAh3ArjnvAxD30zfvn8tDZXXRDGKiaFVhuUTlPd8RjNh36Q+jC7IXpjd+Ls2ULlvCicvdZJr2
p2B+j3B26iLGz8QlLvhtMRBCeb498HaLUr2kayvQoL2nRCa/ARvliP5jgQnMLntUFdmq7OS48O5J
FEXMJCPIWVDMnz/CWg4nLqm319GMBex8vXp5Mxz5jUFSPnSrUHNWtnkfCuiuLNnsF6s8/9rW2R6k
+4hVCwB2ibg8f6LCkcU/bCuR/duSDcd2dsRCNgOpFgS1vMt/owabe5hPz1ruhoOL2yPxqB6RvzPL
1y86dpthDy/hRNBR0s5Ok0NWdNxO3guWGKloz7/g0+E/1ujN4tNaqVz4DZJc4Yn+oAZKrY59q+Rf
MkvXo5ICrjwslEt73c3Pk8KniaYyQi+hIk98VHwipLiZZTwd4ORTVO6NP3puJFFYYZXtQYbe9pT5
UgitftqH9beNxpfrP0E/nGvAEF4BAlngnw2yY1pjil0y2NKH5gsCXskNYnGuk4SwaRnLyDPdVceH
hBbK3NczskZrt30AWHLeBe3TJnuhOyjadvuO2XOxsBkmKjUTLxVOXe67ko3XMIFXlSGcvlAsVhRH
VroZVFZ4Z+Ei9wYNutAslPvDp6jOL5MLUqpLHSf9477jjIT4Qvh6o5phg+G79riW5gcn0Gp9rUGq
NHPoKol9el5gXgQ8h+vC93rVpEuJZoO2bFB0WnbFWVHkCGhFG094r4CwaFppDaLq+/XOqMnFJwwj
VNEAgl2J6gtP6CFFeK0UAYMV5dt7riwCqGzmGtAt8qbF+AGdG1lBJwUmFlorbEwzm9kr7aM/3Tow
OYuIcTnZXgqM/ZGylcYNzIEqdABpouvh4Gq/jlEgR1iTHfFuUTMBO2KiM/5bYspAfY28808RfHT7
lIg83cZHzfd8FfnIMOHS1Pu6Vru178CmiY8psd5VfMkKHFZGmErQIo2aZGEuwWdDwu3nBVGWpm/H
pnQqvsxAYLpqs9sL55quQTzdYbIFOxpO8/2aNilG+RPQEFcuuRfDWIrPTgikkNgpgaO895HGwRpB
/R4FklauHZ+0KlikvxG24s+W99oU4jWC+MP2Mnh9CuC+DM95Sj/Nw5cquPv+S9lJQyceCUQkpgfl
X7EFb3NzZlOmauTvVkwvO2CM7DAntThB9oR0HUniVe5fUBtmVsQE5wg9rMALpgyKkViq8O+4djoP
+VRQpNASujUDCmStADspH3RKlSj9ciyIxJILGiVzFSWRJMCsLsZxysFLN+gEHf/Py9h3AHTHoZ8o
Dm1F/hYnvZaSWiIFFRHwmKXyU0kwLi+MY93pKYcIzVWk9JW9hLOMxOfyGEoMdtQF+3jP4uRS5nd4
GET9VaD0HZ3PeRbwHgl2lR8uHVRbcMa16xsq3hhNN8W1LRVon04pCX7lsxCJ1cug6Um/4mugda4E
IgYrMbz0V5z+mgSY2itNmchsOAfCVExcrasHPERXqqeoHDWI/fueVww4arJTc5OAu1zgbsetOys0
kzJLR5Znz4QP5kxPR3k0zYOl2GS7i6qejrXjoRl9I+SawZr1caVQL5tO7nFmcBf4s+5GzerYSzTg
cqgvgQCT8D51naQOzVwaY6fCYHsiMpkEcZbJHJCf0tf5F0Jxtb+JUsU+isdkXLyKo8KrcPmYSrxM
oCIiqh9vLdDTq/GsA/0wPh0WiRk4TjHR7QPKDb0jt4fKeaAZXZ83R7frQkVhYTUYO/Yhgk+FDBBy
VAdVS2BZemk0BQbZjY0C4bSErRB7CdSsWujJXZgVy/Bp6IJUdZDaiC/JbLOmTfl7Ze7nwcIgw6it
qU9Fcwn1dAlw9PDpAExjnX7zJxJk04V6lUggldQ1mNn/E7gt2KAcH+dtYwLUALNtG7nSSugX81UQ
JDtwIXiZLixG25IqE69gE+D0lREfllHEGrRFu4tCOEdFVsugO3wZUJIWQJXrdWuqM+g0U/OboCAo
8zNjW1ub5FLEGXCgT/QEI16+/TsGF5KRt2xC/Duub8Ch65O5gsfOY3zOBRx1pdaA5PwQzDAtlhae
sLBOnfA9iPTG8fZcUz/nq9UgF6haN4CUXwB299SkKr+HVqVmVfM32iTbKrimtHy5oXDkmjGOLRgH
Zm5cQc8903n8xZ5w/ZAe2JAyA8ckYqoBlCub3X7tFX9VNedcl/WKOjdeSXFXkAEGlBFwYV9wRVx6
x0zrKMaN+vuJI5k2beR0JVurubLakL3sOIJJshglX3GgRuGrcyhd306dLz23SYRkwJ4ctNoACP1q
HA3JTLqLK+yZtp1ezaoQKGUqAf+I0JPrFcg9HVbl5/yfw5nPOV1Ix833O9cqXnRZAz31bnRmQ398
EtirPyhiCfaih5wXFUKoiGUDLSxF8bL8ZJVQMfICQhC/SSda4HBf8iKKUlyuWD2pNekwee2NsUXC
P5wtJmMCR+2QujPEgrAYamySC9p2VzknZ9hFMJasR61bTv/TZq+quU1p07+yG8Euloy3m+hDpbSB
C8vgWoQOTQewjHW5Seo2GXa4AxUVC6MVoN0DUl1KQ/tF+Y61lfuAF1KTshZg9TDy1iDgWJDYA1zP
nFPgijNgqyPmTjxwS5WYKFzFfp4TJkuXA8JS027p/UqfBIDhtgGB5W1QxERs1+KLSIiu2w16EdeY
JujpoIOYC76M5cC5GYrrwa5z5gSvar94/lVw8oZfD8cN+hJ+RhF+oDHOm1gJ/jekYy8pHv6E41Rw
wwPX1D2VFyB3sNS+ZiBFg6IV5eRLkhctQYSxY5NmAHSPHoCWJxhCY3ooBhwMFsL70/pxTCE2IxlG
ZKjC2LWAWjioaiB+aDJIaqBD0rgCQOlaKLbYozY1FJKZFPOYtACmln2F1bXLuuT6hZdKLbJ1IiYZ
jEYfY3r5o1N5RfM4vzyxuwfgM8fcImf/GdwA17GJWZkxiWta4M7RFIVBMbBzi0vrJ7NYw7GZ72/R
ObBc3aSPdL+6E2TSuNW06zY3qhwPI+UbW5VKUW+x8FleXP8bPoaCUKjm4hlPcnjPugCHV8csnXRk
W1/43otAt3q2ouBt1PeIMbm8wwkKj6DiXQzS5lIuKeLUqVE+PYV8Q/bxZfggvCtOX9cMUifUnZOj
dZo3Bchv7x5NUUys70CP0aFMgpxkmeoGNnu0UmtBSz0Ht4NYmw5I8wX9xaGT7eGL6I39ho7o3fbe
b3z3MCBnpn4U267GxLixcsstSnFfExfh83lScJZ6K23kdCMNVmQ2VJH1fDFXfohIzCMibkNw9/XU
r2vbWBP9x42hm5RP6xDby42SQVL7mxuVELxcvs09Hz4EV3hiAvTQPMyLudnfvIpc2fiAQnWGS4wQ
eH2z59S7odFefel95/ElmCv9kSYxvUs4JOA+C4RY4NEyYYFbXfo9pg1fdQq2HlvWm90YSCCMIv8P
tJy9LQGoSSQsOCebSXMUgTgMdQlCZXcP8SKW0zTbQ0NtMTvhLu0Nvs4q7eYSQD1200AnpLzYM//0
a73D2LMOTOfLS63UuljVjk4KgGTudgNACUh5fuO0rDi7oM+kixB8QRRSc7YeaeO1FzKItAWJdJ7O
1pKNPS2mTW2Puwf+6h+LPFpJx6ln6fNDGR0y8v5teivtQZb5TlMouFJGzX5JVyXOYORUdSKZhbhb
0LMNbDQL35O3mL3WS93zyqTxpW9XTYy3bo6pj0L7S1daQ2QnGOZ4w6deJyHk32AMGFhoimChW/2t
Zu3eAViWdNAdZ9Rp6y6RaqlnFsbKiczgc7NFLC9PDgovGh7yLnd9Rw6AuQXdIwlAVJs8sD7JA+lS
BaQtqT+oVdcPDdWp1bTkav+zof1jqCK4+fEvn6i61UQR/icZ6UtxvYJ3nWlrZvx7t4tCS8X7Uteo
H8u+MSnnmFK3Mq6kAdOzs/83it3hpMHcMGGypHXINQvqRJ979fqb+euQHXTRSjt2/ouUUEm8BEdA
4bIPh2Z5MhuiyVHxBm7wMVP5YT4f/4OauNQHuOpLHBXGLPRYwdxLSpaE/sGHhPCi4A4ao5ZTlXMZ
tr6aUu3JuBHETuZrpcrSDinLB/o1JounTN/niOM7dQqKcoTmWGH168ec8T8AIihxtATQ/iD+F4jr
yCRtnE4ysfj4j6Mz88+82Q4TK3u7/2QhsEn5sYYUg7fhKIldiyp5p/YhFDLJv26CWBcfUnUPs7/R
ijGqOG9GT/BOFi/iG8FmhiSNPlOYY04Qa1HODS3hc61Pq5LVqmN+dsd3ov/lUBaC4wgNFSK2G/jx
ibaqzeLcyc6HmVTOzEU6pR+X5/A7H79crK0PgWWWKMqN3o71GFt24T3HMNxZp8JF5p85KWPbipD0
E7ZPucV+JKqD+FhIum6RDpYZwCpxHsUiEKQa+eFcPVXotpmtLIsRMb3qHU9UcMTnmnECH9X3XFBF
McOwXF7MKioITJ9lhm3YSlXV/pQp0HCPcUH8RMhOMew9vskcI6AKb/mfCiXmTHrSo4jY2cId+TvB
3ugz1FF47VVdGWipAV/Sh08AsY9mI1EY5jRlFz/CztY0Cy3cjnmHPG3uYYn4+Ky+aaFSPN/ZUIP8
nQPz+Dl6Uixyrd8eo0M8pwQKsleJqBM4pqtotUPTDabaHoRUhqvHiFdqr82b7Ta/I7QWycW3L59c
+fhIUvlbP+S8JKJmJtC5EuhtMWemtZVFBiJdsjVkqHGzWq6Ok+VyZVRkIDzISWS3yvp0DC5eRhjC
iyEZHYsbK5hfPLBK4xw0LoOwzts07qE6u9zklt+atnr8UhOHyiPuLiWSg4CY5McNmqMcLOdjGNVy
DK6LIy2+EJQtyb2qdPbAhrPrVEDRi6mZYXaIGtwdKztC/nDLXRUSdGVO+gI/jDXAxyVMJlj/CEo/
hpDRFM9JYzU/C7gQSPR35Em82EFG3wtonqTguAIIF20/HGpImTIDdzyxR8hW4cKQ8ZQJ8qeWLecw
kl1iMT6WoyS/jnBOBeECKufnl4NVAnzFVEBZsSDw1/D8RLdwPrAFo+fakStaHk4hGve8soW8b3tL
zZRjyMJj/4TO6hs8JGYGdWvghZcfNPXWwCHAsUMNs8Re6iz7C1964njA2U1glYJrDJtpkGfzLDJD
D2wY9af0TUvy7xYVUtxjTkoI/v7vpG4E3i2K/uENEUuIYQQ4qnyBgTQq6lOSJCgXuPsk8KRQWqrU
aV557iDQO/ytBWJ+uL7WKHVTwXDaZ8ZiSavuGD+7DweKeg1/59zayxSmtz+pAxfawUMbWsxzqBH6
HRVOJ5Nsr793fp4Jqe54e8I+Cien4NAbOK3JSaNnM0vFGdeuhmy2u1G+XGk8Sf/H3oyevLLJiLp1
WLpsAYHikVjJXH/qzHIvd76+ke1pfAvOnasAqvuPuD8MovBWc9v4+eVJF2gCfrWz4n/n7e6cxSRQ
cMXUQ3b13PLoxMhm3KYpCcf5tZNUQDHYBgQIvjUMyIjPE1fOyQabhJBmagX9itQCeGrhnmrXrlww
HuqNBS2tzHOQB/HRUJvpyKZQah0cJF/S0v0HXpmvnUGejEjzEspY/GV+vEphTmAZvN0KIgI+M+2H
wOpFxszZ0iSmVzdyoyQ1K9mfaDTkKk3ZjwvpK3srTd9zhnafBycQ6HjgzB1/ZbGkHmGIKGzbMoEZ
OxBFLYnj5kByxUW/mf2Gw8MHUEHDAt+z29FvCObDxSaSuxrJ8DhNa9AvlErvrbSclhpuigKXGYJ1
8t/QJ/df5DrBUecpA6s2ioUoRZW4rhbl1TAbZ7dxI7RkpEsWAwrqdD7Svxzezdiaw+1MsXd7PPp/
4GuqDF+EzmKS/rsx00hBEwQ8LdPlUbl/XwJmeYcJFSkeUncYASQz2kmBBcO3/4FmfcMzYKHVcW9M
zmqSP9vJyFIYWWAx521iUwhNf7l749v2p+A7S+PQ/uA3ZFuxqkg6yNZX5pGU/G9hyLPjEQq7Pu5d
Ys4hwjEs+Guiagph/fEcpKhVrRqIMQfPtXzirRtcVj+jb+gGa5KKM14QKHxbkvT/iL2kVP3l7Fm0
YSJ6LkdvBxxuEhA0HbgokZEJJbpeGwEJYd++XuM/diq4UwmV164xLPu4axg94lRfYMrMGWkbW5te
AfY80+2YpNBVdNFm01eL+vow0A8H/naSN2rS7ehzY6yoghJ05Pc9uklAprrSWVrqx0g/FQ5Pl6B5
pQSbbH8lITdCmvhi5b9Tii+BsHb42w3wYB2gztbPEPSrgxfH9KwYaR4qbF/efbAnOHPI9jWt8W+R
QkmUF685CaA3s/HOe+PhOIXYLMSBuvT2oWmb6xHz0yPf1wHwktn9K6nVKmh5OXd8Kyz5Y54uWndh
g8HvTIGki62ewceqYtXR6Pg88FPjL8Bm181LyU83ZUeGGdVoA0nSQs28ow742JzOhMmqFBNK7FTb
pC5LifEahHKGPAZoUcPjZW0SjDGn+NqwhDdtOrdKKbUgELw9UseS6Mk2EUv0UQnvWADv7q0BviYg
l3C9Vgx2o2Foo6tBpkzCcPrM1CVqSOlqtfUEwNqGJH1DEbaj8h6IsYxsmwL2j7DfRgRcAS+6EXt1
oaLVCEnA9wt8AU/KFjjaoBnFhE4n8OeQjrglYL+tvCZLrJa8wOonPwzLtykWFT9vWRZI9Plx/VMb
hw+H2eU41WVpn03RyAeO7d232zcw+TpNZajNm8yMRf7M0D4rDDgQse95G3NTaVQ0DICVyRmfKPlm
do+ITVpbWFvjvmJzASqQ4Op8KLNFYt13PtEaJ76ZC9qKLIMn3ZWuN+t/nLvjOLFQmswmYh7iALZJ
ZAEx+dgdc6FdLfd8vrfuE33g5qWIgeAsfasglWMwTT2kH2qWLl0Sx9Ysxl7u4+mljxK46mQh2BxP
RRujttO6PRDsRcGg7pHnCNe3rEkU9gjPPWh2QIswLRJ46K4wECbpg9431kUWP2phBVu1HOY2mNQC
rfjpfBk2YJoxFyrl2W96pTURIQ6h2SWVcGdLZA1YJ3ynJPKbLCoBHLOvwcgpT5ad9GqtWfCs+gxJ
KOXXYX+Rvw9nBnV9E+GVC6dqwgiMQSDAtZTGSx5JjYL7cxlekjNgH1YQ1x2tHq2gbsEhXspqL/cb
lfVr+46BGCgJOPsvqH/WxpCrauVnw3Q9HposIjRuQ6CLJpojjiuNhvbAhDaEygCu8zP9QPClBsZD
jxZE6Wmp7uXORFmO/dGm8naTeAGWwZsszm3TjjXL8nsg8v1616nNDHd9oG5v/0QiKOl1Slc0JD/8
wTq+5Ic6YnsS12TXAj328SlE6Cy/VuLHiuHgF+QmMbxfV5N21zr6TkAfjbcp0a4iz7tWUs93OqBJ
sTW9nPINDcq+qg1GjAA0Q3Rl71bzXWh0Ion5n3OcukhNeu1LSUBHicMF9+Y037bZT/UTUAWfxXAx
WUCcOstcopldX8RB3cua7nG3+G8FtDEjZRQMX1fMKAeRqwNuntInim/PD4He4U4A4MvbUCU8vqHe
K46fJMM9LoHgCWdkws8m/eqSXgClxuhT0qsgvvZ/LsSgbCYIoVsopAUUaWjiMTuz6MJ2hA4eTS0C
UzTmA8/TlFUDkCJjO86lCyZf+xi+acNbuHD+3BGCdKPg/7J5ldjr54Q5v7HsHK1HE0koh89ylbcC
H1FbR8LQ0EbBCL3KI0wR3dS5XXeNMihynPQfWba+Ke9eBvUy+kI1abf1W871n2irxXmV1mnrdB7+
/WkO6I5WDGmfBxH/CVPSLdBGUMos19eiMITp4eRRTqaZ/y6g857ig6qg0/D/LcTjuBvejv7fA036
6gk/RvE2wS4HC6elyvpljaWrrfAW6xHY++R6E9+iyIrrGPfkBilSA3EadpwA1ToM3MVrObaz+1az
PNtJwzIdzSKyZw0EnlmZ/+YAx8afGAZGWuMaoKUvOQCCSvfT7eW2eUDzGfCrxv02feIE0zPZCnTS
JjaOy3y7pV3z/9fIqRFc5jZdNBXNdYyrSuUvfpZql92yDQHlJXu3Pm+VQ3nTSWlGcBy8Y2B3XRl5
+re/adLd4KJJV7RRQRocwwJ5vGQlLRhvdli3vss0ijiH/d2AIcEYdtq/mW0/qUoF6D8u6INdptfQ
LTiLJH15UUTok2OwTR9qM3DNSCphHY8QzOpDeV7tcMEUnNhu18RPT1P4ebIdMnQ5D5rKscjY79q3
b00kKCr5nJE83Z2gFOvGCeQ4CBLXIqaUsOY4SLsm9fmkOg+cjyeshhy2+icxeeJgp/Fb3U+ZV6wf
LDwdtBJOoEh6Ghi6OOEj03KgNNiv7jOJmTquwnyka0XZkrFwLbdAK9wSDu5Z+RTLxL3bWu3h3Tqc
POsDGzRoUVqxB/VyNDOPdBhZp76ZkfYFEWWXZSdQExPtbx2GTKUCo2sh4/KdCyoHw/vAfKQ1tXfx
kcG1yPUAXNxJPTAJxZ7JtsOKsHPekfSKS4hp8LpTW/c2KiAPkzHDYy5ZZdJuEli3sOtN2kwdZX5u
HJ0F89n+OvV347I65UMsurI0cC1XH92mhYxFlluYcZRLM0D9b939ib4Toh2e/5dXi/141XwLoVOL
/kGU6nduXV9ei9jistyCwF3wVugJPqzEImdsOPD1bMVymb6o3sN1IT+mR9dtrLvN+Sty61zRW9xD
PWtGK67Hes+ip7KMchipEoY5teYi+MT5bd+QsT0KwnoxAL9BJZ01tQhLgqryaVk5BjdNY3jncR2G
2CVAI6WhzdQxHC5Ka3Ja0hjlRCc3J7F9SmJAq4k5lUWJj3cI8RDm/dePObVJVms4gTlKY9M8768G
rT8/tqwo/LmCsnah10rfIrzMy4F/qUulpoes/+v+hSH4VdHvud5M4Wob+5SmJKP/bk1H38JgIjl4
Roknpcjzft1/6d3M4POv0kb1IJdt3qz9or4si32OmfgmR1Jpqov6ScGXTHOcb4dlQmzip/gEmB0F
Cik6W3Dlmtmt2e9vvznQD2QrEQxSfciC4R+ujvw42bi42HBRHxUsgmU4Gxetau7eeLoKcpW1RKow
8G8Uoev3JEXWvRGLj8iP63NtvG/E9/UB5r1aIsuYEjhr3bxokt7W/j0KSwZ0O5fO7VJBeY0bmrpt
EN/xLyUuqnQR1u20kmzGKrABBFM4aPgknsht75t7rsu4Hjku6e116BdVthq0PtpNwlc2Wf7xhhWg
gz5VmU4s2NuoXjltXHUGx05B6Df4k/tuTArkif5nRb5EOx0hvF00J5QEFe5YyQz57HzoPFC+u1Q5
ALOYZUZUCwMUjdiFmA4E8kO3ySIWAtjpVjkQqJgs9cX3LVEfj9hiLb1FcGODa6HV8US4e3EgLT4m
SaZahHg9wI9qf2tKDeHtSR6kOF5Ss7PgdwVFUaxN3hH22xDjQ644aigd47vvuaqAB2Syx+1WLHG6
nZomH1zZYhol1+LNeGxJFuxRvbGGjisQbInhpehow5BScXt8pxYsC0JoWgfG6ZPkCpfYXmwE9mx1
bL/g6ATfJOQeRoF7S79C8InrFb0oSjxv3M8iKRFGDQst+iaVqQYy2HigEzctYege6bTb044iLsYE
7a2HThu/G7nyrlniZnxo2Z5uMTO88oIiGbCHxhgsIABcahM0re6jp3EmY6vF+HcNwkPSEAGwMlA4
l6LJHintcGRur4J5rcNv3/WiPBHMsGUhs5bk6+Mm9SNed6zxaX0auNTdm3QFwaqjG8EJNSkQWhHu
O5OdcVxazSzHV66VN02x2w9G/XtnkBTuzhDFpa4dAD/a0I3bgEJjzKBu46tTTA473DETdKfY4hpx
lBRpQGIq4oNZCBWQfn9Pw8hMkgFfr4dm3iRudyCbePf6TcufB6G1LrKIBKdC0zpb+FOMntbZVvXy
dnbcWzLEP2ZDFJdftVWrBTdxxqqG7UF8oN7q9wkZDBYFBPkDuCwi58M+d/2Cdt4Ue9YeHS4vRFKl
I/NUMANd7ttz1TlKGPl6A79hbRki4dsT6BRMe+BdTqxKS24TAoJQuRfcxnHDgAweBY4/iahAGF3b
a1GUwaBnHEDIeEdtTHbX17AWwGZWeEMWzcuPu8y1tU2dogIa1cKkKZ0ythWwLhdaWweuarnnCNk4
j1ftE4doNE4oW8rnm2ouAbZ13tvluE9Qfi2ak+fKzXnCEGw2uMnCG/KOwfpYFypiuJVisRiVFknC
F7VGvHHcrglljZCoHoibNybBOWzIMzNzDIE3cUxXOVI8bvOqordX+EA2or+NgJ0SSJ38EZ69DbNW
i94FDeYPht80Uy+RmvEHO6BrSten02L0n0NkE+wyW4vk84J++IVz/R12JwgjA0KYTyepnsx0WdV3
XE6shkHPaK9pA+LulrCqZGbpEZY3Z+xK0zEyFdbipDTmKJmhhb2WPAmJif0PG+dxTaAayuC9kgNk
aE+yH4RvV+SkutSkn2q8CEDzigtXJ34dyRDIIJt7fGnLkGmnl751ZtRXAvyDhuR72DKs/AAVtABv
JflvNLzR7C2Y7jDLYQqA787BgkxBjNK+gBSisgQJaE/u+mpzSPm5StUvMvsy+gBykQz4zg7lv+5I
EVSOLAEtXn+kHGnn/G/XMuEe7sknDT/EXQLkCULtiuw35M+iZMrCp3k56OMCFeGkaoPijtcsHcRQ
AbCwHTFyiOcygelfhUxI63hjuuXKqOIjAchWHbr0QNAU0FCQk4+o7NoIPOY2qYFYgI7wLbK86g8b
rVwzlsghVf6VYxunYdBJ1aedtwW7vaTI9Z7HLWpPADRqLPbD5ZTOAUxJKSJ80WKLdSKFCl7nuZFb
bAlK5T3VsK8d4Jm8vPY/yRizf4SncT7eYbHDA9y4L/6k+RFmrVLrXBtwQpcdlrYgNjlRjVloLlTW
cEq1EGoDjVhHugH5wlZXnbS0wCDubXN3zfrS8kLR04lk0oGDuSB9X549WwO8QPW+5bN9Wgr2nBoQ
YGjQNePVav0L98KGRHORqK3Gnd1A1w5BU53MAjfKV5dohE5YtP2yahe9mQm7pLwIW7IYRAUnXd57
YxPxnHBPp9hTXV/0g3xqNsmgHHtOizDhiOwGT81DbCH4rSTyfyge/RSLYgIOakKZ5jzQiyfwmElz
xyDOgEfLt3viFRKJKpmvoUqIG1i45vgRgrK+nzHDj0D33LZvYwNhz25IuqReQnNSj7OvCJceFK1X
s9+FUXjnKraX6GmjVtpleFu/4I+llYY6e26bneTHToBSZBWnX4pitBCjzEm618oGDmihDlVB2WHe
m4Pyc8W+B5sQJ3TzJIDPGtAZ0PEclYTFWrxyFlJ1tWwXIgHKVR3/8Tg6/hE3pAI+MeYRuyNOdF8Q
rMaUHrxFaYlnvtaQuuB9gAGncxjDTyCQct6dHgRWJ9ZgpfcGg40sKgQcYewa89eMzKTud5c/7bk4
6oTMVRFLx4n8Id+cWkRSgigPm5uBN4LKDSpEjX8dVviuFLXbNcKGgZtibQMyrdMPDzNqkvqAyH3X
i7ljvoHjZ27kmHaF5piY8gusYhmEfitQWFpeEHgan6gD8tmApKutTNUyVN1tqerO9oi13ZekxXqX
tXj/2EhPElhYwuNUrAlQvebIK5WsNNEsn20n/QaucN75GHXsM6O76dxNctOVuT3wPk5uDWrFL9BB
XBM6lEkP2AQWkt6LXVskPtNBJ9BbZD4MOctSc542A4Bc0+1xUPDJbare4kiGMSCoqk6Ko5mYkuRU
tbJb5yq6lFLVUNEC8HP+ppH+8fB8//pljA1lPlBOScISCzXnJdqKGRvKBvNitAhkkh44GO6UaSyA
wCHI3fPs0WsX9ZHh/TPs0ryCRaBUStTUstk0ggKDLE2bCR9HpuNfMl56STSd30bT5zroMeztmY61
AJGcW4vgoj8sJDgxs6viamc5h3YmXKeVJMeG5a3cppiEPujRFG4fSIVjwBPVstgN+ETwYDi5Ieqn
nc/C+6Cq9zS9jauwRcM0Oy8MhrwkSzBm1Z7ILtsd3+w+4ub0XaoCW/1Rw+08dlnD9hZCore0MxxJ
paDGkAP+xR+VuMs9jsfpwT1k7+54ypJwLtMYwBGS6ApNoVpTdxOY+ZB68LrTywkdEFIYOtMWQwBn
48aZj9OgZyENTlgVaC8azwzTj/lN/srY+aAXux3op5ewBtw78OTmnDVYo1T2gbw56JieLXK7RQAY
D3r2SXHRRDArej+dcoWBbeZlnCaks7rBjoPq6oXwOGmnUSt/QPWOeiLpboaScWKGCutQspORIOQS
lZ08AaEMdRz4cm4cFD1URBHYQIwO0sQH6/6bm4ix6beAH9uS5LfknOaLprZFKZBmtj2xrOmQy4Yq
bIzbPTy3yzMfOGwgB+ozOKrjXi+KcJoQ69/psf0rOZDbJgPmUDZ16JAKlz3QbflhR97l6eK/cYtI
D9lUBKsIcq8cnZgms9HvCKFkhduYYnCBQF+aeCtIkEZJMIy7kAR7zU1jFsOBKsWnU8iq3Cd6eZB8
+J1yr91xLwHk+jaZSSC4mOzv0/DKsmaZ0KhXnUBPpHQ5nb3BfGlgvoIUOgR3DszyhorkQJoTgOAN
8NTwl49IMUkg1jAMFg1de0wSTa1rXUrn06zvLbMauBsknp4WXRKltBLvjYE4oJsmNx9KSRxfGvik
NFxK/YUvUawXgTpXpi7d+txwfXTNteTkPRIT+3KLdiQA4xd1AQ86BXMyfHGBxwnfYhvS9CuhN+Vx
npT9OAiVziKtLyn3erAFJ0T8k5KkhhWLDSU6HF7ksRDBKFLTP6e6IePYhe4PLfKWQ/FdPFQ8Ehuw
I/Do0IwOCJoqSLaRtBxAIaUwAqpRkjDSWL8Qm9V0T7o3cV2NIhZoG3konkV73bvsbbBJeWTg86oS
/4VkH4BZiLu68XFsDDY9U0d6AY8Xnjz5Upt1V9cKTAdD56yi5/XG+3u8NRwzb+iWhmR5PGy/QWfs
Q/GBjEg4q2r8/Y0j99BIhZ02tsQPbf1ViA58Zo4vRtQm6kuBvd+XWdTO4Cn7PsrLMy6A78pzQIU0
ChHr0Ng7IaT4ToQQjUwJn/9Nl7t2lvQjEI2QlZbltXVC8QZbZyObXWo220W06de3RilVQbLfpzW+
0B3Kdp5lJNWX3BGV4mDY7sRbktLTQeuOA2Ar3/1KXiWO14S/zSwt/vGbbSU827ZDGpUgTTy711F6
n5FyivymRoT88T+yL397t80/xqjNuxz/w3CSv0csrxkP5ccaGIKEY849EkKIwRWcagwl5AjQAvmI
dTN8Q/zliU+SkcdN9GC8kLcDlFNy9ACSG9xCtG2kTiNcTg9HlA2LOoQkO/hNQMt0yxem/dgwWqlw
i9dd3rUtXCm/D1ob65/J1qa9wnM57IqmKg9fUEES5AZ5F9GG4q0/UNTm8+PdtLY/ZST6de0xLTru
hThg1sBGq4m0M+tTYSXT2fqms67g//nsvFJMIgVug7JogwBzHZKB5nOcf/1weq+YXEwdNPW/CWXS
g8F9vvnwjtBkCH61/XNX1RRuMSoeStdzUwQC3mV5gpkZrdlX1A4iLE7S6/TQDLLfE39Af87rxy6p
YdqiRiVzZ6Caqf3AjYxeG1VG58a6O4Q0Tr5DoXxxR0jdZKLv3Kg9cYCMq4GGSFW0ohAw1GBMRgNQ
fa+JrJl6ezvDajF8KhBQUwfTOJPfc5d6VJOGVbS3iFjSsaGYDQ+L30dPGSm3AUVtR/UnypdIClVy
LShiKDOQlusudpgEwO0urNRga4K7dHkozsPIaJOOTlDo18pUAoy1YW5uDnD1zqVwcKn8obCRIF03
PMZuJOW9ev31Srr/6u3+TnJE0q405WLmbou/UzhPXlTmZuVJrDnSK4Q+r7t4Qo+DYjdHKMeBDM/3
wGokuNZdVrp2Tp9ndKH7+411X7oBWLehxxYNjwXkc08YoCNbalHNTScDieWtvDMV3GaKAGhT9JMP
dDmUeRv1yD19S5FqZYSIuqzirHRE1N8ENTQI2G4PINaT6o0uxY+exslGVqzTchChHH1djIHXFAAf
P503PDOtXLeE1Slk+ZxhZfuNo2K9UtUH18qDNZ4FtLF4LV72EhWmsIDG72IBvQNrzRIDfJFDoYoh
vMaQPaHdQ8et8lJ9pnb1q7C/webpLYZ689evx4p5COWrZq2IIcMx//1Xhkn4xRuCGYFiqxQuAXXr
rvll4HyB2Jo0B+BUw3pF7Sc7pqPg2sW3xrzPwS+vj8kc92z9AxlOnaIc/CkbQZYo72+f97HWqGBM
W3u9eMjqOEpuIpucDZlobPhReko+FLF4nu13HU5jo43MLhqLyUhgSq7PcE/6IaP0RNRqx8LXnACP
s2kbFFWZhl6EQakpceC4MNzV3pZCM1seMej99t7gmiBIYOqEjEiOiDnnKJviu+qixk2dtqKJipsk
DJqtexPWlYuR4e7FRJfSfZxaJP4BWN8haqNjTn1H/N8Dfk/R020dVdWpa7qK9nsuuS6WEVO/CqMd
UzgCcE0iGm48elR/+8LQKZs48yV//kw+rjglFiL1+OWH6/WZ4YIkvm8hHswdxfh4upubgJ2DAjRH
UtS+a/xUfhr2yMwbAh4adYamFfIRTC74E0XLLsDq9PMbR8QVi5YxIpfMSgWddg7Sy9rnDQ3HdPQ5
R/ZE5NkHwK9cT1XRPNedC7xEIICJwCMG2P3EaoG4qL19rsQVJKt/PvRLoKc6YhC1pHUnXM7yB8vb
aIhpseYRdt29EZ+cA0VB5xbjLBrLIWjUTEVoewj4Nxh8Iq7VjHKDSqgIsNSSay1qpyfn7xKObQBt
gxaWEIvm95le7wNNvFSDtktslqH2fVipQZW4ZSn10AKIRAbdljyIteSkLrguyxgj/mer/sOGKmkL
56vlww05ZwIbQ9w3d0LtDO3MEl17Tos9I7KXbSZrhb8b9aoSr79G0r4DUlQlnZ/HZ8MVZhOlDjAf
kEixWGtkXp1o16lQpnZUeCghddJO9Wmwi6BZzb8unfCupYJZDySTTVRa6DqK3vIeh6t0XtFz9bgl
SbZl5MTqmDIrsX3cl8GUVrwIJMHpS2y3kX/lP+NOX+wjI3yEENzyT+imhgorVwP79XQZITLTZ9nF
jONHKA/SoSS9c/TUiWb6zvuFzjfhfPRA2MnRXm6hv1Zc8lKucPUQlTp6gsuyEN1JxzCisrigcSu0
MOFATnrtj5ROtFFQ4BkEpARzE3zndz2o9jW/8bXj2NHoeLHfoIb7IzNkt4jG4xejaj8bu9qI2dhI
iJHT4D2jrk4WdKDWA1bW+ENM0Tgn2FoCkuqh6DIgmwwG11/hKxMhre/b0uWA5HcP+aUYXmZd936D
2MHCj0rNtLWic6NuVwctkK9quRNJjdQLgZ6F5bmAnJTBZQlvcgS4BVXQcx3SMByztJ7SC3nKm/Qy
bo/zp9gGhojyS2fWB0spA8H1H+NVE8ZKrtAp8DBrBeKGiqlITo8tK63QZN24NCkrfpddRgLL5KBd
fYv68A5cZQleeBlo7h7+oI4iZrbSLp/rDSBfcBy5+3mDx+VCZdzOFFSKYih5WCHACYDdshwqbNzz
/rx83EtozuF+9Wh48mKoThBJjXXzKh2Xf/B1Bd7wWLy+XB7oT++OgIHcIotii0CeHa/zFaETe1Fj
tPVPmFGgpxy/xaXvDXrQ8WXIVuWvYT8kL/7J9/wrotO2Kg+RZTNx+AFiu6UAlHaxXdmq/kXIJp1e
lp6AgfCIuxeiGyiju/h55I8KJ14bL+qyIpOtmnI97E503oL0ws5PWocevYAQlb4xLPIXxEgg9dv2
HEkfZ+n/jvh3AHGh6Bi5kbCn0omLFNj58Fh8H+rvQc5KeMHt6o11C4i55cDsVulaXREJy5nIvp0Y
BAzMhhhrRelRibl8wvwRqf6NLPNE7ytt8juVOPV/N2z4BdDRTrqsb1OsS6j03/E7JhzlzdFvLm8j
Sd7MwGJcgEXgH3OdmLJawKzEgk26+BDTqx738WM8GJesRXRHJlUXzJnmRfodokX/jmzHIgflKguu
AGrMBEJ37VrdMNhpa8uffsbJvqxOxf/mei9WSsEH2fPnz+VmgEvh1xr4vHmih9nt8hT1hSQ7YVyB
9DnIFKrZlfEPH5OL1Jpznc07phVV8AYEm+yLR4C610kfs+QDb0ClNSL44IYtu45zlckn/3KKAhuN
0+0lOpM3u0KgxazSZQ8noTfX6cFTQn5tQhyV/AnKbnUgGy2E8ae8MPBhqWQTrw7lgJqc0G1ZjWwG
/FeKsp5ADzVPu2GfLTwZhi7LARGz6LJmaUUMx1/R+oPlICDhzv2nAJQ8jNVjYx/gR4bigiv3K/Jp
uMxW2DVsq5kPHb2zsBPBiBKHdyWM3EyH4M0phxTi366KQTHTPbmMUSbwexkBfud+0GYVe1CiQ/Eh
iALfZrEfqGxWf82NFvVOUhV4gtygjqB+JFt3BTUV38edlnJpgBMNxfqxyBeqOdt3q+XVAZeZWBYm
wwUG6QHlISoCBTOL9gzrp/WhLk/wJDHC//vn7pU25Etj4UuPwop7StyS7nsLKCDuQi8eDccSFTTj
A7ULn8V+ZcHqszCbkW2Wt+fZMFtwDWsJL9lk1lByAWIng+oHBLS0gH21s9pOCSNO4qWRAcerJCLw
sQVDFUNNLCrvyRI/+TrObVZS9lgjfm9Q47fWh1A927MjJTL9du7encB6MzBY1KwgA/RkCO5RjYsg
j/GdYVUA1/+hdU/m2McK+vs9PC1ZcxM1M5E9Nzt1mxOHCpnFwja5/25OxbfJYSOMMMK81y+uJ9Kl
sBBlYifxMXE9HPER7SQfqDHV0FbaXy3v0ye7TIv8WdxEbsV4ZYtAp3rysXjf7dsUiKHZdPfO9TrN
0CKRtHgm5cmpzXFwj8TqBeJ2M6O8QajgV4k7qjQL0EqiNAY+zWDOyEZ63WAXELmeS/XSxiJE0Eng
t6DxtOGXC7N7/19sUcJegKwy+20M0vJ3FiRzvvFiUdb6q2wa15Lbw1ES+S9FmSytx4cWGl3GmFe+
40i2GUecNHRUtGwBRKn1B6urlrERAOI1sjPv4YHTptjQ4NerZfA3yc+HKB8u7mk6va34xBu1ykI7
YNUeE3z4s09QRuSeQ6SzcE8bUXEdA3rXmhhjJzEkpfDAAKeIFjgGS2FblnbMkowznqC8XiDjEw35
/7OYtPF/s2sOB9SxhDAsOyJvDz5hXC8Z46NYr9AVdSguc54afXNDlidhWcW7W0pKy/eAB2Vwp6TK
nEBEcU8U6sLKpT+0+JuLpTRsv0azP/Ltt6gU56CNPOboMHCyLjH2oxO6RK8FqK1U7vdLiJ277Lnd
/c1iaOZp03UoJF4X70jj+owQVFFqC7fMvQqHJQHLHrC6GWKiqw2xstZoay+oNmau9piMZ6TOB+bz
oNdJjmvot+a9QKmFVf42zb3hYXgEoipVDv86kg4pBGNU2ixh7oYUO7Ih6lp/MDReUPPVa5MqLVjz
3TF1f/VDHpEHIhbIer5b1lluNMG/zxVcuzy0QZN0UTSdjKJSlhacWt7yFdnquUPFqSG3U71WmesO
sSkAtvoFYRvcnDHnuaIDBqUm8I4hOEBK6Hh3FA0QEwg3IjDtXvNIItfpvpm0He7iW9nxJZZIrgXx
et3n5RUjqDmJS3kal/x5xXKjSLcvN01qaJMb7FPlsnzDSh4fNpXC3r9iBbII6vGC+m4wC9bF38az
Zv/a2UxzAEzXGeAioLnrsRKeh3jKC7QhgBay5SFULKLvfuHvAzG+qaAwpUQ1f624SJFM8PNi2T7a
50I70MNu7T+On4SzmOoHawUoATFA07soeabuWpD9z7plrMUg8f0vW4SHhYJOPfjt5KMMbWiDHQwb
2/EkXWfJVCiGh1qofFE7g+n4LcNC+unMpoOfu3ygYzYZ+PNQsHth3qHXOSxqhOYT+WJd/AmRszz/
j3a1j0565VDlAShSQb153FvyjIzwT0z70YoYsFCkdP0L/umpnzzNHCDDaedF7bNc6FgqT0G6Zvun
8M3HvKFbhP1Y8XijjrPpbZk2B9ObR3NuBzZj9SEcKkyaASo9mqsLmEvGtSPotivSTt0wwKO90shO
AVYqN/gbkeIfC72m9MEBgYoQDTAL5kWOk1wMvAUjVm4H3QV3DGSGuDHY+aDT1dfZ7gTpNWi4J/VS
fx552ku6rquNnf7LvhSCICLkH/HdC+zrK1Zm6b7Oqolw49l0f3E0Hh5cNpWGgfdvUcGqDxPp0cnh
ssVGg2OJi0nRetHBhE8fKwZnoIjlPSUIFFRToByb1U6L2Jz5/CcBIDyEyxBEG46Of4oQbOY6m+6I
qWP/NxgpqMWh1URSxbRRmFhgwSa5shm2SmU7yi+hgmR0yPU6gTSNLUUoYgu/uPScS1vp0xsx29HH
0PY1wmBq+8JZGAxy2GR4zHoAAKkVjBIHVBn8wIQvf2tUoDODyvEbnPg76bpdhChDjbeSOsmXgSUw
yjt0Z9+ZFrCZ/6UHJDBD5Ti/ypQMnF59Xs1YB41Chn0va99LwSAPii7weo8JWqaofwveX+N2sQwC
HPdrOCEusqAXG3+cwdFiV7mQuhJm/iA+KlvYw8MIHzQn2MotDTNiP42Aex+JFzjw3VNhGr47SRnH
PRATv77IF2qyQPgs2vluZXAmHpqZuNQWs4ixIrbQtn0QkJl/0wymMVGSFfBNkhx1G6gpuM/vhmEr
RqNftSy5h6vIh+kQdbsn0PWv6shqotIvhrzINFLQpxqkNwYwmYw4PvoePC2F/KMVBNwBFzR7f3Ag
fWVJxkgpr5t27TGANJbpJXQ/H2i5fIOwTTD1m9YbZt3F3ak8b2zvO8UjcqPAffr+YMfzLqm2fDMm
VWCUahQACDbpZv0Hqx8oWxx2XcyopJo9PmHUFWS32HAWPZuQv4Jzg6rWYyqr2jGqotoUPtscupwf
33YXwxEedroET1xPX+eDLCWjrSo5oI/+baTxXORd2tmfI1vkA6dmFXJ4lRwaBUvV4H/2Y/1YJ8IT
s1wL626Uu/Um9WdInPFFjaYBbHxxcYEOInDY08NyuneZjAJETqbos5ZyIm/bKvisgx0xy8c51m66
JX77FazRw+k8NzomFXcuXW+0eNeoTv/ix2kt4Z9reBhbiqMEdavBr0JO5OXFwfok1xaYgXf/KbaQ
q26h67HgG9+w5feKq5ZlRw7d3DEgp8pOaXIxur3Q5kCjlM7wjnNtNiquyYPtqYdgy4C0J+etBP2V
m5xDF+4WkbUfQQ9IMsnxSXtPpL1bYgXpRqZsNkla2qiiS5keH3QGQc16tddCzoMFENzyFOuh6X5o
pFu/Wjj7eh7aCRjTdvaoESIad7khCacByt3xBvlJfOqBQB9MAhXN7qqiXTSYro0CYVwnfodTlrjp
JDCjwq4Py9VjIiu0xyoeq41KnQz7CK43YLUiQw899FPWzZjEgtjszktNLmcM9uxrvGFOC6hpd7sO
+r8ALytpX5nWT+LZEpL3uFx9YYsiWJqlKMTcHxcFbUbqzmB9gnQMVbVN4fbCw5k7mZHkCifnSUkZ
ZPe80h6zKIR4xn9nveoSImG7QY9LZkq0dR5SwDBcRqFLPW9pY9Kuf6+08frrYPhc4c/vCfsyNXgB
pCA4oxg5sEvxIODq9XSwdlYgk5PPIGoVaNtV6yC6I6bLFLuq9yjRLIi5fDKUJBx+3YnU5OuLbErp
QsGw8UFYq4xGtxVI52LbGStws1IzdsYPIp2xfK8xtMym5EOSG+eTh8qVJbDVyBhXm2Iasy58Ox3q
qdVjWAjNccobplYgYcNjDXM/+3/SfAAQhYcXGH9BZt0pXZ1Ix2wPH09dfTM+pboJZcdBfzXcLuIM
pnbOlSXElo/V+uAE9l7rRsXAV5gVte0xCirRDaAmS68W6Royy94WX3hoBXDHFqpPZxQvW0tEe4VY
xrqXHnkUamTXFTMV3FgKZ09Xpaj8kKXP2r/KWSaxqemAtmny7qUkrGpASajIZu1pWZ4/jLiICZOD
MGI1I1Ys4LI/rD7d8UiQSMpqOqvMP8VTnqj1Dw0lLno8S9f91nG2kpI6Czl/qEwfwHuKGzwjjeah
rMAtKJ8QlqE5KRjhW4sfx7HF+KrqdLz/WpAwlNH/PsPo/OceowJUFIkDWZekF3V8gk8DoEIMwJdm
6/6owbwFYXPUIJ1Xda+slfYNwTCyoXYXQKmR/MNNsbwANU8KeUWjPgFaWP4TvyodEh2eur4M69Hl
mleS37eztJZzhWn9h/fbCjft01pE+PaBa4jWZofMppNE4dvz0wiczXElAlFMom1ccYc0bVlDVfow
Qy/CpqHZwz0E4cJDEdvXQXXiTXgWRykZ5w9rkSpKYuWp0hpDWTmuxqs0CWAunOp0wPG9gHHkpVg/
FemtXXV9Bf75sdit/J3xkvM3lglvQmeDQ+D2mGfwdUG9oxQf5dxqG7prxwPlo+JkqLwBAfCHdkEl
bROMRqrUnxAQmyZxoQU0HowCJJ+VvnYDKIsU5I4QqwwR0KXQDl5yE+EGNfpGirqD6ICKo4bAsRNW
eYIjkLJqMSgIYQ3lCdzAafN02KUT6wD5c/ZepLXMa1DCXcb6ayHGyt0guz+UgvJowXhU/gXM/qWe
ywfToDE0cddWXHVgI9odUCCARbdBYPkuQT6DSXz+GvWje7IfW1O7fQTDXn+SWDFT+JsVKpsZUI21
dytCmMaXft7nCroFdLKh+4uH3Txq/uMUyEwk82EqCBA8HnPDv22lyk1vqtONWt2lJlYdVQON2gS7
1kVtnJNLBN5f7CZuTjrPWPkBF2p2veBHw27O03NxQ9uCbb18YzKQ/+CCLeEDvFsqNls0V+chWMxB
p8SXIINhKfqW6lWlMx7mvLTR2r1xjzBn9TBn9BN58mxIT+LzOIVLo9pt3+Xmlvfn5PYiZ2BxmHyB
rivHtg2kMRFaZfNA74eXQ3LFouP0RbjJYBpPNQjmFcMTIh34PIdiFCJ1vUGdef7fSPwv5USFJNkK
pQT9X8ULsDIKmDXbf3Kpxv+8+K3fC9a82WkLibktLUkds317iiuupk6liDgg1d3eF2F3UDHKAl+h
u2i8sWCym6L4Jbi2R2I1y9vYTSVP3zV/fLRbeBXMh1/jKyBT9enUDGuM135R2ipqsQCzTRVc/soI
uTB/V78PPmDQFonDGMhSLP2ffGm9eXShFUsadEmf3J0i7f8a6vfVe4tSxX59PRG7wb0SrqkApg42
AR9tBjJnxFmBxVF79yaj9z9uhgW9WdVc12sD3iJShANFOu2xbACDc5th2Z23mnP+5AMOgl68tx58
VS3S/U99gF3zRQGt2DJoV5Qpus8mfIpTH9D2e1S9tVWhoO59Yi1An7RtNB5LA2BoSAqnI6mbjJAw
FfctXs9vx/HuVcevsnrqkSVIub84Nxjo5PiGPVT/VsEBUMbn8Ok0B9tq8n0aBETJ7Pc9lOh87WQj
o4RvfgKD9lVN/0e1YgUR2BlHyqFoxGuFaeaLssCccFRVYFsjenqOSnzedqrqN0Sn0fo9i0PacxWu
XNuuDS4kZVad7thHNkBAv1/g/FMJcOCUxkoAhOJoHWgKgHe2uyLxNG7q5Kxjionj6EgJ9qgonIrT
eg18CC0s27Rjmqwbou8X8uDXe4ALJkkhxQtIqmtzcLEHLhtKA8AfxvBTRaRE3IFR/wCk0LXd5uT4
fry3s7psmw5PSDzu9QG8AEUA6HPBZI0GcbxlZ4wQdcx7SQO4wllRnzvSyv5mhL/bZ5IvSU23DPMp
iGKorbe1QjYSQ8sfVMMuimwF9/AWV5FdCOHgqYbE13/X2SZ9gEhUBLdOg8C85dGChWndb/26nWd5
3mB7lzNlBOKF67/dGfpcKQRz0NNhIZltDvBYml1GpbDxD42a5yfymcyDqk0wOwzEp0uIaIIpuZoq
erurQ0MQsAq2QZnrd7Tay4gRK3reLfLFaFvtrJQVpjhTtsnkdU417IglcV8ZnDjIfTT8iTAFLxyw
2VQJAWZrXF9xbH1a927Qto17ZpXk1P0vnqGUx2g/Rx+bhlnjGjhBqKvxapLXzQOWIPeT0T+lc1L8
LBWbyVYcSInvkpqtXGwmIIVf35ZJgbPL91MI+IIS8AFrFUv1hg3concQdF5Pzvrhb2pDeenedGYn
gcdF5cZqFSv8SJ/KlvLMcUgQS+tNnLm1mpiD3HkqRp+yhyoE23e99jPDoDmRwNletZj6fsh1Hpzv
MOEmEIM59U42Ruc6iemUOaasu7GcC2jnIg2YSZbGX8YPH1K3hWb+P1pwHzhqp/VZaZ6tp/aDuBrs
dPGajWc82EIdhot3IFoivBcN9JHWYD/SqGJizEGb6Ppc4bxZHXNUauZxMqkDvxhZDJXwW0EpbzYz
sDCkD0fOWHzJ2Yrnyn3ZO5wosNOsB3ASXfhUefgN0O70B/NUWu3EoiB4Wa37sGoE0lhRUcK4BHVP
aXEKL7Dk47EtbIIl1JrIzwnwaZNIJVaPCwRu8iOW387MpBKIDxE/WIOpG9OfiLZ9AAJB9oIYyc5B
/5GTdKx6dEhqjadHV7CSvGSBMsSk5NGnQSnPZwVsPDsWtNqZsFDW0wk8MgVewcr2aLCmFcTraMZf
Z0eEF81WWPTwB5G30OeA0hzNhznObJGmToRwe27cNLXVaSVjW/DYda5niJ/43dVeYHLh4Pw8QIYo
485NiKc8AOBcL4ohRiQ3So2efg9XeF1oC4Y6p7vjjqbHDwTzHpLuwAfkljyuBoZ+LF/i8ABbFtzT
BQq+gNTH5sCcTSrgHzCtZ75lNfwr//JHcrB6BbbwUWWOiFFiOMhv0oKSn9YU9h9uxGKkJcfBlvtr
rksxLgHuKMkl3IPcLXkzhkRgaMn8c8E7Mw0a8hI4gJBuhfNe7+48R7ZDOk0ziQ3qewM7ZzXVfhNZ
RDYjVpOqy/iyGGkgVzA2KzO5yxLi+3m3zwF2oT3sERLBssrsJ0fM3QOIw7/Z06kidi+jK8T+nn4R
q2tfQyB9gBlYpC24bwCafJ+CsP3rbxnS8Sf41gWftk3NuZNJi+pH5PHFQPeBn6XHMxbr+YShHLvh
F01wzJ2wP6yQNyV1arm9Jaj/dyXaAFjYOL6jb15xkavP5uySa4DE6Bh1+bveAEooB0Y+TutKh/t0
fo+HVRgf6j0yOUB0n4QXGa81jzHO+k6U0y+6mSnHv9pI+HwBfV7K5wQCJFXX7ekPNHELt09tuaPr
urjyM4I0eowL4OWX4KWrlkJsftQTb3wABpqT3v6rFW56tMm5aOC7rX7duI5OjsZWtMm67UlaY/jc
8vOmgqjkP834nh2WqG71pTSxdeEnMjtUuPzeYDZykID2HsssW1TZ1Ik9VROMCqY+e2HwiZS/wJmD
yVWAWzYWkD0nAwTb3K9rljO9ztFjupaKDwS4P4xbAjuAsWYqmqmvjWKgbQXfOC0NH4KDcH8Yu/RD
6OV+KkdKzm2/OMMOkhniG/8JaQJvKt/iiwGEPwqGzswyl+ACekEavWHJIdhFQhSOFU/FgijivMCu
GMdfxPHr2hwseQKl+EaMtva7MpAdJoyBlq2/6+1TCUNn37e+RILG5ElPY6oZLo1KZiV4AGhdImCF
HNCBBoOdD5NNb5NsEGUhNcPFy5vP70AsX7ksSsAjsn3Ol/4OXtHSS98ECK0YrxCw/RCvk7VLfldb
Ry4EMNXheKfxzfdQON2rV5ppLKv/6jvq3CCtx2Vjspp8P78zn9y6u8VsU6foCfD+bFTXyK0Wh5qw
UUQPHtNQVx+h+tHXEduICsnazl6CoeSpi2AT95FzxpwfeXh6nHBhhIHM91B8mDw4Z38/Jb2/+6Wx
zliemxYOfhhFMokPLu1WaZJYoVoQVBAHMmy3wUvMGKhdl6oMa0Wnu25vBVldTn1XUMlCD55i5uKP
gM2PFV2K7ahKD0IT4a43r8LwzgauEO6kpF2InUgJZy4ojND+0zbDLyT7ETzxLaKgO8sOyDe6sjaL
hQbEvhEoE0ti2v9HUHpUqInR0PHy63fdXtOl8hNfMFPnYw6dZe6Oc91qQugWuFMfD2WbmZrL43T7
dO/fmld8op2+BgrrrilKS8lZjQdifnpbGwISaXmKzjBIa6GJOYcNzrLp0/MC1jAIgcbK53QgGodr
ENGiCJcKui6F7Q6fQyNpv+xvqF31KSaaSw7feV+K6Q/ObalId1a7LNp1AV/KUW9KxPEIplbf3lBu
Vx+/O/G7shga3p09/t1fXtzi77JV8iCPoRaHi14EEb64cjsP8do878vy1q47mOky4t0X/6s5sZga
NdTLZFZpy2b3DGyImDD6ni/rN+ZAEulewkd5d4fm5Sp8p0+O+5cGCDsUx8n7YfFk2BINvz8C+ggH
B8rgvC6XMHVIFWGLJr50vRwT62AFT36tfoFF8IHUQ+NtAtkMsLTmoiLyptOOBEKbTPOLGq77/wN9
xG0s84J7MBNMTFWsDmCNcs4iwr4mx9us2CZ9mEw7o3oRjlH4/y9OsAL+VyDF19cHBTL39uMgCsYe
yvIYPednw9fndf4VGzmjp80JGFJOu6xa1fprrp+B+4L7tLnMYUkoa6vJK6HX5a2fCzfOMP9OnrHH
O0yiodnpESznpu9c/HcUwH+9BqfG5Ibs5O2owyGfckVI7aKQlaDLWcqPUjPDJHXWO5SX5Y0WZs9w
CuHvqbrzdjK4IbljeA4ZD5+yPlwpliT2VjxvjNfWyfh4eJVCOtHkwBHo8fd9fY7pEkSdvJcW7qSs
MIL5H2MWg7Xji5/7MX5ity8hMH/luO4aCDymXYBRRNp91UuAWpvOI+TW/VGMP2zqtrHL/Tb5qEUo
Y8D1vst5LHqp2DAX2peQTu3wDRAf78nafZ3JkHCNBLKvw9E4tNdfeKeUEpIJ+7FBnpEibZ/bsszz
eHuwUT4Z1m+1UHRybPSwAypSIHcFfHnMlY/RsXHBU347h1D7GQiz0QDMe28qbX17ln6+PwHIPY/D
9Zjxju6dMg4G+gIe4LAxCs5+s/dQP4D0nwRtY8YTTbtNoz+x+656OuJTpL5NQ6CFGTWt+0tzv1aS
h55JsAeLra0DdMNhi/oty6WBg7p3oRjrnbPlQETdSjV9RLoZZxtw+qKjV+J9cMHFQx2nDQLyFTNt
SnUFAKERJc3HY1QpAhmUvKli0uMVLw/o6ZBmLRvrefwoMG3jtg2/MmtUoNJt/qRHWi5hefDIxriT
yTUNZCCnd2zoHP78Ilz54VacI5AMApYqIdCxvM7dVmcTfsXIUPZAQwDN59qcPdOp83m4qfa03h9A
t7Y4fg0JK0p2KnMSdTmKf3rNw4gRDROtnOUYn5n7VAmxZTpHNGYvjxKrTSB5tz1ePLN2jwYryfMI
Z6n/zOZBxgKa9ehiVVbUcEdx2LpR9/lD2ruSB0PM/CGFDKfQhJ5UZrxRP3kzqumpYuFlyD4nVszU
+k4bohOWcNKxgxYWy1MF1oOBUyOQ0zONfyDLc/9Hm6H1+anbTNpBI4/OyrtQZnihC4S8vE9ZJcEB
zHs0bUogdLyRL7JoTtgAFAFAo6Evjv1UDALkqhGfpIMgDR+Qm+4WLF5urQFww7S+30fFLBU6bWkI
8a4wmd5k6aSqIAmS94rvmSdEAIwTIs9vU2BxIUjvzwJABEJbUJHAEe2hXY4DTxvWnEaIHH6NYWYO
8ICdKcXDve7mMY8xesGCvfwWWk6xRG5ISOjQ4VknvUslt8k5Txjq7crAHj6cdlZTEmRi6y0/rwKN
7egyP8nnm4TIhINGKlZZP2IOr2C/Ih0Q/skcb4gA2VmJnGl5s2cOg1rs+0rvbKPzibGJr0LhMXan
fUDNAYtzpn5bfNo2TC5+PbWpKs2HUDgReVhpUCk6NkmUxbhBXApq51QzE0JzayaWxfJbtiuO+kl/
1paRHXIEnnIPCIBJUHoi1TvWawy3VQWkQdO1ADdYTez5qYwG2WzfnQiePZmjdFUaXARR5xOpnifa
/yzXXu/BS5vm+wQVxCFLBgWKY3qe8f2yYpu1+LEuVimANEY3JFRt1UwchtLBPqDnAMAp/zDTzxrJ
+pTc4jtxVlsiu7o4CEOl7hBD8+I8RfPGzOGVruA3o/uy5J0QLuE3fI7FwYzk4UM2kCz1bon3IS0f
GG5jK18ZLn/yMvnmMHcBjGBNLtTqcU1RWBsmx6zi4T1UcDqdbw4CYp+gQ4Hqk7BPALhzvwPC5FsU
hN/KIUNlS5wYmAKyqVZDZOeUJ8FCfI9HlXJHqwyK0oI+T0/EotatBZ7qWiDp0Q5aqnNKEl3bXLP3
rC0t5Q3zHRQUSlhFbHm0kEYLMYTNAZu71E3UPBy9LMIaoV5D+NQV7MA6Xwtbc4rxTP4Z86yVeY9i
1gZzar8ZPP7UV8i1s5fPTTy1oZgWzhwRmZOhB4hWRF9I3aGmrjNPuA2W3BtdWv3Y7zUEnXJ3Z0QB
RgQYoRz8qzPsUe06EmkCMxZ9ATk0Pu+a/Sue/I3/cw8X1N8Uqqbp4BqQuGkTGNDj0GnSvIgYyIkD
SNyKth0aZmAEe0vjRYbmd3NxuM2AFSh1JZwoeAzUe6g7U5a6ta3Svoa3Wyj1GaK3TWbA4ZTa0rA7
oDH8kGh9gShgj8YDoMr8GQc0umQbcV4YALw3lTlzPK2z2Z1TksBtUPUNC5QN6thCL0OH+pzWX5JC
sq7Ts3tqjIzuDY5J53f+renAbPvavzAaQXBtfNfzVLp+ONHPO3O1hcU1R1vaH0iu7pZHQXqMj0ia
ANIiyfULcyDXYzSicLQOVx7auONRZ3ov+1QIM0EtSSjgixkSQT9jte1SGZJ30I0ouw+PA+ETGMFZ
41JK8edeU6gDafcZUcYTgacIP1fsPTIVwylzKMtQsA1fkX42w631/0Pvryoz7nk0Dgw/SjPCKC+3
CH3kbxU5eXAYl2QogHkjfaWjD0zPH+DOTKLTKIKul8mHkHOFgAI1C863O5QtP7hnsZGkL+93ggzO
o2ExHDIuKFkWvU3HfjNipRacj6BSa3BCc+ztQci/4woDQ1nx2R6FEvqR6P1D4/yNBDGU4+f5pwa9
3I5qDH76bzthiDd0ZW3NIOchjJ/xK7OGV1dcasfnz8l5/sGNpmnp6d6ZUBjEJMlqrGM+S7AAsl4x
GunOdZahDAOTwNm3/n6C6KR/Q+0J+XhQvkJuRpQaSmfYqQuKkWhh0eU+mbx47Af5ttmKZevsHJXO
zKUnql78i46DihgwQIkNCannH391Lch54tmsN9hYoGFGfwzPl7IfTSwlwh96nv3SuYSD4Wziz4SM
Uhon4QE2CSN3/VhUrd7FtJwVqfUBk5PWCjWJqW6rzLGe7mZn1tF/E/7OiQvcyyclSt87MzyHjI8F
lSs9Y53zJ23JYQKZUfou9m6uujZCMrzJkDb3EnzkIBDZcC2U383T+SfYzbsNtK58LBHNmebeTGcS
qRuDfb7EJTrWI8Ytc3i4UxyHs/xWNCvOc804bo1QWILsdmw+jRpCxivkZLbAaPI87fjOJQyWcraF
NPg4AYDZTD2V2eyD8MXk/VNDNR2mkuJwvZwySrMuhu0jjd0Wf7ExQ+NZIOYie15ZUVfDir3FSpwW
Lxnll4aNxLneQEJxR8riW6ZI8O2iL9p/KtPApfCOAM1Nhgo2IKJUEz/9fP7Tz9zpRmqD47ETxKzb
qt4yLmayvp50Wj66x8rIPwIm+Nt32grrz4qk/hHxotcnO3T5GgW95tr1tfU1T6fpVXlLe9HrZFTe
bSm9q0r04hQwWdHZ2PczCV5ew3iNSDTVE4a/d2DbHiMbNC4LykMsumL0mb1iq7HQbXhk1vfqK+je
gbTSBLmaGlhUItm5cseylnkrgOPBFlyh5reXT6bQuNoPlIffJpmP8+vQaadEubdtMiaEfo2r/9M1
U8Hq6sENO00QhoS9tTTX99of5M8oXi8A4UEZSjFJq3djDuEsNzxc+ZNRMyxTJjiWAESCUXJJRPc7
fumc9jNqYZ5yiuTRRymKsgbxrVAlKbOcKzjwKUUJkyPAVC7ynhcouip8YrvViFFMolZGD5dYcIEF
IsyODojorPTvsvnwqSmyunErQWuNjrlRFaRpUrfuho3H6q592PyTOC4EL9IpLKswLBTs3rgNZwUP
PIZPAcqEMgOo2WYf9j/oKfaj+HToBmy309MsO2ERzYtON1HAaccGDrc4Pg4zcrbv/mP60OKSOgcr
Fk+a+vgPm/M4dj0Q2MCYdCwosTkezRNaaCbf1gk+guInzSUUlSulcRDMo4Ih6MK+yn3wLM+FOeMv
Tjb2wGiou0dK6OStQv56+xzvxD1kjPRsJE7gSWx1IH7Oow/3LHoW47ptzTpzY1IlY5kCzKveG3vH
oz+XOGPsENpddHSQp2cEEe0UlATQbEpmRuqkU3SNa22UKKl9ZdYPWvHHg5OTQoVkEQPFhqtIufms
3ufZ70ufwIEBIBiOK+1fzJrPhBw2dJHPjz8V4haL7STdQU59oNJmQyF6S9dnAT7XMDKiNU+7gIOn
fsVxi7FR9vrbCINEjECsaOdcD1i2hIcl+Vg5ewTiRXHp6kr05A2iHN7RD/P3PIKqObUWfFgrJs7s
syLgziljDXxR5xJQjvd3f4wJ/JhVkCPCbRxz1Et39xKQ6Ub0YVbQUpCsGXoewZs161B17spEcnNI
U/JCgdDPctbpqP2RTJaooFK2IUszPON5bR8BsMIvb6SSRvfVj/NJwSayYI03uLemrWDzF8T8G7FN
ms6vjRveMEsQHQG3SaRKgJwg4ENNlRKqFx6ZYJIlcwMQDgLegO8rks8901W3BL5H+JhE/zZcbZSj
eUWZJ+eCSvc4KJGF32F45nnCH1dE9u1S2F+qHV/WPk1ic7pk6um76R8xiFsr4cztMAbNCbp+3T1D
buiyso6Ks/oVmkHSwvYmuGH4gGRBafbdAEj5IF252Q95n2xwGldgHHnU5VxEwgCIFjhKIW1fpfn2
JADiRIbuX+MDNJaDDl8m+msID4ZziDTlN9jQ/GZyh+HxHZ1o919CBjDKcEXvneLLzs40/mBgSahL
BoKTvvNOhWcnxiFFtWjnqfrI5sjMPuW4GL3Zd6kj7SAJ6xjMJF8iq/Isn1llD6Sfl2Rs6OHWbUib
JMAjw82maI1ARJKyba0jEkt8DTW/XcGG4jqsOVYI5N1m5P9TcyDPo3AV8qEfwX7IkHaWk1DC4vns
OkTydNRuxYCb/9qvqCnXgfVM4l22QjJoax0AGJ/GD2+jLqPBc7mskzRDaRba3JpVTKVMTyt373vp
sbboJLQcbhwrMayy/12MIxhiEjV+6S6GIwlm+xqE+wgilxGPTiIuZRPEem3TYm/IqCymm/z2DwpJ
8ULUckcSu8AyZglDdFZD1eyrW7xuEGMd2lGYU4a1IZoVAwKPAA4iV9DMqCHahJ2GG+UXu7cJyzdi
qmG5KhHJj7Vf1pn1pE3QFv31LpzfcDMhdlIhNYXsQr/I++Xv6AQ77VeVeIVBiQ8C3Czun+JtI2tQ
60GC2yqGXDw6VNVpTiF8n49GN5tVH6K2b1cRvDsreTR3c/7ZpagQMm9YcfRoU1d0Q8OryzPIsLQ6
jzLao/OsdtTLVR2284TiAk8I5RDeleoGJiFperKy5iS8WWZewINd+EMWh45wb36jk4LWx3LZoEy0
izfbyjg3xget7DHD42OYjPbwuq1/TYacWUsxwc6yMiy4RE+53figgTTdCEdnGjC+9LAVF2w8Y9+J
mtZQuh+I81QOsyVx1VuHmFapZEJk6vT4avJd5BKrnyhJK7POL2pz3RlVtJuAoTybL1z2YSvhjNSK
D+EYu0HFRHxfOYwIN62CpioPd5oy9Q1VArAaPykH4DWHW4jsRr7W8DFtkt1sx4Gcqumt05BEYMbm
rvTKMIwCpcQVKfWaqmwFVKnRm5dM30WgMZse+m9EHPB9vrzWrrb9SygeMcHmzfpLTOxDxi+QRlgs
L2FTNWra3qk7QQe6R8qS3Pp3raEPQKUHJBkGm98IsaZous6ScZ83vgMgqfVGRBYuGsKRxakICO6R
O4q1oeK1+/MKXPa4lKSNugiMHZYIRKJYApJQj4KpNcW6cU3LEZWt24/Gbp9ExI4hxd05MFTC1n0D
eaqT0gli2lN5qAzJGQz5oclIn723y9TLQHMUCMefsbdxUqjMLtssbsPAo6sv1Q+z+WoxnQcJQi+t
uMi+pXlq/h6SAddkQCoeyVMrko0Ndv6uK04PwJ0Dugzzv754HVWMLGxX9xKt4GjYwnQ61JuLQgCC
niUd9zZZuh9mG0XwQFd+vS/kNGQxIjyLcSmEM/03r5RzBcIEanIiT6lvWNWt8KzFUmGGOHuXm1h5
D2JMGKkfulDmZwOa0r0WXXiVyfT5/qJIpbhBsrI2HVzm+t9Df80CUeGQZy0A3L6w3qfphAatqim8
0A8eUoM0QxIU47/4ww2d8b7QRs1eX+hVCEFqKCf3jFNJj8TyHf28mOdCbveYdc+BH5pryK4zrmyr
mLYTz7MWan8IBuyE/olimM1nmZdOs4dKc+hu5pM33EMvwgYC4Yz//LtCoVQrxibdgblOydWqaEkI
m7Wzk8yGKQ9kvsUykyoqekMH2FczbRpRk5xZ9co9LQOZ2KNRX2iv8o18IGpz4AUM6DQHuL4rTkwx
b114Q38GQLt0xUxfOD6zlAP9pBL7kxfUggaohNbM7uDTqlLNzthYlMZ+643AoMjONmnV/RMgPx1z
+ay8NLMcpelENAgcIpGTzWf5N8YVhZU5Gk2mxwrkX4AalywBCXKRToRydMfjH5ZJXTsG2gSHHqjk
liyS6WLxZwEyFg4OdGa8oPd1jIUKZqVsMp/QfVFcOjJgh66F7ks+nRNNaRA95TqvFSuEo4K6hRKs
J9jWGoskwpSYjUzUhkSwqTql97DpKMVDuSj7hKul2jxXPJ/Uz2p1uOYtAxNyJQ/0XTOSKBDkq9lY
q0OD3uQfsu+3VJ6o+xTAQwPQt53jmUqDtgNV7kXFyucf1JkpWIsa8k4ojLkSIwIg03B/ExbiT57R
MVeKvFandE0MVi+Cbrov7I/quG26v9Dkv9ZVq0WIgaoRRWZle469jneAFvA43BFPMtl+JGzRCmwR
4e3wvmQD7NxrK0BUAoSvpcmnK2Y5bVSTBOcd3pl8pALXJT15qHeGBDVckckgpVNH3z5I5ZqTCaaa
QYt39RMSeGrbeY6LA3nRfabp0zxzx/KathMdLE+Lo1NMzcesoot4cEwnyn54h6HVGsq6ZUFLFQJg
phSJ9O6FoJP68afDwBEPepP9kZV5Mr7XP1DjDEVsfcww1ULs6vJ1UAUhgMY2oLmb42qsedR63HIA
VWvzSK+zYVgu+AX9E5hduTMCkHH44jmhRng+Wrwq8hT3T/w4LNlDUpWbONmM3GbzrEYKUsMFVPrL
oCLkvdzrfcJWmhXN1oGx+Xc7fFUYpLjsTXdB9Y7DUVsLCKCJbDXNR7cPC3nkpNVSmp7iNxED5VR4
VmGLgZGNBFY8cLdtIGWMZN/rp4kpVmV17Hx7oMGbZSYcd48b36J1rbc/NrplmLZHC2L2AxDuaLHl
KWNGRdKaI/Jwf0JGLPo4vBpY//C6h77DPGGO9oX6lyZOH013dBlcS+dVK8bjqIBb3IWOnVx78ofb
0u16AV3FkkA2Jwo6HK0wBsLeu6TFIHdfJuRtEMZH5ja2v4pojTjDIMDXJ4B0jJP72ZlsjWZAoaLY
RIWCm3N6y17tw/lrxVN7qHNHBtmu7o9jZbBcX4W/K9PE/xkYoQWJ9aX+3VGztB8i4BJMx2t4Ikgm
Npf0myyRdjCqp6Tj+H+ulwKNwdFOTRuALX3BVgljRbOkT/lGXABpKb5kIOg+oenGKQmUFCP72aVg
q+1q2d52rnqpCA0CeorJKaTFRUTGrP80T9UXVYbDGNqC1CZWrkoogG3xJsAvbafyX2HNq7yt3oWo
t+jAcybqJjjP0vtKjZZVgLgWk/De29b+p3SgjnNEY40S+RXFUlk9mE08JzWhZfnvSwpyLPIISZAT
3KwQDnAmvfELiU1ETkFGyX1lpgnlzEUAVv31nDUFyrTu5wJ//YsT1lGKXgJUGjdwnO5wJWK7xPyt
U/6Us/Xin9ylVUcyZxoIS9sThpemL/OGFQoaUO8xfoShkvBLpT3Nm1ZzJn4wvPL1Ml6cwnZABaQQ
6Uf2WMU3TS3M+coIof3bfjg2iVsnw2GgXNVnSHXYkn9tQBMZ0PPmk3wMTxqcJbr3p+DYGQTI4uzU
eDyaBQtXCWuu4MTbofNNVLijhE6XT58qLCtQkRhcH9gtWA7jz4xKwqTkxmXlj++OVNThexIVmHZu
iV0bzPaxsBf0qDHV6kifeEG5qJG1ZCO1JTJWd5mLHqQ9MOvxJrYOxs8v6P/Uu+9jNhWdEOpq/ewv
DJTMIKvYhXTyCN2QPytOHZlCWnhbwfm8yps4Ix8A96BvYlEs7rkZ4Sv6RK8ImOFjMHz49a8X3ff7
92tRcta8WQeaDFMUxAUOAH/S1rBlr3FsSjLfVIDzwZ5lfMR0+QxapsVayn464fSQ/mMWs+NGuTmB
NMAt5xxrXcrJA0abaWv/LrRXr18HBC2sEEsiYziF6dxDNNOVWCtDdmlyqRqiym49r/mD4o6OjLkh
gNvLEkleqIupLv/nN+oX1IqzrRnNQBs1PV6kmHZ5rnhWmD+Wm6kmcxQoyvc3IV2GQr2C2RFypQBd
HQo2thZrAYwp68q7tCSnmW8qm4ZN2tyQ0vGyBaePNErfQZX7qKq/UrJ6fqPgWI0lJTrQVc/D3qJG
vQLzoYcqjgbMKearEMtvLoRYYUf3Xj6x1KxdS26PEDkvovTu2GKbYeywhwybnZfC9KYzuMT7u/8U
dKmD2i+qJUIVf7p21qR8DVwJW/gpcxae0xSziUu+ozO8FV7kUrxg4K9Y8S2m//ek14V4+dhgg4/S
84wB0ao6eg60GgNdscAQLJs2Srw8SK1Eo7XHRn6z5JRumhc1OrcIfGIjM3sD0ELcgXOXwWLTg47L
0tqJOKpUZNscex1tocZhUPZ7189NrVaQ4hRmJ9SZKh7nP9nyC7HBTKqELUHnMDBqzq7uz56PQ2IB
6h8gnvvyu5xSZ8Tdm7Englt+DIcvkZHRxNuGLauNKhq8364VOk4yhnmnTla99krrQg4Z6V+z38XX
AXoYuSO7zN7P9SoCYipLXF6brwuELbZLTvo4mc+Rqv3io+1YEi6nNOVscPsUnJ/iUWC8GLMoVPHc
DFyXnDHxBS1ohk8GX3qZf46YbPOzhIVP7Fb+2iuOwUMYG45dVnPI7lZmcIFj4XE5Vawys8duOFjc
R12h9CY8td7Or3mDu2Uk8uZzHHawKQus06ZGJ/g8+T2d52nu6t5dOnIdHhWXn1u2CQ7CuPwWgtSU
73m9MNme/QW5102MwN2mzE/pnRqXRxFzhNfkRmmZWkItTK7uFJba3qhNf+3hjDPYDEZhi537zQzg
KdCGel6kUgSTOcdbqDHTidJPOcUetCvv77/KdTgQP7Z88uFBsfIoTioI8uWURrV0/U3Lwk+tKigc
MFsp/4jdwTEz9TQm+w2/7RxsbjFrR8NNbMrgTykqECHcZZ4PCebZztP/DqnY9HxLTI6wGZTrScOT
Z3OGJhS3lM1wQ94fr5J5sD5R4iG9FgLYu59+Rz7Q/hfwxhGT+tIaDlSprpysfJ8JBpr0atXxwFP/
49bbMSrmBPJwKG1axaBixHIxeJK3YWsjFrCnQQeZ5D61jk5Hboo7jzYOSZgsoGAa0jMsAbEKaxD6
m/fA1u0dWS4ofJD5qEEqLhBmdrLGxXWSOofvpEEkwnoWI265jAA8efNsYkEHwHNO/Ot3DjRJ2oZt
ONLoojSDl7qp0VxLN64UP2Ba40BQ9gTTkeG/zpjQQMdGKvYgzEWhd+61SUY9DXx52U5+2n+T+OyE
RXrYjBQ3aNaU8smQmU2rBbdxQ7koJ3ilw/RWyewTHfg6WqT4Q1dZchJVAGtL924v1DL2HGAW5EGo
eY2bdJwwjbXuL/8MdfVIDbL/707K3MR9Lup7OAKVYLrbp3oLotSlM9jachnbnh/CA0m8waTzmfdA
2sFt+2yAcYQsVEwe1jVvyQiinZc0upmlmAC4SNq9Oo3abPGpQS+N2SSXrl+cFS88DxXWB990vvm8
vINqxxo6QLCnnat778gODKsKWbkHbUqHK4HlnavkKEdAfYFO03erT4pTdvZycia4UYkcYs+vmjv6
5NIy/yg2LpdyrWYME86ph06yAxbJiVwFyXOyt7sD3F6XdYIOfFk/g/VsHEh/doj4wj3EO1WmKOyY
+IA7gAbf7I+3vPBrsfx5d9VzCpc78tHkHqXn9SUGXfc1vMs9spXFBhs7pPaSgQ00flRqC86nN3cy
DqvlFi0btxEEasZfVgd+t8P3pFLQ+9o1hfxc5CjtYI90INSSapTERnvuYj9/gRyNZiTtAZW10Poa
y1S7PJuotdyU3giIQihMZ/lZsYdYCpuPJ3gRcZrb64EKEV80dJEJRBF/cQ/rLIMFa7ujfQKhjWjM
hxZMacRDcTGKe2sPyPEvTLyqq7n1947Z4bSOGirpKcHIBfabGSk2wHlPzvl6Ed9AdRMwhp3fRDFJ
5qbIxMg/bLNtpQmNtmxC1YRBMb8rcNEnymbeAW/ja4G2rtwx/XNqxeEztvNO21VLRwzDHpflwUcm
3muubUjW6hMtiMLktt/X/aEnWjldzsE0d+xcHAFYtZmD6t5zXsx3xsEEGLseeEOBbltJdu5ff7Bj
OVVIfmPIw1k1XwMyV9fjDPxrFUcttIbVfkKkL5iN2TdItG4xChGyT1zMWiB8jIbbpHrza/rqVKym
TRPbq+4xmX865TalV2DyR3ZNPh+tS1Hg/Q6D3ymL18lwq8yuOIhe9FN5plI5uoiXwBDA5bDJ4xPQ
uCAd8z3yWRELLoyj0O/SJoggbu9wtMYQwPbYxBZQrozNQEP/JIE66LuOu1cPJe371jX5znVLoFt6
f8LLHH0vAACnW8VxUB+tmzx/LHUdlDjoYqpBTSpLJwhNJHxGEaZ+zSRaTAnYBGrCag6L3oRIxfMh
tqEGauVRBk4TPGf23lnAOp6QvlHEA0CYu1OwD5tUh06gmz/dbL9MEjuGn8GNkDel3OWRH6e0HSGt
g7jrlPuhd7TypQKf+mzZtIdE2OFDdM2bnBPsSweYF6sXN2Ej7p2rGzxp5MNoIIiXUYgHBfE7Ev1u
5gbtqeH2MvmqhiXFbsOqsKoYbbCjpxwpfdFMgYnBC8K8uyC9oHQp4BfrzoHsulmXAO80EnLz29TQ
FseSoTxIxxoSSGFG1whcI1Gqp4ALyWmG/nbohAkANW9N8NSYmYw+PL1hWeOTpjjr6q9J7CE6VHIs
Ct99E7ZK0xW3slXEfIenaVounayA5OTUliZ+cDpVyuZKWOnutlWZwUooiWy3mCyuWSfoACy+YcSv
fQ2kK5Sz3p7zXoeWRrFMvlAUV8ZC3Zp36fbiqh8kSHmZTShCM4U70W8ZpCdgENwu4cXT3fEurghH
JeDWVjxwEtzyyDwDCEAaOoma2Onqb0wZnV37gNUhoiwNrvZWqyQO3pQZS2vc7XNrOl5OggH/zGyL
4TdXP9vuhR76S+/H6hYLj7VzdXOL0vb8lHzWZMY3IpGI20gqoZgt+3EtEDYiv8vTn7up3Jx/JVbp
19JBRMPpC5hcKT7yBvmMCNPOWTiQ8KFNzSQFOVc1WflVgJzkZ4sY5ezRkAXOQa3Bo/bp76ReGPmJ
tmZiujOpleN1LNvx7VJrOLGG+FEhwCEyk8670NpxGNxXxKtkmWkLWjQsI7i57SAbStthvP9h1Qrf
N+OpGUpZdzfe7dYY0k5V1J/raODvYlZpNBQ9W6dWso2F3GM2dXcOHouHnvdbfVMTZXOmW1fyAcp5
xe+wGi8fibXEm+vT/ouzYpBu3o7o4agaaawXyMyIQSWM15t6kIIzYJjb9SsfYcLqH+sJ0QmJhMqW
58SXFX0DKTJRBQ65hSEBXlcVYJ46wFPzmkCvKyZNk+cIbldQFWdfXlrSxOg5ot5vVSW9Ew8vfGn1
XwHw6CAdokJTEya9hvalfPJy4PCZm2JZW1sC8FsaQoKq5u/pP7mkIijIYOP4C0xc6CUKfj0UnAUG
q5OXpIOpgCYmCg0nylaLML+so1q8NVwgKzQf8VVcv0e7hz8UvZGk50YiZGz0771quwciXiX8w+aR
tufexCJhH7SpzEax9GuVfftjmZLD3W9tw4YH0FcZUZiK81pgMUhikRwrZvufpjIaVvx+xVhA93+n
v+JzUsHO1W12wRwp/jHlVuJ2a0XZ/6LT+MHtBiUZ/yWVgsUpj9r5m9fFx3AWlQtmr/QanZIlc0zw
dGE4174hL+ONsDrp6sMu4k7/S9FtEApzyOYrFl61rEbQ7n4UfFCu9PRXJ042kFZqNGpu/RxyrAt9
XDnnx7Ym9hAZF4lkVXPZRTL7LUVodhs2mv9dDx5TFxCkHqNV8gcL5MmKY34/cJeEcXRbZZ6Je9Jm
sfQZsT63jLU1F9pKZTf3868FoZtBbihLGPlvYW3iXYDTJpo5McKF5jPebgLQKYbh2LtbGZgq2Qog
eNi6aHafRp+i0wiKDpCTNo+rhksylUAbt//8r7bztCJg5hx+xEMTNsRCVMOIukiujLWlN6k3PKFp
61cIHbb5Gb/j9IzGeuJ6d4AF9yL9lMdzZ4GJuLWVvUTQdmnsPSQg0tWPH/AyC1EEVoza13vSFoyX
vdNjZziesOsJXDu0v6ynwaLNqljWVS2SE13FfrVD4GX9OYadybMyyOhEbrrNkfKnk25cpIYe9TR5
lFPq1eBK9igQ5TuBECKQqDQ2JUBKdXeWXCvUc0hAYbYQz/6LhYkINLNhlJJO+ddk7qrZHXi+rIiU
SF0wGNrNmaSk3Sw3XIjbFMAQZLmro/403y5slo3+w4jL7bTlErShsYDoeDukluCMLB33CUXKBGR6
C9Kq1lPcLzQplvQMfa/qYkMfXk3hT4bua+wiexRFjfWwfrxY/Xg6qahzFIE/LIPqPiyiY77AhlF1
19OSrUp5Msc0UCpA3oBljWYM0qXiGIzjsIxHQ2bVVE9xxTAHwUw/q2lePYmfJ5P+60WXvtnDfWW2
0r5u00DTQkg8LORiBc1BfR2antrMVJmoOo6bWKWBpCywNr7LgDupoQgF78uukDwqi4wZdU9PMySi
018rDYkaN2uSTByutN/uD4pnfblsmTwYARhnUeFZ5q4sywv0OJ6qtW1QzpzK2GBciG3oIILijaI2
twH11fNS4c8SiA3/2Dnax6KAkJioRzDnlBznEmzZNN4JhpCa7QrqKYhjpg9PQUrOtloYi33J9SkX
MxelZkX/aSdb6dljQQ61i7n4cO892yoE8PMTsQ9zzvQerqGcqUNZfJ1VIsZzYPJ6fnkC6HTT0fyw
kf7XcK0WYWhYgwdIbPXs3g2aqcMrMVTdcpq+SJplNXqvYXUdrOJmHs8Q+HGwFbXP6HC6ZJPD6kRo
JnxAw/yrUq7DWpsHM1ae5uWJzKe1Wuq6j47BIA8/XW9n9TXAPrm/54xyvrplIOxdHzQv3oioCM8T
b5JHpAmjqr+yUL40fmrPc7zP0WEDZ0CT+GcEO763qK+rl22pKGfSbsw5vM0r1OgkPOdwCWzowFD2
ajDO+xKIkOtOL4SCiew6gg1AiqCquX7kz0YoqavGCKx2Hq6dhvk0K9zbKVPXnPsAsS09B3aIJKgf
6KpWMhz9wYQgllTjaByHl7vd/bAKLuqAm3kBMrsAEla5E3tZV5Ijze50/pLTqVnQHvjaZ528EjX/
oUJd/VmWKaTpD5NHrqIhVbDpBTLIMGqO0YCemWD/ks1MCeW3sDN2GrRR2XijgpWfe4JENrCbb1/N
nCKMre7OqgwuQS6+qXdPvzWWpKlKyWTJTIDNszTvj3JoO3i+kAMB7yVXpD0fRa1HrcaSCV8AZAfx
qamZZcRLMQPNViFjeWoOwbezARMQ4duKgHLJMssJTmwbJOKvJggwJE4G4BZImIBy3ItGiPNORNem
rW3T4tkH3ttSXe1GH43vFMQEpUZp+OLsKysbNVzPV019iPA4MQ8jl7W48WsURgEmqDzs8SZ0VOGq
707m2E4C+PmxpP9hX/6QI7gabk3Vr5yp6ZNs7ZHfwfxIAzJ6tEamQSugpBxxvfwnFAD67HAwicUZ
qvFxVNtYqMeGKGa+d1kkBg50zwQjYyw0s1yyLV7XmgAYy5rg3HF16HNc5882UsWoX5jJEhbb9n63
I9nd+RjHCu8mbE8rMkMV2aF/qpHzldXP4C9BsF5/ZI3CgapBl00/aiv4+kxyZxlXgAEkJMvedAQ8
riSm4EY1fziuscdwvjV13BEkJevxHRepRNeLGnf9u6jxRgnAxBCbo8QIr83X7yDuTM1bD0LIMVYl
tt+JshwOpdHAAcPmNkHiY0QURw1a11NmksWsGrCSXdiGM75sTVs6uMTTbcAExtuNstnvdmaQMoDi
8cv5R7LPMjyrj138H88enpXyIQu8m8yDc5JelI8/Uq2kREucd9EUslm3bbLbsIx771RD1FsQ+U6O
RGZafic54Z/zzvPxK2qB0Jp3xMTW76Qe6bObdObwyruHaRXWoFrWVpkZv61hNZz4JiO1+HykMU3S
xtOTqUmhpCT6bNzNL+1HxobCwU2WBOolj+UAZhQvUbS2UHi7R1dhEWj3bZpR1UT08yeF1d+5QZLS
JYibWgITDZPenLNQ73TrmKFERjTkQ5p2BjjcJLv4WCMswcXEGqop9JIgq8cCPvrrsHpcFI3I/UqE
FOXsBJ4aMfKgI+gYMcB70WCFHeWDUeWB09pxs26oXQrK7RXluYdTEwuWOoSaHnIGFWNZ/nCKDVDO
Z0bZC04epb/EP2DvLuzPrxWRp6sRDIYWWOvQjitJjg4R+QWxwymQgruNft9Xd3T8wYPmk7l4hyGC
HciC32j5fzvQwt5Uj2vfPxUEDnunUM5yWystOPMpSB+zi3YvKgcbvmm3ov2RibdyU9W1+3Bj82bB
9390YoBusl1xiJY3KDaaH8Vl8nXJwq4mn2Rred7n2106ZPgm38JGP/LYKsnIKlOq6QWtDLXAmqfj
/KKqIYWycuLpy0srJrv0Yzh3OKfZqk7p27IvIXNdvGiPppzrCmb7++7g+1RH2TEvPPRrHfcZTh3L
G3hroG7LNEFaBpAkqjsMl/V9oh5p6HCP2knk8bvF1fSwOK1SxapwEAh6j59xGJlCTXllp3arIxu6
30eOwiDwDT9MsrpUou0WkFeHXXH5QIZSOu+VdtXrlSlu5s45E/bCST6Nvr+1XXZFWDaUn/lxfgdH
ZclOHJt0TZeyxilRxy9OQtZnVsRecfogQuzLvZRR8h67E5ASUa091lA3o8gyF5B95EOjDugPFHw4
0LgkLePaPcbGvywjdLIJDN5zUWV21DuLXrENycS82UpwiXDX9YOS5R80dFs4PHAJJudnH2ayTknG
lh0Em/8/UilDVquTTWKbcfgM+EQk4ZBULVzSQWQjMFqeA5e9/DQVMeT5kqkOAW05T11r31Cxj9Yn
KK7ebmc+Lr2137nK4O4EjjO/yWUA4/pEHDnSDpNQOiuc92cbGMIv1cs4twVcqO3PMEdffIB9qhCa
6Lmd12nXLhU/EDrecGp8dQt3J3kl1KAmmBaCimPdoN43U/n3zBAtidtBg98qVZLXI23rkGb8sh9y
oVyCL5eip4CZQibaWqRPD9hCJzT7s8JeuIbj0tjvgNjufN9ujPTasMfKtlGEtv5xRyIVxvMbMPJa
UIkfyqkUaAW3vP8X9X25TnAxwpNodAwWkETi+d1XlfLRZM1C+HTV8sg5cchxWN4+jpHfkNxFiV5Q
uf49bNAGZR99P7O/IektkrfYPvKI1ADf8niim048lFAh/pm8ofTD9G0R60hhHhvn6SvM84pZyPhG
qrLPsi1kkScteADbpojM+ytJZcyx+KKIT/ZFK3KJokuJhfEX3+d4VPuQ5zeyJ/J5n69VnrQxGBkm
f3Z/S5uXIQyjJUqlBSgbhg4jeKZ09Ewq5CdKxykjls3GZ0FuGNMy2tPzHOFH4F3YMn2vUF+tf0Vu
CL5ZBrl6Zz3+uws9hVHyoujWVBrP9h/c9H2Q6V5zrCQKOB7R3+VuBnpz1rYaXl/QR63X7mpO8WL1
3x8BDxem57JDaR3nBHxVJYRyNPcZyB/4RdqMSUcwwPU3inDBru8NDSqbSB7LcY42Vm6/ACgrvDNL
7CgVczHu58gl9Cmz50YcBuD2stA7YL2xFyN4Enx+fsx+igYPJqNHwT3zALou0R5TpW8L+3FJA1fM
KjwR9om65Btge977mN72s+9GtHSu0RkOTZepezBQg/boJ0xndMBTi3LicMPfV6H3kApGB79FAmWk
7si/MEo6i8omDxoSG+jNAXaIFjlIbrlNamqSheDtL07kZWD7k1WD9JxJC1P9SRsodCz8HLsT+XJC
65a3XFyE/otPgJoXITBCAhyeqiNvkgE4hhfJzE1E4oNHhRo39ff3p5OF0h4uk0MFQ6eC/dFWssz2
BSM8k59ZFVhM3iIEcTAhAZYu6+gO5vlJqy/uDFdG4/K+m8tBA3iRJ/cKWcQYjB76pa6k9jlUyu6h
t7XdcIV5R15LAGG6zJFeQStnjutfhDboNBycnVTv1r5R2spSC2J6AjM+mhT0BEGXiyYD847wb4Fn
bXp0J5+in98DujvQ1wl7dwEj//S/g1juixzxHZ66byewW8lvLJIe0sIKT00VugRzmxfPfWtRF1G8
CEOF1Y6Nz2mOIfaZWGotdvd60TXIosQ8EHqBfhZqOE6YHUO+OhMfaKnSqnrWJzh/uFswWjvAeKxl
tXNe8lVp8z38GW3zlhtwKMj7ROl97wAW8lo+DtiT8bfVijHSKBMXegKMNri1GU/Q9sywszi65qUe
fhzZP9xvGerMB8C/K2TpiYcZcfDXSngGiQkN7c6hkLQprno09NQ52V3Oiv/EpgXtn4uyrNieghIl
FRX5c4zlB4VGBBtniGlo7b0/dKYsDi4ryxz8cj4phcX2ijolcd6C2nVxGxvXEOFufK5fwgaIDwGX
bIqdiabBFXhoBpuG45MFkOwZVhbPN8CHXF0W6Ix5xAFnFg5I9EQ58B3+j37MU9EpTxjFS0C3P1d3
WulR0w+cuAUV08bau/iHQrLBvUB0DZQpxYYR8kzGdT/76f0pYC8EOBPEf122YAr9IUeUHJCb9i1G
M2AIvhQuoAPdSRVgMb9YtNMbDuYSd96Vp7MBC0AcC58ENT9fdUtMj23YTHo9Br5X5cDHDPWy5ND0
7+z4Mq9GQUocJ86LZPwpbi27uBcW22L3zSiAeVIHjhLdlbY6yM4BekFGDr70vj2rEY9jmDDPHKvh
8N3KYmIO5HMY44/FnOb+RZ3zF32ike8nePv4EvLBaMe5Isjro7PDOZjKtDq/lXbSMqHzA7BzYOdj
pNh+m7Vg9M+NbyydPQLDk8Jgj2ZmxWpK7g4XjlP+EpAiF7/6il2Xn96UhK7lP85epkqQsrfs8AvC
aLG5BRLnKPmHy75+HF1YDcR/GPrwZIzW8V10hhJfmMpgD2ralHA7nJwngdGA7+Xytpq0pd9rmPgm
4vlc4Ws6z5Iac8quRukwJ4Sqxxj75fIenRDA93GXoK0MTIKyrVLvEDPRro82ppG6ncY5gyr/IGlI
+CCvMkTjx9nvkWd7XeWMpR7QD+mOWN8dz091oMjNyUG6xrZsVJCeLUllz1V0b9UYunrMTKOW40EL
zUfcsYXepvPF5HRl270dFb/8le4o4z2dWqtuxffkW2o2ypQfBJghmBMsmHvINwQHEIVnwujx2USU
G3uXoNgaY0KG8KE8GjZd+ROZDQkDRlQ9HZUGgNdyWJxcB1hy5V7rmJn2DeBlnqDBxWL51uIwt2V5
x35T6RkuRb1ud/b/Xe6PaTreHpSx8Mij3LgX0DrMtdBuBEZjU1UdLhaanTHcVsU2Y02hxb12u2jn
HBFrqdMQ8EAr5AiAdJbJL5DecLXodJyFBkva6SEpcd0qWMN2wUM+gB5NvFxLoExatvINEopWLqAp
AuHPRoLt2Q/AgYqBFNFzozFgy2XtouPa+1ndjagnuD9012RllZ9nLivq55DaB/kWit4qTPpu3PYi
Cv2bi1+j+FbAT54wEKilpBuj9uChR7/LU5xLQcT3WiEEuhXwjbZ2sTs3vV4/mqaQ2yjVUdo4fKMm
tFd/J1owQ1NMExR4Z/cH5Eb2fFNp8sxvL2kVR29MW9s14ERLHkB7UR+fMHpVRQzdwrK5kmW120mC
6PMLrJeaGgf71W9u0l0ycf+izisV2+JSutpGTUwlwHCcLalkdI1mnREu4BpTQzEsOPj+gXOafDzz
YskkHqqPMZFvB7F3K6ePIQ3iRb+33d2nhFD9w2/kFTzr6bAJSN/ivh41fBoc0ej8PhqsgcT1Rb9q
MiG1m/w0skc72pIwRPuXRc2RR+es/HkCsoZP55Hqymv1raObU3IYOqgq0KZ2oLJ+B7+fhQyGGblS
oeQnHBGcJkcKtYN04I75XHqdNxQuaKszAUYH9lg6z848yGj573EoFAKba2Mph2jRmQ3PEX6FhduT
5kYOPsJTRk/UttxzYIEnXl4MwONseWRSo/g4pE88xVo/EBlB6O9sqaXh897VDMXg4Tmf0pcgabu0
YHQ/hPyvEeNU67wsK/dq8E0YnOtV1TGiBIFEYYTn0EcjwzG+On4NGWqseEVjRDlBCacVJtj5lkro
zg9SIgOrahxLzVSHiC4H6pTdkhv4qvS7aLb/Wwe1Ug6YLJ/gyMklyoGiPsfxyGEc4EdWr+WRI4hc
LE8dFTJDNGpgFJc2f2Q+9H/g+b6xru2S/NT1zikzOFTHwxmNQw5BpiS5lEtZmmL9+47zqjv5spUi
bKXVjZcE+ynT16jLRsmS7t2lkYLkV/GrCpdlTZa7L6RZ93i4mtaRO++LKlZdSeBcmFKwzdKyZ44b
2+czYwYyUI/+LIbVZaouCqPKF3Eu87eAAVNOGd5mFUOuBthp8o9B7nuMBWeXQrGnJhxADAjWwbGL
9rXP50GSiMUHYubZAnVaOCCuTqCTCr2EBpsfyjFi1VFFojE6swiKDkcgRWMX631cqYtPILaAEF7Y
MDNfDoX8yjuRAxU+Z/P8jGEB6YENiosK2DxpZWvxufRacabTsnYaZqLKtVE0MbPbc8crCv+UdvIW
fY1+Zkc1UwiYOv4P+VCwRzS+FQqtx0gszybr+5Qb6joBgFSk+tFALK4rdNyIOv6ockwbxqgEtFnB
yzXxveM0uvWDgsPxec9P6HAXF2yb8RAL/JdC6oSygU7K9EtTFt3RHdw6/LfAoIo641dC2oW5cZPQ
ZIeCfhOSJ2i0sFcVLqp7Q5bG15f0SSc4mRPrYb+4kppd+C9/kiRrs35oo2XfMlQNZ9Ihu/9/Nrnj
C7F8phLJk5GGOhk3r7ww8jBNR6BYJ1XWv8OywkNz6WrlvysasvYyymTJ31dy4JMAMcWFlRGMuhF4
77v7q3b5uaI2pz4MqDukfCKin2ecYWkH3AjPlTXeNPSmfOV88/7O6Y9MR08ufmBvtbOKzUE58jwX
hyQsYyzHrMRyVGT14O+ovM/lkot8JIG1+feYBK79/uDI5oyum6G95mWuO3LqgnPoNGDwpJ2t6wq9
JqQiqnN1U/4XQdEYqmgc7ZSiYclvWF4PwBC9PaHo2MJMZorSBkU2vK2/uWiBk0cTeEWkJMcnwfnP
aPMGvGFGKC/eOHkMb93jVjAfEA7+C8oa50nN47cfEOd8M+9wV+F41rnKyzPFQl65TylaJ2rnAekR
kPuccvbOhpDvGahwchmgIH+MEJdrvh0VRvq2+xCTRIRszsyGq8zh7rQvUSBPvG78A6WUBlLKyg9w
hnedTdLvVRNUZCXNSxVB5aedlEJswA1BJV/7cN/y9oieGSM1jMIpiOzCgiCuIT3fKwU9K4lduHMb
u8WDOv5N/boBIQpp3NOhbMgzXeVjNN0pZg6jd73VqVKGKVfzllDmgaQpAWUe5Am5TERFswFLtt80
/HWfyYB30pWn9/tAiYSKrCxazg2i4qVJOjnVadbwuZAHZdIwVDeCWkBX2C4xZ93b1OItkSKirdqX
1ckBsjlq26tSHLll2WQq6Oic9IKRr6jknnjTuPt1jXvZ3IA/id2iXSRFw56SQdPSLj8MsBG4pnIP
mCZ0GRZN9rc/ahhn0qMuFRVY+UkOQcQlguPjrw26fSTcvtKWpf6LOlJBQ+qRJN7YcWNdRtjnk0r3
CM1DSPGsaS+lJ4B60AABCjMFj1HeZG3v+TKkf02Vad8xjzsQ5E6R2cN4VY76PgPww10ABCPmLX2W
n8UyUUlwAZUXH1muxSZjA3aSsof6gazgeADYaosAP/i63IlB3B1AdFD18Y3MV6JYEqOaVFut0ngg
porc2P6MsuYvY98zso/RAvXMUfY/m/KFmetnU+DgBWloZLSIoMIxiJ6yv7Zt+nE+snkHFBeyv7kv
zaIKymd/cMrx4lHAxa1XfU6y28+dJmeo6COqKCMZbf3NiMBBi6Zt6IvLYkdUMtuHDkmCwv6yWKTB
dEFDAbeOQgl7P4aOcQRul8beO92dSi0hBHJ4or8xRh6n17BZbV3VJ0nDfavv5X9y/MdpjTTtppnZ
c/9QzExmcrXHqsWdJyeNo6+/k6s1qVfzHPalHzUtiJY3QIduCwFxhv3t74NexI+TQuaXEFX+BDDx
DtYMstukAFZCzBoYHPv5xOtLub41XqOXfLi6Shqg+P3QlW0QKZigxSeOrAv0GENqxLz+k4a4A+Yr
19TsPj2r34pOWFOQDTQo6YcZn/lIS9paSmlVDkGhRdv6A0co25Io+J8KMpggo86nMenVwkxWzDep
IgyAVa0vQm2xt6EMcXHumNXxK8nP4oVzyT3huQ5/Kq1yuVU37dYtdT9HHk8Uvsy5ZHar22R49oYu
YAw0YwQLRt4ynFL6XphKufyn24MXZ3ZjamgjWQndhTNkzaODHWmVfG362NnSZ6sn/uGWjB/R3Hpl
bHrTn6NhFmO1xO5CymQwcXYb/zI7nArg2BdpN42J4A+XWmpQDda+MTGG2MJTfSVxP2VfSiNDeXj3
I+9xMUNzS1SPeDueTft5Gz1ES8LOJfvrg7FBluWX60OwB9dXhykKZeMB7XbNCZgc7RanYUOHL5gi
xnN5Ok0oZveKCZP5c77f69gbeWeFV77UFoCVh1jCVlXqdeI6zmaKod3pVEwOjIeRfoXkqmQVPVo5
uaY6/JDTZQdnP/nEwTLjLJcmxmnUi+rAz0lSKq1/U5u++GeTrt2tAROd7LYv3RDVuC+IyBEPzXZm
bAhOh+BItowLRkDQgEDrPpC/kRWVvQS3xZfBluYCDMSo0EM7Labgo3xzRqfqXrWaGz7PO+3QL3fe
8m25MCudBFwYN9g4Fc9BdSszUsfzDQYJ8EdvbbijxSS/TBygDQyrMFag8KeUm4qoPW/Y/sXTkXM8
Mb61yj9sXqsi4CTO6UfqPKYcnlEP6kCRFkoWjAXz+iPoSfvbmhQJZrQHgAMuAPqUaX0XcNxuPaG9
0NwT204p1jbFmWseBdeH65jrdjgZWXH4qWtggpeHVk24s46W9/ZtmVgOa7JQUxLHbIhE18zzQFUT
EDMXuxKZ0i+PJ4FVPLTDu7ekA4tczPM+9db3NezrBaHt0ua7uDfeCGBZ0MUTyP6WTS2ciHTuJmzK
WHW4vrzoC2p4ekKgPvhk4qc6aDRvKHaqcOZhAS8rTx4crNzrO6iULzaqoQPUXUe6KEA0MzJbbrl4
VUo791gSSDcTHs8f166cuLg7FKUk7kwF6dfybdxPuagt+Revpee5X57Pd269Jdc8zCtvGGTXVrAJ
Zz9yPQC8ZEjpED3e2sO78W7sP60PZyv48vRgGb/yWrv7Y3r6YS9GWLgXwffVKaimOtcESECj+UFI
62PvEyHv4wUvZPSqJc1zbGa7j0sf02F+zXI2pG6I5PWK/la+7LlhjU2I5x7WBaL8LTz9Ar9zqksb
R/Ze8rfIrMUF5d+2LqqKCjkXUc2Bviwb3zJjZzxYdEcAf5FqTCqB1LhxKmHnMHDWPhhUgJWJfuXd
ZYbXLNdqcrv5RGQ0PhSyLxoR6yQBtiAEB7RZeY0F7ydEObEFvXQ+1iBSIn+D3OTNPD8RJheXKeCF
b7VniC/AK9myAfSVWINJS53KDwNxJgcrWvEFpwxsgn14Hz8fN/xdj0HU/Di45mJcDov9u8iIXYbm
e9H0h8tty5Kklukoy2YuP7A2UmS9Bj9hfQyn4+FqWrugrnOYfsBdzfIrh+o25GcjxaWayFsfRx6C
Dr51m7SwpEqU2lw3CzBgXnK6sPuCWo0jhv58riPt5eHnVuWXdOQx0YLsRX04dE7ZG74juN0ue42x
bHws6nOQNbWvBHIJLbtmCOUL8Z6IUuTroNgSlrPvkRwkQfZKyCngP0QeOIZNF3XP5dai0A9sbdyS
+4UhsnOnS1H42R8SV5rIoDtk0Oys4ztLC/TIGr0g1jw51uZ9WrUb4+scUKFO5fzAF6+0QCLumBa/
0A2grTpEwO66vxAr51tF0+nEfPm7fdzXy4pAGZNlspPPXCuhnKFbvRmk1CzTXnCzGPPmrKjbpayJ
8LnTaxNRS4sbu78i6xkJoEmxsmUC7F3fYMftD46SkO2fFaJa0r3ARwjU64H9MowuRia+TB+OPRy+
I4AvLQQ5THFypG+8kOwSxLMtUnPIoiM3PfKsaXAAK6qVTpLbDkC1S84LguRugLbtUNPXRAGjTqFT
xjSxkxX+6036Yt2/dSy3FD3amxCNediJQyeH4CyWp5i/XBuEtYef71EdWlb9ahgjOz4sT2BFgF/V
xItqZZfpE73YuA7SLS4sickUoirlBJxNW0L4M3T4qL7V3Td/hxTpBxCOCRq9L7scTr9gag0BVE1r
ohvRPeP0aAkND3J++1S8jbEcNQo9PHvxUsA5CiRSTJe3EPftoW/srBvSDKQjuRIW4d6+YBgCCBMN
7TadbXX1hn/fxtLVZkqlw2dTW0B86919DGUBHZaJcoJhCs7prtoWVGnnV5lPVLGO+Rp34wj2W/Fx
psMP38TUj/DL3OG6e0dknx3DfOW/rA/PdmyJ8XztFlPYWVV3c+LUQ0PWzo7ZeFyEVZNg2lisPLgZ
05gvg0+Xg+jERtt39cUv+Bxg8FHHAqCx2KRfr5AA/lpZy2J8481UyAUB/PuuBKM+8/M9nJfFqzpC
S5+VtgoCxdil1Q1cZ8A0g2p5ToQrsXtSZVOTOBtFANNeIogtTlK4xvM97kjh5xJ7hVQs7xYN8gKu
GEpJ89XgtjPfNwNOaOKpAZ2JAGgHOu+Xe+OHvHdLxJo3SqgevSqdavbFOUXFSq/O2vLrzlpqj0pn
ktUqkOqoTVeBV712zThPkYPaGdsPWneJaoNc3SsaTwiVmQGUyk8hDdHK7pUHUmvypKjtZ6Ma/VTP
XQDa+8no44+/N63p2roUkrD9ZNtI3hi8gcwktt8APZmQzhwalLUB/KFm5BT4Rc0CVZVVQFaDo3L6
8S7zRliBT7vJNY+uFIliiTiAkOfAG/Q4y58IoYcRxS3UXgNH6YTjBe3X5O06zp52Tv7M9cS+KlPe
SXb2IEu18UQ57H4Jjh/NGzNeyr2Ii6ATButg0jgSQ4LtFFlcqDXldMPPG++sYWUQbIvlgTywvUN4
Po+bON+j9q5Qj3By8mTf+9YgoGkBOlAivAz+CD3Kpsd6wyaJiC9W7D47a5aB/AY1YIh4EekfkTum
IxG7J0wdn9O8fggxJec++4+yJFNio2ga3oM6dlJ2Mz98LaZwFXYLfXKdaCcW4I/xe7uuFGbxjyxx
nKf2/fr6xOAADZARI29sPGZPZrEX//wV0vNGBTM5yF4ibgCOxZa7KALtiWwyLuHAnL4y0fMG22+3
W1twSI3P5HkySX/wdF5P2WjD+dA2/9gHAyFPYiQqagvjZteQulj7UzZkcKM+fEjbuUC4N0bgNDVU
h7a5guWBLWs8YMABi7uumf0D+FNoFDMTil3pMfuWYa3RqP3Y8KIsgHXC64QLbboPEtpyUqOixS5j
6uqrqcETJ7qhyROULXhJshUg/llLEJ84DtO5qeIkBsYW5a4hy7I5GjCMsM8Dpk+oSbYdxaGPqNBy
ctFvIv+LaDDq7H9pfp8AI1XGsTMNDCAzFc8DyMWAWdOfYKuV6U+QK3CPBXmMblUq8x0aN/MaPjj7
18yLgBEkF2J5kz4mKJO5829+BIEO6E6TFsKqk3D5JIgxHtCWkljkrf0Gzh5lIgFZIrI4ZQ3jdLdi
ZpNVrih7KAlkzv7sr/2pBJR3JKGM8sw3O5L2FOb8DSePKeT1Tl4EquMFyFe3cLB7TW/LjipC5kvA
cjssDoy4t57G85fQwA1xR0mTahYiviAnDRb+/jNnh928iLC9wohyPL/e3E0u1r6ZFQsIUlXApZx+
2OJvjn8tdfaBcC0WnrSQcZmz9QOiDvYdWjKD0mBvLLuPVnvgEKJ6u0gpdPLzWT/nhetLDFPIOazo
WGk9+/g54REeH37e1m6vmOiDojZzIDW966V0xFXpc2gmMma30NQ4Y0HFDd1J+WM6FpbnJD72tKaP
a3EMzoTv0T0sp3X8SyZs7PlwNWI4MC+9Ut67pWW3CLCBVHGQIqtEBmbIeUozWSyOmHA6l29JSfcP
jMJZ8iowuzNELGAaW0a8R+lA6/zf8MnP+pZ3ZrY/q1syYeSQtRThaYSZKSTg63w5EFIX0GtsdBWU
JCKUsvqIcPff6zqljcOq3YCS/9/C3rrj2VrsVU35MZGjdjlbdoRRx3uVQzIx0lCp+h6TqGiFRPnw
Woyi6s7eNwDFrCJcCsIfFd+cTshyYDsyTCli6OJmponwjbjw5PnOhRvRToOg3BMHykKRnU7IaPGD
zQ+3sdgcjxQ1QI/ZC4lemtQjde6WKKnaILVGI0cpqTY8fabCblohd62lofmsU5Za3/m6QQ+Bn6aX
slJnTu4n30PFimHZIlzfEPcoytnSjT3g1R+p/9VSp7OTSvaZ6d2IPC3Ge6pUrw/K1n3t9HatDzE3
UZcLBa0Wc1zfPzczvBfLJmWX6f2QaKYLbfOZpPTJvaW6vXj1hBCSrdPou2q6Q5OAiu/xk7kQD8xw
GwM/iw9LCc491qT7pvAPmQwCWS98hBCy3xusmwNO1YiFJ6DdMCZRAzcYziZwgIoI96G/jEF9DQEs
lvoJjrovPCQZotHDLujRLg5rbdDsOjVl8TIb3WYxWJ+1AgsJmJyzIwLtoMd+MD+P0hR3VXENG/07
9va/c8zr8kI2YMRwNarC8NFJa2X2u3R4GVhIuNxi6aIGJ6grFqkhjZDT8GJst0o9hQ6utIv8Gc9j
pacBrpbtTszzrFA+rjrLvfdZvhdeVyVBi/BuuFJVAKnc5a4+lw6lHwHjCo1wa+TeEX7iDt6F8Gq2
HL0Kp8Qas1GhDILRGYrbi4KgDKArgRW/b2XN0/TeINHO2tNzPVtVs/xL92fLP8VLLwIZ/IxGu2vy
oRdpYEHlPoJPdgDcGkdUVpwY73Gj54VOwB/qgepTwGBhVFoq8bhFC7ExHjyn7As2IkPlbjMwZWDa
QWMbX3uxaJhSIMMWYwV6xjCkdFCaSDk0pljrwmW7EGalPkD5hLvY3tXYkNH6eIMdX31aYVEi8f6N
bxIwTWZaBTHsR42Xavc1Y2guH3tfwFSMHU69di2yPytahIhZwdQPZmo83VdF/ewMPs4eVrtddZmt
0sdcx385Ho+l+D8mzKcJZvZzaMuBNom3zNovtXnDCbhX8gs6i4BkKLChEOaKcBHByY+8HCuuj7Y3
/kKSipRNcn8ii5Y9IZr3xx+lJYi+4vBc3T5dv+rRHvcNNnzZdSP5esdy31AK3b25lQ6kaY/kY4SD
NOQ4lpf5kfD7lS0+kBANd9F4b+gAGs5tcyht2VtHwe/NbA6S1PAeqBzJ6JhsFQFKApAYWAd3PgCe
dGIJoJmA1s01C45m+4arwBR3pMGGce/tHrqa3hgBRseIf9ht5LvFBuE84fLEHt7QyXniooRxuKPY
BessAO86XV5t5IRdPPkx1Bv6Ui8QpG1Rpi1Ra4b+4kfdZPKnKF1M8J0X3EpYWyqYNaqj6n9qged0
lwuIFPCaH/vIv2LW6qQ+hgLDf27VSfY+mAngOS6iUH7RjD5cialgayTyeawC5Oh/VkW40rNBTdcU
6yil2mjNKwAeX+DOKE5n+cgpzqhEJnxdy77qkPBgXVkx10k/Hn0mxjAG3+dQA1JPYRYGFXVxgCw7
Sel+TAUyL17FZvoGpA81swEZfFJzF1yUbGFBTGntLN0T/BNFoDpUst4ISu6SeecB+FC3WCqEirwM
sfn043G14FHx/1Kn8zkaDsrx7RMv179e2Lj50zwwhDHcjsbvU/yPWjFcJzH8pwy9ZiyQRhka70Tq
YzNbqy5RJ5T9RScmHDbYlmjHxDq/6GA2/34OsaBaaUuv+qz7KBRcqFkZLMSCW1WUsHvAhsH1gHuS
kFoYgSNibKyJoHmslkS8d0Yg/8y9nqyUNh/M36EL7i9zY5h76LfMOjhiIaZaJfsLfyauHus7VkGw
o2zaMxXmTRR+3N5UkDHyRO4E6SFpae5IylbTeDsLg/sR214+T+Ei9XcDnA2Y7bpA1viX9z5jazyx
qW8QOSzcGMtWA8uISfL6VAHc5fUKx+fB9J9j2qOX0ocNxhpsq88T7zYztLKW4YfDH9bSAWt8ht11
yugcENQXX8Tu3gRoJy2gU1casmGxP8qEwMzzUc97c0+S2iJhQj4aKlwjpnD/6muvVn4Dal2cL7/i
XKzAg79CwbWx2WSEuNfN/uNvxW5UcFTj8Ee0D6tU7USB28mSGijQ06e1vL/VsYjspvtinP6eQe9+
bxSCI78/B3/K0UViffda1icFO5xAokEmDta1eLF3HortXnbsU0MJFRfu6HPTDJY8cT81Vzmhy1V8
gOyCfNQs6lmhVxD/1NLu/Moee0rIeKrbQ/ofW0tmqeOR8snLPz34kYz+sRVt0WDdtQa/iNxaWLor
ghcyZPF/RSkNPCOYrrLlERHZA50ejwtRJzPmrBUsBaa9zmd0IbZLHmjV3G6cKF7vxanrNBqdmbXo
nNb6jcQuK7S7XV0u5CcV9oAp9pOwUOylnYAs+YlMV7+JjUK07+h/fyX59tDlqCZG/vXIlgOnR1dJ
AerKx+WvtN1v9bg+9iNlguuFXvX5L9X0nWjbklCwHmM3TTixXzvWRoHylyTM4GbvJJZe5QCn7Xvh
kzBjcXgP6kf+ObY1Oib1r+x11cnZ3hCTJlYBVxsLsL+jW7VZUh1TYzbXpnZ4wAHOpdYe6HSCdC4z
L2cOq9+8R4ukDuM7vRg0YB80csSTF6LLpuldJjyf8RBK5FUj66C+gIoXhRj+SsNhweb5grCGWTuV
luNL4s5JKmtzGeYcSM3r5xljIoq/DrtKFSWO4+8AAbBvx8r5G8Q/xALEZF+AFdjKW7iIiTo3J8k3
yaYBV/j9qh08L0HMPKw1lwbrwQU0K/VjUg/1KeWCZbg5rHFdd8qnm5kW63wNCSGKCc1H7FvO+Ivq
eNhGqAEnnD5yDFpxBvncaCB+iC88ItNI2//o/kZoSqQ8YokaxHAB0bq7E8FndjgthsNzBU3/uwSI
EoupXiexDcHG9YJgE+yO/fCkCF2l0Q9h4uK5XYzjul6Mj/fH5hiZe+BueiZJTaLISE1boI9y9Rku
EsVdipyBhIRPTRvcQ/zrf4j4B8+j7H64lXe5UHqTpWCceBPDcvK0e8bjreFEzwxl1obyJu2eT14T
OW03ArTPswJwvn65pHZg0AkBxzNzwLPSN9S30pwKyj4d4OeHzWDdSilNcZP99iLBg3Bo+/oZ86db
CZ5Qp9HjW6M0qKFxcrg0N1yeLSGUUn/zFziBApRfp2XZqFexqZtbtzlVizVcH8LnrW48HCv9/pj+
sgTk5d2VrVXXDDMxryLsW5UFkxMhQUpSHKZP8FKs/7y62FSo4JfTs8/U0tmBFfGcOp/sxnH1OWLF
QITQyQWNapp+jVsbgTFaJPEmkoIcRHbZH1GPVvPRTgx6ugn5BOTm9JZSXSTIW7/ugrggfizeUe73
KglYzJmV+8onfRXaXnKs/PASNa7hXQ/dPLreXdgVd27CgIKB0pKc5jiHGrCshHlRSzKcIZVrKAeG
UT7YkQvPMGp2dyAbtj7z2mu5IsY4aU6xqerjx2+QWz99aXGuNOFcKzgg7q8yXMxDS5L2s4Cb3icw
x8doyS31plqwqj7PuiK2+gk5zwx1ETxEqrb/kxZP9eErRcx94MOm8/PECH2US8DCBXGgV9r34DUV
ecjYw8Ra88cuMTqym46Oviifn7yGtiD3r/FYcGLocvGEt9IDvB5VPYg1KmYZqjnTrD0A5+z3JK84
E5Z0lfntmOnNm0mwLzUm4PdkUsW6RMpKIRtjkInxWKs3MjWfHDJMrPPrW9vRmSUI46CPeeGe27yZ
qWIBVh/ju+ofvSZ2XtQwgierefdC/BpY2l2kYlrB4QGUJfH7xaMJprfD/RxGviJtAUw5zqgXfNOI
76JoNJmgKDrVoJpOSDd78ZBB3O8ipa7dVSSz0mUzuAeKxO1sbiv7GX3kjuR1nn38W2VjdSDR8yUa
XheWc8wstSMkqYWc80VTJi80W2smcQ3eZN0DW6Bs081Y5V2hVG/tgOw1Fj6BYynHEs3Jh7HILqjN
YsKCv/51ha63WBLjgnwtl0hmn/sdRZeh1jrbjGqwUB79PUGJtElZkYoLxSWhJDBmgSNps/2b8V5G
AO/fSpVwzfdnWVBZRtyCbk8Wm5leQC63d00SWkf/3Eha7yhpGFvRayEwtNSPCb8BI9wuxHuiIe6P
UQCgsrArbzz2Tq/coVwB7rJhWFoGDp3T//btg/sSue6PRYm3vdVj4m4Ho8wCFJuuMugR0yESk57D
pte5YosL9Xv0EF9nGf1MZrL2GWYKuvNilNPnkr7uLT5kPA+iC27viFTxH7jh7ImaKK7Gz1l92N+m
UfWwF3YEEBoviff0fq+yFKVsFmDHRWf811xXw1tCKFqPPujH6lpPvyZrZjrso6CyrY11IzJX1QGA
+o8K5pOq++lh0Y0/olJ+0aibmnrxaYJkOtLUTBBUWQ67a/9drgXHu7pDLtK5QzKaslI47G+3tlri
6o3d1jLIa2Xg9KN2P0hSGISHwWXxOPppGu6x/DEBQyJagecbz+UOWl7l7boAlBKGLwB1BT8fpzD9
tcXds5wIm3OrYbv8L5yF5yisU+wX/xFlDHxomn0Oor6c5CDPDrO3n44vx7vPhJqq+xjEx2oBlRVf
jKieqdiFAIWq8fsI1olJ6Y9FseLsuNaNlSZqGnqn7PIFi9oQMA13n0RjpKUW0etGBD5+rbCvKdNs
IOrgu7hY4l9Zd3AU0hPkwjprerBs+lMs1kpZqu6qmoxOFKpiyxqwwFh/xWkzo8y7WEezFwIXhzRA
sIT5AzTyPx/5/UtndV6iIdxPItpN2VnjrOHH+K1QJT/f4Y9mXvwXKNvYLw70uXAKamS+Dha1TyC6
9SMNvRnhBoOto/WgAsyw2CljeIwo0XP9Fh4+Q8Ak82QwXsFwwBTgg2K/CcqqEiN6K79LZVcargNX
H17v5OoHFTheQvDxtPV6X5AgOsbw8wCOAIXTY+dQG4XhZ8yoBGRoEtu3vGYh5pTNqrhcvxdowdZd
4m/elheSxQhyUKtwWbUZtWaDho0nZDcJ1I3ajg5UGbKywVE/fY74ihtnCt6ov0xjzr+BdhKrbJz/
rQHfshploCYh5oZ5o5dioagl3ybXSFdGr+qVix0X6niS826rmmXY8mOYE9yDtaB0mRQ32AdNFYy+
Eu4xsTecDNEh9hgakvSFH0j4oqSoCw8LvP2irnDGZ+CzZHRmGa9fvSVtNdsYP9xDmngn3HVhJaFB
krm/G92QULAJPzSWnbC3SZ5GMMpYsi3uxab3PNmvDMGQm0RvalxxOj0BkDp/djlHqQwhmxwL6RxU
arZn2vAibAQh/L4dNcXXFvwsDHq2mOE3u36maII3eUrntFGvGRuvi05cBum5kmrIwrNHYbmPPXDu
3pYHl1ltlot05UJ38Yv+M860QMdvZoSOaRs4kqNwDI7LmoLli+aOAT+Mv3HJWI5gTZqJV1va0eU2
Jy6foR8CCpjHOIYck7obj8ApoD2QPJuCkTMn4ESF6NR+880yGqNZm8tB4Ntan4cXaWWeSOeXADy0
rxfwGYReIGU37v1sCC3RrY2LXftHoLEvHFSckj2VrKm0OCftnVhPbc/I3ezmVXuZq3B+63cfWSb5
h3S60hehsLwdFw2fMdJ9q1KNXunMLq4qk1TcDiWEDq2nYdKisuWO/9+16+Bmbjdj5AR+3FB5T4f2
gAk1WxccB0raHEfCEM3UVNrrn8SSN5xOK2wuHstxeVMxi+MMl7oMYeKsSegobtCkHXRxsXlUIScd
UmHGOdhRQAcYob5T77otN+PeYkDBmc1szzArGM2wDdeQ70mBPcprAw8+cq+ASsBOV9joC4yO4glU
RvmyM106UHPYBCUKyhJYG4pDP0cAu6eq0BZ63M60GRBSu38Mf07ZnX1ZwP3nEiJ0ERlgKQnyJIxp
cGLnYhKgH73Us8S+U5INig2EzBxbpWtLTMeRWLVrT6BVU5KIpZEwvmswYcNagbQdcKdh+XuMoE21
SXf9w8hyTxPRApM6q0DuObhcafIsz8fLMnthVr8hjd5UeW+THZNXhHEmfcUhr9kgVBznO6MjMUWt
Is1VhtrUu2rD2kFHadp4Gn4hr0H+TS31/X0+/MTnkN+/cl+Xed/4QK1P3e7esY1I3gqgNxTe3Uw9
/7J7AbsxH346AW4F9YQzt03uELRY89FjNdA3aSWOKm96uxwK20Ic1ZJdKG8mMG8h4q+twzuS0VFj
vbDGAVhWkiFSQV5vO+ZWIkJgjc6V4iG0qX7CTxVmWpPTd0B9AGK0pb3tWd+e5NEqCNKMhs3qYgNL
UA/A3DvdX9GUpeo0JaopqSoe0CIFElN/G5lWu7vjHKqh1rFuFTyd1/zIUfzWfxIuPEs0vrpGbiJj
j+lsIRAG1AY//w09j/0UM3h9pnP2+qUKNLIrO+yM2b3O1yN0go48iKTjy+wLiOx+xXhPpnSqcEkZ
oS95Akpx+fQCaH842ldD3Ct5rd95Zq+ePCCDhegusuCDJfsLpDSJJDMRjFpvV8Grheu6x4mATnOB
gbCJ4WPh3Zc6RWq4WBnRzwC+uZKfZbNl+pgvcfAUpl6Bk65v14jxuEEK3/UZnoBOQPsVmOGmIVtQ
O65MbsoOeg61eB31K3aXUlvWkpAZB+gc84OrdBhKyF+2A/iByWdbM9d8YPhVsEdAaTYwJCayVZ62
bcjKtNB8G59gVWC5deDaYgIiJcoGuxCGAJY/C0lLRpCAZy/s3TrMMQx4ybnDhQVxIcqAUIjQuFVu
cCZeXA1EMkO0m4Qw1WZ1S1ZR7BPMMdFCuThUqxa5OTztgO6uC2voJg7zMLYaSUALKhGwBGRNOnqC
TzZgENdQn3dOwAsvZ2ST/LMPi0tlKOYCIVRK+BlUQtlNcCOLYlbmopa/RS5yan10AfBUOCtVDp2E
fbqNxBvC5woCAimIpcbpQx6ROi2H9d8F9PybhPyS3vGwJbhAT4bhMGgA9Wqj+sH2kRPSSRieiemp
NtZ/yhHOLTwQ/vj4WHEUyQ6YjSZ7KEwQ+uLRC6UsrG/6tdQweDsnxbP9P81Cis7etCLEG9g+Av9W
UqEVbKv5Y8Ys9qcGLs1Q/3U1k2+TWJMih7+TyrdMzH8Q7O8PWKu/4ZeZRWh3Ta4jvoQ4/DGrU4h4
D1vcEQbh5Bg7UFqva3zNXrkaAxd+zvUrktVqJgmG5BRtWeXE2+/eNt+V8TKIV7LgTyrRYAPDSXUP
D76jFUl+7AvgiVj9f+TAiA028wdlnCZZXj3QIB2Q4lypKQqxDrwh3ptsC5AzMRO8EQ86XIpSTLDU
WDmDDQY262e4eCnD8sCn+omztO98LvgG3VX59gqYw5D7mHy973wV41ODK6TAaYh2erj+LwXDSGtV
dycrgyDv2CqTknMVukznVz4WrLkv22Cha6nQE/HvAiNjw34nR3Uc2kpK+1Wcz0tSWfu6GgD7+Zoe
q/Cv0qews8OPTKJhwqdJ5IkIKJpTTnNSn08V/7hRC2ppnJaXCGot9ThTsQMawvQw/7qMO2yCIPZl
nEiXuyz7OhpVloRYR/A2scE4yUk5zocT1Wqmh1rsjehbUq1h6nvkIc1moRRFl/DbaNwD1L/b0ytF
vkKSVmXrTdYSz3JJeUDvLQbDIy6yk4YNmVVu3dyd0nYy+Brod0oHn6y6gCJ71yFrWygnbRPQWFZd
TwhjA0PVwBfuvSDyUNVTRHrYvNfcwZBIbmpbW0ZghF2mv4qijK+aR535W7TX+zowZizQykv07lnf
jShc0n1VgJK26VXOewdz37anc/Tz/kEyNo9lDeL1k8k9XbTSIXbY5/28NJHxlftATpq0rfbifhLO
Q+5Ty5fIwqqo0hXL1rZSJ89RYUL8K9YqA6KRNY7FYPSittYO1chrXQMOHzLhGoTCf5gtZJYGN253
nfcvnu4N63p835h7+rjhuqvyuBf02ZhdfeVDeq2AQGHnaKXOR1KvFPzSdhAWs/KNFA3B9+wtNqVE
eyeKiJgcyeAx2yfaPauAGcvBvy3cF8kUrIJ2iJIZjorZy/+09ksdn+/JEfXzWjLrUchs9e48AxYw
nvwQ1HEpLv7Shio7jLnLaT+95n7G79SqS0fbiPqFJ6qJsVs0GCkfimiIuLtKqvrAx0YjSLxsFBUQ
glozmD3qZP7A4Vt+YCg3BsOPoU47ZsQ/AlAskdjD3I2JAy8GZEvk146VsvWTiRq2uaka6S4YZWKi
zYULg1NKO964D2X3bq2j823bZXqOkYoDfu2X28BSbaJCDiUROal87gGXjS3fhwAnpHS19IsUZvKh
IsWmtTFnY/YnMwEDsrTTlMlRWSJHegoOzpZCue92/Lun5jaP3AWpXxhOYCZ5ASCFf1+vfO2hvLhj
39qoZug7LU2gSgdi0WebZr3rSF+cEHZ7PuM0XBq8tvzhMc9YFFU7EMK0SoRGMeg1SNKCcaZK5sU7
UeJkx2P7GgW2MOTmBrh4TY19w6hx0mxCDcAs2CLazUAYEGSiroT+7W6/deUz9pGhL+N+Zei51kFy
I5fbe5o/N2xIIQA5mwua4nrAXc6Dly4P+XR4CbJWGsWxEMChr8Grc9kxCRjU3Vi8OOhHm7weNRIt
C3fa32vdIlPcoVOPejE77qReEegYbigvlUGGFj/WoxSgLX+qp7tnuSbbX6xkpyHVA+A3p99zg/jB
C0QP7Pi1RyKaair1179TKCNA03keOT2yXvdRHFEsRkZsEO7XLESHGBl/qPA/VqJ8ivKVMiJVbiJl
MitGRKRoHEqAJugjzAqX/wxuiu7D53FJCUnVmvUrd0sF95SYWidEik5T5rJN5/aocGqseyFMecVm
WN46sdOR4rg6jg+d9/VpZEqadRWPX4SfFg458uhTa+GJ7cM9KQD6OptFxc5Tm3CS+lNmHU99M/PE
g0Z4fJEe2KqKmWea39WT6YYz9pZ+E7kn3IDgBIGkQvlFpUq3rUjjpthh+VlRmTHqOQAuadsTFrUE
QoPgFnxWo3tNkSV7I4KZp/RkMmVm7u+BYxR6wIaW8MrWMfFpwQniD18D6brcr7M8kyVXllQnecPP
XCjaTWps1xELyRvbS4bShEiRIOQ/6DfLM+vMKMjN8EzccPeaBjB/dfO+o63V31DvO29VCPPG739J
u4quhHnSKYUVSGnQjq8kn0/bfkgt1AYieycyawPsS1NYZxnBVXjNrMIvF+W4t6CXdXqrv3jfMWTT
6aWb37IfmGoITXcvHBFjgQD3NwWPlwie7ncN9GYXia2z/mkvafg3NatnBrzg+Uuv2rSeTSRzCUmV
kwoyEf+70SKmkT/YLyVVo6poYc+66LMyT9bqKj1s7sH2WMw5FqpF+5XHfdrRHr9hv8G/KYiP0fKS
/aYlRMI2S43PYPlm+W2/26puYLRFJjOEGv88MRYwVG0TD76asDGBPGOHEf6PigyspVgS8duazjGp
LzO5IUELPIPWtc3a0PxkQN3Q4O0Xi9+Grd5UKQGwOuqquxLQj00tsCm39jpMjK/zk9MFQvGdEDhX
ICXajHenrQ/NfgEGcqGlcDzC+k9eieQJRH1BXVK/vmyElh6yB/Xdw3XuF53Q6Jbus8N1nPU6cWqs
46ICXsXpFVGVeItztcQ3wOdYfg7Rast1jUg3vJiue34P41kp/h5wQudpITKMUbvZLH5hth1+WTXC
NoXJdSMmFYl3ZCOEaOlV+sFUR16W7RiK7t78698IDyPtLSK8M70n3j2t8wy48Xwddh/Nfvlozqa3
KPmte1BvcAH167lsBnE5lFhI7yhpXvq47H/0ZXVhLtH86/NtvbHAtgS2LaFQF8FdwJZ2FpJw+UhX
07ngd3qRgexiZvmoxuHupt4we5nQGJzxvgojd2v523PQlZJLvAoZ6tEmWrk1Ry1DmxCgoXIimSYm
zM61CuTvkvk0VRaGEIhZc69ARhgR3NHPXOgCdo/C3l79n1Bi6NeWN98r05dgb9JHdvqI8fumOluZ
Pdwu1mGHKPx/9Jdw3f0WTDhY5HeEHuHESyby6qf4yVsuLBET0C8lXmV7DssN7nRmnzYNKX/Lj5gf
KnxTBCfdMVK49zai9jkdXIgnMLkhYmLgomoXjW4Ci5VODD1pnKd8CKTcErqN3fPyww02dQ7ohdU6
lQdBB4FfGYRyh8MP0zOWNqhpIsNjA+yZrh1iWO4eawrqgYU5q+fKq7F4KYEYVACpejePHs7jZFwl
cA1f8EiW2rvjKlE8ojXwdfZjN85pTiRnJb4cy8Xizrao2lGZOHFVcMhrkA3mqbJRRpk9Va6ZTcXf
QxhkMhNlgVUQuOSFWzxyy2/5jkLChdX+CDazI+/dUtuazxDgvJwK8oeTOrLf6z+DNhF7e3Loxfzz
78AzZ0HUGVQ+uTd3M7H8Y9H7vTYsoCE9eua9O9s3tA+96yVNYDS6XJTJeJxCqok9mF4QCIaq36tF
zfb6w7Gv5M8PkTf3+l+HmCHKH5nzqZgwY7AtfH6qPZTpSLL7vBYlj+pQTDzo3law6z0FfZ/cadWp
pdVGT/4FCATeG+kjy9rVbT0ix3sj52L7tS8YrRsgTjGQUZSeyHhM6BO8YxJmJhhfvTb9bV+NAkPu
LoCtsDv4vJ5pcvx1/YM7brkdGLBU3HuWVMWZJWjsDn6bKwmIlBpfsWWpyrftXZkPwTBL8pqTzy4G
Bi8Rw8mUfFUiUtgl7OJAVb1WW3lP/oKQJVcqxZOiDmcrKXvCT9GTg/OtAMtiEFlaOmvNq7TEgWUc
h0qqCIlDtwQQpZKKrxGmqwtI1WHMvpzt6vZBZ3BXRqRXygXlC/yPSjA8lgflkcHGIwegXh+d+zld
apOYpZlHGXshiFEaAd5RAmRPTJU/0llqQ6hlg95/YqqU+iZ4gzg/ZnQTXCE8GFwJQlblLTfNiGej
pvaoduNG1rwjEx4KvmxJeRQs3pTQQYExWIzVQpmy5o5/awq6TlGQibuW2Bzj3Yplv7HlpKaUa+/t
+hEoUe4s/radTA2a4kMqSaeBbgZ9RhG97Zrl2/M9L4Lau0bl2ALd2jLOh3MT95ndXGGhskGONi0z
mjTj4G9BQYHl9HZoJq8as8+g1mbLTT7d3z5CBiAM5EiGSJyqP2vGmF+RIcm+JqMFkI/vOROhHJoE
k1yYFkddlJ79JjycQmy1eelBDSHnUuXRlv4SQ7TfPJNAUNCslrLqmOFimn1sXvQ7OxNKNlssEWrm
VYJdQCOZ68NfEDOq91BU5tKtO/CqNQadei+R7sFF/G4mLy/p2GBh+bZk/UCK5fPqT4hEuJvfPRAK
ULxbwU9SxOxvgvRpk9hVIuF8jmrBq6qEdvYDnYByeERXrKuDAAP+Czt/SslZvlg0Uqq4we+whre+
/8Q9U6/jhk5mPtSVJ8gDAhxO7ztkSvVIl145G90SHEeQv7pleqb6ENiKCFEkoJmxyrCG3E3bOIY5
z5+kKkVGrzqc30BnENY3UTnEQXALVrTJx2VnmaGhhqSIfNG94CfLG5DkEIOAP+xxy5ZL1a7g/XZ3
9HY/VGFCYr01u91hMtxoPAL8w0HGI9EoZslUBHQGWoxPQ/wrqNieiOFGyWrmLzGunMqDq6NvRufP
aNEy+2rrQrBf4T0cLbDBr+vVmx9G9ZVy0hfqDY+OFTlU3t/1GMr8IMewiYP9Lq9ppWZclxale5Ld
tGG6hoCJZ+/3rgEtBediqNqIJNGKD2bJoKgfn0Fj8+jCJzM8dYEyShsSP+5fTBzywngrQkV/T510
zOP+fUwRrcRlyNBx8wAAJEuP/YX6NLhK7VbX+nsWc8G3iyG3/ZbmeXbdvAI4W8gR1phbSjWPC5fL
7eCMo3oTsT+G6Dzb13e3msIOd8D4hD1gU/jmn3Ur3yB7Y/aDiAgtbf5YLrQFbXGsIItFd+rJ6oLZ
U7tU7ptwfRSujkn2YyfBXZ94gSiRPIm9bFs4FeOqJkND7t3y33mGb2GOIvQkTMTgLMdjeZqn3xIj
Vd0Yw3CFEDSYLUNl7GsiYS+wIX4R/u8u6ucpod/VCNtJcW6QuP24vzTZahGTGSROMLyiRPdUG6W3
S4cNGIPANIuPjNWGvnsYFp37vTcBmcE0slNb17uU/9/J7RY3J+nGUxAS+jEfSfDO5T6LmLIER1Kn
Fm26O0u2vyDvlOCijzj6nx3NdjKlgAG/H7eTsrMCqEqS7hzHd2iuSZWuR9bz8HJETrHQ6DxReLf0
I48/AywItymLSpd4934q/7U6hA+w6Yr2pgRjqt0Ts6PrshdzDWH/pyDlxVSgANoTp6pAe3NqWMIZ
vRDv93jkGGZKMy3Btnk4aZSm09uhSMvM0Le3idJPw7iVxwNnGGaQ29ofWZ/7SnzT9fSEZe1wJcHH
2uS+8ZEBGnWXY1Acd6r4R+TCt5rrc6LRg4yoJSUnCpcFF1Ahy23UIWc9V/WJhWHeQ1NiAe/obgsj
pF2zsxHA2RAQ9FDvNA2/J9L8shm5qMzNN0oX0U1P9cKVhDxmtbW1d257ZYCeSd9xquCE0DcNrjz7
+EpmOBxetoh7J1Twmvt+pl+mLWLcbd8aL/Me8t9K3n4yJKl4RVKDgkPt5OFjNZ82eeX4H43OhN/G
o9QOF8/u1W2njQ8DSola+Qz30Q+JA747PgVw7RObPXM+WiZ+sVltLLgARuELvbweix0OnOrhNRhT
PrIX+V4j5xrKNSRQ/IhhAG65pNaiTFgiL7czdn4TTE69+Xk35SMZkeNQR5vmvLb9ZQfpM0rvPmYu
gQmSCURFdwJJjaNyaNwiddJ268EAHuMRnudjjQ1EN2SLtJmCwkOX5JP1Ws/VvSSIUVeq0me8dUn5
+XOTmfM1VjiGVaz/6ZaQ7at9wvzgdaD5qy2EhrqlhjQtDx0K02PdSmI33BzK5nTO9MePShW5EBOS
BWhbQ/Pf5El5RAjCGIovD97K2jHHpduCwBS0O8aN2dr0NYALAKYkaj6avktNjVKfQ0RT603v3XB7
rUP70sayzDweufdUzSPINAfflykKilf7zg5O5HjYiosWsnewHxZgSVTMgY2bfOn1HwnIxevaSdIh
7EXJtBNBefDGnGYP0BHcf41p0LWSf85+Vq7ioa0L79zrGCJd5kITe4fvAR5XHfxNCu4UbLHg70DQ
mKreJbx9xCP7uapWvJKDghVo5XC4d8aqpV9q18oA76n90f8MTCudfmK3vp4J27PX5NvXtpHQ17Xd
KxCkIzDDulG70XEydtSFKm9bS+HxIYMyutTxcWavbCqgwZvbatBA9/zo88f3HysoKPRXsc24oj7q
q42bV1RY2I61mWmiq3H6vp4FK2JpOsC/DWI5QB1bchEvHDoz6fj4DkTHNzyNjpLO4/EkbIJ7pijA
sDeX1Ta7oZ8H6Q8FE1M9a/l/5cI8KzP08+cmPUSHOetUUgrarRhE44/Lymcrs0xy4lGPPuQGCWhz
2O9WHkKAkDXEm/4Ju2rG4Mpt6vopmZCQi6BhwEkMPdsbayXizRyt7br4EGc9qzWEBAG8LfYxr23n
+2YcV/v/dSzpbyW9mK4BPTpergoGUUQtdhQRq3ynFsbBFVmoYouuQTo071TvdCk4eGEMTWTQ7Xwz
tqqeA+bVQIuDjy/q0SnbBSxPJYKtAwsT7apCmC7gW4IbUKDp6tYRdelkLydhEDI61B9hbYBPf687
ExbaCnQ0D7/95SI2XFYEqARlIKyLdUvCwD2IU8xSGiFmgtG7tkx4D7cxCxEjZ/E6RdmLvl9QRnVg
v+DLccGl8PcMVCtR4mnbwHleWk8DRtI/8Kb/Kk4HmfaFc4FvDroG6+P5Bz9O2krPodW2T0tzc8M+
uYZRwMHl4H7G7ZDrHpR+kOgk6AvD2XLUeRiR1nAjv7y+v7dcC6ccyaL+BmtMwDfOKJaoV9tYy1zi
mQPX7SgVNRpM1iIpMlIvTXCpqzl6jEXU1WSnvbuYhmCG2Hc7MHGWaeWU17bd5Bdpxf99iYprOigD
0ZOtHvP91WkLNIGJ2+Ogm25fGtjp8xHWbkqpIbGy8g2c/QuK2ztCQT6RqeKt1rdFWWkX/Iyb+UsG
2NbVi8Q53sgDyIzz3k1cY2TA0QW1nXJqyZtkp6oL+fjXxDnUNYSuUEj8dQmGfK7x9dFbPzceR7WU
kcgHbHtdv95G8Z9zIRuCwKsg059zNlSxgx5azdd+JpjBlYjIfhkLASTCMn9Z7l4vBFP1dJNZEaP/
5O59GYJz7DVi87+T63gRqyFnSx/SdfELG8azkFN28BI1hk7jdHIP67HD4Kp8S3+XbVtZKYWc5SR9
tYA3fxrLXgq+oUJ4S69HAtewjcTxOPGnOz2D943Vlsvor+izF8AAfPVwtQ/8Eyjr54/bRu6vs0aK
9hDdIsYr79YqQUbi6/ZI+L3FfLz6c8MWCE6gpdyGXp3BIXT1OCqP0+Hfm3kliMjNC5NRCdb02mrH
+B+x6o00pRDFhJoshb9WY+FkDOsVeYDnLDzEPRKrX2BNy06YdkPYmtrZe1JMAqpZDg36iAvZwFeT
YAUurEDBqPRbcCP60VH5Y8u9h8oDB/aTzWsBlmCZ/x0770ZOL2RkQO8sNB3WZRqtpmYB9wts0Zxy
MTcN94auFqMgQwboBTPjgzo3ktTvFRhagL2wz1ik/PZKEjxkt6DdS0yTUOIsG7SU+4BviOxytChr
Iz7ipIEoODNMlZdtSfgUsS51+2h8jwtvzNFbtASOpQc4oNEEc2g1Q0YPJcImWCFinUQAhO4rHyrv
rpzA0l0+yRhGCWH0DZgGdJNbzXpKAj8pMAfFVAKEZWlMF6mRnOQqZ2WChzVR4/EUckWOQTVniBBC
CM2OrDMEgTdE0zVReJYKcuBPMflg8f1CdrQykBAcYhkte+fuWpuV983v0B8Ne2b4rqu4FOfQjDef
/X7KFMzlkIpFjcIPwvcNC9NcucEzLer7le/vDY7VKZ0fRtHtuRYo0n+u42mB1PO6TyEwyeFbTnY6
G59vA8toiu8pGSas8aJoFIBNSl7CkD9i9j6ScBPyqnl5WgA2/AXJvOaK6iQLjjPXSg7IMeGkgabh
HQD7vMF6zjlWbZ9cTZj64WKFtCy2J+1YXlc1XQLNryWbsrroOvNoiKk4CpOLN+Uv9hEuMnzV+6H6
wB20ptaGK26FTG7dI8UI3L7AwL6Ytbj15MS0/8GoyTYgugOF36PouY7WZBnrjD9IBwQak5on5M19
WqJzCLclbzJIcm78nEBOTzsCRIf6OpI+TBZlVq1iJ4/fxKCcHZOxm82Yrz+9ImXbpSppkaeKScrZ
p/BOlquKBNjBtD0yiTlaV6NIQ5ekl1YA+n2zSj+qV0xCsZ9YG4pugC0sdRhr9dWCpJkFSygM4wQL
hl+89f+7uM4VmEZiXogUnnQWy5U1p/DOds3s+A9VEi2+7blTsFIUX8hfxXXYsOYkgDnnKMUVA4C5
YpvzA8Cc8nYo53ApxONtn8HdPq+DclHW9CmHZXS/B951gwaS8MgtU8etM634SFhqwO0gvvqALtwq
qxn8uwsBdhWmBXBI6tQobxE1y4dX6VL+5jVuu6Cf88nw6xpteIJUb5WCEuyNPbKkgDgBN4zCGEBZ
crOKQdL0oQvZ8Kgjhg+SxITWG8HGRMn3Y/7PjwmYsoEyQjXj7NZ0yOHmS61DScx4DDpzFZDWMpj3
JckxLGuo5knPCH2F0caHOd7BWDv7ARzv0OGzs5IB1jLSiqOurRxzDENkw3kzrVyM6MUPbtJ6Ti/7
vfEVNJAtJaXLX0N5qe0gP5gjxduTigaWVItzjtngfuMPBJyDunWefB3Y83uQHojfbBxLuI3K/YtX
GOse5/yfLFCijcaE+t9kB/238h28K6DOgcbCvo1UkhU8vGaTBFoZ4CJ3LG/jtqE980n1IA7BoFTc
4B4T6TKdBkq2+inFgMI6i4+HpFmp27mtSkTcNta4FBdDn9U8mpPkXj3Y2i80pQ0y0h3lwSgwBB96
kHv7B5cSCFMkeZg3CAUHzLw3rI5FgwOAzzKhOgZ8S9LTmoceKJARm3QClSEqn7w1rbwGQz4rLNLr
FsYO1hMX7aSYTTqTZEkjQOkGmXnsguLJ0EkCgz4s7WPzdHln+N9JmLOFh4ixyjZZjE2D76MVaSkW
sYj49yrgeSKunhjeydnKaMmoeVeAMxlRvI7qfZZi79TvICCQxhJjSq9p3yHZGcVwOLI22NE68qNm
LyCyTOXkRY05AXrQbzxIjkTGc+HIuBl2WSmIttZNuev5fCZPiY3hvtEQVr4VzTyyFCzykB/8kYTp
qFyYhhA9mIM7PdP23tws9YReWukq/h8N1WNYd19i21UcB1zbF2U0vbrzj0SqFqpuUifMBlmKmo9n
ZO1j53H2cbeBfuZwzGcRhbH2kyrXZ6WnPIrJm7aqF4p0FnfdJbeCOFtDKZdP02fMSKNBh/VZoYlJ
/ao42oHOedQ2dzyw349mFTUcIcuY0Q1kjSEm/oVgWlwIcOpByGuKsFYgDPlvL2ZA9/9obDCOYg9g
u8zHGfYZb9I+LpWhqyLYkcet5/uUfAyKHvocXq6afs6etB8dcb2WEaLs+iH9pqJlDOVTx3quIXya
jWKzsUrOMI7mTB/tJfTkJVfXk9pkTaNXvPD+0nfZtcpb+C52k4q6peA/eh0DJcSU6cjvLRYlyNKD
aexJDAo/JDg8dXy1d8809wr3BDtpdtLDpGTRp8P9xT3mFfjR3OYkwTeo8wYTrWv4ZMXIGlQBkWEN
/7aVuu/Y/R1KG3Pcvbt7gB388opq8I8Af69wnMWTuJuItM5/63kTG11/qm/IUddz77ilzpxwOpxw
M3XDUeNcF2WCRdV/N3CkY80E/3MuKmEpZOC6xyjdbbYV+MJhkAAOT7MvkcOqhE87ARvzOk4lKGWK
7O1PxfN1yXD4Fvf80lLfhusr5DUHCaUsn9nM8GEyx8u0bUZiH0qQn5P8Uko9aMsIvBKsLRkYi7gP
FZMLlk1ELppYHOrqse1DBGrjB8xZGapM4qMvIrBDYqC8Z2fHZMiZl7nAHKychtFrDc5iJhqTDLMS
dngH348ZWfOwcAcSOHM6mu8F7KmPJRgZOfHyseYGjNcwwUYzyvIaLaOUXeUfnH1aHp9Mxk23HDEC
OVN16ZGGpa6UiXSPDYuggHnVekVWHzalEca9OOBezdgAe35gdq0x5iW8QN7+wMqAeO2Y3GPCOogC
NGKvbmbXyYymCEh/EL3uBVqm3B65dLTiVV/3fJSVuiYS5h50CkDc+HpbqYcQzHX/Fe2lytcOgFL2
8lUKiLDZsF4Myy5FPPRxbWUet0xanEUgnD92cce0lNss4r7Z05nGwfR92mlAJR3pi8E1b+8vydit
FBxc6jRknIxwXqIoUNzBzF+czvFLyAvRuOeioesxNqMFcKNXysJsBYGH5x4hdkdIqcNoSYCWELgi
Z2V9hyNgA0VrelZChl86CXZhs8iNXGNHrXMXm+lZvFVr5y20+mQF9hJdXVZ/e+GEUyCKmKVZefJJ
dk56oUZBfLOsLb53GjgB6MknD1X/aTxL3Lq8qtWjlMJr9j0nk1Ip3X/rfLZlFeseajfNpvjWnKok
y6AqbJ4jrMZRH0i51+OvIjM/qRXKbFlPprEr4JFM7u277KIU+UXmi855SKjEO2RVxF/tBqZhMQM5
GNhSaTetU1HIKmLQmZ79ZC5y+ta/bxhd104E3NFsCcRV7TrkBrbqXYtOZq6vHaXqLbJbKnXdydWB
gk2saDdALSyiQCx0MhA1vSfVJRkb1GRDjZcKFo/w5g+BtOo2fiwOW2ALvxwuizbDcxWh0mrpYM78
U62PGSe6ucLoZRlpq9eZj8SirQNSexCfNM8SoCJiyrXu+iNxsa6AEILxQB+crUfKqblV0NsoMuI+
ojexFgPN+H+IGVx/qYldbr7fT13JsMxbrYJK4YCBpVNAZh9nduP1QtjdgRKTN5Rgk5CbP9CHCmzB
STN/Fhxf3suBmEygJTJwHfFJkBSUXIvgPgAoauRFDqjydLRuA40RQpQ8XMziJGC8yQW5IIYbN/PP
RZz9EJEYaCsVJFNaRuNeA36nW/bwsDxSxOTrXTAEr2V7sJdx+KW3qKQMYd7NuBPYEG5yE9aWPtNT
P8NKt7EuiIrHtW4V2IkrqglHy8+Lb2TWeOMDvHhtgEGglaZnmihlYVwxhmo4yfqjmDG+0rB2d6JC
H08b9coAnPalrVCRm54pLeFoAB3EOPMUiLUp9hR4dZLt30YXbZyrgBDPb8Vl0goAyAunj515QA7g
GaPlxDtM6TdGnViFJQslDTGDdo8IX4FumH47sn5vYI1LD0EslbK8eJthABW+YR9NopU4XSm9DC31
1w/8hVj2BwkKT3dSoBa6CS3vA6C4BHWU1cjMTnB3WsT2c53FRLe2Y/TbONjatYcrKV3ZsmWpqT1A
pDMLx8LCARj1Y+M3wOoSNmLwPI4bDnVJ3ua5TQvFLu4B1eij+5Bo3jxYcctlY8c9Q9QbMqiB+ZkL
5wBdVOUw3p1dbz3/IpWU7V1W55eoN525desxtan2nOpZtXoAO9av9gDrM7ErbTfxHZUYNM1hmJ0Q
lMSrfrLjgN1HZkcawKmKfh7ehaK7hdtTLvtt76xIhCIRNjfgCzKXE/bBN+4ndmtDVmLaJAUNAxqP
cEcDEKshXq+nOSPtLROhTlF4D3czUU16tJNLiw4bsEEHeHnvoN2i1bfZr9THB2N3JBeWtVZQQiYU
824o4q7j9xCTZBQQ9DGVdSFUHYry8KMRI2CFx1fUUG98EpfeOJz7nZug6WKXvYv7p3fuZwuBo/ht
k+uj86Diu7aKMjfhqFtY/cUtHQymmeC4A7HVmxExPhJTdD3zJ3LqfoE8SioT1B2ul6ghKtOWFkEm
L2rEj1R4cFb7wlaBS/rGRjRCzaU0Mq83K+WrLPMJUHop3kt9FRdHgguyppQx6UKq4kZNc8k+q5Co
LIcU5CEUzjiFqRBQjq/r+4Pgx23UAqhLkoYC1Td0Q/jM008HxR1zFN4A5nys9+BIk8qGR5WTWRzZ
t6c8QIkM6E/5p/OLBHaeaIIO8N0Bbjk5wcae13tYJ8lMyW6bqjvHERB1doAfKbTlf5AIbD7P3Q+Z
7hTXE7tcq2lMSU3Zr4lBVkb3sNlaOf9Vsrm1aiIlYUJ65kZs2KzlQSOJMQYyfyb3WC0ajgh5urxc
WYwv4OkAZMdkF0Qdx2j2B360mkIw6hmmDgTUr/fMn07A+D3d2heyX6eYXeehv/xHNO7FG8S/tFk8
AYlVYUYnRx3nBYvv5wIO7Pb1KVRMqfxGxMzis4sCgZ6U5GBO+wWtjXc7tYKzxNS6DL+GmzkYeYnj
MyN31SFNgOLIum5sTCscfftwASqGCkmt5Nd88C1qVbPo7N7SfRyvjJSHpCyN+2HdM4fLAY5H5G6y
vb1uzZHx2DDnYUoaLH1YPx2GDeaZV+EgtY62YD8GkGTg45G+eEh++DV1G6eassDdUIMvq1tSvxSM
hDZCChP4zGAhzzTsGUlB13YlaSqdXbXDaTLme8ZI6EgFBmdSwYyMmt43NkwGKabYxtp1iuL/gT5t
HDfTSGiVy4oAc4annEIjwHA2kGcMA2ld0JmlbMYK3tqJtH3srPpsW+tmEjqcKJBlCd9qJEdAzwIr
QhNhHFuEi3mQ/wg9ssjGl6YSF62oR+WAgic/xE3FJl5ash6wTtaUwtAMRgorWt31zOEFRcp0KRUx
zDs/KosOA2tit4fHOMp4CsgTnjIaU5XSIE8q+uCEOkIkACb/yF8AJrsPlGjCkC7JEY3A5nBHd8hr
f/onv8iQPTR1g6gfrIL1HFgFJnxTqVeBQhO6eL45/nT5AdgxVdiIY+ndYeA+pogXZVDoXSrt6zVv
6XbiRm861ziLMwr+bbb0chfEOHh7YkTUIO6AW+ySQgg7EetP+au+XGWWalqfjfjsnOKNyWygwNsA
uY2z1jxOL6Tski/g0qell2DpgE5OlDHp8rsBpwQvbCDEhseiMhjMnnFFeAv3jmA+6VZ0XggtHUae
DlApN+SI/cAMFRXwYC87qpgMvJdyZ4EXUcEf0kwRBDX3GHMT3LIJ+cbxifQWsmNuR4iPmDVWGpT+
ikAlHJzdG5CS/2NKmRQ9EE9z34J0qo+fuIKR2+1er/qsrUcJTFf0bcpzmF7Lb39EPsftQuhXiBpn
mtj8DaGKfs4NognCXfVpzlFLDB1RcLv3sf6oMpjST+BOgFeUXLUKZz/L32MWP3t/DrjAFTtIUIE+
FH8Bv/50F0BwCV2dz5wZVwP27gTwjUo2R4XwvTyXvbN4b6jqFi7Ub70apLDYOdbnRrtUWS3hVUbp
mrorPWAd28oAjtTrokA1Fbk7l6ldKDriLPBQHt8vNBHboO+KUjHZDCppEQhTEHSVMIiTPOgR7NX0
9WSgXE/pdihCfd/FJqkKz1EJ8E2F1iM0OmNbUgCTPgQf3jUrPi36yWYC85it+8UBShQtoVv4wGUi
PaywhLTdxPl3EZurB1RXjlLnnCDbt+y8b+Iv4CMz/ioUAvrCte5FYR6P73t2t7GrIL2yVjLWM0hG
PBzxOdPgRGTH/zz3rfXNpHfqoh9qisbJggC7ALC6/Kf4k9Rfb9dGt7tiyzK59So370GPMSdaNqOA
3mHIaSTTzQf42s2U65en+TuMs5pZtrXML11Oq7pxdpeblLR6AcUavrprLKAhzCc3n62mrJx5wndd
F1DFZqwD+MNeDedVjwrkOk5s+paGp6Mcx5EPuR79ltn2aGpPyPOW3froacRXP0akbZXrklWmcEH1
bPjmLcXsnCVRnku2DiG1Xyd31HyL5yh7YQYeD/5IevkDfaN6n8qb2+c58H+9qQSMiWruetkSkZ5M
APszgC7d1suiPrjvaOLOD7Iuf+bnv2f/oE/am4co3qj5ZEe+/UHS4+DyrqgSh2fh0/d/8tkEf5rK
tUmUdyKV7wi7gvgmGal1jeZ2/NCPhxnrdK1bFXk9s9SFAygCLJbkaZU14B4sPuAnTPVDvsqpXQkH
dd5POW0+FjupteNsqL8YtHyLgbxmlnt1H9HRKnLNhHUP9iMPk6QrKPPuJCq00U1vbi1XwYD45jd1
SZ5mncZcpjgk1liSsRwLfgLleSg7tQv4Jp0/T0NgFuN5G7lx3k4aYB7AfVLgM2XiEvZUwc7jZqZs
meP2MfInVzSx7DVMNnT5vtCKaOu4B6FesTYs7hI2bN7yIcpNuF+jGPp2VLMs+gQBckOU30myO+dD
BgugbLnU4KWJZLWmSWrRqvDbtgTELNIw9hjLWY7/vtnhdWfyJyjm7oDvuRGcc8jT1hRuJAyaD77L
hC40J7hRKhYjbLN4R+UnBRZ0wtthsxEwu6k51mCzhXEVnh57VPDl/+iUqPG6QqPACCMeAkK25KFf
x96AP2ndEkaD3QShzo04g1Esgn3iJzH8ftHM0YE0rnbnS/MM7qbAJ8T3QvMSmWn0Vh9tfHqGSDnn
1MHOO3t7ZDO2zRGpMRZ2MsbdIoFCS7WYuKB4NiOAt4Iu/6XWE8f7LiSqldr54T5o6nZg199dw3JE
zWU+atomW/LgTJHWxuYkD8Q1ZazTJlYjepDxGYVh1zbjE57jHPzVTf7TRYYO5H8WDBTEioKBanpa
UPhV3mDErCpsBdl11cGWMH9werGN9kkI8+tEve00JfTCWA6Q1B1h7c5JlSNVxOTOIt/3Mr0NkSZC
6N8EeNCx6I2aVJCv5gNcAileByJ6UPKX2RcTisgv2NWpjuii8b6qFLefkU20qirKzj8R4tj380La
VObg4J4uzE8i0+WdnacwRQogftvIzZs1KMQKbTQc7dpljRpOSXVTKC1L82Gkj2LfWtAcrR6i+e6E
/S7IqRKsm9MLpMAueetOz1Go9MCYYKNJXge031IEVgLXUGxkToKBZd2vqbJR7+qn6W3w4dN3vDGM
RVwvrfLy0jBk1Ew2JHJRWh/aU8MKquUv+266aH66ecIuJRGFuwqAfuKYyHnu4aA97PcgRdnUHWge
4Dz7fzTjrLWp86ePEpcyCmEI9lD/SvmW9XXuFU6X41pHAPrYrSYzjaqjWENUnUIq5HSt6MZhAogU
84B/rceM0LpKyG900R80rZfAFAXTI2Yhy2N1W1f9heqzjPKlHskSMxPDutemAxgsALPjbebOujrj
KwHlUBFcVVGz6XaiDfiWVUG1EaelDNerHpXLpDV1rpXPb2d1ogccX6w76rJNV4ZOjAndzPF8cut1
wJ3Jv4ACZKe24q84aoGnw/9EozFGzIDF+bMo1x43aXxapFi87wyINixhgapZeSFLnuwiBhHSNoa/
kRU076Zh1WjhHGeRyE6RXIvQLsFpbKjzlqXl+mFXLliZFPPmeF+27Nv/G5JXjMnlgM+khg7IeQLL
HWROVA8us6JYYNqsoXDmB4pxL98HgAjS9hDbVgug0C7lIbjR42x80Lsua8P/h6D5N60Nmmegjoyr
Gc65hna8NEzXfCVgX0ZeDIuZyP5IKoWda3BWu+1acDeqlTURAHQwFveM0C6Hykf984ljpRVwQ/R0
ACs5arhXblAl6xXPaNJOHSHyu+bNYX6MMrcEAHZeNbLwwjMvU/W4iswCNngnKBo2OYOqnyrtwU87
y6MIduV5vavx/bNCkH5QsEfg8md+L5RQk9lXpaPUSJR1vOF2+fVYalmfxUae9zHiByfv4qZSV6Ct
u86nY3BOu7YwoiFhmOVHHCj4rFEVhF+hRgCd2MuXjYp0zVLRFTthFopm11A727u7In3EjzUdGVrf
tGljZJzvUa84NSYP4hZ+4TlRol0NL6JZCeKV6dJKsGXvRWT0pd9Fnspz2C6rs0q7OTkOYdhupYUo
BTTXIREtOMdFlTQyiU4bME0P80aw3nuF9i7NkSRQ98qxONwtchmaoaDBT0oO0TY0kjzUF5jA3ZYS
d/1QnNaLtola3/O5rmi9Z0tTR02dUfSJwUWJQCFE+tt7ZO5xOHnx5dNj8ItnneOKFyIYAyTEwQE9
TEpQabi2dksHArJkEX2oY561C4b2HdLtAf6h65wu5PtmmoEWS4ZUXtcu7xP1SEnc5hZGwEQU5GZ0
BrTJZI9WOIODV/bT3xcDanKkCkbTUilQZz7SWkzqd02medG25DyYxHwSXI60ksi4pdmmG20PW7Vf
cysHfqujq3DPmB8BXbHteUS3jO5fjYl85BHbUGVp4OIlYdAPPJikBSRy2K0brc9I2wDqNBdb4eIc
CjMWv9uQRhe7KzNCvdUkKFaPDY6wSSuTz0zTN0RQ+T3Xg1D7ftjE1hL5GiWEB/3jzlmkIgRmkT1b
w/JVbxyrtbivVMnJ6UbucIRO34FqGc5/S2AVOcT9q4/FE3G9qNbDKao2EqBW4ynEeZBXkDa9pSnK
B8CtGM0fLZNRyshimFLO4bJxNSLxBRluYihppmc+XSEcPz/SP6741Zxt15UZYTRvSbUm3KlH77Hk
pEYrrSuFLPOHy2M+LJqJmr7oY2yi7O95z6hfvYHS/QIeg0t4VG4OfmY2N0/gVEZmKAIde1650UDv
hT7jR8c9dsfR0u5W9AiPialE4afxcGwMUvrU2dsZDs69c6pfLa11ue0OqxDy9V7pgOwiUJloilot
5zDLKA46pdtDF0zzB0JFapZUSprReA9eVE5cSFVfUlmdcjBYzIqHiJrZAfpDMMplH/F1ghHGc8bw
ss1iSjKHm8VDskTpdLw19G9leLpadpQAEs9yoqH/uVlIl97wRUG37OfNpCM5C4ofnZY9CMmSKvRu
U2d7QOW8QeKOjzUoCWXyBKpA64hWWdcN4N96N7oj6RxpcImrTpH+zDXVMPXJ/S6LDhqO09aW6CCw
GZEIuLVOZgAtT/NRP/tfFJuURiQEYDfP7ikHZeXfBDyrXkgHD/obLmLP1V9e080ezgoQAOwKg+Tj
XhNdvnY3lhzrwBy0xWw8TnBBHpW+nxUnYMiWtG8XDR5im5ihWDd9vDqk4c/oRl221Dcc16Lr+S/H
iiQmzkoIUDV33xzQd+IlcPd246APiFBz4SZEcAqDv94o7HKe2oegqK4jQeT9mKRco7vd6vqtFbVT
eOkUT7xUT7knFfZFsPcUhDwkOuemVp1owTnZD4ZNFSYeNxI6z7gs3+bcXLp7vjyzXdTYzWlrsll1
loFbHJ+ysfe9W9yn4J9XBr6j+IWA2U01mF2bWRxqHqGA9EDyOWbm82iKb8RcdgRm0pNNga05mB+q
e7GWqMzs8bBmChVZZxbG7tle8z+Ez88Soiyv9tq3WgGLWOVopjCuvmNyYeH6CZMpO5ikxUDGUMyD
7phJWzeskfe86TqVvm5xOCvg16vfAZR763VPRK7zw24GOjJzXbTlZPUc/e8e8AEZbQob1AdoMlNF
karfdNN7AL3hpbuVINcMFrf/DhCSfzHP9hHP6IfpHff4l722fK5fofnl9ycZ7fb1GFFWijkvVpAo
Tw5z+nF8vuQd0Dc1Tvi1sdspjVxFiSuUSb34DRN0uxNnTfvlauWwOUGDR11hsZ/k1d0XweI6h5cv
XxwDLpyixmdZlL3xe4sTwxrl1mSZRQAcoaf2udrtY77rMu3aiz9aVSImvcGFZuHCfhXdAMz7L9jr
kfH5pH5aW8wQeZ0s9yWILaejrJVk0OoDGt5A91KXllTuW3WL+XzOJ6mDSG+2AAi1ywmpAD+hk7i0
Q7R1n13dmYEuyPRNGpYPsvRezA5LuYofLe4OHefqlNBgJGbvLSs6GV0BSsRTj3qjNepLQi5Z9eHn
2YyF2Gl79RjH4/dEfW3IAKsRjrqCohRZV+s8Ra08eSF+fvFcpMognyVY1KF6AwE+6A8Ktdh56juy
WaZw2RbD8EWUNUpiikztxHXefX+kB5JqPRi4Xn8/FVJYgmEvO50Zx2WfF+Nsmj3RGzesGrtZfKbv
XlgeP9RASWmcB2PWUHAhpcmcBVzVLts0NKtWNOrsEOEdknGV1GF6r6fUIGLjIB0Byavavkarz/CN
1u/Mi9RT7MuTUA179x+Sb0F9/wY+HSdOcdvB645sXthx5a102Etyu4ui8vDz1ROJRh3cl3DdrZrJ
PnSac5dNfa00Bg55VLEupFjbRa0SANSXcAADKPiPK1m/OkGS/VWm5Jy+Rb2BbcXJ4/BgewYhCXUn
7L6reiRJ5t8Fr8zN5zPeSIcuOQdeh695LTIMU7m2JwrdUV/91Fe6DchIAu0vvzwY88TgOgQiVo6Q
lQ/7WEFnlK6x0uAgARWBX3yZXwN35f8vhjaABR1xvyCCnX2pNqj/jWWt6si3wnytEPqz81AdwAHX
L0AIfTg1zeauWPUzNQNr2ZCrFBIeIBfJDZwtFWeE6PmhKjT3p/szRCp3h/WcHydY+cNH7/4fKC8t
7nZiYY89cL0jomHRHG+1/JzpAupGaB0VqswLwa6GQ4Q8ixAQQzzypSHEORXLd/mb6UH0xk2cpDpb
ryRfdT453OfGSwGLx17jqMtUzDKl3yqJp2k6pQ2fdf53G9Qn0EAQmOZzcKahmjsG61SJUHOtpJNU
K8iDFrjraihrGIkTifkBytK3PM1Vw8/s8DqTcTGUL+5wLnD4GWUu5GM/2hblKAKx/Y22yPrvrw6i
iDRW3BSQCrnu1q3SN9DsqxnuBRR5O7Eb4r109G7Apfd1UVEfUeaRFDhpCECpFykViyHMqAUoCUGx
xJThBh8GTr6OsFNedTiblCIk9LCp/8iVv4ONxmue1J69oc+q0SnPPc6Gw8cxPqg/sPVJ0CBBflhX
K/JrlS/aYrqZTvvLL9JVcxVN4ID2ZYir7lQ9IlA0J6ETG8/8E68JdzLXwfGuKDL1nYSDq5Kq8xP7
nDgQfR0yVRzUh0aMMPS3ORZ9lojKbRMyBzMJkOyUI9znSr7nkwEUphxGP9R5VMfOUtcbALyxIy8t
/IhKIolyT5IsO7LouBwgNMato0NwOlEbi+njy7NzUmQWFJvTAq+XSU2eoRjvch0Q2pFuOUl4QvJr
PGAOsH0m+s25SAfSCjKwCdCZYddf1+7t8nkTffGZOy0eCKJ9ZnVZnmk6T8+IwjN09Iy1A+apz/BQ
caDyYYl9T4Jh5/ilxMaQRFxbxdRK4cxQwMCfCIgZ+ptZql6XoMjVq490mky8puSbdy/Wyq6JaLPR
xftxjFe2KB5Owv1RKEzCy0+Tq7w92Ws0fyDFWRdaiMTZHopmh3dBaR62boGPGl3huF9tYTGubFaN
XjDkBI4ibezlAkqHtTQTebQNNd/pXzWL5NF7skBFYLqm3vVliSyU1z6ErmUpQlSSIFWTJ3DiVrik
usSvRSC6vsv6wmzQ0JWSkELqzoSOW2Qaq8T42sz9KCxJ/TbIdfsPMS1sJhxNNcM3ibSF8wLNWg8q
iM9RmvmOfn84o5koa3yYCL1Nb1p2OGM0I2HFekDuHIR5Vt44M2KHacBj3mui6HKhF7AHX1JTX1j1
SSEbGsUAfE8LnyD/XwbszYWF928NkhD+/e2T7x4dYQONIOXtC7Qr5XJQ5jgtOWgrmrPQjvBXbL7E
LW0Z90C2UWK5yKjnks9PHfwVWXMjxDE3yJxN7CYbNoYRIjMtT+atcaamh4ywYl8kfL1pNzORMiJu
HUdvo8mDblqW45BC2XfEorN+qkxYPkRb8bWaSx60QAHrAXUdA1LAjvwvrmE1dk/T4XjuMJdl97nq
g1FsDrmAFgXkPiZfKGLr61RYWsQlIEq8jNPm+avEzEC+1ZOxVLpt6JM+4p1/qF90ENAV8BhrOmv8
LgYh0vC+n3nxjugt5nNvnsrH6OJ0aDNo/MP8UtLHhvin5AH6im3g+Dt6E1ndyowix4a0ZTW4s0JC
EMXDD7L83ZA/gI5jEOPb2U00CZFgP8ghmLcjnMnEgI6Ho6jVzDO4oe7biVUS0B6YeBtO8Fqmho+1
7nfIUPMjSDMt1BYRcrpLrM7Uvyxopmtx9qegQnQcOQ/MmlLR6S1SJtF7blqfDLgfndQuRHMte7uG
Ck9T8WcnWhraDZZJHt9Wa6vGhayYlCQU6TslvFS56Uu6DxqQyJpKcG962vKyGy7pdaQJU5zj8yrD
HzHwUdxrd1LUeGIpv3zTwwURcpIs07gydZUR3MFu/mDJbcO5gC0f5CLkBUp3PbNwZpPcPchd5OyB
GSukR9jw3m0UavsHK3IHC+UhF1T8pYmHYLikFlX5EPCL4BWxvBM2bWW82C6B5Lj6hdjHq0pmGRp+
szZ4oexwhtolOe5MFN83G13EO7YOrD48z8Avmnn3XbQQyHzDssA7x4vKnxLwBPBXY5PwDTRSnJ7v
36VKFuvx0xpVLidsRPnN/FzuJi+3msDO+fiOcL8uaW7HnsATenL39sieGCj1lWtv5k7wnezwk0/4
woGNtZ4TtvaCvKcK2NtrgIQpECc74I2Vcg9RJ6X6AzklIiwAtNnXdiV2WVZVcC7YopkkDpdycEki
DywYlmsCLJV+mQ6rQinww2ImdK7M41+pxwgRNCWf/aY0ic8DMI6WPkfPF+di8DLi8dYlDtM/p/zX
mICFUk8PYn2434EFfGuCrEZdb4mcl6VF3zvJ5XH6ShGgWtWkpgk6dLbZAS8/Eit3HNgveb/g97r3
DIGxcuDoZBHVNB3ystxt3+2NFERw2F732JJjlQFYguiQO7trmvH3ZduR2hdUbwGZyUyKh0c6arIB
f4+K7Akfaet272aY9zjdutUeh86rK12fUk88TJD1QJ1x7f91/60Qi8X62pcM2XSKBM3cuAh4X5kk
Wg5mXAd53nVgJLtvZ4wCTrMNZMmOm/edOOW4mQyhBMPQEl0M4McHxF0K23+WJqJx73TsmPISeYZU
NqCue67Udc+l4LkqtV5IIfeoBA5hMQlnvyICNU1FUwR+NfxcE9PtaOZ65CIsI8tJZQLpaUgb3qFp
i4SK/DpfFH9HNKeEexbBvD7d0A4QplrqWtGVJ2DQKdpoCjN5VCyIEgzczDiauRfQDQNYs3zsNEqZ
BL4JxLW1kJYVEDipsw8Qcx0To/w54EXrYF+tvIg4A3bconInw0ARQ68YrCaY4xgN+khD7a5+67vY
dWUyOr7pSvYks4BegAHZLv0Yl1XtWCcC77mI8E6BUL7Apqfw1B1HyL03EKCYaxU73kTlU1VupWUX
W3uSC9lyt7qNOdSRomcboTkXZGjluna0QpMMXMTnae2ExwZ14lfkmcSP+/7jcc34gn+BVAwmuOyL
mFT22yIUAmG69454Bl9QV6irA2DlNJphQ7J/xaiH/DBgfqls55s0DIbjYT0M/IvEQeXJkPWm6qNX
uXqwVG+yRwR05+gQZIDIADAULxUYg/at+QjPWQaoJO6VG2NaYyvRCaE06n3nhaGYx2fHkE5VGTAc
2pMBFOqbmAMoDVXhyIj8VY/Q1z59BGG5ydqEN1e4leviYKC4FX989ezNPgJAqKW30smc9Vxoauup
npkj+Ooqdug8tPVReDVm1mTgQ/6c9HGB1N/+3fKUu0YHUQGUvVY/0RTMR5VYtc9A4Mp/ZJhAChBo
82gEhmd5gAuZUvQyjcRb34JzAcwzhz9QMf948as3ttM1MiYvJC/MguY0xYDi6ZaRnWBq6U9Et4/Q
7K8OED18LWSWnFzHrc88MP2R9Cr8rmeCzPj4XICF6+b1HwuSP12aotFIc1dMNcKyLzJ/R7OuP9sX
mk6WRklUeHuBs7hyDsoSvYrEKujjk93RjckEZzFu9yLVyBwtMF/gAsjNMm9+BDkj8h+FTMeOBamd
Dvnu1DG15n0gXfYeeKTI1mFLlBblMqCTKGv6m3rdDqGwREzv+c6m10bp9ZXG8rwSqndmfkATEsRR
Mp0Ib+uyUhV3BNLcZ/7+FCGsO182O1MLcxNfydnNN05Rmwwd8q7F5Z2KVnQEH5n3fDk691WNUuCV
76DRsbq8K9zQ+25wMr0B2dMKV1l8bfxYRxzvJvmkPremeJgBleKom4b2Cbr3J6JEnX2Zg+h9yz/L
PJTB0UUtGOUnHxROr8lSxbraMimP19HZbs0Z8n74P2dqNY+T84kjmySdmr3cl5Vtr47KAavQdHPw
2aUj7SNMIeg00tstw0symXiba4josT20jgJ/CJnWBjgF4tJJ+9mgym7iLCmvhStfzkg6WuzNQkoB
/b9n28jmjcY/eACECXidgbBVFJGAi/z+QBAVPxSy2sC1eU/6CEPu4qrTlISuErCVlRYd5k75gqOR
fnkL8aS2V7m+hOH26zDSPnnThmVyf7K3fYhfl51EQnU7LtakQhkAEUNGDlYGafD4gIl4OICZ2iEM
do3KXyAvXurrEQOsKT96OEYU7ZK/v3WBouFuyi9H8saXuJCU1OJFpijgYHhdNO3Ekq73/UCXOVRF
NUhSWKm4D+5I+31/ANECCWkowPfPTkqFNyAg/g/5P/ozZDMnsAI3jqSF9IA88opg0Zzdks7ME9Ih
ImXK3Peoabnl/6QCVreN8zGqyAj3oLZkuwvAdXsDjGg8C7pqFMvbBroFjZGNbT2E/eUcAD9X3RYp
vqiScJ68Vk5fz20EHjSJ6Ht50eBf+DOj5G3sq36KO2Qq8xyK/eCj37dZ2OU+RV342aqPdCKuHnbf
R2BjXaP5K3aluHUNhezaiZ6GlAhBqINS9r2Lu1eqZgdomm0xpGxyWA0kpljv1F6gIasDDxsdLnLF
TUQkmxO6qLOSyf8disq2Z/JCXnazsOtg2pu6ZJX+qGA199oQistVfcxH2CNXb2XLM3bnUjK5o1GA
UO8FHk45BrnINHlUksyyFQEAZfDT7SJQnG6aWOQOwQjAipk1w9CdDEcOmToMf2myDbPvHI5fNQU0
JGRCoHg+thy/DeW9YffE7AIF3TuB3U5lSJaqrMCYQKH3+fuaRzGWR+4n2kqp+s380UvCKewGZV4H
8bodFmzsRU7Dxt1uU/fZvNjMywnSFb6dYtt0wzvP1Ffe21ewTY7fBez/Qh1KLVr7cWlDhlRHZP1z
Ah6JmPLK8WKN0W+L8zB9WwrdUJvfSWmuF8QATh6vSzLSxE69PgZ7uN+2QNHPHrkKWGl83jZV0YDY
asCgiRzmKosZlmiuYRIOsrMy+r2PEhXcTLGEWCCXm3HZaw1fdWDAIHmoeMrRMwYQSkogHc042q83
Wb1XyXj9+SRs7UJqxl78snv1rt0hVHNH80W9ncfcOEtY+02r1Brt2wDPycufehYco9RYUWTc7nKS
KT58AZuPiGJYwRyjrPfFlssLvlHrrb70bO2U3wNU4jU+j3AnZIlFLKSEoqwomMGOTDQ/Csiki7o0
VbBKUqAmZkdS918b4fWlYIb5LOKQXAO39LJYhkxqe0QnmVyRe37c5HRjUzO90l3SMI8Ew3YfDJt/
3xBUpauwqQa6f0aFVUa9QAA88dNa6atj/rgojXs1cpE/m0DMCaXNW6jA39Fzl7AUup2eCNsy7WEJ
JsEokjLRxBwEBIOJ/4tReWflF0japgKMBWYS9g6+/3Zkf4GNtNSv0n9D4e2y28bwWDg6ZFCWTtHc
pCIiFs2KSxzlt0v6CHuAL1a3alvP/YTLbmrlc6LADEN8hvTeQQsHBkqdmk8mCCe8zxrMeS5UDWRZ
XKx2UDpgAhkydCNo9d55+qfTBI/REuRg7MT0x1AxVNxINJhkoc87cn3Him2F33uADS0yEpO0Ntix
CUfwQMmrYe3ZwC6b2NbhG1GOpXGQS4dmGFIE+7ZMVpsgVZFMLwXQBphjsgsAhfvPRxT9uvuYKuqR
3m/hBJ8xXk1frdD/2P3P23yWrt0TRHp0MiCpU83Oc9u33v4NEjg6FX2IQrf/p4S5PUJeSwb1o1MA
7KbT0PG5XYsMQmSLEEqv1Im/w6LUvbVOjEQ5tS9xWpSpCqU4kE4qk+Jp+vSpfGctMcoPuDIe6ihn
VUQnha0va9tFSmt4rD9qto6LYYnq3uudFMEqBZyC191mTH5TPJLNoDfjxT2BygLOWthSCaKryfeb
OSThxI2aIhp3XYOIUQ0mQHm7/8t2k5z/KVdXxISeUAfozP9uvAhb2yaQel9CfidoZfvNqz0PC67m
o4Yu783ITKyTyGuJgwiw0Xr6Y0i3ywD6aO4NVdY9O5z5fjr08Y1cp8rXpeZFx6lAoekwst4UxEDu
+ll5lu3TxPdqlD2nbeV0kHHjijor0b5HD0WYLswb8NAlJ3mNcmQTTl+ZtUM8GKdNdsw3hJFYKnCj
SYz7eatxUV5TijangIawneODxRnAyMPZxpKg/BkAA8GTdKexVBPxB+1TUls5UMbnWPL0AFn1lZQE
yUan3wyvqUyeZ+ZxfmPnGS7TINo7K/BX/Fu6/6Q7A3Z7wErP7+wOS8CgmWglxirlGPI2bRuiDTcf
JM1amqM+TVzcE3X++IwLrWp1WIBVlVKjgj2xEYJif76ZchriCx4fXGJR6osGjKuy6xcxylUUsnv8
NEfxgJZuF6b8Zf14++W6EWiNT/IRMPCyvx1FxI+C3JILRd5vGgDCjoU4nUXmLpsXAV5qbiGRghfK
BphDI/cba6+s22AyHNhgtok6vXUP1uK/gEK6mWVl6GoDrBS5waSbe6v7wpdOy3fuj/oUOth36U7Z
W1dG6KQP43QSgJ38yijIZhbFrjyK06CicRXVCwhB6p/OQBPSwsUdnXIKXU7Bo3775+gas8yTkz/8
+8p7KeAcouO+Ne3cli2Y9DHgBtMXKdji8WS1iIGnGkpaKO3xCf2ywU16KfRLEZXsipLR4UaiMc1u
fFDwYjGY4pbaCzJkTM/Gg2aaiTB8WCrlkUU/bDXlLc0Be7gzRdhSXComIUHpSac7I504xBtJqpTD
3NUlepFwUxU4KqhyC/4pTjYSKfQ0cCeHL5zsTFxKCaQJkOxmiR6nd3ndLIi449wmdIDQ1jV31KmH
e/PlYyPR9JyBFNaoGWn8d2L1sWxwFfWXLG+tHZq9YddImz0wc/QDZxU7pMo6h6ETOIZ0UG6DZ6ap
tJ8I6rNrNXnx7JftoAYedax15uCJa3KLOe/fkvD5jEQau7sJxLAYJXVEdXS445Wg5n08xCQvdKM4
JvtLHTwwEwFYuc6DZQDU1T/d2Ce1pe/U7P1SRRXFxNWejFnWwfz/2MrR6CbBthPhIgR11NQ6HP6M
Z9gpR7F6PT94K9jqcKojBporYDCFZCXezHN4yyd3zpL7cvPkYT2n71wBGEhMC4/pwQU7rqWwGIkR
8knDeEyJoSwyFPFqIkWxyebiW9GS3Ml23lt0mX7UT/K01r0oOrQlsHXXYLLU1O6LmqsO9AHNrQUO
gnw8sw7r2LQwcHISVSzcyr5wOcup+56+c8e924SBNJ4QzmudiZ+9RowvaFnKbfTysRrbjc7nnXRq
iC80EnYnSBFhMcaIEmn9YBVR/+agFhiHKe1EUMYrjVE4GW4CRGWxS9JWA1+LP88/k5buNA5I+x+2
XPZCjqLzNpz1BIJf7ytaCjOmsSW3S5INMHPjuBuja7/8jqZu+sYtNKXHaElSDgKTENhaJdbieRsd
X8bMQjVxLMnkP9tyc7eADsPlH/3C3mxLLRD0pjG7U7Xyql05khVYjAhCcl6aLhuCOgD3DTJo49kr
E5nMr3bm4hl3imSu1/Ji1vvBmrWRGx2O2oLR+kYwBJZh10ghLuqxhM7BynUEy0U+lsE4R8760jyj
5g3ITRg15mlARrIYy1XuCuedvGLbLvA3ji6rVATZUVCR2zko+PDKhCy57+zh+Lio6kt7ClcGHSAz
7Xv+5REh4uJonlIsTDXjty30k5gYi+gW3nJWPPrRoS+6//Yxk17ijVho470x9rag9VzvLXBO1EWR
Hcpu1J5SowQW8ZCawxw+A1XQraKfS8jXh+AvaJoThVvvEoCAPBulrbaLOoFKgjoOIWmOgf4igx7I
zyooCm1UmpZKM/0x2fsl2bFwB3vt0WaW4d7dsv/6RAG6mGwybyRkg3KLUP/MOKkX+qM6RFMM4yHT
XYTaWdXaRvlinDeD1N28rj8r3HePRq//Liq/Kme02TK48AA4KWbOpVPPmOTXPNw9aQApxXH5upnL
1kEXizT/uhQuoJJ8HCKZk1oyXe+SdeMVa04rrq2PntcGB5CTqFTE9ZSttRlbmayvfAntX/xZCBld
73ns1/pm/p0VHifEjLpe+nkCmUAJR0G7SsKOrQxydOu9baloz28YuT24rDAZgglKqz0e8QoBnNS0
YnWtZOcX18AmzS0JCHPzgIk4DVK3dbuT+ML4cGZFGC1RfunvdHT/QAzn9VuTmj7Rzd9ZtVxgBdkc
J0VX42xy2rcKxtJ2Sew3wAAIWA4aE2tlRCes4wt7FzaWSxxajdOx5GgrpLYI92cNMMC7wASGuNZ+
D0MijO3onH5WPjWqRSTvkDmK9ARV495ghSSrpomFzwYEUtRCW8QiV0OmO6d2fqYZrQTJ8pT/Kipy
xlTRVKsAQxWgHOzzswSBwP8TLMItuJAU7R68I7HOQhWDGxZ1FXeZcygtg3QiRSM96JQTEMcrESpj
i4qftCYGu8ESALd3bkB/2KGiZCBznt3rCGTys5lzslLVOwVHHl86DVH4v9fsC3npfraOJSaczt3U
e0RoAUKqFuwzsbz2111yMlNJdQcX70jn54/P/LmxrY16sL3XzFSaA8NXhTIexXUn5H8PH3t87H4h
59NXahu87ji6fAwLuCozZq7kQn1RN7jCK/lacYy5sXjvy/j+NFjEsng9nAvVAiiVS2FS0ypPbXIn
PgkoGPEwE6cj8i60SRm/A+nTGvol/AXB/1H1ngb/tZy+du/cwEcvWW+3LQJbdO35DyrwGFjufxK+
qO5rin9zr0sVArDikO4rsRWHCRgOZ92cg0jankHj+/hIFT4D5QWKVZSTyWz13YEQXJ8u/lPx21wp
CdTPTNxEEN790qsHUs3cHjrYcEu8pVZ0/grGf0jibuE63s9cLNjOpNh4o+OcJ3YZtjy2WI5JCQIp
WvDiCG9Bd8/Pt+F1c6BJ33wyZrFXclqnK2EfP3fzl6+qbXXP83lZsE+dU/OKoKD79y0AFb2EgRzO
EOCP3puyWNvO8LMJdoYicX8r+5tQ5dMcuJ10tT7ql8Ay290RY8TZvj490wpr2bokUXigZ30986f0
eoiCKFfZDWaUcF8vYeUiaAnZFD7+I9dt63SzdndoZAyIdighhl9OWIMEpewSaBNlcyCy4YYbYtnF
mMtlTluU+fBqAjlzBPUy5Wk3XFcIw9aGqtZ0eIRfrht0bMzdRWm5tQeVM7q0GHbcGORCSUlgBkY3
jwk8tW7HBpqIqX9pDIpQQdrlvi+gjEjO5fDbqe0W57REVUF9XySJmHgP9VdO07R/O9d2CDd7cGUK
ADSid+v6uiKV2tT1PvtuO5TsrecWhTWG7rPwJ9a6pEOipC7cOE7ydN8qz5UbApN6OF3KHasUzfYQ
NgdnWAWGtpY13UDBR5KI08BKGAVR/s8ZD991n/ldJNi+fRpH28nt72QgV8w14bRyg/iADtWYnjpD
GgVd2IzT5ZzfR5cafnUyrDIer0k+l4Mwzp3sFJoo0PfiwCtr+sq26SMkh1SFXJwogZXeX23dfCQB
BLgRqBrqWswsGzt56IbLiyl95R5z0cQaG2FMe5AlmMlUjNXZ8hFDHPESo+D/TSXXUF4V5GpbhsjV
0inG35bScWMUsuzAQ9vXv7Ub8GBbH9lmy67jX7uSm1+2NC3T5mFlwcjeP6WSnxlCeLFGRDmOXi2Q
bZXO9eeBbDVbo3x4uXnI2jaspfSqREiGimut17mlxRsq6hqOFV0NCtbAlehqGsD5PNH9pra4jK6d
BC8jnEW2h5DAu3+sxBT/7mIfKH7R6K352+cPN8qlYp81ZhEcIUv+0dPoM6+R/XJ2q8+/wZjMR94S
oiErGSdM0BxqYQfdtV+3SAMchazn7NO8Y0BvzHIUXsP4FTsJupwe850b9743PKX1XMTzeHOLagLb
kHULHkqauc6Lfj6o/1lTgB9yK2GNfrYp2PtkZy47TkFxmeZEO9ubZQGx2yepHWgq9poPJml4+fSn
q3zljiy4UdrMlehNWWba+JJEI62H/0NCFtvEk55uC2HGuCh9D8O4mPC08mFTt3FRwIkbznJN6P6S
1VrqsT+Ueo3SvKfF7S9Uno3/UbkBNkgI2caQcfBFHlxa2iC93pFK7IKTaGJXNsBCZpEM7phIvVlH
qraNOLG3CALrfVqALC5YKoYHtZyOgSFarPfj6opVSqSgnNjWF1pSXLEHFb+2iirGtIXGj9cQqqU2
VEN24mWUsY5/y+ZJ1kTE12bjHZyirOzM7tOsjUuRdKpbGY6XbIKO2Q6ekT0CaV9YtWyOP+9MOQ7W
xremgk+d2Ol9qdRvf9R3G01Nd0Yfs5txZRhsvMeHYcueHk3H6/u8F9u+uEWV42CDZV8UYb7sGDcu
dyXn8cl4mhag5+uMddou+RHoTHhz4PapOI+EKumBHf3FI9M8QeSuJXLJ2c59r+DYDI2tXF8aznbT
M/FK09lRgawHBaJR0wElQ62PVwfhcHpSUCTbaWF/hGAi4+qqeES7bWgzOoqLoBCycafPemsL0swa
g2feXgKDGqjnIWSdE61Z4znF0HGXHwV/xWg/vq2KGK1RjJSGGOwaZruDCX8RX5UlIwmDRxsxsucI
ZwgXJcuq8DM32karBx8Z5Yj5pMNkHqToMyu4kO0TKMddFtM9Ky0X7K9JryKk4Ln1Ji5ycShrVA6V
THo701rwrlcsXSP2AgqE3aNG8IrQgyQEpjzFG29tbU1WBpq5n8dtF/1wWAskLLbPvpjtYAX1LSjH
lZ5lYHSJpZ09nr4A64/2/5nZgp3f1X8JYF6FolxLleGA3HOO8QqJqd5ohqTM9Xy79aD+ohjzCiHu
XTvvC6t2/q4cmW3SghDS1LBuaNcmCrK19mtO9C1kBJ2kh3cHdaEobKUmNn+PU6PdofP0NF2xfaQ9
a9tphNQ6hKiB0sLcDQAWkLJVscu216U8Qj1d0Y0J/h+xaCbJ+7hqGdHoRc/12jkOZhcdB4reWTGw
PicuJoTx9qtlDQ4ZHvZBbwqkXjozZDl2k/WRgCjVpgDE4FakEyBGisl5Qe+DeCqGKqE+cxfLfwdC
U0vRCHPGpjkUPXSVWWMIOVgNyEQZnzO9WhPenm04onN71ePPr0YQqFwustMlFwKqQJuH72c7VrND
+0BAkdns63quvKAKxZY1UzQ3Md5NgAXqX2RMEP3LI8UOu+00XLapZ9TH1D/OdhoYAiHZbyzgjDST
gfjk6Q689X+dnwJs1FmeUgwd/A0D8Ozl5NNbyxH8zq4eYUvFcGbxBgmYWcE3N/MVDbx+eoRGH8Vt
cbVmoEk+cG0HG7SnTsQsJifrP+MNcFHIPptn7kPdQyydQ66DJG8ROeAKqhzAe5irZpCN7FcO1zB8
73hNYupryXPCiW6G3ehtwfJqTH4ehZ58ldOGsoeSize5G6haQuOjKMTQSayYDH7qxv+laswhHWQn
64yIhKRHZ7izHJZnxxDjYhuz07qde4lYUxhw/T/iplY2sKloEcUKGs9Rhq6MraalvWItMXB0nFTO
ODHm3vYxJZwtjQq54Y7Q09rMU+nOBG0xsPKeishvjI1G4etLXl/n4jja75VqPRW28lv3LJxACvw5
YqXt1hQyFxs0H/HYa6L/hXyWWfA6JDcdH6zZjSyyt4iCHw2aU3185PG8ht7Bp9WXcu5GL+4o1LXD
W7AkisA37As9dWqtNt4kO272XVu3ldix+6xEidxM2Dur2BiXHe+wKQ+m00drtFoKkHuf61BSVfqe
exFnoOEkUyXFifmygNsLupvXwun2c2prqzV7H25xGLtd/yDgnv/s6z55Ck32GBf0iM10AmZ9Cqxt
nI05l+3c/q7MOZtWvx0yI4NNSdLcW5xg0QEQdfZPZ5UndevjIe9IuxoPWIYUE0j6yxXLXXo2lKLf
/aSsvJIy7DMbHqBgcGF8ZhC8O9yTjETJRZQcHBK6u1Rtls/BTwhgGC+9dUak9NzFGO1hJJG9QDs3
vlk6ykxh/k+/qOeywQBv32omNi5vaCqypFUZ0hRUrGPDtWAWPKc2WuZmDBFnFzfTyDR0bsrtpa0A
2M6fwZvoBEsQvBZLNYnjvlrSFCAGfquWHsuNccGXEflem6fYvzb0PAUwtizj+YozMRmRazCEQPmR
U4DoYt1ZWb+TwS6AAM1tbELaUXFz6pHesBz5iGVQnf582jU98/G4BqMsJnh/KvWDLjADjn/Nvuxg
gTk2YpXNdHbGGMgyr+IbNbxzklFsM6qHYJ6VL/kc+xusavs2tilMNGvnuGrDmvc/O1o0fzVgPvOE
Rjx8G1Dq/1yaUxdf38EEH0oZaHxYgDyeC9EDFO80e0kw6wW6081NAMbyOUl5gLSZHgtN/69OsyCW
oyqHZwDVIKdwSLTPg2UME2oH+Zrr0IDReIJ/SgpQ2Vs8cOMu/i6DVP7pFuzAberB0/sGnCCtigX2
WcaCh3rsTibh0OupMtDpBjb41o0Qr9kXkh7vqYkwrUTObfqhfMCIeQVBh2OBF9qKXvypiw+qeyUP
mKb1GUpc078+D0oz9cSvbTP+/uU6CrmzTPf788V5XK0Rrwr8cc1/Iv8nNSa30LzTRPOdIUXHQRyw
pBp2LOfxmKUMm3RsqBd8opNxbMtHdUX6Kh0Jsf7XyXRexuwXHZYLzHP1ZSKhTvInNEghv/6gRdgn
XPng6JQqcfjOR8DmwoVtX8ULG4IYR30PiNs2EvOb386eRVycTp0qKTxs27QCBb9/YBQIfp1SM+Sn
LLG0G+ylA8774d+NXFb0PPkF3DF5zRkx/gY9e6JtQzW4b/3UesXFJ7QX6SY8pVU0dO24s/f+rcM3
BP80tYMN8oAHCEHhD/FK0miJPeLHElthH6d5plrR+7HKMcn5wa0pMrbxAeU1/OBDS7pjQQrj60gb
qSR8pgTYsODLyuW5vcckUaA+GKYpY+y708X8JqjtgJ8ORCfbJdaxvvEjBZ0kH1IhSTQuZggs63Cv
nF3NHZJ4xdg+NvD1frNVU4GYvuC478gA9RZ9uVcv+rORM0/rSOcMOY4/fMlitGF3x3tgV42ORIFO
GPkWmEMYGGPk+Dakve3vgjVF1v61+Xmg8WGqYIxtKXnInjEIA6P+E1ADzSUtA1uAjV3LFHm6V3Ke
Ywp0A7p7NgfosE/R1WiU3FLmjAXB+XAbzfJYTb9HFp0MorINMHF6HNdHgHKL4h2hzFQoQ7Te2KBn
r5nG7eLOyzm0tQ5Aq/7hb73pD/7oI98XJTdsAKx5urG2TEQFPqJOvQwu9kq7/2VxqJ9qcNVv6fIf
od1crC1CaJsqxyX9hbIWX9a2Uo6xJJ57o0MslwSBpRUcOCPMNJYpIhs0FSMvWkRZGVzOpI/dYPxM
/sl+mqkpYxmDgkRl2RPEtLZeZwjiw0w2deTY03YC8NKExsw/PVz9o3FgQn+GZUlWpAcjeD7e+nUI
lv8OLnosYpIC6KmD9z7mM5ibmouBt+b4gRzYb4qexNyJlKctKpVfg/s9CdQ3VPifm2Fn0da/FRt/
481gqu9R0iGzOcb0try/YTucI7t9Tnay6OcasORZGCX8P3zDPniXWqyaTXSPQNhXh0/MPe+Cxq3U
Rl0n81/VxY/o90aGCIkOvOlR6lp3YNbM2ArsYB9dtRO7P7x5URAQ9EBJteOWkdrRSPXfmtVQsQqu
tY07o+HXmTpfQUgHiTfobeL7juh5b6FenWX6BF4HuajZgS8v3NJkU1n8LaosLqUw7W++OHShmevW
RLTbeTpoz+Ika5AWjcJxlbVShm7Rwhd+XJAJUC9Uf0dqx674U/PdXO5sHqAMh0L4H4TDk8aCRn+V
3mc/Ipp65OaKGpZjX8vBaM2iRxq13RdxkB9vp4frJvw6dtPQY0kyv6M96heGPQFfXKh1KBtqpK1j
l90BKoI00bpdF9ISTYMwkGgNoroUzuHeli+NrcpoXqzoK8OA3/BDnUjzgii3UBqf6bunzDR36OTU
eFy5C0CMgDn16wbTVD4jB0UXTcLhJlOCL1Mv3rezFoG3tmB5g9czaSikFjTCLPTfSYW6OzCkzfIn
2SGcC+e83cP/x7//3zK6diUr8HB5X+uh0f94M0ibEn23TqqKG95M2cFEQQtCMhimsPUgMg43q6tk
9k41P+m+EzluBXeITW8TB+MlD9J60C9ZZjIZyoeqI3ZEPK2ebMPz0MypXXhamfPM6LXNvdeqCfeG
L992+Pl7aUJ/CaH16IValndw9Y/meVREwteBDcvAphZDTEUji4bkomGPGfAHZMNdj4eMwIfq/aoX
V2BA156kPySTQD6yqk0Y/BsgthL+2KiVGSVNm34tX5iyVXzpnTCuaWlBxd4VSMaVSKkortlXx/Gi
5J5BxJgQI/yMpIDqEhBftgpQ76OF1JoTkY+jrpjq8eFZhDsUvuPyLEb/xw7WAuuKDQldu/OathwK
fTqidpGeRNcNX3GntM9Tcjp3LLQFRmrqMNZl+Ke8rPjYB4E9aU9Fjiis3FN5yRymROzn4Cz6M1Ba
86/MN/EAMpa8wm4TBsRSmARJlz9xAplUC/5YzvSsBw6WF9R3jkx41DbXR2UMdI/T8DPJCy0SMoFf
wckye6s/8jQxaUa/ziZL+ZSnn8BslYMB96X/14GuFrwCKViPW49D+hBt8cIMRNUYhzMN7GKgTvMH
j7ur3uoA7OvMZxy5gn5CHdc6KnGFeram/5/zNE4J8x4heQaHKqbeA/IvvF4o6Do+UTmyBaSfEMI7
PiFWyKWrV5q99Ki+lghmsT/v/RCCbruyShnR/HjG3fdFvv5PHhlgq35ZkG53BwBuQ4LQutQ4NpXE
sEApBCGllW2UxHY0zTvE4YbAisagff7wYHwzvBI/h/dtyiJCn6bQbpcjMXxq3Ka1mZzAddJhRfro
NM+vzlIbCapf/53PnC6SmeYAWT/W1pHa9abpDGmHFxqo4u/WvbKi4w6ptCFX/lwmctxIEV6J78KQ
uR4HXrJ9hpsCXtzzIvt0YUCw5hFjquK27anffIRkVcpQE+NUymXqMrmR4CAvCC4ZOH4607DNuZdb
7Nr+ls5lEkjSFxA+qFRUeh+wCB7T16JeUEzY2GKQwllJN8zkSzf0vY8HY7FPy8cMp5zCj+DQddU7
eIOrJmov/3408Aw2f2jJP7rruFLtpxhz7JvzlDLtuk/Ue/ac9HJ3LF1UpZ/AwyDaM/37PEEAXrel
7zIPk0L4UEIT24IwixFeM0V2WRrgX7gkD2P64KzFfqQkJZyjN6CKD7c1Spmm2cxjF1ZPLVyLonHD
3lWjBfjUmP7gCbBUfR954eDAf3cPdeQWL84h7ipQNFyUya8im0Rpx3couXYGsQLLyJd+6g+PxFR3
RTTM7J8B9skcBPR3C5hCkufc51bDOV9L3+/MEPPK6Ft23abAH2HBXj2mJV01Sq18g2wwNMN92/Vl
z8roQ3d9VAUED4Nr1URBUihtLu9YwyQS4qDWi/XcFfIJnglLGh8QmKo/JC59jO2/CUO7E7OXlSYa
8GQqP4S+wBfA6uO6JmxEMfaRdxas6mZDRDIr6LrnBBJyCyMEZWGe+cX7Dpjuuqa1URTBgC35kdTG
wFnv17lrPlcCskUm2jdilYAqFTzG39lBkR0XymADbvI0Kz8hw1QPY3P6H4SDDEM1dwnBE7Lb0u41
BWdJUa8dA5LEbzMhXixi4ewLheh4Oal43BUFEraYFoT2v+3d1XmUnGEP/Du6MFrHT/a2hXqb0M6C
3w8gi2MZ4NFFVukdRfo1zt0P3zLxnzq6j3pLMztcr43ytAAhUS2zHih1weKTe0ek9jAR33VaWcl2
i/HcXMV6XNCbZwaDfySMKa2Ro3cn8WI3avMukfFj862YOoeCrm7Kam14hPNl2md68igJVaP9EuoV
oRgDxFKWqVx9kvyjIAGtNBlLUaXO3gzOn6DwAOO99ZQmtRnlaG4VaDX2ZZ+1VeltlXvF+g9BiCu/
A45SXrg+8wkAaW8/4Vy30aAnIlviyjJysi0PIUwT2LVLYn0GHO768g5Kz8wxxjktK1iif6ovIvoF
QsGB9y+GbcWascb/32/rnPhRbrtv4Ti0L8JDLYd+Y1jGlPn5hOHKsi2/B0vBWETaCpa1YHrOMZTj
YgsYeUfuy6+VOO9h5X5n9cQTa/orcwQeLLmriA8lpuR8s7BMjVEKH6NI3fO3iMI060t1CU/+znqE
48FtA6KkUbTAo/Fylwi0bACl0+vqNPqq9iq22TOz6R54Fg3OMVSAPYXH41mV1wGPhawkB2VbEvdO
hhR+auWoCyOMiMnBU6MyVFm5LhlZcN9ACxwitZ0B77eJ5sSioazIZULUrmnORGyE1iOJKDeKz5l2
FGYVIz5PGoC9q6bVeEOhmLRM4jYL8fVRnIKJyLc1dDO0K/6UkyLLOKCAWzsnATt/u8hSUrajiKrn
vznh0mOq/o1LFAsGdcArXwZZKDVZ5LAg+L9kDUL7XCC7L+4Onre+CCmGGPM/B7TMcGaWTp0u2hF8
7FadkeK4DfWxyCR8PgPgncMVIp/Y0VDiy9MRkgdsdVZg/zSqiGIcIW9nrvEaG6027eyVT+YBhnZv
pOtTWKSfZPJPcQem8sHvHjf1EwwOVZQVZtuZ7yJ5ORNVhtfooMSQHM0pVN762uwIJn6HJ8oYmdNL
8h/SRjwK3TAGTxyHfdSUkfDMtIwf0fzrstUejxRQsYP5pgv7j5Ao+uB3sQgZjZXxhv1FP+k5sNza
FNWjLiIroU8/cqY7IobakPc67HA6NdDQDRLwfEpguCLllz4HYPuOk3VLh6iURoLhP9eidAJvMRSp
PofQBN7Ib/8Sdpq4vGluQyo7yhSch51Niq51UmvVbfPf7f3urNQR4XH+ZRsdByJoMH8A2fnZLPcj
/ADgMzPeniIr78OLz0o1eZW6XpU4UmXgWi1vPUINprx34KZmXca6+64IR6Aimo60B9Xf84wT9ukq
fSyXIRuCOWNDypa4heyMcLifbGVhI5Hrt0ZzMOSB0trsbGFYeTLY+lwaE26i/iBqZP3JH5dFv7n4
wFsbszLB/MXvryBWXRTzj3uf5CCyyWqAqUoECwtEsyXnO3ca4zOQ9s5a/fRro5BgK2qR4EcZWH08
2kHm0jxMnvejXVDbYKil2oyetbV4aBw+bDh2zqMYFjNqfGg/xZl7/T6B6p3FrCtkoTajjswMK4x9
adyqNA+oH5xye8pKbimhdQSb1RVXN6lgFsTXdKkN0eTPR3BkXkFZwPGQUKSmNQtsdL+fz05PKYle
jTLC/ShuZKYyBpZz70Np1iDUyrNaiYitLmnY4dmI/bk9GFU2L3VIw0vWCCux4AZCcVzUg9OCsr7i
8YuT2cReDKZjRwJX5oAcpJ08RRxQAOpv1ikQIuaZtPLRBddtspDgJUmSUmXlUJRt4ESE2O4WwEx9
so9QADlzs7EYZ5SKDkFBt6xfJGXoxbttT3TsTL/A62n7l2JizDKU1YUQcZohQuWRRsSsTUi9TSXa
PyjrrLoUQ6pCugwnL2e1W6RxsBHRTVU/WTjGeuue5cqsEZUu8hFSlUQidkdG7aT10UjtOran6E20
G58gE18uhpxPRS2lf2mTp5lM+GudOZf0iOD9buxYurVfpYKKUA8Z63DZDRcBCCnNy9D+lbYL58/j
Ctx2Xc/daXjrrRVEXqLDIm/TJDPgSfd8Ac/lhlcab2888MC5/h8Zkyb+tQ5Bv3ccsM1UxNoiEk0l
VUC7gvUvtNpVbi5za50T4UV/9Q+SsGWjrqE04Ucec9FrdgMpESD6Mn9yDCSFMIUuM8asYeG0K5EF
rgIVkEP7DJuK0Chbvdh8YNZ6cFa2s36MLk7qH99wGvuVDZXWKv/vZmMexARbSevdTJAGBQqDXnQY
kqx0RGm2b+C1Zl4A3pWb6vIUTThXDfmEFGdaE0fDNVr2cbdbvLMbJZEmlVMSrj5/RHdZXfiKzV45
wD9ExpCvTcJDN0OPm6xofG3bRKtSsOuYUeeo1aMp0hMkhMyJ54QIkqkg21scki4ZLzNtY0LMyZwD
To0hIOw5vG812iu98XGrg8rHNt9cwJ8dl/rn0QzSxHBkDWnvKtPlGGWXPcW6LcMHAvmiUYHf9hxL
uctTFt/FhM1Rai3MvouJ/X3mk/jdNyB1B9I1nk6OJpIe7p0ER38RHQm/DqHjLMfeMV0wFteilYGw
V/KTYa10mMmrYtl3c/Cg6S4zycy9EtxtRijDiIzEt3kXz/hbfazemc63jwO4EE6CLJzemC0FKzzZ
3a4hVDQbapmseT7TL2j/+BHLz6bS5cz8rhp1m6uXlJ4N4hu3bfAjAUzjpezUo3HOkLlfkm1sL66J
AQT/0u068rx6QckH4vTieZcHhyYN3fUNK1Cy7xxURns6R913zGO0FykBiRF9OH9hAau2iJP29sdZ
tLKMmnCJMwy0DrPwp/icTWItDZ0fzL/C2pWAmKVNjufsSOntJNPMXuYsPhfsvxYcsBJWtIASY8xC
TUsOV0ErhOOZ8C31LEbV2jDdj5WtJ1HChRhxKoX9L6mtn/sZnh1CQugjKr5CrlipClGz74MUwiO2
7yh2WlshmdZY3EVZtCLXuQz7cny+nLal2Ft2Tg7JnFfdd65sasToQ4fUNq285968EdhCXkwL3wNK
/st+E+G8MHlKLU63lrI5rHaMxO68AuZIbfhUCrR4W/mXy3avUBQWbOSPKHtMGp6/0GrRUXlEhaFU
dQ7LOGGOqlV2fVKPk4B4lbfAmJPEdmPrrBFRtwXvVKSi/e8NWthQ/TzH7tFBEums1YkTq5IgQIS2
gVgsPUoitmvWEA3XXa3y4YFPM1grfpdo8/+HYJGc8XLDCvnAvaLyGlpfcs/QNw/SE/J9Dl6H54cK
3U3CdLm2cW5zAYNBDs3BmFUE7dKObQw0/Q1LIy7DQSEh/vhjrkmD/2ePoLdS+I0nos6NMgei2BUc
BNVn99tQ51Pbq0nexuGUQoFUp+DSqKnGyctkxVXCiMRL6lxtDfVrRkD2jFIQLirS4RpMs1aaCpCB
GgOlYjs9P8TkCSYt9x6GNhMFAhJjBEK55oAVcTs1GLg09DICFMZM+5lrUck7tJlv9xVvoKqrsS9B
7lyo+m780XiLJbggaGgVge9g/9lu8Yvk4zRAQEF0XQKuFcX7V+roROmIrX1MYDgu2eHzgOAyEu7F
XqZv/2v4tmRJli9eDkOcwkxKsZ5hl+VhxraceEm2Cyq9C5Yly1XitOqt67uxOG/IWvvVgSqrvKMu
X/M3YZHBt0iT/OBd+8b++U5HVMlVOdVjbROftrMdHUCKEXINKq/s0Tiou4A+u1Eu2sSVt2mXOgi8
yPVAzOmZZc7B3OYkerAc+8WtAY/vD2n7zasqgtLD7y6Fbj8MyIoy4tJn8qJ7qiiXYF69JdILt5H+
cfe9GfIdan4xyUc2adT64MghvciCXnI2tzBCt2x8mzvopNy1ZDoHnTGunizP9DWIj7X1A2IYs4Ww
eOS3vjYRbos39dSTVrYXXYv5Zt2LZYeVicgqUOQ18WTWzU22y0TRUC2o8hWaK/3BGhU+RSK3oVlW
VJemTwMTShUBFHAAB6GW8ZYFSWi20ErchMhKrgTsuUh0xnzPr4Jhgn4+aXqePA3Xp65Y4FeKw3Iv
CdeBrTgeHWpZvSvlC/Z6e19/DSYSz0RigPWmjdyr1qdaiSwsCUoQ906Y903hw/6vAHP9YjgIMw0U
/INzNdu5vgNjE6b2Co+tTtEOO2UC3qK2lUODRqGK4L8t4RAuGMKzHKsXxl5KEl49ICy9cibHbWZi
J0yDim2Tawt2RSvtBpD1wMVDn/MzRKwMRC/glLrP0OlbdTEognHwgEkv6dgpaqHP0t7R2gU4nR1t
psYD7PmD+iDaC/xofoNwNItBuwFFPzYNP7Bx01Dgdqas9iSBj15+8pjsrIfUJNoTVnoiWCWDrpNP
f58u5+UOULs1pTYHajK8avmocRtYWT/Oj0d8s9Pssh05fuBRKE34xOdHBxUK8nyOqTgOS5dpfasn
NEpamrPOOvcv/pm+RFWCJ1ySwMr/jt0M6iZ8dzCpEpSOBp9iqWDDiLC3HYy/uWQyU1R0W2DNKaNo
tRLwYl+9nYkq6GTOVqem9idFSj5aDt6NzTcoCSskPaY6g1+03hj0WBloxXjzpz8K4hQaqtNz5UDy
wGYAbt0Hu3HlgqYmk25ERZ+fySJ0kBJMwSkcs/bl9/cNX2GIEdWnKcm2yqsFMIezwBAUj3Wtb4pL
spTWujyQ+/A8FyxN5zWG04smomCa4zojmT/vQ0Ik/r98cQD+81YorR1t1cbJKUaM6OhZAMuCb/+2
80SglnLFhIQLMFEAcZA/7qaK/mezBaMt1bVynaHxM21K6652liKpw6fJe2sDscKbvkZRMB5OXyNM
wp5c3xVN5Gslnd+LbLEG0Vy++I0JEYT6Phpqlne9nXrdT6DYy7keFbzRSrDpQDGGRfDTFjxjEgP6
1lSgs1yOOJ5bqPd/UNaymG0TMlLUZJbjUP7+AIvEG/7eLPGIWZSdtFCQh3vpm9X1syEy1P/nSxAg
Q61VAhTpPeAJNrw/Tdyic1txJLKPTI8J4JRNmaSMEmfm9LWkChN0oWVBBfWg1rSdxxjT3V+6WK9b
kdDAHBW4gKBuLJYbK2LGuTYQxp1zdBRVU0o6XTQcfyrMefj+38kwaw7UNrrva4pyVQa5DCJ0IELK
i/7+zI/NNs/DUlRmP0rTz/M+TK/WXEjoTJI0FgJvAK2Q/niAsmLiyCx28Sa6optduZkIfsvqPrK9
R7iwSr5TrLnVw5HGp5GLB1/7QvUdk+nBB9m1pW+xzyfqwhvLOQhxXL6G8M6knI9nVf9ZPB7TzJgF
wPHCI5iSRkZW4cgStYucf8nVUK+R6ILsfpP+qWnq5BAr420UR3lXQ3y+AcVF426BuvDWcGLlyj38
WYrKJi2tx3HfTk54RJSOMfqO1d06YHB3UDcuulBumFHJ/LuJA6LnlkxAI5LNTI4PdyFmC5/lLaxx
3ukdC38FQOGBsy+GQnKaxmfb2KEuGB78JPQ2W1oE3MZp3/XxatIdaK4kL3F/mwRu0hq0eK6Tko8r
PqFmfRomzj9mSdDy34SE8IdxR8rs2swCC8VXap/pPva/6X8o0lDfcb8hrtbVZntXOiUtUmCCGhAJ
cP0BHb/j8Q1LbUKRZM684k1FdMsoniYUclkryv9dSEypV7y4T2Te6UtQttmtSY+j0ZjUu578oDDw
hdoPNd4MYGy0ktlAv7Bw/FJQLvV00JpYiSFJ6KbTgJpCY/KneMxeEzNyyZZaYsfnPUcAhd1+foS8
JKomyNOXWgjfCeSYUHXRtlJ3JAACiZ3Z3XtsO61BH87soFCMZF1owGlZJyyhjx2Zd7076yTwabhh
FdbkdYYdMQdxed7s+GcJ85FVoJVg7euQnfh43ikFovohofJkD4oYrxoW/z/rkVEmZvOghBRyMOlE
0460caNKem0+N0RoFbpYjiSe3wHpZNCWNpLdPVfm2m84UfKNMu+nFFTxfx5hw80BUkJ5rTPHSlOk
8uHss/GGYHQ1TyzVVhLBWYq5eFvPxAMGWo4DndVNiFKLVA8Og34vMu3zRhZ3KjxWm9nVcztzq3a0
qselwd9BNZTRWMb8iEHOhKha4P1f8MLB4W6NOh10ATEVUgCufUlHddCsQZ9XlnpT5IFKYs6a1p4r
Hz/IdjhblNloXtPqT3NgOX1nkdfMBRgUCxvglIi8owMm67MsxYyflizMNEMpZ0Tywj3eQaJ3zMoD
0vcLDjmwdna9Uc1BhMW1SWTI/0HFXLQR5UW+YBc0Abl6qEQH8PFKkP+GxoeO0AgYcdRWUcFps+KC
UIVLjElla6WT3hqV0nk/lg+A1DxnFFkyk4KNG3joH3L4wm7FAapCO5DTTsj1aoEBHTKWCQ0QtUHo
FoM5MLGMHceBXGMJQgpPuMx9/u45UQpW39HUTjIYEAmg2YaVEULUhhvZc7oIDVD2ogN8f95kRBf2
B40Gdjw5gr5JbLzlPwLr4QolGBfBtu1d42cl4MCG5idU2sCx2hoxjXqCfG3FZQD2/40sq+Z19gD+
8Kr7AyVitfDjrBN0U0POnBv87ZtGdtNEpxYWegRTQzY6npEHb/BwlkJkienbMJsx+a79yNOuS6Mv
Li97m6lvW0ou6Tt9JzpITGpVSvACTdX/H25G8y52dXjFIxof+qxj81FcUprXO0dSCoUSxKSCgNuk
Ooe/Wc18VO5hU6cltex+C7K33GKjorJ1J70FYUwWPrVzFV2NVtwJ1xNhSI6v8NHGN+ygb2K1SXo7
LxkBc04jc776Ye+cpZnzCOXnIy7152H9g5cY0RubHlizKptmxweLuu5nrGffw1ZRT5JfrjCgON/h
4TOymUM+FWk5rcSTKG1efDbagkgl0ywETTAbUpy37kR5FestyXLCHa11SxveRBcwfT4d+s83WdJE
kKiPHqyfCCywNSpCfyF6preu0Uft2OYDKo35F3w4kBYlJ073we4tiKU/qO2wxiusHHXX0XrPuvsL
/FLPYec5dlfqbP+n/bSAuBsJ9FpaOIvOhqQynpvk0LtIAPxkIjdTWs/fAUWi+9wvFBCWTtQDwoSM
5/oAmXJw22E1WO7x5t4NmODLhq4sDvvjq6CYyLq5+ahAxarQIu5WOS0c2uKJmK1CHw02zmXLYml3
IhnXlzGOjL3oszCT+13seIiJVLZkMxF6g8dQnSWSlInQ+BP/l5rXQX0lAnEk5/uIU8pBTtl+GL1O
MlPbNBROW1qAkwXGbCyYNcT4+wjHpU2yVkj36urxZxqCnY7pzoCSJlgdxXwp58HOveMKerAvE11p
FbRR0ogyxdDrv5B86cbytCFob5uir3gbKNF7rVPYftijz8pxFR/XfctVnOft5podXmB9QqBKuSIE
42ABjcySQXCupYhpUa46Sz/MgW23JYE0EinNF9rJiYdwC5EV5UWHJEdPFYCcUC/qZm7bBYR3oGKK
PqJl5qmK55vOlRwKJLlPxxgybMTdIJ0Y2yrVUUaxEqP6GZIf4U0fk1WpAbYmOz+f3kuQnmA1tO1z
k4Wi+5xGAJi1ctbL76KVDU5DMRkzJLXUGREIlkgwG9AloszLYsnnhGOO6w3SxFganalnUJFUL8+i
YI8gKwVZzD3cKUSxIHvc91wm3SIdZwao6IK2EbDeN7oikmufsc4B+KwNi2zoGXg5vgfwlWb6dphM
JDp16BYdTPfKxcLd436fXngNjN5jMhBlw4+Dv4U+26105rAJgbe7WEONvkUeq58WtA9ZEVYKOCea
+214TUiTKKls7dHutiLDurz1w2Z+1I6O73GdXz+upzDV2oGamFb8Gk/gXkfTx9vxzneDdvQM9fH1
dVtPb2ORIiTLy+B6pBkvklowgJh134v5Yk5XkISQeHQaH1VNuYN5S/8ICL869NbZL1hw+Deg97cj
X6PM7lbbf21ccLbclHkAC3WXlWW7WnzzqqnVQ5dDkWxEJtjV7sEGEt1AeVV7f5c9Hyn9bwEeCRJ0
GZ5DUH+fzj+aZHGoOwGdjOOP4S5DGJnZ5tz+XOSH1rZDiJ7t6jv1Hn0yZXpZpPpdrVjvlYgqPmKt
O0+64QTQDlvBjGxQseF0Ek/4Tiqcu0lSd6aSvxzPOwj1+VxAtRj8Ld2WlKYwxw0MWL9jvQLYhbft
/X0/CiWkj/nbqGVR/OG5mhd0gfjoV10UGBPoVDBoW6peSZn21JHwUP7SznIZB2TOPja3X3jJTucF
LzJYUq7UMPbNbtED38EtHMkv6bcm8iHJkkbEfIdKV2/KmqwzVNKHT66pSUO3lQmsxz7g4MOCLF4R
P9qCKStitcn7sjIHiguAHmRbOaVHQ74HWT47UPpb683C8XVlO9zc92/QMNYfwDTc3kwHQrUfqNcH
+mExpYjICQfuP4x4/YmxxJLO4wDER/er/LQbpnfQUnoG0gxhmbL27EjUWgZ3AJTaOWje2WKBF2gD
yAh2QOcTXWnAWg/ReUNvozNHVkhZ7JyaJisB/p8/XGbSfgWq59V2fr5IjB1LXT4MyG2J+vgOoabW
MPgYtxBNcg2Z73zFZrmCM1S6sqwHnomyOhyu/lYYT+d5ugZVEVnJdyynLep0POZTETGUZ9dVAk/I
Mws7Ru7X1OmVPsp8GmRhK43qwOga+3EsMSKTkR0vzjHAXK+wZvp+VSpGP0RLo/5K5fFRZB+zp1Rx
gShwRoiNh/srvEt38Lg+2WAhgyvbPAZFTgUJPSoldOFXWIXkFy8hk2M5eFKpz+WulnH6L3epiwZp
62w/3Ny4cTb1r5J+v4lGRFsGvvrNrsJ3qwvfkQSoSJ0BGppSX4Tyfk45Y67BYEhFrcgc28bAlKwa
XtKvt3YSMPuGvhPYPQggK38Y+PBqYZwaKOiMPexPSw07XwNEEQCCgRfwbvP24UJxe5joRyAuJWsn
2rmm5lHCPliW0EyQpW2vUb0rTGP9nyDlU7jE8vsPCAT9li+Ff5ABuGD4zjRPVnoGPofFgR0lFqHs
UY+rMduZZES+qRipdhhPUcsmqDVCy4PoURrB7KJWH8zmNuZ2mVgyydBj0PpdWE5DfaQdnJX2IpIy
Nstt475vFToO/AyRF3sCdwPTn1/7zFJSnWlqw+Ew4rOWCDwsP00d0LUTePv2gqFMnq5RIU2E5XEF
rnwRkH03sbHBSrpqT4G1d8+MS8NFSuDlQVZ2RyKj4GEBAyPAdTlbMsqgKzCyeEX5nVZxH7jYoasS
sG4NQLELBPC/kFES8RqP5lVvE7yavg5u1DRE1G8fB8Usl3sXBMx2VJLjYi7Lbil85O4s9uLr5Y12
hXj2MweJ2tc6kY6ReIL2x/ZUhCfHWbFn+vcOtZ0Jfw4Yccxmkbwp/gFsdtqf0Q+aOvfXyUOXhZAZ
sgDALH7tvZqe32MPAvwvDV2guVN+blpY66cDyXFDII/5cOIi+FhgmPAwPc6XQWGIRwd7znhqx1MK
FMsvc7fY4F48ziEaf4y+wF0NYU9bGCIG2dxXMIvTgMzYh8/hjYMsOuWIiAQw1Y0NuN8y/C/u1DFv
EkREljkfvu5xmfBq4o5DNaVp2OzJCpUircCY7YKgRw3bDxcoNFeEwiNugfJN2cPFlapaE9R8xDbb
9iioZ95QtdKlwIrVW15AjLx7etWhRsBUnffy3DAYP8v92gDhM8Onbrvv+myYy3+mFtsSOTPVmtCA
HG6sQbMefXkbd7hwvJTsZvA2DfqiqPZgpWIRGNyIdfL15jOwvzdVINL2unnhl6N58mow27j1+GRi
+g/YeWiWah+VpnQLLBYoZRuVuFjP371Aou1zjRqkCDyhwMM36X+tHRyix3d1YxMC9tdZkyInpLRP
SzeOxaez9eE8eLvCH5aigNyjz9o/lST8eHyTLiwfPUtwyPDOqbo5OFOKqt8GBVJxV/Itsa4FN6Yh
oAqtR25X6RQI+8btBBQAxAS2fjXtbZE7L0TzwIkudiFeeiS45cNn4UxdwpNCHRBWqD5vJDLbEfw8
ojHkBfp/2rI3FN6zS5D2CgMZPepU+pFBnhLz+lzc186UO3OzP1m01ZYT8uR74yHlIOg4EJRBoyED
wwxaW53Kg87lScutq/VhOXJleLeqR9fOgVIf0z5FF8g0RDKMNc7M0FjAxjWrlgk869Dy0la0P5rP
7dnYsDUQaoWj2Md+hu75kCYA3JVlMOEE1wj+1G0a69clWgCQU2SDGqyV8Biobv+k0HZwZKNPgSOP
s7o9D3aZYX7eEw3htdO1/si4ZYKAgygjw462iYgSZAiFBXxUKZ9RCuiY6XeVSDWnOAp+IzL2EuDn
hJ2zr/OOptZxGYvw3mcwtdiCKm+IuZpe5bSQf4DQSRuchYzDN+ZnYfXh0KNZQ+JP+kRIu1TepWHd
nijlaqMiVFhPiXsa6MAS5xrSuFs7ScihEaD7bNo1FCAdCDh09vhIngeXH3jOeRqDPt4yAwz5VsiB
4UBLL80rsxigjiQnQxuEUCDmgFx+VNNojh8SQCC3/I/HkqEuoml6Ny2shu5ADyRRST9U8PYPoYsL
3BG6V8ZGPQ/fiuI/ci1A8Y3Xk5wMykhTegFyZ8zo5MdkaJ5nwdeDYaZG3bV/nyxe6LlmJwBzgvET
c/iXWBnJLsu4hIBnamg16JsSttHJm5LZ77vjdFqsC7dlWLrsasIxfz7q5dtLV2a84x3ppuByHQ+v
VknTWJsDUhgzXyxxPHCuyA2VK13MmW77ha8UVaiGZ6aMOhv3w+PhLbirIXH6Hw2g3+DurWLWMkPJ
K+RGtUSMMW5RRw05DZRVljKvruQw6KFyJ/OXIFuSXp4ejrvjglUVEv6KttkjXU9ns3OsrznP08Qs
65XhYNcykAwa71EQjoRvPVEfSpVd5X56M+trcSyjECs59OaHMz6LVVAKVauDPctNjYW4MVcTt5lm
2qezov8N53AvDkANrHv+z+ckzDsTa3SXHSCHbZwZWLKmH6pipvJNzQEleecS63Hz+WtW4xJgsJPo
+Fu40YhJLwr+gEGqUE/yRp7f1atLscc7k8JetVjNsoyUpCRApb1N8+ezPsmfPrlzbYpdrrCy0YYO
6CK43i8r5wGNQA8H9ykm2d7muOJ4KuqU7eN1MvnJLDReow4zgS3GWAqLXrQFSJX5IQeLeP5rWMVA
bxg+apobg/ii1wLUvzvKeS/nbkYSgyQHzdQVBueVQYT69vrIAaPueF5+ryltAyin4Cmp3JaFpHcz
a8xYdUatQ49//IRzkFfhlsGAHhaobDilHpnSyHx6QaWfkiwgzbWWpeM07RtpuES/1tIwMQgid7BV
QBB7552711KXqtef9Bn/v1VhPOjEnK4CxMcohv9weZiPzkqYCeehINTPGeI9EEthenkEpOm9kx7b
/iy35eV0eAEgMdCa55LFK3DK15o/pvIYV7XKLSypTlT9Xm2AZ8oZmhkv58qoEN6/4/iUYUAg8dhL
N9OHNBsr8oAzaIbB+xiG2pc2XEID7tP2NZktlU8wdd1O9qh/dhgu8jB4eHLpx7OWXc9TekWQX7ri
9gPc1eNCDgshjbn8ejvOYG99ZcUIJa3PLnHx1MqrQfAa/+vz+LWDhc8tsuXxVOIoYkkg8yzjj3EA
LuL8wuiPDyGzb0MfjKysY70ykZqsoahPar3kU/Mo6y7auDVByoxH0BJdYa5ncfMnpMPUD8YjKkxX
fc5KzDaVr+5URzDYeiZCq5pK9Z+UtNKRh2IR5gXW1I5lGVgyBGgzOqDahPGTTFnG6dFl+LkfymCH
kJjRC9oM1cIaQAQbw6SMllvi111OBEy8V7AoP3vklZyaJIhIVgOQ5kK5ZNA07ds/lWIWzJa/6CD3
BYkJOEfLThWStEEMdSH2zLbIJLav+5uvcHKjCfHWXK2V9uz5VHvqT6n5v7heR4k/5jAOU3uftS9O
vdU9ozlt2hMF5J+QtZxL01VdwB+wx0mhNXzpYkFTRZGL9edN7J0t/7TFwyfMEqXYBKhU8luIncOi
wbhDzbgmescLTE62s0Zu7XziuFf78FxTFCbX/UNfPxTx+r3EtWaCOStkEmdXwtnjYrl4uI1vo1Vh
NqnifoW0ehnErGID3uL8G9uqEHTpGxEGuhOBM51U+jfNzFi9S03sdJqagImOXq+/Uy7iyWv4Dlks
iIK3i7e9vz4xbHtHcF0JyHp/I50E3Avnt+sAWoQWBDQpApkX7LQiWSWZZ72IR2A8UWW7Cr8gPQLf
wg2VxBbhdp6qwuuxR9h4+7TbT4Wb/5kHd5R8tsKDlTFmq162VfaSNgzdmkcFKY2xD7T/HstAvekU
tSttEAne7ei9u1Gws/MA6SkMlmMyCH10TcGbDCnBXsl/69+mxBFF7fiAkW5I+PjBfU06ld4QEdL1
tITmAoHH9E3kJHxKP5RlwL5pQPrH1imC/oxD/kCQJp832c/7qSvH1+kuIdsbmSR6ZAVopqnMiiI/
yJ4b0FeyOLItPhKPIaue/ZLKoX42zG26KL8kEGeF0JO6s2tB0GpExB2Jni4cr08/WolDf3JNCUF0
HoWDQ4aoyY4NfSvorQ8bFljChVcBZJfaMVbz0z1GQFzPuu6gj7KWuxHy66RaVCkiU9mp0GrVUgSh
DEF48hNPk9YmnwiY10PumBhv+D7Ru56vx2xmH/jiUGcre9l6tK5On4cfg39DbqTVzjoIO5dG7yYv
hz0hihx92EOf58bPoC08nL4CdmXF7e8OlGf6JFqM3FojfR6Ov59AkvldqMCVM4LWb2MlUGa0wdRW
JZelqYnD5LjHcl1mQr3W/JLDZenDkag2zDewPQ/K853ngsYya8KxkD+qrecrb93SM2PSBgJAPPkE
4dVVxwRJYOsZP5Fg/hjes2Dz1TDw5C/6Ksz5Mo5uArfg6bx0v8z2RuYnIv6HTuV3WDYIPTqOTCdO
s+8ik1EZJVypOWrwzZUOE1iTGyyPhPNDIKYfZplwKyjfaGuQMaCSNX5+p5ZB2Kcxh9mmD3LXvpBm
4A0aMay+o9YDeu+FCQu/sS8oRfWIyvhdWC0Kb8PjNo7UJM0HZY7LN5l9Jsmw67vmWdPBynXNeGAQ
OmmrNJ0lW9RV422zIAJdJhQRP5GEhdMf5oJI83U+fgpXRl52Gf31vjpCUeFiyPBsZe9R5JOr969x
ZhbzZWCryRzrf1x3JptlyGDqs0toACJlij0lls4hBRe1FAdRIMMQf6byT+1cYpx0q3o+NhY19nnf
dk+tWgGxmOQlXrGqJ8q9/rU9tLy+CI2W1d/tKLUMDqWsFjs70dNwVsCdF1Ci/lLMlBQWLLVTnSul
bEP+3fJPe6h0Q7UTAcx99uMdbTfb8Xl9Jkr+Qdl/JfVM0aJsQj9z9fGaUJgwslWqij6WRFyAHub+
L8PmbK3aEYtBCmeYKNWkD7+r7UGFTUGn34+yy2ZC4sza5WYvg5QJVmuztMnicKC30KYK9U/j8dRZ
JWRUZhdhQHU0LuhUiK2M7lTCSCh9R/uruUBIQ139cJsAyVY+lquLP40Yg3XckVMypErXMgcMSepq
Wy9Qff8Wc5FY2ITYaXt16Vb9Hr0hjPfsFLNuaWqg/FEONSPGMx9/Te1NYm3z5gEhM4pTZwKN3gZ8
9zwHsjHWy0ySciIRDQZ9w3HwpAmnFla6/eVtFjbiR0ec1GCsAGacZ89RPAu3k+a40/hOhTFpkl9s
C/cYLjBD/AhLR741bXY3WBx2O3WLjOam+OlZVTFO34ATLOFXz8qJUNZwtaevWBFgWDYQ262Xa0cR
n5bbc07po4NYhryrC5Pl4y03imrprAWkjuntMwdWe2jhlc9yrsL0KaPwaLjqUVhW4zh3q0nbaRzy
7gu8upgdcXoJvmjnb7z1GRSPC7KSCirXFYCkuOL/1j/pFkvYDFdSi+1WXozDKrtgHZgT43brnuW5
xRvbPripeHwqTekR70WxgB5eQu1CTccg509ljILkiDA4s39XrnCoCmQMDoDcaNEq8Hlrvn8iRBjk
3RpT54r72cZGDPPzGk/SctczP+kU3840IGFBCgP3q3WToZl/g9FaeEo62hHdoeiGoo6k4KnATAH4
T+uXesfdEbI1lQuWuTue7v1ixUf7haxHFW3uz/j2VqDoWoWc4vPDMSNPXKF5iU6jEuol7UqtjDaH
//MwsqhvvfiD+CZ4fBS4FRncw/ubQtoxgTwfGXlRfCJF9y98wydQ9ZaYlTGru80plC8JeuNdKoFo
+CAG1+lI4QQlfOofeDWpE0HbuXSMyzEvQVohlZAJ/WF3JR1Xx4uoLJLy9h0xTGtLH9qyML8bPZdC
30meq3bwN0W6iTquz+SoFo/i+wFy7APOVWGzDK+LhWfatNg+b25lAQejWa0lvHtucyPcqEqwp1t3
vnDwIN2s6pPp4SbxXp6fm/weKXOaQftN7OUh3OQmcPcCSxzHPovmR0jSQNDzczEQYubkQ+1tKrp6
9meIXUpFO2EEpdL1V6p6Rm+2MC9J2YnDa5ohPil0lIxTTWtj/Gv1zZrNLXU50DswuDxFirF76Znj
UbtdXvjab6JUl+WhEQBSVPtQdCFv45FTwA45KQxoGnrCGu5bcdKUZCyaDvz7OOzCAonYBM2bdQVI
TCSWx/Fbkpo6u0pkAz92WT5nJBNuzpqTGTC2n8f+3r8RIlsAReYaTlIekSaMWunZr0fTXR7Pybz8
O/TVEuKvJM/a3dkT71RrBFuI35qiZncRbYbQbcVCC/a4x3SWLSMTV151Eunu1bG7h8IY6TcsUcyy
Fq6td9JIcKvEC9CbgUfZuXOCJJM/CBeTS7buvvD0oF6XajQY6iObSES6XTO9utwe/DHGechqJ06V
N0G7MlqB1TsXbshkJWvYcaY1OwgnQzq2D41X3rPzcfEX4hxWuEuzcI4YmUnF/iir7SAZbwFjMFdO
zC+fcmwZ0u8+uN9eYofBjYYlXEo3n2UoLjCmE0YTy+Vgr8xKsXmKqqn9ykeQjeMNkoO1XUr8ZM7v
3Pi2/JSpyYAX/xrt+fzI2ZW3MoiG5avTva4z1VnCoTGhUk8/2H/x5F5so9XdeUr2GyCz8/ELZrug
nENcxpPBKDDJKfLsu6lGsruI5PUzqwnQ2z0T8GEx+FhA8Mx43RUHnnGhmjyIQFkzI/novuzDhff7
5oHTJ51CTeCs9wKXFHW73M5x/07twXMEgg74u264CVy9mDGyYBymwsGflswFgvN7Kudft5kefyXo
R1UMBetJvBlOMB5oh+gMvN56E5Qt0x3oIINGWBIO74qs26MmTiFTEb8XLBmkGB0nPvLZFl7NhViM
qEXmAWl25xcQKKlLEUW1xoDNe+CAgIBSy1osv0oUSRDAFWImhz4AYNNM5y5ejRzMTSBcse0c2jai
SOLovuQKjTXFz9qo4vXpBr1ahThxeMJHbgD4XeMo53b8W5WEoqxkpSiwbZ+2IycWlInu5IBBADwH
94aFq48SiI0ErV0nl7bAFdrRZHIlc7wSxJ8VuH6+3tRVsA5MyBwKwaG/9hIK1pNhhX3U3LW5k90V
qqz7zTJcgQXMPZBOigi8Ee/E73ZsJ0Jd0SZWnDpwT5XHGa0YcuusNgAAJsYv4KWSf4l5DJGDN5Q6
kadqkjlCTL3e7ZbUol4zkJz3KypKUmhrEjV+Du1F15mRHMS4MuX6k+yWf4evy6DXpLu4i2EouxY+
t7I52EANCbWM3kDP/En0smaV+BnZxUbuuUg492GoEE6hvd3I0ZruY/bz4cPj2wG/XObNUlXvPIy/
VVlRDSPGIZhF75XCu3s2HHAwcaGc8rEMZUIzAhDCRhS4+dy7ktCZcUrgH1J4gDeL4BhsTIds9KZO
aP5eVsYDKnysVEePx8VHM6GyRPV99xqgi+ggMUL5OuCJDFMQpUfzAqLYlU9cxVt8998zlZYVdI6a
sNtI2HQ+LPCZBdNmBPPy2B+vkMb//Esh+jLsgwuvS/yVZ1j9eL6kIzlKKYuRCp03av1miPBWptAi
hq5FSu7NsPkBgourPkamLmyrNO6C+kodrsR+jKqbg+Xz90P9TiVfRvpyWr7TcMbFr+ttG/iZx+Ax
bZxuUrY/Tw/bzGsnqrXBW8sJVr9t94Z72hOimA/mzYEb5SC52TOMvWvpHVO5Ehrabs10/H7aa4mi
gEr6SEvndT6OJFymoMe/Yo+aLUYNqSaOlN5M9BYGIwWUx/iqtXzHM9Rue6g2DliTsTiA0gOTUr6q
0vm9g7SoaGsyzmC8yY66/zrMBJpK70dvRsceIWPzFAb0vb48fH+DpE+OZpy/oz92w3NIQVNbI9vP
XKJenpW9Qyo6BZW7gTOr0+nneB+98AbGD5I3XZys5fLWqjHeCWgZD8x84XuRf9B6ew0DiZX07m/z
ul/TP2Vl8USdOCnHsLkfXIdO65LWzavX6GPDnaCFiFoaSvpMzWHFgmYmSjj2rqgdLynfO3OsxYPf
lqaRxVSL6s7uD/MMHPC2b6PRmVWsVsuELXGlzdIYZ7H15K1seYm+0CR2X9VD4UsKvcqOH2SkioTQ
yBdioJw1hp1aUIy7FnUWoQt5aZU/IJ5Z9BvUaVaNiaNdFMLmh+vSFRMxXS+OLq2K9zRrEg2ORjvz
wTv83/7s5eeG2naGS9CL0Dfm7rH38sLuGCMnYzTszfOD2aMgNxbm89aEkBYfGBjQeRvsdJAafJuy
5uVE1JZ/1JKHns4hdBbgWi2KHZUks8Yt5TTj3l2ZUsEHlrJz2ylzuRFVxjziFzgVre5/N30aOdhb
vyD6qtsKgnDhh5XbsfspMnKqkiCfH5JcMUQ3uIII+WgJ2XqDseJaLsVno0rKSqs3C5WL3zP+CkBY
zIyUfxqr4RWnizykmwO4AFEk5b62E4HM+LeZGU0xnomSp0H6QBYDIQ+/qJaN4qKcGSXrxuUs+mmf
jSzCtkUag+U/BCxcDpF6a+pNUs4nTrtS0L5EUUSjLKkBL5Jyijlp1qQonjvSBYt1PBtlUp95dnzc
4FvyiH/qAB5AL3Pfjw3ikNKtxE5yw7fcl5znxYPER5PivJ/GHi5qSiEIUXnxFjIGbZaoUz52gmVi
pgNAchaT4O0Fajh2647QinlHzIt2ViADFPBktn5pr6Dlfd2ovFU39kl5IaaqMMAH0d0CBCT+uugH
6inoz1+kdLAN60Qb+D3Kep3j2bqSS1aeVtQeYMa/1xtHtU1n5pJHYW2q/MI59sENWBzlu5Lu2tkE
EN4xqevyhUa0bw3Eh6s2fiEeTHaS0kbyhiJE6MQB32t19t3a+PykJF6hHzmV4eO6FzJnFDDwUqUM
jzbCsdY10sRc2EbI4+Py4xFJP62Zx9/jBBF52KGiJFV+WE1yNlHBr5y7hcnmXjBerGwKnsDqfMJ8
/W7naE1ZweDnl6kqWdmSatwvRKL16Mrh1tGU9JHQmqB0RC0BsVJxSM102gccEd1K407KJxoY4/9K
GOFa0w6vhrA36qYbr4QtjPZQV6MZh00MwKGDr+JgrdWhqgdodWIkQ/K1oMtaYkpaStQEEJd6wiQ0
3KOkqMGhBgyp4cvf1VNn+ukQsQKPjjel40tUuJqf4OUdOOLh3TTzaFOotwUmvbfNis2n7wuXomN6
EME3skuQbpuS5KQt1ZHIxQCUUBOop7XOu9gv6tUzS/O+sJ5sqRbgsTDdUO5Mya7tF3UeruasvoZX
lkr2pzyp/5HeWwuV3bpc7iW0/wE4wtPsnBpml/+BQAVFFHoQOwaeSDBHPsm9AQIvrz/IOJI8p5h3
Fd09073KKJkP6rusJ4Vm+EG5zJwjcOiJVvtO5zDtLC6rla6eN9YQw5wiRFg/wTg72S8azKlbxTlf
XqoBIOgomNIrFvlj6Shum1t+vwofUiTKvsHv/N1ObgPwQPRq3VdcSwifLt90uP9AjtQweC8M8yo2
DRbogVEdBzVM/u0Ox/XAqQPXRjEDwqaumRHRn42d5D2pvKhCSyJ3cYGdQ200plsWqT6GPwyUcaSE
2OHPjM51uIBOQmyeTkCbacOV/mt/5eOUhyyVDxjQSCbaoElTpEtD35FUutj+Bgx758OLZMHuSwcw
UOPlG/6ewaJNow9kXZVUvcDsWP4v77uLtgDwIsPuEWhyG/1D9DtNOQFQMnF2+a4dVhHNEScz34pD
9N2s++jcmE+hFnlxYbRQm1L4HU4sf75dxBE28xZnIMBGZo+tGN7KqtKhYSRGOP0oZBV0YRqddolU
+6lWH7LiLGZZbdcY9MsgVOFLeQHgVhUhK9hmbRaHmUTHgX0sRDRNEHXF25b1ZDxejAtouvrhEY8g
7Ed5ga3BhsaOVCUAq+B1Qx9FEl6UxztTWNY21+N7KU6FhEdrbN+xwVCuafHxTB7jbdqVkvpY17Bv
1Fvwfvp19zbVXp/nzZHdNr1GVW9cfLHC/H9yl2WiNmpB6EsHFrA/DLGcNC7dJqoBPUJPgeXiWcsJ
ngaVub4wWNdnsXTF2PyXSThyGB35KQFohn1TFsiI6ZLU35ROoZV9OvOUS/gkMOqJiedFFAbNZ4ec
3iBAjv5VDz69+wwlcDuEskBjtowm3iY6B4Y/GyPZZl70KRP11AgSLlG6CCLkH2v56VK2M6sFF/dM
MsIPJWibQqX31KfIkWVstacrwGXKWOMQRytDIQAsZEl2mNSJ3geSyBGPaYPimBtnWjUPgOnDK2xX
+qltNIbGpl+hXKq2jWXLVhPUVwN+2Oh/gKnafUHntjROQCYw6qq776ivB4T8NcQZ4/lj4EQkjjkU
YtLia0rsoOgzI755BQ8LIOE84wxr88zokI68rZqtQOIE3ud2OvjlDb75Y3rx+nDAatqZeG98XTc8
etd/YnQmsuB5MNVdAxC8bwYgyd7ogtcUQ8EXBTvqrSatNO5z6rYfDdoa8mK2rRuPAJ3BeZUETURn
+rOQ+yu6X9wPUUUGlfknsBsWd+U+1Q80LftgTL8Z2oi2xHd8v0jbb4TqGbDUNfgkSeV8s1iUReIr
Qz14t4Fkb1d14Q/m2CT/esO05r3LrM2YievTIcmOvwGB7Gm8sWbXdWmyWmWI6on5gmHGQC0KyIqz
+g2g8nv/I12tgxVa/IY8VYPyEiiSuwYuHlJwxajZM2mfqY1zu5VPu18ntNbxZ10Rz0UBUnFYum3J
ITNoRX0oIoMG+v0i+nXaSzm3Vp/kxMZK9Gqj2xB6AFdLQaYi/yie5eysnwACAxKrK/FHMUkEEFEs
unwX2GRlIc5b1pu3emg3K1V0RlSXz54/sd0DnTkSA237gN2UkcTd18JvRSr4V9+BtzAi+Y7eEL04
Jvipe9Y2l6aI2dv81WDzpwCmzaVGBNDX9n3OxMaZI5oy3o8ZJrpAmCUE27kRFZeh2+/MseGLWUsu
PKwIBUQuXfXb36nQcCphJxJgaqTqcxfPb7U4e2f3VL6FirSOPtp1CLXyYaNLuRdx+WnaLBJZJIA6
wVmOvtkU49AWKg70XiG60TgXVwkDYbPO65N8CNcgXqyyCVgBmucoMHQGwn20FN2TSxZ/NS4b55V9
r9vbraGtg70JieyhGh7mWpguVT4A/y5qNO12Lqm1UiY+LVDFqdkZIvkRXV+kKphQ8nDSl64gysub
/vw2Ddds/6jK+lOc85EysCxIR/cnygZWOYqRXguCzmNsRdoP9r9SKwsSuNiSgPesISyHtpnlDxiZ
Moc2HlWAJVKI/qth5A7685OAbKywO6VlcGPuyxqrIZDzQTXBkKDZQadOF6Ct7x6EIuw18EWxtEZG
nCmV+JDW+yQR4373zDvnHvPKXFoT0TAre00KmkBuc2OGi5mBIoEGwnrhRluelo6KkTDg6QgWQLXd
BF9+v55EldyaHJ9D4aUB83x3USSSunZEQ9Mq/axRLwxAo4gx0nKXjiZRb8LFFnpeBYDuaQ1BQoUw
vzuDgYXhasO7R4nPvDlhULNzzGB8RmqOA1R/wa+6SQxaL/aZORaLfBHE8CuClkwBOH3OzIcIL3yu
Tm5egPef5qIG47th0czt7L8eeL2XrVtb8cpHs7lRJvDI6LgciYKC6os59uPyHYesM1KTVWEwVg98
XYMFZa41mFAaccR21MkermwBTsRlM9lQfiz7Vm1+gr+Q/Pp16EMivFmhu+EAHsKCCxg7wirADZ0O
qzvtf1z2iG2RwHVjp5x8dQc3y/Tb/Z4R2OAyc0yqp1nSEpVc7yXy4/tqqpy7vCvLx4dg+NonSaYw
Xw7SGm0FFJJZsaID1dkU0qT10K/zt3ZlxRXTfTWQcHOQwdXp5mJw16qmLObWmAOAQvZ58ejaHMK4
/eTfco/SllH1PlIHTsAa8o27/KkWJiAdK9lOIJGXUIORibKmozWofDSSDRrzaeDN08Es1kczImuc
5sPzMglNTEScOy6cbrAqB8oPmAStrh7h+smb7JaZS914tRRAlYc5Ai4+ttrAh8v9rnIb+5ogZL/j
S5GXaUOGwNjpyM+wkXWY6dqZMA6E2RpT0opX2V+hJGancKsBCsbGMYdePWszehbAoEVZKvSEz85C
9xavJ/CNF9TPN5+KsuDTskv/saM0/3RiSe5FF2mzkX2lyC6NPhX5a8Mh39UU09pvSKkcgjIcGW2E
fJy6bzIEnrS/RcAV7j2kano78BTdqEE5Lu1cMh0RjRH6kRzFk6uV/yw3dBrHzZPKrRpQjkAqK3oT
m9L3EOOf5easrCgUwJp92vvZxrrYiBfbdkBeuesDD1hmJEmE3zwGpJRoEHtDLGVgJ0JHa9mzDWyy
Zw+KAFvQ7KqN3uxGxTwdMAwO5vW0209w6gf8Ve24oSUXLHoYMqdF17nxUIH+n3R4WqyAog6EWnOa
9w7BI/wZCS3VH4weP9QhAH5bhgF5EOQGWxqkO0fC29Bpn6bUJgPsEcQFZzckLZzmfxEaWvedDvT0
qfXOs2IKN62rkLtJbyWp2WrqRUHh+T3Bk60dBRc5mh0FlVIljrGYO9878xeXIsPSa/rrwpfIGDpE
UkHdqo0PORtoIoS9T5HIXLOCAtaAgmnB5YTAHZO4hofYlKTj6wgXsxO8MKsST5/riLoq9LspaEqa
IgtXbc7roJCbnlHZw+SVv5Nmv8w2Lg8Hg215MDS2JIfEO0yH1PtB3nnEdo8TPBkLnteyoflfq8O9
4z38NNyIn3a6anb5yCJ4KlTAEe6PtmTnf4naTg0rLpjx+fi3hQ8rE0KlxRbwaRCGb5uAmBmDmDOX
93SlmpzpmPci2OIkQXHBlkL3uq28mkuRUfjQH+4U5iW3FxH9P6Bs7uiBqqxwXdIb1vgTkiXvYHSQ
78+42G39+0tOq9gPAkn0dc6yeJkZ9TG0d5Ctq7S91dUbsMW07ROfvBn9nNKydKrWlApnaGvukKFk
eLjM+yBzCfb9wpaaI+4OgizZDSpkZq7m2oxDN8nFMMy5FxnnEJNx/nU066G3jVWCwe1XBDGV8x6t
tsv1dOYeidN6/kw8qGnKOWgK7BOlasOfDlLPbmm/qLMbSIfd3Xil+H6842lAZCdgvU/yyMx/Tozs
AgRdrOEBkSUp1f/I8DRFN9xXdbeoKzxf0JHlt01crAu+PftYOJlSHb3979fO0nEgjCgypuh6kIKo
jc91JnlUazMAAf6jugR6BqcT0DEcEa0edGEkazUsgSdJD8gvOUkfFpfVoiFNIUyc198oZAp85Pxk
WAuBBwkhZ2NoSxksv1snpuHmoKviQDoXEexAZtsLXiHBdmg+D8o98EFgbkPWcRKFPSxJhmuZdFgn
DGUGlxOuWcRnn0MWNcrUrB0McOAG3Nl8Q7ZTB3LIEBGCVcl3qgp+ZFTvhJ2WGj9Eu53Q5FX4c2vv
TEROrtAjpqRpn8h/rdyUeHgY7o3rIbPZK31h7LJ5HNvnURf921eDE2wZ/5eYGRRIn8PnK9oJM7gC
/4jiasajQwGZTsdPmOVynToN4uIZzz5ODnqieEiAuYUoMir6rKlSoiPMcOcmhnTEybl+z9+cVrJy
Rtc9skTVQF+0g0aohYeuQK10MrWpXRvau8S8uKLMaoPPCUDU36RNG2Rxgfo4ObUEQTClFmGxaJZJ
ihBMKac59pK79r6FCM4HMwJ/N25Od83YaffxPChIuMhCc196PXh9+h7g4fOYH8a51oCZNjlb7t+k
nOaNvvRwEgWkTOECN9YE+IQo3zyqcUoE4i10HemyP25AOvpdAxQ8tvhNQGR63CohhmQSC05XcRJX
eLo2JxziVaEVfpHSIsEU0a1WlIFEmUhylsllwjkJtdSO2oE12lPVIPNxELXtQc8IH28d29IQPqIp
JRhs1uH48MXFepsD33pPUdEY8RFD8TwJjOdIk0vyxAzMTVSS1l239VdsOzARb2BZ024YeRcMqAXe
NcRwXfsjFMkZCqLX2wvCYbdeX0PSp+w/mpnKKboayuchCjR0MTwNFsBGQKnZ3ekVh8NTPzmlZygS
V2jQ19T4O3HRoXBefobSv882iBAFDJN1wnpDtdSm8V4rHIAjD17xf3GmrTdW0oRdX6iUVm3PQ4ve
noonf5tRJPDZKh5xIaqeodYYQg181z3YY09f8QFqfIHxDAvIXT/cM6y7Go37s72lkgTz2hGxVCoB
OQoX1f4nGJR6+Ntqzb2JvxNqZe6mdEK2MMD3fN4VC+Cnu8d/qdamcLG9D1aYchYlev4aQR9rPR88
KsbxIQxKDJI1F+zv7IB4+EwBcuZYm+TXHgzsKfwQJ7YaTRB3hju7xqVv7shlOOZcHpTSzw3jrXkP
aeuUxpQUoOkXaCSFwI8faQsezDPfpeSh0eFvXPG10Vr/Iia/bF55j3HF6/KWU/sxEEMid713Jc5H
jkw7Y4SF2+Zp0vCfm15DAR2iqbhgWTmitv9L/rixu+pjQkd9JvHm1hBPLtf7m4PGLa5EJcs2dBZP
nLH+0idZO3uIpWq3C0m5aIqXB0fAZCw1nDMN0m4QTF3pKJudBh1ULzkgX0IOqkfORZS/22w/UwNP
ji6q+OSkPGy3XITRwe4IAabqXkSfI7ekJFMt9jQbUxFMVt6uEiRSH0d4gtaGOqmhQpUwy7IEk1cL
uycupCgCBahp4vFzdwDeNYgsFs+x6uxdfSjulCX4uwEgeDIkWCcfJ4EIRPx4gZUbRtKps5mzdSL5
FHwPZbhI9P1m38sbsucG7bO14JltEDNhJDbrcJEjxMqB0LKumWaQ680Yl6+szPXpq5pVkVfXCFlr
5q+6XFPuJ40BRL/ZoVq1mQzHg8R3gPhC5xe61YLBTDK2mWTajvhJ1w6gzxRCvDF1hbObtqUOuESy
IWaKHYMd7afrr7jKQ3LEMXxC9XlJy3EYphdH7Wdkjehi0qSUpd7nPSCXq1Jj6s0I/t6kWareasj+
NbFCGKcZvYsN3JUxJgllsx/I+B8QKm6zPuxAhMQHPutkD+2hJUicOP+DVk9/AWUQe2FNFjFB1dna
Fp3/ng6hZJZZi1z73IbGYoZbWjp0RTZTCJ5mrv8caOurYveIibCObvRQ4v0LSsW0ts1ZOiZ7Jwe0
n/ancZlCD632uRvfeF+RfIcHWoUjFyuXvSPqyMgq8XT8wr+9jIYbSrSiSLr6cK1CSFw5Ot0iwq/d
8cZWAhDHC4CJLsiA25ogB/dab3XNlRzVNybKjhFL7EFvqZJsXrZyOBf2sfeqNCDtc6UEBRF+RZnw
Ov62xYrv3GAwH5mtKKgzJ7/XpdVrpeSbi5t7bisHkXLCRJlN1jVR1em9ivBOsR+FOBLQ6TxHHdfY
4KmCH9u1/m1RqdhLwO1295mVUDdmLC7lcTzw0RQK0f8jicbimo3IqY3/3GZI3BQNSLmSUWrv0I7h
LZJQxtDa6ZahvZJQjtPl4NnNmmmHOqujNQg3ScSPDmZXuQJxubEKM6+UPeSKRVFDETuBV2hb8fdP
4YL04OBi4OzRHT8wbG37YlvL18F5fJ/TEc9kTnnRo/fSjkbdZJw+70UrosQxQgzZiCa9E8lMbN2s
5k+OlgNthkYCnxAaVSG6uEryw7vPZL/hlLXtE6zSvsiDGN+vtel/7SkMnXstTtev+O1emHt4zE5c
PmP0aRiG1EJ68Ai8tIltXNbrW8VgW/8wspzfuM7VILzDK/Sx4CRirDFX9/t/I9E+RsZz08YKAXaS
6ATWEjMAXPqxPM+DT3lHbgM1rIag3JByLhLzE7H/NESEUefFK+ie3LqtrUIDhe0GnriNVmFaE4DF
Ma6I0Z13cRY9yeveUv8Ap8X+9bCu0E50PLGIjmaMQJOtuS6FJh6ph6yL3KADhx8LPnr1BVJglhYJ
4aqHwcaNU92Yf7VrNgK9ahadlH8iIwPBNxGK6KKPwpMsbv1we93hhE/vvA3bcId++IrsuE131jXj
JCosYmjxev/scdrhQ2itA/wxQfp4X2sb2OktQKPkoDsXpKwvq8eOPLF4wqnYwkopTdBMUUAiclwr
V4CH/INGhvJKncgzaESL0Za4RE1Jtd1sttILrW93rX5eg0JYVIdSdGoKmSGMlOxsZT6GlHhnKuFG
6LloThAGAc9WHkBKvVYNfIPt56AEqxbzuNCtpCFKVyNFUoGO65VG2qqvxDk9YSZdVa6npgvsstPQ
92yFYMzZ0Zpd4r57pbow78RpK75IV+wOCySdykSC90mOAvYnk70KZIpympVk9fH0DwWjNnGY1TWj
eDN34pAhQYO4CLzKLlJdcRFtFb7lvDR8Y6tL0IMa7+z8RzDYCHdHaUiYmlXlXrJudxK0HVNjwSM4
w+H/d3n+l6dI2mymWtIZEBvpXGU0yC2pmBVbLOkUUAsqEETqkiknNoSyDqCfUxiN59sAMpCWokk0
2BHzS9dVJXiU2uGU89UFRlJvKpyxxkvtaQZyJNB0c65eI4kx2cNLnbnBaO9MfEe2eH6SXuzghESj
bKkj3vAXRA6rcTymO5e/pE7uKa1nzXwqQXXPKviDMptUobESfI33DpDb71SGlYwoV06Mv4HPiUL+
VavymM8zVl0gZB9+RQWcnchLl14LblsWkX7XYXMp2ddU/deXt2hZAWfomOjjsUKnOIES2BEQT/DF
7mXSVrFukqokNNq9mhXilbzOGKPNi5iaMu8J93jksD0pMUUa7GEJsDyd7SyS0nX7pYa10cH0o2ih
XI0U4J4mJcTU5uCM0KsyP60OpzHje95KApp5tfLHJi6kSIHMl8VEuICjxOyQZXgREVp75iNvdoIB
6dDiQJgdKgC/nT4+fJCW0yHJ6x9Z0Mn8/+cClQFr12LZuBjdqCQkME9bhBaITJQGU3PjXbsr7xv1
Eddl/cukKQcLXYJKu2kYidwOStCSZpB3CounHNkgc82f78ruGdp4rmQFLFiiFsqTlom1Xhd7KND5
SFvRtEThWssMzd7mZL5DOhdFnB1WBPSSLpZ1wqa8sc44lbKmApFaXdgOkJ+MV1CIovMimKANwyRM
3VNczaxjjwjRox8YPHgYJseKB7VtZIYh0QQavnoXEayQSEjUG3fTR8S8dTnRvOt9mAp6oBVIxDwg
IlZL7YrrZFG+EVK8CSYbHwtM/6VdjaFqnSaG1ZZaUultnIkyPwEYQC2mJfXafUiM1Xu0AsDYjCpI
2+Q64sT9MnXw7IcrqFmMQ73PMAc4PwB4v5WHj3fFMEMopyV9uJs5KwTAexCkxpQ+k3CNvtMO2UIa
wLZcSlKO7P3mO+Hwz/Eo1+H44UTSHecOarIb+UwL5eTsNcWmvzcj6KmQQllSDn79eu+k00F6hngM
UvgxfRH4xdmYGiPw/4vEJCpG63gKavkFISCv2W4BqlkZS4B0QkbWm/+J4TF9uUdHfR0umVqMf9V5
ocDZjxTJ34hvN8IqGc1iYR55Krxbo8qeDKEZlT7fqc3Jv1fvzQ3ludUGMJoXXoXBIRiOuT1Nm2Np
IWNQnMSO/kWxu0kYqQai0vvS7WwITTOWNaIg+YXdU8TVCmMkneXAnfQ/vhfGOxJ/7huVaDHsvEgx
GbDdCG/X/rXHVopam2tQyGoVOxYK4WnN7dc+Smxapm2gGP7LKRcfcuFgSdWB64gFThXs4DhyQZOM
zK5/3Oijs2+49t0dg1Vh74i3sShV/lR5anM4TEUl/ymU39IsKV25dUnMVoArty0g3QoCSTdB82XM
hMFvpQ5Jl8u/oUSUZg49TmgmDImYmFHq1OJ0nfgvmzChf5/9K0eLRj7Oh00WBI3u8ZWhD7mAKvqJ
3ieuUd+hQpQakw9xSN+7u1dNvvjzXosMpitZ68KLPICK7Q+euXfKofJjxXTwCjBfWtRi8bv/yXcr
/tWjPcfLpacyvD6qCvP9K+CcGcx7J/QyWovckFLqAaETTTQ1utWV+egrDH/l+h7kbWu0NenplmKO
PJwG8LgR7sJnRZAU2a35v9kQ9v03uDKd1x/tN5nmy9pyHvCCl1XyN8cZWnNepkHKptC6ehRHzLfr
uOLe6cfn5QfbMvJLk0rhEod+Rk0Fr9/l1Vg8rHIeZ28FNPNlowWP67lZrJs+QKvMHBRwDSJALpdf
ixSAmg6zYHSiPPmlPPFV4qfYczVtSy2kimDpyFm23qN34A4uQUTG2P9fXt7JNzAfe2uMJeVH+cKP
ehAA26g3pR21TZkPBXbaXeU7OyQN+He3YvpjizxZP2WvSKom1sNySCCeHYTk4gtiAg3L0CHSzgOf
1f0v7dgLnhwpGJe6u3wLAxtb5lp7amjouVSXNcAVqznmfbJ3Fc4yENm3yeIkwuJGLE7cru+K6NdB
wZKh6cfJjcBqvdLMamjEj4mpeKEl4oZF+JXBDSF38Q/qxKruEMt6DCTNlaj8+wtfcg7qSUplpTME
rqRK29DScTKCVhsxEueU4AUlPe4Z85/V31TDRmKvbquGTd0BAvfBAStd8b4xbTi5L1Ap9dFPPrBa
YE8+gHRxqfZJVuYRtETI7LI5c0DLI0xVPS13TN4kDOGtUVvvc+djXo+AhyKBglU54sLqxVt55TBc
LvMa0Ze5SjjHXDIhwpzV0ImMjqgDERRdX5/AVIYDDjnkdTlnjXder2BwMmExjkmNzuKVLek83nCP
CNqpwYyelCeOWsy0ABrfRn8dRWQUZkCfsAPCK5Aj0m92Q1OFjvOnqjClqe/2lVxMQB+qRZjp6nuK
PeuJh1TXRpVk24kXkAU1Z86TfU91F4yb0JPpkvoUW4NPhxXcU5Xt3ws5LXtiU5uT6QSa1Jy11fpl
ndBwvaUCD72+L0W1PM+aaLIq1kDldxD4zXvCNCm7VvegvVpacudee3WCJcDVFCcovRUdyrpRV2He
5hc1OkjrFU09BtufXIiUrmsiaXqvz17zSO20C3kb9Qv1PgmNuZCs4vYCkeLPBY6cLYNyxj5Eu6gO
XdQ0N3hihQWYvSkjXTIdYcLiZiKS3irPd1YPCV1rxfzTxkg681itobdCPjAN7b/xTQ2HvWIjvAjs
/gzoMElU6pK81tDspl3DV+0U12atQVKeaCIWJC0Qka0/UfJy4/a4I0VvEcDygkudh7NXt64znByn
R6/LTDJ7x3qjkryxTqrcYI2mXXdwboAOhVnyxvMSP4ANc3/6FFENBbeHncMD7eYlZIsnbsGpm0GE
jbzPK2pf+5tzmL4UdquelNWTL5UImE5b9Oinrk7OtHPVBvSqXBLujFqIClF0tGkgai8vU8xqNcqB
x2o2FRm8vRwuIphNSypQFdYrdc/geiHN2Bq3Y1+FqB/LtquntP6k5dXVOmsRrPLI3zKJnEtssDFv
DuNUbb9oTmSZr/gsWDgmOv/S3dO+9QgtKvrZdAsoxduphhbqnWcxqbZmkb1Y1WchS7IugXcBe2+u
1eTdNyI935HbJ/X+L6E+QFrnwbiskWr8RNZKFyXCTqFfI4fhMNSCekxuE5bLtFljYNQKEHEvR3Dc
nxaMkNGe8HJQju5071lKx7cWxHFfIG0pz3p2rp7Ucq2ncYH3zFJfTzBqTOdDiLVN6yJTLI0grP7Y
CzQaLzBj4YMFWHuNGcRYR1Dq2v08CkxcfdIRtDrfmWS4/JgZzubmEK6yS7mSn6TaKwcGGk922vSl
p56w9Ha9stPNioPmo8hwp6CEXsf+h4SJm8vIeoFo1bm44ajGKazFXKxmkt5YurYPLusWP/2on2xX
En6NcQHZMvGctR8q4PDgOj8Stc49BVf53z7MwQumolvXf97DND0YoZZnZoB/gV3Uavt1AQTC8cFd
iL1zcy+Emgl2WFjTYNWeI4zcfGMy6ZXhWQcRy1s9Q3fqs+TQsBWFogaCy4I+FDMD4AUERmYCnXkJ
E2TmNcf7tfb2tYzjOwRnoHUKOJBVrisqLtS0L61pLXsr/9fHdMVQyrG+KGYwIZ9GJoC72lQcX3M8
kMReLvae0E7ZL3h8OfI87haGFjLWiI0efNkotuPuX7jfeOsPMaMYor/HRPcj9So2/Sb87WZ7X/C4
camrrO9/0pDi1UPoHyZNsGZPO4M6geWGhA+NJldbDYtItQlPDgllr2pOHEXrnsV0DFPzTibLRmzw
ZuM9ouan/N9okeO+Epr5bsbJiIVFPKMdAuVpa2gVSKBcwc9deuJFnhdpkqQSMWoDrU4NgFIyoS2c
5QMHB5PGd4f5UqTiUnIV5gFON/PAWmyD8EEgswzTGdtwzvKl8xBcbYpwxst4J36wWzcVQ3mYsqIv
jwFS8/NTNNRb55tpygbx7fUz5GCpeJoHzMpY0XMs7lZ9o9aIFp8NsjJXMYkSFg1Km9qdQbDlT6Pg
1EQsYxwbwKRIEncK2NDGYMK3QUHGHmgmL+GOrJanvCZZByfejsTHSFiXH+CX+drQUiD4svzjHz34
XbozU8WGK/KzgUA4v8kuXAZEeU2zLOIQ7bIvCNBCznJk4FV9DLO4hL0NhYJrNzj7NqGO79achRwz
Kiil2H2Mgo6doxByh2+YYz+nfVRFvSPsU7E0KaZgFcH7GULIkvBFdRON4EpowmlSMAC6u7dlySzl
p/3g2yts7UX7vpXvabqvRKeknsaY7nKZqGuphEp1ALl+5qmJXGnyq3MGpTvDq38UgSeeZ9r4bfjB
B1aKCwIpZolczEjjkWabrZnJWuIt+GjhYbAto5O2jhYA31qAOYlCEOyu3QgrjaeB5duPGfS+n5Tu
o3En2VwU21bTuYDwk2CdNVOMoCKPJRGICIH+0nkvmmYq3tBMECjCGWMWn5JvwpFW4gr2vVPhpp0r
M5x0piC+JaCxmEO2YeHdO7vTMcvxluJ1Avf2Qyz1K+Ewo3aSkNZoyaVYkRKJvqmrK33JJLhQAiVe
liega+Yu33COQJzSRTD//nlAQIp+p8e/TM/fXbtCPMvFdZlFAI2b4XP1opL48ez8yybl2j4akAt9
Ad0s+RACFmtaFVRNJil3tQKN8XuMff846c0nEoJ3AamsoMmHPJYmHJcXdEDLckt8fkHMBmJx2T62
4lhSTzTZKa3wWNhjzuIWDX2uCT9gL0q7wlxw0e7Ax0rseH9nujDiQJKu6GL9oWkgiBA9W1dlMOU4
98Y9XUXpCTH5y+c/oi67Ae6F5Cw6unWJTVVtsnLeq5Ye4+1xSdnEj+0IbhCbqUVZMc2u6Vh3ATg8
h/RWDpxrGKu7oI61EZr6KR2sULJlrF81L/269J6LYhHlWu10JUv3p1iOBZmEV64Jk1fFCoJ/9YF2
fb9yfLRXPzhXVk/fu5RqMDHuFxNZqGE7RT3nB/b8kzX1fqKmXBO02Kq5/r1XxQeMP2b/Y1qhu1vT
xWkNvz69qhN8z3fuSdiqNue7r2KO9v7SnItDb+dNhkVtuGj6QCFPOSs869eFkyKTludqjJcvf+n4
ogLbJJ2bFc4wEMxKV9a658CNQhmlOOkb9QFMqO7IL3x6zhLn/wJdRIQXrvwe3EhONMEjR2trVZ2g
/QyNgM8wmJcFcbmCO+RNzG9bN/8Scz4xISvIIHDl8qzynOJNVroALxVVWEF3KYbSOv62eyNtAeRS
+aFEAYzIdgg6auoRWJjObQOU2sS62NhS0vREzYZV8Vo7q335oM0JzSuEpkFfPlBrAoUX5VoVFW36
x30tAZz9nrhR7rqIEKyxca2Pzj6hLav7yPLM8YFrbJwXxYhTDp75rHfGBxjrMENYLRX3SgKGT7mf
IPyxnx4ENbFUnhz4UUy6DPdq+4FaIVweLuUufSxxx+9y8thNesQlGBAqkys0meswwN1aC4C7fHGC
fP/oXDiA5okkUVGzVYuT0PQtxVoXWVgiIBy3Xl/snSu1i69uGAPlRSXuXNyIyOX7B/whjEUKWiRi
jWOBQmuiTzdMglv5LQDwuS4rP1y4T3xljv7UT8ZHJ2pkmmhn1b23Plmh7Yj6k68QEsH0bwbMjTvn
lQFoGEFTIE3dNNUKM07rh05VUpHfUy5fX9VesyzEmuAZS285SR5M01JY3MTSrp/EvR9GUozrhGd7
DjD0qIOLyadF7J/Cdw3JoNEtmYIBZeI44QH9GYom4iWRJewgZaWYbmttlJgWqVuan6IqwiUdVUIH
3vNFUqPRUqWy4e13urRfMTpqLiB5rqEyjxrmsEorqyzouFCCouz4HwOjD89cg0Up2w1rulJDyRst
MpcT8Zf+2f1fAKooFL17nzgE6tc3+RfGOuBmSXsCGIbVoZLuxm6DYayKOz/K9y3Qc0ND0yfdbylf
p/kAxyZZHF7YrNmcMuliDfrXZ8mNErtZUeJz7KhTq29AN1roYTxMEeDA044xq+nAqjPDrpW6ZgXs
LCK+EokoK/EZp2anpyo7ZhF3IsXcyU0zEX2zpRMeOpI/nksIXrraPrYU9Vs2oZh0liJRJZopu83d
5Rdxxh7/Xfv5wjf6DYcBFqFn0rXXI4tdeLBOx8mRxHlvL8bXbVryuVmDMIwJ6DFO6T7gTLN1ZQ1u
uyi3AlV5fEEfHdUehTVam2+o/Bhg3whm332FndfJssDEGb3hsMzo7SMzrSBh2tstxZMytOHNpuQH
9wVvqB3pdmlVR0uJWsxv8Uz3rp+Oq58oEaAhZoZ1AaWDeIgnfu9qCPw+5aX3YRiMj3KowOmmtchU
JlZelV/bIMzCZtOZ/8wTzwSeLZjkYQvMv8OrSf4d5ZihklYwOYbihUieBcqJNtyYuRBkyW8B8+/w
7hw/Yw3VTgzhlz1mRHbDu2hk/uTgXOWEYm+7Jbca/H3o+2GB+iOtf25iHucAZbvgJdevL8KRhx5c
yNWt/7E/jN/cBD57U4QWF9aMKRJgf0fnkxvewya/0PAiT5EMNUWcL7hBdc7EcwYmgb4qXvqi61jK
LVIUN9JCrH4LKqVj3LXaO6DiQ8Y0eQz7VxjdZM1LzsUSq65HktYgRPuBEwu9uDOQSTyFTIe0ccFr
Vetlmlf2t/KvHbwBb2ZCYK1ADRESWw0wWWz8L0oEkiTJeFd1uC0RkaqXgwwwbder0CAZWjMXRTm6
QkgJULUTuvYKqUGUNrn9acJVyT4F/4e/nNTESVPb6CDAFiBHdA3jyEJvqXBROoO0PWtI+lzxT9yx
YU4pxibVC64ArwswmomSDgI3W9nHcLDpvS2IG93VpfkchVMc6xqQTl3cDjY+AzSfjosZ4rGz8ud6
L4Og4DOZJ7c8gBw/3qIFAyGQHuFYWuox0EdeInR8EHuSu6tSXtH/Oq/aatnLvTCT+fXAzI2SBi+S
qOEkpWREN740X96Tqa4L2ZUsTp9fZ1iTMzj1SHG8zbbF3lteXYwgvyQBDIXZ4aFl8oKROUPPlOXa
AAd6A3C0i+Jy3G9GkI7bXbQvSAz9u6V6j11gHZtFiJOoX0kpSNCMAVYpTg4an0Onc1OhjRC76+Dj
IVhBwXbTx34HAz0BDyNAYf7HrQXt0Phl0+4O5D9Q5GU0RtaxBCrdwtbI7sX8rg64eWwOlhU9VZdO
AjpFQuLavfUe86zbGC8+uEEu959FDutE5gjHUo7JIdRacexFC2tAIs7RSR9Z5lnW+ZveMapOhOac
oE80hvynvJ6ob3UQf8EAg8O1m2a6TVq+f+PT8Ck6jQ1eQClsm5vB0T97f/OAivkbNvMq7G7M5sZk
3v/H8HKZRb/8b/NqzN/0Poh74YxJat0xIx0cdknjLn9c0/IX/er6lM8gFa7DTTwuSMWIT79ygBCH
3pWvkiPELt0d5SYr0SBT0hgu4gMmACnqdMikIz4IF8UNOLw0+/1y0/UQB293k0mzBc/LPGOC8g9w
u0v3nz5bUTW99pihcLWeX8CzbvfID/1Efbx5xJNAaBoL2vfS6rIa67vUNbyG9vM+9uLJzI6Zt2lr
5CAY26j1zbsRe9bqr8PGP4dHT45Vo+/0eDzCCm2HFV7COQCs0mt1NeahnTfezDil2ChP8B7w/GxQ
Hn5HvSdUOiYBf2KyUPEqpMdNRpBRmzhujkZuPPdyJ5mzjNLUlY8aYOOP6l/9JwEqMA9BB3dCwgDd
zHJoFoAUgTfn2t25hKIp5hpFsSV7F5ouj4Sj3inFxGPcJMrf54m4ubVxKdxK1tp3BIFc4V5yu4n7
3oKkZjYoFDWJ6nEv6MaMHu4wr1X2bJTfA2cENhCQzAIAoIMHmYzFjDjthRQKlddHZt74pYtiZMdC
k0jfWIaAElFWN4h0GDGAHY9eqYGunUAuu/A8FgOecsPF5yHFXEFTKtn2As0sM6T8LLqANTTO5phh
4eyFy6jetZJVHb9Cuf7WiH0ZO2VnmrMRgOkkMO9ypRZJd+E0AmQSzgiGUaCZiUGEwaUfCgZB2I51
/xzeZ9cQGGo+ko+Ri8q5r6i/mxhMqRo5BhccP3EzRHOToOCorTL3jp5KbuPbS7xTvb9nKhYwJG0C
YhzAKCoS/CgC5+iXZLspMltfgxOpwfvhjBEO/4ju56zog3kVr8LB0hPKNGPmAni0TofbuCAkoRUT
8iPFRN2HoE2fvW54wvFHTQyltIFmTIME0OnGj8GoPix9ZTx5NzTIIzXuHIdrLH6d403b7F8QGPr3
lNYfysYfF5qkQDCiJfuIhl0Jvfre/CbmMrF+tjQKIasyjdUh8RUfAxydc+HpzkIYwM/RFvvCu27g
gNALzNAulig2wcf6FyIZEsK1a7XESqFgx4EGj6hPZNKZK1C9PQWegCODF2fbiawwODskOLm0PM8n
aEG6WUJlCyGzezJxHHhpj7YuOB33vWTtJ/7WVKbnHV+Etcg1iiPLAsqxUmhcIELveixH9GDTa3WZ
WW4CVpw+lEvntEhE7wQC06gnl8AVjfFCnjExxALKNNmjC9ZYeTKJxcNJSYhddWLej1kqtn7KS78E
nmoZcKh8Zt1ewvp5BStPGqJWH91ywPkb9CDKFdAg+3vDmmEasmlbwBkPl5Kt0nB4vYBfv5oesjgT
cO3B71NnKkodHztNTcnMeTZKHtD6PujC7q6IKQN+5B+xF0Dcf5Pywx1d60hD1YXpOI2rsKwYXXhh
j+6aAu+wxpktTg791gMZgfxsm28MlXIivEQnFeyPScypkazPdZTLqVvRqSaV6jzus4JGXflw4WRh
HnTJN+dJmeowrqqj93LzKl3QxBJTbh2nKf4EDjZegV963+LoRpDLDA73Vwbxowk6+JgBWD51l8vB
d4wiQ18lHvun0hYCfYGrZSDJCYi3aqr2LcKUca/G4Q99jAYqA8oNdt3U/AYdqvqtQbt5FT2e030e
4xi0XnojvvhTFT+72i+aY5/q60KyQ3fyBtfsjUdHtX+qfb0+dirKbWzQ0Tozgqj4ns9CnamC5ogB
MAUvixTNh6TdJHqUUYUrvdvvAhFKKnknT7ByQE9bgjDik+7ypA4+gRhgle76XDrZ/Q35moPYj7JE
wf9L8jTbdT/Ts7uwOa92+Ifd8SMp3gQ4afXMx9YtAbnJaKOACFZQhnRHoBtabaJMtTPElju0yhki
E6m3yAqFP99ow5Oy+O7V4IUCI6TOqwO+RKOkancLJwwYH+4uVmM6+E2k2MQq2NLrmJ2KH1ROQXlF
FrFR7RGNJcjG3tW59T1pzNGsxEZFa+irzK8FZcHmQ6EBjg54keTE2mFO9nRvwnYK5NqM2L1q/W49
Sf3mH21RiJ4HEWuMpjxG7USb02IGIXxJaBEBIZsRQD+9TNd2iaoSvgbOzVENYLwZjBuqnKwwrtyN
kmVl/LTD52v9za9pLJPSlXlP+HzNMxQN0ul4+esyt+niDtzjLjmNi8b6PaZbHAcqfdcOZpZF07yj
+fMILTcIAaIgOPtZgTLmKuKLTevxZsI3xwr9rebQQva4L2XFKCt9dYWYEe/AUCDJFtfzEoBttA+5
5eRQsNZDOcEVCOUe4n0pfeWxUZT5ObCtZlwW4ZQD4hRY6RYdxhawU4X01W/VMWoURZPHORtIxaKV
v4NtgMmga0LB+BT5YpVtcgj5Kp9iafOtfQr1EM0B99VqkMWBSg+zPRUPC9XYlfOTbAAMy6OJhfm6
8RP6d4scXiQAGytBxJ+6uj4Em0EKW/Mfofradx1EOX+BAlm3jkCK3nrmngwJLUDflnUgekQ40Bfy
AIFjx7y//Mc1f3cw9oIirrDyBfSyfzQFiokmw2F99B88P+XZz+YiU1K+Sqy4eeFIMVyss17ieriK
AcW445sjw3oFCYAZhJPnuy79S6+pBmc/Kv1CmiLV2FnuwPF41ExlFnVjty9qQoif7SMNDFPl3tGV
X8NjP1L7EKLQ3k0nL4DkCbt0Ss60rpQ5jNanNraSIFyxeYvvUNUvcz257YZRVNUvwwBATM9cbIOg
1MiBfqtC1ZS9kVc/jL4WdUoq4X9qszFHN1nqKG7XlID0mN6oH9yXw6nfRW7ITA3T3hg3kajlrKbX
dyP1xoIAUW4GCRH4QnKxf7o9+EbblRO0kY+25L8COrmhpeEp8Ces+InnJAafSxIBDGJqnHAhkftL
FT/g324K81yO3eJF/QeovKxCFN04YMob/uGfyBmbsz82yrEdElU9Co78LqjI0CkF3tXz3w/jKZIJ
LvrVth1V0avLdDgM9SttwS8JeNO2pyjt8lU0gKaWBt/W7n0faBehIsQQUTBPFpaAoqp7mkdYkcck
oR8xx9KQL9NmTwYsv33Zu8yceG6hJVrKLcVUDBc5Rz7GClIW4arxjUyROn2TmlXhaUidPRjy5gEG
LoYux3QRdgOky+EkQA5qzLxZm9gOVy/DwJWiGkU148RXaFCnqyYGdfNpsAbzT00rL6n9brxopgUt
75s7ywPSmZ9FfXhFwmbxVN091fjn/2nq4YQFOa3E5xK1N8Nkv20JpRGD5+FBuAYWV47oczEHzor6
fQVLUSLlsVwWxhWEa+ad4YV3FNp332gMvxtU0/XuxWT++UdrZRGE41UiydZTq11bMBgBtRLOZI7q
zqcQGTV/U3y4RGL5Zs2QmtN+bm3qo+RFmoHAkHt4udClCX/hJhJNsPw7rdj+n9htLcg1pbNGcCyh
ujIHy5ZugOUJ5CaCK+8HLSbfc9Lbj5R9jAZpwQyVnryUrNQRDTNEHhmC8/UaVT/XK+gFK45sxfwZ
Clq4o4PqQgMjuv1OBGU4O1egicLo260jKUwT73zIiBQatLyFEfo2rMvdfDQSQ0tlgOIjJJ3cJN2M
Hqg/jzrWe3oK4zVCS9AgpRPgXh3GjQazxkmAXpK7Fk4VrVD/aiAVDAtEO6J3YDgaleIi88BUijFW
OWV+OiGjH8olq6PggCdryT72TBGrJsZMprV+QsFfX5C0BZMTS14FzG9TlxYnFS69AfV7UKPNzGPF
8NqP+NFR3art/YvO+4jyKQ5eMesTLb6Jq7fBu/w62pQIzDmNudiToo55alTEcs3t0/s/FEyVrK6u
6Njuc7Q0ZhChw31l9WdS1+LwtO6jSEuuFhdBGxwUAV7NUqv244HyqiOgIvEbva8AY2dGDLBhJwh5
+urAMbWUisd4wMwFkvGTHdM/bNw9fid6nL2oRqQyjAnY8cjC9c9s2O3yplt/ofUITF30CFid07dq
0YpCAep+n9ozMpCnN5Lrl0SGwuovF2vPfRsisC8W5OGEPKNK8P0Cc9ALM+K5CCTIzR0VwP6MOUw9
di1scDuRnMbm8toQW0Wd/LpYylhEUqFj0KxDAmsBTAIuqXqonHsveiE2mebxaiV1rbTcG1TtHbhg
VNsJfY+PFN6UBGi9zDMJeLJgbXkoJMMP+pl4r4ZPiFFDEl7IWQCFE2chKkKmVpC3npnMyQx0bcoq
IGXZ53Y4/BsVDX8X4HQEFGTZUkPCrIRhjePQbzTXOx6QUnbYxOK3FZGJwrHDFLkZgUPIkXS4+Nrl
4xIsNwd6Zy33v6VfTZAvOkHJGd02oaClMMZRXDRF7RgnOiKGh4i1e3sWGy6WERwfK8fbz39c8Y1d
QxaG4P0bWhLQ/qCxijNLhSGkW8pRbGHqr/EBrBEunzvgibDrrUxmglEWPtfWHAu6vmx+O7bFhsgt
k0aKYoPPk4nvtpEhn4pcw0L68eZLf7XXvOhgroangOXYGHiCqUbBthckTIYLM0lyjC5UZ3nc4zVG
5X1jniJthd59bfVguO3D/NaF1lENvIlyl5ejWR9WKO0wkl/3SsDF2qtOpWHtNzjSxnzwj/g8GnFf
T3a2Pvk2aYv8e7yK2sQGdYMYbc0V5hvvLRujbzincLBJfV6ER39etx0NrOKhbTKYYdMq0UivvXOT
IZBKFyxZC2Ftm/lUj5tbY3snPpwIZ4KQkwGmZ55Y7/i6hjqWhhkYFBQ3OvhFpo5aIOhnXs1VF6fD
4ksmRVu28Laa8j2Zb4BN/0jd3wFV9GY2nnr4qOZtZXIqfFIcNlJ8QBkpF2a8hXPQesKYSSovQ1BA
/EbtNctaWRNkdBS+YBlpaZWtHJaHUPUcLIu0E6adDwL8DQQHRxV3DULywU/F9rsxpSXsdvE4cy8P
slufajNpU+DhruCz/ula5Ef10Mbs/yMefzcO0pU+cQ4otpJfwceBJUpKlfB/Fos/g1Ob5dmcn8mI
cIR+BNhcvkB0tFOji9RCaiEY4SJPuJD2ZC8VfQ76CgbXpk0JhB1PHKJ8oX0lg+Lj6SWPpbUdh6JY
NSdVBPsz6Ac2PBL+hcGWmqh8jpNpciiiQ7BrZU3bUODe0vE6XkBDJN+W3yhuZTarHE5o26fRytsI
mFOJyRCaqNwE7z4voIgDdUp0fPeuHPOTMzUrwTw5VqFDqk4LD40S+s/SS9bqf1R2YB/Idceak8AL
0dv4rxjJT3n5695uGwQcEaqn8Fzlur08iPYxZsYTJkZKJ1BAndTQEY0udILuy586KkXlHfMjui+c
Q9RmAEYhyNVDUUGmN3PbuxiubEorKp56ZJ7ACHMSsiRHH/mBaG2bFAJp426vzLx3UKqPHI/n6Kb1
8fwEEPwv8fUsCjvDzvOiVLaaPRRihhD74Pn3GFzAzgOAd/xUUai5w+Zh9AV4VT9rAznG8nWmGfVe
SmZyF1B4BEyI995hTHQtgC+X9tEwIbnUR/X4XO9Kcbm+8hScVpQOANb9OfPuJHFIl9r+e38CZpW9
fGEknZzX36UxoZ7nk5Gf14STE0nvtdNYP4GhsJx/+JprAxzme1KJ1MKLVcgSlIx44VRkWe5dB+hH
xoyaShIcUZksmKESi2+Z3MQKy6dYqooyH+L8XLNvGtdqjKVPavdLq57ec/8UMGtOTPks4cLgtEPC
AValMo/XxMBV5HO9jFI4/Qc5wc4QRjtU3QWhqoK6UoNp3NJr/cghYG6vs1tQfClxO/23xD4OwStL
iuFxKJsX3zwdre/fEEgOVCftTAJ8OsjrjEECz35PCBJBmPABxkuvtlDcXlP0JWWoywSQjCbqZAfv
gH/zo4c/Ck9wHGo6Ja8rl6cOET77c5K9AWjqSeKL5eQRSjN1mWDYoKEnwOz7WyzMX2NUZo7McKWw
dfXPbmpFuiBzbB2IAjKK4ON3rfQeEBMTzLrz9gXMRcP4mL5op6OC13wtOavr12F2FUmmMCtR4gWQ
icnlYrwSxwlyeJo4It/uB1qwtaBj70t5/o2S5fwMuqxcjhqnsFa6MVcjzt5CuFPvugt4pPagUCkD
j9eEU4SZsdTh6HikjU0NcOwW4kV2HhMrrcUN9nmv/W4yUBK2yYxZUyfmHdFco4CpMRGJWl3/DIV8
iAUWpR9QFw4HsDM5LHpjB+2W7Pn7LvdRVbpkvWLf0/Q/eoKtRRjTSTNOzHJgxPgaptBEL7c6JVz5
u2akp7290YbHgPQCkcsJWc7Qw87ocmQY68KdTWBvaUET0xWgzBpoekwegSZ1d3kkq3NPIPLfy98k
CLYp5etYPYoNEHltH5k8PP3C7fV9VgeJCLaM15oaC9TYSWKOdh66AX5ngVLks82UqT07hIIQkv6c
WCdgeYX8Ro9JqXdX10ji0YVV56+sEJG3blNUpHDVdfbF4lAingR1ZuSjW2BUl91Uk0JIitpdkXuV
nBatnyeTFVy4xA//RrAnWVVZRMpDObBhmXhoKChUonmuoo0obO+7enpmVxP1MWhmGxBF3lntjVnZ
J4UB5Wq4H11nI8Uo6ivQs9/XqykHhJremFuq8HznW/kKZlZ2gcYcQ554qCmRO9Fb2wR+OF+bHlCM
xjRAO1o4N8qvk3C86dMoj7VJRXXCjgGlCMKyxO5guFZruOZUL5e8Gkqfn/PYo5woWeKwvXbH2yZ8
eJaNAs99Ms1hJ0bCiahPVZCiEq71mNroGnCIJIzOKrhwQ1T1+rtif8rKdqfw5A/MzEVe9n806mTE
bAiIa8hQ7xWjCY9vKOf7Ya5drHPcM3c92aOY3mYTwLD0pH5Vf0UboZTVS9SRr4/IcNX8QlTzLzmC
w6VFm1ikbHiszZWW6fL2dERvwKwPnEtkAJ5r1SqDwLQ5Bg6e/9xguoSt/T5YTRml6wy1cgAGhzbV
hG7k8OQCMFL9wo2E/OsW/5+2OByZXSI1tDCW31EKeEasR3weY7Ce5C5CwvoGNsTtLzRGSSKqj+xE
NGs3cRyDeCPKoYvo/JQtEWKzbBAxWq92SEwjQFli7kBtGdstL7o/as0urYfddbcRxE2dlj4OqfRi
fFtGFTqcZWBXVa2lqIotbBEnvuq8Va581by9hYgdzFKnory0I9vJGPdcZS8MlGDpVpykgapyY3ca
FuT4lWjFhYdve2xP2Hn6zLu4b4TynZD3/DpYIsrE4my/oLiJUh/i7WT+ieKwcP+zsIHAj3AOzMS8
OciclOdEr6NMxwgp+c3TdYfFrCMX9FMhHW63n8G0ttUZSr2fYkZsXYMyqS4wrbPIdRCCYXpqFPqN
t9frOY5JXGfzFkrTVOoYbUc0iC1wMijygqqy8CtMMhox+ixu2XnXgbvp+l48XuHF+4M6K5PF5dFb
KI7Mk20BWjqLa6jVNQuPo7BPnCAC37CaziuCYvabuLIHsNr1YELPLBmK/NMms9BaAnZv2T9iDWTK
asxmter7PX4UAhOOuYFqwHHXg5zuDInMw1EFMtIWRShfEPk1sMcfKPxiF2YUIbUI+zGLTM0VADNJ
jpZEau/kWEoCdghgnHD0plcvi/sQHJuAVPPuJ5oDMVSKxoyFT1bDbZVlJ+wAXfaLkck5YlbBS941
kYqG2Wlp3vj1Y6icvKYAC2qZi9HivwBj9DiywWfrqAHuHMwQxiAL4RqV13a9VRoHhtqzv2+OiV3u
z1a4ANlmUCV9y/Rxqxb+uZPTpvIlgDdusXZetS5FYzOsNK0ecl6AH1guxX3PeLMCzHcl/P2i8GOE
4ZR4TKp5iAqL/hJehRlKO4mPQZtQZNyJh3Gvlx9KhhFSvXAWM5jF6rwFQDBrfrcBB5gp6ufgfNC0
wE/vxEyyrq3zgCkh4xIe/cQ8SYGgZAPRwhRlNFFvkIJOMV+7FurgH9Jr38k1Kh8su4hum7e55gec
42Z8XBjQiBadJCbV5927Yoc3MUqFDBT0Q4gE5tpIp4t/D/IcO1DvtizJD3PaKf2G+9eiMCiETdRB
ArcedgiN+9FetjZNhxZyIB6UNYxZGjztlCpbkegD9pAdRER/REflT5K0kFnLghgbdx6oIuovmzpR
hCVkerxWBoJVdeeRwYUeKMkoj/wdxNWUb7NhtRZGYtc3Uc+NUOZui/OU+jweKlnotC0e1Az7uPKL
bTH4a5Qbxd87ZM3vyCRCR+PlBMNelrQZ8MUiN5weljwmtgtuL2hdfg1wO2kpJH1Im9zK6QIi90zd
g+nrMwjRkx5gRrYfRWXBA7xYmp3IQX48m7Z+Oja8jrpdks339/x49uqWrpF44PchdbmFAg09khNz
vRN5ZDMPRgF/dVMr9SMZlBLHhE3/I7EYiIS4vnm4GagQZ2E7LxMiTG1Aq30Uh+VyU3I3Hlen+ogE
A9wjanwsrF8n8nzjE7DdGHXhbRfq8WGW4Kzb2N+oR4ZDwKQA+UPzdebJH3nF3aYwCy/jr5cfDHpd
i+S3h8NwSUXUJ3vcKFgTJwV/MTYVUNq0Eu0pNL5INZ3rDfrx2g4InU9koo5Bc18N5L2PNPhWMIYI
uRWPLjn04EH+gX3Rm0cdXwGoXNGoYp5W/puu0Oy1mDfd3bN8OhWMnxFebSBKNf6NWvxguUlw2kvP
kp6MADdz0X3vK26iC6WqKgnX/0Y8ht5J4qqmMs+30PN6fa3BFTtCIDLCqQDyNWl9NkjhmUkk7sfF
Q5+K4+LJXlNdJeEbdbWYPmCZm2ERVfkNnhrt4ujZXbwUdRVEHT8h7xrWxnPyXH7zyiulM8GDzpv0
EYoLHoc1/LvIR8zndOY0hQk8kCQLI9bf0te+USB75UJ7Ta+PXhmaSe88PWcLra0n0SGX5Jz6AUVg
ZeAQd/gUksB+FhOCt9bqBeM1dX38IC2at39WcISMRedkXN8LpldcHr18JTE3NSFF+PQPu5jS94Vv
DHPRWnKPYJ2pOAddb0Fz4LdSJF3Tfb4IwUSgaf32/GLsLNUt5cSqRE8uMB1iFGJg0ZIJhyzX/uR2
GZsJ8hv7ozoalOcLa/krjtHNbTeLvYVSISTs1I3RVQLhRsbLYB1X97NLlsjhMvQIwAQfWneOrEon
wHtOPvoBJdUfpOtFLb87FkQ0RGWsX9BIEGcRndriOtlZq/kxn6eDljASYHjw+4TTStjo+t+tRxjX
+ncM8XusF7MHuvJ2qnVfUJOSq14si0oLXsFYItRXtXtgUvdRRQnUBvmkRplteGJ/CbDBghM29XZE
m3H9j5KQG2IH0ZZNMobXccWcUfx7TV9wXrB6UPr3f4A6yiika0YOI/Y2zRPbZ+vyAZNfc+CyPqlq
coZ7gQOjYoy2zEXujQ/7NqAIi33q5dEpnYx/kEZnGzMX/JIMBIZN/IFp8ojjQgvmhCsUpZMeb8Mu
EGyqGGW7BBFpli76UY30kR0UoMTMQ3lqAmJOMzxdXjiLKodZhCay5jXa3JZrNndbmMGjfTTwHCi5
GrsxA3K7YrjvrkrnyYiTMmOjD/gIXTycmJytOEbJYDWThY7vmJhWR3ImOLPFDVHBFCbQf91lX/iB
OvAoZK/b9Ux4L8Gll4fhfjKLUCLwiEhpZ2S+7xe9meMTbNKRWGA7z0r6WccJWekQuxmqCvtjef8E
ZwKT1LGvRUHe1sogldoO9s90Kh1h/2U9jw0rfhyO5O7eWe9cvbm5S8ZNpR3dF2lRSnulJy1N0rSn
+3W5sjr2VWGQQ8V9wYMepsUmF+UQZGQ7T39u1P5zMR3C5tNkMySUIc3XFOEIQjwlC1Gqm8jyrxYq
4mlakqCnzCflB0NAtNPQYISm4oRLPhjRmyt7Q6dDZFLXOwylTY5QybC/oSfWALsJZrp3nWL3LAzO
UXfI/rdifw3ztpHMn+E0Sh7dThAA52R5c58+6g1sZF5jFE5LfO04hn02Fxxg/XpfxrXDatL0y8IG
Os0k8R2Kx3dMbug7OD7Ixpk21S0tVULK5VyWudGXexP5pX9wnPjqNBkhIwi1wp5rCYvKtV4UA+uq
DkFSw/LG8qs+h33PR93r6dAqgkjrt+RJrwoXO7x7rfeerdNUHaeq3xexlg0NW+GrkEYsi5f5Q8zC
RYmcBfPLGYndwXTE6Mt8qW1qczEpWWUoywgEMshMdYL1nZz3jkMRiDi92extUywHKlBpfBIrIcQr
bUzWfEEkflzbY3ioUB8noNhdCqBQCc85uh5A23VkZEaNzGVVWmFG5Nl9ngLXg3mHOJeuziVI/sIV
bX9VL4r1D1d7n5FtLVv8pm7OFkCvg7w+1LC2cBTWeGZYk+BTQrGRxw4k9svEOicA/kIDMHUdTP09
lVPwRACxL6zKWaDBDWDe19/JhjBhj/rGvasbA4ZzaKN3NKKc4YVC1I6ICK13bFU1Dd8lhkAWOabn
Ubq0+P1gmH06bG+hy7fVxqwsANKTsa1yblijgk9oSmUJde12IUIyUk0f5FgyhtkDeCbizoHSuNQE
V5mY55+PmvwhSCB5C5kRQlMQOSsb/PlgB4xy0GTJ+0Bck/10lLPAYDdSv9VsXOzG3FPHZvBbACyK
Dz+jmRKtz19Gq/bOOqYQKi4QUFVpDiM64sYO/3+29AlFit95vq5tEVRjMAPbTWzuydK9mvV68vCV
otukonPiUthYRDRYm68Pmuak7Rytgn7orudgnuFhOfSd8tAAjvUrsBFAe4BjjWUKTk3WmVvnLLeI
dN9AYvSmRkV/L6OM5raPVr8guOCh/mkgrjIqWf8vrMGhjirQJUj1DGEZ+YsGQil12xMwHP1Wss0J
KxTI3qRWmRoykODC93jnOWqAvx088ZQIDekPy5vDHZA9VL11K5ONQGuYZ7JZ+uuD+vWVSl/P3y/j
LKco/etu7QMfbsNoykI7+qVyI7Yl99ePlB2RRwVsVNVYRgj1EDXV2vIS8OyhMBnrF8SzhrAnICZu
DhrwNJM/zFozvUYo6ovZE8lF4Ng+41Kp9CtPjiKQaEfPEU6wyQlmEV34GH8GwP+PHuOmK2k+/EXu
XoBrB2d5Yt8OLlxezcj+nnMw1Ps2QHMRWVVRYu6kJ76Wayh1tzHfVmScCMnmrV0KvzcYPjYgXxQD
471jwXida/5aKjlZGQnyxkNvyKsdNgbpRFetyuhtDP9EIi239fv9SlQyICkCv84W4U3/Af85Onzk
/RhExHrHsPln6YeD2sdS566doRotFofB22IV4IzY545QcAusPUN+COh3nGlHlZYEezk+KtAanN95
D964asUVrIQt5eQAZ3GYah6T5e/yfGUqpu4Q4zRLjI+T7RKvnND7mObXTfEXoKMA0XGFpdCyUANi
ZgW/16WfgILW8SNIwtKetRdG1RAZV4xPJnAXorlYqHzuffJODwnyurVz+izRtHo7WtW5jD9fHpXN
nf/lvwcsPaHZuRlwE6ibHHtGKHdznVyZK3Io7YixiIbh3eapdiJ5tBag1/6s+yQcLHiaOmnrdSr0
bjLo/RpN5/+U+mDMXU7PrDGg/P3CGiWwV7gBD/4i8RUaLLLJ3O/dhvqeD21gC6+VptdgU3P+MZEi
xWX3iFOvv1Mtbn76EkbUn5yaOawOhH/QA464nq5L9aridveNWB/lzHUmR7upRBK82fNHrvdpDGPD
jcMR1yfDzi14aArTJl7nXP74w8GdMylEcxErolqNLf2Y2ALbJhMjXpomscUt1DhLMLm72LaAsr4j
mv5tJlnbuTC0uV+bZDF7TwWfGd9MX03dTJvB6Zba/ntRY7NRp7B8mIOE4/s6ZWH+wQLaPBYZcjyj
Q/uldblz2bf5K7uEraPR3AfTvuG/zrheJd/PtxNjbJKVfq35+s9uCSQNCi799djB4wIFA/P/yVXT
iEcQgcAuHj2Et0+IZdsncpXNsY9jSoPnL2Z8sZb3Z6f0VTKLvYpwf8aAlV/2m1lWaGtUv2VJDG+R
l7Xe5KtcwcCf1c4gfzR4PFv2qyK+hXRh5Ot678EdOZ8Td2jitbO4ieB18sL8m7/cI2b8gdL4UDZy
/6iW/CmWj3jlRflG8lF60ASreXuYD4lAen3qIvtl5E17Df7f/KNEJC6xZzjIpe6KIePp+rbOZl7Y
nu4uh251GDq6UpxpVkPYX7oxbxY12a7mys5YORzYs9mJgxMRI87HXOfQUA2DuDlJLEseP/GhhYr+
pFMdWEsWOvzOw1T6aucQikviWARJHE12lIYdbP/Fjft/UaAJ0j/joY7er522l4upQRv06lWgOMh4
yzfhXQDtA26omwaE38hhbCJ+ZYFm1Mm2OMmO7IWKXLUUGsFpPnn5WqSqUJGRA7vSHhmqjXI8zkXS
/fGEmUAz/DveVq0mp/wrgtpHbna5dATV++bR2lyZqWY6AOUJO36mHqcc7XiSQWMk8A0H2Y8DRIwr
6+xp+xnwNmbfn1o+WbpdvQ++UL7BmjTuhVxpQd7nFLV0LJuSwyT1/lTjBNsjTM7F26PjqSwuDn9K
up+c3aGBXZ4jC6snSvDZ+D+80v8MDUe4yMCRAbTsIq6H/3E3b9VQHmesSpQmu/z8xXzVxZhs4Tzh
N8xCRLB/5cWS3M3UbKBAqr4ZiJlcp0bzw5XStuX8QBXs3D0TFKcQijkSw7/sORdPLF3b5U2AjJJS
AsCPuIbyGuzilUg9W0Wad7VQZMDUHi3EkMih98tdx9qAEt97cLzPXHL0B4oOxj4DcuCmQ3eZmvW6
7ZnUtB1vLhpcTVW4rxGoc7aUMWUsG0P1zmwMA14qgWKJl/d1J+p0DZY/rJCxaKGKA6JqYobGKjt9
2Dn+Bq6jZ57D2eauTAEPhZeGehzEETwPTPhojuFgxT0Gne97fe6No5eZGf0Vhp0sUA2TQrmC948a
HeoJ/Nwesu84nNWMB1on8VNG8iHVgkSOTnN7NtwEWSdc175Usz130AgPJa4453shUjfgi8a0HRql
/cTjQGoerSLglIoAL6ZfPrj5vI4zmOvQHK/D1KPEFW+cIRe+GdBgEmpSnbri/wb7JMFncU3YNnib
O9UAFinErXinRHZVFyHfqsMHzg7dpGqU7lizF82cLY5W5AIuj8rIbi6bnNK1oUF+6CUKy8H9ey5D
pK42R1rG4bCtkJuR66TGbcuwVG3hbpY86OLRyyvlUn8LvkJRJhuwNcdfpsaA8tHrkYYA90KxpJG1
YBDKMyM2oYlv0rbvLiN9BRdjXVyDSI4gBVm12iUjG+SfQcw2U4tsNTghPxOlLVKSLyRVEbL7g7+U
bCjM3ewUQ7kEcjCxFEwWIX59ZOKWxFAhFWcIUt2cIKSkNHaOtWv7n/ZMRL6Ow2eNbC12ipPZLpn9
k1X3Lf/1OyNA3FFR9+F9Vxku+OmHo7wMTnYOxJH8klmUfe5qb0FD54MfWzuKoBh8rXuiLK5YF46d
mlY9tuVh5sYDKW8RGmN05EFwJZucmZMguknBMMc6Y/KRUEKn2NduFL6alToHaz8bjDJzjPYNdwIw
0iMdNpU2j8MxIxo8Jixf8s2ypR3Kj2yAdhJ3iL8VUReNl0jIzP5N8L1HpdYXUdM6EF0gqTzc9TsY
Km5zhX44canDNWK3GIpVgy0ZzPsqaTA1mTVrizIv3Wider2RkVTgI8DrAbVFJdx4U385EFUipQIB
WkKPIOPzHXEdmwuz+e18SwWMdMBqUnzMV1Ltx1JBzo91ykxPhmItkLlGoN3Cqo69u9vASqHtOtBL
KIs3lmYBxMGTFf9DL9Cz2zVfuV5bB482hkNsqCzD4KYzUiJeY4nwGbr6qCkw06LRpUVUhmKLS3bZ
zq6qlqu6Ia4/jCm1Nj2KVt8oxO3UTO9YqJs04FJqQFdjIyihR0HZLI+qWe0Vs7qyJZsOQ+zLVl3E
i+DAANxZQ3NnU8Iay6yxX5+XqGjxUg7PjmvQFi+MdDmuhaHwshuywaPxXwDbxlJZhBS8A5TQbaD6
1XlAXzp/sZAcB0mhKPkvQCSsPeVI6WostqW7QRBzr4psbhRBVs3+dEA3E2wrL8v/YK6pgx4g1vAh
ak9oChD8hh4S4FY8lm/pNRBaJ8iTXC5NWZYYqEhAXHNf1zL9rPaHykpxdLPYLj6B7QYPnZwcPqrs
7bM1bRqd5laV0kamtQcF48s9ahg52a6BCl0m5QkSV180VGUm1MXiC24I+vk2MpT9D6MBFmAfsVGJ
USokgS5HYLjy+9AQi35LnIarFKZHODhMleLXhthLnbIbFO2hKEm2PHid/waJyiB1W5whTvjOnW49
0mPYeS7u5crUDc1v2IgSAWN1XkEPKE+2cqyQpCfARFYYGblawSMkTxdnvYEDcISYb9Hwso1vwHxR
kK6DoJwl9Banvfkl2SFHe1W3hAiyS8f2mB/7j4wU7bIl/Rmt7ScFya6Ih/hextmCNSM3tzmXjVal
hqL8WQGLihH38plHKmkPpfcOU0ZWUmNwUkv/OBdAbwu6LFF/nj0nr9DgoYrGEw/2pTithFXfK65u
CKQyg0GAHJYc2/ZraltjydhAltstTbO/p3N9zjQbZfY5Q8dSLoywrvlYffxfM5PfvMTjMBR6IXD3
2RfmKbH4/N0zG1r65h1jvfvN70DFXOLW7g8wFFMp3xzd3+s8jUd1Nu0fNrjJ3PZMW15x/levTPsC
toFjcdYiKGNUsoF20G8VjDOOKNMdAb+tGoho2n6LxzlJ8xtH5UYucY4p13wVOwZUUmKmGNki+9OC
Qp/365Za2Vgak2qWKoAKQheDYQ0sMusmVkw7PMu7yMTXI1ZiCpazytUMzzIQL04DN7+ZUiItprrF
aowRGrUHQfEt09mkJ9wAdPSXDf43dzznMVRqFLlxzNNpIYD0oeQbvf2r1XdNPjbe6tnimL7Szmjo
VetQRLsMpk4WNe47Uk3IHoiGyYqP9rkNzRGEFHfRAxZe/2zVt/mjgGlHxQm3LaGWrEPhSG3ovUm3
eeiYDaUIMjwT2f6dM0qsn//B5JUQl+29MHjOgZat6/fx9wyMPx9fNqJBJGOSVwsUSC18LQEBmJJ/
4zUxsthAgJTlRne7gCnHum6rHVleJMC+4LDnY3E76aPMbJioA/iAKXpEsKgjd7Bfm/niLh/ZAF+R
nd5jqldVVyNiIbTFGObziCKd6FSnjetgG7YSakCBIpp9aIn1EoCPxZwqzqjHx0G5MBIAARP4QGwF
zp6yolVdSqWGo/TjWfjSfWiYRUwbJgQ73i0uCXQ6mzNKKLHR5ZznJyxElZp0d/V0csTHoOw7HnD0
4q21s08nBTF4pjTzVXn2qiTyzORuJPteFQ46oFmdQ1D7OYkjTFpWWiFL2UtWG7G70gK+KlDGli8x
k1BmZex//6caqob/SoH5zdzDM1/IyWyE+WKekDagkrHy0PqMzxIaBo0jOXdFEzOksMiWQkYoHVjD
4xW/xwCak2bdqC1JZ0xsWvyM/iA9EhshM8GWzTC2fczc8XjOuYr+UQxgLNNLaK9/7ygHnqYWuram
UcK12UHeCFN9wiDZREeZPg4d0Y49WW7ZFteaejbEsywJ8qVeoMTVbbGcTmk5nnMZjHfMD2pDVt7Q
oDrftxsPdFIUiVtXA7kJg/gvx8AvTA2wP41isc1gIFg6JvD7MoMJH/JSk2ssRw9Z4sjvPE3/JUpN
xNTnZNAloEvTwA2NT1asQyvQsJ7WhTLo8J7qlnxV/VnbOy1UuWwkMCDfEvnvakpadTJvgxZV7VSP
GuZGrMdLuDUJ1LGHseyObZzJRyi82RsGqP0ynowQa6dWTxiac8DUNwSeinhYppD38uaFA+9hjIEm
soLl81Wttws/e8ZjgndSjUTV5EXLOIJ9pwhDyQlB+rJF/rhSy/NPbLr/foO6TVAytdQ6gFB3G2dj
EXybPXuz56AgaVq3+PFgGSxe7UFDS9ohZa7cvA3dG6LRb7P/D1CK2nAB2l4TxHTbjNne8ibHVqj2
5te+4jJT+1oI7cptqWKxI/T9EmkHCUPHj5UTN9FGpvdCuZJr6jcf3wZr7bx8Q84vrUT9Xswa3Pp2
vm7boFgDcUWMuTk44UT921JI6dgz4yy2FcRALRGBmojtJ8dz4USC7feCvkyL5FWtSvV8jgqSB23k
uiF7MnukRPgGpFVtJtAecBGb8GYUZ3whpwDGxHnhtZIqrxFi3foqzaniVt/sHimCw0vUpExeosLg
L7F/SLcHfwh46SL1UrNdscBiwoA+2bQ/mYsL/L+w6fL+8OFDgBfqZpYUOiOI1jGnX44puNGUQGd7
lYQcep1asGfy1BM8KLIjcGJvNrOKRqP/enh/khpgSAWvAjBYkKZtvDxwwFZIJzbQTFdOFIVEfiCc
bsnNaNhyrxK0LLCfIrn92SJ+/tpL6o51FnvOdNM1rYuP23zPP2epRI9JsWyOQdNfky18u8Qq5CIQ
y8kLTnDtyZ8Y5WUvT/u15lsd7v1GF+EqeNbQ5EQosZzAIdoivUpcm5NpcTQzk/kqv3cSmHgaWi9m
kzGM3KCm47kl2tk+x+dIdFEbhaYCdZ6EemcVkCdE+Pyv5EgRKOup4NMVQHdjNVg4ofFUk6Q1Xya5
btUkT0FKbPEsfl0TlBIYOAquCDvAPFF+OwT9sse1xv8aE1HafKxRLUn77+u62smgYXWBS5LzmW36
8AW0d+oEyDM4T9Ksvj9B8OVKdBZOA8VCghsVtMOzheaKf9msTHfcPdzof2ocI4wsz69LSwy+sJEb
WGQuwGvbQeH24f48muQN9Mk3qKcEvM3Gp9Pjd3hMIoa+j7bGMvkYwk2/i0zlEY3Jp8V1PEDOkQuI
l2+xLJzXbmtLnEkdXGvqyW3sFA/RIHa+0LlhAh5+W5ej2sllCx39PjwBgdUInb4kn070+t3sOYNs
chxVQbJP+VQ26UxSvwhcEpsgSxQqFBblrsWyQqXeeBMbmKSrthJqEhQIf8ebuVavkB7BYbzthRhI
XSdwAhtP+G8BicSL1o4s2ynD0cIJcRHr1cjSVH41X22o8CZGOb82VM63jcjXKnks35+BYAYDusAx
vtmJpYjAMzIeyMaoJ0c4QTNGtUsWmZJdHTU8Q07/+6dGZ9XM8bvzV/2V5pR6dDp62ibpTBW2Kzdy
d3Tlz5bwM+6uU2y8o2qqgKSQQc2xFfM1sOXMOv+u6Nhsu1Vc8Fx6fcJgVfWAV+os/yGUycjLXUYN
BMOVqvZ6f91fIFk2TYbYLcYlilwAH4M5+nS32yz38uIoAm0KvP336YVLUHBw0eCNqFO0O6nA5ZQL
DxIJ/VWImRjOIc4OHRDGFb0Y3gj4KaE2wQJ1wSm436OxOFzrMtOs8PDed4v986eFgNvsCe8RNqHd
riCGhDOE5w3JBuebuhpRvVpXgdsdL3WL0ZXX/yJH3zIZINulQuoLm92CfEkMgue9/OO70ZwBzMl5
bqj2/dmlPgoBO9nEpIDYETrnvxlHlZVr0EJS2NNm+CS5FWrBBhzgjk5EonSkKUkK3rCS/9TQQxiL
NoV2a+u0gQ5BV/jXHfYFB0yflBfokU/Z9v6l0UKcgQHBjwCThvIdkPkyaL7dJCGrhBgsBrMqGMy3
azqIDviTsweJz2D0RBC4I7tML2aAFm9kF53VQdeoND+YpVwx6r229yNiXwcRG7Ez+5RhJIRvWcjp
kbw/PgIaJv615dkhj/MgDnd7Rqt78WEJjTxbC8yOI5/zFvvvs2muGycIioE6OmkfHDFNulLtf4fi
US6h02uBL49OIU2ARcfAub3yrEXv0ji5wqUiDxONDlVxbplVZy/ZpIDyrTOrb+/WZmnj4AR+rpVn
u2ZWjduqwlxEaNkI/lKM42FrbAOhYBb/PsKmzEpI4sENHYCiBfYpP6ZTM2Ketfxt77kPQ8rjnsTL
6dTR/oIftItwYTmdFnTzzZBHIfO2+IBtrggftEuf9jocMAIozdoNUXGUIyT/LPe6cMKLmlocxpVC
J4TRA96rrZYj9G9bEBiV8kq21/4PLtPVvkWGHbWxV/h9vA7HCZ6M5em5Wvn13DktNVc0dME2YR8a
b7RfLrye04ZoF70PAigxX+KbZtm7Ek2+ZCqRZ7Tc8DD/UC0s3LIx4wIiP+B0Gcrsg+qmJqO6Xvcp
UWsV7ZFs1QL7MZrmVYn9bQpeqXqjjKrjG1vaMC+CpaDDIx4sZe6be+51Eg16PspGmV5STZtWZm/R
YQqEYTYDlIOvm5VAKm6JeXiKvUMibo3f5Mh2Un29rQCN/lFnmsOxvz+eO6pa4GI3WOkS1wKL5105
EUgINEFEwFoikAvz5SU0MPmsGq6Loe6mvSyJaDYaTRifnQMW2wUBkQyvg4AwjS61DQt5wUjMQMZy
J6zui67nf1LWbZ8qUvNPv04DisnR7r5D8ejVL6J8JIXPRwHpnO36T9TJZd/GrtIuC1OEFIcjH5MC
NfabsRx1hJsh4ez61IRVhpvL89byFMJp2Uavx/H7MVjLf4q2ykXtuVCZzWP2z0rjPpr7OQ23swf5
ohxxF2V9T/7Nr/p/1LNyBaP2fsoc8QjS/nm8hPSIt2Aw2uiyLf76KbJO+Ruu1VRXHL/k23VxWizj
ahwm+4Kho8PYSGPqTmf35Q6wsU87BLz/9IWVXR8XxFfLujKgvWuaYfwtk9uW57IfNf0dE1N2cQXZ
ue5IcnoM9EaJaKX0avdJv1bygPhdp+MQIWnFPdEObno84+slFyTQUDVXTHSDfDg50oANoJrybgUd
geWmPouGRRiHxbJBXqz52H1PldV+XD7i8Xdz8IdleyZo6G7GpEpPXwyqeDB8Oml+VLiHVrXqI3+k
xhdHKVCyLP/PBF7Ju61OKus2gAE5Y5zgF9mic+1mMifa2B7LptES7iPbHmitAGhNZ40obmGS7uLp
r+GA69vx+Vr542TwLT2doHx64YowFKYb3zCYKkfOj3ZB5y9wHS7lW7iPP+sBrMUCx5tyoAKV+o8s
qxkG6y5X5pDh4hV0eIGlBdiUjvaWJxmQLuQIObo3XoA4tEgMvZ5Nihvvuhr/DRFX86zPV9rQ07P0
16zT4rLd8oKx62BFhAhAdqhw7eeXIb1HOZYQ9RhisSKycAtBI4E1fq0TyA4UU8E35UHO/Wenubk3
QHwImwfKC4cC8GSe8HAuHsT0dVlXVtQ5rM0GG/9rdbYG71ENoMixWWrOounx4SWw+H4p6U2xo6R8
4GcQ2HWCuQY+4V6iOoAyK+6bMf7Dxl5DRgt6ywOSPJj8gVMHP10bRyy+E1O5/LuQSMMQSNynN30h
F58/oRljuZbONRzQoc/xn2i13TvN1h3bUFE/sy9/tVWRrfbwn5XA2JG/NJk28QLrwFvozXFRp6jU
IebcRULCIx5mwhGSD/nkBtUsazb89H3VbLv5ju6P5D3NLmuOdrmtnpQOQWniSWvvbnUYl5Dhr32n
yapM2g7G9xcfihEq7wawZeZYWDrKx6OuG54n/DWjyiUy5tpkfIDnNSf+4IwxfbAGqY72KuHFK1fS
eKVMeQHTHUr/vi7wU2qooiMocG+KuGSudWLfCUDuwCi096oyG+4L5grH7+KYyNXnkSERzuIG/Nt6
N1fKcx8HmPrZf8v/b3n3WwsjLcUVTzsn047lQZxCLimyHkhxPb954ufbwwRPfxn8ZuYzXNUDfMmV
OC42gPKFUFIFJfVXl+ryPQGP9dL93jZDpHBwz/4LvMqF+a6unR4gfx7IbLNkXiCHdmrRZGxim/cA
4oiNsXtKIMs1wQ0fWgh4Sds+gRhP3NSH8I5lhBfbl7VzRPFypYJvmvmUh/TYby9oSf1tW3BELOim
IFQYCoiGhXWKFJpxuMUMj3MDl/fwWSdTtyc9gWMpKNE23vsn9uhcqotx3alo90vcbWyHadnf7DCY
m6r5UqWFidFhYFVxF4Nhxc4oAKzNAN0TR8dkoh5wILqi6V8+pqSvLnnWy4FneOGDwnFb8Lm019Fi
XEcJn32OwcqJT7HLEwdYErNmDh8kEX0vjaii8b7Drfc5Q/rjneoXZzdcYNj4xx/rVypsRqT2hIQR
taoGPQa8uapM87s+ZxIgHz7FVcQYvTlAhweyHtzmPatBgjE8eZHx4EeGKcLcV1sywh1wXsuwdqtF
O5y9lKXTsLxnNRWjRiyal5u6dEgMNuYmE0YsC586WDZQwA0kFTqK7jYkHs4WkbreyEU97jPh5w4j
guzTtEgxkv7ER9HLMk0apaAzqQDnwoi55rCoiYsO3mcSEzaoSI7A1wxdjqlRKps9mZrLMqSV2Ym1
MQG/y20NBfFLRHFUq/gnFXikb2fs9T6uLNzQZAJZjSb3y6z+Piy0wNY0awpZ4tLJ77TZqvTT+viy
CV137nZ4bZcPGwyR5rg2H/6MsW+hJk90eF3bT/neguDkdgKpvulXlzwOBJHpeqMKHLxrVq5w3AWY
svxoEpTJZ/I+GXuF+wM8byqLk0Zk5IDIFhO1XcTkX17IlfOD+0ib+KtJcXoJRGX8EwLI/MUZqFTJ
+uFXxXGVXyUUPbjBRgO1FO4Y/pkRPaofJvQhXSYT5FXApAs//gdG0IYmTPis4SttfcSQi8ktCWAV
JRuF2zUBVmTJU4c9RQHGBD0+Mffz9L96vLkbOqr2OtKyVkOfEZM4VbglVitar7R3U1pLIEXPEk0J
5bp/+WCUHfoKAs3Y/0sFSDlkzamMjUQS96Rma5YqXr7X+7VxctPZTzIpBHznSJonrqZzILUA0N9t
+AvheosH9PcEL2NF3L37vurR3OeZdSmM4P7EkBIRoDTKucIPD7/nIO/tmhPR4LxAve4HhDlqTCI/
p8FxpprX68l3Hntw8SYBR74+CihkGSf4mKzmaXrecHLmo23UDQjonzuDHLWUXJBiJ4rjFftBS1lI
+hWpza/oqLEEGihTNckyGI2mywfXw/cgMM6wFvwCKwYkkVHifCiVg06no4YUmLWGMOBg4dNNN/+d
coK+B5IdDz/j44nX89ibTA0RTmBx4nH7zsKATlJ0+x5TgbHSL2RdcDxRkuEo+Wybfj7Jbxj/gHYL
blcyzn9WaLufX0aY81ahs2xXZR1RPrnZtotK5R1eH+fNJewUQoNgLRn/T/XX+RDxS0jY1JYLG3sr
LWuaDY5XQ34t75ZfYBWP5wC4qgdPq82cJjeGcdWWHAZ+lV5ZrL/fPdj7qXVV2B4Db2XYqAJraEeD
qHLphBliDwilWbcUpnHpcPYau1pHPxtJtaFgx/Pzx5PvM3IORtVBRTDOjcx/Cbw1flvQyR9F8ov9
K8sRGouNdxzgEVKmlyh9ltfa1xfd2JagXdiStVg40Qd12cc+QBE2M8048Sac7U1We3G9DLLKs0AN
PaNUVOSpVdP6fqf5oFRradY/mfxgTtkwSDK3KTkor4O69pLhh5LdDXrA6YJimjzhrmx7rFb8/88R
0TTDFh5T7uAEbQxxPJHR6LERHao5RHZfhdkmvHP0ACuGKaPAV6PMkkQUgbGbwiooP0iuN7dfJU9f
lfrZ0p40aUw6W6QDAInseK7ORz5Dk34gTVeIKe7fVg4VXUAsOZO3IRnagwCWbyvSbersD9rCMn7o
AnApYBbwNo+e8wCfcOW2t/eFxh4CqTJ4pAQKSawnIo/SyvNS7DlQEoLj4pU8OWBF0taRT7/7Hcyh
LSOeOOHuKOOqVtH+hQUv9hKYPI6TRx99mCf8F2mLGPOE00rifDMni9FyDnJ+eUVrBRP/cieKDZSY
kco/1Pro5YA5golq24FAPkOidcrP8kLpY7w8ssDgHCZrhkVAblhNj2a3BRDmOOP2UEPb1/DSjZGq
74y0VF0v9mj7TTIs3TBRdaj3ANCfrkH7V7WpF9ADf77B+YmgRTVbZIu1FMFVyJVOgZo5b9HQj2ez
lbP0KjnXGEHr4OZZBtjxPkRIBRCwChuJ6BF8D+ouXaWcB188bM+tXOwTCC4ZnbPClRVhusRX7De/
N7DCb2DxDEPvwALW/eDG6vQ+/XZJuXvtHxtqqczCOxMxDPllcDKFxieFpyGc381xoNtwyP2I05ZQ
QSWhOZLnVhulCtpP+D2OwHkEqDawZrdl9WxhJG2e9qsnYCkCFnoZ2VhqnS4vlYzRbLT5gozzrpSQ
R5tYo2MMQ7CKpcdrs6d0GXOTi80tbL4n99Cb9NgTwYzZg/yE4N+g7dneer5kMxKEue3dvdgbwl0n
GfMEj5rNJiGVSeMQ5vKgap8gy2+im2KNo99DZKFUiGrLlHqN0oMAaHfR8KUKL6nz1AVPeKQBAiPE
5zN2KFhyJFavQUoa0eYXi4I+/rqrw5XFJAN81klsTnaUCHzvKo8NrNPTjKBlmCRNn6z7TECu7DrP
Gl4Biy9wskXofQwXP2WZ/d3x5LhH6coym/kjqHuX9qFKRz1icEQuF6ENDxMNmSfV/qIyVCgBYgXN
A7u/85wreeql+k8Ozn5E+ajWaQ7JiyqDIKVWsK3jXtVnqYEy13tRpz4h3D2wW0psS8n0w2duQCUu
+yj/Gzb4FXeJRNnjpq9xN53wcihUad7ZbonpYLcKJmkpNd8BXvw5GXePSj4tx/tu/zshaYB10cOZ
SWDZewX+LLxVfvwha5LtKJ/YT1jKZLJUomPVfNcOI5k+DmUKxq/utNYsb1PU9i8rfq5S+EDsLIG5
2JAWCNSB2AXhUHYkxx1rYXL97rgiSCu64KZlOc1ONw7irdqEfXEQKhvcnLCs8ypMhoyoXTVMjUyT
vdcfEMpQnmtw64V2H2jzIsh54O24cUu9px0HggfmQjPyjkgbfjA7xbCDU9ZDfd6ZoPLAlgIr/3CS
t7QJsca5T0b8cbk3vtDJ46uzfxX62GNt1DyW8XwuTkFibmKXnQqvuvN7VS2NNqJ/wcbbA3sSohUH
ps50a1r48KHJBmaLcwXIY65UrUvpI9I5EQyQSkeuLA4J+6OGovtNnosc10TfZYEWJFnDbJtV6Xwp
lRMqnMNKVx81SvvIwHPZaHT2EmhNbEqaYegYNkwmshKXxf3MTCpP7VX4VVvue1umYyOEFSaIvqhL
SyUac6Z3TMsMPWrCLG6d4jeYQXW6Svjyz/NBA0rPW5suf7hDTMkKx9NTjLoStx+X8i6VFOnOx+hw
c+VDrpUzUjh/MRAuOcZLszLQHpZq73DzznZsj0t1HWYjNC8j0segPF7TNeJz0beIEa5ZfoVNk9Nh
QXHa0bdfkObFwSlPwCfqvAnC8cM4RDGQPAgCMEGOCcYgQyt46342sCFnpTgJod58AHT2c39qn176
d7A1Lr52oG/u+VnijPrTdwhccf6gk0DqLN7LSnX7LqiMzZ/LvG0I4XE9WTXs8P5S9O6mx7vZTxYI
vRTKWma4QG0Oct0PRFebnNJ2t5LUQcyPiqmhcL6/3R3SlTDnt3cT8dWG6FfZb4fCzdkPKYTEam04
Pqsgafhxo2kZvASb4WfdsJXUzlhzOnS2e44lcy746S5xaePQ9SHZwXdianf8c9w3qw9egw4eTwEn
Y/aNqPn9Y2TiMG343C1eAoJzXA+N1a82rNd01ZBlCudsumO7UiV6q/s2qdgIEKCypFoaqNn9rQdr
dGnQOxCyMNPG0CzWeeaeyjQbuENZR76a6hgfbQN7UMkZosuEij4ZsufwxsO1WJuuDKpR804DEcLL
9ZunTSbZAGIwYq4pK01ZndEBb2EekAZHF7ine6xD9lNUWLfGCq4IYnucJSoUg+sO2ShCFS5vKwil
DxvOqIEfNoTKBAdvL7YIqdFVM7s6lAEjoxzFK3NJ+eXMPdvwA85pfkhhEW6j+7FX9u1Hp4yECzyW
64A2F8w6udHZ1a2Q4JbSzTQjmpM5zh7ULkR7G4Nc3Fc8x52bLDyXpU5inY226G8wbP/n/3tzXuT7
yNHvCYgw6S1JofbFEUDV7hkj3Yj/IquM07u7IzQ42tj4BgDwp3ar6NIAX3JL9OWCKSBudQBhAISp
cg60DpFq9OwDJEcjYTxjhjOynHBG7kDjA8znFbfYAyg9ptnrPKQcAyE1ArES5QEKPnqNj1ADpTG4
aah4T63ForpDv5fvyhpRZ4POkElIhzwWsQiRGJBbpTy4B9LBDm1HOTu/OEeanKvELA1JNyWmof8Y
DbAOitijEQtpXfMfhpuCneWVFkKpiq9h48diatFVbJLCRXORzUPWJer7TBSSPZGygzUUwt34sxg8
2dVwV+uTQ/pVzxPJptSfYsBx2x7g6/S+1GEWFL/gHc+aqJWppQvH1TaTmPEYkn1vfjRpTkWK+hfH
BcMLQbirfq42j40JQtFn9oAlKmEa6da/U0SzvbIIGcaoa/YHTZP946SaF4eiLZ9gZUDE3d3ByXV2
B/On3NnxDQ++bXf7eCqFUNhHl6aVin2AFIDMfxbwaC6uijpP2dblPCcA7p3+5LuWZm5KMMkoazqs
+4vCjnJeMHNEM0FQ6vq9jvKRagoT3Ytb9DX6SQ7hJ1ayCwLO695vGmCAQrerBfSm/Ewoht4h2jNK
SXEs9qDx6PaLkZlNXxjWeDG16Zwv0B8J2phgNW490gF3kkosh+yD8aAP3K9KdCxoe65ZqwuRWv0U
Mt0tZxKII2U+7DdGjwucsFQ49+C2pxpFhZpjBnirWccuoOvNOG2Ur4n5CXL6Ql95EmjcGvHq36pR
HsSckE/4BeApNMw9o8Y+pEbQNgDIk9ktvPzgIHuIes3LOk1tLLGz5nbRAo8DC6FO3d5sY0WFiX13
EEJa2hbGQmSMI56Z0XSg5iIZGiR9NJ9CZYFXNZ23F6gkuHUsbm9KKO92Mwc+ZfgTBDrSCM4dKrRa
dOHqugN5RUsfxKO6lEXp+mQ2+SAw6JTRnLh81hTEikuahpKBbbEraae0lToocK6/4eMGzHULeMBQ
Ri+NC8HTva3xQteoqUoiyyAINr3G52qFca5nYNAG4HskFmJ7Fv/hz2FpWvi+FF2rXdjIp9aY5/QW
Sf/Gu/9UC6B6JHChkeqCapA5w3b0sdlQsH9yOyaiNSSBEAs7z2Bno06pWClyxwkoncgf5bK2sY44
wk5WZqFMt+uSfBQ+pW9HsXFM3fs07PJwpbyJvwRNgYr0CV2ZbBipW7T9E4Q0ST7oXC7S3EHuZeKs
nM2xrwyKmqicXMRNkiVqrmxTtFD+1tlXGbGQ4WuaDoXIHBQbOWkTrRaS3J7QrGwFdSwqLuDkO70B
xYI7H5mpbdFwFjpjqHJo/N1q5zXOM9oUwTq+OeOCN6FpzxFqQkkjPFS1TLvfD1F0/8YpiOqbAgM/
WegudVEQMRQv9Zz15ZJbQmf1grORJlAj6OfCNX/+5oVNx1v33CuoGz2nvyIWyGoJOT4bza4VPNzB
uND6HqTy3ydFXk48ZQThqmmWG4FvS4qxiLFeabmHdojGCHQhcUQF4b2xHdT2QE3CqNXeZ5zkQkoC
YnaMzzdjHZOXrz0pXhUqFjN/HhtxQNBpGRwxXvjDsk2Zmk8+Bw8ivjnENMqwk/phOcbSCG8DY7OG
FQe4HegQN+rTS8+MrvSAZjzz92Xtbsw3QfcYxMfWsjJdMmSIa1D+IQXAQDy3xsAFdy++MRIFcnxx
Uxy8YDh4PPhj7Mmg4mEOF7Vi6A2c/XouGbyFgmVEkH7Cste4eT3SfuXEi92VRs5omTah7KKKGx/d
ioQDREiuR2LLrs0VVrvjbTtBEcQVsXmzBLKRjvYPuN48e1fK1rxpT3D6ZhPPvBGJUEDFrEcycDyP
oetoiV5AxtJ259VqC33+G0o9KlfenQZOCoLgCffNDPbxIskXyKBw2yI3PXmHyTFEwO+6C9nF3+IG
LJHxqyXGvp19Zf1AlTC6rDaWCt7ei59ldOvKBibnzpkCj7WQWHYYvgQYOhxzlpARkQ8DHoNJCtXv
YBdI2MD2coassWi9nVkIpzs2c8vqekcqzzgNjaHoBjcgohtHiwLTkONmcCHmnTDSIT7pHFeXwv0r
6E2wTjXnCx1XNPUmBy7bUWdAuWi3GyNZcRxiIiot0irFlkCgiEGJ7DRBq8MzQt4TxgqAZPy4Djot
V+lxoc2DFZNJ9gwS6lqgWQGazdq8Ts0oPgQ3kFfnzQqldiQ6P40qWXv8JkuXa4lnM7raIfPFY2jd
w1gFQ5Fm5q7SoRig8WcSkcCfBJr8qVu5WtyQ5lHeshTSilirPfKJzhQHXyLqOGDivwqbarx9X/Ca
QMC6Sl5yNxXq9Acu9PApx4tU1m2ZTpOHSOSthyGiu+tCKILT06hBsJbRe6t7J0thI+exoDU1wPXY
Yzm3GbSfZd/GhnCduB61uDIF4lhAjwJ/EgTREhUFwzi1jxzl82+TtpNPDTEWggPkvihI0jM3XvxO
EQGIqHVar1cAUbIO9BHuPUBk5SsEKC9H5eIbXRQ0AbcEVm5bDv3HcYsqzevFI1T0krrsRZj1b85x
5xuS7g9X2sqgz4wQcYbUQoLS7Jf6Q5xmiCXVwbJT5ZCvMsN3hSK5SmivrxfbyD9otniTiTq0HQPc
jbn7aFFcFY57ZlTBob+MzQ0G7HyggvlQKEel7OZCH5/2keRrYbKhp51/czZpJ06zMOo9f4n37Ogu
9QAfpi72lRgAUdFfQ/TIzI48V4Lg+j/pNKvInsIr4WQRr0QB7LsZy87B5LMsOEVCPfURbGPQaBGI
L6+qnOvdKbnVaFR/oRs92ouyuKcPOnoA4DhZx0px6Qsy669DfPB3l8WR093Ng0HKJDmfJaq1uAKs
AEvYs9dvx1W39zdtbIUl8Uj0CARplGoCzMeshQFEcA8lNTULgUHjZmNHsZvNjuX8Eh4rtGeQoOYN
VCqS30ILdnYsxruYYVn4/j7Yq7s8Yox0seFc1yiYzPsv9YJ0KhjIYZojjkayfRV/r0h1P+K176lB
Aq+ZEMlHiigm+eFpClL3MCrK52mwqMm5BUWfz9q0wz5z2K8QrqFncKKwUphJsv/s7k3A6nFELXgS
l8TmDy4vlkGleusbziJmTFrtYG1QQ+1lPqqsnVj3wk9gvsDQh5siergoLdUH2ZSPG/RPhKdZjVyZ
gk0IokTxp7/Li3eaJ0pxjfKXtAYIcIqxOV5Q1wKb+ZEVFVWGkhnWoLRxCQ6oVsxc7CNOuqMvtgvj
R1ikUS6i8gHTBKGAx7gN3acpk0xER36w7odLpr1LT7w6lmwPu+tUq2PnE6iYJj2ap7HpCqmWJUJZ
vuxbVFUViybXpeNqoSnwS9gn3dGDw80FO0b+1Drv96DxpyOOozLQG82SCGlsIZxo6vfqPOHhNb9e
c6WtMKRmxsVAB6PrzGvwyE6irlFs+z2xg/vT/H8neIZ9+aRbwA8PdewVsVARpTxNh04MBJ7NQN9z
Ehs2xz87FlU2in9LqXoiDunpMGGcghs0g3B0+9KyWZgnTRA3tqXHqvV7PQDNhvMMYCwvBnYjEBg3
boLj77T/BUR0MEvjSdzdgkuQTVFGqQpAxI+SLViucZVoziCe+rOOyDN2/SEIjdyC8TBq+tfnb7ul
NXqFBUu/8ARTHYZG/iKEoESoWYuArResrNCCoiKQLp2k7YldhJTGzvN5PaPZ1Yir1oju8VEA5Zti
MF3PPhT5sIpCry27uWZGWhTV32oUHOgeSi2ut2xTNQ4TsXNfsvcyionuhGIgvu4NikJlekIQZq5t
WRKVr8oh8KbvRrAHcoO1Zp8sG2ErO0aOgP6FQqssz33bSTkRRAxu2hCZKSS+ivMeBIy6WsDgiiMq
AU9cB7WF2uP1FY9Md9kCFru8gb8sgCaQG0LBN6kK3V72DW2PR91BGachZuAtazL1366ptGO6j3AP
DzfbfzYnWk7yowgSJEZ2OOmCl8yvVf6Il2tkP2j31zCihCTVPUnD71MWVvZ13ay9U3GqzL6k9yO/
rkNsuLPSKWywcqPkVOjFs6gOy0rWvLL1bWlP+4g4bOR2DJ4AAFzylBPUVt2T0h6RePq08Fbjd4a/
PQgcPuAKx/eJvYU2CftbTw70KpGd1oqSBlzs3wKDh1MOPvl/mGh2sl4/083XdWY3jDH+lW6ezfH1
9UL3o8nF2Amh8HkNJEQFesoc/H+pucbGO0g5vfi48WJJUVNimpdThsziAyxCOwyfQC5PByIil8oR
t0EUjsWEFlLoUftM02/Lrf2MhtIa9Ik7rZ2xnyhcmgaCT8pefymomEfim95udENrAPT+iNUnhR0B
pALJf8byTGUUzdCrZzxvNPmaz93aw4yxf5t5l1D2MVz5sq8nOoKGt8pQOGko77DJuxKfsotPT4/G
EyD33Xj1OBClyhiGqvuF0fZjsc97wvOnEpCRvNodr4f8RawW/AKSfMOjimFUgd8xMo5uDSA960Kt
utKdHY1GbHymIz2I4B/kT/0IowWit576ymB4SIIquYp4V5qsT0yjBDwmcmP+4l4rVypFUif5+UDW
9+9A+/XppPkS5edOpBWMusIixIR9BafKxqoHml8Tiq8CGqyUB8zPDclnSJ3Tz+x24qLg4sy7+0wB
VgmzhjP8Bb2Zd4BjVX3aPCLLYJZd+nxXRtr8moiZ/D216jpK9J+/y641G8iXluXgrUUiN4dhaSKX
ALOm0YgN3Kmf/cnPnjXkINiNPAm4yojy2WIoVtmxZ8Oky1C6SrC7QjQqShY7dGBuo933KYp52b/n
9JdFNwNsl4VLhHvpvjg9f9aW3LrRn4HNutYm+YfSn+M0P2kub8o5YJzdHP2kvnkUclAYP//49Nb8
LfVsf1dsO1HnemF4PIxchoFE4hzILUaaCuhixq398xZF6ALim8ZuF1CzU36WiBbYGs+IUVGRRYq3
MahZhRPgQxLWqiukR75q9FcLGleCQlmmNu/+6hcxQFar5ex5Ntt/DSTQ7yojh/FEhu7uZZTbZ2bv
EyNxwG4uuqJlJlbNP7nFK5EGmIR5v2H/KQcxkx+nN/ubBVRhLMA0G62pHpxzjq5wiSbhlwQxWv5o
M9exosHF5tORy8iZh9EBI7OGog8H2ZlNaOFdpTmnXGz1Gqb8Yb9BJPjexrHQ4YKh8oIyIcixN5s4
5Spru20X9kNyHRf45DuDkhkB2e3/Ovjt5d85iwjSaYHwE09V+ovm8HaROF/aETscc4ZIX2R0y4O8
dV8Cl4X/suAyGegUS6N7eoIgQ9sL9Tlt+1T9ZpzCPvKRHjk9YS/UfqP4TEBNX61dWZ7pYo/+MlTC
PyrcaOadxKigbUYEAxiNSSDt+EyBvdwlNZmmln1KrF9InVJgRD/6HMZkL6P78tuO1oTgGdRaCtcf
RnhTouV97zkWEGQwhxtheAPsg/ee9PBReIkJxuwmf+LwXWnQDt150TzygGg5ogDrrZ8I86/8qvTu
xoCQVhNP8RwAFOKYlpa/+by2GM1Ff9HyP6Fq0YVWuncBvseVJdhervrAEVizlR+1j7mZe+Ye5f6R
bY0yxTBhJX/6LmAkqpMsNEUvVG8PD8ztZHLee4SKGQf4nczsbqXnZFuzj+RyIUlYRCm5gvFBMZOD
Y9UdyZQ7YhmaQXM3/3P4H6nzS+L9OBNAXmBuD23klX4I9ZKFL5NIfOqltRje8XPN2ODhNgjxUwXt
NnK7924bIQe6Pku4Rs37P8cDN6aC0cn1Lxyi4hG3bcaSXffYvqdsDVRHUN+EVSGOuFjxqocg1b5C
bX3EFyq36X4YUTSChXAGXkfuAf9HLjYI3+0OXDc4D4wO29QKQAw6KZPyzw0gmgZqZMwQKP5wdhEj
dNPlwywLMBs5/voeJRchZtICH1BqOXz0QKi1phDsSOkp0AH30RQ20xNSTxUK5A03+5W4Sl3hUBWE
+BGagcG72P4ZTcoXJYRqj2qpajMYivOm1re6nyYrq2AwSV338+1wg3pwPeG8iQbksGctGABDGL6Y
FwEi6MYNuEtMpAbVtcIvgEcdX66AMwhFfIpcZplVBWt619XQyPGd/3d6DZ127W4NjNyyLjDeex4i
5VefmwO28Pw+T7W6eiPqfF7Vuqt4aTbbVLnLXBzLZp/LI9Lu6zvXeDf8upeaF1VuzxINJHWa0hVy
c/C12RfZEXe/cczMeMilBzpYnXKmED05E+zQ3bXK/X5qgguQGbPAnHBDrUdHU5aP1YjMCfsoqPTk
CrtR6nTdJtUtCwDtAy3IhDcJe5ieHZXGYtjCgbwaW2CgYlALvsw+2M38VNGVRHAsQao2W9zIVC7/
N6xXIOGrOhbdgpSyYSJPU2x5ZMx1PteTdMREObG0ATClYi6inPEXP07OrkLrfkCoToJlGi0qm96x
V3l6IyXFIAF9rbOL0+Z4M174Aq4sGiLx4pj+EGs2qoCWgmLekisRXQ2fM7W1SZPdyNIT8xw4yZaJ
LpRwOTTULAkwWTAczCYsEFsHTS3HcN5nt0zo5klP7yLRGqC0esz00lRd4QYQKeSJBXqI4dZG8j2a
9xennHOgQqU9mNA4Xr/eXK7oveJ76sLapCUVRpZugtwQxBiEdJYfx3G/MR4zJCVroff2s/ZOIjrA
2f0GwqgIY+ZhT7DZGf5GacgnZ/LOxxkjhCSUm/qF89/zR92oW2T7ZdhxRyRy+BTHeVYecYdyzHJD
9bMYAaFyKAxtyme3aj1rnO61TigFgp80rSsr3IwK92B6MzqNdWdcNumbLEhUf3CAz5JqDEL5GxMT
IAJ/w9Gt5BSNpQOEnf0Jt6g6UmehIdX5DqskMnyYzLaOvPJSCEX5Lurt6eLs5KzrHjYyJiHiYbBI
6AKuz2McleGUmNF+NGp1gXVkc8N5vfdSEm23NyJ3LnnJi/WImyoIC3vUk8oGIw2+AcG/1CcqQXM1
qK1s4N03WPMvWzmAECu7QX4Urpd/lZ2wmvEhNICb/UcjWtcA2XRIjq0/1QEQeHEoA5BJs5GB2t+J
mBH4BEAV3kQXONCq9HmfuwBpjh6g7q/A7mYLP/dZtRR6u+Tbnig8mbZkFVnOYU9GYTVeXu3Byis+
fEJC8rLJgGGZndiAOPCH8zojNSIfHJngqUl7y7PxTSgOa2Vx8BVSYrPGrnNiZI77FKXc1M8U+VXX
VZ+2lz684N37DLfrOK84TKSc0RZkBsjkNjhqfuoVZCGVMFnPT4EVZuYdjSIVBHuQfREOCv5kkxV5
9+T2XMBrwtaZkH1w+dF3H5sP22ST0+b6D5Z1ft5auiGZCOTAv5a2XE8MFFYnNrPjxb5FJMzFWkAw
rGphzXuDUX8TJywtEtzFD9ZfTKQZumW7+78F0IURrj1ZeWqENU9xXfFzVkAm3ADv4D2NiJR27YP6
CLoCFp84Ekv5SAwsoEblpo7wsd0vuVcW50gnZ3oTJvSKZQ4EFHalCjDEZGGC2+s2UeHSNrU3tkJy
9U1jo1hCO9+koUe1vfSjZe0B4+HwAEdeYEvzjfq93xr4Zjy6ptAKtO/gNa6Ybm+5hYGYdqW5JalI
jG+s49fG3jjoNVSKXyqn3uFSPYW/uVKrBPeUNl/MCXnNhGYbqgP4Tfsft9np+9h8+Ft/y0tKOlQn
Kkyy6NYJ+DhqhjTVS7Qjg81gnoG3WGra2qDIkOuRLyvT2usYG5svyRCxP7Puc1JmrewLNNKx/ElB
LAHFpjT9OTyemW01BCnb5MPskRdW3NRTaF316SpyISAW2LiSggrYz3O1VCzOpEWUOBxXiRNXJKFu
SFTN5pDi49mnX/7sqWrc7FqwZBlSLcrqydWHNhMPAsumwi3w5y3GexzEWr/P5v1QOaaBIBL3HWXO
vanBsHuBZx/WFfJjmagBNrh6oDk82aSmCBnfvdyG/YhTS+CRJUoYn9nVWu/NtZ8sXPcDbqZXtbfZ
S7US4epkxmwdZX+8TlxxglE6Qi+ISY3gnIoZjXZtoog55Hoj7/bjLb+7jx0lKx2Rkv6KzQwFopxI
w1gPZ5whZKA8h4PrSLhhmTKYBqb5mUnZ24l2Ogcmso7pZAnSRuiAIe0CvVF6NdrvCvLgxLSNF409
TOWaZdLSqTZ+rlc/WKpRch0Vi0nPiWRVdYxNh+6t0NSfGc7sfxfPgMZlvvJJ7nrQlVwuMCUN+4MP
OzVo3Cb4baIY3zXCjmr5HwsH4BtsJ2a3T/DsN8a1+uFdgyzmr0xCz60q6EoNnbZDDOqWMA7LMzZ9
x4uqp0TElTSJNW0ZqYj0Qg+dkthOQhCw7p0r4C3ALzYrSGlBYKcaz2cYoTLWHWMHUHV7jnJRGQpZ
QxmAiOPpm3Adb6i4x6b2p6U1pAZos1Qzk28OCwubzrrorVgT/KmJEWHhj2hQaciv3BYAi6UsEpEJ
fHw8Tq3FSTWd2XpAu6M+Kr9pGccXULTJlfaTDG42dh2SLlkvdl2YIXIjFEMEI2EvxM1fYdifO7tD
ibkDwIUevcyiHOc94q6y+STE9KqjDIswWAnDIoWG0aOqQz1pqbKhSgK9CqXR0TLWIhkihr1zS/5X
BGgfcsIfQfoyK+DXl4+7W2QRxtPV6ziIXzYGkomiB/hgwNh3Wy1DH/Optqutdbuk1osWvhx/iTHU
9660le1X2tQUySqLKbosuCRnPn319Ux05USz8qkmvtDNbSOyi4aRViHbXxAT5q53yW2bBUst6Ihp
3nnvukxmV6ZvxYMO+8jAgXsVv2g08AmnJuX17PFwMuqbJc9hDFuFXBeFZXWJxD6Dyvdzuvfoyu7u
4oQzghcF/DeucgjeT6a3UPEspyixG/AZQnekR0hl9OQ9WfDEpzr79BiZ7YHvIcDVWRA34bqFvZWr
+kQcIeN0z+AZDKsxp4SErrP07lK1BA3DnhbY6j+GgsWX8Dd+J9ErvDe9yEuUNYmLmYr4IVwj5ArV
X2nMyxdU3cXk88Bo4k0CeDNLfFy1n07Gfb/sNMwPKMjjnp7H/gQtonRiF3C8KD9Ayj7QaTl3UyAk
fKYktOt1gI17i9DQTnUPDi9QPKUp2dP6SyYFZM8aNoN/yaQjsLipXPlmqzpXJULi2NqK+LT/5cvX
58/SJ+1zKJerYtVhmLtL9vleGFNDf4RIo7ljSAnCeT0HLqNR+b+OthY1UXk2wy3SqWg+fZ/BACA+
OUdVBWw6PrmQ1HHfspVnVodjKi8nJG+Lj/FqxR64fZs4799yIJM7XubRKznR9oOmKXBgwmOkD7Ad
s2VLtEitYjoHxUDpwGnayD9LsmmV8AlRyhMq5v/IPBP/6wmaIBQcKNZdgQSdkunIiknqg9k/aYLy
AQXvzEPxbH1IMQSEAGv1AVglKOS9S5WechGCa5yMs1/NHM7ZwB3QMGjIJmOezaiLHCbP2050yUjI
xEg/GGtdVkHonU4FtknEUv1XVjQDomvvpSKkhI2VWHTY/wGpBl72fbDPYisdvfdh6Cwd/q8jKsMt
KlAETz1PfdHTiPZMlbqDYSg0aIWTt8rRnz9I0R3t/exb3MIt9LpSOG6U0h1mPjuVGMHpzFPTtCiW
zijvFMJEp6Z+Wpt9FUayVsRhPYFSvM7SJFN+yd52mEal6IiWaUb60+dpeHff/++LY9fVB1om7pk5
MmDM4of2ERVmEwe4/G+eIfAQmFnpTcIznSDS/RTTNGGih0Sc3JKeJiExrn2Ou1zCOVqBZxlo5PAE
PkltELgT0TcBJFXZKUFEBnNssBJRkB3u7vRYWKVO+Eu+ePrWk4g3jYCQLtt0wCGdijhTMbOnFDkb
eS6dNYqQ0yYvTPR3mwgRNEPYr+Ov9kuLzFF/w3f2oua+IeTwbnDlZTVPf2fQreZBsLhyR/+GyZKJ
wVDG6YNRoYTwto3SMm0BQCKrPp7pOwhwnI/QJ2Fk//WvcfpjgWaDAWeLv1oaw/K0R/mYMIYtZzMT
qEuUS1Z7zBXgK8x8GsjRlXawMmELISpzFF58PQn8H8ou5ySMAMi6zCCRux4FozomuiZeyEd/IsCx
0mHmlAEZmoZzYQopRyIuwOIwBmVogU4nsLjgL/CEgNhyB8TyX/4IPnBuEHl5LADJFB7S0DjoN3RR
gb2rrO+Np39o9Y3q+M9KfsfrnqHOWlXNa2sy9Cn8YtN+kFW03NorkTqfNdxLuJ6xJFKQTGrOrTe2
0tRFC+qJvjrrteW1BbvAOLhZdJ0vDlLM4lkrMRbrLTFP/YF39SqU6Ynxo6tGciUwW+HWShAYOJZM
ozZG+6LXYe+u3izvn6gLyxzum2yMd97MsUo5AvTupilWgmrxPpnMUwFgY0nY5oFlfH38p16iU//K
Sa4QxZ+8mdauYyLo6JI6jQoahUu9n2/Ds/ybT/AfZi6gEgUPPfhbpR6PngtvYUQnV7MJgRYtSn+j
itMu4cDuEv1lwaNd6MAI/v7EARgo4HGXfTRIP5vTkU9DJJhUYVCLtNlk2HSiMfXvn2HVENId8SBI
EspWMFg/7U7sC5MxVtT18W4dO3CrqZ4Xz583HbSV16tVGOwJr+kDcxGaD7UCjVQZNi6pIP+MMc8S
UKN9dUUa8BMkiJurOwwpyJo5VNNz6xWzuTA0tJOwYvopWt3patErpPy7JHaVxui4n59+OTGyZEUc
Ox4PmGsolKoPrWXGFOhE0XRB0iIVdmSwD1o3wIWKfADImInTgULBSlLbDcZ8Dy4lOnbdDND/FR8x
syIhm/SitvqgoWL8xabi7YjR8Dgm4ri1q0v5b9P4Gg+xzqo1+LlAtAhj7e9xCie0ALDzbpzc2O6F
sbfy/fcEV70ucylpv2J6iTXeAmK6SuwcIckUnlikswO1g+xjEUnBzzVfi+PQZmcCDue2+9gmW/g1
XvF8yYdfMpzzKAk/RxZ1NDNs/nLt+lXzMcJXf7KF/sDGFeE8y84SL+Y5TuNz5S0KSrrLRbvJuK/b
VuwFTPla58be/JwRoaC8YHwPvVuXn3MaTba/Pn6UDadOkJiK14mTfNuwBs5spXIxOv/JWAMt0CWA
11Q52yLGQ0/B1PZJ1LINTRO2/8LOs0K2srfURIF+tft6/7EUnxVrHeT5zgIypv5SX5mWiqhoSWAw
Zdlr8rP3MljMCsTkRkqKtW2ypck0DfBWHUMLubzygp/6X71RB5Dt2wvagvF9O5bgyrVmzlZQTTUJ
KzuBPwgz4/9MDbDLze7lWCOrptUR1ShECObonlLvpTi7CI9+pncmJmUXXRi+eTOFBSZDdHT9MM6F
J/kEopxnjqFHRMkWVO8FD3tB9VfIsssBs+nL5k3v4/yDMMdy5m8zVhBk1NGPbgPv/OOvLIDzvbdD
cDEVW9wqrpT3RzUz9Kz/7YHvd6bCESdAobtbEBRTySFFXSfvJSPIS4EhF/EYC9m+ve0EBtRvjUPz
l3wkrbr4Q2ZNqRdMHh7XkAh/NEr2FGWwGlCLBrftIE3eAHppo3WXca+u0O/Q1wHjAmhBct5hCZ4N
IU+QOusUbPxl2TYA298krBCsvr7YxFDD9RvYj+q6HYjtEHRsw+QNXh95kAQWC5KqlJ+T7vlvhJlG
JcS2HXruL/QyeHKMb9wn7BjM+TC2fdv8poprjMf5OjhXcvLQz5uLgGVtnX7xBD3cZ5yUuXkAN1gx
2JL70H03qaCNf23jWTn+j4ktBkuFTgmpm5zVrYyvObBOjVSeYZYqJAwd6CiA2zO4PKpj7JP30o+p
k2smshzhdiKQ8mIw5zZubKuV52ed83xANyKfIilOhXm5/4hZwwTHI5m+L/HK2bP3oTGcBG34Dd9z
55qoI03J/agcMQjpLW0hvnWLncW1R138ueZ6af3p1xj3UpIDqml6614FcgqBSodkZn6eaLczMgMC
mV25YbuMK6O60kKPswXk9CtfKDr8VOG5xHN3CkUkowP+ltp5FFSUP9ftpNqNhTj950gc0UR5WrR/
jTWwxq9/OgSX3fQh36K8tUG6aRJPZDkYoOaUrChsaWfdkCyn5sGCTHpsg/bQSq6wRIEraup9/Gwi
tlFcO+5vcuLW9SgTBuwCmWWFUer+Byrw77xo8npw72xG5NuAYhkKIYmxpE+upsrVBCvGa34WI6KE
ZXg2bBl6RUXVgBKOnGViS3EF0ASusMLXMNJQtvMlz7fKL2zzC1HBawH3CBOVsVN5l6NdN+X9iTek
2u8YRaCH9TgFZkobksZgUOcAsRmhL12IbHcYS3rG6nozqOuX298Rv0wnWiFKOZ1F6x+iqPwANxPa
DQssjbiS9kSDGTS0dz4Kx6/v7wXsX5Wmo6Z69uj3w6kymLVQvPUUlgDpDjHfPNWZt9YhGs7DVwBk
/EJMtXUMcnubQ/xkYEQFb6o4YxhMQi7Qtau8T+O+MMAcwfskvgYitOxqk81jG0H1yS0UAZ64NZOa
5LkQpC6eJBv8p7ioCUgy+0iPh9p+xQ0XOGATEoG0iB+i570g4VX7qWi0r5SO4m3ca+9J4gviKmGN
gW/sLb7XLkHnHEkuA6I5I9g32E1NjUdnkVMmnGBiK/EkWuC0VgltL7hdTPLm5kjOo5QKEFqMY/fF
N0HM9mMthWzu1aG2XTnCwPKQrDINqbR4Pjrw1h9DdQkH0g+6ZAQuBqiwssNPO9S2oWK0vKzHQr0z
vJf2khLMynGrAk0gSy5edmEsbLUdrJjBIX5BQGHGd8S/Ii0HDfMWD180pdCRdXTRDGEe4vmVZiSC
QgFNt5+l5ActiaJHkvMS781mLi5AaRSxVjB//T9A58GDHliM7uNHycaVgqrZH0mPR85cNbVECERi
qa3fHq63IoD/14A17FywM1cnox6oZpDbaMbNrRguCvicZFo7Li/zPTpd3CACAmOqkfujJq9+7Lar
nw/eHHuFiJhRmuxts0uFTpkgOfNBdkd08yP4TeZiF8T1qLLbuLH11pYVRD+mRslMgl9qbI23Q/Qc
s2ZNQuo06YSFyzWOTvKEILWsUvZ1MUfqJCw+Mujl0Fg5Qx0y4+DbjLOUx20770PaJDO29jT2wwGC
CV5mQ0iMGvcD40pO1K0RKAGZp/pvzcbq9kddyG/XnGj2ztb7IK8V9rFvB/9slAty7/IPcm4fjr3O
ao6Wvc04TZeyfESLSE8uSQMt9p/fdMuc4eo2MKpcGWuveH0GuQNaXUFKl5P+dHsOjlOHQi2bZoQZ
z0R0C5CAn5QN53x45w8WmzDHboEOA1aS/WpFPmV4dhxe3pGfpDHtm69LX+GzwQ4dmEvTG1kBsyCE
brNkSn4oQsP4ZJptoh5LCJDMQqcKJ8sodTLipHUBB2hmUs2BnpZVpJj2kPAca+CE+sK/l9GLXEYl
cHX0ik5yu5uuypczzQFIH9DfrXMYzRWHhlhHAADeZuAqXx6jQJ0+ABGI61FaEF+lRf1yzvRVVWRZ
PbcfdTXLDGcGara0SLkAKOBKBqC6r9GNzhT4F+cgfXkoPvy7Sh7nUnRsAaMKebetlETNgC5Eo0bG
z7Ehx3B2dl6QENMghY/ONK4Tj77LJgPi2yyMjuuhjTF/xS37FKVkaavywHN/mL+iwdYdD/VAH6uw
QCb33iYXH3lXW6TE0JKuz999TqSH92FroDv9TknqQBMXE0LBXlISJ8Uj+GYks4GPP4XllYk04qcR
6oIa/ALugPW++VO/Uxcs/IpVh8eblGUUx6WouKWF+522ij36MCKRZR0EZQurnjItYUWOMw6PuF0k
IYWA7A2LObzczFplZ2UzhR8JkFR2Ss5BoBGAeJ9r6H3iTEILNQ2lmE1KZqVkl/ThugGdS2M1Anue
UwDbGNlWz8nzF9th4jbBGc4k+e3y7VpF7+DdzLiSkcSbLqUqL3Wua6w6njX+CwTZWGgiAaGSVd/0
ay2AP3mChfjTdq2bxAzwcGdBe8i/ROMCyi291oj6Y0Oq0Err2AWT1swPh7Wd1mYY62+9N5vOeVWr
vmDq0ebeptIMkx7QJmPO+vSQoaf/J0U12/9CLPAdi/SVQsozR+EF03syXpaiOn21ccaQN9u5yA58
ffGQG2NvFLRoWaBnrJtaSYy/k6bNHFZWT1DyIhUOi7kRODGq1XayZd0LSUqAWTHsqsn5Ts7g7HJv
4I+pF5jqF8EQmcTPINu/gZ+CjAb88IEiIadY5j7SLa7NxiCh+20UozJ1aVbFNtGfxfRevBUlru6O
Zy4gE9ikaxf3egq+07ZIH5xPOudoHZd3e6wW42weRGZYJaYk2WyjsmPEgQ4Fm+Ji2ZmfMoqM3l43
XquPy7aD9xKEGeNsmhLXXcE/SSm7FFbtlIrs8hJ4dfmUW4xpRcE+0nSM0Hbybby2wQ0m+2wSMqoW
9/+B2EqCPaKTxywKtjIyQLSr46sv/NRr7WcgnF21gj9NZTTo9X31ABmClTTfS2pousz/4HJtDQCN
9S9CD7G/4s5FrW/42k7ub8HaA716PNDoAuuzfaDSaL5o4zE4eCOL4zlyP3p+8XC+JTbp7ObkOz0c
1Vl+cCBBtfmcwSAcpN4CQEYhik7U9pGJ+D/4Ie01/CkN6WQ+FgZuo4t9tWNXcJFiM1XfTrEMmJbc
2Mlfxm1g8Lwb8PVdIXZdH21NFbWjg8TagyjaDQokwHSA/JcieQzhxzEpU+CrCBq4c2TjYNhavCGj
u447TQG6aRzz/8ksVuNTDZylv0u07xhQxTwR9F+xkMKL1qBvCspyWKIfZwKKCVaMS+qH5YL2YTH2
v5Vw65avMc8HtFqYi0hWiDWwlxmCiMJtUpLlMsIWLUy89nXhcZVhV7OKQ+XNCYvF3q9oQxSQbFP+
WDnHRYxMMba1Rdpb9UYC2Pnb7+1L1PrvwgCxLEzfqVbyKxqCNzZDrdz9+MweTfFCeg6vi1PRiiF0
Uu0ms92Dp7Xxo2w0LhaJniP4KUxuT3DadbBNy7ULSDUR+TS/kda0r5aDUhB4zrGq1yOzMIDr/zKx
yQpXbehm3ftG9RSOX3yAPQE68Z1JA7oq+RwAakAhBanyBVEHISDcSBw5FBaa76eoGcyAYoFlbKcm
YdYwEiGXmzo+X1yDlJDDMlR8f9hEUg3YVtJ5hkuvyarw6WWEfdi4bJLuzfVWG02oF4j/KvI1jXo4
f7PbIg6p0xJf7yFi9ziBFuixEQNUbTEcCyi2/8B7AYc7FdJW+/Qv13yO7I/cw+XY5Sp30KsWderZ
bNFWbt051SATWRFwWfPpEadpgr5Brkek6d72RyrMU7nObrjQJ8tcMmCCBEkKRzOuuJ+AGa81QAGX
y2JYgtWOJ49J8FsbQj4izKdD1FEAP/BkDBnkrV4ZDbXBbmYsppHxBtoaJ7pSzNorbxo0lTO6BII8
mCZ+pmXTibcp2NHnPhGHtH7ozD4AjEmM1zebKRFUyreWj09lZSFbk/i3LcEILTevV1N2sUGtaRB4
BnJ4ZsneTolvW/Ew85htlG4MG1+JNUtKrP8W42qgA+lfuGSN0OlHLB+f8NLZIXUDAEUYe29pvcDW
ZBxlteVLKBq4ZGNA5Jej6OCps3L4JEHTgvM3TvnZCAr6C96SWVQmcbRVZAy3TltDJTHRZnp8pqqu
RLtHIra5i9YpT2iaUgrrgchlv6s7Yp/nIhqm+FePgWipx1zB8OgA7yLa71p+IFnKqojrH6csPz1X
1yKGHEm+MQXDWqbEyNb1NlBxFmTSBrd+XdpEikSdun/orqc0X8SbzM5x/1woSWaL/oNrmgI9/UQg
cDOAwZOU6z6HILGwFDjPyRomKJujN+DbfJgnBPob42VZ0ZqU6Hk4SROJ80niQ7Jn5L5UpGsTbo7j
RmHgUAQOY98xFP8BHuRpYLSLww3rdwl/wScEjHsFtU0tUnCiI1Jdg9oNRNzcIXxxX4RMufOzBMHw
5uO0jHbmOg8LPHAAPMoeM0oecDgvqkRXBR7w4nlvEAWJCXT7XkDF0Bt7bXExUiJcHnO785fQ5Idc
4SdHTCnZ/5KizoCdnWTfaZ+f4cmMR/yK1Rye567ABHoJ9mhutoYM6sFCZRjMSpDYUm1AiShYSssd
Xms/uf0SFBnPqj/IlHTK1Mx/TY60FomVcO0VDxZTE1J1hRhox5h4ZQvwLHhVEs+ypizslHH2yFuz
nTChZuvY66ZCT+/3R7yzWRmwkXB/HuEhG57ZOOBDxQPhy2AHvwSz2Msm+Uh17gXIJOos1SgnQJLo
XQT5Lc8AiYyXRnLJBMC1ktIx4vqVEQU+h9vjYyCrtdqKfo3HmmFue1BRZ7IvmiN+9bjqN8/s1NS1
L4EJkK/8BatXGTgdH61NLjnCY7t0KHNQmDgP6UnR8AzNFZ/Zk3keF2A/7JCRySVnNX4AMjvozOMO
qI6sf1UhFpM9lIB0iczDhFJr2u2xkRpAKb+fDa+V5bMyGYhXy4LWtLF5K1mNnyTS/Eej6i81ACzg
Qbqt7/L9qowi1LZhr/SfXs3dFFHEqfy2m/2YoiM1M6tgGph3NITtZiyftCP7e3PQlVUp5sMlqaUY
dZj7V8WTD98kW9UfaTQ9xbFc29Nv2i+WjkdxjwUr2tG9QlIuYoT7FpEsUOMsjCv/IpLJWkygaFGx
z9rv4l3lqm+Alccy9bNbkyyPwwPFut2Dpa/3mq+rAyOvVCPFIiE+iIgy5qj9JJjpOemp7DC53xX5
3/6QFM7gJewXVYZLxdDtkg28lVQ6TpuUNCnrdmhU7+yh5HMyIu3ehG9ipYbTJFIPoFWAFbBsBtYB
cpBhNAxw1qNEh6nhz/uqWQ4ybhTsiLbXjlIfv8Rb0zfzg5rQ1NLMa+w05P/ms5Stzkq+QhfsQ/ZL
PQkX/cGaRZ6AhpCv1+lpihq1FRjHLlbondvxNLA+jackADwpeyK2AZ8SgRrzv4x2Oi6fxEXsuUq+
KVpyADZQLdjopiAHspQu2poi4iD3LC2KFwBEZBN8/rflRINmxS31MxZ1YP8WTEH9DfE1A7PchKRF
z5Gp5Dwv1CQrdmG5qOPJRyTEvbUoWKnniNtRXifjd40P7mAwjwLQoInyfuEpbZoxf4LnLmqxAMxY
ddFTATH0Olesxf8W5j6teaESVMhWFvBiv2t1z1SMUmHbCBrCcWvrZ5nQpqPKuW6mP1fwxjPM7rs0
8re8Wb+Q22XoqKaGN2c4tgGT+CgpQsUuWHUwY4+KVRfX/dPsPaJfZFAU1CWCAcCdwOKILageGiHe
3eMGT0FnB32NMnEex4itu29NuAGNKRxEcdhWXSUxzINW1JqdkoKkBQAMll2OqZ2kTRCchztRd9P2
basTNlorJKKMrBm0WaBerFjzB2gyendC78iWOBjcv6iiw15GIjVPwFhWkIuqo0DtZZitWwS/fP/8
372YA4bo7DPL2/hS0amIwvzOyV1w6Omzj7NYhuAxVQAORpeNhK08a7/eCrPHpM1qqQdZ/ZaVZhEn
kkzcxaj27xVvKpnsXhrA7DW2t0PcjtkVFll4gmz496LG50yoVnqXIGdGn7523iqRPUqWsncRTODx
B39rHF6buZGo4FHDNo4N5M5fSGtOndG+5KM0Uzfft7VDeMf43It4O1Z8rhGBhUbxAnT0jy/0oSVj
afpoPokFTS5Z7wuwoX/dhzG6xMEggU+C6Rd3rG18HdfvSPPemOIxWWhMPPGovp003p6RFbw6abO2
GhC74GJc1tWrM2i1mGLRic8mR2yVIH1Uvl5/YJM2rRj3QjSpOkAz0UzHHj8lqpikJIKvEjMvlD6b
khIznc5Uwv5lkM9OrP7AUmcMaqKCAFHQmLD+nPVA8gp86Em2PGEUz2JWffXAjs8/uvTw0R9mmNn7
OWOTuQEXae7GR+ED71od+Ko+8b+JrgVuL1p+NwiXDNnu3JTlc3PzDmAQ7naE1lc0YQu5Cibcq1u3
eTmpDIcVbNvp69Nu9cK9ahJZHX+5KKwOPgaAXb7oVMHJqX+SrteYkgIhgD2vH2zAiUKTDIYSxwSW
ine3tsW3XmLTtHCophaAmNU+6AVd6muBJTtKJuix/T1IX4nrnnuWzW3Zx5+0NI+1X6Zbvc3EqAT1
CN/Nm15ZVjAdbFOrItka1sC8yMhShuLWZixOw0fCExIkOEFeEJsTJPiXs6FlupdSdBWEPAn0XFlC
U3WyqVlFV39ooBzdf5lY70cQfkFkILJvYukHn5VaEvcC5hSuz8wX6pg/OcX2zjFTiO6SfYf7/Jj5
f9Hf45oqsR0he0bqnoi+PjBtkvORCLugooNS1hMZDvVS3JI6L6nNFmS3rHlDl5EnFZQbCVyZOQAO
uLWvimOs8YkQ2CD9gR+89Xz93f3hcUe1AokjTMeiZbD29edYwuYGamvlngzYEf2XycVO6sAteCPk
eq51MpLFRoZxrBquiRQoa0k1/5AEhAOi++CAN3cEUUkbt2CP62x41TkAna3lPjn1ybdmloNj/gou
ddsrlt49kp9JxbBlbvKLGiTkn6o8eZYv6/PGMx39nr/EEfgACsylUHiee5iyTPaV1IJbv/nhSE4O
vt1L0VgqKNXv1uwhRzw5gpuXnIwIM9DuY0bkPn7e743IiRiIxSdaFaCzCwdOdx40TeOoT8dShRVO
20c6bGiDGJjQf5GJWBBX9Ctp+YPGGmFIj5m7th8k7kd/a86ZNCqgd3ErVBuUdKYkdJeoT5qrIXIJ
zsT4n88YKltufqODA2Adu7yKJh0FWtNQZid2DRjPNyF1QPft05EBUDxcbDkiu439itPHIFu5H27g
net1/2ZDwM1ofP/snHQ5MBlx7qLQDuUtZxGYY08URE2I3Cwh0xf+IY7v43+R2aqqdMCW0K2oWI2n
WhwfGIuRWK2SuGAQ7pYuAHxJRds2ft7bYQd+I48XXN+zHQhhd6Ha7uOxjBU3Oe/9hOF6EYpvE0Ls
AWPt/bbPQbvl4Ub4X24LIU72nlq5Awq2TN1evSWPNE2dzbUg2S4vf+fG0v44rmOL2/X6c3mWnm/G
ypFwncTePpmgHgf6ZIiNd1IdhgHn7KxXg8NFDNzPAesUh9xRr0auH5lLw6BkRbzGG8FbBAJchorG
vEPmYVm2u8PeZO7AW5eERxIDhyIrLdaD4G7X9mFWzqu9zbymgayj80Qtub3lFSNy5Qogm048cckD
bgtO2TVqaXhb/Y9UozKKfLV65V7loI5N3rEfYf37Bz0Es3cjX+ZyivB1aOVx59Yb6AUcIDZLV1Nh
+JHGa6HuSMMSi40WjtUiShntsqrkGv2NO854T8dGV9wudrgN8ve+pG246b+UQzZzy//HNYFYZwQQ
Elm2NJtMu3i2ovf6ikqYQ6aU7ogqNJVbwZIp/IC7Q+MFBYkLBl2n9dqhhwm3kxC9de1MtyKApjRh
QATLDlAfjuE3byEOEqSvDChnDCUXOSK4CMulTuRMu1QFqzRp9dg6DQoshjK2uTnULnQFxTTHJe4q
SD0VZcB7Ht+0rysJNWbL0wcsWVZA35qkUQoKtGzGs179HgJs4CI1apWcQR+cpkdRz6iHtTA3PXL1
AIrzi5mb4Yv63AL/jshLG/c/SeUHVWTUOASr+PYAlvBqVK8poSDqZBqf8xJhZRJ4/ZyuuNQzchje
+/F1B0xa9QaZpIuaZa1thOOhHxCjBTZFjClNERouTPqKaAgm7aDAP5lWs4TZ+u+sCrlrZHv4NLj4
Ae7M9NonfGhBdAWaBxeNCsPhn9QGw2xbSDc2lkDqA82TnFCHKxML75EcvZbZO+JlvajT3jD1LZDQ
7UKTGO7ijl7A/HIahuwpsMqtD0S5+SaW7mNtDSN8j65cuGSg44oyYAhm4a7fB+5YAcCStBKmY2Nw
X7C76wjNUYLU5db8ICy+y1xQIlKMmYGuFjqCQ9oD53r5Wyh18DkIU4HXooh4nvTYzQeSBYfPLupL
tIGqceBVnLVXvY7zFgjCCSivCdtK4b5ezaurhiLwOCcdB1MDPslZzCvkcO00gvYPFrjpBGlc3weD
Y72ZRzHkzvqGJHJ5xRso9VmJuc2Ymasvv0VGo2k/Pzn+Q7elrOEPoohdNUJ140snX8mQyLQQXBYH
cVDvajyJflRH+XxJEgfG00FDcEtgqb6wWmDIGtYedez8aqV72WrXkQEcG8kZnF+fJPX1AMNslatV
uW+MHv0NNUPbl867d7ySYqWPTzTaIJDZDOE2ep3i6y2jN9qNK1PqYxNtMuibD1/GmUJSreKYlG9G
qXe+RA09mkLvgUVEwhg1KyVsLUDf+IR0c/DI0rrf0ce5B3RsoGSIMBOwj2xTVSV3pbuZhxhzi2GE
+WA3HnFAt4KwXap5jgNGET5G6KTimfT9O5IBdlfmmJPQijJ485JENmDHRn/YhXvYRh55dXliQVuf
uht2CI+NdAcDJrYIx2Z3gUNYmc/2CH+4z+NdmLhf0t3opmbS0MuDSjNo3eEgVbJa4+UCzr4Mx1my
az8H2GTvDP/EL8NOJvnFwqs/EbU2CyJdmo76aGZVc0lRljG8eQAy3GFGAWaRzN+BORhpvegFgHDs
RQSZ6jWMefUyn/MoNI17e+DGne+58jQvolgJY1t/uLwgbp/dYrWajFXvx5KR9WrRioA8BfxO5PWE
Np9FtZf2SQX3IyEVvU3hp5VqhQFWo9tKJRp6EVNFGFDyCw616XXu2MOTjb5YC/zz+Q7+X+q6JhWY
pcN/0c7IroUELMGJI01CYXcSzcIp2up2GhJ7bb2aEYoOI4knvx7YY7vqzlVx1NYf4evOvHme01Qd
fAEmDpO7n9fnhb74LZ/r+W+a1lh57yUurYcs8+hCTU7s2TkcadDu+mU1zwt0yRtowKyKox9jpLQy
uS/2+4fWFh6yNJwl8KMmBBOnG6/nZvlOVzrDbp7UJJjrNTOAbjEZoZg8SJ1yNj+bmPpbpZXpSVnF
SaUs8CB3R+g2MDkBQkacaRXkHV8yXIPJOkpk0YU03eS1YOGNgOSx2C2s1vDbPhU7kDkkE0nSYDzQ
3rtAwnJF9DMf8QuqwSzjobMAMdklKIWJsMhvMVj2dXzo/hj/fGQB1lmIxqHPCm+GKz+MseZpDv/5
QoirbIbdMUq5UJFqs0Xfufg5Sk+2u/azmalbQ+FMOvbHDdGMbnHqSbB8tvdhU9vkbyNEFy91rG6/
P2NTajr7HYXtWDqOi3u31xBrQRDEQosW9pjQ9evOApWOL+L46Us2UqoPbNghRnqHpzC5AHou+PmR
PszCmdqinrbOdZIzMkcDDqkwEsGhCUK7sfl3/uUI7ZAZ6+MTi/csRZDtK4HjpwQ8rnDMmcQyLUjc
HANMMblVd7fI7qLHJSPQnSkAoK9RfdXTjIGTV6WLC8RgxxpcT4YlXII43FFd6Xy7av9d1W/9kSni
X7RBFrtU0pl8h9VaLVKTRMewg0YX1/R1JuS6H0XBrQcDbKy7BtbhvPWnnt0vUrk364jHo35F5bfY
cTxEkTiuLTgdsqxd6JzkYc5UpmuaBBxv4SfAc94GsG9GWGKoBDxLB0Xr01gxU8k3HmLhOtFU4my3
LLoEbJ0qKZ3R1TbKDc7iTiH1Lza+8dZZZ40tiKoGpTX3XWULz/gJ3k6Cdbj8oY0cmhsAD0HygrF4
Yz9u5zdWIENeBKulDenj2JdfgtzzEJNdGrvROqnFOENUYVwudCWd37sDl9z776voG+ikjWh3sqcm
UFtvJUFKBFD32W1fDXCZP3JvMA+sxA3dmx4iY7WibiHtwsn6a52NtJnztkId2v1zMPD5bMHFN8Kf
f78/vGAarWrdOGuewwmWUTuTk8pBILXifMESzYwL43GAemGU//CpTlpT0aDG1QZhpYIFHFh7Mti1
hRcD1ZGLi0F5EKvFGNNuS9UKPs3YVXND038EisSG7ddfgQrZ31BCkdHLynT3vdUNgkZxkoI+8kQg
hzuN0xRVTG6uT2YrGUJEMJNO131qUduJXd1Cg8X5QL5Rv1XZHFu8/oK9Hu7KRLmWeVdIX0bo8BBV
IJddQE3EEBnSwDlZTMSoFMBIALxKRQCgSxW0+z3ND2zY42eaQpHOQgTnajqt93Mue4EKJ3b/DtEw
L5MuEkjbY0clqYz7Jtr8qqJgbVI4NaO2X4FdGmXmjLcE1H0vNq5FkrjkYrfRyXP0CyBK0HYheihE
pquy9g7c/knfi07eR9VTGtcW6tAr4y2ZFGEeb+UZVHmlB2AreGLtUTl6nFgCJSZ4+gs+PX+qlBEw
HLv/mjXaH0qFcm+3FC/fcLerdIDzglFOZNkMQsNlBDcrB0ekWupc48lssBuNMrKgvps18Ey9Kc13
v5sNXQdIvOriEWe2xOwr/D02UAO08wRE8Y74qMOuZXFlVy6+j/uQKTK5ApRVaaMusPmnZ0nplhXo
8MnStpu5rZfqkKen4eG+Ee7Oe6Ey5rSgJ1hQEGqalFUseMFidkDQz03zO7tNS88/Nbp34EZFlMMq
pJg7Ns8wiNzOVGfQJ8nQoiaMz4P0RxGT0fPpIaCS0BFKactG3b9mgOMbAA26GCUGuW+ZwV2VcMF2
5MPQGPsLpx0nX09GFa0Zc6cakK76OGva3+kUhhntvogtKv8yyl155cb8Sr70b0xB9e6culbBaDYG
xhmgl87L/fM/lJSm4xzpFuQ0F5z6P2FecjWSsebV2ZVDuLXbxNhx0g2A2xECn2iNL63HBYGb+yr9
W/AOFTCv8aN91ZhG5gnFFtTmEaISI6T9XCaiEZOXtqB8HNprlTILW4oO5bwqfNVZEnquvMEzBbR7
GK5/62BBvcm0jPuHThLzHPog6Yi+fQR6mMlnzG6zVBXqZiktyo2Y5jzBE9Ed+6isuYxmoPjIfi9J
ri2DPfVm6UDWzWiIREml7Ihe91qATiyA2jgNjgCkC3qQPjItIHty5Cma3mobGE3ZafvpRzU7pQkK
FWopyUpZl5hhzNoJ+0jinEaASLOFurVH1NoV1sdH7E1q0UP/mibfUbGh2TDDrpW5cJsWOXb5fXEs
AFJZXFGbP4vPHsm7s6q3lMbkBXWL8blADBP31nVMLtLB/jEHG2+n9tO4AUg0E+31QVxaVNlTmiE5
SiqxJBHUuqX1IQhalE/nMNYI7yn7uKn3XTifQyNer6oXUTzBJcZD2n0M/y/UVUvcyD8Rd5RPBeOn
DVIbTMooMf0FzuHLy/V7V0oxkY9N59588IYskxVoaWo+39HzrlOOtz0hkCdIDKuet5TyEZIu8SCi
B9OrdI1YOVJ5H3wWp3yviNXsxf3giXcVqpQbzK9pdDHWF7Ua1A8MFWxGNh3Elp77LmX9LBcM78Tn
AsWMStMnU3dnQ6vcPlSleGyMsxnsxekK84Yq9+FlfBzzTs8achEwdMTvAmJG+/82deMHrz8s2mni
TSoqmNOMCNseMqDrXG88zIhJfIglZzFwVZIMAdqBJjVylJlA/NBKdIdN0R+9u+s9VkB6BWZIHVuW
bJMtdt/cAwa6k/b7der2XIjodFXvb41yaRdHrMv9tQPdi9K0cYeb1z/I3+eYyp9m9zIbFwfjO1RL
818RfN4Y5PqlJFN2JlGdOnCLOLvgu9Ylyy52zkfE9dEJfky+0sPOU771X8i80W5672OqIf5immZ7
2vxFP3P60JbhKCX0DN5jflwomFOGs3cGHgts/oxBHm9oT2ye+j7bngRWU82uRX6qtYDysGOQH04d
Y98dD4+JesM+OO1YutprI3sf9ViSILcOk3z31jzrrJY72edmBLh8w8XCZhbrhjFmpqsSrTJuun0u
YEW4V0eEThDvFZcZWTcd4qZnApmyxJxHlPkDwhlim7w3gRdF3bIMLSGgzzAaJN5LfqHjPF6C8N/7
eD/QgDmyqUhTNxV3mm7zCH8N0sOKplgLWnOwMgdCwlNqH2tHm9IWvnCrJh3t61ox0Cg78hLO7FzJ
6NkbkRSJ42xQckXnB4gQynEILA1X5w4lUePjOgm19TLT7aYofEb/DIMRVMilW9REyrMJEA83gpqW
OujYrUVsuIXColul3yrVCUgpvffhZp38u0bk3FP9n6sBTIPYugoMV2/y0qP1yBYWoywv62tvlCfl
A0MV/W7A68Y1hZoXfUJGlQHiF8A1aYh/VZfTBx1NdufZLfM6FQnSeiACdWNov2hg8a4YTwUr04CR
KWIcVykmKmC2sG8L0xrh9+8angZ6HqGVn9emZwa8DXavLFbOHhFfu/30HvRDToQSzKy34naU1CL7
XOxKM42Mnp+X9BUSFjjbXJ8D/ghXBFt63xyTs6k7jparO4awVqBZF68jjtrd0dj551M3xlqIC5aL
4td2M6A69aDwH2KxDRl3yR1TNpIG3GVad2dBo9aoH2s1CCS4Oc7mMWRPS/5zakPTu/aNtpJOsV0h
9dfx+aCEdCj78RFZXkdNUEnLVcynHQ5ALIsXPpej6sssx3kz07c/iqCKS7Pqrab6lrUW9nyqUrFx
zSzmtlDDXud4RoSqfWZ23XIqWxV8wya33yRxwd5Wh5+H7Oh5+sjGA1zt+wJAyCdy+lWg8nnuAIpF
j0Jf0y5UB4ybT4sx25hUHrpqxar7mC78yVTSmreGbtkFKcMTodVh7vCc6Jd2+bmjOCYR1OuhSIJg
dCS1n+u24ITG7eo/E+xfq3/SdBv+AqDM4v8Hjwo1NyOUZk7p2tzrtCvkFXcF3w9VDW5k4GyewRq7
So1ug0N8e8MTNzRtw1JbLyjogcAKMwiyRKf8qxmkbHxJFQ4x4ptYRw7eBcKNfHvqYzbMgP+ge8+0
dhmaagdljzla074pkMQmHQW4twiM2rH3gk0qCWaoBp9Uql9+VSdKsFuDALYSb/eVjBU7KKy8Hl1x
N2pnK2L5Ji1+hXYjCaOLz6PBzqM2HF6ZtNomR0jsh69DzL+w2oMyNs89FIeBXqTc7rG+rIbq7TCK
94e1LeEhxjEzk0srFuqNXbmxhhlMBbkJqm2ZAMVlzdRN16deEWI1JQk+2amPeaXusd7hTKKG5m2W
kDB0DLKKtSgCagZDKnBWNysl/WI+d0aO0vWzGC3fnkjQXk78NjtysLR/9wLpFmsj7CFUmzAD6mKN
FTefSNnCe6UF9jMq1+ZIqMw6WdNlwRwnBqO5FHogYoSmceHVjAk8q1+xhI9qGVAum5fv0cbWimDl
IvM18gNJRsGHtyjINefX4N666suUmL2a+0IQi8eDR9Rbj/Ich2MXkXV6H5qvYRqS8buMr4tpYqO+
rxqf8zaVUvlVtQQxmQnR8VDBGtmHp1lkZAVNzsZOhwrokqm9WnshYIW1ku6I6p43AYXzEIai+CE6
pMJ3uUXYfpsAu7V42n7OV7hOw/9KOFocpHX/NZAL79HcLVd4dHwMdOiAu7WlLuDg077O9WySSy+e
NI9qVAx4MrAaToK8eYgMDqmRntHbZAmiNKQ8XyxX3R7tubptfG/kWCQ4HVFlv+oDlkTyFkSNKQOB
xlL4XOlAMlR0NUDipmlrsvxbkvL0d+EPiMHEHA7YrexR/gktONYwlqanZ6uTMq1YTywHzJwHu8sc
Ivxglh4uWg9I1qlaDLZu2JEAuYaR4MqR2QD8PmXI5VLAw3RXpD3/WzocSwBIlapJW9UIylwoUAle
XRY17nMc6Y6NVEgUgyjIStEz+MOuwKFoU/Xv0e/AOev8WoHjYBfcoT/icteNTwnFs7BUw9En1dWv
EqEKHcylpRhfS1WLW0VY5W780CHsLb5Le+yxercBrY8itSy3IK9gdWQvEzXM3QASy3rVeqe5PuaD
C4ZLxAszCHag9Nw5OqvpJRFWUYXhd4c7kRNwSL4DtPk44HDDf2JYhZmpirOKgYaqLwRaEFxG1l3y
odiu3I7kNbWyfscr3y5dzINNqJ6s36IbNa2LxPP2j7Nvdzcmfj1kT+24LprLHJAAAWxtLjR95HNr
u0G63BvTeItWt/aBiQTpqN/E4bI8kviqWaWpen8rfEDqdnv9l2V3r3dp5aXVTHbG/sOqc8TxAnR2
JEShcIJbk/ClopePSNNUwnxS8rex7iY0KLJXj6C4ilVtb7Pz50nRQk+vmCIxxIxu5SR8HJ8l1OW1
hGfJsW4Pyw1Mzgqj5Mi8fWqfClTu0iXwpXzJ0ecBCI/NnvA7b1vVV/8Q/mKqpvFocZuF1aiOscPH
6A7XXYiE8KwdU7Wscg5ZJ50+6c7QCmQD10FIWShin90J0yijhe3D3vuSAtZ5t4haoQY1Vlgrp2hP
/A1Dcf4sNbr9TKrq5WRtms/E4QTM007mMF0Nvpch3wuDTZtvpu2Evp3SbfXQ1ZhsrdLXfk0zDmsf
GIJ5UmA1XxKqB39mqfQ+MEMfVw4EoOt/Ef/q8cCikZKNLCS3eveaJY0MxpWEG7Vjes+XFh2lWSWP
yW8rUje97MSqazmi9pNMVuB1AuWeNnetN/lyFqiQ85Kfv4SkPmON0Cf/3PUmIACKYG2vMTKM/qaV
VRU9elJR/36yWgzRrT2PIjfBWJBGzvCwXtc4a+UfUhErVSwASdbLhEp5V6W+Ng1H0Y/1H9Q5JOph
Dbe76d+FFYHjtvkbZWjh8kIiHxbR8mpFhd7G/KVjOjHk88zl64jbN+YhVSKnDCdrsavCFATwCovt
A2Wnxr8qyjLDDT3QYOAdjJop5SMtUAngftl85g46U3yDppPx7/zOyrKT+ZO9AMAlZIf16NhWNO+q
pSF3IPiMQRJ/DxtPVxhmKNqCrZdBkDO28eRZ6Sdz2Ia4/HPFjGB3VWhS32IBtYmCvrs8j3oaCqas
OLSCi9N6KZXc+NnNKlfPUiNEb1IRTnqOhiSqei5Yzv3Eta9+xe5pva/5eBp1Z4/LxZcU80/FAt0A
1hBHVkqTVaUXBIdn0/OAHG57Q5KQTNo2yOd5I3uCZBrLZ8qT/cmNwvdAqPP4BLvq2hsbmYVqXu3e
5Oc3vRPaoIL8kK+vYiLj1+9g5/ExHMkFp741wmcTS5y8Xzqb7HMFw2D2UrujcFEKsBSQ424pfdBr
0EfYMSj09eS3hGHmhSkW7HaD6trZL4EvGRldW+Sl2bxIEYvhH8ARV0Am8vMle2wY/nCWQDTs3Cl8
+wSnmm1fKRRNMLMuYh4jfUExcqY9JDoJN54Qo9mwVtIUPNXdWFfpSqm6ndbwqg5/9JWZlRWzd946
Jj6u17vd4ORNpDyP/9+xdTHed6qX8WHlsNKE1voMQfDZojEMzjSifyR4THTh5dITHy4vf9eDA8lb
V9ld/tJeRWfQ+XbONwzY79Z7EpgBwCiGDTKAjsw4z+XI8ZkBp6MMlukYTlY4g7l+2wOzjeAuCxaU
x7CbwrUPeGA3LJZ8/mjyTJTUohUKpLFCw2AgaecdNNj/w5T5ncyFacyK6os7/T4YVrqEDRBvbX6i
MrWZEZY55zsY0CPNkaXCUCXVDuTla4F2V28sP/q0xEM3PSrW3K4ntRbmmZ63agMoSzH2r3u4pXXA
uyVkuRLymYEP1WvWHhxg5f8CShyqbVyKd+2KLH9KcEaxqnBqrz6qdjUlHP0xsJqRJczYQEq1S/Lu
H3eFAEbsMWnCcheC90jgr+MLYcFmBrXRlFCHceIFuuUnlzay3/kVAeklI/+AzIUTFDMzP+bJSpzv
46wjYb7BJEgGYJUUJU1CtlUlC1I7maqY1UsIzDfGKR5aGjBQY0aXI3MdH2Y9UNZJ4ThbaLz3tBzB
nuWn/3DiTIpMWJbc+kyXxnKR9LQzycosXuztQIxesno1SY0cS2Iz4OsgH3fxn9AnUA5/OeN//auR
XxbKmqQfdATWEEfuYRQmRQ2Tg3BrRocMIUYv4JD/c47LUevGWqnpUbbhqjmMP7Frt0f9Yzpfh8Hu
uKqqg/bJvbxjnPq1OBjdTHfi8VhgxUewzdKBDlkKBfTEweWggKEWD4eYmNzFbhLK00OJabJFUzPP
6hhpi5ZDr8/PZG0qkv9a08rPX6C4328BFiVo9j4G7VqADG1JA46JA5gUF+rpLQKf5D486So68+IH
KYASyo+wkGNCl+0Abn96D+hlF7/0fTItMuemD9xi67LL46NLjaPzlJ8SS07B0rzVmxzFikYUCUyC
HDujtnnYA2mrXfZMGajsdoU+HDsP0eBPc52KeOAd4LAir1hW/n1s3jb8OF+75GKjrTtCIoJtPXvw
iux9lmqZ5ZLq3TcAc4PFrxRD2MG45HlFxSM0Vuc9xeG8R3kUmZb5nn2d99XYAWv4F09STTgrkP1g
s7WMyIo5GgLfk4PpvA8hl2dFfpsVSiug1dEek84FtRmUdVZFQbTj7x1aMkV3/6TpiPx6PGRjzqc2
qoT0iqPr/z6tRTD+SRXJw9w5IvwVj356cuFnF0As2Mong17MtmMuMjEixGOG7oEpj0r9Lmf2Q8mG
I/fFC8CzScvMm2caGa//YBWKm4RPjd58+UzKfayAs+Gq/kB9rb0VhKF3MTDk0a+428IcDzHyybdz
v2CH0+pIrnJWbeqOCKQVupVU0n66XZa2Gdmw+gkGW3oDS0m+2pzRFPEPgp6EumeDeyY1Ts6JsAoT
GNELekRxE9OzIt1eP2/2xa3dPm0WorzLAhqMQs7r+jf5T52dgbEpz4jvgJgwmsgN4UuLAqN04Hi3
DeBIXvqR0BF2epz+2GIO4sWQGtj1S9swELbNhE8BP41NG6X0qp7hN1KvT5oTjJd+6cVSTAC5bzCs
6hFeHx64dnmhGl03C5z8ZWExld7dRpQFgjV+a03kakDqMxj++Docx3woaHN7Mk3LMxOQxtvcfSJT
QbD3jK3CuFneVyG6w7vEzIMoy4TnoRsfMr2qz6abZSNDCIStaQ1ceAYmYUpJ1mzg/HqGVih7zjVD
Pu5l/EVmTwNVM67a7L6ezLFIneHcoJHnWWZSAhVikMxlT1bqTgxT1g9LbZ+Wtxw7IQUKSHLeyYUY
GcdgI+w7JD6iAZsi3/S0JYR2VvoRktMIHXwLFO7iLVYcCqrzqfUY89u7Gsvz6ZPMFapH6/f/e2dV
w/KMLx+gNFLBRNTPpzCuo2RAJLHJMGsI5vw9bUwWDmS5DrZTM4j1tf9MON5dcdxS/2itbNZaZ+bY
29P4ooUvXXyPyZKs1Rb8jBTsPEVek1qu1JHfjd84c395OR2VMvlLwBVQJrP+rSkDS8RFemN8qMVS
lMART7bhHyHR08fbp1QcNSu2a8wM7IsD7XY06icngyMNGYKdl162vvGr6pzDBwIX0bwHXs3gIw0g
pP4EHNYr2rtx6iMEPIRKe+tswCWeTTAVdjPvH+cNJJts99SR3csBTeC1VOxvgbIw4+wQBfwO//I7
+0Plbj0OrsJq7099oVWJzo8MlyqZ3Lz5RNxnG0ybQ1s6uYyTOajPosP+G/BbQQ2MPj7zklVHUv7N
gPN/aTTSwXZLlm+3vTb13oIpGAGOEd47RJ9R8B2Zp6os4pBINZLU3ge270dhfnU/YaGMGvVrB8Zx
gz4V1Tp+hAcdgSO/kX36C4MLtlO02CZtM4LP7cNEQ5wbNMMd5LCMQcnbct/dK3NEvw/4JItBrxAs
hZ24tIn+YjAmZBVQCMwkGushotTBnw43p8krwiokfsIm9nrYPIPh5oK8pVjPBSBmKeYj60kzuko4
KVDKnOBjVZ1pEX2Llmuq39i3WM8h17tETMMIqdeOZqjP7l5uCYwI6gxthc4L0WlR3d9idMbFRIdt
CFcaKAUTg1T8Nig7N5IIG1auBWso/NUgbmb+CQPzImlRYGljRThw9UY48ytTQiehBVOmVyJzIBpE
66EM5OzjWu6MtJST0nO0LAi6Gh7VgbrCruxe4D7XnMhO+wBj0CrWJB1PT9h2Q70a35q3Xly6gWSl
weJIzqZ21FZ8KCvbd+kfowQ4yAGNNeBsGl4R8PDke8iEm1e/a44fs+AkEsmTdIw0cAHXFSAwDGCi
YRhuprWhMul32gXQBwej3YKfyYxQvLaUCvExkXFKfzbmrqwaVuU47jYc1bZvv33GXAr0DhC9zEYj
wE3QRLS7MOp0utPSUXCrWrYWdJgdWFqUCylgUagHdBdJ+Bwd/R7G3G00Lkgz48aHu/3IM4on2JS+
yU/W15VCSTskVmC2UGb0TKzh95EWjKoIoGow7qvL6Bf6pcRf4vJQf8tGOaZqOaGDs/tQAAHrBn9J
y3sWAMbaKussT8+YkZv1GYbvWCunFWU8G7IAE/LzAD/jfmxY2zxdmbAc6bWmzvJyGq//387+KA96
xKY0IbtFnBaPhx1BwfV5nQ72cswuzMQ2iTNcv3TuV7lU2JUUcg37sNpChD0L/+PcPzXjmP3/1TAe
ZnHyNyupzfvX9p37NI8vkbnMTxS1YZxGZIEh43LnYe2XzzZ8JYg647zXRgJkRmLqR8VyrEeRCWfQ
d40Xv7RT/GinrX9S67bqoe1AOY42So9hX9PKF4qngeNvrd8kaoNf4rWcuHwV9kEYvjKakIqzMIP5
ocNJ6b2FksmMbEueUNSUDwWZmO0dZhin8cSxhigD+ZjfiCk99H1HpC5xXwXymhBOgGam3rbByzW4
tdrXcP5Tn7YnhlGnSWFelasV0IkpirPQtkhko7szf1l7Pa1hjbxdjr2y//lQRS2immG+WwyGUzsT
ZjSZG8s+BKRG20O1lZ3h18NNOgpE65vP7J/3F2mJDcDCW+ZJSco4qWPkFTKfBrIhIDmgKw3x69/D
a7i5+mGn0K7/kg3sSmJSKYAUFfs+KTUrYRgjK6fyUcfQZr4ANAEFJmydr5fz9W7FZ/akaWoYVTfd
hiem0Td3YVisN7tzLvz2DInbA+dr6Z3Dv+MHzbiQTDW/9qMf6WKV67zix8qqcw4Iecc79JRf0XBB
nPwNX01sHx3atXAtIFOQQebXcvFqvdocAcQYP8x9U3B9CcnDl+M4hlQnFcadh9QaCbBQHcQ0vm4Y
HuC4x5WU9o1nG6caG50cxa2nFVFrm2yYn2IEmiDnsemxr77RZwt5yU8dQaId/MKBxHXkK6ZX0vD6
8uJXV63T1VydQGnYASUGonSBt+jnKBe+QOmUnECl+hdrZIOs/mW903pGtfendExcY3PVokbbYhrq
+0ZI/gfdCPibr8FppdgcCrlCdW0OiNsZ5Q1UAppsjuTSWes6Xz5W4GCLWuq96fayYQeoKVHUk0jE
9ogiu7xxQ/z8k02MSQ3mkIoYJDQ4mirM2cTmS7Lpfp1z1do/1EGb4aBhP4aoR+P4Khu4iDXbbPAu
D2i4WAlDde19uXW2nb81f2+XpStLwsLJ2AjU0l0AHO65TQIBHHQz4vNfvnLHq1PCOj9rD5cv97R3
L0eDHAkN3AnJktKnmD84wHLXxe5fcB0PfREXEFxpzAxrRinzAdn1TOnutCGeMHuh3isgV77PNL9u
xAbLy81xm6NFQoHPkvOdrTDtMiJcz9qIj/Br9NFkH20aSZUcn9jkBsve1+NxMOl8OGHyruXwI1ov
pL5pMcONkKj18OkVKDb1dYxedFRhzntPqD4jj494Qh7/UckV0EHt+iMLqMs5znYg22BKIRBfRSGJ
5E9MLUblL+YtCQUXEzetf9jkXzOZtEQMs84IQCRZU6aqot1CC+eaPl0ERYDnFq56jxGS7g4F3RjQ
VfuKmJTvSB5zY3RuBU8BDBSw7wDDCR37yl7y6LBwn4bHc/0nhvlQlgM9voUEhRcCrmAGj/4JZc+H
ehXWbJGZRJ71HDkLSjIajYzKkc6azuhB9DCcMwrHHoJ8KlRZQTK7LZX3NM02J6WYROeRa1iDCdiW
vg7qUd+E661cHVBLBfPkhDpNeyMWq6HgfsLq7VKTyvCCxLYh4VXUvSGFHB+IXqQxmR74HaB1ZiMx
6J6hRI7mQVzntz/INK9Xxj9qsk9lzhnMiyV91zjGXD7aTOjPwAja1IpSrL3VTPepciUlp+TcUvTG
1eeY7ikc7c7ab0VjtDFw+D0Atg6lC7IRWcL3oc/mDikmosYKVdK3FR1pc8eYLdZOuwgjjJzIyOCd
z1hbl6aIkh6dlOEcyAy5mEF7nHSpA/wcbTYqoYovvRt5udiZRdl1WUwlQx/gsawyNudySuvclTl7
holpTEYA/FrT6K9E5PNhRhXUSR6uE/bQmOhLCQevbZBxKCQ9217CQcXvKuc+GlYtx4SislvdqV9b
soXzX6HnCwRJ2V1BIgzqsuXVVmWVTW6JkmspyVK1FVnoYUC69GDsl/cOrzZLCAsIJy+SEbDXMG/8
rFkYr0Tb7Sza0ogviZVU0TyVUwGIwqFSekso6x3Zd4Awu6LvVU/2LKmWkmUhDgkStc8Y17XIZyy1
eFzNTy/nxbXZMBHsjxBoY8jjw8WELMVvcJcTsYiCH3bL6grLYRZ8TtHFA7aLmmCi0DCxUL/Y8X7F
0wNb9cssJykrrOMe9H5jgtn5mMH76KOCZxc6Z3Dwglapd/L2/XGy02p1zW7O1kA846wVsGWx4YwS
XKjZrXOuEatCnht5z0BYcW2Fm9NdQvqRAO9J5xOEb7Nph6QfLoBE9nrIdh4Cb5fn2G/7HP+dGM2J
8O3bftI9ftWqKsngT0SNR+1XxESkkR2l0GXvPeZ/avZxyDjpi8fWYSmfx3foCfzgl5yKvOMyqMH8
csIhxf4+Ys+PyqX55z0g2RCOlPcmzj24kMwsHq+2MH7yGMTVhA7t+0L5qIcSpAHK1AeVRnaNQKRr
ofwi+qAPnXU0kIqxcrprqGjBk5HiYvCRWbrR/Ui0tWkI8Lm/oRmIWeFcR0/2/sXeG0xf4SaAJqKI
0umhPyjjoBBMbF+PwJ0Db8eMVyHGB1Jgvf8vzxlRfKCtnenGcgb1f0BEffkCekD6KZI6OXBmUuIp
DkOk66ZisZvxMU00KOhokX/b4m/mm5x3mcCuvSknw5WEVK+llW/PPC4I8EvelJHaq3aL3CoQxN9O
3/90Iripe4iyz8WqCJ/7l3gevV30VIihG7fw9AI3UrFJC8YD1uUJEt6Y3jCnwuB0qGx2BnkdKIbg
+YsdBWYo2tt7dqQ023YHdJYwxDTnDQN1WN5SzHQSAT4HXo3yW9K8ijLstzowox7aD15gISgtF2Zt
hNlz9bZ/CawMstBDkOdvq3V5zXFYqBRYhHYVEKEv2bDULoWaibWJ85UHsinsPH7Whi5nusJzbKIP
JaREwjjHt2LaLfhwkD6IScioqAS8PGs3shigQvHot140kw5n7wiZAfSa+d/bOF/k/ui65jylVVxc
OyLvAzE34DQh/xY1ae1+/7otti1WIFepl/msPxTBN8B6RDIxSdn0xXLR2yujmll7Mwv40o6eaHYE
6Nw1RvjRp67cp1jwsE5neObc8aEytNEB2INIjfpfPPkbMqW7rUcHHnpNdHMF2v9kVaokGLuMVM7K
V0Fje5kb6J21c9orVaR0qJa5vExJrHCu6k4847sOHgCcE7l1GIiqxGcjLWToorfhpOoh21iSY9kV
6HEzMSV7lxxZpdNnOud8KoBdqWUWqgr7MeFycWYv0UmxdvrEo0cWF/h+KtSyFgFhV65TDLWcsjoc
hJoopcYwx4MhBmUKVuoqJR7eM9cgH+v2suf/X4bo/4xkKnblorHtWNR7W33NR7eNMbRD73N2OjQk
4MA/CAvhOdonMJwW72Y32ltmVjC34o0TP9dsYy84fL8M+gHnn/U49pPxdq1EwY3zb686NQLS0D7p
HfvVMepAc1Ls7NGQ23CFf/AZuLhl6552uZ+v3YlcETyNlnfrcxqcruSkF7yNoMwIKSo0te44doPK
l5/QvfbR0Zt6FkQyeDSQZ3EibV0k22NzH6b2jLBb7qNrsvgg2CbUmIcP82EvSQrtEqTbAewMPWja
IpkpSTqUsd7N1jVQhQIvcjrvYd8xfznoNxlFsrE/iDAfeFrH5R+HXtUBsf5EVXR7g/O8EXylltWI
5rW+WffOgmnxNbZkXLMKcO5twBtpgXgsTAVtV0j1bwvLhkJOIiVQGhOt7jMnDWkgu4WSktHBjDJT
P0kuhAeKUAKUJTZL6hfWMkt3SFmfBvLw0x3sWfZFV9pF828jrCEWNKAP1H68nLHVoSXLgvipSzjP
HlnzC4UDkzD/T23l6r6GTnARwQe0KoqkV7HvyiGxHriDYF9ruKUJFbdj9mijQ9kmodu3S8g/hB97
fdXk0tudIxGc7TEEdviEARi0pZTqBuThJ5adb+CssZJJeclS4/mqXswfTFp50n13m6mqA8InxMBS
28/tb3PcEgUbub0BCaw9w+H76fNkVvhHV888mNWMpSHO/tNIq9nuHiDLU5Uy86WqdOSF6s+0nj6C
DzvPETLVWePpFUYSVIF7016Du+wZklPLrk4hiFVaz3r/q/wrMhR3oe253EgqBjIW5A/jInQgtYdp
DAA5zIH/7+SNjSeX8HxGAjZyiIu5Q44K82avkh5Nj+O0pswoEiUFwv4qDckMpuP47N9ZHXqPh8bx
K/3rBYRGXF0pXoHLpKOMHmfwcVtl7zqWO5IFWX63cCCO2rGBqeiz+VYVkT9uvcl1O4ngtIl9TwqW
3f69SbMAdnr3dxuSShYpLcvk8FUCO1X3J3UMjtSCuz6SGU/ShYSY3QV4ZrhTe6jgusIp2H/WI43l
nm1NzAv5OLSa0N94dXm95LfEruxLGLW/nzhcD8cSNJcY8uvMSYIx2uzlO3TZ5nda97za3sxc1iNL
+xquymRdLDDFeQ1AiYwmtZZHtSsWyRMCdR4MIGyP5gS9pCoYT6FEpxMOBTxY3YmJybnc1ZWYru2h
bSzU8klQveOUuLDNxUyf6z4oQuStDQUW7on06Fz6aEyRU4VRQHHu2XiyXSezJTQZPFwjb0cnmpTj
kM11Cnz2wOTQ7S/vD1YWydt7YMYww9UUo0cZA0ex9CuKbUUr9SZAS1viVShC6YoaiSN+FZJQf3aY
J4fhMiPt08LXDX82Ta1MKjezBADKZ0I+qNz6F6jTmOAVAODmr5M6s0eHbcSTlzPEpzuuBWDMND36
LQl9d1SYN674Hj8yePm6Du2NbeXQLAlEFeygPCs77wc4ZNCX1VkiPgeCDcHj8wf8d18G9CMdBYdY
6rYwo3Sagis8/tAG4ku7h+tqMJoCdJuWqOH5Y6xEFjxmbb7RBh1xqPScA3wxdkwmjgPa6Xr6Bz+f
qG7hY0wjUX7/6XRC5vOQepcGiMzIVhpvHjBkL0Jd4SUVfiFGNJy+rnkr6IaGd5vH9GyUEo9776Vc
urBsIsrt+8arwEguONxEN3FtU3F7z4Ij7JCy5DKuTixS2xDCmvV7VDBz/RJeXiazQKtrnWw7XpjL
JrQsobnJhsUc0Ovdxo3FBBj4vT/N4bXBgtheb2/qn9qY2uE+qQtf9Pw4e8EVLsKnMyuzHm/k0R09
2vpQ7M+AiZsqOwOlJeAayy4utycpqg1DwH4OSQcjRIOFvPK8zwtWYk5gP96ZEi0lF3V4etz2uuld
H1eN72AWp0ucsPx1kmM/GkL9f3Y+4ZPVcePidZjVebnNiKsgWSfL5RRGGz77LGsLPhB/QfVgeUPR
4KPooKmLRB0bTZx83Wo3WyajK1x6nveb6lJzgSGUFlvFd1cObaAfe9NGkfwJYtFHzA6xwVdfKNyS
gNrmkmlP/+ZiNO3J6SKQAmmygtHQjAYJcWdnDijrkZ3/wmpiZ2wDfikGVnKmW0T3UtNu4CDGhah6
zJXc7QNbUCnOimpI6PjaPDmV2Idev81jl8jyxefdxtioIdKhSHlCiuulB13XnDhYB75krFFCdDaz
9rzZ6CpgjTHVvCNeU9VUBHlEasAOGQ0bK0WutWSdQrcVBsYnUrlROopnfwjsgLF7icjXh2f5ExtJ
Dsb1bvrlfka9PdrMTmtjO8NgQy7KZQQXiF/E4ZUiIN1QZejlQE0vmg54Q0St0FONRATZiG0Ir7J1
Q51IWGFNfWhccJw0hDj65YBbsIhVkoF0WvaHefFJM+zlEl3j+hBCxrtBLrUb0uTb+sy/Wq/3lEy7
L6PJRFTCOIGoNH/FabnzzS+H89S7LO2ZFj0GhJTcrREesaYKITVlOojiYeopK8174AbaC2qFLaCr
OJILYRyWg846oUDlSqnm1wCx+7S8UKOqncjLZK/NgJY2RuwGNUa51pU2cPMT++62MJ7VAp5ATq/y
df4Ukr/lTRWZCip5HBY9VFqEThW9Kdzs37R9LqPz+YTNWPMcP8TOGzRHO6PhAcEdODr4WfG5qX6P
4Zhe5efPh1B8Xz5WfXIRNejuRzx6wBRu31ZwGH5KV4xaNtMYL7lgsweKkWxQI3W4KE9ujYKzeaKY
I89kSGAhdBLWR9AvqkYHMxe96DLaqk/hiM/uS59N82mpscGhcZSVDWf30lFGbv2tgT8xbPhXzbtX
VLFvvs5ghJ0naWgnIvbecie6WndWM9Ra4vvldYNVhoTxDdzCCMwU5HOdvBRCEEHDr7tiBWg90aIE
36X4sUXdEPJMTNP8d//V3ycbYCIqp5ATW/kmti+70rWwdAJ+89oOMXWe+I3zSBLrcEyKEyTkMidU
oRxrR83C1sf9iI8rJbk9lTF7z5ISQ0uCEkfJmdJaoEhLieJDGZrrc/BReR6l4NRyC3PmaEhFKuXR
hjGl2iplGop2HQdmM5ML8tpeYMjXdGX0jf7EA42AbY3NWXXp29XpI3mzz4EqUAiKJGWXj5TH/PkZ
k6hi75yV2YY+sIDUhUsf/w+WQKTbgAHclBm4WEVGjLstUgZG25I+c4p3qFiq1LdDqZOrpAl7faIq
DVXrfUsgZg2NxuX2ByY3B3hZ2GvxkWkAvwiFOTDDBN61Y4k49hEiM8IMpCXaiSqSEWsfiWdQnvh1
LqhUUqJNvuHiecG9twljIY4TmNaA2TPfaQl4wL+54G5VfDeN7BIb/JsVk/kaYt0uSwo+nFxwk0gW
ZIUrDE4e/fpESjatfWJSXgB3z5eoQw/RZ4MauV61f8WkQteDXN+8ku4TEKIyp8hiP8fEFXo/3WoG
0sFIUtAi3I9/DeGU6eieiXQ1AAa8aGfRneE184ZA/xa3tVqn9egQWYJKWyQrEeqPLsOtxm3gIsE5
j8+akLXSbcb14zO0dlraDT4iwVXBCcXSRcmXSlxQwvtiIzxvmL97Q7U+D8HRrVFht1huhvVGZ6C0
JA/xG6740Abx7WD3ukwSh44kfVrBqlOCVX62mrb3aa1PqB+mq8qH7ghXv5oNay4Mzf6p0bhMXRrC
9gYWEPmynahztAfJKBDWG171XYK43Np3nyHNUJlwLmEsvOckU82JFtW2/Uz88y1O6NdH0utbTxqv
Im8WmHF8slDXwUEqBrJWDHjLxhZJ9mT5OaQnrMCXlgt9P+HH6bBs7l9yMv2/ZT3cLvKcMxcaeI+n
DAYhBZH6i4/vcIt5xTL6Ir5s3ik3dshN3xu+LupGJU0VoiFASI0RZ2A+9YN83OYLO0VSfky92Z29
uFz10mYGBfxTfIje1J6x+pEk1T0SRmfbHAiYDkSQZy18kIaovfA9GBX3DttJesEAKhZdVrPbLvf0
A7MA6TwKzBZj5WBp1wp0dUyVdzaX01FrkXNl3E73HBF3JOTWar4fqe4R/RDBU22Xnhmf1/aduro5
jQBXF9UmZqs/VTQ25v5VCeizBhT4oehqklpYiFDho6S02YlclSvO0RtYxv9Y7jveLNs/Pu7CoHfS
PEBB3dgz8EOaU4wOJjIty/ihrYxaeMJ4AdbPTcj/++0Vqrf7NS6pRCS/wkv8YkXOr9h1JKh53unq
uRvL8vC5pz0H5k01W2Pkq5+GbrPv6hoV2KG0ZcSqH7d+hVaNEYSNLcHlFVzck8C/U/EHRrmmPnlh
OauHb0hOqmyTuHCjuX7wB4f0Pr3D8IBcFoCWHe0/QzmJTjoiONQGsN2VS32l4u8wRxuBN7KQfz5Y
Bzn4T9nl75eqK7t9HW3meLUPS7eDs0MdjlK+9TSC2rI896PTb+Dhe6xv4iPqUM7cJKhqrArnYVdy
p8eRcEL3+tnjYyEo/psXy3MKerVx9t8YY8+NaJySQvaZT2koJqvuJKda1weCWc6yZxQTSLRguuHP
qN+n6YzrMOYrWND2vbq83YDMgw1HgXmJDW1ToX+tJED1uGPdK4fpifXKjWGd9ZG1XsukaKa8wlQm
DZjp4i3uH09C3zK6Jt31tL81soUcR+8QVH1hEv0RYk5FdHuqnxwTUGj7CTHC+mrHSQYfdIpWnBty
VEwxckuWoEYK/nMO+mvsSmVmSACmX48p1/AdzDycW+c41EJ+7x/77LFlf9OievhKPMS935k7SMjZ
+tAQeAVf3+MH8YicNXDA3tGcprll1GbU+EwnTzScZqquZTOsPKCBNP2hVl1c05cuCuAc8zq+4Llu
IXGOCxW7gbkv+UXPheBxNmGiovFZN+8+iUSakZ+lRL0FmIAv3zXdrpQdq2PEBP7vfOiNUn9S7npT
gM39+BfYPLoVrRynxP3Vs6sr9emckDRBrJyJwJ88Z3evV0s1E9w0oJdo4RrAOGFDDPwP0LVUY4MM
0ieppJij4wQfelTYuNX1aWJrVmfNPOM5jMMoYFrxQHtOx/zb8wU3YUbfobau3UzPwDlApMV4xiYQ
tZsreByd1B8n4yWYhWLfnVnUiy8lK/lBf93HyguD8dlJ72K6EI1cG/6dWBJdwyTMFaHuzKM0Gexu
HAfCIp6sgMkUBxELysZcBV0pnDONvIti4ewetNRdy3gw/dfNd15D6wyryatNjZcc1ZlJxL9IVYFK
83TLs0HFjjjKU6W2fn9doC16mjCvTM62TApT74oKaunPfO96C2T6aVL27vA+Cx5XXAow8Nu2PZb3
WhSKZ/9yoBwsRe1M0foKG2foCRy7D9rizrdnLsgLt6gbNPWctH/TqUp1udIcBoSvO1FCO0G7FusX
NWPHbCBrV5i1cjlJoHyMNHB16WyNPm0PPF38ZZXI7Q4pnKOL745WkIZoofSvEgUP/rx8npKWigTe
NO6APQV9uNT781WpuLvosYBPcIMnmbYGfrwxa12tEGCeKyT+txag59qkbPhwHB5NmvY6Z2/0nwjW
5RlWOtb0LDhyozRvE7RY83YaM9aYCRaQguVUhAIGoB2tLg99/owp03hBmbQjXxHJQ+D4DW31ZxO/
EBu5A7STNDMQVa/zy8hIMxukRTEcHdO2B42/aQDiqy6VZMDLBio/Z4BAkX6t8Ml2VVME5ntomN9Y
AXuDduwA+BPWBQfF4rjOSte2cW1jmBgE8TYVbTgwd87lRWloFiOTwrTX+OBkEUy+e7GQdpvgDBqB
rllKO5pCUBK55CYM3lyWidgJzoqyCOmndW0F/WxuzM08ViLkfdwxJeGs+nrR9bGmTRJalGLyjgKf
O+gyxWaME5CXasGQtsT43oNS7cy++6k4VGzeGBr82iDaaQVbNqq59/CD4w37Odk+vskvTEm61hm4
Eg8Bx1G4KffSn6wdaWGZ1HOWlJSvuk4huRbCH/UH2fyVQfs5Lqt2OpCnm787xWf+FpX9JBf1RdNy
mVx7WjcvUr0lxLbbwvUlGVIiFelStFIQjapOj5SLDoVkXlTHW8eNdduyKlTQUjf0HWrhX1M8vvIl
6eCqZSoNfHlk09WraJ+2hu6iFoiQHUUMMiwkPQOc3tUKt5FWBE4kULctMx/cf/R1cgODohBXui7g
8kh+5TiUf30sHZ9PIQOERfapYUtaz+aqzZ9mjZbjbReJmU9WFm/791AhdSjzauCVE+WRsDgXR+5O
pd2z88BZjoitwXZQtB36BqpfMuicHdetnUS4hZfXxJMhtvH4zi7pwnxR0ISjgAtitzCt8VODv1AD
8sAUXTYvuIHPmzxVWuBIg35wpLJV17gm59Jdt4H0YdImxcHgMfkkTGKwG8bRV6JOfCu4tMxmcjiM
qaGXYsWooJK5SuqlxBEK+GYSreF8Jt25E3mxhhS/lxXvmfnZ9xXDOwC1Ax5P0jITdynWaGIRHiaE
fYzdTJ67Vnm0PB8Lw4XhmfZidlKnLzebDncUUbF0cfe7xZJYqcIXm2KyLMPEZ1vlfYRa2/yzYlEJ
Wl1UR4ZtG+j3QbGK50coPqhm8HKIzSlkuPjdPnmMbKLA5Zxvl5iWgfazsriZaGau3HbPjQ4ocg8L
wZDyFUK6n6NBjx8+iHgyXS1V3JXpaxN4EmATJMAqDk5NJ+XdG4UibKjunJRu7mdTwFUK9wUSM5s+
7GsswOgasrl05+Brvex0m/bIaMfRMmVvyqEXLCLUTjTYQH4gD5h96qAXvl44YPaXgB2UWV/d9eC9
XbTP20qndjs/DkoaeTViH54sH3H0GDAXGMJF5ZoBLmCC2NQoFfDrYBMvU4v7gG40yLD9z6o5uk2m
4elbhSukodF+ElaFAKv0ThcRRUNYRRtyY3GqhDawrALJKRyq37rKXohvCNb7TXvQyKkt2DqyeQrA
RC0ccHHNl3U8Sz81ZxyJKHrJrKPaDRQTBC+fkZOI2MrMqrzitXfnyJWbUOIqtVSN+nWXcYchlSex
G+uverElVa7s/YcdBdnMu21EbrSNMBTyHSKe0BoHyBWsQNGxwNWzWsapyvOlRyYxvQWWvKIf6K4q
qKL05nWuhGnJzNcEUr0rfXPcOKbuBMYXpfUfD7BZTWzjIh3OQ5tMVKnCHu964+9uCj5NmR1goXVd
1yneZhwhPlP75B7pnqccYUnr/3hcaJ9lA4WM8o34wBgwJ1wUrXbjPeVGaU9i/Yxgp4tKkkTuE/nh
avpt4Iogq3KK502FkdWkufBtGphgs5zDpYrrgc33bsaQL+zexOZDBZ80Gn/ORtOAeAjtVRXJay7t
fT1V2P+khQs55CMjPJK0dZ0Sz2JZV3A7r57NXOZqQAV6W2G/obH+LWjH2VYwcuEYrY74UC7j7y4F
mWDJEN6VlMu1DUTzfvWaMwcdB6favlfKGGPn81M99LLdJ3EikfuRu5E7MlNYxlytH0vTC9CSWb+I
OYBMwvXi8uFNMezFqV2a5nuZHistSy6Kbvio+Y8q/uo+fyZogPOGCOO04Scfsr4KbYNCyJ27AMYD
GmHsfXknuYCPJ6o4LkHEhAcG79H7YRX4F2TAPV8QrbIMKt3NqThhNqNErKNJV2cCpWW5r6cw+MHu
tVjkT/O7i/OYo8C+rdEotIWMW68ASi4LIQ0PdvUFOuTUuLuHQZToEaxa85GItCl+wJMFeg+FPXoy
JZFzytSgc+nY5p0Idzw/sWLzZeU9CF4LmlzmLULmeD2kt/yYP19DHL9YXqscUCgN3/q151prwgGp
gBCm3EjAdgaotwy4eWdzpfdk4jcLqB5vEKx5hipo4bCLnPs5WSaia6PStBOvWjxjp+EJG+/s8ZgK
7nL5a/LgjSLn3v6loBUrNRQkIVs7KsfVA3EQnd3mQMRPjMjxD/onzSjTztiaXfrhOyNqGCbeRDLk
NIQlkdEOfdR7CqsQ9qxeqy0ndn9znasIQHpdeB9mh5vZHQIBVcji7nsMlrT9BCN2nJVNhOOcniIO
X4dcAjgwk9vsyV5pDMhzB8z0xRQjThuQSRI9277k8kQCLgQGhW+M5Dmhxxu+rLwPhSNOApN3EBGo
6vFYKKfA8AVHURYzpmjjP+dHBU0EmmG19WMn/8XSVsQ/t1cSghlQiz1jojr1yQ6gRK6/bVGCzMiv
QzFjca90Bgtc0RJbjzwGE04KyizjCVBiemq1sABLZmNFflxARhWoC6WuLMKpJWvMS1dwoScDJS7i
TQ63ZoviBZEDsMEXD5Tz2iik13dcp1nHPDAOIr4hDlAGTdEvXkKBfYzi4x2eSpk6D9BWLqT6LOSY
+KEgjg/gDR9cwT+Q/pAntihI0ou1Agb/DK/J+HHYHKwk5IxK5urCLeKek0RevHnBjKXDJw8L6qtg
kVL8Wa2UgBP8nIacHboV5oa2OvQE47X+4trpHJRNsiWZVxxbowqci5A9jgCh0K9bKkRyqOOkGe0S
GO/mpsujrSY/e5IIMOCeTj5ol/LDCpREwHuNlCV3FhsMI5rUyFabIwh2AhVObo04CG4aYzXt6wsa
YhuwJfE0ySiiM0b9ks57A21uzmROzJCA52TZO+sDwxzhMdm/XD7ZzNhSTKu3J+y1sgs1uByOqbKv
WGcHky2fKFdfT6HeA2juEIo6ZsNBCVhFOnHye30DwwJxyNrx5JAS/sy7g77RBHFRC5/wWJJAN3A+
+oRkNkHd4XXX2tMnjvFY/S3/UiL1v1aauK2Ul3P1xVgo2yYVk6YpXLnQfKMAoh1AQiMmKEXf6wpp
azVV2uoSv46nVqZdlOgiDgZyAsV8Ib8Y6COo5tNQdmLlDMUbhpWtut4AQJwMmfUa9tsnuzBnyex5
kH2FNNC996Nxv/1o+oBNaxxWxlC/qm5ptvmd2asSgQ+VapJ4RfGGGIj/jcpv1/mKlBUvBdrA8Aik
pVXBeEAvJ/GijToyfvOXWsQS4qKB4hpNmxMiuKZ/b29TIpTjP+U7iGpJjB4nnplgIHbEYiS0lj+M
Alo/e8udqe8ZncQCFCI+ARePwv3t7bVBe04ikoQ44QNFHAzlDJvWOepAdoouox6EixavDhXeR1uU
Nq6a08i/Om4H64NqLdVOahUZ4cgQ6wGqhm2nbu/4rAhijco2LuXwG4DOrbsmjyPYD6qXrEYnf01H
h/Onsu432Rzz3M/QkAoDWObHPptCPNErQNlQFuEDDOxzOWW87jZmB9gQMUOcTp9bAAMMFHEZbjIg
UswlUpHFpx5s6wZbU79op9LMzyQFNRKA/duM4OT7bAIddQdCSXZRFToGKQJtVMC0/BRofKBr/SxK
lLc3nC3fJqf1ySPYRUZ70mTW2Xnb0ztlZjSo7hIFsqRFOZFrnCvRwzLgv+ZklbgHak2uHi3IyPq4
v/WbnSNpa4S47pVFD1retJfygrgHzrpqQB44I/6ULh2/JrRUF4I0nY3h+p4F9hDs+o+MoxDj0zFj
rSzTrnN25uslm7d0xbCpuM7NL3Dqg6unovFNMMMuAKsB6F7an8Op7UXpbw+RE8AO4fMfBJtzurO7
cKE0PLjWaInR2YbLtqPj5UFRKa3SI/HoHLP9XrxO7GWSdTJWe0OZ/ISdfS6MFszharNPeAJR4DPG
syolwL0gVSAYagxwTyznZoox7j1+adAlTzqY/6/qlvHOghkV6B5Bi93ThC+slq5w1ONDG2tFsyDU
vpyWOr5QsRmo0F6SkpzzIyfsqUacPeU2noZna2bCNWTZrYAeJcOIkNcG/OUPjKo4USaFf2RcHEfe
9LIxYkt8Uvi6ntRU1DaPtRrlsk+y7wjfTG/a56DFUAXXLd9zWugdC5Tup3vGl28OnEZiDVwtUb8+
eUYLz+Tj52Lr5xgyB4aD1StM2TR82pueamZ1y+zKBnAB/5I9iaicF5c88Ej7XK15cRQTPXSX5vVg
X3O2voCG9o0K2ZkGS0g/zS8IJ0OyM0UzYaee3Z2Qfu4bXVLrTNfQAfLiqH8JdC+kQSz/HOnL+LlR
O9W3Zi9g6kQNcCWqwI3bHuQJ+DndUw5SFU/OKvWQh00e2WxjWX9XxrXjxT2u7Eoekt/36gn13qKo
6IEvJ18p7gCeCYs9Qk8Y/LyvBhWylozwLPinuJ3f6UbuZ0aq11B+k3uVWKqdzwRxgplmyvNqtCCE
qFpwunPnr34dEBdj763mIpSrfd29DYBzkZezegKiltDDPiQkig3cuvxaqd+oZA0nCLWJNJhwsNyf
p0xALdHIlT2Xdjtjbx3Uk+czA3PeQI9Sx3xmBqfJJU67KiJf2rVROXHCQ2R0HPaHK5Igch5cXvLq
h+yMW9j3tiE7E9tTc4oydkR2lfpkTBqinwk4wwlMUkG8ac0DcU5mFX/CWMZwqXRabU8FF+Iju2wt
zDMZxO8fwo4p6ctT/m9mmJWDDLPi2NdFP9XkCOCJBy5NH03dWa0IVe7eAw2gz7lb5s4x3a7ygPuO
umi8K/3XQR7exu5bFzrXa5BnrDb51eBNg3imgBplgt+/0v35PhSEDTwj0hjjQAD0AXkdnHhwzANj
WY7csYu/wT/n3UsxYfVz0m7wJO3VZUPlpO+xDwqrXach5xV+0uYhQn3k37P7+7jjZX/agp4J7P9V
CV54U7rzaQcBFWxBkJb69DY9tXXS2VmcgjPkuh7mEV+d/YOivbwQww+l0z3hOKhEZOwIM8OUi1Tg
n4iImlUE8gisSyO9st2Z1PVif8lbbrbwO/1ZMpbMnpRLhoEWUl+kEd58+g6JLZSKa7ITbI2vb6BE
ESNKQblnwCgyFHRGapyKsl6kQNtxCFvmPXZ6zrIB6TpVL+Apm7V53SwJBN1b2v8306iqy2dbCQXg
lUifACj30LDjCcvqQ0TVISlc2mo3ElWIFRPPQopEYa1YRTyE/ardt5Fvo8RvMA2wnUmQPgdxvMid
ULf3I/YTPjUFUAY2SnywW/RP5w+lzL0oZXIq5H7Hz+H7lLu4WF3vkCHtORRIakqzRBdCHjxthdwx
dz1Ht2MZC8TOkV9AGGIPnu53NmMfm1KRWKVp0RN0q6J6vf+74WY79e5Gc+Y7eYYyGimCFyUNtm4h
yz6s4UvialINv3VtiFqTZD4ViKmZY7wa8UTdqprIAdtc/gX5FtFN6Z/y7UNQdQmkA91Q1j0cEaMK
oSHD+p6sy3KxLZGHSNRTZW/zF20fduiqI8tUqRTUmh7DYASFRFFfNpyf12Or8Rd+wvSpkiknBl3+
2lnH+iamy9QTj7KEyQ/c61oPp78/aTniRThwzJ/lJ+SDuF1jD7L7wm4wrsejXxKyifYD5HMGZ5B6
ncAJFczsJsAzcYDvLt2wMQTDYYbA9HO1Qhr7Q2r/dVmp+tWGvndEyvHLHO+DYzYo/sXJrMgZisIV
QuLgHIwN8dsyBb7+PBnsfaWlsJzrlPN9c5zQ7EZCnp8EJexGgezxjXHuiBDGq1/FplVieiMUtEe5
TaZtXmDekJhapgj7y8MtRmmp+ram6XqVjQORS+7+pRY2ASHJrEBKQYOe7W+WIg3o6won/t2QuqJ/
pp0nkgRdQdz1kTW+TQM1p5gp+jLSb2xKNL4Y9LdSFfXVEUV9WpMFR7j82QCFUADdgfV2c5LCejEp
ftaQiqjLgmHF8QJJhqnzpyd35swQRlgJ+h/Urnhr1ZPGYKzl12WS47ORc/qfe6o/t8+hXpqCmJC6
/tVpjJMsfjARpiSp9i1ODpUR14r1d1517o6aKzbMx+0z76FlntQFE7xD9ve8E5gE/Tc21jXR75dG
fbKLS9zRqGFIH7pkwUU52ZSrUqpsto2MWEG2mldaIGU+uD/qviNhJoY563+CYVoTts18zAzxHoDq
oNR0Poy9FnaND7dw0hlQ7KXDsTepbzNSHgAXYVgnEQmbfBXVfTmg2LpLl/Pi06iab9ouuvdVN/z9
PmxnvvI2qW7oydVl/c3q4w9BDwTuXcmU4wM6AAoehIEyUWhYQF8+uqPWxF0+L/GPl/TBCvwkuKNT
gEK2K8qrqbTOxvBu0xNBwUyGbLdOh8KwapX6vKeUNE5FXOpjXMc4RpvXuPzt0z9eNO/PPiGQPvO8
n0EO3+ugVYjd450HfTyANDe3ZzY7M2p8ct7xSxgsumhuE/ExzGcwuC8twRR9FkT1g+Pkfmgbogb2
M7mGq2/UZuekN2UYOh6JKuitgrKFRIAuWzn2xv6LjRwWUxqpZOFQgHue9lnsI3XOrBAjCFETfGbl
pQ3V/mUb5uVpvCipMBOraI/B3Gan0YC1HKF38/Bc2ujHvLbevlgj6WHdiy+3gTJQEwWTAqM+RL7D
uy7EiKofFxhNCcMPsoW5RJtoIkmodFsP5zMRgFy0gsHSGY0CdEGwQCKBSiZB6iatmx7QtB39QAA7
usXszwuKk081obRRpdvHVdt9gueNaC/sa8HavBgzl9jF68Ff9eLlQD73S7PY8Snhj2UYknt6vcYg
YNF2Q38U1fDt0abyh0iccSzmywCT7Bm/nCVWXU7jWKrjCZTunHyDb6AnEr+g//6QIwq1/1/wpuXx
IU9G3ztgTr3FNYY1I/uAJz/WRP8M7ICJS8EBBTe1WOijP/DJE1k0h+x5+bUpPOr1m9TrRD/xOYWY
xpgh4WyGD4R8738vyGcvc3YTheX61N4tyXKNiNV5yzQyokZltKIaJH/O21Y5b6xmTG+ZUoVIsNUx
23oVC6lUg+yYCYdxpYnwC32Te9Hmy40Qmyih1K2emOYOT88GfeJeASiBMMb+7bzzOdNdJceHDZe7
hf5VVJQKkfPlHp7XhtzwioWdLU0kLDC9E7JQH2GteQlfDTNWnI1OFZqeT0aB7jcuAk1Z6vOr8Gjb
7p9DXLFnYsSYOo8P6lGKK+q5PjBLhy9Zl+piGMZTLgtSKoEU2RmB+FDKvF4S7LcEOSvgOkiUM4mT
owwPgT5JnYfTae6MXZBSQmjNLcWYVJYypPhyVSqHe7x/QFljEF67v99ZNIFbn08REI/H+HnGdlnH
aoa7wdesnc5XEHxtgFr6mTqBKmVGYDeJwyEGUYkTowCJHq/KCcm+XHlaiPu+pWTaMuBzxbHRl9LP
wihUC+Osu3IwzXStafGupH8V5hcHfcGycuMr1QcFHdNMtSxf1KQi0SROvso3vL07Q/oicou51BIJ
u0CrqE/18HTtu+TC/0meTyjPIMxdDoY7OISCXtHulJThEpRwDVcTNxt/Cmz2olf8BtE+kcaGfvGT
1m0n7+v9fI2Ksg9VDYNVFFpgn1Qhe8IETNSYRqZzw+or/VeH+PZ5PdQXmM2jvSCqeppqqeA0QTAr
wZ8qUdhrjVOKnmsgzpCh9Rr9Vqr6t/n/EwjuqyXBNu61Z11Hvbm+0dy5R2k9kEZRQ6jUl5eJma+F
YEzk5tkjtC05OSyLugNeyu79OcTxcha5a8IU8ZpHKzoDIswPgeZi21fy0JPHFV9yN/eEC0hlWMRV
XKko6+whXW/6Dao8jYCLuCLXl537dDY2i8kKr67UYU1LEY5iBBuW4+u9HBRcg25UXQaT8tpAzOJ7
sZmWa/2R1uQ4Y2fu2pBQPVyxObC5ddU1ErzBNdMU13a7/PPMXCNA246YpURyQ2AisolrxqMjdpw/
F5H9fSYUfH1fC4Z9UFVDIfEbCmq3XQJ5Ko0E/SRZqMJ1R6RsZIe9M/7rktxsdYw8OyzFd2tQMra4
p7SAphA5ME6iI5i8k488etVZbNfxi5/ttTiPhg5QKlrR2EPlkP5bQByhFgOlAcpFyTgeoKWDGdry
yWCXWsqRhKFkkJA9O8EsFp2uROrgWfhLCUJJJ+bPi6EIlxgf9DKNjiYlq1RlvkDzhZRgsZ/tSLGe
URffa6XCngYqXopuM9a0xSZka1/mMsARjmuw4sRUU0NysJ/fnB+ZjHLA9xUB5dwbdoM5aDzaJIGo
P8z7Q9MHvLfrjH4S/EXEnOhABimNWmFyzrwrZXxMyO/M8rr4NkFS0b0rySmF0r35lY7rqlgoq9dL
SRla1bJLgs6Ol2ascOVg5mzvLvQl4KcExwmYG3cWuY7UBDnzKwNZaOiG4sAD5vJejDa7Narbe/3m
iQkpWzVcp1DnUqqmoekBReWuwQYjkExDb0THa8StStUrw9QTlij3fwXMnAeDiixcq461wZe1Duv/
tZDtxvda0aXSZiihH7s6Ro6nKgVuHIDYZjoqHSprTmmD1uk5UbOMiKDVouNKjwvGfKkB0+9xIuEx
YvCRJw5fl8jAC0Gzxv4T2fpx8uIO+39qy1XazjhJjZZ8fqRXeYT5/Qs5fmnrBFBbN/CTNFCYNWbZ
biXNOdFyCRncNgrtvv3QAdi0rnAI+mwNHaYFok3EaEGjQoBzACsEylbgqF2E9dhsW09Vegosuc0o
kXJwdAxVk/pw72GdGa7JEj0iaR9BmJxW2BhoiYwR3oiWLYCmnBeUspQLInQc14r3oA6/aVAalVQu
kVUKlhC0k5cRxwNkD2Oy0kpVycklqlYdyVW7k1a+ezoqF0EiM2XNaGMVdtBJUyTcHIUSA7HG5eZ/
46PkpQsuGP8vqtAFjOjnPKueXkS2UbqWX4vfDOCqVG1e/L99I0U+vi19yFpE8f4erurGHoDfWu6F
RRkfrDGsZGbCh4uJLFW2XjngcFqW7ON0ZYCY9d1eLBq6Ti60FsJGQFuNXNXesMRvch6xFda7Viur
86CJq4vqL0ccUGSBJE2kjtSyfzE5abPDS+ebuKdN9/Leg/66u1xv7Lyv/9bzDBIWu0bJhPFBnO2D
8x/Qbb5qFpIn2KQ4n9neRlqP7e67wfaql1jxwhTvLjPZw8Ixq/z2JRkfQQc2vHjIDAXdoIyQIsuq
4Z2C6iLXRCH4mxaWey/m6oKc91NTXbCHDaeZSB4hHJJTnmklQFXFgB+2qhcwrDHNLTmcFhbk/fB9
r8WNNv3GONlOa2EpH77oA1LXIvB8Sblzw+a1p5LAl13FHRBk7HuSFUIrz9eY4w6TXmeo1xIyppLP
WegtAsCczxJzLwa2xabUnnPZc9dfA8PbRcPo7OBWU/kclGJKhw1WbL/ZcbbtniL7jU7/NDIhN0EQ
lastwxX+qn+XIQUrf5VD5FNyqpC5jkOxumjjHayKg9gqzQ7d8pjjl+ErMN20SZij3gAgIiv23Fwu
CuevO13V20/bMJk7g+ehxxCDc01IpeZpYaz5I/F7dD7bTvIB075bD+btgGM//Zm1P9vnOWmhSCld
PzSrfC3EX+YQnK6+5jYPh+vawYCx1SWwKUqEkMjAABGqx/sYqQfs/aZobOr4aCqVRB3XlzC06rK8
VFZ1BuLjvkmT27GVtPy2PVnVNXkMv2mSzdio7BQ46ZjRkj7Or3LuQLzxFHz0A4nAJ8jwj5UDhvwY
iB7msev9FuZiDU7oXWzmBH7oc9/HEHb172hUzd+YrAUm6EsGox0fjrcV7T3zILAk8V7xnKBVyLi0
UA7sEZ2dZ4mAIuWK7sYUMHw3ofobU+JNSsEsT82yZ+ny/X1Y2ApuATr0Kk3EpU4yFVH4rUocIj+l
pboDe8FxyaMXxzU8k8cqzVmBgquY53AJ3d0/Ug4hixnMFOPRdPkVfgmdjzuDQmbhfhwnTnokbutX
SFmZEnM4QBnwH2EaHWzLZfA6xASJ2VeMl2gB5cmX39IGISVKL0zlETb8dXarTS3CzLoWkwDNwsnV
x0bLK/jvbbS4qm9luaSI2QknegVmJBw0A5rqFgJab72eGfOyBl2HhOdFClaaNqTbVsG+8yOoYu2g
3AstWp6BFnzwxHjH9viJuyZRo6VEL+l+VlDX5zLvA1kwrUl+Wb06aAb1yYJB6aVAbRjI25SA2CWf
uonjIEZchz80PwJ4Kk+/CItVIqRz+21iwK0KlRouAl1kxPCsuqVrmPRRX3fHuNhJMq5CXNCtyn2S
FpBpNXDCC3zy+mofSuD6aYdmVVgI5xfv8DP89UQeOdFHomC7vyhEir2Y8elexfXb5n3ZllLmGuA/
2M5NdYsmVvde7U2LIdjWGrpRvpksaZQKpAM+ztqYD7tyOCiO09oiJKbuxWLv7WCvuUaZRMky9NjN
OyRv3fbuQZeDIFJ8vb/gB5SjOtBn47BTbaTkf3oDGWCy2q4ahFRz+KZdFGAhHhnnB2Mw1epbuAHG
cdA+9cYBronulEwJCaA8o+6Lna1e7045lx91WB/H96CH6FvATI9pvQb6LUclPNWgs/eVwysARe90
dsuLRzVfA/y2VR/lZ/kMpHBawV49HgOEUTRkpWz5aOnqefCz0VlV1wKuUOChaH8A/0QeLwqAZs87
S+e5bLA3W3zfLT+6o//aXFGV+jGLBJ3/uPCcD4ME29dbKUUzHfuNaBlr6KrAXZ+1TXm4KqR3IUP1
B7yJAWkUa8M77zACRgcq79CBcu7gE0uMyTOCjiZGAPSn+pH5ZYVSkR6PHPeOVwuOAz1Z6PC21z0C
d9wXDuqyawxODlY2lnT1u2QBD5+OEsjrCOYqrD0Vw7lZw/NT9iGIi31z2TOan6rpJFbIYamoPa+P
A+VI7BHwLKdpWjpjaZpvitpUQ7yc0zkjIilx7fPjE9WDzuC4A0/Z3KEBFj767zDtgAGtYmOMsFim
424THUM7F04OMTJ87C5BHDzEBeDB57roskjNEpBYR7y3rQeGMuPNFD7m/G6v4eji9V4w1KwqrgCd
nD0WZ5SBZyKOSHIREWRhEXqbT43QGakjGrRs7YVE3sRUbqsSHomuqRLtqWM5ac1mvrlV7WXhZCXZ
jRxPgjr0J8MNjfiVElG80oKFi2tjKLAn+0VStVvFhuhXuK6eQdCeV0f83atUIUm5ZgX+ly8XEDJo
wefE+RLyrqKJDCwE2tjABshO00nISoaDAewXeJvCjDUhhHywWdI/EQnGwNR0wOFqTLBGYUdokkBY
NPAXZ/uHv3u9cCeggvRfsiJiPMj94kKXJaBf+36yZCXGR5HMPzaQhz7GOFRG/cEB+ybuFJdf5Z24
/1rehJsu5+6NYCF4+Xnn16HzX4LKy0xn4l//BktBeTg4xIvD/DqSd2kEU824xXJlOZ+qPZfMNf2s
hn0KNSDCcF39fo2LyAhQbyB8tGA6LTdatppqXamc2eLuJlvMBezlwnd2AJv51Zz5AwtytlC5C8CE
IszzQjfLEPP/1A9/oTcgBABCluXPz7XQfA7SauRIlFeW1rKMuIVdeHw5SBMvVeIQCB3Rq+8nxUHo
HeySKlD4l1T71rpSy22WGxTti+S22qJMwY1pA8VBF9Hyf5gTZDn4fX0CcVgPaLcYznm9e9Ni1k+C
BNA5adJ5J41yKFkG/W5az2eCE3+EtJDPFWAZCFor+66fCQNjZt/gD+GGGuhWitGnvE4382f7LDb5
MiOjW4i1z8bG65qY9ny6KaSsqdV4JJy48EhEiYeOjDfsoOfS5gSQmoYERiUgSnSYNBCLaF+G4gpk
sbpYUk2lnOFWEaarszt3HGutK3AAUiJ6gQbOeeLTYULcceZkpcnlm5VnCScHeES5N03/uKKdFV06
ck15h0yytMD4eYYzmrkHD76Sj87i5BSliz5dWss3RBXw1D2WNr50FO5QHmx11EgPffFDjC6bwdI7
SBLHyerkKxlgyrVHR0tLv5Swy5m8fGrbl9y2cSSfZxnX1WHuh4D/xccPmsQOb2C8q39e8uqeb6u3
EbzIgwXwMS6P1GxPWoF0mBTYCYM2vzyYzU6mN0Hf0QyvQanCMUrA7VPMzJkOt7mbUdut0F0LgRTx
WLi7L0n9NWrQicpQANFu5VxTE+zr2mQERtmDVHJhl+y7PUgI38gWSBhhSHaXYjBRixoDBbobJyZB
Hlha6Bmh9vtzhIemTkMcGmzCpv8GHYFSdso76145KlwxOIihUzP1IXyV1tycOkbfbQMC9nqysJib
BrRbvjuFpr7s2S+fQ6WMERVNOETeqRm9qcp8+bf5xyS/mBPpyFv9D69nGZlsqGX+5PtOVr+D2LUi
wBUtOXEk2aTCuhq4mD+LdD78rtAoOf3nSuesyEtlIBkpl+ls8jN/anwcLiam/Aoq6BlEhJFes1sb
IGTlR15eSSbG/59P+BveDwC2k6fENDhLvKMhV4VA4eBRRYazJ6oKnQSph7VGtLVODjl7C4gJFWxI
chJA8WUftZPXD1J+9Vv8EiKOn3ezOlkTTdrGikSg/t8wGFzlMkpqCmQN+SSQm8RdC/p6wdqShzjj
BjakAAu8epnulmOPfQEebcCsaW7lRtF1oLxd4D/R08/F6PPzP/PoM6a08gVE/33D+l1e+6314n+1
t77Vy3zmTDSQ/3H54AKA2htFxXV5iMEGCEigP9TZE9dOtFgQ7QJCP3PMa6GykWaFWrx9SRa5krP/
dhkIMK8oiGXh9zupiVMU2+6E2g+kLCAMToPW0VoQbHXOD0k8i2LaLYI9gwIE4LK1u7Fsp5lboOCx
0nvRMF4oLHqds59LjnuaXoCsB89PpEZnx8KCjg1eGT14JS3TLJ9YUOJVV+Ml0ygAcG4hZJbV/+6Z
gdFGrVWk49bzhDar2uKeaj1C+X++lnNuPqMsJNKFWaQW2/5qip01kZV5InpEd7wp2yLfXXfoBDPH
VfujoUBAxcTXBakbOh+K/MiLsz6/P/QQyiBwk+An+0/DYMAf0Id+ukEqLsAZQc74v4fwv5Vg6YFJ
DyMv8JaxzABlKb52/L56Q4pWZ20BB0R4nqSLiROu5+pFMKnryb/Lw2ApbJC2zxaqrro/RtIDxeEV
ifHFZVs8bz4dV2U77/G4r5XXyFKRjJ0wrdPQ8YdK2EnEIG7tmaeSPAh3rg5rkzODN7+D2EbwzRNE
jM3go4htR8SJbb4217YN43AJuY5qS0B9gCytaTefzVTssURLvvryZXJE19L+ZyYhlQ1kHg89FoLV
ESJxknXKmzJfrF5tBA9su3D9mKfiaYBNDmdurgag5ZJ/ehxqPdWQZIqjPBeMwm32uWalEC85sj2p
3CzlhCX+t0Tt/oEAcHM4JyDKyadDb86DKUCAeVS+3HvFloUlH+OWsgPiimqE29UgShLDvBdR8JXH
hh7jb9fXMl48blfb6hr5pMYZ8kS8SP9QWSRNyJbSlX+Vp25u6yzBFrvtx8TneQOUP5qYeH76D+6u
TBn1WmHMeWCEuxR1mcHPYq7yFIDWduNZnPSgTYhLfwVV55ORYt8q9WM8rGVGnjrdJf8Kln0xEJqb
9M1T0IutiyybPafMXthCKpxzUBA274tV19msRGH8cmiJMWD8Q92tbXW1kriZvJ57KXl+aCxzdLO4
mkQAxUa1O93NzUDcWKAtdGYcz90ZgNWhLnXdOi3TGjD/jjwQYlPXll3BRhX/1WX37dODgcwC4ubH
CD4l2LiPzj7VOPqUTi9YVWtndxZy6vMab+R85yi16tbP3oz56QEB/NsHmqoksphfmUVIbuHFHbMF
y54/srTxIjA77J6Ej0OG2Mltby33tDcvGqD9PWeaG0nBzFpkhV7lID/wSPJRYxfeK4yadpDPb8hn
WaoU44s4y7f/Mnd/WBg1cw2yR7ZFTW9Pp4IN0lsddQ0GFzMDaMAsTien4HHsJ6LXPStmJ0iT+zYU
TP7dODlZL1DDnxF2enlKf9vep/HzZXeV//rNOd5VV0/XshnQkil8Q/BFGYupwRpDLP7T1SD/TpZh
520YO9hstRmRvuGk19dQkFTbfEXF5GsEysC3BTh1/paDxesbk/ofqMKSxhwVmznr4KZDfGOLxYAW
4QQQo//dIUaUy2unw2DehZNN+xoWTreUug4EClyH4KzwVfSBcOqzjRSKxWtf2msk35+UXNEPV+qU
eNZ5/umfnjt5S8iGohO85zP61piQ1zCnE0ilfy20iGdfIGfLViNe8piyvkNHzQkIbjlE4OgG6C/m
1Pa2FTdzg2WjKeam/teyca7QzLk622BH1dKfaaCsvept1QZdf54n0A/uD+Q8Exf7wSx8HvjDCYE6
WXfzhV8ry1JkbMr5g9IyBs+H27N53OPLvisV87F1D/ZYQqgMDPy6YnHh77kl3EiNm2B5vUyHBDO+
y19Dlwzt4T00yA+X9c/3NAB0z7zrfV3KkC752tDJ3/WvnsiFL1NWIO77FYqQ3JnFPyW/YMC/Vh20
UNGQ80jaRLztAMamJwjgtecKEcELwVZFKrOEk/pzYwH6e4m7gkx0bEEbXkeFqNvZOw7PAQ3T6r3e
nBeGGBQ5uwilZl8K0VQYlVbWU6ZWkRNawT7KeeLRL8u4l8CifDJtyKqwT6UegoeBxGYH6GXxNWiD
T0ZDi8gu19pEH8O1Ze4epgodzB6g2kzWH1RJhqrMRwmDtLsshoIhJtQ3v+ErZe6jpMweqwh9uEEl
7pFwdJYHUFmxR8v3w+fZvxBWagOlUiGJUKSTNYpPhx1KA+7laaVkDRx3kF30dvWHUQTC6CsR8isd
AMO6m1YwfUwJTNaNTa+YeykcrKwM3Ksy11lt3Av2h1XwRWwmtdRZsLoDsx/T8CB8BUqy4WtMIuhk
4pRoquN7Uuxwd9QjmgGmUTzUmR30IDNllMyiFnUFn7xj9ncbNs7WZ4DrBPV1vQmAdgwSdmXjz4Xn
s61/wgEusC7zo2gz72Y7ToTc4yK/BGPeQ4Mm1qMvwi51Hy6/z5z6YaqUlFno9rSDYamNRbV5lC2P
kT0aWtDA7OHbmLq2ZJdngHy75LTD4q7qNl7kAQOovmtnleMJYc9jEtXPWw1bfW4OxC02P2vEcLUu
lB1tqYtaBuABk3rt1TBePiSHg08wzF2oKhL5Hk0MRgaMHDftoMbU58oPchyjIHRyVorFbrhUPjEX
nQrvjzaWtN2ZQvpobgFEs4JRuoSEXBzmoX0LMjo9SBO0GwYi9UM0mhPZrKAY96xRd47DjvxeXSFV
CSxSzfsoBrlbChgVF1gMaL+aAKTOdUgJE64iBikS7ocOzTjMjbgjbtSQjZA+IgNbUD51UwwVS/S2
N13FWTC3+g1ye93wl7xSYXhjXh0FPTH0ZDOLieLwBGoIqiWtYG8ZN9o+9MOD+PKTODUeQQHsgDrP
c/xqP6y4goxJjZlI4Ku0PBoikcm/u7hDOVZ9d2XJoZcw8XxJQDAztryUIXwdsBFD9zPWLB2voeaJ
ViNlTrzOazy7ElBo59nFvA+9yfr/HhrulMggfMFy1mqjTxdcXu+RlXcbLNUjjPTSt2RzxxjgVn6U
lTLrd9ZyR5eSAR908uafUBAiEwvAa6dQKzizrnNlkXAkmlJ8w7RFyLCE0rCrNRVz6Y/VErEyoaii
tp7XUE82vUVXKwW6B1zYHDTp6CHPyfmXjKPGRnFVfTLCZ8RiYfC7q0PdlZ50Q5PqmoWUg8BK7TGR
zCrmyEBfP38SVnVxnujhZ1J6qjmfiaMmCWuGbbGiCPx02wMABgMSFwhrWu49cNmMWrw9mgOQxmHL
Hyt/dfzI1HjRTMopv67hQ3r6vTDtHupbP0MnDKJpI42BRN5LsTaQ/n/LD7xbKYQ8az5wmaTS4Afj
FotMJ/LsYdquiT18+AC6uNIQuEcC2hrGUY8zq7+zAROa0KyD6rWBHqt5WraKmDgxj2b95SH5w4JG
O6VnUVg4bUJPyFDIodfhCENBrW+NW1WWZn1eCWjrDxVeuWoUv++X3zjsCJo3dZwzCjwA0AI1/HNo
UGdWCftxeeR4yw6O5cjv19ZjNRp2wJVA8i9j/WE837cxhCp8vsrFOYpJqbYp/2FYfJ+xwhJLJyv/
fwTd60ZQzQe9eX5iBbmG0U754sJbt6DuTLfdVKINZLxBJ0C6SoczCAtNP79p3gY4nJoyqdub0VCy
iX9TyMXN+jhPGE6SmBDm7BHcOWpqRGDYztuXLV6jUQ1KG3Vkc1HnKZ/j+XT43hhf6FzQwmZsjxDn
Q9V/i0vWQU9sNLBG24vTu4AkHAy+juuxNYMmIJsAOK/t2bkQ9OHo09PdpaM/iayYXQsU/7BFSKV5
4YLKEJAHFeDOX0UdHNZtfWstLkMpMeHHCT5JMwzrrI9VHL4+0RSIfOOtEjnLic3agAlWGyGtH7p8
tJrPeTLf3Z8Wqw2mYHdvRIwB+LwQm5BF2MgQ40Hbak3ZxmNUuTawrVLr0y6vbQYIiivtcSv55uAG
wkDOsza5xVAGEqhEqzKSj3KEKB25u61qodOo0OU0y+f0aSZ0jKmU+UbCzPex8M9HeHaKXnYL7R1z
qxbQLCfxP2gekbsnE1nd7mVT7Piy7Iu/plYLyVyxOKsVJwG+97yMUsRe/mbJF1tVd+9AhEFHHNSC
AmZTm7p5vQ98C4RxviwOvNPCNI5RUFvWyFzGAo49i3H7Et6IbKBy0rvTPn/SV+wtllHBDF17cXsT
3kLtP4Mcs5ZaDNhZfNGsEltf9771QAqv1JsaIkRdAYGrxHk4gRIVov3VMW9EaRDW8sE/l1Q2e+lW
x5GwDKEzMCbjd70r81G5SnpZe6XmqeiY6InZBAWOdCOGU0li1yznB5+wVpSkoRh7eF/Vg8Qi3E/9
lvuK9XuYPIJea/XoleYtF+b0WrewLk6Ywf2psFLRtXPMN4Exnt9qidFkJbpHyBDsh97PJsDbhdBz
kIOjDh47z7sFoze2fiDNZcJJWizQOC7AdZmBvGqRTGtamfHDit022lFcGRDd4DE9OG8eVFnFCmyb
CmC4XwX1SESBgmD+d7bRYg6mubff2hjrYPXcSW4QWZmldHo0K/b1kL1dHE3VN/baLLwZ5Iqf24NO
Qe8yaO5vdEJWm1fY110aiEObFGscVk5L5N6bnrVnPk9Xn27urU2Zmev+p4gTs0rSNdvEP9jTOasQ
3+czwYqQ6c5qXSNs1FaIBrTtdM1IiRR4QEPDli3gLH86pthk27VlFCVkPdAv7cbiRNB886J9YQ7q
Zb84m2knfqNd/Hqiny3XQ87jlWek/b6pqovjCpKj1tYv3yOT2ezGroo4AQv5bLnO4MfY/EkdkB5f
YZ232PtGnG42RciamcxLeha7jkGR4wkxAWkmPRbzhoILEvojjmR9qCsT2K9M3tHU/FTgoeYEevCo
HoxvUVf+nhNJkl+hg8EPRrT7wQyyiMiZNDDXaosXrODspsBeEmQWGUl8zmJMW5IkBctlsY4U3e97
ab3V4c/7DeVOz2Vk/A7+FXTbA4BJ6H1AcJ5Ggx9SAuB8yLuhnj/mUjOtWmwsdcacogpmWO7GjOcy
ec3/HHlcirb7gb6ojeu2+NUzSPJkCAqzXH2NoH+oyt/zl6zuz9Dni0ZXMhe5Ck3sWWmrIGjdHSyd
8ntT7mgVQs98lwyr/rDE5xROv+FrmhjR/voVKoVRnPFd6K22G9PLrcErx2eEFFil9yOqRzLAONTi
xFB2V4vM7a4JmCRjm1g7D8sHrr1OzdlmbBPt/M2zLWa2Jz7SutiOpI+WCQqlftjMlaBgn7gqxPGf
E03Tq0fXSufwCDtNxh8AhRxA1evJqxZYRViP0405QE4n7XsD9jMIEPUWF2YqG4J6cIDikKAVzwsj
ITos2v+MTfWidToES0eP6YeqqzCErMzcItCdIQBxMQYR/cYGKBQmWO9y/y83jzB80IqSFwd4cRce
hlqQRtNwBfRgR0PJbTIF/wP0GcsVeG51LnvKIHXg4LixIT+Kba7/JcTbSbqHD50I2UctjM456r2+
n8NPX/vhqJ+AYDnfuCnTKd0spzwbsVkeQhGMPwBZWC8OJHdkF8kWdmQZne6rd48En80I1z5zy6xs
CCXvwvGxjkbdGEEq0W+jClLf+hl7WmIa3s9IFeKWGE0i4Lxjams/u+cJnwIBb25I6t+m4W7+dVg3
fmtTeatqgC78JnGCyJnFwYUchJivT+6p2y+qjZzF1+6U7pMh87FqzTHF+baRq8tPKBFKGsf3M9ix
FgoiuAIWzlMVcM9CcuS5k0gHUMDoeRjYF//PYiWapQSNfLB9R6JafODRqOSxfXTagD7P6lBG3C8j
v4bFsDKSyk+SfR7kpq+s+3Lc6sWcqlO5WtbNG3GJrVASfbtkSl9L7FL1TN/3DNQ8y+IJ/g88+sEs
B9h105g/6WrTSF8gj/pRfrtYHvOedByBdNEHjyoMnJMg3HnhWgLswAfjh/XpqaCRCUESKZH9bxAq
EWLxk0L0baccW5gtQlP1/kwPxtlYBBByP23Gv2f/BFDgOxMg6CbMREwaAWhl+y2vFJN+5biVH2p6
x2WazZdZFax3/WlMLoy5izXTwV/3M7/qP67mxyxXYfhWXDz9nsNtXDGIvi5MK4f2XQSnc1UHqOO/
CocHwcOWTUaoebBDh9GkRKCyzDQGNr03TmxHhDa9b6LSEK/fnvoMQqxU5ucTqsiOYIIZv0RcVwR+
iAkjiqQJjgF3vmKCrfnQFKKT+E8HD3P8jIpUwlsBmGeV93su7hVpD81mj2VTw14oqwEVjt91RDtQ
SnUoTTUWtSDdS590dAhX0RoB+p6yAA5Bqa+jnlquJCskPd4O98HSEfpoe9ifVlnVCQbJbtLpgb1C
KNZkfUx13WfOEsgZyYxX8asfbRi86yvtzy932PZ7Yeblt/iS1O7UWPt8BlwCgGdzsxeE3RDFROdU
uI01lO1HFIPJLCpmSN/SKLLKI5d+wqLI4z5t4HPDShxH0O1h39uaD9z4o57f82Q0MB3ino3J5DQT
qR+IVHq1EQeEDcoeZJqKOQgtBdh64Z5ZHYeGBYIq3646p4if9/SX2gcTWI++xv0To3EIguWe3zNi
NZ5+Ls7sm3kTQkNbJEF6AqvtaZADaD0rewDAyr9a4/OSLvb+JfYLiZFPwh7H+wRQ/fWS+1Vn5Er9
GhdtRqDc55PICMVpWUkoBVEwoCMGL2uivKVM6bdmAg5SI/ho/DjyBIHHpnpeflhXOOM16ZLd4eus
o5Xzn4k642hOGt5bcHOXAKzlO0gCR7B1SBaSMXDG81hm5XTlDiRpSX/q6q+maletEUdipqrsvtKg
DVBX//4qbcs39XmUdF2w3dnCygGDnIH7zfFG6TLog3HtFt/CCzLRfa2FHQGERFAr+iFZrt2pmaWi
AgY16Nb+Bt45xdxTtcDEst0BYa+hQkAi4urYEhfz7iB7nmIajLfNS3gmW8p0eGVKGiOf+XRTRTLh
Y0QKI6VMUVKXeqWIPTIJa993oxFuOsrokL0U8UqYvbN+FTyNcrhcM4X+e6PCjPPz4B4ZsYZKYj9h
wyJES5IvFY/0fbloM6QXbh6mRSKQyt//HwCctZvdY0iSunTKPON0t6VZcuWdV1f5V2SGlK/JSvsx
Z7tvYl5s6wRmzQFSs71Yel7hXYlHDMp5RW5ZPrWBF+WccPaut9LTW4aXgNHucqEWTed2zbC4kfdi
P9lGAN1iDI74yFwBjP/8FOrZUw1MDqVYuTcx29I3LYFYm99tXNyOdk2mZbCpWQwQjq7sQ2NZoH0l
EMDPOLpYrsNpXLqVdXMXIBOcWneHUYcwHZJ/azPXnQ7f8WjYS/UJpzNRP2exkfRkEcCFr4Nk5H3C
ER3JM7MATExaEm57SFHYUkCgcU4eJzRcRz1K8lVgqxp1Xsbq/uXo7sBb76Opq7ZTqsjNzucmfh75
5hf8QAl7B2Ia0rtICy9PGLLrs0V036NduAwDnIFX9qxBqHMWHPO6feRZV4aoK8K4wox1LFwpk40f
PFFoRE7lQa0Co6VciBLMaFMF0vvj2YKsgFNgyo6c2qT8iYz8fwJUXucTtuWhfdTe/4eFA19rpm9m
xIbe7JXQZ+bhz8iC5lOAjLrwQtokUlD/Yo3Bku8bTfQN8VGRtVuWRLQTcIRuoZsj/yJ44JlMfezE
N+ieyyo0R+k5sv1HJJdL+llBNMhWqS0m2Hp6CeA9SGDamV2whQeYPlnuPAQ8qpWQniotx+QPHzfN
gUhXWSfocNsEUV12J0w1MN8g4tgU3p/6ECCg+uQWHIDbIBm6PxFqshSFOB7aIxjQQ6gCSKkCG72h
P0ftblR69gQZD5SojRZnKHjRjfDWNnqulTPGeYzNy+YHTKUxn4hoid7ZkHEvEabXv8EfModwJ6Nz
V9j418UIVEMOWH3WLGnLyja+DbjK3DQjRz9odp/pxurmCicW7Q6GZpb3KTFZ+nfuuOYoeac3369j
+Jf7i2I42FvsfJF/mw/cN1QTcEgLwSmHG8y9hZ1bljQvK3HHu5eZG3e3XRf9XdLZuO/xqgJe3UJh
wqcbvnLIYiKwSRMDYM4ZuHo3eo+SacB4M+ZTX7YVdY/DDswqhvMKY2/4LswZxL/ExHV7ZLzEHCmj
nIY7p+Yq6AAau3D2+P27iQ/BEXCYbNAXkiLnHBjTWaKtjNsi9Lb3Y/6qXQa5Pt3uE4NVbOoA0XdD
XFQHCvM/UbgX8o7J+YbJCu1hVyfVpkRbpd1Zj5QO7dC+AcpBHTrVOuT151E+bT9Fy6Lgz+ZS0MBQ
q8aKq6Wub8bF7CISvOZI4sCZvf6owsOEaS8Cw+gBJcx/Y8pRSi9f5reQj9ZDOOmUIH+By2K6Oejr
+7EXy+oap7bDOkJCLg+jT4Uq6/eKLd9NnxXVzH8ScStfqerFySiFtfuPu3jamh7i/tQiHs2C05Au
VeqMWi9NDvFi6ujieROPqZVkbg3mONBzj/Pqy3RkUhPhb2fKpr4Jy65AJP501FGdFvccmyMs5Kvv
XwUaZfO/7qOEyYe/NkRpy/voaPRV9jQpcm5a9xPal+ZvRxzFHEQb4NucxmlHtXBOGsz8+X+CPQAB
2ruiWn59byHo0HrgYBsf1JLgCLvJuMoskgGvUrZLGyHa38oE8wCLRvUILJE1/C7dKb34HwOuQkQ+
pAKMwIOTipFOngPV00zL1ymkL8RC7PcwJVvhMGdZNv7r2uuZ9WV14dEYLSDv3yN2c0MsFoBV+nej
wAKg6hfF5Z90HffCS03+uWmCYB7uStOULmGUGVrTxBuVzJP4CmtTkxzZA3Mu+1/EsSHQYLaYOt2s
V7SD+WXguaoYiGdZPEAAccYe5OD01Z4cnMxHgnLHlqDgmm6v8hXxF+wctPADbrZ3p+JKdViFGLwK
OOMqYckRqnytpTFGD+14gkhlx4oU2xVDmNmCaJrAG0IVL+2qmIQIHr7GEk6zpFBJv0UO5qthk4zX
FohSj761tk6NvuqSUGJIt6u18PAM/8L9FbkS8Wd6qREqOFBuLXEHH+lLTAwFspF3p7Mmmc1hZt3h
2bvIswWksKasNM4nCKWn4aNLk+1O1YDHHPYLZXhiurdf4rWIXPABV5o7oms+22jnvKraR0NRwgB5
09EfBVHa6uy8ZBptZCycc+9p7uzW7j3giBr7NnE+az29iYoZ+svuuxp+BxFhpdSytw9c62+jdx1K
pw/rYMdsZPnRJmbDoMVWHzZNcSA4lnBCCDJEPTNNrEwSUQS4qr6ksPjWiK9GRgZDwa0e4SjDhBO0
JZQPkTdpYSPa417oQgSVWi5XKCnwgw1FvbSvy4/JF3VwyykZLrQxGeyTSH1+UDMdN74SSe50jzXf
WCQvSJXDm6d0SJ0UjeivCxJlEl6In9Kq2keEnFg3b9Gl75rNqA8yVNrElU4+PghuTSsEyl3VMCtm
lgrB9NWOTqdW8UZ+EXl6G4aPtcjfsz2ZTWFqbKMksh6cNY+Qj/KvpBNJX4Aq9fzqQLoGhVQrSIfu
qO5Kp54lUJJ1DgfrKs5VpLq+4koy/Mzyb/j+FhLw1os1n1Lvu3QVLHZHZwXVup4INTVJpxqU0HL5
tmZjjbnoHrnkh/14j+od68NMcwQmfwPwDD2U6YNvQh4ybPob6jD0gCVzRdKOiIuoSjsnHKqhR0AS
ZRCNvaYpwZzOoJBR6ttJq0e/tMRt8SvQwt21XCH+bboyBX11sTQvFcQtWPWyc5AEtMDZR7a8AYme
yezpC0/KoqtggeeIGOXN6LQrw5kW3Um6I+6hc+XD91QBiyl9waksAiWHeWxZ4yRJS08qQk4GGeMT
1tmfLoL+T505E0qMoNXFOdBjZkcSoKTsVjkKMQ5L31hhn5bXzKIVcolTzwzpjJZe1dwrvgcu7YLh
YqQD8Q2tN5lw7znNNLf7q4uXpmYOpVWqtSdYBoIQTa4LtPswo50fFn+Ty3WqJT2GV+CU22w4ogbl
Tdy+kmOTjrf6hKlUjPlOXAHYVAA2MNIy0NQpwNgWzEasvvpgHyGKmN/u88p75+6DGd6LOpKyb0fv
DO727q+35Ns1PK+GkAiHj0VcNWTP1VbSHMxGPL5BP3IqFOLI5fG1ujsjoTTRmxvd30IQgYeM20j6
quf4fQEt7lhqsMQ/Fwwrfe3hieSfXf5pZufpeOXxG7RAmlWHISdoj8VRvK+REN+u8+iKpEceo6ai
Xy/RXBgqLji1RcAPDgHbwEfvneuEFrLTQklLOqgoCOSk3S0k7wd7QjzC6YkbHk9YASfmtspz5wFa
iqSJQ+x2HAuK032DholoHtUhooTGnfoEDJpuQJ4y+WOyevKpSTYHZpl9FzclNnhOiX/OYOGDZn1n
cxTunG2AhQ6MzIRaHE46VLCY8+Uv1vRlQvoPrB6KHS3fMeB7OUF/xrIlzJn89+1mNxOthzS6qjAS
ooyeM6fMIcZwn7kyw7yLnzRn6JyJFajSi/Xi7urp7H/HBrAB0Xhk0rIGw97zRZIK9/yM9Cbkbm4x
+o8ATI0lFziqSMqnKm54RSx+SIqO2jlyeqz4ZBZ+7KyjwzB6ls8AhxhMvR2YyqmpjQvPd39K/osq
ZRecsaSUsxo4HWQPLn+aI+zNH9Y+iTbr2XMXbb8Gf5ecP7Q1IXTzrUyoAmgA/gSWVR6rhqH6Irne
7vKoNBPrYEJeDj4bKRuMuKDrNtSha0AQ0exHsl1hVMz8GG+0Zmf8+MfCUFS2SenvaVPMuQbxGFV0
jJyIG57IkgaQ3k1TtOOuici4JJ2NM2Gi7IOq6gaTozhMKKpMm2EhKlcslR6k3SaKVKR9G88Aib6F
kmL69ZdkJ5ma+m5jX3xV9KyrCscG3yYpkSx4cOXH/l5wkNLy7Ugw/MLmraHLEjq8M88aEv58rTCQ
tFDVDG8COq7QaeSRETLssdNtECj4a1UoHLcilEfTclUB03FtedQ8NiZGI3LhiOkVPRxSU7JJEOjn
gCzVEr3fAethO0MChRgMUEQgRI2jK4EVaHFhp2/ftmZPuoHcceDcMssE0r5fHqjBROhkY/ZlWN9H
Qa5UUwknjjC0GJpyvoR78x178lLcQNlXBeKq2+/tJ2Rg+fphyeoolwQzH77XiSYUlCjMUfzi+TvD
Nvu4CEJDIKxp0TaFULioOMKTAgi5Z/aB52rS3LeNsuKMny4Hu8rQUm/+lOSw231bIBqxSaZ+s/qQ
/CxXp3YFZF00rBayptQ4OEHhiJrhqNyBckHe3J5I9geB85ylot0gSkX0E+wQZJijjggFDjdnpAfJ
d+iHGhayI4pBRhlzuHR+VU87cL/AidedvkuL7UIjHyTnNOpGcwE9xulFX4+FZRgM45Ewk715FE4O
/SChVEeM7YEPo/sHUdO8Cj+cbWupLl62IsbTfDgCzj2+52K0uTOZzQGNQhELs5lQnpQ1ogmHZDPW
8ZWWkGXF8sA+EQ6E4l1TwtVl7y65jB/YIMI8B+y0UIJtOx7OfHkb+h/+RsFV0GmpzS8rJXl6hG1z
MHhfnFe/QwaQS/llanVRvr2FvxH/BBm3C6vb9Enj253xBQT27iHPFcgv0Npt7ys2kcjcL4sMAmhX
hMvmB24C+T2jX7y1+MCXF+xSjW8HhhrU//XwuGutIlQhXkSSDfDBKZYqH4Txn0Nxf3PNbj8EFuCb
+P5lrGOSlkSY8nmRI+jm0jDSyPnql/3/rJYcKQxWVwTDSjkCK4Nm6CJCpH4F9pgHSKA32IfCWjDl
uXQWguHxoN8pty+wNI/SmAdKQAeCDLokmrgad62Uh+wuWChTujxNQw2ZztEa9v4wZOuDH1jK8QrW
zgeubC+/SHHaBL4hesBEFrPu/Yid5j0TvL2pRL52z3MEUtnpTws14Esg69FnCAwjEoThvrQmexYd
y5l8OZBmsSJ1n1GeoJuE6amzbS28rGIniKBI2mi3i0/GgdgOdTQH0xDgta5TtXCSta+ccFK/2g3M
/xkD2XYG5IDmfchBxH1XZmmMb6+ouACiJ6OTIhjvHL5EmzmTHmDS1K7Ehd8NvqAsTygM+fVAxjX9
2u+zle0jqnxH2cTMtpX9W80kPP2ddJnvYAIRlxnQRJGOvdSJqToyeUC+CaLRnVyvjMn9ujD6HkSG
TITlZcoas369TFFdS8dyaoOs/fOKRFtQx67AYTQkF6v2aCv8It1WLqsDBpcmPh3rvnpNOLgTLh1E
4GCZACe10Z/Hpkor8x4qzzT7CnYHMD45S4DhXTTggNgSE8drHiqRCsKfOOIBG+D5QnVcmar3Kefh
Mm7XHs2M/iKd242Jl5LyHZ5Q8eEmXXeUjmLg4teXpq1ZPR4iY5WromrIgpGWcb3FJKpnHeBQsJci
9aijQKsn+k1UiIvHiqxAOkHeUjUQHBuExPpenpPCUiE4eTdyVxAmwWa0yGC3psqnZLFgjsxjl+Xp
Qdp7/azO7cGLgRXbO5anVX8D/QJUpz7PzpbYDLFQKP+jwfkvkViF6MrCuExg+6h78S1LLoLlErjO
7FoKsko3/UIK8hi9RN14nVgWAigosg0sWG7ugXMUW+quLGPMi4ily+mm/NSplaQZir9gGCbsaces
vj0u+Jc2yx4UokzsnFJzN4eXR5ip7rolVk2wuBrV7+lUC8Cg/+XKfw3SkEN3g+6LkqNRUMxWhxqQ
eSEZ9wfe6e95f+lwurrT5ixHu4U1H4sYqkwdw6qrhq4PYhG7MNhfbdzNVCuJWJvijudRNE98WSYT
VAAAD4TdTLloOd0KauIuiI7vg4mXVzKeI2cCvIpEr7VAcdHJphCCCZRKxkWQTfPyczxOBl86nOD4
90gT/5FVSW2CvteAevaXOkbQomFaTNlDmaCLXLPX5djzqXOQA77kqRpFYx9XTNKMHvKTcahEsQfR
Zy78mxe0+pvB/bqWWn4+DwvKBx3F7EXK43upL+JGHC2CgFz6y4Wwa14boxs7P4HML7VGhzK5j/a0
8+dZweBhAnKtFPJ3mwJf50QRV8xNaOdZ931W7tj43Os6U6F4WPq0yZhSRLbpUF1oztx+rllFSuZI
+UiKBzuo2HJlYv+mN5SyE0rJFxj80PWZ3CDX5VxR6Fu2abB/g04eCcMBTyLLqyAdg0hb2ODX6wPM
eYnpLxarMuRF5uSylcUvM4Qx33JKZOg81nzMnteED7ViVXLeswR/VPhLkPVLz+Hp1y3RIrlkR61I
POcM1wVU+Akrnmcg7zpwsrpvZxA/J27pelK8L2PFCBxcFi3mUnqWgF9PS/sRvlW+X2YNe0WRj/+t
gKkYMbbLqbIpcDAmggRYdBw6wZ2kNJR9TQ9cjY/PewB09szP8D8QNOQLTfGKGjuqy9KGiJTfCKCc
0DnYBr78rlJRntwDDCNCzqYVC5GfScwX0is7TBdQRdDhLVF4R/ZmuCyrWjqWQhlukkaxJpjENqgG
7HoSUq2jmUNIc2RHUW6A8uIbV4FTWHZQwjkgkRhZ1h96hYy58Sk6axjssXlXXX+NarDPd4A3fq8M
d+Pl03Z+xgC7acEv97lgaW6wQYy5Ud9CKCa4SndbAysYVn9NPghQjZZNV0eNPwjgg+NeEpveF9E4
7hHz+DOqmSENXtYYtDn3hmf7W/J/nhE5TNyphOO18vU3e8AHTr4Yk9Giu8e/sDeArbyoBJqGgKAo
xhs7wIhDNjMIAY/6ZFwUB2TKjqf65sGLKqf7oaWX47G1AXL7SUPhOx2JATtuAlPbEQ+dV3+jbZy/
XoXxatVsGLsAfzonEtCh1Z2Sazz8jbWQ0csYg4YfgVIic65OPm7p2/8+N2xhXD0ghJlNcETeTgbW
GdPOrQ+w522xb40/dl7mtES4ENRV+s4cGIqdElts20aCooGFgUYoyLXBvrYvo2m1x0kGueEGJL8j
Ammzd2XM9U4SGPjLstx7WMHeWZgJP1adyJY0hOmfZwrUBzTRp/mBYhrKX66qREyKYJecyrQLgPfK
6/c53tFpHJh0E6N1gferNLYjSQRZFkMjr0azLOZsZwoesVuOjXM5m+UKzzY6df6rU/UHSC4URlD1
Bp1lqvpWUJTET+4F7myR/QwGoqeF8w9gXF4tWvkA0Xm7RN1IjCB0ZBr46G6YiEcijgn+eGvJWQrJ
tKbwpvlCGtsxcdBCsYjuHebX9W2tk4+thopEi+ne3Ogbz4kzpJ+mX15WGWxHOIk76AY9S8KDAwl+
/Q4yY3IwISN7ombstNhpn0N/XHzZM0Php7MCp6BHApI597C70RL2+IuJqB0urRjTI2aDSyjJhlqW
ZFld36cThtNIdqn1EXmaU8qJgw+03wkFUrrmJvM7AqX8r/q1zuHEfB/LS7ePmN8JtPnqSbmOQ5M/
5IsNj0XJeQDfpRnIy3ykpsp0NBpZZqXEl+FONywRBnwsSS213ZObGHb6X3hEjm05ucgfQ+6UfOSV
O30N7Q3wrYkL7OMGXMEL16jXzDq/zSGrqeNEcLYA2XuHBuJoM1S5f8+KYpEfHsM1Qy5mD4wWnM0r
IKmT09ltMzOvQGqaGoFOOz0xqn9b//a/AaTbpYso9DkBZWFcu47OPyYv7xHoBOArvB8JFHYYth9T
lxHCaezLTN4B6Usz2CV3H9UxJIkxZUsUz2Jufzv1o5bopaeI23GImDVkQHIE2xMbWR6j8MxZMk9W
f6O3r0YZ2kBEagL14L1sfgH5VToAkAsuHaxlNrfgYbooprZ0aCOhvjtaUyG382w/6Hooq5+b3xqv
ntzw8miSuNyIofavfANk9ypqJrko64jenEl9RKRnW/CTRtGLcXablR6FN1rfDgxp6c1yPBE6jIJs
blfYGITltX07cIIOMxEdbrC/4Hv2U3dvfY5eju1aIuoMw8iHOU4bl9kE8butUj8Tdn3BFYSpfw1l
kSDXVc68GCnR5TbPZeH8r9ZoJjmoUONaQvspq7X5yM1gcequzOYXB3wEOEhWtkbGGtIrhX44209e
hhxggqyZfyaZTVt2OdXCWmHLIw6FmSgS99LZm87JrtHXP7c/6CZzg6vAEgIbVtMRgOuuXBsfARXI
iQbHjgYys8kgnrEWbmkJcQNEWv9Sf9xdWtIWzBU0bhkadELeD+OyEYtDXbWWkp8m1HjBLI1+zPTT
v45QLQQE5fUjaAyNLCW6br2G4jW/tamCSlCXRJZ1zMSozDkyX1JZrBN6fQm9TIw0F/IQm5S/wU8e
vXOE7kQHgA5G4U46ptr/G2bnMxmwE7bH5RcUHUFx8f/tr9qTuQFMxBou1fuklAlmLUJRy/EAnGUB
lHDpy7U5SorssN8yJDwSXHFqV5uyndt/1tlCJ6i6DKBlrYPJ9kzD+zFkZ9lWGWG2M2dJ6EvFti1n
MWeY8B3RpQkEM2wQhzcCV63MJwZcr0erddGckeFRppd1vo5vz4jxjtin0ELoV+MQd1SIS1/ej1LB
1hqoYAIPb7bPka1BcaBBO6FEysOv/2PDLASzTzglNY1NESL4MmIKWqyD1lpYli9LPnE+QG9neD52
j0DihTbE4XcuhfImCynOENnlKT5QnVwB27dyuTbt1Z6wj+qAbT1mbcNAdbB2lpWI0gx2biE/lLhg
s8LMCqKtZ7TZQohn8HrjMaERI/FA4s3gu7p/4VBfubUTAukkliHr7jBtLOJYKk1c1W4GBTjLMgpp
eeqhx1z5vY1Db04ML8eRekF7b+BG+h6+L78TKSiIuL6wz1HywCe6L6Gwiozg33DWthoeTGuCBgyx
k7eNCQLErQzM6V3TV8vLuPcI610av/6r8Ohqw405r4aLQZJfEmEMtQ7qWg2gN8DrtueBX8RGwFw+
QYvKu1fFX3fIkOt0emvYjkSVDJXmMbi8Q1qhD6sEYCEhjuDbVizwJBrB5UnzVUiGoMKrg6BfVzOG
BY9sQ+Nb8nPDRMDNfGTZ+t/oOyPMbNoXFg0ScTxQ/HwVV1xlYebagQxKNTOQOAmMaFhMIDU03jmq
KwXQM45sfgyf8sGvcSynwt6s+IPvQz8ib6QTNAskME3mVBV0YP9Hk7oTamwd0hyhPOwnq9PsgVR3
COm02J4YL/e7QPN5CMz/3u0J+Y+Dh6cWppUCYVfeAzXPU1Im2AORB2UF2CblLa3hvkCxMVeCeRd2
FeDyJgH8cpYVUwih5LJm3jHDCBOK/5FYlRiZ/B1zO3U4Ov8LK4EOQHtpYcyj88U4Ewd7Y1xykaDL
t7cbShOAt053w4g5M4d1RDO8s6ptxMrO56GlqB0P8Tmmol3dbjgWTFm+tlm9tMT/LathhbA3PFe8
5HjZVzj3iamJWS92Xu13Yv40G4kLTM0R+LUHFHvHnk4OwnPPrMoN4IjF8ucZ/KuUaRM45OLy2jSW
RWqeJDVz46rnh5ROnOkHc/y/aDQF/XpZj3V0JiKhj0gEc4dAx2LscGqThVQJAAsMphn2yZNnD8XK
B1xaaiJ+EsmYlaO26E3/xk022frKfAJSapnpoEbwivGNT4ANnXkUcbpBi3o+zI3B3EBa0x/Uw31r
YbzZq8s2CoSiLvJLRlnHH0DT7ATz0wb5c0v1pqszp6ZClFrHZMWkOw31+BXrfw7D+KTDnipyO21L
nZUGS4yy9sFCQ4aapQfjmzweBmmfnXZllFQnYLnVggTbqJyHdeQ68Wui0op4JiEtk+QrXprD8y7O
XtiMPc9DZMvcR43SPbT5dyjU2iYAalSD3CLLaeUwFIKeHn8Z8MmMofY2BIJQs6M+N0TGmsJg8C/p
rsKC2EHDJDkEdGj7GHRCPoWWzjtRLcls67DiuMagtthrLQ4ADepfju6Rw0496Ra5XRvBLsP8T96l
uG5X/WUUGDZCVCoi5Aw8NgBRXIP/u0TZE2CA8zGrbhlyoDcJWshlePK9BIyfeV+E0KWlJ8tBFx5/
Dq+TgNAoOEIZS+NKgUEPNGnD1A/KLwVBDG8xe38GfYcaJQjuLMXMjtk84dugf12QmFF5yViBEnyl
HyjzvoiKq6ZxyGhRdivNnJIzylqSCwJoT52HS5/iSKtlJs59Y6JSRduU6Nsv1vVGhtGMwL7TTn8B
eROD6YPSO6iC9fR2rXV7vBSbqcK9KChamexuM1q7VLo3nMY0tD34r7+pvPV5WLVSvefQCAFS7Zse
iuzNh8iff/hLT/qRmUtYQIO1GIu2Vj08BPaibRI5QDtmhP1YoDjGWUXNwTCi7RnDrB9P/ki9lVm6
pq2GUJ3XrEOiCgzdfuJj3O5p93L9qVUKhNntvRF6fQ7VjVwp7FLqZnhRbW/yG/yz72V7J+YqTvju
GHmemq8KThuU/4EratCBNUfY4pbpthjG3Lp/0p4jugDLl96BYg1Df/ar7Jxx8OZNPPEILwhy1ON/
OnP14I8cP4LlIxy0/r9MxufXBFXcyCOwN0JBHbFU0DsHm5wLvNwjSv9nVC8klpv4vzlMyu4+Mr4I
E+wtfEFVHL8bn1/lsv2l0LIdNY14wrjyz51K5p2R0k2+Iokjpll6gO64KWsgCIiM+uMkst0kJRad
yh8g4hZgeSa9J3g+iBr1cgD+Z14xubPCtfV5vT+ANStj+gijGs16a1RZlMnGGs73e7sFAJCrzsIv
sKpWcEgA1ug6d6bXWXYpWlO4TFzWpwBfQWhZyp87eH3SFeC3Yw+QQA9w0ITmuHRSIpwY4rS7XbIu
2/KH3UQCIWRt7XHTiEDQBcAeH5vv4vRjXjLX0FbIpJEB86s7G5DOcqlOw5sjgU7tyCUV27Hhk+BU
syNX3uPYE554iGp4uhJqsvz6yNlYyjQPBtBdCdJ8scKz7JGUCYNDycHbmJAhnf6n6/Fzp23TBeUO
J21gb2Uy7jMNYhsYWqAgIS9TJl19ROOB5DnTQuobaAspoIMqgTYfHnrshqrt13u7bqBh7hRjKJTI
PbNsJsdQ0oXH/bSXa8y5nBHAPz1wS5E3Efu2qdnHTg0q9xAuA/Z0a6EIEvZqXhjHzT8gAsUb2u1e
LjoE2XSyn41+ZA34NKaGQOkVtLVY9qxiEUYLa6uR/R8MAc+k8OVlLkbH7qCNJQSy1EdHOuQyscsp
AsS8roe5nnpGBS1pTlPyAFXB1OTxtWX3JB734+dAfp64ljUVKBIx9SKPxqN7W7RVhQ1Gn8TT3V6h
RMTsgkyfZFnyz/FHS59U06m8f3zK9UYz/BbFJIu05IBcfS+YeilYkSvgBmUPq8cDHWmdD5tJOL/+
byhz4nqyy1ipl+kIqdEU4L8gd8mAlVMj12L8rj19iTRNDggUm97xxzYnB4k8MEcdJ9//hx194f0B
EBfwDNWVV1n26I4iF5jaonz5hlWTsMO2T22arrux4hp7lz/iXy2+NMvdikUNlDTid9LqQuaO9CxK
iqV2uRr3bsko/cCQ7kkvj6MoA4FXLyi5diGCOJyq6kyXRPzePwtHnTOfyiDHVzQ55ONAs2lkQCEc
5l3iQzzljqN6YWya3sTQ6g3ESUd6bacgSPEYcmiTy2qHdF/CL6XR3PuR8sfND1TwKqzJX0e3SoLk
9A2qrd6L8nmcIm7dM5ZBgBQW5gBHHHsc33jBZX8w1vLtC4AOmoVVhxWi6VEWLl43WEq2jyApAdGR
8tGyScoaZfKs+b1dnJPbzunELYVE+gFXR+MRzas1dxuJOwl8SFe2qnyeHTquBO0JrOoxa1Vh05MC
0KP0fXzvMNQMm0eYC/8bOVilT/fYBrM94tDNic7qKB2S8wT6pZ9xjCc8u4Nzx151+E0gXXEYlRJl
h5oAsCHmWvVQv/RgPqORP462bGWz8Y0kDgQWs+8jrmz0oMXZG+fcNfoqgJoBAyjlXRt90ZNn0CnH
ePKi6k1QlgZhqeqneHaYr0UYt6mGzYepr4ohAWnDjrY43hKsxJWX1cvvlIcM+rJXlUNWT1BfYRg4
xNnB31nSukoI0zD3AGxzApihusTJQfABf4TMF3cB3K9mJbCaU26uRSnChh60iJP5bLeTne+fI0gM
GUXbHpNAQN0F+yIEWGnWR9LoawKWbIuAQ/TWzaIE/3S7pYwuhLxfvzPMMR5QdrJYk8NZgeG2vuT1
iZGZWYpdJLZIUJpnfnn4BhJj1mytQY8fjMGeY8lOtsEmD25cBZfbIOJLXxBmxt1fFIz0rjilb6cE
OKzc4bF0rcbfmXdOYqaGgvIFFIhy8QngEddkM8igrhEEt3IIx/yFKQKKiYms8q/U5DulZNDbVbse
nNp7ExLEYO7AXFGmOO45XhRP0k5Z0rNc7pto5QlN33WUwofp27dGSFE6VTTeJPsU+W2PWDI539Y1
e3kjMaAPUmkFyKqi0/uUt//3XiBha9YfkY3tg8fzr0oIIcA58MHUC3b7/nhhINkWtAdPS55BkUU6
7KBsaAJormlaB3jLji92S7VpVkt6WclACClDE1YvP5WmkFpGu2Ixj9ybGBMT9mnj/qWw4ya++0SC
U6H4bHXkzpweCv73h3U1v12F7p+8JOktXg0y2uZENKKmb3AHxiycENYUGfTJET164UkwoItojDsA
ka+rFgC+O4H1BYpP1qsXP4qYantGuxQygs8keN+ZThJrT4LvM8kigQyX/dL1LSXCG5YaEV5GuYGR
eqxzO0xyG871JVSqcRxSr45JKyFiDHokf6C4jRZjEK2i9vqLaWpw+oAgbgjj7ZWvJkN3RUByKyBs
niDw5h6sCIx/t8Ttlce1JC/G+E2ZD9qkOmE7LxryJtPmUXjW3Hc/KobyKqEQQ+nDR0zvlApHEOGw
LQ/H7duFyJ3906RVDeMzwBoM6CvW5A6fH19L8m3pwh4DBSvem7/vsi9XrixedJh5JOVE2jY+C7ZY
/Nr9RFBDPuWGtpNQPLHcM8BekF9X4X/EFIiOP12tgfx/JDiZQqcU8LwtNYcFsYRygw4SQh5e9N4u
z/LSvL3q4gIFbLDOO8AoLU0QnfGfFTuBTnqgTLs/p1D9ZHbVZ5w2b4YKwMTFj/lsknz/Hgq/K9BP
x6g3CU2TIHn4GW4H++/6nvbROR+4DDzUYJEfsDrthLnCjs60mBeq87zKNM9xkf91xENd4mlFDj/i
ICwpxHNwwJ4MuSY8Sjrxjb5uHkoYEL23+X1Q3Ftv+HVVIs7IsXuy2b4mUsNooMJoBOrQpJudXK9p
F3Xglfgpm+daTt5jukxKE9dDHO42cxI1uTO7VYuIJyI2/yHF7EdxMwo7sPAyqy8sfIaSRbXqG66m
HQt76r/p2p+0MmtzHSUnJQ4bx/hgPK518TQcCbVxw4T8fMnXVIjE6JDx0xEdYSCCVZphJ7kMcBb1
ApXXktpx2WsjNcEyE3urZG8O1kwrfESooWy8pjtYHMM+e9v9aFanH1gzUYxnhdqoLc3KMI5Za04m
KAHtoByWCVhLWkZqsx9xzOh4XwLnJlLtuj6Ih/P4eIvHwf3VTrQ1IHD7GFaOXtBYNh/609MQMusq
KMkRZBiZVQmZp1xt+btn1EOUEnRYZJiq2TuIn+RMf5n9pxCVAScuTyizyRAZjcGkCKPEUve8sDSy
wfiqUyD31RrTDDbpsvBHheQblqG4HohiDjeUOhm8qYbVNMHiYzhkvZLbrtBfOG2vkEJRLNZ/I9Qt
4yuqYFtLZoCQoVj+PXsnUehBCVy9/rCDYffqw62dY8ygPU1lbcyJZDuJoqGohOFc3B3WQkdJlLuw
WwOds6HzbGoYSugaj6K4BziFhzA0WxDR9pB4MpK52sTASrqV9zDXJvA7nPLoPhSscJOQUiGKzWeU
X3NWGuojadufKRWZvs0khEbxb6RYeRSuG2YOthGDeyiK5sM1zCs5Ad0xOGK5Obwm2I0VZiToN+Tv
Acxh3ncSbAypsZzEdip94ZcSmBdnyI5ynccqpu5ZvJbD2fAJJFLyaabR5fdkHpftqckmSNHHlMfv
QMo+a3dM5qevmNLhwu3UlpKimzoG5GQxApSLm6kFc8ANNGqdihWVBZRwVM+YfjQj/ZtKfYo/0Mr3
D8Eb+VyyVrX9HSD0iUY363T3+akeJsI82x6RaFXFKYCdI/mS7/0lPuGmqI9EALygytLSf/TmoOTc
CB28WqeEKb1/NEiadVXxkXZfPWiOq+smlINvZ4Y2urtsR2GP3Rwe9r483/B3NJILii9WpR702LAN
jcQfc6AHuJHKGSpqULNOZGALBAc29PGWssxJ9zVo+P23Li+5dWtgIReyeaginhMuk88AoJPZVz0z
kjxEpyZqY6V9vOcl23JVQNHeJaPJNkSTmygfulD7aTv2I+zFatG5leU2zb2ZIdmOg9xO8sE6RkMy
G4wIxfTDmp36kznQvj/Bu3ZRFNHMbVskh4eY3ziZU3oZ655UTCkMDhk+6MUPDsxMRPsyMs79ZNb5
fHcki0isGDGBanBX+ZaXDGzIWsQA1WKuQPboRoOaVDnwo75Yx+DBwtluD873bOAEp03p1PGoNmdk
YKfVoOXLfXAHL00rjaRB4FRu+ouzZ3I2UUD8BsIQlRsneY0xkMWmFFS3TfwDJb1V1FyJfodOut8M
ogSBUuAvXhX1ru0rX0x0+euvCKTQHOjA1iC0qAAk77j4jbRJkOioBjHwLGTbwo7vSKo6XBHHGLoG
YuMH7TSEx8f7taKdBmUHUJLax6NfXJm4/rXIHkJi/bbSQ4ZoPZr3QKITMbBK9aK88XTjLWDSjYgX
2aWWvsAZwYAucAmPWu2dgplTqOMZCvJ2KtM6KrAco2zf8Xgnetfj8hpBa/F6g1E6FpN+RB3g24bk
jQ9bqCf4QIyg/agZm+TPFPEY3LLoNioJ69z0a9dcXvOJVgeIakbWFMTRRjCwemUGQ9fGhvvTPoZ0
9yB0iqr6DZaYEE85duDnBGSpDNxAIOwbzbXvpOaFaM+YolGCgf1MRmxFSy1lUrC8X4pHiAKT9pna
E1LfDEf98Qmp2jADr0bU9xonL26EBjnCjhN7sh4frWB9WApEjmTrhIe2pz8nqmiL11wdynAa0pLY
xhu8a12LivS//HoqEDqlqp6JNGlZqzF47QrgOmTkj0vcqaLZhIpjCyfFlv0XwMjSgNK6/MQ50LVS
vKEvSoYAqP3E2e6Yn338Do52S7TKqM5DnEZ8oyPA/pbOIAj3I4BIO8pUvSNrD3gfdyUzJN4pbbOo
1HLDfpZFB/pmi5iF8yclWeVVbcpHf8pJN3u2iecf+u6sTY2gpa+pie13TWgTmKVgtn9NvsTSDRAw
xlqIj2lscnovROQK/ObI5NbUn4NQtzH2ApHEHYtrSqHN9W+HuoZF9N7NNNTGP79FjUVOV7In/bkD
6Ta/ZOmRyPWGylr5qOAS6I1z9XiQEcueffY/sYDiRpTDzi36MCBc7yPBM0Jl65Tv4MaCKHApJf4W
aJEoxydgFOuz6kZT9hUL2aBviDBsP5ADOdTLdf8nDwBk2aPziuynkp+C3UqQXr1pzl2qj4u5LxvB
Kiw+6+g3OCuaL7pkmXonDkqigAROTPKtZj2X4vBfSnk6OQsfYmi3qK4DK2GihxAiHjVyAxOtO/VT
awzaBSZlTVFH31huCbaY+Ebs2QUUIjzZd2/CwHiR2etpdqhOt5SsgpfuzQasFEzwtWxBXjOZfAcZ
Zmpf6D6oZvKhqdc+87Dtfy0NxFie2EW1pBv2Tf4h8pu4+Jj8tXOiACnhL3409LUMDDkKT7uzsDGt
eih8tZmONGU1cWhYkteDv/zYFW4ekUA4aOYSwqe7CGlCEnDVrWeZGW0TPTroj4YnKXwT9Vfow+vG
YVxUIfUcgAE6NFfmRtZ4BSzYRyEuLvBLcjgymJODUe898AUb14CpSOzk6GXuIGXJb1loF1lZum+1
KLsBt0xveWOWmo4Pk76u/kVgy5eko7XPsxsR20cNm7/yROGcBdsbY/QaHLvwFJbJVuhwSHdDiKZZ
/GCyKFRoyuOU1lVdNGnUE6QwZhsgFI4uMvbi+QjXU0mYJIlZNY1HqLrcHdmkNISHyd6XwH457IRo
ndkk8grGgZ4cAGq59+CwN5jVeoIj+4Cul5b61wxrbwWU9QhEBCGVQ5FJvg/5cN5QZwTI6WXM3LVt
GC2bY9zjAxwMxSdSgW9UaFN0cRrXYz+p6iw1OPTJQaFdltmpPWm4NUU7xnuEjV218YmoJDb/xtA9
04buc5Q0bHQ3k35AX77yQFp8CoAPN0z71MgALLoOSBuVYV5dH/+r120PjOwKP53pUVJtU8Mqlk1G
O8sVt3gY39GMD/RMOywmMDFA76KMdArmDQcwigTfzjL9KvRhONQIhHMk7bvW2qD4b7GXKlQS7s2x
Za93fNC0mu5cyvQQsO+pZ6m7NKrgZxQRN6gUYJVzyLi3+7ZWxGVEHcqivJDAZbOZmAprG/xFZ+wC
dB30VVtF0k7LIAyGWZ6J5zFSTzQ5D3huq3VqpCUkH9v+EX8IeqLczV6rZcLwbX3OfUrdfEHJ6M/J
NWEMLDfmbYiGjZQsBJZn3a2WcHWC3Bce+tZlxmSF787roaF52F2gnJtO58Clh0CrRQG0qx3Z/a9j
k9yGd3t/QcL/BPqKq7LzSfqz4mKephLcN6r2hDh3gl3CdnC1Jx1KBJkKcfBQFia2265IKMrQyJX+
Tdl1fH/ibtJaRhnmW8juaHpQLX/oirS8FYiZcE4/HIDUse7oZPtYylBWTXEOKAMldW6GfxntNPVg
hSZNsb82zuDPSWlcoy563Yc6T3bmwtHiLBGD+66DFbjPgcYBaiZmHCPtsZ6suSOLhnzKGFTDdclm
TE9/3f/yKxEHzzvusxm8rqBaAiS7LWG84OO+OvvcA4EMVKQHuBWgJjJUtT545p6iWJmO4ANJ16L9
/wLq7BdHtBK6/eo3NmWUqRhbvaLqYnB6fBlvITuUgguJCZjBE+5lxmxydTuBOz5w/3j3g7//W0QL
FdHGQKn8xLZErtsQoz9jonFY4HvHfWxmissh0CjPcVUZ4xG9w+Unsd/SVcM8TT1ddrpAA1NY6VM1
kR8t/4fZnCDNvpMVdRDxBnUh0cc5eiBSmKXlkfBk44yBu0oy/zcXgNfjqVS/vMpoF7jmUfUv9mZT
ktg0y4F2dAfSBBQaQRSHqaXK+IHgAWs0SPzx9YNvkdOcQJNkt8k1AHTr2Yeo2ihzlp8imLNd8jV5
H4j9vGVqPwRFbAquk3aLq15cLLSd7aaDpFvL9UEw4HaZnY50TGjPRBzoV9+U/OgK7D7KxTWW9ebE
3FFlqlVm0M5i8pgzhkrwCd7ojxI8pBixMNmpHiZeQk8N/DMonwjcE039G2XAS1BA0++JEoNMHML8
YyT5vGybSA9IO5+7wV24+soyR1XSewLegVbtWq/Bn+mhMGAUR0vnDVAGQE6h2/iia4TFScRyHSCl
5K/vQKUM5lj7R1vOO42Koyb2xcF2ZBcrAGcz/NDr4v6g9yF2Zlh2jRxwX+Zp1oWJmz6N3bOBuknY
yNcWAJwqdBYGTXDRJhGmNuYzQlVH0eKnZOCwsKAqb4kOMhjRq5JChxeD7bjzXe8UamEB9rnTGjT6
6QyCTPdLXnktSdaLAVgckjQXeuWfaeoUaMhAgb5GYYaVbhP3RlBMf6ov/HMSGOlG4+sS0cp8CF6V
cTwcNCyp75rGA9Dp5BFZy9fod9i3rmwku0fjhWG1pMai+nha/zK/vnpxaRaAIP7CtBiAiXR1RExS
bWYxpaT+RReyXCYMpoVwIymF//I6HeR1I8fyraC7bUo9S2y5SR1FuoZ/KA+W+CDZfxd24iQ8YJbo
2mpkodNRfsyB2TDRfWLALrQjF7Gdz4DOnoJ18wuHkAEd2HKFewcfwy20KbYEVwlrdUULvmghvDbx
QtsyfNeqO+21CZDvKehBGEldm/anr4cUUyVOlpgGoi0yUqU8VohiGF0OSTXrFBG+L5EI5KXUSAt1
rCnxS7vMvcCxZ9wE8wcLOylaaNAphulzElZBwOhcALA7vSH5eymmBKa0pL1lY9eqG0i7/NnJInNK
kieyi0/x0pfJ7/1LiFiTpbqJCkERWcnN8KhafAz37jBRNS5bRa04C33nJG8cy0tKkppUTSBrJadv
nMjAIePp8wxaShU5EcR7cUkjsvvxqJbNz9tVE1qNM3SGEGpWoTgyy7q0UFJQQYYNumy7ornlxRdo
+zYwW5EaxCRpb+L2qLkGtKS9X87hmg/iDXL7+hp9tTYPbdpUzj32cEavZhtWNDvm+CJ0pSt+1waf
4f/dw03GmBpWYY+G9EQUodFtVEP/c7EYfBJMPTtlqQIdeHS+EDyNmuSn+9/a5aVQMA4t9z5e6Hid
wIwLafR4+wZ/8Hav06N6xxezaxeMvMn7FZI9vz+1LXwa3F6Rl2EHG/HvxTSx62pZ7m+g7oej4fMX
YNxqEqsuxGvGk04PRyLz9QsBifOHv/+/kp3w/HUx8T+BqqzPgFM5NgbcwnGeFcYBs+ZZUSbbS/Rl
BNths+piMLGoaajd/UAob+IlucVPRVY7bydyQbQN81fbK+7GEcS7ZzooxsRcR6Z+opyxJg2U97wA
G9HIZowzFN7yt3WgBxAcM+z3smn+hWKb6JVS8fnLnDtrB6ZFRkeKtCGAmQxquC81pCCF0YEPB7jK
ikIX+U6BQuYLsoNHSMCZPD2Ab/IAL/OLqO+d7B7bv/CuBju2Lpkv6Ucq9NKPsDbskEdp6eGPW2t7
osGrZWt7G5Vl4Zm1E7rdn4Aws5QQ6C0umubbRhmGPPiueSXWqu3eS4tz6baozTbW8cDfqBQQjido
oS3wAUqBVdmEG7p9VAkZpZhMH/i1P+ojuOV1XrwMAldchLaHINwOOWygxtdAidyqgMRnq/vwGssY
cKNwxKQLu6bWwCh9cgL5iqWX9TodktgrlP5YcyEFoKNM2ow7Rp2TzvCLxnH1E8MrVCQFgLtQup6Z
MulFQlPaO0O9DYo0zcBDU+QX7LJoPAskJ6Kc/3IUueEcrDVofOvP6svZDQp+G8wa0OlYD15NwyEP
Fk/m3nCYdjolpH+uVEQmjDACiRUnD2EyhTUVWgKLIxIpla7nJj2myJAohoF/66dO1opL6f+EpvE8
tw5ZYn3DizjSdmQBhCeqLTwnM9/5PA8Ze43eM3T+WtFEDLOBT9FJ3r8SOViT44v3HKfkmSoZn02F
49QuU3p/FmSRuUt3g4gc4MEbkgwhd6rWKQ9bfW24mkgij1DcY3Km/+It12aE7yAmJTQii+Yq/DJ+
C+WrzrQakM7Xc7cDHgnItnphOXHP7aN0sISeoPfE54AbY7ym3c74QEIPvh9x5MemJP5nJteKLIqc
XRBbD0pmd1ezuW0O6Z3xAtlDvH5oISljBiCVre448Y5R28lyalKkLfXyQQR2KTYWc9j3ez6JO/8k
T/vVp89OqvGyvs7i3C5U5AnHG+Qs6zCgEqULF6/dN2wyMQb8cUhrHO63gx2tA8uIdjjelmYre8SQ
GFWnRfIQE70jwTRAKKzKe6Hspcs079UEMPd2BqmZhoCHZrvTK0zIMzYrgA3phtp7VTfMkgToS/rv
T1Ip6TwD3B/vRETRE+UoyMncMXzQdj6pzBb9O2bdENzI7+aO9QJyvU4sXMtgtyjGvz7CTD1IAPal
+Jl32FlqRxxG3NOsDzIQjDgd4w6P/HkGOc7Z7kyLsiNtHIFiHgymTAflq2z7RCYG+Vqn+H1glPX5
OHMQ1YqDxetL2MCXHCcmKegKWvwGarJWIDvS7KzoAy2rOwSjFGNCr4z7kD45tw/xgLbIOBzLyuZn
9lsg8Ws8Hg9lDqDcExtveQDAMUzUV123YZ0Pnjxk/Lm0ANK83gLI0UYCry8Dv9gU+f/Uwg+pH2kn
K4hf2yjbqnXRzmisBIjxjfWMu7SAbsfBe39EsCNKQcLmHzH7Bv2HmerahpAyXbwLCjOx1nCQqxzY
YUsVyIKds+KvjFp9YcMqtANnyQz6AFxg9OtF8WqbKoSMaFe5twkjBlWdCuWBW7SNFTlY5puMiuOE
7+wxz3W3iyLHwrvkqlssdJXISzv/nR5ipB9Gd/iJRtiO2JV5OfOBKU5+2xSKFdIBi9zIFFwzytoQ
r/wfxp5kSW0OVanWPTsc8v1SJxZk//08YfKfRuD6xDTyeOkTf5psskrO8m4kjhdKIQw3jVtZVkBE
NywpxSUaE9cnqKO/VDcSfSyWfybqI+tv1hkEkUBNHasUcT34e5KFmJuXWGmRyIjZq9DAMSP/xb5o
e+txkqWH39EqBghzvJmjNFwRtKAg61v8gYwzA6ziTE3ghA2kAby1yKIjMF1/egOKxMqk2K+WwX/d
mcyOeJs1IYATLiTwIl+WMxjdfSX07gwSfhnWjnce9tp3MExxCkFvD4b+2sdh167LagQ/NRwkG4U3
mAKCD3iKAQ6Khmc23pRbsP3M2q5tlLfNvWk6xLsvt90quzP/5y7vW0TGoG87zXV8utcFxjJj9SYT
5n1491hVIEYwvsMxrUkd3YF2Ai64HOnbr7OVQVPWL9/1YbEa/5gqH3wKG1u8kaa+UA1GVKsy1rpg
oQ+t164LNUeqzrHxQNkxGxrPZ3wshAMZq0aANXgWrP4eSOGhz6neSZ/X5N8ZBuBhUieTvbCrFaU+
akXb/5nkA4mt9Tc5l3trDX+i1hLu1owqrsFnV2ehURURiFtfRdy8L/ZkOR5Zv8poIwEgYW5icwkQ
2F7w0mSXKp7QSbp+EYMjdMsL51VEE3xYd2VSQAne/S+TgbOozG+eHWQppzQLaYr4Bpf8BRaYCrIO
wpZoPrxEi/SbOQc02DWDVvJo0luwI/3Yxy8PazAnMnEzhVbbhURyLxaewZFckPduDGcZ8mZKeGA/
9LRuTMPBlGOyNBAGZe1fKL0uPiIrwPrVbACW0tDIN33bzd/kbxTrpl2DRYXHPpKCSk7bT1jJok1H
+TUOmIxyGGhbuB3+dX3gQjRIk8qaZtOMjpSFzg0wkRTLZzEpe5DqR5RCsHlpmjKN7hnH6RSlGIXs
Ifb9Vd6Vpk4UogF1YSG9ZX1px9Bkm9nBglYjFTbT4F/ZWy2EP3y50bbj0x6fWrbQE+jKoxCwtnyC
mWqlYAaCBmzNkVwJIGFVpsFtYhTadozCgXFTJ93R7EBBn/WMDV5kZ+0fb1XGxwq3Rx/phjrh7JAE
wS6D7+f/lWjFh1LkzeFPRVygG72vzN7QrkP57v1e6uUbNvAE5eCe5mWkb6uYM3hpITxyzP6AMvEP
sIlsm/ouNv0YaMu4i+LfgW7rnMDt0Lwt8Soa53fOjjeFaeQ7AqTh/yz198m+UgLNIaZJ8YgTXZcv
LplkPtmyKCqR4zOXIkSp2RJfVbzpQzXa3IrHYH34sqKNXLmNMNV1FAnuqTAnZgiIVMhSsiRtjG6G
vrm3Xh+Y4HIk01X2T0bJ8d7klfLkeN9ROHqA+urK9p8WdQm4jINBmyrWByc82ENoGfoSp5CcqqEi
g9UPzRH2xIlkVCziNWG1ijBJRoXmU6kJbEgf2f3D0x4QviKQ9HXkUQZIPp3XJOYjrN2N3wwBnp4P
DN+t32LKCBb/nXqLB8BBd1bz3/hOhsPG1fA+NXHMS71V2EHMzQL/3BX68B4t+2ijYhbV9e3KUFcg
DBk93u/IZpEV/D6QOmw2n95YAbbsb+zeVzXSSmXw1MSQQ87fpmCrOa4WufIO4YMAUoaFr9o54BP4
4fouIP2utSAmJcovFCg+dF3lX16IwnXH8crk7eZTHpAMs+fgJB72kdwzOUDGP5VPUqH7JL6W5BCm
Cm8nzKU/F9cL0P4pnWXmOZfHRfIz91smZ7HFCoX1gg+yk3PAfMbTy+1IHus75uaZiotGrYz2F3Y8
qdMg3DJyu5bLelvJPz4zWdvR2BZEJItYaxK4egxkZnr4/ZqtlIlbo4BwKwpv0zyXcd2XU6nIc5UJ
sn2hknOxkSQ4FXqZ7C0cSCPkutPp/tgeC8YGosoeBuxnJvfnpO1dYAsf+1EIw5UEncobg+ImL6sv
+PB75xVLFsrD/aKyfuUF6FVWUbBw7sCkRNOufvpdFhaiyGCt891ivECBfW7epPtENv1Mkhd4M2ku
4e72hL8MZv6/vwyUR6TFBJVW3TdmzMMi04j9DmypAM7jySbhtBgKPiOGAp1T/GUd2h+ym1q56cn7
N++IIhnJ6sFkaEQ/bztwvpOP+ts2L4h7G/KVQ6QLP/UuioPrYdIOV+MKlNd0FFCG3ZNCa+wD+2t3
Pte+E7HPu1HmNP/t/6CflvN9WUlZccQ2s8QstDd9XPztY34yK3iO5j2lCsgUKJHq0xei0CGpJ4Ab
j8eErgkFV17Il06VmUITQ6lzS3ESA+9QPgTT90A0sZuXV8vIUGOGqu29k0WADXdEBZ9Pn+3f7tvV
K3h6t0W1RHWVg1eZIokdHQZxTJpzhwSVA2Zy3y0mnW/hzYWAkkIbDn6AHtIw/19EePEmqbYYicWJ
KjkEj3z1fBWKI/Wx2FGHVg0ijXyOed62aUocQtrkQFx5bqzCugz9QMpUQnC2/uBXPnruGBb6ynC6
rpQyid4a0Rc9bLLihTjpKr68Qgue2Y4/dNWWyHooI0tG2UHYSXvrUws8chpSFvE/RNQyZfnG01tm
IurE5z2G8DIyyw03AKZVvsXZSchGCEwl18/7w4LxQ1YFwOzWwjOFgel78Sid2Bmq5JMmNwQJvBJ0
EFLzeo2L76EiPu9dybxkvhFnnz0p3GPYoTtdcv643xM6BuBvfTdy8KxEZLSqa/X4CQ4XP+44G149
CmTb+M6OHIv4xxSxVbSajEfFx/vpPyEtYFKfiSwo65usDwEoWKZoHPqqeOoTNty3vSUQyopYhnE1
9Ph6P/rFRZwYuQx/XD06FbnUU+UhxFqghGG369cP1K7PsZgvYf2HHS05Gp40k97WEZhLuKjih2af
2K6BgKkzwTeKDxcnWulxJTmp2gSVCkXxfUl8tqYhoNHccrWxy2VcLPVeJ9Uj3ekw2y+B5Q+NZIy3
3kaStfvhcKlRskJupTbQLdz+YF++/t/kWA6WlAD599ot10Cg6KpyKKR2+YzBG6iy5VeGewCsWdQw
Tr5zARHB1H3cEUABJ/TfK41FoA7GRLAtXQLoRUaWXMhW2iiamSAnHkdlXSrvB+cXc2TmgpoUcd5h
DJpTujUeZnr7MrTY19g2WZQt5QhZ5FXo9zo43R1T1e7xXN0foTGNJVrwXA83YrguzQjVkp8Xjnk2
5dtW/jrXJw3izonDafnPEuFXaoE6qWlm5rORFsYwoDtSNPg7SWPJC3CMZCH2zeoTkfXD7PzFCJsd
EwtfIEcCwsxsfIL8e1wzbKGcfRhpDQaiJFrB/M+X8MTmCwrol15ajOaX1LEil6hhvP7//CBIMu2f
RAwT+/2sViSL1r2TjkTiOVVRgOOaEuph2gFXMQw1VAUZmCR6dcPSL34egdmsbxAXRaAQ9Uq6mrUA
Iin1ZMRTDDctyzO+d26OkugRlOGMPo3EJnFNfTAY/dKhtgSf8Nt+66+oWnOKYrLsT0O9/2H3ihcc
+CbDgbb4XFjNxyxsQsae5jKWOM23dgDLKaVnn7sJ71PmeV3TFgYc6laHQh8t5NLWQwG1KA4Y4QLo
oynEUiWFJct95nIpUrCLsi1dZ51m/zDPZ94dCM26MI3XX3svIerm2rKCbVeig8eU7Z15MjQuhqxM
25Twwa7yHzuDkVBaUAgPozx4HQ1sNGzKGqqDGq2DU1DIrX7rCw634pJMtOBbEth43deXklxIUKla
lco3N7xtp1J8KpLiGLZvcEShJsF4mpZxa2t1N2dJd4x2bODPlsFjzffCojIrHYsVZnlfCGw5pz6B
rnW04H0mJ099nyxLTWYVG8SuTi6nFH6aWBD/vOT7njfdqKQYEwTngmPDZX1ExkmqYypjR4WeVLnK
btKWXfURdKZJUQ71P9oeu6VOkWuAacYOQYF+F3WGZlYftFElik+JnvUABzmrXhF7aL8YMJB/NLls
lXImgPFtlwamdJ7ZAFCyegnEF0po13bB5K1A/wKJQfYKAjazKe/vDnOx2CzE39aWUXpoAunLyAic
f4xf/RGyp5Ktd1bcB9VdO0p56GtuZ1Vq465NvcDPyWJavbnuD1JoZPTc+wvYYEk6SPq2VkOmWpyj
vARSj5fi/e74HkcDP5Pr4pTcbkDBBqsJOlnCpdWPO087Q82q5AO1d+0Ec4KJkcHE7CxxhVNgGN9B
AVHWZ0aa1uBR+tkdajaVWvL5lwMMiMh2ITtpIZ8Rt427DldgM+HoWRB2ZIeTNsBN4+nVCxSIsqiO
H6w5eUkTRFU71jOmL0AWyS7D7EsdI2zSCNPLato6XMViCN0TMxLfZ6KdFEYxok9xPffKxgiaWJHl
LIikgiFgp4XgCbscInKRCTsssGBVdFVFQ9M287nesE3wU8g8T4E5njSpZNXgAIKjpJ97xrzRp4Fe
jYC1UTuVK1RhvAcwdBDc6Jgx+5znGmm/gW3X/5BquZMbbTKpkzypBhjfvP0FlZTrsjA89Hfhpg9T
hvMOrxSD+uk5hEsniGJ+ihyCen0oI4ktZfLIBaK8uS5vTvc/3O4uKg0aYTSfkgQRD3qMbB4eu6yh
b11CckTdY3uQmXF4Tg67luedPH72/EvhTdfcG6p+R7GA1mdseUszy2j9MgWpI0BjvMzagl4wcFWN
2LHRf85tqjBHJIByjhAYtVnz3EDE2+y1bTNH1XTzsSVfMpfN/zffQXWZSkus+JyDVgA27xhOXC6F
eGPOcB1MZGoOIH+HTCe5TlPYb61+irfNFxYhhVCIryvTHQ9b5tXgSYPbGiJtnGXJUiJotpfDNdCR
OLl4heJandJ4I2BB3fi2j+8I38V1csYhG/QccHb7jGEBXSPxQqWJp6quy3wI+tpY4+FZiqm9loHf
002wFYxTF6mSfKhjl+BTTKu9GhfOo10xXi/Jrczkm0FLlNTBcQvOMlCFsu+utA4SRgmr/lGrfur3
P6pR5GhWwzYGLmcaT9zLeBOXwAwgjvXRaKmLw3GnFjsFLP9540Ew9nmjbZH+/b+E0a8O+KtHEpfm
Bf7TKu1R6YkL0YAeqI5fduusq6XMaNrr4ZXLCZSM88S4lxg5noxvG17oo+ykeUbCCHYQSSSepKQB
8OzEBNfELekOrVj1nHOzqrwZSWijBhtfuk5WRM9JmW91uN5JKCySwrsq+urI8i6BXqZKq8PMofox
pXAl5Z6IJEMB33Qm4ftUWUfc1v9HjpjyC/EMPm7VTd4W8R7vD7/6RDN2mhjxZmMM7keqmAAq6LWr
pEbCNDe79gk2wjHkXJ5d8pgjhsoxKf0CdWErKvTLgaHf8QJDu9nq5vUkVTQQix55LcDO48TI4ZvL
bBP5wXnPsIhn4i+DB5w5YHhOtOysGav1DUT/eBRIEnquN+MSsHJRrXWC7L4qYJ3NO5HX6hzqKRDJ
7puVnSVEcNxsYQTO9YSCv2o36rvSApJGTUx67PSAMyaKvPKTHkC+ezySfap/XbhekyAdeWc566KH
NMRxmu1VWlrIHVKZytl94q6xKgaNv9WQsOB/9mxfKl0aP4zEs5TDBA+Y4EqBJGhRQPfavnhxKdfc
B3hVICgrP0SBJ36Xl0wmJ6/nKkqiqkHHZOTQclNfvEOvSZTg4ouW5FMz6GfBwFlSXb6z2x2OVuOB
A3a2XFYlHAvwWe4D2pF4Hl9s/Grgs+D+OiC5UBp2RVYRuDd2nkZ18rq7pYXz6ETdtWzn3W9C690/
SbEhb719wlh4QR9LVfRo0OPla15K/nIdVp6rBcl9ZdUZSuTlIcjOHGybYdFA7pnHB6e84HG1J+0U
BS5T2ohR2ozIlHYcrKw4Fo2CE/Lwp4Z70F5dhN4CFNRISpK1vpLhtsbNL5r4HtoQj6NuHMMePW3e
tQv756otW98gYCt9jvXIq7w0/kSAXUkpSU6PK6MvkLpOsZosYV0a+8C58seqaWdKRdzt5wpOHCNH
VJcIlcP/tVE3DEmR9VIEHaqpFuki39kb2ODUOGrH6tFLaNgMUkX3GFseUwYG6r/4/Bc4g7hbcleF
O0QndvJLGBDWqOkkCZYrRhpxXP8CiUCdSkqYWSit3OeKUoNhjNKmlU+LQNowWbABcZCtCn6txyxn
+0r+v2zxzg/vVQ5xQT8X0cYdoEtk/j3qy2ynOqL89bUsk7DeOqYMHL69a6KgGRTWfUNWX+9lzPPm
41ohOA2FuR7tKSReAcUN3QLURo8TDCg0qKm+GAnqAjhtFPBSi7gQHn0p8m1ianslxnS5mNJYDPIQ
LCzJGXq/L+X272Rhu/YmAT122pT2vm8J0OOGRPLAnDAG1N8qRFgOu9evGvzxTltZjrxbn2KSCPWw
Gx4q6qcmxBpvnb41ZP8Qfvoq2ZZpStG9g+35MajHdzVAiQonYeVkvuI2FaDAt04ggRktPA/iN2xU
G2v8mbiU8jh2V0u8RSLspk9U7UL0ZoWPzVw8bbpEk/n/nyg9lITaSQIE/GeYed7l7w6lAqmPkikF
szqzm1TH/0bpPnvlqoxH7hqESL/jwl/mAfrdDAmfx86uWblNJ54lZOSX3YR4sjxGMMtSKuiUsbQj
gJqxVJspWp6ArrtmWCMHqxQ1YVmI7nzU49GUe47dIzodUXrItW+MGLsXSSCeOvfDK+t2TFn/cyvg
fOFxQMuPeFOaTFiFlIy6gW8clK74xC1KTu6KP/t1Nq3JFMiqPRDvhBDZuChhQpl846CMjq0z5DFX
EjUHBIkkSO9Rcf4bQTBK66GREDfhv3/rzHbxkn3U2wy3eTvdxo0lQrxiE+BuCPG1O37wJKj7FzOJ
7fNCvN1a+B3t0Yf0P/fGVNPZslxoZiR7hvgi5pYPQtqBmM6ksYk0g6VAjlJgY5n78Bx8BmbtCPtu
DlQe3Z9NswFNfFoyF/GZMmTS3garMFtDmJgpU5agakvh1QTCIp8rWAvMIUkD2CScHHidBcmuk5YM
ra6oUk/Eyxugc4ucRoNsVwteihKZ+jRkTmpR2hhqO5cI5wmGfFcZqq6gC0OWdxtJfKTXWARi/0KB
pYk7GZJ8TXIk5NeNIGrTGfnIEMqU9XAQcLP9/COKfDCpPTnXdCsQSgS0fn5UF9hh1qYkgdnajPjE
dQ+YAw8HM3CUH2NGhczxWG4k+mHgkyw0hbXTrPiYdIa7ivfe6NJBAA35qN72zXqT4mqYWYdy0bqE
ixX2GCt3bMzqT0eW7MtNGDFtQG9ZsOTDbsdVr3u1jiBOoPEDd3unt6CQKXClQY/mmTayBwBGd5hg
wUwE2vtu01blqmpUbUuEUIN7W0oDptoncPEiPq/C253bLunEboWzL6SSus5X31XBgFpzvB6yMC0r
ylggpdAW9QaPGlwzPe/wdUDxL/X2q86pFgP3dp0aUmxQo9m6SbwN9XdU8m0/9E1a/IZZ2Ups/1iC
7WVf6lQ0scp4s+9XIb105+58q0BhW1yEAPikNMd7OdguvgOHp4kud9ylq4RLqO6jaPd4NEUoJOR/
1EaPauvsZllUB4bk35v2z1itLVhZKM4m2vdloPZvSFfv6q8vyOxi37RGTmDMAg3YZmwMOJeREq2x
BnhfhnvsjtbxkbMzpdxBisImjAez1DCFZThPwitf8nwXuYpOzoBl4f6xAkMKfXxnkStLHEavGCs/
ryAqOgxijs7YcOW6ZedE7cBnOjTaq6b46ZB4cifvBJdaQVHjcpCCErZK3szrd3Ez0ezogfmqBTNV
ES6dQlilP5fL6veInD7gWt+Nvk4/bZs1P9l+GcKrZ1Pzsa0TKQNsn2e9/yId1ETmz2nwN+tavT8S
AD8dhAkDfaLVa+V7bLTbNMp5gv84xfbNLpiKCjKXiLvJbS3DH3vC7WvR7uaYvPpdZ5KW0cfUFypa
UYuQJUuRZj211M6VvfNyC7WmjUTb546LDCVXOCOtsZ+K4ivWLMvxEiPo1n7oJo+YNqa3ic49Trlz
A135yz8xbVEFEHjZbbay3J3mIfWPKIYIF2PwB9irq1L8HgquXb74YMAkAIaX2zeo1VBCorF7uJ4s
PwLVkIeKAGuA9+aX+gBASGCbSyV1Rxs3xD4MlqP1jJjVP0/LZMLPfBYL7A8BQKuzOmG2yZ3bdDY1
nFoxyFrJhnNdpX5sC0P6EgEVlBFSar0bB0o6zkAsMLiqUXABkumwRq6pwzv4ovu91lPx8XPWUzIr
v6AQgA1Q/8F2iscfeodQ991I/legw8FdkulviLQFobcNA9pi4PdDM4pBGU2oXEEg8/uwzavFH6Me
CAh6+oiV5U+c66xk/2yyLGREUlZ6w21KPXy+7BA8x42mroHhLcRGSwpo8XoBEUX1K5xUNAYRFKq8
mJYb3tX/XpOILXXqlIB5iUdKPknkwo+3uEEkG+wsOSUPyaQaCHXlZm8R9Fqa372+dU9TrBw1n0h8
BU5uA/4xK8izpXyTtbW8CsMEdmmuDReWZPBd/OtqvrET4+ss8UZD0jmHejTx18RYGYY2Nq5VDjRG
sLqlkOZyANRyk6K1jRcEh66t5IYMylHPN/yZZCrII9Jqf6VIeMGPHGN5USkTwrbOJ9fbdXxh3+Hn
hfhK+4ew5H2FlLSc5GvVT7/sqlp4nxQKpZEQ5yNcgFlwjae1c+MsJ8Hv/atEMRKer49GF9w7+o7w
yZ4XV7BmkhhQKucVHxr7WQqNQCiMTi4x7+ZpeaHDnUfMq28Q+9Jc6g2muZlBBkLrw8JY/eCKqH5Z
6uTIkfHZcMxTvMlXJWX7ieHAGu7YzkRxbE7iJC5bHvcNdvt76BX0Oy0YNsX7BUZ4//4fKf3ei089
1rDr+JiAUBGuE1wvH4KO+t57/TMtSO5HzCgFCr9j8OxERPUXGiWoV2J/7KOG/kIAN4i/0Gld9G4y
CyUXtswCq3fC+/+saFiT/ys6q1oJuMsutxpbtWsTK450aBIQ5BLBG9c3QeW/JBm+edcnd+DH4CWh
IRl9F1UOOpYiBcGMGbYRDzYZPBKy8BJBxaeO2Ws6ABCaN24ueXBUcqW3eZfYm7fewvegl0f9I3jp
Izt6gA95oRkcyB//dzZCDc349OQzqLOY3ysHIKLDs/mDnqmb+u5Du2+GLleXTIzXVKU9D72f8vqa
ddO7B9XOOcqoVztCQP9vvUPvDLqqilp56Hywl+QpIPNdIBd0jIUXxzj9obHf/4JJIVjNRi6Jkzoj
6v0Eq2Tktl/4fKhfpWfE2X0McnM82sZB8NNldWI/1/UozPMfbf0vkfYCAyc0P6JKJKzV0Oo2Af7q
QSNx+vaRBgf9akWFc31S3sUMUm39xlp2sSayQwgcKGoKRy/jhPHRVH0FRkp+pcdCF4f2z0Z1GkGK
z4JE9XVptgBvW2a+4zXAgx0JybWhniL1xGvLW/jpKSLdT7UG58yGA1rPn/bxmLL4dK42ZqIMM3sP
1ZhQY0EAU0kvurL0DgBg571vX9I0Dr0KbGUep0tPocvd8+peUn078i03ID30FzFx6kY0vvZHOnc0
ZgOIHcEvbbKccLa6K2Jv8Jqv9g5vAfCiv23Nhmz7WXqNDrsrVKNyI64rzHFkBV2nZpaTe50/IMc/
LAafSPbT7NkkQmyFxp1TkEGOrdOMDqHboKKvj1ZFWErjbCdNaYPlELxUs3cxCX4ybLkoudXC8sab
L7DWVtdKYMOgXgeOXWPiJi2NPv92nxy6IDzYKBVNt3WzTAAoQ0uphQ4TNh6DjfRTO9z/HP6Tt0YS
0mNZuPNu05k4GecH6nWOrmaL5MMVYG2njCV1VX4PBGH4msCGAHe4qOFaLUCsBNvqEi1K0cA9HjN0
b+SRePZ7v5L3OFHZ7dseIV28AyleXCjlM6LQysr9PPc5yKpahHQPfUO2oVKcoQ1wLCBdHS/ms57j
YGwnTngzUYXF8PKIH0ve5bGBOIyntAJMHUwxzg3kGi1O1WuTNlyNmZ5cMcBE7NP6smTv1jtIgIx+
nLAV7F15C3YCMju0WdUgQmVkhUKvkDtgDSUBzLw/Sp/aY2Gj+Uzf17lc5wEIyzE7nTkbTIrdJ/9w
PTIFh4t+eGoUCq14qMr+d39kJd32JC6NWM9J32JcPfQKzVyTVoM7fy6Rw5S5TOm9s3ImOLRLy3+n
EAXXHN4HxOawZpjNnviVAT7EvTPoLa35NdyxuCWidBxloJAKHuFux2HFxC0zAvxn5Yhw+h+hHFoz
bBHDpNIDBemj2shclK3s5fMHK8WOJF1BSprnx7oZlpk3BlXPrFgF79LdaZPpb363HLgtL+houeiP
qHCkcyux+ZWxcWXjf8nlUQ8svLLIyFEVf95vS14cUwicaI2dLIeqG61c72jom6ijj/LkNGCs9LLq
iEOEjQPNDF16wSxRwV1uMWagrvAtMVdDUXQ3SNI8fhq88DCC4R0vIEbapqmbi5b5Kz6nbmmVbjKx
a6uDmZW7au+SSng85TBv9JSK2URd9CBP+FKdgKuo2Nvyp0OzP76EsaKj7VWYTL1zC2jWOL6WtWhC
iKbmu6iLIp2LCIwrxWhH53DbWgMvyidtiFLy9/j0j7yiouvoFM7ls0E3g1iLi1M5E3MDu21iG3V5
0tqXnmU2kUIfcGu53ae+36Wzd8a/bqtpodPUdsidHse+EJhJk0EMOx36w5VLk8NdQbR8vjfT4P08
BDEd+AzMiOfTf49lIT1Virjr3ZdBhWhZWt84glruJMQWQkpPfCfAZoZmPcY27S+ZlC9t1+dlUG6a
FQ4ZY5wS8WF4t8XCd++ku1ag02kROEOu5DdUF+O5k0kOVyHQOU3haDGQ2lQPQEI2pdwrXRarVxdi
4kxf68xDNA8tG+MVF3xQH/JLhnqn+8UpPSKmmRaOPWpqy5ouQESKeaQEsIwLk8ew7/bdgP8Xl5ff
G81xrFFG+T/63YIay6uLVRmjpw4wvBcmIKE1Zu0Kno4StvNK1PvMKhxxXRF4soF4dVH5dEepFI6n
EmPCHZHCob/fj9sNFLKAnpNT1K6rlWVvo+aqZymmFf9SXh4DrPN217oyXFnAA4Z5qrPzxGt3tj0l
vexSSp/PrtGmYviaK1HFskYBsq1O4ERqzsvEKwhmBh03IFV+fUvliVWPqOsN2T2eOehKlzvtPoHg
8Ckucw9O0Ttesz6plF4Tn83HHyjELmQmz9y7u2apWyAWM/EUIi/uqOGGtj7XA1UNZGcpQi4JVaFQ
E64z0XvAeoR4JwcfmWxlxttl+30uAW24sLveROqjDdGVDA79UtneQZ6jQF2gl5U5PMTYHpLGkSsn
ea1ls8ZjXNkU51d88grnCu+nJP5zJLPXAhtrE2JXp6ihA2R/a7oRQdaGBLVMKUGvBt+/59ac0RnY
XA9sZjK2D/XJwTgX4I9kY4HhECiRpJNR+WsIX+JgWCBdOdNjJOw1FtbJnbh8uCwpQLxWT19DWmK8
4pWjZoCr5U4KRGkfBQCkC9SrSTS1wvP8LlMUaZK9fLEueSciFjBoDMLVLS9AzULVz9h65Iu27yvj
u3jBjrV3YT9fRuRgeVKepEZ5s37QSB6RMxVgQJ9pU9RZIiXMZUiNM6X2NXmuGkKiGQRKxXy3cnky
QAUXG6R+xwO92ZS3qkndAHxQ/JDJikx8cSZPZ3aYijXsc5laQ3TcwogsQbGJ2S3Se56YPNw5uy4Q
7np9C1P4A8ZAy7Nq4hLpVl6VgZ1EySGa1bj2ieJqMa9ETMXkC7dvOYqC4kCWnC5T1YolACFmImna
CnIUj+1VFigBxtiLs412qaEb/M0jFOI5QwPcOXET/zpcOEdAR4vMQvR6s1V2Q2Edi/e+nHd2VwrV
8D+mW8OF1xtJGewDObwuswVwzIc6TtWUOlh0X87uCFxgIsPGHOvnFKjY5UQLV5NWu9V+WIp0dPb+
DCXgh40PnIh+irVarWvE73KZZAcf4Gi3nR8Pa9uwpPBQCSWxaRHduzOXgjfEvHbFjjhTHK82aZRD
VcXs4SU20Ni4AbxquIsaOuZ8ntQDn1FKtRK+AHq6c61uPGwZK2LENukrlvXYHekKZ0+oGtkkTgBR
trGslAqB5amOSMv9MAUDPMIBW6iarJ7CJHFwrFXEEDxpZmPtdnxi336tkwE72IabaiMwrQSfXx6O
XV0Chc0USFNeZI0/NRqLn1mSjmwWBBm5blcLnMYBOOcHDGqjZtCdS8jCqDS8b8eM49GN5dm1MpMK
AlJF4BYKXzvvPWjvHAvznXdj/iqsOjhTB9IoD+0PcMq4vdEHcWtYPVdjnho4UbV2GSiViRB4yqtY
BRWgT2oALuUJFFBCfCTjr/mTd2a+Q2U3yeNCZR2yL9/15eKV3cizNvo1JdZ7PLUZjkd1bHGNWZTu
Z/KMDqgv7i/AqX57L34c6Pe2B0NBNXGc40oAp8Fg8U3eWzta+bwQXN0qxeajuqHeC8xhi0z/CVYt
/7tHrhAA20ebC98mhU3c45fECWDQQRHWQvRowlSm6PIy7YTqWt2m1mRiYrcUQhzuLU7KBudKY+Tf
5Sdbk4+tIO7LkTjhOaW7TFM2Wk/dQP2QoywakXren3kfS3kWV4uIhC4Ta7WSiHcGlACL3Y/b77CQ
31j08jmQgG2vpTclmuW0hNZ6uaG64BSyQQgWS2/HvmVptcVnCMF916uU1L73XCAQE+6hC5qp+gjK
ZvIk6LnGZP6GdbSSd3LYhkqHFmssA96cI9hIkFPmIBJw6QMTgwgqDrDlWsk36DyGk5BI74TO5LO3
Ifr37jK4eD213FE0Cd0yejEz6+UH9oGH5/1l3SmSMvswGTNPT7zu0l04aGr2Goo0n+f15LxjvMkj
DtOQlBejXn5GwjvFvZr+c7Fogw0gyqkaKJODm8sXK56HhY01zngM76qnTHDxzaG5KHt3OB2uhamh
Ep8iSPSTzqp/7VTmUXZIew5eUFELNLVZEgN50Pz+AVj7ZxDxTn1C322RUzqRWi6vfKzahnE69A3E
tjLM5HdCZbqLwr2cHVYsBuK1dvfojh08IehOzG8Pu6921D2wU7K2/KUzo6xrCT0978HnUzn66vW+
JLpFklao0TTMqKIND30JseFVJ20YmoSlfL0460ajM8BxFxIMgRIG2/HMGQFwDaFPTiID/+8k7uBK
47F0pU8b7If4Y++QWitylLJ/F5/MmHvW74gn4Z+CqSwi2gBogfkdc9sL7qp45yGpQl8hh6xYo3wi
C1C5E3kvge8QgQj7gezugUp8ViZk9jgwhXYaTVPVqSWnr51YKdz6Oh5uQt2D6DsNUGiUq39OmxTh
qhtLQLJvsCIcfyZlIwdNOBKP5HJvUZLAgzdn17e+At1OhqjnAUcMtZTPNYsER6L/UJlxtKCVDhJR
NXmHlPdlIUxRnNLfHd8o6l0Qn9sh4QvuJh6ONTlb3EEVxc907ouWEAEtGyNlyz76qZXPGegTtzfx
IuzyFIzDlkb3gDok3ABidm+eD6eaDt/ud7rC5+yxs1KOOlQHVCueOeuOnt0ySOXEGPZxfSJ51dnz
uR/Z4+RqT9YmwJ45GpbOvcWprXNraMxT+34WguZpV4DzeiKoyyc0Fbemw9xOIOB6nzi5Yz0Qf78i
RhA0LbMzow5NKfoNGqAC0jnLfuPa8alMsTs2CuNVTn8EwgKTSBqWOJcADvfqqSKprVF0YXG/DtEb
ceNzgjA5JzRdHi66gO0r/4IDpZ/SXmMnOgxOzyMhRRDi1Fe0TpNVv0YPVTcU+kx2CxbvPQ9nX2S3
Tk+eEhZS27iJ84e/cJp15zyROVW7y/8aXXPmHYdENR8z7RZcy82dF4QXEsvy+sau/9NeLkFy70Nt
K5itBm7mUtbG9au5YkHBRpMUSwcYUtqNAZZdKCjqgZF6fGVSlKhQsA/aiVgSTaUpiTiAdTGz/Le1
gYizjO8dDU2ExB/EoPbgDYsZSn3Mi+Z60LgrGVXYraW0RLR9SIwPXZR5g32Mrq+Q1RPlU5gsyKay
HJiskyD76mSpNgrUmRK8ezhGBRi+LeyS5bBlgxiP/iDzLilYo5fsMi631otzAqOAcXkdcPC9KcRT
Y/ekNHIIrtsexVDkpZZMJxIn2RkxWhFBAyglHPb89PL+MVt4LXDx9NKo7Xvnbf/kVjg10UHQrgKS
218eHRxMDxxSHl+xCVP9KrIJat1KucwJnEkM47wLOOIMOGvEmpT/m7FPP47aTFzp5mGOnDom+m8e
havHwLbiBexzz4gqoyhZyWodqO2M5kFcu/VKcjSTM0IqHdnvSeCofCEoZNwnG9BtevB4XdXIjDjm
koitKRPiZlJ6XjkbiyX+GsUmEHThjHGKL+Ua9K8is3q/agqRO59E5XBDT3Xaq3lT4+h3GXYDKF7g
ZHStM/4NNo9QOYcdOvSbcKM5UWeYxNnkDma79G+jdLRRpnqDtS7VL/91abfkiqg9yNerkSBzc5Nw
M21tuWRQfjDNoB+lb3HQk90hhDWRNeGy7+S/ekIsT5D2i1j0JPMtSYdkeRth7DCfTT5oU++rVlJV
SWWDEEXUV5F86MHoQNIeNrQcAImdCSiWFn2wG3m5Go/36UoREzky4jwCxuwWyJKsBLjPjqUq/WHI
uxxNlV4Ul+ynJDKNhdkD5jnMn9mqbUbqkseJvMbAj4j9+RUIm5O5VLgJHjmQHo61+r8G3ltOAtzW
CozGQJH/R4EfKCcYkFnx+oMi6akxWkrq7sGkesGF/5o2bl47SUWByd0Cq7Zpf8UaBeo7vGcUBovW
Dz06GYpSgYPAbFX2IKgGKESru3UDb5LDG95IdhSH3W9hZ/i9I1oHu6jv3ooEsppgLcfM6KhMjKdq
P2KUTjWjP01DEwHL2/WYGUB/A+ZXuIcCLF/+bEE6a3sTsr/MoklX57sFXN6Nbn9xbt0uxG/OW27l
SgRHIm4c30/2lrwCmXs5GXeFgOsaD1bskb6ITxA/ICFrkhKwvQvWMrrgLUfKiZhiUfejW6WSyIpL
vdx5K4bT0mtU+mMvfq8//7c0xH9q7fIMD05EERPIPAY2c2Ac0HS+TJESVTTwA/BNmW1Cog1BL5iu
HywtUaQmse+so9mUsz8nekeAD13OfFsU7Vx+XDyZZ8zWU1+4ZLaa7kJKDcW63q8WkrfFa7/Lr8xC
7+/Yt9gJdwpR7cytqZTIJoO7g/m65HkAxnOONke7IdrxmHxpF/37S//0dC8Cf1UfvI2upnX7sPmU
ReopCw1naqhF4tkAMt5UvX6dpisWZmV7vq3loK7wMBxP5pSyJFW1+mSkfpNK9GVd4SYp+JQanEn1
ebcAkuG7lbEVU+HRIO85Pnlp19W25MEiCP40iQjyXHFYF9r14RjOJne4bkc2G59HxLzJ9pHOyke5
j8VTEwYGtma0NfREer0mDqKqdp9SjfaellqgsaPazB8GRXasApSRtqVe/Xl1PQUKpT8iinZL0GcQ
AIBVd8e4ZKWxpycBDHP5oy7yeCqpkWuomMryOrgjtOPcP+2dWuCnYN4v4IEqxf6o95l+1F5UTilE
q9oATX2/rUfEgTAdSdJWAFpZ/BwmLElt6Aheu/5m8Vk9gewHu4bdADW0az6AhA93ir6CT6YHwyTH
v1HA2QlzqJN7Z5A+FSVCkyOsLDkV6S2dVurLVKeWd6OZ0wSYOTdCtF1vc0Ieyn3e/PNhcgCqsj0+
rDZ85oXJdxaRoUy/qL2vdyAh7zBL27zsGyIvTNBMx81DEe+Pv5l64YJnVsWAH8cCQcXU5Ji6iwgp
5IVa96u6/VtT/NUlOBcdSUH1kWCYeiJQkQXigDg185OztGwfYwq9mxNomFApSgpFos/oNzN2/qN3
JjwTfjL5rn8/X6nkzS2PCwaBz4NBoDbK2BcEUGlit1acKOz8niOnVLwHODherzVsL4fhMzTp6XsP
6lVfyBMR7RF2nH3xyvrB7IX/rYcyVMNbjxNDrdjHmK5nK67CChODde8C5pZ3cez5q5xaoBndmU0g
jlyZOGJClPF1cA1A1UQf0PLfUjrFzMewuV4ZN7Bm1wrj2uZa+l3ZGBdKYcJWXG4/uc3DN+7dRekt
wIw7ilzUD1DoAXFISQjQ3V4Q28v5UCVWSZsCGW43QzSr5/EhZj7zjhdMAMyexQIeqGLfrSj/BXSM
9c66eXNz3kXw0sIfi1xNTUdOpgbs18DPQgsEXkKIo488sejllC6yfpuPZTF23Uurez133Fwup4J1
NT16YPfz5AFt90KcpJvraKDBeJTpI5inlYkA3DA8UPhM+9G5pX4Jg8V+4x/PEYqOe16m2qkwHgLW
Zvg5sJifnidJksa6vgg3KUhUIgi5SUAgE5Ex+vEU1akXM1QO4KT6QolLDKBIe5w+f2GAYJhiNnrH
4VnZZufEF2Tvbp2VuRLQn0v4E9kCHm9SjPuV8cZUucDebWoN32i2q95Ye9yTGcaGVLs16zKs4L0Y
V6bPCKMxLB5MK/R2hp6qmOygBQZmsHAtmPymF8Yw+2ixUqY/Ftb45j5xbR2kyEfCvcGE6z2V9hYk
6xfvKExE2BLA5NK1if+e5LFiv+AmMm78xJwdlFnVhMpEfpsuVuDMgfsFPd0b0AgJyO0MWn5xgRa5
X3Fxd+pLRRsKln4LknsHVQ9aKggnZIfoseOEo2ns+cxAvwrG/Nm2ENnnao/FBSEEn/U78MSGJAc4
uMkZdXn90HmQWZvYfmxNnO1NFdj+n2O8D2YXKXVfi+vJeGyTOaquKTcOBwXPUMXmz0GomyvHuMYd
1nOulhcsBfPFiMDNCrxzqznMbEWLWYPfdxd4QPM7SxmnMzMUKlCjptwGVLBsDPhRWHMFWZFElnoG
Z59dseZ1DvG6U+7eaJuqfxmOL11fAti4eZ+al25k1XXFjJJ1xrVAc2wBXF6hzJH70XdklthdhlD7
oy9J+1BrZR8aQz4XSzA0wvxnhADKP6s4aOKXLZbGxtIB2N/WA0jceyDizxTsGMW5UMVwThJ/Amky
jraQqQnnkUPmHv8jtoqcfY7kvhgg8J5E7z7+Uj8rjaAKT8JZYU/M5plDA6DNqygWCj4/bNZjkq+G
bToS12ScfFd5TrN4BURLQ1pIJ1aSdQSkW604RuCdWkZfHEabgkJO42c4bNz32n3OjRNVR9SfUnbz
od3L0av80Li39etDp0rkhn7z4hfXtP5OXDV5JzOlSgb8XDcWkwjE8vQLm2l8KDHY7G26LPzFe8CR
ELs7CkmUDOQqE3RrxxAw+z9MGO3iHsxh7p9e/jcjl9JmnTXeNQNxmyglfeDptCES2+EuoRTUw6Nk
3W8pEqZwpY9NQXyYVITQC6Y75S+M+Hm3YXvhedEpB+sxYEN1HzLca3z+ZV3D7yRz7rLdycOWDUcp
4IZenxcnQKcjgrPhU3TjCcB8HqU1jX7hp1KHGXOpU6jvjO2LEFId0MVr+TAGdxOx2rP/E5WDd+ab
YgQNZgD117y0D0C4uEQAazofDyl7c1tST5JRCKPg3U7ld3pz1Doj1DAfno2Ryy4Xr7yCYNHN938+
zgyWy+U75S67Y5Xd1wZSrZ2fsO+u4VV3RcxTgs+XA4K8+K6/LMadaqbAncu5lzVdsQaZa7FrgcMt
mY9l07JeTbrnz+fE0ubO62YIk8hnfbtQcDkQD2yzQSMj6UE+Zz80jmAFUf+6j1nbW2HbYj+5zm+d
sIiUz1kXCYn6Af+Cf7PDy8GyPv5SDIA2CxVs7p3/cEByxsVWoq3jiAmoKoWMrPcRrznAbg1LqnPL
qUUGrwxz/7T9bR8/Z/p738I0h1j1GDAHWf/B6eIrUS7wyWConuQczYOlfiTFjApd9taG3tK6Ik8r
QHMpgRPh7AOhKFnMsCNqJR3Hbl5mWTUnYzJ/N3OirTAKUivdlxXrGEK1LxRpRkehCLsY2ceE0Gzg
FH19Lxo8U3/7kyknn3ShfeP2QeuT+w6QgaehfmUNy2O+AgyGmwcVzXaDTBB+k8ASlQg50CirheLB
pWW7s0tk9mdlevT9p6kW1WWiatNTM1rcqDjFCkStdaA1bp8BTGXup/0DQvFwRPsOqTskwaC5+XZA
392KNQlbQScbdgRNcae1TBbnzn3PLmckRZP6t9kn1nOEKqN74858s5n287O5u56MkqwO1u7N8vE/
bosphHRI8RCHN3UzNt7KYiNWkH/I82438l2vfpzxGuUEMY3Z2YLNZh59xRfGB6Q0f6VSjKjp0BYu
bCRzhi9qwt0OiuKSNYrbRba6XP1SInHD0g2s9ax11zFLmCkAlYiebjHJw3BC9CdqoJZ/6mXuHIqd
mzbpRvaYN8XXkWwe2rWzTRFd3l58w+6nHuTTl/6aPRBqybFMKiToVcWIHQym7ynbWKX6tWvnu1r0
qs8gVq8fw36ecUJhSsyaW6x3tkaOx4+JmAiaNCrwGkLcTiHQwGPolAoVTnXbvbIuKE/vy0Er+rAZ
a8AtG5qpuxHONzihuCvRYrw5BDw3Dz6KQ6AhWu/YhxX8i4qbsD2Ziv32zu0Eo1rNZfGmSWX8FF75
k7+eqLj/SddSvwg972IUolvc9+NcuQT3ivgnk5IBD9djMJ6B/ju3i+oeilRkUyzF+cCwUimIpqvD
XURO8GYgqS05MlCWhAOr3b6be6C89sREqwR+cx1Udce0+Z3XEd6l6f6OX8v2CfgB1zpeKzR7ly9V
NALE+VA02o1tgideEdn7A5HxcgHzUchMc6BSYhhCkt3yxBbALJ/fHlusST/6bBBUCUvKpe78R6AZ
r/GMFp8QrSuF9t8BF7/XgZMpV/Kz3GUXY1gkHYzZYkfJLOxiHOveXUgdOho9sMfr5Zg9ECSaTA3p
sEf9KppVhmevCZcU6aTpdmB1L8J4k7cC9KBH4gbLWWmg9nG69ApIn7/3t7czuzdac8faNb+yN9Um
GHdBdz79kqOBF9kPup/6r8Ye6NdNM83bftrRjS4DJA9ZDO2xB9kjzYvw2Hi1IlsTNA8VBe9farMp
jEyUvjX0sYwb0PXhGqmo4CNLEq9B2OvgvWS/5lMZ3aNO4voGH1w9gZCKZ+kip8MCAawhl1ebB+JO
qRXOH3cMMaSRumH3FoE7FJG45qWZjzIMW/5CfPIMheu66x2P6F1LoCc4AOgYOIDHacRVNGXXTA44
PFQ22Qr+JKOo6cmPM2Qvz1fEKYtyOJ/LBqZ3mlZ041hukvxALhqmJp/HiFOqX7N1fDe5jxfErbRH
XhHZhQy/h4flwZeXb+mPtbVQgtdvuJVnS7nIYi/HdrxRlBPm3pKz+OU9hBRwTrsVNxXJbBjk56hz
K70Vf836/LCFR5kpu39yq0Uoffcqnk5quDChq07ivwqg66xOz6K/IZuI1T6Vr1Htnx3ACDHhqSpu
tWRsjtF8ctJozLDqWHwkopPcK6orwzrl812NVLMY80wp+egfcJ2vpAbhn6YeEfsMicyfYwRKvn1m
ZDmAN7Nf1tlO2T3pmsXWqHiT/nYsvPhJxv5DjK5aeLntN3/ZEJtijHiqUHKrWsCwyeyWV7xUKV9p
XbU0HqfRx20va/xJTvLsgp3nypFLC4WyxF6KdZ/mH4GC1cmUkZMPume2gUt849Ig+enlD444fR/k
R2wx6sAqWIbwaILye9rpItJwkV4HvMWg+iHjl8RbMebJYSF9gmfeEoOOpynZfLXpjHaByW10RMuG
9iJ95TM3XWA5aag6UvELUCTQvrjLuIdGNteYo6JElcbjBVTGhCE7RdjjYBA8vaUY34OIskEEiWpf
dQtaefBUcd6+ReJlKmcmYUP3YTKtaHqtAUo9wELOmp3Dk7DLxG/netQmCUZlSdz/o8NcsPS2xr35
l7/7U2EjziLRuCK95cuIVlIOlbx9PUuilrbua0QuWeB63BriW9UVnSQKqxtanJJINDb0QYMI8ejb
rkvR8tOjFImbZGBaHLwU9heMCnanBW9dRSFSWuM5+hxriJdugLAXR5rOwg/HSoL/ez3tHpggWlAW
vrBza0Yk2BgcmfjXYEZ5U5vr+6Maj3ao+Hup+1UGRCVsXfe6qcHu2FFNLIbAP1X9s4pQN5fQpFHi
DKcNgyq/y0e88PuUNaBqU2lXv+I6sK1/SGeidjHDn00ZZB89DNypQSU6wqPsWKQpWOguy+W8ZAuZ
pZxc77NPz8QaNV4WHuhLZaAScumr03hJCwzyQbwgPsjtGDGX9qblsRDjYZXdBHkq6UcaPVqtqSsw
vx6ck9+jXXT13jXLrZejz2Be28WBrgNJ56JGdySq3/cdE4PmRh5yBLvYKEGsOlvQBG+ve0V+T95i
uJxWgidm/rA/FLihM2yvJjUlZn+cgPC9458dl5uyIIBSS9w6v+nFvI2NIWaDg8Mq3qR5JF/2R6Yl
qxkTwhYez9lRRyO4CS30nDQ8NdFdfNByb4eiEQk40m04buS5saEZZPs0XCHxoPr8wI8ZtWcRXggk
TnYeomNa4J27fVTr6mhbuu+M/HLNh571KJmOOyFEMVewQluT7SCDzxJEMGMiYSPVLK5EFvNcM7zj
JzmA00xFOSPi7FVILxekZxPpSeClospQFSbOj321cy3Klth3Ya/hJubwah5Go40QuiyxYhResmqL
mhfE/ytkM9HB3/gChhqdumKgCH7ACnkLZTme00MVSPf1c0STv6kcQz6rcGYrscBANi763eK3P4eE
i2bqoXAj+XKiKjI1Ux/GcF9+2HnEKDJswe1DZ72OQksv52slQft54y6YzhBvt6OCI/ba0dP2qFTo
N/83/hClvTcdauav2Oo2mRoFVi209LC3eM1MpqjvgQQcdQ7Sw8WCEQIlh+oZulDvNXYjpWGEJM4g
fCl+QjW+hon1+D0DsXznruKE9ZY7orSYddatw1NvahUtk62F++BwjYfbn4O9ATIBjVDjL7zpnY8C
JkCzUD9M8I27d/D7fO+nRbYng0Nd+815hxRKLndGC9dx4zDBNOziU9loDFL2R2SnjqaWyxxG/Ga6
LeMU7RX78gg8LyIA4y5YNLLW276xq+70aJT8s3aDZBQJeSnBJnBn/PqBs7acGPSJINhJoHBKpYbL
nqVmcaxYCa93jRBlDL+qJ88meqIKXI5ZGxTmzJEuus4LvC1vI/jWbr/G3OoSM5z8NJXGXzFiKH6M
2M7a/fVlx4dAcpGVs5V0iCmQB+qpbHNwFOx3mejmYP9S3U6owkh20f5LsjQ8l7YyerDhU0ysHi/S
+AGmNc8URyBuKbBxT2zH0j3IPMkictTwPiT1feRSKfkHpPCVtJpsUPYwVIagkZ/5xZCYN3MP4OhG
h0pjiY/0rkKCQ8p/FoJR5ozjSNAQzZd47bo4sZNCLRf9jaNr8remNKnb1pxjbjlnu7YrUBb70tKP
ttBqYum19dGLclP29rqPe68X78nUTROrSG0qyq4Ph7hje5ojJxfsWkmJlkX1ReafqFYtRFGmoDFA
NpGr2gFFmYpdIOY1UETA9P51wQtgrq0N8QQ1kH2bgi14lQU1cnxYrN7xsFUiJ2hBHuY+Ft6+D0xf
e03GV8aT6gc65Ftt50bzNKHN9OV/j95kO77EwJlHxp18f5zjq9NzdequhCf1m0+Czm8l3cat52cX
9CW3qik73OVlrRs/4c5XBL8crGvD/x6KHes/83m/y0w9LUPnH5VthaKUBXvH0RGxO2RQ0B2lOWw7
njSj+YfSMADrKAAFDc+Nr0ztYPhs3QuhHzaHylUF8zDXol3gAwtPy4zLqVDAXO8qFhPBeGjlnsHA
6hSIqgCvft3eaX7SYtBggR97/e0bA7Kf0hKXJiIpgOwGdDdjwAHksOB+4jwwEktoYp2ULFRrAKLs
a7806ZYIpNhIb5h+3pBup/ptEHjaSzMtAE7TYdFsafzz+mZQYKanKVVRtk6Dc3x0cyVaHDhmEp+q
rrEQgChjspFxyuLbavgQV+0XNSYxuYIfVoiXbUJpQK++KnAZ3UsfP57iYsqhOgiJsYHxcHsgjarT
avVJhSymJqSVvfYpe1utX3dMw4plCDsKhfLjhV1wiYLe/BLZs3I6eWsIl8fzfe805+8zT0AcdSmY
aF8GiE7ho4+/MVRzTzpwSywOkfV5OcWRcVdJO7RLNIPgM9jlM2O2w4qiZ3rwo7FcIA5ks9y6umfT
L++Nzs2oucCO3MqyphwGOv8yd5BwqF8w2mtvu3dXcVerzPG6UXjpazPu2UPzmzETglG7/RXTz+ZT
FnvCPnmLfIZObqz1eNqRTfB2NHsLF9emz/3l1Wn/1DwEkzq0m4rCzrCr3PXczcsFIzoGh4EmfmD4
qDfkQlhgNYHiEutZMlDaeVuHVk/OJrC3cckxh4JoTiRTe97UiV82pR2DC5euvTPDAlvQgmDHlkQE
AOXPyE69n7WLOJTYopjFYdLF+zHClv86F5H8KrMcoK2osWGhvLJFnUKc/q3/toPVATHPxijZObPz
n4aU1njZ4wmi0aCJgthrNKdFEQlUE4LjLcfNaq4R1htoC9MI1GcW2foaLcG5ovxLREDfuB7F0oMS
JoxnwG1Q3NfBUDkIVFkmYiJAcjPGlnCy5gO2Baou+4ldcQ+kmEWwV2luHD55SdvlXUPW4GDSj3l3
aVwVJ+3dbDvVJICVztc/efUDKN6Qb6SgY2t5eYvb0iCNC3AI5rd9z//HtSytsIAv31lVLVHxLF1L
vvOSugtQxtFYKccEkAlF0ZpxX1BWuaWn/EvyxSvcNmV3vxXxwj2hchg0hamTBJvq0qEGQFaRmk8/
6EcPv361ocAFJN8nqTD9TSAvekLE7fT9TLUXCw/HbUPVz+KjUxBgkP+kTuOAlUBEqTH6SCWFZ1r+
UEsBug888tTpd0XwzE19DPb2MKrHzeSSd840f8p/TKG31yeOK6siMdRXn8u4XcMpEVWEOrO6CA3E
roNns4f4uDE2asa63tdsCOeSzTkXycl8NSDoR+qUQB5QHLEl2CeGTwWDWUucXwvmTKDmtqo16s+G
hrPIDF6ZEh7gmoqHO9zI/05z9Eww/upUwvrWE1HRBg49rP3jKd6IZME0F59VBlI2J3PRgnQQtH3l
SDvAPOlN9PiaatWa4x/cKdDLryxi2IirFVF1dKArgk5NOko+4zn3Dd40kxncD98o/pu33y6i2qWh
aiqp1RBoz7NZu0q4xor3WBJRD8yAcT+/4fNtm4qElxAi7YmgGQ9NYWwHZ1oZM/5prHRhXBaoSwob
35VSYE9dDrqtzk0EYv/zfdkzfMynNwQuaiM8bfV+cKr5VwpLlDlVE+0zEX3JTUHNZj9YVW6migTq
/iB9mHAb58eFvXNEyMyD1metwesPo67EUeIpJfBFLNbhxQ9NCCsGB7Jn+8v84gylPedborfw1Tme
MydPh3SvgqgM0s4AcmPgH87nhgSfkUoyr7eyAhXuQ0dxY01ml/yTssh56h93z0vfN7gcjJEitH8E
9q6OUvBKptNGY6rJxmguJSHDPH4O7S8pQpQnqKqsKZvG22wUmLSeO53kj6CIaUISQxIJ6lak2r8O
Vw2dI30anh/y8swNSng0dCTpeqZtdGNB7fq4KbpYKsXrCvtC6eeEZQywn6HbCGxl4YW7AaOvlvp1
4Zuf+Ymn6NvF6bVeYpsqU1NiRouF7JV1uzEmVMOBlB/RM+XBDgbk3aQE/mbkxSyTtqY0EFVTZjch
QzdGbsSR9bAzARrUS5wH7iWAzfwzkdL/6xqB3eOPsl7CdPyXq/nthmRQs26eTbQ5g/UsYINXwO00
vhyu0OA1TpC9Y1vypvqCuPedZncIL3JIEcSzeZU6xCUzTWXXKPYis/zBJkK6B48FxyoMaEG/75Mz
ddg1AYh895Bjvh06Bv1NmX6pITzNWtBmmmPuqbTQz2TM81OpDmztlkOFCR9VmQooEO7anQGTsCWt
QLLJhnMbc8hD8Mw+17+268cYKOIj2txHVg3N147ifH/7a6MBmT2b2GLizqz3bYO6EJP4LwgWwBzh
G3e2rFNswh9jJslDzyHhEnKcovQTOu/i0DsNc6IwsdFMMriDp9lWuqQCkyBgc3PyhrvvMKxzSSaY
gE0bTiiMoKSPQ1gcLVtokIxJVNbxEcZwPdA6BzwLhZzHaq94xFPtAk9ayZJ+ATthaNivvyzua8YG
dNRLYF9zkBYQiczmwxyIImEc3l52EdLssCdVHaYMZOhpdBaUPpinTYIwhpwfY+SyHz02kfdlTL9o
WzNh1oMkA2I/pBK6YswrcF+YFvoeuVNe6ykiN9Cx99VVQQm8LG0Y7yWgpNUE+ff+hs8/XIiKl1qW
JIy9FYaloPjpoMG1UWUJqDJV+UDtSpoPrlmfycy1uZyELMrjTOu9CnMf3kPVsohL+loqUtllvm82
E1SSEBAq4BxC8eUntR4Nf4SuSul+yTV4i5vGPr0UEZ3mq/lvnUbuKnl2IUFx1xz5RO9LHZvC7Yj4
DA5dJZCeDuR2s4TiPIT2+ej/OmPf9LyaHUtAA/PXJVrVNlE96H12dEMImd+RG5W6r50/YJ8t1DY5
UNOp8Xa6RwvBf6P2toqehZDZFGLZMm8iBaekk+aHAlzdAQ0wBASQMhpRJVJaszLfaqF7n9WzKB9O
7uYrCOx/zHn4znx8MC8xo5N33q5cKnF4IZ09aDGgznIPHW1N7DXS3MuhON0Q+zTpXj34Z4BWR5oT
+ONo0LToKf2x77YM76kYc04fSekdzVh89pt5e7sypN2roGO/b1AdNBqv5QSIU7j0ga/riZt8sG9O
ugOWzkSiqKO2Q8EKmg+ZA9PFVRQ4xFt5LRgWcb/N9X2JwdCK0mIZViLVjpKiIn2AofzeZy0sj6P5
uJdCchzMxSfjWzbcQCgiIKFcqtJLZy47W8tdSt4TdBgQQ89Pxo8yplRy3TdgjOHPX4kyEyPRRPRz
e2G8KalKVIv3XEdjVTC6PnJCy3wASYBE+QfHXoZYLU9HKIk7qcoic8IWcQaMQ4ZoBHkEI/bB+JrY
AVm92oDlA/sx580tJ1+3D/AQVozauDwaOnB/cr63+WcsKuXt5kvJDlOx+bBhp3FOR5bKQWhVTMvn
d+2las7f+cByP1eR2JgE4IoSwlJNxzS6D0gPDFUbMmoByPxyaSLECLGfJwb/oBlWa0TDZDnDd5g6
glU0kpt9m4Fl629AhHhccLHDD3fJF9hFoDCkV5GzM4Gpz9xzkH3X7A9/21i11o3Cdk04K8Ks3ukG
mIiv0i1R17aftMvtjw3XF9Yt/rA6/0+LBdPZFtugr4URtDjkwstUzs5Oa8RlixmcdZy1NCBb3hXq
IHBE6fyEEwmqmQ3HaAYLnnrOpM8gjF+StrKkctmF3aUdvz1hyIrzZ+2tHc81++YWqc8oU5gI2kHD
T01/Wz+USQTeTIpuyGfk+Ynm92Uj9j0HFF9VTDGqmeC9n6eZdA4aufm73/WKMr5/9JXcI1HlTkf9
zWOZzjXcKJaEarYde9gI84k5nySVUZulfWVV64kWk+9EE54bqtLbezEY07Cus+zErg5J9AWy2Lw3
Ll67ZZS6EzLccrgSlSqZHD774geVYAsFXVfZw1i2lUNvYpv6Tmer18no3NOrw7b20MDKoRDwqh5i
rtm2QivYKXXYCUCajtDpwJWdJlqHCAtwn5S2CjttGk6vGBX70ENdj9VwcQmiK/KCWA19FEaqBMtg
n2wOlj6iky/IgtR1Fvwh0O4KiSHkXrbd/9H8lxh0E3fhFDx+3YZYcq5SuX+69kqxNwXLTMykSOB+
TxyvYSYEnj360jSpu3VakZogoFqxnTjKSqqXBIU2fQUVrSaH9qP4AVlT1atPROe4T28icpxKS4q6
lgAtqmxPcmSniJlbxNfYL/mYAJhkTD+x0Py+6PgbPiIdmQKYP2JLIykXIQt/Tb4+L6kiR80u+6mK
XAluG6OEswPj2qYbVPBvopGQ55ZHRBMmnvQbBhJWKv+SKpzBBjH8soKmk/0wnfKRxILmh+IfcLP0
WWlOZ80jCllvwfS/GWiKRNXkneVitqYRXIQ5KxGmriw/KNHrCKKjybU2oemqB2PEfdxjr74gAJ6a
vz3/HnJ6+bnsEYLPmFBUAmJaMntaYh3zk2r1mvPXv7NQjwwvMDMoAefphhilpHPu+AAAXC7MwdQn
cxTihy6SXRunkPKpBadumTDsM4+VQ9060Ju7DGRK9V2PFN5xv/gydqKW0G2cE4ER2ruO6Rn3+VBe
HP7uLXctFiWHHvuUZ1D1p9sGjSjXlKPP0OuM6+0XzRUDgQd5yrKhOVEAR0U/PBUxXuxz2b54cwsg
k055pcfsJA9axBJFBFtWUg1ReZJMMiHh5rOmCjptNddW1053CFr7/nXG/ynvUDHyd+ZA1ifIsGRJ
g1wSM2RwsRRan3J2Peeaha1LJjiLkIDkpCHfrk6XfjK+UvkJOlCVLZW3ceFYMk49AWEiwpgevcbT
5xMPUh8n3i94V3zCkxQWb6+HEw0P32eBsKlA0G5cjAphx1mxSMzK8aqn1/ycplVYS4LaknJRfdhi
AuWKGfXIV0L/Zu32yZrpNruoHVH2UyOXW2Y1qbr82mf515s+ZJOgFezvbeEDoS3OUUaufg0hKB0X
zhmtFc9y7LLyKCqE2zUzgcyrxTULmKTs4A7uew4wEIvIoVO4S4B2MPtEgzh8wrUiOSHycQ4ArvxA
FWMpyfe4GRhGktsic+50BlWKpN0CwqVd9pJ90DSuGvgWlg0EY0Y5EIlLOoGici7PViQy4Oyxq/iq
oIGyoTND32xupL8sMxBq/tOCjtJxFaeKe59EfETKdfjSO7nhCl5Gj7cRuMdTAicZKi8zUD5AbOkC
w/FPiCGiYVIpf7fvEh8b4YOflQoVJtKaD/iKN62CL3Xmhk1cZHrBreYRtSkdL5quYVrp2fXYePQV
JmVBbdWY6cZU0lrbes78XtfgLdG3g3eYKvjwBnC6dAxYIrwpodtpXr0wy6Tyb67mKnvORvbfe0BT
A/YCF507cGGSIM7vXHUS5mKdfQbzQ2+AtUbjaEu3pfDDCDlW/UsC7xxM5cjXIGT+Un27vbACOqcs
pgy4uheQkaiDYK5OZn8iVb7+6AD+fSPmXzEqVH9/3Y4G9HzLU2039FcWVLsI5jXYP7dUsaUDVnWW
5KK2HxM8/SqqhUYCIsGub5yU4T/2Zw+RrlbeQDij/4jTmcgZYCqCxtuWHvlG0I0Z6eliEjGfevKh
dVEgSQHkQ1BzYLhonxBT6k20sPQwjD0riJSgThXA+Ero3vRF0jupvlgIKRmI5tTLzbwfEimzpLAk
FqcjhGSm1cvkTTKNxXNf2SqncJemBgQ5vTTDEQcY9deVKvFN0a1w5awObVBtOhPf878EDN1YNqK/
gfBEtQ56qisBRfghMLKkMY0zLH82E/O+DlqmAcczOLm5FlHfNbJ78Qbes/eQ6C3aUYHj2WavPK+r
vUhykz+fuveqIDIuO0bVwr1ujBeoRfDj/BGdZSyWPA81yAiCpfYma/yEsZ3y3FzNoS0BtHC4U0w/
JtNKgQGdlDY5ztWGfLm78UM0HXNZLyN2QTpVfGHTGUYFTiFDbunUXpPAc5kcsEPgujAuhgY0tu5Q
Tlfi09wbnXp/WZjLLixRMOayxLwCBV4WBYFweDLzkVPLvUPnYBnOT5K/ySoEuJh8syXGO10RWWHr
WjeJ2lS5w2h1/nNItDNFBoVZ6nk8LW31R99K57shORA00o/8/o/5ve5G0+JcqpVxK6LqPghxfx7q
fxxBZgoF2V7zB59bh6vequJwXBMSxaD5M+ggaXiyiQg71MNYUKS23fPmQkj6gYShIuBwLfdT0X39
pqCIjtm7hyx4nkzkX5SSOtV+7uZSoM5/7O9FecmNt2TjGqeWizYNRXnXQRdLXi/z+IeuXQtNfO6y
emf/c/99Gel/Agb4CrCis2+l7u3uMxywZeTuf8hs4TzB420qvAWMgYyNLM99kK4W2esGoi8t/ZX8
HOQWKfleCHKL0CbDdB84wKT7u57q0PwPEt9sWtc7zbBZTK5GXZLjktvH5dI5RMHg60hVqU2GfqrP
keJM9AKm+rwAJU+xODppZESCqpn7JJ05DuM6Dn8op9swdnswnK6jf89PJwIbv0YY4Y4JtED98unU
Z9ss6ubStLkOaRhGq8PO33KUUrxstyeDIZs7nkXhzzc6aYImhZvodkdydYL/VqFoEjcImUmclZu6
o+JS6jxFbxJfEuh3DPl6ei40qfq1CzwK5CFMvsI0Ojxo2walYhTdxQkrd8tCnq1m3awluN58kcBk
OAncWUMopaDTp88pXBWEcAT4EJhG0iasSDUjvctAqPv9628Ut6WmxTAZenDZeoHnUN62XVgn3moU
kLzHDSmxI20lLR2MYJhXTMAxvpz9jxmbPEs2AimcYNfqyB3yJEzme33mZMxNGUn4Qq5QJYS98nfT
gQUi1zKHR/UiLq08ImahYfN+oX21XlYDsMy1lyQcvTLE7jeGlZm34NhNBy0jpjYEFNbqbYxQFYC9
h+IK3T1TkybKZY2Ie3HQ6OIBL4f73OGm4XQQoe3ms6utdH4TJtUkLQRDhhEH3nTNu2KHnXzmgfrC
kTn8yxY9L9mlnwez878hdC5oPQ1OqrO0uMY4dBwJjan7D8/jXGAQcmSFTKJgr7pvlOn6WZ88lmnE
1x8w2Jtbd87pVfnxlmXEJyuXgfPRI1bJFuaKCLtsoTtMvuuYTS4ov/ZzZqsr90naxQMiQum6eTiW
XnPVso1igGIniyi/Fm+QZwKXvxRqmvf/Nj+xW7/ntMik5mms6M7XV+3QDmYWLGLD4ldWz+pUMnJn
ihCUwRDih+X1azh42KBDuhSCfu9HdLgVifv3TgqmhK0WWYawOEmTv3z+us31Mw2yG7+zfwdE2aKV
O2iZs9EdRqfrKAafltdrvnS1l9XCNYoyHm5LtruR/9h+2rJkVG6SVosn5KSxqCD1xlDGXWNx2OKk
rGzKBPBdZtaj1F1CF+OjgTqXgI7Pv1r70ejoNOnoZGfKhg0l2NuRZkAHwUcH8T4wZwxsf6ZZtlAz
qe0nJ/pf8HS1OiAFYXqDbXaCpDD/l1Dy61R1MTISUb+Um50AkPI1QmjR1fyIUOPElZALPLi9vO7j
Da69Z3hgCBkbk1BfbdDfXcZmIqYV7fQtuCzKkzDrQNIP+8Fb9qDRmYhskxdX2KO7OXHN3bA=

`protect end_protected

