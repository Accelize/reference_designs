------------------------------------------------------------------------
----
---- This file has been generated the 2021/11/22 - 15:46:18.
---- This file can be used with xilinx_sim tools.
---- This file is not synthesizable and does not target any FPGAs.
---- DRM HDK VERSION 7.0.0.0.
---- DRM VERSION 7.0.0.
----
------------------------------------------------------------------------

`protect begin_protected
`protect version=1
`protect encrypt_agent="Synplify encryptP1735.pl"
`protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinxt_2017_05", key_method="rsa"
`protect key_block
Oj1QNbwkryZZeOyhvhV1D97NwXvr880jaTZgvwjSRzYDZiobXJ95iLFzC9S3a/hF2QaPCwTQ0eHz
Y2MJH+v5SDd+f3k4YhbWDKVSU72dDM2fBuPvEZQxFsmMUPlnteSb04KW7bkgbOYxpc4YnioLKDQa
0hIGeAM3KAvVDgULO42bw+WvcjQl8go2gGKYGKU+OHMvnH92+eOkcGy2788oHBBCNjke+ehY/LtV
L6R+INhq3uMpjqMl8JwJQpBQ8WSfoGDuioZRc5zyu9ly+H87dnIUP+nQRZOfp6t3HroT/L63nZ0/
S4sj27ugdeY26m0snRxx31/nYbVicpL0visuIw==

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinxt_2019_02", key_method="rsa"
`protect key_block
GwOAuD+wk1xlfTOUJlKY3l0ULNKppgdHW3kVkGH5gcWxCJR9cklZKwcETu4eL2NRaB2gQdDKv/iW
0c4DTyO9DuIf8FuxFFUsA2K1H8f6jIFQHemo9+4srL5Cmtfy5xY6vELiOOQ3qM5WWm+tbLbf3KfR
aZ4spGmpjQTiWpGrJj7gBlDRPNJttgtwoVnmbKUmWgyLeFdpCLUz2sMZUQ4F+TdSOCdetTm0wc/4
KJYNJLRW6LaUohAnjgGOYzFUWtEd+P6pEvS/fjoXTvLQFUzf2OmZyQc73LH+GXpNNXBhJc2JVkaH
krbL0IQHWdOvq9efevRWa30OtO1eDxF9OoAy0g==

`protect encoding=(enctype="base64", line_length=76, bytes=869984)
`protect data_method="aes128-cbc"
`protect data_block
ncWSZ6d6V5EmkuC+MFlv+v9zjBurd9MM54EFpCqJ6alboN284qtyQt2u4T6phIWD9sQrWQsUl8Ph
Wl8gSYPl0KrGduAuOsFXggQ0+rRQjvPQyJDnaCke586Veyhy2C/kTbN0pNuLsxPkXBKWtzfUAkD5
e2vmDY9CGKLeDb5dWwIugmcZq4Dc4xHMu0Co32U347H6Aoaeses9YRa49Ru2A9R+GomVg6Rwjv7Q
5N2qGFP0Qx9LCOSBzQj4J45LU7sHKTTmjDSl/cR59wkKgeOIz41EWuZVGQ8MHt0AKBJG9Iz+oNXK
7YD47+TwcOD+hzpoSFeGMG8/Hc540ijUVQvjCFmbL0PojCO5enHvZu1BHVJDHsTuvf7lRPxDeGIK
+hW7EGQ8KZKFUrceOQi0zh6BRS6LYLx7EkMxEv/dovFwd0Cx2eywWl5Ep09vcOwtO8Wnk6Ypm7Md
uCkyrTFcKFCQ5LigZ/w1xC6iFTJgdm7rwGqaDErktdIp/wEi3gGAj59lzi6EPUHCN3QjpxAcVk9S
e/eMeWzZMOOMVRYL7434+ULQc0J9INFdfadEJldCBt4i8CZPhkVnzQXSS0sYxk0oZVW9Q01Bos+H
ab+bJF4q1Zl1AdbEBXCrZzpHg511wL1Ry3K8lUuLnCQw6KSODR3577ktt9o6Qp9Yf4jDeG6t/Yfj
WAvqzvHgS8TrO2DRBUXMEZeRqQa63m1r5tES1FhKVi3+gik88tZ54HnGMdaR0qUfDFPSRqfynmA9
kn/wKEVZ8JiijCNGfLMyjV2ubfRW3nC689BxXCYPl/QWd4El5XfH6QCSXga6NtVFeBnErQmVQrjB
049P32/nK+A45HxO8IIhH6mCfb8UB50sOa6EsGy7R7Re1DXuP1lUht7a7Ix8UJZ2gciPtEHRktz/
bLYk6hW4PEJmB2tJg5eNUdXZL5ZqUKQ1ClUdA0/Du4dMW8K+nYaQgGoacTL2b+XjlUJZydbOTuji
/qPNbXF8z3e3wM3cy/nepsr1EeyYrWQS0uqqyOgY597gzOZOMhFB6l+dPpdW3WR4XDcdc1TjH4qa
4Zt8GD3fCSSvZttGj7S9bEUW94tgVpLGAII4WcVnjlK+0a25FvaJmHmcFvitVj0E4hTVP2bcnyFg
0NwHQCJcfWp03SaweDNRDdsSOsiDPa/mQ4vLsMJN0uKRbQl+tAMNVDlV/gxnkvpDyx1ca3pk2+2/
jgHFhqZTOQp/f3HpVXA4OhaUQbp/Dztya84A7Ky+MB1SGyJZMFl98HT65KJoYGIlWaG9HghHgPJx
FCGzeD8Y6FU+iaVbKMVMuVdVZHBaxGAqPhcFdJ+huKdqw1wD2sNFSA6uXUwhkXL91OuLUVO4xDTB
YYmmNUNZwFz0QNJ7kUTSPKRgXpxnNL3YZvFziMARV9FTEB6iYzqcwaoR35hUerEXuhZmflCDYKqG
p3K8z5xL8vmWJSEXSUyNMF32N00kZUHRJhZ+751+p34oGlvAkFhrPSfa9odo+X2lFaMBS6bYyvi0
2WkKMS/PaDg/3Ux9mJXACd7sJPM65tA/VJnNNeKh6ZztDSuNe5ia6g7zkEsEZfTfDYzwB7pDCnmy
PmoLXoASviPRfR62qA4EompVV3Gow4aUBbWPZUdGzsCctARhEsGi/I9kfLKMTp+3E8Mkk2K1A8I+
YNYMKKo78IYnq0i/n+iPbaeVDpHs1OAzVFBRPvm+oJwkv+sqMDar1eXGj36m6mMcRLKBaO5SwRhB
HP7828XV1Rgxl1KiXl1iEueTyqi/gdccIaLw6KedVdSGbDiWWUohhFWrWVjCz/JhDebwJVfkXvzs
/KO2T4Tf2lkjKe9D2m+tfjnVvRjKQfxvhYnk/RTF7hOLeRlXLQdg8Iv8AjVdR29isE7QViQaxxJX
Wc0Aa5hau9fJGGbfU81dpO9FDRjDIym+F7kOlz9kplNAk9zrjA31dZSYWGmteOPMqORFR4xwaToW
KYVYcQyHb4urdGEIYEHZ16g5PqbyqfxIK1MQfnn0nis0uiyjLXBbNWo+NKFOR77prBoCLJaUyOWF
yh1qkCBCXRiCUNczO5H7XzWtCv4N6vAxwIHsAvphRxIHxvPRbziXJ23Er4aMVO4tZc748Tg01BaT
MXPg6lMZ+IZY71OAODfc/iY2YxGBqapdVRD0keZcJ14F/N7if3ZvvYobdMGK251iIdHtGjWFJZn7
1KbcCfbahEOmqty5aQwL9Yjc/cQGVxedCcRcVNh7bNmaIdQbGGxqL5BQMWQXGjE6dGCC/3catZss
nqHyFhhtV2/kIK6c+IO0y8AloLnsX6W32CyWCCpPklq2G/VZObb/Tb/HPjJbcO9stR1uNq4ZZqq3
sTlPmXeR/YCIfe8H2KuzQIde+PDh4bxT5jKpdTZy+DGw3+THoCSVjB11tXJDCceh4oUrNHVwWbQ1
pUvzREPMn1cqYBzlFFzeAPnO3cboYPxwD9fE3GbIGCokl1jAYmGFY+sL1s0HVL5zMqWkBOTFawbK
zDfTVFRTExC9LcWZSLV4OiB+3nnpt8f7Jeddd0pVuBzDl/8VA2ew1gHBemBWcC8szNgy4sM0alyl
QIGZCtz/AEYh+dtbOrWUOSbhCIJrIqKkgmt+dBt3uU3yNZwWfiuoGHlZtC0IWjIfPJGARwBTWesF
DifMP2k7Qx98wNp5YqFyFkHifIRQzJ1ynHZj/ltE9ajCditQe0nqTV48tb1aRmm/+nseMZPoQjaH
8k3Wgu5y3IoTi0u1oQgTOygOdlqsiZWRSwWM3RLw/rQzDugZ8+XabnY45YWxigCXWZQkADElJ71G
DQ3iGe/bGSK1b7ZHbYwF02NbIb5iZMERrYI9/AFzx4eC7q6QxAcqc3CGZyzpQ8uen0LCXYQCr+kA
V26Jdd1GGPetXqZa/4lZrLCXg7bme2RhI2rtA8QJDvIRogRuBliTmbA0iiPhBOr7MHH+3e9eFfnC
X59nPeybehNXwQIHidJZedt8WJFCkcWElbS2k5AAo6OgU3DL5HlQH83jxrohrcPFwpeYgDiwwNkq
EmwlNgsbgTmu/tqRBMqqACRsNe/v3C9SMcfyW+b6VaetuilxxWqKeYU7D/IKbXJ/u55xd893pj6s
T6tINujvolH/0r9KH4mZVxnrjR32L+2a/CRS+nWTvyv5X1GxEOEWpwdothZ6HbmhcXIKn+b2mkn3
nzOTKptGxH+0OsBDLliANuchLGmQsxB1qPBGPAlW3OZITYzbcKtPrL66lkak1XubcRLgumrbivtx
c8MTRNuo6fLUR89hJ21lKxRDu7sxFPi4Cbej86tYVnkLRplznRHHIdjXX/gkLxok/IxzeM92ZT+W
xqyW+sBbO5h2lo5KFXnR6rUprp+14XWgZWrC7FmSAKkP5T6MRBjEhXfC7BPffBVqL9a2jMLTpF0/
rfZa0M353+SilbT4EacT6PdGW2o4kCyPFKIBXfsv5REVeueqTK9P/mWsWnDwNfIfNXSjrwW/45X5
VI0dIUyhb4E7vvfsHNY4vWEchFQvZen4oWeK4OvewzX1mWBU1svOwrxFB3ceA1K92b/poxKthjo9
8bjDwAEUDGQckvJJ88kjVQ748XCMHWlPVr9ux6OwZXlO89axIPwVRkw3gt0k4zI27qoWNblXTKb/
G4nSaUVtI9RKWkJWXX7a/ZEKbAdK5HkGdvkmTWhdDeeSyoQGRqLqx4/cU5RUNKH8ZQL+mOI27jJj
de09vyDcmLio6opc2wMsPo5dhhWZEQNe94eOomamXNrsZXkniadJsuTXZ7shNSFSc8B5fa9iddvm
CN0h0sByakeEF5YbHz4b7BmANXlGvI0IIlR8+lPBoesexb6Eq+FMaU8U8U9nk8h0ESsJfeqXKYaV
ro+HQlfsjiGajWiml/qhIB+cLg01D+JVz2/Au6IS3yN6CVwlY4jUKQsA/pWysIqxlquYjQwLFhUN
soxqMIkbe4KkF2KqzOvRSDxRcpTHcghnvO1QtJqcgnZAvBNWxLAL9+pCJZsgAeqlO1G1DMYfxWe6
noKjzIM6szVlGjCjf4nEpi8gsoIpSihlRsexopjkdPG41VsnBgypPXt2DL9ETzWa3t3aByzADGw8
FAxajMpJndlqnAs0yi4i8z+M+FbqCL+B4Lgg+srpOCOeXAuPjAm/RM6Ls275cJbeOK2dktlxYZtv
mhxSmWf/vzg5XLzw2bt+L5/6y0DbNI4qHmSS/kLyh1yCAuqbZU46BnZOYvTjfSw/bsC4ddH+OEAh
TJGynsdeKVcHB7prRI1xC2A+I5s/Rlmxx6tEHNl38Fkx4DGPya7rCHj51iK8xFkzdAW2567wIKbe
ZiMQ7QvTUmLmsGCVVe5oazmFhTwBNsOYmbRGhPHncToikxaiqxuHq60OaJ77/4bV0dHdQ+l3/Qlk
s/r0GrMIOiJIpz44lPpY5QLlmzcL4SCDeughfE7Wy3A95xlUnuA3ywHojapsQfEuXyr8BlNt1JOu
GT9a5tb2rP65se3R3PllFQSEF30UA5sZ9MaCGZKEXbGm0rTvzpH/tKYxPlHJjNvZ4IkP3LhZ7AGB
sxOOudqUasoZa4mDcp3m7mgtK0oTYNUDYy0f+j4mKm0QWizIXk2HMZ+xe5UojdEbjPAnRjbNMwK3
8aJ3E3/tw2TGqh+EYwRQ7bT9L8+A4YgOoxGMEqEu28tZ467+m6TWWVyVW5A91tcjRhXn/Uc/7xmL
O24dNxVLqP8zZKkN3oKsMcWjaOBdu4IYtBGPu1y4xNnMx6LIal+B7uh8XGkVBdDVLoHq8IZXn2+Z
5mVpswICKk5YCGMo4L8B6YaoO4HMdQQG64bNewZdkyOz4TgGEcPvR9/5N870JtrHgIEhtt8MNzDb
9Dd+udVWwiqhb2jG5ADqohB6hZyPcWDDfrnXYhxU+h241vtnbrJAGdZfX7MPoOg/SVLnyVhW7N0V
YCRnkYqPl1ETFgAOOh+/oMlp+iOIIBJ7hAP8pHePGgzLF3fuERH0jGJphU+z/b9c+Zd8AC56Uxp7
VYtHhjkLis8Wic9s43JCjHIZQbz4dmGDiVfAiNV7CITcadZQP/krGPlZfPBoJx9rC123jGAqNLHn
BL6XVs2Hz8SX7d1QfIOibf//6ycLYsRpXTnEzAw8c2cnicGM29/0uxGS3Ks4tiDotFdJCt/Av+nu
sBu2bZg4er79M/APWeoZ/0/sHITJ2nmn1jUjaGlJZWD86xHi43rnx9OEO9w9Ak8y8JEcep35f/rB
bL4yeWWhPiSyo3kpQUoiRE2jaYigsImMcSi4wXZ1OBpJMx+3A7yWCRbxea6W9mQdiUJQC1kzSXtp
TM5E8FaMUPMkX9+HbqVhEsE48vtvYnVDJeMb6Ds9lNHMc4DqzYC6UOEcxuekYkVtHCkT+nwbjaXW
bCXthpr3KKj9FUZgsWYJxChq9Fmr1Znxn8WhD8GUJJ2PA9gH3F9Z8tTRygkIT6u5dey8RJKKJtWU
E6s6tg6BmwTHFqHnALhneNHZEdIiB6wpKxIXkuYRovQpBcycYrl2hzeeJ4jaAdv7JF0AU99BNutL
qikFrTpcYxyxmiKGllunX9or01y2f+E8WfiW1eBKv1i1SDzl2MvgYEj8aouNmvfQAwT8e2G7A5kh
DAgoxgHI+I0+OizbLPw8xxwd15SgFAju2lZ9uKqClrNqmig9mdVuoGrRnu8SWx8UhuINV2uM+3Q+
783Afo3TjsUUiv9XUnk6wgAB2tb/N5M7wDjleeHrdm2GzNQsRSrbB6Iq9TdE7b/XKM+Sb8QA3cUA
sAIIpcPFX9c5+zo1g06bv9S22sXEXjp+OalqlEMRWnsYnfKVathcni6vAzcyY6F7k68qA4NpDj6m
0zHDV6OZ8VK7QbWxV1lX+ymSBHcT5e1jdGBwvz1uUbr4vhqvEHz2MlaytKeMIvEJS0VG7i6TEFtB
tFi5wYB5tuFg8NDb1krgZVdyXORIPcM+j121clgGi0KK8QmLvhHZFuJF5Ko/5KzDR4aqWc697IbZ
7PG7gHo65NFYK88ybUNPYVIRREm7Ti/y6+ByHTbPT8mbfD5FGmgrRHMkHY2OQpB/6rKfWzq0VmJE
569i6Xbbj/WW7Un0CTiqU9Dfwah2KEmPaWU1bMKd85xPbUgeCRVY4uTOFg4rwcBEgIoo9TlEkDKK
px8rfS1EfnyAldAhlvUTVlxLB7XdB1Lr2lTLKR1a885iN3a+NIeCAu2ETgfPJgqfRvIza33irLU2
K7FjWjvMTzLYgTMiQZAOKwOv4fliLeeelWW4X5StCSi7bReimFQ7qy7vpAeqjyP2UkSlQlPgUx0J
7V7SqvzbwxliZx4i68wUOJNwvJbseFzp2AXh8G8xHoqQ8wyvfsP3kg1jtLy1oTs+bVT/UCTYfGfI
1wu6ZJN/6zfeSoA0RXwRslCj8DP2ySyd7JdgWkm39FYQcKrz7cFwQZ3opKA2gxAcrvLaTymL32da
YbNVKyf6uINFXrmlLP8nT2c6JjGO+g5s7h1X3CggEZrUagfJ+Itv0ETxWFmGdftS7tDiLAdULpFT
JOppUz17zRqofzz1w01KS3OCYUl8K7qm8aP/Hq8c12CYMYfbS2EnS6wzYTlTUK84vuVcYDNQsOJf
EHPiAch4oQ8jkfP23S41Q2yhQ+BY1bRxM3bQSyr5DVFY5S/1HIStp4gS388seYgLEKnMt7eaD9J7
zzmcFYOb3nd5VmM0rllUZ2t1lMUWKIuu7I19it1tpbinj3/ZeO/EA5fRsU+haaRfyIi5cwZ7Qzf3
HpBiOonp6nbRP2ClwHyAHH46zEJh3GmzYnKmuxpevQ86eo40sw+/M+G04e8BIcMm3nXvP1YiY2hG
7e7y33+UxiZUwvhcidGDJf8nIdI99t7hMjKpbFmW83mF1CZMl0wTGUYQg0mbUaoyD/PAgP0yi08W
WYxNILzZHamsYKA0Tc5uXJ7XqwHyJ0WL4wFdDGOMfLlh4bfikjxw0VDuZSo5P8q6vRHEwBgQgHJB
Q2XVSBj6WuqQxFsKMx4CrgcstfYS59irgrKdgBjfSUYvKH1z1mD1FDCXJeM1QD5Asj2dO0r2W+6P
loLStehVs2umsOP/UCTci7IJGlVFbrVW7IgCSyMb18F1iWEMLG3tCUhSqs+luKNqgnFcf3rqcx0H
NYfDATFUAmYpYCneZ1g7UotVLYfhUSz/IF8hYiVr8C9onY36ksOlTQiIfVMPhyO+vh0sS9QKPFNx
adCCwM0DCP9mUO1owRIQSztx79eE5gZs9wrrl4r/eZsoz842LXieZgG9UTpXNq/kB6SC5uw1mOEJ
MbgWEO0Su8DoOH7uWbGOYv3f5lfdnHKrL6VE4CrF7Vqd578p0wzNN3m37RrVbYGZsK2U1V52WstQ
U1oAOiW2Hkvzv65wf9Jge36caJg3GDBEAaU7kQfM3y6oyKrlmHJMzdzfRS736W1rP3L4JtzZeglN
RrdM6KcMYYSQ9igHPO9jGIc9b2VpminwPqaCzzpLjsax14v28Ex/XP66qfvd3pbLd/igpsGbZ38q
1z9QiRwNMAIiWBTysdgv3qLHuLO1U0YwGb5430j2JY32YE8SepCYdQ385L2CNGjjOV3O2b9qvjha
Do7Xl9Bhg/G3viCO5GOYh91FCOYHxm2nwzrFndwc/Uyct6g8QukBlh7Lh6T+a15zDtfHx2U7Nb85
RpHOFcNBNNvZcdq8vF7BKsXgseKZV0Rwu1aZHBbJsZS1NM5IgyzjkTSjZt23W49B/PONg5XnNH2y
kWcLufP+ICa1Ihu7pyvOo4dQVNlW7E4ULyxRQWWb3BQKVhB9oVVknAe08idWQgd2nUbDDnOa0qhu
zjEFkMkmMlP6TltTyPeVXwE4AHsu8gEjethU6xrU7uVkgpC4bDPSTdgMDVyB+QA4kHoImXDDO7Dm
bqJyzKY3nxG/C9/pZrNGmX0As8W4IE+N+ZG67RAh4Z9jXjsIb8VMbspSzaOXdEFaiuA9x/B+6v4y
GgtMA8LQSws+5OKHRxXdF2iXKvPgGUVncWE+CJoYSH5QG+lm6kwb1fbmFKQk6lndzWFFAMRe1rt5
lGOL4ATQnPegV5uie2og0VYiokioIPkRQiBocLtPweoMipqhi+0OL2OerRnyCI4x3iZv93Cf4FWP
95j5qlc9zSZ6YB5UI0HLvGGGLtzEsoXCtdxBFCgsY8xSsJXs8sccg6+O4hu258s2tHCnpV8/BK5t
1+Beylrk0dvdJCYawkN1f6D6yozjfuuGQZvdJMkOBGENodo4e5cxlK3yRwX8cZWEQnJllIo7ZsvD
ETFEtt6FAYhh3qiO9mxA9SgM7BvpzThVYoa6SwusNlXWrX5A8hcBGjlknpSxJgFiiKcgiCFQNQGz
zFw3O+LJp45gDzE3WEd6RNRxYWtIllOR0hm9rzVxNZGVqmUXId273YZYjL4OG2HVDpHUBiNM5pe/
zHU5ZtzWfWwx8y+8nESFWUheR4G0r02BnhHatdL97oPMhI9TfHu3AGrd0UsuvMt2s+wGSfC0tgaQ
LubNQcGRplVt9SNMoFsEAxaNgJAlHhnByPUeL4aEJiyJPSLEChluslSGLWOkbZxHnbzf4cMQDusc
16TO+uKp3+tS6gMknLDxGlzgHKZ/lSC7ffNrQlVmtajN4LPrSVGRa2VekXVwUZIq4qKlcQfR48zN
ww3FVOoqQHrvciNsF4yH3ewWbmIg1Q8p6nXjzHmNmkzppU69/90mrk+B28iNt4wiUmbtgd8WuqjN
1/ZyVXgVyXtsdsUUTw84ZykJ6a55fu0LncRVSu8pINbLLcUAqjBK8+WqL8uNQrUE1n9dCBCNI/hk
UX0bbbhymfBgROwANW+GcPwCmNuVIUTtI/BeG2hSqiD9GNZTOeGg+OOmcDGOje1uxrHO4G+uOjVu
yQy/dpZTeTKALzRzYXqBnuzbCrBFMer6orUy7u3DFeDeka0dWyXPZpm6PhOTesrK6yXTnmK/OZBx
yiSBknISDtH626LB2+HxKUAIhQ9OTJuV/jZOaL7f3nIPG0sCXIuVfmQrPJ5Jg2vvUtBzFZAdXqrf
KEFA0swcFWZp3oulPo84VMqj7ZedbtTzN/JCOWPSKY2wZNuLIg1TvQMPWrVWTQIs5eyZeIHI0Jln
V+MmxsZaRZhWAKhUhcykbZ22IQ+dZzUli1AETHB2Nhmt9WIAP06ljbHZbclCz5MUgolLjJNrvA+b
mXIJFu2NANHTBvVRM37/5GVS8AUTNXfy5WOxN+eaPbWwt8cBTfQrmdy6Gmy5qbpwNnzx/zjg9Kpa
EHhLc1HpZrfeWemK4wn3XKthZuCpVWT8vRjFPb1qtKBl2Sad7PavQFJItocOW7mXossA337AAPYI
RcbbLDMnUPU9whA2qtKJn6soU2dlFmMjNdPXXdH+iggXr9r+D8qPMdyMXH/R+AQf5edHi3TXvnsz
DcLfGNr/s0v7tioaInOVVG3NoT/8AZrPM77upJKH5lQCOSg5tSMYIOkU5caC34k2fAjscEBTNNoM
BXVulHRK7He7BZInA7imFx5BK1RUY2PhDyPVWuq+Q8uyw+iwlx7g3oz4AtjEKyHGIRgHBR6f5BFr
ZRApvsOsHwYgP+SUL5AhkeQSNjO42HQiR67ybXgNjxqH+sNjlBr7oyG4wpVixGc1SuS+ygq8HTfc
LsD8H1chlnKeVBRV29v0XQ8bOoj4YyvdyAkZAffQc3QLeFPnZ8uRgvcfvZFb3djK21MeuR4YMHO+
quAvxwUpBGxcoHvJm+DKEYsOhJ+gZlsCnT6+JvmO1mEx+ra0LdFTJAhRw52nzgbwq++SPZSh8JhE
6yOjRCukNd58oZVuNVhASV6a+2R9Wt7GnwlTekSeqRV+7KJosmawMAu2S++0Uro6wP6PBTDka9+s
V5RK7CXahxD6qxKMMB460NV2U7hoUmkP5aAiZHEs7g3x0+PNtdFZWroUU5QNZQniEmLDXd/0pqzH
ep7WhdmtiQIRzfm5OIPZ/REJ30TSiXbKaR23FMGs5KnpWrv7HObc0gKQL9TQ7XhoT0kxWUMtfyH4
Zmqqb0wa4aZO4orYx07KqWCz9K3hnasYNMDlzY6B4/aHxIpgI4kBZKL3f5/i1o7rW0g9tpYsGSuK
8djpFaSvLUb8gDasyc87cTTEuh4brLmdVAvsKHrdnwvo3r4KsmA8bnXC5SB2G44qMUdnj7c82Fpm
BaQ0rgjtfptJZP3ziiG1Ovi5uUeBNDLalcMN7rLJNKyWmhxjOBqYBW0G0XVlD4ChSlwQ+aMLAIoa
qeuHgBc379O7tPq7AoeaRBz7uOl6Ind2RrSvi8d6VwXLDDBjjgOV4dwJUVPRRsx1TCTL8BrzeFhS
SZ7jZOKAqbrND4mSJB1Zk1Vga2JbSwxlMzQcbE/A9qNZ2i7sdbuGWGmaZJM6Qbxldajpo+EfXgQQ
NfZb5Glrk5TocO9lJN7vfFpK3fBOHipfJ4kPuxFepRT1kU1C0c3l/iRxg7l/jxi7+HicJT1y3MkD
0qZI8SGHrocUwDMC0IWLPFR2p9Vg2TRPHmBIDcHhsUoRSLr66NfUF+Ks/W2sLFzRO+qmoVUHT4LE
a3jsOf0EAamgWX5X83OK4N975UM16NTy/zG7id8niY+kfUMDQVJdB9ZspL05/yG1iMdTSbve34Rd
ZRX7Oeq2nrcCMxkSLLXecjYM9HJC/r7P2mzOW1EkQi7i9BYWg679Q1Za3soL8gohAEyn8EICiIdb
VuSO8SRSON7nI9zunh91+QqY+uCsLMFw8GYA+xymMZcDHnrMv74WRiKAnOwVX16ZHLCN6vIGE5dg
8qCWNL3erDEVRTMGoAMJ1X0j7zpN3B11N8G/gMjzjOL0woi80kKsa/JKhUbUauHwdD56VBfXq0qe
AJaTKr+a0eZ0RrUezosvb+W/Z8t0dx21zr5KMAZD4M+7zZdf2wvhKXDjMO2kVCUcbG5DDyB0FuUe
VLOjhZS5+BFnHnrdcW8NO1Lygp5xpXZkaX+kgFQwbrYW40CeADfJKqLYzWLY82TjhoXdmLJ7ZSJB
dmswY1KrnYKwK3BLOrHQaai2PjGWkjZTHMi9XfX21hm7fW/K2BTrMcj7EzRH7N1ru5u/R0+BcNPD
f9VV0YeSdY8GWQqRAO9Olr4/TOCKFWieY6gVMAUf5kbd3/zCS3B04AHanMndpky17/qv3Hh6Up8G
REny7trFEJCCnQ5el3Uf75I+rFBJ8iJcGAORswuZh5vCrq/t0Tje9tTdz2wfN42CYKL05JyWKMop
Ua+dGTSu76ApLx9YFwHaRFLBKRH0GA3ZRxvuAu6y2fR0nonRw7fkn37GjNLUz0TDBQXpIIwIlsuD
CPzfuvrkSdyVXauTfd5EVvcuBqRnrfVqCTDqXteTN2IvcH9KS/84xoKKe+SVfyUl46vMpnT59mFj
vQs5e88yMrVDq4XdoJGfaRjezddH3KeA1jFWW4cBkKO3xfFCOqkABQ+rvzBomRuOa5H2eB5TNt93
c38dLYufUEdMJDkSSniG0FU+kWXFIEUer6X6qWzE9+GQW9DexRBl0k4F7rHfk3k+OVgHME4DOTeT
UV1Cwks0mIOeenYatOEb8G6za5dZgv9NfZnPQuMIT6Fins7ghYJLOy8zpqE5/MTOR9oAg87EFZ5x
tlr6vNpDT9TVIk0sUN1OI/ZFMSs4+7Fx6IctOr01DXzDRF2KJzDceQ0G3vo7A8Ekvy+KQc7wL3gV
qLOBqp3e3Gd5XcktNHAeNCEcZo2mb/jUNFqnhTYjH6nOFjx8YPM0qOLQehSxxmvuTQvHAYRKIpiC
PyW9W3mSOzCMUDYWIvEtV4W7bkW6Kn24PXMMQHJOh/Aq99U0iDQlmqBpo88IzneIfnJoQ6e+PLVT
jDQAX/XBoPWd4yzIO0lmMJNuYBYyLl6ov4B87+49a63T81PjYvihDdY3cgTYmYx5rFgbvVW8u3Wd
LcsHIG9jDqsywx+rLb+7TCRbwlyjnSYeDwq/uG4FxuSQI3KXnSeJZCbSv/ZlTAlYRL2sCmVSY9O4
wBortd7NIqEr7JwEHHo5anUi9g6w+5C6EjVO32r5fSo0AqHRcNKGZWXK31qZkSKbKAh/LFSWdBsF
dSIWsIUvZ7OqhnNdaVaYILpo2szBp/ktcWrGGpeW2g60JyYeR1spjTrGrmehuUu5PDZ2WqJ5i3Lf
jA0H/2qD2h08nk+xMAJzQCRp3IMwN+O1dh00gkHDWp1GrRcqdLhQyNVlrWyGCS8dGfxSzQLstsnr
Yvjcvw7JPiW5sWshhDHPSLecerv8jdJgZTeRxUMhUDNW7jSxs/XdNuYKqd3PGC4tLSVyQYdNBSfL
OFWPIswCtt7hF/GBJ0rjk4pqxAWzcPXuPKsekGbHnyp5EWCepPMkUB2zaYI4OVUIsYX8dhIiIj2O
gKQ/3J2KGvgDGY5xjR0EGO2qGncznNuYmBZgtXgZldMeofOefKspDBWuKYfsTR+EIZAo9lsyM3MG
wtlXXmviF2WnV3isgAj1Y/gGHYMzCMEbVo9KNzCKntL3Nh1clLyBYnLWOR26MY6I/+TSMUqP0CLW
zNlpYbIqzkOMKXgLj8qBMerxLSm5JfvEsEldhLZJSpTWtmnEkSfysZ9DTg1966xsDZCwrvV9SIeb
AqwBTIlq5Vf1YEpvsalhAoidn4Oo9y1oeoiw0IPUUiLTrgPQORozdsdj7mLSvDpNmG/+t7UCY3AP
od4PFmEwGrgYtgQt5yjtB+Krwkiyo4HDMye720pXQpp/zBY5MgpLuRohpcoupjUDxn5iQt4FuVdy
tTFo0lOyanvlcClGNACdCQPVaAHzRYdkrh1FbE2jOWB/jIdLfxuPRGpifPChr0JfQlH4zxDwTNWe
HP8tODmz/LCT2I6fdTJP2i/apoYE2pRyOZq3v45M3f5S7KqDPMhk9m/SSz0Mvtrzmu1cvvNEEUOW
Uw8+zs2FVpUt60xSKDFP0nRsSmBnTnUzeUJF9bZNaDxFoiczdxBFp0hBNHlG3v7tLNj8ZScCKZ5u
1TjCH2peFe+1exVo19TOCZe+k5ZfKZFKjv1ZCQp+U1qrHDxf4e+c0fQaNjC8c1M1ZKqLm5CGG6sk
npTON+Rix2NEZSCR/8fxlekqmtJ+aH5d07Ubg6xcWeKxnjJ9Nqx4rBI05fEi5OhAwEeDn/hnWopL
zmBO1zO4M8IvJBLclT5hHim+r0OOrxsRatgos/X3Ygylq7nN16DoZW7cSWL7nryWfDQx+4rntP/Y
2SjF6HyDvCI6Z07kTw7jWBEDvvwSEzw5qilu6Oe1/InEAMX0IplV4KfSXsr4IDl0HlLlYw41sHTa
aMt6E3iJMqYY6SbsS9FCPe3DQpShQtvH2e4G2B5l/h120zsMV4gPBJYupfFDPILcrTWaNQGlHrQp
x8apKjApIFJ5UESqqblzkV/cBDyhBu4g7wFp53o5DzDxauYNIWJemDpaoUAdRdHr+iKqPtFtl4YS
gxxX59AubRierlcPhewCiGD/Pbi9jIGQyM5m0VK0rw54NYBMnJs9aXecULGcg7/Cq0/SZo+XGciQ
6XVAspCyEeQNnaJUhrzju706rgzZwsp+WXfHSgyk2KYYSrTqNG/WPv3cWsHwSYo1G/kzzNMEV+zI
lu/nMTcqeZAptqF+C+thsKuR/K5RMkTMOJGxkYRRVoN19QoaeEvalh+6hkKAy0Wo8219qFr32k0X
jwsFdlRbVGHfY5Q0kU43aW827f5pHdWM8ynv+IKF4dameSp2e2vorlJAdDwGlHgyk63Vgf/dZ2qz
3RUHtm2EAlHffFMXxecGIM3fUoHfQ6MplmKBq1Ob3L3NFvvnuP8Wf2t3qyNeITGVFPemq+5awA1G
fOv+cO6qdExwasyff6yK9TvbUlgNSg0oiFA09T3xrfMKO22eHnz/49tL46Tw5setoJvPhZIP6B8O
MNxzmqKL2J9GmfUtoUVEnALqs8PVeoU+GOd5rG1UtH6bWoYYW2bDo5dtEfGxWaob+DGjwrYoTA78
YcznPm8Yn+W2exafFIsZ97a/AZ0IY8nzS+LXPXv3AobgT7gE1APTzgo6luB4pKOBhWa9ciH+IAvE
oqe697cGG3qAJUqf42VJ9SdkPqeuOzz1p5UkcaWObjQ20lvjvMG8fZcy5oAESDbmWG/7i22zGOcU
SVnlFt45GJzDrMP+n6PYtFPN5IBtQeMErYDCP7zwq7PYayZuIj0L5cVEuz90sfH2WRgWd8v548Y9
6dGXYeLNmG6eNGR/6gVDCd/HeriAZHCRErVHD8oEvq4AGvOlyEcDHg7Fs53larZRW4BDoCGLh+L5
+HmAgpcfe8MOJOAK+HCOfVwtao1DxqjaZHBb7wofiPlTPGN8l0zZ/YXj8IxD0ynM8WPaIMXOfHqN
fUVYPHMCaEOrIIIoHiP6DFdgYJATZnj7Uf/cJJlhUTTYn9mEFZ4S6sa9KLCYMVkkKUozcAkLleEk
+LTw/+fFzsDpU9M/MgbvkLZqXvJ11UPSvYeqPHVNC4kenmq3Fta2sy4PCubWGE8lz9V/4wzf0hf4
ed2Lj2Hnjq9i9u0RVtgl9BZAQY2JNCvbKOMRHRnudiKq50ointPTHI8AmItGuPIAPP8UJA4VOGjR
v7i6HEfkEBFoIuRQhPcOE/hCBC2AAzGqG/ldgK0xLtTZxC0K3+roXWb6c4146zgvCn3SzgUxszql
Nlw5ZQJ+xOxTgdG+Idp9HXfSkStYi5P51v420f03lt/0IDll9yAUZdBULXdSN6qEPbDYFutuKd/P
aiqtQ3qKiIYZGFKhvk/KSent5Se6SiEmqblcBPnOgBIEZPS72hnKQX8QGVsJwRlPV2opW5Eyrowt
OtrKgbjEmecRIOgHsyLpGMCzHqqtMGTctodHaOT8PnivT83grvQ7cGU+tBUJ5OcJrAfOxHEzL5om
uO9vX2CjgUE9dHoF5C7q1swnQftdKEZryErABAqxjebAch7W6GVYvUnqIQNzS1tNe1Rp89WR3dPL
YGpSA5Eq8zfM9y4wUDWGLcgjR66Q0lq3mP8kQj365l8Jvtovz/rBLKCbnjjpyplSIKkbjKNeo+NN
uzpPMpwP8jknxnE0wgVhdMG4WbKlyzS+Ajkiv/ayQUGhNwaYk53bvLnoMcMZWILI0aRu7gBXFYAa
HkqdMnWGmfua80gX28fJle/9p84pRqKNO67vdAMfsPBZhemL3SQsHnuv5B02f6CDHce9qBUiriut
bXigo5yE9HbcXByonPprLmY6EVKEEaFrbfqMX2cyeAcARCUdvm1ZXHaHeih9eGj31dKt2FFJGSPM
c6pIxoA3JvFBpOSZCC8GheBt+PhIcS2+equWsvhYm3SrYNlY+4w9jSZyZTfcisiVEHGz2EASdJmI
UTcC3BcYQK60lV25jWAaAYvEeUISsEMasBRr8U8/jBHwvThmDOmrMLQ3VkmVtLCaAkrs7e/tnwuf
6HLIpTcJzohR0cBUSwcMc4UggdiYuKdcG4tnZiIwXuWLtyCdUeUCBG6b07LUZIPrmtMgbBd/6WdP
VpKVbwvffeF5ZHJzCASJhWTmm9oJYnNuCoQl7Dnpwhyh73eMG0fw64Ntx+KjhnVaVDMjyOV18jIq
vOUykynB/za/zjybeXKAt6XZMXnD7k8qe19dF9sgJhLXXKSfGkwCfvDO2VwqBEEBkIIdO78/5l3A
kkW7nV5nir9FcEyhLClXFUVfYDtQxzanlmU7G3U3DIINf2p9nmycJgQ4N/tRhpGk0OrZgtNMnj9B
DaqDB9wgzH+mwj5oUPPDHrINj6i87sY0uJ+Jwx7fLzAMC6nuegkkhTFhChwypMBb9mlSjFUtTVF/
hS2M5mS81L9PAS0bbEsIDM8NOoAcCPPqi6jN4kdsvlJWdJSH87iUZ9IrFnqvcf1m0wsMUl7R1DXp
beMIEpTxD9W2XuWOoRmLBwcP/RXKHzk60QZNqKzpvzUkQqaq2MbH06k2HxJfFjmtEEDIVP1IIDFa
QNrw4A3cDVRwZ4XQ9ONJ4C5Ujf/f5/FaN/dK9crFyl3b0V6Tct/UxvRysKtE5g7AXf/57Es0A8St
qD+21cCm7fP42AZniqjLvXS8Ji02B9f8yHGtGIqcM87V6b6nySWYOeDRde3G5YohvPVpRdBGiDs8
ZGaeIXnItR+mo4Vx5tRewETTGKcetMgRXHvyOm4P60K+wuobUKs5Ubqiahg6lJDPFb+hY3vZ0r3V
B0tIRI/S9tLHrVeMYqG660GR/5aas8jVJEcJE5mjGB+xR4E8+ceFU1qvzWUswN/WGlWPv8hwN9mK
zjZ9eqQD4FmnOTjp463okLbDIqpSI4BMuawNddQQ0F6HNz8aofg8W3sTsAlanbnAp2vTOyl/Q5JM
q/24GlnpJ8Djg1z3UerbsxCqxInr0G0xUoQSzR94+bUbcP02jZuCxDsUkWCTERHBwxHXI9w+ckmd
jLkCheuDghqHbpGdPxCYzLe2pwl+SeAUwGGAanj8T1y8IYwEh6FgHdOqDl7KU7EpU8m+zUeLKe7c
JmOob3Ty9OdSWJI5ixrOcapXeBT0ps8CRCbPM7hkjfpPzwl23qTZLeDrcVbgmcLLG5ArkIDC9/Dh
/Hz+ZDMg5HkLTRXrLalxp+gC9ej4b6WBokCmRSFXtGrh7O3tP6K1295Of5Z7qMfoP3SBMYpTtRFP
OmU5wyHnaLKV+j7cGRrIG66KnwMh7Mm++syFnQ7Orq2kBmp5GIH0EqvozsobD/OxyPAvWLl4elGR
pFNWM8gKBeQP4ghDv/e8RYm0Qa3HKc8PfCvGD3CokmBtHXJDf6f74flMF8b7kjw4Wfbj4XOIpgli
N4kIe4NErwIGi/zLv/zTNBuWbzRNCWHKzjVZkrLENNVEhgk1Gp9oTqDUR0vx1KtC0W0Ohqx/Mvu6
UaZ292Q/iale6EyesYo/KHp+x94LS2gor93tv88cAIG368sRWjIMBtZI6nSWZ2V1Ta/ZiXLj3yVY
0dUnHsBGZbSmXKPaSweo58zFYnBGQXQTjY05G3VpYJJN6Rv15syb2n5pUB7bYP8FePE+/n4wXusI
KJd3Shvf+DuUkamq2MmNkEMQ6t147IZMuM18Sdh/7gs3SStf43IzOoZ4Unr0HjdHPlnuPUpxmoBe
dRlR5rCzGZe5t/nN6GCyqFS/ph1fUMXgCONLQx0pG6j+/w3soC75++4bqQAdAjlAyB9b06EdwlBZ
nsgOOa0YPWFqfXdqTY/lf1YGoziDqXwm+xG85ZKXEAV4LLH7i85fT488xPfiWNTEVj+UN/d8tHmi
+kSnWs5BOlAYj35urCKTRG5SXY7sCwTDITOhVUJbwdqk81qAs6B78DZUbqe0lRW/Wex6XCL6RNvk
5HCPh+G0lU9eYv4Fcmhm9Rk7iWk1cy+gv3hb7jMpK5X1VXKA2kaDbJM2N78HNs62j8OUz3gF4QAm
yvD5UYsOSXW8mNMQdFBsxLwQiJVSfaqAUITtKVjuWLOf1j6X/vQxl4NW1vYrSJX5rXyP14DLuWuH
Bdew28WWkaK96UQfDJWJMKRU0+TdnstppHPzmNwbLdHAxo/vq9yob5gqW0s4ogwGVTg4jE/Vsjcb
I+QceGi8jb25D5Xe7Asgp3pGBWlKyFCHeibia6qWKuz/zQ5PBQLHCO0w45pHjq3Lh6zGXUC+hwex
wgORtsQrCVT/dB0OXmv1xEgHJaUsO31rgXH14wy08SsP3HfuAliMOfPcR5PEJFvVCL6EdWcsrsyV
/HX8ijhLOPZ0DlAv2cx0x6H8/CBS0tW9LK8+yuZMvXjoyvmdg8dmvaFMkB01r8n2DulfLWY9Flb+
YpTXAEpqTcWmDfNT8VcVsQoR3eEaKS/2Mf6Pn+jKwWp7xTq+CBZoyNnAQ8YyQMpfPwWOkDSaYVUg
tbtcO+aikt9CVA2WnSGqnwWKMWYq4qkiqHT9bXndLQogLlhUoHGoH/1gzyr+To6nk+/Ha21wQdu7
wEpbH4s5H6hBNGonBagDp8UC2rYTwoGMt/piHqOOgX35pbJR69ecQC5yrOF2p7XgTGbD9QZtJxIz
0dIyarmTFYKi+1FHwVQcwn5HRJ9DUnRcEFo94DvHzKOEVipmazjPJmdbxd8ryQSYF44YM4UxRK8+
odtSygxS1NbFmdOwxAyegijiNdyFHmmM5tpMsr0q8ouhc98jlbN372tcSpvRLkrn+QfScw8OsuaY
da/rTlO4D2NxbDGc2+nYnaGyGui+JKGZWNSBSfrGiDVLYbS3NEvdh14VfV06NMwxYiqD9x5VN1e7
HTiog1Rl81+JZ7Sy5z2b80iN6m3L9b9UHTiybdSeIg3NFdK2lei/7diEpuTEPrie3rlrO/c6es39
N1ubguTiMj8zN4C51X4fVDlW2k2EjIF1R1fZ4heO/zEPLKlZ7V6RptAgz7Gfykd8ODSTf4YD73sh
idmgXe5T0e6QXNupXHHyGmWN6BNxWuX+rK2NRMoebkOoChNrlAdPTPXGwq4laxPQ8xsHRDjFTeoa
CtIvZvbPKX4QIDVUdXyTtdM/0NbQ3cseBN0pLjekq8xOjX+QFkoHNcnm/d6xanTnfMfFsNYEJwX+
giVd28iLM761qxKAJjTAeRvjdRJakDlFXAhmi5WbCUSxXIMij4nWQPHQXG8mnA/cT7F6Dxay9V8B
jUOLxsUHQAUudKdC1w9jDUQv4dekWWXc+dRaW2m78YUaIGiWKXnd36Br3OiDz86TcWftvuIWGWYP
E4v3tVEvDrm3XQ0KpZXvvS9OYSmnMZGzPQlSwdfn4CcZksEwqcht/7hSlW9yOCNNVRc0GQT1Vy0Q
yVKw/gBYTW6e1dZHIvPPohdRn8kWEMTQWohUgSpXN7ZKF8Gz/eaHiTGN+tCaWhWxCbMDvsw/dHoF
WhhBovxpYSAGoUp+JMm71llP4J1Ick766lgHWlhx+XuEtHKve5/Wgiq7wDupoiv1Uotst6+4c4Rt
qFXnn0rfEN0cboOGQH0FK5ZNKhtdAiid0iKbySCLdHWCvudNELdym8wYvbK/u+bFfoFjY3F349lA
oTJTZpubEX/KxLLYNKSxynqMTTbZWiyTKfvgXWBVo4G51Xfc3BPgPnVG/+gfM0af3Ml7dCHaPeAl
ckiadQpemx9IhP5O3z3y53eEwGhNoCmE+LmLd/zsTuSqiVFigt3MoGc3Mceuwl0WMlJazFQtJo05
Mfg1r6vDjwW33ZnVHA1Dl3IOjiIUCtvQKcUdh5w2+SKzOoP16ZjlJSr8mV/32hVEYdXwItLVhH6T
BZkgpSyhJims0vyIwAH8xS3AdTGenZ5kJpe2BxOH04SKTivFunNF6cLVwPe02wASxCbYg2A7rsd4
pAvh11OGG4vQIo8N9IXze2TNbuhSaMvM1GOHhNLR0PupWRHGbOGkkaYBPzdXLeJ7bpCWlGCF98QU
XtiRVFqG6NVHKt/0MdeI10TjOYVdPJUvVkK/XfykIr3gTpmGxE5a+8tf7/9ov55Szftr++DZ+PEO
D+8rJ1amn/aw/cSIC5E+6qFx0836qQMbYEkbH0Q/ImxrRHCymOUG3okXpYsbVRyd7zk8cifA0XRw
Z0KAxxlF8B7KUIxvQ1rKwQCDnr7IY1SeWCwbPgH99m2sr26QDTSh/xw97LsvtjecI6AHkxgmildV
YduePkvLkM2Uti0pAUTBsZIdwSo6771zqxCIWQfKZkZnaDFRjMBFd7/wFXN6DyxL9v32jUcxJmY4
mmkIYnxLUiknMbY5F6074ZrZ78soMmDpD9xEfdSkTmG/KX4LxJ61xavSoluxwjfQgjb+oKKWtihP
6KpvCLLuziHHqu5WUoBtrrVeik1md8rElXX7s9prChDCTZtX8UVxqomOI5Yed2sUsdDaUiMfnhOJ
nNsHI3pYaud5HjyZ9f55kE5qf7YgKCl1zYF99RhtzIMa10vEtxpYPNfbMYrCzeNYcvFnZ0iTFp9+
VTe9Lk0KVgoJmmMSFJ3+53Ck/E7UbKloUYVUpJb7/bQT+KYTp/gxTKgHKWwTz8EfOdxppIqo5/og
JUeC7VRW9BS5YQ7T4yqryOwrKrDmvGfyFnsF6bFpnTV7Rpgs5rdzDnwGsW1bb9Khtfk1a+7aGKbJ
yN4YOCuSK6eiB3/kiCqwV392H+b4uBZ9WnVbAUdTXEm49h56Cp653KlauGhLEOvsGQzwtkG1kHk7
pk0lqW+1zo5cLLzYCxREc8Kfk5UQ5ZqNVUi6OFWdyYYyI089+7leE1Y1bcNrS9t28RgSGkEbJyxo
pgAx5lgNCzTmo53mLgF21ro7zJQFjmEvjSSBaRlhPvfSe3Ni/u//p8NjMxgUnI7p4ZR5N2cF5GwV
vdl3yVz05KX1xxPVyj6WiDuU9JbmoWwpVc/TlcIal4sbavlq1UrKMU80DNdNX0hB8wfUcjrktX4c
H7wfKvhig+WdTAtylW9Ilxi7GmuOyeb/+DyJV/EgH0TOe9Y/qYpDjURlB+lJMsZ3S9DiXNrkyskL
1Bi2nqjAYhyxrzbPIHpf9Y1DbI0Z0qemO35DnjE+fMoKiEt9WmWuCRkUQyYZdKTR7Js2dQw/zAra
LvGZ303FaFa0I6cuP/t23+Nzx+JTQMxz0C//7xZH9wLKTQW8+7cZBBl7zEz25wz9yBLfNBsGQRja
pnJzto29RmCNpX0e0sAfq32g0bKXxgoIcMU5uKpRjKnAo9LuQ2m0V8NRPzj2XleAOLA0+2YEi3jV
1/NCuRwZop0FpfP/ygkuCgcX5MehsBM4ZFB4Y4IG92cleFchCMD24o2P6SpUHgMpZFZcKQjx5RLS
GkKa0WzRJEQX+F1Lu9TNjLG6bw/pSvdX1eP18w7dU82uOtgutISR4RgiuOVhbMUUYgNPHtXLienO
pLiDSLr1a7D5QueEX1zuEVxpfY4FGsHpM4qpwEmf/7YRm/eX+D416IOR7r75BDc9ueJHneojeoFo
Iu5JVcHtZaYrbz75XUjK8T4EKKlPDH5hUfcXys8solHXJLnpOgtUu/+QYbBCwr0MGm+xb0jL7S6P
uwKNXuNDpEhlaUnzwY7/FQPGg1zN28Q1YJUDZDm58rQ3r1s/BVqnQgcVfs2+RVzZHWGM7LradeiB
gwaNsQUlCOEqORiTQxNrqA9A3TxpeoSH6z5MdVyg9QK5p/4yph4ZsVE147PtzTHnF4glSFxJ3E+A
RkVgqH4sJ6ECLJXe/lQetMhZYJ1eMCjFhqLj9GcoiZg//ErBpcOVf8d3UF66GByEFqfhD2WCzRxJ
8N/59ERO6x5BbOfw5RGwUivN16DPoM9UNXrxvETJsYSTVwG3bLjjdDJLAPcQ2V/VgLMa6rWlV8Cp
aISgoLZ2BArKqLwLr8C50cHGDkHPaI2XSjGpAw2uaE1r85H6ZIjKbjp4JaB52QOMx6/MwavF+dmi
XGvWg+5ksVPUdDBWkxKaP8bJr8HnuuYSqK/Lf7KnFfItqeQgXzZY3dmYYIU5LBUPGxnB5rjCkTMi
iggAamxFGVcL1gwJR7DIfJUHjFE3An80gK+O0+sQ1+tkvknEg7MCDc2ZqGFuZ0/G5QfwTbbF7i41
JR7l7khXeFNozTk+gxJSmIC5wyhnWbTD9bB6DNVHZ2FSVKKW8FQxIbzPYrqAsZtCnRGVKSsoBFqU
XWF0e9sShD73t/he4eV0T6efc8zMUIiGBFu0LG0w6nEO/uD3DFYu+XSXC4M7Ol5Tk5PBRgniTIi6
rYtDyIhh68tcDmjIShy4Ex0wqHYvpf1DGlaCfkVnQ5XIab3GrfRf+3h5ukAXOvI5dK355EmHJ2+M
bSHqrSM5QV8xb5tY/GcJ62uCktmG2LF/gVu6ZqItRbul2zsQCWqRwfM5bGTjV8jKmNxVZXd+/xKW
xhjOzZfJ56/Tm9qfJUtgAy4e0m3IhfyzMFrsUZOT6O4pbvB9+F2PkbVpcPdicim8P0NDgK+Zzii6
eUJ6pa9Z1pBKJ/4yCczrQdQXCFqtmuhc9hZY5RLEXnNTDwcpK//DZTrHf3T8sBQZyAcna4bnzOqb
I1NXO0SQ8VKL91nD2yIVfRmomdyQ8pvRDpTyvNL2jHtQykVXCOypWP6rcpYd23UhyTU7SDD1kLdC
ClmYvTsDvnvL1EJc58HNBxVHbsKwSSSTv/38Vh436/d3OTgc7lTH2hnddUpJEkoLAxZIqFInB1zB
E1yUhW1kfO7VG88JPZ4XY07eVZc2ofNUv5RpCrVS/GlCpEavB9sA7ugz3ICA4i8cdJY9OtdLs1hg
Yw42dpXvv7lHiVPP6B3FLGk6Ty3S9X64bacdJObtb5tDNB9Wb5jQt4eW11du1xXS/LSxCu6UaAXG
ERm6tAuYbafgTRnyozZ4JD6VnvJt/OD4jV4YltY2LhUz/SRuszIk/QvCLxGa99n0QvV4I4GAC93W
rKRoomjHeptlprt+/AyQ6eH5xWmqknhGE/XFtwG+2AglUvf3GFQFlb3cRrpcwl6QRhcGHe2CfY9k
+rALBDCseV0Njf1mJNM+/kUA65Z/oPuLAVx8qGvU5sVdcVkxuoEmefUiaBMjZ5hhIipLMUcCK61d
yWgKF+h6P78Xky6z9KyQyIFjrgoTCHJD34as2IESG/0+f7ikk5mBFqArDciClTCB8tl0GnwaJeeD
jNKMLb0KG+VRdeTQeTibbnCD6nYZ7n6FuC7pyrRCZ19i7Re50sGb8NDMTfkIzw8KZyqDf50ZubJ2
Urv8fIVBeN7KN2GODkEU0nKPuAHlZ5wbap1qIb/HgVTLythoqJUEXgXnxN3lhksPyIEBTg04qCU9
sfw+inrZQjNOVI21Qb6m+zVoEsbHwqDI5W8OVjCw37Vm9Y0XnnjdzFy4Q/p6lhy82s5MG4BOsjoL
jmpKH0jE0Rf3ubC4BvTVVAxUypiBYsbA5auFCGJK10Vge+6IypRx0x7WLgCHy63hDBSrw0ySf4Iz
L67WGPi8POKC6ymjM7A9i9QPmewW3E/hXVjyg5f9TPQs3IPsrGHQBbQE50G6I62K/N/xTXneczBl
8+Y8EquUFEUdOhhozns4PIfgUEgN0WCAe3YRH35W+iXU02f05VPEo4USiYLYW20zNi24oRab0qlk
4x0Sc8ThXbAvEjJE0AjQKpgJHVYqd6d5Nnqj/mzJH8B58Z2qKyYa4mDPgGqZpalnxrLGetSNQpWl
pSMn3EVzgVUl63PzjUekcEVgNZIktrtz78bAVQpTNMSUjvlkyrtBsD+BJ8ij3N+pJZGJG4k64OyD
Ntt/IM0XdOzdxqch8NgH+tXj7z1rCdCVW3yCbaCeyXLxjX65zMPnT8QRYjPst5tDf1t1aP4Z9j7u
Xaa0UQwR5+140uN/4/hLFp3CKu4HasRsyOnN0d2nn6jNVFH+ROCH35FK0xd5AWRIj9eD/v5kTM2o
PbE+0GuIlQw/LEHbWUobKKlvK2QKy4xaD2qC+DjgpHRN2hW6TCQLMcgd2b9A29ym9zgWnGsz1Wdv
BZLSKGKvZSsNrpItSWSye3Dj9i1p+TxZcW1kq6ajfN1JjF8Ik+fjD8waixvb8fjb5TwfCVXM3v02
ravxU3gxhy/m12qz1ghjiRdnNVRae0F8bU4VJS8FL0XId+c8X8ml3fJVf7lBurKBxfhclfx/DURr
1z7LP4SuxLQDFVumDtCIb5FPjCyaOI2Txnpao02HAIfvksePIShPiVZYjgWcwQdBWAPi6m7qZg7P
OolMjPT6ecYey8NaPEdXfwbxgFVObXyr36ZmXk86SanYpcXl81yIXJCmYDVhHCX6/Q586JfW/5ej
52WckFudWE2fcgy2QYRatF9n5OAcl5cHAt317Z+0CTglfuoakfWS+43MPjF7DgE2ISXmNOudB/Fz
hPLjlA2sqaQYsVyYxeY+DMjIVBadDAhKdEiuY1csQJuA6kDXkNBlpMwHoM31wfjr7VWhm3vzMpTo
rGmX2UZ6snU31uKPUiBnaSLKhTlzvpZstk1IUIJL9oyngFBr8tQFSIzqO1wIQKCSUqoEkhAYZJKw
+isGw14bjPx0fMKVa8q7QdErwJ4tJuZCJ7HJxhXBkpYMVUnmjYaVm7GUe+A7iAw+2dhb7kBJ7kk3
IxPUZRPVuAJYWfSau2a/SFDQd7AQcqeA8AdzgA242OtYfJrU1WwCLvsSaMYWc4O3JyAApQpfCeii
3jQ8uyG94QI8vXJ1ctuA6dUD9QiWaZGklqEW4pbHeQ8ATer1UEYGmVlSsqVLBJdCLcrXr897hV9b
3W1pACMWHU5s8wSnMRKt59rIer36pyRmKDri4kIG/oL9zPassfje0s1vu+nVM3HBnCz7yXypSjB0
wqLA69L8qqDJpumYn/BwN2iDc1ozfEoDLY96kiDpM5cVlap9JnUNoFPavsEqwg2zt2zRK75JrCnO
3zFOn/H4U5ohJ1iJu/+HXm/gvqGSa17dbv8WBypOLrJjxLnyL+yv1SWPzQdAx96HTy6kC8UqEojD
c4Zoyr8Et6kpTafIo4DPVy22YaALhvNmo7Sk71OzZ2TnU+w7B8VveqLKJNUHjkqm6eaexsacB5yu
0ZZ6cM4u1++ap3FhevQfPMZyGJiWl2kLLu/UXci1xkkgG5lfPeZVQ+14vQ1ieBrUicXd1yvNbr75
A67sJDuFctvigWgoA1QPjBXJJ5yz3LxIrmPCUt/vXkulZ086MrtG0QpBbnCyyoASdOF/f+4/QFhy
wEXyxmvyjgtwO6bqrZtNnMdAhpv73aW75ruqBGlnCX+1HSkTCuB1xgbKUj5saPK+TCAeQFuIbMuz
54kjg0jelLKAoNdqA8nP+fgtiJW/txdcz2L0TeM3lSL6NgXngsngPzsjYZ5MFOGD46iZzB8vV/4H
ub0ni9QCkJFdsGzYb7Krx6eIoM7wkZ+KpAt8ogc25g86WgOOluCp6P9hsIvGc7xjQfuz6xVhEf6a
gNYHngTUTbrN4PnSQB9hjk8vzzl4KtMpVwZPjqR+5WSGhLhcH/w9czzMd04IiFzXrJYM3XgFQI7D
isysd4PUKf32kk4LmUEUDQte5BktmnuM0V+maSJFpOO37qlVu+w44LQiUaJD+iI6wOebMKjQfQYG
b+cPShGsKuY0sYlmGeQ8LxRHv7saYi3DWw7Oo8uJ9Yl3IzXiAPAAYo7hPEuFKgoLIvgtbI1vDzRp
2AKS9gGExpC2A+6EZDp/8wcaQKYvcVe8x6YrxDZ0Ir7OS+NwtsGnE3yjw7zb9VUHcdZvVSVV4nSh
Rpun7kR7gLwRt2qeCnMMbxk0LtA+BEpwXd6as4BQDzHTCdmSy5aL8rRQEoYJCau2A6GW1NFYvWqY
WLWw7x2e2paAHIuz6GIZ5rkzmIGwNWFJPSmmJfOoU25T5TD6xWBSpUjKrNRr1eA+mQ0eonmzhPoA
SHEvTY/aB4448bMQyPJghPsVviDgs/688s1NIZALNVZ9OyVS2qAYrID3gyBhz0riqly68il6hAUK
nrWrN0KPX3iPejYAcPvpFRzInyANR5wQCo/3Weayxsogxx1o5Y8Ts2Ws5KL8y741FHJctFoI4Q7I
5WR0lW6mQguqnUyOheW5Spxw4NX0RKrFvj1+16EjC4AOPa/BTYo2BXo8s7xPWLyyB7hfCT50xVLg
rR5ltMf2KUqtz3Op1tzChddC1hA4PHEAR4Loe5J/9I1ZgjCV4hnfv2RGNifik6y1CyWWFPKdEikJ
piN54+VVLoLSsm+QcGAgx0/bW0bIIR1zxGsGGVGV/EcJESGvXgGBF6Q0n8YfHFB779IRQn7iRVxj
eRvrzAg16qHzFmuqV9kCc7LuFuR4Jc8ub97guB0vgGqwIMLOpqrsEySmRsymD1PVC0+aHy8HchV9
KMWQvDXW8gbIXdsz30R8F91rZnlaK2TVqPfeLBtvWKM9rprwr2jA4eV/F8P/4Ou/Epga6iL7zQek
0IoHl5mzMP5nqmM2Aamq1qIfwWBaGQMQxQj8FM9delliI/Hb60mms3HtiNyv9kN/ioTSK3jUiweS
13dRzSXwpaw4nJnr6ephjCV011ZciEpovClPBuc+3bcQgKpA8WxlUWYzYHnjwdQyaZFp6KVeKFwi
EM4Pibgvg60rP2hebFIIstLYAc6rcedIio2LIL84eSRVNeVCn13c0fmcg7aRl9KI868WhVWJ4z6o
irZ6fpeLX79bJAMlvN6XJCEBgXwmLm3l2kmpsYX5iRozdD6Sm1v/Zx1/kuXsbszs+oAT1DC4zscr
9F8jJCMEEEmnNc7rAB2BJQbUFNYSHtm/81ydip+WTYfs2PnHbavnFWlVrapr6t1TqnJCu7JId9IZ
/wxzPFWYUughHQu1aHjk3uHgqItZPGKQ9+bD6o5WW1BEv16c9McN2gqG+WuU9gs72cR3L7ZS3Oat
LIoro4Xvp1wA+TDIEokivG1cN80aKrwsEPCPDuNuiwZ4rZsub4DCBSOzCFK5CvGzJGw1u9+7VChf
b3TULhSqKEHyX3Wjyu4cv1GK1pa8ui7Qo/VI6azbe8VdXEKrqq8DeuMRK97LR5NZrkfWJEwNKUbw
QSktZE2JaliVnlN4DS0nIrSvzkKz482BQ03vVFnlwlG7Ue0slo3kIf2qaSLpChuUzmcxh/pdHh1q
vtxqWkcdeevvSvmdsrYf1Y+fIfLSYBLPY6hrmaDH2HsQA0d3+bCLiuK56tYpV/mEuf92l9+chjxk
sO4YXmfKqL034xtpBNUIe1PDo1pPlY+LHrRNwzIIMy1qcPIyOTanv5LM/V61ZLz+HKPzr6QgS3j1
iSziV+YcfJRhWPV+tFb8QUmT83++SOcx6u8vFPIYBXeaZfU8CRssP1z1v/LxybLAGqChpkJxmBZp
O2TpUIvESDld0GVO9iPEuYuPFbtcof7lcmecvyibMSWTL7zJnv4OnVIi2qlzY9xAhjYTeJ7ssOPE
ZkBRVw/ua0XICVtPtMSDPKzTEaIc8N6I73qOQWqWxdGphdqO5O/yjkKojAxikfiX9cSRhv7yeVYB
WF2zBL53M19AdrNRKgrCTa0KdTKQGP+jq/pqDEbRDNCwIzimtCKxDeUjp+qpE3TRX9VHmnzAIJZh
LUNye1WU7e8kJ48XPLuzoclLMzvssIPIzkm1pvcEloTi5x8I7f5PbLvkSwQ/RIyrxkXmfLu36dzR
TO3bJ59AD2kI+ff8lWmf1V2rkHXiCEB7kCai5x/mji/ECA0Y6i9KFSkKwZ59OytLQ9tsl9mOxJyj
eGdeHLYTpCNz0MJYzrMBhThrgX0YzdvIN03PDqaLDfiddVrJeTjxkIfu+1EJEA5ZyWpz7siSuFMf
KNPrgx4Ao6ciC1gOz+4kC7CZMryNqlBDqVef4ptigIogDrKRDbh4+7voUm6s/hzZDX/b+pnRVHmq
gWgaf2BToxD51gtvf2T/cPZRZnNpyBTXNV7UFAnKLysahLXfI2EZY1Xj+i04W2p5q6U72NvtkFPY
UkT0HXi9p9YYsHJ7SRnzw5szBrSFiQXd1DR4HkvJy53+biZJ5RZC+G7Ys0ZE5l+pd3J49DvyTdL1
1w9beze2C90fCZdyG+S0DfC5lKiRLdX6VBCK33fdlVf5cE8jt4iqN5kyLf7FRKa4skHc4YbBqFzs
BRaPN7xhWErxbw6Mo5T9WTCE2UhHHArQFEkaBz6UAbFy79p1bx2Gvw90p6PgiyVkKqW9rWC08hVb
ISFUIkfNTmpwzg1vy4rjtaQNUqjZQjxjkcsNMdr49IvF51mPijY4YVoirWBB1zMCkEyrKBO7iAFM
m/nYuOIZ8BindbOp+88OPFn/6dYp8CjhXLtiu4RnaikgfPoxl6OD65/EfzVtrR5bJPn4fbydQzPq
WMVwdE06RG74p+Zd6PnPsBCX7rxbDQiahndVSaoVOcFwQJrAlUeH/7rnfunWGB6AKlHRU2m7n1N7
sovjcwzB1LyvdLBszwJo2O+Qm9wD0GdN6Id7Knlq8uMwSGo4lsy5x9QuHoP3/ns0TQYYKBmwnF1K
lZ6nkGdSOs1tsb66z/diR0j6kS+a25ONblE/RPQ1lE/rrx5ZEj/g0XiLqJbjU9yml5N+nDsm+uIO
D/kdgaotyrvOpGXmtSVhTphG8jtq4KXUeQN53EiKlPGEvnzCB+ukdh3qyOMkENx7iwkzvfDT4wpJ
760pUETiH27Z1o6bFX1llmrrdkdznO7RR5hRArCbjoYe4qa4ZWcXm3UwhOEJeF1rdqnBgRrqzHrp
PpcA6BFh3TksSJYMsxj4EBDN2BuhSCHx+/OGxc98TOQnLk4NAD8uAZYF/tTFgveq6uXes51ZGP58
+6LcNDW8jTuan+XeKwskc9n7kF1DPl4Hpmgn8bMaTePuTwwwp6ava8gRIznvpn957B2idrRUl1YE
/GQeXKe+WipD2oEzt+o72ejEO1sBWDRL9rZXLrrUpTU/oYvmL+A6J1plHITDxjTjJJLPBBnxeAuG
vl6QMR3WGSKiVc/eKypqxqmxzzPhbUVw5TPRuq9mT3BpCXxBnUKHcOwZwP0foVJvQZELuuu0IDzT
a1W7PRIVpjOgSoEFMdAuwe5sz7mBov0g7IUsW4AP2MW5hhJwze0lAZBoFkyfc52HQft7JHQQxKDK
/UELkZFe5Ldd3xEEtZ7cRRtyGKjVxc9d1rM9+edv8EOrYW58WLI43HWHJJ118N5T3aKa9BdkZCVk
+FMD667GeLbc6HGqGSrTvRyxggGTtRLMOhEgkKF1zRXi4zHyGJykd3CZU1kthbuj/A0Q37Sidgp7
R8TZcGIpMH0pz+2Y1pIO+ZWg03ww20A2/s1CZVgfeUGXKtGa+v/5Clo2woVljqBOUdPfcLmPrSM6
i172rW+4LA9Apt+q0T1HK3hU2RrMu2UwgGjkcl8sdieLpCmzxCrVNec4m/Kq/dGTe5FWekbNvVY7
heG/wevNC1OwiRva2pZ/UjEusqVb99sQN8R4p2/ihC6hG4MyodK9McoNDdMg8GfcEKdyXzTJGfLo
8sRLJPfDj/9p10YKl9wosc1YcZ65kd4cTMKN9ubIYrGUBSeke5A8wGXhso2VQAoT/MR7hcDbUC1H
CpDuuIwZNTx08IQ3hzxCjyga/eJeqU787tDBOugyL40lIOVRevfKcVxV3qLCLn2pA3xSN3ekZxxE
bAhwTwjzNRd1MTOX0g4nlv1ktd29P39ZwvoM5vGydFeTDiOnf9WYnsJglyhDKt7OT+efsQC8JxBr
VVMmBmhPopbgZPUmfpVv/9udflXZNICEYcTZTfaQ8aK9545CkVX4zw2LWo0oKVNrWRY6UqGAwu8N
fLuJ87kZKG1kG47wZ4KfcymCGznrEoMbVt3ifQiMwhCxWRbQGIRHF6+je7O3puGBPXdJb3NUnPFo
7VcYOeBo81bZ6B83lAZJ/OLvRlbMuhVZvwNN8YnEnFfX1RtGrkph/H62x3ZLn0WRDX02Som8zWFQ
9rlDBQfnQ5VwpG8FUUIv5OumSGskgdZZ58RkoSmPhc+tLG/aislAI6ajiA5zjQqfA/9rHVvpGPFT
AL58PiyqTvWNn4joV12dXHjA3btALVCGCBt5V+4jl1SmT1D6VJ/k/XqrN0F2shee2eE4aXvCQluu
NB1b1vgO4zBpPhmrzu+SjGPcBiBQbNNj6bNzw88S1QG8NwAy0SfqbaBlTX+peqDHvaHap7E3tVEt
/bAOEhXFr/5V16AtXBQuJocLvbTeFq8cdnQhkYj84KUT9MI1bPypKLCW5SbdPr4puVrUPfTJC9wY
GeuYZQciA/L6Qbx4B7dEb0oaBlcdw4MyIWGNvbjUScuCHyTTUXy5ydRDJq6gg5Axb8+rxcN10O7x
lAm9h9/KPF7sngyxo+9K/EEVn56SPQ+SLCUx2TXNsOo5/SNtYxSuOcCLOqCy1MfmedbQXS4B6Wsi
tMSH91snTMWzHndf309VyVDoJ1vT4hgz8hn8mX/M662cleFHzrzRCC0ABWw90aVOCenLYnSCtBX6
kTw1acMpMQXHEkjO+MJDtJ783inT8rnNlartxQMVtbUz/t5FcAn7kp1ENovhfI9ICYos4nF9pqkv
/LEd494eYhzK/45J+p0oWzktjy59HAvnswEoBJ63Sr793tyKbzg8k84FbXjhCcuyJrhQopUzDbU1
BuwVW0D5ofUTznFdC4pUgh1yT4/L3peSYe62lyNh4eKyiu40209bnpxUYdmN5y1O7nlZHhSXjZYf
/CkCcHToSg0Xyxk0caEm5Sukbq8kPF0Q8ZOcUaEIhsOe3WEcAk3yIVqAC4zYRPABbUFNysN8k2dN
/EqI43o0HS7y5dXCvL80Yz1fL9vhqhC3eEfl9/lg3/mmFTnwGQv1/qxEdZ618TXiqnpUlwk1pBAx
/RnH8FG2wuUkFoFKSatxeB2djg+wF4AT9bIwZceLPApg2ir6aTnUV5DkqW1WXdD985FAZqc5IGJx
GoJgnIazoZF6i97Lqwr7C0X01E2JvsXadM2IEXKPDW6TWVKIfhEusUIOZuLXHnaftViSffMj1l7X
N2Jf1cTu+PF+DbqgGrCE0AkQ4eXBFwxcgGNKAw6mwgOz2zZMGL4RxuL/CId/0/FBVdKESj1EAcVv
mGoyXtrgQRtsT9cEoliSR5befl6qflZKDK/WoXdWSGbuWLtaqaLRQYCtT1LATDVDjSc+Ymlvno5M
ifXfkZv3f8ZJgZfGOUCfSYXwB9r0pI9n5UvNxGRVPEQz1WcGmN0LxwzlSPP2u+b0h2YJgkzDwll1
5JucpzgPtPwK866s584q47CtkfGkMP8ZzKLck3oKNjNCEJlDydQn5iWHPL4v4y/62K9ftX8l+/Cc
7Dw2J1ZHiwPW4fgxG0ppFtZDngEYo4QFbcHViWdouyQ0aXoa+a0xZmc++Vq9NJZld011A/VnPbDA
2UAZgjuOYaE/NcqglMWBJMhwSlrPFQAruoFKY9hoTl0/9O7ckjM+P8gIh7TSey5QpxgCZgY5pSFo
7M5Y2UHM2caAxdBm4VaFseVxdwNkXJbeinPN31tUkbVFX6GrxNQ0ovNgVmDx1y3ypotmPgeKyL9E
LLhkyjA57yf/xjJt9Js0e+/Nqy42tl8ofOrcR5TElqvRS49g7Q9YvPTlHLYLKVLJFE54LH7Gk8jd
+FXACuzr8gdURGm52YjHC4KcFXU41BSPyRkZjEHVdix4zDsVqttWRfB1IKLk+hsNPkt4ak1Dp3p8
WIQKSJ4U7VUDO6oS4ySNbb7nltGz1BI3h/o5smeT6L92rsS/94cW/CH9cHRmLiXGk8qku7T2HDEF
xNcwWqvJ7H44jJoZs2jqe9Fhm7iwDw0xS5q7gyWdVTFWeamCKQ8iPv4FnzJS7m7TE4bNTpTQdeH0
KzaMBrd2X8DfgAyTLAZjQuItAHdameZpbX9Dwlm2EeGAI+pdUG4+jYTalBjUpcCs2QOlSBAcbh85
esTyfck1eIWxPf5C+tfRmV4uhcWYuqp/LeHu83dmPT1dApgk1Tm/H4tiQrMxkSgzIvHiRJUx2CRk
OY/3s8lXudoceWthzV7P1Qe3cVjwON6Zq3a31nOdXZP0GSLO1wwPe3B9WKIiiSwf3fOYneznwvAe
usz3oM5xWPG/ANSoeRuhqj/hKsnawn7Z69cZtkcAPmtswEUSm7j2rYCdBzj5iMuXnkPQ42jK/vMD
gWYGV7iH7x0VJDJo6GQGzzMoYv3OZm6Qe2QQR+rReXvFcYB3MrOSJpb4emEJJ39dgEqi2+daaqn9
SHvV7jFBlWc4jPjp9tnISSrfJgU1RT1MHY7J5bWgo2n/Qhifalk5TRVsfxEBRDQJPRtjizdapXCM
XjFipz1SxM3cP7olij+yfcqc8w3DUrAsnV0iryJlXlTlWk1+TLSheyc69EfsFLnAWHradc6wPXFL
DlO5kDoNWQf/6qqHQJWOYW1y0OgK7+O62nYIw/00699ZmEp/jdMjMG9k51pQOK52HkN3JbE+U3C7
vGpx4e4FFRqG8wq0fW4fyj7x/KQmvMMV3lqVdXcy8NT1oqlsm8I+aoPojwsr692khKJb/JhZfRw4
sYLDfIlQOnbQd1fqmuFEPaHIg57ffz+F8+Pqfcs6OKgdOrBBydr9lpEA53QGI+51j02/DISFLzpA
dyN4cUuOSkE1SCeEkwRk+9GqWA6O1TBfpnd+1glDp4P+P8gbawDazkF6Ystt5vV5H2jWP8sTziHR
LUAV96iAqx2nt4MvPtOwXVJM3M2TrAbayioyYCKB/oBGpCSANm2dc3eRmarSgiYvP4c0j9jElYCl
vUKhY25e9YYMF04iv3quzeO4XRqQJNQofjznqUo+p3cAX/sFEJt6T4O4B4i9rCKWvvAAhhwUg4Bw
8E1+ztbI/8fyrCRaL6itGgbeQr4RlfKutzlXQdreXgsYWG0zFrC1FLHvJXvpg0bHJav1yZCKy2a3
E1EOo0CWjnCSN2BH+9VV/t6auqIrD24xWJQd8HRzh5wMeRuodisy5BN1nz3iOrnFCX2nQCpl9y/q
ejBuOy1yysLQA3flwJdUyEozFVbjYcVHh7Dq+86psc/Y76Umt3Q5B4fWP7cxEH3C4rmiGsbKyhQ8
FSoCRt+bRO5zEbXXt1TPw1JkXfCmn8deY+U/26gRwollduRNMbXo4SbPNNR2dOarIFX450ql02Pz
UsviQjaAcTuxyZ4dFk+jiu94zofe3SzjDI1xdaZLDEVE4uaAQHKT42z1snjt23VRHZyaq781ZQlX
+lk/48S5s7WzustNZ+BXQn+WMxtNjsS3iQkR2rpSy/GL/eEf0Wd1Yjd7UT52N6d3Z8IbuH7rH0r5
Cl+fLjakHh6jmiOHU8ujNEz1kS001GOqS6PrrelmilHsEI+ByBosznST66BtHCpxr+Ppq4qaB/G2
1WVR1mXWlB4gcUl/6fIWcc0WFdJqJpfKWzajtEuEJF8hg4nc7VwSUWZrLLO3LcVuTZ7HIcIk0pZx
OXD7x2xZ+xwyVBdgSkT62D1MQL7QkDA+4yZDGgHrBiJpSjGO5NPp+f8miWGNmZJgVFvhL93J4wF/
3TcwMHvwMOCvuDXx9YO+cOCHLmXBhu3sTlehhL9FoEonBaNnlpPtYn57+MduoqKAHNAui4wIIxvm
3vouY+uTIryJ+ocjqqCYlcCg6TCORWO+HxyMxrflbd/61K8pvRM7CzC1x5g8kfyWoKKzp28bBBOp
WsFldOkAj+9j0608DlsoFfab8gFkos18DcIxNFUyiDdXoTyLTsdr+HYoftfG8YtZYKkQ43ANj+yA
1eQgVq1R2CjQWijhw1FAsJlNF1tBzKMs/i4zSDDX+E5mMKbXdW58QrWv1bkN9v789L8AMqRE46M1
EwruINp4hXBqYNYbQZe2ffjUKiTEggduLX5CLzBuhWeJTrucv5g2uEU7TMqLp3npbFfLUgXz9v7l
Ro26e5nE8ZQNPRl61OL00KH4/VZn8UjFoXmAvpt1LQ+EE8s2Tx/GMIri9T7Cc2Q/sqAGAkANfOpj
EQIrEiyszUwUWTQ+hAb/9ZJPm4fhQWUdestbT9czDTdLNC5vr8PROYhc1txxAI3m9g8i+aJfcb41
HXN5a9EqLVu670yw59idG4Iv1kzJii3fLP+ehzO1yf0MQEsKuXTnRAOo8629m75wCDmcPe9d7zva
iQH+kBZXHPAFRA76QFrxLNpeuDFVUEA+F8Z3G/3fis7unsADKC/AoMQWpXg+VRG35mw0aq5rotlt
IcRLwXQwZUhfISWZycQ2rtBu51j5kLMHlNbKxZTMmXq7JUXgo1lfHKn07fbPwx7xwJvovIoKPTu3
oC3EDQFT4y4Z2BVTMjcT7iOJgpnlqutxI/DQB8KKUbTUewXXcShYI7fOaNJfdxURjGt1S0+vEboU
ZAe+3VVCL379VQpxkCO9saX8iak95DE8j+XJr2+CwYAeBMECm0a5xuFI3mUKQ5TUmZMBlSY/RlJs
8aTIusN+3JUNrsaBLvkL8xjHj295CebHMwz+clLD4dJ2gbGZOhUQdQBWnWPzdhKgoqTeMZCpYPzR
O7yHcO+6N28zJhm6Vt+UbV3EN3PD28YU5GoHO3/FLugpYqaUGDLMCKPCyoTcZ/IAVgqJblP01Ftk
cjieMWNEI6e1Z1r017sOJCdwLdrc8clu9/Stai/PUiIIjIlIR5zuRGwMZEmhhWsaUSHNpYnCiGNk
FB3fix+28EihnZXSsLzWq+tgmbpRx0wEE8cEF6hDR6Qu693MF2eSPiwa8HAl+xy61wJiuvQbM4FE
sAeWZoE8EXNmHRASjV5jS+hmI4baY5vfvh48Gh3+CTGl8XPF/c5pW6Nibc1yVyEiNLlHkP3XIjIX
VAzchVOkU5menxRCQMUGEpUtzLrFs2OlpIuJ5tnZ8imFzYDFz/9nQwLwswlkIVSYoZCG3z+y5GQJ
vEtNZ7hh2DOwEbcEIKoSHmUan58vF4C71ivcDSy0/cJV62b1O8cvuWbr5Qqd2mnEtQfxxAhz07sK
kSoyBTH0a65X2noDeqDKnpTx/IdI1RKiiU5hsm0bHMM1dYDomsxis8/pVUV17gkcLGLTBQb6eie1
W8Foi2k40UzzIAxJ43Xi/bgBiq7rgKJaOCPV+jGmYbmXkl8xgAoU2sU6fxKB1geRTUKfK+lZ+sW7
TeX9/FskTXjtZWoCg3J72cRVrFS9v1g4tf0gR0ADCYuy1AmFFYF6iVRJJ43VP9IeOpputn6ymjDE
zX+YK6JIiND5z/ytlURfsEjOIHfkX2S6I/ys2diti+5kirG+faWggFLn7UT/K+KmKg0/0OJCSYfX
AJGbPpRXchd/EsNPPN42/xjwCNYUe5Kbb1FYpXPnUp/rPdOysiDkRQHWpkHcQJd3hOCmKMge059m
yERRZNWBQz0VX7y0tYd42soVmjlXdK/S4/ojfK600M71DyGUwd3HSgrOyAuITYkcD1e5W23OjPGF
IirntuHfd1U5pRzMnnsy26aYCU9rgdXunsgYIwEYd3NVSetEilwixY7Ix4GHgEdKd4FCvP3ZjAm4
GGp0EDz9Du4Y18/JrfsQJ1J6Y35bxe7a44iVi9P7xmEbYlus6PMPo37Y/eeh5RKrpHmMmahJSZye
bxEdJubzYY/kYL/q1tEXck/FQuPRW3NgIaoIpeh0fbEpg5rFgXO5Buh5sRYNhfYYggOzoqFylKF8
le9Ko7gaU3u7sae/MHI4Zt0Y5W5eeAfFczHaX/AGQ/N0By9W6s9o0T3z415jJuBMnBLZaylgdI5L
8yfBJgLKdBgxxefgZ4P75HqTnxgnXkEOWRoXJm1uFYc/SQpIqpnFWZ7RH2mE6MpSMG/HP7hB10if
k4o979KmNMQP2Q9sBd3vN0njvOXi9HaPwzrv70764Q9PywBi3mhTDvzrh0lvR/+D3bzkDoR3JUqg
EN58nzr+EHDihRLpE6F6Be6dFRYyFkqmDQbqfxXeVkfUzvK0Gsbl0/+NTWA/pKDeKE1bpaAUtycH
jOrhKPmIwPrKUG/FQFNnzazEZnC/QrcndANb/nMfbnEnJbYPOw9ig4HtQiilQU1pjOAehF5V2/dy
CYwLxQKAXC7X2vsUktwHN5UUU2Do2G0E1K6+Nk+mHDeKyvbi1GIi+mrl8Bwa6CWPXcbOrabW2kn6
9RC4O9nH52nUrwJakbCLEJ5uhKxa9FR1Ijmk0FD9N9ljTHmUunBWYneEPTQOQAsx8NF4BpHNqcDt
7GtXKv5hh4PN1d+ANj+aYKKlCwAG0HjTSLs8nR32sf/xoW2djDdMOnRlEayXHtsnoigM5XgIS+hO
3shgqIObj05D6fNadiV135tla2e+mPRKKUeU3ZgPoItytE1z7SMHt5iIdzRx+M2D+MHQa0S/RR5A
YRQf7F3PiTccZ7ZnSWu+nYbR+BRzjM74o4vXSYKv2iabzLLepcjyz6q0weNV1agdRzXEoQ1wr3qO
ybGL2oeAjkQnXVDhePHnp9ip9LwWs7L+4vx1PeCMeR78GfhpBYI04suoUVCr6Xd+y/zZEL03L488
6kPaIqxddzXCWZ/ugiQLAyuufJUzVcw0QtfUtbukgsJRc+S4sa/euf7Le4xDchowWsjrgBd43Otg
S2d1A2ccWJK4mKh1oxdXWlAJAtxK1N/FKxy6SN6r+vpI6RALkuG21KFBSHKS2lvIuwbh7z5Xg5GG
uFDe8hErSDRHqe3/u8SV0sJuQMb7bLzwU6wbHYcrbkok+2r3r4DKKoFiz1P0VqKXK2OfcvGpQLr1
UPeVVVPCTuTsT2la0NDRDQjs6OdKJUn9Kn6cy8bhgXgfHXjwby23fOnt1LN26qkga+Vidv7VTPuM
9o9pDlbCnZJYMDr8IpmgnCUzG645XlnO9ikrTCHQKzVMvNTdE1XF2G6SiInTFEbcdfOKDxW/7WyK
vR1PKFIZDJ4oExD39sVKsB8/t8KqVoBV0aPFynGj5c8hdKM3GipLtfgtwnnO1CpIbsEwYQ+ADPTA
jaqmlezE6QrAEm5rBb8rcw9BVbivBVdfodUmFXUY8v2LN8Hrfsc57Rb//UgHDpxGVZtdqLUrwWSQ
GwzDKAwaigTiQJhCBu3/baNXYnqCzAAh1yxNPXFlsYyrk2F8JFUajzaehJx7xXbuWsYX/O001fzu
pWv/n0HXC6RkdO3NwEe2GeFwLhAagHrWH3s4Tk4EV/jW1MftGyvWh3t1RutqwdZkC8rfBUmJ6YY7
XvPspGJrSMEuhp9YstSJpgKiXTXPFBGXGsHxEcjc6xIGKyIeUdkb453P0/xITBIWQjKyBS4CrPaw
cqzmU1ypQpF1IrqI1pHYYnNveUh9UFbqBsV2oblZ6vzeq777kSU/iWR0yxSLBF9cEowgrsN7N1RS
tgAfAjGylIPSjHkDvuBIroXX4dFNXUYXP9FlBg5opNgi4XWibr3YRLOk1cK1lLS9BUwH6o7O+4ie
IwhSR2mi+0QkiG+7zJ8nCTsRyxEt8DJzY9NRpzzsndcEZRaKApiGOY9ew1OUtiSpUj2VDda35ePK
DeF3Ab0Iowi6V5Dz1GqcI7Oh7lktZPmFAUutsiTUlKNVOZ41nRmlHtyoL/aF937HHfENqv0+0Py/
ejZ+iYcciJd+2B6lk0DBLiVji7tb0R0NBah8M7OR3GHFtAC6bSdoVyXkWKskgZSkBNbA6oildzSS
UHgGl5843nLexh4LD1FYKQh+L3dRUXG6bwoFkkh7fQTk0NsEtZandcxhiZgtwVlVm6sIH1fgPTpd
hL+Vy7XdooiUfHtPAhtA4hr2Kx1WxpYxXIe/D0WIJLl0p6e/ypjAejTf4KMmPLLpDMRUmWQ0JC/R
bx5y8BNl8PCx74mTklXSG6X/xQn84NOp1OmEajec49nhMRiDx1uMVofY2zKz4yN0hqvMnOdEzpQg
rNl4LE9A32579/TSdK5kZhYsiVE2VUcestSUzB6jm2lihziFFcsT3x/kKrNGPsO2TVFcBO3bT0uX
Ez9tHd+/+NAL0W5SDnidoqyd9zFX7KZCiEY5sBE8JOS3Ki1suh0RRyvp4IJeU4/KO+V1Rck0v0ZX
vH81Ffwoaq0DaSZIQ+x0n41Yd518tmdoYXhFa8RBwGMjs7OOsoY24GmdD0V03gf2yyWSaGYlZUOV
vWsLlhvLo3O8nyIuryL/NOIgZTaP36NBnorGX5dPrnYiFoavJg1W+mcLbORa5chaymaRvwHp1RoY
ymbgqZj3Ft7ExdGflFNBjxL0u0eMQQbV+GUJF1zNIBauiNIlEZw0d6etcTLa9V60m0EaHFMQmFnx
TqjHenUNYVuHgGoRFVBZZItrnMDa287RW2lFJnQJekt2xOgdgWeQAwwDwhO8n1qNGxNnqY7ny/4R
mICqiSbSm6yRjwOHU91508LYUF6XdWlxuc2HcS8sBv8VI0miiAUWuPjEqC9I5veSoZnTzaUM+CIW
mlahSRBKw4VYx3Nqs/7wuzes3nfsfsTwX+R+WBZBVEnsCL/2X+w87MtHv1dEhdhqUW/t8jfZE7hR
Xim5PIJDeZr8p+5tUF/FrWDXvVyAY0IZfq/xRd+swa+mk9oMLFkHoDoqG7Nv5jGsxYnhMWvIImZS
kG2jRL7+lknfH3Yw0TXxd+YmMKjkzP/+YsZsCNKRBP3qvvBeFKs5fKYaNST3vd+qIN5FAMtCNAey
YtQyvaTGYEZoh6T38usPyiLAxY5SpFvl5y+hHQYSRFqkILybIjwC0clueKqheW12bhupTQ0KPqiZ
KlKmiF4FX1lwg8kgCIz57uOdv5ZEyMqphJzyS0ZezMm778nJGLLOF1+NxT23XKAfoyP2H5b06ldX
INqXdYJ9czWrdNAG+GPhSk5y6JiY05UB+5Vu3QI7HyCidSctxqspOulWV9vCS0cHdzb39+ay2Wpe
EpFNUw0VEIJcV8BxZ+JguBn6LnHtcsVBt5OUVsQlJUlmReySKMOB0ib+LDMQX/T0CnQA630q5yud
mBPlarWDNuMNZWtEMCn5L+JBQFHYEBpmZE2OBhkWRITtk9YItB9c7GLBkPxSUKjioM2NY5Vk7hlH
VZoTeYOkf01s4kHS06TmYITly3dLrAqOGiRkP6uy1qUoQx97vXZWvj/Bs1+iJjqF/izLrNE0SooE
l/E+VWV3Pch5QeKoU/QYwDG1CO6ejTw6xrDzLSqALcgz1NyXjw63mzCyBggE8WIgjMOzD5XnkVlW
2gpSl3MG2ojIJK0Jx1xln8hnHH4yR3d1l5oBK4x0zsmcgGkPIinPcSwrIn8UzJumkhunbU3imMIE
2e9Yw6mMm5PBy4/ioaPURM7HxX41WurAAtcQuu+XEaY6qALnP0KcWsy2S0FIGa8y0rWYOqXsVvLr
YLeMOsalaxc/1hBegoTlIt32wlXd2bZFBU1mcZeWjvx+is0ym9h2+lPUazvHb5SXq4pg7yVp0qmn
HCI0h9nmWBXzPASLPsJCz3evnzmS5a2aRTp9wbTAAeI2D/g+2QxrdC4B/TNjLF3QgLKk7XJ7IEAe
ZcKzgzHk+FwPLFtjZXe2pIR7r6/ztOnVbMa0rej5G4odMVFDRwyvqv+9J1GYbJ2XREH0/abrGDxL
3lu8CH8L9Oom1XjWLwZ5TeVaR4JJhpKJ8AadnXV0DRp/yhEChriBFZCDxpOPMusyGURCI8lmIwxM
gjeQ8eoSl2MUUrDYy5DuUEpyQFzAOuvbF3YpkWTU3QAXXXGH8MMF4mh3fm779dRdMLxIpgas8L4J
bHztAeacsV8swUcqwV6IW5We4DGc5573EQRn14HEF0kaLUuXlhTJF2gmhvyc89DkM9Frg4fSlEWy
+jPC+EzFO1aXOPHvbxl//wq5tTLhEVfVtHBgPIWgosYrEUNmBBkXCQqO3U73Mek2cdVi6DsCLL4G
0W7CJlVaRvGs1PPAQE5cb31JTNhRRzr/seuD7G+JxigxtGlsLMuEv8cGnXr7oxsbNtT3C/nxPa38
ZRewcX+O78baPBx5zxeFGBysliwgKeLxbpC/n/SX+yak4FKW2u2kNWIzrizXaI0lvV9a0EVzo82P
0fQdThq/4D2ZRhGB4tF2YLB7vSnR9QkpQPb0AtwCs1SwKi5HqeNW44mVcIsX+03/Hp+5v7V6PSjw
GsQR9XXRsv0us4nFLKbab6vEFGJdb642TbwjnMg9Bp5LmpZLPq+Wbdzh3q7rsLmlqRxtG5+EBjix
7ynL7tOh9Q2rOKsfSWqdUuPqJIIJpn7g6XoiM6hUDWrLF0SSuikI1GEwOvvhxx1eQcqdyf26j12A
GypQDsiJ1ZSwwDQaWA5vCFuZFMT44mlwgUpK5hovE5ak5/840Gyfjy/XCeJMO/6mSJjFxycKjJ0S
vw6fAy4yg1R7qZfugxJdFg0ztxWhl3tZpyRtvuD+/QggcPhmb8l1s6C3FCtTFO08ygtXcpZXUfqU
dKoNbvrQ5lD8ZZrooanrrr16SzWs7uEuK305P6Tp5RYr9S0st1F2scVau7JSvMX5gWwQkOzEftPG
EVDm8WewsIdBW+sLcoDUpZI97nck8D6OXX6l6o8x0GA7zGVgCOgI0FLdS5DId9wgO/4AcbZ5aHiL
T9Ih4FRSg/Nc3JSiq6Pe3mI1jyeFX0tCDsqkvse57+MLE2BZAfIrqmLYDQR5TWu2wHZfYa87QHM2
0mHd1bOqXkbOsjkF1AtFuQk+6gvyHA6V4X5w1Q/MwYgtDCZ9sZPvoEV+aoTrgcYNIvf3LOWINpkz
YnVPNXuqYhDWLMKAjRXSwNmHQ4FH2xwAobn8PeBbDoWB+1nA/AEW+Mdv9xa5J9z01VtrifZlwyNi
7doyK5Gz0v5mG34QMnwvVi3klL6oV8LXq1oSuUNsFlNwODFUCCiub6gQjwRyNl+BT1kJUVowzE8t
IAu7yyuygZFK+YKGG+JC5EfGXuPhYEHlJqb9tjf7KkIP6O8hAcXDKj52XStUggdwZl/7ip8SMibz
11EklD5EPPxLMhkMdwbwVrj/7jz9SlFgc8XLN4hjA0BrmVwnKDpFMwW9kwU4A+ba+dV7qb22eOzO
ZGAx9dXu3sXwEgFcKCpTQDuzcIzA0ZJ/SQ4Bhs8cFzTsbfEjtMo0IVbtr8WvGBb3Sf9j2tsyS38H
mDhB5RQNmtZV0gPAu9BjmkFRkeycug3BLevh36aTuojkh1YYAY9n1HHUY4kql1b6BIrs+u5/9sUz
mBB82PZIomBtwlUbRkj/ZvcCLs+uqa2vslH1GCGUWOV/oPYi/RPb8Vs9BTL1Giy8zq7sMKVipN1a
/aGbhr6w4tRCQtkXJAEGJa99DDjxKWf8ESV9gyrC3t2k7LJOwv+HlrvE83cT7XGlNr9cY+fVKNZX
0iZRYHcfxit+r1YAj8qR9faY74GK1jtRsqt8ImHiZnkq2Xuvfh4iwVYy4REGLk1lnmwM7h4xF370
Ef3U73ZJgkdUbeaART4BjOvhztoP4nhVLRPAZciO6qxp8zywkPSnrizSxeIvpFuhAx1Fqp0GppqP
zZFMJmd7TINzfoS19woeF48UKyfPX51nw687Ie5XhJkPbPhDlcjsS3ufFDMc89tnSePdcvs75Kc7
6aQKFYAuNcJ/uMRqwAksF2zIcv4kxTiQNaMC6O+baeW3pAX3t3lGhovzdu+QZsGvrbenR5KdWXso
teF+DYkUdy4d/OOoO5zATHyMKYCbilcB3VA5RzXq+116zzVYhNZMynLw29ne/6/sopDIRPIWSeyL
4uGkz8btTcCdvAV/QA4w0ffteLYXfJz/1mx507sg7oYRLe6aVhCo3ZquLARZCQFuxXyVbCXKb7rh
/A+PZySzncKwGFrGAzdXB6mVXQiSvFg+jtAt08d53Em8HyBQH6JVCmfbZyHQXcAQPq5h5gJyGQuH
9zCBp/gisfOMwE/wYHh61JAUqVIDyOlIdifs9G5w1VCIFMCWnckpPPYDmfooOXSgpGTau7nVSXST
H6Ec+tGx4y4Cl81VUvcg7LBR+mKINnDxnn6HtynOT1YARznQsVxSjVw2tmQf34TZI8M3qLUwpSQY
/breO8tQO0vKhcGfMKqJvLS1IraCtN9TNsaqYKNB0PfLGnwlfoXMBN6d7V5gsKpypr3lwIzwc5dM
cEOBQGwIiuUY9386Q9dCuaCjMObuJLlssAGiRHwezU5h7inW34VKzVojAJNoz7O8NsuBrRehvceI
FMxA5B3/TVYU+nWYzT63NQ0vcpxywqlZupdktt6RNxPTOal75yIazZ2P0FURouY185ZwHvwAafOp
M7BVprTJlb1idfduYDl3+8WrDJWbfDJBHQ880eaMF55T2HZe7HIv42FEOtfLhahzwQ6i1dMLTH+d
uqsgQ2YqeptN14pJdDqJEO4aiJCC6BVMpo0huiBnTalOtn5rDdKhKpaNrBRhNUU3KLObqILHUQvA
Cnt5iiIm5rydJxMXvC0q4ZPFAWmjA1mQBUE0TsP7U3v+qQRN9qapRxD65P5RLScaLV/+kUKlVR2F
ZJ2Av3K3b4BmEpDDKU6DZNx42wGL2hNN+NDIPLRFAXMAHd4g1BG6kYZKikpCBJ7GiD8o6gMcn2BI
F9dun1oB93hiNhmRiKCsighEcLfd8U/NbDUkmqg26GNm3a5jpkBeza69uMraspqwnHvr032e2lIH
Q7VX8Um6QN+ntIEVl2xN7E7t56cquwF92Kuowm7bho4IL3WRsEFHox37C5wJL42dVdZt6OviCcyF
U47wlPilKYwCelZKyW+sNPV/BCu1xXtobkoHAhMpKXb7zI8VJiKxUh0muNBhzcL5O1i9GT6tU6jV
a7gbdLjsYIVkd53w0L0+UOfRkufs0AmtEx7zDOOurJwyR6Rrrqj6rSpYxukY3L8/DosIjxStkHS+
7zMpRMs9KKmft/IBC02tdt8Ow7AQL03dY9+CdOXxm+Te0im/HAJLUfMj2LYcPog+/2ogyJCcTXA5
gNZCFRq7nzHiVYNDhr51uzC8xer02dUF/UT/0ygi7CO+8vAm+LU21Fo7h3XC+lqL/E2dhAU23W4F
+qV3cnOfWKvxbWy9xa1NtiSt5gi+4z0fmBnARC/c6c26ecydeZ9uky3TYUhtfOvemavkqusDZqDz
jKXC4QuAQBQjHMaItMv5j6VG/gdt5qWcWs9YVLuK58yFbm8HFFdik7B/RqI87vB0ILHBxi5cLXwz
QHw8IwB6hj+kDBLNRx1EYkImO0Cfp1gOzTytmcGTD+0VmEh6wPwpNMa7cwRKnF9W17OtsAYvnl3/
y2CZ3Guq+BucslY6VIU3rdgpj3b3dCfnfgULGE+BmpDq+s5qMjD2B9/HntAP7RRj4ysMoEOFL2tQ
EbolGajRStwyuMu2DwxKzTmjM3HFNqAT1Z9pTQOm3fE5EwaR+T9CVLlcYZlert3oBFTXu7tHLIfu
r2eiAkDNbOX+S3t0XAgAg0PNO+7qA3JUfQpBbBygX1UIaR7Z2iiQHJf5Enn5DBW+5eG8ZoGZON6X
DdkPGIO8eaOAgQVC2GewEbzwm2mqQz8Sm5J4mvgM8O1PDt7pOC6/HP0v1XVnpzPFOL+nsTlQ1aAr
C7fj/zAiHgLeeLk7mYGICAmOUrmyTovp9djjPm8w7PXyfy4mY4oxbaxbnoc7AvbwiZWLq3s+MIXN
uIJDfVt8+UmWymTSKdH4tG+wywKNyD0XYoZZuXr9s3zspx8toF9c399wfdAc57R8O5LBJFUuneVq
07re455klto4pLqvR+JF6+uSbyyu6m76ozokcs8fXLVdNoo6GY32jqqK2MQmE9k4f4Yg+j/Grcvh
yVq161I/Oq8bMUHXyCsi77SFCG9rRLlYOxRuWZBUJ9NOVXBNW3DR2+OqKnqaRAgvz6B/PuJ+OzA9
QX0/Rgz/JxK44h40C7jsxSW0I5/jaCOPWhD1ccr1P0MeDQ4lOergBWBttJ/oyxIyzMYCdJX+XZ8f
W0vmxsaZ8hyvflw9gaVIbATWAbrJjWetsnyj0HDLPvGf62Yd2rGimVtN8vc8dfq4aIky1wx5uSma
4CcY5O5JAm35F80PVVU0wlBaA+4BzI7Dho70ugpQ1xGkRndrOTMMUKukjJtkmuwi5Yr/eQgvO91b
MmaRcIOvFW4yXtyo7dmpa5zNXmpv+u/BqkGfXhTOi1a+7AD2+Yy6yqMftbTj+xA7BBoYaDNWQRUz
8X6mmsOxqstoEFkdMjPkZDL3I2K5VaM/qjGzWLjMXPFLrkaQDeCrzzPWmNtjbLgj1bJoB3EHjZjv
i2p2VM7ZHaXF5MWcIsRVpqh4kzpo6uIpXG/kdeJxrPgdKc0obj4lN+W5/spEFlUFWCL4nbUmdifV
dnJmKj37SbLYWeVCGJztOmhZVUIaJwWRPWyjdAWb7Iyt+nQQOpsFgj5qeaJ+mbLkj6z8cHG7PmuJ
1m1MJcjivI54Bp4ntxgDUgnhMO3oRmT1n3E05W5RVjTjdq0dp09W0ERGaFWrybWjcDyDXI4dcycH
LcTAMxFMElvD3LNjhVyFNM/EaM60nyf3jYBEgcmvUn6R51VIZ4/1EcJt3Ct9jgRKeIzFSH7fiyHG
5sxDW8nadjC/STwOWGr+H5HY3BJYXk34xhWSXu87N4p+CRH7IXH0PbzLsFy9CMZ5afiV3fAYztaY
c7n/oMRHiCAUD7uVmzyik9VZRziSKqHUcnhM/Jj+SVduhs/Gr87zvWUQ7ey6UtPWrHckwrIr1I7c
GMj1bz4Mid0Lbs5cvSFollSzqgUZGp03ij+T6EMGyiNhyqYbSb1t9cgBE4mud782p+3uf44AUzyp
JyqVgrz4zv49oEDZX7Ccaz2b6Q3NmwqFgfbP/spn/x2oALiH4tzRHdqhOsd1qp1PIQ9n+8gsC3a2
y1PHt+mYtep6Dr4XZ+i3g9GNGwWLLlSO7BbcQvibdGmHQKNUGBqVuP+EKrGVtKaLusdh39Csbe0s
1w0V3gRSS7lPWHpwHVL9uy6Y/dg1uP0eVZOFbrd1F4IPF4oAuuWgsQZpoo/9+EN3FmKYjPDnaBX7
4RE77uYie5dwQiD8Wty3lKrqEdTXgnJzP7NTV0HNt9LoSCBCWIMbMh31W/8Cnrei5+/RCbOiApvY
RR74jSfXxnJvn6LSZctLuRBAfGk4yjaf10kHoK+jORzMZu/o/gGFps4+I26jaybuvEI4m7fsBDeY
i4pVBa3LCZ6iWl44zXC7bp28EUM/tjZv5QJTMksmVNaISoeJFJOrQfMvWjQhAk9UO1rTPoF5FTVf
bc1FoPfLfDXATm26JIQZWGdKsrnkUf8gwGkCsRzVVUkg/62m16P4Cgv1Y6SQXkZ9WBW5WkstJyvW
7EW4Ttj2BwE2pD3dgkikPWEeQa2svfbFFzsmrPe4UUUyCjRGE+GI0Kzb1REN/E06cKoAJdueynNV
9/h3JH8th3jhDJ/gyt3J0z876A6ZbGfw39HySX8ZocqxebMgLdp/R+shHN7nzO1GNdyDVHpIjDeB
7szp03xKM4NOcGoTbE4C569eCkDnSI9W1JoRRpBZlg6EoWVzfcOhpdTaARDk0GPMJAdEti4unnCl
DMl+9bSbd0gv2DeUuq9pZ3sglOO59lqawaRcQXMhBvZjtuwTQzTruFoURu//rK7SCV1XIiFKIWlH
gjjZvDYTnV4A804eDtGkRTqr/lU/RMlx+rR/mITB2hDXaIa2tVbpbBO6I64fw9L4EQWx55iu5h0Z
ITFxfz/PDMbN/mCqsnCcE25YDc40SmKvPY8ClT7eqhVHB/u6EkjwTDp5pBP3FnQ2eqlpOtSdcp8z
RzTw3/7Vf7CND2uYWVGwjSWBh8ZNvDf03cl65VrJklQAKEvbg8pLMuV1Pgb5OUn2kUmVbCDEf66T
lU6HEDD2idtvRsXUz5+7OA+QGA2HYf0/v7b8FJTVexWcZtWUbqdUQIznJAx0BOcdeS5YLT2U1Tti
QUjbJMPQI1kUzyRb7te0b4Blt6lASu+cD6T3Q/vYvRvLGw/mHofwRQh52VTE1ZHDZqOv7mixtrZ9
WvwWYkSBmstRJSxPnc2uH/rNOFPVceF0i5bRo6azj8NowNsmFkZPA2i73hCoTYi6S4Qd6fs/I68r
244R6ufLNFZFlDg5xFqlWjcdteB//i/15xa3HCt3ric4KmpEUAjjP0qB2tmvIXSSYwPODW06RHhY
iPEuxPodAYY8OiMRdP+S0IzJszAMm3fqTyIHKa78V2CePQOFOIwl8h9QjfmbK+SZO30Gq62zHvY7
NKc9dQh+L6ocnl9AKx7KpCIQZZQ2nSbh2hzx6O7gi2W3JHZryxNwV83+UMvnrsmkfJ+v9pp85k+r
UjMiKTjxsaBiRgS6R9K7pUr5uBQ1G701mksVP5rw9nx7IumaTe8zBuxu3TYa3hOe4bzdoRp4OZZX
Gh4DPrHCu6XEn6F4eFnhWr881IFjBCIyiK3u2DWDpskX/utEyoqbDGcbndMtnLLVZYUVEdfqPMl4
gFQ7lLGCkFseHCDqNpMEs+90FQisEhIN/NZaQOwdzKuwkYEn3XVI6oXsE3sfXrhPIUt+g8PO6Xs+
kX0HegnkX34ntB/exs4fAcANKlwBDROPNudmaCj3mqXdO0sJnTw1ByBKtp3gipd2I5mHdFRXGgqL
SOpT9ROvbm3pTI/Yzrl90YSy2bQYye1pz+Uc6TGCs0jDHYpFFWkYhbpGlg8WEgtA4SeZyFYsMtKQ
/gnoV2gRCMy2XT3qRxIAwpFMS6ird9IkMl1+/xS80Di1fA48EglZ8fL3EMJhnlTTFeMG+dCbZQL4
5djlQ2tG6dkiC/7h6CpTIyVrWo2B9aQpS42cTDJLkO0ESAilulymqNRq3u0qwJG+oQzGJO0qBBKc
VWyAsiO2iTRLtJrkGA+/8KBQ6tzdkaoGPupLzXBjRbsqsz8U1gC8/gzD0314jraS9fgFKLM4gHze
2MK1G1pJuDMacbGkzqMFb9+e0NDeBvXmFWEeqr0q+ZO7GoAU12p1hv12gEJNy6t/8HRLX0qx4sMf
033GNgWCVRZ4RLlhDwb97GOm0h+CVpEoSyDBc17lE9aN8wi3eH7h9R+v6zzOk4Z6UZTyXlhvhdKQ
5upD2HZyVQVyBfxSAdBnLcyDwOr2snQIk9pFPLy5Q/NrFA7ShH9t85HoeFXrgaFJxrMheH31Grnr
1xxcD8rfyMimr9dbN5pqkzQov2i6Vc9X9hDGmqUnWrF8lj+eAdPF499ZPd+QDgRgUpMQldXdxaQC
5VqvHuYgW65TyDC3hx3S4x0qBCE9p/aiRU9JXv7qCuYWuXIrIajJIS0uUoc9IPYr5c6rT0u40Psk
Re5XuSySNt3TE/N7eSETYJBGc5fPLKzwQ4ffze/CeQfJUMhKxi30lP65x/1+l+9K8sJE7k3YaS7e
qGj8qO6fA4WUj+6QurvsSlhqenAv2n9hdvi3tnXDLU3WBZBke8Wri0MqwCuMWRMQX/fmvWrsP+N+
7nZm6bihJzwU5XyPaDQPGg0OmoLcNay6TpjgHE9uHb0RUuTLKRR4R8ASEaNxsoFIZGEC8WpK2/YW
6pOo4rC+F6HA7VFaWA6YHdJi+Lh26CLLIAMe7a3d6ehaXwftp/uNgzcaTeNUocJWYe76Rtq9HxWx
itnxFn/roKk/Aj/WGL5gXxBN+AhOnR74puHwMOVxOCir6GdhNlVRU0v6B/36wh+YYd7hk4V5q/Hd
h2VQowE/S3XCKRVsWUSP/96eAna0LpB1w8FhkJMtE3C48Jn1O3bWHLkGTFmutR/qrB4MCElLca8P
0fTXEKJF+2p2eaOOFSnQJjaeAvqE/CEHDu7h3blnjVIP8ajSwWRmGy+Dzay00LAGiPLQ6Z7IXbv3
YUerve4aYVcvaiyKMDYWhYbrNh84k588jeXvvWPs7fMz7iQGK1KtMr4l/Dzh4rZUcNIi0gbMzDty
ce/687gNPRXuy973IvyIrkzb1QAvUP9YfQFiPKmsFTX+NgGqhfzAktJ/vwsSkxICXS3y3eqhLu4u
vO/njmHlOZ1rqizht7+pzfesdN/VX65SRha129OJ9bZeW+FMUWozOerlLzKsIEQ5WSTLDxBUraBw
xWFt/nXrIJGK+A5mBJ8V6REiKEO8M1CRgC/m5yEuUOQ7a1VshZeV8V3UsGFRa5Kn07YQ0u5BI2E8
S9oKu3Epah6TKewrpx3+xokTM4v1QCTTxDv/RPTzFlkUwAoJzs6bRU7ALUfSDtvQ42hQpz03+QOA
5u/P97QZTDd4lhK5IKRnqSNwMe5/asYOzbzc0wDsFI9pg+TRHf2CKPl9tXCr8qvFPSH8kv8BI5gO
4n99aUHsQathn/nPZ31SxrUZzxAjRPOWwfmg3aNBP+6N2sDpHleU+PviCaPJdTtip57arHiAl/Tp
CIDUae/+wdTkCAOunwSe8i/WH0ZzStSza6Vjq/0jroOyNfMKn/Is4Zhzerl7mdW6EUcD6RUADK/C
+/ODD1XgKbcupQYWBfpgMw9AR7lXLskluT70z70lq04P1C6pZ6qpZmvos+hajkdsT6gW/UkZy5PX
SRVjjEEgmYFVakvAxNOHA52Upgr6UTLclfWJD3X/GxyR7BU/vWtaabwmXNuo0PWcDsTaowVLXPAT
XlNa2nGegP5I5x5476ft7yZfcUc8o/3pvO6Q4M2MQnkha4n+lACpbkvHK9juodV6LdEfGhrVBIXk
RZEU7ze94s9BHpzV8Pk31EYDMYOzfS1vQB7TMiUuw4+9tAvkUX4MTAclwijT4ifajRH4pCilRT6v
eMct4bnEhRfxEKIzSK3oi4DWV1rmn2Qycg/qK/TbLhzqrLRqIZddPavqgHCHTK/An6CO854DAuCX
dYhw/XNzz4zSD2VMw1uNUFfPdBnzLK1fuHD3qlGHlbhNdd8GzcWDOGBBSeiJ55Kb1blX7i7aigmr
K819GT9CyIRavrzNaLwwih6bkMWBksmqhJQgyPv8tRiQ1jF+mVjcjL/7p2zRFsqGA/thNZAnSjdc
gcyXC7wgazcjYV0QBAWcYqo7BZaPpq0cPU533hiV8lyQPTCZ1yi5iVU/gGzx4KeqwVpOrivR+L7K
RATBqObyRO1kINCO5ykZKZGQA97Ch/R0q4/gi50oWVUnrvDi8HCYVXsVUHNHYpgcYdVAkvt/gzGN
C0twgPkXw/RPJEwPxBQ8/1I3M4a3Uv34DQxIjY8dQo3WjG8jGtEw26yhPk6dYuhUcZw4Z2Wu6eiJ
UUOQrbNfSPlMnHvBW+o6sts6L3tSY/Tl9YSFpvl8MivIDHm/9PceWxmJyV6zNr0lEbQgy7SUnmBV
RBRwpWEI/U2Pz7ouN3YFSIqUMCFXwuAXrEkGgxf1uwXFiK6nZcW0MPsFIR34gaGqrjMa7wM1euA+
XMnppaUjF5PU6eaan5RCvQbqpDPoBciXg90vOPSsC37Rh4Qws22Mb0IP7UdfpBEdbrh8AVqXoodM
HlhfOGBSeltCM3YbSQBsfr8cSMdAjWqPTKUralwJ0nNWwVQtZMUwou50J0AszvmYfspfWW9pMWvx
S7fRp99J7hl3ocLcwZPFDGajvnPUZQvia74gRtzdYIZ8n776L4mvloJkO4YR90ouUEIejYMC+nfC
W1jnNkJmXdGy7KEO0jiGzYwtdrc7ba+MM/+SFLNBVbiid9eM6nCmLshU7qn55z3ZXp2bpsUY2gZ4
o9uj+BXRM9SslLezu+MGSAQmgwjTF03JRIEtr0zcgaLQpj7ZT445gAGjDS0ZReeLV7rpg0seCfqR
PcqcB/xbQPM+8TyNxmUBdI8FE3QEAgkBWekF0UfwiKN3fsPqnmDeuDZ07QyBJF0Yd+ZNZoQf6ykT
da0gxyAt//KjTt9nlnvDMl2t+b5H8C5PFrM5PFx37QtYTGVUjdtC9oEa+K7KwutVYDmYW0rtmZbx
j54UIZKd9ti7x+PJ9Jd2B+Dk6vYdZSTiaWoD7PN4VIEi0TXKlvOJJ72ZDOz6vII3gMnnVcWxUlCm
hpDUw0LYCN6uHZjwzWind3Om1FHopqy9AD8eWKs3GYJLDJrgnYyA6lYDiicsI8cQvVYVUTVtTaQa
9HP1ZTxvr8Trap45zE6xMxs8zQB7Xz+WjnEBjE7vyjay/2qTNFgKDVhnCQVFKWVWDaN1MhlOE/Sx
UfOJw62gl1B5ERltr/V3tB21UQ3idELgzZ3yylnuu8Kwd4A9EmGNczTT28QV4nz2FO3+Gmqx1jJW
MEIntV2nTuI3kCS+lRC9LyBmPYw/aNpupcQ7rUjxhxc0/C8U3gLAsVHeRU9rq+lmyQLaIkj98ngE
O4ceuUlnM334g4oxjAzNqLbOhOzdW0Wop58anVXlZQspb4YySlpyyeCrDYiA4A/n0Ig8Ky1KCiMT
GPeBNoy8mMkwd0fAc7UIfdKefioBpP26+Pz3FRb2JgCLVQGBGdlThmJY3ntvkYRrJqn5iEPSp4aV
azFXZ6ZohADTD69LUjgQPyGtFyLk91O/3ntFod/z9wfZZ6I8j6MIzo/hwvGHiTB+eZl+L0LZqIo4
o7+T4OMjGkjfd5F6wnLYZgxEFhM+EBVRFHehmziQOvNbfqfTPvQWTKDAqffLRjjaoc3SKrhDVFKl
VUHv2hMChZtgwoiGf4Lm3J0IgBYRXDSsGV2nrFJawfP5VISszyMvGT/MbWD6/+cDTlbc7E4x9Joa
4Z5X6604kFZzTlebMWgZj91ZujSpIrsKvM7CVmmvuUYuzcyE7pwaEEzypsFDi1DFfweCix4m2Q5g
Fc5T3L4y79CuvEWq4Krqb2DCgzBNfKJ7qauUBZjFjRAKIv4OEieRXIC8S9DSHb4GLZqGCtjw98Pf
lEaLdBgUuKjQsCoaQFFGqkOw9QKnOEmJ4E/2UbUTxV2PPmhfK3YPLI3juLaohPeokA7nJuLlg/ww
eQzJnrTHlIZfOHKbnsjybkVpaCioVffBhYNT7LZRY4peEcBMDlMGFXePBU/2r0YMuI7JiX9mbE/8
ORMXeyxvA8h+UruM3F2o1RsXaYSiENoEphtlfJtziuu1ClCHuOU7DXK/1DAaCkKAy+zDY5coHmwJ
wGI2gMtl1gzP7fhKEYpya13KA7HAeo34pxaqBeJLwRPSNRbjSDnZtPWfhXZpCLo5jMnOKx7Qed9f
PV7HSjI/Pc3XRL3E2eXKkVCDEe9G7973Xz7mUT/Y0KXEItQLfJSHRMV9ieaTlDI6mNpLHOhbjj+U
FLoDqzUfbbGKOeU2JW8djkJ8GFl0icGxLCKnRCyYhpD6QRxMTQmRaKl8dbPvKGrBcXd/nLnyS6Cs
dIDU7QsdHFkldXl7dyFvEIsGOjRlNGDzpstcgLAripDB46671mnyB/twp+mwvEgxaY5HTZAZ22g4
oOhSd1KRtSvFs8vZxfELE17DE+7XCuvY70YkKLoRkWveQacMSYyZWWU79sJLI6DTJDM2Gdq4nm5Y
3+8/alwrjdPfJADl2s4gUY/IVHWBXeM3oV1EZG/qhUWSiKDuve5wGy8OWYuCtac9WpazAoArFEsT
PyzZbnOaHCk9ufy6SmBR7Aqx97BeHISFBCZKphNHoQh//+AEz8w2i6dwlH7CxbCpjFM1pqkZywP7
399akOx5bS4oi1T0DNILBWQNyzZ766krhW1jXzNH6oYKnDr/UYvxtLoWlACjZYye2v8wrAf0KTAM
U1c8cEJz5MqyqWSsu84oBM6Zbn93l1JOCt7gMQYcZYT2zQNF4p849km/UyrNiWeS+jkQMV7jXPmU
G4xjeRjLGkHK5iVDOnqaW1Zhit2Th2n6I+asama0QfugCeKb4bbJT4IO8G0fmJ1XEgEaxoIFzjpI
lo/ZnUo0+u+vA3DC2XxpelVQJkzXkISpojF669QTEV4CLpMRI3ZKk0iwHLr6ZAefjx5QRDzX/vH6
19rB8pR8DWD3/9PFz8Ine1v7B6ygMxe7MvM/fLp4glnXU3/qWwQItk7eh5LxL1VOrQqir3SQjWAU
dSwJ5K18YYmg5YvDDgTtelELEuk1j4MGF1p1cJU4qmeE7Ayn9RAUHwpFlTyETwQTNc3tiUVfQZ5m
nkt3esAYKosAKrFK5Qvebb0zVDvSlsPwjl9l54zR7zZM3Xg8tid/qBrhV1iZoDFTAvyH4KkCsf+g
Ir+6qjwLtPKfRESf6FjKsX/YAYn1Q3QorCTMNbbKHecKvdalkTNrnK3O7zojCQ+wT7t9GWakv+wa
daLw+LRT6qsuOXjcyL+CWFj6nALn/yCd9VlzJrEww/Ge3XIUMo495gfj/6nU6UShej2vxc1Gv/tF
TF0bO7wKealL3kQpRSLfOlxnWn0hSDa+QpVrRaWUGENDJ54JYWV1TeMP5NNe4lL6VICDLzCMORk3
2W9tHszS/f0U3B6TRT/xunIARZY3JOPMBFZSvd5eKJwXCmSt4VhSZf94egKMPpkEVYwym/NvCc9+
uH2OVen1Rp6AEgYfXAvdCow0yC8YOwEWuHG13nR4FcIfHjmXVXftOpRxX8B5yf9KBQfpsAD9ig4v
xm1QNOlLwJPJEW8ZS61XXL3PZof07LkBoGaDlcxGVimtpRypxqOljRLrXuDIe4fESH7jxkjCewkU
/l1XRvSaNh8GJIY8td+tpJo+00P+q2o8uAUa/X91QzgwFCKOfEq/uNekkH9TZzNn2qa15vjgt4la
PbE8FJqk7s/dMc9i3FTUXsh5juiSybk9hxOFMNflc5EeHgbzNXB73Yd061bGse9VV0n+9qrGubLd
IAqv6VzsOAmfJ0VNM/cNVs1ofi29iUyGJ9agnxcICs1vUSSJDQPRWdnc5YPCaAFpdIaFWPZ69AU5
sTigZgyeFBZxFUnYIzZdLEI9iAD51MJMhfUtD1cwn24yZrKlq97B+O103aoBp8y/nfa7YNsIXYfv
TX9+xC8GXGssVYwBXue9LSyDbmaBqHm/tvaI1YU8Z4FfSejaTrTn1y/NNyPK8Q/7zx25tU+kokCL
8t/ltqQB/Ang52EcJ7vXo2Cr/x6iX/VMzSKVHfN2GOLFn1+m/ebeqEeasPiYmFwDkSw1fw8EtmGq
F9g015v9CnWhR/OVKC/WGt2fUzHvk7vrERnh1lToXpSNQDknZzWvslWzhnaroZJsMP2+hASoRbf9
8x06sBhf4r2XI+FfKzu8/JMR2+xbb0ybQpVRFDXBqNJQcw+Eqf3lx7M9BZqr/EqL1cvdYHQ14voH
n8ZQCw/Ag+GHnmzOite/amgXp0T1j97tHsDlDiWEwORCpvsH82mJkM9N/BLGwUgVDhfKWUlZLk1u
ULrf975c8KQmqo/yFGttM0x9BUhGtBmwMiEC2PitlChRUoBCogxY5LX55gI31cmYIT2694bV1qcH
HT1JQuewfiwyF5asEADqydAXdhh1qdpyliKR9rniaqXpsJe8K/4aUiSn0Ia+m9155mdovwjbwJgA
pC6vQN3GaJWUQKoL69MGnVOnNLTdJeaDEoHp2NXzhVQMzYwZ/S4BVCP0FNVeap1g8k4mzfoX5R5o
+C18TgvLM+xeiLmxuBDgMP2t/KmNxzX+b13oTMclGGe5rdZcni1y2XlSrM2o+OXbE28k2BG05qPy
VEAwNf36n0q4tti2St3UXVpQ80rqSY+Sa11J8EthbIX24NFsdXEeSotKlsJKoP1u4xUCveK2UL5a
RdLqRtSGqEqy9gcIM+GExP3KIjhyh65sPp9QHYy/C3sP8xiw2f4QFOempcdvhhD8jDeYBEYM/Ysx
hl40l+9XmdXKAgJSnmzezEhewLo8kek+JK/cZ1D63CVENRXBv5mKbJo3KjTYP1v2ruRpGOkpUdt5
oginJyQpQmvu51rq81WWarOTvk0dF63gr4lNlexT2doWvfjj51o1K04++xcgrdZXRpJIZ5hLxqZO
QvqDC2LkW7s0tjjeR26s2nTkpmNEy2T9BMT7dnXgoPmrv++wZcKa2SZrm8Sltm9uZKONmYgK1PSo
MdwD14Af3IPEyT0nNAcATinJ/zXhMEoPVP5bAAyxYncwr2Psa6Ei0b+ueAcahROSrz0wnf1LVqbB
2zOaApWpcXOX0Ux0OLkC8V4dSXvWD4DrwIPwYCcHxm01NXxARmF7S1bac2PHsMk/6BImZW3hG2Ax
mM6yyIVY6CNnW+kh4mnQ30LZk8TltRkYFk+nD4xtJHLAuRpfv7WCycoUJ7+7hSA3Uvb9FJTKM2JT
masd2r7vvXHiRZDUt9kD5Yc8QKFe17DtjIJSZOr6fLsqv0tVKnja7FeIPt/lzLvVLri2ovR6G2RM
sfhRqOdzLvJczlQHkPhRImObtiy46f3WUkJ4IQyZEdU0+fZTfiC4tzLZjasBVKZS5Y6KoTVLW+OS
oD8iVEFDVucMUrr6pZPbxygeVcZqajjm/jYQS5pjfdPnJSjOBx9MwwtuAmo3g9RAHORtg+1hIzbs
JbZJJW+mdpzakZDAaboORE0WGgQ/zaP4KqgIjQfyZi4hB/PuHC8ZXIVFr337PRFofZIRJZkqio8B
ORGxZLhCIud6Gp0i40fhELEzuhvxLdeS/o8PjnMwti+YT7pgr71mHiB4uZiEFVvNTB2ziUbDb+yn
S1GM4Af/nPbQXE92XbE7vESMQcYkF/I2RZzvlqH93uR2Ol02iRvHrVC9X7NchmJt8+b5P452gz5g
G7itcoi+ys/xqv8kdKtK+OUis+qcZvoutHfoPrlMdAsnaFMtQIRy6bFkaY5Y0M90UU0GeQ33Xxc0
Mbg+qa+kUJSEyw66Gy75BjRjyANVFLXbA4/hEvGY1+SN8BEfUF6HB27Jrf/9LIG7IWmOuEzLpv6a
8aNquRsiLziU1+LPiq/HHJ8aWfHM5eY4zoiTHCr/8myVeMHFFxTdHlxQF/xg/glOYnKh4AS6G7pf
HVwaZi1qnzXrNKUzmVXZuO+9NXDMWUjotjVmzeoFJsUtUkSo1ZXCVXIZMTiNvTYycY2ooVky9IGA
Gsf3+FJmIHOpxWFOQeAbG0Ha2Gb/DjAOD/NV59s1h3GWb+EfXAA8x9YuQ2lvDUAOuaNw5EJc9SS9
MDGizxH2USTsV41941twrpmQ2oaeaJH5VVVnA6X35Ben2TKZG1HCWWsX/KU3uvTRNUJEb9j0VPJ9
AkclzXwkF/REYPlEFoY290fr4qJd+HbiGYvNgzPjgKPQ6eTdrYlwNpoxeEsHWaMZbY+UzC6wY5Si
xiCqqonofJyQb0CItxE8DDYTpSn9grISU/mHfRmTHTwT+FApz8W5j/C2Yy0AhxF4mqnJME+e7vXz
e9uE46qYhIxx+013+q1vpEC4OFjsDEEP8ztuGtC8dpw++tvyO8Av4F7XOUdjSVbXMXlEKkO3lTy6
0yErntuUdgzOBwWOA7O4wUtBHC+rkyufU25VV2MS8pPd9Zq0G3wsEqIij+wBUBAAszrZaQw8ZuXg
JnEb62KC4cNWtqIluZMw6Q524k7kHPSbxP2xBcsIbl6x1ToEiql8fcx0LNbwbslEwnsUnO9S22NM
Bp7Xgdxe2y/58lIBNVvI+VJH0Dy9egdNBeT4L0u4toR+z7gAZLXgOwqC6ZK5snE5/IN2UHRmQqnQ
Rsc4NOZkcFkyCB1JZIvUuWwBoUbR7uhkxmeJoUGrjcSc7PklT3YkhwdhF2Gx+uixmm/sPdQ9D2I2
Rnp9viVuPA5oDW6pvF1sje7t3gSrtXVU/niV7fm4Qu2gd269QCw13gKNyzkvHjxiWuR+xYGFO8z1
VZgCGgQMufaJBXrasCUIHFy2ZiGjAeZadExsrQPKtoTvbheqzV115Bu8J4p6T7urgvbr0yVRY79W
zy9PYgL/sfKe6k9+hmTwb3pwjKXNzUGSHA85r6Eo2lf3+1bFpO9BU0HO+Wl4UuoELwbe8y/+Ogih
gmq9cpODZw2VxNBkNY2yD/zPA+sBb/PzoaEKMlG/CwI0uyVsDnNckLoFKaktfMZhjb8HlxuusUDV
3tXjJ7cc+evIrgKrBrhvAbBdfOLt8nWxfcRnRHfy8jjcNZCRBqVrUQ6jVBAzLeVhx8TKT92CBSAw
1AU3VgKdqxdk0J+E9Hi0MaNz4/fKQ2CNdJLyyFnTlwerPJErb4NJB3IGnzblMoJYAwizjBQIuzQQ
1lNBMgkCmqZ8Hs/yQv6ask5B0428S0TLjzCKSOV3BAlPoVfJkPXAvixxwRGvc2ADlayBH7jN1z6V
Lgm2hBvLdqrEHX5CkPgHnpvdcAsDix29AQNwrtTV4a+6LU3/EWkPy41W/kxi5oURtr7PGm+B97rr
bpSpRUuH1LcFpArH+jKIiDNyXYS7zEeRejv0SoHSzuqXMiVRy6jd5KtsSUMfvRDqEsbxHGeax7IX
QR6CL2fuN7D1wEkPN2Qq5ByBtkCa1KIMuchGPjQTHVnTE7w4MSjHrbQ5dIDxgrxP4q+2WlakzQj3
5hgthrwQodrtKiKfl2V2QbY3QGP1OmqMZ+qrnx8AHGbohjgzhZ9SEgPIsABT9lr91oMIGEeHQCHm
40oa5eV1ccPrKDWS1o4tBTdQ2KMcLCZ/m05gOl5O4drmp/0FBZYkzIE3ykU44YTL66BcP4Xc5GkH
dxHfJphQS2uCRtfPKqIxO1hILipo1OH6iDKyznmIWiTcrTPlwoXxAad6NLeQaqAVzC37cZKTcX6V
laH2aZXZQROlHCkuLUJX2cXqI4uPcupVV9LkgpHFu75HofzstVlSWzPRMpG0+cfspL3uJNl1X5M+
0QB7qALPOckNxMv6wdEZ1rtb9983rLaUJJibwMALy+2nr6gFgwfDnuj7tn6QecBA8pWyBR/4AbVM
nxNoeHAQ7fegChsemalPI5YkRLYIXvE2pPXoZ+vfY2pCUV+w17Jx2hpFJg6YRm2fhjFXokvVyl1f
L56N37Nq/qihXKsCyJ8TB7gDMLe48LpHyFn1lBONAwapIr4IwLRNiq6LsH2vsjIICiUN5q08QzVT
W9Qi5+kjBupQAFvWZ8oswf4c/5CcXknYIbmoE29wR4dpfs8VDoTHd8Ak2PLboUqpaQuS9ZiY8XX/
+nhEoHEgd/ChPgpCcoUdmT0ZG8kXqsUwmX+xIcDCcJxvzamRCZKZwEVNNbsclsICP1tbZV4DlQpO
sIuuKzvDraWIflbYDfZRUb2LY64EHmxoBQQugKuwQ5xFKPgOap0NIF+vYYxS3DNi8u7IB6niABXR
J4APT9TThfXw3KozdyHqoM3pu2OxiyhZVnaaob1zpdAKq2Z/XSZZIpr4B+68tErMPGdGpSygFc5K
awtQPOOvmu4W7n1pYQm8erX8QCyoX4Jpk2/AJuLgnsyTxWuPGMKz+HL4ZpC7HHAsPwD3f0onNIuG
R5vuPA8n5cfoIy2KkIL1BOw++IzbSUn/C5aSYnZ00GkZlfMlgZJcqM05JYe5ZKsffBcEStQs/7lE
FHa8SN/zT81pxmX8B8lBxNKFygx6Ei8nX4DfW6qpt6q3Wv55MUlB+o/akho9u81m+8Emb/YWe4X6
k5HnOiwezp+gshRdzJRmG1il0qiwxgllvNQk2I89v21tcIxtoeFJkX66Cv/3a0ePQMdV+d0jNIl7
IY2tF8yvV6mcKAUs6jkLxrGIcqdWrXFJ+na+s1NyYB8KOfGwcf7AwZC6xeVgQtRzPExg2u6zTPmk
jwa4HNYfyRuXMjrlSjfxrHD6XX1kZH9+M1ww4kkps1jrGqw6j//6F8Pzpfq+KkCX8eYaI3V72vjK
gxZdS7u1ZlD5h6wHBTmtnl4lHdlYNmej2/O1wlLHfB32TBo36RkAL8LtjaDrJizikxI8PTopBQ79
vdI8yGfF63Dk7pIgAzJME/4yg6NPJhAw3SCqK/NKdrVnH4dYDI+tzRJT9SLLpWeIRi8VoVr0skCz
HeZawsx24/cCDnGRSb9QetDKwDqlvUsYBNMjb5flAMjseUcsnAhroO6wVcrISOmXdnniGph7jHTH
zsw9t+ch3+VEVGrHeuQoFclaV7LWFymlsABOW/ASAvrMGdn/iQ7GqqZgPfwlbaYgTW+juEuGVopY
2y8RXxCKpFSUV2KDHekz7qHKf2xsvRnY+1KZ3/NkSp/fOSbBtaDwNXPvTtSUOIvU+Mu5nXqMGuuv
uZBLxjQlLw6kBwx9tjmIbcK0EUh1/x4JO5kIU9z6clrr8MMZ3tuYu/tlIE/4Kf0aH6Qkv5gBE6O2
TpwLgA17ka7kG72BxLQY7f+zywAgxW8z2L5YnCFZci0Otz04qYZQUALaxGD1wY8j8W1i/CNdbOP8
68LglMW1+IqRyDXD3ZFg/L/AjsaAaG6MWaaDPjGGMXdRzj21T7NQFHvG5JjMqYAg/szYKQQJ5ZBH
cxqA3hcpq03Yihbha8O49PyhJ9Q7GqFR2VSKVai4Am8dOc/dcgcpOH1CPm4yrH0fLKugIuHyJATC
V4lRiQUa38Pe4ouCSihEedNOSXLHnYOqDNixvV3YH+iesVXjo8ZWIBXz9DiFvPB0bgeHvCrSf8zu
6VoHtbqIH1px/9GgEmAb9P0BV0k2pSrIbni1VdkJEcC1pJc/DkACZ9OkkXAPxXj3nZ2Jp/WSRS+r
3PSxhlp5EGTId3UJ4KOk4lWUMGgDHiIZu69mn9TVOpPGqqRy4QKPnsrvn3SlybO3WzADJLL/De0Z
QJ6RzNZaKUlPHqzNb9SgA2EU7vHSzlcJJInDkT/GdDVPj7RtlpmY7rCHnPNtM+YBtt7Te41kJkYo
PmlygXzftnIYuLpfxDbgX7O+ba/iJGyg4RCDH+7Zx3CnmJ3NTGf+JxDwo6sbrku25b/GiH/kALSF
qMe1VfVMoyZh9b/af7mCYG73wj5fRwgBE1VwXRDCqgtJGbawIswWSvpkzbSPsWRRRPs7pJCTTY6G
caqsCqNfDHKBToR22BUbNq0j+qo37Sjajnti83JV346irnwmkxtMREr1+SxiBMum4MR1U7QhQAJ9
L1Uml2SeIN/K4YleKQ8RWVG9wwjwwo9i1fy8DPf7iV6uNOkQvRmxyXDmmKh5x2Ix7JlpNiAz5mx2
mSrrQ19ZzBeNp7+n03c6ZOmmxekU8rS3VsqoV4FmXHXM35Tyif54ub0dhR+fAyHDjntbqr/MOLWf
f3i7WkGRzENNes744i5DIimthxEtmX26mcl+mmpWtAo+ZmAESo0GI97Oxi0vSusVB4B6BtYL43VE
Ezinu5yM+JOyiFwa9SoRbApJ/Y1f4e0dlTiAVcfhTEGMCEPFk5/CXRaTWjl266A1W1ELyZFIMoMM
MYZjALQJQa/QfnxAL5N+tTI0KH0QjYaA9yei9A5fCdBF8EU/nIUoNCkVSNEu+LWxKu7e3+odw0lA
jiz3Qe+di64u/Zaqzt6kcYmR2z5gd+TL4Nn8JTwykOPk6LYmfaRn6E8gEnATTUTawv6fC7OpR+RT
+HyR0GwAIEwYZkGWpahYea188470KhywgOBg9NyQiE8JScRi40LzE9pwRunrtm987KKTqFRcXXym
S2G9anXc4iUOUI5nKd4CwJO+NzOjfarRZXT6dkprNpO2joj+yczpkiPEEVm0qKiZVnStYuTevwIv
DJtPaw0kFsADoo33vDA/6Y3Gm2B2m5lcYIKvsVzhFRzudLjZSzstDy0CisbwLA65b50lbwsrmvhW
z11saEsWXSRSO3PLGJZZqHweepdvgJz/G2KbD0kFXcI304qMc/7POMrbCzhao+Wv1Nx2h6etEwDu
GiApHm05cMmkRB8vSd18/+lmFW7eTNqKNsbolvsd9QUpHpee4bnTKnaIfxkXDB7V4XT7/7kFuwkD
6TWB9OZU3XjyPGKlsSwx2m4uibkpriFP/4R9KuPpA2dDmPeOx8SztunWcJUrSWyZ+faWpQmbTaKb
ll0K5lizZl9KGCplVzbFqk3EhYINATSr3fNCofD4c9791TESd+jFwYvG0HPOnkUDY1EOj0nuJJ7F
PDAkaZHrhmursRs+9+KGxHwJvIxJssRm9WaPRlkuXqCpmmNGL35AHN5rCIjORIGLc4Yil8fTSA7A
f6TQJAKd4QNroPE6TjNYxajbDx1zpacI5QbvZbafqQkWfucnDQEU6FK2qG75jQond/WILg+JSOvF
G9FS45mAPD4OjLGP5/YTH7VlbRt5BmPjr0Vl9c7/IY3Ne2KqWKWiLLdKDMbr+YtlTAK+ApCHJxS/
J/ArVZZPZLEyDsWtsP3PtGSqAJ2BxxlrpSJkT8SSInvOt7whcyVYa/pwDoNByumr2jAzcbHXox+y
43TxVZxfRspYl6M5Sg68eNM5QaBRUFybyAF0UA+7WnjqkemkxTzph3Pj89VcDPfjS9ak6+2fIeXL
0ol3PlvYDQRmAo+oMwosDyoG5NSw8Q35IUJ/k2QTbbAHpjDmLZPkSmivqsp+Q5Pp0nQIlRca6ccF
gEBmpHzQp28iwrEMNnftHHzVKdR8pJvZIeaDttVBTSda8t5DnLli1OsgJOmHw9pfC9vr2w5P8viG
DH7HlSjILRwfdr5c5oF6iRAzV5trmmPbxw7nH1UxR9KChpvOw6WP6Vk1Tpk//toHUbtfLVGmKtKw
ixGc7DPH7VsoR65Y0NwfgXRNBiWcetDOu2y2B5dF4OrLnm4xHocIsGQ3mcW0w9l0Gz1Pcy3xwNwU
YPtghvPngKxYIl58VDkIAdYQysS+WcG64vd5DLWln2E+591XC12FzJG4ZXwsRtqCeyNpJayWSniU
PPzdWtuRreS6wDp1D4UI+IR/2YDH1d4WZNc3UvcJjKCmphJJKK+CqxAE02u3vAAanQaA7VuG/dve
x9g+53wm26gN0j8G7mX7omA5umiesrbVAn8XSHYOoM86aemGKlDXN32+OTcPIGhqCg2lodgkC2+q
AbtMkmongN1diUnSRw3X8cTPI3XQ8OGwgTSmMz91M1Q36ILNoXGzOXvjIJUmTXklLHRdwNtKygoM
XB7xhLmfyKxTLjPZxyqU9uhvopBf7FbupcT7LUbLmckpGh7nBBg/inl2UdVEdLnMkOMe8yCQKYiG
GCAEnsqId9+J7MApokRMYtZ+kIFeBlzKn5bO+P5y57mu1Apsx4KaPDyGIP0BeZxf45F7pOV1Nl+K
BgPj1KaGaRSG/tR6EHtgFcViIhSRlDEqZlyPdhJNHs5MQmaAHBwZKpKQts/icy20QKKYK9ngtwyH
tDUhSgc4TXqGu78zt0sPp2LUyUQTbUP9wuvphPGV6b7m6tRQW07lqW5itfMZgjPZlmpRVh5RwgzF
2dwS/aujSYaMW9M28Q4bH41forS12Qq6F4hsDWhr6WsROX1qU9ZOhzcxLUDdq6V06mfesLfS6asL
2HYLbVmiKNfbjFZqOR1ybzqXmIvMcAai5MWk9CNFmmgWeunKKQ2y3Fh3CLSKDJ/k9XNGJ3hBWmo2
ieI/VLqx7n157xzD1VFNoQcKU1+iIqEqXnR/Ok1rVqFITV5yWh54KtCEwsRwCdB9Z4HvF/q+b61H
YpMtjymUqp8mVfbAyPHKOa+DENJ3OzZNOcKCyrqdA0XOudT9ntncLTv1aKAvZj4u8ODA+fePBl3f
nCiPnaaFr2S2BvQa4y1/FDHGIS40YeIuclMJcxernJjTq0TS7uHTtAz0Ai3Y5LGqItnBiSCwx2eJ
QfVhEl4wuuZQLPuobwDYEC/Gd5L73sZnsOXH1a/7b91Pwb0lDetwDHnYMad0RoTeh4L8B3TsJgHn
FY4cYxIbENhPHB4TST2lUMG96+w2qU4m2NvIOp3RnMEmN2McKGKP5Udvyc99/O03M6+wcfud38kV
uQUAlpOJTasI3aj3siDXOtLdlUDZ9vkCA4fZjVY+4vx0yYUBBgpYF2uE9+W/i/jskEhorbEEYge0
WAaF1kZ0KG+BQDxUNd2Qw/hU3im8qmjyCYgIRAUR33T5qXRZP1MFOl76g+euMftpl1nNptkF7P/5
eFqo2xsQvprMoExC4XZ7WnKalOSvFIVRjrjnB/Mbn+k5DXk4NLjmTy9uhFdjViye+Kt5Wl8VNujX
iD+PjVVMUQCsorBoBVPNs2ilvpRpvgpQplecT2EnyMWLvSNUgDpc25ptuXXyioiKF4Fu0XAaiOSs
Ch95L94j4YNjT4V7j2AWghzpYMXTEtMaJ2WRjoAkZbU/NPHmeS0w19YzONNIPvwHAA8uZWSUnrGf
vhfuQPmrQOEDQNolQuX9IGdKMAxdFWkv6uH3uKD5f1obnGYE3PQB98HbZTLnYnaNCPKdSXFu+jOT
RQ5anxrzHTbdoqYuHDplGCOeXRvHtbTwogLQlcnwPm4c27bzHDUUcn+Qn2+hRkPRJvI1W3oYsiSl
q95Xpxjy62UXqYqRs0jd2GC3BqlO1yRWqLFpN2K6ADWo8DXPUzl0zfGlQERR5O77CvHyOszV2OrL
Htn/sJajykvXDYhHCsdTvKgjYERD3GIEi9Ki24heDdGDdzXtAgXxZzEYO/8YEFkgQYKa6lOzSiHY
Ax51A9wEI2acgz0zFaTOyupjfy/aC68M0dl7sW3598UYsrp0SwTU1sNbjAtueuYtzBRpj7kWXV/S
IELtwHpRqnUIaH9Y7Prm2KPZgJCBSy8bL3vofHNtLki6611fZSEraxnnaF6cFq9gDWKXSe/esmlJ
GkFZO+ZDux3WOkWEYbjDGdB2fQ94yqGfSwVrBIBxy8Aws2GO/Wmhre59thyn/MSjKNIRFdPUKuli
JLhzQL5j2XwEvQmb4Z0F1hHfNMttGJhuDpV7PlMHOS1PLl8vcUdFIbyvbv7PzzELRc9wYQHOCl4J
K5OpML/+6WVc55+x2DOL4nBPhohCfDSJtN2Brg7mfVrz/LzEryzP/bS++cDxM6QYx7zVqWFBgxbr
3h7IgHC47hNx11cMYAeLTOHwuSXeTR6d1COuE655Fq3jRNnmxcIfmiH6/XG4J8JdY3O9eIL/d/JT
JfwIFY8XUFlLNp5dO6PksuogAeRl2CXG0K9zIHZSWDOEjXauO1rKO4d6AykHHB4a6V/V3dnF1DPh
VJme30qpQLR7DazOISiLX3gyBBPqFhFH1aq4xhkcQsqI32n1lY1Qx/yzESwmxjM7WnzjjFEmWX6g
OEbMFYHY3s7aP0Lp9j5K/0acalNUAutBs522fiif2O5ZqD2Xdoym71ZqjmdJd6l9rmLC2c16b3Iu
J+0Q+MNWQ7eDgvehMnLXdZYasgSp60kVhvfp2GfPlQYAPnIQakNhNTKqWiDjh+7x9ypzVkDZCkny
cu6O9dKoBauXEIwEHI4i1M0lrVvzyISB9XF8lmqjTkCSBjxkPVTkF+C8bEMJBg8V5YlzngBiPXpM
QoKNTi+Y/VC67IOIcTKU4Ajb7S8bg7ADElBGE5Q84onB82Ero+3fd6tzGyFIJnqhKZ75AXXU98Ok
90Ctz57wtOtTjAzfB6xLFlgZNBNFuprxKYTx+GpM/UicgfUfYmAeEg5nuZCJkNdmZEOwGLkRQ9GE
QtaS8kVUERqdSXGw8Zt41DuYMmaJqIfE2NX9RsbBK1pdRURX9zJGnGjqSF+YYyXm+nnGCtzRwLHl
UFRes+30tSo16TT8C9AP6Jn5CgoTiZv7i6Li2K9ElxT+I9ah9IGsgdkRIYlkyEanLCEGFhI2nckt
RNBBQ71T1MNpuwkth+Uy73s6BkIuJqn2Gqow9pL/GoKqpaRqL2IoS2/NQROd9E646onXxbTINqAG
zhVNDy2/eM7TJ490FUDQKdYmjR1iKEcpo2zNGXLZF1iKmiTD9E2cSIRo+NrIfUDcCDr/wyuPo/L7
frrIVYAgGgEX2MZcuLy4DPXH9caNvGQMXPC9CqKAT2e8OxYK6WE9tRmydvnTiV3K3LsAfNzxkhyf
BVkKEjiEbC8rDnn5S1OVxcJomkwrPB1LGZlIBbJo0pc97sWO5BdQSclFqq1l0tUuKH2mYwybNgwd
jkt4c3SebPCPRCczMicKpVhr6+YlJKUc5oBfLgqCLlraAHXRSZ4rMtJ57iQI2GLqwzqadEgzJq3N
aPn0a66FqzqXY+mHSjDIXWi80JhzmED19W+XOBAIsXYETot5dICnWqHc3iPaoQiLDwcenIUgI00m
Yf6PqaLKLKUTYIltvrApFF/fpSc3K6rmLdr7h7P3WPXlnRCnWdOt5HvqdiBZXD5859h0f8BlUj0I
ZlCGFo34cJthSCaqPvrfe9AQla8TyDGendaa9NXf//IGEhE79jg07xYrOQXF/6+PTsaH8W3+4IT9
SZZYMad367kNExBIttt+uwjOd3NMfPxUrUlu6U5WcmbFGnyf2VZP8clQ3Pf73lZlFSQzgznRUUVT
KeVXDl43a1yTTfY4Pgyn0UltFgtrMCUaeN2f8qZZ7lfNdl52ejz4QU4jdNqI15TA2M5yqh9LbXt6
xs37bpRm2YHxmIAAOV2jTFNCpyWyxObZ8LVJNsHRPbMnISaps2ZqKVnonjpgemqksid7mrSi8PoL
lhYNYjsnpCItCge1/o2Gi/PHlZ45yIMoYOi2nYAQXtc6cAay7WEDzqHe2kcDPSgSseBOyIrzCDe8
wOIUGrCnQU8Fkk1OIQums1bnCqSj37E1VUy87u/54aiQ81r+NEgUmyHO+wFW2BuOaMebHGZEPZ0H
2Yliim4h4dU6rCqedxJfsupPXMtfTHokR7F3Ni/PRRucKF7mWTq/se7y+haS6a6ycJdARqa6F11s
FaMJZ8NoNrXTkzZTNrNlrKTozo9QiaaEP8ilhFn3WwqTWoiGdT6bisKlNn4FV41xaI3ZHNASJPUq
ug/Orlghc22n/wHLQyImkvis2aUnq+mp3jpIhcTNOrq3Zwcg2KeDr+A9lsPm/QEarQIThdO9CfO3
BV7jWyqDiRpGIaatdSKtUJLVWOgPYV/7GIudtyQyHMm5wZRo5h3PIfuqb6bSc2kF8gT8doexnAcJ
DMjrmIm6AwMVMSr75VrBtW0uaCN2KsOc1XmhoRDvEzncn4IR3wAcn8WWrD4IDOYCCh8fskafpMWb
uNNgCBKMLzXif9/u66vCVIunVHJC8F4/fdAGbjg4Z+qWXlje8q6Hi6Ep0GVtm4DLj5r8601Q+zoX
eVNZoQ+4oGy4mBGxUsPyN0Bfcgc9uieJFTGFChAep75Ex+vYO7qZwu4PYRcenG+c2o2dcZKGjp/9
tNQ1aGHtjqGpAi94pA9Is3wJzt3bxBDvXHS+iIU/+7IFglyfYRnw3sF7npFKavuUdLwE3Rz0F+zv
XYIR+OTkl4rmT/Ybs0h0tAwI2mW5m8arqiQ9TrB/UCgl/ho+NWllWBGplm/YXaaDqWjKWYfLhyAF
iepqDHKWx0YKCKmZl1WLUKpyh9LLPiD2/RHcF+L4oyF2LuyVcD+mNm1cdO8SY+RVNnqsQJ/m6oHt
LRJg5Uj//e69SCy4t1eN8ZXHEFARuUduZKoCO0EwB7GTAchRdm3CUBHw6ONmjHi1zsK/Sp9cxjri
fxfu4EMMo35qMEy8lviVHTBwGlYW99xJ9ljbJns8h/2Gh4TPW/XjmgS1eXiK0qwkdMaa3iYGrXJr
D1/awSjWlL1Lk5+rP/Srw3FieH/FVFcD0jco6F8vlVWVncR3Tyo5fg+XKMuue80yp0pJ0Jec3DBC
dI9rjzScL3LbM6x1Dyd1RXZV7d+CbKBpEBg18MYBhGCgEoOMFXp1s4bYM6S+MghSWprGBRRoFtnX
lhDNWKChdFC1iVS+JQOKdDjlD0hK4Wpw450urrqaGb6OBISnZXlDhEGWpnex1ITtjyRWZwnQa5cr
cawDF71mJ2aa1zNEom+rtThF/kIXNCr8WtH27v0B/aWlifoWEJqMFB6a1v6qCzWDwLHGq3HVgjJ/
GmZPRY5fdO9+zSwdYunznT9xQbC3tyY4IEfOlPwYzPvte91/Zp2OIzUhjvRpi4n/NLsfvQeK5PKB
FNLMmQ/6HWIFU9g6aQNAgqFJnx+RjCD1buGsEsK7VxSz+6oRL1IRosq4L136d0u8LPNTrZeXcAxh
2gLpWPoARB/1IBUsa7xmPUooR7exbiEFDfUv/AO/yMhjyEx8Hkvzr4sRRURwSJmOLIWKS+NLtlwQ
/E/469GtEK+0t3Xr7m8Zowjroduyq5eVyVxz3av/mZLPKTNksZewKv3NhRudyjBermFIFBGaJQZC
iPccPv4Z1zdl92+nmHJ9qq7+ahMgWBZ/qfdmOq6nXAv371TBYY7/e1BNcMi0zgxjRFLrXvYe/oJH
a78Mj/4qjENzpFJBBax+qut216qEcmD3+db1OY61U+frmJiaTFXUQqBkVrzdEO/jsvMuDRJEEaEJ
QsfPAEEU/BUdtOgEFiI/0QG4K3uzJLtLxHX6qvHBlMCgNk30XGkbsVNTkZODNYIldH0UGljr5Snm
YDFfUQ5W/VUOfJYW+6VCmYySaOi3lxt6auGPdNU00vMNDBawbo9eSX1KurBO2TilbO4VVdGvEyCj
wmH0Rh8BvLcZqUv+8cK1s9oyo9qB8of6OiBkN3kNSrb3+KCW+SVaU93Aj/IY5u1/qSC3jrUlgC6o
BN9MryJXuDlDjKwMseLkkqeCrRPXlpImdZY55F0a0G0u3XZ4DcQq2q6V69cDV2r0kuTHlLzHiP4V
+6fVckM6mwij5AbEvGHwLeirMoQrTQY0DSzmdkjiBXFnjEmIQNAJdoite7a6gt6QxGV/YntJamKT
tY9Ok2SB3eD2516PHHNHETV8PBu27TH9ssz7kCH8NoDM/XDwLisr59RgWwBOwCoWhFHcR9hJgksc
sso0dizUhQGmDzu1d+Vu3yzWkSxbe3Ym4Clko5jE10DR8oNMmkykY88OVdpJNlk9YaaOh/Pmi7zJ
3rJB1wYFJFThNkCqpzB+AVgz3zUUHu8GdVz16z2bs2xd4uNo1Gvf296Ejk71MBud63v7Lax1ESrb
yboqtZwnp/KciVBAABO1PY3bpee3+51FwpZCJdS1csZUt7vBZUA2ObPS9lmomHqyvrQ4a/ZciPLl
5M2ESpKmdEAsVrEOhB9RpQ+6R8QVlLKZ3nMHeTgwBGCxdp/M/IAtiziAfZSi2F/RkFdq+lq409r9
gex+nVwgu7VZMhVLN/boodozcKqY4LfPSFGmZRZX5jef9d7dGBHoGI24EHXkTB8+9Kfki4/8ZRIc
rXedniL97PmMU6Nw0qMLKBZAbgUl6OxCtTPFqykxhFamLEJWMaZ5++J0pCK81Z6dUz0F8/CowBCi
cSV/zY+vez/iHe4B1cuYU/bAXFN248PNFMvStucFjGL20nE3fsHcjm3kwvvGgN8RWiCkBjJOT4JX
gq4HKDdE08T78jNMT2gYWSWPoWjsvUfilRmdoUmdpQDzjQ1isK11NAqr+IEfY2qJXFGv1NBJz9Ab
BbHsMDqguSQ6Hq3MQJD3D5H3rCw/HCaGOrKGmTiVFKDTG9tl9cJ5GkDaJ+uYkb/kxDIX5uKNrAkU
6YcH+Fz1ooVJ9FdU+ld8A22JM2yOw7wFdj1SqACVY5QnOLXriUVQKMv2NOHjgPT0GPiopckHcBi1
ZqguliGXlXJbwhBy/7GchqFdk7yAZywNJ7YB78Ji0K+G9tXqGNhPA1cTZ8wcy9BVDl0HSkomZmVw
moM6MsMDu2RR7oitrlu0M7KSKEWnHd/Kh3c0sGCPO6CmjJ5BqW8wzqtsEDdLChnjHXCRS+zZ9xmb
z92G6l2gbKR3OF75J4+Is7+o5K4Xpa8UpPAlAaSrmzsZkyNu5i02E3kDbfTjfZcA6Ms2qmiGDPd5
LrOirO9qnBOwtl7p9/zSF8L7clI+9xTibRbu8J0QoaFoXH1o9bHkr5tppz9XamHzZO+t83WgpR0J
+noSf6znzD0KBxV5PqxqHXHw/1rIW00hxR9zJ7xXDUPz3HhSyYx0KWRcyXfV8/gHsr4PY8Wi5YS7
naGbY3cCqxp7N19lJ1xvazfMomIxY+lp4L3hti56gfycgpb3lkEYCMGP2nWcN6FrbE2OmFi3wRXf
+DR8yJy+bilMHtp/R3C2gbIPJF3OhYHCV/2cHN7ZIw85qs7f9W1H0IoAjNJ7jaiBcHZU142T7Nr6
tIzcjFH/BM3O7OX8GD+drNXmr1EjoZ5AsiE6aqfLakUyiD5OVwFGksqOzbRP8Et1GuC+YvugCCOl
4UVwKz+GGZmTFhUP153dR7LByKjrgtInssK6xz+5TWvRgKi99wMWPXGWQ/3ZtYf/jChFTT1FP+IX
NTQBHckOqYsUGjY0uOirnGSbY3itTsroH3QMSjKz80/SCfyTi2uxfnRulQsdGGRBhLzVUW8oLixB
mQGM/luBlNvtNQlCZycBvNlUlEKC0jOlwgjw/SgG2ZcyHchRoRHiwSTl5762qzFTxjUZEGXZmnxh
3841a6sEJP1Ptn629qNg0Abk9p4qwjJrIO/bIMTMVNYKOMsgxBlxPfxS1t0yh5YCAz3d0ZlWI8pp
XXACfsL4X8lISrzPjJGGob/haI0s+GTX5FK13jbjD6juspH8gicC7wBXovnxoOEx+wJF82A8MNHn
bwpq2Glsa+Eqvr46VNyekKtWzQdknIdYoahTi6MoUA/ATCzDSBLwN7nW+YBzXFfekwOv2hIQs9+l
Gul90fJKwrc+LFXithKfUU+esKanUpOs1qjty7ETmIRyAyVjQ6o5V++7jknIC8kcG6uJqr7bxosk
2lR8t6C2T8v78jfYxsikVqIer7UC4NK1818GoackboREd8HiwPGX3BIW2Tt2xNeeUjMf9pmA6qFe
/MaK3CR7b1VsezeXUOhPhV1Muk6gCywmxpPOXJx4COuP3PXK8y/h+ErFiGGBjt5us+AjNnFHgkde
+9v0RwNL0UsWR6tmp+f4HF9t3QUIzGo1vcjqG9wjNzFmjyiBuzOg+DsGIJrMZLC7fpcbHTMRmHAD
x83O1DYN2LDO5ztbj55SVlmfopIGBZSmUzGV6VJfw1E+d0nwCN+wspquY28dQeoY1zl3ktLuNRN2
0Ae5ZRPJLb6g0KI0Rz3gqQI4/sbBS0vLFzd6PcAcu9kIRdJLygYheO6nYqirXZQokwLby/JNq0o6
uUlASJMAiQZJrUhn8ylHslxVqUQIaRk3mTFo3ti3oooq7n4bI4Sxj/INdHaJBl5SYHxNHtw8h+Uc
3zaUpk5VUL+RREi8gYLyJehS13fLN6K2Un5/zOX2+sIFR1fYtegHNr+/TMhOY1dOSFWFH1/B+ds9
eskS+kwsircJ5GbF3tTnWn33cVVL3pGdPqvhz8xVPlZWzY8xWSPsPncCZzQQd+ZzVHcZ6IFTrZ0M
UhRgAdZ4wB15ub2s8aE32ockbv1Ussyh7pbMVBG4gRGUV+hbxAwf79InKJNKYVElc13RKSQ6wPTi
4KEcJ/QcdwV5eXKrov6J717wE2k8CB8IMWe4nyJquggbVqYk/jlLqu8aaIISQd1y4FZwsnXY9gQz
Yb+/5c2buS1InWEBKsKdqlcXC1W4ncE7qCHsDLLFs7Bp0aOmshOgvNYiJhghlCKV7Rf3HDtsg/qU
w+wV1aqHUXObN9h8BQNzg6Lghq3ncfQjtT/IJ2d/1cXy02YP9oMeXSjjA4GmzjBEtAWqJOD2tl0R
aUIVTPaPkZXuzWBpow5GH7J82EzCIF5TdsEXGzRIqUBtuNdm2q5ROQXW8RNB+bNL8tczaBR6muT7
+LNHCx4W2ifbsbDuJdawkuOc/4iUK6HEKwoNmVTPNtWAi91oLmedMpHs1+Uzh3aar9p2hlLWxlR3
/x4uzFHJqKY0KjxCZQqUg+5fSxMzKFmGQjla/AJSg0bRjEZ2qjKXNKy0/Ss6OZvZnwmpqxb3nREQ
sCzHLV/Fcy5gRTx7FRSZhux28sLmv7ubZpvsZeOI7giwGXiT2oBwoPAeqmLmY3VIKeuJ9tw8CgNf
YcwgKGqAi6CbPUUVboijynyU0N8zH4XBxRYRRItYCDKypfeKrYt2D3OWVLX71ylrhF/67XxOIVsJ
QZETYusnv1+S7PlFkd9GyVxBvRfd5QUk/0hUs+Eb7+2gk9ZkU8DgUgxSp4ohZl+1KSDNkajnpePf
It9eG+45VmPVonzBGXberdkC73Bkz9RwVtgBLWHjBMNVUhwi9AXFF+Z46iD2Qzr8kwU4djdhdWUj
x1D8h2pt4jv9yLLQ5KZXZ885xNr0NBSy5sb/SX/sJ5pzGXoi5doh2ZMaCOcZ+HHTf5e5lDxmwnEG
iF6hdeYdP1vccOulr4TULV3BIX/4IVFijv6SuZd7UPOxGi1l43Kxo5HGwUVNicmmTJR/QKqSSmfU
6IZgO640vaWTsixsiY4G44zIwaCMpnMrskdE+RB/5rY5iy+KvdLT0iKU9ctFgrfx5MbNm/mMUQLo
gOSeU1DWYmOQgjg5B9Umxs36wZ6IOcQNoojsh4KO+01kcVTq24UxF5nrjBDwfD0rHZLS8ykocpi6
ERd+ZAzKKx8sqmc6WE/kP7AXfHc2oa4Y6OZxxQkkN2dytNvGIAp70B+uL7FkKEX3FMVtsmQQY/sI
EupXJVyLat2AUToSNuZAa2TXCHmGpXLdN8l10aJm02LDcXT1YS2ANRSX4oddYZbSZZ0waC5Ygv24
vMn7K1qI1vhvwxSoKhZAh5DZ4iuZSYq+Yc8aiLlWRqPPWPVV5NoTO9bqrv8IKHnQ5L9D1kK3dpH3
8oo/1s94ZuKtMEvLxfnS4umB98ZlqSDaqcCgG+DEw1CAVIVLYmfJzqhuqq6FmySp3cuNbkCqWYo8
RcTz/sf4WH/VOEY6VvM+05yMTTfKqI9Or+tKZ8eLvrE/nrhICyB9jR2LPSmSOEff/UOPrEJK0oAy
0owAOovH+pFm0hbodAMDalYMauhc/Qngji1uL+i3BN950pS/8TgX3DmC0deZcDG3LXaJmNDKof4d
taR4iRFyagAH8FbgXDKZRSLwkUMHrURSInETvRDWtz4GeVga3sDPClZXgPvIVPoMQ0U2aWirLjeP
f+dcbASAm3V4J3dtgblqibnc/VNS7Wl7ke9HLaTbFcNdPFEPG/ch+iu8BPr1+irEYlgcytVTe1Qx
sXl4Rdo4bDtoA8WWe3KOIzrvQlfCHLd61tkOvRdQIsyI9RR7s3P07Fv7Sggk4zNDlk7pDUE636un
KxNLzQHsCiS8Jk45KxC5+0ZqOqeKEYnCRunnYwgy9Jw51Zt0wIBTVXrDGiC6emGkyugi7LEdmA9L
RxTaz5nyFf9wyVCG5ztOlirC9KK7f0hs56msfyMYArZeihfhWOIpSmzqayz0hN2difCeZf+z69RW
xd00iXQt780N4Wnq0/XAzxrK514nDhFeG/oMDlEv8/HJHb/6AdTdiGBoUEZFxochdXSn1PmWh5xA
ZM7ggvNvPPhv2412qnx9/vmkQiAyz9nG22HSmFj5oohPLCzUXu3ahyCRg4Z8Cr3k+O7UQiYAynuL
Sl4euW5Om2SjohmoiLz4AYGlMbesbGWrYc9EKgm71vvcbQCBdvU45Ezlh3bJeqTEHDf23/ztg2Ue
55e8IGH1My86SSv56FYnwk2leIIf776CE/vYKpRbRAxZ+k7x6CqzVHm4U8URNOSV9rZLXmf1o6hW
6kDzE2F4p9UbD47sZxYVHdqsyZ2DHFbaI+//odBbfB8uuJ6QoG8I8QcU7eUH4IM49y5T3/hFhsX2
f5eEWbsy1mkzpgi5jgP6efXz6D4V1V4k4+ySYX1FPPVyhqfc6AVM1FaHRzm0IFLsBGhqWfLH6DzR
r8XNAtAv71EEWUVNQ3zfNrxe4z4IbQeQoP5wkzLcTarKagXo4CrSQsleAdSbQ3tOjl9MsXv5fMcI
QfLK5mC7VQT2JnBDoQ8enS2w3NFe0nEGtmz+jNFqsDDVG9TYwzAjHTN76uKxiOaT/Jy+6ZysQXk8
d6CsreH61wo43PbNYN3oU5LqeNsgIAfyVpNvddmphtHoDbMT05ubqLTho7/Cefv27B77RZ8j54im
OmvEiBMp90liSKoz0JDPpF/I8h2aIxuiIcJXe5ws9BC3z/foBljfuu2Znfplf+pdvyJ+U4NDPjvV
sPcye8EqYJe+eYX6KHWVtWzgE50Yv7PEf3I8X/IpXMeli85ByRxH8RH78qW52dW65jXrzWVUeKQP
SrEyGYB0uz6R7sTLKGpQCRQWHR1L1E2b0tsU0MtuvFjivji5qyPT6fC1kDaFCSUeRBWGJjgKFDsa
uxvT/9b4zRYQSb4ffjcmUUmk8KiRtEOqi4VzWErjz6JYYHtLQnh+Sd6ZFT4hz0z6tR2IJCYFNT7R
4Lh6CFPYvnC3occtAA1f2QARNvRWzadqvusM/W1kOXAHxKSzTfFfkhlvfIPe608xJyoRiG4wSSyg
CPd/0jOSEEqhCttIdwOK+2b5JnAuowV4GEkzTkk1xman3a9kiqgQ4/U6Nj+Sw7KFe0ZpZyTqLari
J5Z/Xln+fsLU332gGVAjTzNE9qCFKeZdplUYJDiMvo4xl/8OjSiqBIh8zXo/qoWSuFEyIRiNmCwO
/+oE3CIkvWb+J2050jJN/WLHxmqGD39QMEGM3JWoDq7TPOTLiU/izeLCfq01/sNKvzqThxJ6kB0e
xQuuZDkS+lF5yd8XaKpey3tlZvjMmo5h8Yb8JzTuj948W2AT14B4AXEGBhe3akJdwpDEMTF55Nwt
6POqvtD6s4p0Ep7X2ONngXrfZsvRVT6ymRlpA2w3tVDWgJYelijVYU/du6wFl2ddosr/X2JF6oR9
H+OfxcwN9OUOxqLhBoLOdIDQlzJqhO2bFwdt8xUlWb3gQUOdWfJrHIIvpWrUUb56vuUJQQH8hI94
rZu+PLOgvJj0eGVKpnusHcOyr2aY42oC/hnU2DPH0HtEE3bG6BHR1vZSRoFUnqMNCuPXKcF5N4/C
iqHNOIMaIOxp+iB0j56ju8JVNmHsex2qQbgFcZR+i1Q93JgkI18EqJ7/wzgTZglh2LXbkiWLSXj9
XtH9jSfOJUvV1XNEbZqY64IBPNOjrR3tQk4JtZbA5lS6XWTRoLszfC+hAv87w/Zc64QMbNFuuEDG
Y9zihycKTwY/2xyNYOBteiNAvtC1mooKMORsUe6QTASC7kYPx0PsY0EH2fHlsIq99VeI7w1o4Q88
l6+rBx0qBqCRkSCPiw/Mcb7H935TkecgmTJNizugGTRRswaCfwYcsaUUDKnDVdn7XpBVTQWoo36p
Eu9J+NcnLrvR6u5v8DgkjuXI8pIBJd0ns5/7MB35848S5kjdFPkQ1H7+xaYhzuBKkYeus2cEZyo3
vTB8oLaUq+2ysD4NZ0PqRmgqFEfhRNEB84eG6kmaE0LlK3U1zl7fkf8towIxliIPyaRsgvTmKF0A
u3PkkwstqzDBdJhqpIk47ZvRlA5stYs8n9bK8Z/omM4nuUU1Vdevg0jOmXarJDwdtWQh9O1KJ/qU
ZJnY/JdW9Y9piJJR7NHA8GlrFDmC7RXrGeNoDmuKbLXvfsUCzkhSh4qvdg8UljkWInKed10wmLlq
fcZhcV8+JGJ5xwHSpJN2o3oELwu3QeAtOV0ENtuhirXRLrmJ95GkinpUYsWNaynZsAsE5ZhleDzn
cxqSzyel9x8bXMjMbxoV5HE7JsTePw7Wp9AeYhW7E+GHiI3ZkWLNIaXo1af7Yz0KfvqJxCl1y+mT
Vh9Kfiw0EIFuVKWvmbm8ZlfTkNrigTE5akRFEFUsli3OmZ2KvfAXE3AJnu8NuH/SbSRYeXh+8b9L
Su/4ZE0MgvrfWaFXkNdotg7wJrxGGwu/hwfRhN0B55I8rfY2jg6jbxdfFbi3oZgyHdGz/INjcNyD
9cbVIDBxinUMYrdt+D5iG33zsrQUZJ1HyyrD06/7dZmKjd6pJ30ow+5Lsbzv4abcJDubWgeSglGd
MhOwRKM0Uw8YHKd9C8A1rTlwNLH5YEmmCq8wxyw2SqWU9RCfksLkxdY/JrGSg816OSJMuHKuDPpx
3+e8wLhk32DacH0flfrULglHUxSDzL0PD7vQy5s4zlUPD5vZUcMJACf4unPTLFdeUu6nZW2ec5VO
yveICpduenVTZpTB+bupNL4ijILo9/GETfeTbA3i9l0L0kbxs0pY4G1fzK2gPBoJHL1QiYb1n2Sr
+Po8ZypzrWZSkploeAK9mF2XKbTDDHTNoEbNPlH1U6mpkJOAjeYodYAX+/EUnL1ymlLcQm2TLl3G
I/81o1l8Qglh8um8lUQULOCDfIsFu6bWX2kXKaaKaeGf9YB4JD6HRINJF4R20jwIBGqikjP1n4Ui
qMIL68HNdWP5+Iu7XsIZ65pCcZvulrcxt8S3+giubTUkp/0V54P0/AX08ZyHPZwWUdBhkvNZ7vAN
rovHN9+Q8WbN+q1dtI+q/DRm/3BtWYgBCbObGBngIvbtDsLfcSfEDBekhOTZnTMzWlt/07ktLpsb
WSogHtcwFiDh6+A+3/aPYR/O80oJdlxwh7BY5PQxxIpUTO8ZNLI6tYS8quQRQOVG1XkQPkvTNU4T
jDaR8bDlfOvPEpwbijJq67uvSLbGjsXOP2YeRdWey//6SzW0iwyck3c+lMpMyaP2+e9Lpqb3jKTV
h+FrsYvvTKlEBjGJ4Do5rs5N394cR8PRFy8z09o/s7gIj54/DTj6vc206m0rcqqsqh0Qj+zx0/uv
SWU/qx5qQrmv3pG6TIzDXKRcHdUsfc7Ickb1+LJ0zTSQvWRUZO62oWcjQgvKwcrdSyjkkiFABuMA
lvFdGJG1O7ZIXo/FWIQz6X9gScdYKjeEbN6iBqnwVtYaPgO8yFcZTZHhastJo0w8pJDuyaJ65Y31
78OvijdXx6bop8XA/MvgZaKHXMcawmFk0ySk37WOncyhWdjLQCfUW4fRIgLK6mmq0hBwhWiv+pUg
JqHQeYhMtYBEVkD54FVKt/iy7hyFV5B0ZfnqKwQ7Yi3HlxjVz00zjZG5UXtNsG37vDgh6flAhvZ9
sxZJl6tpgmbJwycB16ULYVtZdqbi6UIRLfjj0j1hkX0b4tLQmg+LwJNXo78gsqn8OtUplm4BJ9Mc
Kstj/k4gPlK30mrvYA8MItj5Mr4YyGr79wM/kI8J9PUIJWDwjYTBWJyXPslLbTqjt6tR62RrBCMQ
R8lWRI0KU0jRC5gnbmQ3QL5kwMJBeifquxqB8LORvPSg5NxRK4MJAbGvXVlCLAteoj8eDxy90PlJ
CTDREtDbij0/hEhEgS7FsqBthMSLTnF6KwWqc5yhD+8Sv+HZyv9mh83wFIQzYbdNYGmBf8SzcbHW
NAvlTP+TzbtZAWJdz/1bG2CQ0q+5Fulo97Bnm3Sgt56teu0kaHLlecJoDHQDZivB5pM1vBWtk9Vd
x7iWfDO5kOx4Qs1wHXV75gFilZ2oL02ON34wBx0PGJ9+CCacqdVz6mWHbIXY5Mlg+ankatCab9hj
tpl8OHarhZXpu8QBi4Q/50GCxgJrotl9Q/herlEBdf5hg3pHwIn9hwBz9px2udkjPYi+WEIVAKy+
hUhsz3ZxxHbBk1P/CDi1Z8S0HxdPyIA5mAA9qxcoAvSsSLV/rjq7mfo7Q7YGaqSZzyWAT9k4q4W0
x/6HPth+wHJrcEf2zOwV6Y705Z0w9LjcS4qWAPpJNVBzTo7QM6Z9XCgYQ8VmC4Vpgy54e4Q8XOv0
GAU54ylF2XTHvWFe7/YeRxrl858XrCsCjJPzRsqy+Xz/tyFNtwlE+UNs995rdeiHJB//VNgboYyw
qIvrAfv+C6xvWesCLdO/ELRuuQXdXclaoLcEFfRGJu9qsnPKWQFUQdPucoRUPK6JKr1es6k0E8QJ
/FRT9/YUZ9R5AHeufcBb9n+0T440JVWgr23Nw4urXlkTpAnVbU/AGYs6TV42UUQO4g2xg8i8U2MN
4QATywMFEP8orq04QvRtVwxEVkJ/uFo3ZqwUythUSDCglqp3cKk3lOnJoPwLgk0huGyinx10+zIs
35hItyykCc2qWpAYBDQhxSy/smLKCP84WwrwT3HaDVi/cw8WkIlJZ1SgysUGpJV4a61TBBy8C/mN
lP3chpvaNVMgazLpywYo+PD5VsbKFlXA8plXDuKVeTmcATlIwmU+VO7BeOnFuyQKeiYViRGT60s3
+WkeIIy1qOrnELeJH/q+KSbGBitAUpYCrBThkQHo3wgO8PvjdfsXVAd//wrclHEFjHLSNLbIgVfT
L72/BPK9URWLsU4jDVPuOVkcOr9+8tMLdjWJ68UUId+IhKb6dHXA4G8Qi4R1m6f8m1ALvkmTI/J5
+ZvLZJNdLpcQzVormeGy2gG6yjbp5Sa0/GcH//kulIzADfwYKWeHTv2ecbudcEPlfcFE25ysJ6fb
FWqRRZ0kOcE4f8oM+f7XcNJINnc0JANjfYy6qYHy3svdNYkejIHAtQRZK1kaiMfQQTV0pc3x/F5K
oww97XCFCwsd42lP5FYc/evHg02OeP4cTpNcxNj+yg1FRNC3XLX0UX193ZHnHLTL49ycdE0Cq/0X
LLbRMO69tBRsLOggB/qqXyw8GU+bnijsf4fteLRuqvvfJtzA0tXjtnfCTi1fGYNvHCyG/T6ieL1R
2/dmBFsxStT8hSe8gZDidlJS+6gy2tBisQrxEbaUA4K4XtjykK/qeoivhFKvvTmaAQbyLKtKG1hH
8auWgp7HUtyCvmTg/xbFIctl2vActMl1QVWxWvzYtP1i4BMTfAgucQShpbgmnulD9WsZdFiHuoFq
VpoLsHe4WYHI3bl3fwrZoryvSwbM8l+cIwBv0Lx7QjSgq0MIsPyA/0Xy/fH2F4N8SyylRiFjEdoJ
ba4ZMai5b29QfazaJEDTSThlHpSGLwKmTH4XYMYL+dKUZjy8Hx6KmaPMAe6xul1Dbij9KB4ff2LR
8JQ2ibdAC1QEOkmQDtoKsbhEcD5c4ggua1cEkNENWIT0lbdcWrvKLYdggYWPoqLG84rzo7ulBjYu
hLODxhl8n4FKKPH9WkS+2BrEdicuanuqaEGCu45ubVDjqh9el4TeljPpsS35+L0mWg1NpIC7baKT
sOzKgLKJIpJA/5xIzbzWobdgcvXoF0NBwAQcNGR4Is8ZJCoN2U3FauNriaw0Y0zM2jEOAfDjccZ6
Qvxh/hePgm0W4KB0v1JjEWcVFyxk2CON0vTz35UjiqrISvXiXH/2FezLPcOnRglkzWaEJZ4+8pAO
MgLUqX1u3r0M9rGpeEIH/vyw/TM4KZOH5jUboDjdpt5GNRFBtE6QpZhvx3VijyqalE3iMDnLcS8w
sg3hh2sMOmanAjicOzJIcz0WHsAQvldJo3ByqYvoj4F7fNpBdGJOb1IsA1rdy+R82fsZHSkDfnN/
Q21pCw6Bg9w0EEipbqMpkScKB9FQdqt34G66bwuzxUjaBn4+yNXdNC60N0WbVSrtVoMuB68wgc/D
tlgXY8LecyThith1yHqQMjMDNqSwaLqELUkMJK1PjqmEjCRCVncFvrdPOleWXcuwesugUc6G3IC8
Ql5x7LxxqT0FrwH8aAKO18kONqKseE/2EEa8JoWsaScNDVkb/XK4veMHJdT+Me+8Xyjl5nHKS9bT
3c3w8E9RMBmOpXbNVUwdusaO+2R0dKoczsTX/aYFJpWOL3wy6uLB1mtdIiTII0xb4v/Z8wqLVX8J
qGKA5oMaCZ7csa8CZeqS/XqLf122Fi5cGVP5g84/z73lUNhKBgAcRyHGKJdXUg8jdVsPIigtiTOA
6aAvGYVUxusquOpZT7MebLnUZD805CYOIOZxlh6T+GHSjalzdti8vmVVmKuC530GTEXPWM4aMQCe
/ut99Vjh3PdW75vg4yMYzPEiTqoYavXr7UJKWTafmmPBCjL56uD32gMHtnc9fOeB5taINdIwIjDR
a+QgbVJ5f4uYdlhR8APG0gQleBbKD5KN4qb5SEIaEWaGFe1OMv0K+Vk7j/mudFI0fnnFjX/Q2Xrw
W4bw7wN0ao+G3QGbnnc7/jqxfBwa3L4WyswLTd7YAygHcJNHyhv6rY0pLBd5Q7GCFEw8GhITlldB
7lRCjkkUnpE+Ygyyq8cEnzyfNGEsMuQSRwA2MOpHzKU2gl+rXmIeZ6aMmj3MJPxJps9D2iNy8PnT
32omLXslIa1VFhZByDyTXVHwvTLQAPM7acy/igCf4wb6+bZysC5OIQxSojLz99dc2WDgOk2n0nQm
eS4lhqY6BQ3zpagbgNhwgVuWXsdkbzLeHdEkOl1SkE8qkR+c05Vgxk5vrNd3btk8KJo9npmDRbY6
HPTBV39/ovzlPl22G6jPxsOlgmRJQipvujNIy0uvagTXSObugAN4FYEscUsYorFdAtDfPOFZud9i
LpphYtrV/arHt2h/NIoTyYBZoLuSOLsUCcJ2OLe2A48JsdnmEp59rs4HpnNbR1lOp3tZpOh0CHQU
wf1i6v2kcQOU8I9QosMF6o+Rx4sn0LjNq5IyIEoU3Of1sVnTJUucSR5mvoRYhmO14ybJdDsJC0JM
sqL+E0eRxXDDl6JaLxkqRXXtKDfoBXzxnhGIrxVR7qTx/CjnV9dBbbiVhbzKkm2GvRmxlJrDEv99
+tL/XVOXXo6Hcp0E8wM9hMiXibBwnyYhFtOhDJdEqhVnc/HQsD9Gk6AWikum/scFiAkEvXk4elJv
Qz/NZbTSwUH7t1bBmsdPExt4/U93TEKkvodVqP0nNLpOgZWilr0ipkpl5KzIVp84uy2jKZScQI20
hmO1U5GryON1awWrITnn/50BHcZj/1uDRMO+RUsJ+rZ0MnYV6z8kAeUaCVeWuEBDP//GnF898BG5
7aoYES8kzr9Yua8qjlPHpbXBHTSQdorYehR50mYF6ZSgSM3h/1VgCkxkNA6U1l0HJrfpATyt8DiG
S09DUVegxCiv0t9PLxeNc/8pXmsh5l/918pZbqKFST1Y3hMR3soWFOKZRpz+e/axCegp1xx12b+Q
LzRDQEl1flTFD85UFY8XOsYnSekrGDywb2ijsXMsnkYw15Z0Mt6Wm7pqwlZ0AKCmtb2M1brhMupG
bYfD7+1TQl+U+csrnZ/QojY5nOWk5tc295J8ftgcZwtBkujbisbSFwidNCG0vP9ChWq/3MoIiuS+
nzuFBGauboYnqeqicwy7mXIMiwqBN76Zg+Hpj2JTWuybstq09jUbnyGEf8ApXvFiybhEuCNbikJ1
0WDovMYDsSjuwWKc44GVGilz0CxL1GuIvjtqBiiVs0VkWY+GPRlNft65b3e4uckb7SED9UGJW1NR
wt+jqecsY9lC+yemV3QLJexvOI/Tb5XrvmwLL5VIv+HPvmMJ6Bl06K+3wzp1nty/L/qmRU4jsMgc
X/UORICFQewyqdTh4WnQd1m9MKWkjkAF6K9E3pActPwWhbke4b2FjkbXk+zext5efOYhCHWOvJkV
BbU/UF7CTj/aN4rHLfXs9XH/joaS0Y2+yee30awxB2NIB6rWLWN7/kx2UTN1YA17MpvHFzjUDZ2Q
nqmlZSq8pS9KimNugpRsI51gzj/gjfOyfZdyxDVLl8GbKN51QuREa3s6JclxfQ1oX7BVrAj4QjuV
UI/WRCg0Fcvwry2lhgnDldeQIsHnjT0kKX7SjjljuSQdHoVCzBn+z15Yo/3iUiueqzGorslaOJeg
b4DOUMH4K7IZqD+C7EP6NeurgpjCuQ3HbQO8z9ICAxurt3NaJSMxMpQ0UhUkuxHYtEsAFomD4gyH
s2UTnRcQ0GBOQiTZF0PB+WmQKxVIZVbg5ZNE4B34YeIw7lQ1601YodmHMUkiYBLAnGQWHoiyOSOE
oAiWhTLDyxeR5Wck8HNldCJGW8lCsNeNeN1rq5amYqsH+NfPHe0T3vJDYhh6JTR+9eQO9j2gu7rZ
Ooufd3yxyAf5sD3L1S0qiqMyTJkfZMw2tQe9osXFxEPnJtGG43ckRE8G3q21NU9AMhAbi8amyrDO
QCIK9Mf0N+C+SKGbu9CUBlDQkoXvcLjO/K7KO/hzFuh5K+rt9f8kTGNZFhmtRovNND69wxN2RcOB
kszFrVT4cR949d3ycixayCMC5rFn5AHy4QwFq/WmiR5AUykvuLuATVeSvrOHsC0uvY0nldS/UqNP
/Pdnvuv6SyyU00vK8L9KqgJXe9V/4y50kXC3IsAgljxHM9o+MpHSr+4lHWzRnmIaAxFQjY1dH5r1
jQMXsZ9wmmK6wvvyqpmibrhCeUIID6bgzd+Fbx1fXMK9ecU1QEa/jkfP/d5uZg50PXq2vioqBRnh
z4ETdWh7vJPz5vRN3tCfwv0vV6QU6Kuuvbvk0+Vkwo+y5loTafYNOp5vN04lVjTJeUGS99IuoXCU
B+nX3K7RH4CjkRkEz63J5dldLMLvpVUBHvWX2Ld+5pvwmoyULE9CtEGOGSD0zzBmH8bdMpX/2803
ZedGP1oZ+cO7fXuvSX93sHVvwmW9rv4d/9HI2wLBeIGhWn0SiEkpyx6fIRNCDbayDhaAXkItK2ko
LKRkIqFlvziGEt/fH+wjhFEQIgIvE8RG1X/78vdm7oikfxzKDwHVhoQxrHZ335VszjKCyWULroj+
1Vp3a864zS2bMkZWt9pzGB0Rx8ScziTp56RmO1IuhjU9X29nKZa7Ca3q7bcUWwe4lcakbsr/DE+l
8mgLMu8ntbqVQliItJy2rINjRAztBk4eetT0GGP88rgY3nA7WCh4lhYshXcimq6j6LK/WmavdCA1
920Dh56L3MdxIYuyShCNmuBD1MqrntAyhPfHY1u4zPkP/dDbLYxjzcyA/e+crV8DV79lIyqX7PWD
QViRid88T5JXQREpcLVOzDVKT3pbDVawcPWtvyPp0WHWXOS8F9Lpiz/MtBPMWbsX+S/bofewOsF1
xNsLujWhcGYnGATq7LJq2Fghy/xs2HC5McKdN94GO2/Mb0WSlGw64WU+iWPQTyL3nBnJ0hkhNP2k
A/9mvos6QfWxz7QWcogX6Yey5NRwZwO0zk80TaWU+T1DJJsbJP4gMw1t82opDvYfUV6Zz53YeIlK
bZ8szy7VlXgnW2FT9otWRIoJ7ciTsDh7uStrbc3pv/j4Al18EPPq8Ld3tvlL6FYr5++mua5S1KYZ
DLfFoLNp32JFtRGfNhCkXy8zqpwkG+oaCKNHJIo5EyHU42cdN6Y0AzigL/Z3W2bk//kzEiDEWomZ
dojecG/G1m/hSeV+4frDy8wjI63BwcxY7AFmAVowltKRCW+lpRk9bfRtB44Gn4RzhZWGAG75cASP
17MFkUzSbm5OrCgQNqaZbopg+g0wCSakJ+flHNxGaSO0C0/GEona8aA5CcfEwdaQfzr2c1BFyQGD
KMHY0F+iD4m8o0Y9ytfGxamWYS7lyh8Ta9E0WJMUjc71lsnRLveseGm4V1y3WsYvxTVdO4cipYYM
9J9Z2GzGB3mtYJFuWAAJVTpTnNsOjDZuHQP3qmz72HIYAeH8FM3eNTmLYt2abEQjrazdNH382Muk
y/tSgRtuRL5oOEIpPKd0I4v2LEw5D7gG0rmlAOHnpViuSlSrsUoUvKtyoycVWtm378PUhf3yZyq1
vIbjGQ7XT+uZcAk5Nnk/lWn6ihLwyp86UJrINl7uO7oAsYbaX3KxszXk4dUo8lER46H0Cs7S4vdf
MOf8LEO6HFFnkAegMNKYXGx2007Ek5qpPhHS5RlDT6MLFz5ltFrO8lak1EaG4OmtLcnA8yh58FdJ
wod7VMengBrmJvSzdf4ISLweZPTpc0qk1352XIuMpQkkpLROyA1RqYoeND8Omnh43GoqaSJcXo9q
CUDiptIo+67lXnw/KWTvufMVOuPejwlgQgv7YQvsnuxFcx3x7ej8IR/xYm9Ug2z/ZUSIRhOwytBg
lhpk88xEd5eQWttBdX6p0/CgoTXYa7o6i10w1ohRrrXfCjPk1R6Jgw6GXHKVHD811Uj7wDRHUXbe
hKMWWVQ5UASZvACG0hytIw6AZycD+258mIqOIRzf/eTuODxyiynAYncmdUx3PouSL9cwR4rVp6rj
h6/gbJBbse9aMUuhxE/FXIe6hXjO7DsnOTawdwteX9baDGp2KPl7xEMekdIJHVa3x7UhGEhNE3Um
Mg6XzXcqoV+hfbeQSPRTNtYDzQqjciJ5EGKBQQuQChEUVnjACXXZhmnyTxQHHsrhAfC+vHPw/ffw
KRzp3trp9Ni5Gsw8fnhzNwAfFiFFgJmAzZIaRI3AmvChU2KwXkO8GBO1aLsN5Xo/sMyOfMihJN/U
e5urd6P5bXxXG+83pnO9Q9qArnTu1Rks+eCiu+PefFjNjRtPwYtzwKvt/YOBCGpKOuAZR+0lagOZ
P/QTw/jbsd80+lyyUMF6t1yZTHnmY/5XzTn0KD8awj9Oqw9d1zq6GnLTNCs5nmkBGibaNZFkxIa8
ex9G+uxCfww1poIB19JThCJvnI1W+q9CnD03JySayc3wp7t5Oanw62qmccN+p14dNqaphTV18iub
GASEMFQqNqyp+zKqDNpoRKHVWZByZXLEEWppgcciPyt0Wb/P9yRUFXawi3VRH4nxW8zjJy934VRa
bh1FyLMnoX9XVx7DqKUSfrLraVmoQD0D8CTc5CMOAwQ/pMk0luCl0nOK8KWgmkppt3th/u2otjtR
M5q0DpKXp3FaNyFmyV8nqu12k25FyfKuG3hTlNcsqR9QvOg4WsZcd9WGyTC0uIEidQLyMq3aSvga
kGvSi36HZufgsW9Chy01ofleANqt/x6bCWKB0T8fkc9V8AnSKrQypd6UXlDzw3ReEq2ILV8w1zRT
hFGQQ85OqXY2ibRkytn3vukh0Wo8AmFsDrI+L8NoseDS9BW1Iy8Dc1C41Ckv+QdeSY1MOfCEgfrd
qjINEnc59nVPnbH7V6zctrtJKZm2xawyQdxXBrH9YLzqtVWpF6M6pHTR9Acg55FBI7/DRK4/y/TL
smihrI5UFku4Jr0G8CHWDP/oYbSpiC291zz+wUpnlgbFZhBt5r97bSfr14pgC5ts3cn8LCcIKuYk
Pqoi1WNSixZVPmOqWBvylvWj/aVMlzGl+WKQUfpiQpdYD7GOJTYwW4IQI2wONX5t79d0Q7Z1cfek
xuc3w/FnndMI536l0je6O3MvffVQ3NRZp0TefOt3FV+uqaleIC7jvb+TwpqpITaMrrdK2MQa87qZ
1odvdBzyS/mDC4hAMfyYatQcmKumnl+NugvAxMnUAJyeEhcO5nJP5jQeKgVaojMxL/RWmV5t+5sJ
C38UzzFlm47HVs/tghArycm6EVNRGlgt046Ygj1TC5KKqMTOuQpls4g+7AXxMF/BT1fXzzTvwOM1
jXATQVtSLCYBgmaAKt0H0S5HXNXB1d6FSOMrL0pDOqtnY0+QmoJZbRg8lb12EFl7T2eOppmgJMK2
2LNr2L8uae80mRIHcDm8j/EjvBBpPLizwXuf4Xy7CIwZvFn88Qn5US+gw/E/LpEu+g2MMPJsEJv4
5p63iFT8yeqI3ahY9/gccGTXqepqqoGzNfNi/e8IWXJRuKMfujrqjhWZfcBdfTBhxpLu5tW8kZZf
+2yazaqu9Zlq6m78OQPgpUrqtndu2zYxaKXTY+7q1UqipChOlMDwiwgVSB9ZfPEyeOeMwuXk2tr6
LacoptktfOPS9Ob4jzoIua2NEsLa7xHE353QY7IW4qITeFqUEStW9sifKjAUVsguKYew2GgJ96Gw
qMOxJn5zxCySe5wUlpCU3ibl+CR5XpMBfRSrCdM1E/DAuAk7pV/90F1yziOJt3y+t/DWGRdq05dT
FHZ9G7GkxsPpBTuNfubsKFb6lozjMn1LfTewzLUVcdLgVRM1uum1/0J50r7/2M2zNebv+Hw4Mzbu
mIPSyrky+fd7lHP6kBajVlPfPRGBN/gP5S+1jjrC5KQvLExnTBB2l4aBd5oilJxbouKJWcGy6HzN
lh+ZhGir3BkIUGli/xLw/1AEuqrLSEpwnk2aOMHu3dApxvyzyK1a7DW/mwKif0b99T0mTSti7J9I
7YEa0iafkBhUAv54y/RC9x7a7tCBmHkl2enhCoWCNieUpr8keUpt/NNJWtYj6vjJNm51ioZhMFr7
QpjRFKIAHce04N8nhEnZcaG2Rf/SlZCoMwAtMuuKIIGV88BAtvNIYLuVjCi6vb1eJlvIyXyQUTPv
aUppTfvCDCB6MC6xv5t2G+emXcCL1O8dUp1MFTyJb/ccE58U1EZcYCiflqmmOpuTKLz3U/IbQoJ+
vXWr7fsMekXY4hr6t7bL8EPDOnFvd2J2tk1gZ3myFpbn3ZH1bbS+Kiiui7tisHBdzGKzdVSz5VcE
lLFB6iE6SVwsqsIVv6ngfYk27Q/Pwx+VW3awSrfxMi4HdJ54Tf9pKMn+9cxfpttAinZM/zlS6n5y
m0JRuaOI1eX/dLBh6sUCJ2hff/0J8WRDrbJ7UCsWJNL9ec1skbYhqk49UALj5LfE1W1LSNNbAnZN
YOuNqxKwISp+6ewiznZk3hKgYEV6fY60NHZc4dGBpB10ejZUiE20LdQdwJZtiky71IUfXQ9izogO
TOFwu08DCfs+sarBpIkJLIC9iZJ2hlpHawtBen2Hvj8IXBpRnGlf4XBISw2XPM4VTgNKZ+wNVTkm
XsJdg+/FRBYNYwSFBmwc2xheC2NzePmcUpFKI1T1tBPZv2WNclrSSPxqRfibJVtCvURHFKlgkUBv
Cu7jKiVptQnC7NngncGMQWXRCqtl1YxRB8aszOQGX/NtBC1AC4Lc5TnGlEQo54kgSzOw+I5xU9jh
I4a4qxTn9F6NMd4JXDvvw9XNF2lnYAZGrZKicyT1YCwh8Hjv/CBMN6DwldQBTBs4S0YrgWcgPb/2
5BDgMNanJxKCEX+HCwqypjlQTXMJ0L3lxUUa51cy0fHBmqtW9R7oh1TNDJkhnmNWS1e0sAPvsF+n
KmhDs5ju+W9BKwMdSvk4F4/GhWpM69X1Ko27it/cZZIdg4AXL2ZzsuJmZ2CeApybxUMFs/apJZI2
k1fZCMsq70NVNYf+7tZep3fqavp5JMLSmBAhWYuQ+cEh/byKZ4f7kD8Edt3dU3IraRjU4eWzO2D9
IEAaFm42CzM+py0n9rVrw4LD0iUpjJVKyIe08BveFdh+3/mhd6OfYknGzqtsJibJVYTTyXzJR796
QD3/SUHtOS2fLpg4ZFEc085ZgGAp3BOUBBNLAzkrENUGojUdWZe7bSNvHwsQwmA5XYjA3UjJR0TB
RYzO4EodWwxLi08PgmFzu9GH0ioy4E3Bl1pZhVC3JH64xXQiYD1mL4rffIA4dWfTuSD9zdCmzLfQ
sGB6xyHKTaAKgGvuddufGVO8m66G6ra1r46vR7ETkAUsDCue7b2E95B61r2dQISWHAUNN7+mEthY
gR+pHv1JO5wLHlTy6Y23s2aX7MoWTpe0qDwW6XmA3vIFOGBL1bx3ZVDPPn215SiDWdWDgyz+n3+G
EXLMhKRTp/543Q5MBbzX0jAnE2+4vUM2Qb9GlR65aCe0OumobI5qHy78bsiM05EqcVeIQ1qqPdeN
REPg7JsWWGSkQ3E7TT97E/gjmYJjeHmey2lEbcytVvtpJqu3df9jPHHSTgwRGG0YsgVejmKkyHWY
JOUXCkAQfPXIj/Dz1DmwpExxEyZCs1Xv2OBcuqRHvc9V6scsbfTuIKaEvAECw6vuctDG5up/5Y+p
4AYsgpJnhQgKBicmUh/5ev89jvIPr4VNjJhqjBSyhc7gSiKBWAy2tmFYPBIf2EqS+c23IDFE1/O/
l8gaMBq3gWiQJ4hsmW4fpjIhk2I4my6xdz4fCFYBFyerYAx2jWD6399lkcThvRUtXJ+MQvlEEV4p
rOGtTjaWQaMhFD0BSuEdgX25MwKY80os8NWbFOo78AIDp9mXrrR3MxjSCJRkFoVjlmVfQdv4QY+H
dr9womouR7zbTS762GlxcLEbUoAwAqz0fb8PP87cYo3m8Tna1BK8wHmEY6E/tWDJ4OaOOlotsVmd
kIObxq5NNPTQO1ioI+bFIkpz38FvSpdCKDWAMkm9+EcqjCpPPFt7HMMhVmjdQ1GT7D3bwDKxyZCj
0DehuurWoPpDgC2sRuuNddnJYlVqeUb3SAcniXt5FihTumPJfjV8ytdP0xZepfLbm08SvFaxDLN+
fICVldd2Z5dDu20nUAYyAHbgWIZfCTtq4UEQceaGu5L9lfeHWpzv+ahfuJZN/z36lSeEt6KtPDKz
elKCn3OjMFm7BPh9J7ugTMeiSABWfPJyAPg+XaTIfMNyD/i0PlNGGXAlT7F9GD0vqpZQSCS2SEmC
HRIbLei2eaMZgIZEV+1i1fZSMdJ4m3hv0ufKjuqb3WkD4Y0wjLu5yDlRUDm/GyifIu2A9ymeZPzl
IISZkn0jKo0hssK4kPUgeCXKTiNCcinMwo5FmHMdKvYocfMVvrq/FRtLt6gMxNC8L3ab1/GIrvFu
VQuST3TQ68Fr+WTCAP1NNVmf6QVmme1ddkHjs8HVaUh+DnJhuGlXkavOYBSB6cIvEaaZEY6zn5oo
8epCKjSiWceOhmOmCSDWq1+ErKs8qzM/26WHT2yEcBUvsnLh7Ciw54t9tcxOCcaaH/uuxIPKlXeK
uaw8lqmfGiyLjrVF+pJc7/i8zL89RZ5A9dZLrOB3VCAU4UeQ1DBES1w29GZnUvSTgs3nc9oiU3lX
MkxTY9AuYayWcFTmKI7eHicAaKxRkqu1Cnl8ER7jKSYy0ti0U0fkPtRONUYIoKVyHxwOro7zybri
14w58n681THTTFPm0FYgWNWSxD5hz5PLN145FNsQ1LS41gF3BNfktFMCPXX9JCXbMOwpxnsBMVDb
8/LVmHgvK9KGwE9gmdL87evyONvcMiVjVJCWj30ItfmFLdyTX7LrYuy0wboo1nDk20uaFD7twqR0
xHlkMgPWo2DZfK0qLirkL+VREDRO/z1VJos1oole6MKBArwtOzDYx2VIYk5PqP+/mZZoRTpTT2Cm
ZgJ+H+fxYCLXr1+MeN8A2gRpfEJSf5GsoWkkpPOE1ESsVninbAwA0U1xlKoS/th1nXv6J4WEjO85
I87teuxssXMTXBjGQXk9XprHcN0sRNL/sLfEMtG5H4hKgJjCR/eePdQxAzNz2D3fR5uOJ3Th/Mi0
z613D2RNYA2FI5lC/5sWf/er9Hcc/C/qd9OhulAunssGC/CuoXA3zfoe/P3/T047sGE9TdDG67mV
TsQTOHsvb+J123GEFKSEKssorgprvhNb4cwjdP2icUV8LuLyKn83Vr059u7KDWNDKnxl54lA4Nbv
2ry+4RwzvG85hD9YdyEOxQY33jD4g3vRSnvgTSS16Kx0lH22qEJQmOao276y4IJuHo2+hVQPvy/c
ZNlkhq1JWgkRTbkozCFcUSEDyMV7Af158AZlYz9aZv+PBF5vdFtgnANMTk4XyjqyODmKwUhNspFm
qFASLzyNzTwsxV2HO7oFbPFSW4WMXh1vl9LF1SCTscZc72xlA4/oh8ckVsBnRBPLqKOeGBPRkSeh
U6SxPo3Y4BZ0p1uxEfapyK0Hbrt5UvGYL94lT0nkbgQ99rfue0ItNrZl/fvbxNS9/G6mo2GiWGRO
Hrfqupx/wCUuRpGTx1tiSXBqImK5CZz6AzP+Kmn5r8ngqyiLBRkWb9pGPYAo82FndX1b2Ql4gfqx
LRBqSDXkNRU/mbyjrAzYpSdz+2hzVexi35tacnL6B5rQmaDkrqZxBtuy7G6r5avWm0LCuMgfraIu
9y/AU+Fb/dTaOxViXHPpY5WB+tvWXlVnR2Fbu/zbYxTAElSsvHSHY7oEdWZeG5MLD9TFsc/A8nkK
5fVs5VwzyX2yNAA4ZvRknx2qG+o5SW2yzkj0uIlSvabuvXcMFT0OC2hNjuLvKuqxahe6i8evJMqg
BppIy0hhMhzayZ45Uv8trpu7ELko1OYAwCbp2OW4qrnXEiGT0aE1IGEo5T4r7w+xvR6uWq/NvDUK
2YpM0jwmTm5UMzuGUAqXvqh2xAkep5eiYmrN3hbGLbYRtUWGEZxJxsXYt5kU7XfwfWoXVuTERdjW
uQioItvu9BIB57mo7zFFjeFJzv5solb+XJuqR4b7ccizCOKflvs1W3UGMfFqIRBIo6mlUnxqJzTm
qaoVUk5y+sUeHnGK6C80bLr45VJK81ThtAW0cypBrZS9tTLUBJzmE+RzUlvd71BjwocQys6NRPph
JCf3/gMEr1vxdlHb+xNDeb5lOeamsdOf2MaVOEZ3hrQFmIu277pz5scXVKQBpzoW2NaFocc06Vro
DMwDkZlogP12FM69jXIkascg0Fb84zTfcxTJ11Ze4hJBDe0KSPNDmtymgFsN6O5SyjhB4zSVqO8h
NrhbBCToopW7SyxAtkaD+5fNDIqNlxrBMUmoQ8gua50GTjQXc2x4et5EgI/270nJryVUnXcyo0u6
kafu1EzA+h3si6fMCMYx9WS3G+75G4NlMB3Y8Mmfx60tYRGsXTuHQA84BGxUHgmEH6rsBXcpt6g7
WuQ3qs8KH/XBlQGGpQBh/yi9zPg9qvk5dKjtItG2uwSJQIsIO6UtvhkhKiBW5znyNwMZ84HKenU0
fe3JHayhVrG+d6PwxAFUwCvqJU7WXJC5+apC7Z1WBRgjwEOVjc5eSFcI+qbXaVxPfPLBdhoqqsxa
97bfUYrW76D57gQvWNCx1chLiUxp81K/iZSKe3/vxSJmNxAgB2EyNGtCTvZlW8FX5NXjvwb2+SDs
jh0KNIi0qNGXG0ca6B2avLm8qOkJ7CDSx7F5V4pwnkF7tlzbnNGfdEni7L68ANBrswWcVuXp2OsB
cz5v7BH0420O9S4GuNP0u9ksS2tv3r5k1wnSKfpnmEoygrzIYopZQv6EKSRCtLrLBdGWK1wJuwHT
k2q1GIM4tHHNFNLUN0mn7qMPJbseNvtumDMMNoRXBfwpBg+8iF7/VBTubUgzDH2RWNUKhgDHL6p4
o3gr/VFB4FDEL8YLgdEwLX2s0fTf+96voKUm5GiFVYiLkK+ShXTdgSHZmKNrK732ZqjdGchEQ+xp
mYbMeqVcJT4dRGWObQOG/2q+mq4YRdQf17Gp7jPBeyawVxpMeeEQu0CvxffnNmL+UvzlKPR814V7
AMSyGjpnkAFB4iCQu6vG5SmNkfivV3JxlrykLSiyABIiuNZNCpLmQrglWDeXtedpYkX/zjVKcW+H
fcV72ECNMyyjHUBCDY1Iu82Ju6aoWHyQEKF/Db66h8VsiX+uMTO7aZD2nm2mcMficv9OLSqcdmNE
DQGsHO9IlvivcW4C6CKWglkMctUzXLzjh7lAD3k8M9ByNo8Y9laYiOTJbX15oStaiK6nLH+hxDR0
OWlHKFRJ0MtOtlcwpRTr1WV+D7kdLPHtRXuE0/XtGYymo2S/oxY1BDiX2wmAaSfkysAx7Pd/HFJl
yNj0VWUSMH2hnYPfQ0TQ2zGpvuIqaPzVKVPCtXF6u+kBZftAwwl4zRvGeWrDcUtExbQSVjvmK5Np
CKcJpdsshRACVomNXDPqqSugvU6MBPIE/jSQByE0Yz3QXjKz1V2zDb3IMtfLqZsPOdPi1is83ro4
9IzDHRdWdIUCx8d4eBA8drlZCrqNB/oZznZw946BMQvunfii/F0XJzmqI6fWw4KavO94RZKNclfb
q0qeoS/m1KswrsCQvMl2BQvDfc0hk/x591pFYY1HdOiKV8fJ3PpY1fYnBProltjjMbD6tkSBkpzw
w/Bhd5lOmmyN8ZRcvBbnc+Gq08offgB9UIwykqEl7C8Ygoam8NiqUd+3B5U/eoyknDaLhycCIXnl
LOh/nI2GnglcDPfFNNE7P3wPnUZcTczDrXcJWc26h2sOd6eEFO/49lsNhBsJ6GSkfEWBK8tXJlnK
pjCQQhoTId13IS8eOI0TXBMeSEWTfIRrBu01+EiDA0VKMNWhAqLjHUw+MwokMqz8N/phqYHPZ1+t
DCb9YqC7VaFTgxcleiOFe7U32AaZDCnR3YR7IW1Br2R8PZGh/M51/0NWTHDmk00/t4g4tlKJF4nv
iX/2erfOb0XkXjm/ypdmkZuaIs4n8HZSbWh47w2Xw9jxd59jwumO1uCbrdPclijIgTRMzJNprgEG
f87YWag2eAS0AUtDQHV35bXYNFDi38qL4vKxm4ijYkzyrWSqz87hTKIBDX+YMTCxCGQKBo24Easb
A6K/O1BxOxunG7qtSj/S4Ix4mOKPfnb/k+PVg7VU7he/3Kup0kcsOA6/X9IdHTIp6tqiar96naag
SFYjlxU7TI8/VYxaBLBe+dcqTbe+aG+6rY2E6hTadnRxyZFKeehQ+Q6gg1Zpcsvf7He5EO2fZn40
fsF8umHIYIK1nUjA6w+4g/UO/6rUE2xJ/VsywL3y0nhCJ9cqn3oJcmK2USIoqhVIhYNHbGiZXjMu
f47MEqNxbdWu53j3rkJ8EUgYZL5xJ27R+9lt/7EOS+ngRejvIO0mPYLcpJXO7HTodSU9stFg9liI
0Nih6C+/aB0wz7LNDMsA3JPD/bPH+Q5fUbTYTiXaACpvYl9FRYGD4exK0Sg1BZJWjWvq8mHqma5Y
14iPqp4GO5Y2tCxFmoMNXCacEVxNQE52wVrVCj28y0AS1EnO32UqW3O3daz/xbSuZ4J6c1SkU3O9
O2BflW+sAYhVDB4/3aIx4qLsy2fLXX+MRVlQ9auhDndUeU43Z7/beNjOs6vIL/X0WZDdJyD2wKJf
c2UYTGb19PQVKmc0HdQ0d1gLHZWzGFmTQ/L3wU+cJrL4hCYQQUa4zl5Bxw11AcHsP42q7CgYTcXX
BNQwAfLoWNkawqSsr3ZhiQ8enva+FmD2v/UX+ihI36/MS7hfbTter/Pq0213Lz/sIItQyl5wkewi
DS04jQzY541eVaRHLcmwvSwrtNsJ1DRvICHzJ6ZJqc+ZA/VD6HzKmhugsb8d7YFtfSVLBUZeOTxi
wArNGF1dqG2Tief6yB66SybfcaFX/s7lTOAuZGJ8XGlDoRpToldoIaZnaiqOtfbFbNN4FB9/lh/s
qgADTmLxFm9ZYxCmi/xhF4qbQ7XWvFdPqJbRZF9JRXMjqcLFHhuIkXm1A/itT88pU0nbPD8GWDkA
kUUlSs/TJlWWceyKVZYNPZSD7838I7v9i/SwRQDI6gqemUz0/vyIpmj2HaNcKxVBLPOEsh4JQE3e
hYXAXo81GkVtg354vp+34zoHmSIsrHjk8x8eFH2fT2mxSjQbXd1OBfCNn8Xp5sqFzhQiTEwvLrCF
Kh/euSho1pB78gvQ6VSRE+n+uIlRmCEjA8e+/yxJ/pA29pdwnrqykUtvGSeVsi3h34hQXACxpg2E
33kFvY++Rj2j0lB0IgVUyzSA8y00JvNO25JUJu0uyacXfO70z8RGr5tkGVxTXR7fwufRuIbxhCLb
/seDQy+drFpeYIDHgAzL2SlMsLf0Tr/7LnEVLHYx1oBbQmGt3pH6qqwGbLmryGjy2L4kXcXt3444
50GgEQkWnarEQa2NhbTFbIi/SCVGWnJ0XRY4MvVmJ/dwihrafbXQ9bJoZECR/EOeQhDvP63Qnr3o
FnmrxAGpm75/VPUUSixLSBaTIQbXRf5EMtvoSrFbePfDhLvPminbxOW7RiYTu+IMm8ODPewZtTJO
hh90Z81TTEVMlipSoVpniJ1vISkjF0KF6nV0vkR9Dkqy5zwz7HWkqAbrbqtWkhJgqxgKXFwHk3Am
D4jZCeuVrldHfI262iYxSlldU67VB7FG7WAxknceugkUD4ZZWZ9SR48eNwHg/2NwT1FeDj2J89ay
guRY0PzEYHRt/PjxYYIuQI5B7zbc7/bTCfoX6VmT1t2PDj8pxSvwWg8wOp+gHX0vWOC8fbimi5KL
LI14LGsuo3szV0zWYPFr3BPpCS9rpxDDKpOscUdSLUlx9rPXrbNqbmxXbNPySq2Kdwa5PmXPK1WP
ZVowQ8318pEoBJcTSQjlLNxEcqGa1lqD2vSB0JIZzv/VwVC22lx6Y7EdkPzY+7iTjX26de3sXIY1
C+dKGn+b6x9TWxZfU+BQOSzWMV4MjAz6+Uz4w+9Q6/fABTM4d9/PUjwJ9FLlQwPq0GNFh1KeRXAx
O5F+KWPjoDWVWBhiKSI9sMBsRV2galqs3uJOKmXOMuHMKCoN0JmQDRv7w6evRr6coZvz9tcDdup8
9xEvMS7zxQENpgT60cZUnL3BptwfP77nuE8fi+I+jdglaGhTGLDQ6KXRdDPdts94aYnCO2ox5lLy
eOTjNj7p6bUSWNuWt7DAlJ2frB8mIW2mIl5T39NvrP4cFwpluj3MtlLjlxPEcy0zODvB9fGSWGXE
w8ryEtRswYwaWkfNGNvoRPG8SlWacNrE9C62ZFB/0kimxad1lFWh48DX5DrRmEEfs+/mWsnQFeqE
27QdajgRnwVJ/r4JCjLqY1JtS8fKp0WctdK3H4Wd0JvGOJRNVJ4yUqCQvR4DCdz9MUY/6sp4A16E
dMGIP1S3xzQ0gVAMeraUL8Ria6+ybN21v4Ew35hgtaqytzE1zPhUUb6cRdd5YxOldxOlUYddEOWM
txR+4kgUhY5oVed4a1R6v0EYTpbbasUzRkqTicVfGev01nB/1HMYlYwrfPa6il7SdL8OcfnVTq5Y
Byz2jM/j/RWa244U2u1ZA/MLQwA36jCS+2jdrdc4DBmxSupWSolbTacsROy7zhaGAEiSHiNwFqkk
NbG/31OBZLz6unRgxRtamwRBsnxCd+fdhDkc02MmLtOtW+LKD3eral00ZTLrhgzrywpwYiR1cmOz
x3W1NgDOauUeDglMQy5ihkh7w2LnW5QApESUv9DqLeC7LIuTgQf6h3UalF9RpyTtEWCKSGNehidC
xoMEmJToqBnZsuT867mgDK0a9DjLchLF5NBjS2Qs+j0j0JjX61bCbUqbfbewygTEw1U/TpnImG4D
JbJcfTZ1c/rrEiIO70pZEjpyGaB1nu3EevKyztvhno4+xeQdYb6yFpaClACvXVRx+4Ad6qaBzZAa
a0jijmWo8ZUiMKe3FTkAkYvCqmtOnqXjppBV18rF4r8N1jXT/u8iGF9AnTumEFXXQcCGbLqZsNLA
Bt/PRXmXL1JlpDDu+rT9FtNNZ7w4gHZ8FRPV548qiwtbt/JKuYL+mfAj/scmW8BVqiZllBnppXuj
BnWYWPVGzzpFYqV3cETls8cDh980YdTTEd19M9PbWzOkqJ2oMZK8Pd3L7U5WyVWw7wirJ2tFejvb
TKMRZwPFrbT/UILgMsJ02HE6Xi3KvGrbOVEZzm5RdoeQmztgpkE5PqzPPJdbQydDPPzUFZ7esF8H
aHLEmQ76nYnC0415pgPjtcPnr3wt9ENQW3AAlDOZHJxkMU4ZOIsomLUh1oeu9nUqmvjPaiJKuOwZ
W5vWR+dStAzm1MB3/BN2zYWS5YNW9nwdFGHlqpC1Ojdu8X/8fS0W5iguebdEOC4s821OYWXawsLs
DwFnp/tQQN4llD1rAijZfIAUBU/kBxtPfhzVBSf2idI4vMw3Vsiw0dAj0ugF4GlL4riN4KbByJeE
WTOmZDjxVYS1ozI9troJehFPhzJEx0QEruHNbx16xUdoLPpScAqzcCzZYw77+xYOGoCgezMT+uQW
1tE3JFi5TCj/wOZz5ZFFImFU6yusivTC1oeHAYVy/ulXBNwdzVDD10B+UF746FfxMAVpPlRz1J7S
uyLTjSp1c2wADSKtdkhGbqBmUi4odTqy7bIc7pt0dfERP5GaBbkFGrLJUs20RlQ6pPrQdOR2xzP4
0ESBiUP4SgP8CASxNQmLQ9ffzusnZjJlCWUjkbajHVTSND0BR42AjLQBkzvv6NNWKd+VHed41wbc
yr0wNQumh32Lh1/rgyntQPxcXjewtiLM01GLBFVljCxNJkNgreRX4xO/j6Ep2TjZ6a6vyjziJCr0
x48HgnXyzC9+6hfFkRkz93PuanuY7HLhd3aetwpV8q4aD7/bDAb29o2qULExZh6kf30KxSpJ/jIE
zXs9rSq45FZpwJH3PYVd/wubybM/MArHSeJA3riLfSTX5aWSxAogYljtfq1475huF8AFsaTdS8VL
ueSU0PYoOwqFKLxGmkj3kvzVmjkH/r7CPEAOHC9byBL7zjO58yoEJnlVwaY+iabAG1nRGFcf/bi7
J7tiyaJqKDOOCrwhkdu1+HSE7E5rPz9qTahsflfsOzae13uoy6qBt9RGGJxFyXK/TmZ+jjhjsBEx
FE45KLs8wC6JSE2RzlWQ4yII35V7kEJD5xiw9RgzvDgp63k0nfm/AfPekLIm2L5eX9vjem0u+A1R
qyiiLgzkBfiZNmrcEypLtG8TOl+16tiSiEbfZT59Uf3zvMZxIkNy4f7mKymO9UocV1W3tzy6oL5b
ZP7Bb5iNxzwYKvfjO5X0Oqk23UANNVenPBmSOQU8L1XoI8OhCtpUboOriVOxxy1qfuhjAvpf5NQ6
C/8Pd3C1s1iSj3uYMIqM6hY/7pwIvjrj4MUIhX8fqv4vNBA5PHD72qmPJz0KOTjF+nLpm9tOSECV
NRZ0MMFZAPCmfreBtlK0tzGLci1dCnl499aFbvh1iuAM3lLmkc6h+ZwLt76C1jQnGWLNgRkeWk6y
3kL94ItRFKzhWobsZUYp1NL4tlYfU3F9LVETsK7VmE4kbroGTXCCOinqwkRSTiDqMrzvO+7PKPV7
UAL6juyM50HUxTQyVXcyVlC3oCjjM8fYdnrn/W2QcDHIsR7W02GDHSsHdaPswrCK88COYOaIyUvW
4nrjtBUa13E63p/Uy+ghqS3dNiyOjE/Gyj6Vfn4ixQFfBCuZ2mWFEUL2yo+fXWnW2KREeQuPaiYE
/+EtgX2YjuFw8UoDtdB9MrVX4F6anUSCdDZzCJRG2mzBW1vCN6JUbTFn3SO9oYc2+PbVQp1Oa1c5
FSxCFTitIUuBegfxE06zrh9NZceklPqlRfDqviDCemyCCrlGvLSO3un//5knTg4pkfi+/8oAnRep
c49UUqmujP2JliStnjCSQziLuiMeVdm1+WUeAZG3+dpaaM3gRWg5gVCINQNQSVCdWzwXbpzUSGNw
UsE10h1TOb7o9QGFyCERIjxQBz89wqxrMExNI0TGYyZ358KgBoDKoYxP9MRVhajIVbIQmxNd74xW
WnFXeY2tDPoGP2lgjGMKAVwf9wIf/kYvi5xHuyDg6+Hh82W0vrCJcdBBje0koC2P+V45PcYXSuoI
MInXZCvRp+9frxYTav+x79lvXsQo9gcKnOUNZUCoDrnEevIa075wwmcEdGt+VJ8kHy2tlCcKbc0Y
BoOgptUlq/x0vfBASSiHa7PZ9Bzu/HExNjquIUQM+5XNAneqtxwF3MXKfkZnbRub4omPdAojwhW+
iDtrvivNDzWZPWaCWW2hsBx4VrOZT0DeRsUw7EmTfKbUXKFHUN79WOTB2TYtAXH53vp2V347mKrU
5djrBovObtfp+IWaJFBuoJDC7S4XA7xrG1PqA0Xcn0J0BJUSJn6P3P8k1uKDoun84HHyM+X7J1EJ
1iLDGsR1ToBf+m1QBALDP7WJwz/DK9lnKp0aba5qUwjxbKboUNv0Z3z1DXttWr0DCZveWi9VLznv
1b15QFxA5k7Wk+hzmg0RaIp97KDDNLNW1EXEFsoCPDjiIJcfZW7lWJPXiMcChqkNGDvBCjaK1q1c
jfz5d6xcc1m1UvEIKa2setRMGfN0Bsx2AabZlkkvuKp/7hDL2CG3vUCBaZZ2EZP9mlm+F6pQxZhI
T04nqI0pZQTvgNmbRLdoQ7K2x8hLVyVuGriVDEPzLJLYKYq5dbi0rlJ8vsRcp6epFEmi/O0mflMC
NOiSrJnCVb57CA8qgL2Cr1uGSw8eAX6vMFhU6tBd0k1bz3Uj73/yefu5bhjE4RyYRVGqNGoQCZra
r0fkiPPAtkExo3kCSHQ8qphhbgdOBpr/XM8ObYJep+3R+J7m4XdGo3FG835sI3A8TWbSCjfUErbX
34nMV3B5pdyLwoMnjjP/dAwIfb5oFWAkVMjBTGW0vO2y7VfTyAwfou4a3vMQjZsWHYgASghqEfcX
8Tu4ZpaRMoa/ITY0sfBMSGJ5FRF9+pFSjxcPmTYiAnh3SiovWsNW7DqmIO8r5XOBdLlHM0TMPmHa
+WBnJF3TYG29LNOAKYgJsvIvojgc3nhl8xey6d/l2raSxADE84X9XOng1YIUa/CC/9rVmEG1CdvE
8mCFj+WToy1zGYo4A3FoodTVfmWKpt/ZxHlnCnNQ4SCsMY5dFwYbjpOKB1JHEAH6VdNeAZIfhJjN
LYhyHmuyLgOVEUpng2cLYSWx6P9wFbFZTrx2V1y508p11U6E0FkQWZuVYSpD7tCVKoyuq+j4VOWB
qGiEOQ+0uP7kBMmI/45Sn6tX8kfKU4P+gt3eGNXggAdn7Q7nEEo633HmzRAKkoIc4tbV2N0vgmHj
jEXi/bt5EQWXFQ5UHZVyzMiggvfJnuW4GqGCLkEtlOPUqNETD93FVGnvpI2Rd4ozNsjwmQAP9EPS
eSS4NfmzgurzjBrR6AxX03oefeSudKfyu9ZRdi6qdSV61V2nnQMRJFzZpDK6QNnm85HqOcZEn0aj
Y1KAyICqZB1dEDBgKuZqSYBuYRpOQHtfe2S1w5E3x8YheWd65yUbBaesXnMlX8Phkm8xScnU/3Xs
bj3fWAc+AB5ddSNlxlwxvnmPxh+ZNxMLLesY1478JHXIrWMmvxp6vmUCaPt4WSXtvvFh2QIZ4oXT
FVAsylFoEHIewphLuKI6j0iKSOHqzI8uOQljh0SH+wxRhUAkc2Fy7FTvugogBPb5HfYUgBR5trr4
FZII2x13KBT1gtqJwdb9xeZtGRG3WVbfMe93CBc/mVRwNf0aeRJxO4aXbEghY3C4ZfspUyAfrBRE
iAYAuty/zGZcD9QEkXAnt2Zg9D7ogkVR2Fkn3U9BT1xE1TrwqbKDWuD1MOVL4ZKEqRlkbDyNniY1
sXf8D2MI7AIfFyTcTSI0HMFOyalsMwfCiCWvL7V/a0593tCx/WEy6CJt9NZyUh67dA82V/H+FkjM
QTP3KmI9unEtDjoa8HLFAs7+g5fzKvtncUxrExbUBZUXnmiG5/kR4xWaSZ0V2XVsBBUQ6wVkEGg7
bDps/XNwb1GhYnmE49cERzjMdEyf8Rp2ki+zMg/bpqJLenXH1scd+O/MBqfah6u8AjfDxaSKPLdW
5WF5EgcKFvfDo535UeYbxdx6dLRdWqD75mgTMqYj/3sSgg3VbQnodcqSyR+gP3277DhZKB2L+UIl
ClzjYG4jI6qqt7i+64MYyMYDbCAJ4N57Q4nM7f7LtVPwRKjbm4JN4J+qg8WryiB7aY6O1N4QzWJ1
awjs76LtIXcjAdWx+VEVWDrierw/MBWuDBQAJV/ERWOLjLqic/b3Tfm+C8jtU0W2lvbtO1cZQRI9
DmszDobEShU5AD6s41xLEy8nx/e4WksZ5qSeMIOFOTsM9opNe5I/jvoWSfbpILH65ZVPzjmIZlZs
0K5sLa6ZqNDhjY+s67L6CovOfVys4XQyxLlmNz1D3MqoNrMQHB/Qvl2vojE/wEeOCgWy4gb5zWfJ
F4isRwHUb2EtTDrbLzBibPcO412w6+uHSgrP1DAM6WNjn9y8zoLNLiSUfW55bqZia3CNwr0NMohL
56KkYNDDqhzy5wSYIR1kr63DuGssniIZvvN4oN4Eq+OEKIB6kDX/lvB4qXvKgQnFaaAglkr2rDB4
XegGCJwM9an/kP1/LM3SXbumBsslXww+ycYmpzkvwEGvZs/p6av4XI413+bRRyVrYpHELMnLF23J
XEnyc0IC6Vo6tj9NaQkMtOX4pELFzaFmjm+WQCyD0EPi+ghf1wRNMMyC/FwLVf6FRiS5ZXpb2LlE
Z0spy+o5FU1/M39vUZtB4pRKldNJI4qEu1WlqmV/WZNuf9bU3/W5SOb3pvOetYYna9NCJt2e+NEG
zQ09L9HctTnuX2DOmWwYT5rEEPTXZqMm8ZPTJ53camowB88WhVMMCa5u1WB9MkcitjfZ8nKztdfj
2YVDrXoK8BwB90ikL+SmkwoskTHWNpJOADkojTeoKFUDjgUqIoIOXVWWE+dAlbZ9t7QMNwPrvBvS
pXZ74OEct2JFzXE//312uHe05zfnqJzOqXfcCfrq9l6NazfoS5O1DrnvpxvZiSVeOBQt5IXENg5x
mOiQV0Sn/szvkPxSa4CsefpCDauTfYyopobBQOebTgeLb84vnSUIM2cCOf7WHjXG1KLBkuxu6Oa4
JZVPM5dujHhW13PjlwEI+5vpvUatsDG9LZEZn1PQQs1AdrYSB62NinENxahsPrcAsTNUoh0B9/j+
NomvNx1QXxihl1sgCRec/Bqf+QWxHxOhIeGvBBplS7QhN1Vlcl6WcS6L25II6DRO5NfMYvMEJz4B
F+x9CrgEsuoy0xs+I7hMxlChPzB/8z/Ep5C6K/PbfpV/n8t9TTnrTSoOErueTkjS1rxGmGQCqWdM
PFVaEh0NLmRWQqMLBWxk55YcoX8Gq7dUYLAmQDjj7awGJ9amBPPEU+EU4DXSH5+FX3zjsR1MuvUz
Yqs+rNJhfhLddn6qwVwGNGaZuQzUHprncfrCH9NGSxGGDyN5ZyO4bQmVzCnPqmee760wr1N+d1Xx
Gw5S6W6bndpmLc0skXljBsZyos/lEVbk+K1tn9HjBF9s0Pfa13EpVmew4tjZ88qYKOmBx2DtOwvy
LEK+w+1r2bSgzb9DwDtQ19USr4LR0D8r3EVyDfY+JC2j+zerU+9gkDI5tMDf7i/vb1+xXDplkQk2
OMFrK7WNP2ha1JvVQ1GX8zDkiNI2Fbv0ACj8Vsdlwo5nVGNypSXxL1/0GkKKMMiLbo/inBE4EzND
9B/K9E7C6BpRzrEnVKd6rzCrUiCK4+ZVw6++arhEshK2GzC+lCEahzhik/9RWXi3N79jw3XKmR/D
beldUUZ/93ZzrsLVtvM3iHLKy6sYkIKfAuw8nBJJYFywxhk2s2hSwwkj18bMrK10K5G3GOhoy0RF
EdaPnuyqTqg5DRQAigJRT4uGDQp7oH80Jcv9bZQci7+fC5rAYP3/8IStBCrQgPw/NbvshZwZPcXG
poSqLc1C55INEVpmtzprQhGcBUoeF+KKgQTxhdI4Uhf15IzMtDRd+3L+Y62bVetFo+8pv4KycWwl
/8ZM/Izv6At0l+YCdwZr77/cJbQHChUQgTCsY2+y5L8LH8AH0BKrhOGYcMTBUI+6vYWzPMDF+Hbz
v29uMh/aIWW4zjdrQuR+oz5a42wvorMoQiwG/wBGEfPiv3no8xxD/dMI0QW3luf7M3TUYuhIXU/A
n+PkS7LkDuzgQgJDkLoPOeZnxy2UHeL+ljdxFKgHdHlL1sw3ETiLrjJYXYzNqt3F+LZzn8QeZS1L
AdGbn6zH25Bz5U59qOOnaJ/Qcpj5vIeitz6CJH+GSSmF1FUSzijkFEqmDnoN7BtdHmD0kY8Yfj7l
avwWTIzRjDTqkHl30daxW758DoE8xBWmB86/eFxFlWpTWCCX4GkQl3D/RwDVN4LbITqkoGJh93JL
w0nbduw5vxi6dsBuEmc5Ain2IMLnOSwPYx5dRZS6aTzup/xbes1C5dtJ0nWo3qkGLgTf+xY6bvHe
BbzHLkN32DHO3smZOQ/Fc3EaeW/H7xl0W2qJtKR4pQh7smHuyAOATfUYZV3ADUQ536wiWG03Z2ON
xkKc/1rAZKWIyIXbHoYoG0b+URhIToZYp/fEVMeW//5D1BI5SeZ7fycJgnHqW9p8S4q5M5AV9geA
EyCD11zNMq67/qcKnt0moVAlIuyuH08em2/hF+isLgFy0q9Q+rcQLrR/EUh6e9bRGeZjML8s+t6U
aJ0KYJvNti/Q7UPp8hQDCz0ot5sLwQNzFX8IGF6bHCXxXTSmEq4W1myvGdzJRo/bEhSuZ5kQEFyH
WINSU+ICJ//xeP/roBXsNQ8PdhUpXsTjHSOdw98DZdjqzNLAnO7wBzgvVlwXhLmvyiaLoIZyYCOo
qvR2QuwDzsQwtbrkTvGEfegEG0+kpHnYaDw15fMoee9F5QRKjGg4WlHh7jg8lkjkT5JUgb12BFsV
t8Kba8m8XrNUMpzCIDNXDddOKKd2ixMzJGdk8KcnmqCkVr6c6b7JFYMdKnDUgyLk0hwKGEWOOZ58
05H5K/bJkhtLVBBij4FcrkJ8BCZpkYxvfcC9dMWEc2DwE3T9vxAhFWWKiKoqvioeQdXcUxiKOwuB
vN03LMI8K+/U448FfJHXo2mwvy+6zCM6zJC/hmVOwPHU9kdw3Fh0VDXGOOh3MlkoIRErLVKiMq9Q
hWP5WRplSKGNdmVyUnV9c8nu2nKXOJj0iAXh6Ey65H5sOuMOD7M7MReR8vXW2ZYrKFpkC97XbfTn
J82QU3TddaSvO449tnrpnXChEGr+RUPTr5lNxHhs4J6I1JMj2fX44t/ykoCXFEVxTnchvG82hxzi
g4MGr1WKyp6bGXxGFeM6IVutR5BkM3+L0STxm+HVDpQNwrqaoAoXIM0ZS2RxT7NWxU8jeg+IfYFr
H0SWBBFs/+EZNkoCgsCXRnfPS8lzR42G7rd1h1dFXu9yLUaloL3sUX97p3GOygtkRu/JQ9T/8zma
M61H/sMsGIHtIUzSCPlY3xTDRCy6QDvqt0sb4d3F3FIXgubLHNPMVlNAeUQc8Bc9dTravlf4IM3s
ePrfx+R9f2YTw8Lno328C5XIizJrsy/vbfMUWcuXejbFBJHxGp5D8CWfLFUJH2mVvVicmNPkGAHg
udp2oB/BGuc5F4RRqARLyrhGQIZWqmdt/pwrVaJKjRo2KGi1BrAVMbaJNVetutHWuk/STyb/oRMY
mg8wJ8+f+K4TAR3lIh1MHmi/EkOPxEq1yRYucD9krilCmSfppWnLd1AP+/rET3wI/iyFwdaT482f
uGTkmHPu7TuwwzdoVtovERlxiaXAENvV9FFdVGi1reXJgWsFHPRFZJttAxH+Kyc5JWWOSB98vrDh
rHXwi/Z5TRwPuyWvh6vfWRA2xpuI/yD+NFNZ4t/SS7k2lbvRw/jTywfkmy2ny7nlXIZyzIyP3I5G
hZlrLsP5osg8MiiipeNKQNd79gFUhbbLEhJpMdg9XJZ8MaNHoBaJlPkOVjsQqikD773jPfN3mwF6
1kXIeoFDAQe9OOZmvEQM6aIGxgOeufoPb7IU8q66BDhCc6VPWi9OM7b7s2BXGCQ1v2CoLUUjVSUR
5lxOflRVou9xDs69a8NWnJK/QAi1dXPLRz3AYtie+lFKwyOllZfiRNrIYpcuzyRa4Yqcm0b8gS+Y
fa7G3RsYJ1CrAei+/6f35GpeTKemwhRIKyGAv6Mgy8u7fqPkDMMio6UpYo5IfBQO+PB02P8xaDnx
ycrmOakNRXrSVfg35/px3WN9KSNoLZOmN2YTsnr57izRICz3LFpjkO3hfdoJAlAzyOSSdv4Xsmt6
bqGnUNBTMmxNU6lAQKmXFrz8ZKlG6gEraiWi+b7AONr2DUfyntqo3uoBpjq+p0kP2vhYCTP8jkfA
9jBIdkrN8YcpxbkIpkIBYR1jWjUNTumk/EANtkWk63nZcEZE1miox0xXosCVmwNJPVKzbSK6hGWN
gpLOiLtpWtz6QkpsQjD29OpCYs1iCaOOdWCEzLN+J0zVICVxYpdSpck/vk4y/oJ+nu70Lc3qu7Nf
N1WkCTgh/dxnOeh4tqT6x4hZAO0X/nCvoKHR03KkWxwWp3dX6x3BPSSLSUZ5C/8+Wg70a0YwPzsw
8zVBBMw+4W+cCfpVzsye2alOh3pAaW7bkz5WameGSJptkaKrNji2Y1j8kmk8ow0rRPKsiWmBPSuP
b+45UrfSuNIA2lglFZQpMhn07QvFJub57R3tJULj5WiZDMta1NSFUbr5X8D0XJTEEJfsZuxo4YXE
ifb78ZsJymglWEiw+tVViQO5N8IJOeV1grozSSC9uJQ+c79LkuVgiDUOQIp1hpNsFP2TXCetilW9
QE3ra6Maa/KbbDjnHtep9IuPwyAWuN0ftsVNkYfHwnUc71frU2m0ZnqFBc+JkHBC8PF29+2Trrpx
mfxDRplrhw9AsKRXNG9uyS13w6/cYeso7yWxQ5tzYLJ85iP/c2Rke5u+K70YsHMboH6OJEjzT+NG
aUokjbqjJ+X+KZA8Ecyjqs2vuOEAZmAvCDlChL2Kr5Tjwy+YgM9K+bs8+YolSVVbnusvUdTbnXrY
VcnvIhGQb9EYvI8N2aDCGss4E1IrC48gRi11HYVqvZcp9DoEiQtivLlHJAZHjXl0qLqDh4lqMFTH
4AhKTMxrzC7TXuhPFuTMe8iIu4VXwXI1oF1ZkU6d01YbudGnt13g4ojiGfhxCfEVuQ3O6BmetxJz
9vka4qf737qLIIcSiHBqEE3SOdTSzAkhT5QsPrLk79U0IklblFt9e8V01uk0MZt8iNUo/KBVylh/
s6+Rjecnpmewx39SWt5MOisH8GEpSqKlaQRXft0MksDQNX/wa+FkLyMJmL3G1DkshKbDpm8qFMgK
FbVviE+9h23VLjIilIMlaCTnpJgRD+ZMdiPkgOC5sANOySOGgnp16xbZ3M0KM/khSGodrYrXdpDT
4hSRiodza2VPotrN10YsvRHFuk4px6ed7CxqFPu+nWKEtR1l6Rx7JYxRxY8320w0ki3R2E2aAjpG
+Hp8hx8Nlsjy8SsQXTHvIkheHIZ7X95mAx4dUrH9trlsS7eqSviIeuvbffp1BPixctKFOKu4Qmg3
e6eGkk2Q5oLOG02VK+7WR6KY+sJRcZdDXI79oNMDapEzLi/xlZyN/Lm42RXIkLrFruFwLd5VhK4D
NT+mDD9BnhWdOKWV3MVHX+FNVvk4SJFW6O62aJ9v6y7wMMpO4/QAM5immljGGofI7jQca0a9Hu9L
183nAVGPc4tkKcT88MMj+VnQZ/xl2NAMTylI/oo8Y2d+H6cHb0xgx+vP1NFj2zBcFWkVnzSA19bl
V4s6TG3jHnD5jJMCIN7RLHPj1K/KNWXycwhrpjBJkZA8SneR4OZplMxL6dS6dR3Hn7Dbvy1+sVnZ
Go9lKuSwBAshvYg8eH4k26h+IRwDPYTaNHrhSzEXe0ZBYMetx0LKdv/032jHoSU/deRtam9eNESx
qOLU5MUZfjeKxKEehLFhTKhTdeRg7RW163/DDUPGIm0JizHX7CEJI+dg8m9DjoWHiUrZORXhM9De
lv0LqBf2rDRfzKjxUHP1jpbvJEAsNbr4h6QA6SFv6zzak4OBkwuZ3VnlhJup7wompYNooXvC490k
Vik5G4p8SBAJBo5KAqsEm2jQgvBhASF15PaiyI+VyjMg8c35VhwckSpbPKFWLPes3Naz2cwJl3t5
9X0nQY0zGVbKsrVFpl8zwKpkbYP6yd3Jp8mfK6lsj6SqSTsyjWvj0WWV0JAhhcq3kplLvh4EkCoe
MDyXa63zXUsXXATKPpjxSPUUrndjsN11cUv4YwJjjpSSZA+nVkXXkUj9qiVJ7U1jr1VYEqry9dCP
d4oA86oWuqyN5+vDY5OSEob9whg7Gzi56rLFWJmOgsPjtGH6C+dlzzDJRw4VvxhJKGMRpGutNK7i
m+mEaAIEfdqVgetesUtkAA8X3mER3hSHPsI9rLI1WXAUqVa8LCYehNI5x2kC50fMpHCsRNtcbfIu
zMOcz8qyYjRJHwPmV18xr9geHGqyrSGfvhJnyiNZQVDkC4YrpNl78XW9esUnw9ieMnguQNjN2gYm
y7+C5mXsJSQ+IQumb1X7zDylEinNQrPaLmZh/3ppvTE9/Eb/Cb0aVbWf7B22o43xX3xlTOAiVYJT
/ounwwDkMMRkXs0vPHXRuhCuQZaEIIdraCLsmuz7OrUpJFqDnhoe74FT64NOaYveli0Ir8uAB7jv
duwQk1pX/co5X0XIK7qjO5s2pokfZs2K7tkLRibOCo5maYwsSiA4v0DL1EHCxqHKMDHHh0aey+V/
e7UTedq54bX/NKYBvOYNuCkhRxONkb7VqCSsn6+UG8+w0wqth5toW+jkLzl2XONdu7jGAxqQqjGh
PNFs2eGTjfSqd74DByeF2838qVUcD+tOqE2WBD///+WciCDpque2WZVPa10EMi3w06302EjrHoHx
n1ppXyJsqSbtPlcaOzpvkNHITcwsDMPNdXoMHUjXg1ZKXJPvr59IxVGRnIXcJ03ZIqbHwXatsRgt
tTFSgxwg2aEmPflgeTP03iSzs/kbD1wdPeZjB44AJ8WkUFprZNr4hHlQL8boh0MJjF4dULACUHFS
J0GN2Mt1lszh+486npmQn8EqfEe9niyx7SaIvOG/oB4a4R2/uLLuBqNxsDdFXOfy2am0afRByOCV
SNd1195FhwwQU5MtWc00O0R03Ga0b43om5mvB5XT9XbroPwpB6Vdnhr6QXPXA8EqrUrg2t0E8rOz
o55a229i0NPHn4e9IKjGATf7btbLkKMiQIiuQEF7WtoDAOQlmJ+SiOOrFUvWOMhLNbBO43xBujVp
dGHgfFrc01eYP5b6da00069cN08VlqKfprqQ/vRbfwEK2i4fa+mDuHjI6CMOV4lNS3u9Cwiga5uo
G8Wei6fS+1yl4qgbvDvzQw+oD2KlM4Bj6Zvpm7bwvU3Yzqbm4Q1JsMT/rfUqzCXjFQnbL9CGbOVG
eVdTs45AmTcsRdF9WtcYgQ/aqQUt/ijaIT/aQ0hdcyG2HITNITcxpGBaO4jQ+Q9n7dmpaJJLKdaD
vTZCpxbJyKoPJlktsf6t80pRldT527zsZQeTVN+dninEQPWOfAW/GYjCnMotLKCtk8Yefdo4NRdP
psUA6hKCnLoqABQk3n1u+McI9kIaW5thnXsqu/ptHaLLwyc97YqgUrpP9Bu0Z8+9XBshgW00j8QT
/mjNikdzAaQkoD87ihsRHL95shu7ufihOpe36LjB5NDt4ku43r+Gi++tsjkWPf88j6JLKRaNNdYN
cKjsa4kK9QpE236BcWEnIesNB5tF6mGJySl8cOINpSOz8ejM71yBTXy1f9p2Ei/VIOx8zm9qulLo
9aKAHHj6G3Rzuf4u5QnSNQaf5p+5mWESWpfNA7z4lSweG+0sCwcmxsVYUxYYPBkW1muY9mXMpSqY
UOWDF0wd4pw6FXGJhTQabvlCL5lPieNF73A/kSmz8pOC/qkn4b9EaHjPwL7COkx12qtJVis+c+uD
a8LkbMnHzXbPBoxKB/+gdLdLZC/CdacLd1dy8NEqkdXTzCpDjNX8jRnp2Cl3/agf/vbpTaMTpBWR
Ywj5IODwWv3Ddvg+v1HR2vI2gbYOCa9XyEoz5WPG+14zsmlJXRLJ4b6ZuOyHY8RMFqjnJc0M+vRH
EZKgnrwUn0m/m5vkmN/B9Xp0yWYtF2pLpKKH8RNqioEG1v1651n7eiFoSbHa01W6OYb/dhZsiDJo
mvUKa+V6RRzMgk7TcyKbGwzXMI7A0WFEt0DYBBehgrI3/v8FlyiMQMZlnOx1lTxUSzfdy39fHxWs
O44wRVZto7XngXO+acLennQfPK2erNw3xfzYLTgS8P9Ls/JJ+lw3UqN4FW2RINlkL2Jp1HovU1R/
EKTzRszRAhk2LyOLIIeDgPST6vPx0oJWi3wvsInKAdtby7stBmygQjbGOdF0/Nq7DdqZSELJbNxW
psAMLJsOIPkxLSbNDiDiWg4FsufnHj5iGjXfOj+zfQQTV58s4hzpz3+Y7U7VldsdWWVxOS7eG1cS
HqKjJt28KX/isHXu8DjPjA6pmw7kPV5yoi9LgAs/DLfj8kPL183fK+HJto52ILgZ92opk56Jg9/X
B+xD7mHAnjvhu2JWxge43RunKeUq2A/bumpM/0WxoZuT1KOFGohBgPplLFnNHODW+BIqMjg/8uFY
eOoAASGn5E7OCFSpXlftvy2m6ZckSQ3ViAKBPtuRqZGdNWoKHABvgZAf5t3Pi6hPH+xE8QHSgbDk
mBgbjBHjXFXfyXyAaf+iuH8BBoBADwiwfbzeGryg1VlyAoA8dN3z3zv8p3r4+WEmAa/YCX4DCiJN
TD+iBiYTwFtChlnF5GNA9SsQi4kj9bJVebZFkbh1QHKbaHFvrE/inFi5zd0EzVm4glEo6DkpD78q
/z3Dyf4vxIcaLyOoK12OHoO+JsiBncg3wnzz1hIoazrDdybmVLNNpG2DkipNZzZGC4yEFaKihZXv
exwe+Whi4WryKvRj4kXbJJ6Z/clhX5Dwo2FG+4DSdmbuMrQhKUGqy29v5BG4Bqw3opFGPziQcZZp
Vl6fo6hiHR620O3nJBKGTqttrqOcW464tbor/uEjudpbYsmMm/N2URTQ7mCujmvrrvgPW17zmcB6
IfvG0jq6wdnu4oHhKn9JSMdW4jpT2pJtIccChe+BFaifrI+91idCG0IR1BgjrLnxskpk3UXcmGGq
vL8lOtVZETGmhiW+Y1g3BxDmDHDCJVelp+sNnpGCXKEWhMci7dBcEReF62utl5ui4TyHJZqg8O1H
qrk5zOAiLoWhYj3gt3v3UP4mkwqDJjzsutpcxwnGN4+LrZSQEtO4E4f5pvh2ZHJZqkQH7mv1TuO7
QCbwi64LhOpf66o7r4KN2aSe53Gshr31NE0x+Dy5EMzsmZhQFOd03+9b5P0RXicdIl9GXn/0SM4C
6c8Xu1VIoeu/a87ovGQE8OnxBVwpLiqyyhTPbWKPCLMEdZcB1JMr4jYLJfkkJkRNOboi9JpIbUV5
w25dPZHP3A4EAvlVwFjjUmEk68O55/E2KFb9dTbKziFCWvN1troHPnMfX8cebU4OoPC8QxXVE8am
gqk4o+mURyheOIqjQE0O0EyZv2erqMKbmBnyZ57ilXnR5LOQ/R8TnlvCOI/+ofDDXNT1XharZt5h
w36i1rzwcRyTRQZuFNwWXiM7cdY2NZWIaqhGvYMVhspP+qMtZ3vKkRyKzVuO8AtfF0gwrxpxFgEt
Xgiqoy++qBa9haeuzO3n5U0Kcz1DajJ8lC5tRbI6pybV4zer8XUhI/i1lt6bxQAx/cxQn4WFS5Ya
oyn+BdU0XNEvGm1w+qTcKCPHva8HH+ANa1eDr7qzlvpAg3WRzwHVYsTMWj5h+JByA756WBR/YzEb
EEUAk599H+tqN+Wb4Jgeu8mr69AwYTWfS0G45eoXpi855V1z/O1akHB1Z8UOIUWgHNasDhlB2nfr
1MemVUFsDmkRZ4PN/h64MyhxV8svMeh0PuytX8dOz2s2HCA7OjMgceAzyhhYc1j6jmpgSmSDa7f0
tOIe1CqwvrdYrc+8KITqXzesmYkY2pcJCewWSSjXwhhUFLGDPw7/+QmysEbF3adyYMBNbpl6wyHO
8RkgCVw9LydcwhUSoMw1XX2ZOaVO7FTt92vM236h1vSN96tglelAtSBX45lSIwVqzOzS6TkZpTUl
1Uve9HxykxeUwrz8IFWx6Iiimx70rN0teznElWcjRVyGRao9aBEV3FTCg6EyubZ4LJtBIFilVYEo
Eme/WrMS4PUCDakRrYrYx8fgEOXQu86ikqInG7mH2Sg+QuyMjjpufpyCjHQVONCDFD3r48CcgEVS
ccx5jKLqAYztpshTff/BhCBakno9vvH091X3uspiXJQkd67MBQyNEMN9LEpiCQmNHMf3lkEM/Ro8
kBxiKm0JJqCCtSoRwJR0vMOsIrLFFRiF4Mu9m1vr+FlBTvIr2dVzz7Ik2IGtz3C3VZT3kRMj6Hd7
X30c+8VaxfB3Y5GStvVosYXIpg0uw4PkGe/sFFwl4mTzAngZqhPwDFivy48N1CcA4TRvGVN2cuCX
PaYy7mXPf1jC4ZYLDxga9mh3YT2GL5S+Hc0vUr9xrH1BUEQrtUTaDHuNrDS58O1gcr8KyNtC8oab
eFtg7CjuEfGq4Z0twcJbtuqut7f3HmTxcF3smOnbqPG3g33Mv5aEFjBuQMdu5bAE3WT2NVAxdrsO
pAJfZsyixWadL2L51GMcGdzz2dKHABEObpxePx1oG5CfnC5LKyVU3Pz4xE1G1tUWemp0MPxxuDof
RyOehvR90cCgnTHl90V+qftGkEm/slN7MDpjrG13TyIbK9P59jVjZlaUKgRCGb0DIetXU6WkaRfC
xJmkpiIm4lAPkaq/vDkHECwf4Wn15BjHz08GEHuGB5MrWDjmHvTlON87eyoTfc0xba66NQbWSWP7
HTmOgSL11fww/Y/QthwzB8+YKWyum3bUIBpLlJOG5n/1hQwlCkQdcNOLqNL1EQnqCYIp56gsrhAb
HeDKPhv5yK6bk+BD40jyLo0dGHD0Hg67Ty8bru6KCipMjXpiN4WcWMo7jJj3UprUzrTsKjlNFSfK
weBuBp5bumEK1vODJdsMKyzzmaovSLn7TRla+Mam+SDh8QFm3HXHWh4HPftYwYQLrz8MTmiIVZUO
hF8A0H/+QGcS0dOXymbcoYMVFcR9hNFns8T6lQUGGhnaNPtDTk+sE99J6xp55nd850B9Dg98FzmQ
V30tOn8Nc3LkCWbr8a1CSltRfVZT8DQBSRneRIbvpjULtez6AXSerRMeWkCwTg8iGAtVqvJfcn/1
bj3uP9xxXjxOSljSBxC+flJVZF+hWl0sASX6A6DNUVNfycdEFU2P/rVwb+sH73OzuPz40BS9EG/Z
68u4v2nC4wqPk9ZmDvUaCTci9FoqMNZWohEY9fKO/v7lGJL9gk/l/r5k1XjgW4uDZGZWpOUsab7k
aEafDmOmzC1H3hi3WhAIJJmpmTVbxIi/EO1mfmAKEi3rIMxyIRreIumxVUh/B8sCWHAvkSoTVkXA
H2rPxXMMI30v5/61/sxMQeWiHiim3HtIve9pYwKxjmD7/9iSwATlsnQmYIQqV0it2S5k30PSsGgn
bI4UsddwCChdL6I6O8JxzNWI2tgktH0bZGuN8Do9PJAlEVYIusLfuJA7llWBKfS/DZBAnwW/fecX
0FneN5FXR7bc2mrG5K0SOV6O2lXRkQKgLs4KM91SdLb8rTIpgZljT+PzCfIFBQ4YhYDASqO9AKO7
zZUVIXJhH4YGGbf4vDr9+np1TZzDt2k4nTzLWHsppn2RRu9RPuWqX1lnU3UlYJUmuSbeN5RQnhbR
njKZ8D7xkLLloraxFjnoVIzlcxPypOL90LjQDWJ8K6jak5soPh65HLD9bM8txbbJeAHfH1fNanZV
P37jjEFBYscdTtCY5MSVYUViFO3segjsCHEYjO1oYOd72D+JvIqwVmHM7D3eJ9xrz7wAK16h0q1O
qQ28ME8EE8Nvs81C5pTK8V05YsRbXuIiOa/gDnBTHxzUla/XKZuwNVkS3sPBWOWiUHnPd6IiKY/x
nof56mKdphPzGlLqWol2iK7RTTYkppncKCSt4g/v+NX71JG34auZLxlIO9xCP/whdfsSN2dshETp
emSOVlC0s5npixAEHLewdxuujpWZKYCmNSlE+JM6N7EX+RXfyRTMYf3uUQoFFNHyA+02n9QYDIDM
WR8jJQkrLE6kARwqkYn4x1gwneTyhlsKl5VapNZvdbuesEtuo8v19golfcDdm79gIQEiOB84AXSv
rOb046Ti1rXVHpZR7S/eKEtPVPCL++yYcZSLdUbwdmX6iiMTAHlfA//MMQGqSa00j8UEJF+rRNIu
bmadC5noxAgxZSgCanthvDrarjgMru+tWe9RPjWPxP+bQv/q0y5d8gH60/Om6C8t7d+joY96lKZh
Acfb9MKzzHvJHlKVlHPm87p10QFmIdsF7Xdb1iCdV16IVPc0g8ejc3hPBnDHuzb2fCWsz/DewWdd
pf4GdXWh1/yEFQWKNVCjUeJTveATwGoXMX7BF44sA1G585g5dGfqUMAG5iVnBBlDmcBwmO6GkkRx
wdZ8fQD0NUQ8ZR6ZahyGvp9pw5DZKcIIO5wUOhqyRPaUQhaARouRCIGk+NpAWco+AjsfDWe3aV/1
1qIs/U50a98HLdDGLnPnAEFLk+K7NT84R6fnnxY9lLRrVtvRiptxWRSEuoWBYiW5OahhTZmXnRkw
onmxIBXtdvpPUVXow5BM1E73BRbPH2Odi1KgRKBP1FtyRn9gJrfuhIhfYgYCfztQE+BHYWii1g+B
XE9YoB3XjCbC5uZFfve66l0C+h0QHVT7NvhFXM5+mL5/en3C2LEPyBFLD7IP7IAkimbj5Dxy0mF+
JiBPgNAQaFxnxX+hz6ftLGn0ktkg6WVYoq6W33eRlZ+qOO24TCUZrDEC6rWJej/grDdqcgFjev1x
1ZiCft8cmF/EyddDqF7ia713VQQe+jeJoqaNlnOl4le9CeXOlKLFMiztdHFEf9iGgI3OR1P/sOt3
nfHYgKfS9SX0ppApP6uwRPbbk6UvSqBNpn4xrlFMsriuRYLVulLwalMzNbkRVySdEcPz0vwyKvSh
6Yng5Il70DX6DQla/4Qo603Vwnlzhcdb+kjSKrWitaXQ38O0IzipX5EQICZVD2EZt+Zd7v7oPRLo
Dn1fAJ3KVGkDn5KHsmZuV+yeslzVZR4FkttNbKt9Bik8PKQm6eD3abvMNDWhFxxr+F5W/GEPcfuS
uBYQspXWChZHvrYVDVF+S2wvSKxS1QVQovWfqA9qBrrMa+57Spyz+GXjQOHHE1NxMd1ivLDPL/bg
dEHOnlkgEALvj3ng20sJySZVr8Cw34WY+Szy7bwOULzuk7S7ba00YhMRWCttf+bdh3UMugZHFHzv
7JAnUjX/cFZ1sQigACnfBRaPXhEs+SMg5uxztz9BGx1tUaSSPmNS9u0Vzy96p0STX03OSWTPNcZn
AF3QV5//Wv6p0ALcC+KG7qbus+0nuhjw0OTbyTwBJ8MmyetLFTfkpTwfPxvDXLQpnITp7KHDLhFk
5KaM01IP89vP/+gxnWr51ZY3EUIUw0lrksN1bCpr29cTJvsCYYY7OS2hKRZ62jKAzMKzCk+d3fiq
4G47vUmN5B8BuViiXUnTbkBmniLBGVc1krYQsxR6GcqT8pK7haWuIAKF90TTIppWRBquWWzyoSsz
fmDU4E9YMw+VtOLLjcSv854PeHI1g3F+0g2tKMtPs7d9PNeGL/4dhMyQ1ESQgr1tzNm0d5BqpFSY
3vqoyjXLRj7SRtWEnzp/7aLvYuEgLccItWxehSiEuOX4RUze0X9BRkVGw+wGpFfQIU3ekPXMdh4z
qxvZeno2gbXAUImP4w9GGL/CtQXsooP2i6rHG5itH0b/qX+AMpoPCwHTXKMu/dM71HouyTuHcLBf
jhcNxMZmeXR6JescnRzma6oN+Y/TC2yBya5TehtKFkarG9Fhfn7tZBYdyLKRs05oEF8b2zJnTwlR
87RvR9/QYJvru//I4BdZVFe91b4xAM+mOIRta+Hd8ONNjAT4IGIBchhEzQ2WV7Mr+wXPkVwlm0sx
bAVc9B9csvsnWGx4awZhUyx3/1cJRVMD8H9szpvuE/IbQUzFUycUNnsYrasVhoLP5XxLjqqYyIfb
yGN2xaqyO7batCDhJ9hx+kIR7dRhDPpqCnUP5+bA5Ol9+gj/9zw4hoFI2hZ9uoDFT9e19Gy/9VNi
R2OuUv2KyBU44Da0Gbwm8tA6uuWwzLCG36WKijQDZTrt9XRMmR/ClrahGWO02jhn4PnuQL5zCcMX
D15tXhHGYPvKmb+9yh4bj43dCx0MFLLwnow8Y/KNgZJbW+R3pIufmeN9gAfqCcqyL1V2G9XZjhIZ
7T1Pyr5c8oZGAAIauV3VlZPLINrLTPL1gF6RNWN20PO5OViBGE/uPzD92hVLWPGMFJPbvwg3HiGt
2p1+D0+8gwfsInUVkPeRAINzzfWmRI51ndCrEB9AmukhBg6CjDKmhGYlhPXUR+mBqrb7ozbrIC3P
AZ13yZ7umusRBBTCPlfS+yZDN9+z4GbDi/6rj9qC1LKYb8qzSR0J73zevB6UDyzj0lydVZp/O0xq
nvfe06JXZweP9S34qKB+i1vemA6uztt4Pkr50glFklqkXcIWpyifHYV3xx5/XxM+AGpx99bI0N5l
2UKC7SapIzMeUKFCQHUtieVm9X6npcFh60TS8Aqv0Ak39LaEKchY+uegRNby9k68PuiaEZscncYR
0FbGjkJs+SeGcsTsA9NIxstfa2BwHLW/jVUZ204zXpRU2z45iIy1ugM0R/91XXvTqSYqSv7OkwwX
ufKVSRTTZaotmIQqLRlsMcbRVEp5H51R9RCphfz75FXYTTSDlFbs4/ApQEG5sWHNJt4Ap6HQQuKE
z/49ZixDcTYkPT4tS13Et9R+tOXYh0po+NeIexDIyO+g9f0PjiZkT3FGGncyrUE9pbjSqU9+Kckn
dBMBGaD128Il4/3QWGQKNIHRqmi4ed54u8BC2nxRdzFbaygg09EZL7HnKl/mvvQ/Trkicl3fKA2U
WNTc8ALd6KAzXoiC2m0iQ+5VidgLLC06ZYXenrVp41aDT1pUCejyhqgQNhIy6i9Qn9NNcrl0yM/a
chUbnbJvUS7ganEa0faGHVT4WhjRBKgwXHHYzSOOaHkWV5IIMdRghjkSFPbJn5f9RZq1bxadP4NS
anxGVj+ocw8G8VhIAO+/7yBIQyXW8nD35qeVbysgFW8mHerys+qBdRFOISbh4xzwP2sWHycsdj6O
qUrkuoT2LRI4JwNkijizpn+ewR3ju9qNypVNf+eA6N0UuQukN8GUpD3ZOEnRWdLWMdGnedDDjqiF
3LySzTRpVnKvo4cGlTLVe5v6JwYh2nz3+0WTsrITqQT2eoNQu2GDXuAIuiGAkS6IQteq3uOZyiJo
/n5evtC96P6JB0Gs24sW5GDHsSYTKRKW/Hj8Nqsro463jLsc4OqxNaqrtNOqehNkv0d+RuzWtEvZ
VnElnmgQzs/U0lCeQyWBa2V8djemrvhctc5AiURZgrsgfcctX1P7bS9S5P9LfIi+PLhnI3q+p2A5
4EZ/nXkFAmNd6doVcWi539i6Rw4ZeY+XVRwTXEvRaqu5GKfSKLzaGAPPv2uiqcD1FWwGjN+s/i63
7LAuswKclDQ3gdzqdKqafkz3Vp+6e1B+WnybiIVEspEYM4kVMMD3zUeopFes22s2sX/jKkCZFuuQ
6kSkUuY/HnzrGQ5cGqRQf0dPhCCSc1JU/wbUkWxvLAp90IasuPExh5Ww+q6f1q2PGqDHMV/ycyAY
SwESVuO/vfFbxeyRc4afG8van36QIYEsqS7lvx8bp72cLhu1yY4+RVX+wlCdrI/ewmSXHlWdr2Hz
/Q12tD+th+0MKzAObv+7zxnUmRLotmnCzvB/ozDtMSpKHNh2cNRkQjaJHQo5eHvo6tKGbcrwhfsl
QRxnr1ZiuXOadctqIZOsK0cm6w1m3VdFFwoiV6D5IvVE7+ApNgwfZq+8TXZ/OXGvxoFhhSgz+cCf
3nzUb0J4SNmb4IsdDaOGVZPjk1Bn8yG55BBZudORhbiSFIEkiCsytVDprRsW7bR6ib0x1gU3ZCdR
fIwNnnKvU5eTWvWjSdY3nGGXvU20XoqqHD1eTBiqcfZ+Ij5KG0zj5TEODGo/gmjVHoF0lkQ1HPJQ
y4ENKHwZR1lSbnx9s+Thw/Z5d6KGLxxECbNh2eOhZ8+ek/M//H91LhF/0Rf/9zOgx946rwkLHjYN
xv7D9FCR2ZKTZ8sfuWBrbQAw/skH8vAAbmtcGMxDWeNgBML7KPDWxJSl/4hztwqDgQWqPi3af/fT
qE6fm2QxT5qnxgYZINjf6f3dIFbvTYS+GuvqXmufvUwoDwpBae8rTKwu+yyFax9WUgBo9SQ6HtPx
wMp2P86rCqBt0wl2PXhJlPHrl3K8AuHnIVSupsuSMCDRPYVQqzXm3eNTlt0RvmK0maTdLf6os6GM
VKonavZlDjVubYYmOfn1kFz5GS117Xtxh8XyY9CXAT5QfgpzXvLy9iXPw8aAEobgHpRaWtqR5Sns
fJIxgZ78zB03hb6A4aIn8Xfl0FbEg5v8oPm7EWPiTehbAyOqjDD6vtJaApfhQleGS1POBFg1b4EP
+QDUNPp2wTNKc6rT7KF1kFGptGMJudCX7+6HcLQTlGxw2xZZzxhmicRcQjGIq9z/AbzoiVvk5amE
uyp24jzuxn24oWzgW6sL8e+ML6sTtXUWianrTnEkNv5CLdnitbGeWYa0hCdApOnOF+3w3rhX9Qx+
hRIwnEbrrZ+n6swH2BdWfjT6ps27ayuiVk4a/SdXVW1UjOtUZJXVixpI4N/M3R3TPAnZDnYqUmCr
Fjert3b6O3hC/E5jbchr5Ri/pEXIP2HTbGd9WcYjFQQrTWWxr4WRkhCJH5fQSRBjRs4YB7Plq2Qe
E2I31qrWuBJLSRLWE1sqsEsbviv30YXAD8oKLS5KGEZ3S7arcbPXNLifiiJ/WJqhwbNLrYBaDwKt
soXFVnfdk8SbWcGlAcg4hcVeO73D+dzbGTR8ZM5qWBHGNWQKG2wPA/r2dudWT3qCLjUk9U0VHfZZ
oKtntrEjnJKzaS+zHY6jdUKTzuJ2ZbiDQKozurqzHiGMpQfk9XBau+BoV+InrkZ0wDl7zZS6gSSX
lAQsetpW2ITK4+IfKO714zLjwUiaYpgSQKfGS/1VDiHOI9MslKKoh/fFd0BUqfHkZRRWGQwko8fp
WThClqG1ZwgQxvWDiAiSWcyKjYOsIjZ4aLrrNJa+ReD3C9lP9Y+BImHMzU2BMUmzG3QpTCtUXxOD
D1CpVqUC9/JWaPzyeFGgm7NUokOkk+6P7yi3E6kzqsyTbE1TLkPMp9gaezz8Sk5aFBruBbl1lS3P
rrxXhS4eMTq9KPdcVqFDNyUHE5FY8cyVTWTJM/EYDngrW87aEDUiCNobPoKQxnz0zxNjS+agefTm
R4M7xM7W6cf6AHyOe49ouB23k1KO8xJki/ZeuftJK3BTzqcNSIs2oq5tGBByBv95pr0GmNnZMMcn
IPMGNErC5pFjCFODbcIij3BW0U7WOEydHR8kGxrBobX4P210hcSh5uye6TIsllhgudxaWOB6V3JE
DCQfjd4m18lhVqU1XOylBevk3Mz0qfiVzmr0n4b9UUnqj7fNcriLNatL5EVbPDT2jKBh2lW1M1wt
UqLHPTzBL6h9ugfKT57rEx6YygE34bd7/vWNj2ibRMnipiP0UDjgUqOSezdAjOLoZUKDdffCpe90
MxeCRuXEwkJ8MYmR89kWsKvaBQOMyJxPIimc0gnHmqTIOsdLNMieER5WnzD853a0+SQUL8rzFcJD
3nmVAAJ52iIUjL9PZ0gpXh0D9YMfGkmik2tI+dHN7ZHUgdd7Mg92PoTaOpq3bdVBCAMTq2kTMnny
q7tDnY521QEq/UGYBc9Bht7Oy/a9/P+Zsz+kIWk4GL0/jTnE9HFonlO4sEd1hdNiypxbcVz7CaXa
ALmgJ1LaQVSUOVoo2FTQZMeSZ/2/ohq0kwTPrErSOO4t4pnB0LMs8njAoQ5H0po5WfZS4dUhyKW6
WK9/IveOUODdQHPLhEfi6cxNpIejmtdoUWLpAi+24voVwJ2sgExU3zyO+Ix5ZzVoSQ/wI54YxR6b
s/x+/gky1sTsx2OaJiJKmgM72qmDYtVWPTgKjXv4Sgaj/iwkb1dG3FjvpHjot8xhR4yYnEn7ln96
jGdwca9m8JrY1D/Q7f2yyrhDGiXHaGaRf/H9Imz11Yw10K+leb5WGg1bu+cd2rTkhKtfP92ieM3Q
BZGM100j1voNDwAZlga+05XX2IzBnRztN6QBIlWNVs9D6MPg4bAewKmy3WI7dl8NFFvjD0/6wwKw
/4oWsjS+YR61JViPwIhnqSB0g3Jvd1M6ZDil/Gg3+G7/2n6f4RSQyjpLZkRriC3T4awAmBTjqfPa
b8WwUntxEpYiLkSEi1+MPVd3CuQIqWY9nJrsiIilmbSeyeTVGM7+evnsp8yuVBACpjPHa/1wdSsL
m7VQfJLgo754+ZhbnAxTFSqXGZQ7I2bXR4zLFAE66Mf9AIWBfOUDQz0lAkXEIbxsSrsjFWY0Sajb
6YGwB7Y9ToqO81stoDF/Bf8NRTGY65HV8asqNjxgsRm3tto7dpc5XRIWIkXSuFO8SumBt8hYl8DQ
FUXwCCpsiVGqECjVkjLbsGp4fzY74fv5CDpvCob1q99mwX8JDiRy3ppfPVOcyVkiPs7IKvqQ63v6
LEtqYPkUA6UcxpYZFcD5S2ph0VOf0p0lJghqCoGmrZSOITtpf/U8DgYBI1ZZZTeiGDwNEHG8sad0
MDuXm2B3sVadzUxYt7/aJJYQ8XS1p3WV04DjmGwI8kZluGu8FQde4VynKV2GybeKtRvI6SY0aOpX
2PIwIfgjYBBalZ89EKCyy3jxpfvz2CWnbTdJ5beJ7z8QrOCiN7lfoLJy5V97zGsPG7DoAgWVLPE9
THHmuV3k8dJRbwVjpyPfApEoQq9AAI3DvoW1B0g6LJN0wLQzxBDiQphyva2/WTEpqJc9YY1ZcfyX
OcQXdI6fu3KUOxMqtfaJ+nCULMgl3HXON5G7PGmP5wjsuuA83buYtzVPEHUsY8FYsUEEHcTi+mRJ
WpJ6sIJkUyIuWzbXPhE06kzbm5hGzOoVbMAmSEXfm9W1leBaRkfmKL5TBjN/4Gr4njq+ABC0sxI3
ws7R44vCuXgWSin4JLYQjo0QdhQnNuMoNLZ7LgjR6UXswUwhUyBVXLSTUihzG/z3oncQ2kd/Hp6o
fCrHGb8joYdpLxiy5NWyLxWQ/AzBYhfADiSAOvN717jX4ZPCov8hf7ibvaNZquMVXTpw8jYkxe+G
YfXcj6wSBTlygloM7nPapW/Ep7yTiF6XG3T0Fr4bCFmVM42uIyoWdULQtXflgJT6ZPEhw9miSh2w
nUElyi+ldufay8nYC9esOGkFU5MsEpDGQNmjg0LA0lJXAdXMqfmIVW2Ao+jaGsi706Pedb2BxoiU
jp0RvyGWO0AqLNUFwAZ3ednFxAdxPQeRNlPGrr+dN2fwnxx7aURpQ3R80s6UKDOG1zzNq0FQYqJz
S3wFyY17Kfw2Xw+OTe4E4FU3EmczVyRY/2kBlk//M193kTlobaAMi/bnpqdwcsCRjpyoApb005J4
oz5E1lsnBs+9IJs6ndSOkncjC2hK/FrQMFZa3vMuhZSIszsEO4A+f4dfKvKXhSk5kbJECyHMnfUO
93ZcRaaYpGIivhzg5emcCN1mrlJcN7piy8E7Hp+/clwHGF7vR9XVGFSTnQYwilKsU7YHyWQEhiEt
UBH6hZq1cu8lvHwKjQsF3uY7HBfNoVuXFy5FSFRuQiq/sAHZR307EaASRJeQ2J/lbPWRIgXWQGyE
fd3De0l0oS0Sz2dt59R/Qo4ZlkwkQD60hYwn96GJ2ZLI9WWjfpDM3CprCPkOkO3THaUbDMIofVqP
4+8gt1IAFvPtVan2ZNx+v3P7fLbva24RXw6XnB9fAEY/9PNiIa8vPwpeL0GrSJhsF8zV/uAIv4oS
uvwACeDXarbQfbPJvyaIW4MHv48w3d0rImxKiOfFyUqDQrsLMNEef1X87l9wPgx4ep+FJF+/wKzz
SvtF5DvczBr0zX5fsl1va9owCy1W97drNIXsC+gD1oFF1ll1ASvElBL7fcYSKD4X7VOUd36d8igP
gjBCNdPigquJTi39QIsa5UouNJPuedmbFZEj3VA1U6nyNuuBHAllSJCgkF12eFL8UEuuHTxmwURJ
uKHwD5y2/sY8fjgXfIPGa3mASWYR9umkCWcMNSK5KhJacj1I7xaF8bA67FOglXofHSPVyAh0qbna
IZzd6WlPjYMWPaTf1VX20ZPGHjcvaBOAZMfT0cxCXvBVZkIkPG11K830G/AtOzD8ClZeYXCM1XxW
7MIBFFYOmW9aCThuEtj5yU3PLewZDgW3HzFr2GA4G+f3KKRR7aLhOv0dpXjgt0VshOdKcRZ8Hi8e
OL6ezvANy5IclCCLoJQA3ybH4PdUHe+HjFT1VZWGgpbKbWDwfLabVrziNrIC4n72EOZN3DcH//kC
4OTNHYT8RlJx7pEHjK8FrU2MTEQVliNyoSWtXCk3C25/Hjt8jKMb3HBxu3jwjVrY+QDIZXgbNUUI
NuBFU7MHD1G2z0mZbu2YWs+eVjE3oiClDsT9DaZ1ILOfXctyXZeT6mXzrEUuSo14OeECARjFfIOz
XwPTww8ZbGOiqfmSrvSlcah1cbNBse0au8TYCC6oGfiJfQsLw3YRnhPNb/IkCFzZ+VzWqY74xUii
TOL/YeTxUIAdjf3JQpvN+dv9c3eSvGWkUnee3aOiJtzxt8zukSQyv8N4Mhkbf1aKaollDegqrneC
Iiu+/GBx6o+eftb6c7nSxPkYiW1fZoMJzNB2d2JCCg9DBKi4n52Ntgc2F7YpBb9qxGBF80fWbzjY
p7ZhrJ+chvUmFri/DRGbRu/kHaoN/HR/1CVkwXXzv5zeXfft8G3lY4m8FJHaOUiGZhGFRUx0SDXI
36/jFA0n46rvuqFiBfyfFEgGFB3McvrudJW6yPrNr0zlXwel0gGrpfOrdwh1HCi94CHzRKctakfD
usBw4BZ73ez6l1EPyiC/H3IXWrqFEMbQUwitxlq0V5MfteRtw2U9v6HtXejZtQHEL0xaSm2dy0E8
3eioev5Zrl7sys8yDne4hWdCaS9M6w5t6erpjf4prv4RKJ2BB2p2PlOBDm8FT2N91YKZizLE7ycN
spfRNmIS4I/a5nNChVg9HY45yIiYWFIc2kn2bN1embZwU3EUlXjvfq4OKY8el91cdTBWq9iY4ujm
F0Q7FCXCoC0nMJiZW0aUty5xjAuuzvoj2v/3GPHoBEwhXYH8gvNo405WxwkjwsRDGsdQkHkdLtCu
UfM/f95R+Tn5d2XColagmhoSzOCMKVzopZEvsnP5D53/QyF9QZ5Bq3k68w2NN07ekm2xmKYHweJL
XIFGBizDewqKfwjLe8K6nGH9Ks13kOhbLIrB9zLmHmhXwUQ0yV2HqNnRn4P/NJb5L+Isd1mWlEdV
HA8XzmTlxssrxcnXaVgro5i+nTaT2NephdSgxbjUPBzCg1LNGIRgnco5eWX4lQ+U2sBjJtuk9zXh
e3NaLXs1jSIye3/aQw+GRzxYrX+JtmunCzoPCvnJ+BoxBzhUBzIubJ8IvzSZQZAoBPWMoSDZw68h
yGOQd0A2zArVg5QRQU/wHwf6IbNdoeT/h018pxn3SdWVcH32fM7MirUx5B4VgumKmucCzG5ESbnj
onSu2U6gLJoKGGixF0QUOz77g+cj9c6zR1qNRfXJjrIWVzt0Gxv8yIUBuvem9AGAGDxFD8D2CFXa
RLPCZ5U/dobPHyAuh4Z0FHZcQoLVR2xy0lX0fnNYiU09jTukdUfL3aimltCqKw/CcAEitkAQ8h0j
CrPrc9qp1i41S9PzzS+/VqXVsiCidYRIowtg05TT3pNTC9NqXcJCGfSMUSHhxWAIIBQ4EuZldAcV
AIHzfCmOF+Hrw3jDFFMn7ZoVbdtoYV3EPcElAk39avNKDAUa7A0BI8h6wwPIikm1Yi1vLcJy8tiv
sLagm37KMhwEFjl7uKN7YYsoCeMeSxCjjMCkuB7Sjtv/y1vcBTz9IiBP1gIlVIUQILLO3nz57xye
9Hf6SMJZj9NEyPDyKCI1DtfohlnZ1NTf5xt6tKFIgFL861liSj6d1wsnHqdwqDCJht6tFWqU+DAW
DrMyyjcce6Y8ebaV2zLRRYo9zisR7qc2YNJo7xhsUwsoXOVf9cpS4MHqz+rD1MyQluGv6Lp3Qqhc
jFK3ynS7jOnZxFZPzEuiAHeG2QYKxLmCiWeBVfc+Fw6Wgm5yIj2lakSKW8kdwcTafS0Xy+vJsDvR
xJHscovyDFneM94NISQ/0SLsewzeeBWBtSCVlItAVSPXAlevKxO2370E2ZNUehsikuJONxjO0KuV
zXfptWalgLOGElYqzzp5YF/dw9n/rhKZZwCR19W/KrZE7IklYZ4WDRV3RLnv9sneIcua2I551Oyf
SY1ljYudRUid3e8QCd58J/JSxaHt8nUHTjDTigb41SRHucAfXV80/dJXo59a30hs1bHtYcK854Ps
CVwu4nYqFGH/tcUekE+CybQL3hK7VJC/2Ug3R5cqiRgRo+prrOTK05OwWKbynKS5ZyldwYKBaIB7
raFCwwiJcRdmui46GtQHXHiRquwGZ6qeda4yOsUB5iqDK3y/tPzxYDBTnGWiLkVH5nA3exJ+EoHL
pLDC7SPiwNfIunhyela8hRNMwTLSyzFoj6SMZXkQePUZVBUmd95QEAG74GpFpvLgq8TZ9+XcZ7Bv
DekwI2sZhBrI0b6n8HPJdFdH4zBpT6Xao2aPRxcTU+cgm8NtHGkG84a01kkaz7cMcdk7vDBPBhDY
Jijox7T1d0m++7nesvVluVGV975NklpvHzFCSIiSA5gZUsCWfXLLZ04v6Zj3YYK4br8T1fgF5+dm
5mhDpWeZh+zd584ocyGPzB+bkkv4LjMDmCTyfCh6VSSPOY7ASi4P2qUy1UTVWM5NEPDRl2+wP0L9
bLXi/0Hhr/Ya6JFqO9H/BmqCxBQ+v59w9b0ZesxNBBmQCrFyhUMtIG4YFwFTzGIn4HhaD9bUNs3Z
LAcSM+qqSBDkB1eksvmYV8Zpusj1yktGP++lMtdhFqfcSte90CGIj5GqYjpYb2RO5paoTK8fWtFy
GQtbqk1MrdAbb5x5OUmbbUk05gYABP4wWmJEgwXhAAWXc7SO6euDrU08z6wqHmVfwM2qHyvVX02z
IlcYGVzG9yS1AyQIuKVIRc93lEFVz2GUtyp2bTYyQXMYaWBHjtgVpAqPAvHw5mFSAmAPo8ezwhxT
AOByVVKRrLNoM/vYxy3HrklF0Y43OgZfaoa3mCGnDUCOpqVgdxW0JSHTuPKzluB7FcQDa2fqK92C
x8WkTIN4f1INNVeD2efTJpkX1VK8Opi77lTmXqIy27pLWbaGR8yFEaZntU6vcBHSk8COXBAYhVHL
bsfSaaESsY9UVp/Hmny2jzqo+CF603NEd77ykLlPJqdqZVnAPoBdjsdmuw5yd0yjGDaZHBJgl27+
1d9qZS1UCFFwXp4BLQp1GPKrhK1UzUxWyTuC80e5JgHtSwV5HFrVldzTx7RhuZhaNGT3U3Uel4gS
eFuVRivqGLlCINf3SuJXoidbrhedK0I21H9P23aTebNDcpIweNBolO2wnu4VB4sH4groCOUzqUik
z75uWLTsJ7vZP7ckNKjQ289GuptKryI7bOSJRotUcGuIEfh/H2yWRRcLnDmP3VF0w5bWjXNJP9Qb
gNfq3N35JGRLfj/JDX3pMTSBOgcjoP1pZqJtPgH0DuBbmhZ0KuetH9V75hU+UxgB4+9QB+e0RcAe
2pzbMuxUHxcMUupDbM4CCSz3kdlgVmLQjKGdKR4WA6IZ5nXhrmhjSLvEHyGoqp62FOmZ21pxrKtC
Z14JLVPHcs4JIldf8Vz3DvLRm8cYNxFkxr2bvcqP8gY7oPvsaUOZJi9W+7nQcNvWiG4gr4rFEn/4
IrqLhOLHxdgc8JpzJEeDD9eJo0vp9OE7IjEbZ8p7N68YC/Oiu5UmaAWkVi1frJFt0TM/YT26mBqT
u0CjRXOfS11mX33DW7cW2+9SmTJW3nm0Oz+lqXMwjVnm+Va6q9uqdPtBYhZ+vsGd+uDR7DsJuuOd
ZcsdTZ9JUUts2ry47YGq/0eFMME6KEZwczgRTayBZU5XX606v0WVbQ5Bz3gkegVJQgZqRh3CO5dk
7S4JIk16tsvqucTh0ks8h+LK/YtjviJeivxjn4513Ecnie/EzwtflWNUOfd3rGH+8RExZv58Sfwc
ePRcB6xWrP0PkI39VawBaWyap64ztkkbP1zBJgDYwNc3A5Rj5cG8I68bzLWNImVdv4KdAxiVUpt7
1V/uKQqb+j5cVAqjPLxJjPJheV2fqDSzYPkTjvGBGMUm/WzwLZeuUEalMu0yJa2fCzE3vOZKGJjY
nwig/6050h6vPDIKXUba0wqGS6LScH44McW+h3SWVDm/lBe+8yMn1L6DFRDNTAMhY5MeR53Fpngq
4XvIDO4KyJ6+Gm8AwdRj0Fvcn2T0bmJ5SUF9fHr1P6kecMkDANMSgovR/VK9j4bQDYYQGLD2zFJ+
xPadV9ByprlPxB2QQSgcFSNdE83w1XAVyHXan+sUXfxlO8oT/tsuHSJcc9WoeYZyd015Fkq8S70S
Ibxa/WbqKutaWQQiXWU79q1xuHg/TroJuQKCEx3RLSNDVBJndtvVm19q0LmoCYGzSaUx62VUY3tb
wos/vpbBiQ2kMnSg9BIzHesjcDgtyuHmRgajrxZiba9Fan200VaGui7rekVpgb7GdnP7FZpoeyb/
CFnFE9LLxSy9T4biNDCgzheJHjxw61Xg3d2bBQrtv325FHcW0ZSuon5f1TDQiUl50MUQRm7TqbRS
gltfDRTHkdjKkQrBXmFBD6EMNjO2iJ9JrRwZApHitaCInYb/FT1LQJ78AH6AnSlK/Wqti0qANrZL
sKlZuU60v6DQP23+lUJ0CXkemHnL4ZFkusLnnD9F7/c6nMJeoXOQ75j8z4lZHmJBU4dufcwqzr1F
wi4R56s0xT67XWJW8eqRbAjowwFwBebMkcTheVfDxQDNQa6JV6Jx1ve4EFWOfWLXnmXcSl+W7pen
UimkODUrRhnHK8zyKp8AHWL+PsRk3msnBIc+6CW/a/jp9BHI4qwgxYYxpqeHMJBLX+crWT6gvtyC
tlyrCa9P+JswJznbys/lyEoqzjFF1X6ty0qrfM2tc8WUvLwHAGOtBraJH1Wk2sO0xIuRhMr80dad
4+I6m22a6ZKNhxfd9gupP5Br20yxdgjEqFXU1EExtN3mxepYJXI2WbxLyGbT4P+jZNCfb8BMZcT3
by/NI8zo4xvk3vUVlxVmlJ4Wsb+T9xiBO87+SFOg4v6XevaGZPRhONUVnwJNnQunAVBBO0yySVXh
+ZGZ/3FSHHZ/Z3iG9jmK5FuqHu+ms0VAJKgQlS9jbQ5WhZhYHEVVunTDyw8bs8fRV2NbN972bvqV
hqTmarLx9Ba5gr/hgXRfUOqoIPP4mXc13kcH6/FqmMWexEOw+OgTZaKb5Y5I2I8QbP6t2v6aUgqm
0By6eQFqgOMPqHKZTZDrvqT9uTb87UefaVQr+xjvHrvrRTArx0xJapCYRgBuLanqVSVyjks/hYcy
c6JSXnNbjnQo96gvvoHvJKj0V14EWIZHISrVqUXFcgRO5h00UFSWDvgiRDg5COP4OYa22DLNfU3P
wlkHJbxGhs+ioZAR/9s3VhgZ3mxrvkWOdJ9+dKzoq892QzmvORtIOoh3P7ajfgwGRgy4sep1QP4c
CydIueBLSVIgEOqcqXgc3UiD8++cIFIiOVZu2/820CDucaiPkjcRgZ1pU2cw0lyscw2XTiP89Vzl
DkCOU1SkPsQ5vMdPNjdm+zWkm3zQ+8JJ/vmNLlTe2dZhmEkRYvnbhvivtdJYlv4kawvaj9Z4ioz6
zIM9v8AHqHzNR+fs2UWJWz08KSfIYk7DGRyC9ERl5eKkI/VT7WfaL4gT5zKgqODeK9cLCsyST3nZ
Q2i2FmSBKZ1h0YYShonD7pGQaFX0bofbI6716ljZx5IiBy9G6NF4fqDO3GVVxkFFmFwEYDDKLwRV
4Bn+7CEE2GDXP+ZtESIEh7Uvssi5tUtlfDBYMDG6NhqM9s2rD/A1CfZ6AxbEYmAOGLcfzva8xKpY
OBhanGrvj4eS9Ki07mO/UexJwK5xnCNmtIYTbH70oYjEViqANdPluv65iaX7UQXDHJxMGxmy1+8j
gZOjrlnCIRkfUoF2cyHFI0yJP3bQLaIvU2/K64S5WgaHzXQC11ME8z89weAwShYBGwRQ8UU/nBIy
QuZbAViWaQ24MrwOrFFtH+aV2z/ZyIrRBeHYhr1hXD5QR1z+MCdCUZf13AHVLwUEIuev9b1+Wmbn
65BEBtQjbuIECiPKFEhKbspSBsH6bGF4cD9vsI9n78bbWN1AitJciwg0OQnZ+JApktwcZFY66jk7
uwjbMWJUoaj0TaDU/MsZS8RVYcJNoHTcrJV+vdpEhZugvYw4Zgpwa8i1/i1dndpltn/NqhJESgaL
m4d9x2J77fqKRfbONum6IWLhWQDrl2JUtsNV6GoeWPqYisb9tWMMg8OP1BS9q0YUmtitIfkiizK6
cY7m9gsKx2qDedhz91uGdNDaE8wN/SwVuzYJwf6TsMEbx2cG/QLaVMsSIsgHGr9QhjrttQa1J5X2
uFAjnnwrNlX3NNGVFTpcHZ6bjOAVMTJUVVKsNQBC6v8JGf0E1/8bE86HpQiD5Krvpy+qWI98WN4L
SdOcUn4rrg6ASOFtTNLTkXfUySe57Xnxh57Cwp201HlE6wcTI2zVjMokqdBQxJZ1nXcpi8hEonW2
9ugygizu5CzD79hmAXLiyX7Mf7qjm3/zeasz8f4VjjN1tBod0Lg0yEA64N1GKmbmb+p8guhH2AVg
j9vOU3Wl5ZqMVTxCyC8pNNuZHKvr52tSA3XeWzd29FIx+Qo6ErwmuAXpySzksrW7e6PqMEyx/lOs
vPQUz5sCJaHVGAtZ3014uMU9dsgzCjnMaFRw8BPk7vNHg/5M8zGtsT8PpzNs0Y3K5Vfz416lRa4m
ondSYf2dPxPFP/8c0ISxUEsgICu9+nHmWp5L4vVvFf4+Jzkp+c6JphDReTl4xd2oCb6OyDsQWJPZ
0TohkieLgCHDSQauDXYTeJ9NPws85z31pcknaSa5VtzzziHvmptP98eoz6m3IxUFy3wo33sMquzo
Sno8xMaPcMqCEq5Kk5TSUylvXga0Srisgo6Ufzts8zOiXTOQLv3F/WjV5wcZi5Z3Vlgv7onqQWGF
mbcwdFfmtjivfgHH9Aa/kdBzkhzNMBTLNfxAH0Idkn8P+DW+r81SG8N7cnPJxqlDrWqONvrOLg1c
8hLCjCjcwSSA7pLGIvWyHHPxaNK3rWEqYPni24YVIW7FSHA/ljdgVUOGseIoEQD3OAB12W+6EFfh
idiei9lrhR4Wq0jIGSvs683llQUI8wkSpSr7hNj3NfeUNrhJXUetmqLMCw3VlY/W3seZEb+56Fnp
EICq6XV8QhTHZQFIBB1Vxt778GqzBUymZ68WYBiCCMpxDiWACopkaFL3I5IBC77ArYcCnngxYLLr
vd6VHWLMD8wuHl9JWsY7r4u1JbaBqrK3bQbuoVoRvI+eaK0ORL1JUYN4XzUOenrzcSssnjX0VdHy
ipswY1s9yjzN+oHa6UOdQFuRx8+9MW9PI3uDMEeZeCyuC29BGfwETORCiAspzjj/0xvQ/Rdnq9mg
DdHhQZx7uhvxERMPv7Bgb7j8D7VASAcMnjgKuPRD7/hWiCgLvY/KpWrQdMmmcnk8QWyc/JqTZpQY
z9usnpjd210RQ7jw7EQ20GxiwUhv0PevmtddMS8hclnqK9/ZKTUfuPGrKSaz0y8USOC4/Cgp2YHr
EpEyj4H2tP7UCpUgdOHZR/E0qL3HCO0YaBEZdiUYgG2JTFSv6wpy7w8u0x6q2MACw+2ngkoAfnrd
e5CMo14PT3QD1t0cs4gihR3SRwDgr3ZCWcsPgbEoK1Tcj5u/2eBCnQsG5l/qlAi/YcJRh2Cnz4lI
VqhIExyKH7+5ykixdV03jUWmYRkV3/5U7nKqX/I+4Re4/OHIjZyl/xGs4qFhY0q0yhyIvYU+yE7U
TeZue7Wzv1BZVG8YSAdRKkHZqblDWgDyiog+EipT7307EA069SsDgSlEL77ajPZaua91sauF3Ey/
CgZb/pcJM6+30/wRhNPchYs+FgCBPih8/Yo3ORh63duIJZsX/VBtdfNK5mY18OLQ1nH/ke52TJwH
mRwavl6XKodH1hTu9K7HxCkSDbbwPtUYv2BbHGDvNAo3Du/ndGVLH2Sh3DACcJOXB3sS72Haaprl
8v2SDc9Q2QFR4hiieZw13bshN2+KFMgS0t7KUt/AiOzyBxugSFw233qSKRD0/KQASqVyrQYADHXN
psH3+69WosUVE682tKGD0W9lkoAAuC1VuoNja8dP58MPwaffk4U+Pyx+J/29LlmMoGe3QeMkAE5S
LxdesYvyOWKY5BGmTB0QY3cLNyAyra1Sz5wRwi7fpoVPMl3qb/ADC+ZB30slyqvOpiLuPb3zAlaa
nXxivlkqw6gp8BqvVWNTpi71PNmYJ32ppfqvPkxov+RVeD+VSGJh26k11FPiTcqkkOrakubuEU/G
Pkc9jrgcWHPawe2EYqFOjFgnEFxj1+urUvPM3/L+eF1pkIQVPWwoojkRn7GWw2Knuj4pk5Lu5KGV
H2H6QFR8dF49264f19QNPX5445GnMBZKA1KaPmL3DwNWuiIlmrV8NDBKKDRPfPRLVOj8JGB3jzhE
RSMN5mAK2nAODsLZhpph9/sUOc7MtUHMEotd8CUfXsgOLq/R5UeRG/88WhN4oNh8krujIsJuua7K
qxKT2aWvzVHZOPzmfnTGYt2abLrrJeM7AvAtGSMmM05VwioVTTTS5dec7UWXzz2mkDf9IsJGbQ4j
C9BJA4Eyv3pfqf6eN2plUt/weci34VbHysL21fOITtAUDoj62XPb3xyIbOBxjItabYdAMqN0fE0I
FSF9wil3t6+P8b7T9jVP0gIu59Td8YvLV/k59GBTdQGNvJTtEf7HgtAQDF4AMaBXhEkFD7f+gAnm
kWOEiOTDbebX2hn0UtgaoKPLmKHy8pBIY0athgxnjhBxCxrEnYT/HqVJnWIq7SsTKcvRa/yP50xV
cjDqwPytr9KzB4jBB+HmH3Vgqn5KxtDkOdsVCexyICbp3svnnNrs5MNNNbbWGUFHHYAF+iy8qYFh
FT/Z2aV/Wr4af9lEMPi+OubfM137VwuV5JKYRpqJ0hk4+WGlhrEJAKlsivsCQ695NfmkgHtzpj0w
hGs57s04JJYYorSbwdhBsy1sIUgYTGAsbxjWe5TNxqbK+T6g6qn/SFBIFSeamZXB3og2nqNe9ONk
MvTvquJdvp7AIoSBbFVSunPsAd2+86fp5RzOnwzHE+ggLTwmQ8I0FWatV+jMUj/nHfU+zTqUFqzU
Ipo5KkofBGgJIbX8UBETErH/undqXChEs5MVtFCk5+gF58RfPz+tJ/MMNDaOS6NqHv9a+Ttio4w+
HgEdg4EHNHKRx37ONdR9J6JffKTgD8lRE7oXbnS5JzJIDTOLWCQO7OIzQqq3uBe4/rx280WgZYHG
5EK4fCFMYcIQIIKZg6ztRWEganF/PTSD6diuWnCALIZQ5Ar2Y5+mRPIUd04JAJg1C9CsTuqMiXMf
gCuZ+jD987poZsqXseOMwKYFznnMQYnIn3LO/t5X6iKK3NOnXDfjlHS7jye4/NPqhp7UvxE8xno7
4uZiZwAIht6RjrlUyUsxOQQUYHtKOtVUV3zR4L4fPCsmG4xJVLJ+YXkSXsgdtXpWt2oUr7027Mji
9PluQyLPCpo/COKEJ1ZGwwoCpm2Wm3zzUE4t1xZ3YZTBf+ZywScqUu96HVyvMALio7vC7/2JKdKv
kEA+ET+FfLklKAapcvJBCdFvp1ael7baMOCX7ZzKkALNL7KITCupxX7oiR2lO8mDs94VPCJzH36V
Fnyloztlp4Np5POp8JPGZ7mAG+rh9zwYEyhJsPSjjZYEyb1FfCnCyRhsSz3GHc0TaMXwVI1exUlN
RSaD4rBwj3g609jlQjxoeCoVYpFUhSoDXrwFa+fri5C8uM9Us9SkmTTeKconUMjSEEnd6wGVumys
6b9kO7wyG4O65/K+mwg2FBPWXYyBop5X+KYOvqpJ+2dbiOGtsfXMEs4oFWscsBuH0m2YGUnxyhjB
iCpHY5D6YOZyipilARE6g/eyaFlTXKpzoqyWuBDmN+DqQXQ5xX7Trj53h8I+SCX/HjCiTxxX2HZh
Tkke4OfFNXaNt8kQfACFYBTwoQNyRd+uFiqp/jTNHcyKzf3gYBWTzsQJOPdM+ZybzG8tmjSgSeNO
zpmQ79vYYjjhW5R3BZHnfM4NW+25WZoJJ79dIU4s4sCqCFtJR95QiO6+/PcRuF+so9pWmfOJEf6H
waMzAs1Sme1Dg+PX2uwGQSMj0CnK2p4NIUUsmqbpDgaQY9AF8IIiMnOf8YO/BmEkm1g9RTAhrQP8
wbTn38lr1vrXPXrYBpKXuqc4VOB8Ub3OJXAnh+ZYxlaVTX4wuILz+r7a+U1SRtVGeGwqmnUrkFjq
QqYoU1GPh9Aqsgu5cc5SJgWZ2gPGSPBw4ZwQ7SB18dPLLollacVidQ2pND2IrdT7wQ8l1583BR2r
T+om1PjA8Sq7eQ31HeTtPLOFrN4W5y98nfne+rH2lHHq7ZQ2x3Ca80hnXcbk/s2t6yLu+4pvk8kW
tMh8hHX+Yd0Uo3CqA4yBGw83zHL2o3o54Tb3Y1hnUF6d3VRUx3Fp1kLg5bgXhbP3db7TRKXplA7k
3JBipLsSBm387XnOj2iXITft8CDUQIvmi+TTn5iqsQNPkXMu9l/kHax84gJQ+3QYRWybIPmIC+GR
NNBMpt5aC6SBMxqpsDOrPgaq9gP0hXsdvZaPayeWEz0KlTeOfxiUcxsQLjuVm3szRT0Htgdd967i
0v9XzPniLiOE++g0uSt+4J3hQLxIfe16Up6fbVnVjkNXAnydY0qRqhm4qH+xkIXnWWdDtGsOM1Oa
o015/+KrvGBF3VqiQPlPriNBARK7jtR0Pu0RX/PRHbkpVYUyandUCORQSaQxqNQ8oG/JmVKmwq4l
n9JncOisx8N+ZaTVyv00ImbETXZps+89zlisSR8pg8+yoNDcmtqwJ2Vz+k7qfArp5Z0rf8d447p6
e3i1iLEC2azf9i6N6aeGjert4zlWZMlJ8fWIx3PZ9QRN8HoUmkNLo8qOi/jDqVFMPuCsnPt3K1gC
0zwoZyyBFM4ySrhbR7i2S8eH7C952a2IzEEaNaKkrxVxb15Ei06aik2TDygTpLCrulskUOqW47E1
whGquvQCBHOEFO5iJWf6LWrICuoubtfyoaTuuX03I7T5HpACxaDYrqVGQ1OyUmsY8uqkY0Lz97bd
jBV9435WpWbJtH4z1S5Ayy2+mBWhVoyk3+MgNZ2hBGf3IPeDCAuTOImGX87oCP0D7SgqB2lbQNK6
duDZseqbw/Tktz3JUQNU7r7UmaQ2w4AhX2CVlfsQPcJvVkCvb5AQ1A5Gjpsuzr7VClPkht30OUCY
b3IJXN2itgAW47+KxitnY0VDPvvy6ZILdG/j3AsRkCkiZmo1GgfSYAbQbrwluZcJyy4uetfTO5+2
MyTuG2vhJ/n5VDW+TpzTfg0vuMbx0GFy8atjK+ja0g2IXpr7kUa51o7euUxdGm6MhqkeP7HHNsWb
W41E+YPCGgvb2QOFowrQ5lo8dJNq2xK5vcRPS2iBuqvz073hq0e32GrUePNpwYn4ON60bRwdIY9/
tM2zoBzoyGzT2Z6OOrHZp+eJG1P8f7zteDR+redfm+YpZypEElL2wpX4zZAjpjDUjDAdSn5KyK6y
ZZEYepLp06LvEPc1/JYZ5f4DJ2kgVKSuU3gs1phMB3pbi2hJkW8JtOpjZO7yzonNlSfMwPKSQ899
UO5tYiP6S+A/G2FPN45wMRseAPdSlKr4TvLvqLxsBHN2QoMif/dikWwH0Fn8XzGbIWAdfpx4jXT4
wHlJW/93U4FuBb4ikM4ZnwDG1OeLBNHCmwzxmor984+rkpbfeEGiw0WzBq0f5H07tXtJhjox9O7Q
7jl0kljbj0ZGRE9IpznF/pV4QDw+cD3h53gWU8EJV1jidDS1DOqk61j0ND1ulbWhf38mq95MO54R
Kz3eodG8ZLIlYv2iGIcvcbdzohljT3pfs8YG/EuDrXrwAs+kj/nEoXYV/NdYXgNSIRobjuz1wjjc
Fhal9mSh5dCigHl5Ja8/UZNl6F4Q6Rgks4T5nX2mRgBO7Htvt6kG8u6LKp3doG7Bu5JacVNPtTrH
ADViftnnM6CUD/ERH1xzYeHaZZQ4Pl6plrDN21YR1a54yTJ8LkDdOOsd6Q7o4ZC3k7lPEF5/Pa8D
M8WHM/YO5/GPIdOWsyhAeJiHAWjb9UPZtbsnqpyb6KnIn4Nhm7OVPaEJSX4r91QKpj5KOi+vM79o
WDahd9j2NtEQ2bc2HKU+EGBNPK1EvK4WnxsVdOeDanG/N+yceToxqpKbZAwv4cC1YWMu6C7AmO2c
RBrk+xVyuyukutJ1wlvJD96gGDPyHZXIovFlwgMpeGSCezFn6xZeAjXGVs/XsRcF9HWjrX4n/Yaz
xDltc/hpj0H4wYxxJXqCSmMk3Absh5Y1a1ujRno/kjJL0DkBGwyzvYh1OaP/5qdFIzihL4F3xohI
+UYRcKuAtc1Px09qSjYA4sLwk5ttnula5YIhrOFLXrF/6EbsrOVAFAbnpjTZNWMtMxxIh1Vqr95U
EsJaRKefN5/Um7q+MdairqAdN0F1yEehzWrQ4f9mvNHSY6+3mAoTPW0tcHGvoQ8KXgNcttG2OSzt
Ksk7fv4GMDBpGiWQiDvcm4SkYCPnCSbETitcoMJdyKuo3n+Ziq7W1anTS32VzsdJ2Yj0KQBeMIKT
qoGPtWKtCW0yAZdJN0OU/QbJeM5lZcEYUtG3go8fkvrxhnheY3nIUuIIpji06oBjW6opbR6t4ZsY
r8RyA0TMpZstVwntZAuAVTvNZiitF08A+rfJrlkM9BLtlfBfDh2GWhKN1n+5JEpXl24KvqI2uAWi
maFGGWU5mrurUIWbHHlcih4mL3k1oJnnLJkN/39zBPs150DjXQgE3xolRKscUzoa+z+Mz0J4aDWo
I4O5nCVVTT5xXMI9yZsnfP3GRFVSOJRPFimRxbk36XGyja8SzLQbVH/Bc00XKnW5CC6perUjlMYV
d3oAO1mSmURedSDz2zIVSU+dvDgvl7xaTn9wJ8Yh7Io58q/VNDdpFc1L9IOLQRaCV+VACO05Fc6e
0Qi5uIQjob+FiIDi9BG26nJkvnulIsNh8whquymj1FjB63xvCCNAfodNxCinU/cPpKymAxfNIX0r
x5dkux6YxYZPfb5x62S2qSi4Nl+OjF7CUcdInh/VzlhVHtHM3p+G+nsuUd9gANmmVtF3/fvcBO5a
1aFDIIuNUOrllpvj996T7pIBmJUlXKtL2Ut6AxmE5jeDTBghzhk8G34Uj40t99QcNqfp//xb9GGh
Q+zlaM09JUaMbHQTVKLDv26C4eIinCPYh4FBA5UI8fVYLvj+dV75EdVrDB3M2+atJHgUqlXmBg+A
A4+YRkfUVmFN8AqdynuSnOKXNk036u0ArPLKwANexRR6eshIZgbuBFvgqVWGZW3SfbCDW+ZWPppB
AlmngwqtUyLrUxor703HH43HrAfFHtGlkdYnNkEh/T+xRmIjdm63F/ZjqIjZv1q37RwYvL+Ky3ja
derx/GKKN5q59G3KpxCul0ygaAGK/OsVuIn0xZ8Ac6GsjJBZFmPRSLLyMVM34sqP0yRHm3MZErZN
OZcKtZne6JywjMA5Z0vEtifcB2EuO2uGMIgeq3xbkVJOF1dHEJAmIPr57lDXf2Xd3mMgdwLx5GN3
4yeETOWtaAIQGsuO+nm0DUV041r7m9IeCtQYa85LjulKoUhoLf4uIRcfMSJvfN/asNsHVAHsTcGg
rQhbrXf/LFy7aR3wJjDeNRZ7bd/tpVrO5KzAJKbL03wFPmmQL7iwGfivnzN9S9vSKrO47z7XFfAK
5wpYudzxEebiAZt6nQFdnpGV6AOtcWWXDVfJ8oBBeOu/Fz2wYZxylkuvruwrY5icug9c0JEPUesB
pknPmkSSZrQd6cwPdMMrVt9pF9EPH2B838Lq1tT0m8sH7l1CqguczdMgBdf1+rZFzRs/UDIaeNyE
XtOBvUUfq/iSjFWIsKbS/uqjWTpetrbYDt626ufh2OXdBSj8zQfX9ww9VCqaR9U0HMjav2QFbFoD
1OMoarH0uknPylFV/xN8fgOmdXYK6Uzf6iCvy9qQytyFu9c8n3Rolld+ZqVUTy6HsFCES9UI26jE
32pSZSQsg3wq/mjOU4T/cK9gs1WMbDYbfZo/Mavxwd2KYJu7vdRH+L9Jzi9WdbIEKTyjnWqVXp7H
G1k7IcHUDCCPBVLNBPUSDg704UkBgs04OnZfHOnmHIdcAtSJr8TodyNuXu4y/mdAfMgbQ3CigOnW
0cUU/xTIJaAhXeYNmBW6QEam852eQtsy0vbXLP4+nfoe2tDIzXTb7/PjSHgnVOIwIwRV1DgKM+2C
q1aeMsfmodU5chcjoa+NAy4LjOeNFejdHgIJiE7UMuUAZ0np0k2MYgO2bNe2aTKN/fOA2MfNiKWK
8hKcBjq1cSMbqCDw6bTmb0EmkT5dOvx4FwS9eo6Cjo2PhMA4IXbqbocNBeND0Ns8P6Q6JT7ZhppV
xoB1yeG1pXuya8Sd/L2Hf/TafZTH+Mn7hu/hdMHwQ4SLKvGptnKefPKubMJKI3ZkSePVlJ2j7v/+
+ZRY7fxPvl9NHVA+PPoi4wT4Hh/pEP4H9LDatprpRwyIoRSLlYvcWv23hN9t9RAglnmqTN+dsdQ7
7dJt8yqj5kEOecKflDwVe4qR1QUPyAjuUCvdV2Kvml828PLRq9tUHOYu/KHOPDIV3DU/I8st5v7o
IxPLhBRt3aZOZ1cZQgKAHsh2mc6k3p70bxGiWML0jlLgkzyVxQlxjcRU3CN6S25xmv8v1x5TV3Xx
Bh3BwIJtO/iy+B3lTsvA4XqoOB00fyOeKVMwGDht51r1Ys0z7YXidwzP/y0/xdRWNepGF8G/kUs6
etJ7IuJu49TFwpqrm7IagXNO0KPJb3VqFeGbDUnOY0OM7WMmVFFcCv8ir+ekzqbLXeTUiQHO797S
JBScB84YIL6uUqiK8p77uL4CBi3p19651bnI9HVGoX6UFnwY3J5IeTNOwIaOQVs1yYBDZq7uWlZO
wqL9AOEQhyBNfZ3rGAu6rLMY/FIswwyeFBMJ8IQ+Lhdl//LeC+DUvxegajUBVecpPLzwUZOXmf9o
8WcLUi2/pEA9sbMv6r4nUQapLG2BioN0hAGeelngdXjfLmte31/yEvjsylHQxGezTp8qoaGcUbcX
o1u+bxLSa8AaBEMrvLL0cbOT3/4Uj7h5QLfhYZk0gUrLhdbL4sNt6u8RlWxL5EPi1fvV5KtqJIB5
g8EJy+7P9OrBFJ2IqVMPLBW2v7CeR5WGc/DjhhJMCWsrJeV4P7gN8gI/o0gYRP9Fu9UNj5wSpQ3A
AKi7sNxu92naccS/tny2EPJXKl/cCWYbKG8iQ8s9XKK/8EKVkgN5gbrRA8ZXp+UQ0WcfK+spPnx6
NWT3NmL12qMkEYIeqpD+fivhXbOrTH0VbnZegYE63FaryDAKOUW5KRfQc/odRi32ZNkKC74ROvsK
XEGWIH5poflcRgCRHA4gwrqsLODsrPS49Iq+K23JmPcMPbK73icRsa6CP2U1br1AccenYSxwpiex
VUE9Dl9WGcd4k8sE/Ejls9jihUAZ788hccS1N8QcgaqTz+9xg0i+Q3KiIpC041rj20LPkkZITot/
LdB4Fbv3B7sF2cMtANKbUYQqWwuNW3I33vdK0sHHheFyFCs4An3bOsHJzn7KziowGDvlu//mFXRC
JG+a29eaPDSCJHlytCk7Ykbd7LryzIK73BAAkXMHCJnOrlHD10LbPd04JBMaCzOo/tECGROw9ulU
4kN9NvOFl1n3eUMNSoNdOCmwrvhKLx+YkWEiBC8couZJXiuksSNqh9wy+fliSprSvl/66BQW9aKF
QEE3DKOI/3KmOhA4sR5WUf9zILPvwKvrT8Jr1pSRhqxx93md1ngRzkVVWs00eFD3uDpOcxnCrwPD
eKhwgoCDi3mw/6+fruQ/bVvMgzDEnomL19U/iLWS1ohPUHSEFvhx/86pZQSKtOIsoMhWET8lYU7A
nR9t0nzuySnPxUcWSWIYMeH43ER6hBtwSud44W6CwtmAhvf+z6rDs/dp5Xm+yE+aa3gqj4HsZGpB
NYagJuyFJR1h2GMsXMMnKv0meUHN55O7uzJFnXogJxUCxgSedd1y3qYgAjP6Lt3poTTPIk98XKWh
l7NDpKznRYZ/h2i59/PKJLKbEXZ5BdvfWgyHm/RoPEORqx+cvHoymhiD4ySvFHr8z06TDIMghaIB
9a7qxo7USbE9K0t6stoQ8hyIgRI4ZIJijNfkIew10pMet+/4vPfT2NaUQZCdT5bY7Vgw1y/B+3EF
Bx52Vq4OD/pyqQZ84xhRC6RhnHLDN6EYu4JkuvNj5nscEaS0B6S9E3vFbgWsYsp17hsxxEOqai4S
q+g4et/27BylomKyKuiXoDd8MruZS+2xo/gJSx7lzIZRNfzci/4VB6VH7gKFn1rFAwUyS3eyDdp4
6EnrSokiALpMc+2s38v5tpYNETU/e1oNf3k38ObgWNy1XaLP1+EK9t5WfsT843o0E6SYytDB2kkV
ma96CwONrQaPiBRMmwjNDOsvUiHKA7mhNnUdr0kI7iyzn8LDb5OfwO3GnpDYYYCMozekwl7M68et
mqA15TGI9KtMD/0Zj0g+dmTqpTbzXEh1ovLIrLCU7rt374dh3DJKjoEOwKkFcW+wFvb78hPsKsT5
OcMu1cMGsYE9ZZfNUegT9w5rCBVRhvSRctFmaNJgOkkhEu3pwPg59MYbil2BKrruU2eSHHubjKQ1
S/6cYq0+OGhAwUeMhmculAfgGbuBN6NeLept5zgmp45otTr1h7cbWSOFezLIc3AYXzsuA1wUgN7j
7tnIq6FDsiVKbDOb63qCo1SR633kQa2bg40DYcefwtXjcMCmVkyp/hUieenlLgU2bprI8Of/SImV
GqNDSz/BgQ4bL/eQY5UeAE8HyHol5vAnasOxCE+wOJjlJjGkQSFFhuFQ7jXYB/6GwpKECCXWXNTZ
n5cqtyyRIOyFEuW690wdl5Cz8lHGFSHngoqWPNxyncUJrHG1LQv4deZsEmKjpELImRWHiTm+vUG1
zmMKmcVIbYJQtinq3rsGAu15e4sKHYFHyk27Ik2tuHrr9hDrWrbFBHVodvX48gREpGWXcunw7QCM
T+McrVhUTP+zkXODXcxBxVFvKkueiFaO1pUiwTmc4hzbiBgELrbG11M75sCbHw1Imvq1msh3nVj1
4QMIzOTKC3ePbrVGDse9TddllgUwg7cPZdvR0inx/8fAEEhaKMUrB4xlIl6/KEGZJBT/g62jrMpP
ujQdxaXuJVWonHfrN6Ig0rD0GIrWfpW+MLrDoZ80m3w+7JgISxk+f3Z1PntcAtLgBUE9StPh4onp
xQWUVtkUmuNFXdBxe/muL/+DnNDbi1aBrwSZL5O1mEROM7PrL3MuBPr55Zd/o+jD+BF49UK12VXv
Z8iDEjqaT6P0dQ2e/FyJW1BxjYBpQgHsOsJHkHNPLKqvSdlYwlGSW1SjdmOd6BbLuVO35SwpS7j9
AUjqcx2qe4pdUnV6BATxp2BvlYkJxRrSm0gYuMzmm/NckFRC2jKWZJ4da7MnRrCfxjWOFSyYdtP+
yV3JJirlOW8XOyr+Kjxu+fS/HvWQfQCfpe0NFiBa66vO/fNcnrmKP4JELwRwQyabODE7XqiKU4vY
Fy/KsPRGFiOVDkYaPVFXfJzLkLs3z6LIHXc8o7+vIFB2kp3HbwkeFp/KlW1iXbZPBa3SuoBxujaU
9oDDQ3Zyw5mt1srR1p/pPInfGxgpXxEv5DwnRpiXYFJW5kKtfBLKO7TKst199g5EMZe1bONcZucx
zXBEduPj3meTE2Wc2zlkoQyZ+sESHvFGHK6XNWMVG+Zhl7euagy9uThvNRgTFMZPxtIuXUnWtbUY
Hg3lw72ik44Bv4x+QAk2hKUggMdtUDEJknrkYNgR3Dj16DBjVgvQIWjDEft2L+ap++2Dy5wfE6aj
nf/m29DhxelaRyS5cpMWfcaI+nRZN8drbDLfahS1Pvn/aXB7180ojpXbleznRzePS4oHDcR6u2sF
jHd9SQasPqRGLK8dhb4+CAYWJPt2ltOFeYIyJi1J51HJPurv3OuHstnbIFgDODcvIq7O1tRk1tRW
tK/ESW7uGR6p7te5FvfbDJM7Mery/Ul258FpHC7un4J2nAxTeu1KTTOSFInStnpYq8pLQ3gLCvSX
/v/ssTU1lMGLiFfUqLTBmHF62fyZB30CfqMvN2cbJVrOJZfXI8Dnmowr8mTu8M+Ak32PEAzGgxks
wV3Rv1zy2xI1Fuljh4BUJQvJxyxQhfz8d3GJWc/YEU95myJSyPNhhfNvR+oggqSqIkEU0gXrLbj3
3N5iLH+WtvY0UW1878MwWZhDwogMFSfcj40hQ87mTjFjafGLxk2Zf0pPK1sc2LYzS7FU27H38Aft
D4zDRZHyFRVO0eK/Knd9uR1vrrbgqAwYUdWF64GzvNuQ5piBvtH5t9BcIdVuE7QBv76SK5kF0Hyj
iTpDAI7WQWt1JlmHRIIgiI3ycEd15RFQ8yXzUHIPNg3ElIgL+jKIldlCjMw9os3AxbEB5Q3KZ6mF
jgM/mWEl6d0rZrG+urGZttyiImTbhq0eILgU4/KTQWo9NHUvU8JCzndyO9h7Mb3jy9PDzjBYWwib
EMzDJQ4i2hykXsyGE8hqYUDquVNlhKRD9Fk1+YNPKkr+YnWzZsCpVGy+XofdN62LXVoDPb0bUot9
AJBhEhBCQ7Z/mb9LUuf2wJXuCTeecRHEsWEE0PEDITAx+yXqu0HQjRkZeE6S+DIWP0ghq9gjxJby
/FOu2ADmHPnOOgc128Y9f93Ve4P2M5YH3tFwfVr0gC1A0n6cbthDmxuMGdDUmEWqdkU8+JBPTCVC
10ZOcQ0eSLhP+FRMmeAmbTKliIW3UBdyIBVtaw1v1APaVrMXOtop8dXWKBjJFHoFbUNlhSz6C0ne
V8d9a1+usPeYlLG/VatN/MVJZgC3NFMaFMWMczRHPx/cqB7IQ4KBXheoDzG4JFBehrPj46zrHOuU
2QwymCPAfVWa9YxYjYeys6rxpG3q4IR/HJwd5M2QxM9Cp6/OColSAtGfK4EX6m+KMdRJL9s9E6hN
ZMlbUGYw/zvr0V8LXr61iN7fJtaDAE3oh0qV1XcneP82IAllODuNyZJWgkqGN5aylgoMRIaWVH4w
7QnxVT+m8od2QH9ylawGj8+K3BTAsWawrKtg4Hkmx1dBJP/dHh1NRPKoi9HYf4Kld3WEvU2TQTDh
fgU9IcktUFiJktVekShyuVgXB4KAI40kFZ1rbwJnxQcGGJkF5Yf9Gx5uv2ltTAJMAn/S081yd9hQ
DFSzW2nONJUAp+WB9x0dkIlrCwkTL5zr/NW2Z8TLLbAwrt7BZJsK3w3KfxY2bxMZQnn52XENOHz+
ourQtjP++euAHPw2FHKGD/5ey7O20S/gdP1G81MDjsqdInp82UP4WpVzfz+WnsR50EA3CwdEOu6P
U7HhseOl+egHueyZ9Rbu/WMzL5/gN6PVDzbXyBGgFX9/GxQFBLePl4WZbFsen5AtmhwbLRZr9E4s
mJMPFwvNFkXG53r2es0q6ajkaoopNQ/xLObTMafJH4hhOw2yEdtIqpSMB8+C4vtZepwSYv+GOYLN
BO+0x/FPdJePNh6c4SnLTy7NaU2+SOoy2JFN8RhBXVr/hV35Axtm3rW+vKUlH9b6cmZJupoTCP7n
8ySbm868QPiWSVbI4vzPoyFBl7eJo9y4s0MiVHZk8Tc1YnxpeLzqMjM7zDRNT38ZPl2mvGrTnOtJ
Uohy/30ly0/ZbmPa1eFSnR+Czh+uovOPiMUYhEP8ZbdIc3VHYmF6jBbntzBk7dD6X6eZ5tu++FdJ
MC92uedqo1vM4cWeB39+fptbhLZ+r2v96qaY2PLc7otWwoWJ6NsRNtckt4gzle9cgCBtonqsMTnH
Z9eM2r7qnaZGPZP6fS2uifEcZfMUDW1HuqOKhpZBe60Y/Lv93pMZhkdeBVZ4qh7hDUZ6PrQ4GOn2
xy6zy14r1+kcihp0ju+LtlRkfUxEVJXeILYGMYAG399fGGqXFI+SQ8383rEmAcWPCZ/M7xygwcjd
RphMXNn4lqROUTngK44V1QPJEeoUSEiBBPBEPvHE5NIJOG/5QCGtnkY0PELHfmWU3SaJ1mcwOwO1
dpec2e7iriiLO3y9B63KUasuORSouxM6yfTN6/tDb5DJGQ2G52V9iWo+FEAwGkWv2bGw7NkgPH7p
5fctH4MKievEnG3qD3Ygge6Cy1++ZaqHz49UNW/ClADZoHqTqlA6YBgLnyGLwNFPIlGjClB1whfC
BN0NK6kGOx3T9crOL7RewFOb1GrkDa8somEb0cgSe61y3MMZ1WZM8Jb1okbOfckVWju+BBkkcPPY
NHQGQ9SbWLX7d29vk/p7PxUmbUZgpGrjeKwxDEaV2115wi8S8K/bJs45OvZVzfDBC93l/MZnwnsI
kArKlUxiOOlkO6GZ1McaCu1EWC9RMhxu7f/WRvzF8pyFgmjJ8nJhT0d8d0BZiIHpeQfxxlpiWjHM
p946edgbmMdMM2rdqMfGVOwYY9Tjns9vUkYicPq7FRAVTxzPNvOK1AkdzWMP7wblrJNPl1t+1waM
48ARcoFx/H3B26iPYjUREJyisNAS395llROxnNMuKovy0he6EfbldxVTtjIjN5dQtQuZ5lGB8Mva
q/Fc7OKMKqcznvRkDt7ZmBK21bgaPPWs6KZ+Xeb2V0jq3EJPFBq01aWb4CIHiW1IIsTB1ZhPtrdq
DKL1J3fa8d2sEtPp98x0QoSflWmyx7l/j+eoakXD7spwE+f82k69kfFc4J/KNUAxbpncHXTDN+5V
NwN5PGYcyBYU4h69l9jGw5gQ6DtxksGJ+U2pCaCGie5eIBUYfqIrJY57Z7AtKC4bhYC9uSipiMMr
DiR9U813FgIUIU0Ms5pYI8HpLpfDCALMSq6QJnh6LYorDSVpnALqvf2rnX1AtN8kPcgmPooxOu3a
Ic/CeHiYXVGtFaRX2AFc3B4ph3A7IfQ5xDfCj+kkflrcaltaoySkmtSKOAAKOGKeP7oIqcW6uMRW
qqci/uareU1cVisCz+GvWT6808GT8MtGeOD7jfTXMy7ehREkC02W6kJtrAXm0bitkr581F3g1l6f
Ktim9wtT680Nn+/2xyVza02/yJujQyFMqDKRySF28/ZCvSKVPfffc89ug6s/jaxJpjSgd3l/2Aer
m0xun3AfTMF75XVL6flMwIMhyxq1mF1zhdJMcBpPfLPwv8mIxrrNvPk9AVdu1MvxZeJgZa+w/4al
BiH4xtQaKC2a/ba9L53NqYe03KTr6HOZVjD0qWIa6JOiBDvOVKncmnOpzmJOOxeJSrBv32oUj44o
ysV1Dw1QDJ1QO4KfYwbZazMQaKMDUAbV30CDt9OEmAGN5PrXjhLDvUY6WmpAEI/LByJd+9NTSG4j
oFAajdijPNEBhBAZUXneqxUVmdiOzzgDPcI7G/1MgL9BnhNRcj64dAA+1afsMpZsqVlWPHpfJsh1
FR7pbio3YAT9K28Q08RdE3YFdaELWO+4WTFpszxAHRihpnMMA7JS3/8D7t6nf4AKBQct2kX4JuNC
tkEw3eYgjonFmueOzq2jwmS37OlqpwgI6Bn5MkTixNDKT2WurDAMSuL7dhOnLaLOzoKk3JQw3wda
7QelVY80S5Par9y9K3vv8/e12Nh/28BBfmBPtf/XT4D8uxGNjRmGn6tBj2WomujE5QTJ3AAA3Rhb
UVxj9tIQO3CF02qfQzcbajf3v5ee0eGxRA5wWZzrt5X767fJMKMuYMKCFAzFHhqLVv7H0LI2hIwp
8tjYM3Rd4nWoiT2ovBbyCFlObf2C2lohV4/QJ+WRFTEAvgp/tUjpajkeG+KP3A7NAoXT65Fj4ynW
zz83HEPoWaDdYFPKbLrilYO15kVf4uqqgOm7DChfwAPZcQC2m57nt8oMrRUdr8/CLKvmxi0k1P6v
0ajtEVBTh4mSuSXWBDVgJ9Xc7lOyoybk8eSFjqjmeLRs7aVevxf3OvfMyR0CtHOx50FFH4ccH/i+
8rP0frScMvH8IOu4MzxLthAdyDR3dG4IgjjiyrpuSaDFqap+g/qvPT+8oXZyWNi96dEPGafUUGDr
qg89SBAHZ+8sbt/nVrTK2AwWf19UweCjHLI01oEBdUe7ZrCdgNnldsM+Hw2577DPytBfsME27d4f
NI06xTUlifUF5jRVQhG4WQxNdqDPjXxFQ8oAHpt4JN0YofL15w6vDcNaaAxc2qWIPWVJ/zyn6Es6
5U06itQmP3XrR0cjg8wObcUHr48UO5Qwo62ms30jHfVcjfgI2asI/+C0u9jEjNS2nPzEoeIqxljv
QyNCJ4Vykysyx5Uwyt6y4rVo/UMT8cbt6fpRmUhvXLcU+suTGFFVR6yCiKrFiDoKf+OW8TW9h7+Z
D4sWjRQ+ychYq3THedSZb5C6IVPE+m+eZ81qgJSajEp6AsGrOBnXNZW703fR7PdBic8ht4pTFpYV
wROthRejHC2u9IWmDndWLTi4WAyMjj/SWQfKw4kAOfWnkateUuA+EznUeADt5CWAPIHhZ8c0X0B8
TyhK9PVfNUIqMi9ir44U2hWsGtcZpBae3jzStyNyXWKw+5pho15DzDjvnwLv31YJPgyalSEVKvfs
pRMkWg8FGunaf/beI7tazgFAGRb3d/aTwu1K8izOu/7vZVQQAM00Ns7AMbRD7/Ej3kmQLkPZTYy+
rVXKZA4NpQf3YFV6HPi7PHP7uQx6huT6R9Qlvz0ABavRrRUJZUGms4WalmFjZ2WJmlBnuoPXrPz7
k6++lFmeWdbwGubX7sGS4jckILLm/QnI4B5IMQ0Jf7/WIrfBMOIbJLfoYjHILeF30Q/obP9x4ELT
zjsjAHsFE26Q27+JooD8EyRHW9FgT028ZRbkiHJCi5nO+xmakp0sof9i8UHujdfy78djjWnV+bKI
ZpH1cl1pCLvCDct0NIP7yvoj+pfiqrpBUCnyq70BSEf+3wCikx5nbnjh+dLMl9zNazRh3ouQ1/ri
mN1eqM/9MmPqNNXmqHwJdivF/scgM6hI9t6UhFNEMF+m4MzLKfgleP+oaDlHNVoQ2sRCEt9Dh/aQ
vOqdulqFzJZkBK54mG2t9aLmJUG3D4L/fRIOAQNu/uaHjwqPFWfT2PwBgkugySqU8Ppf7XoXnudH
3b1kmre4qzr+4fcYDs75pfAUqVB8cRxKXYF+7PZl8ebTT4TTbXjiAG9pvAWIxMcRc374r2oAaR3+
WdAzSY3Ff5vssx9TGBNo4rHm3/3dRzxxn4Tp6UXoz2QQFt4TZWfZoYzl7uAt8TIFXv86MQbDo+rQ
HcFGlBBhkaBi1kozcv7vzpPINx9yEWE5QGV+45ttyUp7DIMjGmKIvq/3qWGizTJmV1oS441svs3b
HZRrV/7qiawFeOcxngCb0jRIYC+KMtbzQdVXOc26jgGE0M6RXOAKexJ2mfR5ObsElLMc0HySivzF
XjmZcvV7PmRxvrG3waa7lF1Mm59R7Qq6ooRzs+WniO4LREEBlP/ljiflw6xc+bDHJb0G+TSCtI6A
1aDg264TV3wCcjffpOaHcsCnYAUAiJfjK8AwrmpB/UP+0d6TtSyh4YtIK035Z0JYAdeagjZS1nAb
CBQHN7Lv+jyFszng/HEwJsAsr+rrAsrIMECEUc11bwX7jxRAT0Rp2aSVfMJKCLqyT48TUuH3Ydkw
lEH8XspIXW4yPBy/MFiPio8saGV1DNw1JaZxrtvNBFG0hHgoa6cYD9q7OWgoABZbgwsZagIs0fd2
O88jZQKkxJ6hGi1Lzaa6ZlMjkQJuZBV0UxauCr4mh/AQEEqJ7tpKW9WcOJZSBLQFp1CDB3t10tdy
12lcI9jKhQpCNFLq+Skzn7sdJsfjYM8VTDs47btfeszqDVDKtjVH9kboKidEbkkfeCC21ukIpyxu
o0LBhGFHIFwXSt6DUzyqj+aMEEhUApj39aau6k+jbwsJGr/KIGmRb+ROSXIgTn3pNoCwBwpV1bfr
gG8IpmZxH/1u+tFeB8IwKPloXd8mL33A0cvIMKQbta50AitgQB2gfIiaFJOqGpMP48basUxTa9G0
in/d4rFadu2A9iVwW+JTGyGmnwcLaF30JjWx8OgPH8Ap1qHsGZ1QA70n22L1uO+EUjzFLo2ziksm
OkZPvRSEr8ht58dmRdg45VGMFpvRUX8ZzyhtI2vG1bXFxe3eX52aH2kF/rmYIZsHXRth1xo6e7HP
zq1poh5ORUeKQjteZsCpUpb7iVOT8KQsNiWmL4TjNSHSLgtUXdewv8pOtUWIopXgJ1hCylaBjV5n
5x6MjhAwki+LnuzTNyyT/HBe+xfdnDVBHb4SNKIDlGwkZUUGDIcCJt3anPa/LWZcdZGqYWZ+o+wB
3bipz/iepWoMZBVfiKOTqpu6HgdxPLLMTk8x8Qh5En/f/u6nAq1rnBR5ZblBib/PCPi1a2pnC0vH
wyONPinxFhozOaaj4F+MQLTA76h9+dn/cg2tRl2D3C6uJ6mMRbRQsadII/CicB8sXDjo2kkyu75z
4BYw9M66VO1tCBUjrWbISB6WqUSEP+Hp4kIOXcReMZDpYVKbLmcmENLIZoDJUMQDjQFwAg8d85jx
mnZwQ6lq+51s0b71Ji5N3Ken5CSdeRgFIhSaU/RvUCEOLGg6HI/gutx5ItyDfmmYWSNCi6YxoGDt
EYEKTevY4bU5rbhBApaYnbDrl8Z8IiTvrcJXoCQAd8Xl0Tv+uSAPzEug2zq/tlDjBWQ/GnRntnvc
KkM4ffGZUUarMK+kE2Nhf7uYPtHiRzPkZV2DevP/VCh6wC+Z37d/2bFPpa9Fan+jIR/Z82T1bIc3
w36eapeJDpDxQ7kLlYZbNapnxIlWs4lizmHXYcMH0UBWR4yP9bqQRow7sd8IoOFVqICXl1QxDve1
25P+Tl8S/RDkJ6FsjPJt3z2M0+KAE0Al9YAKXISepZtowGxWLVVOnPDC/MUVGikMrY1Zo8kb69lg
CWL4yItXlcaNPQ6OKTvE5Omnrg6pd6LJwlypTvjwZh0N18BpPDy6DRVfdRW8IErmQx6fROMG/0U9
LvdSNkIVVgPzbiXM2wEICOik+gYgCWpYZnVovOJYGEqeEjrbbYibGUbztu0bUT6SlngPz23pZhDY
g4q1Z8gt3lAwbv0tAS5aUhvt/zC1p5jEGK+tzEKooEVIbgAC71642pFeOd5fRfJnur3vGzzWDSSk
cu/Zk+SrOamR8WPrENPx0KZ9ccY7TBKT1jzNqA/iTqVk58xiUx220jNGD78Pyks4PXZE3i5s1GQI
+EMBSOw6xor7DpbbDsYbrdcJul+p3RrlKqDM35TRkgsHpkhJtpWpLoKeNC4K/3/OnpcFMAsnRFOc
ldImh5y+kjYhZqyBy8saOBDF5swjC4pmKlNebRFp6Dcg43v6L9WuwrfCAqRU2bGrAwtSkOwRxEWG
q0MGABUW9ADpvo9DpXlo1TQUjYLClzSuGlcPMljjOyJJ9PVwB8RW+LSfp02GAw4zJmNY2pAIbcPa
MTSTmZzMooUmuecSBHfcwcVg4bfLmSZCbWhLaIhdqjtJDTn5ERvLjvDn9XqC7nPcOYTf7BjsBnVb
x5Iig2ClYOyCnumbtgDO9/kH2iNslYOBD8VvwfNnUWncyJcla8ndtu4Qanzjl8bn1wUmTTLKxd0H
vCWuX1Tcl2DPVfYlM+Ay6Gh/H7gVRoCdySI0T9PL2h6U+pR5E7SjYudlUPnD1GwxMlGMHia7ANGp
efxXjnwrQ+hohXaq40vpG7JC3HJMEKxj6lsvixpwifCrNc5sRn+JJABbAYc0EtlNV/oYvancNsa8
1n9JP8PR36Kl8HvOuShLoxrXvgWgiR1Ar/X5CAAbG/PI9K5sBtbK5mGprpxzgeN7zOo0+pm7FH7w
IcHaRPSNE9/v1Bxal2/+X+trKnez1fYvGB+7XByFU4XWIo21aQ8AhyEHr6SGzD/ohK6euKMvO/fz
X7Fj44W6bY4a68XsCUhMYP62I9OXCRTXZHB0cGRjPNYQKPwsq0igheHJT17s6kFbk7602R1NQ0Bs
DazWZD/YYLYriCBASab072f77b9S5JaIrMQ1uDaHJ8M9/+AWuQTcKA0nsUl7DVhjTiFwCFRhQTCU
3XHlHRY4DugUUfAF6fisZ5C4bPEZSQFOH4MpD8uKWaX2y9lYJZnbG3tXnd9kiQyZb89wvBEAYvh2
5LLxsCvKjKXrk/wyOTqWeDCKJFE1R/ugbqBxUJn6xcZmH3kG8W2ZyzMkuCGtrCfCXhV8nx/VsEdg
40si7vWfTcIZJRkhsl3yJ0+tUdy5qwF4BGUhX6vwZCm5G9BzAEK7MzyAAIzkhDxvqNPh5/RuiYod
C/1VvyXGo4WUc8OA3YcAdyL3pqFnGML0vZx+zwqX1/o08iSqDV/nSK6AY0bDKM3HudSgO5ptNujg
TsyYrsbijanLpn9A9/95LzUXko6MH5JqOxjOVHy6hnd/KSnm6aLEvPAJSfw/U6SBAt/Z8/LXi2cY
Rey5ThU6oYEE3/pubVFax+qbH4AN3Uz1uSqQdhWngLIP0HtwXv45JJuMAVdfaHAaknyQWk8s2u5c
pSH618P21NOE3aALMNC7eyx6AYDYvhmpvpX5ey4iEx9z3kaAju3FoNrZBos6wxaDobKasGfDvCIN
Yw2CfTswzOrQDqCjX/PpAxpqRHMMDBwZO69ausgjzQDPvmGhOow/rj9ooXveWvjgdPMPBjyiR3Nn
JRXg+dpE6EbLF+M/MsxYEKEC2cSAOADvc26a9VTwDYVVz+Y/XgkIei2PLLD84fJmohYcjK6Gw8hj
v6BcyLOfhLJyirK3ofjW64e3xZFpBLJaFKtlh5mvEfdFW/pg5dZzW2oLrfC5XtZ/eINh+7fjLwiO
0UxsZrmDsfSZrW+jtgADKTMec9bfFLz7j23buKc+YE5JbRz7CrEyqaLu6qP4S23JoUVT3UXjWEfh
dGCkJRq1RZkFJEpvaodqFD1c26MuknD125Jmvayg6owsLcUuBBDkUickqlaRc5KxWb/XjwcSdHRR
gQRmZ+dS2bMeV4B+U03vsT5oiA9+rffvK8czV+VPpXva4qesx64S9nVKTpHHSJJPvpTz7h9nTMh1
XKroDiygRtYI4a4CTRKOR3TSUrJO6GSpY1Y90YmF77ezRRNgWwkbos0nvYOe8k0zhJp4n9Iekq8p
IzWjHRXOVg0G+phf/Xdg+BDJkMZ9nwHk1dKw7Pc5xS7aXu1RXJl3ScwY/gqFOiwI7fDgzHPA+oHj
+9LMFTfTSVGyQhE0eJ74Xc0V/bF/VNqJCHGpm3R4s7M9HCP+4QJI5V0d4r3QJAH3hoxuiQnJ8wLD
9fCK20lXM9U2/BkLFVdg/rMtxYjUIgYrIGxbA6yL0oyTL+AL8TKqEZhVPdnLKryGTOLp+1rN9xN6
YMcVL1GiFN+KbUJ0Xi1iPvknwV9OkLK/g11ZBzinvduh02yWr6P3GpTM2a9tn7eOplDwhjUnW4sp
eIxYgQM3iUaELVgyC+9TdSTujXtTGVOBqDgsEhmjy0Mop4H66emk06r8QaZPNY3MZAgeeSb+EGwG
CFzx3Fz+0y1qw+hMs1QvzPoHXrb4bgLp0zSS6SEu4aFq21rMn/94pK9k12l642L1LjwjiHJXO46B
1jZ/ce8v5iL4yWgYho+eaaLmCzdB6f7ra5WNtVcDUTSZf1oGGKLgCO5V/v9atKTDANn8A+6BqlKQ
Q8XieD/yi0qeQ171UwedRyI/q3abMDIsRbtRwn+1mx6LD17umdI9fCkwMRdj2XcoLdTyXve7+GMC
ukzPkVELP4sNS+K3pUtMHaj84468RRHvx2B4Ttpmt73PTAZ77M5CjyTXfMEHiARsf44mC+P8YrG3
adJfxm3c6vZwfy7xqTuYHVEosE5vAlofNkAUYXVkqOEtXqvZZ1kPRaqMCo6h+oaRdE3WbG27dEuX
Mj3nSrEThFUwmQO6izXoc+/wvb06famUn8nuIlwBaDSYU5vmMyoeOGf7ColJe8DoULKhRWAWYfhG
87KRHHc3kzzFlQraVRvYBjEn4GLxVQ/68PkNB/obu/pVeATTStJQtUMVR5cJHcEXPPRXbO6z5v3q
AquWlxPmh7lu2KjAsbF6KTtDJGfzQarUY2uRU+KxYZIkG3qLFhGQNbOgQqDDhFHD3990y5frr30M
dr2RhCzGU4KGqSmspp9NI9y23gDFck3WG0BwMu++T5T7NfNiVZCTdt/3cnwcfHhMDNS2V1I2cmdV
g5o45/f/Tx/593E5cq+bwOF/uvgJbibKB1Ftn75d8kTc07QT2AV2+HZnD89+vcRLlU0bSIwNivBV
+J3CQIBglXeZZDJN0QvAlZnJEz+UciQTqm5kxODOR/ic0nPoZB5kRMK3OOhCka1f3vKdKKnLbYUg
6ntMV68im+ZULfktpAXfa9rhhwPbPimm78+N3lltW4efwSd3f0EU0k7Y09DDHx6rkWLyZA5o0dhD
Lh+eTJ+/psPIRcKZTlF1tpUqsWZAT9JtZChDrj4iS9pTBBSn+pvTaVABDWlkLU/uTiPIYHmbFphW
OJo+lUj0VYwhe5RmkE22qJMrjVyRtjRqXWZ8vv/tB+sJedR+dfPnxt/yExNn4b9+KIgcW+Xo8ntB
RWDqIgAEFeLaha3rcEeZLQi9Yyf0FpZCZa0J2bUUavHG3H7wUZDCSDPTmE5MNek5nOGWnP+WOMqT
3KRUmcEQh5iyujtkYg5Jn/oEfOUE1ViHleLS5DE84yVrb8mpGBptCCBuFgpAFKzDM4q4HTcCblJI
arAj6fBl2ida1ABWPVshx6XMBuDToK9YzyjL3WYFxOLqGybrxZ3daDCr937o54JpnScgLCe9RDwh
FSp8Bwl5qkRrn/OcFmuQXINcZ0c7c/797A/XNb2S6EejedXotMjbvjY0t6LDtETy7FfgwgBV2pl9
qvhYHXOKn/e7xFroxP0147iu/QO2gNb9x9mmbQrOtjn/69bUeJbzmBsfaZOA1HmVyQfeiuEmj2SO
zM23MNIVUuQp7oNEyLrY030frqA232W0BOOR1Y7rV9JfOg+S02i1JadtLVFn9eyllGrw4HYJWNwW
GJKhdbDNVigY2Omz76kLiKTgkxWWMxW8Uy8WsqtNk/j2aQ91qo0X5XFihNATWkH3y8DHcvo2yaUO
4RbcNRhtMqnDagwpv867RoKQUzPSc5DSDU20Ta5FmRvF3FKGt6/cBv7Uy9if0bf3QLSqcS+NeIbi
0uYKHTqRB+RlXQisAjGjMryNxGRYwZlK1Lr0zgG+oAxW45yPCffnWymasm00L25fSM41R7XXb+eL
ibdEm7Oyc02icHzIIRmcmbOEXTQW/ugeXvheSb5RBT+5b26jziY2jHftAgGe9Jr+xUlbkNkPDzKI
O+jTuon5qy2AtoIt2F0UExEjcLPcOtQpedcFL53WHx6I5oeFC7PKc6PCO2Y5Yv95Y4sG8omOIbpE
BrtJMhgtd/r2R8WBaTPa/iV+3tlcmEa/w3pQZoUbt5zUPwF8JDvXb/UGSZe4i9sMAgAWD5sij+Lz
G46u4jWH5A3ett2beVF9kp6EXuqAU6ovhqeQYxexNOrbrYgfTn9dLSJB/qLgILLdUdb67ThhkBCq
Dd2G9dzStC2J52q5IyH27k6L0QlErsiBuugjqz4iKqCoqQlZIO2kJ9aoqvrNGv6P4S9JbKF/A33s
QD1bvqsL2WWovJELfUf0uaUgRflLC0RJXEUfR/tcH0jB4BywiJUjB/p8x8b6oV1pSlKtLLptsGJ6
MyJclKgWk8FfGGlvvNdNhP4rse6JR0nrv8QVMNIGJRLFvb+Pi/W+grbIhZYtlES3yaBW4btrnvFq
e4dc2yET0xl91b7D6AGcmMEagt78pzaaple84SS9obAJc0nXOjrYkUWYpiWYrcfwGoCKL8aU4VJ3
/eBnnawj4wK4h8UQJ5mlE1iuaiaWN3/H/js8vQvr1vspTxUDwhvuXL9cADkhOtUFHAfrt7X6xp5W
/JUEFbkZcPUprPoFoe6zwo1MoNbfB2+JJjRJ8A2AO8AZ7LgJIg5PjhrenWtt/bgr3DJ3xmlC1HbX
B2E2w5D6uw/VyBNsj0U02SnkoY1s8Od/CXaoHRaF5UCl/p84ixczgSBVc0fWMMB0n75F62E3m1ig
6ySVcw2BgjgJowOL3RZEGB5LX3T8L4rYv80qh3e3SOmn/PH++5CNdkU9zXCo+YklrcYRuiQsbxea
rh45xZCTxPiL94JHmqC0j8fy5jn53voAaDlM1h3/niy106GtDktZrzx2aiRV1Q0TvSd2rgnSlDAD
bhgkJ2ZxDJDpcpzkBkOXCfdcQQEYOT91nLXsMsF34rOygOoKaadfWujEEjY36RP5CneR6NRVU/Fj
HS4U/fyVpU5NOdxks3LBZtTxumOHEht8kiPUN0dFj9eNZo1oF1SEmczega2vmIFymhDJkHpQ5prU
biV7jhMz7cT9e0jkh4uCjBSr2065uaOXS+YrOgnyyIB3TO4vzTQ2ir5c9e/TIfnez+KaPx77X4f8
6QTW8aWdS7CtXvYxW44Doj6djMgtfSrtkpPNEFjGS9eYf1/vHnYFVYFsg9KvuVeLoX4XdQsvJGeI
2XagAqaXStcpXhI6bwe1Xapkw3TOIttTa6zRjgcKEA2oZN2k34jbu37109M20+jPnMbwCOU7cpNb
E/5tZG4KMzQCaeXbHri8nW2N8rFMMfG2sthx5DYxbe0y0kLYMtutztwG3oTJfV5Gu/sO5+zu3r2H
rt/bjuRh3o/BMztlTQf6hWAxKJo23tiS/dNzR3Ww4tMQUvzO24a6eyXc0A1AqMCMAZVevMNfC2Gg
OgpLiLoxqd7cDkzJIqYZB0sDAHO+8NnTMcf+ppM/AjD+uzUd2EEuDmquE3Q90yfMAc7WlG1xx+7m
gwMaA0Yz9KAflQeDvwDhH9+5etcyp/PDrtr2cLn92KW9TmhsKDsiwb40XoWcg3q0GpX2BmGyhNYn
rEYIa2q8CDkt4fZk1DwmO2Fa4+JnxbiJnZ87SbDK7gG4aK+8B8JQ83EHK0+5hGyDAdLGxqrD/ogi
q5msmw4Reawg72JVZahW7qR+ZD2u4FPFiSO8ZGdpgW3EH6S07/94mszVm5J6mgJrTuuOfD7YP47h
NrCeQtoqLYK34RNvR1U+eVrFDXOSeVtf/7mi2eC8ZoRQ7FX2Qpih9mvbIOhYP0lAFbAaIB3E5paR
7kZUjFEKdFTt80d12FpHXVn7VzrH8tK5C8Zf4p8vQuQrQBOGJKDKwLM5m8Fc9TUkOxNWxhR4qUuX
SCryqF0pTwu2aGXrIZZy7v9nQhrPH3ZDglJz8j8G9lbxt+0Cu0Kg266eZN5WWMFfJChnqfIjjt9E
/ZHHYtzTX6mFEyaYENstd6cE6iDvpspUMqDY1W5BOKLU6UH7xwBFIcjedrCfmGgfSDCWFMDm84Q0
xqHkIhKQzySvNCZFlSn4qQ4IhavhLD/yrpYJhS9hUL3wUtts7Ou7dUcoIpICm3tjJ3Wy/Z4k51lz
Q5W7d99ydUC1ktEsmneQtafr4IDV8aA60YKxFBhFHSql6tRoP5YXxO07iPn94GnPvby+EKHV0qrX
N23vS3Eyz80kwd3GGHsl5nNCgDDhrrnYYKmGwOI7mPAtI7/5NC6AmMiLTr23ugLnapzmLmVM752M
xlQ/12L3p12PH4VeDi5VGS+H/qYXxxt6AY8DFI8lTFENNS94pj6u6uplXMRuWW9QIw5lkAHyAsHV
ssJFxFKdct1huCG4XkMTfwXwxgUPJKC4IXD/HCkfpNYhxqZGhYn4j5Neu8MY1BlarbaGl34bzRGr
cqTIJAb8MKot4IRnPwdJe8sbpTh7FIbRafibQbu6vHVJM9fxOBOf9PMgyIKq7RwACeBrng1y1JJz
5oGwWOc58H1g2UUCv3UuKtWwg8m8gTMxw+j4+wAZfjuT80ba9j1ja10bUhYZdNM+9K47aPUxxxMM
a8ohtO5mnLzjTQ+A0YVl3gCTAdG8X2to1nhAIbaj8TzNDQ5xtJGtcF8Y0l4KRUCAMkaDM0uXCPKA
eUjTwP4UbuU2tK7MrENObe/iVYk1+UYXv6MAMVxjUdul2PJdR7Wg/Lq2fjXTMaaqgyacB8EZJA4n
VEXDqI/vR4GVL94XMLKhFYQfW9ii38S2lTH0xIt3qpRb+2+fkHIsx+ZwZxjWL+DRl1xcRTkDBEmy
tERvdT8djvY3mDxXNAErsTl8HeDi+SZCVNZ2Jb2gsDXnMibWrYlsy9jPL9P1HOlcaY3fYh1eHvDG
6mbQht8MiXqGtqrOMDLbLQ6NbSiYEj1aPIXUqzLC98Jj79uzu1isQHuBE/Disw/W5zwFzoxw2uaB
t8LY/8dUIcmKHAGXepWyWl6wIvAywrqBuM98oLGvJ/AYaO7ty3jktdnz7NDIWf8HcZaV5CIKy5Vm
ndoOQmxWqN6rse+ukFANe18/kj0sCc9AHwVd0veE4LFaWntwkJecmZ9pnlDbpznZxkHyz3FUlOTd
wfQ69shRCmoeoZnjhGk7x85Eyn/A3DMK3vDAd2lmINdPkOaQli9shiz1HMIGW8l3XlHEpY0G5+1V
jUCvAnbpBsECpp00G1ykcYQr4eOlpejwsSGdgiqcQExkE3PQ/ftC+kNmIUdRn/1iV6N4f0N2q2pj
4DXP0Xs7fucMfxYoJSxnEtb4A1B7Fcmi1SBWc2V2wFfyLMb3gpKU3YyTWoVws77Kbqfdd5tlxBxW
spQByrYXGMlYzizl2CF9DO4QDAXm8/wbiiEooNJmo5M+8JgtkKo0LWYcEx22LGtu3vNSmFiWCUjJ
jXq3XV6y7d0pIg5kwW4f3o1BRhfaBRYnjQa7ItjDosFj2sX0gXWiJ1kFp2kewlLcCYn6TngDDOgx
rOpr5PBoWxk0Zxwk2FaF2+eVzubgF4TvaTp8mS8cZDJmJ5sDRtrr4sITSdtAHij0qcBLTLVitAKl
+xfn+Rl/k2fBBRbS44DJpP77Oc1jw9eCXCOUIrSiE/dEHzNxJJPDWWZHiPsuTVh8BP+8TccUlRRq
0PUK/GjOkne18tdV6H7sBdgMz6s0ENrNMj+krLdAvOyzIIRTueFdsikSZ2WE4YzJ1desCcdoBfgw
FjsaSXJHsT9I1iDBSPeQuK6IyBF/N6IrcNNf0h7E8h0KqldOiU9GRhHOieHPYY7W/9XQfeaCyiBJ
t01CrMEFJOM3SVejKx/nz//UTkB9uA3ZVcCajmQn0LaxHwqkNQ/SrwkSeZX217KKcIxCTb7XcTnY
T7y6LOCWrLFEt8lrPoGyxYxvOy8hhU4ryeVXJ54aw8a6lHHfPvphQSCVhlItX4/486bVssI4SEcd
WeBOCMKLsoRpU3zREqN9Vt+hHZOh52cDz3/NmcJKpmjoi1FaZDyrnbWv8aknHCSN2RxmN12zOELV
c71sNhxdyuiGvx7D9L7H4GA8KHrtvNovkNpi0z3GmppPb7nN7WCw9N0PjMq4KoUiBIVekoOK7h/i
G3IvGP514JI2wHE5e0mNsqM+DNCj6WK2G7Ax/2V4XL6Vs4OzOXG4GBrij4kUuy/YOi/tTtPOcxPF
+GpPnQAhGkPK1z7vc/RX4hOdyvarEe7+pMN5mI8IQcbhzQhEbSbg+TYI1QIncHudLCmzoHkqciSk
LOit//jEr44jzoda3YsPWPVzW3Ey5EmT5+GuWtGBIfJO5jPbmVSunVz7VxVZ4SdnSVy2VBk6bDAb
ZfB6VI+Dp5+JglMex67QmPz+xcktZBwlj5eyjUe4d2ENZkiCuXnkRC0AapZI96CoihSvCABXFQSB
aIuxGbisvUXlVhcK87DUBTiWmHi1CA1sG+AZbYtyOfx6OPl09H2QShbAAw/Ec70mxFJRd9eX/TX2
RNx622LnTHVkYbr9gVkEL1GoqK0g7GRKyEqE5EZoWbe+4kN3HFFCANR2tQA2Jo80fZB+GpiZrztz
5GYKWy+IjPE/QwTns7RpmDc+H9U8pimuWIRw5lw2AxcdIVnsHVrtXgy0Wi2jRJCGEt9rNVXdpr8i
kCGJ5qcbupljZJISuZHEGH7baHQz6g4iZi+nXkZpQNq/FUWSgbx71y3w8nw/EhPzR7MzTtUYWQNv
AXkq6WRdbHiOvD62t7dFMHiDuW5aRRzcJUfdD14gYheNVusO8BBXA/RPMz8CCtsEm3WlsGrARnqr
LSDTwqArzeDogK+0322aAfF/BfvUMzO7yttQa/ATg+Ww+8Fx389vnszO2qwFeyYs+lZPW4t84fIr
kdLZQKoZLeL4cmPvDO38NnaNrqvmw8ZjTEaWlwUDCcDPAvj235knPkgbc6TyPoKRT2tIht66pGrt
5geXRJy3JGwF9P7lCNYty3uqUw9G5O2XvUBgYZg0C88EofpmVRpN1j4UgG2qT3GsEwh6+DD2+F6/
A1prkWe5NwnwXm5+9li3xDqj9qCdvw1mc7kNoZWcJXxNq04Tsu36cKuIBzQ76AYt1sBXTPG6HlIx
sJ4cq6F302wRxruznUPLu/GVfoVoqWf2PESfUnIy11EOGCmkEGyeVgPRfQ69b20s84hboXPVn3Wp
BYvU5tYkx87JZEt+GEdJRfRl5wqxap1EA8EMP4iZr0pNoFHB3MxDVgM8HE3vBOICAdhOR1Xzqmq/
OfSkbCJElqpYQut6j5Abspf1EvuCwHEbsFvS+Eio3ndAPYjvbo9LzBDfth9i+TMyXmBCjxuKkQMQ
X0hARfSsF/t89P8FEAA7pGDeTyYBxaul9AOlQ/8yfS5p8fVS8Ce/G6pf7aNcxU784jUMTHXRpil+
uAdz2NH4SRQPEZQxwvPewA/CaE7f6sm77pUo8oyzbNtfUYT08U4mPInB0u3dxCmf/fq62gImt6CN
JLb/LB60Ppgy8b2hllFd8WOMVtVFHDpYztpJ6s/O34gmwlMpishVtVBL3U+oBctwIP3zdjSf2YiQ
mNE47JodJ73O7+f+Ut+q7yUhIeQfa8aac5gvGoZvMFyInd7QeZbWPXx4AdW18oXqVAG9ruN/Aobk
I2jU/JlY0hGUJi19bS6Tl/ZYHNvUsYEm1G0cyIeZfZPEcLjJAFRu9ovOrKBVam8njpxwN5gKhjV0
75NzpI5WqisY36ByIU8WSeM+VyOhcItDXcjRnSklhChNxK8hXsWXFNg8aT1zPumlT1U9dVsZSMzq
ik4PdGZbDH9Dzw8+wUJvD0I4JcvqibI8ovftMJkLiIIvJlpAWp2Sx/PogA7/ZJzcXC2P04nPzYME
4SOzRHf+NfRJm0Mi2KT8xEPdKag/A+gqPXzuw3pq9FbAInDLvl4XZpmpANVA665rHX6mUEHD5fnY
kWGssT0SnP++f/phjRidvePs1LupzulRkmMLpzOd0cdR1us+px2xErqs4c9/Cr+ufmRLp8XR9a7X
R9OYi6/J/x3rFinQ1SnswxWwsNwppkV5eCxoHH8YeT9/g3LQFrbGsCM8HmUm9CDR6vd7G1eQBzgP
C0wzkXEhvjzCFyMGWH3n4vCiKEOUtKvSWNCCn+5cgUaxo654UzUwOhFSGms5vTz9JanU4ihtciaW
nwSGyI3kPnXqQhQJvmhXC6fS5/GwjBNy0h2mF+S4Pn2GvybIvPAi1nQrikJYtPGbxtZtUvsOl4lP
/bsDZIfBrNaq5IHyLyyDLAKSomFoGHq0hNhhDHtdpQQuw18HDHAz2PVaROYYhu8e5ySmJ+o08G2c
5sM1X/uP1m1YrR/RNCs+yXPOntBUI/vrrJZI0xXn6jUmUov2oE5DZhe7FWgnFhWiie4AQk/NLjew
1Wkd9AUqBEa3WuqdTXIlXqU2N8nx6v458Zw6MQPx7Swag7K2qQvcZTM6QjS76S0rA46maEyEzxeW
3zM+dhkW/n1t6tAPXNYbdILiOm4IjlEGukv7uXbyoBjPnObcRLXhA9szh20J4BsmXn3ySoGrTB4g
Bx8+OnCOhWI9UaUbnvIZd1LCNd/TFZT9JGPwVnVc+emmZ+/VZGhZnJZkzIB8qPTbUCKsmyOIw31G
VyMLQIWyOwxqs4HVuSwWhJ6Cvk9grYX29MVhMi+YzqIJU88+v3gRH+E61TEo3gek7WPF/C/qeMcw
7X2voaOutuGEzekdJKVboFACxSgyV0kwI8LXD3+9LrASbygw/OYGn5gyaYZ0yO4mSIvpXtKskQsH
Yc8F+nZOZ0nuwa2jemhl/Dxa3orBNm4ujo2e01CHs9Pt3RU0zVdt4mch/d1yGTVzOIg1thQdpuXA
NnCxYxyOfHDYT9Bz+5JZHPqG8Ob8+5BCkjOMH9tbFvMmDXYV1Y4fF5rKBuC1rDRAVVIObHRVZlnL
ISz69o+ae1rXC6gYAhULg5SLWv1m6LiHCeT+dcvqFM6fHn9C0BhdfV1d/ARdJ7Ys25nsNw9QZMUw
SE/2VBiqg7X5M0uPtnzDSS5yNVtq9dJVwPieG1DXVyyQSW66wCtPfqzoNOKMZ5h7mTKB51asnwYK
Tt+mgeT/3Masx+ikNfCqBHElWANV3E/PN7McOoiU2QOyoW3nKLN7ef9gQX0UnK/Lqq78Ctjk8nC1
B90naXb+AbjVwJPdXSKH9PRITAuxFqYPGHbaPZHvvgaPQh5efxZojpqVc1tFNHl/x/KNF0ccoI3O
WHbTljjWfhbO+4WQrQZnTgFeS/PijJ+xCN1U1KuvJaeXXqV6wKawMRD4kGzz0mTSUHpDWC64ZWO0
/lSI/0SWO4q4s1k4N2Vt7XrdOU9ZDskAF9YFM6FvU5J42YRa1+hAQe/dfx4LMUvk3zwlSdgVfn+8
QeC5vzNUkE88hS9arMDg+Hb4s3EvkSi/GngFWam6OvrjlXetzhzj2vB0sREQza/RWuZIrCB20BNG
7CMWnZPnwRszw0OtF85WlilVbGWUxX9S4kI6CeEQFQeFNpMTLXOAkEE+VppN+PB04F5CMQOis4yT
HgC4Rovvchk2yOCrLRGtVhDG83r1zFm/0alpW0beS96y/nhwsVviuhhjnVM8skOp7ml76bAc7wxB
tjKhmm7hEx49Yam/TtCamQP5Cst8PQaczjeeZCyRHrrC0s1yLd57G8fENAjdbHaotmbzZ4xtQptR
b2KevT5L+zxyMu2laiQCy4v2ljSRoznQk/eUtD2/0RRgMmcQRbHa0fMsjvgs6vR7qBinaYGoj2Bq
xNTYNnMyyrgoTD3aqm9yfR3bEAEiVc/sBdQzu4uJGldTaXMO2UhgmL6bqnH9wTAwmjpmL9J0NQvB
W3PMEyOJWIU90UK8UEtszU0QZ8e9YBMz9vpaPLJbyHsVbOpoowTlJwoVq07ZDW7OtWwOq6n6OQNv
qmCj34iIm2UvMAaTQSwtyTPpqeMedslBZyX30v3Q19EHFj+mvHqz8PTl2sb9vOkvABpfhwTotE7I
WWQUEQtz8VyhfuB1A/yczCJSJfMpCtrwMpOQ+JgPzcMDvCZPUyjRF0IYtIlY2q2ORHTsQp8nl8Ql
ehoNJLsoUJpmJawCV44BD8OvL8SM+WSdMNJ8JCSoKnZyp70aJV17IOuZL5HEpHxy0ippkYwLT3wl
jySMW+iLzCNbnrTqE2YQSwL5z8SXDYdn7TJtR3P6uYAuQqH7VzOC+KCZvi38jy3pje10zxkVFcpf
/PoxFIeDVUjrV/tglmQzktEkiViJhs1UHHhFSmc4OJLQOSoObMaGtlRPQZqw7tfpSL0Fio3dJuw0
kdCiMr6pD5P+Jji91C3o3Ue/FEsQ7XHxiIOyvnxe9MSaGzQ/ujXgchrdYLNnxekuA8Frvu5j+gCY
rgXjkvnkc+PyhvTN+jfUIBhDc+aWkZsi8SyugQorCAnf7jGwtwEQReVcc/051hTY6Wuk9wcYKcho
xu3KBMI6KMkj0yVN+Qp4WR82IPCdFu4ZUXbfnbjOfx6AurV0W2DT/cDOecrG6swCo7hxfUl8Q+uq
S1VJrGUIaGewfXK1qx0QZWiCj8KjRg/JIL86Qlx8jigosLDH2PU/doqcwMvrv0PYYPkYgOH3xSk4
2iji/ByE9onjyX7Nyx7pgyc/mO1T7rP3ivDEyHnFeADXkUUz0LV8uBbMg5+PJvab/WtXKSJlkp4Y
86pLQi/YfiYQNWOEb+1L5CXz86MlRGmtje1vserZ4/QXptl72VAvW1cl6WSM5QdaRf+qz/o0dX3O
3FKVsJ3af6LAVsWg1IozQBEdSrrS0Wr8TEe2j6IQ5CT0DTPcEkcqxUgO0zSeZPh0+ASBxS8qYE1n
Sou6nu+yQSjKMnKnzwMr3nvEGQUWICXs7MTZxHUkLGegkic77LH4h67T8mFiklCd6rcRai8C+R5U
V8ii3Rb8VKg4+V209DtPhBaolzfVdQEMm0KfdY0aIiKJ8HgE0/6oypAQN0qb5QkdJjTxrKfsfmgu
aSoRnm9hDw8Odg/9GBqixy0NU8e4KyhELaYcr7NlyxXddXNdNaCvt2DoOFL4Yp2oRf41/tf/kSCT
G90ifEOhDQkn/ylLaOZLq9yRp87Np7s455GNfx7R3nUPfLnTPssgLJGoebV0Z3zgM4H93iB9roBc
MamOCSEo7HdmErsSJs7iYlNvZ7bBSYHbsgC3UsojXDBiyRJ1oFpfKYT4vNfBsGiNdjO9czIocc1P
L6XoHES8EVJsNFm5VL8lrkMhb+x+IXJNl9BdCemnhwtptEPR8nkxu5P0PRqvMdLsxHXR7s7m9or7
gRX1YJU7+zeKmTb/SvAXSkj/rhZqiwVbAl4p/FvhPak6cEba99MUbjod9a2+IsdPaTmFjKR60RRN
Zi6ZATB1O8k8yXR1pRXnLHZ0UIUBcxDfl1FAvAW7n+EBEgB7v1Pg+4HCkZI8BlOr8WRxC9IrTnq/
EkI4RHBMxW0Ejao1q97IQD7X+beAL4vFhQkVnNQ9Kjn+kMDNXhp9Xkzbp68HA+S4h6j5EtPDbCIW
Bm8iBytAyudA8DrKmdx9cmZgkSNY8kDZVTOJCupg2k0hXoPcQqgrO2eyTIscLzgC9CsWwJJxJqle
xhLhWDXaoRDg/N0mdX15FtR+YDUNH3cni56ubT0jAJkIRfTdf3e89oQVIY6+T0+wL+MH4mEtAdf3
rjvWKogo9Mtrdqf4L//JXP+weM2dXGO13rbW1Npg7YkogZyygTJvFEj1rM31A9JxUk+zST1Nqrlb
CXmwbomLMa/9z1DsXf/E9rVho0HIDPCunCxZ/kaMYK47Tqg/cQ6ZJH0bNhFKhGxag6BQB8FDYdY8
IslsgQ0AUN4rEtjDWGGdnRdQV0e5w4HJEmoJut5jfp3CiKgaAkmNpDefRclovvX1pG75Jq97SxBG
7f8yjha0KIG5ua1cDEi8pDVZudwLcWrqFFwyCtPJTPMSqN7ANBAto6OZARkAd9bxZMS8etXbvXk6
xG18KFxtZ3DQCTnhuEhgHr+sRbMEb4HkJoepsIxjsNxj2FotAj4fJY+aEDtaF/ipi0ObXbVJ8HPa
lnwopd/kOmTqMti2wRu5qVXzph33JkgMv9Qh+F6CARBbnl0EoV5y5+9jLA4TwP3EDKMQl33lYVDz
DuCKzOeUYlfoK8qdGXaWR3FnBPtmZvXV+8kzGaCicunlX8GV9qZwVm5GCJhSoP8D8OajrWwFJb5B
ZA0J2Erp7kcPITeveHL3ej+K2xu8c0HZRf5uCckJDRmGgRDTXh6b3ZblYHH3ZRRyFis6YedgFuot
Y5korZq2REX4znSl8umkGXCGyFIdnZN9L3Hyq+K+S42yz+IPJhNQvtruqJsPvQYISAi/8uPx28Hc
tepRakZ1XxIyGf17bQEFM3PTA2mPvdqCMMYBfn9JkQVAP10qbppJUsQ3hiXF68GQQ0w8/uX1EKFL
v80b7sE6Ft+BWtAygSrvIlWTujZ+V86900aPNjakYioq50rMAlZ9mjMlrN7EsbejvYmKjJP3/jqr
vcVLjtm+G9qfwQ0+SgXx7UfgdxJcYVA7hB0tBgqdsIWf6+wUVV3nukQn1H7QcpxwCO5E5ZpClzxc
te8EThWF7vZyu55Dec4YF/dGhGGg7CqoABbUYpx25ZFLml6rVBbIKtciooA3tpzP0FCordMeTRvG
v9ZqXTL9peaSGsFVm41E9lC62Xt9KTjYgD1XRMAP/UCSSgiYJO2Cz9f5CZn1WmwRU+6Wua5WZRwe
VnlgTTQSKDFjgXX1vcxy/4nB0Igd826QU9i59MIhg4Arq3WbCeFazgwxpClag8MnMq1qtBxubkHN
skPtJbLXNYGmLlCi+ATXRC9g9/PRPXjcrEhNp5bipmbN40OXqRbj7Jo3Ej1AXofaTl5wB5iLJfRm
iwNI8pr5bK6Bk8xQEVGRm0JOqm2RMxPBepG3E/ZAVAfmN5yvP8vKIw+mmwR7jAq7b2l4VHAdH1Db
Rr4QQFR4p7Z+HjGWG+lONYA5i+lRngTSiSytYWgW8fE7IuaksCC02e66s5FUE8uIfxoIYCDogrrD
JOX6CzI4NVeI4dICOSZ1muvgm4EvjiluskSD5PwhooTme25OdZIw6LfG9+LI1SRFLYav7GQslLM/
2wDJMrS045hweVSk3kM5fvPfN/B6RS5RokleHGSo5EOAk97AcPWLDjsR+lCTHdxYN/cbaOfvPTNA
jR23km9A89chu1ro0fSIIcv59ACF5u0ZQtdLxTuURgY2/nVMtdpZMW6NRXz7Pc+4P3JjCKfcunPl
KNKXp1CyT+W8Stb6PoaXJHOBOFdCr891TrnMW38vWWtqCWEK3nlAkT0AcD9bPXL+aO2sDcTV1ipV
hd9eWRQe4IGV+xYQWUL1fTasIspMMMwhBbKJ3zeKr+fheleGKtimLYWuuAxnZUMFvagd5Sq85PbU
mzQYReMx4PJi2yUH6uuJLmmAzJSQH9+Aa2jQLDsCN2I2IJBmQzV1RU+8gZS8BfQIQaVPfakzMuqg
JrLqFr1ALNQm47SvuoNHspeaBdBwCjiyIYCI5ot22MAKxE2hX2Cr2Jiyf2VHrojc+f4yh232ARIN
2E41lyejdYjnIacvfkMflTFHZHQpoJEWS693oFK64awx8g5847ZrXgvdffod2B0Lv0Ohcx5NwDEo
aFgZCJpI1CyHpBDJ+NenphSbEWUCkRI766xnfnv88+0yOMB8/zJgYvCXgVPUl+YNbOJvCG/bKEvy
SWCNJk7oDmBVnma4pFpugciGy76IAMHKELBdntWZ6yv4Sg1nrX4dFV26h+XhdNxqBTpRRmpR8wmX
k8V3cf/FqwfRTVqVa8FzfaP5tXa1hjFw1ZDfHQPX3ZRN4Ur+m7XPbjFBMUzpxNwghJaVWd5ijFgA
ETU5eOIXvEl4BWoVVRFe+/3U6Y2lbqYIkTXkX4k0cJFcBpWhg6Thx/ficNRSzmUAen2CdkujcKfU
b6VyIPANdddJiS6KAKPPuQM2OTQfYj+8IdJkpztqLHq+Iw+8Kle5OmoGofnc185CbsXO/ynirNiZ
c8/mj5MS4lgSI4dJPSvgCXhHq0gPIHBVfpZdz8G0lDY629pjO0Ygr1TX2Z0GawKToP+aq8cuo5kv
oqnq6e9fh6m9E+7YL0PqFA2wfxWaB/Iyrz1J1HStgRQhRmJMiyWvsHL/Xpb8ploch4Iz/QbQyQ9B
oJMwI0swrKAidsP4hQ7Mx6gYGF4I/H4vSgPMyrG4GZHEAKHs+A8VD+vzjiNGKjTVdovdTuOcCqfh
mb6LRjRtuwA7/BTaczTxD4XnMCqvWSynnhpZ0f/LX82O+9OujjwsheDX6XB6UHBoyZ/t7EJhLhdz
TweGPHLUdTCOaWOX/sZyG/ZBBdxXYV2ufjrbb8NgJy90iV6urLkLLBuXM21oOyPOuQGI72M5NqUz
Ax9sNJwTwpDYjYdDcOzOclh/DqWvopZoLVBxTNfZvY3RFH/CcZDVj0Qrpr8rOVQ+I/Ov/21BbnWO
N1o8YM/3r1ZEYu86geP4neq/UPrFUmFiI/flNJALDL4doANrZvQf0ixbzhvNRHuIj9jC/rw7+HWt
LLicA4eXHrEnwEEI8DXoLxEdS2hifxr69SO2UUyDkRFBSaQhGtoeaObxiaCyeffFUGRKTiwfCxYp
JiWFiIzqtFDfs/aJFy056KBbJmqOLKik+vIpLdgsPPKvQP850Cud68KcnijZzkXo0BMQPuEKFwCu
OAGXiLUDCiKNP6ofnMWcFVUmNtyQp5U099Y2zOpityxIJ/hcHuA2HBcawhrahZ7SsADbU+WHHMOH
ZXKaGbdU65nFzTVP4LhKPlQ5xqbKAOgvPjzHlDFzJCamUSD1jNUQBQNK2bDCP+w5MuY7wcLB9Cql
bTsKQ5nimfNlQa76kDejyhHyluY/pfDPKE02/cENlSxi7XROx6J7IZWBrsP+FPLwOB/MZJJyxMzZ
eEFl7IYLk1Hw7SjI5IkW3IEAuJuz4/oDhfR2vPC1cdX+UAlxJQDYUqJ8CtKbks1mfOztckQ8+hmt
w4sN0b4kc+zupIjvrAmgp/5z5C0yHlCV5PvMgDNH7QcibKybw6Z1qiHNK6sVZNBDYT9dS8UhNK7l
56Zf1PiFW2pRzXzCEE4AGCL2dt/AF0eSggKyT0kBoMzNFARKyivSBnPwGxaHCfJxE36P/AidL0WO
0tHethw9DoxEnDdP2ok5ubckLFMsdOtX33qLvrEjuGU/KzumZo8KaA+F+o6YPhQSf7UTmtJkr6+R
JSzQvQFdwRHJp2cgBCF7i01PpK8XnecY1ONwuk2ngzAR/2xelsTl8kER7yVj11e6xMjJZnY6Q8nW
6C5t7DGhTuqEVnQlXYJepgokYY0YQf3AaVMXOb5Rp5pDFsZqhWo0ZHj1rk/PfujjlJvXxt4GGVAQ
iL224r1mWoS7Vwf92IfXBjiLvOUqlMtDyb46qQ/sBwPkd4vijNNKchE7O9lgsggWH8ETd5y6ddBr
OrF6UR72Rij+WasL5ydnF4a5nDQ8Lm0WIJ6F6raTmxy3yivkpHLprkAslzZ6KLYyNka2eNRaGkji
ijN7Ifx5n960AOPqnLA6t759y9SrL1+DhWBiDMli6F9CMJQpGB1MG1xTL58x07JAMrLCE5hLjivN
e1SdT5rScX6LzCk6ZGZrMPZ1XMfBJCp0zoFKIf8WB46Tm/bKt+58HMvZBaVQGV90D1VpUbEXfujt
2piKJ0Yl1RFCjcgwq+p32A6gLDPwMaNOt3X4Gqd2GiUcLgjSFTyWq7HcXm3lBvu417sJDDZO98+I
kFrDPuhaFrANF6EOf4xHqhdkbGDpXnXrOrsgoEJvHU0YGthwiWMl7gg0UMvXTmD2TnODlKoVYE94
7bXX9eVBW09tOThSjCXVfkr7sapat8+/xT4Xww38xCZC+zWsbe4M9qHX++8CHOr23RIIo9+9YSna
LlB9IlnenB0gAJZqf3uLkGw/8/Cvbzg/EMLx10mPKxfN+61ipOVh645r500Tc9vTBWaTyecvMBBk
CfWQN3P3A57OoGECRUGEW2g1wBt2yDXUVFxrBGg+TpntI0v/OSmcArnzBwBDe2kF416q9rVhdJ1h
8yPZfD8pUaQdmSt1Id8gSzzRlF++sqN9sWGtgO16huOBvLFKxYheN1bQIJ22Tz4/YSoNaW9rnc4v
FJr1xXEFduQuBJloDkh8hDwhVcRzX0HTcRBjc/Q5hqOZ1q7hYXV+hjoIEjqHpcmS2R+6yMTsa0IQ
aoqPnKTUJ+0Axpf24QEUrAarVCJVZ7Hp1mMw68agY1UmndVitSpXjTt/OK1KoJhFi3SAUZHBMX1N
JlDzW1vgijivinogstZKONfUupxb318/WKErIsJV8S/hkTc4bLXc4W/vkXFCisenAbY+iCHO1GZy
5c4CXocaLcCOCO+wU6m2yD2aK+1QKDKlI8OYEnoN37NyBVUTNFQv+A4g1jvcP5kjmiuUMsdGtajv
NNeeLugauHGV2bj1n6yXauoacM2b5wFn65NueFqQM/KTgb9S8qONuEPdVqdeoANza107CN6zuPSg
p8OvKUOzr3cNVi2XASFRrQSLqo3BzvNlQCNG18UqPNC+opbh89tjLgi2D00JhjFj6jyaxkqkml0c
GhY4mLl3ZFGAyq5aco+Ik6Z3nC2/Rj4gSvCIO/nrZm/vxbs/rpVbOSGLNjwVgnrxwCO8mG/I3lbO
L9rSICtn6dCDrUVcFtygvzm2rDGepQl0PrrkuzB293WNkeKZAS9mNhzEKlnKrIYnGkgSWgxbA/wm
0MucPP/m7E4CEGn2TN8dCcOIJ5N/VR+JZQmXLnBew78eVWnMOc2uHlquwJ3gHOYH+TZViul1ytNI
QYV1oPAxoe8nAQ55hG7AgQiUHCzjFx+JOeruMGyVkVMaLkGECr48HKxKLvgZwycJMqIcVA6BBRL5
NSUXaYRpQWEGor8S+rzIqXXKej0mAdOYwemxUOviSs+00VpQvNgsd3h8E9Se9s2oi5D9dRCqvmL1
BZbbHm0bbXXSNj5T6muhhiP59lW7G5qpP+KDQyjteTUwzCcxjdSPIEXM9ZMBfqUOXHDdPUcVyZ5k
EOu0DUz4Wuf+34l8g4zetNHxmyJOYvspF3DAf7zN8xhFdV7NytEKZT/t6h5PyZcx/LbT4VtlA8yE
rQNSwWD1s5YL9swpSraQ7Eda9rDm+yN2WJsGd+4mfJEAOQk5PnUaLgPa8Krz7/Yu1MCeZG/4xJb7
2DqG9a7DT7CBSWSOaYX/KlCWLxPICZihjJrh2qsrQt5RweZnyCW4Gz6dCR9OFfElvf4F18RE6sXq
/tcP/qVUgO6YydstXnxtqJ28cN9YJY0QkDXFvCtYfR3jBf0/ZGLyipc4DT9M+n2i9oWoj71cMBod
tENzk4DiE954+RG2wtAhgKHIHHdeZIfACXCWzG//VXINNvfYcm8d7YzSpD6h1RVENgQB5Hq8Rfcr
g+pq72bhC1uqqrqGRuogpmq17yHqx7H6Kz7/GaH60somKLhedPD9g4AKXOk9JdMoIAW/Xfl7jmrK
/Bv3GTrNQ5cncZiF08jaigN4FOdl6JW5IieR+JwvtLs3EGfqEywVBlhWngnpcg7mM8eSqzsFbEYX
6DTlf5Lozvbbf6cwey+8Nri9GXOV4kZLaekVUUuNPbkb4fkhyTh8WHbiTCVn8sSZPpuIbGZ3nz++
mdV0Jd7GMwNZuzoUkUCZXtsLC+tSJOqdeILK3CyILS3bhs5nbKpubC/lphuX2k8TJu4Uewu0aNCW
x83xY76zHDr4nBmlPOrtOP3T+CGDZ0Nh/nin1HjDNPpmMa66qWsBGyVcB07Z/V5PmYv2K6keGQe4
TY4/JgR36W4O5MXDoMU+K0bzxiN240++aHm3I6C5/kmb5Oiz7pV/Az+izPRnbIIa39zhxMXyGTgK
8bSbDPqzWfGU2wjSF+JbfZgdqKsAnXtIPsdtHjJXauTf8Bz89xRyfDpEEglu6dDHa061RLRw+67K
bDprWH8Czh7ZnYVmOWWZyEHeXt3ULzveihK32BR0BI9ZXlCqDKpyhZejd7qHPbDG6qkpgNdGB8wr
13DgGIw188nQDo9A63Q6DqK+wbu9aXaYXyMzRvhhgIciZFGYCE34/kT14GPDl5T1vrhWOS2siWia
bbUMymJjYDoA4fCJrdMIdCBqAj0Cl29ut/bTA8NEVJB5slVZsjREqW1RNigTDblaceNPb64Vv35e
wh/gh1PUasPCumOR0dN9a15djsw1gmCkH7sTxFptcHpp4mG7aJi0pFzs3/XMnihbeFO1FSzdEdfO
bXAhzYiKvlun1gOnid80cEK1tZ8SrbYdrCszcniVVcH3oJ204TDb5BK6JesJ+7lxk1eIjNcH/0hd
MDzaAuD9U4sykF4iNvB+gRT9drT4lgA6xFrUAy0xsmRb0Rr5HtpCm49O/Y9W4VQwLufbsAqnw7h4
iEFAtFmluqSL/bBR7y7KcB5yXjZrBM4eloH9JPIRxl68aaZ1Jdc8TBFiciz36sGmalfAMCcFkJgi
jNdH35ZrJCvLbygMpan23eMdFHVtBG0fZoAqIYzahXZxIwCMaIiPAW3uA7vihcc2CPYvRoZQJH+v
Vy+HmDNkmNbZTZU7IjH9aduUA0EFMgpRaB283weF2fnrmelCKB9EKYGdrDCKfqS01Yf11BnT70lX
a6Zy3EPm7sB1UzqoJK1Jq5OugbjsWOySNN7I9YGHsY2FnF9m9w5x6KxL6N/77zRw8DFZmPVYj2S1
2NKz25lYnbc+tJcgqW+GsqbngTEH580gMq11hPuALrltpdxtkzWd/SQIdHHz++AjeE0kFdwGspYQ
X5vFWMtaR28kzU6gnvCGbqoMxMBTiH8Mi0mIsJNCctwyQA+i5/Hkh6P80jm3xsJn83NI8ouZdZKc
+aGTzyNCGyDanZephsMqiz1FT0l/qrG77VrwWPRhr3SmYQTfvt7EzMw5OHHrTlqsCs+m7HnExImU
h1U4p6qbIH2Pk4TbJW9iXsASHOSdc5lFAleE+rsjNgX4IX5YcOGdahGltudSsrMzdlZ0m+IbYsWY
X7OQl7ZbFJoJtuF8KfAnYlTnuVYwynXFG2E78PUMV+RgkyNpVf7xx8gvXvUAsJ6wbjOG1ibsmi92
rnJOqxp6F7mYZaCIUOoxltSB7wQwmIBsc56moAfloycNC2WOmNvb7aLe7mf2Mr6mktYIDGAuQpx8
XpIYzf8a6lXn4SFIRh9ycvbZBMUJKpXkyEa747o0+UlKl0O8AD3MoOET2ihI8bqOP4BO/pbSN8Dd
W0gUho2DxyqhGe7/4zWEQwhDnegnvTfL+XCz9R5J8qEoMoC3B9xHbRZeXgxMu5OsKKf6uU0KTCA1
dFpWMorIjrldksXwjLnhnet0uTsuYtOFM9W2wOwZwHG1nJE4CdajdNVhixYb4gMioHDu639HTs57
ZvadmIJZtcb3PKh9GafQqX3mEOJvZBX9Oz6r/ggWFN/VVQldklhBhZWvvWYyarxISFeUvYz5rEXD
KSJsasUwQTfGn1mBKdj38fHk8auKcXFHLugzxi24FTAQZvrFJj3ebqQzAkG4vtWkZ8IC4N+CyA02
7j3B+S2CUXmxZG8oRMBWJmSgYNL6V6PZ3CBnFljkmJFYXRmw4Phe/2DNpelIA1Z5MFrVqZbkemc2
85YVaBBVa6g6Tas3Ynrvki9LovUdsjR3+iXcciFPSu1emn1E5vK38Th/91zzhBpaeVwW4eYjm6OH
vWyiZY1agK7aoX6bRuX2aP1ylDbCCmgMmVrINwD39LXA/esnBvnyjKe3YoDFZGd+txYkqFIVuTWC
HrW6K03ixc/E3f2U6Q+m+nUnEWKd2Q3qXIf5dxnHG+lJog1UihmK9IdKNBEp8RypjCxEDpoER062
c2eIrEn8Kc1hGUx0mVp0n3mIxUyE3tJDHedCiMIKmVlFBUt5kBQoWbnc3h+N1V0acEG7MN3whCJv
RwSznv0OCtinvNrD6t6gOqc+PJdYi/f1JJDyekxzXNHr/tUUha3pqe2ZSjp+uY8cCpmoAd6Jz2xg
m8hxSzDcvjq4fjO3OVuRiV+Q2/guuC41OOMAJ9GdGbilt3ObPEmbcQvm8/d4l/roc8onl2ytsrrh
r3ZBRWoyD+Z1bJHDBfq6TPXHrI5Erz/Qoq+NGjxvjbzDBdpESeIxxuFMZJiJGefQ6yYgg7Tr5GFF
Gyzr7FFX64lWOF33UYOC6NiD7Oa1GLn481ouqe8oXZwzr8dw8EYrjef+1NFdKL0KELxMVxP38yQC
x4GSTWYTM9xyOYQE3KPKeLH4DCgvSoy+hUwZA5aLBZu8CqvWj9xVSPRpR33gxKAjiNvhl2k82u9W
tMvSSLpdiAvD7CSxCS7+OMclRjcFAL0SogBZCibV/KTNpWEDs3nwRhCQh0e3F/9pGcQhSi0IL6qM
m2x7fKbMuN3G3djanmSn2JZHriWpEsSaIM2Saa7w4Jnb7WY9L5JkyAeqcvqMg2RWlSgdGouJeave
yEXxg0sMC6KGxBj7uM/ctRc+KNRK9uGc2ykdGN7o0yNFmzGNKfb6dnTRMGZCh0LxL0H4rppdzpY0
OfjGVJSesSLRTF+OL/sErwIujFIMoczv59KRZmQrOeXJDDrmWibwm+wv7+mo76KTX78xHtqtPC1g
GFuPfkl5WWe2LeUoCSMRxB12ZvE5jZ7P6GDw1ikAqP7HKt3twscS1Zl6kAOdwkaFiYFyEQdmzQrK
+k4zjdPs9A9l8SuAsQ+74bX7Fc461nSJiFWtrSPjqSR1yaIa4pwXVs4UtDVadjpTxnUPL0BYegYa
SzKJQ4t3skZzmmHi8wvAEVGNJTk3A7/hcg8WaRehKWzAmUGP+DkFVaF5eyhp+dZf6vC0OfT1hLcY
RkGLZ9olQWs77KlLk/UMOZukIUJbFP9kDgJkGuvpp5VHTx+GXr5mfTF/Hbu+Qi/+mfmc4XWCPUux
O2jFiqNHni+HZ0hx8l1DhuKab5zlxmAXabP1sWAdRpJam2uceldYtOI0tK1lt4E/fUE/XJmG48EQ
OgVSQAlpb8U4vyn+GHQgfPr7DLtbIRDer4ePyGez3hhrB0wOW6WOgR6k5sA0cgmNS0P8DbfJdTr6
bNnpvVbRpT2LcgwtE6q6jxfAv8/xmqgxwYYBNHa2tkoXwHpagzEwVx/ldzMraX93mEWJnr5f3tZI
QqAy0jQaZH+OnN93YxvahI62pLHxPwNrXrDWXTe483YRtlO4I4FaQBPI2LpjaGj2zRFz7qKhbqGe
9zbi1ltFYvkkibdbsusOXp1i72UVQYJXBvZjZK63YZJbgkOgoVSPDlSSHSK2cHBaDlX/k6nHmtWF
Mi///ptyJvjDe6x67WWxTmLIKw/2HiUG6vLt0pWaCuXRGLMbXEdn2owueZxdNlh595dyDh2MEVDy
eA+euoK1mXPzE2B3k+YkK/2HFG7Hbn9AGzZfSWMqS8SM2z7i/rczYhX1lYsSK5RDihaLhEEsJPt7
+1t3KeJCxVGEZm6r3WwtdALbpMIKW+N7c5P1LRYe21vKfxI2gjjbnuP8ttBoU4u2xMHU9lchLLw8
AC/QblImYQmxaWm24KykYEQgcAoII+BHBzaNbLWTZwmRgumA/3dg42IX2BWvLX4gPcOG56RFanm+
jOmmqdB3EsdzQQ+AJXRIm80VnSkeXObZmgsGxF3x6jxMg8JvZuCGd3gRIZcJEKZMIad8ZNH6WVOA
hty+hvZ8X7vxdfrZ22HJhOe5Jg/Q7KqA+egns/CNP4WWlZnTZUkn3ztW5mzXlb3aEl1ew7k0ROps
oe1sdsF1rloDgAq5QBkRT6lBs6mabsONiIe/gMfaS3Y89gT1hhNjjAnzWdnKoogwEOIwGaOpAI0i
4CKyymAWK6fLmwqv2JufiX3I6yAZe9yqNcclkfgg/N6Z9Nc27f5ZfBKiayi96xoSLd3USCQGpbPL
cVHwbXzUSp1Tw2nIc+Dyqlg5nNIyR4BBB8ABjsOY73KVBvDb6GSPGKocppxwHlcgIqFXnb15Ta90
7yj/828o1dS5iPariUMrBaNGIB4y/STxQX/AqXQEOFairyz/CeyM2xmfLrKx6y9aMcZjKo0liNSj
pGkluFD2rMn6fmHECDbd2BQ7t3prBYWA36SEp+YIbX8ReMdjla3rPo7dIZx0IGGP/3/YtrG0JZUx
xUjIYstBLTzOu60FgTsvl2tyWwX1HP0DPLObcRBf1Aj/vDAfBe0REXNEi5NFdYJ+1Fb4ua31ajUi
csUaoTMy/1mZ6+Li1Po9pZwc7IuPsiN8n5QKq9wcrFLLnGW9wxsvFFp7grNObTwxFuvGeVqf3sP8
lLDm72QF/LxiatPk9YL7RdIfn4H11pHd1zmEFeBVqQcJQNSZhmgbCxg2lSgRNs4qTAaoVk3Yp/ts
whisFIaBRwAP55Sqi+0OzUTMzyh9rWs7y4LV7aq8HZPgNp7guSFXXY2Qj6guaAJn7zjQOfi5GzVd
VVLpi0EyLwJAXQJFEyj1TuWh944aLo5xLEyiLh97N6CodweTPAsZn50ho6Qd496+1H8ttgPPBBLY
g81D4sMkMaOvQ+bh2N5hRFzHXuDzriItxOv92oVc9RK2OxKzWQ/701AdWZOPdZi7891HIe4yhSpi
D+cRNmy4L7iI7DWLVTpiAQdF3ltkejJTQfSAcSJA0zF6QLrmKQQwCGPYIlsKGDnMobKKSpD+IeQQ
7SXztFCpmDlITNZNJ8ehuZdzGIYMTwty+mCjs3K1o0UvREaJ/I+VLDEs3NnjkuROkTOEKBusHZ2D
Zm5bSWNPUnlq2RVn8HhsaeN9Mp0F4M3k/Ur+46VEY8BUU/yaxGpyK++wUl0mkQOKviFq+m4P8/0L
MWtGCeYtkQL5gDJINg/XZYjDbV+cgPPRLtWxeHU7HSjsuDwJXNebr+SfpsLFtRtkTwDbYQXfHrdp
YIFDFN626pu4ngZRDqrl60AAW/bwvwigX/DzfxtiIQSkOoSb1hcakbpIkun+cgYjsmR0kxHTzFtO
i9U12RQSnJRRW2g1FHDG6rzbM5FIGdrhBfV5pdtu4E+KoKtHJbCxfkpPmafCyRxhBUbIi5eLkwo4
7nLaRWY5G7WoBMb3L6jpDZxnXJcOPJR0dJwrH7I1+aOCCvmVS1z/YK/qQK3COyLppeMwXWKMT+9G
P9wKM7DnOun6L4ncIkSKVyGD5IxYlsy2u8zllH59hgWvbBiFBoWmU1T+2SBTi7+uYa2UBauCU82E
h++fM+sgk8agsBmpo/zxumbMjlTzP0ICIYpE4TwCR/Uhk7trKIkr4kzx/ONxbzwzSRu8RIHZiad8
WfkdIpIVllIg9T5NqgrFMTskm15xgXA94/f98fGYTrbuYtBEct6XI4/RYCxuO9LizPQ74udY3pb/
LTRdHBoeiMG3MVWgDkns2J7ClykKzjPqQAL2rHkEY2Z2cn+DNeqV2PQJ1fCh8BzGtDIGpWcJA9Cl
TCMxseeRgDug2MZv/eooxCWSVuOCHkoAHhzIEtLvqEELzJ7r/7iI/DAalFOHd1Ek8fW4AEvl/nI8
201o4V8oEX+dhqZzfJYqurPAjiHdHvfgdT4yFlpqrr/lVFDU9C2a2wfhl5rQRhXzYQlVxa+gtp/o
dJiS+KuOs8Zha5aNfmscvHJG5P5rc002T8g+bscxKK0SWEFO8Ph8S0rnUEisFnru2xX4QzQzSKJ3
2r4MDH0K/COCK1wnNsNPhWm2TzlM1U3RitsIH976oaJ58vMUeQRiLhw66z/P5AapabAB9I5HXoa/
JC3DFM4hDBfiOyMRdRT2QquEN3xDKiq1kYfsT06fZhcxxjzLcaZlmBEIwfAZqZ9SsyqKXwJeb7lg
py/GEFlYhzb9UryGw8J5ez9I5/Dx3wvC8toeRk3IzvEtUh0GltNH5PNWcdA5pAOW1q13nr0xwjvy
ZOClCYUd7CqT0n0W/isCPOsswKbTnuhqm+WcyGTplTC6/JdsJ8uKd/onNQ+a99ZjkZ+xSs1C+Laa
qOmXNChBdh8sw3fmya+rIEoIsKqZFsZ/feFtEwGWfMaSszBzeH7eDSOoG9sLUqkSYqokbL0JHjDf
GPlQcPvoP+sYs+D74yqc116zZeGGrlPzEb/QEmo6oiyinHPMw7DNEzotPuZO1aBw4sKp/ut1ZSl0
Lk8g+cJbQwwQKWZWBGS+ugKV8/X5gFzyywjRwCIgKaHOzAaYVtnU8CnZYXUJhDPIkKHhMKbbY91f
MMUZyTabtXF0mgDx7CBw6ThzoDi/4cmuzpn8ZajB5uerFPl8gmuk//vHerqKcNT7LfvUwm6NSX7A
JCPw8l3wfFA6Eb9zesx+gG7EU06FULQCCtWJsn3MQdKSmDCGHJzp2HnZeveDmZwjtXeDrT6GftNa
jy1L4SB0AVlIK7ejyGEx7EbcBYTGBT4/iGwHXUEQLFLTF1s7Xxv2yFpCI8/Yog8FDtFnMZsPYmnU
z1SaXLCIHkiS/UuNAEqlKB/vauqhV1lxyAFwZf0xj6FrAVXAfBd53j/t4IUDaf7QmTEsfmVSxC5H
Aczh7S6kywg4edjTHZC6ZESRo4cyCKZgHrfrmLqysAX+7MEFUTv1KwuQMfVy9g7xmdtz5ROQhLBl
WXa4b4Ff4qKEXPzxoWy+5xw3LIs1bFk+Kh6sCcXfrpeypT58LuQYYBbSQ9eQv3H8fh8uGPAb1azu
5hvONnNv422RPrsYo4QEbGSBtx9AslPBcnt+5Fne49hTEf4nSvagEEUUdgHd0I4VxBRuXjUmQ3Re
eL9tRbGhcJ35Rcn5buBzNojZZBKU1fSnSWBL37lGSk5eNXsEXtxQh74Ll5JwW+FbdM3m9yuE870o
nk0H0brq6BC+n2OqY21GwqHshwewASy8BaTZ/5R0gBrJ6Gc/okw7vS5beS0ZHp9CuGtKVhlJbYr/
3Y/IaEkZjuEXJrtk1TotdRDdIUqCRGA97iVINegW21wIRDgny9rTgcjeYdIJSbIFc8FK58qMdfEb
rNH2YriiOsQKUZuJD9xRdYOltoJsAVeX92ZoQPUUioc+Rc9I/1w/gBYgqsR2USd05wYI7/Jd8ZQX
EV7jQs+oqh4Iu49TNCXln5QIXBm4kZd6DG9z9pDcPSMIs3nlC0NcpS5RhgBOW8hnoUoPT5sGZNGl
UlbuA34YOA8Y62w+0f6Bn7atf3gu21B0u4mOamFn4IYpoyf1TOn2dLvZMe6UYlKNOUcBHE0gdy0h
Hm6Pfkw7L0OSKkdZtX9ArOEg31jUHY0oI8aO4iRVe4jRhbkjnDRqst5xnHW6kF+EjdCBYTT3+YBZ
JRrKYTEeK8BBkKeOsrqiPy3eryfitIZYGuqnhiqRuNSgboXos9nsz7GNOsRnq6enATTPNO4XJrCb
IejcpZIgmz9V00xekla1zx50GsOyR17FFw5m4SXPz9ykLeTc35A9cN9ZJhwgjF1+inwNlLHzMrhl
tG2CHtyW0a4/EFGvPY94tzwIqUvJmul/GFIcb/wv5JixIbYkvWRNxXZliXEOIXXBk70uquYy8axw
AapKwJvghZpGLqL5aikDWSgC3gJVd+2WLeagpspUGvuklOt+zWu9U0rj+D7YXq0O7ubfmxCkMOZp
JoRN1Y8bsEDNT7hf6rJqIyrqvJLyjmHB7VIA5ctjhTaCavzywI7HYA2Zewd4y5Vbpn1y0m4qs3nG
cGDvIdfpNnErqx8ec50YW/sb6uDwI+ViVLnk4n/vznDtF/I8fHiQw9AP6BSREMl27e3fkZlRtGej
8ykuLS7BdyRSwq0yPKYrnSQeUdCdZyYGDC1ZZbPaRbN1MX3nb/3pHEcpNTVtL98hOnXJdh1yTa3u
KvLVaTnL3krNVCIDFwqrwz2RtzgTCe5TDDkThxk597q8s3JRNkm991/VKg9B8zNYEWcoCCSDvjZ8
h/1h15d8I7fkPzTX3T66d/iGvhn0s0CeTANAt88DJo+AE6lvQefhJ/67UCBVG9h+GPEOjUqQ+ASh
yMPBeVsqXra2G57HdXVnSnEh+T9mqk4IgDiXA5v2XTQCugkZwdKhGCkTl++zCb8GfWqv2L9+Ejqt
ev6DYscFoN59Wf09e90DAddu8QJngHfxg4QOkMeyfpGRG//MR1h0qK3BTIg0RgzC862pS/gl4j3H
S3R0W9rZAjmsQtHLhZpk29wsLPVT3oRIkFdQuJShHPnRDtVSY6QqE9xCzR5YR9P5K1gUiEh5bEgl
Gy/4I/lA9UENh5bf+oqTlFndyZnWnR2iXPUl3cOloGSLcuvgQTvaOdCuSS86kKO8VOaKQ055eo58
jGIXdzea4CJfZjZe+G6FN7ofMOnehr1qZhIKeB6RQ59BKqNRYMSbqGgrn2SVUkDYIsJt94nViieI
5PxhqeUBfHpLOmDUFhfA4+B3SI/L7SQAfSJHOByIEMHUhXVq0a1sT3/tKvUhwdbR4Jv8+J1uOvSd
f/ydYOu1Krzm3oGOPPe8n4qa0Oxy3tF+bj2VkpDQb3I+S9tN+6hu5omKe/xEuT3WxpasShJbSM2I
xLxD/4SJC6iDrcxtPLJruw8SbXbke9k8SwWVyJXKGaOd3DtRwzDtwLiVlcyO0UyEdja7Yivv49tt
Y0rgy6kaslbz9jqJIS72ZM2PNhCGIlSmsGmuxrS8wMkROcqdMX3dyhsTPcKFRdyy1883NF2EHYJE
Diuhu8CqtjErMzqO03A27EUtmAaNEksyruyL0T8k/JYAsU0HwUQknPrWZ/PcMl5I0FPWlFwX321I
TQdKEw6h9EKajxARxhx4TvXA9oyMBfjTxEcJ1wjeFy91zrUbsvECMOaLt1vt0G7kd0cIehNAeklN
fENEE/re1aXDFBsv/XraHBczFQaKOY+0OeDhrzeaVzlu/SVC7Cu+Mzb86EqZwtuI8KXN7GqkrfMK
HUGaiaDvC+152gyV2suuDCWybxDYSXFTKrh7CbeVgdq/brVEXXQNuc6QVTsoMWB2iw21fRZnszOw
x4G5Gam9jSFEnJSLIuSG4ck3UUdxHHG4zjcYIXKh3GTBPz0oSORLDZaeq3OLH1j7pNI/q8WkdlZT
qVnEVjQ338TVEIeXXf531vTs3vRDhHqPZKh4GHIpq1M0iJay9xDAXzMNHFe3tcczT1R/SE2kZqy8
DJbPFkARa56o0y3ABYu1aOZm9Gg5yX5dtsJmPww9ADZacxw+q/7ZY/ltFeidSbWAjofRpPCn/ycv
eahx54dod7yibXPRyKYsZaHziNxiEImrVgFxQQh5igS5aubaw/SMtJSnTrCho9C778+IQh9dMFYg
N65Yv4WjqdlZprOq/ee20xp5KTmFxB+ZxfYRk5m4PYSC/Ai1tps022N85X1rO+3Xw4UkjyvLAwZu
zHw2SETFmfkiAnejC9MImN6nTSfo7K6pDcUNxui9/XAnp9vSqPq2uZPrGFdPxHz581ODH9dOr8YY
AaPYdJElRgslsU6wi+WiyzmLR5dENa7JBXeNBkfYbRybQgJndMbxhc6bKKYp7D3vdcWwil0Cn7Ot
/wkE5KzLKJmlBps20t8jBouAiAqmcTEA0lTQNLjuWRCQ7DS8twT2bUuf3UXoZdau+nFjnWxkpkN1
W5NhV/hrYpagiY5nnAQFTTreX2rfedF2fpLJnHloaPmtLO9T2m50Sxc0r9trua2OWiae/stR+Iwf
xvCkr57DzlsXuBYU92+s2zPMuuKnOZtXS048FE1cYZtOh2O5wetiV+IKai58sqRIx0SRH+54JtK2
ZJsDR7LWEIC27aOH5ZSr2K98IOTcDqe9Kg68oqETYyj+SPJGI2vbLAWLasj9ySRLYaoktIUPYAeB
fYQF59YhE4C7IFoT5tK1ENxC5rLC3RS/CYpODuv3vRmc78K5jLNjXU2nG36QAgOGvC/qaJbg4PER
J0u7iH8T2r+imwTjEoZfp8GGfXe7xFcIzMjtOlZsfu+nKyINJzqusnFNWJg7DboH1R8mfbdp2Tga
c46WV2i6kImX9Gd09k7gG3bqKPFqm0FXvKCzQZf3IQ7DGKAUMrlrbT3LdQZKDZifDnW304DmWkGA
6tRH1fCJAvxFWNKuYhyqUovYRNU223CaRfL7ieuKyDMH2BC36VdyTOt5GUOdcCXJeu1os0q5JxFA
ekCnuXbbh4zgxcQBUlfS3wmgYjLrEFPJiQLNtZcnLOJ3WC+h8o7B49eQyk9R5rooLo1VxgjmNooJ
6rsvdKCc37n8ZElUozaW5CsNU8QzVb3vo72eyFcn+zUBLBBEbyhmFs2EbhyAWyGUuCl9MfyIDPCX
wM1ysg7XviY8V2mlKOwFDWjKtTlxVnKxmylunDVO/Ve6l8hM1OMUH0Di7eGGjlZH9NFi62azfuey
tPyrY13ZB8RRMYjR7RvItmh0y7Dfvetgl+XZnTseFF7ZkNgOCYAiPib5ulfoeCwvWYPT+Wysy8hU
I68bJhfK+x9n0Y/EMpLsDwX8ygZ2rGMW4F6CB7aTux7OKZo7Xl8+ngMX3cTrqrdoM1qAOZJVSdq+
FQ04TmcC2MMjY2IprEz3Dm+vznEP5AMlYbnuNSLNzNE7/TC4QksHukZ7i9Rje9FFmCu3BtmcLX30
l3CYVFkZVSKmt0cMVYRLAlqo2xZMVMayeItcHjeIYnKS/lefTWbIEbNQ3ZmkeDOvOgibeY3+apkD
DXTWNxM3aFDZ7X4XsU8SDm3/w0CgbBLki8NrS+WpI9K1VrgXpK9x7vS6aG3Cols5crbeVF4bH4tY
3v/ilSKs4pRZDjOflOU9tFq2fXkgIje+mMDmW+vjrXMFGH+wLlLBfxz2tSSRJxzEPEmgx+fx8XQx
mlM3nWAJLZdAn01tULt0wVYPogsaZGQVz0PprEAxnbibqqGCChkPk/9v1qj0tCBPYw+O/isXLC3V
KopjJUKFDlFTw7Ec4daIKdv4cDjJHKrJ35ANkh5WjE+MXspYHDsyVQ1LYoyJtnJD2HEXOb+2ZWNk
12bfqVySAqZzudxDfl7JndzWIqSOQmTS+JypXuY6l0hUa5aBNMrg9AEPNxGnltSOm8Potuih+9WM
0PltvFwuayiz0BUjtweUQ38bIGn9czMYUz18p25W3TJu8BkvbXmqWMeeCw5+tIhJLVhKS2yT0LdO
DnclZ0KXWX/7drCuKNmG6mR4BE1FdLWgur0Ypm2ZIiQiUtswwp1Ce8iLoFbGSmA9boDYljSYG9ks
APWbdDTpHlQQFbths3s5ezD6gIdibdRcSnFYv5w/tXAobusajk+PDy3l73G3ze9K4qw7N4fIiNcG
xGYPOjgpKLFI1sYY1VFcjN1v8GU/Bx1wuUSLgb/Rf2HjmESYR2MANQ9aDPFojKyxWGwBgBdukxgu
naO/CTzfpbR47WhSbVrI/QA5ErV/6lUX4T7ZFI6GPVEG3j/6FzE85iKYJXbK3zUNIOqKDU4KsOP7
HdgiAMHiVhf2M7jZuk4MurkF4cVSXrTAUgJ1YMrf5m+w19cDdh9m0sfR0gAjukGMpjlxes9cUg6u
qGAspv44Cbkz+3ErTvlj9vx2qG3iHBcxSPgmr0oDdFzajmmiD+IqlpvOodl4zQBVL5iRX5nS4JrS
kpDoExl7CybzOJNwe6Ai2K4Q2zbZ/GAyU4OJ9AA1l7e+eCCKoKVpZ4UnqwUxMCSwbXRkLOGf2tlN
q2uL4exHZwpyjlAUZxlA2vH8RG/mHdP6LtX0ECsH3d4CTsUzbdoVbqPzaWc3/bD9KLxV+ezISSgY
PO5hKBe7orvCb5fL9yGDlnKPqlb7PTyWXPucg4BPUr6UAK8MI9ODMT0CReWOQ6IW6DW2M3j0tPQQ
h+M8RM1lmWX+6R5FDSx46WKc3aqB4lCf8K0ivd2RWTIPVlzObiVhOhf7eHU4XDOYuwyxPJ3ygQLx
EI68o9zt86jWBd22WcgfI5UK0bwpQJ+ZsV7ba/4QDWFH657tn/FL+O7FTosJ5AMnTzB2YzgTMvRb
MjXRQ9IH+2wSNnzm5iKTDEgBwUPl+QImU5KQ6R36tJ8j+lZO752MjnzWPgEHPKq5MH71pDLpPGrN
xyeFE1aIWpqAM69b3op9+Ovluu9Cav4yElLhsc32JLKBAWL43MYV2sW7+y+igJazhdo+rcBISwQb
bEllMyE4/5TmrLY5VnTEznBjPdBQd9uPPhfK3wFXw7/L0VtvvUwAaN7yGN5AkuXfnp4OrGgy/379
WWlgFxGmQsEankNWflBTboMB1eg3UzflEmCF1wcLGImhhT5HPVG1XSGscZs41GKeJJLoWhEr6c6C
rf9GWx+j19rix735/gaSCO0kfse89DEYu771LgebqLidc6n/6QYOC/vIEYL+wTR3Bhc72RZv7jHd
p1/j06Uohj7h8YqUP0N7Zz6rEObWOt93yhReLNKtoRkjD2STPf32mUBUBMITtE6H1kzEcDTuIv/M
3f8AnLi6E0wVX4GURSu+mUBq7Ofla8tvIp33qyywopuZY7hDFnY40zEHSpVyEcjsEdeW+JLDbSPU
sZMSdPakm1Nr8vXWVhH8HnA3NOnPyR8y1P6GU/rZ7TON8GDb3sncmJofxgEsHxy8fVF5H6WyZhkt
7nAmByga0bE9AU/282bA04saOdRP2AqNCc0XeH1QKqmPNHprjXGVYX85JMxSe8x0eaCHNWzmKUur
tz+couKVsPwvL1W57PL3hxSdcEY76gkWbplF5puUhttd0m9xX8Y86wkjFIFbk62FzGh/KXRm+omE
m+hkl6fl3JDm7RGNrcB/QM8xg8qbWt2qqK3PJYcQCwuhCfA8fVuuFTiQeH4yxhOtL9PcaXCk5guT
7STpxABxZMJExW+z5Vfn0Huo6eN5+DmB8ykcHD5uEqI4t/Sddpu+m2xykl1WbmQ70V3d2eANSdMd
jhwj/wuxqIEXXZbWIsXjYxHBRtnJSbvt0ln3QTpgQhuioFat7UiLnGv/xlfzzj6Qaw5aQNp4mhO5
kbO/eGXcs5nGir43kaIzlT/uIpqMOaQetnqfDdNO29g51Nrd16ozVBCihNmYcuQPqO/pRD+sMKwV
0+bybOgs5t5ll92BM9AD7aDQ1BbHeTCDseIVFzu3isFIdshsD1mXqDEl73Kb42cXaCNoJOpxR6uT
Ox5qUa9YWdKiaLbyZ0T0/vJCXlT2s30EOFQqQ+CBGUarpkXi5JGmuq1+svp86kHvWlA1nYONA/UL
Zjyuko2OZsrGP3zMexXPO5+ZFOxvE/dAMke2y2sQ9ij57slpM11Mr2H5vOW4vDKsqYPYGutu+r90
EfxiJBZF6Xs+BO9eNz+eWsOG1LT+k11m+wUGjiOS+meeOhuG4CAiGt6HfmL0OgIVLuzWcLIBRjwN
CLul7BTlBkUneIJubdcGy2l8wEkRr9GQFln9FgEpAivCKEkyLukTdo8PVuU6u6TouRfS6g7TbnIv
3IbzEJvhxFSe+4UKVO3sPTQF+Y6DsbgTCI12rnRRIMeTMpNL/wvfGlRP7QXcH9dcECro9z/SNVhb
gpgW8myF0Cn0F+Oyhpgbx24GZiuYDZGxS8LVlbYqIBYHcA4lShLKA6qNHuhgPAtliPF8wP9ppWlQ
34NgE3vRcGk9Eo0xTPlE6bfH6L7f13HtyvfUB1NnDTKIzQAg+3ZtYkzx0+/UIt0E9DW5eE6ImsTE
mEDpNGz3CGz+Od0oBp0I5li/uXAjL4v2Ob5VRbj1pVRvX2u1R8qPzCw0zcq8zAY7GZB/U4qJFwzE
KoQK9hl/dUAlkusYqFGc/b1XYzHkDTe3dnNr9bk6+8lURgP65Hi7Ka2GmV/634RjiPSD6HrWeO/K
VFOvbWieqCxn2DpqrFx8RpXwkafIqLnwFN2gbPXcNEajtQNlFWI371YSQMuib6TTivP4UZ2dCZT1
8l3Wr1jYwqT5R31RtvLoU3OOT2rfkaaOYtCEpuViPkqZ1WFYn9JHT8Y3kO0+D6LBhQohf1gvMLF1
SAeWEoWQk90oBoKYnrYilKoo77B+89utyq63d0LFWI7Q1Civ1GvU9m65NHNkSQP2o2iULQyGDuVO
ENHHfr/6UqfTQdm0ltBM4EukfVjLCpJFx4hjOCIKzLnxUMnvTJZ2migtOF4Ns9qZg3a6qik/niOx
JZ2QX88I1DPdEgDh5oc7IU1IrcvCNZMzPudYPx/wR/utESWIFh+aA5MNwikN/8+tcZ7uWUU+/CXT
WvQC1Q4aKEp7Te/udH2U1mJ5K71iCM7fLaOwo7WaTU9pVxqk5llbNY6mEj2tPgQ/l1dtqmRab7LA
vv93ylU9xrJ5JAUm/H+DKr90r0V/edO/j0FKLmUdBU/B/8OENiXkvdiZgLWDr3Ls9gVuIWaYMzeF
g/Tt5F7QuUyMR+LmdIcBOctWTxwI7hETAWiHI387vAYMH2E2TQZgxBXlSaDxJt0n8nLDDWKkMbSS
4pBXukWuzpDOingnFDm8abG7tJw+5lcpzJLylZ8oaYA9axwcXSV1znNVi7zVvg8MxrxnzyLhBL6y
lTgOLPxwje3/ikCXlweKdxpZiAPH+CJi7Ab7D4VmmLQu1+p7wYLhD3sHlkwqRGjXdD+libdMW5wy
ox3KCRQqgBjVr8mGo2XhWUzKlga0sUX+rRPkCZ2p648mfjLGC4aT9BMg07jR9FKVoo8J+0ce6M2Y
AI6FHx0AL59VF58LHFbXcgpC+3ZxVDgwW71EAEwvOaH13PKH2CiCgjkJn0uaKnpalxLvTXGqu5eL
OXtPtLDZGnZIFypKcmc/CSF+dAWJZz1q3KbLbTSL2xZy4mAKdH7MIWXWX7Mgx1Ksk7euCWWrU+8Q
EKmfZtI1I2ruj+TTqH+Da83uK4I0hPI+58J2DwdAlafRHSuglAwjt9hK4dcaSAop70uE/YcogkXv
k2c1iRzl+6x50DURqg6ccrw+gkkfm+ofaFYpr9VN6zIknwYOZB1/Yx/sUu+WqghAJ7/kaEx/G97l
Yyeq1GVVE+xVMhJao+N0ZvQKjiKQNEsy3smLbvVO3/b/Isg9JiS1hreDBNU04v5oTc4ci7TDeM4D
LgzD0ougulbZSHU0VjJvOKv97GAdKrK4Fci1XuaGvK8I36agZ2/3Uy6PmdOgoFwfs6teRmLWxsc8
2TqiYWBxfFwCUxswOX05Nu3xnXIsRfi1X9apKVs5TECYOPnVHPNDtlQujNLrXhYZRPsJBgQ/o9yq
JbeCvo30A988JspoZ9Lne70uxiarl3aY/8XIzT6YTfYjf/tpIvlKSx3kwCOkl8ppLALv/vyduqoD
AQTrPPjK7stKw8AHEdWZqiMG//sqqfgBvbLeO6DpgB3fClU7oRDk+5BiX3TDBNM1ko3asx3wuDYY
QJ3RkpYIIE6HURAtA2DX9KapHXyqQFuEhfVWxVO7PeiZQ1T3Fjdz9bcbQdvVVs8l1TDfk10PVevH
22rj+5xEBdRaKtYDBB4l+qk6ds+6QLzcojTQ1KULC5KGj/o6CmdnLczis16MJqh/mz531CMemiYN
T6VoC/q1o3E52NwI1YoEV4Q9Va9jr5dD2lpeve4qC67W7k5Bk73DbOe4jwRd6csSkdkxV4D3WQ2R
VS7huHSToZSeoINXXbrmhdz5eFXZrvIhMXrA4dCfcjdB+dmJVkSiFeLzerhiv+sB1ir/ujs5/p0/
ZVJz0iFQooT0CW2oMjoYUaPOI7jugmslx6mpKCiwc/AYK8ogLly3C6mxr+0mGE56DNesMA5tc039
8dUDnysbu7azn+gtyFbiT22ph4wxPGPSWq5oY3CVkuYsBsS2FHa0gizWTuIS8TnnniCcYUP/0zyE
4f9eCPPwTllFOiQe0AlFzKoQEAiuIuRWskRapEVbofTj+CEgPsbRYaHyABjqzN8Cm0iL9re6Wvw7
pGXwxCMMpBPJKdDOdd1AGysg5SUNvyFozXGtqbQAw62ijbUPqvTeCPJHWtBIPAWfjOleLIl1yJ9O
HZXp4vt5gAxcOO/mlim2xPtF7EGTxagagSmIsFLVmxxxheuGGXdZ+6SSLPMc6RcLTFA4PoQ9yN6k
wciN8uCdwWoPANliWwGG37oIhX52oi8dr0bSzdMp2nuq1QSEWXd8SstE6zaKFzT6zyVXtnnsZi7h
OhnBjqmpDe+tGaspwTPIrH2RCoKaUmhDEUJEFTnpXyL5rE1VJestiBvhnZ6YRMJNmiANErElniHR
iNnzX9Vas6OVKdRcjYR+209WFV9NMgSss6iBbww1Y3SCYfDyMeoZCVufu0z2zRkXb9YKC1qE43W2
+vj7tZZ//uPsgNUPJuLp6wj4h84LCLwABcuDXQ+LI7gMFpKYbxsLV9jRgjaGNzjADfUnUFKgQUby
+BTQTXLk73if/8mcu6Vgnc1iS8Om0oe60B5cBbZaL7FIvZ7HCidv4skw8RQqPAr1KwQfl0qOR6UJ
So9Cke9a9pSLQPNx3YJAoWNFAhA47J39uKLmDspx4lP1LTUXlsj35eb1dI41/e5+rFJsPlzMC+18
8ZE2ha9VQ61EcfT6BWGrSIrhAdvOI1ew2QSYWWVFa+v74RECv0qLMr64XeXixh0Vabhzhptpy6HC
FrIUYFSeWXXqB39/UJIOh6X3cxl2gFjMrKG7tCDRCIxVwpYWuA3e5/sXIQ7QAh0viZqOmKHhiJPn
+d6dSdqw4tXEn8O3zrEeUrCHzUXeePXzUe1yVLc24ins4w2WRxzTRA3YRERnBS+Fns0oCHcJ/3Zw
5sw0pBw22W6+q1ogFbWeB03YvPxx0ZW7X2JkFoR+Zt2aOfyqsRR9vKJZ3MXEedTZhlOnVHMzNqIY
8ON3I9dZZTyKyzshW15Q1S2dH62da8TlDSHUlpkF3raruZ+cZiW5FqwWCbzvGPPYW83ND2skWYhy
gyCQbNneBpjlHnRiaVmu63KLbY8ql+yA1IehYlLHSoLQdKiu/cSoV6Ti0pMuy7tlUhDYOdRi8MUz
lKKGGbFRvkRQoMXb5HpvUnUZVVeSmeY0/Vda+GemGaKo4KEY5Mg9f1uPN9qzX78i6x76wlLZg7r2
+JIpMxTA/e3MUVA27O6bqmpUugZFzzAZNS1ogoPHEXk5enpe6RSRJ2yqROQ7BtaEfQd9e8vP2CbL
iyHKsQ1DsUog/p9KIxkxgUmroJw1Oj1zP6urSL/DRUh7UxeRffl275li93BweIGTBld3MC6ODhJ+
XCFh1hrqXmpoaTiLzlUf7nMSUDdJJ9XTpFOt8L9BYVrepQwa3qzjE3v1AIYcfnClS+9Xoh5KyB/Q
L4eBLOS+NrMRllBjy6uLybgfuyfJy7+YoueBtXjXDBUneseygl10eCUoMTCfVzi2WFF6GGRE/Eqp
/4rstNEKNknGw37nR6cAjooKCXXtSIgsjnS8DBOtoDFgh1X3KGuZ5OKAt8DJdDxCzWHDDaKNxG+9
MCLqw8oJ9CtZ8i0pfobaX/0YleXFU5mrjbRb1SPavcPzS+tIvcZvv9KhNTRUw/NmcLQBWCCgTNVp
RNyjzn3lD36LqR7GI1WDGpAFVcnm5UKMn7W+16Jhl7L7oFAUYReq4exub0h3lJAuzjgjsZc7/odh
zKm9Sb5ZgUbRIQjSt7jjRqgpbfXbIKl4XoTWIqGMURmwRllxmtsnTNOjIjVtYj8eljmxou4cyiLt
/By3qGtnHk+Myk2RLf7toPjW/cwNAI9DsWXNhByYWnSL9h11idz4ZbUkayvxUJgniMMqsYbKnLAd
MScTgZTMZrpPAkLSaxrCd5BdO4buposZEA7pQTnpSh/WXOxn8ncj8k9v2isYSbb6FZPwW6l0Y6OL
ELdpRqF18aJ6Uy7CjzcMh0Zf3p0dUVSzmKgIXvTOpjDhqig07oksrItfE3K8UzvYDLIfB7PIgOyF
78ey4R0c3fSB3tZjlB/qHyOWc1qGweyvwpB9OMA478JfjH7tTHewM9r49aryY/8buArwIXZ2xAuj
FXzSsPEnZqNy1IlWHX2/bat2c+J64A/zxoZgkEjm1GpBqYR/t4huxMwlnolrv0r7UX+MbfJ/MR/9
AQV8Z/ExzGVqYEobNh7/o2e/umRmCykRCx5m4VLBUCi0A3gaaqqMDv0XB8T9rIyO4wt6nkWeGmtg
+9Q3DDsSA3cqIwhx4PXEr0paD0tVdhozYuC/0x64qvCSaOpF1VDVojCG8/H8CKyz7tCmOVkRqjS6
UEmpGgJ0VhtEH6pqqGO3I+28h6Eqb14LWDzsTVB4KDpUWZnUoo7mYyFTfSsmo7o7wX/Qz4cep1zO
LD+CuOksTmR54abGjgRMeIIjIedHJeigM7Dxv9p8S/rCtHoC2VdOZW7fOQwagdI3bIxJWCkV9ZSJ
f4odNChj3zYE9PJd76FzjqEiVgFK+zBXHJmGqcexCgOxdjiicKzaT78iILPPC7cSyR7hTK9LB7iM
Y1FakD2LfhqrmfXj2W1X5MrtRSQjPOh7Ydgqh7JYCLEo1iijR2NUVhnsUjH4u50GPebkmLOtgWG7
MpTHpCSjijcE6CpHKykcRj8MpZXQT72bXYyfZ7l08v2XQ8uHEreMaH35nO5Pl/B8JbGPLqehbbQb
nly5+WD4gIHHSp65RtYiO+3Eh4AMfaSCIFvsI+VhOz6N0n2Z5iBw7mCkzQCCAc6p6t1L+meFOX/H
WxTrLhGe12NFpnTfWFiD/Cc1djIwaRHQrXUtYNHp3+aeB8QYrSp0pHUNWypMfuYBFk2b5VVBvuLd
EP7SgcDi0WdAbFOeDoLCoLcHjRvw0jF6wm6Hrmaz+Owkw9hmiBsiDAjTmjXgSC47WRtwBl+xy4s4
rtJZGlBCHzFUloZSWjswctVvXLRWkg7SLjx/AsXoUrq+x6mfRpvqyzz9mKkrTc0fSEmx9CxDyrCy
alY9tJpy6r6NWMIGuTaGrxjDMbkxE76j28JcTI9bA2jvm25ZHyurabKOT/F5j10ocZ/2E/XBy73n
P4E+O+M9Hjb13tikhGsV8oFvdJN6RDeTANPXxhP58RPWHG8Cfe2TitJfrNQYVZKUa1n0DhhRGlzx
91t+fFHtX67gbaIP33hClF1LFo5fnZTyHMgE0/5zwQe1yhDLQs5IJF9k4cwV8ZCjrX0G+6Eowpwp
MnOdPR8umeVatsRLLzO6Z9RfLZZKNad/9PISS8VNQ7TG8MISXnhgkVvxHiKZaMAcG6MWT+uV2pNM
DctZjkJW5RVAmJ4b9OV4hC6rYVko9S/Y00+rHTSowdsfxI1kqS5/smyHphC9cTkhFPqmRriRg1+d
+X2f1dPrF2RjZcdb0YrTmRaBkxosUUX6p9yxtPcDaQnkq2BU1gP37jIBbEbaw7MixrRSehiK+dqN
LK9jyPbthF5M0IfAXWfxCnIqm3jJmoVuWtKHgZlzN8R+aaD+R4ns+lKTaF9Y0SKX0tqt32gpdIVQ
INMvJ26LaX9G1gm8nAt/XxNH9yepzW0LncP0BVRFEVtUSzGNWZtl+ONXLqy23/OD71Gtx0Tl8zDy
gvEVHGc1eQ5Xr+OwojKqSCeoXdVeZUmbqwlid2DAlB7lbwZhhOO8FHZjU/Q5g7SM7nvtAWCn+lcJ
4GrMNdJUX8UAn/XAv+RyLdoW4wb0wiIvLOaQGgDbHPFS2iG4QV+8RRjmAiR/8CykwKOPRvgDY1yv
6B1WKRC0IP6xdwUj/E+K4EN+mdNfXAm/su0ujT1Em1icddyZxtYb73OoQB2pYJdAbBQgOwkUgESS
Vyoluu6W+4+nudI+z4Ra/Y6mgH6J9Hnx/exezy4WsojZNkPWWMJk0f1LWxjg7r2ZPLl6iY/6Az/C
qGDG8fPmVgWdUWFPOJQlkTYDOHuhECyUby8nFjzh/bsU6d/7+ZbQanklOlVQI6plUsNO27qd/mVc
XO+Ywasyw849AitSu/NjPsdA6KWh2GK5o51GW54TXnmETcNijNzhjJCU+KPn0MI9ArFZf63HLIkZ
I83bE6CSxPxvVoc5kdDduJrCy8kFjKCsFSATqriI4m6QI4ttnvGE+NqAbEvqNOBDmytdvr8BKJBk
kCN8o3njH3GTKGqeaBGOKkJiRJ2kzVqbUKKSdDYPtdf48itYuHmsxbN9PavuwxG0JshV2DJKt73q
XvzHSbkJKQ0qvE5i+taN1AoH8aUpEsU39WA4MJn1FogshsIf+O+/vdzmJVPEPQF04Yv5L3sRNTsL
kdT/LhSHAJTwoRN6aIcgelJ2VZh12WOnIA2X2vHl+lcwvm9f6UW6cuzbwGJNv3ekntdhP9ynhqRZ
z/qIYJZG4SJyzzUh5ZfhWvP9prdQ7MmgTgbua/AoVBg8YKmvntV9BoP+4i82Pytrgwoi3T2JNA9S
XaaHgHSAbON+emakqSs2vkSVu09z8o2mC41jDgjzWP0t+iF/gh6EJ7nq2T7RpvwfqGwTtAHaaWpL
lhhfN4Iv9kLvh2sUzPC+Ja8JuwHXOFSvWN/RacPn2GiuFu8vhDYNL5/b1PUSTET4/slUKKpe/CRt
/5eUJ1VXT8Or1PdrfXGghmnFE4l/LwLiRV09IuabKB4w3XKUcGEhf2ZYOg0PdaznpWaMdfxghD8y
HrcHh9do+ijYetIYoeB1XY2sTw9HHW/rCUu8GPuXdsTGl20d33atpKZza3nbx602RpW2IqeC4g/c
WI8lkypWv9iJiTOyJgRs5TmsoOawZzHzLqwhnKGVqaTzUTvwjuVQ21XAa4h3NvbDkbKln+VtDqh+
qR85GEMUczylbKX/wMzMfMCqhwzvn0wXnHcHLOslBMiKLtMvdfxqEG80HHKm7VwQcwjFJcPLF9nK
Flruok2WPFFeOqdw7T9jc2iGXxgW/LEg5zzhuj/CqaeqS+0MlAA2dKus3J14T1Pq/xkhkxqxxhje
Xf58CG1uvOUkb+d4sQQKGtZl8M7zBJA5DkWKH7G9isKwPj35eZY+0xGZ4utv2RBFsqoIvDCjpPb9
d66gTcp8uYUd6EKF+cqsHt/ScpTqxXGRrEvEnWSye4bbqtjL4qe8rB9bc7eepD8DIl8OnCj2OjjF
wnQIWcBxATHjnzgFEqKyvL0Y02ls9lWi+W26GGfLzWSkN3zyOlrxcSBUfmAfYqPtOARlLSZ6D+qw
RKNSMRmRyigV860OW5HRCcaafA77NDFyQwv9a516/FrvyeHBfJKN8uqfCpKK44yRdNIiAubbpoBD
9pqLwfATrltYU4VsOpqGQEZNkBeiTswFDhQ2o1gf0w8GB4/HgXzyx5zqHQlQQ0v7yEOZh/PZjzPY
vk4lnL8YLlQjjyhMHxSB9603IwfX0KqBVSXNUYJICk3lgcryTY/q7kRB6S5OQEdAIrVRSLKNHCg2
HgxsBBf/iKEzdeugfFc5f0imS5UHNgpsTRhh68pKEYSsXG7QEhukcWelXGU+6iLTdwf+I1VC1ScB
BLPLO0om8BzPnB71BKaqROyMhl4pzv0W0QvMmyylOm44IzCYK9BsXmzl1VYUovVOIYoR4t4nD6Ya
M0H6zwfw+J5YCf4PEOONwIlBn0//OnjamQvWjQvdRnMM/Hw7l2+roM7nKft2zNWRSxSMj4CNflTj
KTeuTAprWCeT3YREW+K86rPdm1ibJi025dK9RMxAuCx65e+SWw/Rkg0/G7chiLTJPJgh9ZX167UW
HeudY9LbC8um4BDXUZNzNua0ujWp3z58QKXMPmYb50NALa8WZISW4npe/wz0lHGO++EOjAdd0sxZ
O7RLMKO1fO/UMp2oDBIoQU6f1pdQBah7iB0l4iTKEUDFLpaVDVCWOAsedDFN/TUxczeOMr+jQJMb
d/w8S8nd+ulqmIoPvMQ5aAyzM3LxiBQ8ChjOoTeppIktXFcFU2hQ+rw8o1ySdbE/JJiAgOG+l5WH
o6NTUgbwnc/aG+3Va7X9jnC/eoIrTZ2hOnRUuH4S1B8T+ceDgm/F1/pkk5/oL2g1US7O+x0Txt2L
1XI5tE2B3rdXZqY0uW40ZrBn1QNKATR70dSASfzibbHwtUxRtpqKfLJHUsySUCKoH3FfhdYwwDVL
n+GVM3nL4hrj4z/Scklc0xEfIvf6IO75nRrExRysTnHs7hAy4yzPUKzYRn4piJszPic4W2MpVFc3
SqhZFiPRkrKPPH7IlaU4tkzUt/E2u2VW7u4jOiHXmmdAI8iX6+O2DVTSksgvyCn08uAbss7q7ubQ
FpzObB3SRWoIjvFC23KdfC2oibJR8HIdxmgE8DVljTgIh4j1N/XCxFQvp6HEkdqaNM+LcxE1rdrf
j/PdMUaQuVJsQbglOpbG2ZyYN/OCvqjDz7pn8+VdfiRRSs9gDCJe12NzX1UjGu0GQ+STRLQJiGEQ
Xy1UQnYqh+tRcav7Ew8uNHCdRm0bpMfBUFhG1m+/vF06EiC8g09bzJzlcidFRg7fHPOEFJZgCZxg
UwnWCgiqiyTJI9ES5b9QZ/kjY7DQoG9z03LPIeIak+RHEWLQlVF2mWKZRXkoacebQq6RrvfCWtO0
BpBhKSQO2zmxCESt3G80WTiGQ2FMnKJKxkkV1mxkdu1mNI1pz4ANt3WavA0OAAKOGgRKoy8SzU0F
EnO9HUzzBDo5tsMSQDP80DIXMcJAOtKudi6LxjKZ61zBEqWE/hoA0Z+mip9+0oraCaF3StLYjK0W
s+xUu3dpTKjqR0KX/z868D/paBImQTS3OW5yJfw0w+ehsKSOpjN43orvErKX6eRtD/Wq6LeXrWUh
3esWFda+Js4VgCG0avHgK7XlRVZfs5s4tB+ZM3U8MHvag/AwNtuv06r+TszQTzWF54Y5m90tuosv
wfa3oUfbu6OSxBzpso1QZCyLfuuhxIbXr33GpsewgfSgsIDCORuE2zCvl6GpVypAx8SrogvUVVjh
q5yfOYwhMTqCgYjU7/bzNm4b6F0fRgsolHLJJXkOBR+4VxuexLNsR0CimYS/Npp3yRwf6rXDx2T+
mWMbA52EnvSNJkVN3agdiGXPVflF5hIYqf7dpvGfrvTCN3SFmruCfHS979YJvWXoerOufNUydw7/
YYb/jbvcv4bTjBLdZsS4W08mpk8ipf3stmmGzx400HEHCgfRMkhLXaYhjpwwbcxlo6lqUKkHWUmQ
sWGirKOvVYqSkm3Z6IkdHuGBmlU5/WmVi7y/1ujUzNpP+RNqVc7O3QXakHksym+J8N9Ke8Y7dt6N
a9n+xrNIw/tuaW8Xfb9iXeISVABYgyBN3qGa9OGJwvX8PRMmkJc5dGytDzvCDhUX1wqWdw2UlnW9
dbKewFSRF3dbp+4bN1W9jTMbzc8jbFfi2A4Bo/6GJTiEFsL1qnr/4IrCbs0idElRxU0HiC5feZfF
YVn8Pas3MzF3jG6Na/63O2pKNZaM8AFH5OxplGsPd4WKzXsm7saRn2PfXLxGkiiAUQaeZigZDx7W
12kYZ02YhqNvdklw6ehnz5jKZqRR9yeC5r/Ox65v3LftViozLFxskSLEqSoMe30MMpC903HQ56sp
eoNE1o+cyUZOYZGG3SBF3SyQN0lTI2YZqvhnU3kdOvTTeacfThBmW3F2oBbeK68oiIjBrmXeGoxX
DDGXBODHAiXnuOqie3FpLd3t2iGxWCKLiGcpK+pBvSUjMfDyrLpphrw8Kzw6HfxTes7AmeArE29x
Wot9Irqa9mZGdakwREBoUGXOcfEK99Q+zraP/W9VQJw3mBRjDDta/tni6L6WJwBTv9pxNKWDWDNv
VC14ssjRXrvrGjXC0RNmBQVUBiRgLljd17aack8SGl+ubXsU95OvPj/AdQojIwnyF6VtMzm2WLJ9
sSCURQp7yKzu34lKX8yjY7E7/+cC475NRHYfzaAeBJ6wZtu+hk93CZ3UvZWhNOMbhx1QH/1MibWK
tfV9klZ9beshfkxjiFP3AEGh4idW40CFLOHiBCTN6Xx5i/Bq2MVO9ru5619/kCdv7rCQbSikCDI3
xt0JWDifl2mFVktiLWYZ1IXmz72KAMsnxef3PpBAKnA81GHjfmgF1NzpCfgHdvLqz5E8qmRqd8ms
n4jdv667+f3UwfnVhGK3I+oF71pYzCUmv6dqNpFcCsl6khGECEiM7d9eotOSrKIt04RHl1gt7QR0
4WaQqIQiInqFZf710jKlDwzv+1t/beFSZiuq//Fl/8w2aFU6jfhxuBrsgzaYUQq2nD6oyesFrn05
aWsIs1MkjMuQgIA/hnzuKKns2nm4d+bfLzMHVHKT7O1775r0tHkPQO1rdr0x9MCzknEdfWUWTpIX
D65NYApJZc8Sl+B5vSPTaH4J7ou8Tlf0Gn0x73WyipTnJoytdRaOygUOUB/XEJ3wtt4c/bqurqGo
e0G/kC7toBP855oWgwJnXPXy1i4/cgKj4AMiVwxoOaNO7RQwlDY3nSBPPtHknbLAZlMsJbv0qxEF
h6Ah3dtuG3VQdmgYfoajJ1hrNAczQ2fnPydQIP1Fkrteh8eNLef5IOzNvrRw7Ce/m9Tkq/uNjY7C
6WocO7nYXnBP2P3rfAUxyLj+/8GVu6HVJ6ga4gIiPEEY0cL96ruT/CEnI96CTTZSmAdapeVand9O
EfQ+w2x79kLkSy0bojiOQJ0S8qJUgmwbgNlqg8V9BHQekdXZUR5FN+5BnK/aGahg2H2x4zjHaWjK
vD4vM3GPN9Quc3ow1xTDbloYWXrGiMHFLNAxpW/AKfQ+swa4KKbi7V+iKtJt9e/b62+mU3uyRvUQ
rjMvYfTtxK0Rb6ZQn1X3wMXmytufuxcBwQlxBIYbV1H8an7NqYtEb7tCSOh+7rtfnNzoYdGlqDqz
+TWgCDaRd8DWkWedwtf2dNjHepm2hy95fSB2LGRtBym49TAfYf+JaU6PzPiN9+SYCJvfdcW77POr
g6Kz/y4exEjZAsPJCS755YIOW9dC7B5EOaLbgmu09ZE29VEjNZb4fDZVIBPO5lg5TgKyr1XMOtIg
03kz6Ps5yAajg7xUwO+L1kw751MqzPPuYLUnPdeLMxZ7rw6hrf06d5Uzj6hqdewgEdbNYCvOyz+q
QWj2fmtfgteP9dnNhdX/2pjTF/0Yzc5gVU4HD879mwCrdjEjElMozHkLvPT0zR/G575R+A3ricwx
Xif7/O54E5/t2xjRJ3YA2M3wG3WhXeLAQjAWY+RLKPvGDL5+urWawZ3QzuvulVZbi0LyZQuO/l8C
aZonOMISGIJi/fVEEyK/BESq0ITLq0fNfeoWKkQkj8oKrWZp+Zyb3jvu3zfPsasSGpawibeuDJ4g
PfzO9qGfADNxqlCRZz0b8efoGgY9BHb6/2p6FHngmKasHmenECSKid6zqCBvtRek/UcIK0yPVFYY
hRpSP2fLezZiqdiVA5Dvbu2BX9Mt1rMh2eJV8o7EDb4zqzb1d/l4ynusOGOOPi0kTy4PFbMU4W4q
bEWQjRyVYKEihMBkyzrUdseJ1UNsE6WToHgMY+VL6gczXnNRSsn9UKjhhHLthpB0egs+FhkQIbun
pvtNiPrxfdmhd6aMIrmNPzXsB2hHunNFT4WX3TJxQnbGoxWanQOurrusyttfSMSv8mM5I+4NBzVL
HIWoV+QDRiX3r1Jsw1gq+oLkJP56ov00/qPaDh/O6CTrFAfR5SbFVserL0+KHA0Et+IuqmTKGUZw
8+wdmvbr8sPVazVKC9JuXgtkB9M65vmUf5VYJCkt/nMwz7ZOZ+GSPnk+HQ32jdT60xS9mYy6T0/8
wKSPxbzPXVlkk2L0Vibeyvi3hBgsnKnPCs/mmiu2846XUbaUad7nj6JbBfNUs8KEtQf42yR4KtXU
yMTJK4MXJEmdLpxtot7vhd4TgoH0721n9M9vOQh5K/k2kFHjbdQYz//PG1xe/ZJXIQCIrVxfR02r
4MfRVhxzSsm85rQ8seFO4Tm3z7nLg94fBULsUDp/ha51kf81YQBQJsEVRI2jP6dzZl+zkfVqaKMb
Jqd2Qmolv9W8STVebvFpB3StJmsseTEDfXGEnUqXPBWJNm41AwopU/PFrJu76lJ0LzSUY6sLQh74
NZ9DcdYcAcYygFGvh/KES3mOky/M73weMg4i8SkD8VjFo68SW2t441HxuYKBAjn8jJhM+Ikw5xab
PRbnLDcAdH0LVhEmw+/82RSXliRsSNg8i2RMTDkVlBlsKKkXVZXYioqB/TIvd/anWsHQvzYEFXrd
QJEB+dwqrBxRjq64scq3Ndl+J1AHEM7+jYLEbQEWCa33dK2HBHHEcrKXEnmiFbeGYgGJvOadkmWv
wuvNYIUlH2j6QhDkEojFLZxAen20QX9g47h1aKiEIzkZT4QUys2JXD3Tky2eQuQA37rOlZ5FAMrS
PwYeQYQSDhy2o0r2usRyFVQIvvJGQ03qPpSiZONeWPG9+HkmbPkao8wiToKMrcAk2du09COiR8dI
6bnblxb/rEgnAQnyPtI6ruZahBC0ESjsRol+VDl/N6q3mb8/iD22Gv1mMXfREjG9DONnPLjnpHXD
Z0s8KcBksdyMD+yXikAml/BHn9Pmn4PdqoOBCp3dKnjP8BRdSO8fofB0sp+lwAiOkNWENs2XUCr3
CPiq8/XyMI3EqdBfOxUOfSV/8nRQhR1u7+e6mYK12onqKr8hQ/ycm+oOESUGNA7qS+XP09Dwkb4G
EH2ROqxYqywc5RPiDkE/1SEu/7y5Lc72J3WTZOxVL14bLSPKV19U6ZthSMvz3Ns/Ojhdz5rE4s+W
3A0FMsUijwRcGoKes9pq7g6uWz0+s+AKYX0JlcOAMr6g4yAL06cfQQ4mWGh3EjcuOq6fQxKuDsTv
SUTUi5FDmqsfHWMD2q+8ovxZEp7HZUk1ygyF72bzGe+mG1M/2JrLF5oBHvDiR8V0R1w4RVUd0e+s
MibTgrcres9Wovgc8VNKKgp9gHJLq0r5KWJf1oCsbxDHp6qQ99sF1hCaunXcXsdbe4e1Nou77nwd
q8OrxiWv3ZgBlCTJfGs0WecImJHwenqHUtQY4RyXRbnoJzIGbramtwCZt1slvuaRsE04qqrKmEyU
SvBKIsfKMfnHYGroLwBFm1bz4wGhDMaj7b5Peq8FEpUFsQODKsOq97Pucs5hzX6B/6NJHH6oHdT/
iO6mupolPxFWifCWBYhKeW+9S16yzHk7w1hqeOtTaLCxx5oYVwmBmCaJc9rK7xpJ0m9YNde3tIjQ
PmKGaaTbiFdBCWA5O1YBLConPCPNMD8eguqZ9CTFQJAXQmRaW29HQRKd5vo+AEncOCQljdF9n1WU
KCjTPsq9Jd25P4UV80PZ5RC3CAp1JmtUkw/lb6ivsZ7B1WJZRnpWkfPUTPageq21d7ml1HWxnCVx
nP57PYQKIEoKpHKpe4wpPuI/eaJ4wNS7PtZ0vK/3kZDkrc0XHOROwkRscRDtaxLahUPPkyPIvLK0
JkQKSNfgFrSEknXQaTJZoRUy5yjltFwr7gAvhpe8vWl1sO8rT8rKAwvm0hjHjWhITPjYAq7cY53s
PBj6gG92D6IbF2o6lpbixTFrcktJRtomcmh0tAbrgX/wiIIS0Nl5CfJy6sNRk4D78GVaEFbbXqR4
n+QHd7sJfG4vtmhwI0M7hdDY8QVc/PZficaQHzHmgNz3fq8S42HJb7U1jFepFK8s4N9fZc+bmmcn
JVfO7bhkk1/OjTkD3pPWJv+0SNAtiYItmv9YFu/w98h1OzmRs0LPGchuaAkzTYbCLAifa/qe8nTs
IqzIBlzha9DO4zksgHbIKplQOF171BmarfMXTIGq+OD1uppxdbZoAPP76/ypolFgTyLrCtV4vyKR
Yn5N24ULhuvT5V8OjxLByGcrOCxVsghJbJWNK6sj+hancsIo19K37Jmvzv9VEV7gJ2PztD/Rg644
TuhckGcOI7IrIzHADJxGMyTHItGHmpLMISAnonDp6OWegYIW8kfVRHpy1/RRm/bSFrzPU3GYSjNA
f2C52TX/+oO4mOXzrXeWhnXyZHXhvkTOZYM4ggECR6YKTVPcRe9rtixY6eEm+4TgFYHuJPoMcoX9
sVv5cgWiNMwbiZ2kuAUOLYVnDhcZLZFRIxasgIvLLy/alniX27XjiCAYkGY4ZENe7Wztf+F5kYdq
ZiLQn6JhIbxl1yTVwEAzxRmiuOMWx0dCBvRhcCHD3VMeMN+BCWGVG6kOO5tRuvRB5W9Edqvswk/v
Os9jfExK5wlZIsgNR672Qi6aqGvddBlnXOOTonW5hKVe866iGENwZN9TeYcl/M+wU/BE+MXb6n8u
mxT0bfIVudb/a9vs6JUqIgmZGbz6OjpH4vEm01cOzsZBa8QIKTOtpZZPoRyrEv8GIeUnpmOT8JQH
4Rqw5thq5XH9afMhtI3gJudT/Uof7XF/U3YkqI5qHAfetB2qfXf5dUs8XwJVVh7C3qTzrzrIO+ay
RnRUW3k9BRwiNGANkyPGTNzuZBV14MTVZzhxtB16yd5FKpiki2y2FKWqGo+IIOr/ctEJeqOKInXi
Voqux0sw4YtNwSBm5TRz5yIWaR1ZX0qhQ3KG2m/edQj5w0ZPQ16JevtcozqgREOXrpfQ+yT41YVd
ueSoQrfkMg+WY4HPuq1G6Pzy1599mB13LNVYCV0n4qhBfTZw9pGTNwUafcgDt5NOntJYq4omk9K1
CRzNJjF4X+Et/AaAGIEcONhPEjcrKZQy6D37wDZA6Xczz5VF/rhmokxTj/gULRYiSORr3mB084gm
QP04ZnRYyh90CheEjG4KhJ5gv09XtNBQJEb8QQfv3NdMNnmWnIXd9x+QoxVNYtk055JcgNfa+DOo
Ae3b39IZxS1LiEmoT7jeL61lYOe9pvHUtvOmV8rOrDz9vZPn/JXILTkTFEu+skiT3WAuyMv7sYdS
7P4KOFmVZ0ejpakzP164wZdWOPj/bYUm2KZZVKUKIjU79eBa6YNQtg8QFcSZGxqViJbK/av77bR2
MisR1YukESWMapTGNdaLzJR7PvN8neQbNeGeHk6/8+EdCM7HVa6YpXdfwkDzpLzHJDVIQmA8lPUU
2HN7CtJPSq9g33kJ+F83mUTi7JKEZ1LQlu31zzqC7qxkg2xsiPH5kpku8hJxiQwSG+r2tHGiEWat
X4dTDBo+FyRrwLkt6UckfCFb4zF3S8dThC6+1vNh6r3JCsS2IDY+dw4G4XleNIi7adrbHRe5LZGB
LwhefcUEnufaXy7a7jfSMe6QjLgPd+yF7MITcqK2liHDB/891pnYri+WfBIaUBIcyLVOVVqqovvq
PMPTEn653REuI2Tb5OpNDAIyWqap7UbKJdmvIEC6pxjd3/CHMkfMgGXfopj6i2Vq3U9kncU9wSRv
z199tnfdXMPHYOOclnauWd4OfWNC+9qBxZDMitgBEamIo4nLXL+ZZd5IVahkW4sxqcp3ARAtmieS
KX26OeZKdJbOYX3ObsTwkQWlIAIG+NZaA+GgiE7qoO5pmxNvTVx8hX3YO4fRoEomKHZiloYQvAyu
qTwaZv3y/GJ6mZUDI4ma6d0ObOD9GITs7eWAG7NbHse3t01R8GR/TiZcIJ7m/rMvGk4iNM19taza
xA0/kfr5iHfQYBDxVj/SWLDTSOmr9ofZYgI5QtHVPJNjGvEKVR96hqeLZPe5al9dlNDuqsxsev7q
8MzKdYshD9/Wzn5i4nd6YEFNJ+TcuLOCdwSkd7bKGOyd1in1GFwdcWhzIrkY8k1puoqK0wq//eRl
SUlGQ6i6SZNOsmJP5GrUeF5Ldl4tTFIR+ggG00RC3OHeSWGlRF8Dkg2JsMTWHSyWNrhi6pEyloTY
F1KFr8BxCstxlUyps2+Wn+reo0OChf0ljeeMWlpE2YAHbOI0g4t3+arAn98Q3zWz0pvElXYLtPSk
vDMf+hQlM7D+KIk69kZYmhqv1f1zsFkbz3LRgJTxBw3BD1uDccFDAc54pogcXpG6htTZ2SN6qrOS
dq13C7N5W7vwUDnLWA345K1QYx8JB6PLS34yeLTGcBRVyPhPr0+tffqeVRIxUuQu6F1cy2kfGzMa
HIPSXQlPKXRH83oQI+AXPuwAX13TUW1TGQttQRRcB17rSNfZYlS7md3VsKfNpxr0Q0lNowZYF//J
tzE1gngU/6yw7CqVaQgntTgE3oUxihuNlOI83Vz9Bxx5AZwYgGY1u3N8rs4U6JK3JpM99z0mRP8W
XkjafpvBOzbUVjDviNXdNPoh7B+cfTNU1T2B+Ln27h5WPNLsKb0AC1Es9nxZzA2Ik1fhOwSYGB7q
1h5OYZnJRVrS1s4qyKfNuQQ5PqAl5X3oxNIE4n1h01is9OpUQnNzPqU4U+D/gqpMevZXw+GAETMo
AgHzbv9iCwKcaci3Pom9eu4Yiv6kZY6C5ZYTTuFLrIJD02yE4xVkwc/9WHpzg2WBipbPfHK/INCL
GY1MiBiPWpPGm1lWDah3ds9ocll5HSe7cSDmYDtshXdItyLB2plNi1FtkUrJtOZqf+uN+vLJ0Odu
9unCnf1Q0b369SFaTn2Eh1NH/TCFjHUwiIRlLbAAMQ0HHL7Aea3karbEdrHHTkVY/hhkUEj5K4fZ
ljni1wrjQvHwKPr+fMFN1DlGflbJTtEaCRByPaX/Lg0ODyy8RR3mkRUxNPfuglCmEv9EJfmQIXvl
YY2rnjK/PvGnnByXpLArrAtpGcUzOwBbFMCoUr4tf41wLeWUdv8MTknGPCma/ZL6EkuU/xKJXL6d
CZd9DJbsaGxmcdRgFhmzxPVT/LExlK03oOJT1B7J/x4efUhS2N647/WWR/WvDXHjf/4rFh6e0sfd
NGaH5x6Swm2U2GfgD6mvK82MCo7G+0q1jZxxHaq+5PCy61GW+heMLDXk3vBwgz9b8zpVhAaUN0ME
9/EK52v4J1CscVNrBy1bSbIvvXYjNQnD1LKRhjW3AXUc8rH5m2Ax1ikeyQcKnp4maOlSSSJsW2sj
xE/bnfZ7O6CmxFErOKN/jkwAviuqA9u8mL4JHTVvFHXLm4zpA/rFwVTAY7dcdzjIUCV/8mPhhFCG
xSleHG64MW+FWCArFPw0aVX43/TfPiaxZNShbWv1d3ex506nxt4SzDRHN+RnLofrXb4sxI8ilJoe
CRvlWkStWHASMnp9mxvFsdOcjNy1vJ5JtEiEXxEGD8iAwcwCOdVSTRrTEULxMwdPc3WfB069tg+I
ObL/31eiO/WYA2kkvet6Q/bRT/NYwvlBJCOnM5+5tgrVF57JBe00HlMzbiPfRYwFAEJT68uR8H3Q
P1/bXo5ZxBvCqa8aZhPews+KNTY/q6PbkdDnbfAnPfyrVJcqzz1Ar2AF+HkEicYC3qFIzqRFNHUr
KR85QuGR67mm8hsq+zKmRexTIv+fZ48fzyAAsVBcJpJO8Re4cNQC4+mxFqmlBXBA/zl8XR6lNbz1
9MgiWPxbve3JPu6eKDRtaoQSGsVrw+Kkj2A1I43psm6eQuaMguO6jHh6EQy4ZpJSbtlWSJNM4hIo
br6gBNrW4e559lx/pfxZI5JvpDW3bQaV2qYXbY2nmWReMi5wd80j+8sEt+TRu7xkG1MSvnlrUasr
B+2CXzajs5hnovYpWVxSQqKp1dUeHcN78bb+X5SlFCEHDVlqontaUwE3UOhOKhcxcxeKe4Wrc/9y
U/9Xx+KpLYD27rj8NWoyovqfQN7udSqRS4pY5WmMOvnh/ALnI/90qkvOBV2wzu/2mOSuZHC/oaan
T7EXUXKBtDjJOSjWrP64/m7+HfIh8XNccq8s3YN2cbBh7OX36OGktpeBnlx8Hfmw1BGwM22qZUAA
o7D9wov7UK71c4ZkwwXfg+hdJoKpX/NlfMvNarZel2IKXQJQCBaOVrvePlVCp1RaWAreLLuXAww/
mWaaKc0iK+daubKCSpNGKClClauEG+54Kxg1thel3GRXSc3tLJntd4Dh/VTpCEO0mfBA6MxXPL7R
rUvugqfr6gDddMTmX1WZwnGjdZavwn937N0XC8e4QAwR7Upc8J76Ql5hbP1dBtKlfewdsTzpk13u
cfblMPoJyUUSHCmfAmQ32k43UszpBQ1WAGEXuakBsWkF1KTLhC/RxxWvbDDxICIYF7rZWlVBdMoX
TokR7oQXxx7TqXkMnKeQlZnX7mx5k2BE3eto4y4Zdx/L6dAJyjlzmH8fwt5K2WAeAZLVKqJjouVv
E7kyKdc0GjD13SQ2A57TVcNn2/Y2cfdVSQCebMDVMea+udGCtvWJ+Gd5hoxioLMafPjdG/xAr1Ip
BQr89QZitsx+aClUW80xb2qnoOSS2jViT2bLg37nS3IGzNinJpbC7JDsKKAfBKCma/TYvNxaVz/G
HH+Xpi7JIHYfspT4n0qlrDBI4gHZojPlpSs7rjLxjhjIOdcz8UohKyjuXAxtzfJ8WscnvBO2OeBO
ygW9VI/s8rSxq9qlko+VWdRwDIiPjTjejO2zAkXYYOOAf1ksUW3gdJzd+E714cIGTcO+igLekZjD
H3epcXc0nDx7rGGSLHU9jfX+qZXdRVc3tyXNZoLxUL3sMRJl1NE8/aYfnXfRL603koyNVq58VGNY
sIXbXLFMjwid4YCc0ZAgl0NMdso5OwbOaauhj/3uALmnvyUyuijqSNB473BNyppCgiTbzXP9HlKf
bUulbRfUphi8A+omovNZ2jy9bQoYftw/AcczkvMJ5HwHkCH3L+H6YUmQFLYeO1dozg/pbW0DxsRY
XZvteQoSSbuGY+4Jj1hFomTaX0c+3mEJJMgnVtrXNJUKnVngLPZFj1NN1gNR9WvhycjwoFJtTCAF
rS1XM4Mmhlzm1krzausLyNf/5Xy3YEFjv2UjuilE/VDurim6thwsaaHjL+N8EOZGZnpVpaaybI20
WBwa24zM7fi6eAK13oDMM0yAfCTB6PNudQkNKcQnr6KnmvAs/4eEQhf6gf7hb54s2ekUYPXPH/5u
dWRB92zM6WL4187RtKQhVgG/1Cpy5+blOpqpMD5r3/BCnraKMkakTZTxxt3mZnMEXKtMPSuGz3uw
JKVIyJJ1dgG/C2bvIYhGiPEbbsyUdxEDbRdX/hWVZh8GcIKFZ9yiRvXJQ2PuFI68rT5aARhsyfUE
o6dHjgRO0PCtnphRUkflVgcJZ2Q/DYJb8Ja7GSvnJLIPcn/hMUjDG/8xxcrae2TGWWfcpot3vguK
9yQwGt1kPUvhVnGiEOSLkbBt2EqI8zOxlyPWAehE9iiZWpcEjaSNYsnEEc631HltCP27wPidtfCy
3o3QIE9/GKTqZApeVR2kEtA2SLKEkQjK4lYlf8w/1vvz5tQV8PEeWkHJFJ8CSLsFGlZKnSYKY6ro
QOT89Df5LoW8MFJj6FSbkK1ke9qYURSTqnyl/ZyvIN0Y9eTPQ9nrjrIMaj10CCCBPGhTYIavxNN/
h5OtGAfVVbHR8wgEuei/sUQyf8s5uxTMnPQF3wFTphxC0aQY+xSG8lNtTS3Wdg8CFCZSRbhGwodR
Ey4AM9LKV1rq4az+i25KSU8nlUsIKHt3rvTNjXtBQFOYL+mMkxhEuAoU89mBCtPT3ISWoC0cT72+
/ret8k8hmKyFfO+vN3vyGh8yHdFvNH/S4/De+ztIOdewcCOY4dh3oMfzu0NPQjF0QSsa0xqy9MSr
SiVo8BxQLUrxaic2Vr6e4ZyWE5SVuMYvs295+chHW802oI/lwi3oeUN2WSlVL4B7KlqE3npsjwgT
vNMED1rPz5Zt6fVl0DqX8J+2u8YRMdAef0iD3LH110iWJRJBy8lIPtaqIQimGqkXKFrb2ga/vPeb
UWbzzHsXD0E5BfFvTnc/N9p6Jix5iaEsEhHtZgB068fP8L5erIwxby0Cw1fKqyFCzgH+YmKl+CMM
aXXl/LlcEQ/XJ5VDT1lbqH5wXbZgqWhU42wYcf2rG8u3xgNyGJODWov7jC0jrNfYl/bicR4tQlvf
s+DWDnvDIyKT0sSJGb9Y3iuDlSJoQaBsWweoTBKP5vYsNs3ULTXAkSqXqk3rzpzgQklvhODHLXJ3
iLzRQuTqRWzuGWb6qsh8O+FRChYccLzxj7wHoN7pd5DUhsp3SMuVNuYw7i+uuaGsu7nu3SG0q0aW
5R0AkKvO41KX2kDyw9ABkScKTvduEO43qbPwC5l6eMmty1DcRKlDYldUponFPiZv2kW92vOSqGdH
iFzGe/8a26sPXefcHUvBHpH4e/gC2avQmihmIBWxdaCy/8gbSVS+tYaRp9t/T4FWiSMBdmQ4Q0Dz
Lv04Hhl8duL+JL2s4glhjPCtg4hQk/nUafSEBDYbmRzQ3SAEWg85fhF0W0b0ikIc4sl7ytMXdZBq
yiauv4dspHieGmTwgEBiZ71e0stdTskBHFY60O7k0k6NCZRIkaHRDtHcsU5rAOY5vcV/9zvxmKjO
UVsZWsd8lVfdoD45V+O1dpAMZZN4h2ESGu1xGE2JyhhT3VUGWlvqhxGr1G924M9Wf5C5WJ3KTc6S
bGYm9U/nd5AemV8rNMJhxn/WRSe7b4wYPm9gmuy4tC0aw5iOtCsDJMLFxjUHoIIhJQr479bJwRoV
vfm53Bvtiyu7+SGyTFgl2VJvgXX8FqVuWb6wceX4mcgaPHJtI7ynSUK6iydeA53dAyO8UW2FEXf6
2qP0Y4wCUqWK0gXVzg8LcPMABvAJ9FThf2BanJLDl/cWrVpKdmUBkce3Y9Pf6+0WU4Y20BstIAME
1+xt7ys11xmA9jxOknaqt17NvhpiZaVUluNKLLnGB3C5sYCQf/JEDhtO01UDME1d7EE4grFb2lVa
EEUySQmEZXRgxOCCYFzm0LMy3eOgn9qCrtE8Rw+fSPx8FHEmrAWVjXL1vpzkQQllxvBVznEr9Uya
WKMHUfLt72e6jlAD68PbjjSU4b/dIizuGlcMVOUzGdHXwx/CxvRjxsTzHAdNVcenagjY2MpJO9u9
KHFGiY+mLWgBTrMPHmRkFgSov987OmjQ2qiSl0fwTPX9puvskieeIOgbxMQRGLrcW+LjiZ62xo4p
yYhwB7YEa3cJeVs1aZDijulUPNpeELdxqbC6s6Rcu/iwXMQaJgVhV6tns1I9jklRC/36WJ/PEXwv
KE/XXnpT3Lz5K4ELTxeB+n2WLcSC0APXpO3dbZmfDZorHd4pYy1gyoDTmegeHAWE6ymT4jbOshFd
bz0MrinCuBzmI6S6Aj2HzjLQWBipHnVO6Cr8DITtV6jRbhxfG2MOCbTZ4/rj9vAJAWa6+NjBL0dR
2NEUVT/ebvPnqIGAC5hICk++NJ4+aSm7yxHFu7L4lEk2keAMfGjpiAubYmnHlsiWoQjFzvWlWw/X
q+f/51AspRStnagx6aB0trr8qSZASTlYvPu7yaGEAeYroObq40x8tGwj0SKDOlWYGpCopPcXsLih
8II7BYX0sF1wT9mlRD5EuqPX5+V0kyo+uh88bafJEIlBNDkk7aM4I2rBiZ7oOJiur8wy2h0GEUAh
b8NHdrImwkD0lqHtjlplna2zulAf90GOWI6SQ7RTL/pL82+rOQk5ujBibpsUOFMJHBm+lv1fyv9W
rXTilOmWQ5/6CDUon10N90+skxzkuS8qjO4PgHVvoN9x5tMoGBbTTmOrZyLXgEEUgDhHCiDQPA1f
zvvS/7lDgzbSXGp1hD4N+dWVSmgY1fTuvKU8Gmy4ZgQ08H0tpgzFMfaq6S6NJylTAo2VLSEt3CQA
mQJxl4ZP8VfL4nA/jDQ7ajzCi2lUJ14M/zRfq+F1AB7Enx8TRCU2u+AAIvAWvNcyvScrqtv8QT3W
PphCfvzBQo80/PCoGQ6BRDZbm2q2Uf/KlNzx779xzHdfef7yuVIVQgOWFwCEV/7Qu0JcREnLBFux
dxhkEzmbefhqbras2fGi32zyq05eJKQb/n+17iobWjoemevG+xUcAnCCeznmrrprwFif17yA4z+2
Cc76LMQHUGsu9S9UGnKgxBlcIFDrIeNv2NFkdvZWp4Hd6Y2lkJFn4A0Bp6QWMH0rzZwGrlC9a2P2
T11pjzuM8UPiYZDrAS/nBwZEN/D7isxGHV8SSU/fkDyvWDjmDuQhGb2miDJdeMPjWx7alHOtjVn3
j4ytgK+0D1q0MP5wjUUNH1XW/3DvNjcEcinhKyfECaGyby/OIYo3KyOJdqmSIec8n16bfagH0VCC
sJ2NTu6S2EZpg2Vp8ivdjj0z51lNtKmIGujegRFAhmRPmeMQiG1KwUUkEfpTNJXd/fTcTfCPYlYx
pSRCfwmnkGbuJuxmdqMIM9yNBD82MDtstCxtiIOFY9TGwxFhRqUSK3kpmCVa5zmcwjTF8gyyem5t
LagjhnT2HmpPHTxZVzClXLe3NNdOUZ88QcXNVPdVQvIzI70l0HpHuqdYISJujNcq7cMLDghUCPm2
zLgCbbQGxlEcSKptRETTmWiDxzisYzjTtYrdm2nyfGJnpJriq7BmpwocxLw7J701roHqGyosiH7l
OzGBuOUofjmHy7ANaVNpEA2+S5v/vENi9JBEu4cDYSohsMtn+njDUpJ8qmdcpkYIaP/jOxzk7Scu
fshzayrv8o4R+J3focbLvmNC/T5VMC60Jfr/xYcSZfxK2rxndP/Fmr3qWTZj8M1XEWsxhGhIDe4f
MerWYXL1LB/3tk0MuCtOSbsFwx2IdtYbszzNXFZ8P5oDSb5/s7s9yrb3d4C//3/2d1/nSday9uSn
zseDj+VRq5bStiW1UXXwxj8w880v8tyLBgQ8o23LN66v1BoorJ9RIRi5csAC1I55SUVXkZfTP3Wd
dU1LS7HMmId5RRtACQLeSgwNb8dhZTQtPZtbdDe8KBkWWwUy0Uy70kzYTXyf+EQxKqpr+Jimb/Nt
eFXeZXunDPrdsxP9zlz0HLiyjb3Xi/uQ4m8xFjnPee1WWfFlXebK/qg+8/8f6TwzaYnNP6cWYJqu
z1FKd4Qm0M48DLxDA4HWHIrcpaawjfYHFlpN2Amj6MIGd6jZs6I1F4ONzWeiHnmWeXN5mTx10u1I
aiQRcuY9Pjqcyxa67y5yJ8tuZsE0bsg0/y5EgD4g2X8LZN3qEEkbh8wDTuCbH7BJwYDnkEBMuk25
/HhjgX1CLEst/A0M84e9XULT6OBJHRNpIbxBg/IgQ6OFGMzIs7D8HZk6kYSGaRijFD2Q2ubXClsr
5kqHOgwBHXVjelFq3B7gehlqerD8Mbe82AQRIpGD4P6v6xRXU6M4Zg3ud3213vwoRUvmJGMg1voa
/9SiI+j41loGSE3qTApqpIs/u8t8yhuc/iWRBIXA6uzBrvP2OP2RFUb1DsLzWh8NwFDBxxcZycfr
A/e6mEunslDYSBjI+cpudrBGknFVL6ZNRdd413hVNGQGi4ipj09qTE+0SZRywkt4WXFRVndU8jyY
5XMmrfbuzDW5byDBQzUbYlII97EzCHGngr2qoscRdx+7lspzeLEDZqjE3m9784flD28MMa28kkLj
tbDk+wQgmD3R6BgK1L1INghU2/1qqQbn0aOVVoPECmhLRq12+DP2cTdZrPxB999kuVx5fuNr6SqI
0iIpKpbh3tT5X4rL9643PLtc/jApY3Um9FNKVvGRWnLFfdO8WxSu7rCMs6X6xHJa2lfqT1Z2jnKc
6ITZGVTmiUgP2T/8TkzflzQ7DmbHq1BIn1LYbBI8MWqF3UT3grcAKbHRp+B37I9CtBaOqyk5jb2I
EYDLzAWhjreVEvH7LBpqHZnFXygLSMRBQyDjMxeGQdxbM+UYk3OfVPns3wuHM/h9f8hGfKrP1YZu
xdpJFlHu3kbQzzgc4PNFrUqYlLsrddCMm1TmgndixliN/NJ9gNdRUrd7NWJKnAYxo11+iDYv/AWR
iKtBrtms0dj7ol3iNhfxSUpvRLcsRsnQMpqIIK6xKq0R9Piyk3pu1iO1gX6sbIeUZLzZHBJZh+Ll
9dSO6a+2nRbweo03hzbPxVfnFeXxZs1uZLcGsTdHE3qsKspFsfJ6VsM1E88MsoYQKY82LUUmEy05
JR7rsyhgiqdAehR2RbLq497Q9rRAjaHvaRUwLY0S2FPfS7ET7a6fgUo0aXpfVEDCbxidsLd91ucW
vGwJBs9GbOfULkHrW/oQNMgwu7ZYl0W0vYdpeVb+djhKvxSjLlmGVZuUyhL0pgosmIVHpkPTdnLL
eFCApcBVml5avGRl6X93ozFUgmct9+LbZBBvRy0xBvMkwhVkpfU8/UtGgxfSL9MYaUH+F+abK1OA
sltxRNu3Vb0pDEAEJBuADGBdodw6U03wl3NfZ35Mg85Gp8E0LtjZz2mlpFhsVSOgBUdLGAQW98Th
KZkOFfGJnH5Ile7fybeR3JVe+qqALEpNXnmQi77MUI6Z1VCw55wz8Flts7GLxA5Ka2vfwTMkv3H/
2aJwuZgQI1IinD2mLjZBy2ssCvxXlz9X4AuuwPizHbKFszCwyLI+2M/qHTVbXp/fV+EFE3BbgthM
bzfhPCTa0IXQDl3lmDk2IMEV3CZd4JWLuZg98pJ1jNm3OM2LHGPpbFr4CV89NvFYKcdDGsAcgMrh
3YuCr1lYN/xlp4HqpZF1RWPhETKwCAaj7vHVTFwiLYnnIgcN4vd5tlYo9dDFAco15wlcV3BU0hIm
nBIM+9pq9T/SOdiRlsvzKUdP4hiYXZ6nc9UUZriN29p7fjHSiQT+A0w6n5gmRBXd6633htkCQQjf
zD/oJrmeNQnxx2UYoBFTYGstI3XvzoifDG+N22643r8zUWjVAHqeR2GOo20jQ5dUPai28puoUHUU
6wOHEsxVBKkawd6FJ+u7fZy+8S9lWS72SFfq9kSHOYxFQgBDeliEO2BnCm0bF5uraj6QEKASTXtk
u8Ibd3HpgDWUwpVvc9e7mRBJjYn7h1RrTAYRJtjMlRpsWob+Y0gLkQ2oyMgFLmkq6EYYEky4+WLp
JzVl+2sf23PoDwnlVQKTMSpW7ySZ74hGaET0lBO5no47yKFaKKsU/i8D0nA6+oM33g2O+yzedBoL
0hGthy/9zm4snVhrk+Um77y3AIvhKEUxma2Sg0q1T74DELzcFjuffGDkrpo5xTLfNQy7m5aItNaw
21O1xbf071d8PRbu/qYOI3kwVuosnnoARMqBr9TB1LthBLoYbcM/Qn81nX+QXa1EEBNE8vDs3xiB
0A8T2Uz3vREA+7avCgRyXzb2ufQUIMcek6TU1KydY4h0C9A3l6a0gUu0D9m3397UtAwVcQPMgX0V
CjnKpJm2iUYNOdvQjBJng1pSRvbvuxw1tH0wsK609XtswN48GDJKLYsnWZC9gIHYejD7M4i/hmk4
j33lBqQL55bmd/xUBaHmKfjznDMRyai18JyN4ULZOH9BVsyTluzU6cBTp5Pdhu96mLKJ26hh00pT
78J1v7H9Bm3FaEXS0ZFvLoMaJ9lebZY9TDkYSXvmJvDxJvDL+uvUIMzg27tC0pYh0wq0keEVnFw3
y4giKZqZMdh35bQgiwEp5hvSsN4ZO0CjNtaNo/qbsxGuWnzwoz2I3CDLNPRVKGWbx67uH7xjzDOJ
nJrlIDNOlcsgS1Ix814++DqbqBjYp9/rYwZPA6B8ycwDVV2zzqhJ8LiLJ+XlMnVt3BMmZEImVPda
QGgPT38s2k652i5bcJJ8JnQVpD5RnfD5TBeVcobjoPYW3Yxydi4XZniDgyIlu5+/jGvHeE6p2eC8
mT0QXcws/4JEYuqcdL4uW78roUDBr3Rb1gX95YPh8YCPWdybhbgTJPJWmk2G/B1eYf9RdlFr9QqB
LM6B4aHabUUfQUWpQVzmRlQ5viUdaXC7SQJjAljFY27CNL0QZ+v8LFSF8MQUd+LSO113C5bbsPtq
5gMl6P1Y2Dh9N9iN8yCByuduGNulJQ7NxT+onSZeaPKa5GUeWloQ9+ev0cZuvzESoVozvCZActJF
vRLVUFc5KdxyYkx542S99d17gIliAVsIyp2BLBPk8ZQ84Bd/gzrBIya4qRt8b7w7U1f76wbX6OEH
e1T35V+X7TfpBXeZ2J5ZJEFfDn8DKnyqyxYUfIhAeYE/DPUytIPlkfqtnjxd6gIDB4hSp/qYZxB3
wyoIGsxcFRUZtuAG4CQRaUCFhMgdZR2NYEDP650QeZnqErJhlUEQhtYOXSOBoAx6uImbTTtD8R0h
FUrsSW3UOCJPnYiVivM1gkw5d3w7wEQwqy9rQlL+CMCj3Pms9dfzNOge7LQPGtp+ZIMKDNKGgXcy
UyzFw8ceXOYsRuhUM8ZdEJVth0n9Y+ExzLjWZCls+7M2uBZHmPqKRmwa/LQ0SVExCYo6LlMz34+3
E2o151qB804YVJRdxQmnxIwjU/3HOzT973H/gf2Vti0yPiYEzdnusut+rO+4KqmIcS7pMC9T7WhJ
fTcK5/CocbngtV36+BL06vExeU7T6R4kv9/cm39Bu0ghcAeRQip2IeSOZX8nDZccD6LADdrwkza5
PZtwKr/eu/gGyU3DN0qdmQXyHGIPDZmJsKjJEOp5SyMm1z5v+XmnT4+XmxgmMvWcSX1bcQg2zXGJ
f7Jf7BmPdgVoWMDQfg+aNvtaXoOkUG1St1uuC7zRDPpujhNWdq8LrRL3AxVV5JiwvtuKFEzhiwAW
h717ysOH2s03PPXiSo2rxudiMLWlLwQ0AbnEq+0T7iUwOkIst1rd9FKB1NkoucKQweyfSvnPcd97
FNW1yX/Jw5V3kfTIDDObntBb9ddOxxcA/UsE9flhhc0HASGqfT/WqMcs4QioOPLb/P49xctZQ9Sq
XLmmhD48/90y3ZpU2XBuU6hJhlQFT4CPfuiHgRRAwxdx5kgA/wSuviJNw0cRU6T7aToshjWB1qvS
i4xHZFRvcpuJi066OCioLdC3jgC3LxFFEZ2PESgoK+9hjmWK7Lk/BNnmxyqHw9wCXGuE9dHn+ipf
TWA26gSn3JkR5Aza3U6czIJqGV0i7TLkIxkJ8CXEOU3GSjl0GpENGLhtnpANcoCG3TvFy/spC39Q
n5nUgL8Qr2BkKVDWINlLv+vwQVEQYtrbub66k7x50bKY/tafIB0TG8SfntKicWnXwEmUQchOOu84
MqofMM3CGVfBb9m44Nr1E6QKj+f24R0uMYLtSdFnX39xbI1x8SomY5tSa3vhuTvq/ZljQ74IgLZF
2t29pZq0/zq9kQhoPf4ygLUaL95pg8QofeDs8KDE2sahxQP1Laf2c1QJGpXvm0G/la30UW/tQS8Y
VbBY1m0O9zRxyUsgkMQoJidv6buoFHqpouFQVw1gBNcwmk/OW5gJePz+JTv4/Yb1uE33emPLqcLZ
ccxuVm49jnJ5qIYn9JPDctjmw8lxdiddkxIYVvt6CfqToTef03aHL4f5ZAs6HNuEv8CE8H5mZdmg
0U+vD2bXxLVI+ugy9hO8t/VFy1/CKBLToiRdKzDo8K5555+2yFAxV8UVMjEyyt9ntTixIah6we2o
tWnXsZLSpg/XoovSTZ2HsryWO5NhzHlgrfYLokXMcq9KK4L0ausUWGv2BuIHHEKxKKn2dYUp6HAW
ecym5cGeNrKWQW4Q+lqhINVxxBi+gPe0N3MCguhbSPTK/Ot9z3fLI8mJFj6XCcCLngN4BAEsPhW9
GNKV1rMzaR2NTeI1dExQgQbX7UcGh0XgJ9y0OItV8CcJkuilVG3fyXiOAxcub5bFNMX5/OyoRnD+
DgPLEk76udzePMJA5fgBFQiofUFXxbnudaklm/SzU4xfx58alGcUWLHDwzyqsslxz9DvyVI6PW8R
DzGEahm5UC2661N24gKFHLIFKL/veCcChMLkirU2+bFmvjXzrrye9qRLNhSsF9mE9bThyhvBms4m
3zMvhiAToGrNVCAEzHor4WA9XUjCOgnUY64lOprRzBKxulmpEmH0aAQjcH5XKp6DI1lMmjUNik0u
KWKr+nVwixgZhiq9/6+rz/J7C9kb6/aKXhl+k7WN6RBNJ70+UZj6nK8V5vmkpN3YPHecLjs+JVzr
w/bJ5xrPaR8PD21jM477mX/oXOkzdQkorArvX1La8zN4eZmfAnOGNDOmCazVHaTbAlhKuMJevBvl
+9Q9P+loz9/a/c5FGbqRb+cVFNLfh8mwV7TCnWNCyb5OBFjXCKGq7VB8g4WjwbMoKZGMm0YDTsRj
1+VD+6jmNFdtx4axpKsBJpX5h2Rd/seTSrE6wnLi3NPsd4STbZcaX0rRc/yyMzdTXcqb88wypIRf
Zlq+T9mt1xWakbLhXsTNjGZ25+cRkuf2yGeF8q9UtA/EsERplPkSi5ar2HMM4b6RC8iA5zwFSZmD
HR+JLscJqo/oDdHf3aKcLqnmAG7f4ir37kngZ7z9je/xkqsnyBTj3sEk92hhytLMReFXFYxc518g
IJlCO/UfhZij5dQ9T7wOMHGJzy7AqcbhA9bLc+SlYZTVlKB7i+D/k4pclEgrhzebz5Bjr1m7o25g
JNNUg7p38izcWy/18iEkSOlGE3cGamTAcNmN/CyDtSqghnWzywVo30KMJjQ7/NaowJxeXrIJToHw
x41xLa/yw/iioCjFr21MD09ulMjZmqHGec7w9Fch36tpktk4lov5qPFktoiRo6guvDL7M7YFhH8T
HjLENEn5C0sdc8HA0lkCLlepRQTz5q6CCOmOy/WijKf6KeMN/elHW4b/xvX9uq9ef5I+g8iehagu
SJZ4yLrWiHXIJO0/rX6x2IwalS4mb2Jbqeb+d3BD8msz7igEMukllcbMMX6UtqnH/Rzam4glqean
A6MIUnnwVAwexmkl6Oewh5KAHxiScc9CiadQBz5HL+6VSpi5OViuV2AGkVYCNRPXwN0oOC7sY/R/
2M4PS42BwedB9M7SG60+iA4Is05wjyNDHJwwoDRPeJ7kEY+kgNH4kc5R450EDb3ZHUUxsMatGT2s
QF7vCfD8aBdzYb4NgT0YBRKd/4MXkOi/YpcdD/685W/ORv4gysTbrP2q7BDOso6YFh67ZV2il318
QDJyO3AKezMdN4MndsAF5wBpWLtF8DgWpOLdFSbGGKd3TkEGjBnl2GhsM0yO/9cMrfXruv1ifNSf
5Akp1zeknHT4GtDTKcJY8TZxpcIH1CXlRfvs359b7l5fLrneykIXNedTbHOU1Z3EA4UAkI2YVkgj
K6T51yzejch2gMUJ66ZhF7mPY41QRk+JtNutkgp/EqF6afm+pn2bROIU5kwS7EsE6OYp9CxlCsKH
1QHhJFYKCoajWKmxtFqDqHo3owQSMqybwZL3x8YSK8P4Qst6C8yBs707DAf3WKQGGf0hoEVOekkT
P5FmGhiOstNWnmuh3ujQUq+wQrpZUwCal64f+1KyStSh/UPBupty2hL23VGp552jv3tBhlqJV4Yp
DVFvhaHOQKE0LbkwjtUNkELbqmXzitnJPVEDDAkv7ev+TqU/DMdTQPR3uKGxMfSja1bjiR4kvFjN
MrP+D5XFik47HMzyFudSPBGyYqTIAF7ILpRzcHRxkA97In+0tMVeQZPp7DHpDSWq9yOFubWGBrL5
4ksVhcIisk0vOTY4310+XGk2hnd6SyxHZOPDIHEeP1WmAHOgqOLfV25kzvY1tQyBrpPus/HT3ALS
h6rKJOYPBow7EZW2zz9Y41BShqRvfcSjUM7U2oyeGU9QMYDc6Ij7d+5NMoD5ZEflTA4hwEJkgJyj
ep9VOP9rn7Vp+gjyzmpwZVCjIcxBZDQ5SBzz45URqvClkJnrxx1yGHZiQaKPznyUA2QSScM7GQCM
QZWbxVFpCs8h9jG/fqLymu6+ObVRUU3spqIW/I+1+U/JwDZpIP3APQfPZ2+8iKqTw+XDLXb1XaAW
NwyqwRKQkQJ41iviwXBuI/cU0v0JrSnWmFlIe+Ef1PKl9Bz3Vr0HODBoT4n2eecJaU8dCXhHLlki
nF+0vNpgnZXukJfZ6QN5bOC/ORcaU8usHUswyOwOpKTmBPz2iCtxGiFMjYwsex7RpSaAwpX8XBvW
zstbsgzL/H/80j2Ncn4uZgEJ7dJco+bBuFGRQJik5jiJ7PBQSTVsNh1JAJSsm8EU41r6HkxC4Ac3
XAidPIPWE0egQiR+cDdIuL0cpVygSCHWR8JlbEXkA1/oYYzbzEi8EKm9UgErNq54KorkvaE3rJL/
/2zDsRD0lgstl5mjHBwXJlDpZCw5icWZNVuPM+SMVgGRYmjxMBiFXFMuCjLBdX9VPQWFVltfaqwF
j4QXpn/mvFsMbnEixtZuog04L/zJONYVP0k6gjGL3Xx6i/viq9y8vYs8P47kswZKCfHv+onxjQgO
PfC5fJCkByGcvKGJdAWTOVlZiLEOdOlnl4NbkN3RzbVPcrMNgbNQqUpfo6DhYfy9T3vqp984YvAj
ZlQWLAbUdedXcXyrjzIdwssk/C/CeotGp5Bcv7VvFOAo/9Gdu6wEMo4VvQRG5u0uE5FTxnNnMkd0
2cYcVPwLWXx2ZcnktIMvsihuo7c/3S37xAiv8bE6Wi9IITA1DjkEgqZKSLNIGo9heEd9AJNFlR2S
DZEf9Tb0FQBb5iQx0HAOeVKGTxpkR0ivtKIKQDcJl+RX6+He6bKzuNjmLOTUmwCkaEv+ye4X8CnN
W5uaQWmgvsgVvOMjvxkrxg4dSbjJAdT9msWe4tt2wdYMaGhmSR98yCnsWA38WAs1abp3pmytRcmq
Qib2EohVyOY26ViwiJFCTmgyXbfKt2ih08WAMfklMkY/71oGGZoWtHDoGnspkA+CsWGjiOOogqIH
AbbiR1C1CNU6WADrazgPCHxDL8Co+cwyG/YQUJsWMVcECsY9r5MTJZnzL41hzrEOHROUZ8GDHry1
twbqvLIc9C8jDrVMn9xJNlJa8JR0KFn0eZUi0GfFOcwg+tCLEHX92+FuhILWHVmTIydDvrePm0gc
mHaKG+Tj+pQxjmauwHwnBppRkg18XUXtdc2YO3jDjJ8U5B0rq3GgXuIXBV1Wpm1ORx3cuJO+NKgU
c6ThjbiVXWHRReYGddSgiceb01OTNtyQF4yFhIYofgkvz09K02fFHArdLB/ftHgJ4Z6AZm4M4rbi
p7Nwpb+coY/FgIbi/r67RLPUnwxiIAzbs8UDLgmYtrpiTXU1eOP3IWNLlZtMcopXWJQY5JGsRMNd
u5Hy981NG8PbaFC7mSYM4pJUbcjDmk6vTBm5lr2oBAedEAnmIduXb9AFqzPqOjeI2p4mTG5Ltjjn
/1ssSMGrQHShI2K/v4BnGeYM+s8Vz+HJksD5TqhOvlUmFLXw16jtCXLnp8av6NUhdFjdQCMHDUZO
5G3nm3pvBfDWbs/JmRdYaxEDtfrohykPQAxTUi1EPZM8Gzfg+DcE88HtXwMM6EPEQi4u1hTrZh8p
gSlq/ykPPE6PrTGgHFHKgV4K9SejmoLEZ3h0xpSlxSNXlbYsAlETYTpaZeIVOtCA4vU2rt1wwFqW
GH+v6PqOMhrJSeLvS7Oc4f+2209PpIHLv3XFH4Bz9f4rsdDwEWRAyJudSgoxiKtAx57JeflJxUbS
Qq1su6eEQFkcXoixWRIdDWtD+8LexeXMR+iwW6IkO/NGqu7r+YLroOtnX7PDhU7lsuWuuGb0Zajj
dYwhst7sm8qep/WltnILI37dUs9AzYSYGq8kOh+ZSlUY1r53o34zTGlbQ3aa7NKWApGoyHNQpwRN
aZ1AiSdFcb8NNuNrayZP0QB6G+HErLuuxIzsbcFbcxWclzQM7Sw1yVcFDw6a3y5ZziwK8LYfkREn
OfNVMIsxJYZMJyYnT98zWP5dSPzu7GdwvMbrkZtwoxqb3oBHpfhNZZTA13j4VKi+UoVC27fbQCRn
jAuU2MNkgIBJS6p/Xf6idPZXofSPZUXF/w2+piSYNHuIjSHNtVT+gNtQmlrEZ7+gkHrkHmdDDklo
Y/y9cSMg3VfHc4KNiPLoSB9MhCJuDtKcPZewSXdqHknQiRX/NGE6esgth9+PI+1QeVRn0hRnPBn5
sn6SEIi7i+5YiwZB8RTRfhEWpX8qR0/IltpqlXPtBwSregZgaINIAsG2GXJYnAFApH/fs5gpuux5
K5mloIM7aTJHve/nTpdcpoOanq7FSR2l5GAK1ShalASKvbBIR3PVKxLwkOpNW1AVI3jxXsI3XDY5
TuTo9i5tV4G43kET4d1MQj0jXKFAZE6D06pOnEM8YE7xKHQkKJigiKwzRPMHWaUJ6sqPYJAUKgMl
0rDKbPpdR1F8BtketoUGCXrlcCmjnDj1VoeX9hBGZlpFuURS43ITh2zipNxmsexbClzHq+72wHR6
0XcxUztVW4CqlJfdUBdOBLwdTt6Gx1aXzEjjt2XtI14QI0NYouqFkmWdvRj0B991rxTUv1x6AvbU
7JW93Fme0F1Te1UMTO74E7uUuMciMSwim7ksQG1RCOi2YH2xTBlSNgCDgR6IZGQa84zA67YOKQ/h
H7znARuYWfyodMZtHgjfkLdoVAytvmXchLQ3jrveMso7r074npj63a0BbCZBoNKQNS7Fd1dH/zIw
G6GNEhZ1v1Ilx3S8S02ZGAi7uZAo+11ksBaiH1vCbhKFLUxAHfrcXFCpX3lfe+kq/rA5VZ+qCYw/
YuL6N2rPXCr80QC5EvSL6CqqTfvFUnRiaPKMQZaOcQi+Shu5Z+zPGD//nnwwr4Ar8OItTW71p80K
2EfhukLDkZAVC4vVX5e7TwNS6A6AX9MGOFtDwleoXk6V3ArEQ++6ehMf7RAwHtKk9XppcvQdnE3K
o8r2auN1iLapUVh+2KQ4ABupDJIgpFfRoGDHPdjcvpkZrmRo9MOHD3UEn072K5xKd8iYRNA/1IIe
Tju1FE6vjwnKo8+UE/0672BDTvcMWnQG1f91VlU02bk3aXyFLis+Nn4SaLxXJbiLpJmvVYRtPRB6
QOMPxFWGbiZsKCvg2WZNovZd7FRkfuCY+O+k2tc9xXOiVOgRkIM2aRgELOtqynIesDtXC3kf/htG
cxym/XplNriJIdZnNLPRQgVqa9lFdj7/OD7/YYlqYoocSEOJ0wvNzXgoBHXLkPB3JNxrdjzfFf59
5zFvAcAIac6OsEBJ/p3/3yf1TC2eFXwOoghP6w+1xYtxTwp7Fe4ZzRC/4oblml2OUFJhstG4dGxb
sJEgdrRKDpm0KT6sEzx4rPML/4uxo8dh8yPljh34QRBCrOgAEAFYDhY/ceL6Y+bkTz9S8bLxfIxV
RIB73iJ/re0JoQDryclgVz8Po/9u6swQ7HOoUaOulb13PhPPVocp4oDf3nsNBZ9aeaaPm32aWqK7
Yfty4L+oM/0eJ9V28uoacj7avjzsBDNQikgTlNMhDECM1fnXvr0RELeYmeyFBCGGrc1au0h1dTJq
vUiJexuDw7TaGlz8SCXNp80D3OnhhVa/Dnzqa7gg2NqrdbswB8hVduM4nbBUHaqr7CG0C8sj3d5o
dnx7/URssIa02C3hDsy9ayzS1vPafeMcxS5/B5cyQqZR6SosJ7E7F/49ZFa/NhYQt0hjUkWITmnM
wZ68p8PS3gDPRedCQX4NkMPbQT10cqtOcEt+LN3Hj3faiCkbqyPcwuWKM1JOgjXV9VdM7Un3iUHI
RxFAVqccokfEYVmC6MGFeVdNddqm8luV2490eBPYaMZ57OzEw7YhS10dF3UB0madDVH3pIvHExKN
oHrZM6koTypUi0hMwbUa2IMb5Q6YPPMssYz4I9WBO9jXTAIpVbPEXkX/4vyyeFeyVnxSaaihFS+n
D1O03/YaY9YHZuIPAzDErpjYD/a+O/wRIq6seLAtIQvJk4nMAodeq830vT4DVfE14RlAF6BNLo9g
OXsy8doJtD4xyviDOPkJT+/xJvc5UWt7b6CJD0MJVrK8xIoLTgLKG0T4OLmNo53ZjKIPfqr9kE43
seUlfsEXM2Re6DMO1wL78evz8dTKnSMlLWSn/byU8N0H/xN/kuqWkixTgAIUlUO440tw7SYBw/Br
iguy45WG+k+RDrsDj3JNSm/9WshH+y6xEVG4mJ8PikZhwOsU9PzGk4ROOKl3T0FWVOS+bGa66p9W
7ueSTSHzFUMvWDl/K0kNeaIzRZWoNnh46nCGsChJQMM3BiWUn5JHUEZpXiJ/uK1+xLo7kWY4J/LE
eZT1YCROHh/BcvAtXO+P4eg57uApMgboep9III3Rfi4NriwQwPI+pX8P3s19BkOR0HzX/kNLXuVD
NYHTBPtwH+Fo54GrrS8xCclvxN+PZ8YVovp5ONjy3yD08BW7gTDitzg5xaVZVGwpafdQ0ksEvwi8
HfyquxdrElw0YF3lSSo/w75+ZkDnM9JYaxj5ycKWsQJgQ8iIL4btnVvXmCFWsC9VQWiRTSVdg7jv
RMKGBoM6JVnb7yDG/pWwAvVTz8/4xdM4oCE26uSap5A4sp7Rqgqrq74jn6x2cq3B+v2bFudTkMnt
0liVQKpOOKHJdInUeqSK6511R1vCgbi2gMPUpKd+jIsaE0dQrsBqnDY6r4jLTkPk4huLahS3I3MD
ax0Ifre+3su3yTjXTZ7EZYsjPTZdngxh8ihabr2dB9scS1/o+JOv2Sb675Dfm5POKHSUVk6bScWH
iZAmtJ3wvrXHIC2pxSkSVuNQQgTxJF94z+3EfTcz3H6iUYWKKsv63MvqSbTIawe06jyeQKM8++3X
43fRTeexA03r4OXAbGsAjDCx4p3E/mAmVV1WXQYFRFpWAjCaEN5CJpeHEGm0Z7bj3TCqF/1uz3ZV
/c3xXZc3bRfXZifElPqRV5DuloLj5/DOwC/nSd3wZ6mXtN8mGnCJ9kf1j+W6TDM5rn2QFJ7E5l7E
uXdCkl8KCYBWwqVT/ziXEcrvC1ya1n2qz8HZte/oJgdyCJXfaAbbMA9MuE+jcXmDG26xyHR+h5A0
Qdej4dybFxzV3jbHHbs5NxoA24fwimX30cGgNMcPRn3FIZEOLwOKpcFgen2dmo5KmbrM2zq2gXWV
E2i++Ip/Gf6wF7MVY2NUsdWfG/1LNej7isSB6beY8RP+r2yYUieMXAZA0IxnDMfV1qbK75ColxZ/
+npteSVHSwZju0TmQDDBneuVyj1SvWZjXho9M+VvOwgbTL75Z/x0O/LxnZ2YzlGBGw5DgxbX5SvR
vrfB9nDfu96teXFst3pcTX3DaD877zQAtn8WGjMf07sbrZo2t2XTNBWFW4Cw4BdTDLKPSaESwjDP
VXfo101ykwTquw7z6JSWnJz/Wx8Ayj4fP1H8lW3meAS59uvyEpPGgGGsrSdDt99S+jD41MpiGwfu
jYHvVHOYHIyjro+xxMPrdYtnG4IvIQR+R3GTji8A+UpMnyrDBMxfoNElBtExoMqBjCE2nta8p1+k
w6OocSAHFQ/P4htx9yNdD2LSTGTh151w3VNGQnK0fARepufcxhM1+XuSTsLYEnM9w3gBtWaIUbAy
QxzYGpH+wiwz1vCO99ceRSxkmMMLsxMzb+aEERa9g42e/HzRPBmQkv+KAriC9iKRx6TuQe0YqSut
UARwCCiIqNUywabhefG6TkawR/pesrA4QN8+jOImO2eN7gLVW5am8uoMGWCvtowSyZVn2uaMexwL
P0dh3xxaZtf8qeS+fF+2o5wuotY70nRlJHkXv1C/Sz+01vChqCYEbg7QDxDHALU3+PgGXtpJBqkT
/Jz2uQlO4yBaNRIsT3t7SErZGytX7ZXIh6qqLNwswE4Asoi2M0XoWQFCnHhKLYliw0ZahbMnQBMI
HJXab1JsY9qroSnbG9g10erFEgOicVftrRmKMWbevMY/QqC6c6rWzqYmwz6x4LB49mS+/sQ3ssEX
WgoGx8DZKHvSP26zwKUJNOOLnjJDRna4XU0ViMgpQ6kdn39psik3oe3e2lH10KqRaGt3pD8OYA5s
35Ub2G8MOr2FI9X+P8d3TWb++T7yAEwnjiGNC01GrZSiFAePw/9kzb7EfjtdgMSO6uQjEAnZ94wj
J6n1mfWkD0PbSlcJUDvSzV2mTLicrhVrfkx1UjojNujeqHIUEwv1gviOA87tKPpjxeQKZz7xQ6rk
4BEksMvaUkqA6B7lKS3SVW/T+/rgoU1ugnfherFwRNcbMMaL8PcD/9b5Xnr/358GB7684/MbVytg
ETj1wFZ39fM5uMM5e+tfuyRNfWk8y+VsfKIenLYfB0nAkrhiLTe8y66pG15uRIMDmZG+B/YaoxRr
vFwHNQM6pONbSDMUrhQfUBc72tdaRHLdBpbtv8EIF/WZlepIoFcJtcr895AsEMSpck3v4FnPqF1m
RFuemdZPMMcb9zafYQwknJjFbNFpnDkk9pLAcjGfLGcx5apv8/SgBKykR1RfDiMX0GItleaQeuI2
yUmMDVZmeh0ehQWoftTmurwkBDESMeJNxSm1tmPHbpWjgVuZLzoJ+iaOoK8tg/sUUoIHqLv/oDjI
36O1hhaG9QhRvjvgWb8FFrAGs1baGBiMo3KAqujaAAo/v8wHd4DRtgaXFccG+FI+39tiaFb8mmSp
wVHVkh8yzLKUMPNwQRWbaOkU4jkkRiSpquY3G6cR7olDw8ZGU77DN3D52oyuGwFDBKfznxMlVkt3
FKmEx8KvO+5GJlXqlmQq52z34zarGl9AVsHR4dtrUEr/Py8CudQgKJXe78AsX+HWnwBwGRz+VzxD
Qt3jMtQmhZMV1sNQLcUbDwGqlQYrTe4R2ZgKB6WLMYdQ7Q8OhuNDkKDD2i3DRKrIB26D9SgGRQn3
c3rEQX/0irHRtDoCb4HXTbMyRTWmp5GzLsarWOpZ9vLHdqjQha0aoE+bB/nloUjnpXnP2OLCswBz
u2rs2eIfvo81KmZEGMV/Cf/rLcShiIFTVel9epcILNXsJqz02T3erQOLjmV/hvewzP0qJYFX/nO0
1/eKvzHYkCwDQqahFlo8nXnfLjisNOxG4Yvr3UWOgiwnAatYsh60/0mDihwlZJTlqJhe663LwVdu
x/ZpjBin91JFfE3Uu6V4ETCdFLg/SAK8eVSTAlKyi4ByEW9bTFjAOAaUCviF3L5GXIXBuAqwJfF7
3TitJVoskblYnHmtmEs66dfCuDPvyjKdJewwIUp7qcJwauSx3kQdbpCwz4IcppT7mQUfi8JEYtw0
ghsfKwzEeDUupi0KsZZlY4XRMr8lulx6qusKn9AcP/jfuB1PEtdiE6kTiZ2xtDar8NbywCM/Fn7b
Hpg1F4KFoDE2dra3Oz9AsXnlP5ZbMJ6bjC/c044flPieOCcm4VvSnTI+FRTJCosUmLfRdB2GeK4p
99Sp20PSDGheZ1psl78bYDBA+W8LXC2si/Pbvfg0VOTvOY+o9QSDVOMlFg6QuX3mADeIFDQPYGjp
VXCl+fiuf3QDk7L5UtogBXQt1fm3yVt2JT5ZNYeisEIf5S1NAwD/Ri+EZ16YVSpgD3+lJCkTAN6u
FCSbfsUSBkfvZY20P/tQWtvLRWX/GWVHlQv0hPDvDLOiRWfJ7/sd0Z1GF1Z3uNHyGQ3jHSXZOU2F
2jRtwGOy3grJYMvjvn0O/5PTkdOND9uxzyGMGui7FLo8ZP3Xd+sLSIZ5qfPs9BnrHsEPUiM01Ffo
ivDH3plBUwpKGERPw5BpLimObDlepVFGdxYPoWS+3rg8u90ZdItR17gBbxgCqncC6LKGP2hRCiKe
6QUTuuAwDkDSzPwP700Jz0SZlLHwB8TF9LKSSyeJLi/LWP3KhahY6dlKRdcT9GXFZUFjO93wFRMw
IlVPFACYWrJtcCWutcKm5Y0Z9032gIPicsHPIYGj2ndIq+xAEpwbMiGo2zmvDV6kMFw8Md7chk8A
WqaOouoW+N5fcC3f4Mp0eIWCXKeFkYnIVyU2Kmq0BllXroNMrNlwXKHdvYCKMDhGTXb1wwp3Gdn/
GWepsRqOElDm2Kj9JoLeLOW2/5L2dN/+BpJXA8WLI99+2KW3OBzvri/3mUjNL1c+6TbPMUNmF6bo
X2T2sKueYdebYn6aP7cdk6685jmneC6s4uSFXJZbs1SvHxbYpAne+NaM4W6whgowRs0Ic4DjfMyt
TgdFdBSbDR2kXZSpZXN3ZGYWvspYyZLz1GaoTD/gHc3CsIbZkzGR4welWx7IVQO0RozjTvaC/H3o
m+q+uuwa4VYA9TxQdGoY5Y8MQ6ULQrcAKL+9ylCvsIJX5GRXV1UcPL4Vc9vsLTmvPONIpuujxFJu
9q/KOFARxM61UObsGxthKVUaZ8i3zOeMiYuuORxtcFd4y0fjzfAtivLZt+0y5hmsoIBY3pq1mUOo
pppb8EfByEmg/wD1fVDCps7JIWgg7OuxbnlghlImbjSasUKK2B6RMfdFCY+9HqswB7jhr7BW1RFX
dtdRt6PCUInsnN6NjvWX5G5S1ttxT/ZF+xqRH6lFM2qm0dysOr6NJTVq7v1oU/s6qNF/bBP8uLYF
zcuWMKTP7R1Gn/ZED/TosccCRZ/rYb9V++msobFqrdWgNGEvgxgPATtsKSxBa3jJT8bnC1YYUDB1
pyfFrN3C6DuRfcVUd/skkKSaerkzYwhvEiE2ZWGRGTQLVYMEY83ePEFUh1FcZ8iYEwwWN77VJdCj
gOaaGjRlDMvzw3YFe9HOgzn8IEEwjwZFBbl/tVuQHuXLdOouCRKjJFSxxZNWNWEDC7omlc2FJ0Nq
xIHIl20nLwRk4FBAlzHc81n1C1XLcTK8dq5l6YCCpJjCIX3QbTOaGXP0XyCbEK5czmi/D/hEiFGy
4XlNoKM8hqD8jH6Pi3C4q6moq2reB0qppnuycuFPQHc+HuZ+fYTQWvCTkJoq9K/azh+oa8LDE93f
mEVijgrOABMC8QkmAVyUFpUOQVn47n6kGqcYk2LO1+3GP3soOAFpACdV740RDFA6dRUO1Jyazj3E
ic63mvA8eTjKqNxLL8WwofvJ76kpbbdkB2jFpyXrRiO4k1qH19iewQgIRZWOicGHJvHJV5FtPrix
4zu3Q1p3O833mhZEfEu4AbYu2/pQCuaGFh3w59rsP6ivi7rp6tOnAo7MBEVqm9VVRheGABUqm2JY
qxaU4SxODOQKCH9UxjnrBg59X8lcph8L4vQyJZhjQRdKwzVYKy8VPu5ttHuaW9mF64aVA1pfXdeF
uM9zz0nRz4Nqp7Z3pcTKG/n1S0paqAz0hGHrdEFhPr1oAAbo6x2CjL7xknGiUMGZg1M4IVuTiMnV
4UhcpW4tuAlvIuwOipHbG1xBv5nH2flRWUIygXNwXj3GM5NTZHylwo4obLPV80XUtuoHTtxcJUu4
t9C4kEXGwf9g0lzqN7OR/rtqCo0/7TK7GaQfvgGoKGshtYOE6OWdu3Pq3vZNJ5Mz3PJGzA3p0cnD
Hwcn5p74oN0JjYAJlPYMNN4rzgpzsREG/0YiMQ8zpdI3EvVhZZIILAQ1UJXLDMRaal3I0ZALaOWG
DKLdsZWoVwOQvasE8ydLKWnO+OaE4yG5oP2nT+wOLVydrw48iPEyUFsDrBKxHAzfu8/jqD4o17t8
vOsdw8Us5kNJEb7lH8uXVQimedvJSVzM4N1DhwZiqdr43sXGq9gt0XyuOQzvcMS7O5g0i4/4UVF/
c6y9b6TATxXnt3NNqJIhBIXgx7s/L1poXpA5R1jx33l3mNH5JvpP36VOwEH4Q77TIQG2+fFYsNjj
4oo6eoJlQCfV5AzgJ0XCBig1cWC7y5LU++mNvOgT6AtUXwvr4MoEGbkNADtrzGsZlak2QlJvkrCe
M87V7S5gvXjghfToYVgEGZ1AtB3/R8HZOdqPFmvxSy5EqdWQ616SY3vVPDfUNcTgmkk3yzjlIEuP
3lnP74dSf+FfLStPt9+VaCBEltt4sEixPAtunrmqvy2mskjUnSo+WwBFipCA74JcjKfvC+76plKG
C3CzWLTHtWe2KlRKx54NL7m/Bd2z49Nfa9MyekqWCRXV2VcFDVhGlnPiH/yINImjdn3fF2Dwy/5A
vLVIEC5sgaI5+5R4Jv/Iy5dxZmQg1wffdsyES/pJcM5Pco1QdENAvlBr62t+MEnF8IFljGzKEr9w
OnjbhKQqv+qxL7zzmfdnBVW47iDKB0T6vTXTZyV+5L+f/b6g95FWnLojsBtNPe6YO73SZD9XfV/X
Q4/VbaEEbNTRw6D//Put8MTTwWb3xRkfR2jV2RsmoVVi9/U/a3uUOFHBbOLuwFCrEm9o15T0xFal
Ki4Qk/5ddiLidnO1NZ4XB7ZMPoQq+7meRhaKBb4hTX5GNDwIhWQxrykrTDDrwtHecLZy5huDKemO
GR5cd2Wp6jHt3TA/AlEy5XCF6/AWGztqmP54DKEduujQW1Pclb5SOTse+PdDq1Et0SXyn6tgD6EM
zbSD4oN2dy0fElKcFIra4HJeHnW3aP4jcfGQ/O5+CCQChGO6BJRDNg2ojBFpglsOrpx1tD4O7Ukz
zekw8JSNO8LqJbHJ5o5OguyR8q+Dj3h6hdHxdAsPo2+PtgzXeD/b/qgKiNpP4M1O67lVKAF0Z9om
rVRmTH4h+2P3aLUfbR9kW9gnxdv6clnbSKwr+TaIgMN/7+3qMNnoUnO9PwZeJxGi0T5VeCwPuJnx
GshLaKCD9lsvwSjPMV6mLSxOXDezY961oLx+H4BBO8p8vIXihpHq8qugIkpW/OxZDlUHUzBfa+Yq
dT4+Oma4esgX8Kmg07TB0I0yahVO3XfHy7EBRIVWuKZXGsILRaoSHVKu6rjnD7ZOBpfjBoQUcudH
RJFYa1E15MhnUBgcT2r2qbZ7rrOzKsANqkBBTK+TUXwX3kOQ7U7sS4iSwIDNPcs1AQmt3w3kSoWW
yy0uPddkyeLU1f6/JJQ1/dcyJfKCPEZ8BK9Ne7BwI6YlKiT3Lrm0d/OC41L5LQIGY5HFlGURMhlZ
rF2vDidM69PO5notRhXJ6SxWz63axgXE+d+jXaMTpVjnQRS/sM2IowJzp9z+mv0jXmQW2poVroaG
jR5ZukYOUgDw9dVPWXtMajOLIBxWeTTaFHYiIiiKq48GdInHFKa9fant67Rdmwh85D1pfv4AqnST
mzyon0jr3DoLNVRHhWqyWfTp3+VHBg3sZkKoH+INK++o8M4Dv9HZWetHLO5qe1wZO+hVffgCl7If
boOYkKa2M4zV8qluMEsuKv87Km/uSfKRUb2Tv/ZXWHn/m4EElC7Ygd15PfGBcUrc5AR0Z33hqBJ/
SQK8EE/cQEw3L2DZDux+Q2A3xc1FuBlkqv5OjjP/FA4GEfrKPdrJs2LtfcGFkJl6wC4xZVheYzIS
6P+ZaH6xxw3S9q8t0RFVBtiOokxb9znMSI+oxgrvopoQJxdog4yQJ3FYzqYwe8Yvc1L5kjTiigip
/Pb5ggKjel4KWUfQGjEsUgvM5LpGOSvYZB3cIIsFkK3l6ugcs42WN0zkcV91TiCS3NYu/upCDb8z
joZGtPIZppXN0wQ+KbdiyHQ1nRcLZkh/lbo8zMN3muROF3TUxF+y2vqd2dv44rxN6BYHokW96kBE
LJKHEL8ggmRx4dTtIXeOCjn8FpL4GJJ6qqRW/AIlMz0z0ojPkY60RgNw5fyGqIG7JnhsGq5hmCRK
Vlbw3TiHF5HoQehyMeykZWKO0G9eqnI/O6g1zPXOjIuSX6giYaNAb3TQqAKNgurysn8KhXKMncQQ
a3PZBGLDNaD23G8sOWf7dGSz7GUq4s3pvWc3s3+N43jgY0jIYEWnnnj5OIQvx/DueDo8la1aEm0T
YCI+ZpgQnvPipW5fky4ifvdwmyc8cOTzYT4jGvG6Vu44WU26cyeGwXDLaoMvNOqWbFhf1DiGKWHl
0NzU7MbsUnAUCSPZo5cJKi+QB1m2yTrMsz9neCXIOteO3+Ot/POC/GCVDKiVwj9fH9ZVYwRfb+oq
XfoIMvW3axlQNMDijePseKF86ii6KiqD9BQru87+sZ/baqvqxI/Y98252UsWSJ7XknJ/9+xexEA6
etAKfqn6MJdgTOVLt5Yzb/VfOleV5zUZqljhdWQ6Y3EpoxlI+fAqsnJlcmpQ1E35OpfBs7P00fwT
AOOZMRkzaN5NFAaDsPjtPMHr2MUfzLIrWO05Xvtz0O8qr75ZvqG9XJXTkDLkPD/nQOQ/IUAM8LOW
KxsH1IIBq9X6EoX5CfWNk7R/kh4v6V2vU9K/i4l71CsOjcP/IKTSH3BpFFJsTuludzKU7NJhu2Yz
sQUGFxWKZRxN8wRAL1+ktXJ/6rXZTLSsRyLsYDPAOO+YTetBGFti2uuA8jT/LUW+WHNRtgiKj5lC
Qdlb+o5Qe45q1h5+sLk0ZsEGhw+Z6FaAlwL6bOVzvPbGp0RwNngtrB/YwpSz0Sy+O4WoFvRWTsiD
27ixFGXDaHNvPHZ3Yy8e3gX+kM1tyz90f8ZIGIlcvTTIebxaTP1rmE75SGFYpbUCdC43sciUenvD
/oAmqRAbxhf5pjVZW5Tk9pjEna8Ja8/OG0rMmfcD1JiC8Bi5wLDBHPqcCEkTp7iJ0I3Y5Bc7Bqh6
8sDHSfuv9uRT62SKJau+ZS5zMNEqOp0eSekxhtZF0JszdjxYPCT+W+zuDxILUCHRa7HCvoo6ccWz
FbWmnqLX1F1kzMlzKuyYQTXaMICCtt13v5UNb4rpjbyr6wjN8TxMbu59Dm/y7clM9Gegx8d9eAfD
dSvfkgx7b/td4XZZ70E8uDOtekzbpl/ycGNIrfjCetNcsT0GCD8gWBmC6qQEjzfmbFMRx9bXVWj7
bT7lXyy5w5ZleD1ReSzIUUqpa1EpLs4NBiIkLJZW8R1zfUu1Y80tqnfLygoOaLQrPAyOrjZr41AE
48w5JP5oxiGW51mB59Cth1PpeMItjzPWg4u30svFtHPPTGcSwZCeRa+FWZejUqB+4iOhWeJ6FNrC
C/qCfx3GhNZHyxJdo2QjW3Mk5dfujrYTAOi6HuO9t9qoGQK2caMzF9rNIl96kOCcARrDf4Yi9+OE
s816wNq2npqQ6URZ5yYXoXV1kLBZYA9sMkbc1IOl9Rl5sXa7YuA8MREQpvQW9tf0u0yR6GYorSQ9
tl+Qfphy/g0F4DryDo75KwMNypW9iqeSnRKa9UInj+g70PP0EX3LivV4gld9ru1IEi7ZpSvMFDWY
K4ooWvn7dba2oKnZp5f6fNMXhr69SpdC4NkNFrJOly2i3AupMkM9A0YsSf+CdLxPLpypjKsSl5Eo
woo3FLOAyVRNKIppscQ9RDZxEqciuJQ+fCmpp51qZl+0KTPMnmw0PD08ixdqDfFzJWnEyvvwiEbF
dsHliaBJh843I8QT0ICQFGpFZywIhgYWQAWEOHQz4H8hiMFEBPbiGIUiQSBWdsvzgk36iih9l3oQ
IX7Iz9Jh95/e84++xm7m/4g6UuaFawFg2Kc0kM3iWu/erwMu2X4pOEK/va3QylWFzF+QPg6PQrWu
0J29k5dooqptecpDzVbYFeaeS18A4sZxBEUDyn29Xsw0Wb/XtkOWfoEs4WqP6BnpOeno+wiRapLN
sQXkyOsWhCz7XNdInRafq3gY01eupzBerd6SkQqPM7Cxr9rXskuprYm4fp7gzzXyo6N6sXA9d9KC
QqO8rX6Tmnwb6NvG7FKp3TC7YydYiOmgFsfVR9Up/zMkFyW4j4uLjiOsmBEtuj1iXBwBeTxQmAZ2
gRkJkWiK0r+dfc8Yh82pThu61OwHekMZQQmI8lHG/aHFdzKr1qvyn95ip8u+45VW+pHYwAm/uHKo
XmxqvOthyH2lN/x7t/eXW651vYaZCGZys73PfK3oy2yOeyBLMvuHHF8/ZG5eQ/CGdUszOfnu8wm9
/cij/WuXtaNPEDbrMV1gf8S8DXQRKyeQTCUYbgLdZM7NTL8N8t69bZI/PneqTxASuZgj+LNNw6Oh
mI2ozffIzIe+Dv8tCayotGdRDx/KhR/sFy9uVbxAt4tcpcpTLy0gO4It00tyVNnGWWKIU0RUUygG
BHC5zfuqegXodD8Bg4eXfyH/zifusLQ0e/BE5zZXg497wmv0eUPCKeedh7O1QYcs97Wt9VMsja37
chs/5xtFO6IyhOWvIaVLcA0bftPb0/Sp8dT2/BqlLCdiw1tYYFHuIXuCBXmTneKd5rCjXoyKImeG
KAFFjpF1B73k4V2zME0XGCo/IL94bDpMZgiRJ8+9HlEFZ31iQ3kvYwdylccxhOG/nCvKPiSJ8xW3
qnlUTS6LejfmQvpzgOJ42/eitTWCg1EeD7nQA0nXtEzUAQugIDLK3CqO7mmngGKNaTq8B8Cp55v+
tpwGlfp7841mStVXCoP8T7uo95rV1uBOm1n1ZNJj6HlvgQMz/K42mc4j4IqN7idNKu+Q1HlhDX6M
CYC4EXJUCgKpi71WoQ5p08S9NzyDgAuh8uz/5peZk38Ho2agNe1gpHOqopJWgjUlihiMW8ZKBJy5
PT60Bz0PlLsyinkWpnZR2q7Mjx3IpCu1J0oUFlGiBCaZMTVWfaqjTSRbBq6DRozA2hkL1Jxn1orr
iGgwX2lRiaSpClXq4GHQAtjWKTsfQqwPOdmcruTRjGDVjRu9G3kXpqGfld3MnvetpBkXZ4hKaKlA
ErGbpKW1TkdIBFZhH8DA0Gdf+X1j/DvsMbI+Pv/4deTvB8nSauqXFf/94A5giH/HPWlZbbNtaPBH
NQbM8EIKelPmdeT4mqpTvmpiUfemBhZA+XVM8x6Ce8ysmqT7q3LrKExZyon5HabsJ0BHzAM/lvwH
EGfQs93NEZd0dd/lub9nsKXZMIU5GcFPhXHS+yU3mbArmiwblEn2Jyt6MuOITH5+DDwqSZzSFJZG
nijlsx7/GOSZqzJ//dTtSdEgj+c251BFFx2pd4vZcM6dprlu4Iau8BgHXbYY21Edd7ZssdQCRltj
2/VvoEG5p2zgXxk+lk3iKjYrMzAeuhv9JEdLd1rGf4Qxn7FGuEZlOvhie4QHpwLmtbzuexoOgvMO
C6ZqYCdgInwMz0siv4C0j/vUzORVdyL1Z40vCoYE4aTSq92284XEhYgb4QYvPiidSFmMBNVvlsm9
5Q0LlG5KN/XKGcs+9kr2XM32NissqXZrrDjWSNivelvSh8rGsGj1QPcNTH1o91CEXuFwMx240Quv
R14ic0FpjOoAO4FTwi1R71n3lVihEy6/gkI4aIyynBFRurp3Q8zQQ+u9DjpXAqLY9/8odSnszqPk
5+E1NcEYoIvO9lcWN4N0oQYJLqrFJm6eD0q4HxQaDoYk72i+q+O7LTp3Qq9lBiwNwzvOyC6/X6t0
kBQDz3zVpOf+5wk0K90KP9kqTKLZ/+jd96dULNQbFtBi3Gw6az3n2uD3MvajnNMpS5SHacxQ3npA
x/koXG7Xqc3h2bLWndVMCrE9WiWrz7Z/kcslgayzEum49gT9E6UFotIHmjhaQMRuoOFAvUfKM7Rc
XsORCK+uI90Nh9Zk9y2IpGakYGVJigEkhPx3+TGi9VHdWouWHgPNXoopPtnbjUwSgfZHzXjB0sN9
tcTaWgnqgwcxMJ24z97Wuu0ObuuHww14JM3eOCwFOKM6eoliK8GzqlENdZiF3TCfATgquaNxD7gN
FjONZ35xjW965eWBTT0MaBPcxzLzacfaUEKTJyXGMM8PuO5hwXiUjJUojf/ehDDxRDc+A9A4MIZh
UFuRyWeKqlMhDrV+EYZ1L249AY//vmLLPRYg0vaoHu8JnoLnC3lN40XwZ41f3dIU1M94ErbGwdq3
rQXOUXSu9cuNhooxxXD7kO11JZuRFKb4ZaQymrnUbw8CO8nkjMW1AnHTfi3+SRKMAVI9QMXZoO4d
ddyZ3P+do6yJVOs7MpGXzwLwourbQcN2SjZnGRXTUAkLhdIvKw0zpp9f6PU6o79Sqi7MneFXhpVp
IiDo43IR/pZYkIvrAO83pkPheiRnPGcdtEs+tgqUVewNLl5bz6nmS37z7LVpFIuFsT6rx0wxZx1h
XzdlaTe4Mj0wYMBQzeL8HQhI9JBmW/FyeNvyrGxSvGZ9DUMnDbiAZ9xK2RgHXijCyaLxfrxeyUzg
uVTa3ycHCaDchTh7CjotqlcIfMQHsueGipFqnSO31RJAFaFcv6lICJmbRQ0LjwUupFcXXNhG5axr
3WcP7CyJ+lZHPndLWIKh+HX7rM5FBzXt8XaXua2yOGbfC5BBXALxAN/pc/y2iwS6nfVL6a9n9Ork
HAlJunttwrD1B2K/DOz2WtKOKfGMtjdrtH30Loh24HqEZLRRN1wMKmYI92gI0VdTH5BAg6MkaNnX
N3odDXx1UMSWz4aAM2km72QAHDl9z4bf6F0cEFXRbyD8d6sJE6uNOfL0lTskG2zz7ps7HMzC6fLj
3i3aRSOFTDvdWJaCq7w+19AsTkrzwEfzx5AObBwFAltjVWgxtaSKFVLozoPwoWn2vo19RDa3SbNE
sq9PFyMvYFawxDZLiWq2jMJTEJGwK7D3IMV7r6H0N5K804/tIRJnUobtnw36WMaT1rV2S06Gno5D
hGUrp311urs+xLDSq20SfI6MdJDDrC+iQR2yBwISt1q88eFecw3Xax9iWWfkguADZMHlERCSpWy/
NLhAuEcDz11dgkfELv9NssZAa6isoTJoo63tltSr85Z/uEw+/xJqKeI7mrtWXsrltiBr0h4Onx/T
5QATOcPeYizeRSeS1HP/QA2L9btKg15b0SOoIGij81HcLgoBdy5qSCEWhB289x/PLnowODixlqck
mq5j9y10S2tjAOtMm7yViNQrjoLIPaGqeacllGqGdEmlJwheOVW/Z/Tqw9ZIejZGci5PUSJN358k
+iuVZSmtGq6KY8kZuqNTMy8Ub3Pklw4xdRprAVDaXohlOneDlZzXR468QOrjHXK/TBm9NGVAqjnL
285kHUxuc+60GHScmzjhNEhV8a6625+Q7O52Ip/uZIWto5uPAGD22bzLtLabcBw7m03xb/ORd+97
bVDS8GoJcejUQ+vrcUQQIZoJpPOamCmg7GrOc3qkFOIhOMZcndHDODuZbamVKAAzNZk0WHEbnHlh
+0P9n0Qe+DCI5MJLbKyQp1HGZma4oswbzxbgN26g/2hxQekako768xXhsCk1DugpeLA/lvg4t1YE
wNoMKryZoklWTdCVNciBDHOy9j894SPV/shPyG8yJ73oscezINAVT6QhiRq1EoFmtx5swmzzabrF
wMsBi4vmcxTz1E1gKTXGdSCgjcmbaFmJMONSS8mBPX6/JY/Wj4/QJanO4eIXZl6u//QR+N3Yej6J
HvyFildWX6QBHvvEgTuPDjuTEvmM9ZM0GqzAJ58UivRy9mdgwLLoXnbkzt723jh3yVxgB/CwNzd3
A3alm7aU5DvvEKt5HConZjIM/aAZNNMfONcEKO7xnp/YnjGU9j/CDP4yfLVak217OAzGpeudN5Zm
2OdFqGN9fNwW6v4Ghaj5qrZkCGS9+hPdbHIZ25aHLWk3vAWE2r/CiTqN57UfaphO9FccZCQdGWdx
7wVOFvGTjSt+iFAs+B3xxN2rOZzIKX51mlBdT21rRyPBjjiJEiH5rAOQyNNiyAxA/5YWP0zAJ7fb
z4YePhRqmCwH2X0tTHzWOe8utgoVmLn1pp5GAfE4TdErXxRkNziG0tDk9ZBoa+6kpP8OHv07NvaS
MyOetq22CXjZg2+kN+R9OjZV9xP2MF1Lbrq1j82xMXgpktQ1iRzXntFNKkd94lyzz9AIx2PlI8RF
xsU3BnI0U0tmJrN+t8xkreIhThOgCTWpT8cwGVDcnibUgjJv3S9QJ7YpXfnHOI38qLF1NalB3VJK
Hu3jszrEldijDIjCQQ+C1j/RISWafVO9317q0JpAmIu6YdlJSCaZZbPg3/hk4rGD5IpXqX6DC2/D
Uw5eaZ9cOTVdoR/fZluyKdE0+6bt9k2n0x4kT7DXIfziSq31vFKmaUW0crF350jHCta0t/Nu/pUz
Ke9h7gIYKAsf/Ivfm8vCxfuPDNP4d9ctdb9JI8OLU44q1qNBR1vu1JaVzMygTVQF9D+o/PzYYuGy
p3+i845fAWxvbTWEA/6gshJ7O+IsNpdJi7MkevD4ukiBxZVanOYayayF4jxwqmXaaRAQv9mhjhTX
pFdEEadgIlOYkiZkN1OtgSJU96IWqElDra+0P9QFA41NYGI8aDv8dXosA2QfTM1/bfEMsFJirFyv
r/wEsyer84GQrB2vZfpuY+wACtyWkDUiELGeqPxTf5TXHAiuHOfi/dajN96WA/hoyHF8hfrQM0du
7D9zlwzKY2wNqnp7rH3DM+Z2isLOII1Dxcs2BcKL4HFpy+zgfpJ6qm1vhJ+j81h/FjHMkFVnjCrm
qS1sgP6DY+NY5jKRVyLDXIveF2IXSsun9vY6tmUHYwvHVTdsxAr9Lrs61PQUFiy1XwKX0S2al3vp
kJlcn6UhtyRi9FnZzKt7NwB4eKmi+uPeH1H6hfPgsbhzYlykcepY1ww7WQQp8e5EZQfPVPOPlPc/
adMuzKqeWEWMtrMuwMkG0g3IW/a80rcDqw3i6FsvIC33qdnkZYiDHBMkssqrhn8eX9i/4TuXmfSU
IFd4n0y/lhNf9AEMoySNdpPnNOjSTZjeb/hVTISIipakGlUhWXCCvOKA5Gr7Yu5h3SiCJEeDjiPO
6Yx7DqASHYwpPymouKkiN8gJgUV7AIdqtZkpo1gWRss0Imio8EzFabkOXUDoVgqRBlqMB83m6u2k
WZ6mnoGZFM0w8vE+1ICjxiJUp7cdR/UJKn+2eKhJbkOhBQP/I6tPwr8G1QzSvQDXbdrBaj0B1hkC
iuqKSYdNKFQHEVyVZ6aCXfkClgLv5QpnFrn6Y87VqcwLsCrav+koFwI+JPsrM5F/KHlvyEdYSHxo
0mvWfQRiP4tfDq5wZ7RGwiEJ4wgMWvEu4SF1xgsEKj6BCCY+bbUAMiLZzrajCJYyc2p+Uy19c7jW
1Qfj/9c5dWBxc7y9u9HwxhfI8VQI71N3scXf3h4kRTYdmgLqQI0l/VngEyiSFHpkArAcoDLIhIQd
eB1IuxEhTX6RFHFfclab0pofmi2AQ5ZCzO14EllT7mHf7f8cgOIJHvr5TGmQzIAR5ti6DHlwFmws
y7IGlZMsRlQGu71S9zltT0j2mPH+hwF89Rfgh6jZCSicRVRSlDB0gvYjcArEcW5u68EZhHNLz80+
sk3TIFXZ73Q4C5je2nCCd2EFj/njYm6rdcdpeTJLNdSAOh5bR1ZK6ZB70qjvmY9Scoy5n+ueLK09
ASdcXPilMaBP57oHFh7O/Unsv1xJjEKkT3w8qV0d2/WdFit/skWahX2giQlXei6GeBQMym8D/8NF
CG1zHTG6KAlk4R+1eZlK75RE3izVtooqbRcOjARXyHYE+HcXQA/N9Ea9tRzwwLn6tBairKZk25Qa
M+xr7l9D5nMGuU0odA8EyzR0d9xjkq+pG2H5LUdJa12Y5tW/cUIp/zngTgV5DRqL2bENM1UKUnQP
sEGnMbi9yFfVoPlOCwF8f423vDRjgStwYosi4rpeNwfUaINf8X0yGzknKcKezkFYyxuRgZJ2IVTf
G+ih/Y7rc1x5nnujoeyYNhiWAb/tKdESf187cnpVMHxw9CjIF8f8825lNTUjZxAwDtgg95jKwVAL
MoNrGu+4uAy0Srro5vb/I9VaEBnIk7zoMGzdejARSCCDb1yVeF82stXn6Ykv2BcNPnHWGlMuXwO+
2TUP7tYpw4qA4pQKWEcZU25N5FOAUMV7D+mPtONlHNjDXa3g3LaPTkti4iAm1CMexs1CJVoiGLIJ
y+oFLEqaQmuSW0awS/KQ0+7KEoCy1kjc4LzG3S8OFOiXwQhLgndSR+FJz8Heehb2QwUmOszUWQ7L
Zj7UHhsDaS1ugY7O/XHKfBIZ9oxmRgpWFfN1WauZesCoBkmw9YQpHemwPvH4iF4b5b8HlKkFALaY
Mjw3AtelGr6uTW7oJTpHdMhbQig+NFquI7kHrEKo5NDOk0QY6szT8ud6nPmr4NnSVCrgr+3KCmri
YRuX/1mWeVjayWt3+tLzDqDvR5c0ncwZZKAxd2wMpQfuYATx2MDHT9koSxmr+vocsOE08El0/LQA
BEiFOqP3lqk+sBMVGmU9yCN7weM4rzA2Y5BEWA0uGsiW1rr7bVHWC4ZcmV2l0VVn+W28yjEhX1bk
EOGunceULgnsVASiiPnVeEJIISTEafA2RE7XCpH4HKabfSrpsJetKr4FGHrNWluuRio9yMuM3OtV
g5zx6DxRo5HYobCdaRYeS0D6ervv+itj1FisGqSn8IKrDFjrX/wrQy7V6tv73C8CxXTJcVcIpdo1
Mb48Bcu+OtcD3wDLTByh2rjEMo8pmxtiWawzC9OTVXFav6TtyfBMzrdT7QwSe07xjN2RS7ePp0nJ
bnziLN+ZkGz392NSjkgOM4v8+X2E3cfDJr0n26LtmtlxJ9dRK2iYhMRJXtt5H1YbfBQ6KyYid/8Z
w1CU52oXtIVD4VjK7/lQGFS90gb8r0JiqXDKmpaIQunP+pi5l6e7lR4FPQ7V66ylz6eAvECDglW4
PKphr0AveBhXFRlutIlv+pIRXZcVcjyaCs704CkME40CNDH2LsZH0BMeVMQZ6F7Vm84bk96Uyuin
GRkg4TyKU91+j2Oxy+neonnvmOzgSPkVGCQZcg0Da3EmjSpwaYmckUM7xs50B4AKzK+1+PN3cF7K
zTUCVERO1mvcxZWGFgvcCqWrISRSPStOxgBA0JrDtzDr+mlZadvzwVTW2Q9Nru333moagZySLmVb
9odBAKRGECiZxjoCys92m91dZ2O2le1qQ6hvspt/g+AN7sEcHPzCbzJvLF/SVqqr9U1DFKNQrrfI
gjumNIN9o4fwa4lmjJwD0IltOnR0TsSYjbsjdHzqNJqNRleDg5+cv299xc2PVyuO8gJ3Lmi2cSc9
tqHWUrLOugGJI4DxYKO5QoiZ3FFeoNqXr1g/iCgCLlsD6Ih/5rL1IK3CtU/LOHDlmEudsG2hUsLY
kte+mbqxkpe9wc2kyNUyKFPLIXfuBlilZSuHmEjeFxTvZAqqrk5gKrWRxzV+7J4V2maHq4sw+8db
pEPm3zgknLmMfWPoTmxtcydF6uWRcvOXsCbB5lrigUEuAHgeFsavVTUtHk/UkV8gWZzIEml9ynL3
k0IoVl0Juv2FT/GvO/0eKscAACLbCWrr6g2nVQc8Vjwh2qeXreXlE7kUkZqQoW1iBhPSFECXE0Du
YXG+zxlfnJdbcZW5n/neoRK5aQqdtofASDCclsi5dhlKDxEHGUfmF/IvCq8gD5VcOBMeKbqZwECm
PYWmRDJE+wvlYrNh3niVRgnQbWb59JoFkjRQi2lfiAZOPr8RTh+uGPg95m+YOIiJCyd+h8nNRTS8
PlIEZppcf3dHlycn7lX2bHE+8jDcul+aD3gv/QCtwuSiHhu3QesRraIDJIUcyKJ3D2l2nCHmRpmd
TsYPV+VLuZNzQzFkmo71blgFSo13+hbVpS0/xyaZ+n3EQw58bhnKsbk77zY+rBmQ9t27aLcXmeyD
M8Zs9vm3HT1WQDXtQowqibNwUs+d4HxNQb9qGgfW5O1twodw51/U6dZBSP1cAH7EDvTiLwDL/ZPe
I+AbefAgs9T9MUkAydUzResSBFp0OonxvruJHPNUzVr7QDQyC3nmPeWKamUSf9jvdFJcWntzkc1q
BZDzfJM6rKVA9eTlmKIzcQSHwWp1Yqfdt1cbam/4AdppvOhqVt66IkeSyqU3uyGuqo4rsPICy9ii
85Clzw9PCJDGQXfhzTwDup6ABNRBRq0i4HaSiEkh+4lRVsAA5ktxFqstsSZYdyeOXrDJj917VcPq
DQaPhMrqmvP0sGygSpkjTkCxrv9D++rMOnwBuJNMHaPlB4jqte7biUgCmIecGvrku79kUfVskHHn
bh+H93fM/SBGtn3uyBj36O3ntWbSlgUhAE0sUy3Iu+/2hkEMzGaEIb1TKd2BqmlZ3f5gm9Md5rgs
IyuZbuc+KTG7Vzn2S1NJ1cx30gzJOn01dLHidSEqgXQfMqUQb5/Ckv5ToMlpW10JDBVMCpFJSUwv
5GbjYoEO+ayv594rEUH2dM+g9+cu69ZwLApshVujicL2vUGhATpKN2PsKFIYqkh6fy+rwelJOXrx
/BCLOlRyGV48eN4j0AqaqLWNnRrpvRJVFZI/c1NdnkMUKOeaOF5rfWRuKhM55ST9iP2slsQXV5fp
2xKbOdn2TARm2HFQlS/QjEq2Yx75UW4XN5cH4+wNB7QBDn9COp1Ia2tXgyNbNVmg6hMm5lOKnRx/
MhwqEzugTuOKdk1izMP8+Du+7OiAM1e7Pk9UtknPgEktx42LeRqBGtgxESCHIUg3OwbcDpUMTNRS
UGwnH0PGVLCRLof3L/8bnf85mIjFu0VcTevEIZihKTesGt+2ZeP75LgxVQWu343OMqhhgdgEEsyK
/kZ+HQGLnWJxq5JJ2C5KVvY6jC9/EPbb8WOK2maqGSp2ADdHVCBMRfMRkElBO0eAq4wMhyt7+4ha
0QUkX1fXw49XtDI4+iyUqV0IcRnoJ8Avoq5meOj+RBTYYnV0ud+h5mKEX3f8jeEO9xVMxXHSU18P
fmr3fpDiH/tyADxwt9wWaP7Ui3eeBuu1bE4N88wCwoe/OcKqNdG227ZEcfIIRGU2S7f3l0NK1Z7b
EJ1VxC9DuDUYDLDBf859MqYXDLNyulGAsbhyXzDt7tHNAMn1SYvqqALPtr6M15I7D3p8wnwwtgds
hyRzQ50IEHmdkAVZI0mitNYrTbTOcEnLtCggR/wHVMZdJzWCnWDV3D/Q5GudbnHW5ISXMY8lBuDz
wjPwCIeeSaSxZF7bI3WJLc2lB5eCfX0/AN9+RNcTB4f/z0bqf+S+Acb1QKLe59gmVmE/RnZrvH1Y
5vZEhqTAvZ+V+b9ai1MjhFozMTgQzabCkWiI65j7TGnGx5t0CgG3N1NBUzEF+neKBqMKaZqLIkuP
pVyS0y3P6Ox5bt/ZfEDZmPaP3ufI/eLywPucb48BTivXdNyY1bTbSqSXO7teh2Jez8LdfejU/f25
co4rU3kpTzwz/8p6BHfvPAdGBSTooGA9YQl28ZHuGb0hNN/eB4kOtTI/S/MSrsmR81XBi5QxYH/E
7Y1zjRS5zNk/ER5Pn/RbuWVpcqi1XXGmvxtfJQX94PuEyDfcUw2wuQGsvagkRPPiqK8yxV5TBfsx
rI5XxCaq4j7BBPdfkabCuCFsUp3SfSxYGFv4Ra3HOU64O4LuerMAtQ2UBDZ2nwkBSf/75Qo6Rwvq
sUi1Krk5UfGGtGj2HNdkWpUFgZ/67h8mtHW169THz5OIQu91syzU9umdZj+KPiV2YhHTOc+xDz+5
aS45hIeRWb1i6URtCE8Se9KlZQLtbz3Lyc0Mn9oyOJtaU7Ruc4KRcnXxQPDewCFSdMl8nak24vEP
nybLP+asLLwKG2DOfd0qFXnhNcH6PuhBAKERRfC6fJ3f+W7dqW0mZA9mUvt86zk6Qc+lpzt3EIxg
rx71OrLlo7t/PWHKYgA4BupXcykt4AmVGYxrNe2pWyaW3Wbf7SjR5IVEKMGWxMq7+YXIcD4uURfk
1O4GKZt5X2BPLieitT5EmlgLKy0vYY4byU98iO0vhPxo/wUpFmpsxi9wluDfct0RCbgOenO/0JKX
QbzStxRnjgqsn+ZfZJXnPE34/lXh0D2MBoszr4EJToMMCNSbNv57I1phjgXE9N0kqjkF9haJ+9OV
h57Q0gbCKgPSzHfHlXYpT+Zkb3i73pSC3NaJMllH6825fDKucYpgipxWnIv/Rb/hcI/SNHXNQJo4
qHWgl/FyjJnbPcb945jByZCWA0M+HSJ/K8VvGVAL6BRzXC5FLFFb9g/rr9ep4XwpTJICLi+UBW8T
bBDq+8vEeF0gYg1fJwNll4NsM3MJ8cbxhRxt/oOvfao42S4i4yEVe9yDE9SAUxDgggRq3qQPSwf3
4dKttfv6rzeSJhYwqrCoNpDpzDD9kfUr0YP1tHtOAmypgxgTTF/VZG4KyRZL3VMTTua7UurxJnXi
HsLDFkZdCXHaL5OM67tGbjtUuZs5DnAP0P3b8boJXEVtNoRizywhDW6xWAW1EuYe/x16iqM53igo
8n4zIx3gtzBow0OODlTyygZUUOxTaVhryLpxSo+3rHpbvOKs4CQ+5pHWpcN+u/bCJ6bBxF91dCgD
Pq+NYiCNILNx3PRngnmkHmoU4wOs0s/UWcGupQdYGNWQpYkgb4CQ6CC+WEf+wqpreLCKub64j4yH
Y7DmXPFoX20+yOGDkQd9bF1RCEcpMR0KgiUK+Eh0LXzHdk6inW0BxGZqUmQw0/GZPJhop2i448GB
TKKQXWRqB6Z9bn5BVSbM57ENne8TRvZ33SBRVKx7BOvITLRNJoqa42OscZaaEeUGD/7u9qWJzOeW
sf0NQn4AHP9vYlWatr6NXcHebUzuQYdMZSnhDhYFn619Oaqm05FIlkcVbBax92wDmTXnKdYZdtxJ
mNej7g5jwsoJuNLhgn11JUHSQ1nJtSoczgML5MTngHPpazNmDEVLCvj116F97PG+7gCygLz8CWhH
pNgc/bAOAEhYSQedKZNKi2/nhAyqrqvnmTK2MAjaiEZOGS2TxN9UTMizPM7ypEU1WkzqwQD17DCd
C4nfUZGVljVQjMHpyWK+XVZno6QQdLdFtXre7osApJjgVp4oz/Ol2dOt27t+kH7kgljqig5K4gJI
eBY1TSSmRmWss1ULf0aUg+cjx3hLzcY2CiEdOlmR8LJk/fK9czkWyjRxYan7I+v+PkISlJwkrwr3
mA/hMfbzNy14e48mcL6Bsule7l1SVARZq3QG0mjC1eubEVqIcVXiJvIUaHKZzqJ1L3uknypDdksk
foboTVIrp8SIIlXPqIlyvg7P2UlTVxExkZ0tNwMsvDFScoF/yP9OUpWbyRM+9CVqQOViUiAczmKv
xKASOXMnzmX6lEcORDQtQ5aEgobr/sN/xGLLJrK8bQRo147DX/9ae7UgEzxExPqsOPoHh5qHVgtB
iPruWawElecDR/W6Cc0MRjvoXz0q/HzI7hX4HL97LRh9Sr1Q0+rQ3hakmmmSYUjOTkl7cGv9nkYU
gSPrfTY70tzBBwX6WQZrZsFR4MgSW29BtFIZVypc225DKEjlRGI+/dJEhUTYrs26H55oL5gna7qd
XDXDKPmXPXLrFTFi5qn87dXYmoecF66PDM9ZLwOkvSzKKyL02ic9SWca2l8/PcdhReE9A9QHiHiz
Q/CV/03vcPAKl8In5o1kVBzQe2UU1nDd79SO7PiW0dQMfkPpmwUvXNdfA3kH5OUJ6glt+puA9BH2
61Gz+pMwt/6MXiSkQ/lqDtYI+nhZkrbsB5QT77Pte9kjZuaBghjK59L9B/S80CVaDEbsE2SdJw05
AELeIykCy4zOGXS959SbErn8aFjvo6dogJpJ9zcYn93VJtGQ8oizdEU/Ir/ZPjoOFLU5US+lGtq6
N56RQl3D04beJhN1ulRJS3ugIhC5Khl24AotIc4EHOX93zaOe+7rc4+s1CwLYePimEMaIHYrWO3B
QFP3ELbgt1mufUwgtwDRHaItYk0AdfKSdTHuJvMQLLuXUr6T0ULCt5BISrYFjml4hjKLru6HWU9F
ZfNR7bzfLg8GdEnYqKKikykIAG21TED0IMhjt9FwnRQ207UlJPW6Gbh9T6Pm0XH78pIHDyGqGTPm
i5USbjsojMRgmILcynlmuMazxhH8sKSTDAyijez97UEgL4xIka7aFCMAlsgB4yD4sKzUMS1Jn7/A
fJxnrt6gmPPT8034MLKTfRaBBqxXUe1CIVzs5Gxdo2kI2yFtfQHh76efxkUnBlEzJUY6AiwxNEfP
fDWoMLeQCYL6zc9lQUUTdhdWt3fPR15dWdeIRFmJUiRyF0lFMoIXoOVUpW1snP0fG3IAWzxrE2R8
o+SH3N3NSc7YQpY2npOxQDssIXPqK2PgiFwOcbW8Ef5FI5GmlTwNv158eRB3hmrVKH5ND9RmSe1R
PQxkHaWKwEnW+oPFgB4ogTZ8cdP3GM+cRZWyW2+eEGXAoybZB9XcDz53g0QpmH+gpvJAC1Yn07RF
ckJRxqdP6QNruq6O8pxcoytm1QHcoHLCCk/IPH9tzBcG/KO6Rwin7Myfc6c+5goKZ5y31iUwPR58
DjWTQK12VfWyW8aT4r1dC6F3hmrJblUK6C9P6ZWf2EWHGeTRB833EpF3OuSL0U5/IMaqdARXe9dG
m1BbS3w0/HZTJoIM11mj1u12OgK+hsBplnDifyD1kKQ4zPN6oJqIf6DFlHfo41aCoq6p6BEojTwE
6iNMrFe+tuMXl4Iv8YQOpd+XoNpQk9vzOmaqi7gjFm6rQUtgF77KLhpScJPtnDm9V3Ibi2zh+Sbr
JxIOpfhs3opz6Wv2VIlonJvmnte/5q63Ux3hn6nFSYTFbE1iYkvOWVOEUVMaaYUEbY2E4NJQiMTx
peZsntQJbhyvXP7YSOVKqtSqK3GLGky9vL81Rff9ckUHd3I0s7dpgkzmlplwsiu4/KbBfEpiMo+L
Wb45cqy+CzJyIMiZ+qvTZ2pJHVmdgXsAEndZceEgwpHrYZjNybBiRyJ58SEj0JrsOrQhn+AiPMt3
wF2C0Bp4zwnlMy+gNIYsdsgax9dpgDHfWLJB6bB/pAkfWjXFAADIG+3t3Q9wkQaBkfSkFlP1uxwj
m9WqwszuYJuabXXWwHVnMnqF2ySSNKWG1Wq8QoNBPpUXykNpe/HCTlDGjxY2x9tx8Jpx8k/qUrsq
jSWXIFTx47qYci6RWtnyFLgin2YXRViUQ7eX7YdRNvuIhfvrOdoToEoHKfYNFRfwt5tCEhE+DQiD
qLOc14aYAWAM07nC8iKcNX4G21sEVpk2dPVLptc9a7CssGaTbQAZrXsMq9x68DDh0IqTydhV+npi
GpXD2T/vbme9oT4anwjJyjIUnw3eio0YpXAKlea1oC7LtCXOZy+gipdB9yw9Fogo4poK8MQ3k5wb
jHkupaomUjnHpQ9Z27xjRLtsWoFFtGd1ziYSgnswMxIdGUK5o3SNzrn4mweUvRtgY/vkt0c2ViB3
BXWMaOT+lDUufH5hQFn442WBEEU9LkQvROOMwbB8SzYCdin8CD/Vub2Anov6XS/wZkPQWW31dYbX
D+chbadCd+cF9dpY02qXS0glzcY6mmuCCQ2xaZkEsjHShRpv8RtkOZqBp34B9xrrMGhEZFvvZyuE
y4S3yT+JrVKT0Bo1G5sLOd1weC97Dg6klZBik+SfQLbnccVmoG2c6KYYO9PJQGjh7RuOAUBfvUY9
mIdpHVp4zY7IauG/2i3gUR4NdjhNIrBX+xdf1i8S5oe6sCeOrfsVxtU7pGkTS7HDdyuq59Q5Widm
xxRg+nJx3tEIIMLX43c+9PH9tYoNkO4mOGWH/NmkI339idNwPZDoxcKi1L4JnJ0vUkUnxjf/92Hp
sm9UGF0Tm6lSUObsls+CfsyaMLj7Wj5ATZVLpQYCD6A5LW5ETu0Iwglg2daJWkpQmoRuuQPKLPV8
toEaY1pf19OrYfe6uW4RffObLoG3bGVKAiKcgXNDULBKVlafNmn8Cu21Xc9B64BtVbl/vGEOOwCk
w3SBbucK6hb67oRR3ibk8cg488oJ0PzIRCTmwaZgAQvBvPeghJLhPTKI6OsM24iOhIaB6kNpikYC
EmDCVF53lWpeGOPtQGIknv/1Zqany7+hWh3ym4PFdMSdEv+xg/cvkjuPb7+5BjWeJgatckU9ofWt
INMrUxqEYD3+3qxBo1paPwZHmlHSgV4dlJlz+UvF9dVyN6k/D3wd71hmbYhnGnr2EZYyvtRQaRyo
3qp6ucLBM/wjwvrqC7FiOCtMJ6+bbOCqhgn7yXM3XXJ+A8BlrI/9HsV4ydWxYSc2WnbOGbvdyPNm
+F0pmaqbqWHnGn5kS7jy9hDO6esmRfew8G/JslQFC1lzwFesPrDN8gaWZMM8EU0fEcPe2r68pFFi
TlNtNkNJHVtgSGjxzxcn86QCrmdLFdvInx9DVQZkNkK3IuZywjiDuQZ4VUz2iWZVUTQibXS3eeVb
ckwagGmp7l9e795w3JB3OF238Q4kdthgXnzj5WJXEmPvgWS4EZGq+qGBqA4UQaOqmLJwac3XuLSV
snz5JZf4a2/Ug62bQXA3jOJ/OlYHq0LXJVfZ8Ik8DjsGUrxynckVD08m3KBMsqUoO9EBmda194Dn
Ur3b4Q+IumDS8V0TK/iYOs+nNw0aFRysDWYwt7Yb2ZNVUcAh4gd8gHL8YFM2k8vg/a3/vxRXjOwH
h/Nl+Fh7IF+n1XLHIe0jCpFuszE8t4a++MkagzMhFYG2nu57MKpUZjfz4lH4MTtDi/o/QhIq7HsQ
4a2UapJyYSJMRMXYd3RcBBGWFf3V2H6YSs8J7+hEEoRC0EwziLw7fVXvUpoIFvbcKzh9ze4Blezm
Y2U5aRVQrWlxbCp+VIy6DErmMThagfDjZDadWi+0f0MWW093+7/Z6kyDSG3VtLBVeBVWyznGQdUT
FDuk7j5yA4+agcpQWif/0K++DMRELVfmsgurWhqbodxZ2e5eRJYquvddCZIhkab203R76A2C5zvw
g5PRE8Aj9Nx1Z03kX3ekrjmJf9Lq/TAlXgfvDNbYb6tP9JrBFVaCz6uOM/t+yB05O1DHW4oW2UIO
WPqtzK4ksKAjFV/yyP8EsLKTNM0foA07kdAmN0YB8rTpRHiLEr3XMAi6QRtBbtNV8TeUfu8zHkyM
FFv3XnL9lgO/wRPOotddbnyL7cQhdbGeN88WNO5IJANwTK92HXYIgVz0Fv/NfpHYZmxjqy7ft2Tg
i5EagWXBSr86j5Q8WfCveyJ2zNKCrHhbtk5UXFVwhJ6LoR0fV8PFui+ez/SRfQ27JsoHDOj4G/Ao
g20X5seUxMqZyVcPOwEtTKUC8nsfEkcCa6VCuTDMzOPenqX4IA+0s5TUArjps5uBTS751kwg+2KW
iDd8du9XCMxRGwr8oKfkK8j2mBQowuhQN80cVo4I08zmyO8wOKd6KwDqrTC6H7CkNioa6nRjb5gu
cKu8MlMbX6JFJPZwVzrKOBYE4ksYTqteiAwz+VNM/hJZd3haWuSRLEI7WeGHY0Lz6/z+U2s++OlT
4JlZXd6abRjPUPvPnNyfVkyp+NqtjkhSCi7AX48zBfZzhUjLrT0Z5DBBoqEIfJ+PZ/QAKyhE+/J0
kXgcdr/EFVyLJ2zRfoXs2SQx0w44Z5Tfn23M1NinxrhSNFhCABd3tAdgTA1wKgchjaIjdT/hhLJQ
IGq/usr5Gc5d3xrwx1CJ6bPCWXXIgnGIvoYhWS91TO7s7gCDHgEW56NL3le3YrQCV9qCJ5dZtrhG
5szyHBXwQgs1wkrdQgIC0dhQFVUK2pRHn7Y6oehwNjpmUBPv7Qf9ovtbWsgZzLiYbvjnkBXXP7R6
y0vXKVn+/I6hyXHC1uD5mraTOuFE2jwaxWdgkOHZK6rUqdvZSwH5WG7nbQmXpwlbl3QWXer9Un3q
EcL3hpDpif97bDzW1unj4yEeah+/x6ZSnuJBLI3EDUoxsdqxZv6GQ5zKit+nxt6A9KJwX566pnUz
Lz7nBfp6L/AO32FIx93xIg6NZl6weASK249rd3GLc9ZxaE0p1OeXjYVH+r3oZba0G4C/MU6Dklx5
WRUgflarze5MMgim/0hf1UknOxYeZ302sKLPxdXL+Yqsck4pUryJoRpWaBETd5R4GsjJWbL6QP1b
ag3mE1TdTjC5/4iZ0uIYlmy3LeYeMBWl4dW3uzrYZU2qjkbhfTFPAhXtNPyQ95YQKY8XU6sA6A4H
Vtg8eVDCrMiaLqT0SbC+pB3MzDnUqHXqrqe9pI9YmyUQURYEuUUBXOs8TxQKYsMtNDno+ggQLT3f
IVwZisuXv+5RPklG03XNbnbpJ0wWutmq/r61W8p4wqJv66LnRxLliq2va9OvXjsP0JlYAkHDbLh9
1bO1gGCcqw5M05b+6AJOhCf9JRQIbHUipj3kCFfAnJLz4K0kVKhZ4l37COBUysQf1KQnCrmCTdnY
E+9WMEqMQuAlfz/xbxjEyV7bxE6SLolokPJlZNbx9QepGEXqFo9L4N0v8IX3ex+dvmrMHhfmu7+n
CmaqR3949eDTWI8jkEurLBiHSrNHyOf2nnLZ5B0ZXX1DkAacE+BRaGMAUNt+sSV/qhwgsg1pL3S4
0AonH+v4Tzfg/LDX9Re49iQQoJIkPHbZT2naRf05OR5d+pw/xQd44W88ixXZGBkgcus04vB54nAI
1JPGOADSGN2VR/N6xO/Y+Ex0cuGzDP+hGv5nsxkldZdAJwhBQv4bnyDFpD4mb775zb+6wxKY1HwQ
+3p0JPfhOA2WufBETXms8osmNsGjuyYtBblaFLMKWenqs23sF9Fj9synyG2QCUu1EfNeiFrW2bBF
JbEkVpyxmmvKdFx5DW1PlUiro4rpDMzbAIR2J0q4VUZBvHliVyeEt1cmnps4VKNeAIWIcpB165Sn
QUJr5bX8sp4B0TA/zvu2ovzUAIMoItsBEOqbmyjb89it5DhjtnDQBN2BRizML/jo+Q2nU7dLY8KU
yna/8RXFPv9JQJUKz4td0d6tVR/F4jnc/3F7vkuT8jZ5vjL8ZI2Us/1WUYDJguMMphbY4+y+E8P1
QMNU5jTtHA4rl6mcdFOQXhced/ngZO1XrpA3VG8Fz1dgdp2hPbTrAK2NOHdeF3ncJGmEfOjLbCH+
7lJZ5v1GllX0yMh0MmfCtEBsYLcg7FlK9rly+lslHEMtHXqDa/2eHhjtT63sXtwJC947etd2gqMD
lAQwC+hRktxsJL+vw3j46PxYSLPCmdgFXhKsXUG0ay/DI1d2EKYaJeh9h/IsItmR0EYvORiKjiit
a9uNtO8p6DcwweYjf9Zsq7xxm8zAHpKBmH4nRsu36kgY0M4KLhsaWVeDBPA9l/HDHCWV1evmOfcq
2Nvjk5e8nCuaoqSqQQ6mwQ/R3z4Y913Z0+NQAV0RXdExzgYnNI4AhgqmSHESRZ8FogOpOPa3ljCq
vLdmpBBG+YSSCyLmfjCCDIO4J43Az7NKjCLT/W6d6QtaeIWT/upvK/Dd7DKdbWBFVnCPtbRyk4H0
EsIs45anAe6ab9bp/fhsdFrPtfspSU/ZPiXS52bLu7B3cLhoWnNinx8IM8vALwc3PueXLqDxdK0q
WVYg2iXoweiNy9n/H7CHm6SLxuCgdhCLdh5LvMbG2rwcvhB4pom/TqdpO5twfaLg4rIZYTnM+HFw
MGsOuKbKQdsKlxnunKdjhunmDOM4fiy9JagQ0T8ribiKXhGfR5Y6tqhoLWXmmo1QtT4CGzHhWvNa
dQSwmR44RsmFl+eXSKJd0XrrQIq8YfNTiV1+6feE6GxoNrFBmct8s3e0Cd+SeensftDrkUtyQKjl
etHBHIUPS7n43IqMx5wvAbjODRVgUXo49A3LnKGuGKPH1VIRPJwGmR10tPq/4GeclnemLwguwIiR
vMcE0XHHc+P7CHkDg22gsjA0YGd6WLOUEo2WX/cSguu06PTVJiq4OVs2SJeOGXwjCnbnf8EB1OFI
X8MXGz7TdlH81F5gkbLXnU5ul9fb/JUYjtP5ppd4yx8t2oUfxPHlw0u0bWjTGFi83Yqxmnm4KQH0
6LVsAUak6iNUrNQJyGJglMmWMGA2ARlCLBh88gxHDjmc+Y3Mo2JrKPU9PCOeibUv/Yb/wRbAoY0G
8E1/Q78OMS7SF+vDyPY14Dz+zhyEkxv/3aH/W6FOfXIfPVIV+XREEo5hKmI2pXV+TJZE4fmEdNCd
KgfYloBdaUbVTgaN0dxubM63O2qCqVhYq5QSGh9b2ha+1MUT0wh2ltE80exCexOdeWO9khl5av/8
LumIIDN9czSgJGtY7ZhIFdzER+D29oFUqaUnXjYt9hDexjwh5Jj7aL5By5UrvjkBjOEx69oh1oHb
/ZI8h7+lmFLmyQd2EC5p/BqNyaY0LsU2WVcfV4cGZCCU96tuZ0tpaABL6wm//w+2dpLSyB08iHe9
iHmx0AzzEQAfvOjBJ3KSaHh5/LHV4dRK6pFUxu9a4PFdm6O3S0Ecnftmspu5Q6kfU5r76YpAMWOj
bT5IHMWJCzx9RbDNIl7MoFvDBocdKK66TIh50c5r+3BfrlcH6q2dGsKA7qZ0KPDh3HHT0cJHLTMK
USlJ2Vz123aiHqN/2MdpfIk4hm04E1geD2djHCDBrh9Z0lCuZncszICdB6bwViPxxSIQtqYgaa1e
N5yzn5+EC59glxlYsqQbRtVvSGK4b/g1MNvQRFympCznqOQY6JuetOkO5zlPgq+1Cqp4cSm8u5sC
UZLIkB3P7NY1B9RacGAd+i4TbmORt/PxlHaxTjwo0FZ40dmcbkQijvavi/jCYl2y+ZoiOEZrRqmr
RlvlTKsPI19M890lR0dtPLG5xsJFhss6ijofo6nH2uOmZqA74er6xJ9zDYlceIXejFtSPZ6AqNNM
S4lp7OLll3TFrr/VjvoLXdd4FOoy2Z8xONo7rseZMUJDP5CHj2S0SK0H4b4IZSvTd9Ita3muAR+d
Coq1/2SlIUOygW3hP1W5Z5xw0y3ast7UdoztM7fyzM20ktSHjktW4mp9y7e3sGLnk8fVlPAQVlk8
T/eQTOZxH7F/fQa05i5r31ihNlU8ttBsn99DruMn9tUxltT/Ywfqb4HypzxRdgGsEAj3wI7xccDw
GmBl/XI/T3YZ0ibGFTBTJwIbm+HXlB1w39sJzgSKZi+bfemOiFn7amAbFgmMZpUX2mXL5VpVpFs8
OJwYhzfpBbv1vJjE8uqrMaPQzummUHcPVIhXpALffHKGUcAl/zG5mgz4Ju30Hr+oVXyc+C392/ek
wCee+9rn2GkQ5Fr+uPJKMGu6MaeZmyHcbC/TDYYnFrNaDZhaDuv/gFOJNqhnUMecFrndF5Ed3mt5
EeKCq5EuDw0S/gcZysrIzm3ulICyedXYHoKjSViOvqo3hiDos8acWY2gVumcRcGDhkcf5Q7Qofn6
Au//tCOfXm6f0OfksN4lQQDUosznRGVHA+Ep70Ta2ni4I3wuGqNuoXhwcEhoiIdFdtl/+jUrWv0I
V28j9XAKTOelQ9+nLGdoObxpLNj+o/Y1nSWAIRvBTCKCR6rE6ItwKVdiFnoTBEmNAKHfR6/5DpLM
X/5VJXr92oS26UqxQMLnXfpkDMt/EIxpj3Fn5UAvu0NlqifT/SqK60FzuH4YdPX84tpqYRlY6/gE
YAR0XxewU1T/WiGCUvD6nogN7y9IfxJBrLSSGNXhoUgHRt6nWT5oZP6u0b98q4PpUXaQa3ORH1QS
XLA9qvz1B7er19AOFNyXYR4H5AN/osCcM1RYHiRjFTmW1ISwb7F5apbUUX7dXdZOLL+vt+iGk9ZN
A7DePBTFdAIvgVMSdcbPtXRmIxirV9i2+iJbqdZ3A2T+Edw3sC+AXws/V38o8/vGLqGFFzg5ozt2
55nz/VgGRF1/N8QF90V4hKibMTzqOqLVTST/Sgia06CIJ221Hp5hnWjUE1xTEyqAA1TOqXbPYQgy
R4ziPdza6GVNsXXHniwB/x9yfINM/TMTOvLQHl+MAPqByhWxhGEoTTyAX70xp8GO1pCEX1yCUfbT
y1n7YX4HEWlLBRC9ZzlddAvnLmkqMTB8zgXzIU2ZfHx3uZ7Rr4RJ6W3seG3wAPO5iZJiFQPuaB04
W3nS5kNAJyTdH4ytimxOtdNDPipi/NXF1A3ua++0SrAXLqGsFRXmHrL4P7orxSfQG4tENzIWhjMd
2LS3FzKJ71Pmb8adR1elxHlDJrouiJrzIohZ933V8iWrnX6OhofiWFqNNs+3wzEW7xM7ukH+TIsj
7w50qahXON+NI6K8Y3z+4Uuzfi70jGDtKZEZ4b3ZUNcuCwELAGDew3CYh7t7D1N8V8mfMZ10is3Z
a5dQkAY7Xw7d0uUdTfyJEIR4rYi1UijrM6BBhFk9y24pqAdN2F3Q4LE1dtONdrxO5DwQZtPgr/rn
QGsjJemnuz6024FRe75bMy2baBn2ZTg2S3ao19esr0JsAP/DnqVmdrDC/OpeA4iQeoQ3sMyOgST6
cSrvoXY4/K13OQT7gjLPOn39wmqB06tTJGoExhfCNTNS0dvQmNeoMpceC7a2uGcV8mERta5tQRxW
E72pXk4asXOX7dH7U6N+LYsaHq+iWVkLOtzMRRTu6qNC6TAA+ihggzXoD1We5Agz+egeKJy3j93V
a05i+Fh/NXgf9pANDoWvtf1fztxFlOKGzTwhFKn4U6si8Q7jhfzD+WcmGWqQmyFWwy4H+HUI/Bgb
vvfwMqyNAzZ+c1B40KOqjMpp8UQuaVZWB7epg7B0j18zQw6aK8Tnad9Aa+UWPufRMrgMxMaAPEJx
cLNQTa20W7rRU0q/PfYL5vGQxYnQkdB0XAs0uDHiuFfaEqxLOrC34XAxb6ECz1v11R8DT3ZZPVax
Ff2rKzQGQNwWDUzU7vLXPmjq0u6DbIA35Fb2NhdAALgFUh5n8hNPWzfffqGla6SjspLNTSmtpJMy
cphVdPnw1/5kYr9koYE/fqSjIr5xcFTGznm63FUmjMMbHGxD6b17wCi4VYX8AOtLRvRnq1ul1UOz
ABAaFmQT9deY4/ZFw3OTThB05qR+pIvcAEi1wNQ1HEulJcJbcEI6oB9IeoitcKAMIlDxRbaRMtf6
Q3A2QK+0LnoCzYeiqqft61KVQPXYdN3XbXyI+uZJBytQyISiQhMUH+RNaYCrgEkRNV3Sb2RlbZU2
KR519fMapH/7LQ2rBhjaZWyJTurmxgNz3DJWcURtDjPHkUS9zErAoDeyqz7kfmn82q5oPw0SN+yA
QXu17ssRjOtjKKNMCKBD71StabBCTMyMQ83GUXvOfgVsO3AtRpvoonmWsJggRpV92xd5CEo+jZCY
NgCiXitEB5L1TcydUaGEMoct8eT6khy1vLXzDY9DEBI3ZGPTuj0LnybKYZk3DIMLl1cnNBJiNFR+
baSEiMsqL5+uY95WT1+OeC/soR058uPUzoF0EXrGbkNc7bV47cYOp5uZjA65DxovEP+KqSpCi8wC
fDQJZNSN0yTKjhiZT979Mjjd7CbN5dyVEYZs5y2P8stVgXXi8doLJzafhWVjizd917XeCmW8YJgU
/VdZRj9ZsMINsCtccLqIRvgXDPQciBLFtcafXIGFt4oxdhPWMyT4itHqk9wv8NwBurM//nGszDFB
71a0hQ+xkLkbV/LZODH3z3ci6oKwzDvZU0EpU1yLBafOZiap4Muwo36QvvUcPxnGu7ktziSbS+WR
pwGN+Wge0fTMUuv1djkN5rQHAYbBqT4nVB6QPrg0Eo+WFc6aRm0YvNkHhJ9Y+ipWRLO4KJAabQfg
ormvwhCnzpIgIydfIVDRjbE0MHg9ULWkU9X7rM44N4bCckVO4LTKFGoxTACZMX/ZvhoNXmQhm5gQ
5xcyM5DxazIP8vczMKDA/G1jtsAKi8x66zSuIuuyGyo7Mecx8xg5MAULUWFZOwWYevc8KfCCsnU4
N4sMjKMKSYywDdBmUBxTmhVoKHWmYkrbjleB02YM8vFn0osTQdBXmzqe2BUo+7h3gyDQuclmo3ql
ho3h3zFYJFvg9Z5hsliscDIv1RKNnMwWadOLRAj/VEZMGa43FT/FOz+45saP1hVIo28FzkKyJELu
O/6DeYLC7fiXGy13Spk5Xd6nJklIv/2az+T70CqWvz0WAHBMGOMc6lu0DotLJvX2IotVM+DBExJi
RDNdq7/kvUZ61eObXs//9V0y0Ca8xojE3ijuJZxP5H8g3SJDGgSkocG0e4xV8cn9iglCyqC6Soo/
bjpOQv+SoShreuu2WUjryyX+0wzfiWK2ALLkjZnLA9S6PnuErrxcGa2A3bhI2T6xyYElDBHwQ/1G
8Qd3Jk4fBe7OJAyM1lItk+OHD4Hgjb7TfUNl0WLlEn/6XFItNBUXBGPcDl9Zt9UT3ayIwJ6ckgvv
YFUw8uGPBgctG4Fw8DrykIyDSt27XGl53cT5uHTTnrVi3IevEAafrLS7nhOLe1Hj7voSz19qsB2Z
+gh1mDi4W4uUOiLRay2qF4IKeVg6zzavJuXkjgfyruI2Ebagjr+g/mhLYxU5UaKAejr47P2dC0C6
ZiaQg3W+X7jJ92PkrXVxxxhlMUC0XkRgl4n6JeMl0cakf00RT89LgNBTonIMWdwoBcPxyvo9cihm
3UxSicD/AkOSz3nuK6ckvCNcuHP0NVKSEWsK3uBgevRF5BKm9irhq3Wx5rQ3RRCk7U07WvJHckuU
6tG9aJGJf6LRnI8czDpT1SnOLN+fXktTRIbp1NqVq0jCuh/bK4+X21iS7YmyUIJGoC1/Om1yoYk0
f4r6fmyjpx4HAkN5Q7H7gorBzFWkbfS0fcBQSjy4cKp3fCjG1IsmoQe0JLiouz7wCs5FF7TXMuMU
HbE2JweSKImiE7/roneY20TA9KmKLjH5DtFYD5V/dW/LPibvOxGXijJKYJjjZnHbdBqrl74lCqDu
08RuEKFqX9DsUnvlB0XyfcsfxBcj/+Z8dHeWxNWfhMFhhQr1kkScOizwiK6H5DgYB50ReCFVxn+v
215Qj6FZxN920ju58HZHa1RM5IdhQ7X7yrRFTKsnJy8q1PRP02k/oZvF/7tvDsL0dZV18S3vcXaA
1F+Lhb50fclUVBWUywQo8LJREGwvEI2PchSAFeJncB5TjnPtju1M5FubT/R7QUk05NgP6mAA5kl5
JnNWEEPhUaAUi2vAjNcsHWxml55i+suGQjcvy8Yjg91vLVfdKGw+71zQVf43pwcEpfGGuU/mvIe6
/ewrWq2c+hyWPZWQVoZcaiP8GNLiyrZ4JO/5BHHXTY1QBLI17NtR5MCXDisrUPWvUln1bx5JnYeY
ix1J/6uvM4vbBPD4C7uzd8QhKTSZLf2akPuoBBtQWio56ew6nGnVQqa7w2xbB4Owfum/vdm9TBte
UgmYaB+tK78rBuN02IetS1VxI2/3eam1DajQfr8OCjmEzpFNbEYzD3Ja8jVkiY/Hw0jQHWGbGHM9
A0e/2kr+i2g3usRrxCaGC/voAQqKFOoYU5zsVPJMkgQ16y4CLRJDCE9UXacjy4XTkxSIhpWGMacz
dgLhOG4yDsucsmrvJdJgoQ8oI4Xv50UDRqrnzzOeqWuLRvK4ltrLs53zp1IoRoqAqRRl86EiQxY8
XMbtjx4ufXSxd17WRY2LccWEQRfTBHcKh8Loa61QDGqLEiTr9BMtOkuvASX6DzrUeIXPaFOhuHzD
bScTeOcsDokSZq5gxjwP/57FFOv5LYzH3Y2jHFvCWeIBzxpJAdNPQZXPHoOoBQWG2xq+UjrFHTYf
no9WRbX1DAK7ZPNKaHItiBMAhvtl1KvsYZJwNCfogJJFgW+7LJOtYg/puxK8K3IdwZS9Ph7qWQMg
dpMdULS6wws5m9M5YCVxcPoIZ/McTUL47EE9PFEtYYNNCCGv2tWovf0HxzNjQ8X8mwOjgKgjeTfd
KjjeUhfxo6kB6wiZDvioAg7EsyAkbuaAH29HsrePYpxdM9jnxeFOS6nQWzDKV3VzHNV2ozMknsxc
9exeetNjdSir+IzaBhpVVey4hzKTImZcTYUNBuog97NqX5cl8TamXXjUeUM7VTPXvNJ+slL8yTJW
WkKHpXSHYMaFB89x11ui2yjoLrssVfOe64i2KvfCTFM94A9WTxOG27VvffQqse5jJpRPmBI3opmA
vMM5yqbToySFInctua10bBJxEg6KoVagVyLWgtdbrOZHQ28fCJ4p/l7FzoePiHrNnU6SVnS2Rfl9
mtPldb4HENVSNn2KqrG1SLTc+rit16swleCDBZxZ7gYpKP6i90peek9D8Nlcno2BQm2HEZn7ZWo9
ogOmtDInHvM4+H94EheUSTgzjFc3fTRB4EO8iBG8VMsT4iKDE4QLVBgGq4hrgGrnMftY5HCfj5b6
faBpHUVQWqVH98ugHwxQUIhfFc7jBq4dXV+dWaZ7QaIC9vJYpNSVlD6i0jeSfLKGE6+BnmRzS0nv
QAWaoNoi763Eno6dMYzSSDwOzMbYY5Q60SKnXiA7l/cay7EoC68602qtjM8Uvvd1kJgWtAmd15gi
GtagkHdM7Yq9vC+PCz9VzWD96qMhtqtnYCJ6p68zJ91Wj5lfRt6MvforER9vDiWI9/9cIFssgwlT
iVKJ2gWLIwBGv5Ap77SRosXfWG/viu9LJ6m6y56rajvRJgjNuPmQmEbmuLgLfXt2lQLiMEZfnQLy
tP7TYVNBNkCLIflSzMt+rGIEfSYkKza/fYZGFYCFUCIR87kKJ63wtRNe8RcAhW2N/ASwyXxlWrz4
eaWiLBva1rCmKj3Cx3vzom6gGUU4qp9oI6re5xbeDRzdH3XQCtGr+ZkYmjiVLIqyJKDQcunTQ5mP
jxQYO+Zi5uEgjIuEcl8bCwmiqty+57r996amVbZt1b97RIe9CwTReqJEY4VRaB971bFyhKh/Izax
hbgaCYgJhWFBnOoyGkI+JrlmAi3M3YN5Qh3yrsNCS/djolC1zIqX0kIk+0PCX0D54Ow0daBlc1Pe
Y8kgaVw8d3kt2VEUgoO46dpv1LKHpHY1ULzdOjD+lYjvkzaiQ+NTKwfP3Zg7Mg+2u83AbeNmlDwu
ctxd0+8BSc1woMurSvVjxGBkvXBv3koy4pVyfczfRxUuPSbeXYR7jr4m/0tqgVx7SQ1xSvPFidmw
kauFw2WWB1b288EO9WPsEl7S7jlFhwGAygi4lyS7tMN3cuDT6tq7vIFjJLbmEBb+pPbEhFRCFjiS
pLGeffdvOx5WS/X+X4lF1xy4Q1YRULxwlDTqYlrUvPT6It151om9lwXgaaDlYUzZvPztM9QYXFwO
g/Y+g9g09wncT3pvVQrQ/4KkkZk+NiqE1Fc0dg+qZVu1NgnSdLRtiAHfZJv/4I0z2BEgc7hIZ4nc
rexue4r3IqU9P/xs0Cje9pYtohyR8wYyZ3/hMun8BDK+6M6H7zYpfrkBEhIpggJ082LIgoNlSMYQ
XhADKrGLVj4y4R6vdBYOwiLPWz7tuaKXZ+eZAGFx5mbi7QcwjwnZrRfHCh2/L5Zc9j/U5HAN3PTh
7mCcMzxkGP66ZzaqUgp9/EmbX8UIZRoQeMj2zJyVgMvg6t3JPLT4+ibnuL7shWb8ER49u2xOSpuW
eO38TTiKp9LNjycYBwQce/q15dDyn4sVGJ/gkErEdJZWLYDB6j2GDdJhzQSMMdEM2iu9qsmIKSoZ
FJEZWVDa9P8eEgJrhJACbcHfy4c8Hyzyt4j4W47MLDtW2MD3FQ0A/EMowX3CE5wjFqX35qcYzOJ3
CUswA2EWXS+9pclrSEylOeD5WnlfkDtHLGvtFLzjp2mJz+ymCVzgIz/sESsjFQADFbDOIcm4jBBQ
eiqaivFV0iIuaNBJdirgr7g4a0NdGOWUVS7fOTiicRXTKENWD7t/fcmt+nsZjHZqtfl4VLzm3Bb/
79lFvz+pI2WcErSQEAzseMGeAmLTODRhkbJO3XJGH4kZ1ruRYjXFDadDeVGAZBafE50/g2TRUXxO
bhtFtBQWvjMBRNKHDbSSH0rDApAMgufCXC+DIQO8snINUuBDYB3SFGM0S4zfiqiG+00c4LHtkvX0
416akYK1U5BrRJJy0iwFZ3aXyyZhOW+/Iylb/0b9zEZ3FgX1o6D9wg5QKbinBMSWtfkeKAobIzZC
VprypKGzKxOXTDXLjwu4KC1zszVTc0okG384mj/WMEYGcJu8iG6WxX/7tsMumonNhi+/s7CNhq9s
ooTyeXQXka5Xc+M9QlEXUJ5EmurD4V6j8zZXy64PtLasJVXFislo/SkoC2nUGb/u96WQTqiCKEYc
Gp6iA0HgUVntNUU+A2bDZF0JB7sPBy85lDD8igzlNAYVDjNH6bge561gY8ae8Lz7/lQPubUMldLh
T8ry4rRL1CAO78F7gln7/Bgt9U22SPfgaxQILN1jRm5wH2HziNkP18sPiWWMuIG/lYHqHeve49MW
meB0mO9LQEhrOmWXHGyjKeBbsniSAh4ugO0PH+pkpQAUPrUMHjwtCD7rJs3MaQxORmtD0eHK8iJY
kHie0aV8+xemWryeFmnWvyPPPTBRmantVaN2+adZl/Qq22SIlNyBZpjzXmjZVw4UKWSLktlFY00Y
Jk5k+OmGn3FlRjnDUthRaWI8s9XE9LP57LUbZ4p6+KpxOM1S5BIPrW/aQaDu077vApsRA9jAKbAL
rPFc17wgLKkV5XROL8GOSebU8QDe0wYczS/GJ1N1n77iZYcbQksoINUqPZp9tqKd8x4sYhBmRTP3
xpWw/2uRqpaX3ETRjyC2KaHuyKyq11gThBfffMvU30nIAeoptHrT+n6P8IC8MpvKT965t+qDvYYb
SmwVjYAEEGzZpMG2vbNWyzfEhCgCgrfA83q03WrLpBDg6sA9A3bXBUhH8AiuqBzTfjBbqAD0ZKEO
mxAGHKy2+zcyypRKlrhUch3kLwZT2SPImsFZYZ5AXu1OVYqaWwNFKBYguHB0ObG3AA8GgqrIMmB1
pEnLwMtzNHYp1TmjaZDbNOBpwh48oxh87hdIB8MJklqHRHZE8uoZaUzFmJvz5HYpFDbrLMyDsI9t
FyduvdiK9NYKofEWfmT86OWciJAWqbwK4+uzRUZnCNSKn3wabT9XvOjQ1IzccajIX7/410S1B2zQ
TDagqm/aZ5R9w//AkEBBFOmuiZvXJ7B4Nmo0T0Z/S++2KSVCkW5//S07FF/UKslYodnTWJOOu2zn
HxCwlwkNyotWax0e6cdghRKhUVDKHS/pJFPfBuHhj3QX38wRA8OeR28raVMXbRPaS0IHvfX9BB+n
FIppsVLnZLBdYXsy4R4PnJP/tmpGONSXQqvrtuuz5Fh/Jo/zwZVJeRpL2HLNMnD7h0ArHmHNA4aO
L4/o9FlmxDx2LkWVrmXbPAWxYcxODhdFpbEkTOvPPds5XORVHX2bY9Lh4+rK2hREUwhtzTZBnnQx
DvnWAmZi7Nx/ozETskeu2hoSKZT75lc0xMRCtIJYuud2PR0Veq1ojMpU7rw2ZYjMsWniHB5ewl1g
INxthY4mrnUeD+Jsr+kdw4iNbp6Fvy0RZLSWtU4CZWLECCqbWdDmaAA5LElO1fXfTL3/6Sc3oDvt
kGJx/6zg5LUW4cJlRrI2IIra0Sgl3jdu+LFMxo1TCP5FEqdsldC4iAMGXc1zC2hlczXOxESBllYz
3Mr8iU5gg/O0XrwiSREUcccqrNuzP1mhda6PJNeH/f9jV950H4EDXSigIJn9WLvd8Zy3pcPyq93p
bgFs4VwCVJY6hkj/YEMXq5doQ86DhFXP68Tc8a0+XvCOKqg5QOHLVbg57zn3X/pZdanWeMGQwV1T
vt85u9zOskIDi9eSlPNaHWmKaEZiB43/kT+DhWz5orvKpp2Js+hXlqCC/RA7dwyrjpkQi16PNCLU
x/yhmA4dERDBBnaJziLmMUBVB5pwhZvcuu9Ypv+CI90fVf9QdXDOFTXYDeltLSdTwHuOc55Igc9e
wUQRds7KuPlQErs9G0KqJzPDz1Txj9JPUTwfvskn6bbc3sDbFKHZL4cb+AJn7KWBM/6cOKlqTuub
psqTZDsAb8Dkov1m6ZLN4nxSRhVaiA/cI0BZejBnpKUCWogvW36lFwHOgOyWfTYUlCSs81pamevP
VmLcfG4zbSU+z9ZKOpK7usYg/qNti8rXWdB21/B50I9+OZinIVXPhd+KyUPygV/ily2SDzrZOpvd
5fCzT6zvU+bz1Tq+hMyt71lppvt1PSS+7JYP3TeG+Ab5R3wtWl/WesS99DXqi7yg/qydd3xwbbuP
GTiQNz9b/amXmEZVlqEJ+jjjz3vUU13BfmeDMBqTz+S2b9OGLaIxwAWw65ngdmHJGr+iwD7bHfuu
R7L98g902xDHUDoeFXtkHKM/FVIqAEIVM1P7AM1sGDOmPwjAtp0nMArftt4PGPcDpUGDGhDrFOKK
gSqpXxS1ZX5FDp5E1B14H8BQdEsgFrWXhptfww8p+YA4dVG9jfnxXiJmVi2IQF3TW804zdnsL6TN
s2Pp82RiCvMOHkfSmk8ca5AHw9FmcD4xIA7hE0zV1e8KgWgriGDccdzBTYmFJRtuF9Vsq/qcHLTo
aC8JuvORcRaBp7jXKjAlj/pYq781xTqmd+I8RE2d/aVnQdSiu347zCZ6P1DzPkrSRFPia3gLiHL7
iWaXxeY0Kc+rj41E20f4luF7TxtqkkJCCx32cTJZe34maRqR/gh8QZOHOfbQI8MhwPS74B0xjwjw
75qmuBHVV639OzUv67UZQRigPL9S0zvHltgsbPgFrYmVPmDjqsw/ZnZj1yx3P9EUs0M+zOnCop0p
5E8SGlqPiAAZaM7eq41oAm2O+fCvMlbyXGz138OysmwVvnIu2wLj1J9BroAE6zxRGW0Rgh35HBvX
ECIV7Smvu6TRxnypE7jO6kNonpRlGWI34dOTaBA+bBcT4ekb5gFJyOTJoM087/6cDqrwi7p70/4h
GIGDIPQ1gTmiDZtgIOJ8h0XSh0NiqWPSnpbfs2yFJKvDdl2M28nFqGUHmh4M+f8MsVo/edHoCN35
TXR7xobctCx4O0VVZTXPPCdx3/wRyMQ/TqnBtt7tMpGrpac9JzyHJO6HXVXL/zjvBS7tRHyniOPD
aC5xeLK4b1T8Uy4NLaPSrj81vlYredXumNNiSBvsyZ2sLZ4VtHyev3iq52ExuP2V6YSb8Q7axfrW
5e1H+HjeUG687hr89R9YdMltVeVcg54W3cAaXwXHf+rFAR0D+N7edOCA+m6ixb+M+MgFg/0KvoFL
qsezlYtpAWQiJTNIj502sDwoWog0IMcwojDs/RM73tpibyYO3tLutH+vr5Z7FD+7EnWNA+HSygY8
h0wEXS6zgd5QHTR6S/3Lym+CCXkiA5J+68nNJElM3mxIgPHT/ZbfY2qv9wiRHWTkdzhz6xOK+3a3
JgcTijbe/GcKxXATDBfxRWJkTWzJUKMFPZC5UgD7Fhtb6YWWTGUxecaPlgfJOlw70OsJ6YSAMFUL
YOnE86rChS17cXn/T59GK5vf9Cl9IoGQtSgsWlA8AIPDFmmpXFfMESvRF0ONqOOUUABI7yCxC1tA
hs2tZ5nWnaZ4agKarFO7Wv9N7N3zmBGr2G0kwFwuAeZCC2LmtpEtnxasQ7atK5RVr40WmhFyNiBK
Vf82Lp0r6b0+BzSgK2O8WY4v+hrz3sKoHOjLdiwLVfeufpxKvTKh2CxhB137/2gPT91Dq+54IQPj
UoC2lzndJa07usBR0N9eUmFXlzdwHiXaj7MVmzUpMS1y8lNwTbP6c2xiZZi7Y5t/8GevQKGd+Tfa
ek6OjZeCBhETBJlLsNNr/Bh8RoqXfozT37d/sffkLUdPRUVTlqo9o53UX1cc+810SsJ1ybnZJu/O
wZxIZBm2vQLHWZbZijr5gsfA+bkpt079ZNQGIMbuNrdtndziDD+Vq0f8SQz3hzF7y2pp5doGqF8M
otC6U2wDqLa9eHTl6N2CS/jdiOvdlmO43W+iizS387yhdPnpkECrorYHK71Dcal0PbI/UCuCyMjP
pEUleajVqPnKbCzZGdQvfr5CE8f/lhsMMvvHCX6lgEczBBGGGRtecICbwfRyWLVWYKRmXQ198/gN
wPS8iOvbJNhg+AT10OUISld+LGVYOKs0QKuFEgU/f0Cfe+L+j+yuCiy9KKBBOysljZ6yUTn1zHeo
P+hAWcGYafdrIpv12yposohfKJUb2ER3pr4VN/8N5zJ7L3rQkWLgzEWgCN1dFtwH1eHei6WkpFbz
laUJrVGDrDp3/1CxD1VYIlXgXO6/3b28qSluUAZ7t9dDAFltxzy047ZDUHQP0oxdkjt8vL72ihVm
4RQLyWnmB2OI3JjQlK8B0raEFf5+bZVAsXzvnxQlsW7trOqzpUmAcLb6g8kG5tNT0hxaIRDwSd1R
5sBs06mlky2fLQDf/1wQlwlo6Gda8C87u1LFG6YEFrJbdxR7KnhrdNJuRUbR1y11nRtLBHwUtQGn
uQeJT8NXlCOD5+dc7H9UcRUFRh8IV6hU3y1xjSVwIabClOHmr/0KedFQJ3WL8ADR9KKMl81tUd6b
e7h0QLnC7rPr3QtMP7Q0iYXP5M1Na3yghRdWRSwrAGMzkXvT8660B55QiHvvFacaICHF/Vxpdb9m
Qy2oCTr82vCTgbBylFFJCeaKqAn4RUA6uByOBPTQRrI/XTWXMXc7hURjOqeaLaxXkuKa49obMpc+
9zKw605+iHfed6rSCPgoO5xTIgzLi7ZA6iw4gUK8fIgy/4Hh3d/0KMa7CU6CYUDvMD+EhuP/HhOx
2OZf2kNDVMW0q7GMZ3+IRD6QULaWfaCZ+UzFk0aCHuL6W6Gj65VwlTCKEy99Z3/F8vFHL+xAppzg
kKcnxCicafXsv8Rah/WbldVt/YeKRtji+1MzjwElNKB0ehAtignX2eaTeEAtCiLQ3/FxKqw91mC6
vgubPQGv1lfpGn5WABP/L8oJJJzFv9jcHOO1zGe7kV/8MT3zffMuiy1OScObr3d5+DEBCuYdGarF
0OspVBeM/41lPi59QtiOU91+wbwxnxXPMZQSf1eD1Imq2guzyalFEDitpnbdC1FpbEoAy/1Z4ldB
K0aL1T/webfy/eD+b+2t/C7cLAHFV4uHBcxpm6ICyMu3wiDlKVc2zUFqnv8A88VhJRKkw/YhVDKH
fc0FBMR6MA8ICg/FxJ7huubZ9NK6p1lAHaFJ5v7ue6GxSibF26A7x+7Ujc7k+e76SJohdr9XvQQs
OEwhN/aaiTQQzwENCmw7XH8JrSOjA6Z9UxTTP6olHefqCbspv8lsxqebpbAbdaUwd1rB5mEP+bbO
oclc9dqwP20WXRQ0t5lDm09yvob/RCFmdqjlsL2trSnZ8sGzdVd1jPDbrZ+72xnmgAKyf5m0ilqI
kwefCMqN03GfYBkBgXiR9lun6ap8YrzV/+Y5zXp1rQluJ9S38Krh3bh7FzdlBLw4UdkMKSaPzeI3
Zs+yHI7oP/6EYQ4ZMoV1qNXfRrMD4w3YGvs/Inz/iArfNgnfZWr2Tp13fFAkmppYb2wDPZwqIiz1
b7CLy9D/1FnNYn0tqCoFrDJaNoGwBuP1xe3ZfXsCZhjawe94tAJI6CkFHl5SDhvyD/B2zGWRoXuz
aL+YYDNydC6fswxT9epoAJUdsWmNTdiXu44DjF71o1iAhcqbWD14neF0rgceIbmWNCthiQlDjoUF
G74m66j08Qv4TLrjQQD/og+FV/DsIy1epYZIBgYJjUlqgjRvOTLgYife1yRmiXrDwSA5MUWA0WMC
RzPCUBct68ifw6KiIRwOzuc+RHss6/u/WU009kt8Tlz2G5EjlC54ByvW9pX0Xb/CsJebJLOt4hZJ
Vz4Hylf1/QAvjqGr7neL5oNkQOHmq+JGV6IjVfwUxvGI3KVhO81t/Fgcwd6+TuCHewEc9HXtF57E
guMpVQD8MJwYhjaFlqJR1fxPmjVnO+Bjg5T8/GZCp37ZflvM3Wc/j9qiTVSXHJBKTLA+vAy28HYA
sndIun6xQfQpgr68rawPn6uUKZahNBbHCx5IeyjMnXQ5VsIA4Me8KMcu567giXU4OFiBx1C3t8IJ
pycspy/Xe8C8CcH30xIi5KMMTk41X0blo8oN5Ft5z4uDM1g3s80cGBimhVNMetdMkrwxzLcOW8ng
gsFaRdkyoABmXm4XD2AB8g0HWHdfn74mFYseCDQyA7LIV+1MgUYqTjgs1QAjNyUb0eTfQ90ZpF/o
W7fYEF8RmwOKRtFKJ5DPp6hYGCz9/9rqaCIIX75Ne772WnezpQ2k0x/xJ33jTz2LM0x3MuIJoXp5
xQi6jlwIBiE/zNN/8x0cy4WWTNHG0X2NRdaAE/QPUO6sqVEU2gK2V70bjEE0m4A4wPszGFX5A/Ah
U1gYrU8mUneG68pG5C4ZH9hF2IKK/Ci8+WEqiMGSaziU8xzwxYDOiHY8qm5+e7rROhwqW2NN6/HN
tbvuB0DVBQpDhOkDibtK3OwGy7ocRk4KgdOZPonzLMFbeIixU6X06TO5ugWyZZchdoj6zfIMajyA
uFuxz8jbko0fkMiCH6vDXGy3o25uhdWILQBjAvb1thmrdpgr07HfuC+Nr/zUzamkYPZvxs9H09v3
F0ywe99nj/ewdvKAWepCiz/TSmACmHXfwrNmAZDLjj1hxkzEUcRaFX5C5pqPC9yYRcfViQJArKeN
6GOCsK0YicuU1x4sPp/EteglV8ar0NlYllOTba7q+SfdRy9tgrHL7qTsZUZKo66SrrUjzlP51lns
EWhz+mJgaWVX7r3yBulnQdi5rRtpedv58flAV1NMjKRpLGdGRwuyDM1fTuCT76SYMY4Gl63Gqpkh
IOKGJqPw+p2Uahdk4//X3s5JdyKMbUWTj6yE/pGaTlD/MiYyllFarEImJR1Wr5EofEsGxxAoITmC
ivMq3M97ishGmNT0mg3J7fe86J2M+/KyvPvlF9FEqkx4kQiQBunz+TVxKE0z359z33yGQZ4ax0hS
+TT19UN7kPh9/4h/nlrVtRXc6TlE/ROT6A7eBaiJbSl6d2ALMK0ih78Izerk47Y8EDjcYK3wh0zk
yi+iBDJW3KpVtdZzenfoSDNRcshERyxIpA4hcL07iZNE8xJ3QCzOXB8Nt/+tx83F44yw2AeArQgN
wepzS6Wowoh+8YIxGpYfpUF1aY63e7ag5Umg5O1IUmcwnCG9WbTNopu2AO3GpGOnADfQZFg2TWQR
aaoBTZ5r0T36ncvz90tiYRUu6/RtoEvLB6CHYqyPrClwShTULMuROXOYdkSrLOM6o7iFzkxO0v5k
4oGtFulTWc5Bj68UtbH7Tevx+xjws7mX0T2IA8BYBvnKJvbNA1tsdTWtZoZrhOJJY0fgvMsftLK1
a7urfUH2D5fjF7c38KnveIPGkPUS2ywtI2T4u7WyA6O1oJMW6JSaZ1vD/5dv1yCvcrhxMs3JRQvf
NBMLX7uV2HYDDELaGigwgM+CSscXgJfF9YKoUS9AX7OydFJt7YEmEYbMWVKB7z4sFR6srVIKbGC/
N2s++HVh7ye0UO+PjINu7aIqhzHEwi5PslFOyRLWyd9XDvyzrZRsknR2QnjkS24W2Zh1Vofds7Zv
OQJLlRB7oRGQiMW1dQtiiNtC+DXALI0jtPIMl24Fls7KiQ/Js97esy54LNoS/GNGPPZWdz6gaGzB
q6DcjVE9wMJkXy60nIGjZmv44aVSCaDRpeWLk7o9wzZWedJ8TIRSD8ESrZ1nmnNpdwEIWWrIXGH6
rxz9c/pYuuMLDdjAE7xBqEwTqD/uJGo4ZrTNvG0E9vKQ4DhodHYxIk/WTzMvfqbVkZIyzzFad0zU
hIZuEgJZU4S/QfUrkSnqhP+8irXEiR4iWGR4aoIQ0c9s4KJ7tcub3fYxF2v32Okcc/aJRNERHjGz
gLmojjtfdWj/rzu4tc1Azx9Iwc+/jRYA6jdunEHIKWuZ5UIFmLHTBYPbF/qiG9u/uorT14u4yXyI
BGjJArNrBN+ZhigEjRchEyG8Vz5zZn65V2YevWkcujYMsVjTk/4BD4W0rbfl6eX+H4G8ykDdCh1j
2fJlhR0qC9uxuqeyNhQaAlTeuF7yvchf1luNaiMAlAeZ+QlX8fp3bSlNvSrX1g9Tdv8848qC8aYO
bpojApuON4/JqMwz6EtiunS1xRBbxjsE3XGx2F6iRfD4JPbraYo1veMCLuRqxGQkdklUTekxItJg
JAwn4zXtmtd3Qa/jhSN+UjmPh6ldHzeRRm53pc4JNserRkT3pOInhJVj/tnKyCUTIcQIUMuxnq+y
1bpK5SfSNvf8wsmZcWoH53nxoo+xftKGYLPRhzM71hLaOGDRi00mne6F42pZcTSVDm5NPZrHUHfs
Z/pxO7FHVOWYD29a+d/wFIJgj9vVRC2+XUvAuzfpE01otLkWrYjc4ulMcuUOOnoBucE6F19tefTD
nXmFqSrmAiKD47pWh4aPS1AYg6ZieBrJZ7yU4aMNe50CF7daKwFRwtSWdXMKK2LjaEYh6g6mY9+s
Yh0cwhQZj4HS7c97TkW/w7Fyx+yw0zphLBddbu4PA0oFGMQjJNSFfSKoHe1FCqeKnbukGItaeZ2L
R10j0QWPDzstS/7dnbwe3xjXXz3QTQOKSoxbKK+L65pcAFjaDqpb84ggnhyFGSEU1capDBWSsfc0
QKDfM1sClqcxw/XM91l9L5cX6s2QCI3koCKZ90KuaZEftEfKuXu+HKQfnY2FgeGrKwPwuzF/bNqM
AQddP9yQnDYpiYx9txVX1XWsVE3l9s4sMy7vrRmSbTnoSu6xi+PJ1JqKjPkqOv90X8NUkma+5vIS
aIEU/QkSdb8mw1eu7Z8yNTOZQTiPEZOpbf2fs5+wKDLsLfI+kogT8Hf7t2pwCbZiRakLnM/bUjDY
cEgVNL2DCyheYvVIER7h9sqTNG1N6MiNAYwnAqKhzXSJFduxOWa68INx2TkaJhPt++YSWbq0QCvu
IU6KYYW7/6v4YlQw9ZC35BGiBTqqv9AyqjnKOdt2sCngQseQu40WodX7glSOlNvts1gpVD4lIm1o
iFaBrAEAjIqownwKDAOxRBUpf/qmXa1J5+bW/THq9dDBuoQyy+TnJ/JaqnOFjEmUq6XPORHcTOiZ
fc8wowYF5MeaBEAGFg0MiAfZDvjW1wZdlFfwfCkGrSutCQVBxbg5Ll9ZzNipgG+GX0+fREMWdshJ
/bJy2vlqjDIsnquoQSa1wvU9ZWyfnzvqruUaL5Onu+wJFFaPvBnvLddgcwUGFbnIg0PxHfewOujg
eJM9qItf5+eZM28MC/k1CKr3VwU+1GoOgYXBIMKADdqre0fZiW27YMYxuPNWeiT1MHmvoPqwsALk
ZRYqCBTNIWVauqwzYJjP3BmQF1hiqk8s4Sl1Cza/rSqZ82+475z6BXki+XmZObbBKJux7CzaBtbE
otWNsI4J9XZr16w6JoptHF+rit88kRiVgLCIs/6wJt/31D5EAPXgfT7CzJaRDfU2Uz9Zvu3ywEw8
fqbOsTCB7uVfehVNn82sLHzIgbg9uHB+Spblrbtm40ijGy+eQS5zDnq2s0vL+zPa4ItMhmwvrgek
8kF06v2TnN//i2CSKDWtcpQI/yAVOeZdyh+YZ6qFNhQZ+Q/Ao33k2lq4om7afsRVQDRLDMWP2csl
Ts3uTsw1e87RwzbNOAqnOX5urN00k/BaBnYAjZ+ZJRA9DjAhsWAqxBYauMN3k+q+GR4ifmocwxsL
mJ2K4UUNPXd208wLzDOfkOPIu+/lejYPx/ijebQmz05z2eXr9KSgiwGTB6rRdW2QwN1HShD4bPA8
xKXI/ooNsqF0MlCXHHZFQBvhMdHWZVuLouZl9xIuew6lck11ViuLPaAjJEi4bEB9v5sCmPnV792R
/3B4ihr/viW1j6Y02JYb7SJ4QxSYgXSstV2Zss5LaDO7/1D40XTSj1C6zo7JaltcciAEdfZHd377
dQG0FnuCsh6/qyizdK1NgveQrpy+DsNat5d/F2/eCcyzeTXaHbZTuwmzkCM6tNE3t+lLm09TzoKM
rrsbZTZW1V7UU5dpN24s4yvzG0VF8SjPMtMvsrUhvJFzU7F2xXNNTscdxY64Czqas2EkjrPJRK9y
GoizJA1U4eh6w69ppQ3YIyDbsKeLTEJLAJqJZ+FEx5OlSsviab0R1XhHBZKUyCPjh6VXj6zpTAe6
ftRjYLTxge3hlRVw96lF2aOmL4UF4mk0td91MKPIenNLlATuf3OAHWUsn6diYUI+iYgPAU+zUj+6
F0o/DzYkm3or1cRGhaW926mbONgBVMR6jllClSu/5jv8wR4aYn296casU0sDmSY4i7Cs5W8LN2JU
GaCyWJaC1Q/RxYLU/4++iPmOjdAjdo/InPNsOV51dP7fDe4JGJADMAz91vzZSM2OXsUXTgInqatk
ZgWZ2VP/E2kNKKXX+uN1zdqVesKq4LUuv/84d6eoHMiEsfRCjFMY/unMHtGvtYxTt+gmk/g0QLeD
DMe7NdhkIjwtzXjBSD9iwHOYjJQMVGnEvlLXBmVlSUP/cfbHjAw1B/trVPYckz3OXbMeI6zuCDZN
IKl3YqT1O7wmI9NzM3aQoxFPFdr9bCFTYIYLYDkcbMEckAk4wda+Cp3R9us258ih07wHmOanSV7l
qZVTwAnRn+ipulvXo/tzlo4qR4xbj8x76p1mRgKlkuIhPlOFbQHpRP4sXwf3M880dp1s5NVC4VKL
LdvJbbJgfPX5uu1eAHlVHsjp8WbM1xDiZ9SPJkw2LtQZKtDIQ+cM29+LkCkfG/v4SlhBThO+JpUp
pURjr8UKK3eZBp8cmv6dq/FMnLFRL+43BnPHa065tVOZmnEJ7g+ZSXgVszir7AndpodEPfoCrL76
VEJCDRytOU4whUTOnkIW1kioStvE75PUGH6g4YMIiJziKw8BVbKdFATnOtHggBCuqahVRm61bxhW
5n93o2YrHrhgzneKOCsLJw83U/J/1CX+furLuObWRZO3I61iOA9lR5Lx6u5Ma12uED+3ko4Zrqfy
AFYCP0LjvVInxJGkdOfoBvnSd7lZoCFWOqJXpy7Sf+szWHV+yBA2vV+Zm4pYxTrWDmSRXEYVjEx8
RcvxxRRSr1Ck4wozo/LVwMWFaD11mvjcfxM6wAFTIt12CI7g9NhJuXY0AAutb1Z1GgvMDPtajimq
C7D9mAoPR5et+f3h4MMYnYAi6114jKyipzXVlIAARjimO80MJoU3O61Bc/yOVn0AwQ6SHjUGos8C
XYsoqI5XSZwG2yaluk78uueVtTn9taUkkpX31pf3dAEx1oOEyouZn+RC/OlUGycBDvPSwGXaM8Zw
+qS3+HAFfPQmUtTcOW2xxsnSN9NVscwRFNe71chgGFY7vcAjBH/yL0pPHdcO4zYlmbTs8kcFQX7J
g/mJIEkmFlZbg9eOckyA9MgUMHYYBTYNxmpQhR8iSE/91fVHzBM3gZiaDTNdZd1NI/mfR4NdJSVQ
e7/2fwT5WMLr/oViAhCv+6VqyHLCjiTm7J3TrDHRSLqYzn3uaCOumOnbc7V1JTmV7hYCzIibJVLv
NHvR8RKR4BxuPCg8du/OToAE5KbGdgrwNJLu6G/ErWwoOwlRMgNcVfUaba7zzcH5TlTKHGMxOK5k
fvwC64tpFIaCsz1I+bTxhOUbC1tfq4TN/Q+bxt+6B0yZ0YeO0I0nz0XbY8pgv8hq6AFfNjQnJ69Y
9HYY9rjbY9rfXS1P25AN06M0V+45qBuZ31DQmnAzgL4nNL2SSn60L0qod3MuIt+HsoTiZNRDxJP9
cw6mSZv481W05xjPSQQyabHqa10caJaN+oRMT8VGYn6AZMYATTr1zD4YcsatIuKECIvVjGQJ3lAw
JUCPq21ysXHB/WdtHyuTHMqrmB0D7YSTk2Tgrkiio/unDFfP3Za9JUSjKvDihTSqfEBMEomSYyAW
WHEsdi3ospLNTU8avTqh0JLxYR3I+g4s08LB+k2MAcVNJ44oLKiDI5t4VADk7q/iOuRD5O7RfPEN
CDmjNpXMvbzwCQlvQY707LCh3DMIDvA+L/BBArf9+LDSrQIm5JYGO8hV/ZdSEMJ3e3uDpdZ7cpY9
w1KenHemEWSaVTFj0Q1epQo6KR4AOwfsBTEHLLLFxA4WEo931J7NrJMb71bLFL3ZY0c6EnMGo1At
EXDHQIkGPmgTM0OIX6Crmn73aprRCfDFWqgO1uhmL5iBcuTiDWybHzscfSu1NmrYawwxtFGpL9fg
D1QKE29L5HYuqRgJ/c4Q8OMKszwY1LhcuGDcsr2DQylI+Gv4piO5Ni1vJaOynGubbOeOV9TxGu7E
/Z3tQYWQ45HetW0KpArMW0kEn95KPhoh6PGHtQLEyljVFo/0QTEwdDX3yEw9tiM1gglVUXWt5EBE
11fzhZ3+i8vqz9KC+sNMvbY4C0qDukiwYGgLe0Rx6GLulv5kO7kXpkMe6lmcsp46HnQUt45692qb
mqSDcqAVgo4MQShVS61YwDxMLgI7ioZ5kWmKzq9UNqW66FK331Co44dJm7cJhQQv3oduJ6UiiHng
Fmz/jCt12dbleeHYBHKE8jCiAwaYXTOC0CFB1/eOBQg1+huocbfRHZzjl9fQN/3NFmpHAswLgwqo
ubIS+TIFY6cj2U7po8B9iOUAW9oV1bAyVZ2lvSPAu3XNs2Ge4oRK6n5QTfLJBoRSZrzFpuRYSEbK
xbbp7XOvBKhbTW6Ayk8M/dByIwL2MR0htMNNtcSKVI0PIwfz8wViAGPWYJ/ar7oR+qBUyYDRVRoK
H54oIrsFD5NpViWU8v6BZ6Cie4ceOeBhe+PHa02omNpRgRXYLrd4MWLX9kVUcUHOkJYWWDUX6Wgx
EvDd9s57yoUYaH3G+/fpn26pqF7H0/ydcmhV38bA+t88E8LWfiWfTGojyq6XSAbd74sRaVkVXKvE
7UoWs4NTFkiG3uBMZPbTHKnbWrkQmyGWX+Ntk9rsSdxZ3ID7LO4gvYBaCA6orrS/58/C2w9a+Ybp
KRfxOpxaQr6EJyfO5NLQ3hF92F6/z7+KplUZA7tshS9K3yGPJ5PufRMtdqR3ZFaUxJ58BNgKyVo+
xrsKszPouvU5Rw1q+6V8FkFXDhwSRoD73q+9ykLK8ssn1TlWZjjv5JxOhL/mjU2+rqVHs6Obr9Zy
yH53MtC7Eg9uu39B/8Acc+nW3r3syR3Q9lWpeDzj3a+MPUrAh3FQLRt/kYymvaRTDDBBBbJxC1GH
g1zS1RA87tBlIbhh2Z+9jKptF3fam2fc+GFlxN8R40R7HxD/e+u5MBDi1FKMLwrz9OVBiew89eQq
hgHBu671eUoScSAV8ZH1r+Ch1Dylgnvapo8TZ68u1LssMgFgq467oAgCgbec/uubb+qPyq+afTkQ
XfWQkSQDrHemUwe6DBprDHCm0Gtd4QfUEoi7DuH9Qy/dfiJkLzmftmMaE1DySvycFSMXXh9Ll+wt
PViZgXrK0M7+rHdwySPPsJWITKeg2BTSAit0OhYsNoJn/qq55xrTiggB4LizPdBaJU0H1wBzzWVY
1gmjXviJ3tAZ4BrqDGxcaljKN7D8lDBCVjY6p1Pw0DAsYSyXBcqG/7jQCBLYvDTJEQTicJsAVN5M
Fn4g6AcQkJipxmqli6oXC2Z4yVwcuw9gJRGTp19U6tyHlRE9f2ZQT9LtEC9iS3f8Ran9KDWhsys5
E1BJmMiQKAfPHhGn8SVkB2bdo4CEE9biSTqKlHnwol0Hf0Aovp3f2lIo9hrMsZiR16SP8XPII3Z0
uuM2El420SOI3jnoxrAeU+wepToKQUfDoGtrNzS+0Wo0JS45U0hJmYeOIxtVYJNnk2DVi94ExlEY
w/b24MUtKYgrD5yairUq6pK+oZKh8mJ8dpCoQkPK74Ndi8yWOgRwAcPoQ2N5N9ad2y0NWGSYZqPy
eVHcSdVO6xcYjaArQDWV1CFDb9LKi8SAC7K6C589p1BtCyjVC80SnrQC5tw7BVPYDIm8wYq05evA
HIJTjJp60ZNrIJFDuM1AtJ1LYNji4NtCzQxQnCFMaiZJIi8jdlcNVUf72KOSd2vmeeFyag87FCLq
YA+pDwQckNOgyHEokYNFX5KSlNXqjWRjXfY+FLwrWMz/wF5h0GJFRNLnBldpbAnBhtKPbgbyeJOV
DLqmZW3QsXyJa80TYJkNtfcyPnbWwKL9IJ4tRN8Qsz74b7VS6TSA7roTfLm0MeczqeVhU2REDLHt
5V/rCYcM9qTxjzVLH5mRX94CY5xNbYD2q3Jfo7AoUAmbRyon3hGZC1+uW37KzJXKizJ6Lz8ONvHE
2mkpekxZYPmo3nrmSSbSePmdBVIHbiVlnYgAwmuvKTaY5T0kvV0tK1C6qI60TCuN2clD3Xmg6Tn+
TuCRfVaqP7YmSnpVX/4nC3hoFtJKklloJWiiBzegwmWaLOUoG7OCUftlnS3U+qI27Hz5aPLAduK/
eLSNL5JernSS2SXXZH92ZqdL+gtDTx0qE8kpTig6lT/8qhoJRNeZe/Ur8Z4SQmQ6rK0XhAYXnkon
ucgDDOszv850TrlX0jCwy08frmVlnNzxK4NNbPCr0fq4nFUfFAXRCwG5X7FBWIPHBwIbp+Yw2fGu
dQcGKEmvD18HDNAJvdayM+RIawDFFsTV0uCDqfgKh9CcZFNzXBc4TEOnogDM8BaPZpHYXOuD3u+3
qaJPK3H/svHz51YFcCt9iK0NKF+YzDwkYn7KI4XYYFQy9m4L1/YV/vxqiJXBwUppjdJQucGTFqoY
M9L6sb8zqMWpJnnbxSGg2ZufAgQlqncneCREcM3XzossF1UjLEjjwDkW2Dhr1RNhiZDAsXWDDGTY
UP8KTSYYbzc3aX2lPPCtzogJtORe3+TS4CXSZwmef836kSqq+4b3OkdjWE4lwedVE3Bcvc5etMRZ
MFXrROmsUISoKL2XwT9rPQvPJtrSnTyur4XvqhMrVYq1TsFsnFg2PH7J/u/Hh0jl2terxGQq78er
uxe7LIjlTFW0aR9aBKBhNq2VPkstYkFdeul6PQXz3c6gponzAIWtYpaXOOIqUPLLCUhaEkcJB5p4
ufHzgXgmCHDJlqiFph4JUBNL/5lkyMWG2GdgEElF+B279pYWeN60/G/PSJAwmYdVWeLlBV87qSxS
NKjUF8QRx5ZCAe54N4cd+XV70HYjiPwGSfyzHp2atDCTyy9bxoc3Q7ZnGvlaop2o9eCSNB0FAd8f
SOb71AcdzLa8t3l8YxTU1bqf0YQA20IiOh1JJ8aIZgz3aFeL4IbzCupojZqRw5oIhs9NrPJMmoZE
9sr/VHh94GID5xz4NqdaxhyHxVZhaEdgYlqxgKmUWPSARgijCQvRGu+/8kJNfjGMxZrKoKaBNYh5
2CFfSgoFGJCjO33qlDFlNPPz5L84ku9pLJhsuYdqNFd0RM4JNnylVvLlVTF+FT2g0aYou2zPQ1xD
vgfHyB22zZoRcro0yE8RvWJjeI+O8dgAsLb0cEKAeiGGA4MXWVloyb8mwu76oAJjJzPc2UEDUbuK
9NFss4uiFEkE6jovWZ33rPnwsWINI8lPD3YHAe6SXSxMNRD5J3v/8A1dPtPIxhJZAq9JxHBrF0fH
yeqod/9hOD3osfMvyKgWp+0pqKKHli8CILm5EEhgujsJ4BhKsoR3x+g3hB87jcvbyx34D2Ws08nU
FL9YMa2U2jBZQaXwg6TfuKGcKxiYeJ2wQOTxXJEKdy/Yyv7VSUfUmOuI5FvT/F9xl9m9IHGkaXlu
NRBdwiN7t0+oBrD1ssnLanC0TiUH8tF+I7zCPlMeFlwwkbw5zpJdvQv9Gjajj77GeG/C4oAOi43i
svBVW+iRvgpSwcTBUfo0qa0EEKVgSMsvan81opmi5d6RbbhtIAXby/KJFQTKwQ5sjmGuIPRIu0YD
ekFLy8gOkThKBq0T5vn8A6r4vK8vUK6V2LJdFJ7KQvkJIEPzJwsAw3zmPMeuTWu0aDgPXje5qm0Q
DEI6qF4e7sCkYKBLZy2QtKJoqClTkV5U3nRZAJg8ZfxOMbUj9CPrcMrbHrR+ChArIepLRAyKZwfX
sDuXx233sL2+c3cfKlVDF7RXo0ntSgi75uRaOWkMkWnqPaNDCXeizHagwm54KchemKUJ4qjYu1W6
r9jZ9zdhe6Cl8xTSskQkYo2v7u4kHVLK4baqe4loKcqOinzJW7WhxKnbOJA0oeIbhfKPqe294Hak
tnCf1ZL+kPlgwa7+H8QFFvYzQ3sWuT3OOZuWBF6MfV0uOV1VTTamxXhz+7ZoR033ved+prHO6tUa
k9ukB4P4Y8n43eUl6kGrVaISidKeDoHFblKO8g33zciXgHKRQh8gfIRz548bOiHnmNlrbtfUQToo
6xa0kQ55tgSro8SB0xOaxkixHCJQ1ZyZAZsF/yoVEexp5uMsJouDKRTG7Ctf95cgA6UuHePphCcC
FvKO9sqjTZUs2Vp9nNnHH3wL+3f+5pW2p63/NBtIU5+REL0VgEJ/QE2c1blg/yqM0XfcgCwB0B+V
lmJo/oKay3/oDVf85hzz849zPQtIIsRapkltlLDmisXxyBFXHV6kZF1v9Kbz7R2qncGtA0NJf3nD
RptZfz6/Syraoua52liNmTjQeoXYRFyk9y7gcf/qH3ubW8ztX0qOB5ZejKgzLwVaBlY3C+C3JFYM
Jao7m8nrU68QCiwd8idjE8zZWqw8sN/SsXS81Dr8XcNLnVRw1K6i5LaAc2TTMUDfthZkL/cgwRf3
VeWkTncrP7bozjbY1gYIY8tbJl8Lq9ZNK4LTSWPrP3miiQhOqgsdAkGzjZkGjVMsIRg9W/7m1zrY
AdSXwNYaWSevsxI0kSJ2sYcyA0HfbUuhknlVUrvCGCBW1qS0+m8Hyk5QSppvxeAcUsn+agrHDneL
o9E068INX6yWCQ7OHvS0jp3hSvWZx+nQeXkWsk5jXRYHADEKsxGVFD1Eh4kjuQjKYhqsXxrQED4l
jW/eBJjKXOAl8CU15aFYuDAtFEF0NHpRdQYUlOk0kVJWCLcD1iOD/mZdjze+a+qff1PB8+Tcn9rP
jZUYWUxptFWpcLCPRgmxcnrJ+l72UH3cco03kX9NZSvIrxEp48tHUf/V0iW8W3rd2CuZGa4Q62th
2cv0rtsGtROBk8TA14h+WophZnnL5HmEeNvXVqxgp1690FdjkikHwE//oL96H1N08M7LtdGiHBHW
u1eUnOc1kE0OOdptsr8GuiyjF13QGrmsm3HVcuLa30XBX8dpFXpTRdx/uRSktNSpTpiRqHYmgDAX
XPZPxlNONj2D8tEX3RSuETOVtvZbycxdxaTDnBjAz+e2gosjZzZKE1Kl/kOnk4LDvh27Nwj+1WeK
fkhEnszRs03J/7tRSZ8wupxGUPerzlQgWoCBRVyRw/S88mJJ/ZtYTHvnO6xPkaQMrhU9afgBlVf0
reCfOfTdkTEnajz434tAQSMVTtRisAi7XRDZNBRC2Mb7JNrP5rfuTwxcpin5nvsCguClik2yzM7M
r+zE3ozUHUkUq9yltcsReYMOUxlOHtRhG35HrXQGTxcRz2BJQ7fIYcf3vFqAGVOvZFkKD/VbwpAi
xQoUqEyUS1Vt5AQiNyoIDn3kxycvTpSPwNpLQBAroUL4jOLNIcrArkTsaCFaTIZjoZcIdxLyr2Xr
dDrMlxWx/ukC+q8M1G1H6kmeWx8EL6b6/9td2+GSpji7f+xMJjy/E8vo26x+mYBLzPPA2+Syo8Ig
LUoFweg3dASQFHgt/4HLiryxULJ3Oq0hSa+ad0/xW8cyfVH+gryv+TRxLZTmtF7nvrXc8+OATkZJ
9z1uPu9rpPezRyNtskV57EEV4si1INnW3FCtOKhnBUIRoQ1wbPihY07ZWR0gI7C0XiE70S5c5ux4
fKFIPE60WmF/QOzsW+VM/5v2gqg4VFlUnqWp4s2vtoFbpM8JV74EFueWVMtEMP2OF+rXjW891rvt
Jc59NCyZ2g3xo5YS/R+nuQLtJdw23noaskT+9EGeZub5rX77pc/pullYMPgBz+8xw1gArmdD5gT+
oyM2Brap/FhIzwuElq6n7Y0rre4210G2Ojh3ZqzZflrxYxrb7besaosqYUT7Owjx5aLIk5N2nlHG
bdhEmw0+AvPV1sQ4UfwM+6UiYxurbvkp3xeaeLaMNeKXQLmsfF95J1A8AMNq5TywKlfEP/7GBduu
He5Zzvky6MF1BBNSsGDpxyxn6z6SAV/ciWzGE5wQtwQ3FWF0JtPruhXy/MEa2Khx4ztjpaWtZimM
mGAHmO0yv+ohdWP366ozE+fK2HBDWFcJz6mXJyzX1d3J9krqNxSIr9biIM0sTaLrlLtwBlJ0FMtc
z36k4hIOs2uT/CmgE/fevsdpEZLj1n8KHgU4aHoCve5+Pyavv/q75O0D/SVz3vLmYEFTZOEp7w8p
0braWiCxjCAqd0cwidpqaPvuT8Ech3W5Nme4Fw2uwiOwrV4g1QgLiZLM2Ch1VaeDXc7xq6W9Eacm
x51kZGW6RNyrmRj8I+GI06pV6gxV59srMttXrDlmiyNjHxT+7EVZSksgpP3zGJBZgboBQJaqkdpF
lu6buz1f6ZRRf8FIbAwMGLg79YVP0kCTnBwOiCTnQDqQL98pXFJzqUEmdkkSnfIV9ZjlJ2RqzeFl
nZkb8RZNQ0hMdpOMr09pbIs+nEA5Aw0T5y6ntpO74ZTFMs5C2JzBRAeIZ9Nh1NMNN4r5RLLD5tKT
hwOUSbAhTYPcFR1tDcANGP29AhSUoX955fGsbIFJFnVxp5L0tnvXK3H4v4LaxkfNTI3K1briAP0Q
MLRmmzk0nxTHVwx8SQC8vGm4xTUucqkzcEoAJIGIVxi7l0QnEzruJXEBrK2EY23yVamH+q796ipE
2JyZ3UhAF4A9t1+dmxYw/qWFkvhnxmCkcv8nWwnXY22R3svsvN/rK24GFe5yi31Hcwwj/wHLqMTU
vhcpSu5zwfJAIbtmqrwxPIXafJl45lL/EbGStMCOMEVb2BEhN71MH0QmrqEQZtsATjn/nySvGXvt
DJR2/9ucArtMppu98du4yAGgAG3ium/hX1i+gK60Aa0AZsW1rWpojhGXwAyu75WyJOV+WEWcan7Y
aQyoEM/hamTtX6j+4sTYJQjfy62uL/0nCjsLAOo7ZY8oQblLKmE8vgGJLkNvy+xc06kl4J4sw+20
VTpqo12W9U0ga6dQKhZfZmI93Vb6nsi+THznqN3wLtG71YZ14oSkIPiZa+UiqiFkp3jCx+qoOfjv
g3djdrNFAk6yolVJ2a/lgr912gliqJWmiNNxwFfCfWQTinshcOeR1+L4BhadngHiGN372O16aS7U
hY8PiDc1WL+zE8mR2EPqFDuD53N5oVkl43FYexQsZjOXPR4mqfVp8rjVfGZikfghcMEHS/GFkbkL
O30gJsGgCipjavCnwsZmlxkrWLpbCXfI0yY76/j3xjNC2njqNqoectcgw4JJTbl4HGhMsO5LRJbn
50hHpJM/EFs7/NfA2Bu70VysIPJ2EQ5VC5N1FDOxr0P8YB0/IkZAs8CZDbx0mFU0mb2r/P2I/CFU
AZIZhDiqttlyBchV3cq711Jo1fWSpIK7H48ZoWSWdapJhQQL2SGSLtwSuQHI8t3CQQBdm/zZMEQj
gllltDL4nN4GMYJBHnxtOXOjnn3AXHx1p6o9Iqt2yKPMsVNlEPc8dnVFyCeyKJ1PORM87LaR771n
1CNyQwYvX0ffDvwDV3KQE1Wd0UTc8vmMEMQEuDFNLMuN63E6ZWUFrTWdsbtnOejcqqq/syXQAGow
B/Rk+JqoOmdggK4MBYfkNEGWUDl83B2u6QeCdSYgVSviVphZSa/v71vUVcFo47llRXvYoAMbHdqc
TK7BkyFwCLCdiShPfO8fHGL3AR6ZQoq60XXCTJyOM2JnfKUgeuAkVMVVpN6JKLyfGG3Z6bQpBGx/
v1qYLWjdBexHDHdaQJb23Ll7hLPukwDt1yHlfSqqhsQ18vRfu2fUpNKMdRyymb2WxoxRcLz3Tw85
NGCwWvnXzEzldx9FKSAHR0VRzDGqDonTwWT4blzhIJehHRofRb+xhg4Zm0Vdg7DWZcgP04j8+ARQ
+UgVeOcsPuQslExSFRd3cpabIctYQc64CUUf1UY/88niZieZzQliN2jhUyBG0up++HTHc+JbeGsN
anNIqI5ObHfnPr47eTXfkwA8nODslzU7NSD9cu/3TdA3hhpHQVnSDqxlx9rxrizAaOkszLXZQdZA
0Nh5/K6RzFFbLq4dMPPriRIqkke7vaFnWmmx+Y8RTDzVLzzaDSQlqxCr2+0i1RgqHHdXmxTTghCW
1Ntbr2rCx5oNd2UzvbckJ46UdjSz6sQ6SQ8mLQ5CjdTI6F7nNlyn3r5Jr8C4NcjQFvTlbPgV0FyT
wHWptHUCQUvd2vaTur8RP7ZsJak66Khlb2Xaq+Rq9c9tlXR35v1tKM0/9cRIrqvDk740NJz9WzN7
3Ado837rN4BiJsHSVwLsuq64ZDm5W23UHIlW5lZXdcndR9aopALWxa0GHzx+wYWFYZuwCrF6ABvN
V/NRNH6tAUJS3u3J50BW9DVrFMbhwWvt9TlLhJoKkD/KHarUhpHqJoopTTcUNgeB9TbVvtxejOcv
ghArFJnMDuXzQ9HRBp+nf2a2eLtcJv4KZZfr8TCBLBL9Hd8rrWtGeOMKfER5/snFzfOhRaIhbEKo
gpJ7M/JU40ebgGHfst7ZZVBYoDhZqdtux2dwnm5hpPUadKr8LeYzTnHOdjlOeRuH0ArkMjCrN0m0
r+BJPfkp8wSk22yQzrrvaZuvOvYIPRMjxuq/xccTvGehrnTObCWsnca2xEFuHTD7GFpiDlMOTi/V
nJVgQxzrIRNTcG4YL1EIjM5t7kHOWyrMVw7hE/3weObKnETITkRrtEknAXmKirudawNyx4bu+yLI
1/pi2farTSbumA8RQYeIsYW0uv6Iw1nA3SNYiAEdF3A8QfNt9Wq7QeH8ACvVFuHGhvaJ7HCzl5wl
h5zfCR4DYGcgTdMjexOylim223nnXy2h2wJlA/8nO8PUDmGqMR54YJzMWvSW29zF/8YzKt9/ThhR
JMZJvIR1MelftL/gqjmuJjxCAWmxW81JDNaKlXRoW+dyRLsc3ZAtxjCeDEhr7EnmRr8dWj0ckRTU
GsvNBRoiRHgGpeB7jiLSdqYhiXFSvg0bKCS7YUJlsQ0EIOuxlSKuNVVJ5kgTMLxvd6qiWtAqqwlv
VtiSIR9kLtWAlKiF3yF58rcI3jUNbRXKerQCJ7/Z3WDAgeAv/3JPAOk4ijCFQQefnoHDbylXLGsX
BVucZ5l6F3E95fRpJ46UjxfL8o2Bi34RCGuRAIxOBjbAYKiDujM8Ysi98z1TLslGgj6XhK0u8734
Ss0ySbeADGi3OAA3A5v+TnWFgrwvh1YZBtfxcq3zWd/nRJtAvNyAjvFPgERK+7Ynsp4MLpfA9+75
b4D6gyz8PF1Kb88Oua8Q/iwl9mA7vusFJrfWl64xTxA2ubVO/0Smsbos7lJ1lx85q23jU7Vww99L
Us5POp0Ct5xhXPy5u/dvK4v3kqm6UJ272RafI3+weD5pqHB5nZvzMvjbwhE1OHTKZSfrmbA+ZkvE
y49CBspMwyxnOLENz31EktytyWdoGXvXLuAhTsIKs3ADY/AI6Jsmin+kCx5btCzzT2ORcIsm0ySt
PqquQ6qNqRBuIPA4LZBz5vfmOeOqbqqGKk1WBbDCmnv7O8fmqq3bTY+0BTmgxD1CsfBLuqFHQlXs
7c1FqmonUEeybO/7niIPw1AX9vLRbLZrCDZvDzCQdX5MTlJPrsKg8M9+OZuLZKr+PgAmUcilybul
3iDVWnvj8oNfIRvhOa5gxzJyOjjLt4IRKRUD+Vpz5jyLqx8arRT52VWVLI0/Tzdnm6KHvJuf11EE
9PzOJ3y4kTvIuROMH9+Kc6QHJi1pTmAGA+pGHC7EW48uykqLixxXIfaDp6s0vSo866jUK6+88Z4D
o9WKNqdoSga5qX92CpDZqWagQoODg17YM4gb0TEPK+etZ+MeDduHgDwbd0y4J7nKofevee/0inuG
rjnlWMjxixy5v7PBFj5ktmKUjT55P4Bll11AfpjVySo8t7ndmB/n9UOggtMRpG0uoq5zgKHI+gVZ
ZPIkqrwcUkFrYbPucxLuCgNNZQ1YRL+zO+FHaibpMpa7Dzy658DlS4p2fmpprH74lZ7xjP63aKTw
/EW8yelpC2zHc3jpSOdhdhzFpG9ftFSiwZLnT5lW4SkKERJaPuC17IXuu7m9xdCAEWy9QDBmn2+O
nBzpT/rsxaVkeEBZe1Yn7ErhVrR53k0GHy0Xqs1DAFmdfFN59zIajNRiasyHOoaknUrNqAP80NLi
YZIbI6IRGGIxLOL5wjAxlA/rREa/R+AfyZDTORtJ/qRRjWsqIlNF9voAOMYSm6PzEAzilcdo+F9u
vg4JdHCvHAgQRSukEtt5rPP64d5NsVUZri4oup25+0F8StJI81TpGxv0wuWlfByarrcNX1BUBRY5
a6+378nah4U/ZHrNC36TJfXQKCyF7BKw9rCE4PkD766uu8eL+y9HNY9g9nqwp29y33j6DKi4zDGn
ZpifyFIlyfwxhV+X9/wAPDZJRv0RfzrZBmPdzRLBaXh8m8+Hlc8wnoFsUObLNdGUDCs7sqhVWAHV
A3joeMW5XkZXJLYdl1SzNsI5eQScDrtHuUXcoYAbANh4iCwoZUEGplGGzwNk1zCRrlIvZADFx7PL
MhBypqW9RvoT5dpX7IHN48ZDccofPen+F/DMaVpAToDiH9xlmbAn0H6SJ50NNul/KyAsPOjo4Wn0
UmhipIDqWwcTHCn5JUrpQgNRcRH97Fq+xB6aDex+cLk/2aDmLF4tPk88PEXVU0k7romRXuOggAJC
ngYcUfWrlaIXJuE+xAs4UTfz8RCjZAdrgoSQIMcx5WW78q2eq//4c/Gdaw/XbLsXenSqbaSplG4P
/79l++NOJR9OonehVUG3tPMxURn3RK6lz8IvSegJqUf5MrjzvJh6NWnMAGOqJqnj9vdIZ56QUZtl
/zKaqB7jMURcK5H9VDjk+0DK90EwXQ5wa6MVr49Wz4W769DWIxNSwxv5rYyweX0wI7Vqc6zSdN2/
VVXJjEuEBnmwANQu6ctwujNiSl3KBtZQZJv+MpUuYo722COmkNHawsB1H/vsqyOyRqAng3K9umKB
CKweU7zfMAmOJEQOsF+F1vhvJ2JtCBIjNzjfNarW0lKYfU//ts0eGQujHIjXyyrnwZ1IdIwU8E48
neQBzGAH2sVtcioAJqEeX5V2ZODxrHM8UvomXaoKqEZh/7z+qJ9a+OC3pcfepG11ztjbYezjxjkN
UrHzJPL+u22XAquU7DZ8mL+8NTc+J1hbl41/nMmJkcWEUJhqdNT1pP03Vmy2qsaGieTsFgcaAuR/
/mni7LTAc/hBdQvpe2CI0OgxfY2Sl26pWuya8i+RzKs3RcfFoMIKB66EVMienlKeWmou2QCJh3lW
/6GdqmKiA0ew/6wueAVqrfp5ZMo3U6I88RdZTBzlKwJSwm8GM7aIyPGr/hpwNg+z9PGObNYgo8Wm
BY5fCcxcSr1qfRsA/uFCiWILjCzqIeU2fe0ZIKqHS9yzXAegxCWtFt8FXlytVmARoMsZcWWMR1hO
J8gqC7hMZDS74JqeJFOEmHa5N5bCmxMbsFIu6MlaFqRNPO5H7AiVxDDWLqOHGXLG807E8kypen3s
EO7U5LfAi9WE4N4DyWbzbKKSRLd9hCIXAe6uvjVuRp3zT0KhPy/Sytk2nb4UHF8tMcfPFsSwNebo
0sNsV0x5kSsThzgP0QXa/UDmR5kD7HHPwGLnitZ5cRiisWKI9i+WXEg7ycwvf6um/TNGMXDHH5rs
fi83aiT0GQIzcj3wbKyxNFEp2YQpqpPqVvMdUz8iLT9uWMqiflclDNW8XXkrm6XDsuhqcrJ7FCsg
mFy+TgKkTlDaPxhp1guGU+ZFPxF020Rlt8PaBK8k4L1PkxRBrfIEVPmS6NRjFaZ3enJPbrHpvmjp
zQ6X9pJFi1vXE5VFehlrtGXwSg1EzIGuIRnon/KmgfpNV4TF5asPNnbY+4W2ixRr/dFoUHlc06zP
gvr1BZT+LAg78jsRLUByvjghfVt2Tw4fTWT2bNaJoz0WCyH492aVAnus0T3cKnkXPZmDrh7iTrOB
WOlgEwyI/9X7pn3qE+StkKOBkjb7ofpcmyO+fyuhHN1towQFpvIeSuyHL/+4rAT9CzPJ4ErA5+dm
6mstljK9OImlyfQ5zoub/TJdr4h7jdgEHXjsf+QMamIpOyLqfP/1/Dx4k//3M6KoxpXMMHq3f90t
VKpEj9TqYhAE3W7BUH6FMPt0sLmtWKw9wwbobifsnd8JYToA0OUFwb+Ps/WFP9ec4aCSYai0aQLo
L+5Vqz14CDYksQXmfQpNySjVNsAkVpKp6fwTRgnZMzdgeAIMUv9U9kVVt2A15DxYGT1wTtV8Vj21
Jsg1U7IcBodqdIs+E8s/ZkHhyDTmv+Q/od6cUeEGfVdAT/cLFrgUdP6wvRdvG5OScft9tqM0pkji
bj58/301Nbg3nadBw+5kdNfSWcvSSQK4G+wSuyiIRx95jMTF81E88KtQ7BVGD4Jcc9oIZ6x1biSe
Y0JBkbdt/Ev1qVlTR8n4Le8a2+Ncqi7wQ28Uf6pVD4jAE7JbdtVc+dgSNpTyHGYsDlk7H9/qyMld
pfx5cMLhrbONLwG6914iTtiZzj31xKAhsooxb2hkfLjk3F5V9H7CQi2Y2Dy9dXoS2/CXVWNlGonq
USFF59uWDHz/YMVkD2GE2kCmm4IPRmxZ0Ytypy/BqEkQ2Gg317jAhJkh26nooS1iSuA5YfvrLwlB
4xfYAum6M7+catSEhaDU21G3hz8f/YBpBbEM8BQWBZoD+LbR11j6VSC5a4BKDFe0hN9RSee9rSRJ
FU7MHKH1JbLB9hPcvQDm1EZwO28Lb9cu65Fv0JdOwY0KuHwISRgsos4i7x77EdJVVTO6Qch3tFC6
81LDY7s/ptbWTgGqRnk7h1G91F0O9JeoMa7lONSUw8mB10yZJwCFtkmm9EmiKkEEzE8pySR4Kz2i
5nb9Xsr1jwnHKhX8Y1kVpO1esTDzXVoIquz5fua/NkK8CixE+kpoJyWyoE09mx2yc7nonHObn18U
pJwJgW0M49GrY1Fqx+0ljYa8cBndGBjIUyTJ7iovM0+0SjAQiSpEt+2THpnYHeDyF4pW1jwWkl7X
qIazUiy+lQsz6mRa5TxSjOVfOju1gjfkEQZe/Ii46u0CdnQuLU++HTLsFlT6MkXqF4S26sslloua
4I6OeowNUUNTFVA2DXX7jRN/ZWge0PA+5nR3iDBylVK+xkclEAX31L0J7L7D+bYrQpt/C3AtCWOz
QDRl5eFJc7NSt9LOfRmm2vcXtMwdI3w41Dn7KONYPIZE60t/wJrYSLo8huNqyvULQslhBiJ1aONn
eG7Z+7thYbOzXgZ7P0s8B58dznUY0JOanGf1lMLGhrHQRZE86IHGuWWdZQ2Yi/LzNI22Dr/7SURa
sgZwoCbFgXr6xlMihObVPlom5nVlV+WhYyeeQNf7JF3j7Rd7eTjXUKvUHgvKORWkJMSL4SZ4a6jA
Q5Ihv9hpaNxVGOOEu1aK1T+0BAR3FSBOKDOl83azE0CaxB7MeSSzRm/d/48b1t4cnqhxo3SUXue9
uzA0QJpC2uKOOVBdI6tbXWeMkVPK1imVgRZ26fRcQy1rdLuakpb2p15rGcDZjP9/sqdcPtcgSG0r
ED6v32osPr/2FmDfas+A1MXqcvj2PPQp1t1lUDAS3uNkFV1dvWjp/HoxDnD7RiNXgpP9jP/25rTR
02VMdBa5gukNnmdmyhDygaN8IzNC54i19WCVxcR1z/1vwajj1tqpyd10vv+3NCGFRqtV1X50kANT
w79lWi4Wr+ZmhvLYWqGQLrkFG3oqW0pfuVL4lpvL8pVIcxxTJejfehN2NGHq54Oao61SrYP6eFGR
XHxBfLwkM5Z6eTiMtmun/5k+xFNt6QX6OalAKNgXKLZt7dP2kbuaZCker95CUya4t4dbxDLc8g+b
2PTsDOs8IqzbAZqxiL03lworim6lMHHmx/Mp8Z43CsRa+6qETrksYECgpVXqjzhitn5JKqyCJo5+
s84YFJUfz0/9bdnv8dfZXhEDN49XvuhZvZAVOwI8kgDk123eq7g542GrOupE1D9IUNIMNkuykF4j
znwHlOBcd1gxhpeL6gGXvWn5ZAOyIjSxPwc+NO3d2lAX4zp+8XN18G5I1W1+xSk9Y+fq2b3HNIRF
BUayz3M6ib7dLS0ImAFnUHjiPEdiLY6kYTccj5gMFY+ZDiPRUt1yzDHIK2DQxqxFopaSfzXKwbhx
oksBa2AWY9UDkYwMhNd7QM0N0R7wd959/IjsQ19FMehRj3eJCsoldaSenx33/TEWUkrKpZ/3cJwY
Mzll8aKGuvAXdk3zQNBOc7ROaorP02vQj9WwrmCC5+4qV8wHOEXuzvbpNXykYnHm0jhqqXWMMjtC
jv5ka45axIXmvtcAptWtWmRBAuHTbTS1j+r2GLtr/PtYngq4b0E+MBSeCUGYuC5UUjezuO7cd7Fl
NJbUGAfMPo00HA0jUw4ZRDPX8X8ERusf+HPfXAIC346TWVzOUrw9b/oP5ewFvZ+7uixNnAqZWSNG
KaJ1ZMk/d+n1beVl77Mv93zUn0zoO3GOYBZpZh+Klm0u332wAtNyEO784p4ACTvKVXcpV9W6fnfb
EqnzW0ehiYkydyWkBkSTCBYCKsuKYDxltkd5Dy0K8vgUUm0Pywg2rMATSjATXFQ1nHRS7svcyFNF
mDwRvV7C9a02xnJVSQmrlDkYBC0ROScg868NAaxUpQ11IRvcyuNE96gQRFI9VcGSo+IJWr2SfbEO
Ay7jszXlliV6GJXo9taDeoiWPpbBtfibcm/oFsIE6lXU8bKC1omwb5pJrJietp+7+vLLwdTuIndP
Nh6xGDfXSS7nlOJaZUCfv6oVDUvp1Cy/JKuBXL3c3Pv0aU/GUv9EHnqujbe1APRmMxSo6b12mpil
FIPWUKJrigkEO2kjJ+kSB7qCH/D9HBoNfocdJ/2yHqEQ1D4V/M5mooVCSNDF7pbkZqBBk+G8MZWm
wm3Aqu06vIEqu7Jg6Xp2XC7RB2WQYADkJ8+0MuOpiGkiX/Z5ak9QtP0V5b55SOsHPko0G1YFJOiZ
5wiumPaVgz3+mLHUYT3EswxUTXLVdIilIhORN6xbrQ2YM3+wMsXYVYC5XYW2Kf1z8grpy01YPN/6
YXX0g7vpcmJb/6nAj9bWYSnufKJpsUPt7/qrL0YeT2HF7MISoM7JjcFho4EsPktHDJahLX7v6QPe
rXIgLwIU96BjpkWVtoiToYVStbb3gimHzy3kP9kpj4JCc+R42W7h9P+6pXOtFjzcMD3PP1cCrirs
LWkxKHRfiv+MOHabWU6YTXdWu41uyBo6diRWMApjFFcYWbaC5z8+5bk+LBJ8IvJwvO6FYEYUU9oF
Fu0Av61lqVejMdqiTv8NnYk3CFQcCmpNONjv8MlbNME73OEReyFkmyInJWRkfyz3n2cxPa3TeHru
NEh1LOQS3Ii0bTa8pZvbo+Cg0jk+38SHsHJAxa93QvOzSeJ+Ed33dV7IdNqm03lOMcfFETRUgcAW
23lAgbK+Roa6lzQhUpAF1Ub49xRU38dgVBDkDTK9e5V0I0DRjWElxJFVOojZN6xYQOYHTnv1BvPf
HjBZfPdccODu/m4cheG+JgE+cK1n4nYCEnfU8xi0XkD42wY78GEZHSCeaLvtA7w+Ig93AyG3VRQ3
GXAhpd0rCwZkR1COaNfIEzc1BbPswSIaqZsVgd4kREGzZp+DkVnK1PXp0GcmJWffrNgznjktPACN
UGIHw2qnG/NupZvzzUs+CFbtSlFgg2+d0G9ypG2/dK22s4KH83HqUVoAvCfu0K5Zz30r0nkTveUg
sDHa/TiIrs7iRbjt9PqIKsFR3Xl2NJOgWO9rH70Bk51V590gYtRCcd4pUeuPNjfONNq9HWykhEpV
vFcOIalTPbp/3ac/7z7hf1Qfn/jOFi5YP20I2MSDweSDRehZrFOa9QC64dbIJk8tpBlKJxKKdaTA
Wtut9O/Ra5PMZKjUndT1j5TxRe+q1t36teBxEf9ShelruhOaYN1brhz75+CVFHl1eh3rd/jJKgv4
2pw1I8Ww8+gPYNG0Qg3qlSOUPvh15zbA+DVvs4WCbqpaMP7DNA4RPWBymnRdi29gREUcndqzBEW3
CMxc7NtE3jbVLtG6E8A1ofcq8yS8FTXsirRCjXihdyKPXfaEpRqmold3sSxp1ShoaakLErKZqQzT
jbF3i58aL0P+SkYLw4QECAVj8NfxEihKXKel4i2ebQvTBBuFR16QduHkYLlRrhpMKEP7hrNSFbFh
kSmdu/wwpQ1LXPEsttDxyVboy0zMW0tAEDn4seNIiLLzEUdYLzHcIhlpQr8aeD6QvETK6R7K0gBQ
2sGaw7H1NZJ/DTGiWpjXV0MdA5CqOpKu6Mm3f3DpDz5UEum2tatfsUFIU26JmqMsLSWVxwHZdzJw
Jqu9JnbAUzG0YMRmRTTn11z33KjStokJlroVShHCuGVa4qZIcIob2rlpPA2VcjDzsTYsSnUzmrAg
jOM2Ihf4ATxad/SBasVuxbKcYK913hyzCfQ63kVB5ryguGOGPbfKLtXIZCYpI5tkRCFQAd7qnmRc
/Rj+3+2QUL6c/dPGg9c3tAESsd/LE/gVgudaq2WjffzMnkR2i01qflZnXDtXFPrEGMZ0uVsINP9+
LjXZW6O5jlh8SgUFa5omE1muE0sdBgB6sYaoZ01l9Y3aEaNpz04fUf18DxiywE8qWEbioCRSrTlS
kMdImTBBZsiDq5Ma0/bbbGG+s9BO77DiA4QOzQ12UfG9DCWgS0yjhAyShRhmXLol09XxNkHDEX5o
xycfjRqeVteCEHr4x2YBiYjo6VCudW1kV70+Zaaq8GPG4mivV13cBPJ2Z2UgXO7gU/3ygp9mPvTV
/peLGm3VLGrMUPFIlv/9IhMH3xtt1TnvUZfXwFqH3X9tbfbGGd4G9katDfcBv46Y1D13rGk+v2HU
rzOrpxllIN7M3KzaWinK+lrSQ2uvQBf0/pNaTIdI3jOypPLl+CJgAf/Wq3Br89lCtxBlr4Wp0fh9
6CbUNSf1nIygGOoOKclWYIWgrmrCimpfOEtAlN1NXOLzlbNNB8SCKO1mIDk5T/N4qBu3O5BOy0gP
bE7S4eKebfymEWq8TD6oIWO75zcwQlot2zxNjimtpERzll1X8EqDDA6ggZb6X+16pejOAk3cU/rj
2PWn4dHlQ5pdiQonmqAEyxIy7pasZ1+ywEQOzsbBXU341ErXoIRNxqqLmLF36giQ0LwrrhfCj5OV
C8qiF+E/0gHXQi8bKtpyOAAhUE9+xHulba31nnbFvlTfUGEqSKck+9ZS4zalrkdRm7EqUi6sBAvF
le4JFqRfqQryPkJlHqDPAKGnJByMJtocaIuMBHtZJu2N9NLzTJyInM46+t8rdB/r+a5FZhlGGsu0
KxSd1IXunfcBfLdIlkSgR834BrVJII7vIoBtUTB3YT9f9vVtw+pqUIu5gY1ke/lZOht7Tn0lSQnB
NOy7m5nf/KA4DOMZOU+09sk68J2ca1ReyJdSE2rdGwsp1wvPpalxmCjG0vGeHwExkiKKKoJIK2pU
0/kc9TKZEhQgAgV7n8ZloJF0TLhSjEnsMqo2hVpGYXAw7Qcslwa26eHL/3e5wUS/r7iOLIcH1FXS
V9Nx38LQee0xyw3qQz5B/Oe5yTLdkgsXCe+PigXRqnEqw0prAPCJcHodUHXvl7g9b2TYeL8vK+k/
jm3IUV0Mv1AkSXPX9n4/B4xNEyaz6sJRx8cfY67cWN9NvLYI4DRKxxC0r/NGPoMkd/Id5kfxV+M9
04wlcD1z1AAX/HG1e8NqG52FpEKAYVl9wDu5/mLSBVhNd9wkDFFb515b8IsgPpaN8BZO9Z3tisNH
dpySYdGu6lpID/5n/5Igo8zYsO1QhOGnG/wELasSaxpZEdT/xBcdhIeuVuX33T/qXMbK9UV9CF5U
bCsRl1mPhDN0SleMgbQDAeuhbTZpnYhZ6bp7HQ1EALJ6wsbF0ou7mmPSwMSFATrS/l3sqIV3PCwi
ENhYJViG1mAVSsKaBOXrKQicbO9Tg0OIRj1EFuvgHvCqZjGi7FAbcku6HiyWnDYknNntZBR3p73Q
qnmjH9qM1L8yM+iSdthrY3/G3GVQImnhb5lOVJkwsceo0wGsA9sIy3i68x548NakBe3f93z/l13+
tP07OpzX+Egj5WOu+hr79k4B6HOfRggzw+K42nDanOt0eUbPsRmFDDiFvnKWTwIewppOsdx8XjBJ
kNXjlHqV+I6iRfBR9gLAKcBWIUVej2xhoSXtFcyO7Vqym/BIPqNBzeE4ZWXXYC4N5FXWqwZPpvy6
Zlkgx2nbdF+NuHc7y21gQIWL0othyk2W1HVNMlscb7HJLtWNtJYWrz0jIxXgwRngRJ4VDXWwlgwT
3er5gt2tqOeU42nV7Y2Yd7C0P6/0S8l0ZfCJVOoAP7zqbxs4cLBZrx914lAishCI/ZVsJkdajbWr
agHp24rj+dF3aG792zVZTq3b652IwIx/YQMt5KlN6WnIQRcdkZJn4uVGs1YvlzBZ4F87Y32s/Riw
ubhUngq0Hup7v4TuU3Bl0Gkg++VWV1GjnXjZ202joPSIkQMOuWKknEtTEYc782keSlQSf3qQO5L6
vhSmL+NsObJlQYK0uJQDXGYstvJu5Hhmosz/pKRpsqf2hxrZ0pIxnOpJ/0bkVWQET4Uh0gTsXO1e
b7f89wJXiVBXi3QweADqsKGoFip0bfsseN4PuaJUlQMh+XDBUGB1dzx562PzJkiumcOQNNOdEA1q
Av+BlhEym2VPdrwp8S9FoenSrcgF6Ps0DnNTme3mKc0SJJl0e1GAiJw/XzimKCOdajPq0X1hLIvU
H+dEs1M5MFwjIRsgKdrOEzh864FfjeEGnMMf7ZuDuKrt3UBW/iJvH04X9NCx3KRXrIhdMqk1FU77
jU2lmZmSDMbr7nRDpTM9ICE8GGLtHTachF9EbxeytLB5+hAqe6kZptm9kgV4KAucGgrssCm9o4S7
n7NSKTnMDwVJycEFiXsk4+ktEz2iFFP0WcG658Sr+0TsqNDjNhVk/wMKNXE8QfC7sFxjOfV5DzTN
8N9QNLWA7d8NZwN1EoYI9yKniBuBvdgn9OXHziP74Ozb38Opf5cDhU6N83ICIDzlxNAxcrLBOUTV
rCA6AyM1iBkVAbpkY0ORtn5du756QtH8gpvESFU4Pan+zwvlpW4TCKhoWDTh2hRwHZsnSDX9AeXm
6SPjqqs5WUXzs5L90GCQ0V8uLhMOF5C3na1dBsX8LfcVGTaq/5do/9dRjC09coRHWGHO6Zz2ICMv
uX7w1pSM7RA+2soJzVdg5yYg3TqmFuXQWc0T3c9KATfmgbwqujfANH9f4cA+87Po+mYMkIy1G95f
SLM9UMIo3qp4myLrEOwRU2pYi56DWA0oM7sFjcPjymBqYFcL9nSsKFKbNcTy4FQJZyTPQbnXhaqg
aSohzlkQko0SwUeBHQTym0toL0dI/OJLuPG0pCz+3ElPDgTs3M2lNMhGDVafgagJ7tc3JDPRTSyv
Z8xbTSTr2uDQIN4cC1LxlQ1bEVtJz1avjVhQ6UKsPOdAinXjOvaQHuTdYcDP3XcxZFhoiCXjlUjN
I6myMbXvQ//ZqgpHeYhsHHtBeu+TSqAzET5cWg/FTGByJgvhVuQ/Rtn5NY2tk9zwn8vrmgEp7d06
uxzKsWBNXHJEOuGEVPbSkM7uKD00CdLE9BOMmYT8mQ3krCeyujwy4CUCwkPhIp1tl6MEYALSV/t3
eVOH/Bl/O/kCN4zHoj+KmoM0iOvS7qOSWzdYAlpgu593kIEH65BWpjxSe5kCgz1aukbhGyG8a8rD
O5gsGBi+cSlrh63k4JksJVzEJelxQ+Ck2NG0gpgqOPdz0tnz6g4WHZmxbrCW2rnbjkdutFLT8wGH
+i0QfEL9CjovH5ZRbqqS2b5ENmvt2YsI21iFugIBsdrQ1tsfeXO0xbZm8Z3k2wsgxZrIklRwW6SW
fsajJtRoPqRkWpfKUfR2DHY2mN3ItjZ+nXRIlKB4eEiJ6s2elwXfKA5891i3ijJIjhGNnRDN6whR
Vh1pio0XVO1ZMhbpWoXFMk5xhADB0tGa1pFoTbAcmr23/vazv2ST4Eqns/hxJMq8Yxh5jy/mjQqK
V89D6Qx5+aNmEv3RHyqHl58e7szLE8NhX56Q9adcM/0j6VOWa9fAWmUPp2UC8Ozwd1LIHIWlR6gk
xJiw6gpEkd+Qcex1xYJnoVINLAwI7d0KC75iEGf02n2YnWOginDD8hHeJsd3yrCem8j4EOS9LKh5
ab+u6yvMc6iaXsT+/d4i870muexU2W5sQ0G5kz2J9lObdPhv87nssfriBtMH/61YDgQsaa9jHfq5
7h86Ivea7po5Sa0XZBm6Q80bA6ftUinWdZuQOdAvUBSEE94e4ztGMeYFzM8yP3LSHloQdsE/yAkW
nyyv4lzG4t36YOgfTuB0Lr8om1K+2LRey1XqxrcpQdBfMOk2hahcHar0Tc2QwocNpnRRfiMUsU8b
ThjJzzhV+A3IBVGp2whuNbocnRStNazgsblEyKdBmlVmXhEUyyGksF1ZzWqz9jeJn893OZEyRkcS
BXfxxt9ai+V3+IPug8aK80uiWzLsWw/kZlT9fX3x6ZF7ZgRqk32aMnYDQ346GuDUqwd+8ky0Cp9N
XzGR1+PitOScn3Zn1UwND5LJkZX+eDQirrr+vvVGvf3/5AimylDs4U5qjZ1PgKDaatodJcjKSkl3
wEiKrr9xeMl6ACOkdkSPbpH62WyeneFn0BZPlpoQZsvy0kfAO8s3gQLMHrDCmU/BdWa8wdjFMJOf
yVFEDthLSaCQkShdQI57AnHy9hr+1MBt9JZK+rT3sWp1y9ESGrywDpolSdRM+Mdg4RZMg8WvOZeI
3HpRejDejWuiD0uiUn0SjCFSHcdrifk6sYhi1kiHLO9kyenXbRTzrRqk1OgEaWHGPEf3Qsbmhjvy
Ac2MJxlXp0TxobiUbKoiO9j7ZJMQwBs3NYHd7F6ypdevZ/W2a6NPtkAq7QNR00Qt66vVhoAMkV9O
mx45VHi91mgCb4UuOZVXK2GxhfzKbS5BaU2YfC+CBdyuiiqJ8DNfWdy6R2dbA2D4ys5G9ndlYcuu
J9Jm947r3eP7PU5tWqYiahXULoaWbBMTVgl5IPt3iOGL7yPICpqH+wMCs52+vE5O3x1PiJiz8ju8
yHOVTN7cLGcJUPpJwoAzvUry/WxYd8kMoQtuHHykh97zpEn+btxIHQduOGWuxVpj+YPgh0AFP8Ly
UXp1bkBM2H738pvUH83yhRv8M5v9hljiNI7X43ZH63GaqerlKpsGQuohttjvtPpLL0V1vty0Cr0p
imk9DdEyKNWCZPFsmbyrMJrPstp45bbnfdzALJZile9wZ5PWCsvCCAEHPN5bRBeG15OeywBsomfA
jaDp2fJn4tDrxwuqwEWQ7wMcLMqmoA0uaoqaRNoZqd2zcBySpz0paGFEo/CJzrLXGsEKTWm6v9V2
M0+tZQBqDyXTtrJ4lvqNqp4kZFNeJvsURQy4dfz9G7YyA2fIkSfI0OsaUTNWCSOOJ4gde/+YRehL
x4xJPBrH10YK60Xea/gmgq0X9Dxvoat1nv7gw9yN7wT/Gf/VkjC2A8A4wju0Sxnl4SbSUU57QqoP
78Q/WEX5/76Cwdg9taECoXh36686dcJinJDza6OOcFE06wJaaYW8uaO+ubyPQ24IpsWKQGgrUQvx
JFzWj6hiwmF6qRCn+Bd+eDvJyIGxauiz4XRxngeL6J87ehj2LnZ6YKV7gwGsjHTcllPLINHSfWK4
43kiUNYdi0+J498xAcZxuBpBC5Bmvf8rFgFTshCk5c7sQsA5fRdTdxX/0ua6mvQa4Fla+CpbdEJC
vCzYcUow+V4brI4htoaKYGwSj01qUiEnjkCn4AK5Q7Abk8bvRxFmYUXQpJxMRn+H4kIKT6dO+T4y
ozckQVB6OSG/wXzknGfE6bTF9Bp1gSYA025N/atMdTQV0G0a8m8wrkH4kmjbGgbXOxu++3tOtI0c
NA5VG144/NTtlk+wayGTSAIs45dKK7aaF7dIQyoaYxbaxKCLoIxWqYToAvGM451H0Yy2PYeyQJiR
hj0jKO5VLo+GQR8VYJEOAaED7pv59Ta+r0p2HcAcUxmuNXx+5ZW3yDK35Rcg6hXm2Ls5gKuEH3jV
jHnhToRnfetF1+qipKk8ICkTg8RqxCm0TkleWLCaIWV6Cb7kcr3jm0c6TdI0L+UByRCYui+KO04Q
3Fsv9+kuS5SJuBLxyQef/Ij0KgNSQQXPDZs0HQY6rVujnPZlTmgMNpoIhoEzFj8Jatq4QtXId1n4
sBAkpoSMV75C3rjdbMTQOobwx28bdE31CgmXENvdjdvx2rxICCAL8DO/6xVvOrBCNgkg4aFpjbQw
K3HYyU6BJlMpNuY8eqzDe5f1kphOEEkSdrzfcyqyp1I4ob4KF3ofAqprUHhDlzgbY69n08QVr71G
FKRL4gGq8f0uS+qZjYkAUtWJ7mT3W72e3c1Fw7gmWeduuDP45EUTJ55AY0t1Xyiux4t3FkLnhRcR
xfhWecYzJ+c/Gszwli0Fy3RYLtS80bv/dRVryn/9WknQvJB9g0ZOMtE+gJzxTUhBDg0mbhDyQO/Y
U25kuxlfHfgaJlKv064tcUVo/BK71z0tYrEiNBuAUNJsTTiPqZfyFN3uetGSbC3d65XTqgc6xD3Q
V2OMP438sxKzGPfRHM0xb1ZJru5mI44TAw/981L8fOvqm0lX2p4qf9S+i0KB7aUHVfuWMCvOWAoH
BUcJceke+pjV1envjjoodc8HsdrzXTxC7ibjte8vaGRMwKcROVhsUH7ZgwswXl0zissK2zDw8Tb2
bx8SF7rwDfVEhNKfIJeGeO8vXHb0h/zjtua3pEiyYG5SDws8sceyED7em3gPL0nrLmHiW9OoXeOA
TcS93wmNmoqaqIzDukLhlxA/L5Ni1QsantwYJKI1jp2QTSxzSOEjHQ/UfKiI6EEEWiuURCw/qmJM
HkYWqPGh7GEEHujwi6Cdu99ZdQj1B+CKW0cuhvFyonKGkRSWzvvG/7aT16tNa08ZwTPFpTYJNXgC
A/VYjNGavc/avBnzhPVdbGxBCDtSECm6+t1wSZBEgM7tl20+UFnWUGdb78mW5af2ZduVBPx8SzSi
I08EBBUKa2XgWmtRfMgfvvkevpIHXrkLMChPSnkaP0wJKz7F4/WC+VsJqX8iQ8QjX4yFBX593DHQ
S2RjRZ4YfATsZoo0SHXf3pHn14CcMgyp4cJzpz0AyJ2fK/NgSIGcSrfijFlRY4iyaQa++iQfi0u/
gS4ijQ4geRysVUFs03gCB0P80VcNU78+4D2BE0/3IV1OL0c29A2gOFo2ZLuq6fFHTomzkP0Av5yg
93q4jMbwikVwHooAdLktEiyJYewncUHoSFSFs3L45uoTYV6Ve8Pf8szJDp8Zgp+SUHHHdo3N23er
Pho/U3WMH1MDkfs6CzJfPu83YCBTc8DUeiMkUQ6gwIvfMK6qGkW5CpBsn9x6LOzoYUuPZr0PL1MD
5+EP/ZQoiU+S99ySwG/a8pKAqoHYDz7LN642xGInB79pRY9P03mh8SOrQY3eM09vJXC7ECwkLffr
DiEq32WcFmkSBazGC9cExdw3KcXxmycvrGkvRucmEFVuCeHqVA36ab5HUV7pEs6PxEhzQmKSpc9A
Pz2sbvTUUgYhxSL763JpBHZJrsLCliHVyYZocuMSZZoXDMn8LAaFETQox8mmVaY+5/SQsjkwkTq8
11C8/ifcdIIhLGb213L60C3UxTKISs0qjM9GuODQFmeO9gd/HLgJUSMNtLSjerLlWDKADNZ7aqj2
nO3uh6me7TMoMLz/+sDKBSLMM7zMwEBWAa7AvaphOHTSuZ7vhU+D2VbGYlvE/I7VBnw9PpL2/clv
4rrTkQ3oQxSL/v0xwUL6AQeUuI2wa1OsuxT78VzeI+M8cHAjAQSS+P+doIbmNV/bMGVJ4fczS68Z
eAkO4Yb+x/zcAkhytx+tderv9vrGa5DCvffIc5tL6TWBwoNKqKaYAZek4qjAJ8lUR7RdTm81k27T
EjfhG46Z+W6AGIqZeGaaOQZiuyirPnWMoXancmKxLSIztsUXntnepjml98IlU0Pg90yD6Mtq8cQ7
gVnwxeLGjNv0wUmKBlCqeO3n5bpnNnqEIfbuVt9jKOAeahJeszGoSUXe2DBJhxFPH6ryXBXgIxyo
XFgieH8bAAoJ+sNXavOkSv58q8l8TRfAddhHFrtImJNkLFGR2jKg1zwG/jJ+G+TQp/YZ5Ux2UYYY
3guva+q2vo9k2huIU5uHZScDEuZLFI4YDYI1DVepUxjOmugH0Nod/zjntL4F7asArTaembXSGY6l
lB+NsF12xbhkXcZ3r72AfMabfgnMBxqBAwAm/hm2CD+JZkmcMLG2KtVtp6eDlgwWG277SGSIvx9E
x+Otec930NvHqxJbx+qnriK2gr5Wgs10xXE2CppSL+VhQDswUA6GBpN2Na/z3eJaf34dEHkWr4LJ
qcfnL/iXiR9+Qh649pXAXchDcgwWOleIigbv/halr7826dkhy2W0nyeRUrh9a/kN7IBLI4jPhb2k
r7JvViMImvPY8gZzKYTjdaw80fTs/2btEDNKNI9gJpWntL/j2td7Rqn2hgONXs/GO2M9z7XcXic3
Bt+bZ5Pwkz0W4eBBqKp67QrcJRLg9uY1n/FeVa8XGs4ljD/wA7dQg/EGxkc6+eJqU1ZAI5ZaL3hE
XdVkchn6LHsju3c7RA89mRuYzO7ybope1IfCAc1InlSjkYzePt55e0/Tf5mmDRRqKdjasjyYl3xa
Glx9jYy/kndy4PxyewP2tej97wb2ZgtGu3j6sTZ0pcO+/ifYSJwjkRRUzNi/4P5yVJfA1QKz11Ye
Wa/xxmduAVv1s+q9kudbtINM40M86HC2/44N9nEvaN9gR/HUpeJrTQ+yAXTokZyBdxqT8tfdC8pT
J1AqcqPLsJOiBvP3vO+elBsl5Dnq0zqD/3+CKnoTNtKoMFX9p+X3+0wcurjaHL/GTc0x9Zqi/3HJ
56r4ewfST+TUPeJiMONo3pBJ4NE6iFcXcrqpbB4vJ+P/FwrBVcL60OTk5NuWshGIJZ+CBPh90sVE
i+dGXuku3k3zGNgwdVUWvclo4Sk4fYM3E5JaOLIUvFhJQJ2MzMwCmbMC7SbSkA7y60SyawE+gltN
z3iClIjXambIapfcv7Ax6dv74M6dFUywWy969vJBk6nXN/ubKAJKab08V4+r16ZO3swTH+CXGxeD
HnRiAfDWspI6ezr6QmCljGAoKETA9HZoDbmilWZ/QSf5xuOLoRKbkbt21HKVhoMmjJ4XAmsmu5re
csgYwNaBKf+cXXgs/0JDI7MGSEGEfEixrCdTlKLrakRBGXKVAx6s3E+c+IiuypToOuVoPik/mZCa
+ExLX+qQQFGxPYVaRc9mVihUXHL6F3ji6mdSjUmTOIz6pLkW/3pX9HEOgqChvnFmPDM/kwclZM/4
dh+iD1jetkMGIcPY28sN7Yp7Fm1JbREC2vVvGJ6vlM7WLjJtvP1tvHKocUVwB/Ea/lHyqKABq1fs
wYg3udir4VtTGbLmyFPZMGQfVqB/3YYWnR70f/IjSoxH9xi4W/+jUiMqpdZOFUb/8pBo9iQ+6LK7
1bTuR8EQrdHQTFSn02quAFcT72NWM/EQINK1/c0vNTvmn060bPB3V3Qzm0RC7Ify6Na6mGjxAdyb
z11Rzmxf6q39irZ/9rlmydsQhi4cZq+8aoiHde8Qr+nKH69HoQf6DHbvBX39FCTn9EfeF0lpfTSU
d/UWl5NAGyoV+bEwrqBiodFjki/PZymPnn+wn1+S08BmtsqsA2jWlXkPP7cnguJ6X4wYCrEpnQfq
mbGxvjpSzMxrcq/WViNMzG6DfOfDsnA/tsQ+y+1WamPDJqzTHisNtKLJtw/sYi0bRac/Tf8VguKt
bOkjYqqO2wy26fnezKpb0cxoZjAc5QNF47L96hgKR14hDv9RZlPz5H8fGMkDLTkjroYoUYCvVD4B
/ufVZOfKwOaBX7pmWXyhOaYukFYZnO/Wrco8vhd4tO3vY/7I/7DbBAHv4llF8ruMTqh2XLWuI+wt
9PypvraHG9JaMkiZm9cQE9UghowxYUzQ5vKZ/HTxwanAa84OEE1H5N02PQcslHbFwlMh+eWpfZmq
GLFx5APfRvvbXIUIIcq5I7JhO/Ow/Yj7hnsrJNBl1YZnq2gsHv6Ln6FtCjVeU9ZEzZ6N6+MIdtb/
/n71WW1JcHJpJvRFRq2HS5TNijr75d09GsFbWa4muAbp+90vG8G3xor0tZnfhYdGhMSAeeOacQFI
QOP77PRXZAgnQBAPFYuJtsezhx76Chr33F3XyQeLaBB/33sQ3+CLK/fBt+FZDq7ABm5CrKQEmWTq
X+/gypfzCY7irtCcxp162eQfPhujgJLzbIeMeSJd1oOlRunNye+gBUXxCLnz2nutWLp8YPNoPmD5
FJ/7fxeusFetrEeMfHEYF2EwNGIDryT4j1E/Kv0LTj1cs0byM9k9uvXeYDMX+KFXXpN+WJs9CRt5
jHNSK6Tk7UxOXCLaCdgnnQuTrAukL0OdzcaPOwtlFGJUKRR9qQHhbsCW6/OOcqVtFAZWbOGSwDll
ExhefzgrnE+K+dXCTm8fJI4NILmRjSL+ZXOZtVKCgBqSBgFg7QwalKvmiU4yymL94yvortfSs/vJ
KEdedosiW67xjwYOezjddh1pyoQ1Z+XLGPt5VaNsUZSd32gjg/8ZsIDldGR9ge4nzsgrdo8kBm7e
oPdIaZm6fQ7U/D9O+Dp2g+iqcpIp8/sIoDiilCd6+JmLz3yEZpdFa2Cp3bV3Zxn0mRvT3w8RMpKa
VHpxpGDdGPQEKuw/avYh9UKx9ZQY+G7H2RE7QGbdV5A+hIoewSzTjeM6nw68WJCNHE7fktF4xrLc
BUfRO3/RGaDDpEj72E5r14axNbfxpufjEPcttmROPxFyw/jjH58Cl1yXO2xlYvvNu6PB8EXYA5UM
0yKJJorbT5XO471+ajNakK1TFYjVmvuaXbh5X9XDIkEmIgA7GxBRaHUW/U6pbLEcPi9B9ELOyxp8
di+qhvpeBs0d8FaRkkRtlrAd0cS6+8FBRwWvybtVOMF1DdTjp0bwsvkKKXQReewB9SgQpP5SJrP0
dkvmJsiNlu4u3Uek6ewbIC5sKK/AzW4pAB2dr6K9NJ0e6R4gz+XUqJKg6fvgoVpXeV6lVZ8ztJUU
J+ccj+sRRj6QV0O79by1y1n5k7QmGYIkrlPAzeO9BZEEcHKSCzspDJBZvMM9N57Z5I4xS0y4BiHg
kIXAQT07P5zL3adQSjdS5qV/O2Dx9Q1s+IOLACJAaJB7dLIX8a7VtyKRU5aKzxpVw6OJNC06zAJC
OQJM3IeankjsdBC3A1NVV1LfIgSVTJ8wHiKjRxg5AZNWJKYvjmtyRSM/OdtgHgg6ML3w0zmQ7Bmv
M2KA2gAdvmIYNHgunhlwVB7Zq96pesJLDLG2eCeNhNWiKW5397R4EGkGH33gW6Iww7hCiFwHdOSf
cKMGVyV55U9LuMOYc5cwL3SHJc9CprlN5QEJHwpmCGLZPVEoOZqcwh4zBtiDajlcRXGQCN0GClW9
YVPVPagrMg+EvVNWZ0luHyblM1AkFFJT5jCLmYA2ShGL14Xqc+NxJFYK1oJC7RSXXRJVAvXHW76C
CGE7m4BrEd70eq1NMgEntiZenki7mDdY2xRZTQ2l1FYyjOLmWCl+L5qkHcmBK/2B/NHmb6nwvlAm
ybgzoROuTlWwaKmhCK+JzJtdLvJGE/jxDcM5VwR9WEVIA7Deoka9bQkQpHZE9knhjFdCULgVG8bp
wcjbX6a3q+ONH170+LqohByXrc6Ti9YJsB9HZO28glS28O753xoabrKJ/+H1Xvz9iISwkMdwUR6j
LnfruW22RRYPYlY/WCOmTc65ca7Jevc4NqIb1xIe7IUr6xAAjEwR557zvDjwvyqpkWyfemQowbKF
duGQg95jlb+4ZjZq4J93WMPhbnvnfnDeXI8NPFzOPnqK5MOinftkovbpz6YFGnj9mmDe86pB+tdP
XOnzsKqsuQdSVIpTvsdIy1PfDTCGrSLyr33H9C0Oz3YshPYL0M2jFV43xHYZ1wgILWKO4OoCl2eg
NLTHmS85xWl1H4MqyhqIaRdUoGsqgQkNYDIMAgueForQhoRrHfj1BNVvMH8vSfscMnmodl5wuI0S
R7fzh/oXTLIvOhbLBZ9jFfOATyVu0RmUe1NMn8ibPXnXnsRxNi2X48XAhR3+dbTTAi3yhiPL2IMx
c12UkTrhuQ29RqESLV8PpkRei7VCh7WJ4F3BrFuJhpVHqWxZw4WW9mYe3Fn6wOizkD3AM+2h1OKp
hrdvOo7uP4YbDdFpR+nmr7tpVWkONMraDubjrDC+Rm4VsyBOUmVhj5YmrtDkzY07/P86lwI0vlDf
aQBYA8etYyJEAQlmLcBFL73DmrJRpJz48fCRT4tfrsBV4xUpjAR7n00PQs1bfO+l59wByQ5s4Z/b
4B5L1K4xm6ZjEdNb32saTIazTLgZNKq+mxg13oUMHhzZ6NkCD+w/SoB50Ca7FSJj15B4l/KFtPJs
jyGw9yfqegAGg6ReJJQznyrjONidOQdsU07IvXI1lZLoxqTtJEQASBIkRVdHYcjM9Kp0d7ux6N9t
N+LNDni45seYe6Vm7uEwQkYc8rPovf8WBvknX8gURNGs7KsVifG7/tpSEfodIfEYa8prRYoaI57m
T+hCwWk8QHIztPv89NK2aGrYIy2Y3Eo5VGGK2m8eu5Jdjc+lF0XJRIpXbgW3Ryzi/3Bd2c6zfJBU
HMIQa9vbTgVBfI7BYmOongVb0R3a05Z9zAt+/QMhlA0SqawrvXxOJQ38rNOkj8nOZ+hCBjDsNZ8L
hIlx/bU8eIgB4ftSLg8j0SCRrfM/8n57RLEqaj/To9r8+f36PsEGDRIs74EZs4TjR2dwm5kG70OP
TTMocK3mUam0Adj67EsLQzplRADhDZ6KVfFaYOCuFvZLU4GP0OH43O+GID20fGZGbnZLA6nUG+cj
flrAGmJH0wUm/cDZeG18O5GKJlh3PEBGnHd79EY6QO8wXubezwweQLG5gSzLAj15Q1kLGsTqf0TX
nSQzjLYuN9mTxV8BK4e4mLvHph5C6WgacV16OMcJmy8xDYWxWmK9rSNJ8emCN0ySLVCjmHtioQxU
M71o4bmlCH0u+IoqozZrN7Qiuyk/dAHiaBrAdOqi55piFPynWGkaoDv9hZhlJQPNY0jzIvLvBYw4
8I41d3zkZjDdD5QxoHg+v6i2/wipa2lkLEOjExzuHRUg9SlcZMp/zUG0Z0XCWSO42i1isq/FEZlm
2t2k43uUwKgxSeX3nhWZ4kNy3vFG/o/wN/k3ipPUz4fI4onQsSrvxaTW559S6AZNA17YM2vrWJPy
Qa1tfVMvvoHqM8b9nsDLJaq+34chod69kUxTIpCmWGhQZqjPJcr/cqMaqdy+BJZU9dyNkdFMZsk0
gw57aCTL3aPUl4AMtzInbhAUn+hoBpXJg+llrB75IRK7Dz5zw0BX/1D2gzsJbufCTa3cMkrxSiHP
fLv06UPx1CQXI8UYA5kbR6lX0l7vUUH1G4T33JIhHtva5YTUhQ1Bzj+Xvl+5+GgfjLjmeq5MHrvP
feQCBVJyLE/XTdE25hM3H+AUCNVvhCOKj9URKhKsCjubfZHLxeDWq5Ydj5r7x8fnoz/BRzThXYD2
qoh7ZUh2lYJNpgUDP5cG2jFX/cb6SyceuCsNtOOO2b830PF0ghNZZdZqwklcx32Rs5RPWCUn7PL9
giiH4hj4NIwdwkQSH+AE7Ebj1OWILnLcJqCEcG80BVOqzPlRn3jvIoG3YX1MOC5E/fk+iR6KxFq/
UccBxYXS1ncr+2HBAf8m1Tv8qfzLX/pTw4G90roB8n5LEtY6Qg47/plHK56IXKjw7bllq5HXrqHB
ZNiSxCIqDbFguLrHPp82SAg09XD2otcDrDWUKr6JAmh4itAiEjbGLQRw63O2H7Iwl5UcIZvoiiYf
Ro931wLgf/8WxCxF94gLucoFzA2DqPj6+0p+RwtfnG2BvjqPyNGWCbvBLdxXAagJqD+JkvLKyiai
Ge0Q8/lQ3m0ZMBycNxie1wON6D1XojRTLa2tZ5yvFWqYaiOXWy4q3rrvcgm28fR9U5g2KIBrOUW0
G5YkOXL8vqzE9oZ7jkWZ2K641AlEpwKY4cT5chzj4rUVrKgFds33JzaavnzAnPj/upbyko8NLAUa
MWCS41sem9D6ddMU2UlkIa6yaPOcwlvrKBozzrJTyZOWj4esLQFIB0XbXQKTWOGzxmx2Af0+G1QV
+uPlrViBK49m2eb75IVcj4GuAqwUp2bkg6OSsp7xkjwzGvnjrUys4Bqubs6cJdr6QxTW1mxtsabu
rW933hpuqzKmML4P7LeldtA5oDCX6OF7rXHI4P0/eis9/YGaac42hpXG4CFXjxx4hjyGqXIG2NZj
JWbi2ES2daqvwRUQiOL/JdYRWuOtnlTjbLD27V9ps5ja315IScyy4c9kgPEbI8OCUdMLSm0PlUoe
CnkajU7oBlHEf1lI3xrZinbcXytkuI/UF/t2qpocdzm2UdwQbY2ad/ketRIK7hKyz7HwQbKnjI4I
9V3uPsx4dziY7ahL4vBJLoftKRikAiZG96XJ0Y/IgDxYVM+yas2ck/5aWeeNY/lxExaerKiymh72
s9wx1SX2q1D58mirpyH9Yk4V3K5yeHJC2yUeQ2eM97sLsU0rFqMHbOTJCqnlVFZVH+Uo1ym5lHbM
mUsR3zImybLrbjSLYJiJndnOtcJJEy7yp2X/myb5uSs/Q4V67/ySEXiPskkiM6ndVT9bzERmI6lk
PfmuZ91nRNCncaIgXwXVWHBohZere+R7jzlM0ZrE0KqSBgtpxVh4nCjhVQhBTYAruhg2tpVZ0jNe
JDiZSFGNYO5FKqZfgcK9QCT/dFbDjOBfqLzRd1ho9RCxnoJv4I3QjX+CZepEE2Sdcl7rLIkOq8yU
aUkvpOxxh+hWsUIWK7bGb8ejuqSRyv1kOlabN2aodPVOb6I8MStpdzSYBL5B/pp3gh/gKAdGpYkL
3CWb4UI6v/OZi4KrRRFPbFXwcY4BZFVHrv7WZU4VtuVx0StAxeIXHlpLLXuceriXsjXSUXAULFBr
Ek3nrURjkctwe0tkOOmyB56tXEOs13im8DU1raIQOcDUGRnSFLvQiaSak3g8IV7NugJmwbfzJRyI
3fuElM24mGoOFl+doJ8pRIJo031sgKYvrfZfahyO3IyHi5IEUPPBt1eMTQPVTkqEaWDWO0zWoodX
xqTDRF8wngsnZOc4pEiuSayKhUf10SFNyi68YZSOkQQab8qrGcRpu3UooEr6lyyA731FK3zNBV0L
hJXapS6jAg3pu/kT+LB6/g0KzMuRpuSgDNwKWU00LcZTAFIGYvlkrPs2eee+N4zuH3gedIaY5Swb
rv4PzcwDqkfee+NtGpjNtI56/ETa5MIpL//qhtg6MKxobzW5unvy6gRNhuiViDjvQCVXEtUuF4MF
jKBYSMnMiTu6KdHrwMb43aQYospMgeuz6/75g61x0CtXdPdB71Qr+KaM7K8LS/LSf0gHQ8fP1oHN
p4KOua12B/fRGDD2it+tDnkUeY2CuR4pdAA9fZ8aE/52RerypP78CG2gaNXzl6dy3XTAWuDPgyoS
bDWc9dVFjBPH6hl59ZdUV2eBt/XOeYO8JrnJh59Z8DW1igXZskV8dTHrynpZhKaLlm3XLx75X05L
i/9uXfKBLre6ESpm/40BDVIL50qT92m/QvprPmMSKv2tZQOglhnkUyy9Ab+C3wF7bW0O2r8UG2fA
suCPFpO2bYs8RuOwwcZlpMLpCDKPOu0AP643+yAaKjYa/bhWbwZ/fASIW4gdEv7mNurPLvO0aXxS
L8bg7Z59Hw/yWKvqHUEXZcU496Lk356aUkIxb1WsNzZV+n5+jFGzHCSUDhKWHIEmquEpvgWTikCu
Ar56qvRpc9zSMKXgmx8aMdQ2fXXMtb+YgYD+r7j88p1IGL5p45EAfrm48ozbBPfJg254jBoanK4Z
gR3g0oU0LFUA7z+vobfQ+Yjgi0Ch0fTtsfEEJLzrBs9sg+IupOSo/6Fq9y2ELwNvh4aPc80tOhEY
m4pMDlVUoX72YGYknLNzm6YBR7QZE12CrQgQOLqqckVlz73XpOSlRU3WMheetO4fJtb7xh5vy2Wi
fsVVdhlwfwCTde867ppTN+ZjdPR2tzvsZCWNMS9x+0Fy7R+OJBeYaBLSWgIPjeK/hTg1w358dZlo
gtWQ0Nhzb6/P+vrXy9+hSfjLuIOsHmwE8kGo79AZ8FE9tYFidyxkrWWSynWwAwjzwe9LPc5gG3nW
KgrRz9twbjGMmkIzqASHRwzz/bz/mA+iMy3RmEi56c3ayBCbU2xa/Y+PA71wALJHS3c3LYIfPaN2
DhKUxGOnnPMTnqX4CEjY5i7aZRh6GkvUJ8MKRlNHm8hxu1TZWXqb81+zZCGZZ6HjFvmU1d0JKzhz
qWKgUvlcoJXuCYgOUruY9zs4vK2Eu+asVab3LSss4sAPgZk5RyUlCmUV/H4hy9CP0ETtIism9QnQ
zW6Gqc5jyhM/zEvYg0MSLR57khE7S/pqcVmMsxc2DTASJ0618Vp7jHC8l9yE1x2jg+AAqv5aqOiC
NI9U88zjergd7c8rpJMXgWqSLnDqgBMqR+YiG//7gnpRJrUQf3uckUbo1H4ocWrTYUc8GiEEdmby
kiYDfxW05K3GtTMwzFW+B1dqs4fXApxZ0xvsgQ9NwdBSve94IQsRjyqozLcCc/AmjsuF0axv0cw4
srqf5XBIv6BWabNUzt2QR338i219pVyoj5WlK/Xk+EkIAsRkVrsOj1joCCUAFMAgZ2PN2lFP7B3x
8zB09Xm4m3fxIWSiJmZIJkpHMWe5wjc8I4/+EYuRPscM8WT7jFJMWkdbnj6L02LeUiS1ktSNJ3DI
/ahWJUWCJwqweQQFVRU57aI/ZEbv1fA8Ge4duPXcqFEKXDhbs8BKE/jZm0F41oHx1IsaC1LBXtzA
/kcrWDAkY2gLfyRckgenffLh6N5nks+TVo6ETwBt8CUfgXOXvbNDsgv+kZWy4Kwd/U+m8wh3osYe
ITGs3S8+vLXmjmoxcxgRs8+/MMeoHmulO13LETO6wudSadvyjF51167LSdosoPSr/uWLJ865KMD6
T5CZnG2b2dVdD/yKCsaJxqw04A1+LbwTht7cB1nuqiHlyOPGjIXOBaBGuSamYDs7fVk69b/pl9HS
kheWjfUJg/rhgqhuZVfonoIO/Am4ZRUz+kR+kHb0LbkUTDze2cRl/DceZhij7rdTzhrAKZWRx1NW
Y2n5s0tQPjAIZviBcN54uIfy2BQLxrx5dt/oqJ81pMdl5iJxIFziFnyBuxkk3uPh0wkVbKPZVoMV
eG77DQ7CNnL9lp8jpvTA477fTbi+MJ0+WJpj7cDMqeSFbWRNQimhmhKCleYURie3ZiZw76d7aMeg
t784/iByPA7ATa5rdkhVpD42SKJaeWOxiZ/TnmLgP/WLuYiRD03Brgzd1Q58NgXs3ocKOdYsOKvy
U1ICCGhTlh7QZxWb1+f6Gyb4sTk8NnjXlQOGkhVaw8xOj1q2RFzsI1i4PXbb41nk3V+bQqAkzUEa
TKbs/f/Es72EId4ewRgGeWA3GknTb2paOYXJiPSvkAA/1a9Q4nr4K8To8om8ppmKAluc9Du6o+rz
tNkoVGDBMZf77z37gN4DRDdqSiTP+j8dOb99CFzYePX+RHB/u+rBzm4B/mnJr4gV3XdBNqhCuEY3
pRf3HtlodVSsIY9DAN+oEBXHUjcmJjU70ynVrzf8/L6EBUrmXMIdMd07npqn3E/PgloW85+UHxc+
2cF4nMjxaRu4MWbdEEfLwUHnsoVhObDPSq4dJb4FIidvR/e/5Y/z8+VYVjua5/mhaeiJFhC8m7A8
yWZCRSfGScnLUb63LDMxJCUB6U/JOHGUEEfAvudmlHVi4f7yjHjV/6f+AsS9HcD6lka9oVtxfU/l
WsxnZ1zkCiFkmyRAWqbmyi12ZySGAsNylm2otrp/9LeB0OTzhF5dk0BhqAaBPRR+B06kMJ62NBT9
QqTnWNJq6PhC2qUkYKakbnn3tJwBy761XcohP3P0rPu11wTCyElEWQu4jHrePOWqF3eCtAUQBtUv
Q5f53a+6Nj6PE6eiByj1j1LjWRzz7Pu6QRyZ1gknKlYRoRP+jKb93jBWXU+coPFy2jD/ijUDckfl
GOg0WqPMXPafKB1ABK05U378U4gCcivwkbWyrBkcEMT0nNZs60UV+gB3yLSsTpX0VDJIK4oUxLFt
gJblbj1kOuubgo2k3H+upVxmu6UU43kmZSE5LSUaXZzLSZ618yAdB3aug4iwjmlIPynv/dTZ/g3T
YLZzJrIN0UuPKY4Gs/ihP3FNhF4irqkxA1mEZJImFOrndb3CBStAMCXnA6wI2iJKmzr46qUigUQN
beaD1l5HS44ekm0mXb223iPIbikyrkLbauguDn11KKXsKmoSD1mU2Le0hyuEgBDGYupqQUMFohT4
7vLNFRlNgwoNvu1rKZb11Rog6SzkzPj03oA10ZREZDy9MDgAMIbfZ4H0BIUcNLQg6/hmA19cQO5Z
ZOM58G4lBUhqudg/7RjUJmwDx0Hj+wG3sWL9mo9itQNTz5tdGcXc++vDs4p/oiJttiMsF//R1P1u
k2KJLR/CXnwsMlBHmLH9AnboRA5K8DpIVboVNey8pFAZC3RaR/DqfMbTuIerogF/ANKPP3syoidt
/fWxjCGFqLhZD6xpTPAVJqcTcufDKmD6JF62Jo0HkF2R9XBNrVTjhE671FgA1Mwj3BCT3/ai+ZXx
SI8schFy8iRULutcmt6gW3FCbCI5X5lrvI34EnnYMcM3mv2BYMmFM/5JA3dULXvG/AWevAwZUw96
0Lu5iVffNkcoQeD+T680Lv5S3uwisQLnpVB49rzizoK7FUd87I7WhbIpz/VuMPkvFdsPyPgbJxjQ
uPTWtra/ga8HgAFkmT4iTJ8W2xM7CtE3cYYPI8HvTrQCiut9V1myRkf+bc1QQ1UWayGMJODSZ59p
RP50Qi8xRXMkwXKLvREbRHtEkIW12jK3fHFifauZSL6lTHA5wrCvPKP9KH0MHoRjuwRq9EqwIEfC
uFna3UzYjeY27Oi2QINCx+It7MN91ktV2wUJlSoQwBOlXxrcRGaFNc+lbFhX/SEK+ug3eOPSchGY
dH3O2O6QsiwPjh3bpWmLQPKD+rRNCiHHvwUKTNc6Yl2HPJqMttzPu5pdRwN3iPvanmPZpZBv9j+S
e8P26eDaKPHNOf1t9BIRpKPmd2jgG7oGrayD8amAH5qUL2q4wj15Gz09u2VIx8rz5tlpKMJdapqd
85UD28QspXkJhnLYlJiPiXqgiDDem8DYCNc5y7Q9Q+A/rXAkBu3u6edfmH/T4txjEFeQ4RMgwYcj
HDHI8WgnYlM+W+J2AkxgkH+fYQhqs1POXDjlFa9bK1PMeudOjL/qAIcEGyoR5dq8wI2pelw+9VYD
f0Kd6YZjNvnbLJMk5s2VCM6i5S08yp8qDTeCXdvxbYMxVVKX3x9VOwTMU7pLfgDbW2xddTf8PW9Z
DetB7RltOqJ7bYIRaf6qXhcg/bd4X3nXsForAvTeHBJ5RR/YfTMSjIE0LSKgR3PnUH6HCj+mpAhv
8BsNZBv5xtDHEambBLWrX7Q6cqi/G8Ews7p6sj4JVN2qA56bTJ/QNdt1aEcqbchLIifiMWeYqGET
ttiBA0Ep5ixtN5tSkpxAp+A7tDS9/pDCqMOZUoXNcljgGTZ5ShapBPdTk5k9aukLMV8QcbIJiYOW
ywpoB5H/Eu7lvULuctoQw0q/1/31MOGmW0Jr09iqVhWVPuuJyasMffy1BKyzp4WNFkhodeRoGHPj
WiMxdo2IDUPqgEpVk7iIaXqc54rppwyySq5u7IpsxhiTd8KG9MYXHMg3LsD3xwvdOEY9XfcPQJZa
S65kt82c3TCn72ujJNibtSYo0uSC29R2ddQol3ErOPgiBaGT8KW4xd/j3PhACpPQO2PtS9WWgPsE
WiIJmox8aXW4/btvAJhL/AmsGXJhAk5a0ijNe/v1ceM+i5P/nVkIFfWafI3Cwi0+h2yKp0AAXI/n
/ICklTjo5jsOY9euIwThi5qVLEOI2+9BrkQRCKVt3xd+mrtrspx8Tw50vFIsT1k8/NwHKC0btudl
7fJ1tFxzvkda859jO0RiB1ienQfr259+zb7YSBKyxYk0U5CYe4Pf5JT9K1u7AjYjJCCpMCevr8d7
c3vWKL3kKDrn7OrCXLdb5Dv5/MRhLnUco5inoxQnCeiTiqgwYxfZ+h1NdqjIU5f9zzbyoUyqE6s/
ndjsN1CTiK6XRLq3gprH4z/WyjnzWpkn6lZ466OQMNFf2XmZAV7QbGyjbhr52fPHlwsCmjdhyWfF
SSJkGgY1i0aVOHl4P/WygeJ3J6Gvusrhfl6JqNichnKmNI0QA/7ILqpXzTa/yuRLnkKdf69J7x81
w6xUIty8zpAFpkXdpQcRt4OaNO/ykzaGBmmobpXvucpGZc1JX3p2l7BvZr7vB1k8cgKKYcBmSBND
nlMDa5lMGF/+aOpfQiSfban8nYp/0BEdEB0+3OI9U47lMjE9g3LVdT+AWayoS9biI1I/1i/jzo9l
tAtYjypRTGMAkKB32HuN/SG6eetIyQp4xsIBW18IuCONz/A8S0BKi2IynWSzViZBATr2LUbWBjZZ
t4jvQ+ak01u/Cgys8VQzD99M6u+qi8xEuYJcBPkPwyzj2A7YsJpG23zawdahxCzZyKyR/DUrulMX
TPU6/ckmH7uwLjqs6Wy5fHzRRP9Xz2NiOOOgK81M+vpKyolCKmccFZFDo86ug8DJqyJyvrUPGM2R
pOz7gcgP087Y/eQfk6lQor9+g1xXtAzy1uaoKhLuT1NdRpLLSvw8197xmaqa+ANKckcVxToCd38v
w0rpvGdK10czKXHKkBY9gY5FaI7LKFajeD/c7AXyzBA2rSK08X2yNRYY2ehn/aNfObX7EI2K4/Yq
lqCJpdYFr4vwyBuUIYzSRMneIzG48ELqdaNPjBiqH/4TR6oDFSWH78luzM6x89Q3LPGk7i33KVRN
PM4YV58nLMuyyCms8x/1ShM0He3rkJu/w7p9YqVbUwLzInZkXp3ct24iTRqp6Gls97gQx5vxUl9P
0vbLvKgEuFmEi2KeaxWPzRRCUrO0vHTq4/b7EQUlD4bT3PWJFK5AnxI0/ffOIRfxTwWvfA0gC8Cc
bzqaURN2zX+BD5UNFNtBHwA6i5xy0vcU+igcX1L2H0g0touyOE/al81O5vMosRVvQMmKCTO6noWX
6IsIdUIIsyDWTND8MNMJCcuNz1ZqfBZp02FR9vPsD2Z1BXOBSoXCN+4TDeavU2Cw6fJ1Aapl1Z6/
SX/ojXCUDI3tOcMbU/4XJKimVlz5Q/ThvvOxnWTYaMl3A2fRlsjF1YngQj1i/jGg4PrK3K8PoYmJ
0VuzJ90R68seQMs3RkaCT7aXHJT27nsG1F4CDU2jooCHrec8COXfwb1mZp+1UsUHxUgYwrMLguab
qvW6uDtZhSThcL3zxLRsb66azPgoURbOULth4VK+W1NhyhAyvuqMsAiH7uwQEVGgOXSSqHE6BqXj
P4ZIxV4LVhS2HV+70l/ePvb2AxV16YCbFFkTiAqG15RraFcmsMCA/AiyhOa5DT8kI46UijyyQGP6
qOczU6KppPhjBh4k3SRLJDfT/kWZJ628c2XaU0pO7pkDUew0z7PJakSYbogASr2kl/hfaAuq9Mpr
Dvu9A+5DZVzZvZRXoKG5WssFKCLa9DVTqLJg1ZgRtsMJzfOqMxkaFe+d8TOo/t4txvM5FDd65GKy
8ZCRpDHtb7roBWsCzc5J5reujJ83jY7ZKyU0mMtweufHrluhP6BJ1CG+3wV/BLs0tWe47QSTISqK
zGdxpb1D/1x2u1lb9QQJ4mFE1rpPoAL48p6ZzdZ0o749jJFv0sPqmhHla2tF6twJDHs9GfWHyNse
sJqnh7zBHuL1Mn1C4BI8QXySPoVYMoYlU2eBWs8vTqhUZCnP77BMFzOtXDZP6VCCtrOvgykb0Z6i
5TlWLiGcG3t0mM6UqG7fbHqJLJ77nH3CkqKV2cnv09ERTh0U0wOnl4O8kV21z1nlgpVyNXTCg0cN
Sjb5y8t3C4ASszOaPaB9cbkqkYoduwcHwTJGjV6y9OqDOj+KZvBu+THzAOG0VCFiR55V8ncJE/Iv
CeKDFEthi7hbDa3iSRW3fdhBcCL0HCfT6HdBME4aqmEmLNoByMJM0Zy3ybasrHGbdt8dFsNGVgs4
4mqhwbcNbIa/DNUqGgDb/GBexCQbdXh41nli3/00gsyWR7xDLtPC/FllsByJ1wlJlenah+UFSKHy
WNEqoT3ONmSRyIA/YEggyY4nMHUCQauTMn58u/HJGEXTXV0BrYHM5RYgYoYSeVdg4lDWKOmFC8Mj
503sAUQLC8t8x27f2oNLqPWRSVn3PYZNodc1VAc+VWjxyZr+76QZEZtKzIGDGP/GtE3BhrHBQ3HQ
AogMYSJ35O+BmOWW76tI6M/t1hgoOzn+YaSdCoNJUfdCQza0DWqdr4Y1XfiLYcL98d6jhHNSpstK
DQ4UOLNZDgjOX2fA2MZCyftSme6QaC+qZSIU0tZYXQY09NelUMeD/BEKsnV8jDVa/BRQnzhf1sb7
vDqbAtPGaGxWGHbnnyYn700se6yuMG50JU21cnLqhk3VanA6AKoQukT7kz1cdOwiywpsOaMYGfvT
S7Uzdp8eBBIBCU/Njg21tELyniKVHPzMHKEMoSE4zceMT65pFEM1GyGL3Xy2n3lqmM0G8djcQjTk
+lW0naaB8UWzioq1z9TRiEMzBGpvg/kJRl5JqO10WAl+hyIL2GO5ON9DtGamQ5YjDYi8w1uY8zpn
HI+WbpDxgHIiCtpfXqp9MmXBqq7YM8JO69HAt0mReledgO41dzYcn1rzyZ0JczvQ67732iRoMKhH
MJ5Jr7lb2V0yJQDgeNbmHYVKpP0RyVVO+UrvDqadvGBO67jfodgch2a5Aai23N2zJn6OdGkU+0cE
Lrvv4S4wnr6waYAzOtJGRk0gwop/MjnuQATsOTMofQeIjDQFdw44vjZ6YC66edgJWO8myxQQ4sGi
56np1hxOVzgrovrYic3YGDet0pGr7gL8zobvZhBVnI1FylP9zsgo2gu1Idpxu3R9f2vwXmpKguVA
M4CYM71LiYJXChTVtEAP/H+CLDM5cXMEjGJPH4twN9KvLxGFatJUDwBItlT5tvkZ5K7jU8CqAvr/
TdC4qGIW9Blryke/ENjSmRlQ7AaDACfTy475b6q+oKXsa2lj6HUnnWE/B7zS42Fxj6+8lilV/wbK
Pap8LJcwG7cImU5sA/4qCT0MFP2X395tdQWX048yZMEomyNvghQTxxN1hJ1wRjPV1UrEh4arL20u
M8MyvUY+r4aUmy7hBghvZQuxCiNWzEtiSgHctKW0xTOSsU9+HS6axzWiG8BNln7VQER/79bkDCp8
4etob2MOmHwKYGnKSeFRcHxPrvKhkanysAm9TCn5EDsTJlDvKIP5gVYTMPEBuA4bja3LlaTBL3WB
nY1rLAqHcsa/OeiR8SXT+ZqKFkRJF/xO/nK8UHJ978tR1Jav6DL9omzNDuxOqbijrEO2/EdFoCIk
ZLCtgKM8w74ihm+/T12nM1DKr0RSUcp/d7XviI5shflbYPEoQUhpzphEo2onQYsMq251G7SaYPEO
o50BnbjyEI6AqzGKUmqh+UT9WvFJfBw7fUJ7X1LRA6+zkQ9KoplmVPomQU/pDuuv7DdobekLffgF
acre6tsvKXW4Bt8lHe26iuK8+1WRCdd+3CcBFbbpT5jwzHJayLgh5vZP7POZgXP+OpY+QGOQk0IS
HVpk7+RXKXot0azdZUdEcCofJoYQjOyjyd3DSQkX3cunqJP35TxOqMU0Ss2W6BtILh/RnuEPxmez
RmJv73sInwtSbkKituLgp3iv1kdICtaMbpFFSLGotCRX+Og+d9qOOpcQ13FZWhpJcenndUdEtL5f
7vb2ukueQ/jHL6a6G7ISMtXGvTWE6apbydfxEzT6w5t/6gen2wkLSKvYPu7EYxHl9F7hn2DT8rKT
yzTin/q9Lk3b4w1Pwh6d2huKH40GCa1v9Vrds7sh8q9DzQSin3PDOZYPqQLhsM1fDHvquITTr1z3
kPc9cFF4Ap3vt14/I0h9VWgHh0F6TQ+Xbl7ERcl/4/skHr4q/QVqqyUq1WfssNLObXh8DFbT+WNz
+/ADbg8rEroyrkVh37HyBmCnPdedCcc1kau0nW1PO08E+lZ8XolNe1bz5N679WT/szglDJtz17Yu
ZEMpmCzac+4fmjNxm84qXaT+FnTLYWy+uJvNGPknxQ4b37Cx+mplB2+kouH1u97uypOsNIOgo6Bb
OR8DyGdUpqzHpcJK80TUk1SCe9dZTpLG/gSPUVRcU8ElQjYrER/BBfgcoSHGprRGN5l42AzEsUqT
DVxnb8REkHP+QRvMpsuz5rBolq9h2TzsAf4ZtqrVdmijiuuwUQOTNb7AFCj0ScyAU/ZxeyWIXhfC
/vTtlGZJ1EQC7Ssiszb0PGzVVVx+5CflQkteGBAWUwF2GraV8z9ShC2s61IXmEF8oMdbThFEcWF9
e9aJ87IIt8zSNRAHcdA8gpHmyDcL7oOJI4E/m02M+Zfhdlxc2Dn7/WkvgszVlTViLqg1yNip2Mh7
ZtJL7gjlCvcIgj6GPAeVBThcTQ3a0XrVUhK5NjP4MIBiE6Hae0Y7Yh2SQHnJAK7c6+1LYms80cU9
o4KjUaPE7IbxYQBWayfZJi12szM/H0MtvUDPlwncEaQWp1CWqQWzIW7uKktDK4GhK6MfCsRDxaOs
ci5GmxSWH9eiTO+en11v2uJKQiVnvswbyBWiNGYOGr8fKUMResdGMswcC4GJpNPVogpZpUnhN7SL
9oxQ45MZ+QqbKo9xnnabn+8qzFdDqA/qearYqsqFdAWHOId6qb5Y+OOyHD4r8VroFoGPpfCJ4N9I
WIHl+R3kNBgonaW9IgHDelzcodVGpnxGm5fNyjowReyY2u/epVXcOVskrJEs0dUWG3716rJgafvD
jKNgiX4uju4ugljPfKzYz12wmihLLQtwHq/ZJuDVpg0SbALguZT7BhrykZFJ1lLZAgI81nOUdCT8
JiyW59si6M9snfZ4emwiJAKaQF0yRQaUqmrCv+jP+bqNSr1hg5d7iLFW80IjmfUvgrrDTpMKX3Dm
0Dzc+2rqAgQUAwuFyGWobXvFlxIN8+5t5ata5s5kxKGqCm/n/cI48ZrO17arQCFskcokrYhbPrK5
amKrKBYEQ2LYc9tfHg7TKS3+vYlKpL/REoyqcCh1Acu2gly0c6tATD82+dV9icXSfu2Yf5qU7J+r
HpBaqYTnPVWNmFh7oh6D8RdX6n4kxCgj2VXHFy0mcnx9HY0zNdEc9j6eW41w8EcUQ+xOzYXY/WvH
HOJghPOFkaCcfPNjNsrvwNS/nuFggjFwWicN1defBEKssRteNILwWPAS4hzyfNFgVGCYwvLLeuQT
KOOQ3kaFIy4sR4Dzo3WvTsKfZFGFz6sAFn/QP/cdmgyd+CZvIqmAegeVQrtQvIzYy6HRjOFvU/Ec
dRT8XYfRgDa+ZDwKBY2/3O66BW0VCqPeliM1Ruan0mNDgUZ50eoiCNSubYPqr74MR+j+I/qqtbmt
1ofknU9dvo03Jhv8KhbpSn52Gv6n61NE5Gh+s1FiZ5kj9+VUGMLDjxex+bnDQoa4jxvKO72MfEwl
1ogCkCnoS4iVoU25M9Ac65SnknTvPpQ5eOAL9CnAihQwOgQNvpleQ9YAHT6PZORYwSl8UlnXQUI8
qlqLVvyXHTa83WN58140qEB5jdyh6VsWugv4gC+kON83cXB0C3BvxA46lq2oCBorCG/zp71iVZ9I
iws4mQVk/buhpEtSatpYSIQY0rUECC6j14D7w/eBcSylUpSZZC+ZPfAXnM6wfdIKqOlbmFK63cm4
mUYYLf56wMFXpmOe6kRoT1YMJcW0DUCHfOGo5q9s4D7VRk01jp7adFHnIJbPYT7OgSmYBZpC+zkS
Z0akstNm7AWCv3nKa5fjfk+vt+I80yvRYfzIbP/94phBPxHs5uHc2pYfRbliin5F0/lD7pX6b+h5
0zuHyavGMCy9QLb6rqawxsn0YZPIj40TIdKzokHKMCJsX0CSNSAEjBKmBZ/+R5vc13DoFjnlTabX
WM/LpbLajOX6cJw7Tnq906OA1TCf58QprJOVaKJZ3zET+5dJ8sWBlW9Q38si8fprKZiHU7JV/YrX
NyIyZdoEE3kzZwf9+uWqa4xWjpX8K/Lb6nL3fg4YvyZuIscvwGiprYvDxYl5HB/rI3/l6YoR2P36
4J52llRJvnT9V5q9AwKEDHw3Yh8sESWIwNjAV1lFxLZvyEZPtNth9pToNUhQnSs1foLqa2suRZhS
cc+DqOeITB6Qag+176cBoBIT1s18vm2qQesx8vuq+YLKYJ6wIp1gDhAYtSEMgXu3sa1rskdRa3NU
PST7SBQ3oJ+k/jPWAR01YJaP6I/LWArGn6Oe7hQRrVjOD34LpEeDQbhouEJunmqtcBPaWYI/3c3D
0+niGwIuJAHiIkQIgshyQR69KbrosLWZkcwOwyg20gyPzrdFTbjlN3I7OCY8bJI3k64+ocM0gLT7
j8VGriVxfxyvd1jHPRc0Ipeha44D/L7ezniaAVbhijI4Tom8VN8sjr3DZd9ZTjWlzEwpkohkL0Ny
8gk+/5dzYVspP9JAmCkglvwpqq+jjqgpAg7ewz/OETANwDpjCV9dxalCfD0ECHvcSrru4pvTWWmL
3QXCau0GI6QNynLy8W18asif2xgdZE8W40749f9YrYZsJq1Kj0s2HfJNiYRqR6uF5AdYw6Zhb43A
wpTGtQUDVx7oiwMpDhiJy8La4gZ+IA+1lw8R4jZaaLjS74q7eD/n5SXzjeiG7OhKij5YGxTD1JWS
DW9I08iOW6gLyKCHLcj9Uqf8/GpHPEAkFvabZzPiiZkfZ5xOc8OhH3Evr7BsIZLxj4RLcqep8fu9
xHmoNMqDdk9DAxcRZF5auVtgmBxB5K/Nr7oJWANa4sgnV1O+5FaUlUCu3N5AzY6sbv5pHoaXyRIi
kP4dDtAdDNNBy+86YcS9GT0HXxeHlyzBA3+ySoksMO8QbGvLrXwugUy4EqqgesTi5oc0iQ9lLKg0
JCajsZO5mPrAiU9qs/CFh6PqS9CMYt1CctPJCx2rX2C26vkhOSGLCNpZsCc9K4LvccSnKnsmwkX+
12Z/ZQUFHn3nS9pkhW9OGUGYOdQrU8mKx5KFJ1jIMA83rytFVR7uKiyZ7YVmHhVkYjMTcR2YsyEQ
nHqh6VEtmk6TXcdna/gOC9ZIirn10b5IuabzwPgnjGYja7A91PYEKA38uLTu6zhYfVZogf1XD+Xi
//9psXtKbktTr6GSoBLxYmJ483Uq/js7HbSvDe/sKe1v6Ecw25FbmJDy5rcDZQX5jLg3r5AuYBqU
OfWLFbQ63T8m0w08VdN90Ur+DiMkGNhtcrlh6GFR2B4UBPLxVsl+bZIcjTSVzGcOoepg11/AHkR3
y9acGAKLQpEftvwh3r39EMGZua5Vl1DAFTo1dbLdp3NKxVfrRbb/gGajvy5QoLl12XKknjxGwhNa
8OMZMrTBIKx/pv1OVSeJACbFiZp/SzXQ2ZQwmHiK5u5riojbGfVwaO25Ao2iFNA0u81fnDSMuwBx
9EgHS2BfBaiCRZNRQwhq9iiOKO5FP/mraPhN8Lx48V4V10Jlx/kHnonc8hxowMUKH0JgLQ61bGp6
yyBoIf8uUkg5EnenwjQYYxRm5DnGiVveXPz2vVZG77MyjntXzkhOYtRe5VZiIcgtX3llDoumhSPk
lc+a8rmA+wwK3nFo12D0KaSfUu4B4ojLUGFlbo58BG4UD5B1gTjFOZ3iwsZ3OxJfgKo/Kr8Puiof
Mjh1N4+xx3J2HRqwLuFOXwUXr5PR39lypAK3wrP/n1SozQ2sp1PLsA+CBnYp3BNxPNzBbpXCoSzP
+g1Cc1+XC+phP6vTt3HeF1sDxbD1aHkj1nwmZ1owQF2Btfcx2rVi/h7Bdf8Wh4rAwdUq7+GmObif
9eDnkuwIc2Hugd13JB0T6pBVHDlFtW4nMQYaYol7NFM5sUKuE6L8hP94uDTVXrSpubEALlu1huSl
1NIIZdZIaAoRb2R+4lKIHLSIL9eZztUErzAsV89idjN2d6G6S3aQIsf1M6F7ks4q7vr5GENSap9C
mOOIHWsa56ksVP8t0dyJAiV1Op0p+ehmLEo7eUcQpqvOPHrjWtjPUFLdvFUMwNMTZDKIuNoVrSel
dOx9f/jRNuC68CK4HmmKp0bq/EpB5DnmhTx8rE5KJKw6W0zWd9HyEO9Ky1JQFbjPyYLQcn5k0ry8
jj2DbeYSh0yronWPeKHGKnBRhdSG7xlw5o/BYszWq3r+aR+RlglLabvoIU8IYsBLaVzgXKUsgdw4
e5aQO3Fmcp6i66+YBI6enjNN5QtPDxbhVagDPPMb+RwlxzXrQPJedoxLWjVhJewgWxi0Q8h33dVm
G6aLlSAreVy9Kt5tDDaMEmLVskHugSXHikpkBuxiNuyFXHoBXnMyuUpYBL93pE2U6G0EOQwIJg4m
U99ZWxiU4Q/9hQ6rz5RmG1oP0r+m3rTgmPGB0N3yAQxUgcWjpJ2lkraaDiGntICWktXHK/5YsXwe
VQrcHMr//7JdjhyGGtqSHUYwGx44Q8HhQGcQQiJQTuC7mSKd8H+nm9l54rjrOTMb72GOGiYOxl8T
agHOECkfH6W3i9tJLmbomJWcob2d00vtMrtsThfi9gB036Mj9vNmcYsemq6qFoaFkIC5uC64hWqj
gvwOp9wHhUJA+wi6z7QQ9J8ih1KSQZRMhe3FUNkv930L6Ww2CC8KoPkYMiyLo7Aeg0DOdR0px3Xp
AcWYur63qaLXmmMdVduLb7nEyEWwDiUPa9grpTciL1UN7nQOEzN4RLajUbTfmKHLhwB2FDWDCeAs
P2hSAC89lVoazH1PfGVXOggGLjDT/fTzDtfAdM6bUJVpDRHf/ku6/3XT1+hVBgvq/O889hMorDc/
QbFURRmgp7nDCWpzcYVNGT093Z3+7lP7yb+eklOdcICHWJ7/7TWVMVo5rmOSiLL+nLW6oYdBG99p
hdUiMgXNCBXfAi7MHnsn076Gil1zzh3m1P9Wr7+qcn5SQZsTlTU/S5mwB5OH7XuNbm+s44zBaWrz
QahknQ9XgPdhuBa2CHb4a6+R1VIEL7cRIhNt2l0SgHNR/qvkhhrGXIjgywe8iqm4OC02XnwRnQCc
lNyG9N+/Q0PhU3IgnUlVg97wWnG9yHH/YqzXUkMLHmp2TZHmg0gRqhN+X+BHgwFVvYptL1iRT0RV
Cmcj+Gd5Ai2Ac40XV8hp4piwBKwBwmakPzeQksXXDEQetFZ6Y4QSa+/6US9sTYJqOQulmVVXs8vu
p3tRhnhicHI8e9APxGYfCHI0cr+6VQgy5f5Qp2GE/ulJMmoRgPXrGgg3xoZUxZzZpIjhVR3+u2Ff
jpUjwz2f1Lud4EeHipsc9EifUn8FDBk3omMmkqzPFaaCJ6FjgxmdFxFalbym9FXFtc4bL18wSlmo
6mRlymsVezgg6LuBjmf5ai5sLhKSTIXE7j1X7o/4NnlwpekeQmYe/+fkpljR6V6I38Mw3jIncX66
53zrfk3iAYYkbZqJ7IW73o+ExyU6UA385HnNHfWc+Fht7VnT0hY44y1qbx5cLTYPNrd8hR2rXFA6
sYFqG+aSZTdUQMYOCGM6uJ3l3gvQl4e2W2mC5LhuDVXT6HvlN5CsfsKVKP8a1+3qvIFQEjurqy5b
n36+dEjLQa+Wtczz0j/ox40o/Z8oV0oq2A627gqqGs1sXCN1tA6zzO8x7zGCRm+wu8YWUQtSJpDH
AAU0NdqlGDRP8gKZjDzuja32jBZOJ2kwZPKEuHXyh/MnybNyQxYXChxS5cktH9kuRUPTo2t9IcuS
xsuGmeGHd2AJ3jC2EAqTxkF0Ye6eAESSEYxgmluqzyvX8OzRirGgtfnj8vy0Shgafnfa7amwSaXN
RE5WnWuAIleYkl9Ux+UaOD4jC8YP0mr1U6rtR6VEw7UKuw3VpQkTJofrb5mcPCIaHEs9h6r2ISIW
Oecx8A26PBT2Yb/fNS3qyGVf29Zn97sVlc4vMoNOvfvtnW64bp6Wzkof1Jo9rihcDYP6qoIBMvZ9
kKafQkfU5e+nfs5/PbvpYCoVDnXs/TIvtmMMdjQW0kxZPPVAoEUH4eMghzi/rzCOS3racCKN5tlv
P3lVjSc1XcT5YAWq1FVYaQ5ErE6sLmoysx7jH8PmwusugOGcaTCJbVskPkUvM9pgwGxEeE/iJujj
bjtwz05FhQmhWASzcVetQHFatFywobN27sLa1IukBsJlODZ2P+zT+iGE91ThDDzkpnpaET7UDkjn
Vs0xK7hUPoZNj9GVZF4Ca2ekJONRU/oYTzUloKPHbpW/LjmaMH4nKlxh+AzUTTuuEU52BUzcuZUe
dhgWHreKlr0dh5L1s5rjQVxRNL44LfpkV2njX9fXlv15pZbZ8+rYe6d75JyliASXAAmv5J9dwWHa
dRt3IOOG5HgFG6nveAilQDHj3sZ/8DQ89F4CrNpvo+r+1ly2ap1og8q5cQOEWUaNkIcd3JM1Zz6H
3ZOdvJ70MvePt/Kr6PgDWnkEp1V0wOzRVvZTvvAyFRl84bBIjc2LhkolEH+2KXLZ/jHM5QYo7u2q
TIdq5+07keq1MVqBds0e//AolLPJ1BG4y/HYNavGu195h7n+mMpZoU2a8oUsfv130ACPAhkpcwL7
FHvxvLmY3cBE2KprUcufX5Kno1kKb+gYKuAI3ZYtjiE4eCpdaG/Gflnu1ookSdV1m8LrpOPdEbJV
riIl5uBrLdkie0TOxVWUYQYvXCN06oBBZl/6ckVM7fvyqviUYjkzUFtxUHxXwa1E2B0E93HfRg9w
hC4tBYbrb55EzhbVAwCn/u/VumfA6P4yentcwMaGDXA2hupRqeIpiCOhWjtT3hcXRTiSpNrn9LYU
81+cewBqJmlbCb4wtm40GIF6ZpnFN701qJ6SarflSGpuPqGh91e9A6gIdgcSiAX5oallHWqILZ/q
3jcD000cYIQ0mjY1eJ4NT87XPkstnF2RSyFaUlGVlA9YHCTYncrJcao+ZtY/JH7NTIxix3cGN8fd
lGPH2cES1AefuDHvsEzeG40WtqOjlv+X69TfqVSCFAOKEMQeFMIjFef96kOjKHuox7+ha9MxSwaq
0LasR/G1a9Ud2GLCxAm5mHc4Uq96enFumKVaJu4RVmUuipEDK7+TDb+xelM9LfhnmMwlAbFx9auj
vMJnSxsVzMiiNKnmAqsXC3WlSixOy0pTmsrQr7lFZ0TXS+aWF28b6zuAydOiUCYCVnzVdNFu4cxc
ja/Vw7to431uMWgqEgyyvqnU6S7o19PvH19t0o4m1LF1+If13/cdgZCjGlStof+H4xis5kKEyjYr
g4Gad/FikEm0DORvMJ6KP+yIUByIQ+zBboe/BroyhNGqMy6MS5xz7377D2jgF3D8tebDFEyFp8PQ
hGwMsyxFnCvllQWvpnxNgAfIvEbYp5opmc/6aAzqjnZflRxIxOUM2JW1vYswaD7dFK0nmF74D3NJ
j+8O/4PvY0paGIEblL6tp1OG050IgZ26787SAXqlKuLpxRMusWboVh1JeiIoBcWcvf3mfZ6CX9DK
VG4R2vNoXo6t6TgkHzLYg6OKZYyDGoTJkelFO5tqNQnLe4uZ2VEyaPCfD0zKS3sxGy3NM5cSfbts
awTkHNzIc1AuLuoK6LZJy0YgC1mo6JxYhB164s2epcUttIRK/bk41wepnsTSgeXlWx68qYJb8TWR
Vs10yCohQjxv9JZNQ3qznZK2JH3JQfXKM6Eep9x/ZsfH/hrOmo+1tfQs9svyTC6jiFoHQw+mxVUd
CbYkhTLiQZ5JTL+p0frU+vBdo35MDNFJ2MYkbVGWd2lzLPXU8ogkRg0O87izWaIfOiZjxU7JnkmA
x08g3KaMC1C5PqH+gyZ7bjDCGRUsezFDsiHbRP6fTJm+QoKF1K3uBJyzqDRlA2ktS8SNzj6O3aJB
nzaXR6g85mMxYtNTZckufinmhdpDMYMt+BrONHfvIqqvijElYKb9pHoeZDVZhGpiodnUTo5Zo2eK
TzbNigey6t77rhg2+L82/m/f0HDDduY+tQUrP2PTT8U7UhoFZZ4Y2Xu9xS586vUbK5G/jPbLSRIq
oo11Rn/iZR6SVR5CIjr19dOsr6y51Q/2DwTzdVSBlxUp7b7S3SgZTy0W8AKI+wRgvKB1wLqs+LF0
8TF63RrYouQqprQp74zzrrJjvIY7byKxfE6Zs8CRQf5ciNaVJ7pzNP2Sk0dxP2a0rFbLzTMJGUjO
Snsb6GKG47VtJ4Ynb+b1sIJWluG8Pu56b9i1d3POdKcPnRqqkHYEP8nyeBFbUwCOKcWN+zYBJxUJ
X2IIqtSm/hXqbik6fjFHPJ5BG1Li5pSSC2pPYK9VZD8cbc2ub4pNU+KGsRtFJMU4fbdE8PQ5i35Z
Juqau3c6mEnDBqXvmdOw9JP5Us4YhltxOH56wSg7TA1tdu44DXQYKoU8bsnVZb11e7imJe/B75ld
zgMdJYMd3z4Gcs5jZQaoUsBaoylxxQxlN5LyXw0sgTMOLwC8KZRmEemfIB6llR7anbxxeqJSlmOc
RsdlSovKmIpkw8kWqRIftMYc126yCX5TczGsz0dEl1Mu+2Lw3h9EcOgQrmMY0EY+ekrGJ/8x5bud
jP8XQ1aYOslQvjatQMnFcMUgIukz3/4uBYlIGotCroikPR4XtybsDvs9LLEIq4aBqhxkMP/ik+zU
ublEyGTgKnGgO4Mtr2WZsRhg8bP1vP0ssoxerhCsFQfB6ZM4eGE6WqyoXKDXPZyHi8bsgOuKBBOM
x2YsElTOyymymHrFzxH9vu9fl7ePBljuPM4wAlhbgfQAaThcPM3nsZNf5kWl7Bri3bxXnh2x/GZa
ng75oDH6acGKLwImBVr+qv2Nav2cxn9ALhjdEHHWL7vjtUawyQwEx25GJ0VsReVZWma1QotKOJmp
XvaGk/xRg+n9dXGQj8Cdsadf0pjtsJ3nYXvXI65emc49GIBZWklbbyYhbLdu1Zfu3rDwYwaM1Q2s
ROqMs8sEgyVx5amMpB8k/bGk7g3c9Ny7ovb3Qq8oN+jiEsKedlJh5av/2yW2Dfvy+eSoWA3vMHnW
wpXclgMY6YT6tmJnzDk/jM6+a6xIfXcvunH2zG4zRlOUIdVKfFaATO/lnRYPZrbaiCDAbhU74kf1
npjHCXtm82vDU/iOqpjClld74cTqeUarPB3v2jizZeTJraEx6QmyJaqngwV1wnr3y8aeT1lGzg/y
5G/GIjoYd85ojBFr5nerLsHGVsXZbC+4CIGuFVUsmt1sPerkq9AjR+YE/gle6Jw0wgXiebyoT5xo
oIJTTplc51Z0YOhGpKuklQ6m/I1X7o6RTOotXjeutzhBiffDjSA/ljwFsExdDAQG/7XkO73lUxsR
SPJhSI2QlGkryqUboGJhiqIMXKSQkHWrbcNuSaSq0Qw9xB6pWiD5CQI2uPlis+5ZyZY9rC+4zRhe
EPtIkhR8qnK2ZIVpHBo10s3DvTsDK8LAPhNFGnkmGsUL8+FDn5Q1vu7T44bswFDxTzavHgDe1jyf
v5uvu83NuCBdSlIUZiIwj5LD9qVkxh7EX1J2AN17nXzHE+M5nzDunmck/U9Gzltx6Hk539nGYQCd
QkzBE4IYi9OkIWcRBSEQ2vV0/md7bthX4FAogCI7tvy3zoxixRRXCgickDISHo8fG0+InBZiecJh
UgHqjxJNAFyq59KW5gOCctZpEzecIt2j/OHjdDjAsaHk3u5JPdl87crTPiuhBokFBnodEvpq8Dnc
ksogc5js+4P5+ekQvXoA5Iw5y2CVngFfIg4hUcj2eWINsdbwho9ByEuRXnVhCk5blgnIdBclzCKk
RqYE5vSX5aE1AeCOdpmqYWd35g74R6pGVqG3k4t/tJ4RFbfaaPxBKB8sL5u5f3RjLef3w+lVxJ/Y
U6MN0oJmtcJBkmHStfTOGuZE1KfMaFl24x1L0RbKWKn6cVqFSpYYUKLDYvAISAAXbpcpoMYNalQe
F78Ld6JTSha2ykQF0ar1dCX/ALTFI75GVrYHsrIyQ+yxB21wPUwEC26w7lUQHZUSfvev2Wcru+tB
zZIudNFdepUeSGnAVUFYl74JxM072pnA8MfrlaIxdh9W2yUVN//JWoQjRcIo1CVM2Vg9tBTJYoBz
VFCzMUpbyEskfx/zUPtXLkjBIpX7wWv6+FVXU6mTXju4/s+Fir7saNQ48qDtqSLLWlRF6ZBI8sTw
6yPUJXtyO4flm2jhT2aKyMAB7ky4I9kdCRj8eWaJmnCmY3+LjNtFoVwL61hvhMbWLk8ar1a9JVeJ
bN2F9rbys01n3xhJmL/ROFKCItmNIjFTKgkFOwmKeT88h7N3VERo7yQWGKuUDMd6KGtJvd5wLJ9U
4J56dYm5zx44E+zQYVSAMo5KGdlnVzqvWC03ZvwLY1zyW6utDewJE4jsjRfh87jTuuVTECB5B4Qj
OwR0TDx0VDaBnBKMagoO2DU01RT85S/KkrKhJgJRra6MYqvVk8EoaRmS6V6zroAPjJXn9jZFaZm6
pJPnt0ZQVG9ZQFuZSLTmOgR7pgDP0anvLFnH+JVeqn8gGPUpRFyiw75ZZaiwuQGBW4bzm0OjdwLD
mLKWwoTjuALdyS1tyKrYUAHg1li8dglgwxNwBmaD/2OshgJpUPbJYMwGgX7ojgRB/I8VEBwqQZVk
Yghtecpdg+PkeVQcOAxDKfbY0Kls/ruEmG6vXl9iqFs5AtQtXJJaKH21ZzH0CF9GIgaW5wJobXAm
bcpqJRq6zf0uTVzEb29unkz99KU+ytx086xXHnQUbTSG/WbB3kQ8RE9muyO6bm6jpxnB7VWyIukG
JM9gYPnBTj8axenSs5RCi2TrsYRKOh4HbLq90H6cdRSxgO7f9qHZDSX1zC+zejcIpwglmM6qe3GU
sVd9iJMFw0bnfmoG9uzCleIHeMqyM4IhNabIOkWSa3qYYL4QSlgONZDjv2dgUwDtPYA4JOGAqeI/
vA2xmRVf9SKfKRv4pXvS8G2hvrqF/B8vdoCKyqGDcx39+6tpK9PktvBr4L3hirWKtPbNsEniTb5P
LeK2TIyv0HKUeYWr//hCazDNLw6Ra3BG301W7H/gmI80zYVIwcfBMxRj6tnVjB9i0AGwEiTup0Ct
/w4vOCMnu6+Lzkp/RshXECNaDFe4CbjzvxX1yfgh15YKNgKFrIYn51Dbw6W4kY6KOZPUFDnqub/z
3/OJLO+0jGzp7/GOAbmmQl/QJ89a3KvrK4d4L85Zjx4Y5HriCyBCT/hSgI2DkYDuVnZ1jMFegeul
qSUvLDaafB19SIOGhh0YTqbraFcBIhU7sBEsjBlpywaJlS6oV1lN75Q7BkFSC+2LJXl6qUIsM1wY
3EIHVVs/dYI/VVH6SXD9rHoVBg+5YD0qcFe6KBrC+O2Uf0bGldhwyA2H8ZoUlPEAFesoebeSNPwI
IvRysECy+0og3LcOys+U5d0BKSwTEdiL6GKzhTPZ3wGlTMX/qZ2Ow2iKsgRDFtEM+PZ1qEsv9RYi
aLxZzGMA53pVTWcA5rhjl9rgZOpMgZZ970qxS9QuJwYZknvbev7rcD6FIdAYTXTOXrucdJ+p0AHi
8IrjmWEs4AE6pnf1OetAoipwvwi17+bIWLRZtsiuWSyEJ4D4BXYVvAhvpvNs7shgKljl4uHNCVuz
Q6N/nlIwQ/wsUBssGlpsmfSGxIclAGCFWz62BFHzARheMjoaRZfQI1VnoL0GaGbQ0BtO4KMZenaq
MZFrYnJMzWSiIGFfnXw5zx9EGvLFDjk0EPWMVli14d2nVC61oHzsfKHrpxw+ViFq2XOTmmrKI9EM
7lwAi01+IouiZDZGLLx5MJ6it1KCP2krLkv47GuPcs2zUb7C2uNbD+m63wC/RP7TbDwdLRGs5Szo
RMbx8xRyX62PhFedVZKY1UTsvVEZfiQFx5zJZ8+rHcwbr093mC2aKNqLsNm5IJPJC/rfO4uDBnTk
iXagiFbHHR41FJa1FGhEDib0lV9tyWdwZqnwAy0jU/6oVl1Rfo1cPHBoarDWTnlfFBNscwsWjBF5
QWzt/noeqLz/IVBr7aLr0f4IqS3ElSAZFlwj3znb5Xyxo5PhjFbG240sWurxuFKjXQSwIJFVLEFr
lCddaCilIQqoPnJBFlxE/5/9bn5zEGCIfcLYz7VF9H/jLp8S++UYLdgFLorK7yQXDp0Uvp8JPzOB
2RPWCWNpqYL4PRGAnF6QfZtIggDAQv5B1flb3XjQwlO/KNubTALYHdveYxLvBv7LXp3ohFYiD2IT
SdUlyaYRoeucXdFuXPGZUpX13LLF4N+i1/Yp/X7lNSL+3Id0c4YnVQi0/5UOpNVn4njdfNtxb8O4
lRyJERoNFLSdxzLCscnkozqTOuKZkhlJCn34w7K8Mv4xfh5LZTweTFpZ1WCTyLvqymABNMEw5VOo
V1uej/wU0QDYG4TqwHN/27FBQ9Gib6XsXZMpGJfFBjxfCw/RfgyXn16qqgxKuzpAs4X6NV0DaT2I
1KFCuAuEU/MBMlsPeR3/saiyirzpzXiqLw6RRt76urLQ0amncuEpL65sj8ft8/52ArziaZwqO+pX
A1vuMdshGu9bphSGNEznfqcDje8Fl7+qk//AKQbEnEsOuHLAPCqrCG8O72Tfh3Dygre7rcjPzA1O
BQFRttescO2FMc+tBKAWPpMrwWK/O9ar+rsN3MLN//7Kx6rgNpf+qPsG4urk2lRT6ErgZTRBhGqt
sj6orIsQh0xuvGC3FFF3QZ0GjWo1EPdfbF1o9bVjaMDlVxLTu4h7vWtdoJVmJEDMVHwwqu7L9+09
GMfdDS/ZJLMTw7f0rUdoA7Wh1Z67CQ29nXCvuMBUdCm83jI+OIcGnAnHujJy52CYqytANHvi8RU7
kAOcFJfc/JMlthXwwy3SEMLA/eAph0kePVTcoqr/0EtOPuIK7LVjyP0gAbtGxryeZhB8PnPIzURq
mFsKGfWnomjkCtWnb93d7akLQqHz2foa2Zm1DyHFy4NWV8Xv5w8+5mi2u1NQEip/q02GNHGQ2vRF
Go6mP6iDE8YjOtnO5SCOkEEHsSLMN7O25vWSL11AwYPgdFzNuJs/0ClqSQfCngnqypSS4XirsLbq
f13C4qSjVYDT0/D+3Sc6yQk/5TX1r9txFbOhPbk3BhDXIcK8OTLv5l46AazgRU37gYDZPXuyLqL8
RvHNzoPbIv/h/Ceb/K7S2gn8JwHOFa25BCfj40Eaf4/Th+O6wkamqi+3gjoNwGWGnCFZ2wR4Vl1a
Bev53zouRwIUEicmMVAQBssC2PCzHY+UJWoNdQBDWIVfX6Aj2dNIRTPVz1Ti9KZhkG4C+t1tznZ1
QxbTwFOlXnWS9r/MQzfa0m0lM3xMVTQXrREKZShbbgzr+MkGSZRS5BTlM2q4dH7SL96Q+DSvQwQd
pjxEk+N71ypj3wkNLsJSxXDs6jScbk883I3a38My+FMxrbKHKreKm8e3BGursw8LAu/rmXbWJh+m
gmAlOxMzKEW88dNsSnFwkpcL13uATXYLFTKZzVTOWpjEpPZ4YU30sha1TgRLcMPx7gQyaD1TpeRe
+HobdfN1ZusWCUuMjqi4BDL/1cLseZQTcL1zMob3AMv8IhTm9c9v5BBvuxwXKId5Oe+UQ5WOZTKK
Nbr+S+Ag7c94G4jQtBPJQrjhSSZuKaFVbv4NGoemijIiWbnigtenvoWpS/E2gsy5MsXTCId7lcey
Nr0uD1ajwSJTlDYh+VylpCDXGRU8uaY+RSJGTMLKMLNlUqydpai5nv/Aq3aPG88s9IrdwIvWdxi4
EzMFZs/sQK/+yvw79gxU0a7DbHXX/oOSMLPq7nYXo3zPDQMGRkboYZXcDXIR27sahzt2XpfvGUVP
5QS91rnysxK4vHdG9oAdk5zkDmqZd+I26qAXlog8vS+NBoXDCSZ8uQnQ902NuDefwmXxRJ9E2dzB
KnGVFGI9Nmd6eDRR21CTlBhQG3HOQ1rvvge2YK6iGmszvIi+5Vrbh+RPDiHiCqY6CAfqWb9a0W2K
JyQl2afjH7uxUbG1QqbPTAxDQGaz4DXdh1O/12YGcUzonIHGJkVWurck7EjV0N59xaia2ZqEfn5C
U6ueCsM+ZVnXICuCAub9Yb2zbe9MfBMyRu9MMG0JcgD+uvLLFMdOg6AEOmrnQ7JOxY9GBZ6/g1Xp
MZySeeE7Mp1tNlDYXJwDHkRAhO6uMk6OzxSvt8owSnx85U0kfE/WaGIKTRxprXGpBnhtKooSd4uF
0MBfrJf9Wqqom29wEv63sE5Ao6c4/+6joBgcq7UAxx1A/YjL3kvkKWEAktP9FpzfVWMyBS4C6pVW
J6KVVA9GbLcxdHG4eb3JzCQsA0QMlyl64vTd3/+u3YqY9BRsiUQQnn4lCLtMTNP079+CVNc6pGOo
pqVmWaI2qsCkFwVQQEs5aoz7QejSjTExvWdNBGTa4BKPZD66b89wFAbZps5zoIPxAeyoy+NlqTZu
ikoZkw4H8fbuPijPzrKjVzoNOlBa66bG6IZraetSxcTUWOvNdyQvtqCvaGwiM2Hyw5apjGrEiU/Y
4kiW7oWWudVKbOy5Q/r0JCROiys34S1UKFu6HhlS0zUczJi9uosPiecD9VsSlyLf6CSqIt/BmcC3
O35TCmZLjQ7AY280T+8nI4nmYK9uh8igyTnpHRYt6iEtvNyHEoPTwM/qIwfePwlvo1ub4RdG86NA
FAWs9U6jKUowPWKCI499a9v19m+vBdBa3CV1I681gIOnbMfpZJkVnPcwINt0j6TcsqcAfu6HYGnV
oEl5oV1nJIKWRQsEJDwRrp7H08d11NJuC5crUAZv5e0wDWbWxXASM7zh+jhmHwZ87qieX6NLtNc+
T5XWDXXmgil9dp+9We+dtrXCmFbdIZi4UBkM1xiUQdD7xOy+U+DC4I4/l0N98ZFm9LQVXdkIuV+r
yF3ltn1qIbc3xW8qFXd2vIXn22XDYcaYYyeUsi73ui7ogUYPUYQOB2RzA0VKpwkbw4frDb6PJ2h7
AuCDAc2YeJs5q2K0n6UGmPlPTR6FjH9KnMURAF0T9TQ6FYfiHb4uqzJBGH2n0oN91Gjnccj9jbx+
rbiICh2kq3SmeirO8KyVWwjNBTKbGnjaaVC11qDswuuoQYQxC/r6fYBMuCaCkMQsrk3bnrPTNwNR
uKgghdQKKgtHxz50+m4ZsxJOaLna/58x9jiSEQKVgFf7X/YGA55/R8ZNC1epssjQDHfKdD4u7KrA
Gk1yh+APas8TrkCb2tLSilFI2Fg3twci1esK1lmKqp5gWzzt0EBIbeAAehjewnIzNRjD9ua5CE0r
nP/J2DnR/VoQjurx25KbnnsUzuqJJ+F0GB8VXLbncxgWyQ+AzoWWeX+wPIwQwF9Ss5Bm57GGnc/l
61Hn2XpR/ktCijQ6AXxpUrKWWlrnM+zlDaULJtNq5Rmu3M8DKns4huKWtfJgmyVP3SKy5HZN4SLJ
HpAkEi/sLl8CypSM2UcHm6Q+cgBbUT1wc6dhwG/TSP1NMCgQzG1maGW09CIy5SN9Mzl5VJ0LcfoE
i7Df3C6R9APJpBlz38tiMutAR+5tgmLqZBBuzQoW1eoLbVbr0TjmJzfpfznag3TpAvpi7iwBNtdt
3WVWjUW/W0oaGGF3swrCHOXCecwdKkk3/QpOIKorD5oZZgKoLekBoZrR7WLh3dLNM+2If3LgrsDL
nPIbw+/iVHl11qLXBqvjVJ4+nIN1IHNO7IfWWRRoXO+JKjN2c3ZKMsV7D2kEaOx/SYkeVPiNcc4g
8dwc7nU3a3nEdDjM54Dmv6YHH/+G5FVgqQzwyKHwST85QxDWP/Sne+DorcaKbJp5e7h1UWwxRNBd
+acPfb22uYKA0CXNzNAxb3y5Elvwt37ZbVAl7prS//rh+JPcTpQ9vJ0agjqcRzI6E8B7IWMldhpC
toK/BbKJ592SjqqHkvH3pZzN20ASg0Jp+EFrCxBBpQ6IDzj+ETpTmMuAPGS9DNbp2CCUxu7LTZJN
5GNJKoSJPI4x3iqztFyQuP4vDMV6FQ/hbKQ8cKIH3wSQK6KEWPO4OgV5ngU9fI4LD4VMRuUNdGC3
TFnkMab4LP0ZzclMZV4Q5dUMsKPfySVUCGR7siLtW/Qu/YWn5jH8GOQqIvTA72sIy09EIlVSrr7p
HQ9Ru+LolQJQp5wSReCkPc2k8qbapnnsycQIDOvxX4n/+mB5H0uXq5/ec7dqqkVISe7xaiUQ7u4x
N4OkcLb5n04YJyEuwGEHBrT5ubghC6vp9/bNiLu9Y/v2qpEYnfzXMqUyyLn3rucpUPQvDT1Np5mz
HTIc+BCLsb5Lb4MAr0q4QcYteDPzkNj5sEdD4O71cJthf/uGCFhxnxOTH7/zGLDgXelceVUuUXC8
Er/SuqKNh0oYRSGlWiP+haqOG6D1KrZaF7v+L1cfj5e/iPN5mBueL2s1GhnL+OuRjIMYlrni+VWM
qq+gfYK5S+DgAsf8vxptTgZgp1+yPY+xtC0Y1hrT2UZh7xPIwsEaU7EkYXNTGf9ApYoko8Yd878r
oXIEX/RBUaZNO5GS/l2QGf1EELr23A/FMAc85l9KaYKDuWkwLwEb9tREHB2PrMVFxsr1ikYnYMOf
rGONg9qT1UTR/enN1Rt5CQ82qRjh0eNlj0gpQYfBwdrVY5Je+j13V9dQt9oxiy8haXyU/VtwhDwE
xzciy6TBsXptzbs+1zd7V+IWOeo47zG3nYtCL+Hw4LxQv6KN5NdBI2aeKvGQUnHj7jzQ7HSypZSW
LXB/77fLFjphZf52cd080lwczdMaPXyWD/uPgnoIcMOpydqDi/iCb5Yu888L0sVdxKBGmtU88vHk
pTbGzr+aR6Tdh+iA8TAyTIaaHfbkNwcfoMYlLPgl4D+K9Sl/o1N7f2ArYkHX/1fVJE0Q1qAj/9MF
npr6A+qPMbrOFEasH33pv2H6bXRXPaveUdTIO0QzvGSD1dNoZP0NDqgYqSJ8kxeGAv9EI8NCKlkT
+Wj1nOVOO53/HlZ+lyrzPHS6Gr9lUlySYVVtIpRKSHunEBW9b4XU4oy+wIg1T8XrOCRDmkMVUwIO
pB/b8KJgUvz3ydNjEY3SURE+M5uMxMlE+y3QYBq43rX9EFMuik7q5/8uXh/YiHmDeD9zRB7aOjqA
R7GpP5AwOsf1S581FOxqv3OqM5LNFqLnYkSvGjdbLLRXKl38zrDrQ9+z3luiPQrgv7dV2IV1Mc4Q
HQl8/myqnUryvHyudJTw8+jSOMeU2gP+5IqMfWsTKJ5Ume8nFvVKmAVem9tTmQ9lOFH5iU89K4N/
26Idk5u49f+Hneji7xIjEa4LVcV9fk87b7NwvNu/LLhkBUR+4O5Iu+ORlq2ucx9YNUf1GKMSIm51
x6HngUo11CB7cWtohyqOCerBaz+BX1yYgS9JPMEj+LQVP6KTw3B1JSticcUyr4dXYwinaznAtnBi
TFXRsRijXubrx71vRYxwmp5iLsaeXXS1n4tQz/q0X8k4iWHaVO72h8wMhcbtjm7WU5Ij8UQf182s
pHChTb8kDGYcAXQnT+jJu3SZfzf2DYkVk1Jylu3bnoDjm5QY9sq+/KmxvCDMqtZKz0O4xwnQROCZ
LknTeygitii8WLtQqPVzNI0F/lFOdHJNZob0jQue8aOG/QlddrSzagb5A+iQmAWBrowvWNwgZfJE
XNRpQ9faNyJLho47/kHg01Aw2Bo5GBSzhn6rxYSfUQOD/745IcEF/cghHWRaagk1pUbYeBzldoQX
f5jcheehoO+7olEXknYfciXds89A1/Mgcqn7j4xlH79/Hgbi2xFWBJelFk7KqUCaaarmYhZLI4yO
BNu9bC+51kbRL3dFffdcBJTeAZz/Y78IHJmNHpPCAa/G1ETD7vLLbzRw9b5yCyWy27arf9A4INea
OvNsIfzsvG+zYEfvMi01HOqDCqsY40CQHf++Ek/Stsvo48OEMna+Shi88C1VK5kFDzZVXQv6Kpes
hw6rJcYvdmyOw/Gk/WQT7eY6wfbgv4FyPMkLA4KQe0RptRZtEmqmUk+1/LfX2T19paPAFtcz1N1Y
v1KYg4SvqsMU19ImkeJ1/9SIKXSTbUhFemBdQcVbHLSkMMTPfioHTM5gQUhtjsZSPzIVSDIBViBn
ncw8enhwzYxN2wJS1kVW6+u0MSnpjFZBcQ0uaxqC63Lw1+WOaAi5ZFjrz3tncQ5PMvRNgQ8/cqIj
XP+cUakL6x0bXzk9ZOYf+hnUVvj3+5CTjE5fKVYkIQM898lzO0glWP+gqtj0uXSU0n+/FBHL/c86
kmCEwguQuAz4ZyhzGndWyvssl967O2QU7U7JRBE0T79bmZLrxLQt7x/aCyDnkFSBV1NcNvG459tu
aJaUclOk8OIWk2jG7DrVAjFTxY2KNf3Aalyql78jYhuf/wVAv73brlHk8A6tambmLhZaKcunqpzk
K/O5c6uCGLFQAIKecEwUUbeS2sqY1MzeT63rWTKbtUdeQu9BDow9S1fRwo/K8aU3Lq80zesVJDrZ
l3jBSnuGVJdvVfcfySUTYoR4CJNARgcKsmtsEcVFbNchrduSFRni8KJnPkl1LQTvXrTHBv284OaA
qe3A3xRwfucygGAqTXKdjhzprsJUhM8aW1/HJc/HTbGyTfTQFcoR5ZAlBdnNLy0P6dsteAJmlxYY
uGmCO44udXRe0TjWxHPa4fGfsIlNPBsmdEhnJ7VqsWLNu5yKozR2ewlGVCYUas4orEZ4NCkVxEiF
tKhF2tzv0UkDWv62XjJqyObwCDt7ZGhFQSZDeDU/d+7RorlnbQcwop0jv3FFrsXKILKr2vG/AL+f
5L8zeWcSDfgPcRfemxY3vEeMuUrzjwnucp0wRjrsfn+EAIoiGjHcYFXkJZ/daRS5lBbBF1hy1kqV
ZQ/o9WbjWHs3t1K9oOf7iVveSkrM9aoqWEVPZzEWjKMK7206x+TPn6zZWROvZj8VlpH5E7276DhB
av5lWX8Q1KkWwBexNTXtv04eeyzKwjayjvyBWWeXb2pm0sPa1z6KZWBO/xibnGJMYwxnq0BS6yUp
6aCw7nEFvWjwmyh9uT0IOjskH6blNXnkF4Pn82dOfq2sM15U8dwfqb5LaCZApAGVRsVsh2Yelpgr
ONAX6F/UYz7CKef0sKUQbCT9/GOgV+iNscaM8jS5j2ErQzFiMhHkbxJV5YTMefrbEHeNamctoseI
YZXLDC3gm32pNIIcnZS18i7YwSMM/dk799P2y0WUMWnj0+HKJaFv5fHYsSi+l7SH9Cu7fWdUX1Hi
1xo4X0h7Utu7n8QFJCI5iZefBfolCgvd4pfh2tyHcq7H3smiEcnGlP42XlENpVjB+OnF1MI7Mswg
HbKoRUJ+nrXb8lg03bDPeJIFjk7vjo9fl1zqvrLOZeSNBd56UUTDzX3MfM8HRau7J11Q0rBoT0D8
RK/+Uz/pNcXnsHardClx7URNQqJGCW2cNhv9kZvVn+leHSM4Vn8X8iml6LMs+qwLTY4J/LSt7qph
WRNKTd1S+wB/lab65ZJDMZLYadM/DgqxNkDjxb8WOfe/O6cGa2cT2jNVLg2jKebVy/vC8dPT9SeY
rIoad5kPEKzL1KNvN14mYCHuxkVjMAmkfm3SMYxpAvOlw1IseBfPFkFKBp8TR01yACe940VJmG6U
UJdDTITc3wo3papMqJqf5IlatY/Ve7pUqZNCTYJHX2HV8nHuLbDk71jopgLbSIx6k7IlaeK9umsW
mv4kIkziGpwzs8BXo0crO6iyyFAeSJfTazqxHNHOO3s2TLzE3nye9SEq/+evcSPqcEkj/GWJj8+D
s2tKXypl4jvZ8DeDSoN6Fl4bB9pDL8W15QaGW8ns2vnuHws7NI1b7n+0jez9SokSnbWevv6UOA3K
m8VsRBdpHsq9gjEw3yNID0lNfEmJY3gLhzI4FrrWwAaWCXj/k1anSuDESX0U18gHeyFyaudSI/UD
cvTCwDEPC4WtagN1CtGY8Y8v3wEkFYyxqFCt1l6r4vYQwQ7eMqsY3m7zpzUSHAG13f1jIpVOHTp3
UaFo0GeF78SGOa4wI438OXyY2FeKXqTnAgl9IXNoxQ9Sc7Uy8FQgJNB0qVaWJ0Ay5UpkrHNUzH7g
KEPxOXcqnmjQACjBpyySw9BCoKwTvunX20/+wmXEMouyBAWPkONRdIatXbUBOcyeo5zm7sF1cYYU
47tNNxzG5e7gUna8Qx1Ly8XLOdSWqrudz7b1z+eKPUTC9tsxUk7orCVOpY4Om/wthN7M6uuszXbV
yu+7SvFsP5C+n7k6y/icMUjZD4fjLcXONrPrtQMtFkbiLxFg/OUyN4jnWMvTJ3KHrYuBWWP9d5wa
NdDzjl3+6P7yYZmCBtZ/eiXtdNOFivJ5P1o5OKtRR0zFxM6AbGwB1iak5KIZDc422HzhKz3lkkp9
0EZs5tBiTvbEvWn0VYq6AWe3W/fyJtzejBE5rYVJl9FfKNhWH4J/+BsR4/6BgvaV2V5jD5zMpauE
DAr/+2DmoW6Gl4h+rHIQuR6xFJ5nq66Mi7TGFsmW1bvSK3pSTIr8ljyMtaq54O2tkutGUubN7lgI
Y9G6z2KQfeq96jQmfHJQOD4LwFypzmrZAPAC/1pfyJVfdTENt932voUbL9TRFDzHhE3LbN1OgDwv
8n+SY+K8ObtIHgnUtu5CZ/CHEYKsRXviN/vNUgIorXaz0cTtab/Z5GGWmIoKlhi1x1EsHvoLTN/x
myrL/PvBGUac3nLpxZYBbZyVwrTnxEeiBx8AbLjtiuoFQb7cpL7xcr96+u4xVdyhRrGBFJnPCjbB
xD8nDT2xzyYLafjMSnvXcRzJV29Dn8YSPAP34Bl+fbKoLdc0NjqySLuFFmVSNbElnpYdhZ2a9ePF
cHrXvhKIWTe4JsCS3na7hUp0JK6gCL3jLx3yv1gfuHU1hyc1NMVOSUf7Z5wOmZ7LuO+7wkWBkwI0
3iRP65Mqant45apOZBu5aQ2jxzww5c6M/yfPd+unyzAb/VFPld0LeMsQZUwxDMDkdCP4MHy45cKo
kqzg42TCGFocD9X+mYcNZ2s/E5397q6tx9/DACgwrGFrJtjTAykjq1Lk14Gw6kyWP623ngemogFA
zVGlCvdit/0D35/lZkeMKn84GJEs1PEsHnuGVBYDa2me4eIiJHiTUHHXwqW3ruPogL3PJC0W4cYV
8H+JyIs9/VUXJSJ5cbsYZ8vYVN1s+FkF/OVJpfd+nKq22VghMHm7+qH+V4wLeACE8fEiA13P1W+k
aFcBq6PIK/Uss7wd4ws9a2zYzx5W8yHAz3X/XxNSir3pS6zpZg5V8At6H0j/9aoAzwZaUGdD6Euo
BEQcO6SKjQrfUdTZcx/78v9v1D1MJZCxjhfXKBuM/GTkHt3attUAEBXr0eG2cZDoaRoZE9q24USO
9ogRknXHJpNK8eZwIhfEy//mYATh8ivqJXKrHMr5IfbeR/2Vd4kOoevQM4Rz3zho5XTC2ZGFeYq4
Cru5ie3YlUXVzjpJ0nN0WLRk+VqmQc5UYjOxS5TKpRL9rHvyIGA1+03DR9cFLu9taknAx4z2BDmQ
ISAC1g7bkQmZGPabEFCa0EMmEQcW51QYoVDUytp1pb/b0Un9QbBtdL8B9rQ3YjUfmXwoZjpjr1CQ
QW8VFICFqNxryMopzU+MXU82NITbA/dgKcniCTMFwoMmWUFCzS5g3l7+jmh8/tF5J9X9S6mJaOZH
DoqxFMA0ScwST9oa6/5qNPX/uXwujbtnl452Zl8eMT++BRI+ofzLsYaONFeTFgeHQNWNqsbBagSY
Xn8IfreTJf/cIo9JiL4FlO5VB5wBJS5mUvOePyn2MYT+JoEaz8v90oJTUeimHm6Gki7PPmhgx03c
AcVcCFRuPKLuch0uq1dO/nbCL2gQBaHikH8e1nR9mzmYj1bUCgS0j2F+iAZo90dyOSOYt/P54P71
yj6MVcJqvRRSG+AJR5qIOjxMfSP7eOlOiXTi2eUA24sOqso/130bP6JwW0kCkfaDSnYQJ419ndP8
BfUyVqlGg0Do2b/DlFGl/mzHaW+m519XLD96IVBKVKdWsyu8nqzepXXximcJSWcal7mEtbg6b9R6
udrfaOqYBKfK5E2mNqhq4/UWDYnoZl+I/al26krjvyBcNp0QKmVBPE2trElbQ5PtVtE60shF4zaH
QWZJXcygG5nifGjMsmAM+CitiiKslkvsGiip72SZdw4mo6HaRYIrtu9qs1+HEplx6tgEn3479BDR
ECNvQ2xq/r8041ZJUD0P41fEhvFPVt7sS+axzzE7Zr8sOoG6n0trA2uo3OGpIWIii4dcXOvaEgjY
9ACDpP5VrXETS43N4qADFrPJy4pnxOj01sm6EepUB8W5WAk+38zUj3OgghX+wJrIWSaehKNJOrIg
5017vghv2CbeAYu3xK2p2hl4QaxKxuD8ewcqH9x1HD47U2aJ2K+hSi5C2AICZNwTTNdHLLVL8qoK
Ad3sAUYaYgrv2og80jUpkt/+m4qfK1vCnhZRd4LobdaxDVq5MRViwKRiLyUHl11BFaVyRtZm3t4Q
Q8HB0bBU+ET6ZnUeOMfBdFvWsh//wInXOl1VxN7F/2pttfg6x/qG8P/T4VxcQdFMEUave082m+tl
IT7sjpqvjrRQBM9tEd9aORz0VTQbXcrEuX0UpOKj5trUOvzUaot8+LPNdWPl5AM107xpZECDkhx4
B73Oe7D+1qY9pZzSxitPT/I5Duzd9U6TyqmNtkn9svyUWZWXd7y9EYMxH3RXK5+pd5L7q1Mw8hl0
pw+8lbiU2Xtu0DZ+aZHADMEH+IziGbEW8irqchFim5Rntg1rwquon1sXblCqlzyj0DoO3OZBzp+/
4HOt5q2PeGkw5r4kiW03et8OSYH6dUSFt88MZX7OMGcGLp2aO/cjlYHpiKOVANpWB9NTN87vPh3t
aZp0V+2RqSz08ESgfhQjiW+nPpeSQANvoO67/WdVFpH/mFzR6MNSdS5ijtr5SFClX8PV1n7J+rHH
Uwo9oJwEIxw2tcz15+18yozR5ipPtqODVJFdHylacl7Izgcolq9Yhmu9/LDbvfGyKbCwpeIHTWME
+/vi8/p/kwlg3i6N/fQfset9NSNyLUnhc/sA7wNoqUDltEyYfpHrw2J/I3YbpQ1/98ETncTyDQ8w
i0ARBPCG/23daROiWDsVu1JyU8j66atNhwYzoiOiVtN3oCmW26Shd3p1nrsU1jWT0v+m76PON6Mz
DV+O0pkTsTfjHS/pGHpsmOacXPxWJYBOdyUPGHP5mXHaFrFwJCzBVmSLvO4VgO2R3Z8TBYKJungK
cSkRT04Kc4egoSaI8MobeOHxmoQg6vbZR17q4cuyEq2WzGF2/oDuVgF2XUiKmMjIcDbV1xGGw6jK
cP/jVWhlC+Ji83/saVK82cnnjxAQIWgTCvdHXuFxIyKk8NigaF5O/1ghQoP7aFgjXr81KQYPWS/P
iWJEGohEO6BvxhVNpEr4OoT07RZilNUJdDowu/yKS/qRxyuSZGrjd5X8BRTKMPZAMuXBm2CBHTlH
k0MtiI4zTg5Qm87tfGCTMq9CskIs3hlKd9NDp0PqLQx36B8bU3G2jduQVpXbhFa1aHkBA7TRGBIk
OLb7GeHO43QibH/XnX9/d6XrVC76+J09afL+qSuGv0R1GITxz7lWSylHr++3CBjg4yzNHnUGuMtA
xe60gFoeFpQw6Y+UD30hC5OMcvpmkWhMR3cIV0QFTrjFFRyDGZeweInOx6p4D3ZN7yOzKUIwULTZ
vlioL+fRGC7uLMwLhAj/1ZCCn4FOw/tl67zBTkp3Jw9/Ll2H/oaniFzZzWCJihA4/MAQqY5zfykO
liQwdSgJUqL9U1AXuDnWCeGmU+NhWNIr+vZWIL55YZL6EGpkEeulwVqrq/Ya428ZQlJCJN9GXNhz
CLpCvSWj267sE3tMXeBrZZvfxrRWQCM1IO8Q/FCLkyo/ViQSBGqywyFpc9G6aBBwkGq9kdLOJHfV
mtMRy7ciPDt0Zy5wkZCyaR0lskgPstKB8zptjJi5Ulbj1GqHaKb4yXCE1PUe2Bf4Ap1uqgDChUJ1
+0QcPHB6Q6ky6Ha29OyGlFyq6BQH3sqQO3kLopBGkZwXavJBojKcF7fps3HQ/hGj4DvrkhS7vthN
AREbSz05sEOfz1Uc3qHhN8ZbO7u6JYXtOFYE/giOf47GHgpQN9NMFfzROhqPAbUTRkGdPBT5c5J/
oK47ENwRAnkl8Iv9IXeMFCNxD3iDL/fuybu/dhn0tmmpxVe157h38CqkUnY2UwqnM3ER7Q2CMpEr
wcb4lieJNB5NzJ8MQPQjq494jusaE9/bol7ulPWyELL6LNUC+TGzHXnEpq+efL0iwkz1obN3XkdR
3AeyKjXCwbn/K7AnUj7S+Sqzb98qMj25eYQi3/NAv1bVhjuxViG6Sm2A7MGVz3QBmQHKjOyotaEs
lx0kId6aoKbyhT6/oewk3B6x45YSpKqrDZXPunrpGmsKDaORdjGpw59mtXA/Snom4CT4H3dt7y/K
OPCwezbjEdXpQfs7XnbRDrN+ThSD0hvOcPUrEuKg5lSGR//GWpZHKVYusJe0ZqZwpj/KOCtWEWAf
66y8+fwon71cjbi7bLnWjasnaCzj7pqIhOE59PUhTkpejcwly9cDNJyOc8ijxFmZ7uidTW9KDzmJ
FDoOAY3+brZKl16uGYaI11h5krSkqDl9Tu+enY2uQOzyNMEnTd46cfbGIETuCd0mEZYEhRpI3u5P
yjjfVJNbdCWarvw9YL3h8bGJBRH0fZVEKlC0rhJG6/ptBwQT11hM9N2uMiu4B5fEejFFn3DYx5XV
DlADUx7gw+HqKFdDQ043hB1coU01qWKIANfnHptl0e+tAeF+YB2eYLbqayB73dtvJbENdUDmNV84
0KFFt+dhBTQiJck6ekj5A4pmMrF5TbSo4yN2Rv6ZWEa2ACSBWJC17/gHYNdxHsJNXV1K2oAT2usX
IRvGkzBVXWm+AiLHxCwTjhA1a9hRPXtgtDcli4jmoKifLuYZQiHQm0q0woNAUEobwn9+oPYwuUmQ
g0oMCyQzO5b81CEtslOAcofDD2Gtry0DOweBX+hyFoaB1zBd93E6djdj/GmEMZ/NIY2towZvCDh/
+JreYeUJUfJm/RrHwuAfU6HtL3eTWPFjOLPea7oPhQrjZj9zjrFkG+4YTTFCFOG9OViv9DkCg0bE
UD8sImuyvxxHw1G3pNYxox6PFFK/k6X1yFgyNuCQ4C4v5buZwG1Z3Om0ZGSPCpfP65cDmdayFLFB
KINzMTCw4fpdGV36fwDyC8K2DcqMZoyJl+q4GmDyvYN8kB2zUNL/b6p052vAQlLvIOQbIMn7/Bta
B1B9OwNd2QuhS5Q+5RjgU/o2my/p3w6rApMjTewK6K4XHhli42WFqY44CcgAd96lsgksywZ3C6hW
bQqh3bxk+7cSDffUMAO/U16aLYRMvPXEKhf5M+fWx/51lsLRIFtzEaEaWPy9gJTKVapb5G8T6cpb
yMrXhfu+tJ/G+dW9FIZkIBV7oGo3iEK2HG/Y2FTITsU/+N5o6EHWpOJ1CqYeKmrSlNL6Hj6IYLv1
kk3fbOZFcasMEp2Ya6h1/yoa23qynndilRRDcMkvRtU7j2vjvj+cAeONu0VqNDruLlNpjj4lreny
Zogn47+bzPtQXta61baGq1grhNm2QGCeylU8B3kbwHogcEMSthFYN+lkfmmsGQjhcWxatVIWbwsa
xOje52xBbg7GAT5aREg3Is5in6CKrqoK4tWBy4MXmH5AodJe+fC1h7xKi6cnm5uPjYYdexhXU0L8
sCNDFWl6mq1mUHyoWZ7Y9YkodNHqr0Ubqo0QRTz9GqE3aH3x0NbcbSBYPwgxAipAv7WR2yFvMIg1
q4hI8+vOZe78hbX2ka+6tJnPW7IAX/iN1koXV6RBJ7Ifn6fhISt2osb5YBLZJjV2OYXdVE8cxyb3
eCO6W3n6sUINJ4Q/V4ymKxA4aCPWcYZQ9TlkikcnmiWxH0qPZQ8Pt95ZkhtEWxXLKsOAUgMhGH95
n5R3ZSyfPVhMYZG5Tfd7sk6VKH7gz/hEsKchW/vJSltEjb2+V5UOtdYgATMZQ529wYNwimoqcPJp
NXMQ7QWC3g6mxk4GLZOJ49jD73rTNqoTd9d5QZNJBv+68wwzjLQIDgACMZTe6NamsvyoheU5PSTi
DgKucG9DVzVTjPnRcnfV07GI1nWS586GR6eqGCQDUv7OJ/vuni7avOdwfCD+XZjM76EP3OdYmk+L
YqqaJjWC9e8lRFH9Yd9S6qM8HLwAriYIyT4nuuAcWKv4FwPSE6g1nf2LkP+fJhIPkAKWToBUhh/m
YhCBA+u3eXdfvwG7CFlK+24invChDKe3BtlOKCvhZN1FGes/XlIDLBArsJgy/weHnm0KspugniW+
AMNaZQ8YCykgEOf/Yha8rH7bYBB1Rlv3zqYraAdvtmRjdLebOPcy1u95eqARf6beFCQWg9Z6VYhv
Jpxw9n+vSI29a7RALGv3iZyw8v5aObLkcTReLmfssec4S+T7QMsvNVf7fu0Cczv1XAFtMayc2oKB
cYSrpY5CVD8oBmPDe18lK3wktf3s3/sx7du7sViLmj2/F422RQginghFAgwBhpA1n3Z7xXE6P4Kv
eA9vJGSVTESV/OiT7eOoEydH1zy0AJ+4zwYRtOFdFxbZqimwxgrvo8DD49BjZ+m+ONnoN23LBzix
Nop4SWgR3Y/Fta48gKFEjWkavVlpQ5oOmS3FuXwRSCJVXADyPDqdoIp+3BMSjS+O+1zA2NOS/Hsb
CGVq4vtwRJEQunEs/0bZpwIp+zWZdiaHEkMLSzJ3/gsjiyhoNOsMxu5goB6mcik2KGBPAL3QeRys
/lbz8V2v4Oj+6ZKnQ6ui64A6wrrfqdmYrP+S+9s7G807IEtWgrbekiMB0yQFnqEujEFCj9b4HuNi
eVI/LDcE2VqkX+///D7SSs5qS4/Ds1+xoAtTTEqXZHaYLOSw4sGTQfat2f5iWkFEMnxMhwC49h2y
oOvz5tS3I+QqUL8Le6p91wNtnbYSt/pPQMQysrw2rXdgzpzrrG5wOcDLvakSZOwd/dzMcrJwL1gn
OHf+mO4tXjZjL7HBu/CwzhVg4ZptPimmcx8eJ9YBWRQ0LuwBUENQeRcCgT6RPCNuhYLgUyDbgrbL
yL9VbcvJVl2OT9Dx5QXSWP3SHDChw7tPZA8UVXDVlheraZOJkHiEO8bo4ui7PxSSeBbkRxHfaRPy
g4r7tgxFmq0yToDOcG1YJlYzjgxCnkbu7kjZlzmDn6LHHQpJoG0NOOAZEHcRoYenifPCcVtwpc4w
W2ZxrGWHMuCM2drkD6QKyFrYiXYbloOQpD0LmzQmuvuw/zOlr90gJKky7A1Jm4FpWcqqmnRq2bl8
QGkS0JFDfzQlgG4SzsNoV6zNxNt+QfAIgoF2bpYAt96+LcB9tagaiorlhVa8VzAbp9VupfAlEre5
FRqhfmj1FHNd3s7qvHNjRWTMPtVlpT3+ECiyDV80u19fCONP9UeXy9ss4DSrxsGJ5pADlCil3QUb
Bhs71pIcO60A0u5AxLwplAvMUzgdIipmGeUyKmoCLNODq/551nDdrpx+myM3qTyZbU6moYfil7MQ
hPo5pkqhFySlq86nKMRPTt2tPVWAB7s8vK1lzTNNU4GDDU29DFBE4J1EBK2bHtpurg/3LORFOj/2
yqfOumzDWNluo/edmRBlS/b0xWVrF030xyeKDi3dVqQJJXOCPIKsTKDWRafoINRQAXBTsPfu+WLO
jUhcbVnFpTfE8UfCmHvvRkqLXLKaHFOemG3vznw6YVtMsW/IieUsbPHc6ygSlQBD56Qy2iwq/clv
qIJoHr+DnH8iacq5zWsEDM6YVbEr0fZAx/yoCBTot/DiqHUNUPk00DYcQKWIEofw6hss2ffhlTzN
pvWGQzVcbAr0JbyMB4FuHTKV+ySjA4OaqisbCMejExZwOVr23aDVxsEvEwlsFn/3HxKyLmJAhZq/
sl0e/iOatpPLnCg9EUghGMchFqT3qzjrYmDAe9Nc1o8QasQQilVE9x0Wglv2BW0BAxsf8aEH1HOv
qwTyB0HLjqeEipp/XVkCknrQwF4MxIMw2XA5IQO8BkeWaLeD7wPBZGYuyj0VJCh3d4n/2lrVsVQj
9vBPUjJMopcKPRimGfyCQbqhYkgRKk7XO4ZWonTKP/PTdiX93hhGDGL3av8UtJTd4MHxVdwn9zlj
pnou+uhbYZT9DNeAfFNi1+GcmwUdRyXKy6fQ6LB/Sr3AkFHWsxRtXel2iE23PPJyWZQukhTFGX63
Nal7pnvL5B4e7hKEfz7qwb6yiskMQmURDkTI6o3Q6Tcxsj4JmgjApI3Qr9b+HZwcast0wlV6jDnK
QjZ3xinV7DBrNojAOgY14RIQ7WKbOlB2GD2U0cIcRtmg2ZgRr7tpobEzfgEkit4s0DK557NQcRq3
SYO3CgZFbShmsel1jtURBwc7bY+GJg42GKtEL8NAvn3ChRhPnSeAgcemfVBcvROZbjBFAJ2k/1bd
vSBcQOyiopgNRw351ECQNz4J4bqK6ULJmkFdPVPELkwFq7efO2k03BBg2XOCZr9EiLcGknKLYHTX
wTQrryOja0LhJfY6N6Ugtu/waJWDyCINbEdkpSolm0wuMhMwM1xdAILPjkiyXA7ixopjC8T3nuKV
wj0GGaDqjmtlnKgwEmdkrZwrXNlOqFQr8nRC9nFqjZURKpStF4ygylZxp5FTdhfxOHHC8FwzzWkW
W8IAbvz4eUjJM/xlcC81c+XPw7j4NpYb+c05Nx/AZx4A14zsj4V3vX6eVjF4p/PC9S+GYboqVv8l
lZfonPGiSpzvS+21lx8V9MeI8GZ76PdfJTxD/97XZnnQ3+U2XhfD/c2IL5FQWiQVo44xgIYIn165
vNjDQ4veIVCacvJCnJhNZPFjyaPLkYy6UtvVqN7RKgiftyfpl78QRr1tna64U1PGx00ExIVXHSNm
twP+qX/t9BUcq7Q104bjRNCtOPvmUbT6Iv18BgcAKOwbvTJoqfyi0GcyyHBLr3rf/7PgfsDvdaCN
jx5ySP5g1k+EwSIWrSFcOZ9UUlubZe2xpbguJqnUXYFdOdmwmwNK8TP604ZbskZu3dQ/cyvEr71M
syr47aQHzvHqoEV1oAb9VvW7eraU8VrHOtmyeGMS7IHn6YSUKTMlEGqpfqVV3kmAhnqyqRDASAth
me1yz94TkHfkxL+8sj2EPrF8p4NTexiZhfKaIoadIjIK2vfh0XRtV5yrmper3aYfO0gUwoYU9P7h
Qljtllx5w/Xx7YWCk04NdUHFfwKeU+F8t1AL3FtEmtXY0Dz6GTKy4tajShEiTP+977aXkfOma5TV
rh1OlLlJKnaVcivTtZ1Hfdng5RKXdr0/CwFPkKhU2gwuZddvauRi1Mbwd4rjqBK1uzlKtJ6WvMbq
civEtgVW6m6U60yYAQk5NkWlwGSCb/JYJ4GDrpDq333Fh+f7cmo6Tdxtfet7LtvbbA1Ccopozhj7
QZaaSXz3TUwb1XkApoxe+W+jSf+FYLaC39f1EP15Xtj69qjkP/iKik+q7tZ/5VszYtA8Z20P7CNe
4piGxSH7CbAvH68ASOqdPNrupss/xqYfkHJL7aUkR6umAj+zMZ070lbuDxGgpB64C+GmcRXwb+iT
5H8c62TxptU/P5PD9I49kHCOqHtpUzyK9MHvdR/Cwxpeu5cVdV1UTn2rRSf94pE1/3JutSsmcPHj
xhS8l8A4wTAg4HdgD24Qe5oAf9mR8/BTEMcOJ1IvS7Bx1YVT752l7+JYGuMA+DLYGaymDjVQGLM7
8haGEsyPV2GEHH95Ecbv/k+OdOre50+/9Ua7UDq9Fjd/qAs7TaRzRVfBlM+5gBO+Idth5BvQcF8M
Y1amSnJpPtDNxEvO9DvKIfMiBaW0D8DiuM/l1M4bXiFWf2gRCUc8nESK03wMnXThvvwUKsifNi/z
UVPhkWVAwLntPnkzWhIkgyoL4xW0CxEqph2EV8cgtOmurnMhCF/wx638U3eyuTPOOCuvuiz9mX3v
oknNKUemU/tukOr9Bopc5u5NRBjgNEO1P66qqIf/u46LtdgiYKYYfZwQO7ssTGWCfQk7KhCSzpGJ
Ws5tnAWVIDykoDi4eyuuucCmI8DfXVaDPKZjtzLhd5a35tFx59MVkq7yz6s0YFyYrnnCkb4fchAS
e2ded4HfgxAVCiNHeHr3wDAycZnYX7k09lmhZIOYyoCT+KqilYY6UanidtWA2WAEFKI3uxocIne/
BoJeKuJJF5GIJ/mmoherVFDFpDj8qOG9XosWKE0t1VCumYK82L6QqafW4MwA0pXHtulJ/+TsXBB2
dXOumjtLtXtuzEMyJPVsr9fhmeyI2pAJ2sIGHHYlrgiVhgzHHnkHq6vuBjH6tbYPrXb985UfQyT5
1Fev3MuJvZcTKRb9x63ethVmuFlt4/Nsfld3d+G6H+GfsVbrmDkWYTY3ppNO6oPVgBWXfMOlP5Ck
19JWf34CvpEQ2ntjRDJKhhHFgA2QwVNPQLWA+3Cfu/pjrTSoB1sv5S7HcFesayDPrsLRStHPDc2c
aC0VGQ6CABUzYGhOUM5GQnvSYesiqDsPOItmQtcl4+uY5lI52SzS04oZhmkJmsNOtkuM/v5AACsi
9D5Jyk16TBK76bSxa/bv7OFGt//DE2oh4lTOmFAXT6jiL8mqrHJSkLLZugktIL6sUzTzAG0A5YZw
Wb/074BobEjCfQCE3Rh1ECLwVeJTGPRNXGLFz7QQHCAP0u82ERSx8yChYZNV1WRQ4UlstqqJm4jB
t+FWFcoBDXI7kHG7h1I5VNUadrkTN6feYICi+sPHbo6p9Vtu2yypJvkDj8CBqtmFIJC7E8hdDO3+
mrjW3l8GNkSDAy/KAcNe2g9ODoB9/ugpdKJV7afGg1krHwxg8wevLbnS/aKgLSnM+CNOg3EE2416
pg5k8nli9q9FQvoMPNKEnk/gfVqJCiCQiPRClUNggSu1lotzhLBEk5JamDWmN1cUnTFJPCxI9tZy
onLtNWYVgCKz8cWdq2p8hKC/4inigDp+/SLUKlZCFin2G8km5Gp+2ssRm+j70kcdc/e58ZlUqKlx
F3Wpo5Vw80y01zRozhbhsdpDfGPzcdL8gIqUtoBNwf0Yau9Cn1guCEDwnpaqp3ai15DMpaW6uaGr
WQ2IdRK3FzMg3659CrL8LBfTQDbruB+ZgjifIiEE4HnflL8kBNfFUeZZNS8aipq0OFa2CiY6+b7Y
yhv3mCOzevrcY5E6j54nzOoiSkRxwPTdhAcHegs5ZhGXY7yn9rGw7CtrMJt6X6v1fSEIaL4ADvH1
WxI7KbUfYb8Tg8kMXcqNEVpzEFwxk64sQvI64oEpeg2RxkMiEakHTiytzfj2eU2WJ8K+LtuT/dQ9
ANxi5jSkZ2MPtpCjG6FevvaulpTxrPwKqmAm0+2fn4x353awcNdd/HR+Kh97SALCB4xprvBxpkIv
KysTp3XgGu69zoku8Kah/nizIDqKDkYKfSCXZVCuOJ8TL53eBtuaBVXrqDUUsexWUNtytoXJe44z
oVoNJbPSzeSx+rO7yqguzTW7JEqh9kmE7wqTn91Mq14zao8hxOzK4/nCU5jXvVkspebA3OnDtEK8
wwnU1WLZXAFC2+N9LGN9+Eg3CNoTx3PycH9IL3ddp3HGvtXo1qgZtpbt0Nue3/3x3fzh80LnTB5e
HMG/sxIVLSzoWRO2HbWnPj2/+ns07T67EF6ejFo+jJyT4y2Kf+u4Lwny3xpixP7e7X/iILRQRL/f
2erJlhanmBzoFq/LohMHIaQFAX1pY0v6R86qMbvPjiybsya9cX0bDjEu88n31i4NEs1ruSvtIKOj
g3S2mOPuq5L/w9XgHSD94iIYObYrvycztWz1IV60k1B1J4tBw39Lryip0qoI3njEn5rojLso7XIU
7wf/0q8m/AzTc2rUn5yIxxDBulwTwNjTjKIeGEbLIWA2rTnOxO2NouUsOEtFDgMqyiKrlJoRcJOs
1Fa3HqGl+3gPbQ+MVqTkFK24OcVzT4FKYOJYbdgNC4OUaSHuA2zbTw6GIkN+bUm4N4HJWoScB/Jq
yw+ZcIf3q8siX7oxVDSDLkbwmoDSvx+G2hNQjknMYNHKlisOI+Dx/0uS7LCMWIp0Ed6MtIp6XN7n
U78xQ8w7mnnmRQvHBUfiolOktBKsvtLKzZHpg5NqnJ75Q2vYRfVU9ce03BduaWdFZGAFLYVs6r0q
4oIykUo8fgCFI3exJRfGgn31l5JDyKpai/whPi6R7N1K7Bv5pYNtNNbev4f4Eizopq6MKJetRofo
1cOUTC+MYnqcZWYOUhXY9Tud/x/rhRfOMbJeBypez+gwxgjVXAIsVsTuLTE+MSIFvR4NcjHoqiHC
LAZ+wKDjqYcQu3yYf3zBKYg6B2wh9On55MZ3PtBL9VjUtsRtbvOFdZMHYtJ0r7iKVodrtICDq/Mj
reFvC8+Rp9QEC2mdtcqwGFZn0wTzZZ4QXzEMsA7xfp7BkGP3Wx9DpLgteQVNL0DxUXH0J33/gq0o
NXnSGvCMiPK9k9ZJRoWtCJvmqjZtO1T0UQhko1mwaGtxB9PUbki11ImzNHbPbkV1w1EIq2J54fr9
9cnTiL7zh6O2+ZTNdpknmutwNYi/3tky0i0tsS2UaiaE7A8XHH7Drj94b6RUPmHVztxbe/ZKbjyT
HnAigzG0OiyRBFoGVnLh5Sltao0oXBJyFT4iyQVhRA7lHK0R8TWOd+D8glLbTjtDHMKgg43ZJFYI
m9nD8fEFuUuZPveTljTyUGTY5LbGw4T+TpVlQZ9aluoAzSJxj1TvVs1G295CUx3QQ+UfZtoOn0Gt
5KdLYI9WyEgvik3LBa6d64yPFpW6mXXWDPRs7dn82Cu0DWUIXrN0LA8vA8O7nOT+XtPsJ/DkAcHB
gn4XGEiGkeFLkEEr9C6dy97jC/jNeUUc9hFUZfDtMBDMGfQQiOmKCYJYhQkOA3POpHs1UMKsuHwL
ppI7jeS4U+OyRkDlWHdLj8Ezds0TxyhwIiT4lN9Ioed5PrKO+AAX16EXW6sisvCe8QH0UHtxZTs2
a/LCbHSPBFpx8LfYZ0hc+RpvGlVROX9C+u5rmMiwPjKS5fO3GY5F9oN4t2JxM13VMk/vQjdQQgLS
MyRPPusOAq3tifXRweZyUyd4TvwilPGj8oEHzYgJMITy81jZcTc/Rl5bH6Gt2esrtg+fOBmGztPc
zO6CXgWkR9IFa8kl0Bfq7dejI+vO/AqMPohmbmO3KXv1RcP8knY3CBnOm5n2iA8ZsQJQwdOO+oo6
dTxcKT7tqREWNXkHlssAvgGtRLEKLSjIMlHFu+pSZI45z8IlhDpqwEBohuHYN3LBuVJkUwfCUwNy
oO1N0Kyv9M6xVths4L/fNmDQmUbbK1xBQH0oVd5pIlVBbHP8auor5tl3Hry2DiYE281uV3j2s7OL
ip6FLX6/UW3TXpAEqETjTchsdJ9zThEUmPZk8rAxRcUKKu6mj7qz7MljWSBoE+Msf456kme9bCCu
wyqV+rkdnpkA6NNXPQQkqm89DaUI7xeqN66n7SeNNF9NFWnsTTqLwTEyjHhbvG/Gy662dL7qZ8nR
R8YR0NIff81KMTDr0jt0zSN0xEtjAVnAQThywDvO47IFZULAtrQ/EMewRuU1Chzrf41TYckAc5/B
7cQOoBRn3bfE2DNrsJRiXtGE1hGhAO9RdMgRvM0v+P4JnvcJRmoH5iAgFGI29mfz19VTHVTT488H
Kh6tQpb0cK+sFSPDe8pjuAESqD/3x/FNLAv/Ai4FybhP+cn2sgB2pVeH9t/c+7n7VTHqHID/ReFS
pCLD3HOq79c3aul0IAC0fD/O3Vq6Lvk6xo74T9jsDXcT2A2FQzrpXeAJT9XKNLyqXmjD10imC7Dr
Z/vfv5RGUlNRq+HVq3SFlHoEiUgUuSIkPNbXVnebiPP7tfLWRlI0af1gKyiu21ROj/cDYlH5+XiW
Zt7bgsA1iGUABR/sNKSLDC8KrDnph2YlwpcvUw6x+A9idJ4gE0YCY/B3IoNPyktQJu983YRHLaTX
NeG70p7IwmC40OYNuVJOXpYf/iEFzyRJ4AI0dAoiFZ4ZsRRlrqxew+/EV1C5LM47AFM79ylDxTBP
GunJxmWKP+e9sQs2GJTqRPxvPsrIAoeGJgJ1TmPnwWk/srK7XheS6XdBNbGM3fd2alCqo6HlZeFJ
+1dbMlMb3NFEUqwqstcRYCKnbfMWudTi5JWXeOPalL9RqoUDF2MfND4/Avj6pmtjz7KhkZN20+9L
AutCRecEIdmJzXSiJLuYDLrEpsH34JLLlNYfF3+7IlbNEib8s49+SFjJcUsSbacJJnhQZUHwvXfh
6ixEe2qIaMtQezCSNbNmen8ndMv3/x8xescN7u8XBrJDbkIEunoM2hYl4wlCnhQSsoXVazTxffL2
GO91Qe+sd/m6TjrQ2BEKS7n8euEaHeJG59n+JtFeVitfc1b56QSq3km+R7VTve83NBzrYQ2otal1
jI39mwzKBC2Rp+luebn0Ew7JkLxUAI8f4ea5fnxiZYK9kuzQn9Nk64AMwofWU/9jWCAD7KtKDC96
1j3uZS/rlx57zYUxAlDFCiUO4gBvwnhQI5Z7s6L56Ag9Ps815LjWhKRumcHM+qkB8/5NOoF7w8ty
GT156uncw+/lJVKTAxxekfuCaA31AfVROW5E8OsDWQK4OA25Wppsml6McTFpFJqjypUpQohJfRul
0K312z5BasEj7Bi+4ydTUFzPcKGlXxzMCWSFE3Ds/k7uxVEZddv2akZE38Wyx+d80GzrlVUFq7Nh
m0/At9RftsLZXDN9MTFJUhhwg4JYfP6GThGObl33Nuz2mNYniOdNgvjCsNExSLSyuLb8eNXEF0Zj
mWETyGnFBTWH0ZH0Ws98ANO5Vjn5zdkYxmWHyZe6C/jli8BJyBqEjBX4+ErJbDwoaiQsEFdtPgJ2
a7hGFNQZ+Ketagi0mEFk5XjbbB6HCsmNfzadqnwgUU/+ZoTAY4Bb2jM2fVDHfmyUmOM36mN0FAxI
C41cZJdBjC9IDXjMF1a2M+Bz1HQqsEIOkjF27JKXxCIMCqTHTFBO6tupaVhEWdd0yrmDcEJJMril
Do6se7+NBR8tP5tEzU42BiFC6qh6UNj1PgiPF130caDjpv9y5IROwShCnHvSbiwX+8FstQgVWoOH
e5SNKoEK9J5N1ZB8mgMZkr6jgMT6+/u+Y1Z/L1s+E2HfR/x4/xlGtK8dqrmAEC8vQzC77u/AiC84
8V4iy6dKuYBsCkLMJoR5NNVK/21QjFgtWl7HiwMZOnXlPU8RUVABwnT/EosNTHF/rXGq1vFLmSDF
cODX8MVBA3d9HEOjYpA1nOc6Xa2HU7HUpvGvLGYHMo6BmfD1WPM5/SGrJjg8QA6HXcQ1/iCqiWTl
zrGHN/E42FFmU50sLWhDE3Q90DXO/X/Ogkd0ge8Rns14XwCkYRicMJC0uYo+MbmpUhxyNe045w/z
l+aPb3sI9vQydmJFnK3SwdHbJJvys5iF5RRTAy9B2Yk0qlgcar50+ZRaIE+57qXEOcIn3H2PafZl
B+K95OLnUPRzHZlDtwla6z460/Rd3jwP9AkrKHqPGU0BSSYg294tAet6YvasY/u22y5gfcA4nowJ
X31bA5/kCvVQsMUoHt2g8fYtljhtGqwsyzbqPKvbIhy5/DFNNhSCo/3unlkQiZJZJ4EtSAkGN1BG
9NiySmQ4Ma8SKmbm39latPO1NrLc6bdU1PaWiYt2Ux05i00IwGD4fBDih+ScZ9tr++fKrPkfE7Mz
uVvZJ1hCnDd4biS8HpTWqVudMd9pZa9RGpo1cOiQ8gTdyE/+i6hn8mz5v0XURLQiLIi0cm3E3zLZ
AQZKw0ekTz1riRTZ6+bkxOSSDxviIkXBK/x3SkyDlc/50qY3v011GqJi21vs51f5VE8l+EXoMsrB
eI9pQnBGkQ081XqTx/ji3Wq3kpQrmpnCDKaPrv5Yil1kDddAyi4eoZgS9XC9Zzd6eVDO4ovS9oSE
0PMVIn5ntOuBvTzUNV0+3XPc1Usr2onUCcnG9Bf9I4WpSSbi8S4pBxbyymnV80ZBbfQxw+VeLDOn
jUT1Pex3un2t/zaHImZRM5HgpQvLsnmS8uunuxUbWhzvYhvIZrDX2DmVIl5EPWUR2Cr5+t6J8B1o
uF66GkugJDQJq7plUsm2ir61pc9z9EMzjImWlPXMW+Qu7FXhnfXJxl3s8QxbpMIyyzOxqAlFZo5F
1/doRw9CrHhnNcM9tmxRz4Pycf7YIMPVWTOqplhP41B/Y0sfYzUTPACf22S5ppX7tQXdeAGeXBg6
eXLaWLMtnWqM4TgaN10g5WMu+DDIzLKufecBOpVJGMPpCSE9uvU2l6hYN+YSVaZGSl8IJj6t3G6R
dbd37+iVDyKQa+ejxP4N1JzWjHEosdePCUya9s9SfHWc5aHxP6oWAmWVwGMUrOg4XOuHjQL1xnNU
LKrWNZdzf3a9tNkxn9d1fJNwXzHKTJPTTht4ahUoEg+xObI0XYlYhbXDzojnFcSd9QFR0di45QyN
upuq3A+Y99F7pt04xNsOH3b48j7PMUCwBr+ClMM4PByx/Sjw1FQZkPfRNrn4Kv9cp2USaYBFGoCg
r3mHKCImVXHzjiJwFUxh+SrwjVsomEMO8T8c5IALdzxjqRGXUju7HDIlA9QI8fUlxnyci9P+3x6z
rHfy6ahAwaoPog4G41/a8b4QDuc3DmNEUUzCMmHH6mFKmqZ5KSmWq7fRVNCB9Xydsu6K4JZOCsLi
6pGBN57k1m5hBFGcS9nwe8sOblN3H6dXIa73VLgczsf8OO0LqNRP66KY+w5eW14hVReyxsIpXrtR
fvWjJLgFgrn0hBr+5mkI4bC01ybP45gJcyUN2OpppsFBNh5HhoG5PVo65MRx7tGUz2MgUbJGyvti
WVt+fGwp+hQMJ4JfioaCpnyRBJz9WcIqu4lVDbYAqN0uWWAqO6Dp55m3tSrC8ywKSwonPLoBRysS
BJf7yIXj49nfLJVgwvTn9dkHL8z70zsDP5FIneucitZL2X4tJmXIOuwq521Zpln+1kjCjhar0jHA
p1qPiWn0eSpFLMDvp14Kfqt2AJ9URHaYhC2ph+vxvB9Bs9UZnMVVjQfBwwwaodLoLUIEcJeSZimj
5pkCM//UInsOjcWKipic2QUcM/GRFTc6Nu/sGK5CfMUp+/WM8ScLJvqzOrEpptss6oc+AGEQlfr0
IP+5hUR0iEeAG2HMdjqYFEjLPu6oCl9Bp3W++5uTq8YJDyZRynlnPtrXzjetnl8dvuLWgyRPq8MS
RsweXHHSYXqfctu8KZTKtVFpY4aMokCY0AU4tzDwZSUln2NqP5sja9IyiWXYrv/MvwY2gz0PRoqa
M40XtbzgNuynmgXrfoMFEKjtTqGLDga2oJMa/IlYf1dzo1vHsWJt2AewKDjQRmFFd2ILQJ8ZtBpF
82aey1p5pjds7TQVELzfqZ5y6JGRLRuLCfOAppThKIXQ4teWdNqHq1/lqIqb/YxmjYW3h3GaFhW4
eiu+c6WzrOtAkUsrq2LS4QpCf28ONRDsCbm6MrWjtn7yF86PPvN7JhmLWrUceZQoR3UIN/1VVUll
mRSPHNO/GD3783Hy6Xw/TxapTCQFCwvZkmPxK+NsBddyh0F3aAYp/O0KGNFhixsnMoIbYp14QnbY
a99SsNqPF5O8AS0q+tRJ71Ruh+cQNB0VWcRuIDkLEje/8Eq5erk7a+1DsJBDAhPDaoBaa6xUrARZ
iDHhcZ7xYTJcQ+qLI8XVYapSe8rgToyfTcdmKycRdhV5ZmZC01u/igyXTvRJPbnl4PQPdfMzsEKz
yZGx4kF9Ga91aYJFVGTbVnvCNASeWMFBXSU69hVYso4R6WrlSAJt2iAzclyb0FqPRagyjfd32TyF
i04AH6S2yEdAeBlVCIkNh0zJaQZUTFMD9tgkQFtnJMlZ6YG9uJaV/Sy2kjXH1F9OWPu5n9TfR8d1
siciuMemWJ62pjXLJcByNdxhLNvB0SvZTO0UDxWJV9hvcOQ8hSyQwRgTZAKKvONpXxnTUpQnTa+S
2ojt0QMoIb5jheTtl6WECxNmtfo6kduradJfMf6P+UYQPu65HhTfY/vkzAdUEroKF1JUcypA7Y3K
5rXG7oAkk73oCT0bPDislA7OXw+CiOYnyWslJHXIwEoWyO6Fs26lDbCxtQ0zzy2WOb2PcqbysCrG
Hd/Us6nbKAYu+yMynTDiGhgJlRlt/RckbRF46QN/dy0df10T69VT2lMirbpOpeATyBplpawUR2yw
IEPbxdVWxZNbkQ6P2HcoLLGGJTZJbT6KG8vGFEm3eKTOqiBsXGRc+2y9vyO6AvO+eOjGRruu6gqs
4LRrhfTBbQGdO49sqC/PBe0OXJdZ1/cVwzecR3X8AB+l0oGbOTMVEfOKZouVvjJw+NRhQlKMLZ/t
09i5K0cI+XjwJLHNSjaaz/+ivM3QygZYPECimTb6jIT5eKQ7JZ6+LPJq61uLchbN1TwsTTNCpFBi
y9gwArJGT1X2VrXJywzjqY9p04/s/BfDYDdwvAuj30rioB/keXaM9m+4HQS3vhV2ZbtkctOf3FZc
lRCtUaT+9JTGylTaS5PPTTu4x41ZCva3kd9Q41aNO9wOk2aQU7HyNjiK4MqnI04h+KItvJS55zGT
/0hF7s7szZBi500lchESmvg0wF71gG3NlEAVnp7ZRp4E6lE5PZB523FjTOxHXAfHwBdn54GHqckL
akDxARiqUkhZzeqa7p+y7SuRYJdLllf1/5oiL5qL9mgcVRv7dvplQrUpz0gzcnSon3JcEx/pgmO7
ZXV8xAK28rAwflMZv1j2yVnj9EsSCHqeWdxQ33ggfFgrjlcZZSP1kMxR0LLw7N+tlyKPO3ZS4T2v
IfL52xuPdrEa4s3snLwtp9qsWiZ2pCUx63vd8zfB26lvZ6B/4bmoJy3kTKFCZzqeFHeiwVAYudbg
EwEoaQImFgihMM7z/b2IAa6QRiAA6kbiC154WfxbbLwW92IejYcvH5caGZD+BbiX5Is7DbOMGd2X
m7BqNk8FbvFj2z1hw7l60LWmHSh7vzscMtG6hdmpWrlZO6inr1NbAUXoSo0iszrEIzcNKZGL2Xqb
xqpsC371zIhYLT2Sn67erLgU3CPClBtb4v7PUaIqap47A1aG+VS/pAeP2J3Fnr+i9wrtL3X3GfWD
hXI5eU2UHFMvXQR0PCZT0joBoXamZXONhXgJOcDTun9kIPKYeO/XYwTXhDYppnFzknGG0Au5aO06
368IhA0ABay6qLPotzauj5lLpFNB8UuP1q8SiltIdxOB0+2EO8g2IB8DsmL7vP/VG2npvveyQmpS
PW6oQfbeOAyNY7lU7ljk/3jOYl0StEcHOIF/WAbY+gFRxn8q+Ca5NYughBGCMR0UhZIL37EmR640
X8zZRL/W03QxOAq7msA1Maey9W3ZD9dxop4n7qcUPtX+jF3xKT73XABlK7kOGKRJ+GOxPtg13aKX
yxNcVG5ZjD01JhRd8Nz6bl9y9nMJrtxSU23Gk8Z1tj244ZOT3a9mtVokLUwvHPSyaIzatvMlknJO
442nEAuKN+AvQYI0rIEHwmusYOCJG0tFI0oyzv3D0A8Ql+pJ3DfBAoN8FUbGdtzVkZ2TcQiqM6jh
nIAh6c5NmgAA1IqssrgUf1cpDlfbrXw6jYaNtmZuw57T2pUW217KvW2Us3+2jKFqsSWPeQecFSkc
I8XCDfFIqOLyiMme2p0lJY5SWJPxUlKYcoMLPCpp6j5w57DZ+w0tXASfn9StdOeOy4T2wgsozh6r
9fKRQ8/J6ucxgZXUo9pjjcrOoqhPCq67zJsztZl8COPnlxeGDIKiOAZtnXMstMrPJjDdQ8aAznZL
VgJZo/yEjtoCXaEVeoeqEhHVsTjE+Tz1GOqDPbsRObEswPW/cNxqejKfk4hsqEuyllJ4ZRxdX0ds
8iO84OsnCCs5ifwLqcrdryi8NIAVbwLSgnEtRL+BurV/YDaUH7qEUHSECmjS5bFNe4uT6ucaOlBH
+YJVeXUF6GGdaoWZubzNLoTUfyV6M2geIBM+KavblhdAheO8b3D/xZsptDX/ibt/hTNtfAkA0G7q
ge3oIzTLFp40xYKBZ1hRoLVmTGh1RXel8MoXSeKWvSVsqAv2AM6DfeqBSaFHT/CUiiEOndGXfYRh
xx8c3vTn4EDT4KgS4Ie4TqRkovdYtrIm/EBHrUzsDaISNoDVvQEUHe8mYQVuHOpVb1JLZdAGNIod
XYJBaUfSyK8bOrOHUfoSzZ12STJ1+rh1LGk1I4E+W8dJsy/awHciTAn96wmWGj515hNQCAPEChdO
FYR3tLHzL95HjqK32B75DpiNKzIjmQY4kkmY9sTLkFH7m8D7Ro2ZDvIWG7xjb/T6RuqEDcESip8S
GGyedTOs/BQtomXwPyfeh129wT6CkAbTvM9iwj2LXL9ndVam2hy0egZ9ibF5NeF9RSKWw9xavEEp
4AFSMkxd1wGfFlSM7ReoDsIfV3esQX7Bur0xb3MUFtkwXVbY5GfQn1HpM1fS33U/YIehsQP4x9C0
YCal2MQunRwnBqo0PoZ1okx2z6DpiqQT5k5+t5Wpo+nOI3la1OsZTXneLOxvqAjAZmwy37mVRM1d
Ydr+o1KheFOCaJeXgxPhg6vVMa2rZnOll1qTjIAqYS0T2ZVat6Q1JYokzqL8aWj8mA14qvYXoLF6
xyDIuVEWykBswCJyC6Bv50VrTdXK9bM/w5WxOhJYlSQA2fdD0EZBDQUtXjMIigYBXqDukG/NW8Gx
A5fCfzoiRZYJsYB8ce55HDfaNDiE9KSlHtGPn8wMhqtpv1Fi6SUGqIykVGm+cohqYFPYxldN8VLl
kWLAmtARYXMuTbHWHpL4Lw6MjjrrtgFcKjzyim+j/ziog7gZvRUC9/QePNFJ5mgHqvCXYuFlw4VA
LK8X9MC6qGRfW+djkWhkThEud8i7lceLBAsK34ulXz2v/xAzdCd2i+6bu953ZkLK6TTrgdeR1wFX
KkXnZKyvR6VLxRFuiJ5qPuoQm/L1ZXmPM+DZzu0t1F0n1LM/5ybdqZkB/VmXGKaaPnOSPb/imGSx
CzEF5hhz50dPYiOs/G4gdeVQNG0gbfVDwRgscNf7qKF8uMaqAiRITQVloFsqwKhG8L2OZ8Fb6fMt
p3UbHXmO66qtUhXSPbmP5KzQfHzu2aT7lbjE/zLDaUvSmrBQAGJsIxBJsJe43r55mU4CVGf6hSgm
UjuLOT7jlnwhwGTlHTlmBhP57RHnhDeT0i1fzZ1Odo4IepaGcOMzSYBiidwoaRGGWxhoAf8hWv0V
Bsjl4D1vMPCM7bBZofTOMUofR1bVNtHefai2xckCHGFHUt0RWhVAWadyA7OKTBFMIDRAyEhHatWP
e0zWzTvwac7rWLg/N+lWphJ+JJblVNUahD/1T+RsIDtFjhXV/qPMViA/MLNl+BLmgOdbSpG7Mrdb
5Z0uTf0bFYtO6EzsE1hdLozs4IVaMETv4RvVMeDCgT8ikhnjs0FfT5VoeXMcVyfz/YWxHYGisaFH
TcI770JN5+HVdyENxkPvnHgE3wF8RzIPFba8qKJzbqDbed1faFrRZN2KIgM216bteSoYfjo9Urtl
bDHkZRX2qkt/GDDXlXyWdaFR/ttM19H/rxin/Mh21NcoQbvcrXjO6xckMSE/mCsYCwnIAwJBuY6t
Rr96vrzH10jvUyujSU3o4tq0MJeEVMKxAhuyU/odUAX1tMqlOJ3dpEN9RsHOPi52agDhYRn6ssye
5Uo0CA6/BSUHxQ187UT3jc5AePZgz/m6uZEBI42kemm9WewC6kOMB4EKUxEJvNcn4NIm77npAZhi
jldoVVJtzXRregHNCLrdMfIgOSxyi8f6jk207jOVDgPnERSYJkm2fn4sVbd4Hbxuedin8Ygfm8/z
S+zY6xxA3RWEKKx+1un2GsJkpTs5mRllNFdWb7HB0OQt9WSMc2KcF6sJsWak1At8i/m1VhpRElK8
tAWqPiwqmN0UbYm+3jcd8lZitirp0AUYh33dnuIlXzjED+sPqsj3o1iDkzm0pKfRtiYrTjpAQhVe
q5tEncjLYlxDs2w6mTZFfZN1Z/q2Md7qtYUwrvsVcQqkNrwEvIXJ1VJbIdx/+q0TAY4m82yMa1SE
6kMTFYCqDO6PsIwKt5IC+tDeDkrMh7vYmtEqGFwiFbH5XPZ9RBIofqx5t7R4P4ulz99JiKHBvC0a
6PoHRmvd+to6JhaEKklHbnwGJSjhAkZmTv+Ykvi51ElwymDn7LahBxvljtKpelJXRr+pmMe+Ud25
5Vj8ZuXw4Mq7+PhBnYZjPmgunYeJ3p6jlfNQqyIOuBnyFyfm0ZLOBNFoYA8z7WPlR+ujxLGOy+EV
MfF6iALN9dtRgyy3tet1p0sKbBQvjmOwhUvktfndhorZIT/rXMEHL4RpLTpnAJGuMx1xXshjhhDU
qBXR4TTjBcDdC1NqSGKIkUIvofePk4WvZPdafXZ5L+1dHdpQ+Uvw/K0pO92pO4eWIJPRduMBgdkW
Lvi+Bufy7uZnwvC8v8uGX5XSpk1/DHDjhnyz5DX+pjUKkB7sC7IVgbG2UmT+Ka9y+TcRtKsFyrgY
kRRc4jfcQkZ90zVdi7lyMNNDCF0yOSeeRqC+UPQDrOI5bYR3evhHILIr/jEa45rzWXzVpZZZ8Rxm
12hFlrpHEk4bfughpNXnNokwCmeFC0NNCXlemcJhX+LX+dAiRfgEm8S4RoJJb7dCWgxJRjaps+Nb
P4lMXv1CSSM2UaxzxQZkOpc7/dN4vzmNtStAtXzeZpf1Nlft1CoI4vKdHnH517CHaa1bsaQX+xzY
VNSEuiSitRxESItJrjp9sjhRRZsTeRG186ZYoxO8QMCNpuKJcKjZhOVS5PoQIHQe7xJ322mrqUW3
BT4klFUHO9q2SyeGKSK+9rA+FomCreMEX7x/MUU/aoP0kDpVQYsZIf6uPcg30e0MJU1RkW30o9+B
w0PbFoSIMljHgenR4MeB/mlqJP3R+l1AE9t0XarnQFPFLlmKSUB5vVO9mVBbnhP1ANVAEssBAWcw
ZV5BzZyrt/8H/x4ZjB3f3kAia0DBNFIFFde1PFVjjKtxXjLM7H+H4BQ4657ppbW1zb37xoKi+KNu
UTw/RvkWxNvdfL6MiLaLkj+u2KnI+85yrxCo18olswmAWEAVu+dTHDQXpOAEuPg6ZUM5sO1ZVTXX
90PPmgM5wG0XxeU8dpXvvLNTLR8AA29x2hsP3YVgiPSfWbAHtL4mb6XR30oqiBdM76MNKpVe1nuI
ZOcu8Gt5rlrXZM1nGcN4/xZ9zULic0XCDW5xrhYSQMipczVONjAo1owK8F9ersSLqaUtJxrWEgTa
y5cwLjV31TKop42InLc7ZLQ1W77PdG9ZPKF42OB/MABOG8iWGsWny4DonKaok/9q6eQgCf+k1sPD
io5E+3kMKyPMShSAajFTPyI4uVZZQGWFpKD/hhMrNRoDgkLMj6ShhMRZrMcSlorcS8YWs7avDVtx
jDDcByyuzD6ZpnID2z2uEu/ACizbeMVicQKwSBMs0+uwdvmPtPbiWhAS8LwnxBYfcFZ8b/GqV+3P
dRw/ruyTm8/yb62wlZRdoVLaNGA2NualmnefV7JJYEo6xLTdfkl/5zqiHM2otGN/C9zl4TVlYbCJ
L0pH7EUamV2U+2ColGE3PpaT7fpMO55Or57j6czRct8mmGaftwNt03GTqUg/Xtef7FlidytHQ6xf
s5AyWLJ2X/+i0sqTub6AHyodRmwEPTKgwiGEiHm0QBFMS15a5BYQ1i0dFAstuxHTnGjlJ5ZNPkJi
Y04Ouq/Z6vWT5X590jGD2nOzFL1yTqxzFbsPF2U9GZG8O+Tgk+6hbM3c3dTquNfdgaA+cfjzqUdD
8pRyIxc/XqBqfDWy1CQkBu+GRousQA9XTni1a5POl2pAIP3XmAd94dWcDGdARQT1RM4UfNTHWlJE
ExHNZVNshooVO6fShWaR5U6rwDq5BsyXGQpG0s5O/SePgR1mJdMZxpADpLnDFDjpuG34OswKAcQI
mv3e1GydXqDlM+JZuXRPsryQ/SJRCrMhO60xyU9UTTO1H2yvDJWxItVaKMpOguIscRlGk3ZRqYa1
bBPhAxFzHq7fVASSiumynoIO+XGkWJPywaVG3jJcOMr8exN6eckZsPQ/yQAC0aaxNJEfrOB3BNsd
L3tS1b69/ITm1ErJlBO8Kh8d7yd7CPTgP8lxCVC2ACrL3SfykkV0KsgXtix2Rm/XBP5woWgTjV34
kvCuZKL+XOipBuyM+NqLQcDlu2V2kWfR3y62HPF1AVVB66F6dBl/L4G2u3byUvUlDjGgCM+i9Xgp
dmgEq++EViO5FWuZFT62Wfkgh26zjF6DZSJQVJQrS7EipU30IixpEC55PBwrQPhEts+T21akDTvx
fkJI0yxj8JJsvxmNLp67dEfHpW1F1GVywgdNcK+NR3geVY002Mo/n2E+1tav4eK7n/9Myie7OmlX
6MfP7dWO477OP+F5ldAy8J6E6UVnNtyqpnOU+PqlR2czLkjkzTInmtimTUsSPBgevJ0Kag0UkR+m
2MPQCYoNff7YpkxDFMM7ac2Rio1/piuSE6kasWr08hKDN/EFUlNUGFN2tdjWSD3sL3OO8WCE6WKw
jKhPke9S+kYN3vMDV3X8nYKSt1OsBK+hnQSlIqDE4w8fVNnsX+NXwoAq+e59ebmJlg/riCyzD4v2
vC0jKJVRkVrcPmMJ01XE9HHBYn4AdL/OZHWKMKB1VXA9QtIWQPWMxh9aJfCglQmDmxC7zxj0r4hC
+dNPRuz2UjmWwTzbxy4P4O8AdMp+DqGNs+hANgZvb+hqzqP8P1Nm7z79SrfCvmvu+chLYdh9jbbq
gKk4diuaeFEfhSs2Ql14Pbgw1/dmdMHldJtOKWGHUrcBkE4EKDQyYFwD3Fdzgvhzk/BrPW1V/Moy
gFd41RoDTfgWXj2PnokzTj0xErm3o7DdlkeJm7W+HZbw+Jz82BcktFmQxXdHPxNDQ7nIIe0zhbt8
OktBwMJ3Fqb3Wn5RB50ZqRgq21gzWDjs/9bTgF7X19/MX67xkv7dUY0cs7h+N5eqvTce62pPeryJ
8nDqDnaO8X4OhbIP93sUpkgpEmh363f1jr6kwJO3od26sXGe9an7ZATKnuAt+K4SqwTSR3gnY5sm
FLDtm12ZYFBmXKvPEj5z/pX0EoJy138Ztuaa5leqrJED4CX6g8asf1t2Iot4MEcawNHgcoMYkx5f
Ctl6xCxSEPDtST0EcOxUinimXVDYMndAnhdEtPguwrM2eSiM4Fw66UK7hYvxnu8A9ir5NLHGZ9eX
ZUrPFvpyuJhRALFXQEEd7+JCmOnpSlv5MJxbMpGgm9FGZzrmKog8DiXe9Ar+OSF1d+wTOare/Saf
cMHxeg1ot+TsQvuhzOANLDFK8F0E9BP3tbL90aoZHYblbpI6T/q69CAZQQgWFTGR8df0S+Vsvcxk
WTUjgkPbfosR+44XZH8i+iSH2tnFXireYD+gNc7/5Cz0YPlqU8JqIbZw2QBZ6Kms/f/ivE7qfw1b
202qdx9hr5YerV802JIk3T5ZgZTxnCa0tYvRz4wFouaM0WRJeyH6P3Ojr+vBqJb8KXOZ1/znER/1
bEHIdtmjw2aXdboNs4F97YNfCalUZpoC9UM8s0hMjKndwM3CltdMSZVQM0+mvJmjnkenn0VLNBT6
mo6Ia9AnaUk8Qo3Hklr/ypflTdCy6K3K5hZEZpNSvL82nNi1z9sVFCJGFR+Nth2o3pK0wQx9bM1X
51qDRWXwmGRchHtZRhfNHpnqKZamFAJ4B2aUd4U6IZ/BLfJNZlZoLHf87T/RbvpXm50C0jxPghTB
8wFbNnQ3CO+QV9EDFLjZ1RlARqE63Ur9GXpkhKgHT6yBuHc4+xQirHeR7vvtIwOHAvVGoDHjJLq6
edLvjKr4c4dBttNvLqytv3PRaoT+W8XXIZoMgZgdTbLUJZGSXNBzJ5GUeLRdsCBxuwwdMRLZjmKm
PbH1A9sYP7auJbDIUGWu+wxcSjhJTZ1S0dF2oHALyRc8iuNiERUUtmAeiReUzR42Ro7D4ZnoZ+dD
8XhOKzDzyziSkITsafclf3KYO1Rr187ERHKI4ksEiDGp0qoIhDS/AVqwNCJb45D//F0kkMkXF27r
dqh4+dABAExLKAYVYKVfNVG6kvJshc3WYqklZ63z82Wtn+NCkLpv9b8heVpIGT7I+mZQqtKbD+sN
pOymnzMgC3+eR/0Y5wmZEcxP+OQ6SVljQxzIfGnq3J4KtBRQznolVd6x8rK6lt6PBJHPFAO+VsJW
Kku3OaA8RBtcP8Nok1Us8OQGc14K5ooq9oqGNFGmb/Q/prgdv34fZFy31iKdVg1NCqjvbs8/jzQV
S+ILNGb7Myhs/C4r0GspJWAH6QLl8JavWjCv/q8lImyKxZFauRakcFMq0qwbPt+F2mDPOTOkqMPn
tX7W/BisuXl4Fy3xW4JI7YAcRzS1pR/0VLVIC86Z/p8xTE1PbMXqegqEv/EPxVRYH/ywOH3Yg/lq
MoeX6ZDn9phqJeAlZZWN9q85Ae9/55D/Zzp9vioxZgnTofzU/HrW6yAe9vZoXoJxp6YvLmyvicdM
2F0WwGIQsflCxckayxecZ6DPyKnmbo5A4ufNPElsmRb6up0IW3h+7etz8vRNhyNx5kMBY6nuTDVs
JAP9RbmdS0ldQKN03adhdQEtvZ8zMjzpbw5EFwFCYhH8ujap4xpRXjdvNTSyUeLZXnyVFZJANTwx
0K7uHFIONzlVsfP840au8tt7EHziZr/iz3sAriaeLkte1u8URYWMPn2epOV1snOZod/9uol28grM
HGUSgZWux2Hj9VRwVGGzciXxQEdL7HszO61431Y/XAwrrgEa6elCXEokRsvkF2jA2wJblnxuiTvj
Jj15ftBo6W//ZGhO492M+xvLPDAJRsx1iPFEAEmmKmLajWCbAjsZHP2FE8JiBcQVzl0PZH7vLdHK
Ay/8h51u+os8tyXLeqRNV8VP3YukmoKGB3r5VeGXE7USht7EALIfmak2DN4imt3TE1x+Dk14VoAK
oCcin3bOSwsnrmjs3Uk7QwgRK/OdY9IJkYF+RS1/vu4lOOLWhK7BaoQM0XsS9ROVv/5h4a+qTrDo
lgKIUOLDYApJnPKpNW8sOTkTiyaybaTWZnRy+RBD3h/3IylPmsL24l6/dXogGvYcEyF8buROE29U
Ta1Bq9vfMQ+qezINwVP7nnubUk40DGrwJu7TxS/Kv3JtiUosSavcSinJ2JUuNCTvLF1/cadck2HZ
KoIzSc2ViUK+toMWPu6nd5rRRJFYAKjNrZcZL0KmywceIvN/13tHsGTpFnb2aRAyuqqbx2NC0Dyt
PRZ4NNx/xzvweGjAPIidtUXI/scNt8zAMZ8g6CWaaRsidUY5IWJaylqapovtRXHblPnIPfNbkLJ8
Uv5BNjgwcIB/sXE5fZEdrlGX5OI31QPwyZtwb3zpGJFcD1uKjNnyFmjHOZnBAB3S/zGvTVKI07Aw
BRhzsj7LHqu1vBGwaoG9wp3wOyHo9ztvW08oWi56s/quclUdaUknyaEazUrlT4+xIA4fTiTLokCb
de0lKc5mkgIGXSX2bqKIilcnGgjT1xaJpr/ElJ8QaVaOPJrgFFvaEZqn/IaTvNcA/MUedSg5/n1J
1+N5WZhTcGXdK4n6iIoS3XRVKKIVu0YHzSRQpp1mt01iNhSZfCYE402GqdiF6XzCKDwZSquhNmUo
gKLTrpfckRRhKocq4M3W9WDGA3ghsi0+W7s/eC0ibeHqn9NXZ2PR2P/nVBFhBmI0u47DWd5ce7Rr
1jWMBqJusyo8JT+2SYl5RouHw4SRKupNfRfCAu/Z3b9jFNRquXi0+KakKujZEmD8DYcivx2WO5g9
XsLwOQ0dKSpF9sX+L6XEAArS/ozfYnwVbf9rjt+zEGos2icsI1CfAQlZ2OSJ94u66shzFR6LPd6y
4YlHYuVe3yZm9jA3fqm36wJNzyFhb4Ef5OEwhkAi3X2fVjybgH03QHkB2tR5cIKhLqCUTkUmoIqE
Oo4WFTVwoHQEoMudxEsFh5pgGjYNTR1Hsx6uYCyCX/hlhsd12jl6TEK1nsGF1eFT67lYnj/pcuFs
XFEhoe2ARL8ubmtNXKEL/oOpbE5S/+3s9ZjyqwSMk4Niu+aV4QbTxVB7mD0o6jSydcI5UqeA4rkw
EVpNqWDPfLdzjlUBLdPiTUK0LJmcxlVCk5GBQBJ6kX9/XuYQcpRsx5eGV2K4iFfGBeBT24pF6wfH
sfLxBvYQzq50bO4o6cRLDReRYXMKCm4jfbw3tO9hTjQhJAO6gp0PBPZK3LmcV9EwbsoVbpPWj0ge
sz+Q73dbopzXcg4Ly/5G114H6rldt5aN4KWquZJYNotxnqVzgTV8IJnWSwPJYtQ0JTvMmbn53Xgz
f9+8oPQDRaYj2pwB1Q4YAceJjfwroqTG/DckBXiioLeX9coT4aAHaDRjbS0AZYatLHpcUJ6r6WKY
mECpvPdlrUwK0H1XlthZTIlo0nbYeMy1XHkZ9y7GrgGsp3vcki9HtuwUbppIgE6TNpSs34HrKNxJ
D3rP2RlozslckYoN+dkF10ZvuQypkZD1Ban0WopKR6lbc4bNQIi8KXZc80pGRCQ9bEPtA5vPJTWo
lk7ECY+Yq/2XaEeRdUxeRto6TnDrfByWPmmQansJnCTQZvO3SCCKDbaRN+Q2UgIRC0NYDyhGUvet
ZXnlKVtCMHtMXSJekk1+Z7gqTosYyi6Xwj59q/DPjbo/+YKqRQhncBPamES15uzP3dco2HTIB+R+
S1O5JZmsg+BEVCuLbH21Vf+/WJsoNL/nNaeXy46wv7ynzo/j/7lK9Xil2WAe4XhKdMZthoptFmJc
aSpFdfCVSEx2vH279pizPROFhFA75LP8UjoQhF1Ms5/eJCXio9bFw//kPk3LJo1h9upqvHSCuVTb
0w6ih6IJmySJ6WGnBj7/V9wuTtUhobO/99+WhEZMbkc0JSgMq/lDDmiw9GHckCrdHdbk8UVwQ8Qe
E77Tgu1HL4zZJrDQT6pPs93/woMejbjv5O21nriEfjvUoQGUH/dpPQUY/jpBGp59P/nRO+QlGjjw
UTM3H4p4JHiDEJOJcKB3D8r6YeuEpXFo2wfzU84FBDVqw7o351DWO6K0F+JCa20u7w376RdguYjH
FDcDUmdGV2TH1PK/O17NHXxTC9EyzsTH/VLVdKBc/3m/MMySmFZ0I80H6OYT6fw8pc9NuzhoUjmc
QjFMzJXPA3X0a/OQRVXuONdGMxzzrYdF/EOmszeeolt2hiE/AGRYWgTJbtQY+EiZ+Ab3aAVOqUSF
mzzWruZRf1xOPQ7bnm5iSN0mZoB21/ARChb4VKDCqv5OBbnJDZ7E1aU8Rmtjt3LABaqXoW6eJavC
tWpfyxb2AV2iIAqF4GNRaN8lNbbtIaQCl3JFlAri3YDzNlUzT2WzFvEVxyABSaj1iz/iZJD03sMR
kpykkPAsc3HadiA+qRsQajl134RJFt1roMLemZZQxn/W+hRJ2+GdW+J29WgB6vzLnviEpwSw9INX
EHwLzXlm7FS08C4GvDFBwwhGqtn+qotetPoGPKRLvrMWEHJM6DRu1W/WDMaMgcIGtVguG5Np1YeN
at9m3Yqx3AqsYpoiNVDz2jT1amlgVg8Ewyo6F7pcCz9KpB6FbIz1m/WdxpjgQstUnCvxLZswMXfa
9AJHgI1aYQw1KqlLb8BeUo7GdTUdui3jF3Vxi5AcmifgKEdqgQLOwIbDT2O4jBWEBJkpOCtMOvK8
ED3+7rffvp8+jNmrHjIFoPBVLkyoFcB92p8YBGDFqGceQAGSX5INmOcFL+dq3qYs5YRDVDWcyDLA
9A74S0BhxikkQh5BQJeWsoxPzRIiO3cC1YTzMDVi8yTW2iwPzgs0l8IFOWKbrXzzGzJyYeYMNOjf
CQikI4xcxIhx/XOCDcJ6jNvJ8JZuMvbGCSjMn9ZxKEHKCmLKKizI1ZH9MdjqhtCeJfsSCmWLdZLl
IXmrFhK4/X9Xx3fkfLSKdtVE4TIZbA/SO7Y/NknWELdcxi4+99yhY/6xHyXAxT7x6wwAP9SwDdaR
ieTcDY0MOONAzaDEvFwO1+KrS3ZVnSc6y5OA8lg0uuXcXTHyKY+/d9Y4S8EDsLzvl3vvFkQoWHTB
jA9j4SErFSB9BAZ0+4DeHgxkwREmQjHkbTXP2Zmh4tph25XmWqV+yWgmTzA0U21kCL/2WQWiRGdb
NgS8ib4xwXi+DWS2j7mCyd3LOTYQ8e59PtVpeoEw2ysiMcey/9KCM1HYPwqAu2qrINIzKZ8EiJfj
Z1dqKjJeaih0RvwPU7JqUauZTRFod9VS9ewGZPbA7LAntsekIihm/W5hhO0P3euaVIQ89Rcz4hOV
NBu7gFJac0YgYSQ2LTJwHQS003YMfIdgNnPzpvqtVU2HL7/va4phckUgBggwEOfTeT2f4cHzGm/D
Eckf+cWMSGx2yI8YvrBsGvL/Yhp9nb3C6vWv0UMf5QRzyXyLw0yglSb8IuI1CovkJlsW1aaS7vaR
mBIHitv1lGIJYboQa7QNTCaKqaAqUVnjIHCKnwikJ5Ifu+dZwOK4Q0/ROzwq3a0HNczejABdYWGW
kWa64UWuAsachbQi/oos/k5pF8e/wVfXNDG+TIG/0ZYkIKDbbwcb+VoS2DBPzyCLu+eb6Ee6EeCG
BnxAdgNLtJN+o06WEo+KKatRErLOlsCx4nxQQupgaZ0ryoF+lYTxkpbd/NDM1cNmfQ0IwBZ1qx3v
TSr7kemqn1YGv4MYp+Vv2gXSK4qJP/GHCvBuci6rkY7HhtUtZKvi9ks0lAw+JIEpdfWNu+AEMc4a
7UFbTSX6+00DvAzNIxIZvWYXHAzHRefanFY2vr25QLMW0hbVzjqil/liOMuZnQb3JXckIGnI0pWq
e54B2NDkPK8sqq7oumAUEZ5DlSpndRAwWYl60o/RAVY+ytsqBvD1VVJfoS1iX9aIvtveR2oGaVgR
t/kEuGexrJRHwD6sV6XBDJDAiFfTste0L8WXIRBJ7o9UfdaC7LVmYLhuykTaNJcFNZfrVroqnrMF
5c8WPytdxCatki4RJXJLFPZW16OOKFuuHgPys58sGDtLmANH5HhTrxWx/bdnuC414COtmRmLQ/cl
edRxFUltw2Q0iGeUd3yQSe8kCUAgXxPhA4hmyuxX0TfpAgWbUf9RiP++Qz4zkZwgDolPX8SHA9Ik
2FJQzu5uTrmVKskaAXaBbUVWZ3Egagi3n4isfbqIenqxvEPsSnuBXNvkvZ3XxWJKh4KMCV+0U+uQ
UXfhu9Rp7FURKbQnjVb92jOZb0Yr9LLevXRdAISL1U6LCpmLvtVaRFe3mWKm5Sy1jcBEaM2ZDMOA
nYKhmliD58akW3RZcmc1QWep5/uVLfPOh8nwZEVXEVJh4/SS1p/KgHO/ubI1P/jjva8TSCbQVvV9
l8pXZ7FCHIUDzQb4kJVIA2u5HGGSGdkezxS2/b6tPMKhqCzlFXklDGLmTfemfKPh/Jpy8+wRfbvw
/C12lJay79lK0W7tWrZUsUbTQTDWdifmwgcbkZlWaSteJPHnRG2X4SwipWaz6w90ESXIjZM1yvKP
bVHHyu7gujeM66OEFnYtvtchoPtOwBWHPr5Vs7NX+BS4O3XatnYLDFU8crNwFQZji9SaVcm+FztF
5SRw0rY1mcSiPUQG0D+bYwu6q8g3/h9wG3n2Nzf6MIqThiP0QWeVvpGuDoxWb+3rPtAOEIHKuTRd
7dIgHFa68NyNmIoEckfrnKASva2c0p0QVjUXqw0aReStnmQNnsY0AhdUIEPzX8GT8ARfNrQtBF0k
30ODnl3wRY7+i2lPURelndqCgk4Q8FFBcTM4heitKZ8Sgv4Br1V6kC5bKrh/uNkxwIaBOWGPjvde
kaXhj4HNzMQ/BFtywTB/kuXuAFnrdPQr8lxbqsXv5qFPF5hOQuO2GDQkWe8jhIToNdE3SmgV5wjt
TjxHpBAhitFo6of1O4No+vyNpLYS86pG9aOBRJAYa11MB8pnJZ4do/T0DU/N3H2K4FgrsI7Qw1d7
jnRjRuVclTPsP1q02B6EN/Vyg+JeYMEquvx2G6LWPVXJwOUG07BcKuUq+blNohKswTdLN95YcRFE
3BYlBUeoPzpk4IzeBTo8ULZZWNcNLblTD/MJzqJkEmKNxKdixmn60/Y+f7c1/J9tWEdYWToAV+Wv
WurTSWn2WbIwIY7/gQfoC1bhNJUtmr6sEtz0v7m/5ch2OnCTQnQT5IbzzN9WIymSSA1Q6w8lEotl
a4+bSAtbuWh0VPrCRBE3WFKxnJ+he+FFeGePjajAGOZCX/rgGgiF9ihmZtazqZmziHjmSQ2FbW0/
C0f7zwBCdZcNf0Q8oLVq44hiQSvYWyDHh6StWwVSHmmkGIGKI72iBaNjR7IYalAoXZLlbNvovKqz
eCRA8x6xfKZqjDgwdTQpS6z/skk6xTBxsm+GfrhUVihonrx/z0opdnIiBl6QDtYnVj6mceQhIKcy
1b6THltRsvIwhq0nhS/g+hyCWmyLp8sw6c/Y9+kvOG5Rr5fg1UmKI1Tq0JZrEPiFdmz++AxwlgIc
ojLCMm7NeVJ2zxPGjpxkQ6Es280GJJnoigQ8L6jDX7rqRiwTWzxWXjoxDCPl8E+VXfGiTxMMYLLE
135fBh5NH4fNHsoOiwwwtqrfB39ORcefCEYe3lPz2kkBl19Q7z673i3cflCgUMyGNJd3W/VjGGDG
bY0yh4dCE0b9miayFMtg9hNc4VVKkfieHLm6chp6l5gxY0pyIb19KMA8eUcmZB1kx8EgFGlo/+H3
HXO+n4dN4ibLJIgSdyZyTIAB5m6nTQWRmW9xrRmWnhpeEW2Ck2KZp68MIQ4RpnKAAsliO7BCPjsk
QhRngu7abJfli/uCTSu3CJ7hqCEcJhORlI9b2Sm2/rDTROc4PQqiIFO+guX5DGc/zVdFG04Pm0CH
5mact95PlvfU2FFk9Dt2hV0q3dlWuv58ihLKdHiVyqBSIfkk+YYZnzVKI0TZILXMI+n1LocTH6EJ
rv8N4dCVnsubu2pbVI44fgmcKOywy/mh89qAcz75HtKTYD9N5CprtqpBP7LfUHzjTCMupWFjWhX+
uKLGBtZvXEleTwXtViedQnQZs5ZOt8T5bitxzof8Bo0VAGBAJhldTEavYcmw2bLRPhFIG6aglG/1
ja59+YHmXSpDeE4wLcfWdh1J718KIU3lf8bWjP1d76rTKAx5NYeTu/7+30oA6qZi4rEr7qMxDLL0
9wOk6ZNFcVH9+g03xbhxBiqYto2ceAAbJZ0KuT9zLod6NFym0EdZ9g/hWtd4+7z/pXTqCcu7DwNr
ZT9vbJmGzK55hwW1vr/fTllfElsCcEXUduDIFeOQ6zidxXcChmibzb9jDev21lCOkNVX6Vw74KJD
NoOuTXMJe98jEVJJ4qZPc4udXuwuW0yCsg7A+MYcaT3Z9O/C6Eo9qvSn7heSdKLBMDJP2m5Q9/da
0Ychw0o28RiTMG2aAkRkRVlzVO2Qe6dLvZDqu3fr3P43Trl+LMEY+peOrxKK/P6xL8YB4B8QdmT/
B9aiZI2CZrfP0e4JFJS8127W9LFjFC2SxbswV93D+F7IUNONhjgBybl72AZ6a9dVy40T5gT1HWrC
FU8t2QVDpzTZjL3JeKfaaxqol9hdDgolQoGwJOWG7w03qSHpZPjn8hPMLz1rHnAdWWsUDTmjJwpq
RMR3GXJelkJqCJoQshFffeQ+E7GXNI3WrFt71ckslYlxW0SIugs4e3g9HJR24Hgcf8FZFpAd5odw
sKOKx9wgqeFZ07CNvjra0UuLrtYkbytbkaCIwWY70b/RyhLrOeI3f7uU/D7liFmvqndsr29KJJaC
qBmZo0mwd4Pbo1twLeOjvEZZHns34mipf4rPXytgtaOv9yKOprtu8HFDk9SVu/fXi0PHYZfB7iZn
mFi/b2Rn70YR2pFt8ywfptSAvyDaLx2MG2aDJuzAB7dm4HB8MEMTR8ngG6Ujfn1EvcAgDM0642Qf
Ww217osnoObJTi4y5bY/Vf6uH8iE/hi1g9C2xFINXBt9k7njKasUp06/CsUD1Bl7Eyzt2pojWfTa
MwHknQeZCFKmqQ0k50U1k2yDTXsDO/vEqF9Y5NqBRE6pqJ2FHLLvQCBoQm/jVEO0WYhKHN1A9hNK
z0EvxZGgh2UbCS3JEcYo5AzxjHWgN/b5sxtb9b0QxN0s2xpy5FPhz8+qXxFMU5bgQ12D55Nm+ESX
KqdCwJJ4FHC6yV5riaNayggr1twXr/2LWdFu+wDQtOYRciZHrKM6f69k5tdsPzwFcUfOXcZzaBeq
Ip4kllidheZgyzfe/8HaKPo41g0y02fz18DmTLoQ6BF7k9KwAjjm8/CS+5bAbiXF1IE+sFGrA9de
oziS1zqCo8QRu5yVxAY8O0NzAPG0sWy0Aok0ii/sQ/aRz5MP5FoMdApBwzszIBIi+Pze26+yf59S
RtsgHeZnGzBsEH1FKoCN+KpAEQmAKIeegec4AkIuiNI487NR1glZ9ExcVm+3DHZuGTjgq74XW3ru
LeKNPqmI2fDVI1s5MDt1sSDKY8icziv1y3u/EUJFbTJ7CoNIPK24zcNb95bjpozROWvwdanoiOEd
18IfBuV2OFA1yR0JcONzaG2csZsfDo0zCgGk8NJqsbKINUy+P1+lIcGrDP8SKtOSy2dAWGcBUYED
/RJ9O1tnPS2GPXL5dY0NgD299vj3AlqNkbH87T2c0eY3qtAm9UUgSC0mbEFuCi+Z3C9r/E4GIEaE
XeWJVaZ4KEEnn7gyUwuRk76X68IwJPdF+/URbrONs/u5CUiT4cFKbbJehuh+eusDU06WlchRkxZB
+67aBzxsPxG/YLVxsAH0dJ4nbBLD3CcIr0eXwy2ixCRJCgRSQU7GkMJLPVqb4yHdCSRCmuA2pLIy
3LrOHOqdZqRheKoWvgSA/+apnsKvNYkY6FdjLihDe70J5UD8g1KmihYXzG+4LGhsskaaU9D7MlWU
8Om1YMwj0wNeB7GnwBR270xlqJJhxDqoXCG3AO4qTG65sLDjdVikbBFq1u/S+LHkGRluE2qsXYjR
9d7bQT3NOYOelkGsvgNrBqXtsluYF31YkDG96Xu/9HlaMmqSp7TlhkF6CrXV43JhjFvjj0I/KYsx
Lo2ryvWVznyB4O3cWFpOTw7mpJQYIq9fDVT69tYuQIN/WAUNS3eAE3oG1rPdJnVLgBG4jUsR0c9b
CHZzL2xmfvLGI/n1EStf5mz+6t7TjB9ZJjD4lPqa+Us6PzikpLmYZZsXvF3CGriR6nekKaVCwJ5b
PS9S3lPJRBdiHjQj88yJmXhU3pAyxflaAbEP4mgmiBMsZ+p3BP7WYEiAb3fUP5u7zmN75PM5SnVB
8Liyxf0sYRrqUcc4Jvi3aVPyoM7rsXNgrUIBz9HO+jY/WlIbv0s7NRPW7pJP9dL+yVjFMkyYs97J
9ZGCvXmhX+zzGH2aOCY/5jFWsttKAamhOZJ4RkmYuyDPTZQHb56uJHuyQdY6LFt6YcaLMROD2EmY
2HWzHKuAB7ZJGaZMNUzAWlgtyQ6d+u6kLLR4An/6YxI7odvvmslJtV1R9uhjPNirr8KUdqa6Pon8
jAF/RTKEb/5bHIlP9cZKRnNZrguZtGr5AiDkQWTN4QCxT5OJ7fA2RjHXV8ZPkEG0ZVMB7Hdw/CRi
6+46OxO+i1cAMkICecFFj8hOeAYfv8V5lGu74WEbAJg2daqNjliiF6SA3dXINGAWV8YCSCWdPGDX
MgyR8Dl6O6x0MS6rJxOlTl43TaBYwraEZSV+QfHvcXPRSk08ClJW5yp60jvZLaXAQjQZ10x4r7Q5
XYLvaTmt1ValkV4ShJ8fGEKklqcc7jURzw8kg6LPVQs9EheRi6wcZ3NNfpevdS8G8XSGmaapJXU3
148wGHbgCokvnW/lu6q4BlOf6gykTZvzyBBPr7IW/vQ2aOE0lM/ORSVg5kMItmyTuOB/LDCLqHa0
HnTYT8ZadbH1nXq1iEWgrl3pvPS20quHx6Gd78HTMKl4xBuXPEpCqImR4ke5rmaT3R7pkhgzEJiv
1svJaGuphjiDkTDlUPnmdTTPLiKINFOE+0qz7LACwVnYEamfer71142kZQZj0sOeRkix5ShzxbEZ
rgWf5xzRy6bED94NPLwFTRdW10AI08CbZXd024VIOCXXECwJbntfCKfiSRCpl5MSIq0g7g8wjghJ
lVd08HBsohxNSK3fmldZWANsxUIQhBhhqKPqCTd+8lIsp7W0JFCGQLK6RGtLJ1pNvZu+wWXoNujf
kYpftGbn6xQWfk3d12DiSH0IJbkWUf9GnJb7NGorSGHhLahCHhZ4vZVz4j5C7i61oiDlut9W+N/G
hNzwaxNokaqv91hfpozvYNoxsjFSseXtDs8gh6+TXq6+VN25too1NJ63QH30hqT17JsUpzRkXsnY
x5i3wcbU7mvdzVtdXwgp80vzCkWwSMnUFPBTA678wMNfOLGg4CYF6GI6xXXci9Dit0+YL3ontfC4
vPWXcsXTdh3HwFSY1ez/R+R4Mbx++kGgrGUzKSxBZ4HlDtdntT5JjeEmySEuCfOrSqC3/liZSGcL
gmu6ha6sZ0F5ec34zHq9ipLZwoMAI2/HgXEa1BcN+i4c9Jsxn5YIkxxS8e4e/yRXkyqN4IcUrcxV
XN+K5QjSpryEryh51BNRSfmILTwc0sHTUVCIQlESuGllnIBpOn69mnpw+CCfEHEdn7aBuw/EkwcF
nyKrP0BLv7IApjIKKJPEzmmjbix5YXAxGnOKdB5wQiYgM8fb+j0WlL9QjvcoHGlhN6Z4ANLtaaN2
bmveRv2ErfMfnUO+a2r3a4bUNPRWtnM0iuXWTCljZ+jtwwYMdUw3lb3Shwho4ry6vTRufzvDb13Z
3NFEtYMT/XFoZzMfulP/2YYZnrfsTWojlmUQek6TLIOstb0rOO+KoZl7pU59EKkY+Ld6fAu5Ot87
3HJkDiCj10ESjfTpUs9sJg/2VPvlnLWbfdKR8Tn9v2g3ppRTFxLbWIDz9Zo5+9ZHB3je6C61/5R0
g+rZaFfAh77ml45pY+zVOORX9NifLaUNoKQ65Wxdxku49MMJpHxgsm9S+l7D9CUU/UihGa35LKqw
FhMXSXlihDJNbR8AI14QP62P1oiw55Wx4w3h2W93CsR+iCKowSjwhenZicKxFU/9Wv1lgeqRNY76
glcbOu5wC2zIHMvTtLUbeBR7FmWZJEdpLI37KODjRJtMcVpj8fsrUxImfYAQdXwBr4vQe9yNHeJO
PjjQeJwNIJ7qDFu/mu1EgW9p66xp0bVWW/Lc5djIkaVTkXF6I4kCUAMPMJvT715fRgcD3KPNlAkV
/4FdAecWSAl/O7QJ3WaXzUYjNWZrRrhRot1dOscnaE0knFxg1YViJy9NuGvGjUkOGICqLy1vl52G
uWYH1b+d7tVyKU/JewMqfU3ZaAjCvOHCkVxqTPyxL9T4bvWRaNbmZ/nvdHKdJCgRAnesA4ZIKL3Z
VQK2WK/wGcJIkD+sv6grhbBrutD9WUHzMRJNBD4FXFD6Nlee1Zm9Z3A5XgvASDcBrYvJY2nXETsM
cB4ADx3dHqJn7bN662OgyE11arBb3+m2nBxN0kDKFN8cKS4pROO/hN7Z55JzHnBApvpkn+uSvtx2
I4DGnLCce/rXzVvXLc5RZLFhwP42FnwJQq3Uvv6fxguUngBkrpNhEW3qBNL2bI5Dc39+M93xyDuv
LNKnoWyF/yEedREcuusiAgWJ/MMSQHFW17JDaC0yR/VEKFo0fOVulWfulBLRCt5iSEPUi9/AUmQJ
fxc0zOo0xR+QuOEV+gMOFCs6YBW2y5UfAqFP70GtfISC9okOsU2nSJEwqD5lnicQFZ+PBLf6ogFu
z2h2l1yCJWS8xqmRe7Fvbc1AAdnKkt9NCUPum3hxq4sDCB4OqUjwlYuklzQ3gnlqvWWTgUSWLj3l
s6obFBNxTRpJ4Dp9TnfVBytni5rzC3tkUnTdXxcMxhe4NghQ7cWzWyz9Szd4ai2lblPsxD97MVSc
fg9HmVl8NJQ0gO4+OhlUxvNFoLBzDy+zf5Gh5VjbntyY2EuESV0fTdlwHQFDlAPDcyJIqGTH6lEk
nAuRb2zp0lp2pWl620uc/58lY2v8Hp2exvuUNFggRDL8okbakiDcz4OAdSHrqAPD004aapVendsA
tq47TQaWdJPgAcoW3iDUs74BW+9XQqvSP9Rt71jyeFkEp7zAV6ZcyjYBO4Vp3N3LWwgcnWs+BoHX
ZMneD0RBEdRsuapc/OMRkPCTCtRsCdaIsyVM1V3gWYFbJDb8vA5Aj+Ti9Wro0OZrMPhwchnqbbRP
GupbLJGhlDmh0P6MnLpb8okHAZsZycZPpy42UJSvK/q0U90iNX2JDmZR+KhI3/Nv1iviIgbVPcqN
qetmADkthCLHxw5/GdmaTLu51YnCAZ0+VNauT+cW0Dn2RtuM8IV0XsvVFeDRhQucY1YTxZIhA1+z
XJ4CivXOX0ZEQaLW2TDqROHsblEYT3dT/cL53NnLXgw95bUIVulMC1XWsVDKzAepUMvHfPk3IVkt
9qfKbJcFCXkz+c7f9YkLucI5CLo31+MpnQpQ545vK2iQUj1W4Xw0qMuzJnUV2/OckogtgaXq/ESu
Pqrbi2MN5gu3Vt2Y7JZNEgBCrQeoDv0NrGOXdNj4C9Pjf2EDsGz9dq5+CeFTnMU5CLBuKO9Ab8rN
arKMbta8BsFfKfb7OTZIugro8CxXlBoJpsWXuB/ssZlGN+vmBLVfpSU2Ar+rGP0jbo3ROz5lEz5n
zZJuyJfUFHNYzw5nC8cKAYgTGIX9ULZvdXNCgOLnOoRiHrajZ6J7lmAibLrKHLvAKBfbmbop20a0
ZYwfsCp4RSzOT1ZRXjtCbJ7OumZnEqIadEuoUU1fcm/CFuvSyERdeHbYua/yUxl157jW1pyyfVeW
O9Dz7hrDOKlH4yq/xB7L2MuO3U7OOPZ8ZBr1CbwnjHAWa8BrOxYa6JB1Y5LlzFe1DlpsYzhA43Uv
XQGjx6GxjjemtF9eaU+fSbDLcAWYSeSTnn95l7U70mIfOH2P7Qz/uyZH94W4jQuMrEcppqRbcJUg
GeiR4EFDZredqhgczTCwcG03/1kEUg5Kpoqh7AFhsRaOJ6Q3kU8HHDI62DsBj9frpkEIN0kdgsn2
4Wq2FtBP9qdrJjK2+ttRUSTjTK59sDzXfowsINw/4zcj6iQFXIw+itpWR0oLhh948FBcgL6JURJs
DVn/ilFKm/mO6TD+fNzJmmocXn2MZEOHXhyzOhO7ku+aop33Db8mpFnByRnK6Yh9ZTUzWIVlOEP8
hR0DBAXw3qYXRBMYGbZUWhvW2xfpGM5DJ/eu+C9FoVrFxt1EC3KfpyxgMki5O+xUG0IypWlb5smg
7DFr4wo1AiiCWuHQQLr1MHccuDA1HKM+r3ea1jBOBSBIH9YFKmqzRJMt60E5VQgv1cHto1hnEjD2
LDGew3IqJK5yoXG6WRLxkLnSb4J9NHJXxoaCtIk2t7XRTwxRVA5+uAkUDK010aZ9e+ENUaLZw8jy
NN3KIof1hnEAt2mVWJKzDmdnKEOIADnZR40BcQMot+MNNN38OxDtyhEAflqA0YjfqFIOI6xEJ5JC
zUVPSlOeSOHq8tnX7Xg3TV2zbz/003JP/9bDiW2YWHIrzvss0nT2MdoYNzCGruxy6Vm8lBMCM46K
jAzDjmVAmVMABaQVOH8MF2SrdJMVmREGuWF8itVNaowwoq34uJM6DfW4Ii2AbAS7nJAqdW92PPfk
6qgFdicwNPVhOsjgKzLn7LA9MuNN73/rlAr/tV1kUcldDx3BzOlrhU7tgBReSBoqM940fon3btY3
Kl3n2Qm6FGWu9BwawghPe70IUk5wjWdjW7sYdqN+3/8w7FCw3NFDq0WpFFP6Y1h1G8WDs9xdHl5A
7p7Sj6uvTNW74KaK15KQY9x3sJw5bS6G0zqRDyxgSgp6Ih+p4KtR+3LHRoZSSoIgV9A8RDV+2ieX
8cufSA93+XZzrdRw/Qa/FzT/mWrw3x0+atM9gZrje/cenHxHNH5dCS8MzFMAt+sdCSfMC0UXJf/g
aDkbnw8N50lMfDGzvqKvMs7JBJiFOqoixaqPtRwdq/5JAS6An5EtY0NDJD7OX8tRaW+ynTddTVRj
gzLT1CnCE/lU/lvD43wcOsYsrQNJ0wiIWu6WaqIZMvkmNV6U4jap5oeikz5ONMzBpXYS8yH86ccR
/yoJDYHWkMiu9B0giyRKUjDDXYKAdfjDpcCM2tfuP7ucd7vHVqHxiv8oH9DsYEToLyzBaJs8d573
jcd4tyYrAaC8CqG/mnoHrbHHQq5uCP8bmKczInBrN9OD5nLxK/kHbKrozC+14TtAsb6ZVwzdsRZn
zb7tMWFDYPviylTgf2SSiu/6/t1VOtQvTlSlNb38dWD9xroCBzvPZTLV+7gJBulOq9Uk1VqTKlVU
+pKve7CC6CQ5tzxf93b31uECd9jMr20vHHSH0dZDyTfOQajc1fMIAQi9MiYsTkXj58n3HMSpEt4e
ecTVmP96Of9HhG3vL5n0Yj6yCz8vzXFGBWD0BwLNfGy43bSCBz1wDwUfXfPE/zJQZYGz4H8DsAn7
Y7/C4YuaIQ7zUHOEqKHiBwpDgc1gPEG+YZ2E+s2xGYETnQazl3W2ogA6dE7G97+qgBwkEz/HZ9/Y
GsPqr+lI9CHsSi17Td+5zzQtFXgKvEJykoYHhK8kegl2ReQ/hE3+f5AQQt0QzXEVr0oYj4bgmbH6
eKrKQ2BvzbKaDGLAb3g8m1A0AmY7E8SyKM16TUMX5DzBLpVlkhZdO/bJfM/K/MaG942mlWewf51q
Sv6ai5LMuo5RSx5NPqi2CcwDznkUdwEkjJzpNpOUC1p/sUTNZleYvJWKC5rPOucxT1N1dpaMF9jS
JfC9+v1Msr3iSDN7YlC+hSg5juzd0u6SpaDHb6cueTTtZJwpXiKq/IBvK+ht5H8ZoQ7onrlSfqqM
zq12Ar3pOMLTekiPckin18WnPyQldjrmE5f3KGRbPmP32r3r+mEoOBxg4EbtJlCzL1YfHh9YPYBA
7InO2YSxSIGiX6KkbX+zUgyWS0/dAFZFPMc35ATD5+aH/Xfn3AcDG3bCWWqEibYZN0Nsr4HIaTR5
13wyuHGFC70TVkhZm0D2o1wonNOOeQot+9cyT/NQjE47MmuTWqz9WwXjrgCUseQP3TMCxQNxTc8H
fUo6FxMqgg7Zj0M2HfUnB4iSKOiEUgxt0c8BHq1LgAp2G7u0cPX/bnT5k7eWOyt0WEu2fRI2g387
ArCt5QoirZZVKGHEGWHMija28hfsxo75mdaRFz/r9/f5q3HEjAJSXfFbcl3EnvaN390A8XTXvMLb
1EHbdiqXyL808vC/Oh4YkZSafl28m/9oY0wJhf70Eh9RBgNfM6xuytBzmBr1t4hW6u3ZA5loGsAz
RKAAAWhKoWVSNQ7w853L3oHMFRoHxcO8Tyl9LbTpjqeoloomoV10CropXC0sUKtBDJeqLY4EkbDq
IRBEQVP9cnJcOipG2EgV4ZolPGJfJ4kDOHfqtPJ7hbdKswc/bxIMIKpTBc3F3VvqoSWoEaG79AXH
6fovJDA0gf/Q8IGqu9nV1FAm0C0GV4DJRG1AexyGR6cCOkbztpcG6TQg365q9ca+tcPl6WoH5JHt
PSNJwyP9z4TqfTB9Xxgzo5wxWWhDheDbSUX6FNsTfTBFBjcUfpCjMu9a0ycUK1pnZhzCkOmDMomF
x/vQJvQPJE7rb4T5tc0p5KmtySbygO3+oauaWfrr/0P4Zz/uPB06UMQuJD1GZ48aEgjpXkL6DGGK
+q3V/HzphsSS6i6K9Lw8Ccsz4TjdVAAyxtD4H4oN8KNlv9Mq50dPG2A4PHxgDKKX6fYWKpwPLfyH
eyNPjW1ptt1QMKcKMds5Q5TSj/c5pFnYgcKxk/zNuHCczNHiK4e3gm0IyKkhhZWPvpIwyi3tk/CZ
faXdfpiHjwrVKlZn+7kGmp20tEwr0HEVsR1uoBuluEOBEt2glymUto8GxXZnmaES2Q2V+/07yMkz
pGf4NILyLKA60dK2gu+6qvE4WkGIDnbr5KALBWDQ8ODqfHPOsJ5+NKZiSt2uYLy6R1ZjN4vQZ7oQ
GAA77cU7JOpany3D2tcxDGPcJ471A8md5hjtvBwjfIBDPIHhITQwzHtC4Ov4E4op5zn5lMn/zVO7
19xhhEJYqdgmWM1QyHTQNN7Eca2lITdfmFThnTT4vX0Y93sS8j+P0fjFvIPr5AgHL1Gb7PAsa+9a
OHN9T8DVl0StHKt7ZwPj+t22sjyiq7ZdfxVl24KCYZ1Z8cVdT1xIHFo94j3oZFJLh0J6VGZSdajw
5DqI8xM32gmjKi+TcaRojIHRt+qmcizhewsFxgYdfWy3NgOnDgWPQPXn8GkKS6Wd8lg31vgTxsYu
98USDvUMp7bMFeoO8/tUkD9ZXCn7XVVSG4Yv2yn5fn2kJXqSZgz5L+1C/AxOvnX0f3/txXFh8PPV
REl7B8qLY5CpsNo/R0T7QNfBtBIWWJsgLhhxzay0cVAsDVgX6zQ/Hv2dlJGXH38O3+hqPUiAEze2
UNRjIJgZqINETbS3ja6Zwj4sT6SKqs208NSL0FxcReY3FCmkd9DkekZblq0PwKKtM7j/9S/CoFIO
2nxS/IVriAlOrN/LB87m6FjyzmCZddqnJuVG6scRkZYVVe3R1FX0OUEY4R9KyjXEF8gfbJgqHhXY
6Rvgai+vmkm8nG6jfmUop2ddVem1EnlBPREZRqnDbV0ac13S1PpTcKgeNB4CYCGOvJkftryzyb4/
VM8XiRFEi5O9/fY59ZcPkDah9PKIAsm5IKCbBsSS6Ga+5iWLiU10gD5Bmj2e3WbQHc33Jh8UKJWq
nMUfJnqg7JHuCc/l/7T/+unICxcvwPWh64YUdOTEO5Z4UHDhpBtuyeuO3y653w9Q7DG3NAFEYy65
GyNGZOWm3CxWus28JqHiWY+1Vgxf9+9RCgaiMfk7hRRDyVfsy9kARCNAysuePTAHWbqf24csvRFn
9e4wY6LLe4pzCbZQbWrY+ohUQidfrMPld3tdVQ/gzF/SIms3AQssSsw8C3Un94GPSCPVNocgnslq
RKzR4+p3E92R5htLBo9LLawOVEzG1QUkccyr7uLclc+BbLu81/QEb7JWxzSp5hnq8Og+Oeh+IsJX
eWDXDT7k0TV2VzP08bn0Urvb5X82t9QKwDlcT1cRyEOATI0yVfPYq3WbUQxaxQ/o4ERqWWXpMYNq
Fv3rpX41VjO/Csujqu9qXgZ7uPTxcJijI8/LChh7CiMe5OUNNI/wNbX8NvpOcWNRjhvPQWSo4MQT
kBtD+Oqx0O87TrjzMqa1R3iTtrplJ3iiD8+Gz7+G5JUsm36PEa/G2UuJCwPQXhCQmRQVv8kQL5Cb
QfQj4Gt9ezpiQSTuArgPn5dZXzKdtO3Rdb1tfiEo2eBUuuGA+Kw/hpjfizdabzSA8maT9m8Uwee3
/mFDq1cOwEk1F2oPGEXrK8F3EX3Y5RAWHn6aunFC7BRdGHYY6CzDeHsRVEYNk4df560xayoQ4Q8m
1Wv7aTMYT1SlbdmjYTiqJqEyxcOloNi1/24UPaB97S5NXlVKhowBIu2vF0DqkVzDv1uhstUodpxv
Wk72C9Gov6MVXvKoAwHhBjhAbFAuBQrMioT93owX/QQnKDDZ6qBMMkeudwvgDbG+DytjGY7nPbWu
iZxI5gnbDNMMU7OzqeyzhSa+3yaGYnD+6L2azEYiCFs0opjGwhLiInf2UbpAYxnw5mcCs+KOQPUZ
U8utcbwBiHSrVCIHm/Bt9vqjQSZ0NOEywykehvY+jB/XlTurw/lvpodH2hnUt/ig87OIHznerh5K
XoH2+4+kwb8oKpn9k6QejVtodplD3VAnQBhUW2hgBIyVu/EnTzXQlBYlKMKJJyH22qsitnh4wvkj
6CS2yxvNkMBxfAumzSQWot9VEPeSKgb3Z1T6Gjdp9C3svtLhkwwi0j/gPBc7UnwBavttgtV7JtM7
Lh8rfH3sSuOK1vR8fgZnaA15hQBLZud5fzEdZd3JUyOqqv+sdUSOgLMlSV3f0axgkati0pmLE5pF
w4HUt58Guhl+h89dcB385BMMCJrq+XwaTNm7qCgNUZAw5hm1NyHSToqd+/Q0OjZisqYTcp1FKpeZ
Sf4r+zgYjlaHoA2oLqaSdZj1e9/MC3AS602OU31b2E/pLB9NhTejHeY13cPmDBx3j8Zk1Hydaiv8
WNv+10LDd3PcVLLpPaaWfBw3SLWviaBRSmevpONel7+3e5Q+/a8NR72KvAvmIGvEAZZNbMLLnMAt
iJ7KfwQRFvYVUbP7rc+8c+U6/g/razn8p6T8k/WO0Ut+VyWKGSL+J6KKbYQrqJGkyYy0FmbIEUQX
T9pMryRXWh6bju4rpNYmZ/+YLULWXl1kemxnyGL5DcbWsLvDVyiraik79da7/E8WciGkFsXOOmWB
jzozNdUZnZ1otsiH1LYJzqH4J9lSoXv17zy9S6p/baKZvP5VeARdCXFOi4MWAHy2OO8TGTpnnVN2
uXBb1ACLcamCF7SNqBVNo452E2oaiUCSCCrjYVE16eIzL9s2S5StYabXZqs5BlqTHBZn2CMhiJNV
wGhbeBNOByEq8hFB/EJrSljRDGhJAU2bV5FIcLS96MwVFILdNykm2cMLccjRM5qgVAhLJEkm/XDD
hShPRbi2KNjdIWik86goxaZcIotxqwxIBEENgNqS22cGc7oR4qxjhRKgs0xAqC8NG0vI2eqqR0Wj
bFXpBWq+1e3xH1NSPFgJjyoBGC8mYk4d2SYRONI/KFDhGIkmAuwSmM/Mz3xp7yKBGSyy5hjsoFu+
mRyeGLFUHKBVC+tZPZlOa00bL4ZOKFKzJraWM1i/3yocPz+qXBMLbOyZ1VOxFgOfaU1txS746dIU
TvYSdrikxWSfP8mkWFzoidHXXzk8Zibvg0zBD1QQbx2nARGJehJfYFbYnwctaWj7u2vkAJez+3c/
HW15a1BsSJ7FjYmAiIfLyhG1MkZSgqsHh8VOYCA1TGqxwauPeFQLDZrOK7RVwOHbGNddnTsRipUJ
tHZiFkMay9iUD7y+tcYQTNjO1nbq8D3FagRhBM0NB0Roqupbk64re7QdjdND8AYiljMaeya2+k3M
qi22/FGt6E6jx8YB066SgWR2pTlPCNz/ke8mnB9qePwesQDkr0/jQ12bQRNO5Mly1YLxfjXUNd3K
axmc5A5n2N9mC+J8GEmaUCbxOgpVvrrk4qt5Joxu5mQj33Fc+3Fyx9z2KqYpgnY4WRh4uWgkvl1f
3HpBmNWrpFSxffzk5IPok9LK4Fl2wlxTBJ3IV4T6Qi8HrBUqHIh5L7chDAGrKaXORvFsS5bV7StD
QT4N3/VHQ8jg7xzhVo7MvHgVvlaI+pcNoydqf9/f5M71oeN/Ub+z/spNSxMmkP7XDdSw0GqCazSX
nqf85n8P6R01HvYbu8FBCgtoB77hjaDAnMNkqh7RiAAfgzE5gjz9JuGX4ZwMHgZwFNrnrI6k91Hh
43HqK9o7pHWdFghVAILBs2buEbx/M7Pvhz9JG1Ba0EuawHk9/K5AvLmn3iLjnr54nUA1lvB+sL9e
gk4AgI/QS49F0hmAgRmLnRhaCWcjQ5Jr8Y+2KoHU2qrjOgtizOq+Ab3HnFDy5SQXrNrQT3VUIQtN
vCpbx30csgyE5IVUk0nUjjr+lOnIzQ1AwwopC3mjxJF5oP0CMZV1IeRSlbKANl5VVBIPJZiyKi0z
e62QqHa7PCM49TQO6eenNx9lpX23Asrs1R4zQKsc6VFXtUkxj3vJHwebRwFHEsLY9FTjBE/Nh8j7
7W+eW5XFJU0Zlzh9E30gHea039bHdBN9+3undjuUoszQiOuMUZeyRB3SLUEXS/xcXWd9f97Pglqq
v2u91I/H9CXp9jYvOhxLREFTOYM8QtvFHFb2XPGK5FiaNz7GaIqotdHyVQ40TimUacvlyb489QXa
sDj82+m0comNF9cA4HTfGzomX0scDaOjV1l7kGAE8OXTEoUrDJOO4enkiFVT6X+9+eamicszZ39V
LJkXnK6wehPEWXZVdMTkgamixJdqQc69r0iA0ZZIdz3RWPmMva3NBxpcAy/hjvhfu7vur44VRdbz
ABrgsQXsJQHgrKIix9PjAC2uat/O0zaElH3qu/cgCJcpE2G1tXcDkpm5j1nejxv4CB81W5KIiKEd
DfyizYew8a9NBjtyFQuWjlYLZfjaKRnzs6zxoMQguS/ulw7Hotj8ZtuyEZQvg2s/Un+Izc4ULpF4
uMMY0YvNNr8ZUPh3FOB4VSmfw8uSJfxb8jR0nfIpJyKoDkqgGSoYRCqgmPquUcNcJ6uZmIpUtqjd
Ey+Vy2MmGEbYVOrNQvPV4TDJURK421USoPR3xl5QDJQ1EInh3Fd3Rsk4WpfWEXrWMfbE/rqcdcCe
D2aB+Lg/qGpTsPzYU75FbshhNOhCuG4gSSJIDUuQy4YMraGGqO6GCyJRg+d2OiFRg0lCh9BI8C+S
qbhlKr0nZTtlmvd8qlBl0CrhB8+FfCadbP3NqN9PbG3E+rRFxK5uCyBzvbXjiu8S0u/u0DbgL/gI
j38UMgetZ3ElIteXeYknGCNzUbDw+uwqoxLj9D+cOZ9+81WGEgfslgPCLhFBTHZQdtkQGjmzUUV7
eAWdeMyriuhuWAie8d7h/GYmXnxk4P9J5xMgSdYKNYguKzE4DgtYJpmsGpaWHb9dvjfN00jL6aeo
gshF9bWrYBjKw2sYSYxqhku2UnfiRjDSW+EDa641ISOhUETOpB5wCFFEIBCPMdodesN88xTMJRYX
m6RFylWMYACaERg/X65VV0Ojp5oZ2LWddl38HaMHfKPYK70lvTnd4MrTzvzClC8FVxslWdrhdGv5
xv5582D4xRcuH2uiHWhBHkDBA78wIo22wG85RxI1I4xrTWAwxLBxd1L7KfnrAGBtHCSjaSAlQ7Ka
+hzruDZcN5mp1sxrdz38LzsaFoKsWHGe0FUT5lemtCd74YvVBYLFWK9CKiit96sH8Lw7SEgFRJIn
rYrQCAAXt+du3/Wz3DnObneP4YlygaaiJTs8l2bf2EefD5srdWSAoZIRlTel51ilXLmqfDRlENxr
FMXg25QDPmh+aKqagvo1VHVX2nei5TEQjm/1y3sMHNt5jcMOTbNebHi0vQfp04gkPO7rV/YqWa1g
NV6R6qjhnWZBroh+DhoyOwBd9FNYXpdntAryolCwCPc+fcg4WolWl8dhE0RXx2+8fn7EMRE0R0WX
bA4K30LgwoIWMV9OD45rCDWj9fv7ubFt8+uR/EfrW9r5vsgcuY+/shYI6UxTJTLo8idnwzTEQAOl
JT98oXSoG4+iznb9BPNf/A+mzRRjjq64VeoZjMLEag6MBSfeFVhClnuwKQBTcHjpxoyXrcTXB0f8
sgr3xi/i2PjokQuOBQtnL2vjHeXKaYcmKdOzJ2BT/bjFeKQoM1/w9+7fJZu/xskprNoW9dfStEI2
IysnW8J4fZkXoa3ip4owOZvffPohqCqBSWCfVhSFprYZVVDqNPlk1tLh+ZYk72l5Y5LCgqQjOmAq
5GobN5Q2ZvJxjlNn6KqXv7/IyAI8WNJOFdqgtrwUEcq+G95TMEY/tN+dS4rl3H+Z+zQnnN10aJaQ
4C00qFSP+q7kPyLBPN9VFo6re3ZZkIgSvzBBay/Gg4odmGvWnA63QQydQ3l9BhNlsV3FqfdwRbaO
RTjzGzHkEh0W27Se2g7ng1wuSHImSEZYBBvCnl+PxGHOm3+A/E4+utWmxQvg8hqmpcP6ASGTiuUo
RRioOEzsx7Msqc7+B/iV1lVCPvgAUx04Q3bFECmDjHCUdy9aNzyrHAvrmeEqhOxFG6RJdE5FAPtT
Y+PixunGPB4PoVD0dJM05rEUsh+J+rZX1MD3lqWbZrUdm5nj2T7IVhOGhvAWPl/2o11hxHImNJQz
N6tV8NZrGeZiW8a0Ww54BAzpeLLoyYTlFGZGKQ1s87IoGygQubczHBYnmkchtMaXSG/0KfYQTA1D
iukrV/GotzNMDLdX6ZERVQx/NA/a2Li/WKG0UmwFFu2fP//D9JmCXH+KCI33MdDGp8vFIk9dJfsE
HJ5aIdlLSNgJouyWHCitZX9WWjCXsstYTU9Y9SzIxqtQ4ZeQYn4u+7PbNQiwMIN6PA4o2g6jWwwN
zHW32Wjxddtr1hdPZMILq9a/yL51xNSppTnEE5pTvVKJ3zmwa4UnuvRkI1hab1u5uZr63pj6jNlE
O4blyzGoZ6Mrk3OIUerYRDApQh9wwRNAcUj43fsWNOzDF3W0ef7zkEBCbRaOqkmNXpWa4uhf7fPK
RV8elM0aDSols8oZ4Ueyh89E3aK7NZJhQoapRQ75ZriHEA/LSj9YYfvhVnaFMGbFhQUBoYU2gPGz
rwxpfhMvVk4VMXLu5hX3jZyE+5YzX6tSBpRAxTEnZTuwfLK+UkHpnxGvG0OjSAMJD80yaLKpeGsa
9mLMBr3oSZCKwX1igex/UqcBpRNItliRuVNNYcScbJUWFynWWe5dj9gumTRY+Gnc7eLj2wFk75CT
W21VCDsUG60mCAs7LiJ9QXkmyXlxBLgSRmkzYhR+5E3rGAG+Hb8jKvnk4H7tFyo+x99tuWqx/ieO
110/VD9zMiGxejfcqk+MZvHCfep0xVBTSxfN2DMTmXiQDcCDGkDEhb0912omWcvE2+12UOQw5fq6
2b3o7i3QGCnudjrxT51N5V13fsGsjZePXkBkHl/3iXBOgjxgYQe9JaFSm8vBpeltdVth6Q3axiwt
qa1xOCN6WOf6orroawYlcGpjNEKakqSVtSjZs1mhWbE39LotjbUZYNRWvSmYFPRXrCMeKxCipfCE
g1+85jKVLdmnzifqg5EdOtHzeX2opNvlY4xQielhGyKPpl7xPTNMRDQKsff0K1EZ5I2za2tnpkZW
KVDlNLaE2iQVo0/1qIKRG/IHPSJcD5rPQ6OYRE4gzaDMvLhx22fU2JCf7/ZlyN87f8Og59nNZU+m
HaDIsfkHHb2eCERU7F3nC9iPo6YW0kwxpJKVtDJAFM92jvL/Jbti1C2N9veG+9Jw+vpPihVrpYeW
ILdeYSPVn8MqnW7+lDQ0WUFrp5YH6Tj+43etKQ9lYnQyVq7Qq0qTD/4POQqdk5QQtFKquWMdG9iV
ZE1jZBIH9S2FPzZN78eOCnzwOIs+iknCBgXMRoVfdYbGG908FkXSBNPPh9A1zK7siRUDm7l0NFUz
5LdedAucEuXOEcxopGpO/ugplE5K61vrNjJmPhKAD/iyasHIREM7Ry2R37xBEU9/Vq2o3XTvxhFF
KqorNszIMycuEfK5YkQGf9IDrIhk12cw65EBeLNx3/aFLaAWnYJhjGtq3L/wCyC20NQIPhYTjCIZ
pmMbZaTf64/xc7JMsbrmCod83AxTw7aT17RJmo9UxQI7S+va1KHVTryXgThEc7fuXO/Ngnxc+vv8
t+sYm+BjYJ9+7IuUdMFLk19/2hE3we2ogixsJsCBmi/3Xu9NEvHeUfTvnAbCVmc5zovg6QC9GMrJ
/2a7JG6NBkb5yrMt8mJY/AenYNIKjfzp3SXUKNe0hcwHpdNlZHMMpTLM/izgBvLpoTUIb/gjHFNM
G+AlO9aMaa2j5oik0DaP3QCWIy2fJNfIF4Nn/XX2TXd/gVDks6YA/oboChS0COWlRiO22VZuLryn
js9NXUiz3dnrinA4NPf8k9hjQjbQKH4WwbKnfxuRLuuzXvdeiZxYritW266Dy2rn6hdsBHY4bp34
Snlu1IV02MIJHZW8dD/uRGUMP9CbfjC567pP6z/2B3sVmdiYOmHp9QB0Mv3WSTs36eAhgS6PiPIo
cFX5Lrubxpwq576c/mBoGTmSM2Ib/2jejP0jHiBNmp4GF8vbVBexl2f5u9Pw/XJLb0mrEuehTG9V
H8BhyLNMqfcWSBzPB0ETj6s1HCp16Z+WzgaupS6L/wejKiiHMYGNzxYtWnPdjyaqFyTMChVdOokP
WyX5E4gKoWjOD0BZrZb70DSZnBNIhUdVzDTvKj6nOdsZncZ9FHszCx9iAbhofyF3kzIkkVgMSa6V
Y6+Hf7gVi0boMMu47x7oj2SQrnaWnTNNzbRct0qYbj7JHcSCzsb+Bp+trIxX2eFmHjG26PcYJyyP
OHjwfCag6bGsQisi6CrODQwHEiKUXqe9vNNiSop2GNpDjogmjvmqjXHD6xqRkNf4b4IYHJMCs+nd
M7nuRLmCW87VWhiN8emRhC6oJG9AwA+nAvePxWFAMePT6rWrC0wunrJQu/VZ41lbZ6uyCYotRWGM
FtQvFa3Dbp3AwEV1kJJ/F4b2fihdSfLuN67J0qm3ZA5W7OxDNbaSFv2FbCUh2TFQqyRNaGdWopNK
DMvckB78im5duVqusvcVqpke0Y4vMCwJyQqIqEOhOQxcczFHj5Dy6UcedsQxcGdTUNFCVNZxyivF
rhTfNkqY6huOjTtdGT1F58OQmyooUUuqD6wgdE7QaXSe4Iq81VyvmXFZ6vE5jqk08AcS8C++erzC
Bg4so+9T80/ixrK1l1gOu/bKI+QrTdDZZ0gZTLBdHW5SHByzKfxJe7oVLPURIQD7/S9abNC4b/XQ
6VRuHEBkeu7PKGpOYO7l6aBVPcMQGAIIhZ91qPCEYI23ZlfQMJJ5FhoJIY83CRN7f+Glx/iPDynQ
ysSDUm/XGVKHj66pZ7mYhUfbSFyW46GVCxT6g+EXGn4Cvb2XvGIv7MwhTQEBAtDM1Um9BygNKhZ+
K7+4fO89F88T5lYfZID+VDNz4lqqBAl78Kl+HhA052ToI37KQkjozMT4qjmlyKib1oLfyAKi7yS5
98dAa96/h1s4+PiLvA73/cKp8mzbSuc9OpmD3Ei8Ji8mYQ7OYqYAGmPD+weBCMh8Y4m6XyyD3Ep3
pXJTWRGDhHQMfXD6WYQnOrtKsFxnHIxSEMdHDK4A5M5G+RQv+ohotayJhuw5eUeRKrKKG64QM40s
8qh3isHVNd8i8AMXV4nZDWnYzm2kGCNe6TZlM6HtpfunZ8yo0vpsOyFejuY37zMz5U58Fbvm6Imi
Rcf84d+Y0ohdeU8Bhl8dKks2M9jVUx26JnLX2w2/j1sJ0jVtuTMsOuyueKCpiTZcKOahO3B1MlwI
WA5CoLeW1evTgP0sreLRIn4lmQeEGlbt+7Rb9nUdgX/YX4qyt67ipz2Cr6pwrDjzOv/2RQZIyUVA
+E3/1vcMzir5vVVnF+R/NiTijWUJJHjXJMqqT/tLxlZNFAqv6aJLO+3x55Dmh8RENu8WJoZJXx99
rEqUZ76MksX/ImCOSxrnzU1+LqzmvhwANr58yTzYZfzy/02y35qUPL3iWj6O+Bt31aUscOPNwYO8
q5WvRzXd+MD3LksQI3UbwAIctg+p0NPxrJc2bLAkPkWeggZWdWvkyRFv+uIflWturw/pBDx83Zqh
QYcTPXDZoY7t7ng67nnmUj3n/H49dP41Wm/tkBBpvxAmBb3yBvpFLyE0DxhUYBfmBIB/oaRx/Rpf
5A8UMpccjCVI2ctNHEv3TbX5S5p1O4aU1QAIL5cZzsTwGpDNe7MtpEmJD2ecUedkmjCrGvrSVWM8
Ate+4Jqam58ug+IRL4ZiQsvS/fvXLzwfnp8lVw7yz5rKGL1BwEkBRiDIBlou151zbfDVTMtBWmCO
xnkZolJDvPO6Q8RJpQFfzEks9svTumvE5XC1sJxwRSiDkDVLKk0YAScNw6/577LWS97JwS0n09Be
INE/28f7YT/Tw7YjhM0O7ZkJC8jXQcs5upQalvF4wvhgsZFskCYQX3OKB66SWXRN2XXyv3+3MZdd
LVibG6ZUP5AwOfq122FMZZpVFGnx+rfhQVtvnRX8hCgvZ1N9GW9/6jZXpUgwYb3itpQjFYk5wQCB
0knkEqx5qAlJ0B1oL1k/HgvO4p/f2CRmqhxXI3NnfJ4aEAdljhBN0KHEyQWHvmHeBIfqo/t+nI+y
YDJn/rbguzqBSH2z1QJQYD7eQHhid/Zhjz4k6d1taZpjNoUdKkRWGJu3F48qfXZVy/vkRl3xlcfL
+nMhXaFf/9YT3oP3INWICKGll5sesFaFJHNmJ+iN3cGtAW2522gvS7oNhdY8OTzDJkUJ5AETkTMA
w8ZYRIHHDL23MXearyKiAWDM+u1lSZSVTEH1PHN8LjfXcpVsY/60TJA8qmh8faR8QHUKWyJIrkRg
l9Ty/DVKocrmqmJiaYydhGOy8BCmG3vutwu2/8+8bpn8oieNDvrXfJ1aSaKAyQudUaOoapIMu7zO
IktdCZjBaWsGwCetj8PiUsATEd4XxTfxiYLQ60c0g4FcbnXBmC6C48fcGDJLgojTvRzDW+6zj52k
90nmgU9zhhRIaaf5ATuxRupgW7uvggK8PCLofqpARag9tNd4wdMoBOlSAwA2lWllFMRQEJ+6M+sm
/3jyiJ42OFV+5ef7ZZbcj1tEFxQ6tnshBCRnIX2XCltcHaXEGEar5szqBWt7HDuTRezFCsbOpN1o
LIGD6Sxo1WKoiKBDzMJbYmA8uyRkoPoYjh0Y3dVbSPxo2MVo91rYF4/ZqOLm8blOg+xl5rqWRDRw
0GgDWuc2BBKouLVOJ0+u//w6xM3kQouGf3uk2hm8VzDbAqOBYEyaJUDhJi1ezbWngkoG9bDpT9oV
rFi/uVGBlNoStLBlTLs0yJsrGllG7tpZaWIgVDVH8BA6qFjeMGibaRxQ0ITFGSjf4zs/KS5DHS8W
NcZ2I/KwsTN3tLSrmIlPvXuD0h/Vu3oqrVqVjODit9fBGBoidMuCDXJKxGgnU0uye7Li7hlLQNJz
6WGkhGjQzJ4nl1UiSsEqyw+rLce92iuUYkpHj6iZCG233QzclciMm47fjuW9OnEmOHvX6qyd0E3/
DGLtN5X9tyBWZuHxXCYaxGx92YHRz047FZCZ8LHkYOB0z9hcVs7ks+LH4XaYEoLShsJbfiaE2VUJ
+G4P0I4kl+lgADi/YweQyCpLZaHGAsJ3p3+dLxZyjBhsfPbxiwwTyH9P/blH4+qZlb88RPIo/NWB
Bm6ng9ouxAr2y0IdOQtZgWwWhNnrCeFH9qvKEyWnNmhv/mCWjH52fByXC2C3EGdZ+oW+tGHFFw01
L/Gyin7bTSE8kEfs3T0b6ujdbmw5C8g4vGzEFwJREyykQZ5Oa+cI6fNKMhhsfnjxrk7ZHqEePyrl
al3wJrT3ZBAJDRPngfp1A0S/m6F74Os1V4v3TSpDRfCfL4Bls0Iqf9aHPLN0QLYZcMSpIfDZ7OuC
MHFJVvYQn/CEgG1DjhNasPF4D5wjOGJKrUY70eOl6358i/tX/r+HckIF5+L8fWJWBCjraRLyjXMf
xrrGvEAxs3848Z2O13DML28jOQ/SylmbEJFWFn9+3NzSDo0UTsd0l2PaK2B8A0RIj4qEA1yVepRL
LaH885PCYvjpHKn2x9pjgCRF2427xAbSUEzzTu1FjwsXx6wOeeWyURYAFPfoQwvxkN8/UUq5qapg
7/E7KwHRnEwz7dHxobCx/St8cPXPvNdnjewX3vGGse2B4GOe35BgsxM6VPsg1WqtYatRApms1sxB
4Y7uSLsSGk0s7ZOK3Fsxu+e48J6Uj93la8Ff9ol8LDmwgvhxoYyOSxmS2W63nFHpfaOYSqDfn4eu
bwZ+09sbG8IvPPqF2r4CLD/zz1K9iJVcDAD487gE7s+GXzvX1aXJu+KUjIL/4ZNkxikqIaQkC/a1
nqbPDR0iWWXZ5+L1LgdMmi8S9YChWZLAXEfsooNsdUVrkQHfJ8RuA53Yj+HfeDvr5v8Ax52m8Oiu
PEGnwFJFLb+cCiMihODfjXwcAFF8yUBnUbgRs5LmZnBtBSE7E3umE2H3Z8dnNykOtNaUFjiv4BZi
YL0QJl6LYq3FfuGOsEKeRjNZ4WGGntt5fEVihpzCkVD3f6GfNCHEFmUs7CDilDZIEUrvcRKe+Im9
5QUffgjBhU9i0Jg0gV5Vw+owaabBQ+nWSGkpM87nZFTanxSG48MwhnFNV6MwfDjWJKVE7itANjKm
QYxXW/IUIWaRjwAFr/ivS+R/MaGMQB3HPQMGUEXH+UNV6tiTaQJNKpkDGPdqkVjDkf3VVUAd1CI9
cQfaBKmxURFMEd8RgasQxEbcbFT1VHfMUeEmbDnPxw5xin3wfdzkyP1mzJp1lItVWbfwH0t9C8+x
YD8mqKuhwqrK/0w28wHoyrunkxM/C3fiztlMVnv9VnNiWC6azI24uCOS7SM6OzshUgWonewLgKr7
ciWB5WSXd4eW/0qAyvPw8q0+g90DP1UWLqKDMeSF25w0t1+0bIijj9G/OOO3TCXrrzbOis7x9S9S
rZ7vqE5UnhluBiGU64ZKPzjBWmEoN1v5uhDXYDRAJyBqm/CBvyBrYxlOuK/6UZG4TA+LafMKUR+q
d5gQitJ6IgEztVWN5gwfiv9vL3KY1+jwO7TOnR4LP2qclR4ncKad03nAuuq1FVzTgjPCkqru+2Th
6W/hINHfku2jeYJ+AxGwXOCcSl1ojTkZ008F81QlNhUBHM6lfCbvWnVx/O4hWDRvGhyZz49uha2k
wLXtoLNqaRXmhwc1k7bdvE0GSipA0mRmiwbADXj/J357UhwtukgDaELjpDrZx2l+eJgt4LI0nF0e
R7qhze3Hr/sIghceCUgoU7Uy1s6X468jFpkd0MPZlLy8Yj+NGXNC6rUQZhkGiF0SN0WWhtSK5wx8
4+otqEWyNlL35qsPqfk2/Bkn0hKcT2p6AL6VTaTgHdkrBvu5GccaKWbMqF1hbJHdJJIoOmfiNCWb
FMUcsa4/d2MmKpmhc9o7BpqSFTmpdqnvIaekkv0Ym5IxGRQMi5kKwR8bstbdF+4OGMWsvTJ+v26J
Qjl1lC03Z81S9asu0NdASzv3vOo4JeqzYxj1zCNh+k8TgUi8Ht0GRL6XXCCPPrpnlhrR383KF/C5
LWmuqEapk9z4qqQJqJbSrGyeuYMyTT/BHvYps2GSh5WliVfrvi7L8HGbrQ8Kw/2MfRdza+JL18tR
eDbo1R8ifp9aqokcGZ2tmik/oHN1grMCaEOaK4PvEd4YR82xuySTZKCmwWu5B5+vN2rPiqYIDEFg
qGTcOw16nlQ17RaVYEpq+gHPLEzo94o6bff03U+xu5xB0h7dhHnB1rJMok0lUMv34r9dLVzGhnUk
qfsQbbmlhl0dzcI4HEdslVE3URqSKqwlqgr/Tn7sID1wKPWkjhjTouHVcgiFwrBzAnssjOu7mnmo
z0oJEzOqeWzwO1VBjND5unZWvvhbiWwwGLAxmXKteC+BWL4QXXd3U9tvR7cCiX5lZXwO2hmFOiyv
MS3wvZSU6dzj7O1Xhud5zxPByBxljhUfkKUdEoqQ0uIXcL9G0/0IhtV+nI5Q/XxNmk/IrtT6CasE
eAx9KJPiOYmsOwzHSeLuzGI8cK3y46xvrT+d+QKd8zu1pbtloAsB5VEpZMLpTcBqsiPGIS3axTXZ
iSTE/gr59Smcw7u0+gp+MvtkfVZvq0bQhDfggfbJKjYXgRQ4UwxyHnZQbn0pcXmx7jW3LUhihj9i
PBbvnXMPg+SMNVW5GA3Rle4Gnzv+QSv0lIZS5UU3JQ5nWbSq2gnwwTTGqAzfW7ilS//hz6YJE74a
P1vfJat84PFx/gv4Z/ni+k/Tn2S9c/KOi4mLLebXFz1+qtLoj76mP+IUh0mV9ck11HVz1uCj7lIg
wERH/aiWH3VvZXeT4Bky6oh5Nd5iHeSzwD254Azegf4+N/GljguHT+N4m8Tt63GZrVvJ297Ho3oX
yKXYGuNj0kvZfYBnPgwuob/EOAuIjtnHkn5vn5tN1ZJTlym8kPjJI7fDn3yPDq5xhdWQOnpXKLM8
KSOhiDQM1yDP1szN9E7SBpzrRd8xl99MT9ODvaojhE9ZjLNFYDTsTslamqDJwFd8FIrZZ3QszyGO
hPx7NhgWk2aeeyi1XLrFntXgPp2riXPcI1AhFxmr8agxs/BeCfcYTFU73RISXppmppxNMnU926e9
oMfk/VaIe6jjYq7TJeiki71MkLEHIw55m/zKg/IOZ82lTIQORe+eK/SP3LSxDFLa9mwrvNoWoE7l
CwqUGc1hIKh+NZThzgGMtwnACWoWf8c7WDhrcSy5Xjo+G4HaCtq510isy07JaoAo+tHKRTGgNu3K
ngsYmHr0ht3SDhRl7IflUBt+ER2Yp9Bia/eXmXUKybOCRX7bEiwx/m0F8dud1tBAEVBW315Yj1HL
JY29m46g/qHgMsyzcC9ckjny6hrG7D0aIvPFNaxBVBwJ4YY8u1viY7TnfyPQxKZz7uGhcg72UYLZ
EDl/LFA7tRG8IZs4fHQURcQqoW2cvXS/lW3iNTnmbdy5bwQYK+vvstxxEEtkcJAUsiU6WsbnoR3z
dHpTPCZlEvGBbFw/lblws77IQX2BVTGZ0Ffk7stdSvecVi3vBRGvVeYvTUv3SMMHkXXpmKr/MFT5
6syO93PJTKIyjcwxZhSbvTQXalj+HuC5UzXaxk9WbIti010s3NQ4KE+5B5q4c1ZsPChJhp56aFO5
V0FecU8OyL41xPleYhaBFO7Jv/kmjYmw7EmxuL64PobjOckTIFM7CboLQdrATmBPpdXY31fvmXQz
J0jpG3uVv6M1X6A/W3CMtczQ6URlfovrmVyvxt2DBVSHl0/pu8K/6nP2N4ow0PPrOKmJnSfeoYfD
rSYysSWtaEhTpu834O1RuHu8G6QMTS6mBRMbPG/Lg31oh/MSc8ppPThRFEy4Eai9HKjsrhDOCTuH
ZCEu+u7r148arufFDOzU7k1mGbAjfsGOrPjluRh4m//BdzAy3xdWx0pjpKzdDnzYZcjjwzxqSaCy
G/2u+ev9tJCImie/tRWE08lEcn2Siaf0ARX+OXe2AZ7II7dSXL+drOEBoNis+Y6XZQXaIc+oCaBE
+CQ6J37GxN8XczEUqlSZBwZiVOMvKA59VXZM0z7RvtlDrfS1yj712w3o4tnMitlxavCG2oPGTLNB
OUVfyIW9/cZ/g0KrjUSElUXr3Thaauv9uwIBngKoh/dAQq26So4UDLwaqMfhd5OCZbqwAvMoDKR3
M4/HYCibiiNHgv7NiCesYBE+r6NgyuElimaBUg0mekf4vocT0ANU7FTj+SiaiN2yUrvysVZXPMC7
pI0mKzDcS6Oi+4p8NU6tJJzSyc/bh0Azg4+bnj/lCuvApgva1rgTGLoSfpj0EpgkAySlB7EGURY2
mGIqF7bceV47SBrSK8HrlVK058cV3fm3Hpi25jRI1r16DsYh3fv6O4wLv8vROE9jchLGPVXg8lq4
2j8p8Qk+08PQjvlvScd4Cf0zJdpv43sHFDhUCcA54tyS1TLSuBbzAJkXLvR17muNXZPFTzaBuZSj
kYjzq4PPpXELTMw6mv2CuHPn5Nujr+Fb0GrfXB+OT856l8FACJp1hFReCwSn75WlZHx/tMAMTC4N
bdzPd5aYbaSs70L+HvZdrtSwm3sPFiQgJoTvK6b7UAccPbn2oKJzFETZIQx4YIwUQpcNNb6334VC
aX10aqQoxZa32uN64VYMCserfHOx1sGsm83NGFit3AVIh7Mx1GODptBVERopHGYqX6JQhyXHzLz3
49JYwL/+0dy9Pu9vT/KD9lXWDfoEqBH9eBLmB3OQxWhi4qxftjAezMu8mCOVoHE8yvCsYne4fFt3
Si/yABId+TAsI8bjKSJYsJWXGIqzhIrEIKPrJJRMaz4MSHFuln4I5oQ/Wj8JtsJNcaec07C929wc
3c3DYerP48+L4tplB/QXCBSfonupwy+Sv4EuzcwZz4oPppMEm3+AYmk4zYxdb9vWR3D4sA4yLPCJ
o7/4aAReUyMDB3qccBIUf6q++qWJuQe2wLlqRE13LZ/knqOxxoFj5hiXQxh7+2bEU7eAybjOIdGN
s8l1bfS0Lz2R6gz9DfU8u05PuCfTE/POb8NJMd7i9aWN4kaFhgj/emqwlxQqW3oGnCy+L59z5YdM
FbgMnrJucL/Dz+S5UcBNBg7TSMX5i+cFjR9ZgNoVINl/7N/0y8SnAkzGA95LqO+PrlgjDm7rMqWm
p/fv6qghUD3qas17B4pyfghvCBP2ManMW+NqViI/x5/o4C3PcL2NpXaDOezbp/edpJykeMgI03sc
6x7cYRniTXq882piv1d9mXsYKrUqoluXNOTcujL49SQgorZWoA+XIdZu2dmdhvdFgggp+QFMroDp
nZlnz//Y+aOGLcPZ5O0HQ8sr+2EvrRz60jCo4khlGQhwES2NXBOXHAEZTqrlefJH9Im0w34My8A8
qVac0/asPf6IK1kyOFy4MfY7joeK5S9asBzhN7/bOY2TDXLMu+Y7n17ogSiqvKOlpf7r7xP8nxQ7
Z+059SNhkr9Cmfzub2kkFWT1neteBPliAyStSwm380zFQe9xr40i3jtOVMCZv0VjmZIFaB8We8xC
A8zbtUfBh2jHqM4SIRlAPTYJ1H0oeiJ1Cq1H86JvIPYWOAuEoMk+tub/sOJePB5FjrSWQMAnjod4
9UuXe5tS4Y6VB2vggEfiOxEAn6gyL05VUlCnG+uJcrojOG+8HRvSmh5xiBuUr7DJi/uk7Np3Ce6a
qFOCzHijlZ7p+Whgd/rHWf7q8GO+cPbbVe9/RRVht9qP57r3fQanjh8bqyuHvHFqV03NjVGF4lk6
yGYGDRRVqYIcgG0YdBjaRKCANE6KKmwqFapYXCQDoFBJJqkq9DhBCN9WqDNGkx2vQQO9RemYr0qG
Z5byZ3O4OsAtVKJt57PQLJg7RyWAKCDV3KDNiaZK0BfwJfN76Ka1aUbTY1a8larqsKDsYCAoCva7
bGu24rLL23UmoZhHSBr7pO2r2qzPGMHdUdQIEI2nINy7hbDCcfdh4FQET28k0+NrdkgFoeYTm3jU
VoHQaOhET7PygLdDTC8//WcAZGUJ0OwCih570kMdXNfyckIZgycETvxwpF26gHbI/DFnepTc6nIU
uuQ2elSTNm9SZg9QMIehvKm8wtEKkl8s04tt0lwwEGV+XPD34YkK7dXIJ2Ui8ahNXBxLrg8m+xMH
5WmAKzB8eWAtohCW91ftAh8z4U+6i+mZZ7xDjjo6MHRusVIMiNt7Fj7hwYLrmavKGHd/ZvAEMaTd
r+Wu5IwFd609X8OWWU2Pcg77fM80RcE7/u9Eph6rMNSOh0R1iekoZEw61HxiZwJK3vNBZ0W1CBTm
wK4SXOzt0ngKTGuiO6xkSIwqx54yKF45b/lYE0HFVcyAY2WqDEuBO46Gn/87YFh3UMbwJ+5Yaj4I
V8aukXWnTT6wlH/qsuxBN7bQdXMO+SPrb/h/3BlzM0EkL0Y3rte5JsDUTBVXuY6D2gG892sxVzFw
98nIXWhhHr4wLWLmvTVV2VZcd2wde7WlYZehLJS+399j2EF7aKxKLIBOI9WH0W+rnMkPq/4hg4iP
+NcRWx2Al+3LH/+3LCvS5MbCWN2YsopXWBV8E6s12GpX6gATVf151k0PTe/OyX7rwLBwE6FiJ2gw
+zpLF/RsET2VKQJRktUigezaZXh6v66wN3GnDgBUpAV1qpWkVnI9nobnLIMQ6JLFgHQim4NmhtI0
WMxiMo9xhFxp+pKsdcQ2RX3UlUJ7AxGhgokpKaFiOoklRPnOft0jIf4azTMVs0+yhdwL14teKaKv
SCJTSiZyNUPQxd6QRlFRyG6NVC12nfnycgUudl4WWH7CAkuNXTSRM2BYkyDfvwxFNmj3STt06yAA
gtSYKocEPusMZJhMEn1cr3cFkVLhcEOHEn7i9T5rCG5JMgSsTJH5IaeBQyFZs2UjIIUE3xz8DAe1
U7t6E1CQ1gz4HSJpRI4efFGNL5jOQ0j22U0se1ZNFGB4hI8ZUJy3MtBM8uIKRUz1n5ohS29bd09u
BxayGTy9+pXhCL6cTs1INQaT//xe1vx7pemDHZMYoykG3fyVRHs6JID+3dlcTZJ52Xw+kIIgH7uz
6mpSHwRBjZb+cyiQoRAXbd2eDTrXyT0xcQKxIPVF41sHZAB/iOvlv08CMQpvO/Tgq+gUkWpZJ+Q4
CMCyVzbDCvFuKXEcng8flwEvKmV2Z66YqFPxqNqd1sYZLQhrXagK97CHiWyICm/VlU4Vl0jhH93k
B37Be/3cD5HaNQQFvw2W4pE6avFJSQ1AbYtgKDGvhzERfMzoxCd4Fyo/O21d9a/ZLF6EhfARSIQQ
tuJmPtdAqdSO6iAuFYQ7jjY/B5FYG0StodieL71iqlEiNcvrax8UtbWRnCx6Vu8pzWDvE54yNDUl
RvdwVlk7npA5jZCSzJ+Z7e8TghkFuJ1eQwZyfwPzENkUhNAE+XD7s20caFM/+7lnDfv2M9aB5I/e
QL0Zb15jM+kuzDQJEgX7mZ9x/F6M6HXAzC6LsFXv4W1oPSvEkx38zBxydUsd7i0U+9chOLPhPCA2
BhT4nC3LbrZEVgytW+6AGGPeUVJXM4jlNTll3+VTpxW8GtCdysAAkgeb9SEjX9j4u+BMTGNLovm0
zDsB9ae/HK4xdT6BkdC01hFanxIW6Pn7xwYHu7PgJYrQb5Q57jk52zVvkkZTG9OW6wm0dB5vipRG
LwuTP2Gx/cLAtyT9m4LCb43n5osAqgDCdZ9Z6nSOVaimTpGyqcqDJta9o2W4hhU/1axNN6pMbE/+
Rnr+Z8swcVsv1FxFfOfhZpVBEvZ/QyUx4WpyWpqKFO6tt97uS8jfF6rqpyqv0hl1vpk/ybpy99Oh
G8tGcvX2/E4v+Ny9zCsv1gxqK+TE8Gp9lxx93bK9fFh8NNrLHUy7CfRMqre2CFU9UgmedhVQ7ZnD
zzuSrDqOmcqxTBLTdeUIGh4CgwT8xYz/teHUr7k0tVYf4wHGd+K3Ml1odgT7jqpdjeO/FDldy3nE
WmPEt/R61O5JMoMC2GOSWa+jYCHxoGAImTca95QM13FpUkGjYoFI7H/8Kj6eDY1sjVbjrKvfR6Du
0Cd3OtFhb+PaXl9Cr7PXyd0l1U4CabzRpiE9+eEYip4AorQu8kTcfUcVHNCZW1Np4uGJzXk6OSXA
A428xtsxZaSuUJwWw2ERCWs4Fq5gZ8Oljp4WkA0HMJdYFkT/g7UT+q4z39e4t+ARA5ATpwQJ71Em
N9AqTnqtMI58NsrIPXTrnZCKOIfxZgQ8QtCCQngVrIZkgCD1q1Ubqhzfcc6x4I09ot+7cHJ/sRyv
RbR2QQrv+aJ0Hy7Wz4fCBEB9C1mAxZd1QT3r0MdAdtaLedbIx9sy0y37L3LRfKLdG8+QUtZKyaBa
dtjjLH16gcbD5StYrcr6NTfCdNYv832KeNuxfQ3Pa0knnCmBRWzTwzdgyYxE0iJl7shYNx0beI/L
9fz1aUllxx9A5KAD8cJCg1/zZxV1KIF6vjDNgWlVo8RjSqYoMuoh04Hrp6HNK1dEkpNWCOR2h7Mu
wy0jEK+KPLTJG2C4JiYEfBKNSTojvQLlONxOezk9S8ATg0ivqf3Nq+Rq11/bDC2c2zinYiz5VkcL
qTfyjek+p9berC0z65N8u+izm3AZQsyRuJm4ggfbCN/vMRE8HAnobe4f/NqE4Jw+v+vlCUBbeFly
NtUzeqyvFlXhrcTCwmtuCbNS+Xl7c+8n2W8Kki9RhwfcFclVSN8LJRiD2uQZ8H7tzEmbpDnoPbi8
JSBoDcQZzARKb8501d7Id1U9DphCJ/JYumCI0IfKxAo9GAtnVeveHeVBfx8zvlqaK4Y5ijdX65SH
1651BgcsD4RuBwTzSLMPF3+Tm1mdjcFwPEqEkzqSdXz8PJDpfgVNGHTkWcl+zMnTXlX7iL63gWmx
7ZdKDjUb6RGTKKVXQdS0Egs1lQzUlb2qfGa+MeGyktPaRWt53nkxyHA7oaS/hD24MAQaRo4x4ToH
Mln0dKhcPtGMSCa0Vei5WoiZX5dNa0qL+CHRE8H/fcmDnytTotQnAdoIWnPOhnGKE6kWDAaSOxlb
SydqbkaIfchwEFIeasLPbl9ehbzzDfV+tg8WH3U45jdxgAN1PJW/HsK48oh/tDVOCWEFAchPs33X
/6lRDvyzkjkUZ9pE9AD+POQW8bsBqWdyhOM47AZIDs5y/sm0qqnsRaHzSWfgVWmQUiEy66YtQEtV
gj1jqcwsIvQOo2H7xYzE9snfbZ79fLxvmUBpY4kDtQX/eXaCVEQ4Zjbe5TzYygzwfO4ZEe7aCQCi
Ke6WGQQvY7X05liycAKdBIy5Mn5+g+2P8N59c8IfoZvHLfwjfqiPKL2HJU7RgHHj7XmoGgHpClec
FCaPgxw+EfauI3oagUPDHgSTFXfrSj3G1URvE89xPepa9FuwVCMnvjqkKP+fYKR+DZIyAjCr1ZHl
pwpczgFKMAgfHkGnycDrPdMSiOetBYaV8uVCQhUMjmLZdEHEjKTgnneorZ/4eJMe6AdN1byZQO1p
IkpheoVRh0IXPrgFJV33KK73cfRfxI/HTSxPMEPy6FCEbhD1bGSHd1/2xmbczZdfUGQF5M2ZFTXf
peWAI18lUfsWVMWphHTjbedYD/W6poKtoiro/eIBq+2bp1scXe11oQXVvVjpVhceId0WCxJ1x8Iz
N7z5v22MgPyP64IOnEEyD0MOCA3f/ULt27QeGXBQj7jVVVZy2KZ8ffcJN4l3dgJdjaxcyO/Bo7La
6OdJFb2hFuPaLFLyIXj7p+bfKLp+Rrpd4N8qKsKQqMEu5y57O+eHKl4+joXY7BAABSSr5gOQ+nvx
rC6Obpg0CzCHzgNaWSihGVlORACEBvDIb3PUOPI8FQHcZSUJVQGMlAE8YDD1gqjANuItBZMbg/Bd
Eoot5iJTMGphXT19BkTFgtjjsj2tfGrDyDZ2eDSf0CoFxAwRQlpPTFyKtH1gDyxOMk3oWzQ9pQBU
E5VOFrf7c/nCLSdgVBhWBhJlejDLYoR+R0URfIA8YdfDI979Z8tAr2vxy9mi7JYigZLjJSthNiLA
tokmOKo4nWUorbQjb443OnJiP2J2dEkr/Tc/vG/cfbBO4ncoMBNeXvlTOQBTOHXsE0324RxaNreO
nGAKwUd+F214sBgGbEWIfTGEUtRUIOD0BwPCckcNje12kR4Z91nj8M0HpZmGBazgOk396ZG3DpCM
1cKH682fTca2ZoXXXAwLePHH4lNp6a8ct/PYuUaXwUfycmgxmOzX08MN3IV1JvLF7hdmNvh/BC8f
HgZOlTOs5/IMWfR5ywWRpghd2LOZy9vAeMF20gw+nM5FmchZp/Ney6weuM/ZKHZHNV24yKLRtvaE
0UiZEKoyfYpRQHbWtfaO0fSFAx695hFUKJaAKqimpWM8XFt7oPn2J2UsHrsYOvJrPZpRbznv41v/
d0icEhbVl8Ilv7wSRs9luYQ13ub8l4/9KkUIUXG25K+b/9lX1KURvbKLNg7rN/TA7otkrRgbWGyg
Oyj/pGx59NtKwVKKvlQROnhZ//9aFX26Oi5eBd4MdVnC4u0UO0SNixvdWKsn0B3+qfFP5cGPlV1x
88nxLqFhUHGaNrstJq8cFctkWoSnklLntlnvTGsF/vEmBxMuufYbV8OpQ44kcU5LyxgoFFNXht9Y
kIhs3PJEptlN7P/ycHmXLftDBB84y3U+MVDwrB/ZOxa257OY2hFPYJfz8etCkJCFyeQEghEWutG1
ADTSVKCveLjXe8RAjQikXuoNSbIiuaENizgNVq6auygvMAWdaoRDTZ0R5vgZ6WFJp5C9GTQRVu/J
cnDdJB57QF6BAAk8bTQd2C8y7XcEP+24cfj+8/Y5lmFqO1475AliMIjfyMlHcit5ZswDUkaXFfkj
ZxqVe2scCy2X7QvWh5Cr11IaRdKUy+Go+jM5Hi0t5UZSyROdf/CHGq1mtRNBRVV2Kz+sLB+AHavb
KHDTqMN/KIpKL7VdK8DcNxRPdRM309aaW02mOvFr7vw2lC2qDueByFwaNOvUAylfK9lfO44rQATB
nTzqyHBuBncBIsy3hVUn2+7nmZqoWQjSFLxsNLpGmhTs60HAcEg1uVALJdF2Stq3MOyWp/RVb6CH
bXSzFS53KB+YFKBTxeaakZYxB04RqaTwOTXi2LqWlSEg9eQSWtpxfDM+3FxG/07CUmvmexB/n8Ka
u6U348dG4iE22qBK6YoK5liG2DX0tA1t9+qxONeYTqgqHQAYIrQJBKNpfTPHVwVyDnBADWMOEVcS
9q9FCwwqkeeIqM6G0s/3sGEZAmonw4n/xvAhPw1+T61FswO2M/K7ujvxDejJgg3A2wEECkBQ6HWS
IncLuK+LMyP7i7wpvzXpbBqJ5lHbA/hA2AGR4gWgfpqeuDdQdb929mcKTr6fmF5Ufy5GYP4bDyjz
mq1wKgay3FlGequfO0Q79y9YUcOFp6PerCGdqOjWIDlX1iAQvDmpsJK9SLD3RmVFNo+44EsQN0fh
y+NMoCHenfFbNOWJ9GCEOgnkxuTyYxwnN8J1YJMCxur3nvDNwd12UMHttC9midTbHlgJSbS/gCgy
qaFT8FSg7JEZfJeU5SxSNV7b8q26L/JqY3cYMXvBRPUV+NtswIS0/MNbRsSvJDqxYV1Mhh9TlrBG
UuAfYB+5L+2q/NUXKGClMBB25IvSgnfGC200xv34GDOxwf7QyJEGSojZ7M7sLLclbf2PmntU1pEa
kNq10RFagoh/pYPviUWEwDVWXNSN8+V4r8B5hBJgroYJSnkrvJ92WqwP89cSlVp7EdH5xUO4NdZ9
EPxst9jGgHD+uR3hQQ6nXYxHzu3kQiH/O1ckytf9TjGw1Vt7Pi+/a+bG2LbrGhViyNLMc6LKiD5Q
mwDtYIe2AfZ8i9cReknNp0y84yaCrwXmig9PBf0ceWuY6UDnBmyg3fZ65AV7bApPkw9Wb2/mvMwv
IpR5Swjp2jWKElzsbsT8r4cGBrTJzheU+Sdw1kiHw4un9YSp8RC9eXhXk1S0PKPVah0zhpUMmELg
Ltb/IkZO7i6YseOMl8c4M1m2NPolzJgMvfXnoSADKMgyx0EefEx6XdThSxvSuRL/zHq8erNLo8wp
/F5iHAwktKtMSt8lA5Si998fU/3wxRedTsB4+R2m8ieAnhI7L1g0F48Vx0pkvGhBBvGCMGKi0RHt
DbyfJRiAL00ZIdYnvgnMu7KdR1GLTGlO+sl+npt5RxD7P8SY8P67VgL6jvM4+JjOh4aQeeLmS3XX
+mQwArVJAPqYb+3i6UGadOqMf+rNFkPtDk0BjRLj1zk/cHrh8v1MJVfC8r8bIMewFqR4SKBj317b
cP8yPgwlytM8E7Qx7rhctAWJE6XoO+1wK/wW4FthOjFW471/DWoIxInB69mdmAMJjePQjyoM6/S4
ZfaGCJhcVMWjraIlfNx0Xciut33za+9jP3u0M3lzKRdFLksp3vmCMYNXXjWfemp+1uvf6RsK/d31
ooBy3REWp/6mD0LbKOxChyr9aStQyu9pmL/nCzBGaMwCZYZkNziY3m0JFB1tqX5nZEkAB/hLQTvm
mYJotLCMbsNTKjNBs6m2m1+8jrsRgqiF/NBLKUCSfBBaWvuZf476b1hYwW56Y++GTNahfY9jB9In
gZ92A2caqsxK93ZLVXOCuHcxEBvrPiNH6gmgjvGKY+6tktsHH5N9vt2dpzGOlAqHn2loUGu52207
3s7NS+QoTqcY0TsT2YtymbYhtnrFdYBCE6kGliPFHwJZ38rAdj7CeXqW/oY0Izaz3IuswOEeXDQP
RlVMjZo3XfAy3H0adlOSxQx0czDuagEkaRAMXE/WuJG7D5C0FuIRpYh9JkSZ6V+ndjRhzcqmOJj1
3zAv8ues1dSFMUv3QS1YslAMkN+mwDtwow9+fS5L9ANolXudHPzvY6fbKXzeK8mUAfXo5Xhsj96S
K6ivf31phmpzND1cliC1Z7IWh2iMo+I7NXUQ07S5hc0abaL/p4AA+xm0LP2UhEWHZpSLU2mT1uY8
HI3NGWbnALHpPhwpjL/FWpjuMhddrsMPM8ATqq4NdP0ox+LMwHhHJROBhGv411WGK8OCIOSWUn2d
+6oNc+2hwkTNYhGFiltNsSbmdEC9z4x5/3v4ZObnnyvTLiFZDcBP420+7YwDJ6UYkwQx5t4GJHn0
R/I9MWBAO/zx3iOjEHwInvoco1X9yNskF7NRj2RhWEnyGk95knGcpcKFXbbaBsbI58/EHoJudBj0
/6n5+9nQTCRasFZK/kuJ5HyHub0SDMENEApduYT6NZhSCXC9BXuwZ3KTOMfGcfefIVwFQuu5u2Q9
FErcN5zdB+DBfBnt2rnCamEacx0JbtaffyorsPH7gprbyrcbrP4m7UUTCuPMk2KWSwGOdaXM/9kN
uAGP4F4+kFsT9M4LnoeLoi/T5ts7h3uaPsT/RpHGR4qMw3x/B/kBSk6tRp44YbVgz/4MK+VvxJq/
RyUE4S6GJrD8j2bQBVyBBavXW3cpBYQbaiBvBZr6hXnplPcCV8SsLWNUkbHJGAPDCpgY+rTpT/V7
dd7gErjjzEb5l8OPrRXzcbD7Ys877t6roQKhfluIvo8pyljNhnB+k7JqcAW/BOt0o/5edSDUrlPl
EfAi7/vn3NJVlA8cCtLPm1nTiFePv2oqVxCy7a4mQaX6+2K8ePIuD0rBN2GMsPR5P35dF3319Lt5
EWt8ZolCS1uVl9gYxIYtZol8HCxixcJ/eFHZcqIKqK0MvvItN9IEcoz4cQd32QoC+U8lj+EU9NOp
lhPspl36xfOi1Vi6sGca7kwk1XQGNM4mYbyxYzJSaFQd/ejEGkojFr5ZNz+wNjAgvgfmIhWJONvp
kMjsRb94sjFvYpOiFb/2jn4TQWsO7fCv8zT5mnNqDNNQQm6ys6DxmBXQLGdbwXk2Lj9B/kxvbp/0
DVs/MWfgctGT5xMJEdvm8Ed+I9pY9hlTXpZgbQB9GnPa3ZQ2PEnLWaQfQ9GjhX8RwRRhal1yR/hv
dw2WDHp2yJf+mGDPEgu+UelzzRjsqn9QSdQc1o5KfuVYkp23yLOoMbaFVWDqcp3bX9YPsqB0fjSa
ANEwCjfLD09VjSltaC9jgcSO2FVfrDyfYGwD6j7W/k5KTcq9t4kf1vWw6sL/c5uXPj0OEeyyia03
c+Q6+aPpBUcwLrVyklnaHbM73rLZnSzyi7GE2zZYPFqf4qaF+qcy22DEdACh4zX4NZg5QW8I9pXK
U9bPYvqYTdENsn0neGlSNrC7aR1bwxu7wyneic0xSgukzWNKvfFfPb8PH2kB5Ipu0W3wlYl1e9O1
HWOUkYXKj6pkOBBB1JTsfcjgyyMLJIQ50DDH6aIlUsW4luTIDosw3g713jqG+u6wLPADE9S964Q1
tiWdknMhU2bM47cpDkGop96OUoGinB12Na2VzXNLXh1H68z1tfTHrLHno6j3HE3HzFkZKRMvZCY+
5dQOGMtTB8Pw8AFOWPTkv8+cfutkSDYJZX4dXyes0f2b4KPuAurcM4DAp2BrAw7dbhB1B7l1F2jK
VoNcljXQuIbDlvPVoq/N9UEEBUdS5YHaG40tKo6gPDKaACA9MbdaQsbshIsriyQ1oPB4S0oxbDf4
pfTVSCxPdbT69q2wh5rjFI93EChBU5De5JELOZVOHUz6k8FzdJ4FDONV6D3oEauWkmvKxvXex5Gg
WsCuzAh1WYKYBVfMSokqB3E0GsoFaOcrDg+VIym6ltKJfOz5Sj5cl/x/6P1Y6IKbRZrjJx1M4YPh
YYhlco7WQQwzoyJr4dk8PgpnizNdKPW0yauyNE5xg6E1m8jtijLx/nIJW+kft2bTiXxlQEFsPA94
dkbFw8xZ3Qjt9xvVyOR60NQYHuaA5PhF96eXupCxu6tCuqXGIP35wyMLXn5l0CjTiGiPaYE7Jrhe
aPqG8xIT4LNbQ5Qp6UO0ZODa7eB7WEheNEijIjvrep/EuF54Ef64Xa8P5Ph6WgsoFhGTqkxAbTIW
L+x0oiN2uK+b02FhwK1s9BO4JijVegebW5OyZ15KdRX4Gg44FVzXkn8JYe2kU/WvKt4ypflN9WA9
7nrLmSBVEwESAM7N42gruGF7LHTXzWF79Ib9jifRBZ3/9iiyIcxcGMkWFj/ilj23SXCqw5en72fz
fv445qCVtkBsIuUiOOgggjfMZrs9V4qJQ9iCMddOyn1RMN876K7oKmC3jPP1VoYEU9rs6AyLDLc5
DcuXqB2nZ7zINkupwRBi0RE3ijkE5PQKJe4KT+VsemL6QAfBQ969GLm2MMX/6V3S16j3lfqJJzSb
wcJWoM78kUelpl1jDtm+kQiHtjbzIXiXp4W8/PZK4UcetY2dtKnbCPs8uusn5NDZ9pEn7jrQrwhd
FXA9tVWe2TIFUVEUWWl9WnUQuTPxyCk6VVjhNMAm9r9lK8AxwkwwaPj9BoYp+4vkRm8m+Oyb2/Ns
wVVEn1T5XbFMRHfs8w8UiZP/TdKD8ydS5c8j8vDsF72Xd/yPe06PI6qMMGmZZKpBQ4KHyjcQ8+sP
ogGtKH6AhMDbdJMGtTO4tpr4kn1IoJHupcSaccQt30fK74gsrkuR4qF2w0RWdpDJy4QNC4dxQHjt
6Ouflgy9SsyFGH3PykebnYLiartsXGiXB7AoIHhSVW4DU4TsWyXcWeoHjuBEF5b7bSYYuepQNSXC
RRSoBdMzKtEkx9MQRoSHz4Vt1YwyMz6LB+fVnvti7KY33IyxFDiJ3TscI6zq+8uedkylVbUaLBZ8
OrBcaWxDK7QAhjnPI52pWqU6qWw7XHNJR0XcXXhk6bpC1rzdaHJibbD1+cpZNNduDBJdbUSBdNzh
Pd+gQXMwM9A/qKs1GG6bDqWfbA2sJIL+JrlzT93cDiv7WwtyEpxHLC6EvsqdGSE/1NEjjibc/USW
2fO5X6wD2CsfvOcCHpZGHZCB8ARWygj1xkn09VoXUbKkX1+8XLMZOuENR6tBCy0MXYD7KU/fZvCw
eKPnZxjtWBAUuy+2rFcw7XKspNUXreD1mT0nOk9BP1Z8OLkPG0JjEt02aBM7Uw41fsJk4yEp98eX
LkkWPB0PUMxAbDJk758ZidJdD2lRLtU5cBSjqiLUXO1ej/oLX6aZer1K90VfzNJYb2PEGCq5n2N2
x2SC+74T26vnqeoQGpXfFxwG2kdRTkz/AoSFoRCEiFiTcBO4+f3WEecjztUEO+TUOiN6EHGT5zmu
Lwsc2tysq4BeeJTGjIUKT0PHC+OYUz2ix6+IWC1avGiRzcy5zi04XV/1EJwN+j16gJTRyv+zDENF
JRSQu7O6hAgVN1uL/moPcCHzGPb1ypX1MqY2EwlK1wY++0qsY6vKxJNlkSmNaerHWxlXtJjFEnuA
y3Y+zsonqO6lxClHBC/oT+1uNoJdabjvSwxFtDb1dmv+c24v1MygjUilIPyGNxWIVubWttQJSY36
8Xs/NZO8SwiWPNIdE+3+WU/QiKaA+XTOxlphqpTU3AtL8WgsuKE3xsKXJJCHdQV5YY0DppzJ8MWN
AcJyT/1DbXFdBUzSO5UrFvq2P5lJgadxOi0q+MXFtEfwnWcTYQ1kTTHZOReOt7s5/BtKrSl++cj9
iVRN7W9R7DB8pTAOm5m4GumQWfZRPhhj1qvdUhJtNmrmE0H+Y8mNV1iJ2j/Z4apzgjP8TfBgpFwN
/8m2Ixtd+8G/+SeurJWz/DU/MQELUnnng8EnUuCMNyc07XoaZMwYFWlPgryzGJGBBHiqS1n9uGrl
KchpVJJUXhcFpz1fiB2UHzsVWf9CrQIFCE89uTW2JjwXAfVMYFkXAkbUOd+MxEktaGKKfnFfmzIJ
wIgMomesmOT4wMC3cn0dIRgvtE6P8xSuYNG5xarytpbjzArsRH1dnb9L+Q52DOQlQV1uzvqX3hzC
OUrH3U/uvzgnJPkSXkxtLYcl4uANaG7WGt+Kgsnrdr3jB2Gl91r5tT3VRTvs4TVDshF8A0xG/eGX
fRh4CwwOH4+lTciUDpkmbeWthDUEOrq18ALCKBfZQa56g+G9pp5MDN+qZ2mr5wEOm5UkeK5FRxJR
eZSUEuHCrZB7ijbhBSBI4O5lHNrV3eAmotCFMk0+qUQChPXqtT4yFWHeoJR/PXq4r0gxXIZY/2jl
ro54XqKSjUY1aEgh1iGhSyCzY9ffZdyASRcE53Es4CIIsXKO2NKFRYO4ToBMnJ9H9EWk5X2MjMSD
Z+x6bEIX02TKVxcyIMfRnat9Bze0bK5Z5RIuQPWzmt88ZpQfgqnIfhroB9FvaRJB1mM/eC6/pcbY
esTGzvGJb8iZ464iTlbwsuuPoO+6u9FuP1UXrenUoB0Jg6Cx4lGIsu3mXr9heu2hCGshYhQ5bSzT
zT2q7Zt8pKxzN2SwYhcJzzsLMIse4XvrV6gEVZRhBXkY6zrLvEORaBMFBFJf2ki6y8qsM3J96WMa
Fd7XPpBaKdtRPqkyfSltSfMCbA2mYoggtiZUK6Ola3B1GfVdMv0DWzVTNzBdhxj6C1R7HYtXG348
MacdFPqK1SUrL0npDAsr4BhqPkrrkKpUoqJ+UpXn4BQKfIdYRmdFHg49e9ksG8c5UCf7p3tiTsH3
xYkXUMfhqh29hkLXkH5fS0pnj5xOB8kOQ5jZAEA2bqoe6Zg3mvXOQfgEVOv8LCq+wLQ4e9Uk5xJi
wRy/kdCO4+LKhCsH6zRrwA4pdFbOonG636UUEHi+WOIldPelRObcpUPaXazF3UkUJQmd6Imb9Xy/
MF6QVwkqgVC+55M2MeXVq7mXe3julLmk0XTLhEvLKbMH7JwLrh3YTyjUsLy+zECvhmuuSjpS76xH
e3NRljmKdkUtZJA/gmXKegiOCRJYP344WoKyYFNloCNdcFchUsb1frvH2FisaleWR58NDTQU1FGy
zFvMZMV3tkzBveEcch6D9XajXjpI3qyjGhP/Dk2bb/Pl4eG7znWbzbyxVVPFtgjLXKAdlGRolH93
BTDrjKVTFDoci+cPGSxs7vwGWxsJczTeJer/HONunOWptEtqDGSvItxfUaAJ1fd3WeSuJNOL4QSy
b9tyKmLhurG/i+D1VP5gqAjHEXSet/vHUbA3sbVEx9XcVFbcOlCfD2UCAKeAu+qNG134ZZ5zx9zv
R4pVM87okci3QV6ystxa2vxzW6OymxytIQ+jtQSmwDtUowf9jISJFeoaShqdkPJ/Z+RvTu4+hlUN
h4J5L6M0Xt+VlLCofl+rvl7jDjzQ5FdBezmTZlXPk4pKD55hNpv5AJJGNGVZU82svRmauP9TaNM8
W1TUcX5iXQ6WQmyDI7r3LX17TYYmLMLy4Wtf+S7zYBqQ96uEqZedVLyHMEKGGuEXi5MpsEnlEIwF
AEY5AkkJVhLf+NdNiSBOhLT4fhPulz+L6qvYldI9P6OWJCpjX1jRRU4H+7lqTVKbsF70SyyrIovh
vv6I4FQCBsuO1R6ccR7ZFFS3Qke+wZiSzQFILyz49G8vZU59wsgoLZ3aJyJK1qlxFiYBpNetMl/j
e1nQBD8GlaXpZ+OV6ID0anA8UowJXnzlibME9ukErsQNZC7Cr5LtLplgx3ZSCFdhKcDT82jy37iu
/5ZBuoo98jhYrxxcLD5AOwkAiUSGoDxoF6tncNHv4UM7N8Q8uMDn6a0zLR/K/y0uNPT/9j79Ajhn
Ot7mTQyyPfKp/6+3cxPKQJ0D8L+h3r9QWBx4+ECxQ0qn+jNNx0j6EsSTpvCWyqc+XMSOQr7hoGPf
OCJTiRp6a1OgrPFtOS8/5K55/wYy6e7BfB9MMmjRzzoDTRlIvHVSQpiGIzNipMFdPdE9Sy+EcSNj
OHAAPhH74lD8hyxxMSscQnmgtOR5B8ePN5/Xi4gP3ZsTyqg8a9URa58MrxUyLfmgCDhqTxNWvmpV
RqnoOTa79Y/YCHIgk7wuaCud2OSHWkD4MCB+zFkZZ80JHoj9m3xGXqvHsWfI4QREsQDpJgnIGU0i
QspWdAs0oYSoegEq66JEJY1nH9xZT0CGHc0KgfNgSblL6+xnGEJvupJX7Kc7ZPtqNWdZUedO3TEm
CzgRp3tnyNSD7crFjxdaw/nhsmw9qR+RsVa0rp4nPNoSEN7jSZqc7Y+cnLqYSSLjzdhMxIa13zaM
IXwSIislRTYfl7Fu920mGTbvVuTVIHi95O0Q8TJIlck22ANHsImgeV3vW8KCP2BNkMJF0f2Cuske
cNTuuYeQ+B3svMkeiXYf2r9fTYO6f7LhQ079uYXlnyQSCuA8S4qvyIc+7iy8SBih3nnkon0x20HB
/inkw6XHgLtLYwZvTe0qDibVZQ7IkQRBCXWnoFsokcKGg+UgQ/elVJM8XmrNrZly1OqoHWwM4LpG
xcDe9vFgzCBhedu4jeLSTjoPI3Whe2BmduXWUhRVGhev9ZAypJrDKZLucJqefDYKXmL1+j20B9U0
7UoXSOyt/QGBuIWBCvXrfDHyJd40B+ffr4PB3sUkMgwBSA8rNpFJ+cBwNqSMDVNGJeVQ+X+jyjFy
WMgHhMgxu/LhA46Z5PNienwDB9LAxVf+lGUoS0VBohPX9mJ/q65Yjsb5oqy7aSrhQfNuF/GMlaZB
TmBKVP7LOLTvSNyuQXfY0jeT6SqDkoAWUFcsv9sLPI6wZ1Giaw1uzlvPpvGV3D7NbJ7Q9+meWlqm
xrPxFw4bZcdH0UZHHcnnMwLV38qfJPMis/zTuq8El2uF85DTM6EM2o/3HnrfTLWb54PdU86BTFwQ
/kyr6GLGCiNfpRS7/qjU4KVI6cDN7cLtpzYISTATXXndOk2Ogm91e6hNOVxnPlCU/utYZCUjOX0K
HrH8SGODIPvS2DYyZlnu0xHKs264MWRpc+JN+YxwWLyhGa2HNV6hmvWsFyoAurUW8NhIw1mcOJJn
cU/hWj2In74L2AuYhTNld0AeBVVtMgUoVCf5tTH2ICWUqgxYULP+hbvkb6+s+lZbUXoCbFgeJR0t
6GsC+LhW4IYqFKikMSpiAsJ0WcQfun5DNrLLialgyGTyIn3jXnSetfNT0NlYV+A3mgHAH3FOmGEy
Z5jznR1wNnJwN48nyE3Nu+DUzCkuArPZt+kf4lQQXyZlNlpu45miZvyUkvMUIWQrma2ectcS+75v
fY3FzfBCti+B1+9yS1Nkkq4v5ad86zZMoIti8jCvSsv2K7wj99mFAZ6g7BWo8xRQHnkXp+klvI8M
YPuDDPoAEtp0pc39hP0JL2KX79FSEkc21n+QlKWmdYEpVNiMWB8RLXAJd9B5udux/pOsojMf5urh
nTQfUsLPkTjfApy6l+B2Jyu2YtHmYe+U4bF4uWa7JSTwGS+XcBde34gwPDc7Tm3KFjj06nBCpPYj
4dy7kSbDhN5XoP3maP2kMhIHNcasNZFAw+vU5Ri6gEZAStrA82YEa8ZtZRcX31lg2lLo2DZq40qw
dxpqZWv7g+FiUG3Ua3hNeB5KiVNGDVFln9jRhw/FX9gP0s4vZE4HzKTRY2BCNjXacl3HdusUfHbH
4Xz1xnY6K+VDB4sUeRP0hos6bH9VDTYssc5HLn3OHvlS8hiX3qoLfvUaYC54COCho5Bdh1UssE9Q
48cgWhYxYzZn/nWDYQzuwFP32KSsWrT/5IWRf5dmqWVI11wxq9B0CdIqT8GZL8GM8eqKgyQHDo/K
2V49rj6azUoMeAkWNkjQ4gbC1UxZgQvpthtinCTnnTdvYGWxAkNxDrUbLMWOoo4n3Is0iDiDQ+cd
zEx58mSkIAqgySb6mtB7CLCeqC1yu+G1Gp8Jt2MsEjdXvySM3FbdyfMMDN4uwm+ozbwUB00b927U
TFPelUqBvWInp5X4UP0WyxF0RjnIyBtWydgcr9e0IIfvno6xZrWjuI9zGvlGBvDjFg4niiIynrjJ
M/Gnh/5fTBNREMkNuOH84LwI2KtyDB2bsIJYZibItgINVbYRAemZZbD8OPkz6A9ae/ivXuh2dqP8
OTu6RKVH7WTpmLntlDq+we9APymwIdoJtXuYWJvKsNHwc8TQ+jm4MxavupJzLW1zW8v7jqoOtIis
1VdwLKHX0TQ1KSCq3T1dh9QjdUGgObHipY4iGh+QMOovMuAlajGneqIvXJjo5cxwi99fg7dvx4mi
BUPAlJL9RQLrE8A6OD/QUR9u2eccmN9RIxlLUi3kkCGVv9RMFrkYhulaLIJ92+fFBcsm2vuqJigu
cButqBr3FVpLXoE3GkKNNSg812gq5HWzIuh9I+w/8evoC6cJJyIjRCFwYP6jJf9ol6o/tDZhpDxV
LgeLN+X+4D0atz/FjiGXPY2PGm90ztXYLxSxuECFn3ZZA9bqusH6jp4XaVX71rILJM38yhJGuP+f
cVPwuSJ93qmbL0+RlGkd7dJ30B+YJSWitlauS7WYFB5pZ04kxyv/MtRaxy7V9HtHmuz01cgOhUo5
0pBthLEVFTgYVQ10q+8oLP4jFK2SA/pLsGrtAgCjm8TziaTaibpirzkzrr8BTGg1lvJl2R0VGh8F
nPCRYbEUpw8D9bN9Ta3WGZQjAyGImzT5j0mP3PJE/qIeVJ7KaizzTk6e+x0cTMzDWqgG1c7T2Tmp
3C8KAQgE+2F3Qem+z1u5hbjIn3vj+7Ikudkdb56tZ8zFU0lZd2gW/G+IuCD9cW+yxoPL0/kweZYG
9ocPTCgV1x8r0AJESilht1jzCmj0t1hSqLw9oONYjmSK+F29KADjoqkVfjDhMuUgo0kHwQdnQ1EN
kHI9BeIjs4W1YFzmu0pDjN0wY1LCWvB7HveXnfquT79D7Mn3L7QF3L2/9uIPPLosaaRjFfA7MboD
KBRN31+RVvd8y66n+SMS6O2413zfQPjcy2jJUB5AcFtsOpOsCEd9deYSfREyDKOqaVYC7u77MyTG
F4xT8MC0pBD9ZcfamrsEZVm+UyFST8ObGdI6vu82FApD/p1O4tUxDkGoOozsHnVMBPJkJFg31H8x
fjxus15xNKMkvAaoJL8Up1Z58HHNgcbqFgK99nFbCv7KNEHqPuy3HRZ7i1ktbc6sHu6deDv6m2wq
YJurEQQmzRujlgguRsBhEUGsahSzwcppiqouWj1M6StfgT72vNOqFFjYmyFKuI386X8tQQh0D9io
Yo0obwyzOUv10CjrKldJ2aPHVuWXYk1VJmqScTWn7PVG9VYTb2472y83st9deEd0pjetMqgXwv3i
Ho7JXe6njMtpW7+tjArale1dYflXmbcB4x9kXBr3Uxd15BhYpEvCsaY4UA9a0dOauMlISenhJZ5j
+uy/HBfgHp86f/BOhlnKR7bC/gdNmHr3TWJJ7sZYBGs0B9a5IrNaC0eVH2/EMC3xtBC7YgmdojZl
6z5YlyuhXoCRpwOLinM5UvNS3V8a7hyOY4xiQF6QzpO7P/NpUYR08BmVpCflzXnj2ZvOJdU+5CuH
5OVZLWGtXTHVpiC0XEmOYwN3ITTIWwWdIcu4QKC0NTsnIjQjRTspLQemrsH+5MaIFgKRs2/BnjdF
V23cOX+Zs9KnYDT3Bwy/60h92BfrXkyw0gUIhNITmmrD1Ii6kVd79pmhB8InZN5CJrqfqZL/9G1a
ZZeBuAfy5S9D05bARD0JjuXKzv72vhEha9lWw5veVQZxhGqpjUI89lYiu5mBGuaxmgyARGp9Fnvv
wHlv35OBaa66EMHIR8Y7elWOE11ryoMOWX0jTx+qM7C4lV+3RMkSuI9Ibj8MGcyzZbi0Pw+DCkgE
VHY93KJwiMUS4Pk4bhQg1zczmVSFDDjm9ZuIl5ULUy8x0nlGbr2IZ7eU7ybF8nEDTyDmSxFXHrLE
LwR/SHKezed4XYuK3MR8bQNHM5L112CFgwSosRDQEjU8d0gZogBt8x3sIAjNQ99DSb1+IOgsKEZE
/Unxm1YdHEh0MJmIwb4HDRoIadM9hd5xLEI+Sr+QXwbM4ZCcfVsOPR+O7o2Oy5giPZjnsKbeJA7R
1RIv6AcUsH0Mkf7udpp+2fwG6FTEqZBRXuk1Qzc2CuJrxp8ZZ/rBKJ7hFJcekv1O0spXG4YB/ys1
mC0aORiTbFcNfJh9Sr3ifUI/Tr3QgBvpwp+doLlLynpXQNQlsAJrDU8qk9kYQbv4swoYPVzUvJAV
Kfh0V0SvfdXrd6D0T40cuGFwvRu2IHUaPxnnmHPfkwBZ+DDlIeekqk4xphEhQaSu7It2soCUNPzm
JhyJNXUyo7UqchZn9fycXkmbZBWhvzoOzM+CyTZQNjNHJugFcrRvfd4irEMt3zP3inMk8mpR9QEH
Ckrt/FrYcXawFbLPBB14WmM5QwVvy5yNGZXYC5r/NKicPYEBO5G+RxKvbIylYlW9WvSe2wMe1z+M
MCtQXA3oRT7TCmogawHcthRKf5hH3WWFT/o7j+CpF4WMRmZGCP2glZ/2oZXE5kNCFvNmHDh8/fNc
Zi4EARtK5Z2PKNYq3QKXb0Xj/mwyT3P+b300t5UFEpO7ftteagGVbIehJAeDtBItCJyrF5ykZCKw
/zoboy0AgowvCFA7CiGLpM0DbzAhFnqMchf0KYVUOsdIvZtodk3oL3vR90m9AHKDP/IJPRbToxmO
Y8bd6XawVeb0GWy5fjmB82cVOfVWXIf4BViS2bpdfxowWibryRiOAuta7xhNdacAsJhcf37fH8Ga
F7DJSa8xkKGFbDH2vihypeda+F0a1UR3Mydh+0S2RBVMJ/Pher0o9I/an56wS2eofbamOtCKS8Ea
FFj2JwIkTeU/5btP+EP3ozfVPjAHDzGAcMNr5Di5cEhh89MIQ7pTa6knitlMt79SUBDHq9KdRRJ0
Wb5juEQrwV4gtT6rlkE3Gvt/27twPrRv1ImQa/Fs4jC0igeGz/xoHYxQqKZb8iVUq6nxWdmDUe1V
D7O8GqS2InllNcIOfi9cAvh1bbxcIZqQ5fCFT9TqiYsRX7TFCuoyL7Kk3pERouXYcGSBXPM9P3AP
jyvAuSdjh4/H7D4AU/FvJ2MCTNAgYVyyVJIZY3wGIiicULMu55Qwp2XSBiLIHAZjAO7ICnjuAaeZ
bHQtpgTF5H6Ts+Dc9NX3M5c2FUprovNrhH+CeMDw3fc8Iv/kmEMWoxLDziFWo/1/9LmFoxSgiZNm
WdjrOdNam7eNDO3IH66zyVMRJIAVTZ4AuwTnint/bvS+TYuSHaz+LT+yK9Jq9DRFlR8k+/zmmng/
JcTHTcC6fhOkyiyqkdgVpJQnIEYmKEUAEpN37iTeqADhw+6xN81QyaJ6aB7J8lSYfHgDpINWStiv
LfinAKJTG8nfmQfDKT+jLHwgZu10n4KoRyRGOZdntJcS3nmYJOsfIPRnc7aQeznhTPXJbGWmG3rH
UJU2pwS7YR/oklyVNT6wocvZJBpKZh0sCHVXVo8hXb2Ws8jr5sdVnewtzZl+w+9y8I/i3SnR4RaZ
8onbftIdIxB3Uq/lUOYNEHF1W0pV/kXc6SOaoo1Xl2ZQ4zSBZTjjGAS/KNIEPFiVQnoPR8KZ+mWX
iCOKCOTgOf+WTI4/C3ElsKD34gSpd6ntvcaHesirO61NsA1yJB+8BzoFPalaup+nDIffesMIkmW8
p/32dvw/i3dHAal6B1QKrAFgfX33LpVGJUsyCH/joFr9IGmU41FiTiG/rEZ03Y1j9hP4RGfFjOoh
HyCkU59QVcZQGJKiaiSN1BSqcRaf1nWRDaEKKyGvoUAEo53cuGoRk1vzs9AU4FrwaEGYoiLsucon
BEjwXOKND5jLgmo832rl+dERHR5xu7T+4KGKgOJ7VklfDV90WSAIuz1FOIfqVfdvQOiCGZ1Qf9x0
EMMNmBfy539v5xfLqCCHd02TkIO9lT1HVjFYC/uJPq3XxDxgOahzemEJDiMjWYSglk9swg4/vLFw
8TDFIVVoicXEN8TuPNTmBXmX0/vNHetwYybiFTfYUBCFwYlYZ+yVrH7nZvUVHczkOLUpE+EKuAd7
xi01gtYEjR5rylVvmUqc9azRt8FJM8WU+MRTd/bJ69tLkVN3HV3Tr+Ek/XzsflnBOO9n0LXQirAF
PU0M60mXMgJ0qs/dsQrQtc6jMycuD0CAX0VeC6VUm166FEFSmhFEedMi9Rj7Km70BLF9os7TqxCR
2c3HWyQ3oOADjWeyLOt3BQaRVSR1F2OcdjWFP02FnJYlIK9sJA0eYccAVoe+tXXBvfEUY3iNx53Q
3pSD8/w/CijD29TrxE5UqX5HZzaCfnDkcmO8oWXlx2oxrLtG07shNb8V9z05QpJ92+EK/BpoPe9E
rUOOoosKtSM9vTW0YoTQZ9fNcfJfdHEodiTYkkjRQiyGws1beScEoelcVuvOALGSwaot5SLkx3eS
Vh6mDHEYONsWrpkbdB6dxAYaxol3AoHKdT1njFYk0vY39tg33kmjjjFWLLV1Kv+O88aNCdV+t59S
bWgBC784yu++i8pgWY8qeU6hpjG8MsA25rpoTKstFtL3wvWc37k5fqRSoXumH/guid8K/qMukh9J
BIHDPr8BlWjRALt4Z6K3eeMNN/pmeN/wheRBDyzl1yMzc1Wew/k1HnwTAwY4UosRftYVAxRi5EVX
P8HwLdfG7xKQwMPkCpdgGcKKTYthChC1JUgjRxETaiyZInmyDbcIT/lnA45X0dFK9IGluMMiNBJM
xRjwQR9iXroS+WUVJZnInpd595doia6JW5FLGKHG3vGGZbyKPVNmauxKkSqqsTOcDgzZABSlykXP
ky8Yfj2a4jOl0hNKodG73L6h9dJ50Qq5vBIEjHgQXzGHHzogDwgKKaEsUJX9guSxrvUclO/arsTP
UaVXknsdHL0s/HQBLmimVu48+dfULb33zgeiaYLiV2XrS/icKjtq8LvkAqsri+EXYX8taUrJF8Im
iF/UO1DFhXW4UmPxwpsMykQLZDEmDHgST/8zhrgJarLLNezCVFF0IlH3fmuiLv2T6uj9cFw+J0VK
JxEXl7ESEvQE8BeHXcz39zm3OyuI3uQuf01DvfLwjGzW04uYpx12F8HWqDVuxm1ZH/riOwywzSNC
Jfl1p45TIGHHtweiRVmbYz7TVI7wOmxzQGwDGAN0SbtiULQpLqU5GYULp7jxk6qgdCXR3pOIV7el
TDaiAEUKGvfS1pKglCVZFiKJ1fvJ7Pzg4gMcS0D7miHFH39Q6GJIbNWdM2ZXZ5U394dJ/oCXfhbK
hRxtBNqcUUnlxSPN7E3ouOkpxMS+MI+bRakPmsRc6Prlm48q/Fkn7/njeQR6fmowZaMP7R9doxy0
dDsJCbAxO06ORmmWCXJFFNEOVBbwZdRgCwGw8654Qp/5ZfJG6y7ZBydefUXu9VkMY2KkQVWjG/yh
FiCgOe9spogcMd8VNovHB51VeDVqHf3tuKPBpeRpZaUbzlXZb+Qzfre2+7vPkGnPPBfGmCJnVXWN
63bqOCWyMuR0roeWXVEkcgsBYBVJ9plDclYsydT8wGL6tx16EH4+CF7f0szAeQVZdQ3IhEvWdmst
V2yJCAgHMxdyaGqzJdmTk2JtYPa7WglUqvb4LORE//vfpwxvHTv+NZGRCVA7TiKgx1HfQ7FpMH6u
Bokh1yyJWDYj1EK7rVvLMRs2RaTbn7WFPsc9zzHchTxyeXzboJPO85z4ivil56YWcYsW6HHkQIP2
dJLIb0YUL3ZukU/qQ1NHCtLATwu5Hab1e6GwvSCv1WOrfdNGARxCCHV57Q09niQqbqv6J9vCPLoa
PunNCXuzDBMshH6X4G3KWJWHuJoA+ZMhfSJFGRDrR8Etkbd+LASHW9ISjKmi9K+dSu4mIZYxC9E4
Keqy/wLASSivyehrZNoRvN42DpMJNFVSSDBfNIbkBe3S8YuyF1rS/L/rknocbH2s0zgcRZj+j/EQ
cy1uUWOiDXuH8tiT4pgxNkrIQ1vEn9A49ifRkCt+WaL62O5haFb6rAMy7ZpB3ZEZiCv9dUPDQWCK
W611gLlPnoYNC9wmB68Sz8EwDaFl/n8u3nJnaED012d5XlgJdVPwfEUhcmGwyUK6Bf2G6aB3oLPj
ks32fr30sBqm16QKzoxwkOu5chgWabsPK0/i6dQ7Rx4w1sI43CKbu7plntyT3oajU1J1CsGi/bBS
mx5lHBSghcgXeACS3tMY1OYP9wjUzX9udbz4pIE8bIzFyGaZCFx7474l76Od8LrwWA/5Ze8/XNSG
3ObfSenu4dz4fxO57XnoIcyuTkOYR2b7w1gsNBZ21uq3T3N33jUriewUwWnyviEcbuIP6V99gqK2
2T0ib6SawUMGwrrOPn9EUIzKLdq9RPwVcTRtifP9uaGrISGcSt6HCdKVvO+9EfHx/1C7fl1iFtJn
E1zmFdhuCw1+9MftwTBAH4nPzFf3f9+IXgwthuqOVYRJtKZMJhRHDECm8RH/GCV9pDr1v1uhcONN
0bQzYhsbB17C0VMQOVtm6nYuaHWsVA3WokSK/7LIoobkFL9eLQuaZVK6bzJydCuDWHLMTcP6RXxt
uHarU7FksqTAAc36FgRm+WHMVx5i3Gy4V6atpgf+QVYHAhMxlaPlYeYDQe+wu1utiNt4YcJKUg0Z
dWqgdZue7ivy2UgEBgEHBqXNUsfouz5qAT5iZMhYdhM8DIBzTjkmBaRw9ya8c+Z7xUpVBkPzqt/i
LGy3vtIw/Ff6jEnb81cV1nM5au0SNRHh33wxSrqxibXxAz6d1DU0WSHz1T90WA6F4B36a1Gx61QX
UGDerRpOhE1sSb5vf52dh2mlqpsPGGtoAiUUgfj96WhXBYfmtI6AvT/HCrpqL25ACRLL61izHfd6
m4VsSdPFVdZN+byftPhVKAAVNlJjIGYKwOO3l6qXrODdra/rfyoZCtdY0eGdnE7QMTQ1cWaDfByJ
H/WCj4KzvJBiiD9tRasxk7+rnl0XX7JEizxKoy90sbUwXP2K2HiIism4JscMl6bjb4Xm2ceAJT9h
HFz5zNRY2Ge8wPbEZMQ+4WUIgtImEpGwnSgV4Dbjiwz5TDWLp47XPsNLgTjl34Hh/mvAIXCNeHIw
gcPufZmmUSo7wtQ9hjwlYdsxeGJOaWe0bEiJ8TUg+g5HspICR+1At+4J22R7lZSVygReznA6gihh
F5ZDB3DUe/VtCInM6iBAof/JwoGmDXz+7r45uI1SX1CNifff6nqeLvoFpvlZ4pR8z5nRJY1cqG3E
7OMlvd5S86yPaor0qWlIHDd43ZUyBJCs2r+U1ihx9L5JR6r4YmqJC+aw8grhFSyV5B84cho+k5Dm
eArDqEcc3s1UQZjP0GsQKqg8+2wmlGm+3j2JZJJK5F5QXd9mhbhF4WhKrzVsqgTIWSBWKBzeL8FF
G3YI462g5QltYVDNXdccUa8MPvH6qvVZPljayREScsrIS+wXo8DODrHOFPxIb7E7w05rKXYYLuJ6
2pk9sFQbRIcGaLh2XtdDSLgTFyN0USa7O3rT5fPvnoCKQ7gKcypcYbSSItKSbKt0nS6h4BlKkei1
NpCenwCkC9TLEWnVEicKMSAZpBff3EmPfd7ynL3xzzXaBpY5nQTzMPKCZkZLyzZ6aGbboWynQANF
+oNcVpASlCoYuWwHuqRHfixhqMrrpAm5sa+Zic9xqp5hLBYJhvbfXab3vmfzCXr2VgdlI+NW+BVI
iC5h3WVnsN5htZ3XG2UjzVxO5mEFByARxAJyiOWyGHGiltYUjNPBGwyOVZOgh+mrhrYUrAr06duD
hUEZtIcV9vlABQ2EvVrqmJmnYo1CAuhBjbXtMoCCACB/Yfet12BfTiPwO9L/3qCM2pia9+NML0at
xbQHy1UdnxaLSEO/uMCAuxBQhs8Ab/cm/p0WbPaVJUFPQp50WMF9vpH5PLPllGVrFnbjqao5B3dB
0Hh2LKKgkJOlFdjxvCWq/pRMfuymECaJQl7ghWxMe/aDMikQFVFbK3+FYRLV0B976o3CU3j0cE92
qdGyryqtDeuClpAlKkpZznN5h/nd36hTX+Uj22XK7mJo+mdrrJ2KZIzPcIZxTag9xi1AUte+wK/l
UijafQepA/oos/cbWOdJvTJAz2V9CTejhMm3TfUheDu0LoI0C/e/MFW9GcJgej4sSwRO6+9n41/t
ApXlmdojA4Pbk7eBqt+9nTxsviZtLHlByFZhoRQjW0JxrQmUUAA9UvRHkudiHDecTEueYo7/O2nB
/y08dNX0gxMKxK+sWjfgR3e9NC1uDjPtfqRCTv7X89f3+SmvWnyK3hkMext8p5ER8xknTO9Q0gCM
7MEW8p5pbs+WcOcdiv1pbDQStBSDHP5kPllBqRc0RDIFpbvgS98/NuhGP2nnLxF45+Y+SVmm9384
laFKHRKl87L9N6SRpbt5Ptu+JT5FAt37qbK0TfP2U7eLOPn1pl5p3Jqep/rNORZy/RF1x82lXcCn
SRimRDId4bibrrQtvk+nIrHhZjBo/GSQx3WGDtE4g64ovFxvgD7tQDf6+NmReBoybghICEhFF4vF
EVGz19Rnf0B+snHpDw3N8x7GdRCwUMBBitv8A0asKLNr95OtJ6p3gT5HlxvK4Ak7LkrFcAXtD/6x
V//VzAVjZkU7pNT81OVDXCgz4gVAt/bXWBPSfK2JZ1WDuOU3ShypxRbK79WwIGIjzbJKWg61Nv5P
Y6EOsNrWFOIf+BTKdLPaCwaBLXWZfNgrhFU7as3f5ecSiSZC0gbkymnXHkg0G4waFs9avDY0GoL8
sRnRhTtQLg7vK3C4mXM3rQEPo0pP9rcJcbxl4zV+fgemlLFtOXVu22TAjn9+ivVr/Sx6nGQgvvk7
/zVHTtPfEaLYHGoOH8UTsXKYqBWOVZMX+IWLibcb7bysUqPjyOeRWATDHBSqYJCqYno8IA+F30wl
O5c/cCNoC2rAybENoNGdRXFSIzGqEaTweoxO8KDELrvIRAhNenw+YVBop6D5BM5iJraAPy2iwxwC
rpPTvlChRdQNEJ3rqECNU5qkT4RSqSNb9dFWdo5fNcNJOPGomnR/jVaeKsDgFKW+3kUrkeTwc8xL
Ef1mkdCXotplQ5TnkjxnLbgQWqm2yfAZqMaP7+GQJjKwIrwyv4n2W6hBHYsnYcFLqEjTsuR6jEeJ
2uH2F1bsmYXtgsEonyrcGOKHli3fGjXLV6pL33GtrxaaY2TQv8d7NaQWFz6ifdbDh82OZLRu2SGn
UjCOMrd9aWV3dSuvp3ka7XdVmKPw76kgtC1LdQAP3zQauEu6qP71gjolozPCFECp9kg3CsWveyMf
rdIWWUtqFSTjPA4mrASw4A3dlgWPjzPb+fWO+DoHhzMJt9u2l7smKXovTvvSHGKn+S9zU5v7/R4t
WUhpJZtty/z/0HILFWgBdUoRQaUyUe7iIPcroCkYYhwTS209YdbToKWrsScnq0kKn+a00z8i7lHm
DYtfza1M5er7h7vT2IuB2n0rCkzhcBsCeZE6w76TzGqCWJMMe/rjALulge6Nfr8gMz9r1q22xisU
xUjpJuoWyQdyTeLUZ3SMhmgSKSSS5Pw/P9maTao2jJk6hLSwxZ6gvIharo9UOEogyOhh7jrk1Tg/
yqXIybjsv5YwDLGGej6FUrSy5oPAroGlxF3XZ02TdiRiLADPvY4/Vuizd+0a4Kk+7I+A6SdWIHwP
HB+bNum/ebxNOXs7S4bdirD2VJ6LA8uMUVyILafvPwEljI6+J8TVm33i8CspFitrn/zalSL0lq5e
THOgWux483YSWqQguFM2XPnIwxnKXvxMccFI9jdjRQLMH7BOLp0RS/DlqK8bQRZ6JUD0VktP2Aws
EmatTQaqGRqWdd2KYiEF1ghQE5aNlkFzGhjn2WGDQNfd6AE4WV9FOoH7NB1AX4tmQus2A6iLjqnO
5MK7Gh2qvJOhOlBCVKb/4k7NUzJkFR1fBM9eqF1tQ7rMDK3+Ue1OTZllSRzkR9ke3qnEwI2xDcPS
btkHg9b8rBsDHRZrWRPUb5u7Uvzf+qi/02TcY26J+4l08Db2s+rcItKwJia7uJ5FkqKj3jKisTfi
d4/kaIHRpD/OR9w/h/4O6D4EZrNmRP1UVxsMLv+CHv3mPTxGYyd86TRdYgd5D97YPx+SjMcqhGua
Bn7iQw/nUU9sz3IPBPCS952/k+kSGKwELnSv9Ty3Lh0iNXL8MjkyFgD5Y88IEOqkw0IA1QfzY7Ms
vwrYV69NzyoinOxgOn6OseQ5Fr07Jdp+pEAZKVtJbk6t6YotXPOOdDnyX/p8G5DcwVLU3u/HbzlB
gwtYUQ/w0fzeMRBdrecZzQ1MHob06QwaH5HWXE6mWHfxsIBpfiGsaUjfdwOPDfxpIhOeFix7Nk0L
a5POXqvtVZd/v+v6NkgM2ENh7t6LCTuYqwWhiBt3MA0Em2UlAiofZGl+x0oo3e7Oa7gjIXQu8LbG
SbIfrHJfR62Ktw5C7hj0SiETwf0tW+se4n9jmrgmZaHGoVf1V1PGM5lAxkkvXFsrEgd6fMzrG+Ka
vXq3pcPrf5nlWHLEznfwA3pxWPdTU/S55FS1RIUD9h63xIIKgRXtoj+zhJEAioIn/hCPhDtbMuLt
SRCXhE4awJHZ3YCcZCzyh6aCI+wBE6HTB3qmoO57qAZ5VUIaIV22qRjcngI+1zthrjv9+uZoP1hU
zHJ3uuvqGjdPDIosSrZGthMw/WrMiNJV1/+H0DIsj78LGcypaaQzRBg4/padSBCgNmflD5S8uYax
OJv8W/gSZWL68krwQPaoU0kP4yIpLYu0Mv4DS5JUMbf1h6TZM96HUuwzJAHvoQAwS9G7AZf+qsNk
1lckGz7Jv1iFkCsR5lcPm3oCixg2Kgc63CNyhzLtb0y8yHqXRToFwz50AivP+JecRh6tBHHNsR5M
W2sLOCJ0vyNizNEmcRL1aVmcL4xr8ec1kPmlcmyo/HxRMIjx2xpjMlrBQ0CxdKDy2clJ6mJ/TnCL
xDG966ad0tTLITDDng5KG8zvaGyMo617gCgEpM4J34F+h165qLpsHZQzbj+oxKNWvEV37GwWOi2W
8htxcygAv97MFt5YjgbL6QftpmpYTGhx5DzinXueKYnVUgNtitDlZw6bhm2ijG5E30GcuXWPXwUl
JF6NLyev1Thr58E/f76OCQEWyhUK/uUZ0QA9cr0d3wN+jGbhSw5AERu80i59fXd7fmfQB3yFtRn6
Vou6aZtKfNuMlvYSZIASVAB/jbJlrR4NvxkG7kSVZjV9iyG8784S6nhGX8gw5IWbXA8J7qQFFjZK
Uc17feqlVsMSCfbM9OZe0BE/a2RqSz0ZlnmUNha9R1huJpD5xVg5sn1yNYyLVFdZeHc9Q0r7Rips
pTv/wXMPYZeTDWdepPaCgyYpXVhEk7H1e3waUeVzGTv4gzWrJvIahLvtBpJsMZg/bLs1/g6uhHQA
OUza9QN6VUB4B374cVhHZ1ZqNBAtEBDkak/YUYQA8trbRpn3Gcsa2SOy6Y8/A6ZI7PF982UilJzs
0ADGJSz8R4hPTZKmitKkibVzMQXf9YGTQEPz+LxVvS+73+9nl3TPHpUZvgO6RpLL8ou6WibB1+i3
+kxD1U+b3ldE0iSa8vxnL6tkfZJBcmb1isttSyZIsS3qZJylcdThE761CMeAyV2DPvqkQX3lgd7H
KB+B0jX1ex5ojbCI2fPfe74P2FckfJxg0SKv7PiLP+SkL59rITgRTQNii3vA5luzgZ9BPAXwSdYr
m6IfyzUxaFfRyZ6hFKVJ4UpTOGb6mDO8EP0mTgINqzHvOyY6SS8r2kp3paqvL/uiWTzdyKL/FMOx
nrfEWL0EnbotP1DboXesNVs1UfJKlMiGwXuC0V5RtOBpVsxYaobDoHOiYOO751VHwmV6vnYFQroE
yu4tWptAkzHOBgAuJKYPOxb4CeuiuikIxsXgRGQqD7owfF7WmwDzbC/GqeLrKdzf0K/8+u+ns7X1
/8zk7ciDOpTP7ugTco6jm/FVD2uTn8fqJCQ8sjePE3DNi4biEs/dDW1DLDgLj6RD2ye9kvkINk75
obvK1oTxssKDLpAgprjr/XMW/1xnDIuETDs6HWO9r0elio+f4jUvLyALl3v0kDvLdYc2ivFCOK+x
Y2dDz5/tglBhxYDvSa5+YjsRrFEgJmvTZgCc2erg80Cw5POkpyGl2+VWS9NsjmRYYtz/bzXYaghu
0QoWFdL4utetHJnaEDVfrDIvo0NAyGxg56xyl4ROKL39ZTDrjLFbgA6MG5Zl0a2/FRzlU6pkHjwJ
21qNXfTZveWZ5dgTi39UMUJGGvm+MdMHTr1RxlDJRLMaXwvVY++17PN9L1cjp0tieUp7xP8HgWi3
3DSTgiLe/6X15rix6W4wUf3oAFKOCu3gBk+uYiOQz9nG2QbdxtOwuz86gsm45nBPcPOvaOqZyecr
F4YGSMzviyk8YB6nDX0YEDEbryqQJTe8AqOl3GkidSGUog1IQl3mBLi/dncy3tsi4FiCUJbkDpXN
SkN9xgxRYwQJL/3c0SKJ7LszUAfDO0O38hlODRxsm7GMiqbsOWrxSJCpqJwvMf1v27qTEZtziC69
mqtpsZJ/o5bWznqx6LWKVydycByUIhW2hP9rhinUZo/S11tYzMCNXQV/ox4BIMb9LFPxvWpft0YN
LcK7bsPDQbmcBk8Lr5owLVBYSXOEqIVAugXKzzXYddXWTe1PLP5qMDDna3M9pvpl3IeJ/EtM1nd+
g0dRl2enPPoISphCUr3a//GQzdWRnKqe/uVYueLadupqbu9IxDVN8Lszn3Gu4xVPGq9f2Bn3T2Gp
PzJwqAw97vVmOAnxd6u2R92WZsdCbkK2kalg1kipoboYZg2ucFIf7bSWMCFILUpQBlRad0xz/+rS
ztWKKtUa5tCbcQiWzhDElRwBbAJuSdBr1ECOIC1Eudg1xeprsTKyyD//6NDDIg7h+MoMFy/nuO5o
QR8OUAepTdYKcA53Q7j76ko2z6tW1F5tgbKlt20sMr7S/KcI1dNfY5XLoas8d4yIJFkFia1gTgtr
KUOxKqjgqmzob73uwOsMqk29E9w1Vpe757UnzokW2z7OcSiMdCV24v/J3w0NFnGXrqLtf9WkNiDs
muY/2Npp3vkDlyCy0qUZzexepcu1p1rPsPKvs5EO4yM8xe4qn4kbF8Xd2U0S+Xq5NVFWnS612/Bx
xxJVIHgZnXCKAh4oOTvZ9YHnt4DjWgzlyE5we/8uiPWYXRPU9jCPs1WEdiTURzox9jrI977rTs8I
MTlLR+eODzhsy/wJGHjeK08U17eG8D4H0ttySY67hdftJaY8Hcy66ZLNbOk67AIw/mK9mNRH+F1Q
A9LSGJc9kZN6YwKBQI0B3FHHau7KuIiNyonfsO1pUA1NTj83noajGokc/+B3jQalVFD6kdwcqmpj
59I8M3B+1kWLakiV8keQfa7SgdsGqC/EIct1zOoRCV5f8N4XH43D1JENqQ00OFZSLfbbJVnAYBrc
6gWPE/aWUj/IDXsg/1wz9jl/hb1dz+4dY0A+xGkST1+kwsomj/DSWK1YDOQqLM+v3nMDDaFuUJoZ
lLHDJQWbiPu0uNnA6/z9CCroWC2rg06B6ZQiRWefVYGkPXZ+Dg+Q4uSQw9yiFYt7K3m8kX1/RyL+
LBwBNCpvn8+fhnTtAji5+aCNaItdh88r/wdv0d2G3iMZn3xpQZ/xQJ+Zv9TiEu6F16TsQgqjKoDb
Ckdq75zX3Q+I/iUHhKI+OVN1ngzdJeF2kwIu0XujmLE4rRpcXqYR+KpuA4x44SAzGDj0NN7Kaj8Z
mjy7ASLQ6xHt3crw48gdvxSl3GQpflMoSxY+lHjIsFMWVjQvy/RAjFXYf0311Yw8Wq5m5dPZL+o8
3ge7L9RrJ9KlTg+QQeiBqRqKMrpBstwwmfZCnXOZYsiKdUd8TxsVXnJJdo3l6TWQP3g2PfNjvuT3
CaUQA7dNjEZ/nBrYb6d3UWGTgI3YsZ+gQj4HIJ0Z+5flbpSqHbj6nQoyNrGTzyh2WIazjWMYby2F
1+Ul9Ds7Eh7fNkQd/jp3XKr4fXfZjY999JUXc2WNYFAlb1AAFZNn1+eqLpcCOrOanW8kpNdq9W5a
t4LNxQhKVJNFVrBgMLUkV4G33jidIxdO2NAxKKb0eZh4HomwqRmZM3U8gqSW5YCs6tIX5tDgYAri
OAhQTvzRXsyIzUUj6xNzfINGRt8PnzcunfLWnXTKS/YI+XzRTdp8vW1uLTv1Bcd0Lvb1ZbwxGpxN
fOjBzWOgK7/41HGfW1K+DYAfB+AYp3QRZCykaA6AY7mrEL8gm8BXSXicZFD2O7O3wZX5Mgi5FAiG
PevpYr66eyrVaHqHuAFtVyKUBYgI+q7mOgt2VQt62yPNXMunZjcZNEvatST74h4bc0JL5jh+iyac
E+r171gzTiWzZHWJw8ENjrQUSPOoEky53l3iYpp8xAOQNRhiLY5SMxw/gxKaNLdmYjM/kD6Q/Yi+
zFaQr6wUua5BAhH9w4HW1T3V/OvZ4lLcwcUfXXLloH5zb69ymmgCxsiFm+3OLiuADE8tg4fMrcEY
wWEDDYzkdZhiIUJ/ALq21/HLS0jRc7pMvbf5SV3oyXQLDD0QfERMHbjOvKH+Et3EKA38aRfOPqfF
tQf40COmAl8A/8/PsIHt061SZzwF5n2ZrNTJ4dpLU8Jwen1+AZdPJkm1wX9RTT4Q1YrUJrdonUTA
Jw9Nc5GThSVm7eaUeTgOZnT4YzAjs/xlUUDY/TX1cIQ/PSW16U1g2WWw3AWYrgcUSDxuC+rFEAt5
fWbhfZ6UWNVlpObFble5cIOqiB1giHJ6qbdRebD4Xb9kHvT2rn0BYnvW6f6yhSjGUCyp0EvbFCoW
wpFAtpJGIIyXHk1PYGQ/Xd3dvfNSl+ClNqMStKJrRh7CBWpISzfRMTxpr714GON/qGSMNVXmr1EL
2rEyD8AHCu0ZFgCw+H/8+XpT5ylSEOsEUGFCOwzV8P+8UhTeENLPXJTo2PrwiYe0ykD/9PyV+l2J
eQY7zSYB5tAyN3TB9w3XvOqegRXLT0i/EGoJg/Jr1o8wZNe6kzWDarlC0++Wf4wynZhjsj0ksDje
gR5l6eNKqYs8ynOP35jdrDw3Yl4Kx+Yk3AVs28WeslApeezMerC2uAgQMxW4DKH2HScnTMkZoU2W
lcDpy0wL/23LknWjWMIR4AyUZtLbmAfJXugCI2DOES+f2FoytCVp80hH0MDh2iKZA0X1ZnieHG7w
4G5/WHi31umxd4GutKp3C/+z6j20W6PTqSIICAw6ro/p6yTkbkVg9ZrRTg1foT59TqSsyRV/crV6
R+03Rytx0N3trcUhL+GHlEcHFJAn6prqXsaqwUDAxu6QosuyrlmpaOUPoJDEp5jOmGCC3z+lhMYf
WwpQ81Q6OO0u0Ip/S7sJi77bJuiv2N/RB1YaEnR6omvtBqKunjdnItry0DuNj5pvwQdKLN4a3oRp
aeS5hYVCZTmeCFHu/BusvuYyT6RlcuAM/enbXfwED5/PKdMHe2pezL9TCmf3F67OdzYriUS8NDHp
FO4f3MUhBz4pOrmVx7kWxCr6GhocUi7Rzf6T04RARqcqPGoh8YewPhW2ka7gNWXKAUi8P1xVb+92
CrLkImn9hGZJ+reip+Wz3S/bIPWNOGie71wurd019ox3j8Cr0TwozuESOW3l3nJ2PL8Grq1Ucvt2
72dRsYTnoHVCQQtykU0bwAe4n2+PGZAISLPjoBdLgEQrleNaxVWi7jzVhir530BUhz/aN3MzCwSj
oLGil98FP2wH7P8LBSi9oqlb+RbYs6/RxYnrp2EBUsqdmRTFSEc3d/mw3CfJnQq6A2zOKZ1fxL8c
4hncdTIoO+ILTcGbWM0n3Y7MhyjjK9yELNSBy2wYTgVOD6F7V5/Tmeqc+Jqbng2MRiQDDjoG+1TP
CzJJe1luIhEcPCVHYsUeK9HFECrtMp3AV2cT+gWkcqOkYnaU360uxk1kCMoEvdoHrJr3Xh5ytRkI
EMDiJ/ENKpniqK497TDKrgNJEbtN9c26ve351Y21YwijRdcO99nb/bCmKUkuADq/XAQhsqBXn5zh
DsDlAvDMUEaL0uqBUAazeSm8KHlSPOmk3Mwo4dITGryXjfumLApvTMlIalFKftHPTtfR5ibouK7i
+AwB0N6KN/YMSZBnzz9OkjA8RebpUaw47PlCDM+5JErw2JirC4iH6B17o6PsYhl9YJKpPNQExvSp
l7+nctKb+iumek2FIdvs3S36lop47wzBWcX8qlWG8WN4xYH6DN4fpi/nutAj4ekqvre2IlvRZmGi
4PdQqpFprlncvfHcY7bTrK1cqzDIZNTh/15blk+fig4smnOwqE/g2Ci5v2FgTe7P7wW9+452Xuf4
PRk51PufvCiyiHJTNyxVJxMBLdr5LeHFLDBATpVRTwfQzEP16PlFnzf4C3AjwkxVQ0VWiEIG8F32
rCf7u4GgPCehKZmUu8jud4ToU6rQQEXoOJd8W07RXOSNDErU6QfvVxN1XVW0PqwrCvrenyp+ZvuT
rqtbb4zcNBJw7EXmbDekRmjmQHLKqH4Nsf3eYghvNfkUsIQY+Kf4na8VXvH9gfmJAn6hmMesEwUd
9KNxnF2GuE7YXd23ZZQplH5KdII2BT+85PnC4bFpwERfWoWt+lJkK/i5UMdvmKT23/ruQMUKLBoU
Oq9+u4vqPGgWx/OB1jR+QSvTmgAexOyhTEzr7Q3eHKRgQ81bgUTl0wD4jdyMVngSuzWruagoD+GC
eFOTsb1Bs8T932gZ+NIAw3r4xShF6YdWjlNasBTQq9Lvua5EhSjrbefanlvNGPY8bN0I57H8AMRF
tD/JDgMPlIZ0CqYOy+lJYlxjAYwfqYHTidsKpt9pRO7lZOa4uicEnHNbiizDy7b9MxNmheVcwIYE
UUhMLI4lbN6K1ynKOzLTiN9Ev+NA5bXgA9EbkvhRSXovsHrPxdmP0RtsYFpDi8yDQh0mWy3l9iQF
WuuuOcLcmK0Fdj2oUvX7+++lXtfGm+3AwM5ZfOuiU9ma/tbQ0ycp/1n63BZmVDV4BM/sNxVSz54+
y0/VK+wrAU6ax99jH6knFjt+iD5M/GjgU296jmlZS0FA+SLmyX2VjNN/7vqNakBTqrPc3WkhxfFl
MFYh+E/naCUkZoKr6JHJVpk0mW8F1OYkUtfZPViFz2bhZgEvoSVlLeeVBA+TRvBW4hywgCxNU2P8
eq2snnrkb8XkQLlfbTDxnu8T52/Smrq4b+I/T4kVeFHhWuTmsukjs8d0jJqDMTERmbOYsA+/Rjd8
/OYDXJQ3rZvC+h/O5Iodaf7QXPh0AyltI8ufXOUbt/idNp9AxbJnmw+G6C2Bc35v3zgyA/RRkKK6
yNYHbuSr/gt9NrqM3A2a7diPuU9PILW4kLz8/HoGhhrDgnCQyhhp1xD0hBp1Q/Rh9H0LkSWlHuiK
DakhMpWrlZHGMNY6p+4Q+hKqcvIcMyrKG0ZYqLjyKZ+FNcf8DvOE+9kirhSXatL2iXAsgqTMWEpY
qGgxL94jbT0yQR+DEV0j9ihsZh+5P9H1zWX/bPaLl5whe9/xiVVBa+NRGMSS2XjdVmXiGe4kBpn2
c0JtS3+pSeOcvktpFdfCHtjIA82cEAn3wDBZqLx6YBWH+s/CWSc9JoFz7En3tTwqi2NvpmmVFmBB
1wxX0WunBBoekEoW2ahtlK6Zqi+4K67EhaL96vCD0Y+NOGRHxgM4EGGJy5mwz0dM4Ada6fZnsw0Z
hHAU78JlMlDGG2rfoguDcWQFcww88WoieJzB2yyVM8E4b6Yn9u7bCEsSwG/N9b0c5ue9/hNTAzs+
ZeWlC0bi6m8Q9GZjC6ryHnJnAFQwtv4bYDxtOZwuY7I1FZfonD3KmimXyCt1sxdvSUSAtwjB2F88
7hjClHgAqQSCOVxUUKHRBISobAGeZtSOiP4D9hIII13/3PVvs3G2g1KpVeU5LOtsYHvmVTJxN/5k
cZknlPBdguOjEojYcX8R01gP/hLZ8UYnKZ75Gu4gmrwdUtL4Wj5TpOeTWaumyUESzEaTLJLx/Bsj
GekUboRXpTyh8BN+eIdISkYRQkZjPS2vDU2lxGh7KkN3jLE7RMyn3SJGN7GCfQVpuukkKBIJZAvU
RPC6oblVK1I+369lqZ4BN2daMxJJSbAhaz02ldOmdFchlLBjb+wKXYx6ylEOJK3uVrypL239X3MK
E9KoVau7hDW2IVanXGHJFDA0BwOF3cABu5gvfS63qRedwsyaF/YUk0f5rkWgpB97hMIU9J+IgpuR
+1BGEIMnMd0jICR9fiNLYSfQq69BXOSS+qD1K8XswieVvo4j2Xwt6oVfa4SuxuiC0M11mS5ETlmZ
vnOM1WcHE/c0/qW6B8PgN0TMJUw460L4nftNRasbnD3q7fX06hUCQQy+RdPsOGRFjT6XQ8CTbGJf
T3aP9JdLnOVad2nOOPAEXT7S761ELAo6iddXfZL6g/L5D1DnynXTnqQkMXeWoqFex3sM+AJ3yaLX
bOB/ze2iqn5eY2JyqsrDtYs8KWgPAGWtxRXiaPIIZubqk84N3fRP7kpO48re4O5bxMK+4iU5eP0w
TN40427JPDJ/e4xtM2cYiT2X22oqaUUvD45dtTdHO9Omx4uq8TFancgQller9SufOq1k6WPePEvB
UbqjTKCyAx8VONuwBgHp7whoTiqqOOUgpszS8YTU6BZ/BQXzDK5ABL6sW/9hoI5VdYljNRhvRfxN
MkKl2mxQUG2ER57b5rK2bEWf7ag/0ECOQD2rTSjwYNtSEqN+SBRPPfsBtQLuHAlZx3AaFOcJ+S1z
RIOCHNCV4uIK1jlEaAHoJ7tPUd/vfre1tiL4eC41SaQ/TeCHdmAfr96hMjEcWXut9aWHBPgQFLf7
yDRQSC82TiuCLYCmvD1BuL8mBewgg6hatgA/MYxv+4dzbuOF5Z3TIf4Bf/PFpTJhu03/0GQ+I4lQ
rYbcC7L/zK90dmAvn/YTkynzbu1R9O6I0VUqi8bjWJXcL6upXYlETC0gM19wBMYRPevKUkkK8taa
AvnzeEX8H6HpIaVStU5uCxHIhHj8uBXCabH8YASQRxNfWugaxRflwAHIwPvANQMzREYwB6v4B5YY
0iyT0XqPuYkuc7Zpa36VSsRxgz6LVIIaYrsjg4hQJHBeV9dI03VeHOizvVzvkhhyfpL3P3lyhzmt
WJ+p5PnebMpGtMQ562ej6bFcWiZcMeCK/2+gNxWuCM54xr69AA8FgtnFFwUmFBtYtBBE58xuuKEh
lzDfXzNWWSkpRN1m0Yxck8A9eb3vPdHzxQAsTSh9Huv/MN93mkzEDvgCmV8S37QK61USR6EhCX9x
s2WDIRbebIMRuPwNkpkhTlvu3iPM4gdkfMIt9pwDgHJTK3aGYRi3ZI4Ybka1+5r7Zz29zP2yVe8h
kUR0cw2zfOhXu6JWnoyfnfUmFB1XUlnS96bVy6hO41cUJmL1dI1YgcgWjT/6sVPDPa8YD+aKpgYU
jHoM4bUNMAnQ4tMX02j+Ck7j6v1x0lfzb7EIhv9aElFjeoGxDG4+C0qSuT9tEn86K8KavQvOkVPU
oyVwF2XB3WsHhQbmTCFxIf8dCDRJfGJy2gtERu8xH1/VYwo+fe4kNABJAd3GN98WRf5ewHs/6teJ
Fy0LKSO5az4GZysTbnJYLuCzI4qjp5zP3izh18Zo6aJqOj9SV8Tk1gmJ4ec7hqgPUVdazZJVbflE
jq8zLNwEk5WMLIdmqz6cBjGDi3koI16I+E/sHwAwU2yAX79pC42TaWtpljk31GfdYMUZZv9Gj9cg
D+kBTNpWKh2YUwBKk0NV8BoB5Sft9m+IOLmMx2hewcA05ILW/mnUVMOBbClYgmasR0iT5kpCK2BG
oafcgmknGBIj2bmXyWY23Idv1TbyGC8guwikgrowryIf38mLXdhyWBnhilODX2Nur1t+lFruNrHm
e9G+nul323W0yjpYk782A6Zb861p5ycBxUOdY3o+XbVm1yJ5XTvh5nsyg67PDlDQVaxfLbGBBkOI
NQ2/tXMCSu6fx+L4o8WpIkd96R46Be0fqtKP/c2f+CnO0anMq9JiwI3z8m7+fYuWBwKiUIAcYXiv
DG8/NrLHdzgrMRi3FmDAgGB8v0wmrATwTpQXzmVSzT6e4E3VftfCiXXF2dkfCsUHvcvD9lUjoXQ5
iCVcW2puSTTnKg5gSTQn66tEQMPa+NURbF1D7fY4nSqzxKA9Xs4nBkP/z1Sq1OUNfHW9zNyWoEx+
B/pF0EMMQwXx470xtcrk1xn7kFfKTvanzfZgBFiM4/z+WmrFmj/s+/WAcVIEvOXGLL0/r/v/JTvv
1PlpjkjCLXxpsQroQybejFu4VOcVzhY5VpjdT5EzAId49yYk5OAnD83OhuPnrMr8+LwGQqD//YYZ
vVgMUNzD7rx+daxX54+OCdMY92VcsTY2YLwzUzOgC/URdwAIvBWT1nQfiO//686tBwPqK1Y6NG/t
LAZYsQTIjoO6piItv3d91Ifr2IgDwSdterqYpKQOdR2E72cj59Hf+WGJlah1APmdJqoDdywLFPhr
Q9A2bJcUs47B4zZQl2iqAt43wN57PKL3bLjnLTTigd522KCm67Uvf0CoOUyCXng1uuAVobOBh0Lj
xcwWSlCKtwhSPCoQ7NViRRxeFfs/Ehujs5+wXU43TindVTIXw8zGEA0sI2V6reQlHt8cMDOB4S17
AItmi2ibRHoWhiNJqbGwNtfvw9iv4zJbUz0ODvDCIK5qCMtb/7wjWhrJoMu62cNrI8me1EkaD6Am
zsyw+9ZgucyW7IlV1Cd2gOf1I3j6l8N1fNhtiywfi8o45j0Nb8AQ+irEl4agB1dCIXxm31cYw5IA
eUprw+tND4ltMaDNO34VAUE7rNcs0ofgMOvz/jVS5G5zWWdUd8+dF/VCaYAxTYuLGMX/rI2UiZPf
lskKfDe3xROUCg4vUaGGUez5CrfDU4MvLK3EwHTU8nfwtgyYM2oUeBVZp/1iiyLn/rJuAxBLQdpv
KLw4KPrCU6/n019Zpsndg7O/ocDvQIh6whlxAYp/tRQk8+by/I7XBkZcXUM4fd76EclEffW2N1zz
2RtcaEikyapyoG4Bbuzpp4XT2jQLBkluf6f9hQY8HYN/oK39NDCjClBvneprFk4ZyR1bBOMwUxPA
0KyqpnJdXgvEnabftgyw59Evvhsb0IAITxAepHmmTY5H3eu/iMm1tCcWCYTJMxH/J2M7l/XD1CqB
gdbS4ql9t1untjFDUWTN66CnWmQPsWBGJQuhqPFIXj0bY5oft077aNaZeSdHK/9WVoYLBncbdtYV
hOlzg9S+bNiaxmc9pojeWPIFuQ4vXOa4CC6pE+i0ZSLRf0jFbHBDlidIndGUPQwD+zdgLr1t+Wwq
DAugsSC+EpwgW4gUaZGsNKxSkLv9khWDW3TaaraDVVysHJftTXFnv28hMCXBeGGE36e+fOoqgdR7
4Q67BAQ0tuY71pa1Oq8lii70smyzA3DMq3pvwbnJ8vzcoIfNflzBwEpzxn4YdWXldGD/ClnraRhQ
hQ5kuc54bM8iB6zcesvcGRdmUrWR7YlZRTFaZfFWn/FS2mE1gYKL6iwEgP4hyy56SeIi2N2jUtcJ
6dJSNCbVsJb558Bbb9L095vBOr0rl5ikXnkBwzNZ+ZJzRT8bNKYWAMmcYB6eHvsLLx3i7h44vBRu
aTTs5U31byMzFRuqy9pwLX6EseNwHg4CRnTEIUzVfMTKXCjH+tZAMzpGGrx9XC/vC16SRGBDvZKe
gM/IgXJ3K2mAv6weuq9WKBaHoPSVTUJzKFrHaDOgiDYjZjlfWhVIcW7S5vGjf0pRhGyhqAIMTa9P
9RzVyAMVUCgy+PQ6bWZkmodyBSvnJIg3dHRYhpzCLOpwlkm8Y3zLKOueWlfGzzfatG0ad//6f313
IVm3d70TGh/Bh27Af9WKQZtoiKf1Oedn6vkKRGtttDIYSLaupWiR+Fpdjj1aDo0poDPFK3OvANdr
Cc/yTP46WfAEB6fSL73pjDMA9QtFI3l0UZNeJi9m51dVbcnXkR/QcEWeh6jf5setLZFiSgKy6Y/F
Hb7u5P3wf1mdr1RaRg4zGZEfHY8FnUPp5tKzBBqZu4NHwgp7sV0V3uGFLBWBYkYT+Pn54BtD9nEx
PHyI0iUJG2mpGrQTp4K9WQmjCoAVQXxRiuCkAPfZaECPYotj1E2GhdNuk3swM7N+DDquaOugW36C
ieo1yPBTnh/Ce1Vsz4MfJjFYa2nU1ANM/Yn8IjjF4OR3GJJ+Tx6P2Hrqh+/FUkTg2Dl7g5NawX9S
LU0jGP7yqDnHo6iGakAYAYF4rf+cMW6bV0n6Z2/c5wgbZ8V4kjeWxtaszdWue3vv+J7V6nqI56ig
ofmm496dD9BLr+ORNIof5kcyKvuJvXYjbgRJiuIA7Cvi5bsZAoK+iuGM/KM3MvGzzin72+0b+TXO
orkLLFdtFX86LE6AgOHaOp62gCoK64bQnGylN9J8Q1hVhsvPug21UYMq7FXPVQdeD0aSPJ0Ft1pi
mBikLK4q0TTD1hmaOvagGXtpMjtH4G6+DoIVRVXnOYc4tFEJaLmpSXlUmVlDqbfzL4Ptyj9ny0sK
UGIS6OCZY/Shi7pPNqlhojL/SvTfe6FBBHsc6a4w+zAiCbsItSc2w2oBDSmmZu4dfJgylRfZykCP
5sE2/CLEoglEjGh4ZfWbQkBMAWOxoF1rahpHu/OYAvhFO0fHgyYUr17RZLrlrcqcxdHAWhqTBWzA
q8qWnA99qbsGSxYwEF9Z+nuD7jrYa1usodItGyGvcUdwNje3haCpX84Dr3B92OiFgfx2x64Owt5z
9VixUktlf4Pmsloq6+6SXoXjEftmjeEVkXl9GO4MBBJmHyxANz8UkLnSHdIEU8IgMWuCY0+Jjxin
XHEQKN9N57dnK4o8w0fX7Sg6GGUF19Qck47BNnbixF7qM5qhwXfRhO/IFEpaYjhB5pt8VRNdl8UD
zsD4i7LQEyDVtYKvlB4BgjsfO0DJgEVveQxMERphxf3nux8fIltmzFgzBlWmlRQ2iWsPFeglT+xz
2/XvlTHyPAVKML5b/zJ6tVQ572ai2wtoYgmxP1KdReFPd29G5msgb+YgY76AZq8NdK1VbQsBYwlL
+p5+lDTFTrvfRVD0pl+9z3HWbKFUzIUlL8nw2+Xy+FmMCqtp0cu16Uhijgz0Iy6n6gIRzsCZ/0dp
qtcFpk1H+ll/8mDF/UMFaEasQzqZXmfQNfTgAsqkmdfoipYSRBb7EvA6swjJo/nQoPtONFQ0Tqa4
crBBNBKizpfYSn2D1a5aEp5PG48Muci59Pk2Rv1um+hXCLcEkzDFjAAJ2jUrYTHp55S3r6aLFjUG
SIWu6HYXCma0duBxY5l6fWTwTv6cdKwgfNGvUmE0zha6t/3t2fPoIrqR5TDm/yO6dAj4IhzCBSCc
S8rDPGv2BuBJ+O8DWummUxj2BtlTYu9LuHGgO5QDjy1aAe2n0Srgwuo1yO73wqPSBpbwYSPWauyE
aiaenUDKqlRL/RIh0JzlFmdCM5TIHd7kD9SRal8gVGid8sFDYI95UCuRjkypPwAm843Ia6mGRdGD
wrZYL/Y51lpjkHpNPVCt9yeFxYgZiVrXLZ+SCzU2gszmCLeaOL7u5E1APTrPNS3ulj9Ua+x+xNvJ
30e2xXE4RpcK4NytgVnx6Tgp8XMBX5ipuigCgBGJBqaTdw3Mj54cPixdzWgnty3n3TY4QVjFLpwG
hf6zi4uNlDi2QHA7wKXLiSxQgGvur3Q0Hjx6PeCrBOg+R9d5uhMaaOfQFG02W0XknEWF11CjzQcA
8EMzfCAy3BKIIEYKvAoxSIHgd3G/Gk3rBaHImYSIlR72k+776ElUp4jkpvqlKtFwSPcTM63asww9
YEgzFVPgQ6JLhfLgGCFFvT2ZzgqBbtqgVIcuAP/WCZDbuvJU/vWvrFkdRUN4YcXxxXx7NNB9/NUM
FrcQEORHekFzgGUidtlXzVvWQx0k0x0N++8BrRjGEdIJ9+iKmQ1hgoL96CyD5uWVRJLXKbFevdFw
SRT0fPPQY+MgxWuzm3OenHmryW8ovhLB6tERNylKiwEeYfAL03e41NRU5Pu6Vmwugjr2y4W4Dn+/
C9J10/UwfPxNrPHJMpb8xPEERvuI78bxcDSmiFeM+mMYD4B+i5MFQIK27HjjwZbyPjAlREPYOdC0
zDPPOzrShFgZpob8ZoA5jkUoit/i1DvfeD/UF4BdM3jgasLzmXW5rOE8MM9fUpcZsBRzScaQDlix
a+TTOCJvYB++9n/cKXYUksaAmE8CSpxKVYiu3eurZkNXDXLEmhpR+TJQyH0p8W/5dR2NLXc01E3H
Ke4CgX0YGuzcEzlGgW4PpQXvU+PRywMhFNmJEDkqctj+hWuMFdqkw6hQxNAD64V51EQ6XwfNbDT/
XBtPMoejFGUtTd3+1pYTZ/1lbSZsyPtKxH6IvBW53Oi7S8AQowgZpmS4Zebx5a/m/r7tkYeiApyM
R3aC1+B32k3iJ7CTTTx4WQ0HgCPDlAotWlkITu+PVbJtRdI9zBJxP5z76HdVsZOOXlBBoPJD5vqS
Xy+QgoVZpqHXX+GPIEbGJzZmb/0uT3ZHxu/z/G6CEeK9mzJrq3mAgWJsVWLOO7PYGJnnvPgk0CS2
1zH/xOKfwVk/YvV6O+JpG0/aviaKZy7Jav96T7ADoXj3XpsaBawiRR0UVVVH9jc25K0eivpt/yZk
H8ab+gCPCPvfP6/JJaqtTsnR9MoIgK5NgJXm+FEbR0TA8v1SWyXduIBXOJ8kMM/DOWRxGcyPrNtq
1Z44+CwBPGMkWgnIaqC1nhJShFDEkqCaQVyRzwI+xG3GQcuzhZ90CZie4+KJovnwCyYTpm5sbhTR
oOLVmfbDaeTyzd0gRtg3cStzXZF4CC2y89l9qaIuourTbLNLE/I8mVBGEH/R8rR6pCdxfh/9Zdz5
300mhFKl3XzORv+aqp0aLFsEj4lu7eqg7yf+LH/2mInD4GkmlR+MeWoosSRujfk4AB8jQRnomXHf
fXMJ153wsTeDb/Va6U5k49WbbMLIV4zE5fgD9RTHvTKxyjIm3sa8vQ+y+NFjPWPV1gZW+iggrbyl
+b7LtG4siEJFfNXbCRSvL/0OzNN8gNG/3RnWU3dQHfuB83/OLBBDo6ouGzXk0wXnRp66YtTmaaIu
JNHji8pMyw5yEsukZ29tNv8Sm4oO/vhhWgL91gck3SZwPfrRz4QK3+r2eProSk53ZdeXUgcdYAn1
y7Ypfa4ocYQFzjHpamYxolZft/zIeqyXP4c7dcFO5zO5HqUITOS6i2Z6E8mazK7odRUE8fcQEMyj
N1cBZmvQf92sDg7SDK28diBPPgNlLbxx0kjNR3zVkkkZECwok/deZTzBiWmyeXgzDaj0p1h6oTsM
+sTBHB/+C9yEvSGs4lBMHe19S2io8QrpqUVtlhev51OuckkP/NP9S6i0MF3jWRehbcGInQfGcxnN
wzygs+mnqqlXQycwr2JUsUvbbqkooa/cvHDptAyNzV1ijrbx+A2IuETJVtWWalcGE+nY7Ti736Gv
9Da+lNxd637FyWoWArOsSx+M395bwn0QK9a6DrG3AwFscHR5AMQB9viVomAEbywL+fN3PXCnBHUt
mG2cePDvBhgIl0IuFUlfmR/zPd8nadTNDPFfLUoBqA/WtO3YL2SNTpW+NY850NCxpwLJ0J6h8coE
9UxZv8KvSCZkTpXcPM2p4U0LoBVcNljL5oSGZuECkK9eIpbWPSS0AJocnTCdxruKctJ1RANXRbm7
naE1rxe9AUfUjIDF4QEoRxhipPvVV5Hyo5G+Asiw/FGcGHzYmc5t683/zAe87cEY1v6x7jbvbMDn
IHtl9USpf+mDRsTKnENaS7SPbADNkZsZK9oUavrItzxEMwobhRaRwO7ZCXJdJCvhieVCLe4/rm8J
GBNJ9nO3n/NFyr1GTCWdyPkQ/RU2auMiK/hm7BvUyh4wRsj3XJAX7Hde/HcbIxU8X9XssvZ8Xci1
Sgdlpr37lU3sO5Tht0sgMhjB7tz2ptFsEICyIfhp7JxuQH6g2L1huFzV3BGX+C9EHGz0TBpJSO8j
DzZ/TkLm5QK2F2upvyHsuIS7YBZA8xNPnLCYHVjjI2a8w0yb7ZtEs9RijHMGekhXhKDArcR450/c
y/YPNZJ8w7KhuaeRllHxOwQW5wLIvV73zB5qfmv29Hhw2d8U2/5KT5KtEoUVVhS5o9Lge/kz59Dj
ODS4F8eUnksHPkYVC92Rew8fQQJak24fjS0e/g6kUN6DaVhiwueqI/3nBWbeEfsrA1JgupEDqTZ2
ZMOPNPS/2neVJwFk0nLgBg6wC9DVxmQTODSTegJRU3AY4ai3jBKgItJKJPNO4UqQS69gn/JjcFrz
xA6Ro7/DrHE5oCuXw9Mhy1WQIR9EdW+mjfGu0Xiw7Mksudztsyxlh1q6/tMzFK1KqJC/h3JwkT0z
IcMiEom1vMmw/XWjncVR7qL/PjhcB9aZ/28jzukBUjl3z+hdYsXemlJ2NzpzuAj/qyVSulOKfaoP
5M7iKNQVWZ3K23/WShYfOZO9jsMY1e+lp2Rr/IijoGtz99U2zwBWmzNwvL9lXeH+MSIcsZ+pbzF6
hLY30vbBiy5T6hXD3u1C2l/+sRCqvHkSQ46aAWGJemJxt8t1l8d4uO/q120X9GabsY+BksaX3XVM
BgtXfMQLhxrn1Hqv5CjkugAYyWrCyNxWa5E4zm4fkWAzZkTivBNZWRG9nqpx2sfklYGqwduilHm5
NeRgDufY0eCGFdV9HgFg5EM9yBJe2JdNyhOXEaJsN/YtZfeDPxheiCYd7mrldGwGAoOkqwBK2PjC
57YCiSmhSuY6fCRDKfiKowr2qm2SFMHXdTijJnvG5ou2cWGLEKN9pol49tbXHS+gKiNnjoJ/ZhX2
fgwsLHZ5ToeFL/K1mPmJV1R5qPeINPnxtvbYzcelWLadrqS78voFkfRUoGOtH2P2YXG0+pal9nG8
ngsG9wOs+EHEQ7A1GzW3AvOVs+HZiNvhvFnM/vogxmMy2Yh6dBkMzfCqnDHtM/wXzZF8h2kQfD5w
DwfY/wUVmEH9udnE/caqLvmwj5Qq3nydh5F5gHbrjTrdX6fSS0jQ1DJJ0p0T2pbBvAsV5L33gwQZ
aJn+Zi3D6JUJunvpqNToCaMgGqmn2IUXVfL8zV6UU15J6L8UgDNZhLmih2nFbLupIbeky0m/1RED
ScO5neGWoLVfjcmaU5+Ix8RagAZ6gCoxoiBs3iiP8uTwUuE9xOHIhU0ZS2DpGPtdEjfFhbt1zfY2
T0S/raar4kpvz5OnFxM1++r4EbJH0ay31e73dJUVRqq5zjfwZDSc/4QQepjx5r4nQ3HsaH+HNniB
tiqSjLHRK7Rv6FbYTV93rnzPwVb9uTFNJ28Pnfsipc5N6Rj91M78iIiIDam6VB3LL5bTHlFOrstm
fQ7J4lZ+96/EAYWofFnCIT8WOAKRInDbb8IgZ1VeBH2hjQoeOZ+I4raJTJJMBriBGz0T1A5AD6CG
X8jcCoeWy8D3GaOqNGo8dSSzZmkndbjWm2z55m/uoPZTuE9E2Xy9Wd4Oa2e83WvFO3BDYsL6RoTg
qYNoEBsDhRdlNZ39JD5hNULTQtR1lWPF91hguJNC2rWYFmVMizjX3PQ0aKbOPBb5BnyRepeEmF2l
S8s8C9297wLM3Mm8Oz4NlT+Sq0M3oZdYEV24EY+dW5na85MA+dcC2zmr94JRfVPeqrfPnq7gvU8d
DcXwUNsf+RTefcKs8LjmOJs4vipEKxXcbsG4Qy0JePCkVFNj6GlmL9wPN4df45uAKlIJ+qPLQ+Wb
4OyxnPw9wyJ997xJSuVDjxRspPbWUIoCf6/SHWa2HlSP/OG15LHbqwEtW6f9n/bKa0NpxK++Phjt
2O6SHGD5R9JQRZ0z2xXzAdhA/1jrJf7IYwAd1vkbuSNjQOWi4di2g/JHTmTK4IMhQzft71PLnbB+
MKXwQslV4RwAnsyNXdb8x/Oc3E6VYaPFi1OG7D7MjQ9beVuevtdTIaU6HwrChdLEWfPlsaSKtxxm
3paZ0aO8tOYa4boDi2fEUihx5jDk8qjOS+9G/gF8LqvKwUb8bXRW5i4cgPM8C1T8k3QDVk7Wt4LV
6Udkh5fLSnJ+gU/H9x+F2vmSp/z7UTwJ75/W1CKTPtogGyeHoLCoTYAD1f86pK1J/VqWRySwE7x7
1lsDMtrSDqT+rHglWiOp8ovXvnnOAQ+YjHnLNKtLJLoj92x5DoXXwuzFMY1a4Y40Km0lx+BvsJlt
CAbylo+5EX5NusWVXGhc3gKJHtE4DLbpHN2tb+de4z6X4fiT9vg2sB8WCR50+5BuREQW9YyorfHO
9Sg6llQmt72qVg/qTc6oBY1d8a48nAnYmrsuM+jc/2/rbl5++2Yhh7V6c6BsGNGUiL8wrkVI9Py/
y0K5sntYwWsyONgKKtI3k4VGb74yKbwaXqMWj6/BWWvqbS8ghmhvnpBeWtXvzodrnZrg7D3nrTr0
/cVfizu5rTL181/ooUVdqkzW1Ak8tX/kaHg6pYP47xUJNhAeJO8hrwxO32T515XWSX9L1HN17AXi
lhQbbwHbniFrmFd+vzyqJiJugCxeG5i37Qe82kEsSTuR2SMMyPpCLxZJcKWI0L16D54hKzz06Wxk
5CrOOVV7MuAkrOu8a7/BJXj3dGH1zK8JE6sB7Rc0jPjgqF+dXYBs2EU0XZa58iH2jbsJi2L3IR4x
IxhTTY1Cc0c4cbqkEkqnM0GQxM+wu+E5HTXskrBBTqdj3nOCgtQaXANouYuSULO6x01VyKcZxfbK
DHL5P7ZxI5oRJdDRQkM4+O6NO0mwJhY3Spd9cs4/RDjUjW9KRr3BreHHhpWJQJx4aoAnosipQkeA
JrHAuRBqcMtSqmga850WuXBa4h8Haa+CqD8af9ASWsY87yO5Om1BOvcgXiM9LCPdpDxYY55WxQh5
amuF0s4ecJvrmAgsQd7+7d7OREHFDKgkX+t5/OHQtXyCqAqx5kt5Cmwd5G/64se1yoN3fLAtEFv4
K/vpMpCicED1MhRqgY0ikxVs8I0wy3pi5lv3BD99f8CkpLxWXOfNS6lJKNO2KGuh/pUT6xgA70Nr
tdVIVoDtG6TsA2YNb4Z1Sqg9UQpT1Uy7r14FcsWv0e4dK1Crms+WwBm5BLG/3jg1Zp4aLRZxQsdv
v5M+kzgaH9LLrXaKhxo2fJjlF/eoqNzQSmeJ4XJYjiRS6DuhBGqjrzgqBjTv5R01CGWFYlPXfvZ/
MGOHFJMQk3r3seEbGAxus75moFY+ZIJXgHRsM+Bxsu8cg2uRBvCdgmnTzNO4z8nvst4Dg1Fg5EkB
fbHDCT4FnladQMPXxcNPIdYV9ud5y66H1yxjAtVdkcYpz+G/16mUc2RHrJp2f8C9cwM11fKrcd2c
88HO/jWJYDtjvkBQ/FEJPmkFd7fj7txhl0VNjSfgzoEfV93oDFUlVLrNBdrKD2M3jSCHbfQiWdnN
M19bzqay1RuZi6FsK0hNVZ89EQ0yLjv4hGyiHxQhKTqMoyp0Ov7JV2mJBv7zv/T9SWl4Gb9qOeRm
vl325blcHj9GxPMs2xxJjzh4u2PDAzVAcEq7nrD0+BzjuzxtuZ6KTM0XJXNfiWnJKBbUu+f2nRCF
wp28skZE59k4mkHqGK7O+2u2ounPppFEd8b8oFQP1GHi6ZRsdEFYbi42hXR06hpBmNXPlsRu2B+7
D6gQXDOPb6mWvJLAEXI+a+ig7UpObFFQdJI32cqumkIfWEq+5KoPXx2s3dmcj542dZyaNb6YkFG/
iNw5UzAm9BPFPAy3whHLj1XMIqHXiuh5+GEGLe3hlBl69DbbebnrgyH/r2OMP6HeIfSc7bk/G6Yp
uwCFPKyqmHe5Cv/vsRkX7AdH7Bmj0XerE1aK99/E8gYYfV4MW0e7TpZGBu6GleXRD8YFqtklzx9K
j5XHtF6G7+jcP2hww8OEjDjqOeh8l32yN8Xmafz8xBmbJj0G00uzmsfw5zbTznCbbguhUqp5ST2J
6f3600ZF8MyDW6vtETXouwrDR3mhExv0tar0WHsv+x4FcjLoZOcBjVtzdb0at8TSHaaDIxA66J3w
CzLPRqOwCauR0omZZf+SmInNM4R6/kzraVifULQOsxU65IY8TtxQkTH9lL1jvJf2yfr7E50RDkuW
IphT52IRKPFdedMY4Uv2GOstRubCkB7rnS77PV/1ZJ/NJqFd4xn0yzgOdhv83ohPbR3PaA5Z9Awc
87IuTs93J0JGHYq6dsBnYJDx7+lVnOYhSiqxiDKYfzHMJWTG5KSkf8mH2FvQPkzrse+grc403RWE
EcgdWRpkBM8Njn5yzMQjFM8PWsckdDZwn5ebcOaZNAd5oozw9ZXoMQPa83KyykZmy5jcm4a/3mdy
kKzX4gkvMMLMCzTUiXKVXOqjm4D2hPSfm4FbwIwONuVGCVo1rOSe0jFEtWJbMaNjNakZ8qVhy/tT
o+OekjdSdh79yEhjYC6BB4z9HitJDPPmusrtVHbD8WPLitRZA3o9jNpmtwfulk87Jo2ie+v1Cr4w
GZyvzGoXZiKwTVH+78kPFON/XxF6zKrt9OMmPppWh4PR1yzTr+k1q1K9dHvfgDiA6yQVoNlrRDc6
ho+fNK45i6I2/HxESb6sJ+lzsrCTqHMjyMQ/mfoN1bb9hDdpZkqcok80SQoRScS/b9rjZmoBEgjD
0ozNbdJCuVGfw0TE0A3EXZToEmdL657CyK/y0E1sEV3ULBAv1PWTPxEIMVIEu9IeL0EHL7Ct9E0/
/vUzNGX8SOdV7FFb8IvmPmMoVZG8Af/Gw95gzw3nCgsrbzbn8wl0T9EObAceoVQ60fRiuhio0XQ0
ZyyNCpkEBFKdl2TXSl+HyAR9LcvJJVHZysysXKx0dlLmHWj5dZQrVCTxN3sEnmfYh3vJdU+PFhkT
/orZT878pZUBfAAbDPnDb3CqWHpcNgLXqP3v6lsRn06Uofeo8TC92atKFNv9uMs8ewmIyvRlxcSh
ghocPUzivy8qFNhtY3oQ6WkPOgHkdcfSiV74EExKySRt4wV/fE6AR7ogNYnkNwXoBJio+hMZXQ14
EKCD6LYzqMeHHPXrUCmvgUpzgTvSxS8HVti1TDDmzUhBGpHVsUIpUHz8e6VlfvXdjkX2nnb1JUPK
zoCnHfu66xTD//J+6PXsj0Nytti/VbrGVdcyz/7Nwfyel1SUMszqoqTf3NnwUpcK97xMoVEujll/
dnEsDqkXPh2UElX+lEMJg/SB92MN6RiwHo4lWwGfrh20QIE2Kiar6vmmv7v59UFoCC6NAGuMSl6X
RCQPVemxjoZECjzQ9ZoAOTgVnYPrAJTNtUENnX0fhVm+6B7P0LH/fLpjrWdbhqow4Xgd8fdens+w
Aqc5mIbgv+ZBw1GkarA4U7lqiwGsSvPE7y8CvtJ2NDmnrRd2G46ylRjvc6jN9CWsTd6zhIhvTouj
OrvgjRr+VKYPSDNsTSPkyKxYApx0o3pPCGONKGJG5g/TJUFybWO+C9qWAT99i3Y5IC5vzdeX8qb9
96jVD4VDl/T/Ri2cpMkX9+axyN+0l+vrBXmvn3z6WWxvFB8u2Ca3bx4lpWa1DWKjprXBIiPQnC6+
+TS1np3ZXlu8Kku4JzaPqhTCRq3DeyCJkEVOebnoIo3NjlXrxzcG5Gl4N5i4t/l14NpkfsticSRD
jEbhUhvlg0dqDNIFxvL0b7gCRVR4T7oAddYV/KDB8pk2T22vcoC5taxvkyrtbQI4UShsjn/4uj80
+vEWWCkekNPEgepafNsNGV8TrpX8ME9ZuyElu84Hq1PmHMiUHSPcXHIOL5zhPmXs4+ytM77flAWn
hC2qqbC6dF/C4cW369wuzFds/1agOafhLU4vqlTwvAXCtjlpljARcHcxLSRu9g9w8tNn5P++bycJ
hJ+309Dh1LjAEHqhLF2kgTbbTHdbdbVuRr4JmYkkTQUeTrc6mjWNTwH9ULl3Nxz1YTkFl+j8u+6m
cIQvPI9OOsa6rGrLJBhA2nFSjCVdN/LBIPorbuXPLb0SznQAkIyhKMYAjm+C0LsxCRMyUdr43gv6
8SKJat7Rk10qjF+jJUsBYvuje6XtYQUSKX9y9zdQjhgq/kzC7XjWNdVZPjYKsQB8uZoLL+fueRr2
GHZgZpCcSc8Q6xINJyHhDgrOQFmhlpoSCVOf+x4XEt115SQDWkWvpxCk/E0pjaR/gtYGaL2LPV/B
xSTizfHFzRiKdEVwANYSo0GsTWetwIl/rx/I3g7oC/mQDtV+j/j7heT0LRwGBqrykyKt/WeU5N1Z
VPGNN1OAxglz75qFiD10d6CegNKjLZZp+8EF8DNqKzdggvivgRWsYLzcXXgJ1I0zVjbL9m81Sd9M
DQqo1pOSP1FA6Ld8fNlq+3HRHGNS+9JMIuIppvbG0sVnETN/z4piXiNBTYapz9Vf19yADgZHfUGb
BNWGLdcYvY6qRwX6sE1TbOPdIYCvCBJDsCP1U/xo4btb6yPh9K2p9EDe9Wxo1HVF5swOjyhycM+T
IlIFBMRoYeotZaX0B28dStdzmdOXhavEsvlnodnNpOeYG5XxIh6p6dxhFBm9fcseAC08O+Ypdw3S
YnPtZDiKoYm7MLWfRCtElR7FVnj1DaNzpHkmHwpPrg5VROxyVii4Ew3u9Bd/Yv6BxblajzLpqO9b
PPAhI9nZ9sWdfbKmUy6yP5ozbIoNwPDgHWI1Fdps6EeRO0/3/FOjKY7Vr2m5TbrQqCzWG6XrhtTT
2bvnCiBJt9aQ7YmJUNnsCfosEwN9bc8+IfBR5WfsbSD/1y5//v40ZSSrDYZ85rFtfEWJHgBYY4IK
Jwi0oOO16bHW4g3cduDrLP4xsZpvyRlZXdrZM+7bA/xxj/NVD/cWCecGg8sHVq1vL14UPE0vJE34
x3hUlOYZz0tupH56we2WsRVigvJH0Ks+xrsFqLJsKw0O+9Sd698sqrk89VE/EXRgtIZcoCOVxew0
GhmtJwllxejXkUVTri6EUp3v9d26lDQeFK4Lkk/lZTxkDkSzbhOVZheMi8QSYH+MaGwdeQ+j2Clg
N0aR5e271UiUwdDKpcKUWvLSLwdENVeXBC1Ow1K7iJHziY1Mz1KO5mvM3V3CS2ihQ5EIshnPbS38
fw9e46C7RJF8MIOQcu4kx6sYyJMOym4TSR8VIB8kgaiwZ0VktqBgXTMg+yEsD0yXnAfvrLGtUDHG
8a1dFrVnBbNyef4nmjS6b0JQUhv6elNSnP9XVggx2ERK6RmYaT41fg98u78mgDPopBOa3NNhEJRb
1pZSmyKRikS49MEPYJVLgA9FLiU5lGN/w1L1QLJw4ktV+qN+PL9KX3KqEHiEGHzgLAeS/4e/t583
8GDC4yzjOkdLHRgNG2ShdJI5tI4C4TvEjC4DPJo+8gdbHEenT2qBE9iXVH/07MdIsM3WPYOW/6wN
xhRr/HFWk5OJBCzrZ0WAyEmTz5L8lld/mqoSKKgQ0nwcVH923GXFxBpIR79EUhcTm7oCp30X6Gvi
jIuX8aOyG8A6Lz7K0gdD2K5XKX57Z6Qr+b09TKHH8Cssx5n+6sTC2Jng1Tov9VqGvWBpOYcgFp3x
eROcTCVsoGGKHvaLdThSF90BmD9h1g8a2/xoNQH+oKHRHpwbWw+WUqNZS5w2GMkI9J7banUyqUUA
Oe7kqKWZ4T6cJLjgbt31FCzXS8TBL8JDUH9w9jbXv0UdFifpVLIN7vnGVX3/CoomWn973xA4g23O
PkGkbQIrfvASqQvh5m6Or1P7idDNWxs8PHY6oCMHAhDeXrjOzSd7PDW5Nm7B2kmC6WsiCRUC24kR
ZtXdquY+uaPGsXdQCmoSPMbV7Qa41f3WM3GYf00L3MWhRjjKjbsl7H2uMCuOI3qcfki9ZsQRdURv
8aYjOAULJdW1lpUEUnOvKif8G8DuiMerKryoAFgFp2ayeKb6X2eNUaPtgXlsPlQIBfm2el/D1rEg
H02Ug7spl/8b/4IhvsP0wmYr6UTew35PYT2HxJ9BXYM6pvrTzDQTS0V4U7dIcpSNB02Csvriovcw
Q5hX7OS88nshvHLJyYDhH7m7TZu6nohivbS2N85a6MN181lnNn+FVGpncrFFtyTXADZZ7AZNrqbh
1t6acN6KmV++qOmyFIrzQnMNBnH/BQh9FQAotqJJbPU+MzToQGmtnS8ls2vrqVfww0PW5NkuDjnP
fUpJEmUITioPAiWEYpVOoweBnDkWg0UkyiKO+VE4l71tJvJ3FqM6HWT/nd44bUE5GT/kaU1f1dHL
GwK0B3XGxX7Dj1UGtfEpZbfYtB1z7fBR3Fqpmv/iYPfPKdE+IluFGXMcow9ak6TuVp37t30A/Vhe
3fyaj46im5O57qPARA7WXsQEzMtbvy0EnUh2lF1A+RDruK/OwcVrpopzgdqA6ufQEQMU+dzmQnH6
kKD9s2uQ/5o276Ff/lWnW+v0DOtKH+LZS50Mjz7ph5JB01I3e8wKGby6qf49ZqspiFap9n9rm5AX
fGtFVzxGEc+DF1g1hX0CFdi9O2A3HumuffaqXE0Xilqv6ImxqTrb19Jqax4Yz1Ev3btbQIAoTqmt
EWrDjdR/70cElrvhvyLVXSBn+3BR+atg2rhbv+xbHpM38GJ4ZD9GrXQ4W87JMjD0yCm7x4RQu/SB
33krHPiSAFyJFLF56pAdZIsZV059vXSxpOvvcwizPwdf3affoHbfb9YQrFoi5f0q96eR6+IGNKHo
DWslAqndnqaUp54ZB+Bz5fpQ68tpJLfBbeEcrNBG5FkdmB9smLuN5I/JSygHNCtSgvSlieMng9gU
muR16gNN+amCtuaVGpWsL1Go1fYXDOkoqb68xEPdX0GoxZBlSEgJD7svx9lcXbWsaBkpXoEhsyAC
gBr0HgO/TZOQJTh/96Qa0ZHAZquivFLaM3YZ4G0v5kheu7ju3AYltBMNu65wgeHmbgeVyzzB9OJU
zRGedIQXc2fgwwMpskFtixaAjHstLZiL3JXci02x8nIGDnkDzFLzRTG3U85e+g3OglR5zF2xghwC
9V9vBi/tsRBXReEgrKzdr2jj+Tvwan9DMlpWftrn3dM8YitKfKXC53+3wJlNZMMuvpImiw7qXWaE
6AQK72zPt5YpWF/u3ZhUb1Q3W2UkKl1PUHGDJJJ1YJu3vvQkYDUaruDk+ysS6o6pGd1SWBlTkLGG
xxLlZmnYeCGsMNN38oFt0MuK0QpfE6ie4CgX9AZOuCO5gSUmHSjIv9lpxMRFIS2okGkT3x0MwUSc
15o02XvH99JnjdUXR5t8YT6hQL+BgtKtD2IhY1ct16T42OqdaTm/jXy0s8rd5MCLORczGEkFp20o
nDuF4jL5Ogeal6MENNtiqY7XIp2ezAKRtfcrS47+KlF8YrqX96Hr8+lOwg+qq/Jnxu6DuVjYE/Hh
KJq0JTirt+uHjjJP20I58NI6+Cy7oJDAKfcV4QPRRC33iMXnJD4V/X5ymk4aorsEZzV38AyeVm7r
sTpHvycMbfjrp8RFVOGR4p5WW+zRlmsIHmIbpRhJpmTrJcc7KYPgjcRvdLZYJTrTf4pUbEa9PSDv
jImx2sXCvzuoaYYmKl1+HARvMGVTQd3Blqowa1pTyiqo2EmNnDxPyQ6LQzMD7tT6uLhjHvtH1pZN
Hwct46ARGo9WLCLTKtyB8FZvBbGhrP/iNCIL0/dWvFKAQpTbw3h+nlEs608868qx2x0AhFCFOkuG
oYDYX9ujE2CghYIyiTt+oU2QSd59vIStwL8+/UfeRYjdvhBvvY1Ni9NIFrVAvp0Q3ww4xgS/1LvU
VC68pfBX/KidyuqnZeYk4tSpElWXobEi95LLqfOmJ4lzzTblLK+awhPk83ShLb4Ainn753EG+2SL
E7MN1fXfS2qvuF0XgT5SI5DutU/3BcPeYTmPlrPbKCI5Ovigv46BOErLfGQlCmF5iZJ5R2Z6aTmL
o+APT18nZrkXxJ7j7ZOWl8PnM+LNgE6BXyA31dVtVqffA35WpwojuvTOH6qW7cz2EoJ+QN7A3O72
6I03AsBZjBao4+eWIjvvgRK03Uhv5QWPwjg2O3IyQzqUFhRDfuUnCHl+h5sodTTvlDjOcKxmL09q
WAUD3u/sfzirzNI60xYYaj9+6HuEJhFP0zqiTgbtky4zc1mqA0Ig+Ux7KYwaEBiuWzAIKx9G8fxk
jSU/OZjMrGZmXLRIDW+hYuLKReKr6PedR98FSiSMxQ60icEiRnzaIvoJZTYskAWONhEAj3a8gVVD
4VVAzDepR0x93Og4+LPHZHJwYmMqYClpejn/Cd3Msxlk2TuhwEh0/MGqEfqcIv3PSPGabiH1y5Rh
zG+nmMC/d+YryUzhhPiyohjLwZg3Ka3d1cttdIa9/RfKXe5M1gXXEGMAEEsz8vo5ltWpNaKct4Rb
y3L0OzhyYktdaAkum346hb2G/WGxL1/9+TA5PJfLFoG+pC35HoAs70Dtzv2ULSDElQsDcGdPz1nA
cRFmgtAyaymXfHfDHq7dD8fgVNVhzLserjL/A2h81hes39fIS5cO42kxmGodqBPBbNKc4neaWcuE
MvhlDy3lf/m2j0+2OOdfQlJPYLq/OLL1Cd15JZIhyZi9cFWcRRuFnprwzGTON9cyAq93en3KMxqZ
phP20YI3DWQULIth4HMnCW+KeQPwKgZiAuR1ppKixlfRhnzo9SsdOVN8Dyx3MJUSCPNx3dWGP8Uq
6NU+w3dyfgl38kWydae5j+w7MMoL9d/GrdYD1ZFoZHgjKbXjWXwiRFEKVW4trZGxgv6qQLEx1/m+
UbgpPCbo/THOs32+RQJDnXJJOUvkcDNezg+JHDOck03eruqfoW4PzREUmgcZU9TFyp05dmVgbqC6
6wkEUVuV7K/uRxrOptMi/RLGd4vTH3bAJ2zDf9Nirl32Ug8p3J4z9OEulKr7tpJ8S+qMZTrY/jJG
clqBrCZqUkj/L1isHNpCAu6b3wOi/hwlfYDsljs7UrpuhcZqj+9XK0m/wTbiOZ9vnm5SEfs+4vhu
ptf77klWX2dIi8IciklAR13QFukWFoiRMIffETtxjC36bdHGjo5hjp4RqGgyHYgAWQSJUMpnOfug
cVGb9In4T3gh9vMkjTc/CSn6Jdna5eqEq485hGAH48PtT7tU6Ae8wpQO6v15JOddAzconwHaDLCs
JTRiay1eyy0brxD4J0XTTacaMIOnWl5PR8Rog2MWnW8AeipYvjGqvdnphZqpdgbJk65eg8ZYmV2T
Svty26njlyi9YJ5J2GyzRUDqDzdCamZOvoO80AbAZingh7Hm9ZryIK7dHU07Avg1vioYy63MRBZC
7jFA/j2MQ31C1HHAFVjSXgBX4cG/CV/v38Nl1R8WRXpHXjOOjKspVFfyvmjAbSTnfcSG1/ko319j
95TJ4bfOK1Xf9eJBhsS8xlIgw9YmtiVjYTFbgQCiJZd98ENo8GQISnKT+DJzl6EJFJvWsfPy/qDU
MM/jJ1o3ks4e1gB9UHjnEKQKGHAN4fuvkuaHromfAOp5YeNc/LVkrCR0nYNBHp9fHSasctLTkW21
Jvi1wKdrjjYxXn0u9sd8EmeHSEkbG/PYEwCTvYm26LRgmgYTVqYfHAdsdv7dVAXaQV8ROvbZsMYG
C/5RMUKhs1DB81G77H6P0HuB3kf1Inonjj2SJETdiydjH3GDClfdazjZwOdIdmbAeRsh3kW/e8W4
p2I8LlA5ElBeXzpHbliGcnqoeBXxzDGl1Mir8JxJb2jcrdo8UfLEGB5LHh1gVN3kPHOqnDj5ltpF
P1xvL7RObs9452lAgA5CraKybcO4LAUCSuPh0torvv9p6fZJX7IyZFHeE2dAThksSzcPyaX5wx6A
fWOqcAIaAGcs7Sc5juN8StJ3gJ1We08OiqEvxR5VEdoSWR+knSK1chT2d7zCzRdWT369ndxChJvr
uTkn2M8lBCVHDavJYT+SH8+b97p4118YF8YnuKgoXV6iz2jDPmab8vycSkMOeNut6+a9MBSMVkQ4
lIQchISCXNInKoXHBweNLLzgOlb0i0FfQ/PJSXeZe50hwl71zcgG9NdK1boc5Da0Et5MAER+0Wrg
xApOqCs6Ovji8N6PSeA4fF/drQnKl8p1RX4VbooONyk+8LpuWLIBz10kQQTVzN9wLCFEOGyZhMFV
USp7EEZiv9+9pQSEb1GPpGCa0KdmYsvBjs9DIsxL+kBN54Z/ShODWPRlIbIX1qep2Y2dLxyi6aLi
rVGMwlQ3EPrx7QvOHUlBMeXHDDhtTwCsHV5IOFSoPi5m8qctA7LpphmaAGDQ6AYdrqhbpHIVV9jQ
gZUPxe3ZpanGQrsVMWhFgDC1InuCWJE5s25LWsGCaHxjurVCHcARc1r8Cf/q18G4vjQDgDv+RAuV
0ZIMDeIq37oYIfuivnDErcbqOS+ZVYNNLsdpTboFxVpjpE4JIJ/Vksh5Fedc4VOkvOC2W/X3mJyi
FdoEJSUoOEDLMIalTB0mKtdHCQGBoQw8mhXvLSNcVuzU/Yfymb90mrHUWzAweAFx8tc3Fih9aAh/
MeV+M3em2ll37xNPJ/l8zLTwyxeeHuKxYRBLWPqZOvZCEbsgfXvfsEVQc3cV9sk5tAeG6Ajl6fbS
77f2CfsV4kys3UafZxn1np353HnafIwRlpvPUUSX8Hc8wMNYIZ9a2hQCf0G4xNO3H9Zy3i9JTv9T
6KSMYyB+RooKnYdvMq5FYQdcNg1TdXNCaepfY6hABgYf95G5LMxQ6t8yCZvvPgJ8rfBDE9AE8wSV
VQIvH+xjjfbqXAtqC8l3EGfhZf2Zm2HA57j8OZxcztfyCP4AQPJ0w972yyvBnjv7TwxJy6YL2zP0
Sh45DIrBiluI6zWY8oSNVcVpG5XgsygNP5wQsrbzHTcrNuwKQWGsw/YFg6JlOsBBoTyCTqKo+ZZ5
8EeASzDwOD3A2RZnvlfUbAgcs9oybFdSsn2OEnudiAxHxu4pYdk4W7SZgEK0qdKBGvveUNiYmKJt
FiFPpOW6N5IiibmtdvfZQiAebsPMdErU6G6gL/+2WOAdPsQpbtbD5RHWskw8eHbw+WQ/h6JugaTA
uw4GLQsSJcyBk+N6/YNmyOmfTvAt4UlKTzqNsb72IIbVPfuNmutdHdg2hqDyA40wdFAYtm+wNwUB
KXf85iOkMJd0Onkotzb1m69sWjQ9wzcMkf0khyEsWi+chuzBF9qMkcsY4bmuZAeLHuKr90vJA6tT
5gnVpNtEhxWTarjbyfAGNW/HCGhsDqhc5f1PsoLr9hlFMN477umEipI+Qr5xhIj7qtif/s9UCrJ1
Fl1nyb8Vmwr+7+3HEhpf2Mz2cTEX2W6vki7PdStv1HQXLGe0ozVXvyAdIWjwpB76N5IiKReOoMIV
lKCT+1gHnbbGNL0evVo6gof4NTr9KZ9MzIvXuNdu1tx2R+D3JEmM5XZnhiNFCNrbQnDs6HuK3x01
3bg5Ewl2516mUWw0mPdf8LnRXs9lMI9FvfsOYU7ElCFkPwI52FcqfcEhoW8rZC97/HPisZkbeKFk
V2GgmURE7j+2G/JhSx0AlWCWxxZRFv2e7/rTHYFxYkSOjMsfjCfXQltOSIBFi6hy4R3XLqg/BL9p
V8hh9GVe8NIVvAAPXcRhSJkHS6oyeofex2KymhGFooSQxVNXLEZ0+01E3ikRJ16uV1qdFvq97uHY
d5jKwK1h0POyO3Vdvvr85JjMiz4HR7bQZgSuWGRQOxMTkWxFDADjrajJD+YGwhOdzkPKjDOUk5W7
Fuu0deSEiA74hFBvXyRY1s2bBCCmffcEnqzskCProQxWe7JkGWDrXca4sK2amG4Oe91QjzkK98g5
qA6E8S9BPcu52u943WrIE8NKuTFZasoSS9cFyCLCnxGe1IPKiQ3Ev9VcoWYnJasYBYyXw/uUpBKg
qVrB/WFcgE2+0lyUADh4fSSfBy2ZkRkXFOL0pD0tnOJtoAEVqV3KJumkE132EERCZ5F7IPZCXSyY
rgSAvjyXjm9dPyDb3khdAFmH6UkN5awturgFW2NGWFdbEmZndZERtNWdnRBzirSOh6wtW9+hqYt7
Mu6TtAs9/mRGHzznGjv54cOKs5U85hz6tgnmThfwP3o+GjFILf1hBPl1zvwDkRSWlf9ifbjwKlQW
fcyLRbttNSnImuX1vm60Qk+P0DsBdqsvK8h/pQoKem935hTltdw3fryGUEhxAqdlXOTTzkXBEIOx
4OoeqvjD3YB+X7LH5/5XvUTy4c9Lo1MlUvOuo7BJoRsNl0EmLhgRrEiyiGx/7+hQWHnLiGbeTyBm
uhN4wFwVYL+27BetJpOt7p4g2cZYqJaVUdwy9KTY8RPJQEDcQwVXFduqJVVmgLubmYgvj4/YAn43
VnQZCPxbhko58GMU9A1TA41Z9lqn9t3iL8xqXltM0HZ4vBi2MMMzYqqg0H2qJIukgvSjyl++G5Qd
HT86VGaKbPFE85PhfRsTXOknxILBzcCzVLMZRrra+4oiAeH/cFSY0VFVmkm515dSx8+2VJ/yBI78
EebO1qw8sEJ1zRSKTk11/cYYybgwIAlxlfeYfEFaPsVFUO6hqSYqNH/nmt2lJQ9Ob+11uKjsI0hK
lt2P6OxLAFYqf8aHRtam8L3NnoePFRbETkdTyQe/d/KnOjRTbzafbDJmSuqIQD3rg+TXTvmHa89k
0k+hebm8BtcTYt5ONOPqAW0V9rs0JDGWp/rSLXUE7qP0V+/h3HzuErIHZcxHrBTD7LQa2vGzBQfQ
klKw5STVUtQZJBVch76ctaxHhYxzN//ftrmJ+7jPu4rXVTbFU+F3epQH+KAfwS/sa/cOTDyFumo7
FuZ4VxlR9v9+VF73RVm+7c9v5bO240uX0txaBfNRFDf4kO3MO0Gf5XdLDWljyopbESIaWDkNDy9U
JTCJV9175cHc5EbHcwPI3V1X9mMYix37wmGUpBvecMZOdcc9ObaryykfpbIe9YlQGyGqw04CNO+j
/WP9bSG8y441ViPwha6s6cpo8eiW0WmpDQvtf7CtSk27roAD3+hq7Eu5EpT9kfLnsWsOToQcVTov
ltsZZq2PfieU+4CsauXhZU6khk9VzhJoNmoUIfxZu11OZZ/ZbHTrYE6H40CVwMmvm+Jm5D3cci+n
KbeM+q4hXbs568kjaPNL0QOtv/k6Yof2245WI1W3Z+bKqIgUz4eaa9IbX6NHQ+PQkYSwbzQmTBOr
0dR6JFIdntdtPp98Boz+2knR+DxLDMjVhjobxqsI1/Jn6qr7RqhPoZI7uMzMyrnFpWA8huVwSCkR
CKyhqx1przr7uIp7XB3jwQ+CpnuSmjOQpAuz072gJTM/yMoL5YrhTfZ9qy7OUimTKGa7i4oAR6uq
vCNEypF1S0i5GNH55iaT6ZAV4/vkVCnMyZNWDF+2FH22+C7rGMRfq3vz5Z8ndmKchpddEjX28exk
eXm++mczdj3GQBxri1SzgBI5LqHAIKmjauuSkfWEgCELSJBBquBPTrp453AdLBVeyFMY3QOExIbU
3+TuacEFsvpXJJvJCI39KtjREjRIgEojYJ1xrboKhhGhWxS09jmEKWHVft3tiPthfzRZJ7HK7heF
2Nu0qKX5bFaTvKm6uBekKGSmM2lbHnr0mQj181+OyglX/m14WFuuYr1YLfzYSFo2xIAdcrltbKuD
PdhJw/pcek1MJSWWUU8jENTPo0GfTmjqwjTHCirhjWYrEIjCSIbgd7JKo1A9NldYGjBT4S69lRb4
qkLpuQ606WOWFDtj7s7zvyFZaJUNOXEjaBZchVnOAbSnfrhBaEHLG951ZNwZebLs+mfxolrzRx2v
Qr244mGs5Fuxj752Iq0+Pb0nFDq/MwT/EU0OOnegv3ZXzj4odqCitEnNOsohsEx6nJpzz1yxTeNb
zItvqLbFguXyaPKWC8QfXdz/NpE7PgXsnvRl17ZNoxnTKre4dK3lMIDdSY/ZEKkcLQ2bBw6sUni+
zKH0zye6lCkTPov4SNLkXDkYZpcLkcGIJ+N1tCZpYHdwZ1F985NuSg4iWo56GkB1QC2xlovYBt3f
EaQgyIyDoJu66i61hyk9nxJ4gfkoJKqsPIPOaAHss6ixxlpdB0kMHgM1s5tjMjNIHsoPYs6l+i25
AFUADe1OoB8PJ0yFpClpoWkFN6QTUBQJmPnyYp66/kqoY5ExakGXMeo0aLSIKAE2a7oDVOyrpp1p
2EclUjMUg9qWN3IKkv9nX2bSQNVDAoqAApxLS+eNyxtSAlBGXQib29RctA25jozQShVvD0/BlVR0
cPV5s+mBLxAN839rFGFVuxyfOVdvkspzmwD1LLclr90jk7prnhVedhPzzJR0ejvRKR0Ya3N8ZkPX
8pJTeiLfvNT6DdGOzvF41fHnotCQE5KEbO2SbQ1IKUaVKNNWmzAtiq7Oejw9cFUOGBj41M1mbXlY
k7k+kLK+dTYFV1JGTgB/F15BxrYqxM0F3kDAw/rvlPkWaCvECBQEei1174KajEpPOORTRoG6i6Eh
+2GfkltD3yvlPhGDxSwg4ZWnRfnebARGE1jjEiOPOORtu9tQJ5bo95XscaJll+ybi6JhQE8qQwv+
SvlkE+TDXKSSvJfJZpxxv3HbGtQwCT7kUFad0ZDU/aCcfvKYXaLXA0X4pbI0/wa9Qc6E5pgLCDM2
cXac6Viw+W5HdweCetjQSuKEfcjH7KVwr4ike1WpaecQEYlGmwZRhHehw/VTTXJYjCwDVYaeZc7Z
fjlyAoxOI2Zj+DsR537WKSke67WmkyCnzfOpTd3jkTuxYpodCMqbQb4X+Uww6/ygbvopg12fC69M
vCAQCHlL5PQQH4706/nZ1IiY15C0RmNXuMVzJb73qS870SZLHjoiXGI/d4oTyiAT0JuvOgAzMu/o
oEBzooX3byY5UYB2uCnisrXbE/zSEVBm4t2AhzGFsHLQzghNAvf/btAwB+qM2vrF/Tyv25vUgnal
BAMPxu46gZIE9Yvg0egvlyh+j5oOhXraDA1JEPhsaOYVl+24lqEQpcrIuS9MZf1TsMsgS1klc3yq
jmIH2xlmX2pEGbEBA6OR01gWuWv9wizp65GPcFzr99eJdii3ua4agS+jYT6g8RaSawaPWn4S982B
O3t0h9C65pxwle84kaaeVLIKVAwtruT8yG+xS+sBgAg9Jm8kIBkohIzkRuW+Sc67wVohBac3yDxu
oOqk3tXwzMz1infd5bLFLMr6gxU2tIMztukFzGhptNQql/Hut34wME0TNgwhmdvzje7WZUjzJHmQ
CwdRtHYqwzD38RyjffdH2ZJBSjyufbsojPr/dSgr0tMhvfC+6am6+HTQdISlH4VRCqahljhSQ/Cf
7lFpyKooZImjhRU3cHvVN2Ou3bMiLSsE1YgUEo/zFE6K4CEw86qr3V4eDcwprLtrUJBlCtx+3oaz
zVCDZDOBw6QYNTXVrfhaUQRb6rfo5DzGoTyxKnTUXvF0ZbpH23FPX1Xp/a4VS/oFcqzHMqmuVm+c
JjWahfzo+JB+JWsu3YHfJ9Hy9s37U8BHeba3IyptQkjvlidAG/Qm5T4oWCBkcVXTgbH2QpTHYhJ9
6V0sUzsIuWHXmr3+2o6BE4ILs+bC7T6kNXrsaciH7RpEeerWXVFKCwUXw5AyhpvM0r93JOTj6gAt
muPR0YnP6nTSy9CGd2H18Rg8kjw0AWnAnQAt0K0k5C7h9EtLfmP6PnZZSADLluy6rwUOOS5a/mmy
N3FMnBce5VkstN4sSc7ZjS8W5tIscjQbLER0n165M14AkEpJtx6wr8GSwmyuh3NA08Bs3rsstzJa
8DT0bjf6lmUoIaDSRnsexvL4HZuWpf66bANlUFtZaV8juRCh1LbXXbz08Av2VRU7VlQNkW9u1TjU
gNWOSEoNaMQDLBQUfdwFxYf8Anl32tsTWce1OQTBueR/AYkNtsHiSKYCIxC+nB4I3TNo1zx6KlMS
PsbLylwGTUsFexanST71wdYxUiRXv/r1xaIFrxy0GbamgKOm36byay3lXE/cnUAXwT3fhHXyrDwD
IOcUfY6H/hAWzhVYe8mvSSG50/C7JbOSlp558z46M5PIBJBpjkDCbwksZzQGxJywDUxZR+gIez6N
71Tmhix95SFiAsY0hwDX0tmNPi1QvBRXtNJTEW+bUMAY+WWjuuTHAS1kwFLs6Zzzy3Rw2r+nYY1r
bMMa722nL3h6XfImdSehsfgWUefX9Y7aGK24/BG1C7hKldsZHHPgQlmtkLuPq8+Hu145tYJq8uwo
Xwn53oW5ZolgTpCpgntgU+LGseLa/7WROvo8cXULYGWVYselQXceo67ewPiiSHOajwqNr2cnd9m+
MxSd+aeYT2VmCaAVESmMr4CZ+e5iJUFm8L3yvw7DuJaZiyFCorDvDR7jxFuZaomqseGbitwkC3zT
K7efn5a9ckhPYz4bvmo9EiCo0aGZhTAhAdYuQtQn1kkynrMbdFn2Dyp2yjCkFJRgoSHqnl8Qy59/
F0eIv6l7rvtxseVICSuLA32FS3zzNnkzrUaOmFzQUhJf6sYmNYp0hM7Pj3V86ugoIaCdO61nYQPw
zAerKWuHmt6TsD4zfZ4pPiaFLUf1uq7vo0bdDsVEBAThWxbu1cLNajr2Ls9dWFbToX2IYdbOsLSq
8TJcOCCgTRSkkZdKLAS7TQHAXGEmSLrclLdfp5U5a9RAIY7G8Ist8b5iyL88T7V9ORQ+24xqwYQj
KN2JXPBNjBREwRTBrBNEj/7KvDKqkXW+9QbkXT4tdkcZHzCSj5+mKGZTWmeB5Ljq0xer/HDN7r4U
aWOHvYnxlpvXGnVto/QM/tqvyrzmrwg29wkkTXGSCgeJYuNmCw5kpSM6Hs4B1Dj8PwzesoaAD3Ay
zkHEwVnpzjprXn72M/Zveganx5Kx60eNDw7/1PALgKO3FKqxbfDGJu4IQk9ePMEDVYpICiD9tU24
m7JsOLpm1xRVx5lye2/MTH9oRcwwJ1aSJ22FquwS7av3zNHfKEPXpEPOHp+ymTo6QFJSZ1Chv58x
0i3fWtoCVeNRYLwKzPydrvhppXvZs8ec96P9jHq9JaEJrKvPMCp9yFeoVf3PW0VDHsovhJH7q1LK
cQoR9P2MHwzM7yNqHdYaBy8rYjbMJuchnK34bSiKREqKfo8DA4N2Edx2MJ+53AHSEAs1MyyvMxjb
eM5UITrTUkcIKiy7xWJBDqO8DOxfxbTlp1c0gsZhnn0K5b9m/4fJpmppihFUqQuyEDv7IG6IBu6f
GLmdaQE65NOrQu1+idIXIzx/i02qxzVXgTXUZ+mO6LDBrI0uqF+3P9DvdXR+EsD/FyZS1ehPo+OJ
IFtR6vq0Fyt04Wh1CdIOKOvDFo2HUssLqR8um468l8GDo4dVxfgUGo7TivSYs7XHE5EWz5YnYxhI
wtTB5orI774apsTwkFsebEwI7cV7ZK4SJZWPLtdSDCVtMkLmn2IJOTWY1tfG6q361xIMpFzDFaYc
YUMW/ECbLtiRbBmTs8OdQJP9NWMHro3xhwyppsSLg7fjHWKPaz7Nk9hHc4hWVPn/Fv4zQCevErom
3pCMLtnaU9/c5PZ14Qe6b4S7qK3tThgB2dGqmDMifdBH4DNVy4Fm+pvo/18FhZ2N7qs3yMohWYsu
gb6N9RVio2OvTvmkVSi9ptb3wSybEftAMkLW25vQe00QShl6sQl9lbsPpWQp67KrxOplxzr8dTiF
gKlSSN+i6S/SJ3wuGYRxjMhKI9sA68CDCcxgt5dWQGuF08/OdWZ0cF7nNjMcznxxIliyFH9euu2n
d1PPwKDzLtqH9cRNFa2Nur5QVizanGMcZUnEablJfkW7i4NtycCyUWIF8kiLkzu9zFYKlfCQRb1c
LS9PAz/W0TSCHOV+bU3PZusxCRpHNnB+jrAQ8dMVZhgRuxIo8tOyb0a0i7VlrOjdwTxGFIoWtnNx
9UrhFzGnrCYcuSt8U9ohIcSF/H8xwbiWhtV6OdQU9dqo9XO5F7FRxwnTRrVeTVjqU17xqMyGmZvz
AxB0L7Q7RBoj/XK7gbElWeITGxY8GUeVTWFOFALbYMz+t8QsMAUePCRU8aO+2Lg1pqSNaiLcyICn
TcPHFit9Eafos9MnJj/ygcKLmClWIKK34ZpjhICF+41Gg79HP0d74q9Pk+vrBvnvf0EdQ+jLPi4N
VzU7iJBjUmEOJujevVlvZ4MzmeM/8UEqwya1jAECJRiNAbbI9W3QECii5Zz3rVQ/stFJvjlKuprT
pTRNxbxx8Uuu8BbHRnZLDiC3Dfmkfa9nJdbNzBJhmTmGsSTqFz4FX4NLQ+xqkzVMCJtUCAmDvRwb
BsuLSE7QT3lVkbGJwqtWFcPJnvDBk9vmmQE8o9qAAanhgXChcqe2+elIsCJqWDXcrIBF/a1JUJuO
CdlL3qowQXyI9cNMQxzWFGvau/vRa+bOAFmt8RLgEjbFOfnUw0NpK/pNxmLXkaeRBXW3pAPGTd7h
FJR36F5ADInzORF9XHYB3pvhju7rLkpySDl2lM2BMyMzVLGIOUL4by2EQAYwzgSX0WWaEcO485Hv
O4ibNTHGyzq3HFoN2PrCX2KrO2WbVyqszeorC9ICtk9X5nt7BSUEB3LfUcZ+Ob7PlhpFL49RxZ04
iUKv2xEb/TBdkuyNyplhSIJu7/+CUHTwRX+me8BrBTaCPawZbgP0ckje98+R6ph5f7ePr9CVXeCB
2+nPQ75KIQcvgpSQ+TWdSBLpHtK1IxI7ycJg/QFxRbDnvUAEiXEymP5TfR1sHYtzu9ACVXW/IwyQ
jLfTiLHLvvkvu/wfFBGh6Gvrm/WMsrqeLjhEaS1vGw+/snf6A91SN+520BZ2l7vKvNragypH7xKG
Sn7PhSj5PbVw8B9niGlTJRUHnKy6ks6+yCZZTvWhiT0dwGPxyuVCL2ADukkGP0VZsNZI8y072vOH
Xf5eK7x1nCcXPFpRiNbfbRYDG574wGqd31vquUSyhmLngn4UK+gAY8CUwSD80KPTZg/Klf5gK689
Xjv//MVFG1QGbNPzL6ITnHyvbPzZPnZIqXpfVhLYfb8FVkaMITJqiTa3wYLjqFE7Boua3XUwJzWT
PrB4/bi8A74L5PvnT12ujHIcwA3z+N5nU6i4ZyaBKIxN8ZKiwXOu9KXkB9iR/Xhe39JOceEag2MB
Uzx0uFkymUENVuLteQczMYKFBGqnq85aiJE+fPRbRCs9NvOyUIXb7kHBcGYORpE1ysmKhH6oANEc
Ewi1kGNwLznVMkNH0BncxJ02sEHmOGDETCnxgFupGfVeivXy0CFAjSZsYLMje9zarboNzXs11XtO
vE+155avvueEO4h9kGcVo/BPUlyDvG8DRm0cvq9W+u/90bh4+OqGwnUPWQJXGRJv4tUoPKPikjcm
MzC86p5zBsk22l4gFDvgVXF6GYQ71bvzxzeudE7/aj+8DECEHDoRzBtVgWc3CowL/9/rl2P6CaEP
6imG0AxyS1lkH9H5D440w+DmLyPC3tlrVWg5/qv42lWZ1/FcHRBIGV32MYUxzC4/CmLbfV82CI7s
LcSKbKU+U7lHsoBFvpij5EQ6DEsepkSZEgbLDsSClUCs/BHOCda5HUXnxL4IpOeiWvbEtJixPasz
oiSg98G/LI842iQxmlvZjUIHRy2wSewtQ7rIKFIjXGFseZfVOmfOX7dGKr2f9Hqqe41mUCVTxyv0
27rjOmXylBolhHgi0UIp5tijoF/PCaeKpBhyYBYlBSM/CPeojUMa5Xp8AihtKfdW+c4oF5Iksk8W
BBt+gHnXKmN1d217BQ9UzEFMF3AqwKnXXKBmlsDP7zxCj4Um6RHfrwSgHeJ4R2fZoAwz+4KsLzsG
n7KICKa0OKFE41rzkiRH9vjgmbZZM09hsPbArS3lKR/H5tqqFmCH53hL0oTl1hn+I/4vAopdDfkh
kXpS+Dmxgm1UaJOkthQiAG3KXMXC+kzFGul/O1olA4zLxYiT+x9Q/veuoTkW8Wk6viczzYz/++B+
d01VxL8ZPPdy3CFD9temGt/NSPKtlUd4XEFJH0JT+SwHc9jFqdlxhp+UeSOCwdbJUF9sS0XWNGeT
VuTQmQK/1lhKF+iJDfm9zzG/dsOU6zGOUENHH4oO7Icsec3nhlkYclZM8xxfVH0IgQ4G5b3nL6G6
XptN9C7WuU4kQICGP47rFCRZ1ONnre98WGMT4d1+HbYA1OHNcbL3Au3aYGjm210nXb17tyGAZIxQ
HWE/ltlruwbKxpyZ6m+kHNNWfQ/CFgrzjip7nAKNvMIcN63KRoVGbVZv1HNQPlBGfuX8DejHcwDA
/l+zp/iJuwL4/un4pEyfiflgbGCD7cevvcvsj8HfKITmCAVne2mAqMF+NrrFrZjouanYpdWjsQJs
0pDfs+2fitcNYxGKRAmawYowj25TZyhW8Mt/KRp+YH9VS8nhpWm91090ufP/2LgkHCm4vftzBdwK
joVq9/ZRrnXvBAaC5HkI68btlnoY27EkpkKOlC1DHkbtOzLfdKpGQtTya1RLJS3TuA7lNM600HbO
iyWs1F9uhJIDCiwtlzRmJoOEFP/4s98Y4KVosbvg0YIiBqetEtYRFWMD/OXUx4Y0qwZd1GcjA7wa
K8DJgaIS/HY1pGD4hQqY8bphtwO+MEbJXSq3xO+mFuUjk6whRnJH+TujqfujV5g1FIEgx0JB6qYl
UkCsR8E/FqvI2KmIm6dtwiPX/CMMNF7oP1X5HhWjEI6hDkPsdJ/5Hz69WD8660lgnJL8nY15O2gL
7MFMBIuhgdzlg1mxkVdxNH40TukdCL1090Y3WZX/h8U0YYReeKQw6D+0gAXmL6r+XFrgh44E4aNF
PdybW4eDemDaWFZjZNI+2HLE/CFdsHX+1VWr6vAOC6L7mQ/Xhs71DOVe5UKir1O1hAK10qZrd87L
AnxjyJHWDwqbpr/sv9hET8/WJHMqFejiUsEJpStDW4VBMnXSCk87cSmo4Qj2vBd0X6UaBXGbYcYu
yABj6WbjsP/+r6Ky5TRAFpgcuvktt19iYBz/PKCAXVel/0JZ1xvLZh5GYpB7c3lgMP8fnBlzXiSL
YCPo6+Jx+rynhLILjGeKHpMG1F1GVdPxK8XXwm8j61ocfgrutaawb+vW8d/O+PfVvp3ly+EI4AVT
B24Jlc+oYQyZ3ycOOb6ztGcR+A/yaMoXVY9ts0bQfKkznPpyuD1dLC6Ao7kdJpIwbD5cxdvW4msQ
6Ld7aAOMIb2WsK2+406L8m7IgJl+etM2ntjYjZ3Pr1JBMaruhssq8IA/kL97kttgryTJGY8Peymu
6mRusgBs1nmkBF3h9EU8HAWSNeHLuyKcZ/xl/MTk0rk4ck0f9vAJt1hqdiMQR6kKw4y5cgRMof6q
Ht0qMuf5ViwH3B1H32MZgET4STrwH845ItB85do/gDG+gq2pFUmCNcKfi1fvx/6MInjwsRhcy1l5
0uwghQf5Cbtsp/Kjr0ENCjt9NCT3Wmy6QxMJ9jHLe/A4M41aO4l0JwfhUleraH751cIsiHLJO90f
8dnAX/5/9OZM4eePci5vWpvZPSuX6/swpDte4JW63t8iV5VgYtprW1u5MqEb24rGVfSSGtw68wZM
DIOlrMWFs7pLZoulojSH56N/sBCBlNnmNFHXfbx1rT5duN7dTTihnYoNfosAUKHDmjKkxHOKu4pW
1PsEVtLe61JTKx+EKyPRtuF2v+E2P9gp711KoUttoG4vgI3Qt2TA8XQbPPEVejHcJ1nSmks04A+7
JnqOUbQaBxJkNmFY1Vwp1R6jcZrg1sZpuuucCL0HMhZfx0fefJvsCVX8vNNXd0/kKul7u9ReAWt6
pyyieXAR9JwKuC5Go4ZYDqgrqHwxMLDrB6pM7epQYFStMZLTv++gcIyj8DtkfOqRJtrB5CgJ4abv
KxScQ9kE2EwWz4OB+p67xHOyZFj6+q4AU3GqF/kljHSoqtu8f+lcy3W52AziWCBCgeMt4HpWoHxm
nfS1wl/Gv2LwBwGPbRkH8mfXj+hHCI8oev6HC2Jdlg3Dqe0naGBjrCB1ppLYg/zXqzdlVVFU6IGY
e28meX9D2xx+0wySXtYHALlJHTN/LQoUBJJ4c6QR/dRwIkOX8/SENowdk5F31cmaI53QRBxek4zm
hqIcFPCiwJmoxZAtj1muFVD7CNQUKMl28ACAp+NXHtrWcTHiQvwiGYl6yAVqnRLBSymvOUQ0W+15
kgDpa3rWe4PlenK99Xqx4WoHsO5ajw/vzZRIx3RacGZfb3dhZjlFtrU4jaact4p2Rhqvi+/XT9bf
nnPPfmzyv7pifvAmIZh3+aIKPXY0OX7Dkl5pLhYhNOY5pUqQsmVwnQydZNXqNua5+G9Srwwi1TRk
BZ6yLb6u48+Qcv4tsu/a+vyXHonxnJQZ0LGc2TFjc51ghPTqNNXcyUWiEj7oOJL33Api3kzX5iH/
YfvAUKJvuVftm1EViPb3HZRWZebYNlhN5Sh1ZkjzW0uLRH/11Kh0om0glFOYQJSB3AWKeorUq64p
27K8lYo11Nk19DXUsbAstCS0qof1G2g6Y/xBAsschdnrOVV79HTysi1n3+9DrwOlDIvOhKBBSkx6
W4d2PLmH9qfinI8zdF7XTn7bSTKSiVOgTm/r2iOnxDiOvBWME9PJ7i0qxYqjdiJXZ+T9IiCWwGvp
X/FJkjLiIjOlPjxCq9vy96MAntWZyNPvDWOxNAALq9AI6MEyHzBtIkOD7lKwp0QzPmQvAmL6CrHh
0HbnbADAuhFvodbzBNcUtcM2nttsPhxLQ+5jK7/pg8r7rWDQ1+CbuuQAO18kZbLBY1u6MddEZi8i
BAqboehIQLH9KZNfxhYrsvaxotq48INX8MmXa7BymcaLpvjt41Ay0E+0sN9Ftg92L/UK8HBzyr38
DLVxvwzFTc+6jeSsWlm4708glH+hUVETCtO3VlT5syx/efjkRBgwHLnXYKuyh2qyxf2UsN6q3uyG
N/tbdmhNlo0EZFHxMVjoEMbOTfYhrd8gXPHe+qNKHrabkJ1txBHgTH20LuLCHnl905eUSuNalmnW
lqf1ULZ79dR0ncewrDPpILv3SolWZWkeH0Jk/2kgfdLuC2N9keuzO5phDcSGoQJLeDZ/qQhiDM1a
+aXr8V2xaE7EvK+DIPvi3CgLn0pjUwc+6rE62qvJkNsxKbiJWZUcz71pKSXwHVdvZab320kvHmS1
VA4Sz5kjbpHAigZPSsH6LgOEcDYrZ7A+fVfWwaq2L3eGtPx/aC5TON4ByTyEvy2vf0lfeZByywWE
abHHQWMLzWGNfqSUSltOcYee4EIHqSKXHgZgew5MVvoO/yfWGY8MbyDFQyhblV6krz/ukELZHDC6
vQ96CWxIQgmRHBVNSE36L2P4h2XdXhM+6MNwVy8Uyo9ORq2tMA/r+B2eYS9CY+QV8dN4b4R7+QIG
MDkhxZkuEFUYlqIv6uh8NO0xQyO3MDy0As61LTZ6/t61e1GCwcmrJBlJO0qEduHykO/s8fNlg9ga
SsXNwsCoZyPR6hwO7RPfl1FPGybA5lf38SQ/5zMNm4uOW0EwkTF6WUfvuBgOp4XGgHoeZvUf48mU
PM4m5tMEFQC+JkqB0H5o6FoX08h+9n/5glkOXXDExTRo8CFSezhVyWjt6O17pOG/hvt9/JoxIYxm
j/pEJdyQCP+tp3HbovEqbjt2yrSz6fjcGvXhpgoTaEc4X2HDAplpoAJiB6bs6kTUtiXp3Qfek31h
dweT9T4BQv4oPgj1D/YXFc02piXG2BWNSMEt7K6ngsIlrlUyOjkNs0wI+SlhBnifkwahLOAQtAlq
GKUNAfs2aIm3HLjcpClx2tlp1g4j8cnnBYVO6ZJ4OiC28SkPAy4uen9YUpPBJHdsZt0TdRCtqJgA
O8DFAEvopICgDQ3uXb0+Z63aw3RohBAL+vV/ejgWth1YunTiIs1OPzGgyh2sASUg2IabcsWaf+C1
JzpekNKgfnK7wgdLA3PuPyq0zTTWZju32pWRrtZlm57S7c9V0gIqtZlMR/pe+pshorSqeyVSSAxc
IRrvXwhD2vJ27m+do94+JlnbqbGcrdHWMkbc3EpaG7m0pPALQsNTAFuWC0vW+DJUQmIaX10uD66o
GSp/y3ON9ngRBVOeQgQHiAvtlMOuF+XDQ+skhf31bdnrciNfKh2vBHQbaq9GB2VKUvB6nDcKe5Ep
md3nR7D0jGGl7mJFU0u87jvjxPWf43jrP0w4k5Ar6Ile8CeJRrq/tsar7f8Rn1GUQ+PsJ4V7JKxW
C2lBzT7AxcpuCs72z3PEZCvBZVC3chhy1v7aFp8jqEAL5uo5Wm80XJvErav/X9PEPuUDsu94tpJc
PYPbwTTMKbemqM4Qzw7bXMWzSQWM16svJBmpTtM9GHW4F16/YdEhpn0cGSZ4uI+m4xxf77+5EAam
AzazkMbA0qnonjmnWNzyV6aJKZlHCg3cUtByQFBCOeBXT++s9nPcqhCn59uHdYuMR8Wzxg+qcz4c
nfS6G6KcLRHqgZT+nY6+lAnAZCW00JOLC15Yn9bSMfLKP35b9pdOYXPKsOc5oTe6gAvqWXJm+6DI
bCItBbDqwKawDMSAP9bUnMC+tdEPnDTLoLdxVgiXWsYNE/A9LsErMSI9cgZohncO+QZQyB6Bqhax
uuLkqxeUCxGuxAKouoUtBDMF7SkeK+gsR238rDQ0yQc2oR/KL+pA5bBp68f4rjFnb1LdLqZHkCIA
4HGL6PQq1IVl1mo+HANWkktrgJnQyDUgiBqjE+A05ItWuA/AEinPglyRC9Uc5kKz+w6nCC4sYCRJ
cIyZvAwKOx9HaKivgsOROsOim/rOYjBi0g/Amhkli2xF2xr3WBixFpG0gC+mwS7I12yTVqYvmGXr
riwou/idFz2H72CLiCl3qpcpvpy66rQas72IgIm1qXC+9+eCAsXyyrMlG1jO5DrQrRl31wmheB1/
gyqiisEVfoePcn5LMakrBIF+vFIqP3QK6SdoUB3Dk1h9Z2YYZ1QD136FO248kNX2WOG9uRx6scSF
OrBQdSOtxEL2koTfC6Q/Z7bB7A8er9MnycXM3LO5E8HvXltoJiR4dYqBkf0c53jwWqjPvxOqTtGL
x7XP7Mm9wQoUGjTtbbDT4RceqxHqfLxQhR6mhEYQ3AlJoBATiTFkbPhSLOn2so/zHQm2KBt4F6++
NAIcj5jqEda5ib7766B0/kX6FJb6qnK3avsRq5JPuwaJfuKSt+EzRUWimD0iTpTitBYI9+0/joXa
5DHyHeIcR25cIBU1MqGtrPGxtmgsvNuVTyjAquPt+XESaKs1X4ewezMVbdHZUb8rHTRo01gCWXn8
JASK9nwub39S4q6UorCbui9QQdn/k3qzlSsNnNy2rF7ifJnRgAgoBn0VWkdRB0pr6AECwB4S8M8d
ju/nxVysDf+4hh69kuajrF+5MavwSPSjngYNJcwrmtNV20tznX1u+Zs60vpflCruQEbBDYniUtY5
WFYcWCNu9bQvkcm8WaiEXjEuuu7I6ZqYhYf4kUNmxi3vgvYFkVhNtw1/QWhI2mrGblftzEP1gPG+
O/KeBD/XHswW80kUgWd660+laKfdIxBceHdC4Pyd/vaXHMtHvF7BCXQYj9DeOKsLReruawHqMcxU
+OpyIdoIGUh5lAEZZdUsKRDk0Xv4bagQkoGpu84OXyZcRFRjqH6cK2oPU+Wx+YlIhdJ6jq7W1uvv
U583CuTCdMV1PnFJVk8tmKFnCMfAZdipLRAw0hzaVLfR8Q6kxJ92gsBVYOc/N5C7Pl6Zmc0hPQ8Z
ng26tef94rYJlZl24crFHIw4MeyRDN5A7sjXxzPhT1dOgf49CdksuVeZCMl3riTdDv7NQkAevbdQ
6HDWuYnSuz/2j9dPtsYXt7186X6T8AKWB4r7Vb4xzHttvn5Vef8dnJN49c/rOLYePvT08RvsDMCq
T/VVJxOjqWYbhsRRF9fH8ehiQrTAM3OXCJnQb/JUFQ+DyZL/nlqPNYwkswpBQDSFMxL0PpXL+wiA
l7P4vTYZZGjBihK+5z+LeAk5AnZvG+ebDL+Fg3u6ZWiMYgZ9vecIVJ1rYgsjoQjbAt37inm0OaEq
4fIEX3yRwahoU6/fszQRoe/C2G3+6u5ZyUVhW2Og9BNxf8bN8mvEO8QdDrpA7/osbl94ezqeqWGV
Yu7KJ8nyBE41bWpwRZJl/7AwWDAX+FKxcpquDbiUJLgMSH3Cb7oxHVqAw16x8K4cJubuf+GQujT1
34rljh2NzCFnBBE1itxcZOyzD+SrZIR0xZjs1YBgps+VPEU/SR3Ve7BDO0qb0o4r/rCyq3jalrlC
UUPr4qewG7L05vqRxAnGF+ZB/Y0oK48YiPOEYlhWnQIcr0vJ+nDvTrLXCBKDis9tsG/1YLIBTdNo
X5XOdvO/RV155pD5maUvbidAMdR/PDCSUKOm1mE8tXdC77QO8uIRk2g1bWnQtNKCJQ/VN8a50tc2
aB+0C4JbN+daxS417f1uTkBCMG1zNmgBRzywgRmS5o//Pmfuz4Iv681lLTPcURyfHeeuY/66KjOx
UJx7FjrZJS0r/fnek2FKR3j9eP0zMEj/q3l4nucUS/foZNrPfwvrGdBRSufrO95crO9iZCR6avpy
x4fcjnOIJwoDAYMWKO8zn0BezxxkspAlxEHjcnpeyT8yRpvrRA6+NqfIAgOWq5GWGMXaVJiNyv9y
COOcxM4y8h5KRH/K15IjVzZ8xqOoFW2GVdcNXQ1SNh+mmIzQFRmTMUfylQ2LmCe8wbAvGQOtXA4v
3gKVxyZOeS9f9xDuJC2Q1hLzkVN1NmjbOAQVNNqGa2liiONcA1IHrDKaoCJrf/vEXijyggE6BRBS
fajlUzXXV1UpqS7UgdDZqFNFk/QRCeIQ9vii3cxf0HStUliNBd3OytIJ93Pyvayl45eZXsZBpgZ9
KqfPem/29QGFF6zEQFnnqacd4SYUWexZSEGtsTBGgEFINNh5OGWw3DLTTzXqOmDe2ha7rxClSt9J
UW5WHw4/HyieBgPO1fIeXp3Ez8u+OfGJv7EnsnG1ppnUQoJbJzb5kz2A8ikoGxGEW9Q55xNUuGeg
1q/eQft6wXXoLpwxtc1EdzGrIqX3b93cFflsxjqQHI1oGNkePIe5EpV/krRuOQ6iiOQrhbZcB3lG
ODME9Nu0zUpeNDd4FJBB1u5LIIU/OU+Vsmuumxu9rpLtUMP2RMPQDJMgZbNPxJ03Ty7ZzS6HqjeV
ALv35Jq5pMY6L/oKf/hhYaUQGMW+ToPX9EPKesjk9+jBmPzcCcXPyogbvYk9volnVQkSBXtGSE/Y
Vn5SGe1xjIpERcQHXtYRA4w2SDvIfVASgLRYjtWylT3UEiAAXK7Vnhl2KW4naMYFxcmZdqAiTaU1
8yVXasTia+yx1raUTGCN/SPUnFjFHbLi/ORoMiO+Fpm0qEFlLzDgtR9eIohy3yjDQIcqRYkjOKJH
5PxA3vgkeXUj2R9wM61WsjhxjgkO6gDavXXEFh/WdA0yKGWzTTZUhXPe6UBl43SA1U5nN6zm66Os
1UTVXIY9o1wbhyAikAvH6DPg1qzWCBm0sxfVymjcvuAEfzFhNEKWbhrBBfqtt7eDNIXD94nZuYhq
JXoIpKekqtbDrBQHIDbWQJ/+w5DF42eiyHFCOz08amq4dMKHIPeHSE15iy8f5GeOiut+UFl1R8n7
gjOsZnUATyi48ihCUaj/P5p0Q+uK0NeLC7WQgkT826zig6TopUE/cHjjBfe8hp5+9EbdDWLjpwwQ
SYVx2N8B1S2nIKYODxYxDpqEgq6kC8DF9IUxDeGz1UDYaFE6pNIJy3T8tBHteHDIUgZS2u182rgL
qXbGw23fY3X80stRPsrTm7k28G9J1LVJteuXyZUgmpEUD6DkCIy7BK2/GGwRqyds7G0JksY4r23K
ApEdNtrf+k2XkPJCM/hgLmemH926Ta8xlLcPl9cXbqjDiZaZmbkw2MUBdDZ8UhBNLR8MzAwFbLfR
q7fp9f0LreDvUGDu5kXPGYyljeI/LTGVVr8E68tDKk4ylA9Ldv8o9OR+RYCMIi2Q1DP4sXb3vMLC
+DbfwpUExtcpdHZFvGRdhH3Y0c7YUrGz6n2gLBoTNCSM8KA7ZdCddqY+gS0D2SrqnYeOKKDw4dYr
PLhk4HovyduBnnnLLzt5OPkLFWWJJkAweX+GzSie2sraBvz+ufCVWMfdZpkWaCfiqzMCld7Qj0Wd
4nuhIaVodHWxHok6fRi3nvus4tqk5xSanA+GQTdUzg3C/5b98/w9z9uIw5jXl0tK0fDH0tGd3aMg
C0CPf02PXpWxeNXVjYC7zYfsMbhEYIdQD9Afiy75sUtunASuikqdSzhW5nVINCJjuheg69TIo584
pa3IMmbqdCxQydbAgYeYwCmsajULyaE1Hku7VtO6uWXU4s9qC95dgVnmfmuUjH4yFYeVuru7OXsp
vw7aKClEMsEs74puB/kfiySERtNj5d5iNSQ5LV3FZIFWm5XZqwz8N48kO8qBeNeqsCPuOJLsh/rc
Xa0nEudIkJIoMYG8ioC3gCPe8zEcoGCkZF0F83ymFuLl3ODCZsMZGKj71LpvxdEbW6GfXMVe+Ll0
4SdfoaIVe/oKLEXqYcJlxlVDugs80+tFgOEU8BOj+BKxr6QFVFZ1iEWeDT1DcN7ZWv9+OOZIAFtz
eSBA3ms5Oj47FW7kwDpwBMTyoRfHnTORLPy3pg1mhzFV3a4hSIbIOnC3sXWuapSzsO77/YCTxEHx
Sfl5SyD7h2vBLjxp5TTTIh4Jme2buDUwVx41XUQ5Ts6DTXB+2MVD6ZMy2SEMmArem60+zIXg8DrA
3K4XbyG/NWs9AsOaStip2UsSkhSXDjncif0/5cP9ElBMc7j3NFOkvlrtUxw21WfV5fIIimQMz7jv
Rr7OytB1Aroc6uM1S3p/IkLEEpSQ6cH+cCu1uIOQrI3Dw0FCRvNI53GZFIvJui66aABpKdaxG3lY
POiCgo2qVsL+6f8KC1nUhnhECIBrSb+yMZaD0m94FbfK/Qwu6pSZwDLvKjOZgI2ND64UnsgHkhhy
vnftOtgOuSostVeUFTUxyEzx16dWnA039TUaKQRRNLziYCdcqqtRrZc9veohxDN/T7ciSKCJdY2Q
qA6qngfQXODfduW4ajlK4IbPTlBkaKAq4TjYB0wXwHPp63SppYaJfwABW7IdlceJhgnmXyB67wIe
TszRFdHA6c5wh94YGif53zVtEofSPYS6xFaH5kKpORp/+cztywfUXf/KnKMdbPURHqxvlImpkqJq
syW0LDjOolipiHMCvTigAf5VyO/GV7QsrfLobUcf9ld7Cay4Vztl7pImyT9zud9t8AdI0e02diKK
oLeSdyHapV3bRqB3N6Yxtamw0sqXdmisDzCioyJrSQzlQg4rS25Jb6qJ/YiI/6N6IerpKNqUKfU4
dwI6GWdphMtNbjN5EPObEla+102cKHwujKdA8QvjMn2YJSHdBX5XoSv95ltSi2URlUKuVAiZ/sE6
6bHs0TGvXozCOYNZVmm4TaO3+uWraRLn7fWBm1hLV+suehf0IivfUqvRAbT1pwfSzC++PFIla89K
HqPOruUkoisymE7ov+vjan7xJHlYuymNF0M63gUJgvosJzeNZ0E81Q6e/AxkWyB+qM5xeRXROoU2
6LIW6nJphzLBQjLsmqQMySA1EJv0KcxuOP4X340hTALNW32v8fOtmdzYd94qPCIQV/HmncYO1SBg
zQH9LD3ckrqUc0xqrBC+uDhdbYwHDhg3IbhFGWP9dunk2Q7N8rByJb6f5s8A/ujgPpNqK0u8Voof
Mqtumvprqe5sElID0CEcbVB+fEsHLdqUKvTJGQVF0BW3DQH7v9lQTYgOziDnyw4ctZctkIqyBeNh
TgJQq05CPgvPIpmMs9ThbOHBoJXEnAsvyEK4zs62PHrKNcAld2mi3iPIB4Pluq/qCDUKoXkV8jX/
EmaLe6YjUz68O07kdIxBdKw6EGJ7s5Iz2QaqD/THjuC3DI2KWmh+/0xbqxH7s7VfyE4+2/ZlRJDS
jbEjDnvEaihIjIqYm/rz9KnXkc2DJGg88Fgc3vW+l5rVlPDxAtjNrAa45xihm/E1pW79tzdeBidU
JQzJSCAym8Yr3FTzKZLs4O5sWUz5uSvTeJdw4QJLknOtLr7AicDvFeO9Bdl5Pq7XZx84+iflTK6Y
xVDywV74doETil3sdufl83FvGsvBw22GnJAf7NeAXGzMr5KxDEkyR35KnLsNFX5p5qQldI4X4sTc
3SAdQKsjgWYjcm3z78dyf543oH10uXI2IQr5lbhLljO03AWrxOP0RScxOLcPUOEqn0zHjrY6+pQD
dwuI3dAf5O1yE/yMZU9S4jqQDB8qcvpSZkF6BKl6LnFK1juLJpKNlppvIM3jTWGtxyxiJeGNWIXt
xKgnUD0EZ9fIYMY/v1RwC4qzMFMHRCcobt71EKAWKY68NMsZxvFzTM23+ny9isGGdEisMnN7ZBeE
wSd9kpqpQr/ZMyd+us3yn2EanBit4NukkU0JJLBBvzZdoUos05FHqrHwqiD9ERLhHbuKQQflIBha
9mgb7Rxs8gwAtv2hFk1tjtipOz3XqtMU0UH1n5RIRS+NQoCUMiBwR9Oq9j2/hIAIEukd95efiq+P
HGrzzwiNjXsUT5MbSEqvSaGMwnh9vUZGOecGwBEQ9u7FvCrYd9bwKDmOO3PglnDoXoXWt0pyFzNb
XB71Kmo4n53o3kLWboq/fja787JbfkEUStRmDDiFDO+wuC7KVURCe6kjYPmMahB1U1VuHIbEUS7R
5oU1SjpBBNUowr90dxpI2D1FGWRY3yU2p5vdApy4uNf3/GMV5u72/qrShWeTxiPkxP4kLkjUPgnQ
FIEOFyNSyxbTDJsOvvmraDiAE26uQjuDg6nnBlfnunsrb8qVFCebGb3YeG3vVdzCsVrkjNq0Wxmz
8h4BNwMUOM5owlE65/AowC19fkAgpbhc7dMuBJ02l/n+3aioYZF3KHetTO5uKKLx3pyd3q8NXDaN
txieZW+0zIF02DApRY9dKHDWTF8eT3B+0ypLpqYBOPXEFUuLiJRV2/Pf22lM3CMP6r1GDgy59mdq
7I1AHH8N8redlkjewPDLqeMxX/1gk3zhiSfSgHylNTo8YF0KdKTCy2g/Qxb4PLFA8cOyJvqqdNHr
wSIGtQvErNXRV/beUFu8FzOZ1OX2cZ8n6Vnz59hBD2n+5Nst0xtGuTNAAGGBNaOuaRdcJlNPYH1w
zVLmONkStCI/flJzh9311rYFuEX4i9LilQpM7nIAnfZpymTJ6E4/vF7cHCA0Hm2Nbhr21vyGeG+H
ztmHea4T/eRr0NFNrjEP5wDCUrvgn8RnlX9nH0Y7fJB5nlADmTnvJeNt7HzkYazWlh4DnY6F1pGm
KUUcmdBJ9WqzQ4s5FVb6x3VwlAYfV7tsoR9WWAY4p0YZlgZ6e7ULCsj8mGpkANLklwm/upB+c0w4
trXTS/ti5eMkp+47554Hkc++NUGDnWJRRXWHx1BGCHtzG/1q+MObmfbMtxkWhatwuR9NTNZ9T3D7
0msrnvfBtmhOv1EfO5FaFcOlKVvkVI+wMfF8LGZw1NtGdzzAgo3nJgOGp1PXbgnfG6Fu9nWr1qXV
6FMi07g4jxZUBKQDNaokTb4gnmKc6mFUYjO0fQ5l8GEoJAiW1/TOZNbD9REXTpkUqxjCufEAMjbL
TOStGl5Zq5N/109xPOpKK9TrGMnbmfB52z+MvkhjAoARd6S3FXreD8AWaYTpG81tED+fIxzzbNO6
q3lw/al9K6QE8r8k54jf7Wz0dLA2YtbqkF+LSif07X9EdSQK/33Mvzqkc9Fo0nERR+bbkarlykMp
xcp8+fSBylfCw50zONFrSVi34YHu+zpLFpVEOn/2U/qf4d6zQs0NG8fMemMUJ0fYyKFq4H8SJWVX
WYkKqtFwXSRewhIStYgQta/e2r0RriVx5dvB8dXJJmGV9fIEy8v8+ylE5CgtCJ8YP1ML753AYAeT
dHIHbTPn+m/amsHPXP1lxCkb1N9BW44v/fGB4hwqm3pkRrC2d6W0S3Ef6K1ZepG3F3rly81jLP/z
jHVZDXTJidN7wonDn7lltv1kD4Dsb+0+qUdOV3S3Pr/zfK9cmDsKu07XYmpiRrdXvhOUrZ8bU8N6
1n+YaMaCVdkSjhmazSiEZiHn9HgzDlkdIfovhvE1pV8O2WRKeQLnExSacoOL6oIw/SlzRSlqeZIc
DdvsTAh/8go+Z0D1J/6KYniFPs+pvsyekIfMQo0BxdC1CSgIVK0Yw6kVi3OpFQ+W+nARJwA1sp3P
su4jCwPPOUzDVKIswXf7L/L3mGeB2KMDgNZvXORoustzRaqPdULYCWrCXs06K0ddQTR2ft3StupO
Wpl9IRHsJv+2lqaRVbyRFLHY+cWK5F/X4Gji388/Gbqro27FvceLAH61rFS0qKYnvg99pHJD7zYd
4OfWALM1zqkoNshybmvf+4N/FkKVh3NxNa76M0vh7kTNAWrIo1GDqzci92xoMjTGVUwnh9sv6nPX
QLVX3KvFOyepNySGieIU8Zw6BJYvkGcoBs8RKijY3euWmL6l6wXXp8pdptnL2TF7ytmamW6zPq91
OtSlwMvlQmTvyh3k6qugViBDfemtaqWIANWvK736dnfbTLdQQUxZpW262AnKVU4Kzk7T1+qKh+4p
ry+kXhYsh+iu3+3e0Acr75At/UCV1inquHGGY/b+ztC4deQ8pK4U/MrRU/hgDKkusIKRvJM844/R
+dKQRgjRXQNvxUDq6MLz58PMPOag4UXGWfWCZ5Crw5mRriA59ffgF9wdP38mf4lx6jMI+asfSRyq
qhmZVaWJbPTkc/T3/WR+kbW4s2Uzs4wD279adamG9IIGFDQPs0c3LYF+5XIKILq4zsHA8w4ARq0S
8Y9RJk63BOhFGh+Zv1l8AEp1dmyY2zG2qxd/1iCFbAZ3ZJg8E2pJnUlNz6wqst/veElwBsl3z9wi
Jguto74eI2rJb6JaBS+4H1bsiC7E83zZkqgMWNey4NoukyqFI5XOZvEWSIN3GPvApzx3c+oArX3k
HXGx6D2ZGDiBQYgOBFW4LznYSGumzGYTKMz/aR2EwK1PdMcYcbIZ7q3g7MUDAODJ62PFn2slsAqz
PFgWoZ58j4YOWtCd/Z+HK4H6aOe7v50LmgazIn/4Rpql/fTY/EN+TKxHpWF9Y/fJXXDbUHRSdCZf
WSdH33zJPeeHSRDMtbffchVgnclsDIrt8qYhbFdW4N38YQqE71xYBrnQektsB6ibMcqXfJ+EJn4F
uaqnsWgBIpciI0O1bvsmDQ7lR0BnhKd+3HsxY7hWhatxuoCdYelXMAuNW0UXyqiJH9H/w8fd8o9P
TxABm9LIrHjueslET145eX1k8yNvIR4q4VW3fNh+7g11mny59tQajjq9CrY+fpewHT71bHONGTMT
GWkx+zjXQzMFwLU/ApyOz4vlrO0cuMLtDmoD7H/+HkN/EbxrhIhT3hArcZ3ypq4tNgoCg6rF7rdj
WAeC41Q4/LBsOicRibjmC1jcMGC2u5C4Il2KUqGMW9XWeXBnavl7mj8KQ9bYtUy0fv7Ym2nMgR3I
BjVE4kY2yOdMiXCVN4OiNkHLH7aG2cjoeVwrlckUicruxZ3Bn4S33CV31NKjHEhMW/yr7K751zoo
JjKWgKzCwNpn4fO//FtTrrg9xFNHigPHQUu4l9CwUJ+h5CH2A9SMayzneF1ogboKdPFuHUZUWDJn
yPqKb1TpwW+5w5FeT0aOyTIXQ2u8MO00TTbbAF9wnCUObaoXjEU1KCCqaUdeBAfFOqOsafF0Egei
JfvVCpq2W5BuN3JknrM9Y/M3q/tuBgdwVtruxF/39w88PPXFKS+LT1Yp0eEmHKeHXBcmNsOwy5Yq
NfGhF9UuU/1ChNAW+BsxsIavMpfm/vi2NudJC0lSx9Ts/811iz9Sj2ArPbYdYHBp55/Njj/upSfn
9UfoImrG2vQRucI6EDW5AFx0NU6egrZ3X/4g7lsmv5eFupwyeTdfrq//hwFjKD0cvjDXxvu5JAYR
SVkt/BEgBhxPjfVYclBC1Qh6VPysFvDjCnKq8uEQ9daVk0VKUO+yaSbwGplQhkfPupJ3lXrVG9iZ
gf2K5MYXVxGZgq84zOdUyEsEtmc1Ii/eH/WgbSMid3g25bKKHGihVAj+1ziXTSocVBje7XW1luEU
BvVmnOSlPygGWSPZ6ZYTbWTYQvoI4fkMUmCCBb0KTABYY6ZVQBw+asAm+DPj+fUV47tpiSYY4wGE
RippbDsoD/P8QRNVs3sWFrOHw/qgF/42BNGdTbjAi4zo1uweO/Wu+UvB6NvJvvZuJ5CcuSY3J2sp
9URUF1CLrRib5ijKx2Fe68eCUKcqTHwdkUY7zRt9zWWA949xx7dtMKRWJ49YOkA8Vs02IVSvdrS9
LmN9K+8UNwA+iYLfj1jOsRvtP7EiFs8VAwS2ekOGgIY3UXhtRjMq2Mjq8jtqUy72tgXTPNlSz4nm
X0TBTINTKA20I8mvDurjPdf4zTGlAi2VH3oiAlKwIWp1t8zkK22EasjUj4GU2nfdXEAdGt37H3E+
R9sYie7bitrZcWfIQVop85F2qIEy7PicSebVqOGScChvratYgTPNDgLKtdF3zCY4sUSv9hg2HXug
psnL8if9qQyXfGk9mnYvysNw5fTwcIqeGr1C/dNKIsyTlji9qguTTJAJZXUuAHgHzDn614vKV5pC
JZRzcTFEvI204StjpgwG1xk3g3XITh2gn1Avl4CyLTnaW+3gdjR01ZVhZjBwm8Dxn6mT+y20ANNO
0/8och8+0ltZTkMRKIWbIRzJPtVOG8DIPha6MAhIuhSu8RLK8X6e0VnkHbZvNIdy67IDFyQ5J7/k
5MqDaQU/mBSL3B8bgTWhrL00TtkMrBa6RkrSgEB+hXz4iUFRr9BM5a8QEsPIhUHdQB+GpyxDGKuT
7BROajf4tX39YajqYnznUq90frPysIKrWYag4QpmKWEeyMnSU/Rvo7GdXUzsoonzc/Dbbsv5FWmb
5Z7E+zURpX8Q8tzdedEcD+y5tPzWfFPec7lm8ZMhcrVTXZjx8oEKCsOF6K4j4SxUNPYjHS/l4lRK
2sz4UNSa6strK5dXQKxSCPgFBgpwOb9JSIvkXew8SWve+LtnqrNLMpDOM3RSn9HX7KefSY/fp0uh
cyplQvwGJb3m3dccmW2NJpJ0lX5gKPRR+RoimH5sPfds0Y3VHp/42q6hGhAlmvtmepGTGEBYMhPG
w4dr+nCL0DQEiD15qL0R5lWb+VVUHhIFAVSfexynaUWbVNbY8O7Wy6kGF4cpS6S21m1ppq0MBNHb
fNS/Wnt/NrAdFCAgMHPjxbyIgkxxf9xcGbs9mSvex1TV9qh1fCJa0FQBFTVXCO3ZjLiv7pj89+bh
ZRr5W097oO6r2Qt3FuVydtJ6z9FGgBF25FkMaHpSOnQK2ZdMP6uz16UDbjI4YAlzUiSxYKSfjQUg
7FYqTkc9rr7zjk5qiJBSeADRC4786XuBEjgNjZJa7NuaWScOpKbTpoAvrEyIuOXnS2fn97bjf6Gs
kZSm7ODaTsiWF/eht7kBipvbdQ3HsKjssVMUMTFWlqZteXdvaYZLUfgks2p0iBfOe8Xm6DI9lspF
nm98x6dLrx+9LN6wrIOS68omXww5NGFunNc+2kTSnvGrIsSD86SKip5rrjHpc1lhDjNnXBN/t7Uo
67Ecwc483nYyJxiFcREwUUYnWjcc2Roqq6iiW+Oxnk4IHqiaJeS4jyDBNGR5GNOKT6/DLALm3UXO
6j2Cvd+M/On/6J0Z5ltWEpUWP3AsCCad+VrpoATbSggKk4FGg5SqOCczWE4JD2UDIGw1VR58OTeg
P32ynRo+XKq3w2tNp0GkqRdn4Ozn4sdjr1YlgZ9v0ngFOYys7oyhTWzmThMWbdsdCU3sAZTZys8v
qEzBW5uMUCLg7JuSK6r1kmQHDpnUPkbyB/uq9DhbIiA6onaQgwiV/WYwdI+cj68cEZwdkpSFzo99
6jwOfNb4xOY6Dwf60/hJmqZ84ii2IOTmaCO/RlYQiFw3DA751gz6OkGbWL2rH2oMxBL/NqsqhFqD
++wyS70AQKWEnA5gBg1tvj8HFiUd2597lmRNoQEnkZdC7Q9SxVFg+guuneURTvWA4M36Typ8mbs2
8NxLA8wIEBb7xqM29i8zmMVbNp/HXw39R1bwTL8hf0XJkfnw8wQX+ItO2P2FESMEUjhgm9zxVw9i
yX1AA6eChxhmYqdh8J1KNqQN6GUsGef6W3faOI4f1mbBtx5cMUIAt6xKo/xyEXzcUSPQLkenfdfm
F0sXsiMH6FN7apeCWElzmcYJIzHlvKMXbpZ7VFku+kxglX1rjqSe4ILkTL+uWjkGSnlQDrWjSrNT
DDVlSKTdUVpMxVXyK/mcXM1EIhkX/GJed67ftgjzfhQbKvP2IWACb/YFFXjUsLcIRBsFo7Kwptv8
3e9q+38A3JV3pllGEfosXnZwjfzvkgzSiR8CcsCDLbMj3YgM5xOavtJqZs5CY9YPLQchrS51WVSC
QEr7grpFKaM1u0Gr9404AYGaiGjUS5APqMn/EInQu8yb6TZ2LKRu/rIF2NGRPY3MtSAsKKVz+jEw
w/83Qoa4XcfakhIYe92MeRiuXoXvLIyRGFCbhi672y7Z2HOJPv+K2a8gZPjiyhZt5MbDkaKEP+fT
r2lVJj9tzObQHoRM0xWYUC668Ak0ovOrnKAHD56IORHHFmTUuYEK3Jbd/yEgVIC7wAPQKPGrWXVo
9J168/ICSvrtk5wL5i3dqJlnR8eNSvPeaNtrCF3LjG9YAqwbrMIf1ayouXO6sAwggoIno0/v8b9m
0SrAGaz9BWAvPMfiFnZVyUxuTfjiIdMMlOOZzNB6x9nowPl2XyeJIh7/nt8GzlQ9sXpMie2Czh0d
hBzndChsOaFqZ+JBEFaHqvqx/Ay1BLosNKkNEz/r83ghYYoAO3CDXt6DVyIRtDOHIGspDOixRhMK
9bJEb+MZmfHFmDzOMKEgGNkOia8y7P4gHusg4OWnFEUkcdD/US5icHmjqPT5FzXyRb7sYaLp0RA3
4/Dh+39RaSTICm7IMWaYOimQfHnuCREVa8hy2LXBH7p1lapUejn6fpQyXHSpILmhO+1G9G9644T1
94Xu3v9QBNIOID/srWBzBwvaulYosO+R3pnmS3GCx+Uyw4Ir9/ZwfYxDlZs5VmvWYFyszmj/+MvY
kxZn+UeNfI8tV3VOkIwhjXcvjpD/J/BRe6999beZjnIiURjNctJB+C5Ks3NucodmXIhXxD5UL/LN
3j0SeGAs1i2YxVaRkQlxUZvgADrs6wuxw54Ti2Rfgt1oVkQm1RZ4uKt56BF0cQqZb7l7TYltaPNI
xzgVaLcM+Lj3FOg6S6j1PKld1CKkFazZ3BbB/gpsU4mns7N3LW24hdinZRzmnlpQ6sCp3SKHZX0L
b6iV4w96hzBlKBBf5DezRzxzMisuE7UQaU8bZANWYVjXZkYyiEcOAYbjbpB1jand+3g4yD44+CIE
OQ3hfQWIaad2QDcdL+rMo1GOatQnTXpvSO++sm4ctyDw//xbUDOXrgRwU6vEskKxVvXJ0kbMkhLX
89ZGenM5OkOMlS10slxV6LYweGfmFSeUQl05hbsWK2yvcX5fJJu/SKUWGgv3+6FYOFJwWbitFVf/
hIDCkMFRAmoQjb5x6q+LEd3v2uOxnIZTjRlBisSQSEq+VlytuDsenlK+p2A9P0WQEWRCtvtLZfit
HVxpj91YSXdnTQWYYtdNovbN0tfP1Mx43Bex4Yuehae+72+j+FXxSbeGLaHDjvRxTeejdq5xJU/I
BJpgCOpPUQdUjmX1hEj06QmGrPILNAHUsE/mmZxNVNPcwh32si44LH0125pGch3KzxeSncBr/3tO
gC65fsrxBv4ngxTSExozcR71cQmZqLteDPJXIUMpNRixIoVOK+TcOG021Hq013F2QZLJ3yJcK6aR
1DDf/5DTDUMLBPS76SSGlDrdRCFPnmULIli5EesUB0l3H5mXmbcTfqHXLOEkVSsm1b4WlFWMV7BD
gi0JiDUdWWXubObalnl82as+0TtTV/MaIOCoPw+NeT7a83S/s/Yru2yOaW7p0Zaozz25Lgucay8T
+MMAPk90dVEQvzE6yiBtltVUl1Xx/rcL2LWRFI2dmvHdS10e4YxfdeYymT6KWuPatuHv+F13+Ibw
0OQq0MSB54ezLm7LOOt+ozdK2vG/chDAWL8y1RO0mW7EZRdrOfGyi5+YySA0RfFSonqWomLNGBoI
RitNVHOYWNUTKrV/a0TA+a05zYursYLsjeUPeQPTAiPtU+iMf+OrP0gQqbqvaIL+uC1RDvS79hP0
t+7gmCz4r4YwyT0f/Fj4iBXYTLCQw0ab2VGkRZBPUGN1SVpw4cn50FVF1MSfJLyu+fOH2aYrpTfZ
QVbppNZqrksMeOlICogTnoZr4pbWiQMNyc9ERwJE0eu1qSncJYkv5KIfciJhJ5/TkB6RYVBegl1M
eRzeloPKKgJibHfW73ASDpDrGbHaq0kOZMYQ6HBU548aW+mMEZr5rEC4iehL8ypiDhNnRd9gk0rx
hPRJd0pxrN/32C7YPrt/iaz6d9bJnUBnse2FS7x5SttGJmTSdJfo0W+3NMIk8Dj8rNXESYicWIh8
g10Xk2+JdrlHaIGUdFwApzpnnYDhAFFKLDQd4L5P8V2qG5lj8pvo1/eQC7EonKZWasBTEs3FVbH5
y4j06QCLBQn884slIOylIDs5L0maxCF6m9cW8790//xW3YKx7VxpFdGfwuN/iE9OMWFvRLSCmSwp
pXNZ1TaJatJGhSZeqP7v5HJoWuqh0VbMqNYccyTfFFE88n3pLMTVtgVQyagnLGiHuEI9h5AVaPmT
K//efy1A1hUrNnZDGg1TC6me06nMl14e4+nsOmDdYLT1emnxycqH5jlMMxb3h+G7+b7+ktxGGxht
lFaKK5wYqRA1ueScEB0Fs5V6Oi0n1MqInfdgD6OnR0O7O/7KcETeb7+EBQETCraykHnsMSKr8GqP
emBI/MFkzV+RsyS0tLuQR0RJvWrMlNdjvgox64ahq0C2SKy/iOI58q+y0tuQ7tzTDDGG+YWEdxQK
Or9YDyQ/CiUgLeTyJuYX571xYL/8VXlf1LTF8rm9c1iBrqokUw9O0gv0tiBqf5AdMYXfa14raEJK
2rFkTCq6ZoXUxf7wVmrhy9+aTbqjhxdVdDV19IfDqgCBhdp88UQLLgcueArRNpDUhF8vkCinwUO7
HO+XCSH+akV66OZ5/zum0wBhqq7qYcgneRp6vbXSziepGUurjs4PJsOSbc+QxDOMVctisvFho1j6
N1pG6yuyelXntYuESp9ADll9/fVGt3RYNN921mcZYCuMr7MC/JyGy9OTNuUa704+GsLSkRhnSHno
7PwdCLLBkmDHGcjqb/eNvRytcBXsYJ1giwGd+xF468Z/xPCdBL2WK9cDZCcASwvP5zc+YBa1FQRe
Dsrb7UpLaag3EAXmTqxLd1/KBbTX1TQGq+7xB59EqmpkkCfGdkAtvH0xZ5fd6VBMQ0uSrNOUvW13
zQqAQLYGctRhg8oDqRoQIM8woCEIrZhj8cq9hzncoiQyJJQkpEtfYbmB23ktcn+pB8US1CN9M/c9
PVph0Izo7Oicrl98dO55ZEXgFjz3uAXMtQA5bZmmdlIXmpujbyZ6D3TDDq+Kw6FKan/E1HNRHskI
w7UbtuMx4NanspI21UWlsDZ9m6rEl21qWsAW34K1F5xvtGVgid9lDtA8+fk+yS8XhbD6PtmB0nNc
ry/ZLBWXBDL7M3rn6rEv4DJk6gkk3MrtcHZ1B2cGxr+plQ+Q/8ZfsVexG/lK5xnY+SHGnD11BUeu
/XAuv21REnfOWj2mCX1WvQUYKYq51D0S5ESH9VH6j3OPlKjJuMAKznOv5y5mlYID0oU8+boMH8nP
aKoFaGjk++NlolvRibfOT9Kms2x2dSmE9jCW8A5pVS5KuF9F6wSDLstZw43bBKtR1Q/IC51ujfMM
DYHUijjxFAxGctreHl4EXlmgMag3jtPih95rycyQBnpQhbUZI/veCctX7/n2foyhQASPE0gbQQ0I
tlhT9dkhKeJmR7xYDmDgZ7sQHiaQyenFieFmYgaZXOcI4J7HSFOGOtDLtqChxtFv0QcIv/fSSXeR
FMMGLBGnPYkhS9AqsjSVn4+9w4DwKlE5maG0OTcOyOnB9TGvHJjUJkar79e0dg87MXAWbxkf+Cmf
h/qlFrvektfbC8RsRyujDYQfnC12j64znaEXLFqLIlpTkkcM9d0Ug7zdqMi2SrCrI3GY/CvCRnPc
kSB+SOg+UW7FnOSBdR69JoQOLr9323QwJynhM7HqWIIACXw+MFjYsYGw+qV2Nm7VzKRkYp4+wGNl
Z1Jq/vapCrzTmraaZfu8qRpPpcc4mM0ZT2QZs13MjW5rs/T4c6RDzhiIpYXhx/xFKHPL3g+Z0yo4
a3IVrEUQWd5xOzv9rqowjWILNhtPtZ8u2s6tN6I4hO4uExqD6bFISFgky5L0FgvlHlyG1vX9jaCv
zjnIkL5KhgRPAoaTtzE9a/HJv/vCrqW6LuHpJZ7xQNw65ZbYmAy2BER6PbQlijs2izU+Veozb2oN
MzG5tTfxBAYBNSQfWV5jnnii8CiNatWENCLtK1tY9AUBjC8PjFZLSZ1AUtjtibA28nv1refXsyFH
1nbuuHFnQkoKUPCKUj5nYjIzmMjbiF6paWUWUw25WcacvZbUc+N9y4OKuqgVRCZOE8icQ5T5ipeV
X99xN6VpYbW9EKefLeB0UQC37Tf3YNY/Gn0Caq0dIAYxx4mXdtf0MNvIQAnjU0NO/m+Tr+z+GxNT
tdcWdXtjR5Rvi5w4qUzo2YuRlST1dsOYvwhp9YrxdkEjE4EjGtRO+1OUa8A9E6q46+mEfXUmJSqK
kh4z8MfuTHhIYBDSEPZYblHrSi8MYWGRh8xtDhYWDjOgR2nqiF0Hn6/cVN0yiW6tfgA9mtAWH6cD
lcvDbxOkAvJ8YdWDfC6tP0vrIvE0l5k+q7+9rNaPjo4YKzmBoisa7lzUQVgBUoMpTv6ba6CishKi
V8Z7y4RYqxUdsxKqEj6uHb2ub8ssUEO1IqHqCW/aJt8vM3GyX40HTaZL3Vzs6rNbO9aCbMJZe/2C
KwAW32QvP1gWWWIq8WiVEBFpONxHvhkbRBsy2oQDEVAO/6yuyShOu965vVO1Zx+gIJ9XB+P++8ps
8R1hDuDmPWXxp6w/XaURThMn2fDOZR2nBw/x0SeampIukqJZcszqrptTYy5+3NoTEKjcL2A2N3Yx
hyi5IeSQfR3PvVmKExROQZo9uX+096BxxgKRhLDGxF2qXsIAR+h7s2R3Gux3RqQQEWWG9hBNYPyO
nv/EHAuhUBg2gwydbIZE/zRSW/Ct2eNvFay4GeGsRlKMlGb+nW7o/kJgGRu8W2W7m7fM5W5usNf9
sFg/M6xL9QPVjFD485wkRrbx+5kcepjVsGYLdujxZThg8rb1A4yb0qhrBvBBVQpEewwIRUB73FkL
Xx8Tl2lvcQTx5AVCdmf88aboni0zPdkHtWZQa30ERbEq6C8f1D313f3mpfqAs7zwGkWNl6QZ8Peh
oyYwHyqHeZs+3vALUcfr/CHmjOhI7UQNxOXZAUUHllRT9zf21x6kKJiM5VgPlhShihycAePgkF+T
+z+HuR70KBHdysa4+h0iR7KUqAAw9bQ8+FemKLlyN5zgjWH+XgcG06cif2UcklSZz2zPPGvUYrDC
3lQvkql3pYKhOJN6/eApRJbIZ8Pq6LV654itu1lcQj5Q+97oQWnKMj/etj+e7VuunVXdUsgFFc5w
lJfh42ekwSrrn4x/9/34p/A/jypurWz8BmsIIHf4zRboDCgdACxWdP+4YxRLAPPGPtdPbebwRgGX
1GFqVLAM47WShfAcCM710NV7a1d5ONCkhfHDXxZacDqBLgGxLqRFRmK7Ge2ZHdysCUdpIex2OGrP
O9uWpFbT/dDHGTnyV5sKPiqUe26qI2uVv79rWVBGursMHyfnBSOz2SIBXIIf7doizagsZAuPjs+8
tD2GUmEQiIWGkqCTt74gH+P/q/kHFf0M4D56n3/vfFckcC5f2OAFDQ7zk6U5xzE6DRBK/ZXUWcQG
Nn5bo74DSUvA9WAig4u48cp15/s80qENWYM9ljgDGXECVeAH11dpaPhwJZYdkdCO3iIhb+Tw4hmA
KzWlP9iV4mfprXDJ3Q6P6moGgAVLB68CEDzR3s5q5fwGIat55K1xdDVHkvjEBjZbbt8FQVMjFqNB
Fn19LWMAxuZfHByyxrBQSx+WaqV6oknCNBTEKWYXGeXUuad/8gTgoQ2aRJP/I3SdzQuHV0Uc6RK3
DDo97Tgou4F2enbrQ19PSqIQL4rUBH4xodDW9GueUdg0E4jjlgKW1FxF/jsU29iAyZ/qy0S2t2WK
YdrEOQuDzbEKBZttBAIzEBeMpK1MRYwNeC8NtBswUUGknc0OyHfJ2X75ZlLDdhYGqLWoiq6w8FXF
EiQsKt269Tha6QD3DDrbZfiRsoab1EeRScZ5XCQ8iche7JhdrijVyXBXh69newUQmsWWg6j5qJxO
btCIw2b2+nfqE0kM3lj2C99tpsskZNuuAJqwKtB1pNZePItFCZGZJTstcYoF1tqe6/nTbKw4GhgJ
gIx5a2x7PGaYYeiYud2Rc/1Kz2iPcBZULAySCVPI8v/TQ31mOENbbibV45+D310WqvXFf0ecwZnu
RrVHfPU9HXxRwCdqOhFxCgXjIClJ9T+/cMrg5jJmOz/a5nmHJcMLlhFcVXcr23qA21zIhlLU1N2s
IFTZ5EqH1OFvNeeAmBj0OLYhBryy0jg1NTYGHX3tqmqFbaAXC6oXvxqyxjetYzt5BXB6JZLJfARl
wFNTX5P6ynLMovQYE6GHq7XaY5NCOVsN594ziFldUk2dC+x+9DTcPC0PUJAxkIKM0uIie//pgMlv
+iJrId/ML7HGoJziF+PNypNDMvxKjek+EJJiAJ4Mdt5pTFfB00K+GvofoJ120n/BBUvB1z/QUg7z
LJxvLEg09zidoDWzVRclForHN+xchb9OMRkuD4HDj7/AN2FCxZ4+OpGIQCxXpEybZ+wgaqwp2k+b
9xEDURFJPYcBV/a+P+ibXt2NBmfVB48WK2MPeF9HyqJxY1KsZmXov5uYLAGqyehaAilJ17/YrzS7
gnHf023F9Vxuk1zan+roEWce0ZnzJyCQuXU61HaQ2q3IN99M/Qpn5Oa/AuTpMOnAamPB9NtxgHlj
keDcBwwqUk7tCjBUYbQ5IPwvjPVucYzE8xAvioQp2G5+67AHnRLJj1m3y+L6QmTt+QBxVOUDtLzp
TNdxRQyvayStx5gs3Agb24ZNjsq/E7rOXM1A3ucNZgjdhWTmHYvOswwNgH3mDe5A22g/UjgSTKey
Gykk9KOH+T5FV/5I/x4pL3gB+SX5rK0iwZu82ZMDAsQ6rb5PtQjzqscZFUBOHCG/q3nT1n8gilID
gSwwqvlLoyNP4b602/wESSjiQooQp5mbzyQM5f1e8yXeGJqpK54l36ETHAhXQ6+dF0yR4FVR6Qgg
s3n6MFtDqnQ0wOZ7jHty9si64LScpi8JbpUg/ZSk0YfTfvSxfyOV4raMMznBSK/dxjNglPsWL/OF
+Wz9zIIptwIk/Qhy2f9oA+3SQPiccpkWcRc7W/b/71vsH27IGXOnBSkjeZLyrZjqM5gm3uF28jY+
ye8bgM6ipDQJqrd0iNVfV+AYJ0jHFK2Oke1DEyxRBl69m8B2jB55cbWOVhYQl4AFfXs8UIpZe0wA
Gp0MqlpzTbSymiwv+KxNFmzOPdTxbXHNw/kPgJi4wkKL4/iuePn4dlPG805xE94m0hXUZAlntA77
LrpfLeYYzACNeqo57MoWEv3sCSC0pI4HTkAPOy9VD0B+jDNeD8WlC9kD8XUUSrj0Uxwc5VWJuekC
oGEhZKmuZ7xJPXKGCtxngjJ7udvLiRjz3K2jLCaOrWhazkhPxZddVieRTuksGNPWm5cFbqnlZePQ
MZEkObTQHWwURSDz0+azd7asUbVDjSk53e+X6VbY2wQ5ZyHywR6Pel66vZeauNVJq4XswgSrQxHD
dNEbkUFnE+xO/9qkNWdtEPTCNOKEigNcLulxYjwZkBbkIJJIjDujImf0I0hGwg0C0/ijwetyAE/e
JOyW0OOFCauK6DLGfuGKMo7rU7AuaIRFNTTGLkcIT1I5YgNJzHDjjBFlt/psv3WVJGIMG26yCvGe
GCY9nU0RsXS+QIisoonFy6UkQkaZNAEpeQ0q2E6efSvPdh++cAIhHbpRwIdZTdBHiIC6Cm6EXgVE
XSyduG2Uaj0MlnEIP58QCwLE45X8ovBnS6z4Qs6AKTNbp8kKzE9MbIUJllixcMml7gjYRcCLn2r2
XDAFUtARoaxBVQHDMZ1hHN4CH3At6qGbpr0+gZZmgKsGGDJLJ6VT6YOaEXHel96IHPXJ+CCsv+Jm
rk8PDTWu0mef98oZxe5k1sJimkZ9dSF892rgnLe7350Mq3O6fXQKyhTQcpLt4iu0ZRPzC75bqzG5
bju6r/7ohxCTxxk7JRlfiKreGOxpNf0Diqp/jhUKoo3XuPNwjB0oh9D6vGmwo1AwI7R5VTtkIQ1b
2co0CW4GTa0w0ZeMZ9QIxFtBpQs36ewwfrGtghMeRTlJ6ZAtYWtGkS0RgjcLSVNkqHC+0Cwjs3Ao
UGMVLyXMdokfp+HRCTpn4I0qH+Vs867uK/7NW6Lyq95CpQb4cu3Yhwh5nlnNVDwguFrEWwJane2x
rNlAVDYv9YM9EOLqMQSzn500LqHX0jUpY5W6KzPe6wA1Kq1SslxfYohhonSedviYXtdV/GaEc6xT
eLTdESRyI8yxJiXtJWEtkE1FchMknOrzlGXSFEtIVufooxdhOfJQ2tZ+t0csj0/XPSj7/P1Unm0i
UoBdLIpeINGaq/WMri4RzNV2/y8QDVKJlE50HZ1OpHmnXyzUxL5olSTZTGG408foH43LytjLMlt4
n9UJDSI0sVNP1dvud8rkwKBCxtCxDLFV8afcWI1TuNgavtIF5JdJYuQjIGTsO6M2jF78spi/21lZ
P8DGxwaIIn754lrKGSLwu5cB/G1rGDL1pAsQvyNKJa/LB8h/QPhby0ENJPRsfBAtGCBiZ2Ti9B1n
QMEA3MDErjhQuuuF/m1D8fuNJ2Sh2LCd3Vopiw6MEc0vTrfqbJMMEwQiUIxmuyEqQIcsqnX/IDG+
XfVPontiEfLOVxr6GMgOvOF8CFWOpto0mCzxx1RD36ESHPKEwS/mG+HLceJFXStnS4lEWQK+GSmf
uDTj0Q6tO8Oq4VPk6zNQq7c/OctBMf3vaep1YF6yBGYr1KqUUs7XyvGJhuWnWs+WOR7kNeKDPpAO
yZKJNxfRZvc2pTdqWvMoeDgCAw7tfLC5wHufZXX66kDL8uIcydYBGNQUk3vbZTlSyytc+0Lld+uQ
+2QRD60M3npdvmfKfAvFbe8sdXdL2AyAejOxjEBzbkxp9qnvQSCDVIZMLOBc8dlMWOabE29XbNQT
PbxUBV2TUFvfVkmtUA2BAnZpYsd7ftDZgLCgUMMw+zkyrCD5FjU3Z10SSRJO5hKSr+ygdHkmHuMF
J+Hzbf/SOXm5QQWlYWgkxMeGGbGKXIi54eGNGAYWQFombwXcZzx/PKfmx4ftw51XdHo/WnUMlEly
gG4UOiztRNd4SDS+wfQ/RiLLHKXfEkL0/QQmYL0GcA7zNG8IxymJ5fUCnOpHqSYtsLqilrsf8OKS
1IYIZV8cj0aABOaj/1Y3BQOZSNOjQsbdy6ukIBRjhnMaNp6kQUQi+L/Vg5cCyG5+GohIdPkGC/fi
bE7X23uN5RRyl0yoXoVgNjQ5nARlHqmXlLwPO29xUVXB3/zG0XVbVuwqOb2S0qYpJm2GfWp//Ia7
69PtOwmksvimCajrvegmXn677g3Ls+iWog+Ze/ynMn+Ly6qIBGwIWi5zpgvYaekF+cH6oVPEWG7B
gJKH4htAuzxflG8ipSZXor2v0jKiQoOvpvC3zwv0T4z66XSb3A+voghfDTsp1eogFgTaZdbiDuB2
bEJyFpw/4UpQ9ob8/uEJ0jQZv0CQ2HNWuwQp4RRnssMm4IWoEmfEfUXkQUBUquVkMUXrSxt8VyX9
wYRNv+Uk5IZQm2fsvzT65VKKovfmNlEvnFNGaJX1KFL7ZdHIVxaarbZA/0UGtjoLh0EpUhyQOS7V
Sk2gKN9S5h8DU67E+/syqlWjw2jhCi4lTBKDMWfHgwfTj/wep0c+VFDcjyWH2Tu1egPQyqZhWEQE
yH/oU86aPLMw3F6+935MvP6vpEkn2CG5BYpy0i1RoZXviUaGYMdgb7OYLMUzP7Fi58mf7pWhi42w
XP7pasOtIcOEbw24exPEvmodSi+SZLBJqJ1yblZqGstt27+Uq950KdXJoeLPOtVS1rrDfVnBQnCy
NxW6As0ist360OhoJSQTS3MJGQyrJBGkNqjCZIwFpdDog6TqY2Ep9p9V218mcM4ngQeiscNKHhol
VmtNbYHpFB5ZwtbRgv4rYgF4zpgYtuPx/WMyN1ZqB9sNSt1un5PEt8m0Kr3gWMjrNzQm6QqJSqZK
35fIMTALr12/DeC+WcRbav9FEcz8zRRsf2O1bN1C/XBDRqxg8wypakT405+Ll8W+2/4K/FODPrxv
ZitlREoTvBmLG0RGdzTBtKetybUTshEvh3tfdJ7l0cTptBZjlVY/UtOuZp1S6fqWW2rjausIZ3dW
CVnpJWIg04Dr5MoLLeGzjINjbI1FCwtIegkTlwJit6jHuvckbbML34mLa2Fo44ybp58/rSJzutQk
rQkUaHdHjyzUUOObbYoFEBdYBeZ8aMHZ6qR+JIbHqS+OqiAuJUHtlA1K7GurF+FnJD6YVIj2NbgF
55mBLF3y4Ijx8J9TtNDwFUMv8foJUDNndYjB0FUoS6ecnKLxk6U+42f+xCd1n0jVxUDsbiBSF+1R
mLbQ4PwjUYCE5TkTbJnr1Hkjp3k0LYD+ltTfgovZwh36FwFvRLuifCh6w2OxUGaEbtufLchl9IZi
r/qwix5wW4ti/ImTI7rkf5jZD9Ut4fqijLir/IZjtCwrKHDxhs6ByT3PYUrsHdSdcY/VZboxOjw2
3qdAB9bcOtMHFfLIrlBd3PBLVALwjN7lYl6ITYulMyWmgRFJUJmTZPHTWJzecRPUdM3ZYFuMOWEW
t5/aVVYaiHKFoHKD5aaxMvSFAo720Tj+S64jqYlIsiEE3Hk1I1MjDTze0K5LOkXaXITj6US+ZafD
aoEyZi2uTS1BwVoHfWKg+5toEpfeaU94aAXbMsr70ghI3DOPSIiBJoqScVTFV0wM+u6XGSaQ0nBF
VXdueHIy5yaUYjK8wi+CpOdbkn+o25psFxhFjwEghh0NZa4ZlTgxM8TG4lt/UCxFxYbjMVO6dPFk
HS3tRISlvPTY1G0EJMTLlwVzazZEznRT7xOEKfQr8v4gOq8Wm9DQsmtzh8ttUZS1oriAFmCkYktx
AJE5y+ZvE1D9rv2h2qMRrQuKnNqE7jgJCnh/XDI95MssIFaMjkdO+SM+eKebB+cDCtVMxQPTKkSW
CFkl3aXQtrGRy5MsIY40korD2jlP2IXn9AP3v4hiJvThdDIXAKdFqWKVGhkG7dP95Yt5pglRCZV1
1Wonz/fFR0Z+m00f67kCmnunjOyefUAHCKpRYdPmiIN/XicHFuRTX/mtC7BJx41ll7zGSMKDSqox
48cluDQXQO3gYGPH6bWyqOqR9PSAWndNoIaEEAZiNHtYjLCroyzAwCsoZQQ7wYr+7hyf4IwgmP91
e+TjD0a9uyCBMqtPzhG5mzVbqc+iVHeob93dniZ79WZdVcNQOqFt3OQPWZSCbqPZe609ImL7oV92
JMxoM/wx4RTUJqYz72dhmDFqzRpRi7hxLs34v0MtXjsKME5QS97E354F4qRl+1gJ5qFvYkR3ZxqA
hiXIxldJadkpX3MV4/c0+Qr8SiP3+lrO5YmMsMjanvKk0/ySmgD68qHzd1ngYXAcjXBQspkBEf8N
QXB0vWRdUCkGDBu9oVCTapTMIgCRadmGpKcLssxlCLXcFFlrueA1TD6fYv4KfWGexflfpFVOIBQw
LfyzsevGZTLd7r3vkzfCtGfiS8dxv34tWvqhCSERQ4kRAaf+iGeqHeD9xnu5jRfXh37GA1FQ3sxs
txkMK+xZOEqm0Yh/oait8geBNC8tZfm3iUC6PJOWI+1JZ0GNyodA6uc/0UybPSRj6DHYvbzHDxkD
yQYlHQJC1a/bLyz5wYFv5DXVZvZ3tLRwKGrpt6eaeG+rClWJY+NJ2saKwmRBsDooxXLpIvstRwgc
kM/ip2HDKoWQn0PYH8QskZ2XKT07wqhk55FNH5eGYD+tVn0Tgnj+71+o6geC8YPWpSA3B5LPA5WT
WIbMbzuOtOQtygryq3gDNVsJGMAKHrXjvlNWr3t0QhZbqJ8kLVFKVVn9jfy0is+BSuhbbdYjfiik
qHMq1Tn3BOlGaewk2o9x8T9ugHkU1iQTBsAC4Rm6iaiOqu7ms7oGfBEspTK7Tj85lA/WGpyme5fT
EIpsBCmhQ+0GGMLbzrVkMaRN2/1AMW9CXTY3o4toAZZg7IS02r94uJjATQhQSG3gi+UjIvOQslcP
QH4s5N1FDX+N64KD11Mhh/12sn8XGLejOBs5t56aljG4qLLTNqCcPJwhOEup2myRIiXfRMnNVrp6
+cBqmjnURZmrCxCHBUC0QMBmBTF+jD87WMwP89QkWH8CoDgMgidus/Cf8jh+sc8HfyjbDXAnEJbA
ieze8YrUvpl64UAjfk6ymuC/m7/DTHEWJBoW4ZdePvk0LmuGtt2/Myw83UQGtooNjAPSd9jv8zoV
/v7fad8OIG9cNimLNKikGcsEz1FkbfOe4FPTUbpCaSheBNR4m/ldk0TxA6pRNoJ3drco72JUlYlL
9xKoEYJazTepTDBckQcoF9gXjhIQZaGqlhwaCOIDyFB2fFTUdcBN1vqvQuvzxlOMKLfBvgKK45YK
wHRBJposSONOlqgdjR/12UW9Hce4SsW3EC0Ngc4bebzQ5pE/w/WP+8EvKj7q4BFw1p9oojHAtcU8
LGvq84Y1rXnIhxn2gfoQpl/e5TQsY4S+xVj4E3HnR0/lwHGvhx/Tdyj76RvrQ2xIzi50d/AZSc28
Uf0eKJFslKt3rnt0oQ6H2UGlFtWr2+0FsurvGtVEqkqbPx4xw+nlnZs8vncuyxrz/uYprx0aOg4S
isBBAubejsmc2PjiWhLBNETffAVUxmlzgwJlcJl6S0TmXlnF6CxhdZcvBQA9hLXIT8/zBUPVFOTk
oRSONJGC0O28oF/2kUc2WDGVmF9D6XmuJh5sV7wUOmOCCfJMHX/UjfGjDfDudV2zdcccRmb5z0TP
ToiMs+lNr99cDBnLCVqQpkQMgOKGYPit9SRcuqPyUAoVe95cYpXMEx0+N29vzMOqN/CeoFAhhIsu
PJboCawzzIrl6Y2UVUEVPCDRdGxvLpzM7C2hWwKnDU9Zi5Qjo2U5KQho4IEt4sb3Q6YUV723bHn5
jHnhGNiYSb3IBlvAA4PSO9PgjiHRiCv79KLJuBhnXlQsGeV2vaLiQBrZ9trVHPrUq84OTYGbenGy
zMQ7mrIIlJqLIbium2Vyqo/MdMSAZdBuLGkOHnfgqFFwEJyCV3G04yFaJpEnORysCX9moTIEP5zZ
MREKfgPdtT9WLmW/jb36DmgipLniog5x0qQkxyRbnualf01qJ73hfwweubV3V4MoMX1YahRtWbJ0
I3zsW/ob4bCaMS5ByC52TRYGXgqkl9kwtVkXh3DoE/4Fmks/IhdQ/3SP5BJlLTHUjzzwzrpgPtNz
id5fwEtQ5bmJfCW+ner1cPg4y/O0ro4VuM447vFj37d/CGJzxW2SLOo2uT2SElcvwKocGQiY9cpF
hriahVRj7ULjORjUyQVvP2QgKeVl6w2kDffOHnYnSHL7dm0jL/Y7uYKIJ+71tnUYQjV4htYZHHNU
VrTkgcS4ObJpC3rRYDc5IseuHibkebWSSQmmChBc+fXFCOZD5rGS6MG6Ikq1WyU69jiCXEglE3Cm
YO/tGYQPOe78owery1M6NKPavPc75DIpnt9BirPq5Ms1QO1ipMEkSfiUUPXw8mjiTJ60m6BPbXBv
96Iwo7Fv9xCktxClfQfG7gMVfpXvTsONdh+FgRrhbO84VeT6vHjfexM62tgTWJrvTX41/9sSi5b7
V0Dz2CaPWI3UcFc2bp51LspCwyZGH/kmCHN3wAwp2vZPMWjcntJGoDi1BVTy1TJBuzJ00Sjb7/3z
FqM8oSrsGecHpmhN/IAY8gGEF7t/z/mQ/9jJW3sedgDSkVEkGnBAFjGK3jFbMA+7/3WgKdmgz43l
YK+27rlHEW8onwXt8kDlhtc8UNdFPz4COrAG2QOrsu3P281+ec77HvdBRQOqGd792cBHOtPvA8Tq
WXpdvG6xl5GQKjXZ24uCnDPHvWo3jYri4JOTRNsfJ/bHjd5oIEi3xBsrpItNuviRi3Anly4lh64r
UipHBuzqutIq/ZZ5Chp5GYm8B/jCIJ02tF3l9f6sr+Fft+mkHazUooN5bkiBSY5KonFElUY4kl04
m+xmZWf/AMnQAnhnVx66F7MsC+D2R49FZelzC0HHNBUxrPMHM3fjQGVXjRbvC4efiaL9xOMpWtQX
u3zlaXpS8TuNMyTsCoi0KAPo4OuG+ygc+G6E97R9typLpRqk72cqWYaZ9pHUkLKbpK1JS7WgOhue
Xs+gRQme40J7Ur+nOAsoXuoDjVrew1Hv/t7X4UFIFKYkB7B2EiNGeXnixPwLmJe/bfP4WbGD1Mqd
a9l0qSiJslCdk9Sf6V0JA+rqTM18nfE07+dkPw1qUQBr3qqG2y8srEFIca0lVGsT24nKltHJicii
ACVzHfxR1/v+FrWAyjolhtHutJdqa7ob/CUXLDEa/WhmCHFRkgeBDkmBpQkx0aq9vLmFtlzIuCAf
dURFZ04YIWYbcElFrMF0WWKqG5Atv8gT++STP8219L9GIcWaM8gbBTJizezlZ121p7G9qdTKjS0V
x9roqgHgzgA7I2E9kox1RnWICOX5hnqgBi3tHteTBU00MUbazdOAx5KZFDQ1/HsSbGmhN0KSlDTC
bnXcRPzjBJa0BwRPVzo/29/k4FO2B1DuCv2MIRUH9WtuJNkbBJEKcguhkM0wq3WgOOlMN91YU/MO
Imp4S4NJ8ihxEAvb4OUArBOmS0IRXlccHHrro0cUONRkMAVVpO0sgL09sdZSsGHBDdqz8FkCBZgq
sf07JnbSGWOdhDZxEEq8cCSdmpmFtZ2YAVumG/Mys/JvkuznEXUVCYg0iS7NS4O73D4hRtun4Fjr
olr2tgPqZ+FmK8TGHBlWMfIN/omHPzCgilkzHlJcgZDgy8clwFjItTSqWvRF5JOUZ9T7S7xd8G4E
6v/oEgK1Fc8hqTlbIWwyY3/usa9H8QaJUAYQlYZEchYJGUOxk/XLsaoQrLhfy0nDzsGvasvyQLxR
0noRxrOfjsltmPATrVqQMPN7JhEVcEU695E13407Z83zgU3ZM7C07FomBMuR1MjceioQok8Sl6+P
9VwaKsIyypuZUCRZ+Mte0yKkrC0osyQl1WKS2xW2b8OLm2O3fW1Sx0+JKMIxHvECgHsJX72aTwv7
zLB5wBbxudJAFge7BTWWDtUuR4H3LwN7rsL13LpZXpKx2pgDb1uRc8h6dcC8aVcTYaQ0XRLhmhZJ
kEP3jxUqtWF9L6j3UI7xcf8Dh9dYQOjzxIBoIT811dfGvSO+onHHF1o0keO2P5+anqhRpu4M8/BP
3aoOqiMc/oSDlUk7Gpe29MBROU6m5AfaNPCYOC4MXJ/OLhElCxFKEDtuCtMZdAFU4m10SX+mLE/g
xcjdqGkj04tXCSFvUKCuKHlnktx+v/JzIBnvZKnW4Nw2x5Uv2v5WPl3Pk3RWHSdC2jBCK7Id2eMQ
RbdABms4a4CRT0f5BqXd5s97mp60li1X3f6r0y6KgyZM2Em5J9zCFbgX6zcSDD84JFZ4EJSW0rq2
yEh9kRmNR6QOlxO+2I3zoNv274hOCJHN0Uyaarz2irdQdxs8OOjADcIgGv27iDr1ZJaA6NSyUvoR
1tP0lJ5z9Od+Wm5CHwHWyUy6xo9qZbIyG72UTYxkCoDgRscSL7TGNss5LtfRopeMmFm7CDRP0GxG
DTSrfXfXlNUU+l/FymU0E2f0e28jaMOdwnZeG/peiRlSze9YtSgo/c2qAbTp6z3aqpW2OdYVVzEZ
5angZjwtJ1xCjEZcxFXlV/tetTHluGJvzYDjXuuYkjc3PIZKpIx7h8BBGfTl6blG4TAInMb5/i49
otyfXcq2kqSy203GHHqfsfVcyNfta+1NFRmS253FTANpsnduF2n6/ry4AAVX+jEEhtjHHyeVcz2p
PvnTodgLySH3EWPjXM4/D5NBdU23E5WClqrLdvudNeo0LotlCSnrFJo4tGQQ9beC5tIAGdcKt30D
lSOBZYAG9oXqhur/lMl1+v/YvH9DQ1QAOG8eBtCm0ZoJYIQ+SHOhIEgJxYwmjPdZtF7rgSNU6rVL
18QbAlfGSFna0fOLnwnSSWYgZxcPeQY/JnJyOrUiIj0LoMFY00zC0bSKN+V534jDC33LnNhizuls
NwqyRkUVSwhNBR//MDREKADjiBaFNRgyIrT5ZLTacqNRQue50lebGPSpPepiP5x+ac1tFEBCWgh9
2sc2CWe2Q+9rqMaP7kVZ4APwk4yirJay8McMjlz1ldqc6IxykquDvTWp1wdLl4p9JsYRbOLoi3+m
KwBV1DJpwfy56SoiR5bJIgF/uSGRCqc+NH/zA6mAlc7OOo3SoeNZ3PLKBBaSxppKCQtrtXxU/fTR
8d2zXopDpJY6u/ZlYtcWvEst83LRwLlifgjJC0Ika5pfTEBTg57LU7krMdlvNTdZPqUd7ebt3Bc7
m6PzmpPe/aksaEvhbgDaty9OQsRqTWvpCzSk0g6fC0hyNv2zv93+H4xUTLdK3mYhtzEUfTvHUVKl
iY3OMfPvgRvWJR7dtUsphdXXdZKy84Ay5Ajz7D6wCOxaIDOYGTZ6ovd2zR0L+nzYNmHFn9f7z4Vw
o3nBBYxS1XFIRg3Gdt+VRdSY5vVlMMX/78hJosgziQni0dVJRdPYnpm6/KFLExZSrXl7C5GRl9Wn
pwODOq3kID9RzznBvLww59Up2ranYUa6GuaVqmOSgUNIQk4nAt+YW+6Mb8KCL8DqjUT78KbiaQWa
MKKnZnacoZvwOaU3C2vOHww9hv9datry6KAgEYQiEEN7sj/MdDshBP/J/5/LfIn2TRts9VRQ+603
PoWfQACxqHDjMxTOhw5MINMoKyuz9V/zP39Hbnaa+PBgJKazeQVC4Ndh3TeENr5ww6SN9/vggY8k
fITeNzvSj8xF/UZxj4/iMyoEq6uLqZwDbvdRtUt5qW8mbQFGjoGG7k6ncjIortd3rLALAHvn6WsQ
pLcQl2IU/J1dOPwwatsJm1eMODhieTTsqcyXISnj5rLTDFFPGM24xu669TKYnv9jJpU30MNvpEvd
BO3JUiIujjl+mZ8ArbUiVzR5xZtRaV+G1pYudABJ/P7L+vCOuupIwYpa1nBfZ7WSXqEzv3L//wgj
aEO0cCKi9HnfgOoeMLvTFrjGU2oyGg/jJ+pCnV2XVxhxEHy+FAAxL5SoZ4Kb3AJvLzOL57zd4afa
69bWvYooFZK4TMYl7TaO0zwBaDzIHVGlyBStPH0AsVr4hT1J0kBPxymqqoUUSLzEasS1syOC5tI3
a58jzaQAtZUabElg2m8dQZPVV3wretrdVvVG4ueU/iSuWfIgbhF0jH2PS3ilwtFGfprDz1agcbRx
rlJfsEy4IMaQeKd7RbtaqK7ldnK96Z81JAknbvyW5TUdrtc3anfRSt+bA2AdXW6xh6nHAiOkVQ+6
l/TZil4HvioGGJyalHekb7rlL4CplqFD6smgjPfieuXsGXdv5j/P4jmog1srBi0tC2OgqNcGgQMQ
FHIL2eMeZWd0pHLV+D1Xh4PC8CwR4MxWMqJ015pyNzqq327IdUOIPDojD9/6FFy/Ivo4kpf2bYsR
CcH508KGWvWf1/mU3XMhbzTNuuEBq9pGhpdoTJFRRHBYnO2laOCs9H23BJ1hGwb2QFrrggiDfBj6
xMmALque1fu4GabeTsQwnd55Pl6W9ndXN6iZ+ti8eQCSCtBCFAGCYlgXD1b1IkvaPYZCPDYvGmcA
09k6iAEdU+ztcDiyeqtJmAeQjc8HoOT5SLbbsJubzzLfcJZpwJsTUl7MYjha8Chnl9gWZtUOSUuL
dKa/JlWz5m5EBvYZlezUnVG/ED9UcGR67H7lmGhrAM5NOypEEV4Zt6H9ObTEUIIf6glvQ4wEnXcE
ZhCiH0ijiPqhWQg7DgROjCfmOEk7P20xyEIlzWlMrl/+523M4sEbUch13w2bJwGDWaQ6brwwBwSd
wh7mYnKKKLbP1/w/fsRnMwgX40e5IrhjoQJJvB5khrd2pYKF75ZKUqh2Eh2FhEGCnWbDjxRvNnn8
onT92kavIdSsUMDY7h68z0vs+kRY6zDUSlc7YjE62MrKZOIEjoEUVsu2zdQFLiPnuG1ME3eqpNiE
BCAG461Qe8dJFGbv8Y1GSci78olPtk0aMCS8fubd0MNpR8Uzpxr8YuFftLq+voO1Z1oEHuL9R8qS
332khFKrC/W7kR3ks6YUz8+VBbBCuRuBDHJtKvBXFzGgiQ+3NQpjIYj3ls/7H/Ttiu0jk4uCBF2x
X2/UUVy7fCytnojbLBWpnNA85oj3z62+ylv6JmnpkX9f5U901rrG0iB9D0DNGrdeu72FjxbEeJCE
Ri3wYuXFi3p2If1z1eS+9b9LrQzu/Pdm9Gj5Tdlku+4DFXs2HJgvksm8oePd8QxxxMNV74THUrwL
qxoEx33W3m5ZVaXSWsC/fhAkZQV0mgCZh8+XfqmQvigSGp/0vSO6DkBHNIJ5YYyf1WzSFEWNV7y2
plSZ7eD6cOhmvtrVSYeoVXbHnmQU2PHO2IXygVwAB7fq3v2NU3C+PsE++e+RxcHfNuAqZWH5x6j8
PxSkSuXWYf7a099Co/GIGS5prI1Lf/pYA6OmI8C27NoxZmGdowI2YlrDYboUtSafzNpvEow+T3wI
w5yviajRmomfVcfZwY7Ff7/XbiaWu1DcMCdR+0SYhH2d0bQfi4Q24Aq2A8nZYSDjqEJGN0R6S3td
OSijhQnzCbFCw1X8M5Oz3uiu2XJ7iYIjWHvw1OirHiTIqSjxcETxL2Kgei46PnTjymmGYncHx2E+
KtmGfT4+FWgrkb9dfvaQzWBzv8xps9lPlX49s7XnwBMIn3S9jhfuFJgu+JS8LOCrCUCm/eACdp/c
qiDNbaiKiuAcPw14uyUJSrfObVc99TAsSLPClEeZnD1B1Y1JT0/X8n6UiGG9+8YkmXLxFQpQsRgF
pGobOV6SBfrgWHcrjMQpZcOPAOKIIczt/eBMl1oa/zwQzKEv2XTdlB4fcWcXNiI8lmvUxZEk3hIV
/m2slRfBBMcNDhlo3RK1I7VrfKj8jza52xKGmxAzJgjR4F/U/4yuHkeUMPFS3euQBgAsWl7/ZT7s
w/E1EjaonvSnCEov9GlDiZO77Z6kpOUlYTmT8r8DWwYdSJm5nI7p51hNVzIQSFpRkz1u8mV2IlcO
SVdeChWQAurevjp8caWZVNqoTTD1UVFCPxwg4f1dLu/5hq4SMH8CMnSOOztYT0MNnzcNlRyD279i
mKt9TPDhNZCkdrBZxZI4FerrWQOyL3cBtCjtmCo/t5tk+aofUlOtl2XXJd5C4DIf7QUBaPmfrx0Q
QBphF2M9HK0DEBcP5CidqeMDiixh1gEDX8EAiVxMo7tVQAWfhNA6Zcb7cGHyIfDzdIZxWFoWKtKn
7TLu8KK4LYSUNZoDTOJ9KhZX+bEDxSud/lRvmLWy1skUbsHqf0yrjLyPd2MCbgFTYKm5I0qKkUYB
c2VDvM7THlfMmRyUAwu4GCKsqRMRHr50Uw3CkvVT2UH8rXZBvxR0uUF9QIfDvwqaKaYuXW37pj9M
0ZvloRYfr35lcW7zAconjZiT9s5QVsRdh/EKMVldadDyJNRbUF53aVI7FPPOBoY1jW30wAhiNjLW
jIgkW72iMriu8FeQyQul1ikk6lrBW1PoO7T8LnEFuG1qgBlUAJ7AbupzZzUpDHpt29iV+lGhw+gs
eV6uH6/0wjOhlws4sDWCwPQq8U+zqypSxConinGkgyX/Qz7VSQXvzu5uA1HpjBPWymXK0Q4VKw3J
i+m+FaU7Tqrj4BG5lDKwBv1HNGOtcwnRXkqj4PMCcJZaxPGjMRSqd1H09LtI5L3r/Q3dx4JKA9JK
ACIQzkBsA74hD2LMdRhOsTzAwvDpvlYIzFgdFSuPussfUlBOVSK/TnUpPwwj2rVf2Zk4RgCJqPUH
C//k+KqYJbUSErIVPCfxy7nJ5KB+jdOfsmtnMjXUT7Lra/zPbow5UL1exiDTpjyC4E/l9kSECHbf
RkRvSyrDNUIqQZh12hEey1qbPEjAyI1d6PhiPriR2VhRm3hFUHW0Q2EUbomZUauLCGeOYjDpAeye
8dS3lWM1clFZzmTswfgn9C2UMheOqCAff2t6Xsw2DvdCHO4ui2WvG3qyRyWlkDGcPSuJLR2vNGEl
4SZ0upJW+x1w3ZqWg8Y5Rm9dZIPhRbjqEj4ej2g4GGFVkRfGjzV3N20bTFv5be5sL58S459li1I8
ImPFYO4A7bwtmM6ojOP0bW7TdfAOzZcGZ5NUQmIBGjpObYWEZt/Cauh1GUIXqkOV1Jd6aHIMoU3x
ZiaMze34BY8osSqybmAgzmrcz1muj03eQv4yCIzLwuGj28yaBnJ3UQqSGK50dswxPcrgfqqhsEXt
ao95KF6mpgMJpdXgNtQEFGno9UAJioIa5RLhyX0+Ong5nQ29Biz/d4BbXsTE/ieNjJ7jIJzVYGf1
zOcmBs/TTXX7DKFczldlCTfTC25iupGEoH63/mlOelFv+gaDYtGP9TT+dUGIprS82/SrZ2MhrByN
7wFldvfm9meacn5F8jE0zHIzkODWojM792m/rjXepFvyKbkFirYG90dUL0l9vNCJbFMh59d6p4J0
GlmxpG1vE5FmS73fuY1+b6aDUGjIYqMuGmiv/445O1tSvnruczIc0G8a9hPHOb9W44wl9WtZCOR6
CRU/dlZhv1H1S+keQFVlER7IipXNdYA+wuuVQVyFeN4w9/sZJQRtHXLXf9rOCZtofTBdRroP6pJ/
fqCYLHUh5ut/eYplqqYsIdhwVLxpFaIo4yCD0511mqF7HJXkfEdZ7X0+Rxj/weC6N6Q2ZVCPwctn
DOZkRBPUUcUfXcvM+FLyl0oYXpQb2GhI9DQ1jUMIYvkg3AVwriKRPv1nUWs3PAmn1oD+sszick41
FehRe+I3CpiOWSoAYtau5L3I9P26HJR8fYpDsul5AXLonfn6aTyLB7/gaVgvB2Z90rWvG08q4aNA
5pxC0OD+2fkkDPBPet7X0ITy00QH2yvvXZpEUeDEVdjey7lvE7+F0NlEu8oEUmuFO9KH094/luv+
3NYKf+skuV/k1FKbuFCTyXsVHc2Lq8tzEEDSUTkDnJ5wF5GXUBLcAm4sbl8Fmxy1ci8qw8NUj5Sm
AO1XOxZkMzUZd4aauKmBdJjvtjuztfW+yIn/df8Ino6NjlwnJwwSdAZ1Za8q39Uq5VD5jmQHhqtE
13HPA8Q3knJoHjZFVPEbZUaVM6B/8F7X0P9zn6LhAOrpdjoiY/ySbF0XkmomnNi5HEYSaZGUwpPp
B0UUkg0Tl5Fv2i1t0VhnWKAxY7iXW6O95sWmEd4NyUmHU0nErLKvHWzWTIsdnb8MeTEbNhxL5UmI
ynfw08OvfrVAJEHpW/t4nZjw+Zu3QUJk1pOYIlC7kGa6TXFYMDFgyQI13+G+h26Mj5k393KP5HQp
f8yZ6yKaPbh3R8HLe9FZ/yRRU0mfBO5TjYN8TAoKAG3eciM6A6oC5uq/ba2eSYa9fGhfuHwYhAmt
+XTuAVmiLVMXwGwpe3SuL4oX+rmnf4/tbphh7abj3ROt5aPXJyeJzpTY7KEce/DZQu8SgwDwcFFg
rcl6fBhMPTcb1q66XAR7SLM9DfpC5oCslKT5V3TAj6uqW5CH7fEUKVtekkyd9E710lSPSHY9w/X0
lPsl/FMLR4FfTW9n9PjpbqOk6bzOKmdj90YhaaF18tFoOAOjrZ049WmrVYz+3k+oLTHxDk73pDzd
bW/kvK0co5ZIfcpOQ0hrBgj3EAhBe3at5XYuSegGdG2GQFIaRl5w2vImJY2jfgvK958Gv0vAemAQ
lFI+i3p994yd8LEqVUx2gL8VenCNrgZLmdbvlBeeemIt76G1VuQbAxBkSYFnNf86Eun+iTmbEOF+
Mev7Jn2zv4rL95KVx/zBveLyhMUvGXdurGCzAEnS4W761ktlgBitto8rghHUECIXFTO7SqV92Uok
E7c6ib4xNZzvUDJcrw6DNqynJNgK/GFlB4gViIQ748H8e4Di6WGZz/KFHDRvOTrcjBRfzH40GGya
zRu671wbyvrul2xm6fBigan+YFsUni96s95U6aB1n97dpswyX7465Z/Y4GG8n8/zuQC6XnGyFiZ4
e9vPkWeUChIjA6jTzf6FTy/TOEHWDIY9PDpjhgPpxMfroxahnXT4L5GomR+l99sDjrIUDAmCRCaz
G2jWhWmymuxbBVBVo7BzwaRhaXeBOmo7kZ79CuU5uMkLRHoCrgQp4MINuXR8kmYEw5sbr4mX0keQ
wsWIXxnicFH2VxUQOAuq/anm7w/oiZs7UnpFBouHAXrZ2SKbc1qaovUjbyTjVF1u7yrnJeA3cNpc
/slNccavy+QXiANBNf4VxnOj9oEMML+EvnTUd4Sk4x4hJe5wk3xOFw1+F2r9uy/Vwrn7hQkqebsm
WjL1U5LYs4kndgoJEF2uWPqQU1hqMgB5d0ynLk/MRrN3SS0AkE4EHCJnotCJ6cfpDQqiZkuN4NVR
FqL+F7D5izxZ/oXZgIZFtJrCpLKnVSY93q8GGfagsBvkrsx5GbkHP0U+tcA8l5LGAKSVKv8BF7o9
YooEflioaabqjBe9Yl+lH+otCUanl+PuulfYws+s0ngy4FxIIsBzAmGJs4muSYUsWKEwtEXn9Ho2
P8SUeerRjQeNwOIKyI+/sAxsPnNUKduzrmTyrHkXWcRCEc8OxJ4cHw3uCBp+hPBR+Pj8QL0rFkVO
VF9xcat1HKcCDU5glZ5bk4KsyoMoEy2tHpmbCtyZex/x8JdLEUG77IMi9C65OWQz41hLN3dSpVKD
zXNZ4CJKxwy5TsVb8kgR4iUzcoIo/yxnYFQR0KTLeghZfwKP/FuODNcsLCPJF0YN+VBSyOTRJ8PH
AJ+YJfFj/7wgWhlvWcKvsC/cDdISfrJrLt6fjaT2sSY3S0lPxi6hS8xGITp5N4DSKRQcaxvaOTUK
frRbsh5saZugzggJF0xVfnTp8zJJrvw2C/fQkf1meAhaF9Jsyg1/XuyTPByhZgT2dv6Vdz0rwXPV
rsV8iQsjSwxw6ifFU6KgHq+/7fWei3XHLPfH1y01kGyopi3gZacq0IOlNibP13Dta6jDqJb++Ljp
mp4bVd1a0UUqkksq1TkAVKX6vpO8Tdbn2/NMQkZyCZZb+dplAg3RjFm3aAHeVXu4hXZUgvYhg3+s
ILoiCUKE+aS331YjgtalAE+UJj3+MDJLa3pr/c48Wt06M9fQO3DqyPBq9EZEffcIrTz3KwJ0OPYd
aUye3h44FBlQVOpje+Jl5gEQQiM0/MyxWqQJEKKghulZFLx3Ndzmyf1PpnZv9Pw6lEgWCaKUmmCr
//9xXI10EDM895cMj8gmLlo//0J4pwgQXEtwMsx9wSlrLEBd1gWfeUxEfYn4o2TGH6hIIBfHUorE
RCMtsK9Iqwxx3SW40cr8I1W8jNzkTX0PN0oZ+NMqMGUFHbfE314ahID6Mg9qcYxpURe95w62jHzO
df6bIkcZ84aqPoKSi6FC/B6QrRb4sJu0UiKcV1G6/Qso2yFKpjo5MQskKw2dT8xQSTytajmR0XJs
8FQTILzxDQigbBiKjYhZQTIBrG59mEC0Hi1EEy09uW/0bqzA/BbJS8LlkOZoPP9ZUNU1YiribV1c
0QY2BpKad7641NZsx2MsghW3TaW2XoATMLUIco73kAtG99EwjEGrhuyfQAaoMSF7hfAJEutJbmja
P3QgwfNQ4PW6J2Sjlw5mq2w1JdtTH0keDIw3pHu7rjZcRH2HZxBiy6anSSAzWDYH9r7rB3J6s7ze
onzBOps/b2/8ysJjtQwRrXyCGe7TbLeW8SJBuovK6vvZfqE5VyjVrPtk62Qb6H1KXptwUBct/ns5
e5O3vg6cQ4I5OpUuUqqnghZjIVh5CYYKzz+Jls6nGbtuuRUf5LX/tX8FYk5o/pE8GdmE2pYkw93S
P7GOQGYEGpTaRheBpW9xeHewyDw7oVQHh4ywEkHpgo3Z+CkGd6CqcEYvvdCRW2K57n+UqHQaup7p
brB+6Dz2gB1irF57TypvBXoAsDGv+h5V61QR/cM7TU7whV5b/3sbCbn0nOY4P0mbSA2fuNJ8pAnp
64c6B+EcDBdYmC+ABjWbkk5DQg+6oHfYzXiBOOunBKsZbMB68YQDZqyAHIufvISjo//h6wvDoGuq
xorkVCyZf/Cv0w+RS4Qjt6zOR2IsXPMz37MmET/dPm1ZY51BWCg+gFyfrKm5UokuHUb/ONRhJG2f
WL0SriRwB0SgvJMScy4i1nRKVgblrfROLE7CouNaJ3P7b1BhgBpzdyzhLLIh7gDZq51EChXO+Z6S
o8cvajXhr/49HkoiCEFZcR7oTAfkWuOfu2wkoZ0KU+vL5V2dtWvy33Ix4sk48B2iB6a5yzFloQuC
stKxPQyYoHyMOoD6cqlCHxhcJlDii1cIsM8ToyppCSTf9F/iVQXITm2vOs08pAQ5GA3O3QT46k6i
zRw6gyKqu+MTqdQTzhKM/9lXXo2nkMHoQUCvxHmbZZatJHCY4fBJV/3Alk1M2zkkiFC4O4zSKyeu
iCQzybGtgxX1qGgWKwK5WViksyMXw8/NQB+ZRgXAM1TpIH2dGINTkovaCJzlOZQKIvLVA67pOakh
p8Bxfj9BRy7DJFVDYqwSGTd3zfFJFeB5PKlYmR9cJUBb1OEqBp58S3ag+E/VYpofwRRnURA5VdPA
/SCo/DiWVXokHOhK+TWfFD+xjzNfPEAOCOI7z5ZGxlh/CsMGk+GuGqZGu2KE7ac83dsaXOLASv7L
nyHXVvivMQBVIjxf5mqhQnv1bKTPJ+irLGZKD5UjwuF9pDK4JFdwfmXsco1FLE3aoh/BhK63kA/a
2EZ939SWxwI3pq+HehnH8PQpXUP317/nibT5t9H0WjTinWPxfIjnssOPlBkiEdrQLQMHzHtLwgX4
BXQqONt6veMLc3re4EKd8Kt4XGJ3eF9tzUnJVCCAvkim7u5k2aYCgY31b2CWSFuZGHaiQ836Cw4+
FHpuqQiz2v68CYobpGVPwEg8pCTpE5bS04V5+sS2odhkQGmI/SZQMtnlLjj/vrUwBEg4mlS/0DhF
dFW75LUrSwHzJ/H7HNvVs7AvoeMVNo41ghVsEarPHgT+SyEpn9f+EdTfyUZMNIuz/2/gvi4aieyQ
Q7whuubJ2Qc8C2wt9DiD4qE7/QKNIMpT4G6y6+QHlIlVR3KBE+vZxdZT9nk8x3DSoeqwrucl/AsK
FE2HRAZGPFvbttE5V/WKDIFJ1NqkL9LEOiYQHwolzAEPSIKGCA6JSC8D5AinUjusUKXhuBDJF2RC
h8j6mfUddiwoCxXLSgMqSVDrE/92bafttF2tYd0R86+C1JOUOMiiuIH7mZQxCdj8QDTowrXIJu4m
3iLho1Q1P+I5U9h0ow8CV6kgPWTxAKQ1w+PMVToCv+DO+sBkInboac60/RWrK+ubc4eBqHlDVx0G
9x1622Vy9drD9SS6kwR+URoYz+VYizwG/0L0AJ1BnA75xfcs1uBN4AQZtq+EEl5yn0I/X1Bhqz1p
b3nia+sSIr4baM1AUj4r08avVFStrCMEHRXFAZ7kn86xXeq0ZcwkAnpyDdcyDoarbH998OPdmb7G
F4e1S9DzQsefJCL+QvfYOYzC9KoHykQ/W+W+w6g/laMmxGZNGKg6/0mrhXNEdXYnTw6rNhGm4KMh
jr0TiDB786cyPePcClU4z3f+3vaVYXuD+C0nGriSXPjNSQQZ8vRqUo7dyrzdobGItCfmLl/ejKkZ
9VZLVwz8IfVVtva+EdmAyF7R8mgyzJFj1UpdExE3TZ1lXIifPchM/bulQ1YSkUGgxXZdJ7UrEAMw
O7g8QoqE4nOZ9zOCGiJha8L0oLThC/UiOfUfm0ONtk2r3pMKtLPMdRxvHsOyIl10kmZyneBxdvHq
t67wJv7Sdvwz9YnWnjnnCBaGVtEdwDEr1WqkpEN8fosfI8glP2Z9M9a1kRSaYcqjtcP7JfiovyO4
GkSy9F/uWmUTEZjqy96kPjTUGFUcrdTzaEUyuO1oYnaLy4hS6xH159Va6In18Ys3OGnq1ZSPH0QN
zqNDeLNnNNXn1qmAqK+JYFIgjySAEZEoHY8zIT46LmVrFRyL0drOtUOYWjQ/Y5pCxcm5EH5ZfhtB
PWv/ztNWYSir+0DtKyfgkFJ/ExeswylfY6bmLzA9iOCo/XOO8OTQrX+BeaL6JefCKqB2GXi6/qz0
SqUK0QagPUF/5vjj7zBe7+mANx2FALvCUNkCC2oQKBFJ5liPyIc1f3EeCWI7/pLwrSTOSEkWKDlk
hJrnSQcNacZUWYQH7FdrdJQk6PNfRFQOGg79QZejtx9AqOQNWcWvM5TZTsQwaFNtGb7HZduhEGBv
AQtGCcd1h+EkKfM39yqJ7rzeQoYRVssMRfhRmnzQsGJ5nqX90uwhWWptyS/YyjxvjLPn5+xbZFic
8cNfxh7EMvzG0j6fvDGysC/lHGTiZx8wB1Zc82qTccD+dGbKLLarY70zdFMvxCYW7vzmUxhu+IAE
WqEtTEcHhcFQpIDDc3WkvcROrqmMWReAUoX7i2x5eJYXOEjx5zBQ9ikLDB5ic47VwJexxxWwSuJb
T+sX7eThPIZuBQ7UC62BKYpgHdvrwFtr0dGJkA6BZK/uw5qEgb5pqg7nHc5moMhaU9m1Qh4WSufo
U4o17m/u9XMAP9jkQzvx5y9IqFLOq7q5szKqM+d4AlRFT5iwngg+PWjyKXDROz2uo+26JIdIUKRQ
oEsiCTCQ+cD3nF2JHZ4xiCdCr31OzDx1cbyawAE2gZpQ2tmJEyONScHBuOdKILodgh9naDse+lPN
Hs4OQKk3OTgRYUqtoH+c02VaKSkIDLVfOCWQrbcJJr/VWJ8bnRaZE2+Hn/Y2+ukRe9/06YVJh5e+
FQGpUz3VdSrHqfR9DufvvNbTQgwmGf4R21QuPG7RBlu30dwK6msIAU3gKJwyzwkJ2smUAQuY0Yt4
NKzUuKz0brMSYvZmSy/zwe4etpTtowvrqg7GCN0d6LX2eQtCfv84Ba+cl20XhxcIrPWdUFPFygAB
C+8ZyB/J+zaM7UiOEwAU4j+iqxEknI7ynn8qZCX6q0w0PeJv2XEkiiig6VXFiIVXmI7TVKrXB4FY
RRb+HS5gUej4cUJlNUCglKFIgh5EN3k8IA3hzmxAImKe7WIJ24KJVuCW6S3e+LkSTj9k7/Kn244u
+Dr+sfaCQpmHyp5GIGV4wK2ef0cKx4hxH4ct3rUqcNlR9bsqscCbc44FnlBHudm9zK2PCsN3B1aL
8o4yNVj8MRLLfI0MAbgW3x2iWikwSQqJzSGJSU7YLovVgj4yz7WQyfmL2jABoEo8XFQI0P3nrghf
gH0ITIUSQFjtVBCjsujxOOh01rc5M9PeOzs6Qomu3/6UJlMAU0OdWQGHrkf8LR9IE60JBWHTvPYX
0JKUTpvRpe+o6J10nf+iuCn+nXiVosYRE74mhIuWPUKygzhGElpl8HzLFNdSCw0/7udNUDuIvpik
gjrG4QdjXXkUVt3giXGRhWX3gPsTlYNgJuW2CTqa6EVInCQQ3zRW/YNiQdSCfPg7lh8lFMOUslwE
7YkNiyMnWVc7/sRhcqycxHzEOGXdTiomgQPee6ZM66NED/0dmxaQiZ+Ad+BL/n/4IAWsmX2jvzJB
8ScGdm+jwk9r9O8zOErfonXcWwYDer+fUJB6LlPGMBNveYSGlkfEABkkWWiIq89fnDgGRLF1XKCZ
YGGS9RB6zoXjwLk0Zx7EozMYQ6v8s28zC2p1AcxXTfZ62kUbx+xFAJjddCkt3KqcApXN5Z17aDu0
65E5pyuYuKIEt3BLH7BL7NtjDCBXm7QihdKYYKBcLtycnNOPi0mtZr+JRGDbcSNcep6B2jjTRxo9
hGRoe9KkxIT4SbFz0yfAcqul1WFLDmeZHa8yxn0Z/O846GlN5Aq48+PlhOtgZx4ZVl5dqwxW7sFh
sRJyMFa9ETuXGKHs63Uh1FIh25rRA+Jck1Q7IGNpEZZw2U/FGqsgrjRwuHixGxD6FPj/sSdTTNHF
aMbZt8Q+4Xi9O3LPcjSNOZ4tbzo3JC4s3DIRbO3D70oSwzmSadBrEO0FEGMhcPTuVxjG08I9UmZK
SOo1PmPeZmQdr2rjdAo0Zd36/8iW3aSaNrN0F1fDe9dsJMiN8eKRzw3ve8Mu+EaSxO/2FqS41rxC
bTnOSFmgVP2X7Pl6i6NDmzWTj/MP3R97ONAkqB0MaTtkP6Vt25zo6vDkB7rwCcOnvE659YFsOjDd
2scUy3kMp7ev1hPnL5PubR3EAKq/xXiWjoekHqv+iZbPXughQ6Z8blCuHmVFB+68B59u8kJTNoLQ
8tY3DwobiEnOTvU3D04Vn1gL19rS1bI7ZphqC0tzEJxOKOX/YZXG2UCdrCbE9jQpW0boGbvWINZS
UCsIxX0SJVzD3pcJJ18nI9ZjHvBKvnHW6bc6yGjUonWSCU07Ns7jqEZ5rlbnGAVsa8tc36c+p6Lp
OrZZRWsASWvmj/uv8C8tM/kTaEj9GtLKh2JtZF4sFwCHKGOnA1VUtshzwuccDypUdkh0GIi6wrod
n4L4GA1bipJbRv10qxrsmCuICKiJLRDFsOXeG0hOYzjqbR9Hs4glkPrJgietD7M6GNu9Y6+F+z+B
tlqKMRZF1QRCtUjWdPKR3wMZ4apuCMJfz6p1/WoW3hHtEHRXC5YcqlEcEufK5wo8tvULOTH2w5d4
f5W970gp2vo0/czQN58H+FPLDEilIQC21TmFfyx17EPgcNXvi0hA1NNgE4y9Zbd44Gp0HjdjvLoL
/0pkoBQ+WaHmX46IRhsnBTdfBq/Hm4kDVUt1nYdxT/1eS0eouegGyT1t0k5/OuHQjchVX8JgXFJt
p6CgAz9TSUc9u9z1YEvDsFUayiwoWPR+vYhT4ojqDqanDy2fhkHgBTXiPSOUWiHoPMNXn6rHmJTS
bXZySzW7vuisTn8iSXDpoMzn4bMB4lpzKJzr6uOFZOXG1YcCSdxuuNKMyvVUUKwhAYEaDEEAcAQu
em7FzY9h4TYMlSZg6JVaoPk738QGmiqiggvqoGuvn393HrYKXsc+bghLhv4i87aiS77nT9nCelD2
YWgUIHMG/zDKv6cK0zFYPalexkFTa/2H91LXIXU99SwSppmmw/StqVbyD0md32/anc5sisQDFD3x
tUkhYP4CVBpIEYLydFz3ailQPkyAJczwitNtpxYnPPQd8kiQBNeYyvIdtvnD2FSyy901D1qRp2U0
oM/wzGteqamq6hMG8O4fsff1Ibq3u4p7NA8c7oHXN9Qc6XfJCTYo3/wLvvUu9KXk1VhevCvcu4Dj
kPj4uF7FeAhiGlLoicUBwAiUCOTZDsu7jZ9B3B64cIGhE2XhqhLc1KT+5LTGrVwgCtiXNQGlCmvt
7YtYpobYPd30ePLITafD4StpDqvJzU15zoY+Aejgw0WetR+KUCvt4bnlC7re9EkhwjeUjrtkDfiZ
24TvqE109k3j2njs9odSeIY/607JhnCkDNq2szTQ/lDrfZTtDwbLuQ9O8x0P6mcyKSBwLDqL8k7D
QF0DWZhK6yJe8iw/8fB7C+lMNupTgOGCqr3PDsHXxAQcx0G+mnX0lvh+OwesFWQcHuQtKnaE6nzW
twH/jtUQsBOmcQ71Z2CsmporFlf78r2BAB5++2YDVFcIcNkcUTNHsTl7lDnilwct67CH78wJf+0K
UrNJ2+gqCPw+dsEw/qMEh5JdKMRe8B6eDxYpyYVvAiXMzd21yXYU5Bmw8td/lR4NRmiWmVIHH4SZ
JSdCdr3LaJ+ZmO5j29DtNh+0LbThjpYtDReg5KLSMU5glX+jJX3nSz9OYTxQp6prvboE6+ldHf98
+nJqZzf9yvRysQblZfW5147Whr1ArPqGXwBTbe91Vmg6fxEpwl5W2IUAJBDQi3vNBWzl/P68qavO
6SRwHVsCNqqrubuPmbxHbESg9Tc3VeEdM/4B85t2u77bXwS2l6hHZZsuai+NsXRxE+KDbgnCuYVr
9g1/HCezkQTPRcmgPvOUlzPG7m5E8YYvo+XSeTE9o+aq7BlsEZV+kQwH9fOCo68D4VueLhYmTWXZ
SvGa2zHi5IIQEC1kU2Tfy4Q5+cX95TA+idwVG/NZfYouSj0Ez89JG4y7qcuYeeF7kuk3IX8zci3l
ujl5sOnNnssiuJyKrXMLi3rHK9w1emmsCy9lAmK9qdnpOFthFdLBjmGe5nYlwcrIBHg+zjW2mHzG
7E9y1uwqDuNhzQXiZ02yDljSEITyUgQrKw9l5zSNz3X9sYy16MS4UlvFsPa0jawUjKCR/c3ZqhFe
4pYV9g8FE7rI9eMi+aANb0yHrjWiQYMRc3dRMIo6/1qvT/FC/aZfd8b6KaZ48V/lyZnZov/aivhB
npV0evuHw31ahxzD6UzvUGHtFZRmhuzWrT5aiVNiPB+YhCMsgsRays2dhT9gSOR1YPUmzVbfyCMU
wgjq76LEEVnqnrpZEIrylhFcEgDrxSAs0f0RP9jjDsCY3SgnrUfw/ZBmWde5yfcoHlXU21yadV4c
iQdVgTi8PPmDP5fonWKJpJmvwsGzvfmpXuTvmmK3tE+llarS3pTyD7QTeq+kCDgURUqGXcVlt7Cq
n3SKTlbtHk4+YfW36dK9vmBAETVKRP0cDT5ogw5FfPAgP6NkXeiymWNryWSt6+SHXzMCoYJd7CGg
Y1BswvQ+GgV2s9Wa1et/CTkWT++H2KYQnD5iPNqYKX8YYAaVeZNLNiYCUnVETTNkUV84hk/M7xI9
rCqqdqr5e0SXetzOLGLxCngtOgdQLszCUxMEXiaYd4rZai/Qg3P5WSPrEY+Tpnd1zLZZ8qgcrISm
CT9kMH68tGxt3XVAZMi244QHRrybViKqbp4YbbQlVr+c7q3Ne/PGFLlsQXJix6OVSqJuFRJpyVlK
pXiQL9Z4I5notUibEJCZg+MBVbIyGXNLWmVnvkr3Xx6j/KoZQedJRhNihPl968iN49CX1bPtbek+
1yUJMZ771b5qqocBEG22qJGgGtlL8pESWbvuclEloA4QOAS9XezGh+960L6+M7lqyYDjSHmNFCen
fU2+hB/YUcxthQjQbCVzdB0us85rhm5PvgIk4d8RCcGn5QOxTzDqAMuNA/vEQrVuNAQl0MRJd47K
B/AdBBmXBTsFaflRCvjOzltCPN8N3tHdTB89hVxGbYLoZYt0y4Jhx4XCG/+fDoyqLHdczRK3WTz1
ssYXSYm87xGb0uaa/ENhFS5+eFn0EndUtd1B0fiXPNFjBwSQmwXV9vJQJfgZgjLNwhRHsyJylTT5
PVy9maAcrhZiNTt5wNn+uEKXXJAqCJDsJJ2blkHguBAd/5em4inzBWQVXu7KAn6G50jvG2gHmYHq
Fg+FPiS5mGZUL8xE3szR+vMDbfFN5Ntl3ueD4qwpANtSeDT3PAqdqK4O+sREcBd+zqwq2IGdevhf
LCm5esG/lfAwR3PetOlQsK9LIm02jYVeAy6QC6iL9HLNBO+I2qnT3gqeKYyDXYfy7wteJbhJHzrI
wuIg4Yi8SOK13o//cn/1r55Ze/rCveTAP/xNS6BNXiTzt8Z3YIlPPCF8UYuIFMhKZxQxmsyucfe0
zAwmAhPTEYaaC2ItPm2RgOsTXwJnZg+CCF4sJe5MCozkDp9aV1QtcdCx8+Gvknj8ejVdjgFGF9WM
BZ+jZ/u11JeSGMGCalFE/X1P8Y14twk+j3W4OL+/ng99eIw3SCqc2NtnVDC4CBy4/Lm9tAXg2Otx
T+WjAIPuMLGAl6rWP2QW2mkkY0TMb+ddvhfjqxs6Q/wfQ4lTs8KE9FVN/LebQqQbZ0WpWxIriuGH
14G2acPygkAR7xoqM1KvCNJeYHr5kJvi/gUCg1yMXINEQEe0vaMBNTkTzANWKZjiraGevXyYwu5D
R7qLcgdG/jvoprF2iJ0fHBBgFVxuFQxcMf+5CnM4BHgXztGFJ7TWmyy+p7Lk/0nDq+rKDuNXZ7MW
uhE0paTqoeXa+KvOwHZpqYqygmuAwUfP9pQFDJnlbzpu+nuk23JS3UYNI+0uu6npA/WbqytBMG4X
5d6Rk4DfM1hGMcojqGfPC2lJtv/VQEd2f2oW9nKXhImg0WSDjxoCi0MhtdCHD0hr5hlQ18qHXyuK
AHTa1BGWkLRFkNozROrWLFq22EInEzKbfNBm0i4K8/aw5WcsxzW3u74MbVF1Z0UoLD5xARHnuGu8
CxXkBzGMD9bE/H5/TcNi05T9VLLP21VXTZLufGRqGeCOn1Uhbhw7NKdQOri7WDBSOOQhzxueLiGs
OgGX+3U7RWWVflhKVD4w5pI9e+9iG0YDqRKLztfS7z2q6koSGAHYwHJd0Y8aqe9zX6hTn4K9QRvV
1YAoB24oaiO3uEhCtFeSHS6i0efashTjw/StO1Wx4ZkcVO4AjCZrSXZReoZcPCkiUcmtjuRA2znv
uR6AXQ3BxRkYlmiT91ZXVqi01RUGhbiNoAPKoszRbDwEEh839MlPC0YywS2yVPZ4f72fJKnCr32U
SYeDCQFVbtT1O8H2N7a7wXCb1drtEPaLAc8QyfzEk23UkW2wBmKvH7Gqh9+N1vmkvG9b4rebW2dQ
9JXe1duGngRW98bBVTD1bVnDqMoPlVnbYEZMZprwsCm2Bl/Q4D9C9feHqS38+Z4Q7qKF9Iuv3Eyp
p7YPk1g30JHTaud4qQMnIA37ssC/gXDNC1f16euzfpKoH3/zRq/Xq1ZbtGzpa4lB9vLoiHGVq91z
YpW9OTKcsljcY1DPLO5bqQ2w0q++UYwPFmkXsHTbcPw8Wh0wyiXgLIe+ETs1p85i0b3s1JbDjLXD
T7mRjJGj+MYqwyORG1SrRe5T1bi6UquAq26EokrATmsZBopvRPjuUQs69nvu6NzOuletGNVfz/8c
Jw43QShLQA/A8P+yX/6ed67XBlEwnVJQa1e/KBVlS2JF0vstxRii1Me/OiThnj9zAae1yTIYJFYb
aIR6Vl7Ptbt7oK0AMX+PcmF1kW1foE9422zEUVYK2bZOcN2XIm/OrFqs3t+PQtXbTzgetePH4JPd
S8wUM3nF9mr3YoMWROtfyWtITQBs/WJJovRRWN7DuHqMrmzuLEbY5B49vxj3gmSIGVkFSZAUadFP
n7nj4w6fs8zlhlda/APlqFjdtBwEhd5Ou/aC2qARkcVnlsNp4IY72xOiminpUAvErK13auia7XVK
6kFXp5lmo6UwSRnSIlYi0yMXKKtC5FsdLWgl/sRN+450LbRfbfDaZbJdrotylvy5+/eJFBgsBAPG
pWjJU0HRmskLnrWt8/0ECci+xdGGMbJt+8ff1VJX8Yphd67A6xpC44ac08WJV0Cr8YkJEbSozGVA
BcxsOq+xiT8MGFcFL7RtX7WOvLuNuFDuceuk7idiqvf1TvPEl7MERDdZzjDJ+adTUsHXOlh5wJ1/
DYswn0SHg6PnxXGyIjs5jtgHIwQUUOGAVI88/HJ+n40UFvs7JWR4etnog0wuj76HlyUGiZLXvJ0o
P6yoA/gh1G2f/AJRalL/i8MfZ1DBjterIYxO25gYH3haOyqd8AEkXH5UqMGkoDM9o9I5aBJoYkig
2Q+wHhO5eGXMLSihZfsb2+MlB1mQpvI9hM6o+90sVgf6VWexL7aJBc7Qu9gNkSDDuIYdTHhZqNoh
NnHz6cCHdnDGzP2AiWOgvjUTK2Hmr8DMNl0wrEmVo0KXPdOdaRepHZL+0Eb/4YoRvTJgPnbXZfJl
mHnXJ60IVnksLhJMsWoexUChISAp+qswYPGmwVft7Ear9gDQXDpdGtBD/fKARycJpr8cpviPJMtI
s69rwRSkb81CjPgq5rcCupQZknt7wx4a9j2R5wjNgaTZZgrhwLisMhPSR2PyFfeQ4N0wRNyFph+D
NtzJ2+QNCCHr4tsqT/4qtaIYULiT2216X+NZj8c9oGoabh4y5ztQ1MD/jy/SUvjmJVjNT+BAB0lI
glUrAuj21ib1pco9aXKovG3HhWUIm9at3L/0on+gkhUdjpKyWG3Thk9Xhx3Bys/RbbvW0eh33av8
9F4FSiA4QQqJMKnK0cHKFANHw1MyxLqjZXy8ZPRfq0u2kw3gIZlcbso+pb5sraQtTzg+NM2OgUtT
MiT7F052Wt8LSq9NmQ+W8gK7cDmbFFFkiZQgnkLokay8FA3lVTm3jRkNWmxCYsuY/oLbIU82xJlE
I7JSAn31r7akEw6Q9ZSpOwl0gdgf4Rg5CPw8kFO75LSFbK0czN5xYBet88jE+jTH6NiPPmBJsNDF
0UnwQlIpeeoHkoR1d17rJcVuaz7jXLXRJn0XxS//Cv7ZsHO+bLnVWnfI4Kw1OPVjR/DCNrOU3Tru
1sdFd5XmycwlXKS/QGcvRpXu/97kpO/rUYhImA+LhcS0xQ9mhln0BSinBTwCT7Gcr4j+gZVHChyh
Tk6LlxNYck8u70JLVmORHJ4o2Mti7yMsBT8a2WW/NegcTpEn/H02bqxwjIwm8avq+UD31x6OsRAm
Z1KPVRKcpnssNMnEI7XQ3ByyYhATEhEiLacjpP/ckgjc8X5G+TS2YP2jPXbXATJFRK/enI3MxsCP
oDoURDiBPEJXgUVVJ1AakGLGkiGoynS0HTkR1o9KFfT/4gdvXUKVu3EOyWcy5JZJf8OfjuzlZ7rs
W+eUXlH2TDghubBrz6dF7Rg5DwAQGY/Z8r6jWJJQ97idKyLXB6k/IFNKZ+R97winZVecpWuQD8Cl
vrrph+tI1HeVJOrJ8rE486YP+8AwvLgPDDmzVlbucJEiFmIbTB/CsO0LFEgOQFvPZkb0DPoWD6mp
XQbrm/YLwYXiiMuiM0bEg87Cl0PCds3Gx4iwoxX5wV8/k6uyrpPEKE9nXczO+jGgKvyJ9ohsnoOU
fdEeoRQB3TBBou3xDCAVF4Un7tH7UovKweYrKTdRHn2AZ5sNLphTIwWq4vMEPLX5NMJANvaJz2Yb
FZTPaln+k9rV0eRR1aSaNzAMxSWm7aC7WVkAAyDwsJiNU/dlN9pCg0/mz9zHyeZsy7IeALEdRZlI
ip4h8+3r7gAxonggJxU/HWdW+Jbv02oTCWiVo424xUNtZPI3AbzGJZySRw9BLdXQi0pv5fqA2lhn
zTuqkhweBr90nZfIss+IROd3229eUkXnWzy2M5nH0aDGAOzwLb8VefohPeGLNigjmL2VgNt9+Xmp
K6R3/QNaJPw/DCI79AX9Kvt3z6GVVKXMrXholH2bFI9IXpwBUbVfGKNqzfQ+vRRnf0HFsWbdYaSK
Bw4skr5FtMi7y/Uhtf5n3wWDNJ6zEpQza69YS2P86/WsbJKM7JXpt81HEC3baUlrg3QcxFP2Grou
au9+lnEgULsP3Gjkdv/VCn2DHolVJNgnurhTD/iXrNgBWdx3yWhSK64u3UuN0e+nFmC/b74bTiJm
EvaXFUCilEjjrcoin14XHw3GsxkNYwLETwhDdNAZWecouIiyejX40yN7j1WjG8h8QVuuXDzXbrHi
g1BeA/tYiuUyqvq4qPUVPOpTBJCuWt2kqY6sSgpWTtegPQ7m3nAIKORoegEybM5JXsrYgN7OxxGo
J/BwDfoS/Rt2bMp0t0U3e+wj6mzK5B0n7mG7o6pxlsLRXYU0bnqIJVxBPrxtmzhp8XBMhK13SoLZ
lgjKie2s0RJu3X+7PfIqHCY9vStA25hSqPPt0TiWFMp6Y115R0CxpATdjmDpCJnMtoiKC26N39ir
sZ1srqK3jGo7ddyOmzZRGudfZuts1nsnadO2p/ne8OH1TXnPpp32QzYUlItVZUDwtFUKBBV0eFAB
36j8SV9oIZ4FL5A/ckquOlNlD/FeMZsbOHz7j2sQCORyGHbIluwCnX0oPccm90pvAsP2dbBLMncD
9WfItdOJQu4aTsK88ms/L+KW5n2hQj4KbPIzl3sLBjbGoXpJusxNwjXvbqk3Aw4LMpb+AAjOzVRW
ffVHLhk9dXu8+peq2ob29fkSNy7Fu2HUScYqZtmjoPndv/5NtpjmVSN6bBB4nCctsgaezkLn+2Z4
GKM57BKA97RRPhUz05DdIIiSDkFsj3G6yYlwCwlJA8c5jAfuwiRl5Z0tvmwhCVIfBiCJeH9D7RKz
d4CC0+TwZTWGmCIjwIJE27UvKbPIHJC0Fb7N24FReFIyq1sMfGeIhcuIH+qM22E/TQtvA+KGu5XW
tEqzTQcgiLocun0Hz50jwgcjdmPWANnUC0rDUCRXh2Wp9KZRIvAbu+2grp7M0nFvJoUFmlvczAqM
/LznhUlzVKocujJROv5jKkAK94mkCRunETgPgAaG9LwEddrGjJTSs6xIYwASBxdxK2o2wNjPWk7b
May3+AUg9er0GQoCpPJ+8cmRvFS0AkOeFb1Sx8+amxHlICnN5nZ7SEaT/FE5DEV8PO1AxnBomExc
++zsNdI41sMMirHuPbcEIFp7ZNOwxd4Sx3Pj5hDcYGAUU4+qCgNXi4etuEXd54Y2POEFEvpQZPZ8
ljPpksku2oF+YwUMnswnaCVSHQClxO7SjahY65gmaA4mB0c9AA+NBOmAuCKXFvg9nE/qkojKHBJU
9uermf2aaZktueim/P+h9krBjVGAhGs4kt1u/v/L2ZO26DYLclioOm8firpMXo4X6EgDNnhDMu0k
pVkW9cpXeR9R44Ab2R9/aSW/tUNoxLR6+nROp/wfU/obvh6Mbbb3fzwASg5cb39qfnhQu39SkatZ
F0gnOxtFNkJFc3MpoXm6u0BKjxJgYWvMlWToVwvTlAPJvp4vMeA80+d5MXLYhFlgwhv7aQagdH5a
qKn9zxd/WH7aXpsE7L0u8UCcsXYGdcdPjod+YZtJKoSIc05QFkEOq0CjqiTPVUTD81717Om1BqYE
R4GxgnA2RP1+sxnDNDpKop1kf4JN2xHYvqxJ84kPSNqv7VN9ommGLzPE3T/I5UNQnykfJ80cSw49
6nUN/97LncmSZb82EoPohhAe//s0IpWcVSR2U3WjMTS7yMHJTv0KFvwP9yNZslp1VcoClDEoD0tZ
kOt+1Bh5dlP02gAFn+5c+xjFD9CFsEaqhralMMOp/Bmp0PA/q56cSLt0F1T8YWRbf4nLecKv7cHQ
ERO38hyD4cuHxAwOuYztl7bX2KqG7LU+7DKhc/HH/7T4TjfM4V2t4DwoJpLqGJNvCt2I8yCpEniG
zB0yYnsBMx1uaba/Z3irvdbS4d9aLHx3Fj3kzdqmbRyppPQMSk1+lMpFOm5koqGLK83JrWF41zih
TmyKQJqBwmEdOPkPGZXm1DZRWaWQfg+az25Lo+UFvHuTdnt+XnL/5guyhkF0xranmyKH/4NSES5Y
0D2zGX3CxqX80hpEhiwXMWfEixYH8oopf37EfQ4bCxFBS51zrr6aek4E0pYioyeCFV9q+63D+3IH
Nur9p2JInvHLpv4B9QFrsPMPGRvZr/FJqkaZvcVF5u2KCWB6uRPhjdBaHCNaTq1NlkiWn/+awVyf
i+lCzF9Lb6K6rj7f30zGvhZBAuC4ev8qCTSIwMQT2L29SwvMLqlQFWLmoyBXIqCyEcGgotYjbDf6
OiJMEDn8JWFpvlCJlxGqvOA3Hb8rtNJFz2gEFRoK8YaRMOFdICYnfmv/Nh3699f4y8nXuALHfLUi
9XoLWj6HM2v+52jiATRfUHXBetObex0Z1Rtwp76bSe4bsR3CGAw0UrrCzDWfFegMJCj0ZPwvBkk8
m51SNcrDpuoRwvnPJObUK3UybHKQZdXFBIqj1ABku2r3n6CLOJoJfFLy/YzSDlPrsAjw9hum9no1
NnOD2caxotT2zN85It/OedwCqr+MUhCpko+uRTkcStKF/u98cE485A4z7IRyCOfqQONhmND/5WH7
1Jg9aZMb/kRtavZWRGxsBtU7Or4fmMM60L4i4Hjgb/adurXoqP1WYU+zIRirfh3bs5Oo8YA0UY8m
768iCvfiZ+ZnP6K0X4WrZlrGpqtQpOnKBZvDyOjk7HtcuKxZXnRm18C8Y2H69Fcjzgr3mIqCjjAS
SRb0pFVlsrUa/IZKbmLYBkM6qqm4arc/CS2XsX3R5GEXHqxFNK8vl1qMBz+lPiCz5SJQxTj3ui1U
e8WfsG3ux7IY5Sx0sNsqrEmwDAdMwaxlyl8/ot1AfskQldeYVoSFSIvzuQtbpuFLjHJQ/1OTGxQb
5ekcizsAfgbAoeA7LSqHKNNeihq9b38ASpVHUxGkUU8c/1zuIrKRI+tNQMHFO9nsQGOKjqb4uCIa
Zpp4SncwxP9j5H0YtRtKdNkjSHWA+Gmrnap3BWH0wKf6DSQO+JESPwOCZZNNwD9LoraMEGDMgLgO
kvK2C/R+oeupn+Mn4abdNz9JeDkZtpmG87jx/kDxbRDh28HeTTFLmDZ5ygBNMa2G8AcUKa/Hv1ad
ExbbyIvzLUr174jjYU4gWnLzDA6kj4mnyBbZivBBIHEWNSC+gjNFspmETO0hf6DqNwg2ZQsxQFuR
P+h1D8hdGc9nLyZAgWA/Sw1ct3yxRwsp3rLff7e0P5Fhcsy8kDpKoLKTR+FGfiMHSFYs5mbdfn9T
q9MzO382bdc+Ak86GnL+HMiX7LxkwFgtnbZa8mYCxHqPmdgEzGfddKws6zUC2pF9SQEjGg57sLh7
mEd7I4i07QE7rfqPBOiX39zbmaBuXwstt09oiqUkDBjbk8yE+z5ZCSw797Up+3HHiXouqI4284+R
GjWOa3dNpVjtOzNrCCKRDZzHIHtegNw9NQoqvuIX/55iqidLP7RRynULcQKezh+7y0AdOkz20ENJ
tcTc07jRhBkB6Lexte4N0eZa2BXOIZWvef5MeKEXLHNlGfOJzdvSn04Sy+Viaezajto8gTyUjZ0Q
IiKmNemY4bAsU3CQRTo3Nh7g/7Gu7cmj09gbnBbQWXs0wJpqF2GOhZkGkIfy2C81Vb0TnlnUAXPD
OoBY2P19uyl44fnmJIX2XhKlJBb1k7VikDvYAnUn3XCu3ANxoFZjnEITjTL0nv4SHoSRcIU5+MA3
hwjsGw9hPQvl3oHq/0U28oiDhLqaodKtyyx+Nx3hQvN6nJdoXIujVbz2uoq8TkxSWlqGIpDxBI1J
ZeNVtTo/RpQgl6Ffi6HYzKoTVwgQivSOI+l5OSZIGBlEzD8h5V1qDNP03xeU8Kx0QWpE1wvQ8HU2
0vRBCPwsDNzBlnEDV46/iHVm++A4Yj8HOEczx5/xuZaECN14dqaMDc4vfNFw6webO9XetIPzX1tP
l9p2feXT0jiwV8pk6PWkawCC21ttQjsOtcgxQuPPdRMCJRuNxumpDoqrkw8wcylN2ZdewDu5/g06
CsfFGP3wo2E3QLN4rsexcuzfdb0Z+yZv7styKDJJ/pwRq1wSLQdhcUTPnrdNJqPIpmOkt1gLELfH
DFauSofNG2x7czcCZimUxqAfUU6A8DqImjZoG2Yoc2PrN45lHXdrhYf4rd5qw0DbHT8Pw2wV/iLF
Q+cknOWvTPYtdIkQWbAkVDzhMrzYjKnozndzvXjGcFhLGxUxJoeN1otnaF0bttqx3tYmlXth+z0a
vT4u2rLEPOpMR5E+wPt69jVTf08mG8eGTSMB9BkpsJVr9kuCtDsu8aW8TRgDKAQGceE7fHKPZks1
CZAR1o2oUQ8rM+VzOJXdnw9VZ9asQ6Sre5BEqkuHJJrgWr+AqEmSNu9O5wBSa4b/+Zo2C/E7CFZM
hOOY098v3azbms7AMg23PpzYkc7GoVPXBQaYmvQkqhGvsL50kSO57Aq7JtgYpAXi6oDESbaqTWqE
c52qU98kLJFZelgBxQZuF/Agk6NWUnWctK88hrXxy2BhOQ+JhLem62xup/0uRBbThFUqRgPsbecF
No+ShKH11o6q1pI/ibK+5LIBlJ+h0Z95k0uK0eE/WbwXcoPXn3g7sXl0prAJcpWd89y+cdB8QKGM
yFXSwIsL9FdsVXV12T3bJ1pQ96La13N3ClCHjL2kfd24UhqbFR41igny+GR9tewpoYThietpyT3l
DEH0bGvlINGO53gtFsIbhfPb+7pAS8DK/Eat3HCK2u0TPYWq5WOtAXw1m2+6PGhi9Mpb3SjbNUzn
4+ob087K0iBolAyZcmCRZYj2Cd+c9UVUENFOIISjCJTB6Qc/isVY+8Wl++qHPEt2IX7gfNje65g4
3G68nMjTi15zJ3hcwTcQoCg7OivEZQjKEIiY8mz2bcy0SY4ODZFs1XfPVepG6Qr2Caso0ucQWALB
dhaQDWwYAnJm3JD93k4NY5uk9CvNz5+MHFshc58MSKrTHgNso6q4A4SGn+gZNp6uqgGrFWzDcgAB
SDv1PMAQOHm+2Umrm4fUU1cdaPu7p/ii6uD4LNrkRLCbLLYGS91XAVwYPLh81VMdgnNHhLQqCgg/
yzfeR1vXR+KGtUbPOfF22b37oOAaOY/qvIM9g3W7AqxkL7pUWObO5IofeSMiRtrHcCcIifYNTI1J
D0Y60zweVYBPvDbeN3QafewpnOoaUUXJ2FC1HSTCdqWV3W2rnAUrkTdbtVcUwt9p51FOPsLRCm4g
1brKVo5OqcTjE41orTIQ28n6tTA8ZBTFrUKHWYsTTq7T6h1HJd3AJ9aN2FDN+QoQ6Tsfss8w2DUD
14CI5VoXKYks+FfkCrLt1kD9nh9PYZWM3bEgXcb44RVeNNZzhCQNBmKP1r4xTGb7jSRwVJkgV35T
wcy6GQnuh3afnN4mav2T7/rRAiTU7YxEQ9wp3sPS/iH4IHvE4sR/GKJMCi8xqykG8KmZQRu+un/W
KpcXTpXA1+kSNXKtpYms2e80Ghj7xgGkA1wXLq7Nv+6lcqm8JqwiNxVBjMZuv+D6PWvtieYGprFp
y8jitUdJgwyudEGywUCNEEc/MSXqqmded4LmGqxveHzUmHoAGltBgo5PWiNwMPWzvD8nM47cgxV9
QdpSPewao9rrM6rL6TUbuBGFeDKqJugosI6162nw3lEJFD8ZrQ57Bptw55FqDgH5jZ/WeF6J1rba
E6ND95s8V0TSzfDkkQ8GrNI6AooQkJYFzXae3OJv1PbmQgzSAZooduogEVwjlVPtI0b7arp5Tp1t
grV13H8dN43UIIBjWJDlPKxFe7eTJ2I1dRq/UTFNdGilNlHl2lLI8xTG0aLDLyfJ+tiHvzWMPndj
/BGQAhEMBCGqLR+eJ1vEIAKWShZvuB0dcGyNt+PTEmXD4CvcW2El1jWlQaXMDo31d5TJO9u4Ircc
jxD2LTrKZ58RRzPTcZhAwbEzw0VaZPYW/SlOt4PM+a59gocwMf4Gs27P4eEDuO1RwkmeMBzadJAg
P0NWsyAQt8OFjeDMH06bmsRuhaGIAhyeWI30yRdjZCX3OVIkPSDu2LD4N1ZmwQRSd7oCWcvoBlHy
6FXGyWORw7jiVcHzKzhdkATyfixWwzKW+AJgWOtL5agltiC0AmLDH0+X6h27UhezJHMQTKbAnWM7
brd9eleYTLZU5H4XQ9y/HSaVuEfrG8IXnQSBK5NaxXnbjcgSYBmnE83EPqfUb8WcMzBlYbpy2jLW
lW6jRDeZIm1FEa/FMMNlXyqwnGaoV/r7EA/f0Cz/kVwkjg0wPWOs0LXrPQjswArCvJtasI5qzTa1
vGFPYgKYrn32jutX1rkIAfZRFU7dOKI7CPeUzp9ZsSAFLj6C9FCcQVrbLQwop4LxTULic/k0jcnV
KJ0PBsxHBjOA19bdtjW78YtQIlJf45n/+vbUwAQzcr6eA8U/pxX0sb3Jo/aBSRgFueOl14fLFSc8
8hs5ZVF6Xbx60zmkrxcSBq/aw/ZVfdgormbqvoXEApOOoEnAkJgEgguZtQPmcnz5nZ4hVpBHtIYz
TTPIcZsRX/APguq79CTUQ7zL9apxx7uMuO3rhf59FZ4Mq4BCYHYmoisIAMr95b0vNPljjq9Rj3RC
mx4o+KWq1isdgrGVEen15eDFDHg4YkYTod6tnLHMf6TyamBBJAFp/PqItKrxBE+S5v5BvrbvuMW4
to4mZfxFBlOl+M/xI/f5mWSyxo38rhZKlScwcrJk6m4kg6FtPVvVIFDjj7oaSbJFY7hBefv9h+pC
bCLDs8WpTYwZEJZjWEz0oSz1dfbLjaAMhoa39SNUvaBqtyzjS9jsHx9IegoE2yJgW44g/uN0xtGm
gguggu98Okx88a5USOs7AJz5h6GO2BCoLY1SK8OaMExTwMaARJTto/tLqWTReqsxeFdH19xWd6bR
W+DeOH/D8y8vFcgiX4X+uAU1wbJoT8knEF0wyC0hpdgeeb3/+/JvViXBPLY0bwBI32NXTvel4HCj
gV+5DbVbUcg1hNy69rHNBzSfbUMXWVjq/vJE6Tif6uIEo6TMFOyD4LFZbe9CP4AVjgviqCjHnj6s
Z0Uihu1xnEvsvcJyVsztReQyA3K6r8Y+LpBsesODS9YU3bRZHT8hyj5Ew4tdTVPJUmrJa7XVF5Jn
xNnhxe/TpFt9kXkZrTgTomCW03WlJi9a7zThZMeCGAoxollQ0T8gASZ6fImofoot6BFXexXYuctS
Go83rq4fHNY2WexDUGMolmXyGMPCc9rt2ncij/+WaQhAhA4+cKakY2zRabVcQC/MZ5E4tGm4GT+u
iZa2aQ6b7kp/TMr7hT6AR+yVNmYuNJvSlguMnGQ3JYA7YN6NwQ9HqQmke0EPVgO/iIayn99ZeMy8
M5PMet18qYLuL76SbL2HQWaGyhUYlpb+U2iQCh2rZkNnVD14tVcNfOD8QZFkvM+1inQCaZa20hDL
Q8ohzNtfDXw5LflWAyNtre0p4SRD9GiMnNkUhLlX+qDo+Z/Im7Tybs6tnro9K25xF1wg2v3854WL
PbE/r5a3pvvm2h8C5TAY0UbwbEiOMEwwRfJNyAEJcMhhnluvhh9E57EMekEw6J4d9vXYwTXcvUhZ
OVLq2f+nLuvWfwJmX8Wqv4CEiwauK+cfmf+v1zMjyyErq7UjaGDiNvtkf3TvkqS2cRVpaXExpny2
apAtAUPpNbWY3hcdYOeXPYOpaEDFo+gA1yxO2eLl/gecnkvXez8CNZy9DvUXotxCqSlEmUc4ICMS
+3XjmwR9UCWfjMuxQ/yBJNbsreDDx9ZUePg2tFL7OGTHGkzYI34lTNUiCPpsRsRkJ0jDdLANMo9r
UZCfGh0LqXRLXKQjfNo/DQ7WM9stv6JjRLtIIIURjVC0qe/9+uSYI1lk7wkcqWiMOE3CI+UxWRs3
NnPc4s14/uv+bvBEXorr0Ck8VAdfYFdpuEYkeJ+vAFQcSXVNOWAInIxI9KQxIqUoFcT9eqNsNHaJ
v4FKEdrFqMeU1urZzfnOdT2g/qnUd9w9PnOrMBwQNeWy0NH6NjaWVljPSjeSdHTX1oqF4dBe9Fae
BZ4oCcALrHZfnNLnH9EYhCvNSb7XoA7l6tMqf4btDTClaBnNf/C6ivz/hpz0r9LeuHuPxHmi1KDW
OLGvSdEL//iRbNp+f1jm1+smVYNy5v2KAuMzD+90Ik538NhLJTluf1vd4zwnBHpF/HE0tcV0I+BF
aUDZEaEKsM3PbytjKz8jvtcSQri74/9BRQ+gPWOINn8/EifiqX2aeCtj7JJQ6V/+jGZ1DYp2n+XJ
u+nGFgwbEhjdmr6rxKM0cO8dsp/XGnsOWBgmcGidYPAtKDvRsPXsuiJO5mwVWrmdfl2sfQ3kuNwA
ad5KzfOkO/3mb0LBWK8rQxa5HAoovCb7Sw41ob1VQ50c76qiByfeWY/dTvYwtB1yO7d2ZCrIZpQS
9dzO9mtCIOKGeE0buWepIxoEdV6Eh+ySS63nN6QaFm2M9QQHfxyFISzhwd5JfcRj3w0jM0Mxwo5I
4ANYUS9VvQrz/Wah75+zMsY6vu9bXy6913S1+yDQ+/DPk/fiNxmm+TvRaP1kkv1C0tRqt33R9KAr
SRwuHsgsK4nUNUWa+cwX/t2eGsYWCuFtXoZvuVGg5Ib31Q7M7MQX4ygYztgA7elOL3dAVBuwW6PE
aJMQHvJ5gCJyamzStD2ZxQEeA8q3ZuB+5yum9LL0fxI2g5aKilIFW0xwmrDnHn8jzzujoSZnUGc1
IuowUgM8N7a26Sobxj0NSkTzsFaquk9LXX9vmdMgfxDZDAPuiSYIVkbr9xenMX7HrYeR3krc3dbU
7d5BoC2pDInDxJutvpAuQEqABrAf+MZ8VmsyUKtMKkcxJbOEQaWcEsU2rzjEginnBMaHvVJ62ly6
GSe5y0O4jKh1bbTTg+Iif6qJvlQ0PZV2bTF5d01JIvvFmvuAngxrEkOfQnLFt66VPTMVWweewNcG
bU6wNkbAegkfljRs/CdbjGOwsyAWxdin+vGssmym8GGIou9sLOst7BCASTxtJpIma8wvoXyfJGLV
9EMdTBc00kPKzSuvxCAuhmE4AvsuQuwWP76Rnjk26fURJitgEFEBwOJM0IUvgOnFqSr3JxkUKQOE
K8JYz2DnNFgfBQBEM8sT5mMYHS1H8xb4PCW+JhNzg982Aovzv1hxnxwu4F0epXFw+lEzhBGq8t1F
W4AY8z/FGtwtZX1+me/nQS1oyxtz5FuT8yybQeb3kMOOOmRM3CySWrY5MjdX1B9APQMxAMjCt5Z3
TAq4glUmfMhnP2tfknQk5JGB76CK49QNXwDETQCxgJ7fixyJV1P/o+FE7DL5hvQr/PhEPY9Jzbal
DHR0iDI9l8KmHIvEuPXXworz0cuW0OMqTv/zgoIx7EEhjQ4Gp/RfmwAIcX3q9s7HTXWrV0inPcF/
wpdXmrH4O5xc3IgSmsmf6ynw4XkDd9o5W5GncKUTR1gtYzSc9sTcBdr8AOSYCOVanPMbdXHvCffK
I4xEJFtk8iP1rDNXbrJXddFXqlnDAyE/LVgs26rrKOX3F8hF8UWk05WTHFJoxr8PtHbxN3+KQXo4
QenGeUY2VaYBj1Fl6M9Z3aa7d/rOFbiViqqz68WfrSOCUozF3FrGEtSmnsLD6sOMWRma6lKWBQ7w
T/SzldOmTSlsiVfJYM49NYVunTSC5nQI1qa3faPWY8tFhqIR9MOMBygEGyXNE3BtbaaAFHXCyE9C
WqieMxlKfsJRUIPEmuD5rh1kKgK6S8tAcjpDZZVLr6SDKPw7ecI5UGCv31QNkNpVDNukSY2QRI98
E5ZykVb2/F+1S9SFBTcbYO+X1FBPlUpx9xhN1kHaLz651mCLn5f5DFjwAhRzZkmFwLFGZ9wec4gR
Dpbm9aijdEF7emY6FdG71VInLXUMw8zYKstfnMu7iv8vtOFJ1sXNT3mLoomRm99t1mcpGWa3dT0c
mV4g9ombUOaPsJrD9i9yb0os1p80SDT+0hQ90F+H9h48QgtG9iJYTYaGfXchcaAxIY6wCjsR4uE2
sewAVGbt30/UK/Kljml5y4DQ8z68/1kC5zCtKhVSoYtIGWr0QxWK9En8zI10xM0UxA31ngUnA0/q
VPZ3iB+AjEiVGoeSk91v6C+se229NsKIkwTMPvvPOPM5c7LS/OJCdORBO2e4qxaBAx8VOMmP4iUc
kdFkIgl8MBtO/lVdXNCxHZLYTya95Fgd7b5PnrsIRuPBfubdiS62seVOPW/B6ih3waS7CJ7i7Vdg
q7E7LB9jzzJU6aJVk7/EVl3Evm6WQU9P2pk5E3EXUTgcg4YXyP61z4jAHz2lnNUs5azIGssRve5C
tYXNFnWwgRuyDlgK3RzrDcg7V9PO9O0oGhLiGPrl8kYifijJQ4IxhnRGBz/atzWmF1eic2d6AT5P
Jz6H51L3bNRSbq+0soYm9fH0frB03byNaKYFaFzeTv3zfqPN1/gbM9Is6TRPJHIUn5MbxTr6dAxI
Ge9VVw9vrroqEx1FKR5YO4x+HJihE+SwJOhrCXoyIb0zq0KNWB8dvVZD09SHOcT1DoYXqaD9BRWq
95NY9hNGCpiBen71mNCLAnAle/W9DJVNzzWn+CdIwdtAlFHM/r6Nw06Jj14oNwcx0uerqyNFLp8R
79/QSSjlwFvt1lPuk3GGp0kS7BLPHtdgIwL0OSa9T1qmzIUn8ErPVqBbIBUo67Vu3tsviRh7/kVr
lxvWSRmBHaB4VQHOMBbzAJLZSkDNsjYUVZvmNtrDfcqucRcsvDgs8WgWidVHLShJDclag1P3IMey
8bQKyhAS76QTMIVvI4o6Ccie1zt/Wrce/3L1ms6/Rz5AHf0zHJF1mdS7pgzBcuT5aCADyNfEV3yV
VYvo/YwSOJIvNH1VbzM/AhOLfD/5ZJPEh57KNSTOaPuXD4RLTgqq7Gx5XQY0mbWmP8uGZeiA2sBL
EUTlMkl9TO6UkWiUiugTxLyo+tEah5imnkIcTX29k0bNO+x68lRCXui3ZvfSDsz5QG4571TQEUCK
wUvCrTHxi3lWx5YgCWZFYtSENs7V5EqT62Bc3EIz0uV1o1jTjjocNaWewIxHnvFK3mI2ZIPYg8iK
fI7177yucfesEzaFINBWvzIejY6+QXCXU+9fcIfIwJXfkq2zNyY3elR90Ix8uZA+67nEU8d1KZLV
Z4kpfZJOVCVyVC/EwKbmdZElW91i1cGlz/mM9DJg6GPnddU/SFduRaEAjus5HgEmoLZQr03D23eT
pGtbxNfjeprCAw51DfbzoXbhb5kk9H4ePQsqX1B8+5owzRkodSruzDuVdzrBcBANOaRvsX9UvKIY
UH7noh6V1X4YGFLwO0GPimBtfdCKOeM7LDzwENUjkwJ/49vj0hAyX8Iamu3PmTQCdG7EelBPjEZT
xxCNZWTPjG/Qz2bP978krC2zq5FRQ3qX9v86nGH8EKc5841hTeImM6MlMujQuElIU9Qlj3jqF/pD
BgAH1vRVQLkMLDTEym/fF/vQyNLUqnMuNzgTbBOgescD9VbwdjXT17BIDn1C3oE4DSORvujGa3XH
u2LZFYD9kCw8DDBbfJZiTh95KawkGhIBNnF8qw9LStk+VXHqJBYX7QgUyb6Ml9Av9e6Er27PiSkH
ecYRr/KRoj2ACMOfk8IrlrSDGvpGCvWYAc2GhKmFpZ5IF4ymKmrQYdmVq7eHTVs+rduelgCK5lRn
AzEYCwraPvNdDyQaLyC6J372f7PhCkh9RpBbffVlyUz8aC0oWX8oqVpv6eL9L5E7bY8UCSKn0QQQ
2ii595cVgmYWAKZ7Le4fLSJ3ejo2gQtmvWq8q4yfLeKNtPkG2Z7lXT9itjt+3X5kzkvmHv4rkshI
6c557d2oFdL1xWEXYAeFo5m3mKPgy0x5v2HPJ3/WI+6eiQ066eurxtEKKK/imVW26j2kQfEXchML
7njBYp+Ej1/tDDeHoMobbhIV4u3aa02XD4w8icOKkLwVKO32wj21XXJk+9unIrlfMOJr+HDs/IRZ
dgEhQjbcJ+yA/Dd7KhuQlewZEj9sb/CdkrcTIzLTpGv/iQC/rEPaOPRBNB33b5C8nUi1irshr67L
UY4dnot2W1/Bz0N13KLDc5j2ZLqyTDSY6fItaMhrlzLbENDVgxq2OV9qG7K95AHAmcwR5PNyhEIj
Lio2AXL7AbJcRf1cuKugtXH2jTR15SCFfbdLtUrQpsOI3prMGwGRdDFZo3iPTmPZ5fc8RkcaUzq5
D1Epp3y6kdLxg+zQy0sABD5agrFoOwo07+ERrc0n3t1a7+v199GHJuaOjmXZ+rOotVq2GGYlMY73
/NHrhYqIteCw7lHSY+t4M607asdf7h77p+jbVXYdZ9+4lxHwf9pBTBasTed4Q4w8JhfBouOROKH9
ui9BeJfgaDGfVevroOKevIgcMsuFhmd0Xryx9b3Ga6q14gM8f/3AXD9PFffyov4nlK7A7k9yN6MN
R6iTvpIhDr5OLF75W7RaOsGZgN2QzqANsf0hhr6St7XObV9FaS1VvbjEnH6wrd2kOfK8Kj5pDTbv
cYgitcEh4PSoNURt7INafhX/z+LGzbsshO5zhLnArwS48Z7oIDwyjVp/yNMtFad1SpzRybZFk1sG
Bbubqc3+P7Brmr2DvA9K64o5tOVNyuQCCA0lqQTFwXCHPGW1ZGbJa/dxhD1Tahf7TxsqbKfDPbHz
pksBQ73q0mjGM3p53xW+3lIIdhSXxkEH8wTWUMYj43L/BCeyyHYF69DYyyI5OMVsnl+ZPGMZRc1l
bs71R4dmwo5B5Y1K1XwQq7zePRgYY7FoZn5p2BVogXNXxx/EBWGjyP49mfr6kSCMBnS0ZYJ3DyGc
EkCBeYOdYKOEvs+QSEMRCVyt6x7Hk7QnDoaLapKRL6pI9HCa62PEFWzcWhRPbn6rdvytIcYoHztP
M2SDn/uQhlbG22IofOWlCH5Hn5yH+R+WRoAPJWt1hNdhJA8L2EewfyxWOuvTEy+yYsXRgnXldxfg
l73BHhLrSrLeyoJinNaarx4gAhJ9PpkUjAKxQy/VPfPVpfzo4qgQlcm0bpmdqjNigZrMCaWU7yUX
LDeD7EZ33vh/R6GiUqSB+j8NYG2I50Vc/gPhPImR3nnkUbPcF08mCdhDyCHdLwktqZEuc6enxOzc
reGiZ/AyV2TtZTosaoL5aB7uTqOImFo6wJ2MLaEdGlmBMPmyNlzu1GOcwUs4mh9Tz+NGvhNZw5mI
im7yF4/k/Aqq1p1+XjOPhM4WW8thV/tkWCEfWyPdI6GpxyZ9eQMG1BUFYFYbcx1VowTt5FrsojJh
8XWTAJnx5aLlO/Qov7yiqL5va7umHGn+kZeDhNq9JWnfsJcOgqHaPDL4t9WAFKvLrfGm56ZZZAXu
RKshmCSGALU9HRMwRR5ByXioNu794ift6C0AITf4CwqLdNE4glKMKGCYGbdLkykMxqs8oJQjA3/Y
VzAD3ao8jxo4AucpPWgfLsPMCmaYZbenvjktMKqgNfhIPzD0TOHFKSQrRW8kn70AKoA3oVP/aaZ8
eG8V8pPLo7zkwhCguRDrwsWt7QMRCK8C05UZQ0UwJQ1TSNRaWQ6JBow8CfdHLI7FDGfOdCitVNDE
n1veH4c2Y4iq1gQWQ8/Sol/e4fr/Gh6RJheolADXvuLhgzsQRr5wCs2lU0bbvec6PTLWB97YUAVD
PqLemo7FWxzzZyXaEKxOcDWCHTkD9OQodZ6tSfkBv0UdPTyK6BfNkLfhY48mIwqPvQcYJqqQ0xI9
SL2YVI1W41QP5OsXxH3Yb0fyltHChQp47S87x6mQlXQnh26PWEfHuiCBWE8Z9K8q8jLFrGYAQFfH
Pqo0HSo2QwcP9p1p9uOBT8NgXc2XMqH56E/MGdHBvNQPgCPTf2L6NtpPi3eIF20f7KHBbuZ4tgkA
Vj5LmZbSFjIyOEZp7FoHbzjp/UVD0wGAxQXwIhHmXXvbj4Lop2S21MN0Q6oG5K/MV1VJLT84hsyp
+vFqohZo9FOsAft9o+69wcwf9srCz5ML1holuKN+nwgqu8ceXOWnHe9H5dQmOI3LjCY565go1l1J
KFUmOGaHTWgE4SwBejz0Rt5DWnYvBXStcFVLLPEtVuBt3OXs9p8OiH2ahPBRm2828PItYhgikEc3
HAJ+soe2rIHkHhRSGk9XrmnX6nin4HzmtpeUG8CLe36NQGziEGWa4ThfP2yjasim4VwOqoitj+3k
axMlD1Nz/J8Z6IpiNJiYlku660Iq9KmSPavsDvAJ1tEoxKbrtT8C0aGhkla3bSuYAN1Sg7HwmvUP
ZJV9YJ6mdrodoL2DQTPX0EreBAEvIzKcwUGNOklXorf9II9Qjzlx5lyQC6ttveCWSFhLemQtCTLs
Wq02WdopgVcV1dr3t5kJtOMLrTi2s2UG4Bt0KMNm42X67cp0Nw1ehw3V/weWDvkt7Eo9juak8ORu
zeXEFZ6goYTfq9M8YMBBQPzUELaYMgtlu0eANO5hxdszCsN14/7KzP8L2X8b8SDA++Wj6IUrnnZY
N7TyKm1/0pYHYkVpwXk3FBg/tVZyXmlhKKabqEpsTzxi5KssBLaAna4s1xsP+tqTqqGeELu/OpW3
fgoXMCr32lqBtwd8BuMDbaPlAiBKnuSAsXaoQMZx+82eU0HfzAty8mDJkA/8h1M9cYVM9QPMt+PP
fm9JWpxCpEK0gusFQGZ3212TF7eNFNIIbxsvuXyMbvElFt3/+3N1q6i+9UwJd/Z0FAUZNIo+TAJk
x5TuNQDaG5GFG5H/MBrWyQO7VRR2vjWfg7alCgExAWVwupgHnfMfRT/M80KVUuZHIuQ/VeLTxr9J
kdri9T1swFKmBgMlzsVQpAzOptDKlvzoE/N6XpwQsI9aDB92jmzJo0UQCrPqleYVYVcBN0EgrFdB
EgZ63On4bZXcREH95RtaYsw26jLqD10tlcKIptXgUUEZ0EXYiMD2WhP9O7U/yODFMbkR+IOK3MFg
BGCUTPN215u1S8KSo47dMcxHtVuXKqc9dtg04gf6G3fn1XUcmUw/t/ZJNhAaxWiCf2kVvpQXVPwk
q28SNmUjqQ7T23pfdpZST3EpnhjAGR5T7/nYrqHM5f06UviQUO0JrFVODWmBw5KA6euq4u6scH5R
ssUGJ/2TaiIP3ZwX5N3/Bn1f+88XECHuVmnDMWMClHk8M/Kkr6PZ5j4UwJ6S/zJpH+eqf2wK8Ev7
mGC7Zg3AJc7X/jYdphS+SYErAsivQfLewJOxVFolQK9syR/Qct8fWuq/oPqYRKM2jokvZqWALfjK
fOaBTgVWOX+faqbR+64s42vkPArPj6IQsq9ch3LIb/3YfjyeU768Orv6NxiiLzwSAgaDu2rHU4pY
seoYJBvEO5rLb1XWC81sNNsNIT0rE8nigt9TyvaXKFwwmi/AD7WH49wH+TJfyMUU5ei+y5CD7lsD
fGH73ekx0jdXLtl4n1CdSKAtZrNfg+FSvWab69rI3MXeq0E/LN29ODDoXnjhLZF3R5XIHn4SmbIh
T/tJ4z9l4Tab8zHklUyq6hRv8miotHqclmbZ4zVuQ4qtRPv/3N4jH+yxcIgnzqSQ5FjbgKFDGtx3
fraohQLzFQsdJifcn3XqlCdiSYO3cbx9cAlPC0Bi0pBiHXK6f35i/hKpqZF8qHgN0i8svsZDy6NU
n3V4hIsi85rcZkskLHcvmbXhzD1FpamD4QX+7KP6J0up/Zt3HNE+fHe72MEBsy7SQzTeIITrRKPo
0P+m/b6lfr79uqMhHuijEP5oKLLQtH6KSdaVxHvQc22dCIljdY8+fWj9Dz6ItoAe239ekzVC7QQc
qQIrQcgzc9wJRkGUa+XG2qEKMdIv+DbGzzZWGlDW/Iv4i/xYo3hWfjj5zJKDeH2dbH+XagdqLtao
EhM4VdKrXj0epKWzsk3apw1ZOGhWnWbrxiuYjzcfGxwe9VGwpVO2a2Jy0exdvs00VXfkqlRMOfu4
xfwUSJKMOt9+B0rqDoJ27mln+KxWrbQlJ1JhDmDBJuteT+ptaUxytTMVOTzN3ChyUBJfnZ5Hb+0R
njNiWmbvMIBHfRloa/ocBDrptoxlHS31t+v/CSioG1XmssetH5+il+deZOJNubwVsHBZ0+H3FW+7
nK32Xaib0CkTGYZvfPoe5EVtqISRIeoyGt+vO1hX7GMHgxVJhCYNKqQ1KvlV6cS4o2qa6xUANJN2
I/r+QY7leT5N02qsUqlGAXcm0BgQ4dgqAgFVy6LgnXu22ils+oEsQS74jc6pwlzGm6DpGTgP7cqw
JLtYXYg+AZo/6GdtGBt69/9HOHOqMevMthgXFiGfluJ3DnjLZ7/nriR15SV/lxnteZLVCG0NmV6e
Pq7QTByLg2pKtlccmt2tz2I45vDaGUID/zWSi4JfRH57yc+0taleNI5l5/RCecfYGh3+0POaASIC
2L/n1QYM5GRm2gvZz3v1Mpjey7eAbGJLbwQGc2U4WufYVsLrRE9MJgQyTutD/9BLbmYIEs2f5YoB
9SZdOAZ5hmL93KEfsBdhqWdRs5cLnHRb3OUgtfqmfh30HVvmGdTRAly5OqnO8dGEvOxR1v6PpaXc
NYNCICE5m8SvKeoOo3H1xCeU/o0GiNl7sdgZb+qrIbmUORXGNt1Np5h1KrT4TW+MAJmFS2Vi8Uf7
PEklxUN9kZiXLh4TeFQQUyW2y8eRzw/DsiH5wqs4DMmftJrOrFXFLXYqFVcvG371WQKnsgHUJkce
+40TkgUwFZIax619Vs8YilGiYvE/jhxPCBIP4dSwTm3i/Z0QWFThtzcavgIUDGOTIGJP9tu2UwMi
NlVfpVePrmGaad7us0n5iEw4SwbZtI6NUlC7Rx8koS+2OKCrQBuBlSgZfb/0v4rNuaS4c41q8bJf
I0qcv23z+/PjHYqMcrbTv57d/pODw8efFzNPAIZpSiIK6EbViDBvQllfR9zwCBetw1tQmcMDFYnG
HI754bLKRCtBZ6JvFncfhXvs254fSvbY+j7a6u8FtPi4VOrbJcK/4r4tJncnzxmUAhH6P0JEcN3r
ZwSosfEysc9mtKDX3WOgqXoEPAlg0mnpJXugfwSDveUgPPBw+eacCA5denWH0c+aKFkb91d3wobI
FGpX/d1b+aBSKHprpKAwX64t5yzz9ZJv0u6xj5yGiCt4Gm7Sh9IdwhCUR5Whm4qIzR2PV1X3ieD1
CjPFuQGHp/XiIIwtjKQ73owru4iYefNJKO/VjdyK8xAvZ+Lt2og95wb9nwiSQi/OpyavGLw3wW+D
IYZ+GgsQVNkVH+GUjAhC9Udhyfn4vVGMW1/J0qnbrRopJXkRm/bHe3kKSM+eztfvluCVDhENMALm
62V7/Kuifx3MDIg/8qMoSLAtwlYKDNz9zd2gE9EjaUQSyfZTCJDH2FwWNCHkbPSXaZ/AIoaLDrgx
nGpWygdv3aoNLvhrsSCLm6raW4n3/zUtcUrSHYawy5wcMuaSLggGBBf+Ue5o7+jcXes15A0bkgx7
C1yCMLbFU7la5XXylup/q9SDPP7e++GB53GOqBoHFH2jSNN0qgQ96rjuCQWI3Fh2+qBAuNqoPnMU
mm2ImiXwL98txAwys13ZFYocv6yAg9+1US9rUetLQkfBLk++FFW3STohzQ8w3Ap13Dn5Wotu8/LU
Pjk0dPWUxW8SQSwwCAUDtPkwq/V+W6p3EIbbamKpYLRickeJQMLkg7IeeTeUBrU3hypDlzVJq2qe
bBxqY3u2L8hR0L5WoKNn0us1wNT9FrLgs6OpmBsnadoy/R8FtRGGbcszQT/ZpCWeqjhZ/1sxz82M
nC7z3xmoU9IbEuXhLChd5yelq4AWe+aRbo3OIPsaXBOQW7BjYP4M9nXwh0WFcj+dstsDyg4zM5PX
EN8SUaD+obP+nUl4VDesFMi7f95Z/Q7kjs7/D86Oyo7TkpI5qtZ1gdQ+KorioAn5TEwYDnshiV+r
QWTaqwthUQOAa2lGmhcKK77f6oxjYNApuDzNRyU6Tc5tdT6iIUNs8hoL837+DilvxDuLravSegwr
DjNtvP4/AMa/BFna3kqaBCqxUinh/QK1E3Nq0PiL6YxLQAQSUNVwTYz0Z4yRANezybOxZ2teKV6X
kQHqC/TKfatQ2Dq4XJQZFknrlmSSjcY83mUZVi80P1+6nIpM63rxHlq9VYD4lN/qFiLDev1Zvg8x
3s9yratsD3KPZqK9YHOnkCh7Xe2T89dtZ5hVHh3hBPCWKkjb/uOBpUb6z4K6PcHIoWRF2Lv5Zxkq
RBK3+WoZY7daZFD5sol0e11lharsY5QKCTBnHTSMqzDqzboHoz7MjQ7HKfsLCcMc16MCj2ReH4x4
saWZME/zDBNlRNBdHGdnfirF+kiOFOhgJz2DBEOTpS3Ce/xCXnb1Vivt/zIA8sZu+ZVaSNMFHrcn
if2LKtAXglnQKZewsFD9Z+fFouo1FHpoi1z9F6OKJ39ZXO/liIw5sbvDUDasfgDz71WQQ2z12ihl
xGzJjeoQIQ86N/CPYS1heM0z/jNXLfXjZLSvR5oIg90Dkey9HtHdmE3Sa/LzgPVu/CqSdxLdNkBR
GNt3Og6Occp2iWg25M2anTGSboqsi4MHL4q9NHf902wCyH1xQc23NrXu7etsjIm0FAfxiXE5hjfk
32LZOzAVJ4Q4s8c7L5rfdxR+okCiaMrNvox5cm4w/qmFcdVUzQrT/rpqjaWmwTeRz8JpbJH1CO1g
EyQuBO/10q/3jE31HdbbZHQ7AdDC56IWHLO74kKy+VzM3bsCXc1EBhUunQGkPnnqo1CujhASBGcQ
N5OoE/VVCNFJt1IrdY40mZZvFYwcUG7DsodCEo2XMhWSYdFoUn78p+7tAutRJYGgyXco7UqWC4+6
eEFI8kWqOoQmW95PN6SGY2gG/yRvewlsgw7/sF9DU3WK76qiwYK4g+d4iCyj3jjulYLX6nV2fGi/
WFmz3lPXWfBgo+kCjzk8C2yjanhmn89gB6EWmT7DqGSR6oZv4YkymyByIL4CADro3KxZ0twQJcLD
wvxGJHz79tG4DkrWmfw6GClqbEDrKAvy1pHMlmqkGFdwosiVLNtAEabmenI/LF/IrQv26a309gkQ
jeRIvfseaCFs7fT9rBYgyK6FVXnZmRhD/lTSOtCW2rRFFlVYWGDyA3EzGtUubWi4EZyin9dWKkEp
jHSttpXLDrupw7boWBwp2nlNt+JansDFFaopW92RsLKS4aOo+EFTSf+FpdxRlX7dIe1eoK+/qRO3
dDBLaxeADhHbcep3ihoHwDHddZKtppJBluRsHQrv5L4vhTJYQjWiPXlOtpCxn0JiQeXcMxO0DVTH
bJwUh76Wj/zDyS4BWTpM+yUSlP7s0JRw1LdHUj2Pdu4B/BO5HtniPRwRSbwhrJp4ThjH6dLfDRY1
0Qa0ZWzDcblpteULUWH0RnwbdJv5xlyRZc5YFeuXjHo3mNmm0o7+IrsEVCYe9qmVhAHSKlobEihw
4qeENM0SYw5d2+CeYeZWsrhAxLoWElw9+aC1X0fcCq3paNkkL0nDTqHcG8dQOrFxPN8GFNV3GO6X
Sx7U8L8MKhWi+1WRPX/pk1mH51qrsRrwQ1cQsoOAfkLHPEh3dlRbKtaWcR0rTV5Up/T17uTR6LHP
BY0ekm2iH6JzEHtbw6vEPutTp0qWFowV5sFkr60g6QGLRvMLPRenwQEW2tKG+0g+Du4gIc39VWsC
9I/9nTjj+Dvmbm7+hDpJz4u4CTksEsqgbkF5QZS5oq3RFaD7KAhS3EJ6KSaF+CM8kVPq9lW1KtQa
+ilZ01GGq5im7C7m1WpFuusE4Al2KHLrAVmqVHhIESVtCYX9r4Rt00zZEIwmM5blK4J3ITtxJLqo
6mUFIqzJzbqx3rP6h4Q3c9SS7VxaMKNAo7HsiM3+yzh0Oa2jEkgsm2tLLqdFYcJrmh0vBnHgCRcq
CDXOZpLO6j8xLCg5xnS2Cunpt4vSA0FLdRjgKYwCRjbJO7WB298PXqq9pYJ+Z42jmED6guehuyPe
0tApu5pjuHpibTon8CTWvgARphl55o8TZ77fO2N09TGnkOM2grBwtjSUDvuTewTeOs342LUqckWF
t5ol40HzDSJjart9NJ6IcfJxvZukQFjpoWvgrIUtHo7mJrczP6kQ/DJuHSbA10akL9aVoI4ymMQc
kx08Ldedh/up6/BBbcahdkfn5pggqqPcOJDe9D5Xit59CCxXuvm9KrFraKdvwsoaR0ulDHws4cVD
rzGaC7DZGEEYIirnCfYsC4EYe7nal+brqGS+MXX+/n5r+DZnvfwUOF8A8b76TFghX9W5cyD9eCwY
KMhlrUFNn2w7xWPOXHnAmtdqB0TZKGjYTZlMju4bf/ILHp9LSHbRqPsbVsT3VbywciuC7kW77tKZ
pyhwj822FjwvAeOKOaRYXE/FbecPbZH38QSSBgEKRqbACcjA0OVyItbNKa21jMxHdDIewFyqZtlS
ohUhiSPUs9RySnDVFl7z1DI0jKkS7A4UAovJpabGCGGGSmHoSclHHZpa8bzdwgFRQH4MJ7svIshS
tTRsvgvm6Ti7js0HQJTTseZOhu2OYM7EPHt+aqFWNQTZSA3g3jRp9D2AHRVw3B+A3SybsvK3glyi
X1YijGEdh8JyvxsUnNvCta/oNZArhyxSTgBHacRXxV675YRO9iEo28CkTh6uxx29Y23dj7qTTgK1
GsbwlnMnmGWxr6I7Yy4uLGoD15Qe0khHRYiCaHb13HcH6K54vDTPasYznSYEw709n2OzuwFZ9Hdw
x3/swXEN3uF1rDC8GoSje1wgjIMb+uQscdaG5ylZ6kCwRXzFmm5GrwQUa24Djr9BZZrCGLqlByXS
13dh5OSX4MsS4hqjX6gCnMr039nocfK/y5xSU0zf0um6fT/VFg9LcdT3xOz6W9kEolYOvKlvgnec
RTKL7fD/YM458ibrHlqJUVG7t6iqC26DsXWxEaOO8XJDBsdUheil4i6bYrQZLftAzzHfMMDOjLQ1
Z+lwKQ3uGRmSIYnO24m9rBXAgceNviDaVyVgCHUtXgE1RUfoXKfkrA/OCkfT84kES3ovK3FT44Iv
nmbiHSIwRtoyQ5+vLJeshKV8JkEEPQ/aRzpSRXumC/dNBKfHV9uQwPQ0fMtRhWT9L6BdQFM/JdZ3
/cyCBeI+WwyptWcD8iFpeVh3Om1o8zn5qvjL3AoiyHmeBopDOtpoE6DAf8CWsO0Pa2t8s4dSBA4E
HC6OLz2AaboqKr3B9s3oVjOQVIfHJ+yrfw1RGMtUfy9d9As2a5ZsdzUFhrIDf9XqL1yY62vfUBzF
Uuy5s6kXPs8HmlhxLFvq50sRtXW5bPTMiZtDTNajZCrPfvnJ4il96l+LKWbJTcfEEUcBWAS7tUSU
0doGajq0QOxAUlQsuRHmxcZJZ/cAMFOzR3iZ0Wnw2HT1FmFUDr5tbr1i9b0a8GpyNo1re+GHnaD4
aZLXQjMd+svENetz+ehNyBls8KviT58ZR3OTbgoAiyXLQ9YvgqMmRe+K2FNsrtofLJWEnyMMSwJG
/2Hls//1WW90lRvHvNDN4FduICv5z5gOLajz0v98p2O1OmOBs+fCRcszGCzHDePYTqaf2acESrI8
bBZlIaLmJJJnIYbSgh/QfKxf4XoSfVBztX/xWo2/nVf22+JgxTKMf1Tnz2gmA03P+jNDsdHSfHIO
P/TNqGZYi997GdJe0kXw085G8IiPsgrBqZkdahNmvCPDreh7elE8bgvYV9X079hj29NeytbDM77e
W5Z/imKaumYG/oORP7angLiSvrOP3B90vYe2MbrDrduj9mHX+P1zf1Z5WxteQ30NkllqF7iy0pBG
befkgco05J8GCJ5/6pJL1pabTq9y+ok62IZ1TAde90h/K13EbOUbVcDm7Z3MBqyOjp9spvVFPQrB
tmS9P0jJsM9i3AXdIxQWwP2/6YeXqsdV1ifqldmOVD3t4KVVZIMsn+V+E7wHip/DGCRMOYGk2ygb
ZjaD80ZbyAMH26YnZI5irJRI03inPwDU5fe4VIgEm+HQ1OrJFQI3ZatsB60XV8ihvWi15wH1WipG
9jyKPxPpt9742PgoM56KjG83MzOxjRYcLqpZOL1WnJHRHX2X6anVuoOKQuW1pqiR4QnHmM7lqmNT
6KfgXqc541WQgucE3S82T0EZDI9zQh5P2D6Qr96tk9Gtk5AeH2CPC7FPLTizqr6/PVFYO42IIo+6
lYQgFuT/R+76DlOkvCX2qOZoVCJPB7C0C/UtrI9nroFZIRHmpqeSqEMuMne4KSjcrxgtsTIqKK6z
qzqmdxQrHCjsz4uQL8aEVRc3yCcz1FiP3RRqSoXIyz9rTPrRaD3uZWs6x06dLueKoppAmM2RUHuS
fn/6vvQieWivzdAy0aQ2+joEDHIxX6or20cd7FXCW9DeY7kUwDeuGflPvJbcn4nE5SOcr+I1DWDJ
tpERGtW6/jZIXPe1Q7S1DAKZdrLlxFpGyEjjbsz9+MTgit/ushjE/atMu9tolYqSHriqAFwrMT8F
bEmC6tKnauBhwurxeB9yj9Tqm0hjNBvTwYX7hOXXC9iKJxgcDgdjUvc+EH6wHwFydZu2xA7sfqFr
rZp23dMC3CjxavPzNazHPtQWMXC8dll0DIKiBHaOgqWImyShXrcAvvFv/nK6T8eU7hEVaCxuczR0
f2QAuazjqv1rUW99u6J1wu+kPwfTQgo2t3dswoyYIoWGUvdTNf1vzFycadsrPlWYWNvxV0CZ36Mp
BMS5hvx7fUghhQshP0eT1kFFzO/QySbhpz1yf11xLuCnCtbdCHlBFmK/bmidLOOKOvQNoaWL10yz
D2IK2oCBBFb4WQgOZuO1QxcDGG9ki0xmkWEuNdb5kVRjiblbygWX8tjRZYweD8qkE7PHpo6LNPgJ
MUA15g113ZbiKMBuE8U24/zXyPp1K2rsx3EKOBUFFWpiyh2apJD7DOGZiaS8yRUCndOkXja1rEYH
xFT0yzfXBqTq8sG+I+W3v7muK71cap71EPSC+WSbQwQSF5fVnpf26s0A2WwxfHFLkt/b4OiTZSir
F8Ac1/fE1+IDzOHaspu2y8rOXUXznv9TaRUqRgXq/yajN8wXQz1asXpZ1D8ZE3W2+609lDN+AZVm
tyvCcmIEwqn8SVE+4iW0SPe1JU5PA+rLiGgpziwG8QiP5A7GZ0egeUGUq263KThrYhYyisAZe1y0
+R4YJUemBJd9A3MKcZPd8YvYWAEtDPf7RjabM79NGO9dVs9pq4BxNW9f/ZsjYyVohOUo0x8dYKho
F9g3dxPCKtqRd91SXMg0+unNZWhJwGd49XoLPiMCfZZMdIbACMMytrainBtMIpJeD7LftPDySfb6
bRh1Yf2CsjuCLapU9aAXkEx9Q8WiXQDTevjygNyc7CmmdSB8eSkV+Ijm2NmGl1lUlN/5SagbbHPi
Mv1/teXzDj9CmNtFrYjwPn2VrhC25D10d/rGy0CDMQD8FB6wD4BIwfYiPNu21jRSV5wASE9hvwsY
9srZVk3WkiabsdAaqxbZktDft09f+kvvfFaTSBXX7CkydUxnIXyBLYv99zOtznUvZWvrDTHQF4e1
+vfpSiqj1j3Z/UY3XfJdeyyUDtDh3WpujhtdBKtiLxKseWq3Fitlf7hKK2WFq8by1+RkDoL71lVA
KX+wNQ6Fi2Zb2B0y6LTZMt7nJEOgvW6vix0LBsjo5KQ9rvHBrTIHSlMCX2FSpAOl1t+qTJ1zV28D
vQoksFMyEPySeAUppicHRaYjqZHTwk+KivhAfM62+HeOhp6aFIh3VH165/gdn+F6E5ASVqfHl3pm
drhhJZL+uZn6DtfBweVqxyDYAlQQ+2/lFrzpkX41dNsjRYhf/ivEEkaWt/YE1cxEa22aVo3hEmIs
bt/Bqc4/VBYodqIwUIXEnOGVQ90Gj7FjgTKSyeVK/oEBoUaQXQjhcfh21Qr2ckJ1fZY1DsCztQHN
DINJ/QQ6+sI2/NF9ztc/XYgCtH2GkCDxIkqD8sUhK1zFyVL5cBPZh0kwJYnvtDCefdqRxM+P76F7
cVfWGSTSjakOMXfqX/Gal6VtBrEaW/hhxOOYQpkiZPhEAfE24gMtuVphg3y1r8v9L+oL4g+t6M11
ZAfMvuIqD+h4v5Tc9ZQh3tvoKJlxxy8mXmA8gtKH5xplGX5N/s70LuF7LMoUb/DrHajuUvlQmQqp
6mdNcHK1DrxXORFrn/9gCbFuAGrSTwkQySoPhKxSfHbXetY8NyuxPliHCCzj24TnN80TXr2yc+lN
jehR+y64zE9gk0NlA4RW5F02yRpXB5SWIvX9/Tey4vjwXp10xccbnouYkSwvK3XDrX0fLzrM0/QG
XpczpZV2VJLq9HsnL6XWDL17IRn554Qd8uLsFGYn0XOf5j2Yf6cM+spbvgCrYVqobyLvmvD+Yigw
U/m9A9VDZpvjQkZxrpeuzidkJNragO+5MbVUfWOqdDeM+m7KS3Zamp6k9lYSuJw7rDKfIYfXQmdP
BY1lX4uERHdBOos3gpafBxoNqnT9JyAL/6wlw8azx+ZO5xLabw5H3y4EiGDJYmSsInmfFaaucyQn
bNbMK4hdzsGDqGj73AmlPbNV/E8EFGEDIKrS2DjGRgGi4Mbgm/5/fehZEgwTee9TRkAkx2j4TUJE
/fsmxOXh0pxtIaQ16fNF8J8GB0sK70xra51WzsBiDayxja2VlyKiDMp97XV6e9lnhOMrl7SwKwHR
UNfpC22kNDgVOLEiHNje83LS+ZDSRwOSsrJThDW4lGzNiglv40PGf5Wv9Id0juRhY4hkmWx9Sz4b
VjHAiuga2Juyf8vyTDCgQz1uCJQhh3BuoJAQHDW2FYDAQUDBfx/iVtrchbAN4OwCuV2dfcHHGlTs
GvzgKej0xxL3hQ8EJwpA1MSBOTJAlaMDIEZ/Q+z7LcHqwhtQN+Cc12LqaKLZW2eCBCr6FFVJADN4
6Pmh2RK2Mx+rdkDx5WlZ9VLagIxKdesSVM7CfkTLtz4j8rtvRXuj58Nsd1GeQTn97IwqBxAdhOLx
sLeB/KWIUxFX3W8dy/C0l4SkSV7wpt3c2ydHOsQc8ZiwnVMjnlwC+FdZRMx+z0T0UjxBdjZFO+Yk
fL/Jqnc7dQ4cKhAfl7UZHGo/95m+vZZORrhbzqP7+IG/R5sJzuSq2EtiY2s50USWEGcQ4fjrJgn8
z1xdf711ySlTtD1b0iW4lXO/KGjVUg3H61ValX0IK8mTS/oRmz7X2ipWHW7ukc8ZZrn8VS2+A+BK
+30jAn999ggloUGq/neBtked6AJpNnm2pgmCYAt6DwEhNUtpPhI2pCFkURE4RcfjdHpZ6VCj4B6i
w3ycGL71p6+bTMdk1+uHFfEAHOs9ZQ2gj+/b/yUu5RWHELfGivmZlIbh7dv6/V8tm0V8bRIkMVdo
8xccUz70qvHTpbW1oPt5EKKcYj0yA0Vd5k5BjIr92NvUAbYXAlNyeOxTtrVXcDgVXemjy93I5vbU
FpgGm//HurWAbfO83ZAzKZIrh7PhUDTAxUomiUe01QOtJ57XkG8M0uRSoTkdU/76GLodYQz9eA90
NbTKjWV+Nbt4SMWujjc+jJQn1S61hVZ22h6nxHxRhIUd5t3EJOSiszXdjVr0iDWMcwq92MDf7Xg1
roTRKin9kmiPXcxHKTXfgTG40HHhiwPDulMffl00p7mR9iqCxQmpB1mYgW9XetINwk1nKt5Pleur
n9cocAEGkEtemzZHCXEPRkGdQhvENaUHUiDuRb3ZnVAVgiGR9yF+yPn8QRzc07ta9Le3EEz0Wlyt
Ve/rHHfC9F9Wya6UTgiHVSt54V2pAQt1W+OPyPZJiJvyi64JMcxpEB01a67xQIx6qbeYPdt6AxVf
ZzBhrCuoz+p16B1pdnaL5cDjrrb3i90Frb7U3Ybg3QTBUglv/JR6NSTHqn4ZCC1yhwJmnXDCVn5D
3lutDL14xAjj2PY0ALDQ03uJgYfHBhQdzO6b2z6945TAtkOYLzYRmKN5xMQNLbFsN7xTRTHp6EeG
ITEO+sQ0yM4iMQJqlnaWmjBrqxDW+FlINsiHVOKDIKpOiVcI0bOr4L37tyZSp6+JSAeJMihFA4/y
oTbIDspQXCk/GFU8sk6KA4ff7moK15rDmEBjJPGrvEhUOk814y1RPfLUsM1ICUQeClotLHR4vDqq
oZrz7n2Ua7AVapWs603Ug1jQW5o3sitCtvpPBZ0UMY3n+3vdi8Iru3t8qIT+l9flzg6l+kvJBlOw
Xi3DACjpky1nN/Hx3EHdlw6LwBNjHk1iwh+yupCnFM6trq2rK6z6/PCi5tDgLNgJyRleYZu0S6OH
LVnuTTGNj35WsGvh36HSkTfMcfP/zJR0jYbxMnCuIiLPHX7P+h6aRZ8IL9z+d66WbugtemybZY4G
VFhcKLRRe/O1dszJw46Y4Md5Nb2eD3474ojzDKbmyRqKMIoACso+8EysTuKAUKj4KBnZLsbX+lXt
vdkw7G1ECLPNiD58Fb4faLfd7iSXZP7yECLRFIc0J80giyA+DBQKFUDXFLrs63E3ROylZV6mT0FK
lauvU//W3NunqoHNgXm+r1eFxWopDu5qi4IvdJJ1TVg+/WcfGmzX+fnfDXckQLupd/YTd6c2Ffm0
AWt3mX+CvtMFADcERECDxH2jCOc7Gv38zjlW+QoAouSFIL8gQtR/dTLbhvPOF7dlBhqSdUwtgOB/
ynNsrxiNiSjNC64iT4nQd+ahjYAsJHdXrxD5f2jHn2+s1q+UOac5PejXJEIFZqtDBWe7KhEla79Y
OBV17Md/+oFPsk8LafF+Tur0VjCJ6hzPbQlxl01XK7psOQLlKZfu+MZkuBhPmnVsRxKzVvBPnzbk
vrXloPY+cAuHjR7sbkjVxgCTEbm1s+A496t2UuKHErsx8GJ555YWAZfh2u3chh3x4VxuRrC8Bs34
KDGEMBBORwSpW0/hEuVu4G7zN+ehB4boEW6nTwqpjVK7xw2rxoP2of4UUXErYo+PDN68dFOpGw1Z
hhaA2RgzFdamUsZ3GuBnEfKTSxA/Us8py6ckadb3GIPUqpzmchMTZvOYFziix9e7u1taftb8FjCh
ho8dJ+xagt6gEPLjk2CByllDcyDEUrVbXJXUdHmZadsQStX7X1aQFdVtiDcMtZWH1t2aYe0/ozYJ
ydaUZsA8NRKjP0JyFkAe4SHxYcBvpDCalfTqdH19gCRDCadS0sJ3GBXdBxa8GGSlyKNMfOI5vn/l
5qYYoMcXmap4aO7hpe95ULVX1wgSQjNhjgWYdFQbXSlhMDhFmbx/zxGhqcspfzGBaD/B8l/vaAaz
HJtE0rgUX7Kf9Mi3DgFSU/JK/6k9a2gHeAVxxe6cG36EOmClqqycYLmiDUfxGMWue+CWZ9JXCXVE
s/yJ5PRAHt8x7nFwpgeCadus9fMj8xeb7btMDGGPZJzPgGreValY93jXSDvHvBaumg+1iXpWryKv
YSN8Dt7Rjqc1qgC0c7bEAQMuwAcX3Vm4AAffk9b7HKiDW3CWa7BPnNbwGR7n5OOfXxyQmb7w+oTu
ohVmwBBOX8Xg3tmfvDYPhXwcFngzyEIamldcgwy5R/1mD5HqUyZzMvH+Kz9jeAbr6SDolFmu3D/a
Gvvm1vztN++qYju1Oef+mvo+2N1/qO6jdfY25Vis6SvNpj6PbF4iS0+JFYnIsbJ7QH7UhZZS74F2
LQYEVOuUr2PkX6bNdaKU/D+VnugPQVLTMukTR2rFTjTc/I6ry5NsuevHOTe4L2N3QLGl1LiXJ5tc
tMo9zo8rWfOYI6ATbuob9TFpzGNa5jd2cwWvr75/C+ud5EZ6nA6JxkVSZkuu1fMSVsyQWMH+vmD+
IxDXeLM91tlrmSZnEeLU4FfofaniogkmevIhqP2kIHJSdaeqO32y0B8NE9fXgdCIo1ZvNubmFgue
1PXc3w3LKATpssHODl9IvEUgxMDIZ3ogtRFVm67FTtLn0qJNcuUVIr1qU+16Han5Wo+ypg3sYr9R
g58v5juyVyF2i0ZUujfQR8hc2JqlhnJWQTxD3/dYS3oFml6ll/Wu38oOwA9uZtdh+gnbDZEkwjM8
jlkNFhjq4P1Y15qc1Th5cFfNAvWc7p5lyV+i6Xab5K2+Ms9btpJRSIHY/Ehp7QIRoP0obD8duFT/
PDUGppfCsVLcMw17xbGb7jtoaxL86RhxobwDcXcsq1cnwd3+H/PefvmA4R/iFLRSdizpkJL3t8PM
7SGpAtq96sipeW7l6VjlR50myS94dzKflWwry/ioSeHSnVkRjxbn5xhUyxADTzaZElIr1pEpzEZl
18uHP2XUJ9veBBIY89+IZ/YtU2EtQmfLwTVTYj1xoZ0Fm4WzVQiM66gE5YrlHaDcBbEVKXQeaomf
z2AFFa8vjWnQRfxw3w/TY4XlcHVFgpSrBhagDsB/8qKFvENQZWREcSI/At/h5GoIJyjMQyvr1ZBF
Egw/7qpt+uds0B3/FIHQBJwUzeNBO9ZHxq0rZ+qdtnFXpdgw94khHgdMhAcb6B7W9aWZDokwSgiK
f+MvYVp1/tE0uGMrg+wdvNfIn+tlezybYJJj2oAU3UGiM/WO2eIzsDzFvWkODPHlRjqay5IlRRj0
pK46gHB/K11YCzCuWZUv5EIYzo8MMkccXW0IqLvykc3AaZ2u042KSuaABpDwSqZKIPOjBoMwq3Gt
DXNCKLM4oZjcfdwvVQaPT9mbf8cgm2pvPHs6tkF5QIJVSXf2nVWijUiauEJJvyWPet7Ye+VnlQ+H
pPTFvK0CBCCuGm49nOqqfwwSGcRfZDFW2lvdhRua7nWuzTIRQiszJ+AK338SR+Xw3yKTIRVUFqhr
esyniVH5XIEUAytVO2+YLiJBz39ZvbMmH7bgNgSWPzLZdbsXF7NSCeXECryJoPN/HSh2S68vgS6k
fk3yUxvS8dunkKtNtuOC2ZftpD7YdtBBFwf9ty2LeuL9tefdxWIJQe/CudTDNWXfvu1IEVS7Zct2
076EYyf1ItkBt0NYiIykIKedYJb9Ml8FGJ8a6XbUcjDa9DCviRyYCBJzDuASX7UVSfi+Rq/IZEjF
f1Z5yAC+/Rdbko9nMjNh5aA2DXhWZrFLef5ixcF2isOrBcEKf+QMi1epVqItJP+HhRu9u2yrPu5c
nVmxeRlm1zGoFmI/VJN6JrWL7djuvWfvfTtMzcfq6Ns0ZsQCntqDmeZ/AxKBvltWYJfqNlZ8VP31
+F0Y5RIeSkLTQDfw+e1m8iWwwvd6bKYOhH+CNOzt6CNZLqNWjxDFDGEwtxJoVXTUh+8VNczuTeLs
bmOk0pJj8PpzXjRW2putmu5s2MmyBA/rVAW/0eRAWpKaxY1DjBpSZvXVCWrWfBs4QryosWnmrWIr
iJSzdESycULnKGI7Ag8BYf6gKhBC2LDFtcyhLVY4+8bN6I9H2PCrq4fDvzOOe29GI6VnKAa6OOhz
FWe4T8RIbmjd0BNSmNzLGAK++1o/NUTTAbMwVbi7Ua6Nd+N+3uuv1nprnOKwJAD5TTO16E8L5RMs
wUOqyl+Kx9iFuEMCDLGt/c0m26eE6fLpmz5Ts2qkx0Nrvm+BjpTDwAqgXrQ93W3lUEb1Aaf3Px1U
+N27WEUxxmeKikEbu8eTqi1L76ORTet/7z5q8Yoy4SWru5wmKsThr87SThct7XgwMKahkwRxvg4w
l5GnDpa7Ol5Gl+QKHgCCEWJ3heZuo1hD08G+N506HmIGd5ClvUbxZAIME+hMeaGiWtWh4ugIoO1C
VM2L9Z61I5hcBBezwXatIOs1jbni/BnPi33hzSynQV1ha3jxTSDINgZWYKOD4JX+5VRbVH2hlhYY
9s12teeYLU4XXoVTnIEvR8gRdllKQ8jwSQ19L1KIAKQJ7BPM5xsK3VQNHx/5MV0YcecINXYnR+lK
Q21Tdq4pOD2+rjq7LOohylk1idsF/SqX+tDkVo2DEjOqXUpo3Y0HfZSDJDEp9MeYP6HxwdljLmZ7
SJOmN5aJUbxffKN/4ckRWr+ZKxSRMldQvCp+vKlECWEtXfJAYgHRyIpwjzI7IXT1xWZLpTFjkA6q
y/bWgBnXqgfhNN7vOfAYMgVIqPFHox4ABFrGtCQ+XGmHz5VSQABMn/7MwV+ttSJNF2+FEsPtExkn
eL+SItIZrO3Sqh/JfzT9rVtfjnTdQ/vegpr2bvZb3TxEAYzA1lxy8bRgkrOk81t43d4lh4cXJCCO
iJ+K+r6ni4onHuPTt58/MPcXsVgGPAIwpZFs+wlLgwnwP7xUGU2xtjSQCaYvD+vRaajraRyw0YlL
9JOXwcZPShMfYs5v/0us6kkN3dHjTkBUmZvOH8nuCpQODRXNPXKRLaa2FwyRFVnCcR1IKmswSp5y
DWC7hEWVa/m9P/bFptFjdhVicJPL9s9IN4mV2HJ5t7uWynf6DmQeIy7ALoYSdw47J/AqJZZlh/vS
bjuLjbNo2vJzYuK3iX0m9QJyLd5SC9XwHPz0CTu7Wkz7S45Ix9ELFxG6HjoI0QbI1eOPhAosWcq7
/2rO+6/aw4KqvNYQ/6D+mEHzfANFe6r8udCew2goOvmkwUS5OmxDyr29Xd3qOOsQOsFd82pSsqOL
6+NLKBGa67K3TZgZ/7VDiwlASvyFquAVUBYoe7z6trWyLPv1L3eRLfRphWI70IWQf/xdXwfutZUs
BCk3yTwKfmWxJZ+yG3mVdY5cVZi45vz78CEKQ8RUVz+9n5oTnQjOHoK2Agx6Kg4KYm9TabqUBLy2
lvDuB7JvJZyiWAccqdURaq4AsRUjBzZNC+pt0dkyRLLegjXXPHqCNWvLn4GiKV/zbN3ln0SQ2MBq
K6wQGYVJYo4SDWcNwWaj89WtcTz0Xkh8vIDFy0vJOEmTn/phEwimHBIQm8sRQIB488IJFZZSUZ5b
yBLOJ55mqvuChfPpWysSJL2sTMbnaEiBKPRVRThBDKYfXgMAqPoXzocU8IF1xcskv/67O+S4kTS+
0Scz/YjhZGsx5gRsRM6ZN9IfOwAU0NFhx1RoLx1d+UrSkeUOSIgHDgf0Cf04oExu/rG0H/JtaHxT
7wxZZkGlyfKarp1gm4HN4UyuRhdeAkgQrH3oVYSmNh/dxIg6Jk2ZM+AOdLPmwlqUxyCXqgzgRzNP
gv4XpC8aUW+H0oMubHZZeYKPfit0l7QTZWLJfWpAXHHzPN0F1mNaV7a/YIp4/aNfLOPuqyn2Ub8M
ObA3ML41JaFiomMwItYsOt2AVFLIWCSlAMkjaaqEkVBvfFH2Pnj/KJpGnVkn++AbG73H+HN7nQ8L
k1PQwOnhxBcs5oVV/nmNdxQthj1X0D3TZs62D4UiFGsltiJS5dVahSq6w6UqdFA13b32INxlWU1U
AJ7rjqoMLlY7m52DFKCoSQpxP1R6b9EnDI6JM/SDAIxv9jq5wOre0XYBcBLjecQidETG/6GGxbFp
iG6LeTfjY+SmeXLXPzdXB6HKhBS8wL7xnXKYHguO+vlAfo+HLgdaqu+sw/2dIN3iHLbp1qJowbRK
NKtViMaVd4YUKj7Zx9wZ9RUSCxB6M7rz77DThYHr30kibB8eGD/IH4bixlHz6nsdKyT+dwyvRTny
MvlxyVe5ns87n4DqHSLDT48rxwEyHS7NHSf8x63Ix231VPOE0ah9oXIvtOpZL4UiPgKno+N85XPI
Gzi9oo9/UMKOmaP2EeqwDKNao7u2BwtVxVWAlkE40X1NT2HbgZLY3EgMISR7Qiq1TV5ctFxKnyOy
QtcqkIvoUePbKXxLmsnI6EyqW4XP+RFuq63rnc9uCteBT1UcYuKPrydyZmT4ctgyP3idE9w72JmQ
gtyqm6w+KBk219hL3CVLdRIeGNt5NJJb7DfjzswMn2F7XVHpIvmHql80QxfDsr9DwujdME9oqW9X
KTMGESAd47Jm+1oizpoanGdLuZACLgE2QW1kpIE8xNgbztaAWC80ZMwvnsNTkFneI3BcNW3BNzfv
xwXA4eyX7tNAuWRf5HuTyPb8ejzvX7JHemYOgUzSR+FVV5HF3eDJrptrVjpVPTuE71ppbY0Ev6Cu
I6T26sREL3NEUqstX8yjYUNMjKz0Msky3U/Ra2xRJ6mG7ykJAf/xKZla9YdK+jk7k6oj0IouwUJi
C5MW/mBho7ntpmMrKuLx/iKsAFYN43jA4myrl46abxHct5zdK6l+K71H+ikxMgbmM9kEqLMeKY2u
V06w4Lrt/f5R4YFhRFyjEVZrdTPBzGL7fGOR+VEoGsnuLpxmNm+Jvfipajz/SuioqT1hW0yOzDvx
/e5/s1BZ4ZT4jb8Va61S0YCiIf1Wsr3aX6cTDhuv/9dkzPcIzB9z9YsoseWmeDrZub6n2aWkjDpr
dsnH/19s5RnohuNp5rwpAIhaZsmqJl97LrYHmHGyP7C1WrpjoMscB3+zXBupJMuFYS2/H8/PwLHn
wQ1Z981PkPSwWOOFh+iM+zONostPI15N3PFu8wZJrmLukaBPjgxJklBbz59cMe5VNUamgFkHZy0q
mHzEvtLEMbRDYbpslC9ra7irnlaZmxYHBK/r5QfpX5yUu423dusl4cjHwM9fjg0mA7h6jqD/fbFb
8apLs0ZZ97ft+i7/utJ+aG6gFnI3EMWR28fwDjDRZO5qxY87IALmEaD0TG6YaJSeDjSyWxQxQUx5
DK7JuJKz9+/1C00KgPnlBIqNaDJkAI8N0ZusPkti0rePX636kBintKRdYSwZoOhJUvn/oA8zoN51
PlBrtnNiykL+PEGfRicxfgJt3wVStS0JCcOfk5PN7wzz4R0dz+2QNE4h97XxqcJJAKguPUMPiCJS
BFwn1Z1BNKARsfjCPadAA0RjMkesmngjluPhOSJ0frj5zZA1mg6zrkHwdyBajWZjer/qaqA9iQeO
PZquHEee+ODQx9ZLtuBEagIhm/mPQWwHMO6UpQCiMJD6G/ViWkSm1QI4CykwySnYbRyqwdxFZLv6
OIoUP18OsDq+SsPtIziMAQddibvyA2qV2Nebxaq2J/3JjUNM7vNaMQSmuWIWzVhVoWlTPyahOX8M
VeFpqa/wLhXjdqcNo/UnBxVG9tL0CHtMnUNic2ri+rwFHLnACde2RKR2FTVwR4w/DfFl4MM7J8C/
Tf+Px+QwRDuCAHQuQ7EyJ6tWAneuEPNiZsA1kQ9oqjMHNNJIFO9PhPQiD5J3q38+HQf9s5YL7Xnr
Bn3spDfGM067OQLx2qOg8yAxMfCoYZMyMU5nFPWtXazlLIuWNanW7VsjZmD9LK0G84abXLTD7F8t
xAn+Y92IPzEdkxYQMjRcZ1Gqx+iREwPYILgq9HCL5As3zgvhmwLBVde6iTwDRV7yj1gQacKeWee9
kG0PodOyRHsLtV8sSPXIdpYz9f0Ak73erBfYs2vJi8gVP7OVRr5rG3UwFHY8xPTz2duWybng7o9i
UDpghRDY7XTCXlS8qihoyRUlNBz/Q6hSmbmMauxD4XNWyfKj3CKz85qIK1jFF1UK63ivyrkErKqC
Y3FPMFNZ+ZcNcuU5pZVd30biplAf2CaJ2+eXikX1FLkSlO//aUeT3qChsBMu5n9/Xsv7dbdIsutt
o0hwhjHAyCumJ2CqMYajAkJAW1xcov3ZxYCBa7nKV96f8OgSsv3NqD5E864pBRyM/hPwIBBwbI1t
Z1lzeKbzl8v/AyeAz9wI+hk2gaIAnu0HEDCGxGPs3dsl0yzuJNZpt+q2HPC7ywlVvhWa7f7pzkMr
vFakuHYd/QID2MdYz5vMN2WpMdFPRIQr5u3oVbmx7JIp9SwEgNyvXMvlJS9/D1CcPgHQTOX3ysPO
r8yBChLFjaMgMcU5CTJGuwHYKqLNjsiaFREFA2n1R79DnSDtbI9zlawNkcsw86pPt8qEZ0MZi6cu
4AX21zqlv2BdJh8mWf0CN2ENhcQ/EJGEf9uVFSAbiWLGweDPRpS7by6Zye8uGsN6IBwFfNFKfjVJ
L2J9R0tgTSuY6AeaJlPLF4R2PSI/Ke7y/rVBKy3u35q0pI9ElC0ndPOmiI9dUMRz+ZwzzpQRbjrg
nDiTgCOCkcpGe1PKm9RoH+zhgmAZHSi/1HVCNXFJ9FQRCOBiFWTo3uyvaFXSDTnC1KLMMvuAXsQ7
oTJrlDhKdGvcvwWTp4WFBODNS3BNcMA12jNRm6sr7t4Ve7dGUo/bcWwormSCSW/+5P+pqgj3zh1A
o8M7KPHSqJ2iJESIOWk6JxShUItpMVh3di5TsWVmBQWQaLdpnxUEC9zedAN0k2Vox8b/RnLC+ZZ2
yIzwy0GnRtFe5pLNEfuZyk/ONLdHQY6306KyXgeDVusEfZxpjJzkoOUyklgF1Q7SPQX7sVNCvWIW
3mn7ofBKTDXvdZUcT/VIt4s6Izj1Qlkt4nbxqE8DBsT8Tnilxs5PRt8s5vTykTaHujwzFobys2Qy
xUJR6rP/6+kv/jZmPvf0wHw34tkZY8xxEocO93kJ50SFsE3sBPYrxQ+A5iLgiq9VVlWNU9pa8OA4
aCUuimE4J7AFaPsLd3TBJcNs07PfmOK9AL7cQ+YBe4zipkSe+4X1xKoXtBueEbc/24TgVI/X+0ZG
eXwwZp8t8NMcSL63rRfx23XvDDfc0jnr5kHYpyYDuAE8E7zWF8Pwl/j5KNDZruMjtjxFfm21f8AV
tEPG4uTR+XbT5vdlBoOnBye1Tao/Uoslu81ksq6w1wc6tGeYrM5tB2ozA6mTftzi5YpBTz6wVLC8
gbQj0T2BR+XQptfYXQfG/sI6SfY0jmxQfQmrto/Twxgl2TlXXa2cbAaxqJwb81AeO7KQ9bYfQI9G
PKjtpbuTe8L0k8A9pfjeV/6IXCQVXYxt2mov3oA7ZVXBs+QIV25fY31ZkuFbFL2P6AMn2ONw8ONp
MHMU6yJk+1QlIKtgg1sO2kKlfDMw9yOZBj8kOu/p2dkYJRSvXt/0wt68AObx7+bM6uBKIRbZBCgZ
ZJbO/uVUo2cA3+fdeeRoquQHtQZ1gD9xD3dK6/BLx3lXZRkS1HPDrTxLiGqMNNPavR25USmWcH2L
vgzInTgd8yYxapN5jHmhHybIxDoefeMXJg2acOQLx4h6VVSlibbxBMu2mqI4e/5xWEEkuzL9mYKW
ar92d6w0LGL/eVQPz8WGceHmDqz623lj50+TMgrurKrkx0VumkowjoszcRMznmRba3yVUHl4UJwc
iH68EvxhCbvodHTAjcCoFL+hTito4GCXxHr8Y1fkkVd4Voxqbpgfkw0xlJQBQ2EInKwtACec+3jG
1RBbyIVAJy/ZiSCc5p9lXWVnuxFr4gUlOxLkgrNP4W1hf0PzVh7+2nuAAXSI34UQKjFQRHaDCdZp
5ynLE4r6BZbdukO2KPUx15l3kFEpFcyPf7ZxZecyakC2e4qjQ50q5UyJyJ3dDs4cVv4xWSNNSwLR
6VFnm8MO+Gr4Q3IjgpYm7OIbrMrNbrATHzKpy6nhOHtxbiIX7nAfgFO87+PJLHLswF76tMVv1fhO
ZReTudrkJlMRBTyJL9JNfqORl4JKVTSXFdRdkyvDi7iz2bQlTPjtejr+9gCtvDNZBfHLGKnQaX+q
BOxWP2BxVJpHyF7ksi3GWF4FgktxiAc6f9CxfbHi3YJnAkdZbK3jsM8f+cWCj/TGnL16ALWUFuJK
x7Wuab1v0pq2ChFcmMWqNrgxOhU3PQfpDo78J6PTYI5PmLB88fdD4hyb5ewiK1vu8LD2Vvi0FC8g
OkORuJLY1fJtusrnNlHxGcEEy4JOPxiVMMTOTJUELxSL695t1B/QPVdF/gaI1GKVytP3JcqzSF7o
LGSntqr0yuYg7YtZriuOk/t0/nCKRCO6n+z9C6sNh+OZo2vHxBCbG+TSzbh+85dpbCdaOopa+Wcq
JgnRKo36bTD/MwuUzx2lJUjnU0O9ytdY1MAAiBRE//WHPtwHKU2FlZZg31JjFdH4wmr5Z4uWyR1j
ZyGlTBy07bADAtihIHEvg80UHjRWreaRH4cY1ry5F37uiHbqFf78gM74AJRYIsvtIpxfBCPxYiyP
t0bsdgtBFPdi7Kw2BmNKoFV7xFQi1xv2joTac4VV05PwN1oQbshwcnTe/93nvWnA7JSbu2As78Uh
LjEjk64To5BObQMgFjub4gGlTj0e68OKKW+QvqBGcO3bLRvrCnuhUf5PB9pYyFqSk8s/inJprTqT
b/fzi5ja0U+zIhQ0gikHSRS9Xdbh0C4Cflw9K48q+3wFjjjMkPd8zNoTaDsIblkKc8T7tUoxBYv+
rgh/1hzBxr2LuLjvL6HZ1Z1pp1guz8dbIhSy5vJhleq9IOEM9Dkd5v3lsjx843/WjfxqzTYDQtbw
KUPM4+SocV5lEIUD0KxcljtFJ7rU+o66BlzzifYm7E+WV5cc80rgqY2icmnzJKh68SCTfUa4dG4R
fuSc6O1e8JIZk0JaJewuqk391m4T1I6561TIq1iK8opdz21tlZ73Uoz+UuM8yz8RvPPhlAcqrfnY
qloovOf3kZbyMx0AmnDUuFVrEGnzIFeDIISmaxmG9V91X6w1B2LDDYOArWGK0tl9ulKLdx/gw2PC
x1dJgeG3R0c81gCR0ApYBFnBJQl9t2vx6784lvy3L22YaRZd3HeWWnpu4vK1Kp4VxCImKw3HfeFS
g8OqqVThWfhhdPqgXFtE9Yzsza9yDI1MmUDvNUW8yAYpMzMKI05kTlFHFvfxKMSNYlPN/wiLCobu
2CACZTzn70ZnT+2NGji8++F9U1vArid9QbNwDcnCcqBdvC3EdkNPpv9H9fFWgjjWcOncnmhPvcUS
83oMdyhmw9M3BRVqh0d1DW2nWSyORWTJIgzaUYTAQUSblW5cOVqv/RJ09Xzzm5HrQdyk+1N+nelA
YfYHID5CXxtjsF2YuJqjxDWrQDPFMfxotZJy+H9yhcUFi9QoCVzTOCdIStz8SOTuXYpdfDYNucdT
VGjAyOT7RwvGbkP1JhKTnJfmGhJh8rSub/VRR6dpINKqFmF7hpfWBxgKKr/eWiPayMfc/tQXBhdo
JX5BWcf9xtWoRPQ8Fms2yY+q4K0yNTNPND6OOSfwM94l8IrgZdYMuw6ERgnp0XKvLI5WUuyDGXPP
PXXjAHaHmtKhLU9Rb+l11L9djmlPqD6C4EgbzxKYqUkbrGcf68U9Y89zoToQjlu1H+1nUnDd52gG
IEhg48rZasYkWb2BYYP0fECtt/pNuMWb394AcyJQFtSgqtiIq2Z7ky1Xk7NrVL2DzQ3hJD/MBNoj
on2PaALWEZvb8LHfOO97sGuGXLwDpovkXQrq721Vdnt5H+bDhq1nUpiHXBr2yDpFdIvnALkAlGE9
/KmHFIhO5JYXsAwcFtVLzfknj5CalZDVFgmZF3idjb2EDv2WUbcfchn8bSyJ7IJk8rH/PpxUO3pI
oZjj7GtghSiPsX9KhwjUWMKEu0jaIuIs9TM8Sp/omfq1nzFTEoL3V4zT9oJFF+G9bMOG1YiG5pXs
F8ITkFZNwDhNOYy4dZDJAEhiH8pg8h8OPa1cUjLCs57EzrAl6sTjvMokH7feDMSVqUaw1r28VfVS
iFUcDU1Up6yoJsg4CGYuCO8yjKKSWobnYLBIu+yUR3M/TB0fPpybsaDYjgLwYiw26INLvH0Q8VfQ
T+dmqMPi7aD85wqoxaNodM4uCDJOo8mEb1RGuoDNTkKYU0I2mmup0dVuAupSmr76meFqb/7AHzGq
PuRrvli3zLseIghxDCu34+3awI5nJZquVhajeYZd8dDuQqzVrXv7lVzMEB9jQ2nKZziRIdkJ9IMH
UP9CS4am9j6f4uPf/vwyjFtwWEQNkYmacjoNVO4GkZgLlSomr2oZm4dyu9lM+OBLPYO6OxD5Lppe
5ZxGsrwhnc/w5z4clKjBCb9AMPzWtN65SGD8QMmd9NW+pV6k3JdTZt/L+kNuYjFxzTtEvVtfoVi6
1V785JAHQgwckqn5QtOqw2IOMlE7FIvd3Ck2hQnPUPtyk8NvzCcGePwIyD/dh7lhmMbwSSbmPfng
uPV6AAG6X2vkcyuNYmEqNCVYXsSqlSQ4YaArRSaQEEfpi7FAQds9I4KMO9FsopoWGIMVi5B3Wvn5
o3d50smuK8BPPG7Zvby4qovmf58Vqx8LUB+SWaOCajzJCY7KZvaZ1VOOLeJUAG5Lq4WohMSHar2o
ytmnpENJrOzvuhyIrI4V01BD1i+I4v1VTOSDdQcMDocUOJBzFdlggdJgpnmFtFEA6R6N5toUWFP8
UbdX3c5A35RJaBnK0B+RWsDKAbT52l2DPKUAsV9h9u9CZGvmRPOBsW/b05RO6ohof+mYygj8kgGc
/VufZdFkY5SUhUEqTXD6G64gnt3srTW9WBE/B7IRdxbnQGqiizDV5jqN5QGbP4r/sx/CmsGyXxBV
R5C8kkKQu+1qZ+w3EiSmCQFsf28AoAmsmpXIEJLr/ZV4Xqrt0/iiCh1mxGkl0BLik6I7jCBKSkWd
gBuYEahbQMU+M4KgVobYbvLRu6VoC+dll4ult0CC8bIYg9gNXXqAtKRqHY8D1yKB/G+aA4Zf0Cnt
HEpQIgLO5AsGfyufTRo6Dmkvk6/+j5CQvRM2gR6IvzBYVLko23biMSHeSg56fJuVX4OjqAZUsVyF
45XXLYf+vA+dnesiYXRwnUgIAGj1mjrFMT5pYM/aRaS3DeX2bXhzgz8ocN87csu/lrvCKDGAui+g
4748ZbjSGXqpUQUHRxXqvrsntEKxVb8Dw00Eq6L6EnWXb1lUqVE7hrS7gkLD3CT9pzC8WKX4xE5N
4TEmcsjQtM7+LQUpzS5xvsX/JKYkUa4Thdycgp3+ftfglwa112O2qcxuOaZaFDmxm+BqFxWHybW7
JamTz95qO9s0zioKAvfpTR3E8t/UTVEnAhiamkzETSIKLHQM6gSs4I4i3OZdIsL8CWjLjcui7UMG
1aGz+qX8+hGjNs6NPpoxunvtyvQdH8SPiD0AexggNsM3B7JBQ7gyM6FN4dMNMxDN+hXXutP1qEoA
XptAKakbdowYIjAKREUeKgF/yq0jyYDkleAHNc1XpOVNZIZL6VyhWLSGYToeBDLKcQjrqefTCONL
O4tscI+2bAVw/9vxUeXB1krzZAwUCkQshOZs/EqMt+RkLlQ00SVAyisq5KKXauTPNx3vH8G3FkXX
gjnDGq8l144LrjGfxq5i5Op+m8daqg3U3SeiEPpnQWn+Q8LTUMqHje34SwoyRuzea+7iXCPV+WDh
WKiqpyZt8l3dGjeRqie/LbRDvyDSaaI5U3680ZQ6PemaVEuoJi7pDNR3+vpPsFugmZeQAl1oyG2t
fzITa3QPmyp5QNsIRn55C8jmso9ZxIvXIWY5OeMw72/+ZkliuilVZZ9JMR1Nvgw/5RNkfmynKgBO
UcJZtaTN6Ec+j1CFNoPFhvAhUDVxVaZHiDBgUIXhXQNFbwyHOQnyVmZXHc44NTPjPllQg7xoasH6
3VnNoIL/SH8N7xXNOytRKPiQjZzPdfZnQ0ebc5BGrTH0ELPvGyIjuITpp1zqLLls4UsK1pJ1wLcU
ZoROhqehQFW0toFNQxDcYvUy60u0LA/RVe6KrJ1sqU1wqoLxgRsYKfWcI5OHYjDIr/eKGeryYiYm
R9t2R7EMpeZSlwzhaK5pKLXQR6oam9EqsE0spsylv/m0P3q1zJbjugQ6QBbWm4V7cm5d5M1YZq2o
Ga+Ig447SVgYeIkOkp9tSBrdIjjf5KVcSMqA/beQW1OQU61KHhtQzK+mRjMmxAkynOXzx+NDtBSr
hL1Ok39BDsSD/14vozUFimPcl+2KngjLGIXVQS8bvZs8ZlM9HzUp4XNlhk9H5ywbT0CdINxk/VA5
N8o0qfGdh8ScMhaeboQ+8wl/9tT+Ruvz7a615xPwjev76urV/W2QMCe+jxzk+fWzBA3KBrEIXjod
BCX0EPR/HIipgM2yx4+uyX38BiOTnrNSJ/uGxCDdWq2SBj+z0+xyp8liMkIXLBH0bT9lyrOIanjQ
kYhIP8z8vwW4XzjFbf8YJZpQ0TLtuo0FKHFWs2d9LWdCp/Gn4qiM8dns1WsVr2y/zRxPHn7sPakj
VTNswvfa8mX8m1dyqL4fs2lgcrToec1FmkRJKzjM3fOWZdtt1yMG7SXt0PHw1JFKO+5vYRblLQAm
sZXh7FcvBLZVSpd6hUtu7bY3dc3WSaWwnXW2o2m81+j/Z4DXOvH4RbtXDbvaMb5/aOWh0G2MrJG+
e/Tggq8kisAkJCEct0YVQbLDjgv0Xm7X0bhJuFusXIODew6PFS4e4SSV/z24lJ+zWOrrHtQ/03Y/
/6iVr0MdiPpaGp3VmwLy7p82zr0IZPnStc42A23WvBXj1CGADLu1NM5mVarKukAN0xTc9Ux7VLUb
OOBwnv/Qwd5IMg6CTUsayDe0QwpfqBkEAqlcVp+ILG0WTHUWImb0AmlGPzX2qFt6AUa0EKAyJOYT
FHOpW/K6oa+wJE3ITP1A3XCLjOGZ9Ima1O7NIUbt9uJBfTPLEufV29K34lxN/PCLFURkX3JgJ2j3
R0GqwiSz4ztaShVDnhjjHLtfGX74MEydAJkRim/KDvOKI0I3CZGy2ITn/ltNoT8siS5TDTxBSyco
6DCz5mhJhPAeEd+NoS5MIn3IhMPoflmDa0Z1NDn4gMlN4z9PnVu0PwGlCQjHl7gl9spqcKdN6Trb
jCqEqk4G9hPwuC7oI7JmXCzjE6hv4ZQB+caOb79/VmYFvTKhfpM8cnrSAs07EKSW1cY1gM83nEr8
MmUVHmA/5MPpvQAQzExp5CvA7hLP99W+Nok+IJ0cjuGhnqT39N9KxdjePyhDyskVN7Z0IiYZWe5U
X1oP1COiXOcrxTGVzfRIQfchmNc8dVfX9L/u5uMWhP/Bz3wToVtJmiTCqBCEenTvxpbp+STpyU8K
2fOPQc3z2kKbzbN2Wb6OquJ9dfCCUsTc6soWt/EbYxzyVX29Ghqezgd+zdDVgvV/HSGAJFBVU30N
u5ajxQ/NU2qGVZmkCymHEV6v2pKKrmhszv1NhDg9/kgbBzG94HT8nGCZOQvdYzMJ0ICQ+dfKChvV
zDPiOsXwjGzlb+9/Gid2Wgj++iXddNVbEiKpXzMbokishYQqcgc9uDQDtAEqp73VxgwGvJIfrv93
Nr3qkpKxw5vCrlleE+ZJQ2i5ns87B+ppq7+PIYmoh/ImBv36+LHKwFPhTnkncLs02RCFoxSi4xms
Q/3aypB2yIHqKHjDiS+1cSDtQQ2KRnrF8k3LJjsFIOQhqr+NgdTPfbaiGVeTH8TeBqXdwCKP7m30
sZEisy2sAb5NOhnsBOTe+WpupIRWoKL1aZUganFDJXbGy2FLdGHppl0X3XyajyM5Z1Uq0VOy1Puh
Ap/eCO83Z6CgfDkwLuqep6EB4pW7vabPkQzp2OWdcjyBjvExprppX2jF84p/i9SMiJEykExPbYgl
hxAv5hL54h95oD4glfb+HsPGo41fpbTKSw0H5+esl02F1cDdRUjRMpNn1GPCAZhtfeTEhD3CSboN
JqjmiacMOdqtpJPbe2QLPMjLuoFtGgwIiP5ZCY+Q1stAdE0c07gGZtZFVjk4iIBe2y48GPsl4jhB
AmK+fCGn0R9kHvisH+O/bpWYwXYGghE9G4zosiVVOuHYGnG5q/OOOKJElS0ugR1AFxIXbJs0gn69
SJBey+5VGQTvZzr44stye99BNztaI9t4n/MGhOEjLXxpKdUeKHd584mBrSbjlN9i0i0YCkyxblOL
nIsxFJIP7RScLa4FKaR/bqEkN/1uMx2to8CtAv1R86NN7YotGYJfY9gDkD46ibtuBLK9DCk0RMFN
0/P1worN/pbRuUWx7+rN9Y3TznRZfsDF/i5IWHZ96aXEN2ACduC8O59igOzXyyFGrM99NAIDvGEI
VCzpkWhz/omxMY04t9r5K+4IYkU5YYINlADM5aIOJZWHTD/RG/2I8qgj4HLpXpGPAuiSgSw+iyl1
OdjGRP02r9CPzJi2T2J5Sk5un4S+i1W2tgm37nxW06bz9fTxff3vJTKfxGSsujaiHayHn2GTh5/0
mbxmPEUC8hezqLSzP57vRlx3rMMw3sp5ojuqMGY/ueJW/MprMRloUOtrpFVAjbTJ2qLYkTI/HUDE
oA8aOJfY09q7KA+jpxnaGKbgYh46yb45bGEDlqNso+klx4F55zrgDJ0U6HsC4o7fu/hxqNPyQSn3
ep22L5fG8g1UOFxybzgaoUgS+wAHsF14L/Jbz7GSExJXrUTCaii5SiN6nLoBuBLUL2kEw1Av9od9
IZyeK2HZlWAbccFd1cXDjjyBOaT8kQ3gl92Dr0iSbPyDRBkiG+0wc3pVY8yTq7E6UaT1He6TOSl6
Xf/OGSUlByndIcM7C2n2ntUXqhLZP6ftRFshVXLx2MTW3NcOVEnu1FwjDBUVtDIBYmiE3Fc4nzNk
gdF+C9PSAcXiyKT0z2CyZ7IOWL35ScLD/FvkE+w5ltY0EzFEW8fXUOtajBEUudf/Nec8z5nmAynJ
Bv5AAfnACS7nqGas4MsP202wlR9hgEV9voNYY4RV1A7owBulpj+MIGwl0oGj8IzFm8pYIXQqTVsb
cC7gFUN0NH+M/qJg69VhXnVZfQkkwwOJxwPitL0zYZPT+J4AuEbCyQp9Ky4uWHC16OWMZXcjbYKM
HY7n7ruhY/pjsUBqBjg3iCah/aBOBCydQBQMnX9yYqxY66dZTnjB1RIXnkmkueCi62F4ZW7GSbXO
INA9ct1X58jeo2jzwq6LoyGAyTDGGdXT7iJb7XmrydhaxFwrOLdiisxzRmWLfJXC42AXchyH3f6j
LtiBEgOsqkcqzOkwAXqhM9ZVxIgc9ctH9xz0h6voOlEF+bXeLSHc25ZS7TGUE0JK70AzkuKJgyqD
DWTDLd/MToDXtTSbLvW6rzMUEUOjg/zOIs+hcr2sH6kY60frimoWTB29V/WLLYDIAAUuioBSqwV8
q7U0MTzc1u/xzXgQdScETWJ92Dz+3qLOyc2lqJTjRvedXoBe3ZJZDyEAhliUvdkV5y1Rpq+/xrOd
KanSWR5uZOZvoTJRPRSyLjMKQZCYKdxEOAZpA9PBBp97DpH9/6isOjA/7TwdUjCxVRzSdItvzZ2e
0ddBOiwN3jSYqbGtW4NjU1KBvBLlnSMc7ca+1fTnZfV5toQ4L9OjnSeQJ35wKjNJeSjgWrKFmohI
f1oh8Zx2q4x1iBME1pxwu7mJCsBsRKbre7HO1YltCoXwRij374nJHRS93MvTFe3kGOwWqqF36ztY
rbJM38j1vNILDX1fpN7VpceEFZB1QVwUDM4L69FA910S6GfdGJq5SMWI9YeD5k6yyehET7KU619E
lX5ixou7EzO8o0SRX48pZ9+ruiuN7oGICQQ9mDAkNCMXIJa7N0ZD/0351TGtAFkSQD7NDqTEl7df
diIWQ0I5JTdn5L5wIx5sS2KfK5Oii+jv2pL+2pQ6LPymrFSSeeaj9YPg1/kldBvK3QZZibIsqIqQ
MmAh5/DjFa/pdoDNNnz5Ag7uZM3Pa/6vmJjlZCyiXioai6ulnByqPP8252fKmLHTR34UVjlesi6y
Ryhi/+lBfD8/0CwjqCq68gq/Z3nP2j6Ci+mkSnsLJdFQ4P4UsCochJbAvG9/cE/mjQO0NaYtZEEy
nY41IKHnsJ5rI1Q2vWInzivB9QaaTfrwnxWB2PJQMeJ9UBecciszUpEbZ3Hwi4UXgQb7XOjdrLFT
iZDd4I1d1uufXZVupi3Clz8TkMikCMIOVYALzuqyRKNdg72NAhwtzDJI4emvW3WB79vQw5QfHElv
dZIlwEgLc0YRizaMYSD40hvaI2/4y00C6RAGvOBtIS/CFTH1oBRWy9r0+JvSjZRk9PRyUv+t7njB
O1g8gD+gu8ehfrHtqXD5SAAwUcoOPGAkJtJ3mn79nD8UpJl7oDGg2n641ZicsoeLfi493y/GpYrv
LqxK028/ajZHepu8qEXmPWnWGKYmWrhapGEaC3HVk18HeygEydEkz7yuf2BSDq09hNXSQL+nIgwa
j5vQ72NtU8LPbDqvSaaofkYuxT4hjZX75SWbcBUnht7SA/ZVA5XCZWgBVQ4dzaLZ0VPRLBQXu9IA
qNG4/Xlqi2Bu424LOhfQiv9dQK1grAqzjbXRNb+TJHvBRZjOjqSrUhAv/0BtL41kmG3tvrJSOHPh
9D8XKezbXmqcOCr2WCLl4QRbwP6L1AIhurq4L2s/E7K3/Aaust2bT8YusKflP4TdkZn8bQQIfoLl
dzxQ8VYNH9eJsfZiOlLSXnsEER4cx+vOxM9Au30h+FJTgYFagB3L+Tu1xLgltJvii/czdOgpCheA
hrIMSDuepSpUhb4/70D3K+5rMgSy3wukzlZCzfTmCvGZIVcWxbtPwpUdzuZ0uLdgKByNNx3BDabD
zaFP6AduMocBWbhRSvbteAlsuBgZlIffoUEA3TNTFZH9y4ri5wqa6arJ9W20W8mMqcwZ9mx5t+ae
H99tFgUvO+m3KLFnQfnMoHbMT4I2olfIwQNHi8Sj8aDc9xL1ud77WGoROYROX+0DJhBxKFT39ufJ
KAXpDg8dxRojPp7oYR8MIwJC9sGWs38BorGdLMmnI3IBpmQOgakC5msho0TZ+GVgnNnALfF1N5eu
bssY6w3hcyha/ZZzaxMblcRyiiBTebN7YNq9o+j4+I6nC2dDgXFCSfN0HwvYX+1QIAacjwP2HF7L
f+CNWSD54lRFVxEYyth0fkem/eQMMkhSUzZTVOF+eiG4Ob3bCgd6aR9Tkdw5En4KjVT89KoUiDIW
2xcClxtoko0kwTxvbIG4cE/mNw5diUYQ4Rj1hYeC6NKenHvBHnd7SxtP6yrMbvBEOjC8gPaKAJXZ
JYhTXSoIcRbrU3Zr+R+qR1hIK/i7zvAbxC45rJGQZ6CMRkaOZopD8Le0WblhRa/IM+YBq1fUdmfl
IfF9I8h0cSokIOaFmDrPdra6IdHTQPgcOnIx+b5SqkGiU7cJJYSHYUQQ96XEvp6LFvO6TtiYyIYM
IwiErbkW7Jm1cayL9nsLvTSeRplVyz1sXQUqx1MDL2mmlY03dFUgljOfScs5DoBu33J61FvTpWJ/
SSiGjIm1Omih7uA6ISw1QgSVNF+DK2suwyrULcLbaXiGFTRUetC3oDGceZesivsIiGu+OjO0Fvsq
2Pxu6USZu5pZyAs73NxD31xoliE0FXR5iL7y9/+eVvdJ9IBK3hXTXIF3pW9VEIfGidJ2qP11DLhG
l+0MwCLvB4deehoOkKtsytrC5PnrbH6W0WqFlDXk+aVcIl1dd7EdTEyZaQa2tUnz68otbtM3UoMP
r93scrLG0iqeFKRqsCkcX7hdD1xYTS3+rc9zYQkp4MQgoA0VgRFTidK5G8a3JuoKGoppTuqmHsvi
lhGfcUvoqN8bIm2mMHfSX4EK4L+MqIH4kmClUrtit2RzTxyRxorQfPKzEUq90tqXmYOT1iNSeGHS
fNdHWaSrQbTfQgGR7rOESiWoRY9Uxn7w0sQZBwghOpfG81IE8dgIngjT0t2ZzaBr18LRWS+AXYfQ
Oi8IfPRychkclN18qXhEng1YZRibb9eafAVL6meTjlANH4hu+M6zLsiF0cu5WipA2Nt6ElSdXd1A
eaLWNwZJjszAl4tp6vvxEd920QpPqQOT+uLkH2KO1ck/GwjDl7Z89J4vDrOzwNw7qYAuiX+uM795
EV2fPfcZYodwmiEZsHh6Y2+ClccFuXi9jAvFl9mxpQUuFg9d2XrtjWAnDdKEzYNnH+vbGfLMzBmD
0+8KPPBGWBwxOR88UePFvMi3HzxTGLuT0t8+66lqBif9zq8Oa0ljf8LtOYkeANMJcMTVWqTF11YU
LtagK7JhG58nWQjTdLRuoazHl1xOupawZlf/AZNGp46bxVBA0WWyZNTg7Ld6ANAcYe1N5ftiiKzx
hhO+IAx26WeWenwtO6gQMBf+m//Xcx+PmrmJlTGaYZsOY8vmQJCV4AdhUdpPI6DqQPU8xh+1T9rM
T2kQez57EyvnYi1s+KGfLZqifahPTtafxFqgDMz7fj4Ay83FhwuOHvqrhAFFfjs+bFCupoHtdVR7
rwqveOlQmKs/2BHfYzSQfw7BfOrOdkmz8hLxPkJCF01HTsA4BtY1iusLR2FiCiFAgwVAvSGUOxXW
laf3iHSRwKotFVoCItxfDh5edv8XxoVxug3hILR7zjyrIj4Led76UPDhLEdtgX9D2rkUwJkfUIKc
KVTVCPq1LvoiZ5Az5WtxOGM8+WzwvULaeQcW1rFZXI9McKQ8VWAhlmJeXsighWkC4fo4QoNxaOfs
kU29Uiku/t4o3ipPWVJeH0DLIOK6bru70/RZ2qpBppVnXizZlWFyhmR4DQ3sjVzzjeM01oT7lgKx
ISyAyZjfQEtf2o5IVg015aT6OgREKFDuRhkXbucbkg3oWoB1b9PUzJsPLtgaP1laZ749vAEc1F3/
5nrMGbxBdzi+BhBK+7ZqWEQyX5R56jm8fD/PkmmdRVf6omXKD40FWIfjLXvr373jawB2fdPZEuDU
5qfTpxfuNHwbsfsINuvmAp5iMqmx9nMbHOfIJfM084gyoIfGWRvvt/vJ0tUpamdnBQTbOhbIT0rW
cYz6Bq8SeW5WyeXX8oEWQ2g3KZLk7rny9N676qywOjcnp+/XkJBu9XKtP4u6BGcLPDPJw0wLgLbz
0gdgHVtujZbUD/XeWQxAp3EMelZGyH9PzzaDz9MNfOUtYTHul2Ya2gRavwbP2rbEm5BftQeXDdOp
gzqGkYKW6/OOSLxWD0ZZUHoauFVRQhrZs3ytI6+9zUVDO1PZiy5pUxd+KePKmdqXGcR0oZ9L+mY1
XtoLzZCfRwz8tWLeK+2K6TwtBzAC+7XutCq5zFCC71UN/GLYF7mFbrx4hXkYF7HSUyDE8nsepQ1k
ZLPoAeBeDnsFUFSiHm9Bq7hoyNlbYQ18SO//LuHuFB+5+/5Pfm/eKrqlUJE8e9QSDVMLa1NglcRd
+PkhyIqJ5IQW5qMlMVJwgxyEiAW6LnGJ1N49MPIy1jKYt8eOqDK+C592hfbpqEVs9Fzho2p4h4jD
Nr+YjvxPGR2/7Y6aZQfZprLqF1al+A4EMHDD68wBVbrV9UHtTE/kcTHMDKD8Z+QBGuE676JBJ4qU
crC/GcecDLAUEG1TOuZgQvf5gqXowy+Fzvrp5wkrOtLGfgsoz2OO2ENQpHJRh7DxkoMwr6/X2gxz
hnJYqr+V8f/x2vyO4olxV0t/ayuBhdgmWxebkgDJiHd0KU83+ck/E432J4xTVjC7z6Vja7xeIDs1
mmgwgwjSjk+y11/UKoAvPtPOlB/I6oMQ8P9xGJceV7XCLX12WQx8cJsJ0+jF4G0qIQqNdAV2XohR
RvmPIhmPuCXNdSgGWyXqn1VT188T4zUcex3Ge3OKohGL0z1H8BNGmnmbOT9z32MHJBz9nBAjzsDY
c77s5Tjm5j5E1Sh1U68M8MSXh3W8F9S6BKf44nSgQu/WFc14RaLgmOwJ5hFfggAlxVV68zFnT9UA
0xWeP24Ol7I57jJm3sPqFHDrzUHEjylhUlzNm+qvID5oPjmqwGcKDh0a+uIBNSR1qo/qDP4xcXkB
K+zEN4aE7a/ObsLnYGZGjRxa17OGzgNwBTuK1IkEBzACkItwqpg3cwchKsuUKzuOfAfX29TvZYHQ
dnjUHVMIVVtvu1OGC1Qy129J3TfIiqq9xGBzykQi4kcSy3VzdoEu+P4IE+XnTa5klYJv56/ZufMI
hNNIAYncSyhrSOlfJyVC6Y9tdgQkJXTysLAZ3ZtNuvQJUhDuibm38dI7kqDFMwnRf0m/VYWodHe7
eUL7YinDZ36Yi2MC+OOYRe9mO3ZFbP70CBsnQaaj71Xh6gtF3RsIQsBvZP0oWMYPC+ClYeO1ol14
DBricqehpGZPkAndaTW1PIHuu+3X6iZ22Ftu+9BIgtQK+4DFC/ClI1Og9xSWNIF05dSrP5uCNMLU
7LegixGEE6xm5zbEyas+4Uajb34S4uem8A7mRSUVtg4C9jJyafBc+6EdSNC78lChyynq3MFsubtw
wg6j9VKLfnbNnZ/cfWwF1FVs5HU+QvzPIY+4nUvFIoUiwIHwKXmV5iqkB+u01HXoeO9JTcHFvG4I
sgZjOBlxsFKee8EbC+GRilx9uFutcw+KQzS+XhcrD5p5ez0SnpgyXUS1sw2tUpYAqJzqfsDHFjKD
3NhPpeRI3ix4UI9CulvNXBWqK/fhaiG1OEXsZz0tPmTHDq1cQU9ap8sLAOTYz8UcayLBXje8EiYr
1LGqkInR+6LgkgGXWmv1ribw/3bfTRvsti06Goa9O/vsThwCp8z+WPO2x9NKH20HPVzbCK5FFpR3
yjGx6TlXg8vUpB7nTfrtTaFMXc+KUK5Nk3jshUZWDo96TXbef7cG1tBFYR9xkyLX7SmOmatt33Mo
eKg/7VGTnRIN2ZwqLOJgUbPzFwt8YSZyRA9JFOnI7qOnleiiSh6rFz6ayfU7Fx0ujH59KdzepM3x
Xi0UtqUm2RG773cPO78fosj3RWZrB39qE4hN9LAkSxn+iJ1+BvCJIRzd2EVUlk3z7H09qaiJAyNW
unLP0NzAAUS6sJstDO93KKt8akK8QvV2e2eR30URlT8ES1JC4FdqnaZewYrUrhNmeDkfPe5IHFU+
jl92doDWkcdAX6XfTKcCZMs1O5KM9UvEL0lAXPLpyjVsumTbHv1Jc81+J+Q/q21uwGRCxZEsbzFR
WbbSmXai5RO17j1YKcIBDElC0V2QZ45QEfLZ4WyU0iI3THjp8LHm2iWwyk1Rf2bmnDbjmOXjrMWd
HPrrYNsmJKAGxrfHUign3hS5CZmPi1Tvfm8BHcMXx2QnYwnD5/yQNJsSP0/hBaQw7uYT8bMelzDx
OxL7/FzIQPv8EyNZN7/5DF0y3gecaL0knCe6/KRUZbdglcaevsC0GjZRrPqeFT9jgwe5GL9Okb6v
EGe1Sh7e74kkR3dDXZJpSe18uSFBk7tcNZ3KHL6HCJin7noCfNqddg5woW1oia3rAN/JQWjmkNYi
PaOA2vMUgH0gCLN4DCl/w52RCcBnp0+TmGM8AP5WK2DWY0b+0gHiDWHDeboM1rhLIOSnM1WBqU0d
y7YUOCHC1ZL/HWRluIYaZDcyWX/AYqaHKnMLeEm94gPi8iANfE3Kd6/oskDWaUbooxUZN7eGDPkH
KWlRi6xCc1GKj6UDESv2XGfxCJ8iHv3hpV1ltOsD+05OaRO6BYTbmj+RRgHz0Q+/gZ7qP8s3r/Tc
KCXA223wzFf3Dlqhqn8vGVQvOX4FMHjPv9PwB9CxGW9bbZPIgQdF5cqPLPCL3MPE6xEFcI6BYZK+
I4EmmuYxvhuRdc+wOQoHNjV3HdpQUwTsClf8RDdH8kcl/8GEU4FOjNd6KP5JaHtWLWhG+5gTSdTL
atDiCIIKUvHB+fLVaPYvLSyTvM6+PLNLkGFPdDBE0z6nAYutdHFcjwLKIaJbj6e+52lvSuURbFHl
VP6liof2m/BbkGMSBJkTtl5qpoZb2KpGdw9rwLSPZyN3Q3j08mmH+bJHWryUjzWUoNWOGKtXBdr4
Pc1dgMaTZBZp1642ghP3O6sEsuESydNNOxZ8lUIiAXpPwaDvKTPElsMirXm8L7IKmVvKp2+inSrW
IYAA6euuatY69ghxaXKNbO6phVs8ailFuGjrBnwoeOShg7XlTZQ08Vmg1tCAepTJd38or2TcPlvF
uraA1qaTWBsCs50UHSq/WjYrN+Z00QSwA/DlKX9Z7D0gaS57EPz//HTdaHMFjCf8kgC07AfxXdW5
ry/L8UrRyfFWAGwmyoPTFlbbljvGrHiKm8WljRJrBTrEVhHXBZcsrHQbKaWfBJzweLYXk7/Ox3xc
xW0wnYal18gv49YSSjeoqAm+wditpy5HG6tQwHyVJvVZHjnGoUVEpIHFyYoK/rv6hFgOlaCxwaqC
qscZ7eiNNeqTmIrhUKRtSfJjfsuJWT17CnYkn4EPuQFBylXck2jYd4aD7+ky2zFb/o4X2NlCrpBK
EviwA+4/leano7pSsHmIuSJwgpcRbcQHdnfnNNXDZdrS0Ia/idKT875ycF6A3msIvleXOdQl0K+1
k0C1rknN5G9X3ADbmrFxpdqieHsqblrnbga5gSxzq35rT2fGp/koyVDr1ai5cgIVOR5SMKMo9xvO
JElLKoVp3vPznwH6gWNrqs1h8vbqOCPdWfiUAC+DeutQfEQze839HMyY9WBWdzeyQ2opdu2GQirh
C7+GKqrtUBwnJ7U8UPamYavVA2w+IEnBpdjM0QzIbU6bFXRdc9vMq2QWXesw8MXjIWRBkNRyBHds
KZL+Z4hSUHuIIqMdwm1vtCE2BccQ/QuDAa7N+koXx13lxUoYGVh+xn6Z2mFXVIC4Ps8DbKQyQNMe
egAfp9JaCrEunA8iMxLdpeCgyxm7b90lSyFKlcbCy6A53LJGQq9vvxO5gCQX4o6P5r2dZe0yom1c
n6xL4M3MApE5VVP3BRNWAQ7m7IrbTDtiqBlUDz26sdXMKfpbMGwTd3INQWBK8/G7JTN2jrVdaUAy
e9VRNE/7OP3/ykjROAfQmXE+w1Ff0xVeOD/E0lQR6+zSQyGwSTv9iWqwaR+3cPq8ABUQh40jTpmF
SbP5Yt1V5A0zDgXhP2ijjNfSkz/QstgMVV+iMbvqJsrT4lIhwVQ+ifHC+zAcn7wGubpX4FlbmCfh
uV8iQzh/hJ1sFx35TVqgV/K760/v3u0au5buzopN56HffVdwWg4DU84huA2IiqughZy7rqauAcOG
8pwbsogC6mUt7KgK+kWaES3OAeodZIUeGzP7XeOos5GyyW0klU5VTKK14k1NnvIS+lmPCm66ubVf
DtiGZZoortUVA6VkQGkMiCZInLs8meHhxrof/HHh6to5CRjcg0aQjeMjrDPEa3aiYtvvTiU3sah4
WTv3/A8Eh0jT3lMisP8+/LM/OwAXahUewH/pxPT3VrYnB2o9/imIJam8uW7+n3pB4uTHKSIaV0d9
KQQW6MYqh5Qf/piUx7PUg6GFEULRTB0fPSVGVyic75U4seegzsXQdDMoIhF8RMj9QLpkQCn88cBe
KTxnHpx5whClWNLi0l/L2hjVkFIKS7yNjFgT+Eq0JTTREEgO2foN5cBJCGnZqjLBVkdo7oE+gUfr
OjYgbX3Mjy/NB+ixd+AlPNNUDy+kca+Td26ZuYG3zgOkHTucirGa80hl2nS5cu5e+AjToIR5O0/z
SNZFlGI9yu85rrv31wz+U5y2d1bhpW4L7bvZGdyafELTRR/gvL7mE7K2eFvNfoC9MM68qdKU4rjE
cxwcrLP4E3S587eqf8NGlScHnh+doqheIVdHcJT+ljBGIbgg0pNYhjC2mxMq2ZiGUfuou+AmW9ag
7M/24Pf7mG3qx5mwxzHNeBkKIdu/gOnNR5AlVBZpOWmsiOuuKF3qpN3VX6wtQMgTS6+kpaT9HAg6
cZyFeewuzTLwpj88sVRyYU6ZMcEvTEhVCw78hVs8qBeBCPDb+tWeVxaBL7iYppOzqwdxdOoDu8xR
Cx0MJYLygB5LAtKhP9C+BNgvi+rbznvBsFnAVPaInl8CTuPcDqHyWHiFPfTZwCZ+4PaO3YG3qmxr
rAagpydGJ7+u+dWa3coAZUX5s3QJvJcl6CEy6jaOiampcEDH+FgZ01RQFuoz+5XSrZluDymABR7A
tb+EijWHTNXZ8CP2+msQd25BW7eRgi6ACbWoiVHa8BVbpNa5V1LkvaAwVRMr2Ldalm0m2O47DIOX
XiCWqZTKV3MK1LColei75qhfVdGqx7+4n28NqlzQKI8beYLhaylPeHV7niqQCdFqWLEhG3XVF6pY
UULBmyvYqTOMqO04GT1bvsmoYkV/L8P4q3qpODMxx78NfC5s0u55mlcVbcYcFgUE6GHG5X0TvhbO
3ke/fmL9O5m1hnaaQIdrH5Z/yACpDbjcZMvW+jAbzxpW6RKQ87dPixoC5j+1pMqHSDXMCORGVUiP
f7wANbOSxbo4RZT+Rt5J7NPB7YJZRC8WqTPkOPnykuzd4xi1qeBFPFVIcdwXeYVpcervA6IfHV89
/I+FchIjdqozJbD1bsrffbqaPPTaBFZQdJSS2bMPi8Dv5SV6SFCxApur7pQRAN2ZfWEWu+9hNl1J
dz4IVZb1LcC1iskyXyIXq/L4L1htpcV852JHz0TCQNvDakQMr6XbMt4+ugjWRyhDpso1eM3/3nUH
osiy0e2yY+RP3WyrbohjvbKu55Cjj0J/VZ0VNsWroWW2bMbzANrz9Ou0NZ92n7/MMuBBL50OhSK9
QNoJ5BYL2lixSAQrHd/MHA1shzv/qgoM5T1+fJkO45VUiOKsRNOVFVg+6dXH9HipZK5qujfMw3aM
er2ZiuByNNKpFoM5SlJkkhTc37li0vmAH9fVALbWh8WfVjRcx4HDgGC+TjqD34r2OaQ+VPkqyOz1
EfsfrjaTIZlTeBKDzxemSQs0YrlP6j1u3W33OwXj8P9LnEtrJ/bX80msbA9D9q9uTmFBM2YLyF8t
a1jAzrk+iqWqQQZNxsYgs0ISMds7S7lPuXQ/JZ9R/hSjfa9vDozcmKhkOysFbzZ0b93tIVBKOlSW
Mim17O0iA0DeH7xChcX9wuWVfyIgtvKAJisl6jP8xS1seAYBj2y3aUxis1X71eNv5C+qtkyo5s/J
u86TEL9HGPmlObk5AdL4h9JJs/SUcryiY9RIzPi/w0rS4qrjl4no+K10RT9txZcEV+1iIgS3YqSo
eJb/39zzuD4EkV6VfIVuLeLCuQNV7wea83OmOnsn3ogClq6A3ayQrOlH4A4nY8Bxzhb5hkRCjva4
LQVJfqT1WJpDgUjz+byYBswmIRB7d11E4OCvLsHWnSMsxWNLtZVIaYQeBCazmRfMeqDQRfSE+zNe
HDT3FQUFEUhiRQAV+SshW1mDVQXmqFG2/cVcHFPpYbZqIRX8q6JfvvLyTUCam8/kZfVtS5raODMU
3JgRdPAzE3NqG+QI+cJCr3s56UZCm3gUI6rSBWCDRwvAbqkOCPrYbkNqHFWcQJ3YzBGpdzc3Nd3r
OiP0CM3uFpIemc7v7Nh/2XVV6KQ+vK9eJHqvV3oD+me5GtDNQdgqcitbekslvBDByY0kjGQuC4yt
TzydDFhSUuce6DA09placm8GM8Le7omvTRmheBmZbWZJmiRyeCUjXmJKE3VvIUudZPjjkUa+1d4t
tdyPaP+LUbKAwAnMJ+XalsXwF6T7ejgrHkkZg3HPWnuBzwbtKWX27sf+m0PXNf8AAOoskty/L956
I5PhyLiemlC3mBt8LOh25tpKp+hKNGQf71NEwMu5xpuM/aYPGxs8f7jWLGl9//cenRiPeACS5SRZ
cXZ9Eloh6nuKYYqqBj3O9lrBvxoEDU4Dm98LT907vV5xZbikdNdVSV1CN+EZYc8iG7V1PsswVHP8
J5WDqyZpg5PcvinjLecC5qPmuBa1IKr/Lq3PT92n164jdHWb8R/m4vsC34/zIkIQvs5epW1EDjKp
0BrJzBCsLBI3v/nAbrFeK6AOq8UbencikWODVwxa+pdMz0hLO19fCRWlbpZfap01oPvFRlJFYqcH
gBMdqcMGcq7aLJ2lFeou+OSNkdGmTCaYHzNRilO+emUtWCc4uGF/nqZSnRBrofPkGsT+7tjhxK3q
eww6ZipfoFLO6kWMHEjmbh0hdcFaLlWNso7RwSawg8jKW27bGaDgWTuRgXvE4mD04NqI32lI4nHH
heuxWifZpJcHWAlgmN/VMTQ9ZxOlE/xg9w5VKQDMuZQyXJ4Mtk8UFiLhB9CiA2ywK9gC9bLnwfbG
m97BBZG8ph294Ik1fwkylaGYp7uNYN/OZv1gRQTomd2cfspAstTxS0vM6pFkXUUAbNR1R/2ILVcN
qTxwvVU5UoS+Di1OYbaBK19L04dAwN9XHlailLQEmPGiCURDDnve+Jp51ZI0UG3bgk0qs6rpHOBT
+4CQZdKtSoWv4eRRNj12zm393J0JRHBtubTjFlETchNfcWD+nwi/mMBS77SUqWLbU55b0XElcT0V
gqmLhqw/n2fJeX5GSfrcxz+ZHpqJqDOSAgpvcOb8cs0acZ8CMtRqXuqjm7BJYUY1SXah+IeLwcaB
BnmS5BnZG6PhY65d37hZZUh8BZ6ZQjrU1B+GnbJCt3nZ0crRERmViWiVlM6uV6mhrSMNnKTTDQlS
wYDrRdjc5SHcIrfe72k5l/c7YRtx8JQhY/5yzZNQ7F5bxbWDuBuhYsHE2K0EKR0Z2DCLZdu5O3Eu
aNz4JD8RHSWEeHyrcTvk2o85EkovrUM8AK6lOgBeWY0VYnY8rc6YTTW9pTlwyet/90LKQTy+RefN
XOtn/FEMiAuGiUFYudwTVLHBR3C1RrvLtQQcMdjrIhWeuOFzOhQahk7oro7WFyjtPSZ03DRq0A5y
JgmKcUmFpBrP+KepoGrPXM+jubyhhOqyDl15BQFyV8v6Ysb4B7g8knMe6e4LTZ+wDBVw9sSo4JLq
JZIXoR7cv/kP4le0hrzIgClSlTeMPeQojCEmy7y0UNPEAzSfQEiN84HQcMmBm4miqXSzP/wG6PRg
xaIWYH82F4KY3LLWFdPeuBRrkSRP1BOGp2kFaokxi4kW7JFd26o2fsAap4KswN18On9h32yLMAg6
Q0WWocbAhvj9f6+cU8jW1FeT1qgCvfjQvAghI4ua1wGRIuhcfmg9f76CeK4OqE0jwNUvCw68aJFr
3IyQQoRIh9mNHGjpRgJAyB6x5oxtjE08/+Wd5k5doB2Llyeuf6vZ0KmvruNKf5908g0bAfrOv2DF
RWUOk+jyel4Mhb8yKi/t/w0/PPGZXuEF5V/Ht0D+ku2bCpJ01m3vqTuGpA/BcqnDHffTCrWk78gV
fKJKYvEpyWQBVvedu0hatufG55ziGPn7q9IWFB3++aPSjyq8KKs5cXapOQeBXORPr8l2hlwDaDq5
yHshIVtzMb1Usy0Krco9EgRql37yiRutcKG0+/EjNLXjLbaOSR8KArQmlnboXiO82nwhZubWeZmc
rbp6lmbWy3sTHaru0fJwaQit3MIbzA9BmtbB8vpSsoI3DfMO9YPVpi1LWVebGKX6aAAs9t0HpS++
0BAH5sVRj3Ctn0+QEXzoav6iHmu0Tc4uI3gr7NocofRYwJFkPST7gmSlKx9qH4u7+O+b3LrpeVtZ
VDb/ozTUWgqDNpaOX8zR0iM6shbbDJUnGjmQ1Z4BrOeY4db2z68k7zBtPTFn0MjunmqojttuoWsR
3yXHd9jrDP2XQY9hqfLTbcRFUGM0eH3b63QOnw7RODtsVGg0YXsfFlkM81W00x1pd0x6eCyNe7og
Vrz+0nbrmPNTNbcUXUarcfeEorwXiFAvR2maqINdLtr905HwsXpfOvNlWBDvgTs1X1Z7ZNE2dy1/
dJ1bVweUZvQU8q/i1gaCCHL9HX3fS/GSj0hsM8upQ9h0crO5gxQqWJX2Oas4d3kTKI3AHYdcKkku
WhHK6nI+L6/ddGfJoOGmcpl9sXaMuZ3Bfl2as9eA47k3siHOkfDNl4Nkd4CWOR6AT2aMN/mA3t4q
9QpbIhRO6vrCP4mhuqdfpyES03lclG5pxUufTpwxvlFG/aA1GAP/Eelv5GB5AlaNTBbytLrkwT/9
huuSAyz+mfbQBPFRtF03KOCsqkq8C5ifLSn8r3W3mKGY5Pbwg+Dhtg0disRQFjCiCCkKyH2Ccmrh
y7Isr1cfqeDlZ6BKsDspCedfUBQ7Tktn6Ftk7CajN4HBqGNl0SyBfG6Zu9cZ0uAEdTKObKk2SFFF
XgItx+oOkw3b/3IcT8DEAwGQht0qPnNVMf1Uqs8mwyOF/Lgv6TC+u31lVJ6xm6MJEKItTH1MiqRU
AV7XzrSYP71HSM9pZmHpyQ0YI0ghqppDNYXmMEVr004femt5s8e4ci9E6ovGa3PhigpIdDZ236GV
G9Wt5s6M93/aSHuRnVun4f4KFOgqM80sVxd0+ZrZbC+NkiAbylmzSCx69gji2ElbiDJV+KEH3PG9
v19zC4aN5qg+c0xT4uYNGeRP/Vn4qYnkRz62dSDsaubmGOXLfWecWaj3yU/laSOHdZew8lDW2/c7
lY2mMsgeNmQGyxGdPVdErCgWY9OpWrkdy+3BlaUYcQIYdG0XDD1XokMeQ19+NuG7sqdSPTCzc1fD
YLORtmjLivP/B1K3b8gEK7/5l/B5uW4f10qXPpze0HSAfNsJDfAzU8UmrRIX15Cmo3zsY0c1rA9u
UnuU7X9QWxQO7JWlfHqR1Q2Fg+0Gl8oqkjmXvdzXGXVxzKJ4zxmJOsmG1At+QiKd/oWlpEva9LOv
nZ2dlSOzBgKg1PVtHa7t42syCu83J/FWLJA3ujwFpDuVa8ZzcazjdEJD1Dbu0TdRPLCOVnnXaOkB
6QJ0cRSxqrOGjqaRQ6F22ZY1UJNsaZwGjOD4Ba1vWTeTJ1K5/ETCcmaaAuXPrQk7zFYuUWWE42AC
VxbJrnjNpSTKr9kfVgFMMyHOmvQzsfaRs6o3RL+2eoxvBsC/yFUsxDMamVPYgCmq6uje+NMhQ7gm
mnkxbMT1NmjFPSsYKe+K3ZWGp50F9Fnlx+La/1jbmJjXOTbUAxWmYdHLa5RXeBpoB3ojpF3oayMl
S6UFwNizF7G+qXxAAoA4qYpeZnPK4Cxk7tGVm9obYhcCJrFsJroDeSrOtvBr/YR2SVvPdfTaKsYj
v2ViqGL8fRPRG244dZ9vDg7MvEZm3JfdqfMHXE+6PsCZ9GXx5Y0nrgq+MzBzia49K62qCVA5nRNj
HfE0s38Hfz+VrmX63ixpwrzVRZgP1wgBrK9LmVVj+hYt+Thx0DBQDVfiwOpM5npl1SY1FvvRSmLH
XIwEEv/kWKQExIL/F7IM57NS9uYTz5oIpS8Zs4+jG8pXCXomc8eM8ThLoU5SQ66IqbWSWtdghHpm
UbJpmVDUNOFpp0apJ1/WP/Cv/QzDQeQ5VTxEye8jXsiqjLxkoJubMZc2YVwZn/A1wfFQzS0Gwnyf
LXTlAk3mwJaIEqGQcescvFT3fq11hR8aCjCIcpOuxr0oWCsUGRCy0WfvKYP4pHRDnT90j8agxVeh
AsfN8rTNQc/f8Pipy5fENdK78tLklnkkvp4zwKNcXbN+nwbOUMxgF0vBp37iv7L9WTEkcvmMXRFl
zqWL6KmiZh/PvW6gavR4EoX/uAJaflC7Cnf3aLP3dQfDCDEvzKmxaFTD+wnz+V6ulSOQTNNHMKwQ
qK+GuFIQByuI0AlTGH0lPrTbA6eo+StwHdVlZO5FAFDo56YYWLY1jLRWxsHYumMDAhf8eSWGBDNq
UjuOKaxRHiG5kMlBFaNeNTokflyzpjN4vEO0RIdSziZXkrLdEjaLfg3/cAqT9b/bb1Gw0cCeqz/Q
wkZT3ssO9P7+rLmGXKJxGBnZX5AxgtGK4wFLOOaYqc1Vr6DGH3zHMR1VdGBYu9E55Jv7gf7ipNy3
gfLaD0vO3lfWOTR3H3w+LWF3T6ihTYEgiFNz5bTTT1hb4eLVVYpDxNRvB93tM5CaMQswUFOFNAoo
Vw/SmtO7vhEqkADmiiGFwkv5Q5IJKUGMdeXWBYzMt9g7QLgu/bF9gOKkiy2Gb6HNNeSLSKeOspUZ
nkNB0N/FWg353rfTx6SCJZOySWxXW0/MoNkbyQQr+pHSCSlK6s8PaoRHKfeb/L0T08d1UcSoWBF1
qGXb9Jlw3KmosE5dLtDcCrzyJF/ZHDtzzesFJr5wD5ilvTqUY77ov9iU93Ic2u0/c22E0yUKrLZB
Zc93IGpx60N4L+58GKRcZA+tSOSEK8jmBmgzP9fAMOHJLW9/DNxInLYMyDITwyUWP3hmjo65jBIr
s9y/ZK28tG0Isu3dD+kxWmwxip6wr+lWsbcVTFTWR5a6nOeeqLqckQbE3AfhSUEw5S79wZH2UYHr
29MpMmt7tSEbHMrs4ocYwqxLrpeHAD/ob6EEIEcyPuvQVdFvdQ+zrmnstD08dAvmUo+NU80Z5dWN
iSZ77r1RqcbqYUQ4GG9BlWdGaXPrc0H0kujmo39zATjmCcBzHBnQyNjDNWuThFp1kHXMFLPvPNy4
CTsswurgWX8pzlZyvyvx4wzqkdvrPikfuQ8L6El3oi3RxV4RuP5NpsFTNR6gqHTKmXiAr152WQ0p
y6gH9MMEjM4xcBclIHN42X57t+iY0yvPvc6eGkplY8jekwR/N9qDiC698GEAPQcqehOY5Ue5qZ+x
+Vnr0Od8gZ64h0pFRPr98RgJGH0U53Xcl8o5Pyq3uIOXX7D7DpDJm5Gjtl1cNPZD6JjL3gH7AiDf
pa48fekWy+p9hjaJm/1VWCSloSIkWBnm6GawPHx4tZrpUWy3I7mgTE4yhoIaqvbNQnS2ktMt8Lms
2ht5+JPcA7WH3A+cJGyzjvH7rpdoPs47JGo+9dHEB2EJ0patvUd75YXpDnwhOXV6UeMttVLSoX3e
HFGFxySfEqbcqQj8mHx8CANRu2fMH+qn+Cwse6p60uATu7fGDr4Mfg8Vn9kSryYqSNHjeALzFKQG
t1nUowqgLDfK5OrgeVj/4orGzwn6oGIFyQFhL+FcPrU8ipWz/Ck1Bbal/LQzPqm0BwNYRoRHVG0F
I/50pcCftrKMTkarrig3n/3KP7gCi6mlUUk/wvaRNCljmKOAxR6XnoYuZkqsjJnnHZlrLaoc4fEd
XWxsbGyfRMKa/IdkwJk7Ijhgc/eVjCTkHaHE8IpRtEijvEAgUfK9rPXC2dFcPzBhL4TeLsNXQm+r
UM28WrKmWC8lbqJKKWh3OwF3h+CQj5+4Yz7QN2VWyjenBCSJ9hlF8sNoyJQ3SlKBHVvBBHqV7r9W
OVeQTJZ/WKNoGRgwvgDbGB6WFWhFGPtaY6dSNvyx9cu1VM6Ea3DSm8EICVA+ea31IgzsVQLwbk3v
AkTcEV1EpxqQuIn9Su5xiU4o+KwKlxjfwsuktiiACajYD3Kw0twzKosCIf8aKAPP2trjbi+7dWtm
IpkbgxOGlJrHFtYFfeD5zH7XBugGRaPJlyw6fnNipOCQ9POPERsn7PS77TklM5inAogfjP160215
yHlm3J2HwQ2HWkkmgG4a5N+JT4Cwd5gRSC3/BPC2WaC1js956f5iSG90i/fwguHdVJW00NKyNGr6
VjNX8x5C2Gkg/7u+Z2Xdt3N8n1ALzkIiJ7rHtRKV5k0eVuLOOwymh+QWVYHEaeQC18ptdBu358Da
4L1tvHOBjz7GPudGYdGplrQJmbBdQMrWrms1apj0HkV+kAgkTSJHOKjuJGGq5asfOl4PIpPD03NY
X2VdbVd3O5xTLRPoyyt5qlfCeZDVKmF9KLXmqgjbqaLywofopjpH8p9xopPWBF5Sebxm26+o3uAE
JGId7PHYL7ifFCxnwG2NgMQu+m0mNFTgNpvWa5xUtEyiJaN4ngPGdTwCY3NICs6iwmOswT/SvoAZ
chgbLV7Q1W/CwQhyl5Qf3GVGWQ4T5kQyqu5qjdYwwfRP6+pY4I45vgyjXx+T33u8j7Bx+5xJ30Lg
GVXTV2V6ohW36wgLivRyifZyTsVuq8nvOCMmKiGNxwb/5YjVyVE5ij1WKsJwuB5IQoFUJt0Ph6Jw
h2noyGWO6aFJG1IhnxnFACB3R8TKMt5i0PiXza9+S+CYlgkj8+ZHRrqZ/IxMnYAm+fn1dlTaibQy
R57Yv1XoE/SV4wboHDgWaV7PdRHhDsc3LQeHwTS1E4W/raCdzwto5g6OvECdyk1jQlCkCOMWtj1W
0TeYaLfFkPY4x1kCqFQfGo2z0zVEs4HxJCcsuecTPpWvkboo65XGW1esdza7u1082UdMJ1LAT0aF
iLvyVoaBJ+kq1A7iN6B4tB+km6oDg68clvfWvG7GDm+6iJM8OlUn/854NRLp33letmDaWGP5AoWd
UIqYaozCdoAaQZ9dgGpVvPHUjfVgTQ7Mv5FrBQoDJxvMQD4mFv8fHL6cVodYlbu4EoYdlB3yv9tW
fXBat1FrrAD7c6GeD3NL7YILbptSuvGCEUdVQP26dIn5iJ4sJ2oCdox8xyz0LBPuC2HnVynQ6EBA
aOUvCUz1oFaV7yDA+N6IHYfhap4WDCH04uin7sJpX2t3+pVexCWHHXFBbAZCnMDGbU0Ekyyc1Iq3
IlW1EKdzPttQZWNOHQJBxv2e0sjQdDSwfho2iYA45eAOUFI1FUVqYYgrw4ucmkxmx3bnLzJnBVez
+6AJymy0zc8tPg3DjYRtBcfYtu3y6QcXnfY1Q8MhH0FCsbqlZtJH6rnIsbfwxyYC1WvCZWA7eeVB
BQGYh3bfnK4zukgBOBTJkiOqNnpQUt7H8s5aLGjou8x4V+OozZyKajJtyXuaoAGPRpWi2hXXjF/F
XNe2JrOathSv3TV4+3ki5Z+31HTnqlSfRNiyWRZ2QxuXGFE6BRNTAm+bgZinRMMSaHDtp60bRcdd
QG0ZiBnyg7/Mm0BQHVSRYDTnqcTHK1cfPBQrZ97EC/TnqWqyb4wzPv+jS29cGrIlVFxFX0LaWIZJ
q5S7VYe6OofSuxfb44U0xy8azl7SVao1ELK+pzNb8HRe/0/Xzpit+bJZWadwwp6/v9uOo096out2
OQ0UcXYo+a+MpvSGU0yxaMDPdSMsk1lInV2UBBuq2fBw0RLAGo81ueIXPwbUth9QSOOuLtx3uqsZ
zTTWVXr7r/TZzJQfnj94s9Hk2Ilxb6RiLqbecZ12WN6e2+J8YyUYMqbbkTwF/MHan6JE7LR8XQNs
/1yltwIGsK71Uf2Vd3iZsMQmyfjtqikCch5kuRxKnGekg1dCg1JboYfi8yCzP/TqHaao9E+fiXDa
+rwdFP4kQ2LPNldagCJWi05hWrMF63ch4g7eNuD/4BmgDPoedWnqNYVbOKLeXy6PisRUI8AeIdJS
Kuu1Eb27a8MbW+G05dYA8k1x+e/zaeZBdu0mMSRL4efUhPZpAXTnZ4A/o58N8lGdf8X0OTJTZICO
4qqFAjFaFKLfAHRBqKWxzZLlEjmQIOtEOPn11ZKB8CFwjdqWtX6GA1jtC1ZcY1KYs1QdiLs1+UDY
8qG2b4kEFhxnSMD5hJKrgN3XREOE/k+XELdh49yLzPAPCkBw7imaSC8ENe72a3FTuDVmMVATqUyq
hzS1C+BFjMSfRHxcTrqQYFxrYtF6MKbzkrP2c5EQhqw1fK25T/CbFEaYREty+v3gvLV89e3ef92T
BLBJgcXmqxIgKo06h45A+ZfRTvIBhu6uUt8bSb46QR7Qm/zIuiAHRrg3NquD3r512iO7IQum3Rms
HHUsOpefiMkZg7ESdJm1vp+d2GxZ6qKCQTrLhuBFI6yB/y0yIH9kqd7MHMDxXzuFAKLZC+3rSgml
SpDCT5ZivJK520FPswyFZaWLoxCrzD0TVVF0kck/7znfEWsle7YbfZenQexJ00kDwM2G+HzWqEiQ
jQKc8JyGurmWpFnwD2mDUXakntXS4dJDQSVSl2b0XXbwuPavW2fglICDb8Ha86PMNYwvg5cX61L7
SZRteCLaiEWhI5ag6cRi2S9qFRIaaaZ/c49Xx/At5P0mOeBPg1fBkeUEkpRG8nUyqlHBAfU2fw+i
fanL1N2ZMv0RU8wi/GE0gxzqKFBhNSJ/7i47tSAYDJ85O4QE+Lsn0CR026DwXQPEUH2cDc2W4+F7
v9qTuphUnlCF44KFdAIgmHTOi7Vb9aQtJ0FMt2kPyyVuJSVfU8YrD0nJEx/dRO0mgbO/Svii0f91
c79O4KBCe6Lsk9fci9S+BAB5oYTdMKxE2pkG97f/pt1m1v56v2qCzQFveBNZ4pXhZZNErkpK4+ZR
4xgczBg6o9F47LxzirasI180OZIZIPUcd0yFlHzNJQBgiqIS7pk+CsGbn8UXoZvljRCtsUJxPjA7
8snshImF8D7s7ZlBDryp2ITb8laX9B8X8uBQpj15u6XYmMqbvZPHaXxczNZ5gqBm2a6AJulkjtGs
DhnlcCNaKxyYoT14Z/nGIleZ/2C97McOkYZr0vyPxroNEF4OVptGIowYyYlGx4eGdgEfAETzf2zB
HCIFxYNh73dCoYXEkdar7ejUbH+lzeLgKvKLvXTC6+IK1F9IdSEgXkIjHM/bVwD6vNSP9FOesxpY
Ca+5GiYATNo+oC32gxHCQ2mgad1e0mQqK8aKcxtzuWeMjV6rkgmRmJ785IWoJsy56ZUoHWWtLwnt
VRcnGlCFtFVllepOXQiPha7jcDCbnzH/jMiFDUdD8cEX8zPjCLJ0wOuqxUI+ZC6Lc+qD5F4tT/HV
7bVvprRuNlHGaYiY1fjAxH8cNJaY30PdCSw+HS2cIBRmHEeB9bV778ZPVap1uwD4LuYbNW32zU1U
9Knefps1K97i9b4+hpaWggIQ/uTHBfe04f7ILi7onIfDXlZDDU/Qe8WBBsCed58BqJpJtoe1ZYor
6knxw+zatvE9oMAZM65NnXJRaE5zACZB7OnEE8fMMDf7oxS/uPZMQXc5grAs7VUZ5JI5IQYUcDGG
R8Z2qNm1XzvCEX1druuS6Dhj2vD3GtndsgCIy4porRUJaOeLM8ESJ21Af1qB4T37G4c/Dteialsv
FReh4yXG9yuHyM4a0koToggeoKgI1sHKKUeB/u/MOFsRkwqpm6KoNWFCw+xpA9QvNzyfSq4GT6nN
d9U2gTUBkpIkKiRGaT4pEod0fLQ2VRQ+OKnHc17femh3LXXC2PieW/Swza1I4O7KKIajfNelOEJG
o3CXsPDU8/YTMrFfUDtiLvQ/zXZzDKD69L2hDsON1Cqn9BFvSabMaBXf3AGt8a6FPg7MXHY9AuJP
aNM6+AkZE5R1PKbTROyfMD53MoTWPztnUYTvO1/1m+q4qHgp+xrhzyMdpa+2CWsyxMEmZEY75j4X
m8aYZK72TQ9XIB4/fJDe468TO/w96zFVwnMPBkZkKRjmRZXXe/37mds4yX9nrZgzsda8xs0NNvuC
Ijd3v4FjvCw7O+DKrl1MPASPijUQfekxbMgvWiWwxdqSo3GBco+K3PeuC8GADKfo/QNRUUw/7Rwp
LKFYmcQiE1ulq+bzRaJt5ACq0O88+5ec7KeJa1y5jFgmhLMzdZo/ypdf6LNMbo9iumeHwYoXElZx
umWnnpw1ZwuJIuIRrkZnXS5IuKsbaAI9FHh6PfeYhBYsF/UvSWKgqUw+VDyPk2YYs4emPvtJ79+m
4JPCizcr4YsZX1P7/a+mMspvDnhpEAWsY6zcHBrfnG2oRdG5ANHA++gLnSH0sGJj8KkRS+vHGlUM
2PaGx+rR1SuK6hODr73wWW3fV0C6Co9+sCanIZZt7kPKmNcHLYwcHF/zttuGCxV1wy5baEnTatxM
FTqpX8aoEKmaDaw3gDJ9YlixDzkf1F3fwqT5Hyia4BSSTORgTi46Ylf7paEwF8/ufJ7IS4iS706r
vevJcJ802wBMjS/Ft0K6z4Q9ooZHJUL6aKaNnfGmIMZkJUUwZOBUgpTOvsAk0Ld9BxmF0+rZB/Ws
HSE2TesydzSI7iNQ5vRSexCeHxShQl/g8qwh3a/tLfz4QSRCWu4FJHLZ4qFIyxRopyJjVVmqiRam
Pdi4BUUqfca4q1gyw3j3j43rOjecQKUI5yToOj5eaqYmgdza/6bl20Dyuqk4s6h4ZO5b/aoUNwMC
f84deyRNDqtahIhvBEdha0NFwTNoe/mE8s4MZnQ3D896+xTmO6sD9MMrVMM+XZgrNqD69iI5Yupf
Mu+FFG9wTYCBA44fJzBIxr41UENbBzHLwoILoTR0qhZR66Y/sN6ivvSAnqglWqAZtgeaBF+UXrtF
AGRy45dwhtrTQJOwnK6SYzIjo1Sv2P/AtLmP0TFTuC4PH1sFtPKfNgdAumArbHJnhqIiLROF3J8E
LU+RYyUITvmswbFXuqHlfW6C1voMFaAozoLp/v3tdXUw2rKdRwW522JQwuDhkSx63kDMtp2t7nUM
p8bg8IGjA/NlgV8iidNC+Fy51IZiYiQrUKluvpGrUHozwTFm6jM7f7ZbFcH7gynSGntikZ4I13DK
ixvAymVEGWAQGT4GX69PH1RVqeqttn9CRNantWM1VJheFacI2gwz9x645ejk7XSHN3FGnq778ufa
+a/FRwOp15Xvzxevkq1Txxt5b/YSybaSaZicTZoKzyqBBv30wP7MbSHDChvweLAUN+qGqbV3wbcX
CB2rzwxPAGjQhxpP3pcdiLbQMXqT41hTt4c+4K7abqwWVc4HCJQ6FCzmTVM8a2GfldLVL6sjMPD0
wGjYlPcnUZbqCk/Y7BisVCZNaJ31LF5HbXnqLdKuC6p87pq6uIEmNcDcvv3FfTlsZc/yyS62znnh
IPl5Gxq6X5N6t9BMwGMocIVw+mWx/XXkCq7qMzwFuAZTGTXPPr1Z/fmYl9zAkDqp+sqEEUPpOQ6s
Ydoqhf+6zcxmTZMPWYAQ+G4SyOueLMbka2mxmFQmGQDQsJr6DqSIxmDmty0KWEp3N/MSVjRAHRqc
PhOdT8g3mOJ6zV1IRtDnbeOehYKH5A+uL2E8ARFCInacpjNORkW92/mA2jJ6AAHY1UfAeaNYBn3f
Su33HaXfMsrF0Wu+mJh1oT45Q04tYf4ltqadTZrEIQ9UmkDafOkQPzrx0pcFp+FJbnAF1HWbDFKz
c134m8eXVWQW32M0K0upg1/j07wsnq5CtAqEyCyTvSIsRU1ra3IKtOJlKMEv+NqpDMzgf1wChrda
IoWlzF0BTmaOHm20VotCZTVOESho6h2N1fh+ePvJny0vPFioPQ7fw3SQiiHLFTSoG4pB7SHVSwaO
1CdFWO5Tm0Bi2UK9lXQ1KfSptCeWk96maWM07pKPwU/FO9i8fkPVZW4Dxb2uSw158rSB47SHq9dJ
96H+q+BJSO/HXM19Z/sFpJXboyPAfEGXcln2/8b5OfldGaBRE93OHxLukhiS/udmNu28SfLH+m/C
/thShrnzTQsrV6dOa1PBSuN1Yu94CCbYpDppSCgbHBLb0tNeXn1PZPZ3TD+FT99gerAkFjZraU75
xBMAPzyZLclFkk6HK2AKrlVHxQKZfemWbt3bCjMk3uRMh7SJHvg00ROmK//XF9I+jg0tz9rUxJ91
CbFrmPfMT70K/Y6p2JHR9x92VjsmFGZqf9zeXr6FXSjFQsS7eXePdzOndYExv8mKkYidUK8kE4D0
yUhA6dJZKP2m9AuWk+dQ1M6DiZh2oJ3PTeeT5qH46m/+mXCjQrhGJvLrQi6sabxRwSPqUzmt4Tlh
5dp8OywEsC3ukx+3gGRGuYZPR+jGHMzyBMrTpJO55LoRy+AQgq22T4lnOSYmeA2zKr4WCtQjn7MK
03zFCWc3g3Hw9DE3GLp9FkpQMMZS6V8czaNZuDk4gRGS3Dft/E0z7QOPLNb+Gcjsj+i7gcL8yMq9
Mu3DOJ3+YshFtFuFw4xhY1KRFhQmv95npQo1w/jJQ84c6RVwTmtiBaBtr3TWB2tjcwDmkG53QnaQ
6tYC9OR8alf3lx3Lwxrp1d/VCg92Ui3a3FJfRdtF6M6b1OjNO+bI1r1W+byi6qTjDyRosaa4ZuzE
AB7+446csjLY5YWuD33Cmq5d1iKfkB9wwEA0dRYJSaYuS5Z61Vynia6rnOHn8+X4xfIlc+16jhPR
3DiS8sxJ8jzQkF09x9Ysja5fzJY5lZsD4e6Q4UDxm6AEVhUWWYtBUPB3wYDjZqhpYa5eAZOvbga6
m8BGvglZyWuBgZibGNSGclnU2fXD24xq0NhBCLA27iX2BxqM6g2HHUz3BOIOBUOR7amsjwX2CEpz
2NAuyNLtTVh3weFgo25SFjwsU3fcGIvL3PcLsCCEiXCbW/VTPEHgHlJrURhJzo3nn0Y+fd15S4pi
8oN90v9Rbh4bQ+oqVlsnYqIvT+5BebyT7uf7JrVgg3Bm8hCfL9iCYTWV417I7GUw+9kOjMMewfcE
ZxgAO6XqCVhw8WLv/RNSidgnOMmVo4+AtLOExZABjTadlXQqnvcKxzWBT303ocMeg63kp0V21ys7
4KvlLKZ3FNMHEPrPv9w+5Rb0rQZOaYTuuqFfI9ISAz0nGRU0r+fsuRIqfCUOPFY3L5VWqhP3u2Mu
CVchBxGgf8K8/DQW+Ih1n5AkWTLfXM4AG7ap7iuIpuBh+Y0jA8K9+m7eyVCZLb/Ec7b7Y+vPgB9d
iSnM5Uq4aMZzznOjPHgn8fOEyk1lkXeCXbN8B/x49JjAmKtgsAUCRgiJ/ghBjLQgeyVYKLIOmgTN
/Y/YptyQFXgen0Z3vClgdqmUZomp0IUS4P4A0y8nF6w4yYQVCDTAaGDgeaAVsawUQSrLAlpLx2r7
RkXLvV4hZ1FSbnz2q5N2I3DeaVlL+9zro0jitOgcYLOE+yHlKBhqUGeqLi2PaPmrzx7Gtwbq0gCV
WxoFOL8G/fdKEYPt5K+dabnLt/tKUX3gCOI70r1yLo0oa5qvNqQdVgv1/J7RmKCNipR3RJArMWgM
oLbi8dThFMz3p2JVpiE5FCgruf3D9QdxA1+AdelUiR/QBmME00RsUwVysClii1xWv1U9sbvSnozn
eMcATONIMGMkWS5koA+y/qORdi07sNmysdZ5D0UCU1W5Tb3cKpES2olFs+quqS32ML5m435uYBxb
Ql1GZ4HEf+1TUSjnetRoQI2R8TdBncWaVVMpowJqvRAq5GTrGDD30mJ5BLRzPj4hrDBm+yQIPdUj
yt+fzFE4ON5fzwaGhUN08sJCC3TMW67Cm8/dESnDUGFG5PtbrLPyh6IvVY+IZiBKLU8krErecFJQ
1eSj1xHuf1ACiqce+N9kDUlriIeDukUCIyZRyZFPD90oeadfd7g3QqMAslUDnmKKd02Efo9FP55R
iKG8JSTRltpX2mYOqZ1FSkwhMbls/0pWkQWet8O2cPOI2Bna+JZkPDnALwkxOT7aTw7pEQi11EDA
N9Rv6Bgfm/M5DdTsMtdZSq5a5VyFyffwhynaCZuEDMQrMO2O98omhwqtzuDyHdnwtvIEViMJdYgu
E8KjsNJcOCokdH72HZ1jLpSZftzyaDya03FgnedTk2ZR7Vf+gt3BHbp1H5/LBvsGH3XlwsDnZfVh
xPsv9t2H5AWOHhQJUqaGUZnTn9Vbc4r33kEyTZRlcQE77LDM0xaAbEFY7Ie3GDlOphzSesGKu2NP
geUnUMJIi6JbxOVwocp0QjqRNAbva7PML2Ns5xF6cG6rRhD7l2YnqFjfkd4+ffbkmK4iL1wh8kwT
GyBJnh07R0awVlgmuILRc9D7pzAt9Bl3+cGUNuPfSIU2CoUe+UB1vzfahY4AxvXrBoiPJKAGn0tT
LOi0lG21tpdi20/oeGKku2138JSC4vmbzgI3jAkYxuRg9WmBPXt3THcpDaijVbNhLq5Apa9y3ugU
Q6BlY5iP7E2cdns3aeE5GeuUtTy8XB75Jk2uoyXHCG+g2AakrIOIQTtWy3+nwEYB7Sk2vcjs+s1B
wLakKBEvRiZZoVdyNBKBd86H6LwOquINzmEi66/sHjZXT/dsvDt9vBof56lmRzNRUnqbV9J7uGNg
62YjKmybbevG2OOoYGRuQhj/voaaFLIZne0Pe0HaW+88LK0BDB+RbiA2FnQzXxySL64q08Mutm9L
doUc6cHnuB9iWSMujx6xs/oqi8xp1JX7BwZjSnUzpEVrvq7atLgqFex8DV6Rl71N1zj0raLmktsB
ntB4NADeQfYBmvNy3H16jZh6xkSvAc1c6mXCDHlSe6Xq41bIMxM7GzQxmi9rRPbWxENxLBc9hTfS
uVMAV1K3PQXrrNQU/kxMn3rrXJcIsv0r2UM+k0T+N2iv4LDiWNy/2bWnIU4WHXz4wAoV6vOGRIv4
TqSB46aZN3A90d3N4LlsUT/pldP6q8yWbzmGfyD2ZbXcz6jbnUAgKfE4HD5h6WTHdKDBdUw5Mg8T
9/Adw82w4B+pp6OVvk8q1VbIL/19E6qeIrfiQnZmPI6MgEfulIQozicBdUFsApI8cO+GWCoMkN0s
HoDMXcq5dHs1t530g2GdCFH6Zv0eWxuVh3jiYHMxXt5jzHYStuBxX2vKyF1ThYRp5JWIofd6RaOO
LEnCC5xDjvl1dCX14x5sXdMpg1pMHJOPuiA/td7goT+Ft73WARflisTEES0E9UZ9DrxebZidmR/A
yv4VT+1CViz9lA5H/eEFT/W3rW+Lc+UvSCzrvRtjfclWs4QMytd2NN9yQmNyFTcPuYd51ba6NiY9
PTx5NoqCZLQEJBP8IugSCJ7B8LIC9tyZP9rZzQ4U0DeMfymPueIE6EKalA+K6rI3QXbaKqI/QyQg
1mfyyO9m0j7H9tI+IaS8qP/myfO0k4Ao9lvot+Hrf40bnLgHxsloIplXD4P9qxy0b9GVKSriOW8k
bmiqjlV6PKJbAVwC9eYxvuN63qiNhm+OIzkyLPtzCjSfBFciFeUl9dIY/kdRZqjYDP84pRratO8K
oj6ncfbhXA845IcvHeV2Zqf5ScKI8ob7sIJHRtStZC//KgA6Ntr+8qzddJQnfjJUnRgpJcWnUouW
BxuZRhBMWnqdhA4X8O77iiJLwDYRiTazDtgrdoONnYqdxhFd6aEk2/5VHBelN8YXrsV1LiJaT7bW
cOHEyx9R0f7fkYNyetWga4A3h/+mvbYccSK1hWDSxxamvIfW/NmOjqt5msbIxnvs8g+GdMVhwJES
aVu3lsjolZUM1lmlkbdHx5i9mKZYzgbjA4JilYoAz0WCiVTjGGWAAR9MzSif2y9Au7cCLXOujI0f
eXk0K3yOM1IieZycPv4Wjazl1bxdqIu5ma+X4ummihmGMYv3ncOlw70FC8LutNr1QgMtPaP5BxhX
DuZ9aR6+81gqO62zU+PR6t1IjRnAdbl7wTTBsetMQFt+lhKczzhGwQ0exTChgUEp6fLAr/+AYUyD
bV2g7YzYY+gtPRcSE1bZHl6QFVdGjDxBgRf3GyIxOadLN1hmo1QndT5BOqZfHP2iz6T/pWVLCtNq
Q/bsO78sv8IQpm9CtUoELMX4/ymkIncj26YQ1IBqooxPKc4Cbe2NwiK7LQALa5y86a9ciWerZY0+
Y4mKrFyOAt0TZhN+G4Vw7J5m2O2nFizBJ1LqIFGcVxOgHyU0wBbl3Z1aH1LHGLP1X1JhKu9ui9g9
Uki8NJM9LsLipd0r4quSjmywA1csSQrJUrSxOOkejJSMGyRHrJYIu5Arr7hew2hG1fx0UH5AV/zb
VcSWHU3tTZt7Iv0xNVcEU6za9gX8Q6zXmyh5SWICJli/5anKLpYaq3g2JqKpRS/MpoVirZbk/luv
J75xPTtr/wZ0X5c57OFBSGC5DVw9Syh1rUOwE9N4lCR4x85TBZzlvg2bgRgIMZ6RosSbyY08Js0+
iGtbeux1hBHuo4mqR3yDmMjFhuExrndwVHa6uNZvgZy5WamiDvzRj4fKqSEAW2uxlLzmGIc0lfSn
JXbjPDUF9le98R8LYYN6DikUwZnMZUNDc+mKp3qxJmJPYxW3ppYhUhzZL4+d0TvAGTOB6Egyr/t7
nCftWsSmo4YtOnW7Kcf4l7laYPgBtwjIVaJm0gr8F231tIQMCo38Y26xGau4xXX7L/P5F9eUsDaK
KnmWY43Nys7DZkDDc+CkYIULYUxKGZaHRix2h/LxoAw7hy5CNsr5MGQhnBV4k5fm/QwL6MqjRu1M
zKAdbghPXYOibR+c8qYX2HZ34n+qXutnrfyUQFGnxhYH/KohZ3KcXKf7JHys1q6qjpcxvKS/yNw0
yA7oTzal3+MomkF6a5Bwa/NqEr5e7x0v6NAQCOSMkBj0Ufi85YeZDEZbCGwBkKzXVXpY3QL4Y5FU
tUMMPLl3ymfdEoqakVMHKpYuD0OD3j3FYTM+wHLwA5X4rqSYJNTor4oy6c6RiE9wccpbEej0He0Q
//U03mX7nzSctGqulHJTvAdX2MUqep7FqMvw8fdA1XUJnzJY3om6MjHeOSz5xGowPuma+0IH4ExH
EJGZpa5Ag71ztCEF/7DWlzNfcIhuGEk+a4jtlaHVxm5JWNvb0zJkmj4EFBeumkqkdN2/9A55SACX
ydYQ2pyU904ZmOtb5Naot8hFRa8N3vUG62TtSCXemtBJoD9wIqHWYCuEpCoYE148s0VZw8WBekHV
MLFB8ETDWrWnuSYlSXPUgEt4LrfRGaQ8l1cSV8YOK7/jIuqWrorxBqLzfX3cSgyHlhVPr2kJdIvm
3qAiMr3t3Md1bRu3NC8ihUvjG4TXWnZFBY2Oc2T5Urq08OjJe0easnqlm4xgc18O2V3ZytRMycV1
KxC39k6JRhNmgwk+5jZQliYBJr55j/F7EbT1jzVz29PdOrFfiydwLYDyDPRiGZASC7DxxvX+X1JQ
RNj1mX5j2QbhxWVifsyacUOrOZz/2yfTjONlSx3xiJMx+Bz4NZ40Rt29pok969+W01d5eOYSomYW
dMYAHUDDeIR03Z1DdVE7z3mAy0V0x4evEOzbQNBREJuYGxkxyidTwWOMpBJ6dAexEPl/x/YLMnlY
jfV/59eHqtd0/t57jTlA0qL+y9harrlNuq+r9lV1iLY0W0l3uRPx8ek0QcoM5X5EkxJnZ7lqsSZ/
f72El7aF+MAFe8E81I4gijOgYYjLywy19VAep42M9kG9jh8TarJowG/v05NngOOjtXB3zf61buPe
fogtSrnY83lv5OXdAslRrOJJgWKwAqPAizO+Pjne5xjRaCTm3tIAWXTtfb/KFQhOR94yjONzpoxj
VQGUnpiH7bGxLXByE6oAxbwLx0w4iT/5NyFY9LUUjaNsCViU5xKunKoZGA6OarcRdXi40uIKPamM
Qt+Q6iigPaj5sSgtypelOCA5dDHrqA9QJXyxhQIz04W67bSoChEvnjY2c00XWHNxKQMLl+EbDIhr
obPNE+VL+BwgWrk+KcYu7d3ZIY9kJ+nyq1E74a6BvfQTne8kSHfwyF29oI2duDX5s5uZKN2G0hi+
HZxYW6x8GrAWU5zViG6Oq2+6649ZXh7t0I96avoEpNlV+JFRPNAXxuIjPJ9/elzBAGsgeYbaWe5Z
qbI+x9qFKBVkre1WkYhHhNDHUP8mS8k8a0lqDjfLNC/lF644PmogHyt6sgAr1MXqo0Gxn9m7Z8bu
irA3RAuWsuA8DwppI1db8yyml+hiZVJkrl0rNeVtrMeCHXFc16phEacliUIXlgsSA29BpCrGToHj
z9RRAGX4jx66icNsAnPzHgWMGzjryS3lRQ9Wy/GyNO8Ze1iukLgeypM/PPSruUNJqMQ6zvQlWXYM
N7jwRrB11Ox5Y5tAiDfuZrhd7kRFvA1m4ERyyBRVD6q3CqetHXJVl+wsngrMKZTNnqyNgw2w42Ep
xH17vmzmEEDPxWJjtq/y+6NLijctBZG3gXp1kAVOHO37qpZhOg3sh5emZgCktVIEb0qd/SruIfCe
NMZJp5wOTKo57/yOIUjyfg5Ko+QPFj2JO1qr6rXKc4ADR75LqVbR4hjBPOHQ3ucIuk3sbfUj9+aV
Y40Qb+IcC8u/UMowzoiqFdfb/PJueOFIXSiBFDAprN2BDYQIgPojwHmpSrZFIj+RF37f6TUyo3HP
KHtWcIKHzfzXhy/0iuTWg8c7aojKWmW0fXXAzuIAVpOubhlYro/hSOi8UZptqBemUSoX3hhn4O7K
a+hJc94I5lQtFWrVVaQKhEYtNbpGWLy+xwJMIYN8efylC1Q9xHqfoxszkaelJrE826d7iEcwCSKk
E4n5oUsAmEcDNniDWsSkHudF4KU8DMvtRTFhWAlngVSk+rx8MMLi+eicjjCK140fC5A7WuzOn99r
Zdg98ahL/s7MaztiLPQfJoIhwKKBD4TduJd4bAZ9wkI8Q8+s6Gxs+yjVhk5flMFvA6hLOTJDc7qS
VSb2Mgb6VjR9l3VMmDtmFPzzamoSul/gq1A4Cx8TLYOc4t4qAeYn3HctdzjmkfZNQ+0I4eXi5Ifg
bp1tmEr3+CDAP8AjDkqyMfqVSga02TTYurHfj4XeL5hEnKeCRHMGemy5AqWo0bLQEW+ugGy6Vc1R
zifybEPpUOWJNXjQOK+JOSXuSOJotpIKxGYEOBN26DQI5hx1xShqfp+7tuofF0OTUzALW1m1i6iM
J9PWmOx9ZAlmpXh0CWyuI0VAuSXhxO0OFyWnI3d5jgqdWgkXq9zY4COAlVu7XECZ1+OGCcbSgkVC
vRx3WQCwQxMeyWoBGPA3vBQTitykhY5ngKEHd8/Mg7Ujn1A45pmtFwl1kPFHZL8jba73oNx3erf5
wFJUXeou1BxVShNT9T+yc1rG3KazO30tfbnNCuiCx7KXsrI1vNKo2F4FOa13EYnrtDOx9453kPHV
Ga0So5tIgIbz+0ah3s9Nb2Yr6SOr9T0YVVWqQOXqVgI+DoEmcrG0Oi+EUb9qni0X4r7am3GI3yxQ
JZImWvJ6Q8nuDpXOLB9vM2gIe6BL6qS0+boSQ7BqZUxLYLFffTpcAIri3iEnHvsM6rLLF+BvnX+K
ATWahOZvdF3+InDSxso7NtYuzqS3kQbcPh2VRWa+X1FHoUAys/+pSDybtTrCA+P149ymKXipvpSu
VqxaoXOoXu1FN1d8cGLx6MfvwPhs+iUwChNK+3bkT/bPvK2NWvfxgwHTAH33RahooQUDDcaJy1k8
pt8zJ4iaeY3r3PeEPjqCQpfnLH8AsQH/m3vPaCWOG+IxnC1T1InBh6o+pfB9KCr9PZXSW17ngl6t
7R5LZRsleB1ZqvYkwmflkka2haEhz+ky1b3GqjM54zONgRl0x484aYEGCF6rb1O2Mcwnwjvcb0ex
bbpqCr0fPaXVFYtNoyHYLns6ccJLYzQPp2nbT6dU7/YrTzrKaBdaebm9vPMi0GAslcJROW34JSGy
j5agja1tnHt66zxbShn1rlPvA80PY8DU42tmzQF29i07ncowVRt0oPf/vG+eac270HS8iTU96CdI
uxcpg7TnRyTH7L7Wkxr00Zl6zxP9b4UslFMvGbLwWcmFXQr954kES/FGeTJJTb+eoiRukmwLTUB+
ZY4YnA5MUwSOaGi/GfkoSKiaDRccQSsQG/P8WP01BqTaiU0l/N/u3gStNi+vNbbfKSOhiF4EGCJc
ED7NTaEMx2GtBmk2PrMdbJBhUC36axPn2h6Yqal/G8s4QYn73996cPxukMS4KMiMg76tqmotkwyn
naK7wkkoQpaZTiauPA3x4wFwFvg6Er6A4nYuXoaZo+PQCOrOyk8ybeXkev7j094L1jK73cvYOnOp
mDyhJ4UsZ8fYH/ix6KB8ZIxy8aU1LclSUxwyiHzKd7/s8tG7E3Uteps2AT+G9bDvAS26YMSCPxlE
Obk+MY99bI3HAgEkEs/F1KAJsxKAiRZ+bCMXRnEIwLwM58EMyZD0u0qox23HItQA5MTB3KP1TjR0
EqOGhG7rkHHCa0cg6PLS0N0peiwYwIO2DFwGZST75OkbPDfFFFrCcfS+cuUjIHQCSuHMZO31Esi2
KspBQ9UbpNNB4ERzoD18pjSbFeG3QHYFQdz8G1v26JcakbKQW0160GWF1+/ROjTw3uQ+LUo5AbGa
bM5xe5Z6K+oEW1dr5xrzNXYB1SYA1UM5qUUU0ZCBbgDqUCQa8RjwPVAeXiGxEtGwMPLjKb9eiW5L
/1PFjrQrc7Xs1ldrX2H9+IdzWUokCw6roxSFsNmdw3BB7DcPJmDHU7VFFo7oKNMVLF0r+E3/EuSC
ldnXT+LAW8oo7hpTvtBNI6mQRxzGpvIz2UJyy2DIIhkxKWv9G7ZKCP+sSPtzYUUx3rJnknvrBs/K
ebnBfqPbnw8eJlSN375MAVpzsooAxwzjmf+aBdf3xtXdlDN4UROkt8ueKPVh4nmKEE8oxl0kmafs
8hLSx56K+8EMwEJk6CrTKOE4Yy4QObUOqyh5FoJ0UA0SXQKUlyPfafJixyJZ5WFjCHaeAUYrnsAe
Ay5scE2zQJ2KTD/Br+7VTsfVeFBxj1x3UvD7e3jcdBxRfcWVvGqbuUNVr80sSeBPg+TgsTqUbU4b
IiZ9Us540wjTZEwWTfEl/nuiFyDRs3QVSpprJ8g0jWjXgHuhWvXnKf+XtUOEyZA3oCmvuE+5xulk
WaudW9PawDVBzLY6HayQlTDABS7DKcq+BaLCNnilddmID16Z4T0wmkKYQuN41ej0KS1e/WkNxt5w
qHW4EDOsw96ZMDSKaBYcRLjsZaG9TNyL4uBdicm5NTkehcZG1QGrYTsN3CFAQUvIIe/Y9RwhbMGt
Y7ho7oE2ZgImmvmP04sOl8sCKKXKMdIT/EMzRpssNOtAKWpPCDTJ047LcUKh8SF+KNfZk/7O9Aq4
QphIHl82T3/vmrKlCUIS8uWiBFoRpZpuYtMVNvhntV+fnJggzX6vBuDHj24STpFzDaCibOViPPyY
Lb0YKCscCH4cXVpJpuzm9cW0S8uhg1eQdr0Q5717aSpqSRRCAQlQCxWpFl9FTg4YpmpRwHLgR2ps
1IjSHXQs/zCchRpfeXTFRBhn3m/BKD6QVlzefoMx3ClM2tTfwUyJhiIBTyw6cV3RSLAYOcPssTcd
aO/3NGv9vwK6ffec/TaX63UBTxxhlNmuFJ6xIZ5P8PuHzh7tDCm+LH2BSauRYcIG++Ut7HeT7mih
2p+B+2GoIwtjdW1DxJ6qI8XA8aS9b1OcQ85iCG0KvdFwpo85VrwdVsYQwZsZdnLmhWvv4svR3k+d
Pk7wenlSckJEUl6EjdHSwCkL9UKPykfylBkK2XNXuEfAX0F0glXmDHS2sIICQMKMgUQ86gno6gKH
bZmndCjswmetjmCW0AFfnXUplyThn3txoXaE9JijEPPregUJIEK2aQ804BYmmBGGcNaJ658+RzgU
Neq6pwNIHIfP09dwnzAjLRHeXcZszh34QBW3aPQCoJpKDYv6YSmZRZ9kFyLHXhiHjVmJTVZgY5tT
AbRQiS1K5fA6O5qd5tWnkgXA9pQldnRy39Wj05b3FQjOn3JLj8GV24NbX/yBGyBAMMkFnFAXA2XO
R2OJM1GzGE5D4YrPaYRmz1+v4oJryA8ARuFmb3D/HVcnpaY1Yuv7d/qSU9YudL2A2S2xWT6k4DPg
owTL1BJ6XK1XpzTcRb8zy8iX4gM8QRgWqeqIBIcClTYRqrACJrjNUSmkYMg3oCKYCE3qVEd7nD4k
hg9QFWZBNZqAkCRqYwl9OJsg9ryVSuVrvxKJRqoraLcw0MecMukhDikkaFDUiCwXByhtEJLDwjIN
GzrZqWK6ghWmd5q8hO0jB/Wn3L78qt2wIJvZeiTYgAqSR9C630bkdGMoNhI6ghSlTEDumRwrXvq1
llJtRueaeXYpFWaEwDSI6uRcF+4cUakDCNolrmRTzQN42KzRvtM+01w6DzwNfaqxU2SSsuOI5KY7
ze9WkQSYlSViYkuhhuS/xxA8NZZaG63E816StQWnImCqyzJnx0g2a2Ju5oJDd0mJ/DHSB4dlkeRa
cF6qFdcMM1qUKMBJAw9WAJxpC3erOimV06A/RG8/yf20nidaac5cUKnjYZt8gFjXX0AR9f9L/ISh
XRjkl5ekH9h2RsqkfegHpKorLQQJatldQq6QDpOvU3ATdSXDHGkEnVh8oE9F5V42lJxNZfo37Trh
1IxIiaCzI0ITVvDAB/uH5M4+Vu1GEasWENpQTLO7dXmzpQLDHY1LZvfDxOCOfRGxwuUikssaXaEn
8uyw32EBvOE51YEKnfElDl/ba4FE0xZqLFesB3+mJtfeC00kh1pccL65+CNeSae513Wf1qDDZe+i
YHdPOXxzII9bHXi+F/HQPnaa+8dBxcRi1iY9PzfR/Dsu2AnZfxUHFPTbprcENXjUcPRrgFF+Cdwj
IZCv61w929K/YCdzwpv8qTCHbCqjJr+xPQmWQ6Nyw6lRQDv8LQbYrFJkCIZ6BHDF5scjjl+wKmdM
YTZ6ZbPoZRKNNq3m2cRFQpkARJf43J+RgCotZU9GcAtowRlW+BpRpkon9pilj7OAWTiUb7iJ3Ky3
rac6g8lWHPqTZFO2plIdOmp6nF2Ums7EnjdK0MnWWlEzaRgxX1/niD/uM3ZHpaqBKql5ZbVoIA0Y
Oo5T4Bw9WO6aLEHEJShzItdp0FcJDcPCV8HRJuI5Flnludkw8+fJ+UcyXs5VU6eeK8CgfBPqB+vS
Uj+Fw9C40uQ5kaBSJSlpdQjFHqIDjTHqS8JQUnQdxzB2FmEulsrBwjiujwtaV16ZbiLGZ37pSN5Y
YHC9f30988P0MoxyS93FUJv6HeiASjfVZSNmQXMo+idUfQcYlYiSdOSLQCoZIMfm76EAUDx1FW9H
/Vi+dbDsSWWa1LF2GRYfl4uue4veZfKC83r8j8TEXXGrdHO7KzlrwcOZwSX0MKSXql5dA4KXv9d6
eFzl3bYmh+hEXhFYrFl76RXVBXWnI0wm+ScR9DvWb7/XKMuMDEEU1d3dC1LmxJaYz4qzqTgpZr47
aqpT3IpYq3KNPaDqD3XLDQZSfTKp97jVh+zOMh7lXcqxdtOxeA2bRKuXLxIC81V2nzIm2F25qbTN
G/fGWyGVx4LVBMXpS6/c4mi4eNBDsDDOOrC1VIixl864YlomVsObG6Ingr25NSzA/LP2GqaCfL/V
TXkGdyCzjgzFURXtcOy2p4kOYsqq0DTdJcOCDYej493YgwitfZKh4dQonOoYPJ/4dZLs9KD6euKm
KDYAYuB41Bpzpg9hW11gJJyekjfkGzoH8ihr1nY9aNTPpcoIXdfqQq8tJ1KMzMWsqpRQ0EEYYXHX
bdFPu1EW88T+aDQWpH99XOXQBrKz720hqh0+Ws1fatBymaLvg2zz0CsVsKZgTakNCdH+Pc5Q/or/
icjZCKCpxNRTBKT2DuMiwkEq42SRgMUMcyYOw1mxLBW7iDpkT4TgpsQc8rLuKeM6OonxJ8QvVirf
qncq9C8cvggM3c8LhEhhXvZGzNNcnNJtpuWhhd+u6kkbfFhyrouvqv+Qt1K8B+ha7hPKxaW79x4M
m9oJMH+m0xrdZMhGdh1LYFHxC0MPRTGD6rEJ/0PBm6DSIk7y16sftB3zdXS4L0g3gOrpTdDdtm83
M5KS+RplLafZRSBpgQfHfNwd2+iHH2fLnltcTOxRrWcJoa+8NG++8q+dddXe+MYzvTfOrv9jRmbv
KEDTUpfmmHqxDfL0olVTuWacydk+910Rn2DPYhtFSBBvOYkvwHdWSgQ1Kwn1x3IW5FxNYPlhVGa/
8OhT8NwewiOAwXZYhl3/t7rzo4lRiy9GLwzIROl09bGHWqVt9o1S34kP6C8ntNtoVhgOoODZxPDA
Lzx38Q2+lC6zWZSvJHBAGr+a0fT1Rvv6iLqXOyGZSPxVvtvXGpZIX8MGFOFzN2+yuA8SfPvq8BDD
hMIZ1Z2St4vZ4zXBApBVGjyY0x3yCiEYLIU/laFi3X4dhLzmcOhtovH6RjdoQr2h6CFrrcbZ6Egv
2HkuPf0Kj7U3eHnb+nKOz4E/teOLWSRdAGv69t3862rvyuAoFvJVdeD0SZI1CapUVa8CK2MkmLrG
S2Ep9eTjWL0G1Dj/vS6K6BGeX68dm8e0yPHVOh/pmstnzzFpwO/T/5AyNPlyCZOyHPvovsRR5m63
0uZqpjx2h7Ptbp6ukQrKbddJtdILZRTFUAJIafnO+R5vPy6HuxOeBe/bcia3SgL/OesntD3OQ1cy
Dz0kYb5700w0skPAfuGr92EbbRoRlxC9Vr9mJg6RcA/dtxToXL6XFQbO/0eF8qopb78SsZxjpaqx
mmsz3C6ol77perT8W8KJtf2owD7VvVQkEo4j7VB2flBDQQ/YpHIM4lx5NT2HQmVj4ElT4/QAmFcQ
OUFYPEmpwCdPZNClRExgWHBz1o5QAunD5qh6CH67+ueQGIUh0tq4RY6a4BVaFF0t10dJF3S9aJ9L
DKPmGOQyItPkI5PPb7xhknis8cBHaA1qTkIodDwKlIGt3g1vhal3cVV6EwSZuiBs+Pw8rBRcByhM
g7KwVkmw6sNtElxbVzcwTOS8ifhM0l4R60SZrLMkDJjLb3P1UmBY7jKTXHntkzSGyaQD0Fm404Lc
hniA4TorlCPd/GYf02YdS/lI06FXZ5M0BOZxS2LU9TfOcvIx/OSqRuKw3KUYMEP9haMEyi4oajRa
DSngWR8/eTT8S21oF9HOwniyPfbWw9zj8q6q/N6Usz/F9KINkN1KZ1H3+dAhlP1zEQjkWvg9ohCS
ay3dSWEzgr/gJMnCEBMYdAkbeuxu26Txqwr+eXlpaYwi0VcbgnO/WOAEazEwdhrsgeVy1N6SINlZ
fw+WwqB78AEWloQtFAfIOcAnOxSzoOsEo80yEd9S7Q1t/y6it2N7E6qrMo3S1KTIJDYckAC8Gebv
Jo9QxGcYFrJsBfWDqQruR87FdIOLURAughGRjVYn6e9hKNDvABO/lfP0BeimZNn0zNBtTfweWsrq
chNI0atP0yvZ96gy1De2wOK6/UiUaIudDv03VHxEIekUrp9v/887Cwzsd9Gxhn7FcDothrNcDbXX
d7VgoKgNfBNgy0RE17PSWFzvFZq/+nkgDypXTQqHbqUEZrkOV0ex6vyW8GMz3CMLIrQPfjWB5QlD
K0RBdEGdUpsmvF7cDzhfX5qc09jD0nGUIrqPFUul3RBdw3EdCdJmjYzWEOKXDOr8lNNIsA+wP+ZE
CO31Hj36LSBlDdxLmAh3Tc9tYExprtFuph6TJ0o1LcSWB+yyRSYEgNB0N9ueN21z1Sw/zanE2YdX
1J8St4xMzKldAzuYYauMSYJ53u/3dfpLLgzJ4fC2tyyS383U1a2HHRa3KS4ZGhBKs6KiKG+eaOGu
Vc5bYHp+ze+imVEB5IFRSNwRnmKksOkBTA2auwMGsL7dbOn2/FpMYVTgMTK5T5hFSWpLu3M3TwDh
vJUyRaRMmiZROSxehfkpeVC5xXKN9DqkgH4nxY2Hu4DeNtu6VWif7shru01GGw1TX0x51ajhUKLa
tTR3veVaceM6o6wUcaxX8brgLOVvQHSJm/yBoBFlSTz/CsWFV1L9FWpDC9DuxMV6FjT/ab8ErmgG
gQJ4uw05lW+JvJHQWm2p2FXESf20wkXdMAMoRAHc3mdFPrlQ+INNeZni6P+uh5Xe1xGiXGFdh4Nc
+R/VdnQHS5DmDouHs5qUIuRc3Nfcmfrh81oAk8m71e1jeLJYnNJSO7b+mycOS9LO4L7+gzOC93ju
ZK/xmQEMXsDdeEP82AFeGFV6LupDIypdBhBxTVhX/zjhpLOWLLu/LP/WDVN06X0jNQFYsW2rhbkU
WPovfcvSMcB3Qj8tOXBDDQcLwkLU2rZQdKSPoTdSwJiuUfdEAOq1amRUNQa1Wb8cNYxe75IuN/Xc
ZTkqOa9cYwRSzYzAa3foqwc72OfeTOrnyPGa8Cw/7XYri1kZh3CnQG7mIxQZCXg98nMz7tef6fx3
1xp79ngyirSPHpQFseBre9UMZQ8JjAysC6qYIMHz3mdesZSeCcIn2CMrceTOtyATbMPteVihNUdZ
o2p+M7xsq71t8b8Q2iiPFYb8Ja/zkT9Kl+cjdS5Nz7s0oyvjqed4JBFvpLcJZjhNzoruJ3V2MISq
l/HHExt0DgtWkFpzKjzAhmMMScu0mAxeQ6UjT1F5FY6scgzBdFtnjgCjo8oPE2rIOdeQEmh71Znp
KjWUVLv8nN5peOI7uiXMXZFLyod5wBkHtn9RaXJIDtxxb4HqTryf1O+Leadt5oEUV9+VOIGQmd7M
x69iavS5eUIC69ZelDdu7CZE4UlbhZrAoZgYSYwr0/e/lC+l0kfJiGBAJCJSpyGO3OH6HY/E6slv
3oKsswKiaTgKmvbb798dh1UVN9YuRz3iqocE96itBJ8pK8jr3QQ/d5baahcVOQOOKQTDDI1xwjlO
YA9iVQ25S9b4JUkV82f7sTc7IXzKztMmAFz759BBaNlbqSuMuVZNkoLfjfKdOvFtNtNcdbezOdzH
sL2zY4Db1+4u/GZWxJUG1DomWsJUPzkAaa1383qv4DM2PQLbM7UGLMgcDz64GcIa3egrgGSFT7Vr
e+tIXrja/+MZlY56RnI2KQmIWdL68AlCSLbHXJprU6/GqbajRxIKo9ygSfckuZLOJgVfx4CQUMRw
+IGQXLM2/maGVtmKltAj8Tbh+VqWTQDJDiNP/ZKzMyFVJWg/nGTrMlWtuvfHON1pHREopQfYKgr1
11Da/K3s0jDF49gxSYVmHl1sys1otCSEovD8eLETFoJ9mOC86uRB4v5fo0y6RQWMuKS8blZd94QS
A8eUY9qjuOq7kIVELB/3LcjkmEc5VIP8Ty9VA0XSZmzucXGVYVj0d0xp30V58nEbNJDMG/FeZq6r
GPH52BYgiXQi4K8I20n2XDpP48W0J1gxoGg6kl6FqgnWKdwjeQ9o7fkaD5QVnsNr9GxWTXJpexkw
dZOqAOvyjABfNrW6UOoLq5M7ftRbLqyhWQssVUxplQ4Bs9Y4jPc9Q4edlVIrq07VdnjaBF99qLqv
oN9qzZd1WVguMLlyAmazEdmEhn/z7SsbE8igtvFjgOAYabvxSzrSKMvYNXndyTLRIusCTrYeh/+5
CmUzIr+Of1URIddUeModgc9CjKDmiDfpkZIQL3jiUEGELyoNUiq33OXCM7Kj2+R3ApcFM0qHzxro
jqg7G8TNVUxRtJGIscpbbLl9XMkPJPgWCpjgOyIsx2JmFI4nJstkHdGfw6xdGnhtOEBDVpuNrkke
oNPF4CnB2x6y856/E6fosCCW3Z+zs1t15U42GhQ6/2PHYXoIx5G4CqW+HSL/AL9SwvlRwv5xQYTQ
2jC103PpnR3Uj9wtrnb472kqeL05SEwo4vpYWtG4Qz5rMi71ElzJdP0eEAQKvUTjzOWu9OqBq85h
a79wHf4Qvm3Kwmw4OfrOSQFJ8nVAfiaFkA4W6hfGVXDgWSsqYM83Khatsp5og3GKDcp1J/rPxYXb
Ecd+IZzr/Nj3kg2Axu7mLlRzK7/MGo4JJKAl9NabXbY5KtsnyrtdDK+QtjSVwIp6bZLGepJ6wm9l
pl+BMxs68JspF4zgBAJDYuBLaLlcquC0nCROcr1AeuvLLdH42RkXUXfqMt/nzpJdi3QgxVQDrod0
zKR19he5kN9mQ0QdNQfgn8dmz+pfJfwtHv1U0++aDi4YHrunKOi94W0aPpJQuQweIH80izRkdzQx
eF+oZrCM1XRS3Ts32LpfaANSgXmx0ipy0vldCwTaJ9NAgqW2963Ba/33Fjh20vtJDHb9Yk/ZsHMb
CUFpOfy50OXR+5VO9fYLvYE9/wySzYwzvIQhdpkBJW+aYzsqjGfEIaJWAO6XeKt3DH7Vez9XW/N4
YdYiQaYhRF78uft04oG/Rnx1qfGoRf3u1jaWTZLUrNpBrA9zjOgorqPOscloKI59s1OYgdpmhKb4
czfpGksht+YOjNkwhGnrTscPCs3WfZ6fXldS3ujSIOarLly/zk4cYY2ctXQrBhOpOHjtab2D38Gv
k9aKOSkcXENGe6yyWsLDi9dAgZqInt8VuBe3R1yVi3KL/+tP09gLkZWOVYcmrpE0tKsMMXgp/UNK
k8RTWMqia9aLMrFGfwSiLRQTixi5J83BDWrksIsfWuMGMdr9lXGWVT013W2T+CVTPLJxSi3iTpPw
TQb9IV6WIF1fCN1n5awuwJPXTs3ZYQ7IRUYbZ8U8B/lXwlEhR00k+YoNqYvWM/5BZGzueufSxJ/G
H5ulrYewgJ8a6CQtVzuAxMNIcs2/9Y3LAQ8gekr4aQ6aJWADS0g02R74eU8gaGlY/7LAfqJfA96r
TEM6G5bq9eafBUGnmGAc/1omwvakspwNiZYZEgs7xkUcEy/XoXnGcXLNIdvv3ur6Xak3awe/MX/Z
rU05CttbM36OQ/LJkBIoqOIYSNPHBmAnNgoOn43Tj4LVyHQVuNwvFDMvnN9orX9uHnulxLqWM2tu
66yzVT6gNFD+tJysA9wGak6E6GJXsq17FiGB9pFh8y+OaEaxe47H7ZH/DsrhnFFoXmARdFdcJyoO
wRVXJ/obUM3zYQzRn6exnowv3em0WBoFauVhFWw7VgNdvNw7s9iB1sQ4uPaBE1eZbgHe/oA1Ga8g
tGNQleeyWs9zrTjXw7zFgy5wdkLlIxiDnib7IWMDj2oHNnSZ4rp1wJCKQNhaniUp3sSmHufXyOK1
G8lLLxhvspU5b1UfBID0AftnrzByBrJ13BfnYIJTtClUp8+n78yNQb+FVFdHalo37BAP04IqZFpW
0JafvcnSyPCHyQNRqANcQ+hyFQgxXg/glfWoXGMIQBmbXi5T+Z9WgCtW2zcsRWyZeUSOkBYDSH2K
TJJ/cUCQc2QwWHB8G3kMU9rWTXNkv+y7ew0QFB8E5y1HivhsBsQXdECBM31vYoni3NMB3mR2SAeU
yN1lX6rI72P6Xho36vQmPBYo+0SRfbQkRgJm/ALEPrt/RRqRPthrQBAGHF8HExH7DxzqPyoKf1Qs
u/yTqqV2sMA5IO1SaRwBUByXTQEf7Imc4x/JO5DHsE7Pp8vd8twT8bCObB2as1oCithRcTT1UhhU
sTPEBI1JWD5v7Y7NZtOKQXdx0V8m+JjLq41ItLv9gG04JJtKrfVMuwH6rSq7vSUgudYQbX3etq5Z
cnSt/+PD38nTSdd34pw+loamz6vTZ6hV3UOqYY8T7vzVMkFty6X0Iz+UtK4NEr/ADjNZXxMPkj1C
MwxKgUL9gJncbgvXkU8Ygy8yN76xSY+CKx/QDF6tr1zBpegVe3YPYa7R1IEyfR4SgWNtwLZgbHMU
nCiZIeVmmAGydvfqeeXwGwKMHyaK9NJaWc8S3weLITzvLmVPyLBMwQd3aRdsrt29nv1Edy9Ekj7l
cv9mxiaCft2I9tKGt9bpazQa69CTakvFfHFPyjoYRyYWeh8EQteUMkXu/KIeTM2rn38dwXXBwUjm
v6oLcEVJOJEp7CSwG4dVsVvhPqTrJPQQiWy1boCHjzxZadH9pXu0QV6fVXi0lh0WbhFWcjuLyBH4
hh9bTX0U1Cqr/8uea3rALTZuFOQrPwAMiGHPJz4oxGERshcRQW3pMwhiIFoKYVRsyz91CqHO3F54
MdWCsec1OD1TfqUZDzIjN69wmikunjXgtYJMNVI2W2nV1/ty6YUtfdrgwxz4WB2axtUHlPdFlrLJ
HjV9SYFwYBa3baMEtiHBrKGt1O4x7zJkyeX1TfO0b7EvJOdc5Awqp/lbk63xmB+gwcTajPHxdDBA
kWuuU79g7dC1vjbMrAFY9GrvPZ/5Z9Yw9IowbS+PUAW6n98/19Twvc8nI/lTJAf0MCRpWVHtgAtW
daUYeWScjwD2bMxA9dyB5PAsRQRY14pJ9HpRfXzmgZpsn1/f90xrui+s7JbcEq3PIE8TP3Z3CTqN
0phnMupVIGb1TMSij3sRGWbt9Um6qv9XLIA9GuMCC93Cl+V9GlALL9P2MFytK+MfvCxgqDTP/8L3
ZNDdS2/xf7nFlhlPSPOEU/MvKLvAwg0wfC13rGr1/pZM28pk1KfON2LiqeCeHOSydqkFWlKy5KBu
faBJWNDxgUlBYmKaVlqKXct+cS+Yc3XGDom61SeklssN5Dh6sgQOkphCWSh1TdC16r8LomqbkmuR
3d/kXYhbAWLzmemsmRule7CqCFo/NCjRiWfZ0RLQUjNblk3SvRxB/LbnVm26thRLJQ8m0OZMssHa
W9y5vGMlHA7Xat8D470kSnhGXTcsQojAyCzWPindvFxpGqnZxZhp1NgAQLMk0abue0aSCtfGrVGm
MCq/nLeVVZvNiFfEwVBtxcWITrGidU9MCWWMVqu6ru7k4oDqYZlXwW8AR3AQlPBD7dESI3ZfABCK
hWUb0qaVcGg/54X2POKXMiIQMHHx/guRGa5P6w0KWkWNmwmFudf4ufUY1SF0DkZ2+tfGDYWspThY
6wVNy6kbtFm1rbGTyrqdrmGQa1qgoj6RCqIo4Uon283Ko+Y5u0YFZKrwuo98WdqNSY+PIqaw4yEG
nQyi9XLAlH36O4nlOEsBzodQwd7W34T/n4QNLQDVKyolMwOgDHe+B+3D8TFKk1U4a3QcTr30rg4X
iVKrtj7Ar546rcoE3NveEzRQLVln9+bGp1GbnHoW08QJJ+nYRqxFHLeLN/xiqTVzKoyX5g4P1g8B
HFm/I/aJZP85Oi8TPTqmV3iKW8FtAU9NfhtLk6kN/ohPJcjUeGfMOPT3Wqtrpy7HwfCcreypT8I1
mXKaaNmpulvEtQGCAPMqGxmZTfoZgTXgvPy8FicKpUwnmHn4Uq1hKIzNVn0EvLej6Y558SGRM2HR
W0ceOZHM+Tbu/Krvzew+FrKdMaw8cKnwyEKUDs/88FLGuJTEZPYqxVz028Gtq77Q0uxBq+ZzeXWm
CNT00E5GaO5fM3C8kHtP9WvGh+Z3gFwHi+8TVkZZmlKi8MPzv2HFeYUjVYENlpvifsc0cqroca4v
xmhPI2NOKcSxhraBYrpA2AHj4pXc3un1/zl9kEqIBN0qmJ7gLpJ5eQuoEz8G+/K6sGOHrW4/OnV/
ZOT1wfyORv3ONYn58dS4IiyHSMkR+oXyGvUbi+0SdsRnTipBt8XYdkLnWlVFi81bhjf0NOKb2TCq
a9KXcB779BHm31A+Dn9AwGc4XrWon2cgfqMhUQsW0/3xCT6m54YiLH2fu/Ns/lGHXi8U2ygFWifB
UGkhVCFCxNgB42yH5eSZFsyLN96MvIR8i2bw80czDyVxvfSWmU2ALzoa5Y+fOaqdpNUgkiRQvoJc
CkncfW2Bp5O3VuJr5/jBDBg/piz8bX7NEZ2RJp8cagVbVATA/iC8M3nLeaRaQfZXna7XPorlUyho
wJ3dhFjmF2C4h+rmIpMeHvB7QXJO46JUBpBFKvYzx693B/yskrj2Bab136Zd02ZNxD7j6J4S9B3P
u72t3W37cMQRDHf2fJOBg+Bk/0TZ7B6yfUn/HReUUGmcbbdtyhIOQoT8vS1cU8Di2FgAqUEVQIzK
C+a9HOaeGIeW86o99NTaPWA2jw8mRKxYoq5zuuYOuMPvi3HxjQzuWoQ/4rhVMZQTsH1jjFDnRFiV
3P3kBoedsWxTNTxInzQLvvLbg49bP9qHRz7pKJqy3hDSfToN6/x0/XFlJavzbSTqFfaiufx9rv2U
lrgiOgt3BimF3p3e/LoK0ACaiiDs9SB6gyNhBfF+hrFo576YFStORMqaVIC34s+4aAjxYcaaU6BD
bNpPb/qsttm46pZ6GoEQFUkOn9b2cunDNOvCDVJ6y25p8bq1lT2l/0zfXlbPe2gpCJZ5wn3WcexD
lzxJWla3VCBJRn6KHxttWCHIOygLg2Eb//g2ZrmBqA7wHNFRL/T5Y6Z1U+2S9BD3IKroX/RPV63e
QDPvY9OIeME3lTcqPRVaxKkUjWYpBd6lpqYziZCY9hu2E5pxEGx4G1LsJRyhY1bE/mwHNgs5+Jwc
erNbqf4peqM2Mc5ewUvsgOnyX/J4RIpZM/faJwWpGguNlJL/4jHtFDuSdt2l3RpUYSy2OQPZLlMc
4srPZYLjpsw8L+YH0o1SCySOszMU2iDDU06xNKO08q+lZz26CMsrmQuxLN4WXufMSFfKQXBnXyDn
Nkij50ZKdJG1xZZtpFOf4WdCLeNjBdNpVGlgMGwcPMKLv7vIwnsUy5EzWhyrBIVU0jIJsE/BpwWH
/zwe3RyHLGmReF7nTrl9QDmxXeF6uiFIaYnt4oasqZmmd2IXgy3k06grHXtYuM0ZzNr69UQwOjRW
KdHwgpgzASeECrU4so4/kyT8+O7pv8uoWI+PrPX3t7JudllQNPwGxGw58t8L+1TeSq/EoTLKUWBG
8LCikPoe23URxUcbi5fz31VpwdHb8xgAOlJn/Bz6bt8dAoGaeJZC3mxaXdaqwYPGzILlGowTK0zE
HLXCdqdnvMEZiLxQfA186tP05tutNPXGS3RTK/r+Y48WKSQ5WNgqmTnw9/bF8xxBBl3P6Ldi0l8P
eO8oShJqz+jXgmB5SIkQSJgYsfIY0CnWQA9+CAKVpG6AC1qtSuT1PUx8CqEThw5tuc/QgVzfYXMB
aK2/zOmnIXtVllw0p10O2J+VlrBFTdOCZokASDN3/SrJV/tzHXzpRDBQuq/XIy+cOwp6rh2X+pGJ
K6QkopheS37/lrdc9tMxeFFgUjOdd0AmuuqSRfHug/G1ERhGtQ6Km13Z+M5RG6VJnlGgaJI9uU5E
Ae1BSs6jpm80lNZLuLSVoY6XKciPHEJYNlrTg8Lyd4ONFlOcRUQ68b0zXnHnDymQKKgDyxeISjBI
ORQhQfO5rS3dakAz4XS2cfGT8dKEIGIFyyj7bHVv5WtnKQGuG6fkeotmQrWdeGf2zVjGBBL14J6w
ZHue5jBUsm5U9ZepPRA4h3VwZVzCgUYl1+P09zmlit93ItQkJin+pv0cgWlHyNPqP3xtya2MjT2Z
uijX5kAf7fpSBxtzrtVsObJIWPUcHCs1ccVJjpX1yoy4k5uu6MNCa7t2bk74z94tWbzQEwGONSBk
3Os/arN5nz/4zCdNqcXDzjOkl8dPkN49IonX3fWVIJMbvGEmQL3cmMmo2rvM/lerQBfNKwkKSNFO
18Q0Q/+xusBg/le2hPhEFp9W5yTxnE+I7FJHU5iJOBOFr2bGTkbRBt3xq2oD7t+dHMu9iHuRqXFO
BqS1np01oNtz3J6JlZOERkeCH6u9BPxKlnXBv/EoIthjlOkxwjiegXSQ2Qmx/+MclBqq5nNv5LDL
szJNrwK+I7eMAUiw11jnXQ3DE60VLhx1VCyGItvTD1z+6ZKRlXqkNlPuFAozItlJwDz97QshsQCY
+Jbbc06pi6fg5Heqa+25H+d2FKEqE3kouU8EmK+8DzHgsLhXJ88gQI+qLpOLeeftvkWMomIhQdF8
uXrvnw6uSEet5ftgLQnYNbABKEBJI78JlwqYycEbskLCnaFXe5hXhy1lE1fk/5YLVQs6QC3l+mw+
QSDG51SGb8zQjDds2PLirUQ40giyE7SRdv8XW9kgkppsRjRdvTMXuvYVh1LWOYQOT74jCGdtDWN9
KmOwSEfyhWTt/gZeaSD0OeVkLr3TLuNy+mlZoxQbBOyD+GuZi3b7felYThBn1g7z8fDD23BgwdBA
U3rjmPKBoNivNtWA7hWhhBqXkTpUOXWHERpEScrok9ndCSdkQMRlClektX/WzmHG53Degd/cWHfw
scI1qi3BAvAMWvSYaMRWOdS4yKirFXE/5Z0FkRUn260g/Df1fZfJ/EhyqdG6VEcG32I3ORTCGERZ
YhHdatBCBBjA0KlI8ZnFI8dvvUzT+tXGktDSXghap0RH+ZhW1tbZAsLfXiw/A0FddVA+NjG631fP
ECTQpfh2QdFSVvuPQwYzEjIAo7+QMxUxx9ICsx9nNLOBvAjeII0ZfQlO8jvELteRjzjKurnzqzKJ
+RpL5XarDTV0qd6+qTjw9utw/3RB29r4iA5aeHTFPwPrQTQz8Ou3MZ49EqA1rrYZoP7fT5JZGuCE
x8rh+K79kbywHTvtMXgwMsnx5lCKleKTzl/+zJRPD9sNUCrcH9kkCtwc0yuAAbt/kip7zlaTlAW4
Nxdk/jLA25v4A3gWU8dld/WmSKcthGHk51osor/Yp3z5Lp6nM6OPOZe/vU5qi6/eFV8ful9GWzJu
MDX9J3rU1+pFD4w2dB+I1SVtV2uq3k9rgYjbLFe8chiOHdIn8xcqpbqRoqQo0rq+8z5IKZbsh2zE
Bqd03toh60EVDtYCOvbuYCZyIptbiGUUDb9q5o11l1FSz5VlphO8EWN0BKDB9SFwKtWobxU+ucv6
KfOLv/tEnUeCCDLpnCLY8j6SmEwSW8Rd1CIuS7j8OVqy4V0pva8LnXRLY2nUA4jLh8OomyMZHJxB
cRT+hv3bifg/S1w6Q9qfb6Wyg8kUivyE+YMQpGIAH1kImb/1NXQ/XuFIe30unaGhokB95IOxzKZY
TNDPDzbh05yAocw7t9gfTQ/7gy488tIK7J8DWDw9NraHUdxtnR+SwaiGPUo6CgN4ycbOlyMW52Ce
GN7jtXvHfR65qU/nMYuHsuxWcJdVIGDjUsqx1Yu8pRdWIwk4lqyXKm61XvYzte90T+gWVckpXhx0
ZrbgujbxtnXvEtAJuWw2oPMtUp0G1HPw4l95l7CAElK6so9F2LxMfe+Ynkleas4KTJloy21z5/Tc
LsImlvVA0bbLdHiH1G4a9fTk2MsP1PIevWEwC2TzW+2q2UCnYW0qNBxUsbxmKj23m70aoVp1Sr1s
6UWoFmlyEodiZ8bjkCmfXvNmu/lbPgSm8VsAfkGNG404n18i4Z+1qim/fyU8YKqpyxDLsDNkZUID
iYQFhBZW5oVIlD88GqjWxVfOu5rGwRaulr9KXMsL6lQ9UWjB75a+g4nKO3dwslH/+gXp32QucSIm
TZ8uofQa5Pxvaw+HpofqXNQlAjFebosHBzXc2SJ51ry+Se4My6hvmTdcoxIPklqCj681uSA6g1/w
JVhGr+QfeHPY3EVABIo1QFQ8tp+RPyo0VX5n4wEbrdvUJpnW9mtbFX/oSlMsPkWIp/jDFK1VyJms
va7FdsvseVHThkS4d/R88yttMjn5pLDzY7gbRSyxH+tgwyqswkpCUfBWlhZD2rp4ikIa1tKFDyf+
rM/9WYDZ81tQ9Cc5vw9IGqsik1ilNONulkMPvNz9p7hVqrCGo/f+ClinLD2pnO3/bNVbxPeOat88
1Cocek5mtKZsaWj8SW9L6DcGp+Rq07vjqdvnRoKwRPMrm78cThqDF/daVc9EDkmpY4f6j/Rvsw4U
hwwQZnyooVnTS4QZxu8Yd7TFSNH1wwWiTW6puXm//dTQxVJIFl9CBf5up/tQjVlySzDUEJJcmrXA
LEyDx0+cpYGyE10ZKEaHRm2YCyq92CnqFLtHz7x5elEVJuO0Y0PNp2pRHeuOGhDRA81Q+EyKRHCc
OFNeiP6bvP0IKmY/syebBaQOFKJa5p4dM4jYiYAErvtsKO7GNK8Kvmhs7q3kTA2yWHD0dyCO8UU+
RaYXJiwcnHVoBhhbrKmXVs5uxovKT7zXxmB7O8g/Jlu9n11jbdwEd2odzpGn7XiA2+c9DSg/DKGN
eT91RnSdG+7lmlnK50oGIWhL/f2MdEOuHOzegSR6P4Dl+48LzUmf2zoGoGxU4CR/9AUW+/IksfBh
Zv2pJTG01MHNFFY9fWUfzeTuflj+ihSgWrgDFulvz/HObnWWkMHhZHS70z2wuplZSdlwwUrnX3Hi
xD9glT3/cOHdZtt5bwcVHpCoojSWdP0SSiTt+3Tx7o7+FlwrYX4wz3dcP/YikY9iOucK69RWMU7/
pxzjTeHaxEhMWtDTjVx5C28RxDUNFeTU0gy5wbW9X5CMWNRTWIKnavuMrKsqjwKO1knO2zoHQEV3
SqVQf0QDLoH1jITnocD60Q2lcZyHU7gI67EZyD5Fgh17xwhgnJb0Ocwut2jSuGtfgtxF/BFS6D/f
8xXKa8Gehy+ExBhts/Uh6smTBKCW1iKokOiIEyKFAI94Q7uPATvhi2Pb9GN6j0QtkhJQSoIc+fJ/
NpXb/OKsWUr395clLS3Scl83va3Jhhcf6KhImsBqXRnCUQV5GTwaGW/cMevLlcJqBnFz6nsJ97SF
TKieKFpJDglVb7sXOu489qyJf54nTye5Q7jVV62isNWeKea06M16jdwOqx+sRqF98pGV+az6fd+l
fH9tEg/CKkGAJTNhNjxnlA8lBfdk/QxO0FpDqOgg6zt40wq6OjtOAJ2Ceerufp+d6pEfJjaouVM/
+T4Cy7h+i69/gesX48C71yjfi/+ZZAdf2c1EovVDp4uD9yOwT83tKtbn9ZaSALjLzgUYY1e5KyCP
ohmAg4PKoljRHbG99vcrrqSHn4vPK+SZ1p0oyLeNyGNZr2qB/vZRs0AZGcW0tsD+faI0M8xNKhej
i/lBL9fRSYfhti25ASkz1wWGiKKRzt+fy/h5kxB6Qq0xEIvcrh9LZTBreYEWpHeG2zUPUW6QuSXU
D5vGXfnrYmmnk6nU/D2TMbi/qgImGgQagvjSilnXbGB9c9+ztRrRa81Dzunu6dT30LkbsGhhtT5A
38sV7kae66uXNvFFVO8XlppyzD2K3967MFjrhrwiy/d6YBHUBkokuhCaE6JNdmbvOXQt987bwGzG
pFKkZlorGEBY0bYo5u227S6Wl8dPKX5lq2grcoXfW81yu10rNxGuteM6aI0gYefbRK49tntus4Ra
gT8CXeRnEc1EJZpB9gW0WMSRv5Gd0mFMJY38UQScYewjV16/WRLINrH5JjLsTHXmo2NM9VVccSwn
gb6TP7WzOX383qJqm2Dkh5fjOUI+1tskOtQmdMKj0yHttHQbAjlXH3NbM6ww3IIBZBG1J32J2S1g
d0/LtyTebRD7FT44Mo5PpAf4e0VB6hWDAqnR0WsNphLKNrTSOwQeRiEGBInfNm5qcMIuJYtoPLbq
MKYmYyc2myu+d3o/gti9ZGP0c8mjCxMJwxGxDy0626BfE4pgZAJ4d1GNQGmm5yRmfYzoJDwngMGp
6JgZCVy0r03hW26zsJ7vOuGPczDAqJ8XCp3O2BLqHtJEs/t7F2r1s5IVRLvJwsdzMZqqoeQBj5tE
dG3nGca+Bgntzc5+5GEiEDLrCdINH6WQ+9S6YwGjfgROqwx/FJnJ00HSSu1IDdqM0WuGTz5tXgkS
BHrQEosYkjon7+c+r4tAxnlGWFbJa/Ikn3OqK5t/Z4h1/NKbUZBP2sd+o6cmXWA7Wn2EnTJCOyAt
saq8PyDBAwGXN0xDina9b+NtBQWNmYzkdJVxiNajVRIhfpGyiim56F6pwU0A4JEwNjSh4Zeq5lm1
sAGdZSGb8YQxPGak7IVGGU00i7u8Uf7WB54aBcgGezdcmDzsRBBlikc1NgWQto+ggbh6gXZEvZIR
dtGfAoS0y0Nzk+1MYL0Y1vQPsoSIO8wOIP3qC1oJ2zj1ra0gY7rfKQ5eR3+T3EPgxmWnsNA7RpWp
hrhdRE60unoaB8ASDbxO5CuMOSv/UVwo3pkOYSfkPqH5tHMLIHyhecVJ19663LwcKugolDdSR0zv
AkS0EnFwoOsnn7/Q2YHyC3xej0BOXwd7dmAIsFY3IxSFXylbV0Nv9lkVG/Jalym/MrPE5wQ5YKCi
OUBb4Gey9n1KxNmCFp1yKdcdwW99acKw2uC5Ia9BZDueAEulrGrXS1r2WWL4svFVLNymZkpIZNvv
XwnJuWcc8Dmp1WMIkr58Ak5tb2nF0m78mrwChN1wYvTD8Y2yBj5EMFmoicOMM2jfAeLEfUYfjxlH
OMTqrq+e2y2UT3SwEgoi9P/E5H1NcGOjthowQ+y84/fay8IZxjSXuRuNcsxelIGwoNrf/2M/T/PB
MSJqL2mVIPI6DpvYmjJ6FeNugZtcFk2kWhvNpUS6p3BBTXl8B5K1CUe/90Cj2jfU0AQRK+9hTqq5
siDhrNC+1GI6Vf/hlQ3e5OxQKi81MobFDDuKNB/EDGpUCQtloDTVZyyjjSJ7esWRLALbWa7M/KhJ
OPi6xtbpGJE+v2r051P2goAQYQ48Uo3jxCQrOkJ3qdseF791Bxk5448yWWzHHpcxszKerYrBEB6j
ZJF3kZEQiYIV4Ap0NAoWoEHa8tvb+09+5D8rM2nUj+KLavzbM9X9ojQ+5SpbtfTZSj1GR5tibmG1
IiMBlb53jBofOAxDifLa+HSI8vHodAVDYy5HUN/gYeo8isBoXTKR177XIzj/btqn3yP/XwFx7jlg
0EK68PWdp/UH2efdI24QOxICDdSwaFI32WXFdV+oHInTxRanLrlfpl8Bj+PCwjkwFN6gy6fwuKmY
HIrq9xhT43PRHEQ7rEjaiJQTpjpkxb25oH2RVRLASxj3ZLAMfNlO6iiKX7JwhItad6FBVhG3144t
HslhYg4ThYsX+J2C8IvrchQV8X9y/XBGkEVzrQS8J20Vm8msuiQajirzeK3f5Juo1WXQWrulZ9zV
Pcxw8ed6wl7tMJu9L5jyZROTDRXBPlahlfluwSNZ4fr3h2Xd7dYOplPmJcAN8ZH5hZdPiTMrxgXN
PLXhGsEJwHT0xYqo98aK3P7uEhv6YsGhPN4SEQc4Y0WZy+R0X0/6ia7MK4evFL3xJcaVuZaxmK1x
Lylkpa3NQmE1DgZPX403dh55/yBFjHhOzcLORRtRp8cjDu6QJs2v1qUzhW0Et8ByuO2WnLM/ccyB
1uyUVml3X/mHJm3iiwu3xGIdaHd5PJykomBZpHpCLQq+DERsg3WEsop1jOMgUiQst3tUxabyIVeH
G2I4xJkQXesK3Bb76Dj+t45V5Urk/Rj1U7XyVMFy8Cl5JfyuTb96Wxq1h3jI2xi0MrNM2m53TAz1
IhttNI32OzOvIsCjcEc8KrhDqqttfiGPyinOEdH2d6s4yujloArOpux+htMOTrPrh5A2KRvO6lM0
pG2avQZz0zIIjZOBgxcSaCE44D8/AIPiXq6CJlwSDfsnFWhwcRQs+3zLu1N6hoIDzXyl+Ma0zgA3
Um6u4J+EagUsfmzPY9WxbhNub6EntkgIxnUdoe5Fo56Qh3JnEdtXYEWQcEHcIsuN3XFPRACmQa6B
jytrq8RR0sY2MDGIiZHx24KY1GPEgZjxqUodG+ZccYE+rHEHleQSIAZkAm4lcFCBILbvxLfPjXcP
oeVj+z9rMAuYyybCmRVBYzagL05Hjk1urtHUdoMq3rm5JcEQa7tZ8RHD9SdSjmjTE9e5aZO2r4Pf
t/Zg2nBO2bXGKfSWHMs1RH09LODuIQQkaF1ojvTsVoqdSSEaOb435D8P13tmMxJk6q8KxbHylkei
X+naDFODs1B7Ez7WpFdOtqhasC4G4SHZ2dOaM2mbsOggBRMSsPHPuGiReZdtbdg9fv7aXe96oAYr
b52uG+hQay/3gVkr8iPViuH8Z+6I9YKGJWPN9f/25UhIP2IJW+PA+b+DvFqHge4rzsGdGzJ2ot9i
+Lx/OGYg8iIgPXpSZXoRY1BTwX4xuEhdbstLBi/kajcLdvlNwsFRTG2d/gkCnX7qp8kv9rIUGpw0
expNS7q3TkJzvR0MCIT/rZTVvLexzmx3P7JVKK5NaJKo+E+Ju6uUzBg4Zda11iLS/WPoIeV5zX/Z
nONni7GGp2ZIlfti3c0+cP1WOjEKpDUeGFRgZVPVij4tqBDYOYE543Frch1fZXX3jVHUFw/S6QYr
YUPQCbydsxmItnASbkeT4JoQ37w1Njw2c17OyOlMTUOEDsyWWoBLhvxKc6FR6F2Mse+9o4whGUpx
H9Xz0/Ficsyy01xuDlDi974R/vGGtRlyYwxHDj/qZde3oUMvix+2u+kdtTvINrunRqctF+5R+Vmy
wsdmFoa6G7Ky7ChchOfYCsqtgt9zhFQbbPmiNhnMjU3NQMcBIHOUjXqLANVjmGPAO94mMc4J0z6W
9rVU6LWnNCd/DpJeZ6v1i3TmkgPP5IwBPECZ1G9/3MgPlLaZfdrvXq2HhFZZzBE0AC6D1IGjDl5j
9WgxPTvGGTpXdC9Kj8IATz5Gau2UuaLAu69t2rS5+15IrIV5/6ziAXchoCdogVMZAeo3biDCS671
TnLf0YcRTGvzPyb0+2LkXiN95Brf9iZ3JmS21/5bT5uvVucfDStnSN2knTpaOs3vaFOQQdSKQZm9
lrL+Fi8FVufy8K35BEeBtx4in7z3hPsJnLTNb42nvfdHlF6uqCM64M3sdQfn627FiUeLxfmTbRAs
G/ra952wXvN9wbC03Nfk3G/4RSqogMhWGni84UuSUBUaBdrirKocDTu3kE5G+TyKYAyslEGWG899
QhtZvTSi0w6zUUn4Md5rdZu5bJGTe3Lr1wEbeN0CQcQX9EBXsnThUNpo2sJBaTmDjVs+geDjU7F5
ImhpNkkZF/QM4kswZgTh99nY/UmiWnZU+4AAvj/FDJPP1BXJPbTYB9c77ncoS14BIPiPm9CH0NLj
UsxDbpj89x8PQk9NVGOQXsh6/eDMj0QU8JCa1hhyEoEKLrGeJ5ZPOYwvg3LX+78xIW2DhumtEwle
KVuS7ANor7F0iKbjSUlbzY9H+e5YfdEcUUVb7tC2pY5y3IqdMnl0hu7agF81xBRm9cxKKih96WGd
0CYG9oNTSChFObMl9rxCLTF8njDNWdNtBH1ZdlLK7jZIAPo629+wUqwqOiqN8PrWQ5ODr3zb1KMS
isjIBzKxxYSnqxLzJPceJMWu7SCGB60pWIfctURjnRqllexjgdxbA83W1i+VOXsdg6/RhUrFXtP8
qNfm4GTlcGPGaRSmkxPXkk8lwlBUk0zIgj1C+8MwuF3QhkjjSLFL0i0IwDVO1Bx2HlFpycHdTlfg
tVyOJMAa1YOxkllI61kGibcS3ExSXaK+1rbDFC/lzcPpOWJqeWvDsW4xd++i/ZZCc75DA0VOZ+Pq
E6AphnCROtXyfrv6nhQX7QAu/8xDsDpf2q4mcAMhMmDkDbAQgdJ/xhwv8ZmsDSBANbNwrueW081q
hAFFnANMBwMfw7aXlZ9cXTCbWapHugG+/MBjwZF8iQb1h22ahELa2KGJ35cSK+SjYSVf9jEGFbS0
C99sDySJ8EsQdMRaTc7XIrTXI0HZQsp8AdDV5nc3UmWyTQTqmwCHwrlWZ8Mtkb5NJq5qP++2yEje
p+J8y91kfxFHGNRGfmCqIw3wgi06+DutwzKBM1xpdH75oMBOWxDmK/x44wl/SoNksqyWh765uoE6
R0UOEweR9l17lsEaCsoM839ZSCiUGsaldOL9Y2CRvdsECl7ihNkInJ8uuod2jUuwO2tu1aV9rdpJ
u4cPfR+CE1/mRvQibAEIqXv3xJK0pPX7CYZAdqjiHaA5sKZXhaOmI/LoiPY9d61N/hZcxRNzKkSy
iVSAn76S3r0QVOcIOn5CIxsIcryEccTaigVl1mUgbyGR3ivEc+tZw4jiuIz82JUT8NlILUgZ2Jtv
IMeDHSO7Qvt9KtzzAlYaoeQ7kVuvkwFbeQGG30nJSecwRy8+4L79w6wIOEjh/w0ZeA6AEymvpzPv
dsIEHphyGL+KzvAtvKcgm2k6UqXGqXccbUfRGysCW+U+cuCLCeL+PQILX0IEBC9E5lHfGetZShj8
B3l7vyEbCRXSVYQOEhWJoRpu35DTZ5ZfdETjdn1MrdE/SKcTyoviq750CoMbvvMbozTDF78fwQ2J
eN7gGQckc23jNwwm9KtcXMlpegOtY9X7SzjEWVAeNFlTTv+FNmQfLaXA6q5atbyyv2R4Ia+czder
Bm0PPzd3QG0UPcjRFfVGleYFi9k4k8EBL402HGLNjBLJBcvGX6gyGZeGFq7c7Oa2wO04NY3Z8mqX
YdG1FUnz+Scz2qA97sFUx9pVMnfI9rpTO+yRxZUbFJqusWtYCXR9lK92yNBZ4hWGRfQhQYLHuRpU
P6fmd+OEKznlkuz5W9p4WY+kU+oGuyhxyoiUftdLFqDj9SXdv49kAK/o2pIG0DkSRSz3SWsPGG07
7PWPWycqWgjieBjxQp7yzryfBng1WRnpZWrE14rViLbjm6FKyN7qhv8ohVNM+LY1/H6a1WQzCh9U
jV/2T74EmnkjBV6aGicbhxWTzaUAJ/+4C7/8NjnOJb46LFqrfrNUWcIrzCEKKkzKEkauiE69zTnW
ecwVmC/aUSIiNE5vnq9vkvV/UwOqp/Yvn7GgoaFyGOIhtAxtdy19UTZbACB2Ch84JBP08VAV+VEC
c3G+w01uu40upr+WUQXI7E9z7CRzm5dRzzRLr1+MzquDx69rZpOaZMdQ9VeFjCmfXvRggHN/Wk/t
k8cahBJ5otjEV1ou2DLzcjf4KGn2iDyX43WJFXN2OeL32pKdPBP2QlgCS7RTI4ViurkKvksfJjvY
6+pSsWhlbga5AOfliCIN5n7BsoiGynQcb2qaf+oYcAFsvplLKsmmbROeqwXR4JlOiYi3DPCakwr5
XRjSGY1WJRSnhoytzCskjBLSFDp9vW69TaFExJmhZLdYw3NtTuDLMmm8wXVqREdak51/xNQfa7m0
XcKSFWYTsvM9gHona1GWVqWkomMUK1kKeb4jTOIJaFuM+w5LGyARO9pZka/Pwww7HTWoaMaQ3JgB
+ZfNv8ZLYSzu270AwiJEcUTVs6CGITwbp+vyAzSsOVd5g3n+NqiCejDOvpE2inlF3lcH7hJTrWPK
hv1o7V56lPefTdlUg04GWUI99epL+PQPzIi9uETnuikYM5CW58Nr2MX6GplyiSoE+CmujzMsUGnn
gtFnod06NYk4w0tXbpowkajOjhavz8v41H/tDpIGmSOZLDo7jQe33CF1rsf+7+SBlIwBwkkDMBdM
remfS48r2G0VQPpzGHEB6OdbxYHPNVTRMIazuk0oVthUr6ty3+7gRYA2Vd2z3VO/JZLQLpEm4IVL
eqNXHRvpBVIYQ+lOQZJDtvl/1e9W4QhZ1JcZMpP597FDStFIB2NagXK2upCmyTxD+Tckgf40ypqP
gDPBmqs9C21khq/YWq7GPUZz5yfPoVcP4y+Lr24lLEZoDjI1Kxx+zRfFXRDD+faT/CBF0x6FTmqm
L42cPWuXTyaCAH4SdeM0nYnNyFYzXFpvdYdj6iRCRNZOK1n+nlvZ6Rh4UTMG5DaWtJnyWOE+xKQm
j15GZKmqoMpbxmi9Pbn5JpuCyNA4+FsLcnAr4lYTyuS0xwPUxdLWHn2O+tFhmOQcWoELLLWIeq7r
Bm+FrKBasgjIyhtxd3NyKxp6i+iv5uFFzpnWRqpx8WZvGhm+l8zcTHkbmhScA2AqwkpB0gI1VebP
YavLVnFsNXiHU+ifcJca715TO5PoORTCv7dr1Jy0y5xcZ2H34J96R+PHjfIVTGiyyPuRsLQvvpFH
QcXyQqigNKTVVAFRjuCJo83/eXMM1+xRNCFZlrNUKh2pznUo4gOi7V9DBt+Uhh2F1ckJ8AwSZtU8
vEepggI/uxNlpHvB2wIjR5+X/rBcgn3eREcuScu+Vwy+0Gb83SDqGkqG+McsihzIgQEYvWSS9xo1
XajLwbo4hAeXXC20XCfQs2fouIUsuxjFn3KYODt2Xb7BXlH8I+Kp5L8tCmN1rFyCt7U2n6HRoDIu
Odv0axaFNJUf9WWsfXCwS9AcxiODx58bIzLjO7ekjGbdfKCkAUVTXmg3v9v8D2sPCpsmw67mxJkj
NNm95ZIKhRwLVYpEIRTe1WryPze44NTHESw5okZpSlu4frOQPnhET7uR4T+E02v0ayyzA7kPqCcL
zfEllZ2XXAAo6rn7uI6IBcOu7n5DWMDb51+VuwUTGlHwvEv1cAhGkmHmci+YL9hxpX5F5GznDj5n
Ntr0WHIExfsQEsBDCWuZzuzXmC0iaRb0R2vLr19P+tMcvmViuURjY97oZOc8nezb29+t1WUZSnT1
nkf+1tWvTMQIC2bFQEsyw65Ea0IEqmbQk1AhyF2/0TphM1dFosj9HotOnkRiLVVPMhXjI7qXt7ZZ
GzPcGLNyR+x0r9Rq6aPng7PDvTZN/UQROnydlCOaXHYJdDS4TJ2cD1+IjorGqa4+U0LglFdXqo2l
VNnfHLAMLFATzchrGbDkTBcOdP9yCbPM3TKfyIImRIsu7sdH/Vzomjg499aZGTpalDRLOOBMP4X5
8ElgO3ZlGnW7CPqFPZpFVdw1JvmRF7o0zmCJzctvNFdt2NtUXlAP7q0oOtvTfJ6KKFfLaaz/m2s1
070yPvjVM0Sgym2OIuc48gm916W7GnMBif309iCZrmEWJMxk82MCSMmQo778zUT9CBtl9YAn0cvR
jQL6HY6U4NDzrLx+M5E11ItuSvfcFWojOeJYhf1ej/z5JcIsreDA8uS7geoicPf2ZDNrNW8EY1I1
/0QFE79doYSHNEPoO6/lpy9zU+Hcjq+EdW9W3/gX19JTki9nxuLAANRWGYRX3SdRp40N10yLxRqz
4Vh+yGa5wA6sm5yWBuGBbDUWnJvsK5lI35ioYlLLl9dPinn+bwHS3SZVwiHUzesCDQK67GvJRJtt
KJ5ootLNMn52wl++RBbFcz1ueX43/LMI1NZ+LKSED0CNRWJ9FlTN57b6ahV4C6uOAj6Ye4JjIp2U
AbjbyCrIuSXsxWWD0WEYpxkxx7deoGv/PNp+1hxS/jZtTVliuF1Uz+Gf1qedlhws/iaNOPYr9w6f
bRCbYoOrv9MHcDEota7oKu/Ax9T2p9K6xZgptEN5mBkomsNZKEVbRAOqgDvpy4q31FeXgMOZkjLv
c8LqoDcPHIT2SxqpwYbDsk8AT5LPsq/KDTYOqpraGHAepOBx6Owrd8/DQPPOla1+qNgguoLJMYfE
raM1ttqUdM6JLNc3bhTnPqypu/ZI6hRTp0Cgi6GZKmYGU0DacT+l4JDcjgT1/AkqA3MrRoZQFv6y
EA0TrTttajrXfLVbIImrC5ZGhucRCSowSLwNS5XVaYkJOlFgGG81e1oqZbjHT8i+r/T6EY3BDtob
rgMD5SAkgJyyXgIdZZb17Maad6PtLllZhuyZpmJDaPm6Dpo+sXbPjA6ZJDzEFpc0qWILxi00yJs3
f5XCUnAgkkO5nmQFJzOxQPmrH13Gp1p+x89YcYWpRiT+ajQjbPa15hrsoAO8h30rg5v/1oC0GkIU
KkGjTC4LIDPWJpVnuxaVHYEvpE3Oj9OQoWEZ8tnmBUhYEyn8xXyn1zMnJIKjq92ZTBGAEbJ6COQQ
jnmhY56xEtdP8UArGLaOQ3hSUtiFk5iF4jX7pppSP8UvRI+Q0r3l7UG7mHw+CVl05p2/v5n47Ro1
zTg2nRzND+6hcIS+CTLkcVCPn5nswu1152MuvHSRApcY795BB3kzmgPkiYeBGWtZDlgfVOFDysgC
fMBCytqt25JYLTZyxav0+Lyt9u2xj2YtbrGbFtsjhBVeMGs5WUqGquh44RstTMte5P5iavPjpcMS
emwCRdC7Z/ScsX+exnccOpybZavJ87AoWh6x8YP2KLwIpJTZXDyKGdzLukF8zVjJc1j2KQ17wUpG
/UGpjxB7nG2VvF3KsMDNEL+u/S6dTyQHdydkDyfi8xMcfhL2KVnLNt1ZIi7fIPLdg4y+2TwEXnCf
DPzg33HykJ6q+uqeOA7ex30vfqx6De/MZPC8RR0B3BRrtVcBUPneGgSn/PMWCmIgwME64x5IWHVS
+Xn+YenvSERu5a76zJ3MRUxBLep3Six+R2FvEIaY+ziFbg+AsgbSi+g1K9dXqY/LyDo1y+YQvezd
QTxGICfxWZ/pMorXJJ8t2zS2XSwqcyHb9wcYa4zOWSiIzpE72pCT26pgAnxtMZydgFo01V6AaLpB
xpfdm+o3YDvy9DQXCvcSqJlrmvSnGnCHTSsduM9K+CH55d52scT4rqfKisv6xe7v48u8rLp1KQkF
ZHy1svNJCGWbABQR8f5DQnS72aEMnw9MpJrm3EaugbOTxt1dOSS9w6a60k1pT/XcswddhLdZ67sV
i/1R+j48baxhZISovak52M6b+Lx3w7VUHDl/Dc/2V58dZVbWDbFklGNZ229x2VMpBFsPMxowUt/e
7DXqDG2quXc0/ga/xqKc/9vvDwC5fRbbrlKrwoBoDuXwBD47WUSV8rPQxXw0bdSI2QHwYDeg+siJ
caKTTiCI+Klp46yW0tSbyr7kji+B4Te0xToy6Jg5+iW/je7EkVtUBUchPf9O1UczDLLCaunzArr8
Vm7XAeis0bW7Y3PzIeM/SdEjGr6sQttAqO17Q5w/Dhp4xHPccUH8dY1KO6fHTy/fiUOyLjVWxIIz
XcY1u6g/1KkduQQ+4gSUNdXWKUhGCKPbH2IFc9dvi9cy9x/rTVL79+ZtISvCRlgZHhhBnLo4Z918
WjfODxit7YFD7td9DmUdKGeobzWwf+3vH1sk9SKVzHgffgM62AQEMzgUwNYMOPCbIInNsCUAYAQV
KWoVF5jntJ/AIW3cn7g/YPaTzdqmG/b/cOGD09BynKapdkegb/bItLfaIm2DxYFgq41PbeodJVvZ
Cr8iQQOov2zR7+7EvHvmjhqxZQtmdar4fwsic90/9HVFe9/E/XbHZftCqZSsyVDky88JYpscBm3h
tbTXrcoruehyggpvauoDjNlx/mF1gkis76FlI1KprOeDe/MFyKXVi56RTOndvejDXrhlXHbhQGGD
PmSSAVWNNCbBMMRcgRjj7Xwo9EEcjVmO2u6JqkdrpLBs1VoTNE97PfcTFDt/SvXFVnWmpaV9SVvG
FaxwCZiPVi/fYkgU3Wr7wgE6w3N+mI8rbC0gtw+ZyaIy1fR5L5nVglAuESl7ERf005fF3mYyWwCj
WrdTeMU8HID32ZNnINIaL8aAbnbJdUDOjQFrLznr6xJLeciMI8u/ah63x+1Qr4e4FsLyHfwPogz1
d8LEzbJqqPTQqbnCdeka4fv8ABQnyCZgTG4KKr38wfeEWEcXHU9ETu7gng+wM4x/c/f8g8HvFm1D
fhfazFVFWxdguSqqkXr56PecVDNPjpXwciH4QnTssBjsD/ISByX6ApBuinYFydMltGJXFqDVKZMf
7SyXTkS39ncmkEwgzyYfrgIRN09sANeGOmZLpsCvqMMKpm5jDabnLnvRwRKyJrviGGe8I2SAzGb5
FtYY6KCQ5K73H7d8y2F5BAaEGQs/zQbzmqxiJs9qmGIWL+zm6mZH1Ag0UUu5rFhjH+T6YnAwskQO
YIUaQoZGPGUJD2KTIGXnyW+k4HfKBqu9LEjmyrVi7guRmuFEMRbKpF2NL2AMhOkMrG5CFve7dX9h
G0YL12wr6Ajgm5fSWqH9NUfKmXzwNbCz2dkx9/OXPQZJxCimD3HipNAVX25zLl0mrO84AuUAqe7X
nMBOtiH5Xh269x9JNpuTtmQ3QVyivlZLk+iN2hanlWdZG2xazRWaSovSLwLe/XLz4+189ZpEP4fK
fq0Li17GWOpjBoxkpdg+knVIcJKRCy5Bf3KFcF7BESZzM6GFNw9nS6sJ7peL5PRZjCLtO0NoRQtk
mEaHNt8DTiRzbq/zwjXcJFD5PX+wtuqYimZRujryCrayG4T0g4KhtkrchdTutKuXTmH8w1Klsa1s
FJE3M1eFv14WmbUKbZid/6g+7RH5L/20Sjo+E9Vux+YnyyWrKHTXZhaZWh+92gUs6Jv7yucg/S2m
sNLr+0+ycRl08MYp6UAgJ4u8dcRvGx+3oJCRcrXgCCda8/IQsK3oScWQ98YSbPL65h6DZrl1y8jd
vtTDq0wq44AVxxp9WdY1WuotT1aLKWzfwsLfz62bEjhQUfPIRVhupMBFP3NpNyGaWI/73XV1jcJH
P3pMgq4CbhV1Bpo9H8i7ndxUk1oHkJ71BPNUF7euoI4HzsZntyCLmR6CCBQ4USq2ABdpNLlK457t
EWmuByY37bo+Ajknsc5yBrlJGslaYXJ/+Gmw8CW8vkIMJVGLcLoG5miomrpC0y9sAIazrCOVI+8N
GCMrMbENtv34Z+NgFdknpX+6yF9vzxymnu82F1NC0MiHeSYDZvESqApaUFp8IpaiuYCaqLANoUqu
0zucGggboeeELBQkFKtKcm0no6zEQVKJ8zHTuxQPsSnCpO1wVnLuMRase+mZbhfGADwGSqbHvjNi
ulb6NZUjt4xq/F+fjz9X0r+MaBmPR/ZI0tWPH+bVNOYBqRFK2spbDs6DI3Hee0UGM44BWoUfcwXG
izo6pj2PSk6om55SCtMLOAA7bcxPlIoFMp00MxbyBS6ho2rbIMiebLmkdkG7aeV0RHU4CofdAANJ
NQb/BeqqCIucMVu71Wl+WJYHfDdG/2+tXQrSgbw4taP4OE2Pu6ZNt67wiMxjDyPDoXBAG+26R+WY
dLvUMNGbtZ1IXYnQWwWN00Grh6yeh0HePGUApQcCimmk4ogcfBRvp8CDFYxp1rySzFea+3YrOv9z
sV9xzEcQ4isdfYxVy0Z8oYrGJbpTpu8KxOzfUlF2oOOJn8EP93E0ZxE42y3+WxukfQWPgdra95qA
sAbU1O1m5kBpZn7lWsRohrZXSaXN+9LrqYaoVe8zeCBBikKWf7DzZ+5h129AXCSfPXYO+r3UIOTh
hSi63rXVBEV51w439v9BokhpeWXbvJEXkOzigGZzWNlUq0gO0STpZeOZiwXYUyJBHOuDNm4lmESX
/8WgiUJegLXvS7yfygjvFa/GLVkcbGMsCVsF4tN3z/Ftlf/u+dQRA4Vwt1YHJJ3MK/PvMDMKvsHS
K1Eir8Xu7a/Il7DfS/SIQd9WBtpHTlryRR/xIrWUe+IEFpbDgja7hchvnoDCl4CL/IstBKSgiP9N
FOM8qNlirS9vVMjDrgbicrZ3RTuGpFlz1xngDgUgJGvLK15piM2IBDq2jj6xuMXyuiTN6IIQXlmd
33VjFliDK7fViNK4MZF0FwrOIQSiIQIiNuVtLNguhplLIUd7mDeXHMKcC1+CJosnASwEVQVZB9ob
bKxL+AsHuZMs1LxdlL4Ynp0IN/DEV0psM/oo/EldXYfqlVP2a7I6GrshbttRwZkeDvNs04WeBTQW
+MAJ1wbOa4lLJz1YhuYcY6+WWL2s1t9RuhY0MGscUKAFPUF0XSFejqWQe7DfHUSgZHMPHlo118nw
cD/LHMtXW1NQmGhKdZE6UgD81DQ93bTFoMuEGO/5tFVOEi41LJVp1UIU4XkD8VtcwogVT+6ql9FK
fRX++LF6ZkrXLOjjFjTKLbeeBXpg5FkPoyVg+xInbcusjVa8x/v8iLYZZH9PDns8OROobfa7oYoz
86wxufzcEKkEo4gSTPoYlkW4RwjBIeYBkK3UXnY7VoRJF4jbDrvNcHWH5ZAt+4IjYGwKihG/kT+s
MiStcEohB3PWK4Ii8lKRjBuOeMdxl0bsqvxLLQxToVyHw2L64vqAq6iJ8BpTm7McesV46IhTnI+U
hzC4HTVVw3VQh1rNNvE7/K+Kj3SiU3l03cfqup4zbx2aq6M/HziHwjVuiM9uhCz0MBqQFKRFhxKr
eTy3xREmBivkMySsITZvqK7buFGa76ZxQ/6/DhVrD3xcv47OhY+fRfW8sgapLQC+k5m3wQNQ89Mo
DOiSZpDWqjU8s35di3MbzO1mT4/bYDUeH/o00vKDIQMoM3v55rNo+cXN7RS00BnuOCWYIOPzoPaE
6y1tNjKX9SumnMft+hbnJjzCOciX15957HAq/8NwLZROY73ZlGCHCw1MTeYQz998mypM6edwv87X
Y23WZWf24jGBzWSvQyxXev3vKXkmVx/58Vxy7NkfBH1wPV7jZlgozlDWwD2szSqC4RfY3qHWBSm7
J2hqmq56wiq3eQxBqV4UQX4E1qiErY1SRNaYiFKfDbFNHYIfjGmTytNQTma8EwnGxokdXmGBNA3K
jjAQ6sI3aFsSpqBOOo5CsUa0cPCyBups1no22EXl06feydZkTTUvKZSbD0tZRF2KEdjtRI22JHnt
0To8j/eKLQWqaCEi3t1yN89ti3450E02UDsvU2M8rPSBRNeWcS4h61uFn+coJ54q5KZ1uUsa7OV2
38Dzf+E3LaIs6/xTjhElG7R3M804r5Ck01nkaj2Xvyn+D4TmePiLv58JGbNfLpRluUMJJxbvZMT3
e01e105iwyG8RBtXsRRwOAJhdGzch1B7M9FOuLz+ti2xlXua3cfskm4intVQKN+TsQ54W80mvPXj
ygAMdxLubJ6NeBe9BLaIlg1lfsQoAajDCrpGH2CAOTbJXCIAW93eDDyjqC0lxEpr0XybOeor00VV
ZeAoPeasu6T29wcdkRxsETTmwQUrGHjfIk5r+L0Aeyz1D+nQInONdp6fxKPAFjsAgcDCYzGkgxSh
UZVEcrfxAOtyD4jmcT3EdzZ7VR3Jsyg4QqRWxLrJ6uV5DbWletvXK7PDfizgDzd0i4cnAxAvMnij
BhtiBl3J/S0AtT7bkKgpaEZP5ZOm662ZdiFAVup9CQPiZ3EX5k8NnAJZcy2SCS9/33to10JCpOyG
zKFneY9JpPy2q/gr6xN6sWs6NTzXmGKxXXVmph5N2H6anMGgNS7/QF7dWmSDBnhSpz7EEIjUZLax
PpT9S2xCA9G8F0PKD861aJqIFaAC8xCfgdj0k7a3bddV9QmeSZCYZKC7bVFYI3yR52Zx/05TCB0Z
S7YtfoJVUmgSIXCz/HFnrrqVY/QfgrUsJQcCQ3cInCu/mDcIwgphGmbLSX4+0rhhipSUkRTrDNs2
ML7GpJJlLSiBnsw/ejtKPgq6f5tpj97X15jynW6+p1ciGF9IUb4U6+6ytedMjacvYHtlwvTWV/OK
LWa3X40ySgVNyYNue1JSgP5hr4+80dZVoUO17NJyz6sPb1e1UM56wY4SZ+VCDVBBGW3s54tTBrXw
wyNA34yZ7sTST2YJ9MvCdre7bSIDbBcyurnBv5PSTqfD1mnoly6pYMLTh4NBT4svNMCIyqIetVTN
5DxZuAYZLoVfAgk+KqfLAp1NIms7YkUV/fpA3hQDC6fJtHv47ZyJUIHVFloXGy7t3IRW0KvnKe1x
iMDx7lwah/r65PGfrNebQ6+n1A3lGltvYGXFurICxPm0/I+AKMZHuPaAgUocksAOJgk0gPpML1wA
epARXcfgaORYODleM/XL5Uwphl8ZjDbMQzqE5wjon3Hi2TVd4DKaqrrK5XAfWv7ueqHz2Hntu2x4
Bfg3Q3DOWqPWs8Qi0rp3G9WcGjeTC2Z8wt6UVsMJjR8T96CCtSOulRrAr18P0t1LMrSnsiybElxh
zbqGt27OdjzoVPXRetl+bqnKFBkY0gRIo7Rybuu2NMYIJJ7BKDRVSYjo7GSAxugMMV7TW6vtoDy6
0ZqU+MpLAde7MfdBSCcXAQ/sbOpfBqJZzRVv+jhBClVWjMAXYaWyabAco3SuyhcpfNYSqouWh6za
4Xh+7KrDpwTtDTtOuKJfFznDdSz1jePB0AiZ3dLoifkY9jz3n1uRP9HpK0fETeZTALWVMXfRLp4w
Kfc03PH7a1c/EWbkEaW+QxDgUthnVC6U4Msw41QiRas7ji9ve4Fr7OTBJiBjJseOu2cIuJCRf0uS
4dtR2k4TWyBpzZtON1CNApmhz5VWSOb2HDYymYcXqncQkFMAJhkEkF6n9G6wxvXsrMd1F2rVJHSE
AOyIygU4X5nLGeT0fgiTbrA0k9nELetAqXTSyvJkFMD09DxCZdioTI2z8sOJ4kqoCtGTb3/AGwUz
Is3eFjLuQ0fpsm7+jC3Y+e81STUg36ZQxiIe54zTdm7gPdzuJODpdowZkkq0dcSCIbC4NeqT3h8x
2jxZbHIYAR1a3AGaDqlr1UVqmLOjqO79wlfWmkmNz5BUEEMZQ91ZQOUFVG/cHQEwpaVEYZEsARQk
d12VJzPp3bQYug8K6M5BueuYQkN5eGI/zP0HMLnoinBBf5+hTEZq0vK9+6MM2suKXWyJCjAPNEOQ
NIzQ6aDXB/q+/S8uBGs8dq39VBJl4Mxc0j3lZVnBotPjE2UyMnAsylACARNEfO3otJs5jwLR83wF
ffFRxk1U+GRZpV/Sue6JZDARKQLYOi7u918kctxwsrWeVYW4FOlD2aEePjEUznrovTIQ4z1/017r
ReBOEia5QrK6w1dE1sp2XdTNzZKYtKCmwWSJITHmNcZiy1YbvhoJV5xM48AoyatgnY87MgsUZYlm
2odH7DKXSu2hATGlc1dJwlrHGlOvPrcuRg56BJIcUQmWZ36O45XlDWGn59bqnTnKk9exJovomwc4
sg2WNHiLHuWOXn7hrrVIPgoPNuknND3ySbBe56cTEIKVeLcnTjhwt94HbRR573UMx5lM1X+ODP6B
LbMQXzGd/uh3mmjMNe9vUMad/kHfsTFJtW2YgMYv9/S5/4bM0z2KY+2jLJ/jNo7Sn37l4vGUxW+A
Ub3JRFJy239cNIXzqj4h4gajz03/cE3mzgXDkLnu1JoQn1C3XXHRCz7cYSvZ+JyZ/ROhqqqMeJq9
WeIbkLOYxkGTdU5bu7TVgxCmr/30MYrDyeEZxugiU2E7IIgyUlB0Zp3hDb5ZgPM1yjZZjutohTyE
/LkRwS1yqyYNXBDhJT0/OOpXnt8tc0dIHyNL45Zma8QgcCh9kxLSPlABTTLt0/HmHxDH66ZKm+8s
C6e1jjGD37M+W29lPcwf6Gd2Ace26ReUMS985xt1IZaunsynFCjA6Q2tGNgxk8t/0fq5lcsdGQ10
7Iq88HK+X1jNDc8Ahzcnrv4oxo44elrRN+IuWDCIrU8lrcUiItciYLd4MnSRNibpnvhEpkGTOd5F
q2q9kkbQ31dzQIDJSePV087G2iP7tELnQPJK/CrUp/OGECwzzaviREgoFm73Evf+NKsdLUPHycHZ
SL42O/XVdRCVuX4iIZL/8hVw9rVBDQkVnMoqN+9fyRYAbzqaJk/XYQR0MNTqThG0NOEPbwCqh0Pj
kE3Tj4UotKZw3dAHP6hn8iamlcIu8KRrR+9LP60N0Z+u6HeCHoeD++EBeB9kGY2w9iBvrCO3sDAd
oqIk6uj6VwjH047hTrjqGP6TzQnHJXgfgPSOdwojNdz0+lGpkx/1wVUMOOUPINhKCARTryVEOZOA
hXYDBVEq+zY4zc5qvaeljjZBVgwCdmsNwb110oDlhDClHwRRCaM0PjKw7h2q402F7ZRmhd+ctcL9
rhx8JtHrLnXmRMuHiVWhWN8dZUNyoJgxmP0NmRlkz5vavqcz8D7wudAp3nrMtLDl6N8W4OAyA4dG
JwbO3FcEj+OHn4tg/iJnXZvgzbAsuwmm3yWpOhSAKPCznZtgHU3wLPzGu+M2wtp2ncz3wHiUJf/5
5DgxpB1Ko9KtlmkWZcoxTypspnnSSmsdgfZe5WgcCMgeGmVRlKmwQLOqKK6LeVRq8VcOSCevV3wq
xN5uC55cFz/Tmpl/AGPR72d7dgDaUv008dRzY0yLgOTR1eNnfkMj1LzX1dQ5AgkrRebjsfejaxZ6
hfx732IwkpvB3Mo1OUdbWa5hNtpmE1X0KN1/k69k7xU/cjEVfIUjwQy2AwqtxtYW1ltqYwYHKWhX
IWnAfbhcBVq267aRQdVBi8ve5WQZqUoTIw9IJ2kGWFIH5fctOla8y9WUcUqCEfCS7dhAdTPteO0I
DQYq44Y0DR+4WHG9EFlqegIjN/DqGoCMMKbUHQmY25HJZ0EA4r4LRDa0Etisd0dxX6w9VWAsORle
p+hp+Y+6YV3qcNMcl2jebzcv7llemjGej2+BQB1WFhaRRjCkwJA8rak0/r5gpgbaVxc4qMAccqGu
eHX2qGLHbwXTYq/g81q4T0znmGfiNFBsp2WH6Bac29bJ9lTyiplX/exHmYjjMibTrLXdszJzJpX0
/h/tMolvNlIH22CgRU6GZJPMCtdYAy7ZAxP4O/fYjwefCcnhDS41kVXO/1JakEo5c8t9D7+j73TS
KZ/0HnZnnxgMHDtLen8ozVkJBS2pOr72YPT3voVthVshVA5rvsVKB6daHI+YjWEkHnLHT11/6gHH
6JLrubEqK000SbUiMbrjMaamOdamJa7gGxYIX483LusMQ8pV01wk96boBL+NKJ1lUUw4wSUWmbwd
TIm1TatIaLBjhIf5B86jEdLiA2/Sdz07DeDLaI4Y17YogxWlyCWAd2FH7t7Cd8o2ysamIrb/O0S6
kr6rKo62fkd54tubqCrjQYjYkqeRpCgIV7JOYD5oMAUwdrNtUYzXN8b80vptjrmyfiZHKU80dF5d
wxcVLMl3+7gBHMzUbLmftjwEW4CMml24ZaV3wkA2HGxGSYHsTvjkD2Htb8nDpOsijG6VgSh4lAp9
Ospb2d8HnQ5+IlczMhnAjN+2tl6mBmI5tJhfS6zAeqd/XHUEy/HKwEvFk2WZzJfqjxQOtdY8EuS4
t0w4TWhgT8K9pmhaQAgu2HMrViSY8bjI+kgQUJNv5O2Z+/36iAqJxGEH7IOGWHVfsDK0N1jMoDj5
wR6B/EJW99r4mSCyXE2LuhowqNEF9kumLUnTIrrDQ4Tj7mkw41LQFK7sfZKFNs3YEgozDChMyGUF
Wl3R1gRKkaxSPKEqWSRz83IOEslYQ4ID3/DaP1ukPvAVYVcLccBwQs7+3OoAyLp4q9wmXwjfCLhX
ox9mOYfUpV6nIYxilh1q4hcOSW0Qbm30RZ/dNspSaGGBVx0SaKrETPwW+pgvB3HjLc7oyPs+H2Vx
BDDnLGNMWvFSkRcfMLO2zvxsffJ1RocX2dpZHHJAY1wIJg2W/k9vr9ZZI0Fd9X7AjbrcetC0SG8p
aVPBzj5zr0h2LvK7sOeeiaRqQw3us4UTQYpx/uuzytHAGP/H5xqPNiv0qYs1nBrbxR/nzy79Xi+d
H3mUxhC4ofu/ZzrGvFApeVYzevbHGXOxChE/wrwAIQAnUn+I6HU+iWxJ41lw5lxiJNwHyJ59jypM
fPOUF2uk3GWrsogmjI0xT3p9hbVMFpoF1LIcPlGJWgwujeQMuAZB09BVIC0jAYtjmzf+TCbi+NMG
EFsD0B7EkbVyt9LsZTO5nA3T2Gg/gX+xBbw7PX5D5nIhm5IHcUMuRBACK78SlWqF6jlhHpZIu2H5
iCqb/1/dGXcfp/YBs4+vP6IEpJz+U1AMPE3oCEN80ZT8reHUwhZJURXYzr8iEKpvn2Lo8w+/sW2c
/sgeCYRKRUwohmjY2Blm10VuDMusr1W6uFQdzOV+XthKViIDigKtJQ0JrdarxJccmZ5bVwCNwX15
W/qwxcioMDvdPAordzuFZ5RPyL0jj1VjyAJHV0ZIVvFbx1ss6cK8jmKlD6KzXVPPh6FCvszzvLty
2n0w9tcRQB+wEhmCPuVJr6U21hpEMJtZpalQXXbBLaYQ1AQ2T7u+uaazv/uUAtOGvFN5FSjV/xrM
h/gNhpZecCR+Le64d1nhcUnm5c6H3mEBwEctKU38TOgQpfvAhlTjzMRf9ooLXOhknXJMuDBCoyR2
FwuLbXezt1uz27QXcirISlO3VOnM860OaYykXD5BLi+jVXTMjG3dGz9aKqVQJSfzH9OrACUfXPui
6VotmvjzysmzHdJg8gEQbr4SvuNoq/CjkJBc00sHJYYq59KvceByqf9/S/S5bIdr4FUaze8xAExu
ofQXKAWJYMUrCJeo+KCx4i3DyVJ+hjpwpkWrMs4I5CErkOQF0Sf3Qn6i3pC5n3s+i3oO9ee1GeEY
VIv/kzunElLyxlcpU53wkPlcfLFC+ffbK3J8hLQpZBGRo6iH7BaW9MeoNQo6A9yADvBF4dN4YfRC
5yAiBgyenvUVqBT0qx9x49MCF6l9hy6HL9yz2SChn8SRDc74W0qrVVPHmgNnRGAPvDbKoZg7F2sG
3hTt5JqyBf4KxrLDFOJGg4Bf+QSdtevRpEzgC1OCtTyybwB/PucEiaOeGB0VMj4ttEUb/IGbK6s4
gSitxrht0b/fFta6oQOF5bbC2uL50rJbQBrUjJmGt6yNqaxX3GD3d3v/U7iUciBkipowUDeWalay
YYSRrS+zfJccJ2dzZ2lizYZAgJx1ygL5wesY1Ugndcvtxa3CuHCPUnbZycE6cU7S35al5IAPqTDP
/+hdCWwrmeQNPGfot8RBSi/l71689qsjjjVxGplADV9SXFCcVfXu7srfq7FbHHB2ICiSgy7E7MAy
QX1OLNI8kBkH1JcZsrpAzYLfwR93yGPU+bOiJeF6wbAhIz2Cl83OeYAiGQkfmsbTp2GJO3YPLsof
b77vt3t4QHUBGyfflJRArqnZpHIfT5UVqbCJ5a+BPdT1bp/xpp3oWPgXXG5di9SyW78cSkuuLfWy
imj0hSe/aRwuPvHR6g47cW1nqppNPe/Oa6mdbzgsJ4NGxqXgVKxMahzq7EK/vNkkLAhgvAYU57yo
Hk7lX84XIGoeXjjnfQvz6xzIELHJ6TlqLdJRixVja+KJ7tFPn2dXmwR/EnEJ75NBqgP+NT13iMzJ
VylKZY4ShpVd9Eib3xnKChnNXaM0hRbQVNgPMBNmGfiE98p1G/Ak0u9C3qt1QWQocnWmhFR87Qf4
q7KE4f3rNf7gtvpoGK44SN32OuqndaP4RKHSwYyA8wI1BW+qB/AiBfYt2724BX4zyGTJMIiAQRzW
2jwqRZGpvVu+FTuHFus3WDsvJAVOmEMt+CiEmWKwEZ+Ys95KBeLPdz+35zzj3syfaEUUh1ah6N0w
R2wcLvKS7wkwLrd319nuGR1F1n5IlC6GVE5n4DsGUMT7WPr7f8V+b/nP8jZue2WVXLA06wykcNLI
ykcZHBkklVogH97KpHYUyVM0YuF4VIuGqjNBupRSoVnCjmkodOLnmbXbjt1pXaLlxG1ooo1AkcLa
mscJWoZhnHws3Bsx5Tza0pimuWP4I6MYfoHRElKye1RirriPOqzRqYN0qVTkQ0ur+slEDVoYhkxl
wJBkA1lII/M3dMlgaqZ7bq2JVl2vBLSYc18AqmNiEghu/yD9QOFGSxXdB7w3BQqWEupqxodA/n7P
NCH4kb3KrUZ0KiEBBiWcSDGr0GbA+PCTRpcKexrbLcyL5sAFdWV/89QU/sqk6GCOxJJARTpbeUt3
J1yfugibfcjUA6u7IrYc32xGN+/Dz7qLp7kCItdQ1YRWGIIMvenoyTzzfuJ/lwItukoMFVyFhfiQ
i/ZMBSlpFpkoDn73c/AIaRvixyqldttBbSExZlJC4mU6QziZDmYtcYZIRwMTPgFzxGN5Zn58p6Pm
0H3X8wyVnMyT0L2yLmrS550RCqq3cW+S/npY/TNLete/Y7e/KTbWwEhMyE87NfqIxSzM2fNEjKGc
evlvmjFrB32YxMn3SDH6wrrG+QNVXZYddSyhPq5MZXeTiHrjcroHEhIOxMdAMEmsdpxyAVlB00rX
xabBVlD8J8PdDuskVbx8jhUcwl1M0RJ/KjEp8KKjdF6jXgPxAX4xL060uF1+0GUl0TesmDJQPxtj
8HPrapK2r2qSyTJxDomcMDQKvTIYoqsz1JBk08jkrJJzCnd/ecQwyVrLFl+Z/4Fbpdp58nPPaIpH
drqY6T3hZgj8VLToRzdzyz8IReZOkLeaJ0UCqbAeJUDZaaMh5hXs4tM1upQBE1W5I+OQQvCVkJ7L
fA7e2MScTCtx+lWhgkog32rEZnNGW03ajDmPxh8bSuHksvW9fz6Dso1Bl+9p62dRWYZiYRpliWOa
AUuguhMdFucpSeXhEYrVBF4XGXJny3/X4NINcc6YBlbe6bCDdoinkw0AhuWVcWRiClYeEAcACVLt
vajwx+z+PgGeAAgC0W11kLA/ORDccm86y5XDSbRVcWH3NYO4LAuhqhaOwgWVCtsmvpMUZgauJ1sa
UJoeyJDE+99GRSNZ68fIgDBWllKxHnEgNxj30CyC5CeV7J04hu2Ym8l/aFiL+HIKY/o1/i+p45mH
Um25assnmn+xSizE/QFdzOKc6jDJu5cZwbQ0A7oqjUTjbXgcVrDn33lp2+6zLfbTceF/cD6J+3fg
VROvV1VtGQmZMjZAXDocjy795F+hiAiJjxGZrfLZVRmZpmC3afutijiwUwncMJY7DUuuR+k/KgcI
bPpxj7SwLpNSpCcIaHj/b0KxBn+OgLuBo08kpCYVi495KcZinZTwr5CfeoYNETxQamh6zar8HcTQ
TkQ/Rp4U069v/Sl9DkIuRM/3+G/G9kmyljpEwYbsl7z3duI0Muy9d95Z6LVhK5wPqVXCFsxsGTWT
rJakd5Yi20F57MH5lelxBLIQjLvA/PceVZW7q59xmvAdXl4cppZh2T/PpbMENF/p02r0/4lMFTJd
miSxTe+TtyCl/V3HuwoDkKzY0x6QPpiTvW30TNc3rruJvtIYv6pSVok9hCCJRKozzVxQCmezxVYn
cmwamxAGjn5xFK5j8x+KNwA3JS9lsn+4hA9wVtzN32rTqCzBRINvu5jJ0nIyjklPCwiupNx895QV
CTJtx70wnUjhL+4VyxtN5bYZcEXcgmhWMmsUEJugpb85rS6k5Z7V/4LrlDMpBYSfWCjZfkkakvQk
IuNisAoOqb81YMrfsiUChJCPFgVljQxgiD6V0LFrHta9y9Ztx6hfX0Hq9s0DzKQuITYNj2C/YFS+
HbiHUwDchTVNliO6W+yqoKlLzhgJFyArsvFjof0v7riVle323jgnk9ZsC30we7L0G6E5pSM8vwII
N8TorX86gV02d/cC6gd5I1jeufPfCrXKwzF8rvXu+tJdSTED2ZqrOGc2l5kXhJpCazAe/CQlh8/a
VzHeqtuakRXenqvbX/2WrSS2/Cc2pDIJY1avUpU0Ghwr3y1GBU1rN3CrYQnOlbofKp1aszy4kjFO
6H2qBbc48Ay7h9EnwfoBTrDw2plG28UrHENGzsDqbhoo0rl6IN8TbfpzHk1PeZP7hTkoB2Wvizzq
ct8GtfB9aTAPyhs5CGsXzl8vLq8TgVGLR3WDKwe7KV194CRrMx+h65rWAAtaDZ8if7SizMyySNLz
H2sFpoyvpkjivT/BBXiqgH66Hy32uS0L0UwkUqYaI4OwG08cr86l8q9l9Q10KUzgTFNLVr+zTdYl
BlgvI8zFxhxHQvHW/yKJGmUW+ToU7PrevoNB4zpnh0kxe+5UJDWLPqtNygezrdobqRPzh2EfooY8
0IWKTK49hm9a/aCKn5mWjnydCvEY4jOSzj7jypvJiWo2o+Sqis1iwiDl/8npoC1mj0yG8f9aG7cf
Jv+l5LzbvQirXXqwf6jr51C9Ts/SFLIgAsEr9BeQevoDnB9lak3Yk+0yZN9LO0YANtkUV+w38xCE
JLt5vdRvw84498+ophgUi7aKmQsq0IwMB9mMNb8XYrBGj5bg4tRzOOV1m8DEa6JVutDQkGr5efGT
ORXsqtQMaBsZGzlsZEbcxmBzhVpOEIvMOdDGOhCq+LMgMAjrI1NIFi4fCqdi5R4yXE66eR6cvr2o
6Fnh8p1aqVgocCnHwGBewQZGtdgDVX1WZ7OAzBopvXP77b9V51w5IPSjh+q6e9WyVe4uPdZnmalT
QoGQMS5BMtWb8TRKF2J6K53FbxoLkHg5ot5GY9huGqmGEYxPz8kiaIM8HolW3g1W+mS4s+7QAC4v
dS2SLHUbb9ncFH87CK2O3ZvPYXRU6nDrIbdPULMVHKiwkWViVw3ycCXNmi2J/YmfbURRk1B3t+W/
A8ICH/aa1whA79pRol2a4YaQ738DuVRmw7r0zmGhS4ZepOetXdgHPAB0w7LAwP0iIQMwJU7TTXf8
J0Sr05G4Hwi0Mqo8QOgIAnT9Ey4cmvQmxpOtac0iyv9oZqAKdOSgvH2xPCvYbuyVLF67i62by5yZ
Af5LL+gfdHtbREL8EFeUvLvDam5Q5j9tAOh3Zm58FenujC0vMb5Hh+G/UxPiuFQq0fAzaokSZ6J5
/OWP4yVOf9Rz4pOzY43XWi/OvcL6LPfg6YvCu2/rHTcxjtym4fXuPGVtxphCFYbdZ7/LpGQc9dKj
OsPSOBLvHUyOr+oXoxUoL/eUyU05+e4RirTBIHJsh+iC33Gz2cuiAjUfjzMkVjxNq0Woxdt3EGaX
/Y6v+exIE4O493+yujdCzVHgPDvw/c4JkOsLCA0Tjs3SUROXawpNMHsqcMuK5Q895NG0J126Cfhe
FD8MAO8E3VVcgSNAPqaEzBS3wJ2hHpph94gOzRkKfLO4hnQTNpo+OUl8i4f3cmQ473ZeRqxgf4Yx
uch6dNs39UC2f+/3Z92ecTnLA7NzTrqMcu3EZoPJkf+2Txff5MrhJ4TRfV2Q6b4TUDHHWoW9vF67
3mwKy+KWE+Tyvj3Y1PxATsw2QxMrpJl1qigHG8Em+wYgdHlNAR2LA8VNXJ/kVO7T5RYt/gRvNZuB
cutUobFgOaFpQfCtTpRR8ph5MfZ5aPS3sb4OPTIFWKCJH8oWymJ+8uhcCsxhRBOHkVIx7hTjpYzP
xTtNorz5O9s98/W2ddnk3HNAFa8dc6Yj8izobEpEG3dBrtzLrzzlzJe6gCmfOxxhg8Z/GFG2SmmW
ZISQiVz7/Km5yFX/wRCctr1GQ1OfXQhdyZgVGCpY1IrG3WfIal1e0QqoRGJPSphHVroysbAH6e35
axlHzGIxqfHlllVV71Yk/EmtSQkeoLKCj4YTExF8kNXboOdgr9eDrTeaG0DdOBUmMsvHVQmyH7GW
9LhX26vXIVHKlt/4BcbB+fY/S5FP4CqmFIHCbKE2ic5ihPh68x7qM/8lGfPlzakXlEDhLvFaMnWA
gU+g8Sc3xjOrwQfWqQJPjut28tVKx9YHY5/hjOMTqlHrsg+XQAPD2/R0vKrepGs+TcowMzOqliC4
tWksLHmH3hD7WjPkJHMq3UKSpJupU9R3Kx647tRT7H1qNGyfhnO6Gfr5J8Xw6+fetVFdiGxmscLi
5w/pkiI2S8nLApJIzGnrtEK/owSSqeXjZqcLs+ejxk0RujWMkNjjMNGPcPIpR2mesYN4lofZa3ec
QNrWbiqXtDedTAxtfc9bqamJJ+bJcbrm7RNA601bOuQABhD36IxAk1kxO39aEDkRqb+Frb8iAeH4
X+0ltCmNpnmfCAVJQWwGvTKYi+w0wZdW0dyP4+/JH+/D2a4443Ke+PdA8xVK3C2Bo5ridMfMCNCB
uHzl82ArweRHSAnk+YAPRJm9cZImKZ30WgVcwxmdlQStNkGFyrKIU5ooVc0FXtYntNMj83QuqXpl
L+2qlcf5iZFgyFeYB0TBBKZrDcDzJWNuliGZRabEV67CB5mysjtXktglVY8B+s+kHRilEh+SReDR
Z+oGkmuwF7HYBOeOSTr3Kt6vFhTfi7tSIIfp9cvsnPCAKmO1zx77u8aDKxfH8nbPiDvVIy7oWe2G
2wBKTrO6XM3ycfqQtaCRjCGrEjiCGR9BIeNiT5ChTz0ZqxV0jqF7jErLj7AWEB31fdV48RTbAZCm
VE5d5y4J77eLwyWcfhV9aE2IQ6NoPQgJHD2KW3BeGpioWQh6C25UChG1w6Gnkad2aDtsNrXyHk/D
v7rkwp9FS0BGXfkJepZzTUUe3cyAdG2NEMSUOV6zXQ6f9wM9lojmdxS83Eoua9LergPUMvv3+TX0
PO3x1k5i3o35zlTRqWWtbbA/a+ZqkeF3Y19zg7Lc1pinyWgACp7Y+IiKHqxL3HDnKz0FCT8njKea
MlqmbTtphD0lKIjXfRdoFX2GUqQviQB78TnCDVYgIEJPgQTyYBpO8WAySt0wJWobt9inz5yxKrpV
zFaAum8ZVa9SPcggxATbDmW1+ccWswi+D3LOueUsltWJ25IF+oe1d3n7D+/t0l+x8JfLF3+h3lNI
KD71NfWDxJlUomrLqy05vMkztg52rLNo3eXh25FRriZilgbSS624T/mYiOcT0l1Z6VPr44fnqpDx
9kDylwnvFZZj9dcnSp8uyWd4U7U0ql2vffZzWAzEjQ8/i8XBrPTgemRpKLtBgzDmS0af0YGDyfVG
kXqyTdw0OIWaaxfeEDxYYxuwA8FIJtjovmS9AgsE2mbUr2Ut0SdLLH4KzK0eKf4vGeQ3KJKqVCEr
jBN9Iis26rXYvFYON70vGznHinruAdAJ0WJdSb348ukwfcGE12EGNxJM8DLyv6/U5d3RlNMIBLuU
J/Sa5BSsJI3WkW/SqRU7ZFPNdUxnf8mBUu2cUdaoP3RSCUPnflVJg3N2RVSak1/HbQXoriRsaXwn
Lla22ubmhyv/VsqcwFHCWd9WXDCGzGaO8wbu4wPKPxv8H8usS8SfodtzYjyGdqCAztUv3/BqIBpA
irRMXflHt42vVnS58LVwcfbDVsv3CigD2E38t+Mk0AJgwpdbA6ixVdTIeLxpixM6SdO/W+ih4KRf
FetEPwK578BVYq+EJ4IanY2i+CJHVqT3qXhNfP6sPCtupy0YeNFjwiREQ6anibAaxC+ypGXcBMBV
j6jq+PXEY1ovwzGktitNxHsVyMNmRUTWVlIw/If2exEwcNOZnQFfnVZzZt/G+yDNtfM/Jq5dkiLG
6XwzddQ1DYh81FA5zKc+GHHU0pY7ljLXv+SPGSjQ19s8cEBfGy5cwKt10Bgt5HCd+t1/mJooXJP3
HtFpz/HFF8VWl4NxXPD6dQWy/nUgktCN9TtLnp0+cfZGy3tGx0WHx8DtPJkq/dc5eNLSYD5Nnxfp
Zm5Mzovo5L/I65BCVlWMWp+6cE54UkZwCGVK293ugTKvQLFBXk6CuZkgQdKUQ4GNSI3DIfxEpj99
9vJB8d6M5g1bkdIqAvmB1UVGOxitA0hE89ocspgRK8WW+WkbpzikqMml1GGiKuPXxdhlkcq4yYFb
sRdw0gf37Z/iiGXFqUIMazQ9qxuCEDpkL/hslRsQ4VRP1cwHoHQWI31D50wBoplUd0RGI3o4acMV
SWomCrBN4O6dF1LvXNJff62D7EH/xlFIfM8YUVW9VKjJWQo6qBsBJhsPovTHylx64s0rRdL5hdSe
Z50jhBzCb9Yl7B3MfrtzIeMyYFPfFGwbioLA9PzP55O+47M8fkhODxSW5SXZ+YtL7u0434xIYqu3
R7Uxak6ZhnVuTiF3S/A8vONcqhMXHXN8NnWB8FIjicf6Vy3ZJem7GNeuI79HYA3QTz1YY3PLYLbh
cM4IBgDewH4ub8eSRON1jBCZ/yEn5KDtStM6KLZyRYdglzo0KFknI2oXWMXmMpNcBQJ3ReZisTNc
G5XAa9rBl3h+D2nzNbjhOhvZrBDMTg2SqSt82rYaePyR5s0Qk0FMk6aAJvjKxEHJbr/XplT4Bhdd
RI1qsL33jrebNsgEuFQK9q6tX3VTmXQ8geoRut7OhUN08WEnFpQlZdY9o9554es24TjUYkJKLv1f
hIbSUJcUoMYa6+PXJi3oTxcDMhAtPZLd1bkhAR23mydZm7cIZvLeUXqmk+C0caR/Wzxy16BD4E8V
xJG6VRWMHVLVGPShepca4W148sJ0vEZM5nRyNHXpeW3zxfFCDWtBP3hl4RifwGcZszEiVAIjMio1
RF//H65lmAZpFDw6vecv6X+O++HjxVQ5fILD1a3EDCEAHm1slV71EgzVQxiR4rEQZ3D19sfVzNk9
Fvrwco11egXmkzf+2SOaib8pek4yGwXVT34D+EkpbAv1adg2Uq96Lk3Gw8u6EuEuOKioyW6rL6n0
XSg27XReLEUfbjmVkUE1X2MhGdZEX5J7eldvRch+WnKUOf0MhUpFAqRhgWSR/uDIlgaTJ8Qwiqiw
gfX5qXsKdJ5XvqmzQUgbknsMwgLtbUWy1GGZjvTC3uc78/rwF6+AJCq+wwcojNghH6+exmy4gW2L
IbIZo1Ow1N2Kt8KSsuE+Hrq77W9cX+TLIiZW1tRT0SaFH99iUCB4qU/+nS2g4b49K0F0Gcx7CRy4
vDuNjph87NL/rgu6S1tm8rlkQQPPbYXYOcRpxEh6UJHY+F216k5dj1KAZ6vx5nkhd0gGeoXV1EBX
ZUoE4yHkkNf116iDrE0jdWBK4rMOAIDMWsdds4a0ASCf2Y6vFS+LNPRu3iKpG1o1d/UsT/lIGL0q
5VH8Nypbr9vvJTvwB6EOlBEF4q1gkQrblRyyb0FurY6N64+lYZM43YuZeNzoFRuebjqy9MlnwsH4
7y0f2DcQU82mLyhlZrmqqfep1MLR0Bo/CaGdybH/fxu2CGhqr58lHDBze9BkHiXJYQ7w6POFK/tZ
1i3qiNNucZxTmD2DQLIind6Mh+b8BhaRGjqWmgXJ+WHrTBbR2kHHXGmFdJ1s3jORH867JRJaopiy
BQZsiUPm+VHJ6QqnC+QEfhsVCqoAfSlZ1gEFyrky8GYqy7A00yPxR5BejR8QhIVtTp2IWq79q59H
XjwK83l6KIzfBRZgLX8q2fjEEkkS16QrOQf/6BduSe6o/NegOmvNPUQKObcLPa3jGlOFvo4IRNws
bNsJrOST+34CDOmYmvnpMJmduatei26kf36Dzo287tGLy+SaiD1E2nsKn1vKmsPbtjgfEA4F0yWC
4Rn0UhPQse2gtw1KXaJbae2aZ6tSLI6t9qRc9KBfEPzBpgaspUdkLLe9R5E8jooADBPoJEFKmMaw
vCUs9zMVyozRKLAVctfKtLu5Xv7JAR5TzkFxgrGOg2bV0sR1IIz5ZN9uYx+Mo2+W5ldvpwjxQcrz
lhi6tOUE3fK209U8+PPnwmkmsHw44vgY+zseBaYSCBL/U/e2s3qn1Dw4Kl6QXlfyfFU/QIA/vnQN
Dms1JcUJuBCmzPRfq8KQyJZvogp7j7kE6fegeCMA7eEtrnWsSeUjuIFmoKDCo2xSTksIh4G+JzLc
+9WvyFEow3xy7IHKL8xa+eAVNKD19mXxKd9pOwp+Z7+a09Ek6lzFXQdlTMz7z2YBrapZBulAZNvQ
r/QxXg8xRRIdCfeT3jSMtRfx+45/wPn7WVHrW1BYRQ9FAGf6TO6yf73NqndxY4A75iA1j73B4arf
VvjekGfdkGZ9+qYNRqtwNxbL3K+f0pcy1nuE5p1+AJEqc2rYVC57a7PZ5c/GxjG2qUHaTX2w0qQA
F3rGIQ+0Wc61Y/vkRU4qEtNgcOuvKy9LxX0yQbI3vT23Ds4CIxZ/MHFl4l4L+ddMoFzj0KI6XuMu
mQVbqLA9CuykRTo/pQmX5DX1ByU4SlxvXjZ6254fZ5LTl/rkPc3ytSkpTe0UVex6D4QnWsS97hAZ
FAfo2zv5YXAAI66Xo5CrpbN9xIu3ex9w14neyJelZv3YdmGaRvLkTZj2cOfin1B8zCKR6WWvb9f7
ghkvzYiLxDIpmwJhCwnVA0ghr3kaFMap8FAhdJwDag6K887/07H1sC0InJtbspOFqfr4Mx4OGEvn
CCSJpThVBuDznBlU/AB9waEbaiOcfUdn6+uR5kBJLm6G9mQh/xeIoSTxpGMu3rZjo9/5nnmIeblX
VsjF7bhavO54FNckeL4cLZLUjQazG7F9L7eJu+lCZVqT91foGzgCIrlV7kOcmoBc9H6zZkjyouxr
91/KNrcjcQgVuc5M98qa+IvXRvKtmcz7aAH29Bwn9vZRDUkDhRT+9GvJri5Ys/0OBf27HaF489fA
AqyqDXe8tvGTUP2Q/puh4JFpdHOLLZAaXgVJ2kOKwajihjisZXDxE4KQT1/m4tEbv9a+KQJEL9QT
xzPblW4wRrghEGJ4BPhevf9erepIuYVsreEKhULi7CX5yQU0q73lAm/582EFHAFE8NLAh+VA2ocq
zmGnCV6k7cQNOAFLd1jzhAXjXmgFTCigAtIuS/zDADnEn/q//6lrciPN/tPsU5ZHS74mC+AR/9zU
8Ww9cuQA++bv55awgvnUsXMn3J/vIhH/Mu2CPlP1T+OXhvZQL7BU3opCTFFNwb/HY5TQ6jU07jJ1
MLgVmpk0gzEqAnpRt/TR3V1iXuscnewFLx82xxk/33Gf4jLuVO1ltxO71TPFLn2XkYNNshIaUA3/
+4oYDW6pjQG+HI9H+MM27ej6GF7w67rsL/ndab8ytjQytf0WOAKbW4NXQiDK/oVSwB9IUfDSzNyn
XhP+r5KK0bD9NuCjAalMJFGB1e3kMnCnNH/iA2Vf791amybw2nenx8UOrBR9X9DPb7n4Jj2U50zn
UkWrarPVt0HcrGRc1deDPGwp17QpWEPZASUkZjSh/Eh4kOeevZbXYSv6I0imlJ4swl5xH7MYLH1x
B2rG8TglAxSoOzVdXP6bcQ67Isr5D4nATNnap1Pdn4atCsNlHW7FWIMSn+wyooz+CKdyxi/iCvnI
ZL5/FCSnLXPngZriqa3g2OU3XNQconqCfpc8pWg9dLpveqEWQ/cMGyZJUZ7FbF3RQjz7kMP9Xt3v
PxYhkxGLHdezVrdagmzG426TNf/eRThNuBbDRO7BUP9cUJ1qPKOwCmFpxfZ5G0+sa4a3ctYRr9Xm
ZKquT8AeRIeqDlstgSE9Fba6lv/grETNGz2S5+//NbEHKlCG0Xnu9WB9mMEfLlikkQBW3qbU7hVe
pY0LRpXqnqJkc/goixhfB0KTaNmMzviqPF29SH6Ia//v0JXGjb5S8AgXjA6BUMZZ1M7Q4nekR1ac
9btw5aDOsP/lxdR6V3DJoCjexbWIPYqQlTMNNfxHy9TEnoB9GDKhzYqcJfN0GVXdadA074d+PJra
liJG9dBxWC5ZavZ6eZ8UrctnzicmXWQ1S9PPdr6TFV9LvHfGFw4n2eNgFbsRDFnvnmAq9P0y+9kf
DPNRLQmS2sH2kjgCd4VciL2fCsjMzAktutTJ2cyE2szgwEkLlBUJQcc9/xun/lGQB8hGd7NetrlN
oKl0cw/tkp+7TbyPp5F3bIqN5GLp/QzzK92CvzCz1GGNzVWA9z5QKTU3A3e/fjAF8Sspyk0E3Z0H
6RSQrlrcHa7n9MvZst14koUk76oG0L0SkthdeZC2/ioXzzFTt/U1n07dGrP9lidhAmzIdIamoaAg
n8gnalstD/IhFnH3I9lWOix1Y8Fzem2s0WEt9fn5dVhByMla0PfQI+At7KdauHMFc18F91NpIq6z
xSKBJRbzcwwj33rF5mpE9LW5NvndPp0mItguFGzQu+zHuTUlv7be2Q7DmCP5bR/v+zT4OfdzJcel
stppsO4Y5lgJCLX4V0cIJOK9F/RqWJ8QanhbX5vBykNRPE9VwDSEhmJqhAUHQ3UnKBCy0yv5/yew
hqzzBoeZGVZDjKd+BsbvxWgYNbHjH5NA/mKCCxG281yi9KibUfJb4WgfR7VyYPrzRCdYwTaQv1pt
El0aE7LqrR4k2h1qn/hqyC3oEjawY0NhPwZjijfC6HqiD89auN5xtgAODlhcBJczyei5+LMXF3j7
CcKR86wDeKXKztBe26C6rTvzy9zHv5ROYtnFVcOV4y7KC/tL0rai+wdLHPxvtUvi0utKb6mxHLru
PSNpZO3Oks7l0KsNDALudvkjK/+a1KR1f3l1PpvCCExGwmNlpZh8dHlYj6tA4lWf1wpxa4HV0EUt
ggKigA87eM1nfVrnLFYYcsUcIkjjFbho8geZEUaz00vt4lFitAm+yTT4u44c6WtIPhIsVx10OV+9
eLeVJW6iHgNACsRaoW95iIKmNtH9QR8zjkdyVFvmJHi6LB5GPPkq0W393BKmssKF4UntN3ZKAevj
jy/SGFtFNd3NlT6tIdjAlp3aLXmMuvezn5xULQ3TsZmJ7nRCW3YfcOSp8FsyQ9b4lk0XrwikzTO8
pKXA2/PShKhndEiz38FAcpjU2mBA3AaSuUpvW6V3aKH5sFbXxCSCt5YABYNdYfYCsQ9DYTQqmHtG
qKSIlq0NhLITpnOQEzNXbqVTq0Z61/8lOAReVvpUBXLnCEMsyBiOGgtWjZXnw0Uyu08jf92nqIfA
4BY26Ht8f5o0DucPW55qJE+iWGr0coHQoPNe/Rgs+BMDl6jjGt/DQaeCQGFQH+LDwKkmal9KChyA
RFxyd0SMnjnKEdpxXABKhSTFHY0+2wPrz1nsAEstsjFrIjaSHy1qxVjDXH5sR1+3/AcVKo0vPiml
n7JtHNEwnX21IRfuh88PX/b4eoniNGpnFJSHs3bgQao9obSl1fX39SiBo6QR05z8h9BhfjBfj2Fp
ilGBVkyVtoOuDmMZ1WKJ+krPr4VLdVtp/u41Af8Et/RukY6jRqCYwfJcDneklbkGQYpjTC5W9Bev
Dplq/n5dLtK+KOXKenCUnKXuJGqD8+sTo9jVfWo9mo4xhy5s2Egk8tycRxv6vcDbfkJqBfumdaTz
kBxp45Y4EKrX6enaZxMDzpy9b33GGTAcc77HK8dli6IOQ9xzqO3lLmBS+ANlBax8waJTuNRKyAwY
qb8gQf+UAaCv3WTZBKztDWDXqBARFC4CyrRMeYmdBg1B0maMLvSLiD69jLVl023yYokz8FBuBQfo
+IucXnuWjpgKf0F1tDKCa0KDq/3zgjBJM3oHQ3iPnd35L5A8cIl6XBSie+mm1I5BNwjMRBaWrEpW
s2kW934b3vguBq9dL2mMWuflbKbasBzjHGCoGcOU+w+TOiO5sHr+BtWN99yVmn72mhUp+3j4UpzN
iBpbsAnsjOw26t98t7vVRSxONKAH+Y8cYGR5segVnkjXieUNdGMknCz2MjWLpLjYZovuqvGSIQWS
nLoLX2gdUu2dCRCZhjXJNgXZJnkpWGK73+DLAlQkTJ/dDdAOn2VNJ3mXOKMx0psDqN1I4F6MHFCv
yFRqEA4TDOgWSNpzpv5ZOxOayYZeZouh8hFjE7WVaCcHEMXQ4jFGVSGFyVNro63OrfYbnfeRBesj
OSUeQf79bmpekpgt5TsivQvZuPknwyuQfFKVon6UOSKmmgi2J6OBdhwV2eC2tV0Ci7sPRLzjAI7e
OUpkFiQXURzgiswXCQla/u/BxA5mNMgVuTjshNsSY8hLxp2bonPgn9ATKWZo1z3GQJpfGz9BDOv6
c8gB+dmeGbvcYF+AdzGXYm5nyxvoN1LWg3nl8BDuzKt0zu4NzwsSIbcatYghka7+ssl0Xl4jeNls
+VmVEhRRExdps0M6EbBCIffR70iN0B+AqAd0tg0U4FWeb7sL5Otw0BdWeB1eqC4oFb39zBKCe2o9
eha6s5uWKgYp+mQIZJlYfVMlYIUoq6sAF/+HqZuLaPYLtpr476q9MBf7PMFcjFciz4uavCJg7DBQ
+6E9J7o1bGI9doPynr1n39UGnV/I1Oq2AAA++kjjseftuLB5ubMQi/CrW3ht6lj/LpZlrVHpdMRU
EnQ6TrcYL40qhiNHMkruS54pn51fjyvwv11nPKBnJavYZLbh4meeGWNiBPe5IUjjwyhSm3q0MJwe
RIegVrfHxWZeYpSetSpPKpR4l5IRYJdzbeiUFbnn+NbiZEy+QNpkYc9fTFGzgtWK4Z8+NK+L+lfj
Bz0go+G0YeHYJYJVRWYSapPFioVMDG337XNX5lBnS/r0LBtneCu4BHdl75E+3UUgszmcmdTnL+r3
x4o4KRfCV/EdzUiw6rKFw5OBB6sDvgREtf7fk6/c4sqi87b6OJ/SXoNGOSc6xO2Uk2ukj0QnE9Gx
Q8VK9pssAbbHosplJM6kKR/q0+WFDDBGD13CKj4B7CVaPuWkQ4BmbdSHqP3NfNNBPBRVrJR5H7br
8hnJe1qomUVXBeDgGxvYwiK/CwSJMrlW25pjvw8IXUFFZcRiQwe42NOg8KTw3DTE1GfdptndIhVZ
mzFPvLgORDYMrARVoZt3cAzd/ek6R24WQlQXzi9rpTqLlpYXIHjxXQZ/tfIQOmGzp7JOsD4yN02H
rma0YUR+ANxNLPWNkcKCWEJ/hN239vqy3JyjGluum/WdpMIJe6Ui86djsx7PL/ZcxB4xW5uagpI/
bgvbhiQGgmIsAM50FKhT2aAKFrND+v4TV0LvySN28QST8P5VOkiM1kKgg74rlfAQYs0nrNSPyn8s
a20pP21p9i3KqM6h+bv0hOXFur1LT/rmbQKSj3H+jE162VN+soBsJ09qOVC6WJ2NF/tTQOqMdX2D
WTwL6B+A8rs+ES3hXOoU94Tvqi9ySX5u/J6N3BJbntKX8m10HITVZEI+xsCczdYM9U+ffXmH4vB9
Ufkex3I6f+QFw8osY2AUM2uBrmnXnPLUOk+yPJv7Phj3JG6IBpA5bvvTzrUFViUdczzG9nX7WwU6
JKyD+w8whqK9Ki4z40NPyMgFGJJ2h+bkync6Xs6qH/OBKCtbGN/Vmj3Bg7wcvzVWpdwFhVpNFNKW
4mIAMWo+wKVScLnfpJvSklwV5DVLvVMDuJdLdBVyYwDqajca6p9loFDIEb7K+uId8kOeTQduLr/1
gpGMQIIXQ+AiOKPfmknt1DpyFumvuQXlUc0DBWx7Ut+zwjitZ/NWlL72EB/AJIGKDQUccwxpVqhA
KPpHNp9or3kICr+LP2gS7/OMMvRp37QSHf3qpgIWaMhaKvepkjJBg7w2Qpjrtc8Ew3D0rKSOoNpp
JqoxkhawLSvn94R5piY96yd6pO25fHucJAeUuv5Jx8izyrZ8y2vJyqZ3N1vrCcweSbJreX7fMZa+
jGcPqIL9EyCh+rffszBFJXpmDTgU1v0zX7C40AfUmnYHNc97NNeT5a0YS9Wv/5kid4WPh2Fo9rne
H+WcG52Gu41ENnO6a4I+MlPrWiLyPGSesUF2ATe0+N1q+GdGQJZvh5vkgsl+O1u183jqwoAopRvH
MCTebPlEPiAESAAcv9rCzJ2A4Ax6p18QgtNnyNRSKUgxD0tHbpBsDa47hPDZ6pbkpCOnRZC0HS4+
RAvEL0QrLfbhYHXvPDNo6kejBXN5SSYTwrLlapHZERK6604y6OvEVLaje3QMabvsBesfU5GkmEkx
AksJnXY6Wy1MIFdqoGObDy3+PEp0R3B4TqU09OOcYfkOyo6ytxnVT8YeR3VJSqtTnwMl7HCSUuOZ
dF0UTYuL29N4HtBJpTaiwl6AZsTGDrFRCtaXJXtdNQMJUteiy/Nx36K9H0qXpvW5iBFP/iNHgcvg
c2hG5FoMKRAPb/TWhf5RqnbNGGDtJY6DlEj2ABQyH1y7Sz2cdZ6Mn4p+kLLDENt9wYU7aYzjwCT8
BwrUBciCLkJ/m14+pp8DuELGPAboN1bJDm+sNSb+XSeh/CS5c7waf4e1D7BXF2ASYle7T466AXxG
10bgoyUPREKTxSVayd4n9PVSyKeajSaI3apbzdlfKn5Fq3S3oOE8g8yz/kxiRbTp9KBoFDnKptv+
haL+mTMPbwUUtJvjJqA7XWUeMkqC3dSquLXB0LzdCSjuDyWH5cedc+Uh4vY/Ao0f9bFzKlwh9hKQ
J4SFrdFyuAZQctNmotrGXiWc/swpp8Nvaf7NOvySBD+UxaKPMc/t32zoLAr63wQOu2d+kLkqTqrr
O0tpKHzbZNhJRVmwmcOdih0zF4ygohbVBI+npMXShq333+j9XE0MNwlPtjBW6YTZcMg7za25/rUZ
hxEEPhEtY69eAYvpZV9UKsA3VNDgl2iz3lFSn4tV8lj5BOI4eobaM5ivVsyHTxz0TFW34cycQqwJ
GS0FWwnnMw1o4Gt51tEO0RA1RKB1B+cPt9HvEepR2ouW3dgYXE71bpouxAzmq04QhZnRIctL4gXy
tMkG3UYp5fqFE9G+eSZIygGzvbO8eh2yw0VgypCmsEOTtnOtMGgLPN+f7Q1tzIoNWdR6kl6thKxE
yaOWalREtZpkhKvr0tGIZDXp69DsA9ua2G9fDCDQEE22T+xJL8fwavOImfGWbSN7hD6Mi9gIQ2Ds
upmN3Zrd+m9F8Hq44M3+MQmEn9wUUs3WMfvvEn5Vq5UH3qgTM4774CaPsGTBlIEcas808UWZlbbk
8BpowwOSf+7GB61+8dv+eIbCc42YZLtgcYPkDna3TezCLF/CU7SE88+hkf9HCVnrVFDVRaUeZTEt
xz8ebtyw8cyNHW48dUDBu9qy/yqo5haTGXUBd/m7TI20h4W+Y7u/zqKuucoVp25w+wvC1T6+P5kZ
haezTplmJIl1T1jaxtqORosUVS4UZOeYtLQcymfT7FHIc3NE+Pld1OygL7vDzXSP/ZM+pIC06yPm
4WGMPuSiT5q1Ywv21NykGtoC/7ALendhGgJ67Mb8lI695FjCjKzvTXKUVEPbFu7xrr8NoV4Atrxu
U8E3cf3JnZSDBVJQHIguiW4VF5OD3iLURyHvufxw0TIV8NJCiSxpSRkR0yzx3WeifXTEEFTUlS8g
tdNv2O54slefImjJmUAm3eP57c+j4vmvcH/bDimOJuRHiYasva1FnUzlFE3ZaX7PBAvc8v130Jhx
4sbcEzuO8LeTxmF/jS9/P7lynazUHyKxdzglzG+m/5dxnlZw9rmaIbkFV3nGyCNd7v9JbGd4x4hr
RBUr/GEtT+lBfBMbbe49FdSOp/fjzuc9ZN2E+8UMnHaSi4iPjmr1NnPkaRBoDkGpe6q+HsFfiNII
9j+cVqXadk81TKWPJJIL+dp6iZhbYQdJjOXlr3EVECORDRNjNpWRG6HvbvaJoixiXvtCoKQmrTMW
8iMYitdkgUe2mM96grLaU6fxL2nJxPbIEot7ll4fbP2Ngk06yaZe6bIYKJhKU13ljK2nNYe7mZ3Z
zxs47DfzB5eQHCVBSuexg2MGo0mHgnG7a/jm6xsW9+H34HQATV/CdiUqqq+mGW2R2NFFsNNIEu2b
jPky98wlbXmiagfD31l1tOvwy8g6ytB/O2tJOI8th051B7t/XYnONIm31vRFXh1kwa+gyj8hHXfF
xqZhDCE5oT/d/Dcgk6T8CouSXXMwUi2Pc839/qWprYfxXw6ikavj26oH4XnCe8YStOktpO9huSkL
RlXl+pyhAakfCUgiYIKR7d59lgDW2IzcBHkItwRuEyH8sHfZI9OgvZj6p+7fht41feZXW10fC5AI
GwEENQXS5BCg25b6i0qKlu/oVJt/qjFLtyZaHxAbzqbkVM2SdrMtK3F8W0he43GByKOG+ub0e2H3
ePwnp2uwa43jAFUF1CGB9uamNvUThe5M31AmvqzpxzaHO3nkhUOwUP6lrfSFZm8iaY0+hDExu/Y4
I5NQ1emuc4goHQpy5o2E14/TOF3fZrKGzu4F8M8E3zEHiIpmGuUeO7b8NYo+Y/lxMV5UMNfuJBEu
Je3GinAUA19iRix7N8qkCyqIhB23Vw6k6sTY1fu0ZJVhfjo7P6gpy7leZRtCLkHm5luSpcx7prqt
VuBya3IUBV0hl/RagbctAuBbjKFhP5m93yuGSQ6k5dVlNgw1dmbHhipaW7gG7ov/FobVPku4774l
lCSGpfAug1TiSZ2hNEyZAhJhMpHL9MzDhqZ3in8JoX2fKnUhJ5Z0JCWqtisD/42caYqOo0W8O+/g
zHhgrjjhO2LS54PneJ67v0UvbYL91ftVZalMq4hlrTE5mI4lQIsyRXpF5pz8/35MGU4pV9U5rAbe
9wJAFRF7qnhrt65OM9HQr0WHeLizTnB9OeWyikRF4qfgQE3cqUPDuwSTK6wanySWyWIjRKa0atg7
eEDCbJY0mmQe0W0resgAUKzRLee+3Ia3WkKdWhv5K/qt5u6OES/5x8GUW8n6QJc8x7+IVpczAlgo
sf8NmMfCaIIhadzUdrrhX6J8hh0z1VHicPCnCh3j5MreMUUlp0iFYp3SmH/t7RZ2u8y05kgIID+O
HhBp1dJNiQO0ermtB8kIzYn3KyURetMPUHzlPPRdYrr135pmG4m0xqi5dbIfdLCdBPKXRIotabg1
m4fNhmVJ+QIfgHZrDwOodBKNnp1j7+Np/5gYuNfftUUwzosm4EoFDqvohY5jPkKgLIFGTtli+rz1
eszlzXXYlZ9brHYgVRMc0LJHBXuKtC/iVDrMCvp22sbqBr5Jgi3GhcsHTePiEnL1Wb0N7VlRec1Z
SY0dVmeXG7iHJ8PA5b9EM2DZcy8c3q8lCHd4HiB3P0Loh/mRxcsGiDhHsz8zIpa5pSuGMOypPydq
DJNfo/dnjYXMY4+hRZ+T/UBeEi6AZ+Db0d5j1n7zflhoYC7OrkxD+J4mH+Z5r3f9IUGly+rzV3Da
6M/b2dIiOuvmmd5oQoqZfcc8wsb/21tfvZkXMHhsGNWwRc/kzFVqG4zLRTzcXucdGKkq4+OtkpHb
FUHkhzrTI1ADnZIq2HOlJrkR3eb8Grg/enSUG61Yvg4ljTdIRfpmq0sTtZonfkNRghIAPXyYxP8H
B6wofVJezEmZlPmPd2olwmtZXxmbYU0OHf5MkX7xqFV+P9od4Fc8jV8mmyZxMD7nexYMnoKW32O3
BM3kpdaZlDASLX4tLB6LsGERwcHL0dYrsqDLJVZprlPnujR78rGvsaGxU2nhKuGZLT+3tml/U919
mbF4g/xGJqPUXibgyCHBZP0QdFA94Cpi95YbKxZCGAKIETc5p5K0LaR7Z2WGXwsTTY2WZZO93XkX
7vKdRWID5ZkRdDBgh4gHMEoH7GupZoBQEjPYdrxG6lL30nCFwHWrqSgHdMPqgOPk/ObMvepUkVC7
50pu9G2O+tkkwL1UjeIL7sdGCR9Idj/O/ztEhVmtFH0XXXbByE1JJG7U4XuxQw0ztkq+SJtpeobb
KZl2CmpG0Hvr6pLLMKlm8aJpT1bFJhZYEgWFMoNI0AiTQbLXsF4Cx9i4RRg2vFk/NudxNyg9Ndde
hc+4B37lpb7Su1tdm3S6yLx86pp9u9uu9suBvQ4VHcMaE4nlUdkzcNDNbd7GOuTtZ3GZ5CJaTwmf
y0jRJqrj5sap/Y3g7mW1HQC6yTPsqnVNX8naxTd7cs7ihnavhOMj/K6L+OUzhFll/oqTAAvA7cvj
dTkaTuzVCBO31GbfIMGojWxrDf0gtzMkiJmNDI6O4BXs+wzChSB23PagcpoZTTIGbJu/Su6YSMnH
EXm09bxetBHiOC1btbgQUBICycYnJFRizzvryXrnyW++KWOz5ZlW+fRFJcVfawsNf4a231pIY082
4meXYt909Qr4g67NE2Yy7puhu8fPFvklRs9TDkKWnPBqK4pWWcIkl4vTC+CNATyfuiwZJLj2ngbd
StsW7ql7obOa/qngt9dFMufri+TKUCFS6dlFxl7AOrrYBOEUHnvNFdyvrJaeYLzTUV6w/x3JsZUP
Mn+OjR2jmcMN/MnKwVUytQNsTqZxtCeKkN4FFS1CZO1n69Ar0TECTkQEminZalSFHyvdQrgwZyE3
XKbXtucSNs2+LO4T15/oNFznMFJLlxYseTv8uqGYC73t4SRkAyGFBL/suL2Q+tUEtfTTUaWMnF1k
tIOiQPOH+64X+PfJpNSZ6ILzAx+5fxlBeF29vq8FuXfSCUcvFQZRc6p7lIfF0DPW7vRlFC4oI6Ru
y2HTNtZaqArwqnjqA93xVQtLHH5GWkIuM6zy3q+OnDWGRYx4mw4stdPzmiAb7Esm/5y2TilDGSXA
ZBrSY1TOxNxJrZLtcRLUm0RfitVpmZMnGlvvoPN6QXHdE6oZzwnCK8fDFfgU498lMdYi7G0vAyiR
2pW+DA9mFeaH63AueykZyqyCELioK8DtUT77Mff/iMWOqV/9cc+OE9QmfNd8ksYychgnMIm5hwkt
IlPIiAzl91JfHg7n4tXVDEtho8dApE2YGu+Cr+ccD5PEoccSCrBkcHSfAXBzATBw1GWlCk2b+HNf
bn4EAvyYSgGNZakeGELbgf4Me9rtCa/Lhw7mvJE/BM3Gn8EhJXEJ5GO6LqOIaP03abph8d3kceAE
S3AqDQjd7udBehHiq4b8ZkXAVyS+yRq+1CotqHGLvSZrukbGQBT+TjmoSEbQskShHn3X+iXU9LsQ
b63trxtqmI08smpxSxUpapLaGjPBuTE1iy+nLqDiiSMpugoYX7wjToY0MC02l1ZstmPqfTyiugyU
o0IL8piU6DWfTfC1GziOU7/5sEwYvHnmSgUAkM3nbcb58vlL3tsLEztsY4JpF7cVUgFI5YUzqLyd
Jn2wix5EcjbDdMW8HyvJCTMt3mTJVFIWEJqVR70xz3A2m8bZar5fE+xd0OT2z1EBnaAS0zUDWxyV
gD+nsnF25yhNbYKhoIGLSedtZzpaTeLAePvIRZzgIWstaOMHKFcB7i+3S6/UkWBmnH1pBDKPMF8a
CowHyX0+iJCo3MaHKCdompuSBCV6cc2Krgoy/f5z94ab/TJ7knuNH1yzS7Kq8XWkjC89zG+r7XFz
JENqJj6vs/qh/pPyAL0y4lxV1WAYCGpTASH1NVHE6jElc4efEZMf1lztIWuPraoM6z0GAGBorAVE
ccDnGLQFWj/ByPAsTjnSa3OpOfOdNKQTP1xqz7zkIqwB/iOfpJKYrd/AP6zak8nxxw+jupQmWeLN
qgvgOSTKyBwnChIJZZO5vuG5u+37Oc7bJtIln8H3jAa5VHNcFdWm2gQwVfTHH2o+ZcLf7LmwIRlV
XXObluWIvW+d6xNO0ND0XcFm2mVnSlrwXTWyIG/gVJ0Kewtnim2Exkp5MoWphqPa/AtfasekzBoE
iaj2OCJ9Tf3QJxNX3J9aMPV227uu7gYdpVq+CfH3J56JjVD4z439Qs+1wCcN7QGPXmHrVAC/Jcul
fPmg2OZILAAYU90+ZCfl2gFMne2bRpRkKONCkfjgkSQ/56MKtNLkqLvo59CAHZYat/yd2diSEpXT
6sk7COgpwoVC5JULc7nejW4CTbMag+oc91+hpv49k/cyJg/N/XPEK1KW9WMK5ZLQwtURCKenRPrz
ze0Z9En6vRCwXh4Pld/Uh+3C7NlddMxE1OqDV1PdE75EbLEjEKe/AmiVG037ozmJfhA8F4IF4Dgm
jnaAUKhgWtUghlyXrJuP9dGzFPHqOBgIJkNeRHdsBBUZYG0R7xZxsNYpBfAjjeg2vdAI+V31SBBl
u8tIdf0NNeziAZjmrEQ+gyeef5tkS7YZcN/51HckAEELDmrVdMJZ4CDBZj6e/q4+SCGpR1ZDOl/+
B6hEdrd3xFbEj+Lo6KN6oM0p2clcVRVktQnYKMV+NUxArvs0kuXoBfikgln/l/r6DCNnMuZPekXF
rhBT3l8fTz2hjZZP2Ru7nHADXN1fTNEwVAHsfVMgTpYtqrAsToduUt6bdZpIpjg71IPv4pQ4hpWO
P8sMQqDVlyw9/q1KToi/T9+pP3xv6H8SPDeZpn4Opp5jLbQJQjORdiqJeX5dG2ScTUWi2cEf3GKM
nxSx8eqOsiI1kC6ZS+qOYbI99bysCIbuiHN7u6mbjJl9koyerCkPX1iVV6sL3DXMORC0vHzUx8NN
RqKfnITxxnAfQdqmRyewdOcvVEHemfwCoEa2QQQoIHoxyljy0x16qBxxaPccg1Qzxm/AeT8PJVX6
yvr0NebbGO3gg5oxOLHjyRjq+FOEZ1no4YpXoCzGxwUerAahmf1E5OYVvXWQujGobatbzB03uV15
uHLV2PpcSMnrw+SrSTrzAk3OVcIBPrLNNgDjkINqlQTJAVi05N8P22LUFcGX+rd9iP0Ixn/39w3s
xwIheWtWP0YrF+1mpIIp02ChALYJfEC0pq+wBXvNEYz+86/r+pdOLUSYl1wjl1dLPNFpFlXgdbFo
GFyh3CUNgjf9iq9lVTfUE3vKGyr6LBk+KNk7maSSFN1YgEae2zP89hg5EzOeCnL5H+7dTDryKb3f
kQwh4BC/fp5zHuco0x5A2LmptDebmZB2rEHszejNECrU6dhVdRs3kRG3CY9OG850Mni5Xcawefq2
8/Kfno1hkMZMl0BJQIeGLMq6PmQTWWTtZv2piDCveYXJ1WUczn4e/N0h15Fi6oGXIMZGBeNrYlXQ
NmP3Lbu5rKedPQqyeZvZeiT19xPiDWnjnpqWQSifddrzgEt9QBScEgg4nZ/0vTFm7Pf36qz7TSog
vH3r9bEABywwo7uLp/MTJrfqdkBnI0Fmn1+nBygS74MM015NUL4zHRD6TQgNT/2nGZVq+Bm7+aZR
hzQw6GoUztVDsDqFOPZI09evKzX8XlhPE90p8OXY8Nu7Fc+05B8QzQPON8KmjI4WFNECpgKFwI8S
5nGhHzP1Xa0XyU9+AwJjcvik+BIBBtf1xRzAVBSlr+2A8GWa66M0QqYvKwQmW+CRqk+kE3yY1OeO
0vDOVFFNZOv7Dc5F1hHlpDkMJxDR1hyu2Lxh3ZvqsK9R+L1k9uiIX4tjbnht3aUDxBGEdqn5qNyQ
xOj+IcykSZ3fttngvvqIqo1h2uj+WMloANX3oQRHndKKl3G/XodbI2J+zxjLr5fLXzkoXx80CfAW
dL5afbTj3vDnJijau/9bc7B0BwLzv9zXXXj9k0NvcqrfpHLGPW1OMnt6iEDvwpjUNX6ftjYwrYYr
H4HIzNHdvJVpiZAFRk3R59GksiU4dBMQIkhBsM1XeVmTx4uahnGnEQtakDFZ1BiCtdQYU9nlvTu6
UifvNwPWcdPgCTbJY9J0s74IrPWbtoh+qalH8o/zaA17aeMulpPr937t7ZxwnyLkAyjT3FFOI3Kd
BUQ5aSTxmbsAGCw2S+qJadzqeBUkCKBBDMfsLP5YmZgmdGpmZ1swNOST6g9xLuM5I92aNtkuaxYB
2fXVtTgHBcuCLpKfv6pZYZNsxzB+5BzDR6HUioB+IL/Vdsc3JsvRlMwG5Wxml4KV7+WlFgxyrhI7
KjuQpEzGY6r9G/HBOUdgdaqR8JtO0DMeHgghML6s+uXhqBBGBG8I2yW3Y8HDYzUOoynERt63oz2S
1acYmAqFqrjxDjwSh28LexytIDe1sVfb4QZ07RPAE3+8JUd4/edHimY/aip4p1VGpc2riXyhnzXP
WQ4TAF1FDGVrjdvi05c1N+7kgIPWEBvCvorhWyl9KnLggsMec/6s1gT1ogBBFVEl9P7+oxLGeO8b
Pdfc6IJ6HxqLZ9Zw+k94uWSdJO7ZA+SkZodN/DtuaSSnOELHIbUF8JLTADX7MtsP6nIO7+BdH6tV
dmD8ragJGOBrxtRfDOXIHWsxuCgqh+jd0nrwqoKI5bIMA/IqiHvQinQiJMhNeDkYbQJdG9wnQol4
a/QaUQ0AKM1BWCMbNZ4Tms/bg6JEvpl4BrPdZExqma/2WfWPZmMpbucbDMrmBo9gp+tfeolUTLLX
bd8d/N589mamJ54SVieuDJDVr05CklGgNOcLku67FdUJnTKa7R628BLd0O0U1rVyIjXFeeVdEBM4
Sm5xXV//17paQhoAQjlv97S87dL3Fx6K4zW5hSrQr12dxyIGu/RKXKnFk40o6vimUYYQXUVc92pw
JICgvQZ84kOcVG33hRALGGlPakcBywe/Sjo++UYop+QQ4SNTmtIepyMsUEVvpuY+DqnE2JSH/GyA
rFXqCUSMFhmjOwLcwAwKRH3IMch9TZxsvTx9678EFEvB4IDTdrFfwab2217TLPfkoiFJoeOPr2+x
PLwVED+NlG0esCDVHBAnbVysrvypj5y1QIj2s78ismaL0cmYbLfMb+QAINb/p6G31r/2z1uYUyKI
2JMicpEqTSWEjgnQFIH4Z3yxdK0j/PLkm80UJeIPSLDfTYdlAXV1KEW4FoZ/ItXGxfne4wQIO1yo
fYuYrxUPsF/ruXH5ptNb/uNJFy4l5AfzZypIZaSl4KHhZ9EfLOPGr9HQuNzjwCO+f/H0xd/H9Mwf
gI3tCs1eFy91Ayak9NiV3O5UkDdG9ttKOBBin+TkwQfAXxU4GZioXWudJfhWOOY1HcgO2eETc5oE
xCg6MMqq/Sf5/OPtfRl+faDAr4gWnnigPwrjzIAPmdJhaAuMAHYvZIBK+CnzJBaiPFrlEJnDdM+Q
/k3FiC02B5xCKSIwBSblujIGenN8wWreSkKnYo6CVS9YgxwXZmUDj4DF2n+f/ObW+hHofW/hCTCA
y8tuvCpdB734if+Q+4+qz2cz2/ArExB6rVY7wRoWAuKuXUDE9JHtOQR4saXTNkivG2HO/CwBMmu9
OuAsOR+0Y2Lcv23umOy+QV2GYbT08r3DG3fUvce7WrvibwfZbxMBRZaLPAGPZgy04BCtQGOn0nWx
boiR8eYRA9wli820i7xJGEVkawuvgrOygV35ZjIXFRSKZpifkScdLhoPYKiGvZZvWelqlxR3kWCT
AofDTjO/ICscKsOLUL9SoEqZHbHHev4bxwFYsLlepEDQeBzT0AP2HpZGJjm6CRLrvjyPUGSpdgpp
L32R32IwF1Qh6YvSsNcRxjiPDGl3hjUwJ1dR30oD4hQpNdhOo5ZKeF7OsAGUtPH8/BUksIwh6BIn
IHd6G4cLty3D+shGWHsQ6wGLLbJDcXXluagF6ahaOgwMKEWM/vjJEcHTFHZ3IQhn/OANYvkxDodP
HRk1vxjrRC/Lrr0M62yMAyHqXjM7MV2F/WLQgPywAvRwEma5uPZzhXoKm6nDNlHZvoS27LAygJSK
orc75u7z5i1mPFHvKKfEYMOolj+TeuJgQyC4TYbZ1ArUbkbJiFmE+O8j0GDkgui0x4XNlAZAJiMJ
bzUDre6bouH6XiM2MLVhXS9bnQFnRfZep2nX65ld4gwLPP+BwUPd644l473gjW/sNfj3y5IR4pP4
LqzblTdacy4eOF5awvzlsYr3oZTiD76EAhBVpuTmiKewHKaR5pEyvNXHyTtqaZn3cpZI8PUWbsrG
6z4RlbdNY7OaJMYWiSbLs2/V55wnPtMxt5zFv8tDK+24YCelA0yxCsTHyrLUmsH59b+sFp8VieZS
00hBnvV0a1Zq2RyYSjlvvi9A5CE20UZqrCEJrYG/P4dv/7gjhJP0rtbeJctWC0TsqrlE6lQdQaR9
I88fGIQpcGo8yZ08Rz3AJvxTqKfzwwlPvu6UEnAFCQCql2tn9dkixCuzLT23GWctx+AssCSrmi9a
ESMayZ+mzNXrFXOb3FSlJC2lSSFL3YnZN3NuMdR+jFVqEt3ePihPi7f53ejum3tFum0EgWHgpjlB
zXdNOFYJqfHkv2CpZ8lewKcrR6CP0skdEHJEzy0Ydu4ZceBWNCAPa9Tr1sgu6eEr8ZbzEYlM1uXB
jlEVgzfCacvaDLEzMd7RUkxKaJrXwaIxG8k+Fg7i6Rw9ahBKv/wpBpISZa7UO9XH3NbQg0gzlCPg
SrtH1PzxK+ddRdX+NqfB1pqN1kBwtfnNLpcgMvcDUTgDtXgwv4Hgu7wUJI3AwDTUR48owoJuPFMn
zstm4ly7Q0lGOZI1EKS06hJ1A0NZLOmdIwINgU5UR10djbD09emRJpXXR8jCi32TcXij5XFjSqJf
XAgf399qSImnvpZhvBiq+IwXiOWw1KIoUxe0PHoHnS4H/hzPb0MCY/qYEk4trV5rsWalhbTTv5Pv
hMeDJH7CwUA/RlZMXrf/gnsjI1WKAKjWTv7U0dZ6FE3nBR03kFBpIC9dbWPOhYZo3COeKt9tW1AN
73mx69OYv6psuv4415HzyFZ4kPb9IxSLMPDLjHf2txh2mNO94un4JqtJUknd6jKIPL72k4sa1iJ6
BE8y81VpYJ0SA9Xa/NeNJx7k+BuDQNmSJK8dfJq90dWCmP6GNoCnCgzYLzc4+gBDdBN7wpTBb9Sr
pkZqDxI0LFPn+Ao5Zc1I2zstVZD6yxkWEgRDXc9ZillQBNJFvASY13NLfzfilOfY3LlOJaJThU7u
PSFjHHAUWPASVAAEf7z9N5e6gUb91mXijGeHPt7RIcEY572pah4hq7e+0PEye0mxS4MbuDQTn2oR
uoTtipTkIjSsrAzVNkzPF5OuD2b+QA+WbXF5gZZYDT8eScNrinkvYt83N7ioJ3GVFcJAlk8KDq7E
eWIBDaBGlPsY20HmvERNrZvFidXJujkqcCFnBsuJp6gxGJ8eHvdsMVZcwne2RDzu4R6gomfnkmiM
prBYU7cwUVoF3RGugrsJ4SGHjIznOQ+dT88wJZ31dUD3CR1KpzIkorzlgVew+yqzK2CHU17ayWmg
izZ9ex7THof76AfdMBgFTW7hR7gxtdsW1IS/Rh2VAe+teKRXaX1d85GmgNcnFboLsQsykNMhr3kz
8qAiAGvGIcgzdzww7cLRl90JNN0zEzFQIUjjls4+KP9FMOeKKm7MeGJvI7+WFtQOuwuhhF9ylQMs
iz7O2tgm1aqgDKkdK9EtcvjBZVu7kqAisekjyhfE+DFjVctLgxKl8y/OoxRCNX78KUi91EVbpJzp
q2O44yHZEZw7MenlptLicrO/jbjtv3z+uc89n/k/JiDG4nitrBDZTHZoevGm79N5BhHta5N6wFmj
XORR/eHi8YgxrIus8A3APVY8E6HAK1dudfS0MN2YaEI7msz1BUnLfjlUbyNTQ6jIb9kAlcJXi7LB
KlobUX+qNGuOobgj7S3nkwUWN9JAHVzJ6f5GWFjO4wXypUftYXZC0052Ls1bdMRB9cfRstStOqpR
LfslV944JQYTLvW2TMQ2KGQ6V3hDaPGwcyCIbFoLrpUaGiDxFkQWDdhZy77+32tNxNLo9eqKixnr
8mGg947/ADFTdjY24Mq+Zt/ja+EMniOPKM5ylHk25OBVL10nyB1wPV/BJlM6yxXy6Ov2Z9TO/Y+j
pm/5B0jw6t8/uIbhhPBZ2oz4Tih0Yfdg+AP21ZbVZErfxq1DdSHokmdfPZXJ28XyYkQOFTMoHloo
ON5qZMgX3CQtVpPkRBZ8FxrS2ZhueIK3t+tDNFyo/H3bUW1G3x+pvnXKOjNM59OD4aJPbTDYq3z2
fjA32J6fDOa2+89jJnLIjbFIjsWlTgFrKjIjWdESvwSBKt0ZD1/9Peg2qL0TWxuG9PFNTUGQMWnT
FFwdfInWVAQqGa9t+pGJElD8NUAv+izNWaAva/uaa3GtDkTCaMGVwtOFG+E4QwVzugMF3Z5Pe6Cg
M20ggPH4I2W+XPfTgBgWEBHNZ3iFvsIrwLtvLLQ0ibWmY60060kedJiyfravxxbowMKFxTcahdD6
OWiz/BHz5bEOs/yF4MSnFRSWkgQYZdXAwUEPCttB33QkUUpjwihOd2zmBqk9583SIq4cQmdi32cJ
st2Ikazsy+meVA/mqyP/OeNT7ok58kdmfwUumtoB967dWUrO7XNY9RP8e4cXpg/lA+7yRAU/5Dpz
ETmlH+UMIYBF5OyVKTXCC8IrvZW6617OjXU40FvFz5a2EEKEkIOMKHlnynRli3GpfBCQx68coaBO
ytUvaruXifTfl5J/f7qDBQjqTfblfnZUVUJr2ocu0E+hnog/qBsenN9FOv2vZsr+YuqGjZX6WxA4
dfWuoIE3Fk9hIRfc4R6iKgGsK9y50ztaaa3/pXFhWZsuwXUFWUuQAa35hDSXzUVeWIb44ax3OdEh
174swSQr4uDLSEu1Yysd/Mn5Hv/sjroei6T4ddFf42+zCtiF6hVS2SFgBMI161cX3XWPYX+kWw2E
EWdEjLrQH47OO3uI4pZodk1ByFsv/mwUwBxUE2AbBrGBLp0k3xNMyq2nswGAv7+JBBtm+2wD1r3C
4IdURjqmndmnSyppBBeuoLw4VqRgVxNgkLmZqOvU/w+CrUFqk/72jm2DggappPmuG1hmNT6QRx+5
Id5oxQ7IgnLeatJwx8b+IrRW9ZfChBv3ajQC5Hp+EJ382n/nwJVfFVm2VrZGNb276jBSCcGP/f1G
UjSiK+vCxTsGLlvnzyfMDWe9x1lnWk3eMhRF2RSJSvEB+de/eU0Z//4O7zcSLmlrtp3roTna9W+B
8wF/PRdKfg2tSah7D3OhPxV0z7uB+rLVyHlZ2rYcF1DOpfhrnm0SzbPI3khkv4r1xcCLBi8zOufH
XVV2QECYR8GsAUmMkDxjcGV4BHB9Fwa69k9WRsoL9VNwsi/FJ+sVzYvJX0PA70WJrtXkquAhICpR
I9S33e3C4sztH5OTXsU7U+usinMIXmTXsEnDRBGzDp6bHK5mV2AOftmHZT9VOn7y6D3f3kZzgIyU
oNRB0oiLn7jaQqq2XoQRpJnO2vY3ECBGEypFUYELN0zLSe/maNWh6x0TQ/tB9K/aRhawB3ckQzzn
phEXUZl4j84oWct6g6cJTH87R5kQ6fvN0Ae9ciRbXRWZ2bXbV5ORmDx7zGfTypkUv1jKD1nhmf52
QEU5a7RbbXrXGkTG90SXk0jWskcaoI7YeYDBcXLiTk9gc+RnSDIEov9giTrCtj7u3iiP2Pk0iLan
lI3SvVd7zE9VZn2QGMq56aQP9fb7l5dSppuvVBnKDeHWkaiuh7eyWypWMDojBt/17bTNISSZEUEo
ci6UgmWAlmJuSt0FeL7/78lUY2pSfaOXccCybZoeBmSO/tWmspl5zjxjEa8RkCR1KRLv9kjWQsD3
stMZ0EZRA9YbSHDDbafm9el36wusmqAeeOtL5qL7i1Ts7aVzaCsbtLsj603xFtg8ooYeSLvCReTn
k5Suc4Q1zWhwlJqrp8xdrMLWW5gwGeUn7YHfjuUN0mJDf3lxenaOFYrzSLseyks1S9Aml5qDpZpS
XvWezMFHQ3T18aeCwQKIyxXYr8MWySckF5otJjG1uVdoHIcue/BAsWIONcAd2AFenBawecmFbMOp
zlpKxOhho6aSA0KTKHxz5Kd5tUMhjezvyGYnhCttEFNVhY3hHsKYMNA7WQ/otqahGvgWXDMpO0rc
WOfDxXf/ztGMiySCgJ8Q/O2J6ofxWJNIBwga7JXflGOEU//u/DSoYn6I1iipqUhk8sFAfla4Dd1p
k7qQNNjvp8SGHd46EkccvMjnEdFa+4/txJ/OXen4I48gcU3v6FBiWoHCAP016qW/cuV3dmIeq/hS
7Guadlgv07wBkEsA3MzPiq3ezRlJCshcNzuSpl6zoRBxJUPobepG9Ek/D/QKvrUt9RBnlASolV7/
Gw4WAt74w451zLCLDMsT9Da0pOs+bTH2xpYDK4AosDVk9VQVyUd8F0M52ZI1AIJR2CkD9Tr7hi1T
jZb+5ku3QBPrgtdasHVu5M9HU4aroNjLP+TWpTM+HTGF6v8xBdMFjImYve8AntkJnjnRRf0RIsqC
lsPpTqkBy2pFLMj5ZWxBVqzXfseAOhn97M4NhQhCTDV2jnVe1NNBo1sJdCK62rsyIWtw/3PEI/Ku
GdJsmvuVS0NwQvdNxxgsFUMHJVbhWVWvnn4c+L3dc/ZfT06Z6qB73GGYwVNdpxWM/6jjif4E3uT1
3hjJHxUVZYX7jLt8LDfrh+q0zSGctqLQ7NK2b/xkpHJaUASiwEQxUqLD14c+il3roel/BU7Ym7f8
J4bAnmMZRscflDyayNCTFphdTKTwl7dDemg4+sOoFPaRUKU1hxKt2qzicc9jdiKXy8s0FzSZ3NBm
awH7MV1T3kfQLL8pVonTnNv1iFRwKjuVU6rk2qAhhroJVxWx8cpS6am9KHyLkX/iuZoTOHNwAc3P
cHXAjN4Q2nqcMiEs1QYVkS1T1wUlmuO/lAzA83JizMYkknqof8FROlxdU6hYGoXaWcVPMW/vg4mP
qWzLK/YKU7VCzAnSD7hwMnRWDSI4RbXeJ1jwC/tGmF0x/I9bm8ryIBE9HVyUkysr7X29MSzZCs1+
nDG6mLHdb0Hk/rW82gQKvDYYehxHkxHJAof7bkI32Pr/JC3ZCxd0TSG9vBdxSRzTsTjJDl+2VmNd
HqThMAi2Ye4wGE4HnA6IeuP4+5ktC5RqVi+p5EQa4pYYqApfztv9rtX5uRcxCptLeXC/B+bUayfu
uZEcPrnAageznQ0/g4XuMjmbdlLgoy92CS4ZmFLPAGEPwh0B5PenQ9+DVjo0RpqVITEJ9d78D+ew
+DYPXWNuvJVrQPFwBfDCWyD8oMth2QTUbH/fRNHnZq1VUOAXW1hpH9Bz03B8hJPBqfkXU1pJ9Lln
g8QuQPgslwhvo76J+H1PFHNxfM+OqwUVu5K4CmienNSLb/JamC0Iii+6liMvTB9Lg7ILcWu0aN9G
A79uWCfQuvRLwXRFKYiGwnIhkVENRtafw8TfSA9r3fUQWrgFteTIO0zSue9QUosrgf6sYEMIBWV5
FRwkjRG0dB3PsoTmePnc9gQSwsrJlXWeDOp4LZmapYLwaI7mw6zDfLjI5fuwiidzgtSBIoVisht3
LZeVyCKpeF+XdI4b/A69xkbhNWTE2TYfDrkBPPjV+6GpCs3j6emo6qDYrqaLMYtgP9+HLMeqFWMe
JjXkGFkZuz1wrcxap+iuUIQBK0gcGg+qq2hzH7VSaKRhWy/am/XvWybmZ5oYFllbPz1CtJI6K10T
E8jZ4Tk8fgNw9XuZsLitw+P/0HrjTgI1P4Vi570KpBtdDNs748BhGUSr0SVF2ID+bXGsjJg/QHr9
scZmUQr0tBtU0hZDnDQQWZnlPnYcY4jwH2CFE2IPAb4lQYPrlmYeasgOf4W5WgHzqnh1MrLQ/MOm
GUOu8QOpfBhbET3YxSegaKK9wRkSPyp46Yx3XaKEdlSpbDNzON4i3VyguK/jvf6h6TRcyT2NdzZ9
qPwAk9yV/K3tWPiqGItC+zaIBr0cY0i2zCM8e598EbtrRpN3aLmUnhH/30UgWKTTE3k2U4NH7aMF
b3jQo8xcapOCpFhs842Kpy7Xmxf4k/Zm3Sq5SnG4y3gR4W0HvKTBG1dqI2c4NTD0o/6A8oW5l12G
5E6nuVXgMzbE1jy+CGtmqji5ce0eC03g8AJFIfM4hOFtClJimsGIBTzLB3b6iLoRUE37F0GPu0TO
WDUiQZCY6EWyAjb5v8jpIyiGgbYOY9vcmtP3EFw1cRPO3CZYAxd3YCm1bq/jK5mr7P/qi/JxUIHu
MaPigGnxAxcMuDFdABfrck5XxJ7Q0pFfX4HXEMwNXlhuS1NtLugrGmFy2QQ64aO7VFJH1fDtkt6T
4S6ZQL349B69I0h5FfcZzMiDUnd+hyi83AqL6k8Bt6Yr3c5/XDCPRJSnLmKpcp7yuAqnbqNuJgBG
aHTn94VGuWjSiIqpk32kUbWEorBJRwqoSvfdsKMQXG/WnWdHWyNwf++n1de9p3B2lv5QYNH8Xx9C
vwiiAJnLuiQjErI5i4X7l/pLhXheAQ/EUzTOgAY/YUcFBGnKPekoiltCCrVZ4vU2sC/2YJ/cNSm0
iRkPby05dleLXZzaGr8d+jHFxfi3DrTEpa92COloov3ely6tHfXIykeYG+3/Ho3hdeVpTCYxdQ56
lHhSqI3K9hkdXTqpkkAVz4PLDonchhkQFDaHnzMq6VAMBfD7obY192p032t17s1TZsSAOkgyRP7f
ndCDC++8zn/Ug6X+hmW0oqaq+LlAV1yaSkTJxLiga3ulhV+eKTnrVycryG5utwc4iTEJ4JWbcygm
hxwNzpAZSfYl/Rx6tAE6w9A1A58jm9pDiEgkEjaEIM1u+MERHb0mm9ApoW1eSg2uHdx07gZWss4L
koGXAmXUPLIY3kqsrThz27/R9L6281DyWcJw7y6vatwsoFv5PBUW+9GxZj5YYWzDzrF3WWzdjeIn
AqHtpwRt24Ad2SVy6V0TeRKFjAHmx0c+VEWmpFFTuJZUNIaKePSZH0SOBbKBe9ewArL8WEvCmdex
JpgQNzzi3EbdtGNQvGiOFLav5s/ugAXDwawEVCuKFyv7rng4fPA2ifoIVRy9i8Cbhpu7oXNJ2HcJ
uYH6zWrnLuP628dSRGHzPLp7BPrDC9OT+O/VUhfpX9rUpwdsM/VoGjuyby0ha/wzc4owfGF8/3WK
eKFUSstHexMOYEKEU/8ePY9j+xnYXiAfK9Nlya+7IMMcnM9UTKJx/DsUbh+xJV6ljT/CT3OTLnjh
mlmKQw+YL0+NZB4zoCzsb3+11krWSIOQBNvgggIQvOmY2cUTOWfgAkUYG+8S5qkdDysWVknvEc1O
q7GGYM7/a1FTgDzcSWJqCBqnzwbNSWCcKPW7oRS9gMN9NEU+J5uYqQFlxbvq+6jXvNn7mkcHPKXe
VTT+81cMVGipIIO8jlJLkrG1WsQCWIZrdaJxD0FHre+9Y6VNQPMtH1Y4xZYQ7Mw8nWMQAjeRpaIO
WBm8oj34upJb4DpkTSTWOIMtMy+w8qjj503dDarAIxb6c8uv1lKdsJA6fr5jmmOhi0gVDuxC3NLp
+PCOQddjwIY0zDS0nyub7Wrl+lm7W0OyaqFAicVDg8dJ9tHa83IvCtd8ISBHsuwyVJ/NGx6rdduT
HXjUr1myI9F0Au2usjDuJs4kJq+z2ViPgu4Ba/nvMyBlMwh+CRhz2jVxI0joDIzNbQ4HmfgKaMHK
ArK1Rs2GdF5/gNmH2rCmiXIHVuUjlNSm0SJCXuwWSSjKISQJay6S14OPH4SW5P9tslbfPm36Fkja
9Em+Eh6ltv4S4EX1rEvj0rkmPE4TZnPONfdyo7aW8armHNQwe7CLlwBnRPLmBrB3kXa129VJJsDZ
PhFDmKsiY8Qo/q4S6YWPVjAYuLHBjSu9EBYHDHaLM6pE4JgdyR44r0wdB5wab+AkQgHJKrqYHFYm
PJfYvTBIKD+IsXugV5d8pLLuliomaK1eT0snVWOt93M09boXDgGYoPjpce3/rRq9fzCPIQSkROWZ
6ZX9gYTZ7EymHEG6tTf4eoXDN14ROscipy/1ye/HdcWZM6ZWeDiZUDJusT/HoQZElFoZo3iPCuIC
4odAg6KO762H2Rf5Q06YCgy/zoFEzqcuEwLuwWxwc1RCc0dH1cc4kGWqrWVFv7OPCnhAlYVd9Zbt
2cbijy6UPiLCUTeAGCn8LtACNsF09b5YqOhbM50apvkELbYwEZjxXCZI3Zw+jvwCqvWqAqm4flLa
RMg6+G4UseoL/wxDCPtYvYPtbJ17hm6mazy1WahuXMoHyFN4OXYF5ef3sdwKi/ABxUlRRUnuoxBR
EM5Z8KHmhZDJIYzEuSYxyqrXqA48+NFrrLP32zD+ukG5BwsGeiBvcR8MCUD9wgoibBUYvHGWc2yu
Uc8TnZKSizvvWquNexl2XRDwAu1xrav5BJH5eEnPxmdRSsJInerS94fQhFxwSR265d5ybeqsBO6d
km5HeJN2gkj/+eIWhKadxfZ14c/DMFVVc2hFFhI4jd4O3kaCvpzqeoCUEn1MHPxNq4+442eLZzI7
AUk+z37dw2cx7C4VJbuTLuvhXnRfMfWpGauqZsJ8basNZ+W8bY3tLX3W2RwiQXkOC42Nf+M63M1Q
nuqGp+TCETjOTSkZeogSj5kUK2SS/frZNQ7xidfM3zDyycfLPe0aQYVnAdyuPC+AFKMKGCYmxrP3
Vddxx/5CO5jL/Wf3LZ4NBdHb+6DqQC4eYX+F88MD1n/ElNz/Dwm5R/COoUUdFw1peudP9VVR+GjK
8wsmipwk4i+G74DLll5i5kmLE1uibjv91Nz/QIhSVwSyQ+XHpI36taOFo2ZAkCrRFWdl1obmYlNP
aO7qJMkft77PyRR5d+DH6aieWrlDTfjWLiiwM0JjcgFnSibCTeuEwWjqPjQEEL/AhemorAMOGdhw
aqUU4jMS+S6beEQioUxMriO1rFUGlZ3/haINbM1CNbne++mFepW3ykDOzcGcBHXcqS7lMnDnDFG0
U6ihslIPke+1ck6v4W7QKxGQ8WE7QbZzgawraDguTvqQ6g9LTdHWA8Sihi4wlO8EpauQbNBBPxxr
R1dmbw8p7Vp73S6h6O689/9yq9Z24beJsT5LJq1a3pBV19ZMb0BzQEpDGm0ZOTePIJKdGnA6ld66
PGbaAu2PX9hHa+sNrpx7FH8bLJ0seU+SATCHFu8YZALJHvnmOnq8zFkxD2v9qP3EYd7+YaC/xQY4
sVV/XE7bymYiw018VkC2dSSiRzs8r0wQEKCm8XW1Q0Mw2dmYIcmlKUgt/+VfDoy4E6oFJPTls9MG
3pvRvD1UoUq8071fpLjh/STRA+6lbNZVnoVhL02N8Eq6O3k3euCGrrTFuCw4IwBd6NWTk26mX3Fy
69rxIOdY/VyeZmB54wHZ/W1DAxq02DtYU9JSorSu0Rsnr9Ew/5NEfpZZkPLLlTLyEHCa6adMGz/R
q4hhpJc+5vY4JMYaP0b078TieuZJ41EYgoLJd0w9u64Hm3yQ5wvvfRPxYYLrKyxa6+LpZBRttOeu
YVM9bc9bOIhLUmaspNKqhCgfOtSMyeKWSO0FM+GgGhRnmK//DtQ8vSJSHIOdRJXsvnNnAmLSBDQS
ilLsUed7VVNUfx5gFwlygMLF+jfC1z7AMloc/VHrvPgWZ0afRz6O+S4ZDvHv46aNHMc1zcubKLjD
eIRVoRMGNYslzzRTinv4cuxXDtzeF/zqwptRdxU+AVBvqGadt10B6ed8fqGY6EGyWCeO1PmWknmm
usZ6PJY0YBbfh3yxE2mUHEdFl6qYsSfIqVfVrynATi+q2/foF15eimyI/Qkm7aOEGeVuDkhfCgyh
z8SouWG0IDTyhlGJIXwpNjteJKxvRgzUtF1vwgxYrGbgXCcNnDHpHi5D5fezhcwu9lD6epGOOAgF
PNgJ3r6a9bApRQhQJ3hR7LvsMpq6dLA8gb65S+BOyIg+Y277F0ezoOSOeust6idXzWfpgAfuhBFw
1V0zR3vsis++ktJNDWbAw7uCT7MKkHf4wCqwH8UqVTqbN/M6COs9yQ/Fs+lVrSdlu94xfCuEM6n7
500qsOUCDVsO/BrisiYEelRS5ULSP8r/6M7ijE44O6lWZN+a86LmFNnETSJL3SJ4Kcb2ZHU4N1tn
11MFabioe5wIfZVBeR8fbpBUYajBnlY89C3VOljhvRM2VoDD77TlsJr9erPY9JzHbYCrz37u5+rO
RWjdf6ALhWNpz22MXvnaBZyeh1LJZcsPZjiiROTBIf+7qutWyPQarjXvx0/AEUh7AQ3c1VUCj7YJ
vTWdd7dcWj1/hsOl9r+mDOh6KA7LZ1yXuRFnwSchdGO36l6fOCqmfqnOeMyM+ed7FkhAJ+P6SH0k
BAlLJ6KFonWfO1luKXQlqMLfXvR3t0IeZbvx0Jdi3LOPDgkK5ehMYeqgmDnUpx6edfPN//OCjJGq
xQcDbnwbhLEj9FRoabpPWROb2u/Lprt/Pwf/58rJyeYtJ6a/Ub+O0dt6p/k3ped14erJstszpVk4
Wi3U25GZFMZnAKictZ6XULxjAghJeXajyj42nkC3A1zjrxRUPJ21wM0+jNaVCz1xds2BTK9lq9Bv
bLfQgCD3LWB7cKGg2iSpo1OZSeMQIsfc5A4XEtl1td36ifQQhtvy8TixgaIQKyTxR9JJWYCncp8P
z9kyugvayuwm0YA2ZMp8wLtzXMwaQsh8h9NMX1XyALjphyjo7Zt6lRk1P4DT8UIkplmeYLS8iJW4
SXHLdO7OunMeDvHJ3d+4kUjwUU+Dg9UN/51IPiVhv5IRkE1qFdsC7qZp9l3TkjLkjVtStOggGngd
u6MEI10iS6zFoygE5Jxw357yroANfDHzJ+GkgR7B7TKUsvX2MWqZD8SlfP2wKuDJNTLF7fjDU9C0
8FstsJxkydhMMPL5CYV6EJE8XOEpICOO6AZqYZMXWbJSIhovDejbuWCQTKxrRT6S954wDHfP/aCC
pW8eicnNk1d5546YZIzPVK162++Ve6lQSw5ZndGgRAlrAlayMG8LRCE9KhQyG6C/PU+GhFb0tcW1
lg8I4I5YaqzoE7nW7xhL53EqWdMpRoZpR8CplbcS3r3tR0dQNhkSQFYzyfl3byR1cjZ5hAlOQg5Z
0HFDlxSZCMAOXLsRCnIBGwkLIsAvfpVTsa589RrBR1xsi1PgrdlaEc91f3EgJi5jaDD4/RAsqwMh
Fb3aJLOhOD2ZLmKr6M8JSXlfzOKsleLa6o6V4LqYjjfz1Bx6mwHCC6gBqJg6DFOPdSMvCIvYa090
5yEbvMjxQtI+04rk5cHVVANAucAVeCNMQJdkjePxr2ZTI18zfAzHZMzxC4SaY9uFwlhcx6LKmGVq
dJGYY9LCSw35G2EU5KoVduRi9fi7J+smVzFs6FFCYDXnV3ur9uVZbDkZ1bOAXxDvL84WTvpFVuYN
WHPb484nkppyoCRBW+RZGv146WAZT686FU7+Zu9Uj1cnkrG42q0WuN6XFs8hQCtpf0djXUFrA4fy
S8ib+je0VARz3G2sJhYKwY50H91s64FJy/X9eYaAHNBLxxZ9g9OYbcih+7FOXqMcustKvZT212C/
s0hUTyxcYkKYYlTm2rZB1y/kx57D1/BReKzWBzWhtnI4hsIrkZr30BcAS/4tBDI8B+2M/A780KXD
jDrbx8OLzDlPs01z9RgTnsG7JFz3WHoEmPLcYunumq04gKBV8vCH7Gy4C2GmfCtFjI39TFTGElE0
NaJPq4jLlEFUTFEIk4QGVX8UvBwQQ6yPz/z0DTuruJrQEQaFVkbzcYHMHZVC/i1ozrk0lO8hVUhn
FN4cD+cBQ8vqkUYv4enMsWBkxweOlyMbgUzVYYrKKf8SJI0AvI9sORUuzQxcjp/jt3smroCGN/a3
dK+mgCVxi3YiRKSFI2DU6wujXIx9+ikyxcThB09y31k2CQkJkb65Uc0bCzvVOm9VgtvximDum6vh
HdK/lTT0jV2GsKV/l665zcpRZCNtnniolEYPoMHjjxf0ehiYkTPkWWGgcSY1Rf2DuPOGs2m+SODX
OKNZi7RDX3NhPGqNJYcpneBevf6/c2Z/FDzJT6ALI3WGlbYGXalkTafsm2jqMMpnE/BDLIKerXrB
kcLi3FaYLrgY9HcOYLxs+sMU+u0AnZTIcLTHOedWwEPSy9YEjvEbycq/o8tRiEgEIDUqnhB/XF75
yOjKaozlugROXiLgzHsw1ESxcbIHKSjhGrDuv5mw+AoVPhb+AfiuOCzNbKg4oszQjFUyAtf4dONN
e3a1NW3c17TxbFsOT3W/SKa/gL5jXJQB1sfpAsaEcyt3DLAF6o1SDfvtQXMd6y35d7OKTzLKB06K
MLFwoenYQ47mka3qjNvTJSrm9PgXwFMBLGnJZzr2bbEGktZZNEVZBJNM+rCwCzTH+mXdMocGkFTV
Bn5wEUVYNnymWHRMyB8qD/nEO2FrK1VArg/pu/PqaZ0X/QdCGse967PkZvP0h0Er1gstwO8ZA9WW
mjKeR6uFvyBreepWP1ObDD6QNo1BOVcPiuTerjZUM8hnSEB+F0SRzx/ImHq9kRRHWAujMgoiWtOZ
/q892kPLl0QvqSxAENF+tAb5RaOYC+2TvRmOsxIL4KFCVvDQ1l+LYPRps0cRo2R8qSZ1cDwk5azs
TB0quCf+bxrcljto9oYNWbcZNNWTxPaXrQGcLr4QybodgoSog0HvYodDmWkiN1YG+AyjHNXBNuon
TWLi8E4aoe250f3xs9cb0iQqMNgwlFJ2QN4Ddc+nxZ2Xf8+v0q1VRYDvR1XdLQxRTYVgk601EHMw
EJU4cRGSBO1MKe0uDaL4AdTMA+otqFsTJo02e11U5KaBhMiuLGfr/mUH1bJLywPC/DS6F28PWsze
wYa81Ds5l0Ce7/D5f/mhAcxmkQNk07cMn38vzO2w60iYtXziUxdMGsR7Z3r3HHXZUCoK4nNcoP0/
3iACWSr0OKyDnm05t5PKgNLgKvH1sD961Drrwm9Zi2ArRP8b0+MmrnABZxthIered3xrZRa5nuHB
T8m3I55c8UCXWv5pne/08ONPqUH6H22flZh4nBWfpWLfzz+12gP64pKrFPsDHN2/KvgO2Iwza39C
j7aTzPxC/uxP6JJagXLwX///pvvJ2J0eT4EwVR+tQIL0JdL9E7XO8/kwG3c25cmHWwuAG48RewIJ
gkFiVRVan/FKqqTAx/sNorHQ7C9g1tu6Ui/ifJgeqjQPDZihNmVxKcFI3AU9GAxdeZKAtl9ZfYw7
+fQevIDzcUb9XoX6I83l864+L5qm4I4gw3vY+ZyGp0EqScLEMB1XuAWNhYBtVitedWzi2D03tNl4
y1lkuV2mrU2Z3mUZENQrzVa0CYJ1hXXhy/ZX79PH6p+mZshooxgLMIJB864Y0k9zF3EDbXJQnJFz
nEo3BTTXgtyOjZOd6peYpI0Z3f8yaEC8HFjOLHabFrRrnv3o/ho17F4Zi+TDK3ZMOiCQnTNtr/Lo
FNtPdan7cNX8GDZTbZsQ1NgR3Y1w8vrkUaWM1UlRjXPH57bwju70s6edPvr8zwnI8d99ZmxbdIrg
bS3lDvFXgTj7Idhk7Uu4Ig9UShcQHmYxv7VpPGEFb+G/DIIWMXhkoGkWqsRRTKUShwPaZP0yzAyP
4Z8HENomq5aFneI5TLrZOoAokiFKHxuY7fcp7YGtTQ5V0iLJ7zCExtoyh9kRfB77mZbNNHO9pBnT
b8HIrLHR9ja2OI43lroLNpizYwVhMhUpfwcVwN/YqKBLaozrNg/2XRm3zkF6MWklZ5mhLMgobHlS
1etohIwIRmhwmuASdGnlrRMKukMn3UHw7tm8uLXCYhMyKH6pvvsrFzIzozoyo7vb7Zc479LiIhKR
sDh+8btXyi4sGNztmN2Zgdp0xusFmRpavHyKPh4DGWTe0+MDGdK5qJopOyM157y1EOmEc1agoncG
8N19zM9Y95osq+H8Wclv66KhouyWLOh0RMvduteWIjcZIQEiWtL8O0vfXovp2LBu+0q3AIKxgwru
2yxRBd1+W+eOkq7FFPfVhtrk9sdk45OwpvdzJBlGg33p70C382Hwi+h3tBk8UJJ8rnMdXASTzLNo
3XMs9UApGO6dllYP9jbD+ZGfr0Qgoeqa0GCh7nRqGdswhw5nLBQV+bwZRPS7rTpwrVHpIw8F72Jg
Pl4BT3dkRGPzzFD8wKEL/KKQ6TGufI3TEKRX0kSAhhI6pPQ6EIdvl/ZW9qTx3buSnoeWoxLPumNN
Yt8lDDPRBqAHRtp+rTZCX+XrXp5fKKxezAPfAPTX29wf2qaCdTlQZYArR3c1uYsM4qW39qjIiBAm
tegfrFdiV7qY07mtnywUD7bVfkKoTe/Z7jbQer6bJEUYBGXa5x8b7JcvfjLoMT69YInY/AafeKx7
pIUo/NY42NFnTgmvb4EbOlo/5AU2kTrMJ56fH32+qdmN1hDSIrDPfCpxP6FPiJExQksB71GvWCMR
gGpJaxAX4ixCnOp1KosAI9TrAbXfi4JGtex8Bxbs6xNtyYrq4ugUu7u6cm16jjdXCHw+5hWzhVPP
c6Zz2ZYX7/tUcq3Falcq6qhaveTpBMulkBbkEQkuNZmIH6qKPJyYZjxAEo9Tr2veRWoEI8VLwEFW
4T1tENMkPeB9cUMH8TTfw2Lwqz82UoZi9NoBu1Z3ktnZbZLJ7iVbw4U4nJPOj92QFJZxeXem/Ghp
scCCM1WOiPUOsdk+sIcPVllwwTPaDCrplDlerrqkV0zvlgM0WZ++Enwwft4CcOus0NWAwM1ltg3p
8ZydyHp0XMXkzgqwiIlmqFlXZ7SJ6b8F7FMR4ks16sUoJmObMniQBQ4YjfezI63qd7xb8fFWO24t
QaKonBwecJPfeZurpg783e0SWeQXRWvbissuqVUx3kOy+fEiHVmdyE9jV9E+uNCB2ZF+Wp1cjUc8
CBcjdN3KMQ9P7tJLu8utqlBzQ9/5elVnW+AFghAN2eBSDmEq9JWlSI3HsSIEdX6h8rNlLbZipLdH
N5vydmpbJCBvJOfMIimNelG1eyKeM8AcJUvEqKTa9LdtH0XUaMZI7WbNmDwuE0uouEHowcWiajMd
/wlKnQgsHc5vgmHXRbBsK6y1nTTvt52VR5ps7tqLPlRSenSF21nSIumHwirXMm5PDd7CrYcqMpWS
+GIK/N6tEnEFSfBeWUXgPUq+iOdmexFyuwvIrNlKmIQZ1Txr4tJ+x8kpy7o1CDpM8kmzeuEmCsBp
XoVU41IVNW0WgRg7dvmbkE1SMajus2l0gm1QMKRt1AJzvmXwQb9mw/43xCkZ8wR7WaT2xb+UmUab
KPerqKRg3nFekmhiHms3XA2/0/aWK5vdZp1dx9yuLiuFvx9fO5F0Qp33xOhRc26QQgTZ10AGUgMY
WwVoIDXLsjOMu1fkzXZXrEAerbhIhhMcIHcylqcCpyMuennkFQWA1bknmLVM4OXak2Dj9+j/oSdE
Xa7T33WYg4JxSqKy0OiJcNCaxQAGzc9o7LC00FJ10IloeG1N3iEJTn6ozlWYfoAUEgm4jd0h3tGk
N/h815WOTyG21CcUZNiGv4mYzPsQI6baCuAnYaSf2tWL6mk1ZQ2chnhkhy2bZk1JxaRJ1qgUtaHv
oOrASiUC3Ygeg5cX6WYVxX1MVCj/1BNKIW7FYVOHjR4osFJW68FdVD4ZqeGpow19uiLYH21zBhOn
WEDwMg3HdXNHer2Ns/GD8D78qU0+ChbvrONawi8ZNKX+pXK+LIO4yZZ74+snRNMh+IMDzIW39d1C
AdEPO/DwhbZDSx0rwYtHNfB/x3IsN5AHuEnHKN6bIjJd3k2GkKx3E4UKU7H3GFkCVwv+l0O00pP0
fwHO/BMp3T3jBImtFNPvMZTsEc6GciKSMsNXYhpxRl3pLSeW3Ss9dumZUG7i+zLJ3sLHne7VSLJN
9UI1fzd0e9nQvXTisihPgwYInntywTV+BlqadshvIr4ud5V7LQ4jMmgl6te9ZiAekQjWgamUgrt8
9iy6IMcUvTzW7J+uZxy5nDcKv02d1RienR6PR2ZEU21cHJpGh0UB3y3A3VWETGvo6N8QhiQsz8v3
GOsvZmjXEYSWKaPTy7t+NkZRwqbdJNQi1loUr9lwsDENNYmle0x6ribO03gijVi+E9HuKGAdA3M7
q/lGu9y0XD+OOJFY8M0wprot4+J93Mdb9lkCWJFw1+3lyJRm8dDChpVLxhp71092VNAw0bjBfnBw
0QCNGfayODgY6rvzZR/DusEfHABsujSu575MxcNFWP+u/EtwHizvQPmv4nzcB0yrvOxrgOktCpDE
tt42JsK6P7L/IZABMLvCywqrU3Yv0uqKfCIHfVZpacBD4cP716Ly5Xz6Cp5ja6n8fTfqiHZvlj/K
CGa3yO3/q3i62LQz2AndIyNr+z2So9wlpPjYHob/dnJ7iIw9QuDQVShP8v6PlABDOJJ1rXmFxnrQ
wCT+sC9DAf8x6BTn21Ccf5pOt0nKUaP2q8Oifw4RyyZ9v084izIfceYxaKysPtm5WBc3BS3Xpm3s
DIcVXp4asnMztRncKcu4p5aQM5ndw0ZqnvqG31EOCBIXuPMr/P7x+IqodhqscDIPORAZ2fpukq5U
HStGhF1XSDK9zm64T4Y4QlwaastcTTf0uVX+IEexFrCBfZFryKtZBxNRWi0GIKhD+XZUCp7BAsnP
vl2qypTH0dVOz8CxEEE/sOzPrzoOBBVvt0h8MIqxADXVC2wZxqDm+aSQhzxHjh89THyWhnxoiOBW
/eiLdtwc/W24HYboWbRD+N8jNCq8xygNZ6ZGCD8RVxJwEW82hOMLHpFyRiqFkcuV4KI/Mcy0ZJQR
5ascDKjKkPeeeWsOLhljBwmsKd428NuPf28nAl6YjpSWXpD7Yd26MPCAlKzC+hW1f1mNJRpv0JXV
3QjJ0EWPCBW0Gcx0FhW1+KW6OU2bIe+1yu+CXaOhT0EgXHc2/L7Smu7+ZKwL37ksd2AivqE/R1mM
mUsbWJPgg0Gf3v2hp47xMLHaASIbpCJkNz5r4NrqF+fPQvcSdt+iuXFkfUd1QNeTRuQ9e4eBRGmj
V8dV0aKcYynqMaYqiDl6fvQ15xgrMFc3VxSlL4S/PXPtYLmkI4V7Xb5myNg0w6saNDD4Og6YBrDj
DnU5775bnLc+X432As2AserGrPtuV9l6udOY40QN3W2e2rYngtChfdXK++P9Ql+CTyQEHCcPpvo8
gtsVwKNUoIWe3q8igzrmKsmZtFWFELfaKr1upiDqnFOTvOI7Gw9Sc1+m4MXOue2P/qz2rjWhgduT
LRjZK0dv2/ZKfuPqsY6QdXTJQfayZ9id0CWWfyhvacd22tiMRLtGNx9V99QUSnDS2E7CnhgVfzq3
gskLGLAi7yOlqNFiq02FH+6ZwqM0c8oX+NrglcidrZ1a+7fOzmyGl3cgjjy29uaFWxH60PpXqZLz
j7WCA1M48Fq6PGaBmKELsO+p4wa70KfZ0tMlH1TydKrdCEqX3f8DxGGIgCSureKcWJ6BRJ55afJc
YbeF82OOHR0kx5VI5DoQ7vzjjP8n2yaoFrD5Dj6QqLrsR/73+A/UHHazyQH+CNTgUa+1X9NjgKhy
tyE7pSnVA1pR78fD9pnmaYqCjyCcBB3F5NuMKCkR67yCf9dq2AYK7hF0Sbbf4ksXjlf7oDa6ZOZv
uyj3hrRbQ5jZbPF/JzksRXGP0wlUGWIdOoo/Kb+xGMbrM9TatT9pgFJHoS09C1T+f4qqPbgftjDK
025b+CRrAocQmLAZ1ftljJ3/a3mRgx0j+P+h6h7Nb/8SEnwqSmBb6+an5h+lkoSgojrPuYFb2gG+
4oi+ki14bF2MeHYOW0KxgD9gMU1GAjhaX9vZJR2yQzjcBpW8G7ADNEcXRKpjkYrGggdKWznYFNx+
PHvQc38QQM7ygYYqMuvTzdf9Rxb9ke76DzyynjOTOHdRz2R/iyjT/C4/4Ovlnu1xVmaa+6J5O9D1
0dfmFSYB+z3vbEnM/uJ/VpOdzfIibfrfb+pUZ+O77SWiBDBukswaqxZkIZYIK9/KUEWhlniaJp0J
MVHJiyTj1I312A/GZgcrMAE5c0V3V7Vuqx9mx94fp1UXwtD2Lk2sZhPHljQYo4oIW5in1+t9MigV
U7xPVdmdCXs+2voouoqQCbkqRoXNSMU9fA3bMgmLkBjfP0kjp+P6oWJecJC4Dda92jT5UZSC8+9Y
A9xztkHcMDjXI+ciisRLUpXgt566Vd0Tds833Iz+tTW6EpwEQ2dopWyKvKebZuqnTCY7S9zUZGQe
KbIWXM4QROINv4N0ODfp1E/1vMSgYOfKdSB4ik+LbIHCjXvzgEoDIFx5jCKZ772sMzh4SVJBmGc8
8n0WNRl45rx77/Rs9ypR3zEz3Y2nAjFhmh9IuZiwI58K5gruUby0zKzBR6EaDCss2R/FtRJSWyYz
8XBaN4ZBrqymNR6gRt948fNJ8oFhjUkaxyrmENEggNxe/aHFhX6/BKkbVhiN8J5XL+ik17Nk6Flc
Yroz2o1aPgw37nHy5HbbGedIkdRxz4VA+pnavujaNq/NIehGQxfCZxPJTUoEBBUUIUKNSyhQ5bxc
YjMg/Y31ROLBdqujxHHcIh5BfJsY0yMTzNTBG6TwL+S+WhU1Tda0vmIAm1yuF6ja7L/Zm2l50HF6
PmwbMMFnhocyEsBOl1WL9Nzcm/dXpe4iV3XfwW30WK9GZuWjOYFb6+TL3GZcWuPYSTxOsfjoifT2
CzNvQNzL3ilHT+P/4+zIri44+qaxd59bqE00h6pS35tvgvzUJ3PthrauR4i4kt684czRTfwVwyId
WI4Gtqo2eGcsa2aIf4/3ATKfSCMjp68K78ujNQmZiksFL/R2uaYFvWSJrq+Cqi0T12l5bZfOG5Fn
RrHwPH3Saa2Lw3dAUh2iFIif8okjMDSdPWcdggXU7n5xJsapVV2doF95vNi4nMKNS+BoF3+E/8mv
1QYuir0+y0paq7EyFxqI525Cnx5kURQaRKJphXVdOuG31nTZrhpPGrM36BK6hyoup2nMeBSJQ0bj
lkaKtJYQFVwmlXWwGCpto4vCvNEvBy3a/eaVhPrmqgNVwCm0bg62JzB3DaWJ5DFwTOAxtqQ3mFbI
Y/JmW9hCC4h9iX41te8fdL1AMn/NdMJ4Mf3H+CYxsfmsN9MwrA1+ILa7KdUzSsaMiYSHPnQLy1Vc
ae2B1KTn7QvIwmYHphQaRHeMdlldjy+ry/+2yMFZ+YhRbM1PcXVCz7PClPd3p6oPVWc2Bp+YSb4D
3w+jbkUrfBpE8oHFebQ4fDcRT+bm3JUu32cZm8nVavN4ZyZK9leY6MftShEG2hvwrh4RhzaaOaVR
DMAxLI+qG+5VHWxR0Vv3Jrin0QoNLPs7/4JA0yePzGYigg1CGtQdL65Co5+1yj6Yc+whv6XyUQap
AtSfvfRz9koN6eu9GRmtq0NIE4Xom/1nBl6eHusEAZzsByMmH2jI+a2Y21970e+k9tSXoIEkNNrx
V289dkPAHzTd8p48+kXnJXUS6FKDd8O5WwNknS9AYc9Sgoi+OwmDt7RJ1vQefIUjfXNCSKBQXPze
qYG+xCGgzqqxgHH0dOx8Vey+Z9TUw3hmrH5ncOg8lBeL2zLjNuf3pU16wZwqvM3Hr1n4NZxcS469
fGJEpvJ2YBYyMOFd6dUTWZNAWNY31fQqeNlzQYEt44cB1ZYGpUfcDqifeCVMnF/aheBt5v8NUWAT
vzTj3WjOZrD1YpIfxZWtpI+OW1t3Hz1KeWIA8YBZ2HKkYWOsFo3xuosLIEKTYlpq5bSKu1rZR8hK
fNdZpOLs/f8QhEKnU51mJR7CngAlUsnfWZSlPgJxfdgu9pAnRWZUWX5d89WCcIybudL7SpGOpJUx
XiqkxPoNVYG3IXE0MyPVUZEZ86oErP5yFCEJ3yfgzY08OEHYHMbn/iqUsmpGBX+3QZnV5GtUYstO
fIFnLF+R/px3Az9xUPCVeVCWo5ZRIjtXghGNTpW/Rj0WhsKDAHNJkSTsfJvxUNgdbKPMlgB4uaC7
SGSyx2VTRuKqorILgIzT54FPBuxn4o2itkMLf8HBsKrZbKnQVGoXuCWFfM2nvZZE+MRAnvAJOIgD
WtDPZ/hnNztQ0BCK4/FqWrOdfZkrK6YhmzO14KsVwdALi63z0tfMlw5lYU6odrGBN4u8+ur15IB9
T0Zi9bs9jL10BZ9yngQLZR27OCvCRLrbJqMRrv76WMpmn90iD2J/O76V/jAiaKuHQjLyKB4Gl+jU
kjqzuS5eqmi4MwabDfCKLOqSGvu6foNBpXpzgY8ADPdChRzvXJWQrOA1YdTGSSQj2EFH1wQicTyy
dmbebX5WsBtdlGTa1t/xlATGZDawsVmyQCNjyt+PkB9GBXd7iVFnvIznt3ObgpsQ7NUSxSlWBtgi
vk/nIt43z7lGQTMy51Ou3oVJ239nErnCFCGyZMsJlm9m4WqoRZ6eW/aDWseP6lf7x24NocHbbSD4
Z9HdGAo3K4/AbEdLXtNjmm2InAfoTQjoqPmb47zh+E/Pl4rpReCoSTFtX92Hi2TrkqWQnAlCR+/p
+gMd82JAm6EQWJATiQPs+E/KR3WRpjk1DjMPsO9BwhFlerjp9AgD0Wrr4wbCN2M+NH/CFkcA1QeY
VaXjQJPIcIDV+hRZ9FbVvv+7r+EnoNQ18fY0x9jEIR/X4wT6KW3I7s5+enr0x8oeCPWmKc86kXZc
3L7mab5gWfF750cFOMrFsFM2EIGIDl/B8oPzmOzJGHasKYvbjSif2V+dirBxBNcwISpM1MVh4k0J
b62QnXdIz0GZ/e3hBxEvBuiPRt0zG7EiXq1jHNcVOQMK/j1qKijOyfOAYAALoOFcbJVMGMalAv9a
QQWyneq0oGUpDJjnQRLPi5M2i7IhDfmeWeuOIcrO6BbxnwU9VmCHbAGy26du4T+xFsr/HIivXf5x
R9E+boOrKLx4GVgu+uAhcSmzQI17dH52BgSnXAKOMSmBaG1+kaBlT4ZUGM29RClYOTnEawwPBd28
dsn320X64NwgSzJ7usDMWQ4dCzDXmuTNBumI2zQoUMGtERX+o3htKSOUaBs+V/x/tAdrLJh61m01
uc5xybSDuZSxTbd/XjgmLol2l1gDuoVH0/icFYy6gC6jLQZjlooqoPHLKfa2pYYOo6C68QgEJVg1
TspMUV6t8q71BRLvtSbgL6v1QkJl7Rg7xMPQGNqBOm/s1wq2SeMl3aHhS1ILqBykyCxCFfdcuqpU
fLzp+AX346GyLsUoESjrzK+35KbN8/6iHVD2K1WzytIpFDiv4Cy9WBa15MxsDRY2JqDVCnJJHNuH
1dWCB8L5RgsF+W8av6NnmQAiaXPNabJy16+rrUHQTpF3eWN5pSlx9kt7LPZT9jNNnkagqIZcu6AQ
I1nxoe71pJ2Es5u3ZbL6dhy7rVDMENMxFDBbxp04xvsK/LhE6LoCP2yUqSIu74ESkMuB+1NSl+yi
Www7QeIjuO+ieXUlevha0Gn3sv0kTkqYXWds/dSowR0CMInRTdOlEBg6Lee2d3FjJTPBpHdgA7De
0ESU9RrqUGmOJp9SgM8DkpklbTw1aXWM6FUquPBiMdxd0TaW7U7FzBpE0dMyjH+6ImwC0LjNRazq
IkAPJQQgxW2h7/ph1n2ErxeMU0Kdkp1GM7LfnnUW14HSwauCMwYBG4IPWmHXSjjKwDYBv+4NROPO
Uqn2VUq7NJ/TA6IivDMXoNQKPyHAnsnBq7Oh2DINMFexB4rMpz53G7e+C6RjvG/INZNu14Wya9G5
q8B7wDD0szDTdM2onjpYt19NdfuKxJvw+8s/GrCP/baLekl6EVOnSrUzeTP7RD2sAeacdFmbgSAi
/l2ncG9PQYDfJ+mpjYNBW0MjxEAlQNxUILFyceDy+BNiPxZ/j3ZHvdu3BmvCtG4HtEDF6hNIpZqw
SR3H/+FdDYfZH4FqNsOfvRNGcnA6DBop71pr5ewHXKPx4VYHA5aZpxzCzyvt3I7Hx6BHwWvbqCgq
ljZTGFyZ5jV3DEdf2Xzou7BAaISywmjIXBvjdkoS7DlsmlRCbod2dG3DPNFa3wZ3J7ieq060xU/v
mxJOyHXMjGJkb9TyzMufdxwA3XPEDDX+nbU2qPYOan9qj7RxN1mnzHbk8s+iT5h2LO1iJFB4HegD
wskuEmbEyh4x4a07Mde0IEV/U4wccw2jzHzq9H/iUGkM0aGg8ExkFF7m6B/QAmBRM7gdjrxZCcuK
pZnEKRQsQnGvVRZOZtG8LpUeGtPCInRQlQfMRGbtPgP7eQOdF9NUtQN1/rCJ9NLGQ+hqRc5yGvxv
wreYzE3n5u9taaQVqmWyzkpAWf0jpCMqwYWrSdy3xTE8vd/caJnxLK5+dx63DAllIgexr6bXm6fY
jBGX1V4G1FWEwwWzVHaXEE3Tjxh83I6Mshs+O0Pq7e2p9YXLjOlTU8VofW1EtrXmhzsIznS+3ZUT
3/9jKMUffRALLLsnfjPIH5DRcPtP7fAWwrF82ohKyF2ZQHzWsOShUiEf39eYAbzJz8l6C3d2jXpd
pECGEAhaxD2LwTXgWwibaAdHN34p1KtJd+TLToI86Zj+kEUNDJrarlLDLIhyyotrdGPVBrduj8Ce
QZs83usBj3EizDRpsjTG+UI00MgLYsowXWn0E66PGGjFAJeH0Hne02dly8kc9O5Iyyob33qzuLog
dPCZKx/NxMJ1lubNT6NlE72btRXiWACIuhS2MgMkVOs5kW3kPC+Dzn84TdP5M8th1WAhNxhXxYs/
I8hdrsiFakV5b/4kBnLNjfbji0ffAd+F7hIMS6Wq2pgapDlTJuqQlNBZ9r1xjyZbU319XDpwTvke
/9AjpCfnykN26EV/ohPPRxshMmL8GdoLnnP0pVhZqkPPEco9p9oHu9qeqCNDr2ZfUHP3h3rb4aHy
7xcZPvXk2IGjFo5+1tqGJle8zhleAj+NoPgOhPk8QwT7r6TjZc8UfkvD/EfS+bbKzDN/kMVFckFJ
jSOJvJcc1Vw3kfJNx2v8Tbae2TU0KMhlyrtmtpoCo+105iFkCQruHecSa8dSPNstekxiEYZ7dMoo
44JLP+2svNLj9Xt6qZ/eQAWaxGWPDORawkMJiHjLN9pPANIUF4l6TjXGB10p2FoWdu9we/UmTOY8
mET1KL5vaRi1hafSWiExzyy6WHn3sKSuAAVK89iQxIENW0T7mg+NWrm29y7HJrlcrrHqNef1t4tu
kyOaXq3E3HluacTPuSNIk1wzTv/KFCkRlHZIPI/1cDqlKTFsIuOKh4JGJ9n+N0FR+KQRqnG7FoPq
krC2+Bw/G6666Dnq6q9/lhlDKdeTbJ1Eu7cMT3ljaoUDLmMa5bdWBnURIr/NgIbmhva6gQFA69RD
OJ9+lKSVR7cr8Yqb1gpQ+25CTcRM1wj0eRb1blZbCCHhZ4XjMEW73cLFHdisP8qm4INW5MuZpf9k
FbRYHGIycaJbZQd7MXfuNbQMkqm4+W/UzHlBSs2YEi8y14EFu2x1JI2LGDcHu6KBA9bye2WlBTrK
+ygQJ1tvi+gp/FgrAyNv4v8hxWudkeqNWZFv/uVABz4hdp5hoR9MM5ST6CyyYBsyaAU5/GPZlzWd
JP0aJL2Yx3pUvjzL69EtOpiZWA7uQzg14seXT/px5Xdg2Dz5qVkfLXI50j9DB1ggnHBT7TUHPMyO
JFKXktvtaqCUpixWI81l8bu07aIF3WySdpfgHXXawgDQIC428Wc3MVp/KX4Gk5SCUp0qr1VNlhft
w7fiwF08FvLJLbqRVdEOm1Hum2FFNVUys9qTnzqAGD0pHYk4Dpy+9E6eQxOlp/w7ZIDwH/lx/0i2
TwfmclujdcH8Id7aI0nupKGtZktaQ9Tu00O7snxfZoBTRtbC7VyFsL9WL9I7c8L/587XtonHAK6t
p9b2Tjdoi4cA1wdReShx1qwcNGXPwidC/MPXTyiL92ojSVzeVpKppr01XN43N+OxWZmBHjmUWbmT
G9QHpI1gzmz7gUk1mEQwa9Cw7BNqlLlc7CQG2PvWJ/zDw9hB6Wladw6owXh3Y8VCqAycZy8wV/kW
teWMTbFH35IHqbi93+cgUrPnO4p3ZIlpv2AerYUSVCiA88pPDXQzc0H08VFn1lyPeEjiwcU1dfzk
XnM3sdfgYXOQyuOw6z9bypBLDT259AkF4aMBbLL31x8khoIo7WXRfuZFmA6510BRGXhjQDrtVwnl
54PA3BqBh2K2tnU74bvD8b2a3sa8ljG6+L6bWyTh4lHV2VFKudhErJ+ivS0JQRD8YCrjCZCMO9Ki
Yd01Lkn6OVUJrXc2bmKbieVIMNHvblN8uwibljXaPPNba9KSqrMKoFesEvaSjL9PfVhpc43nvcvI
AM30RYPVtYI50/DOVeUsdeV0DyJmhwKdsUIeQ3B9b6IzFKste6tODbyZPkhBRr38Mpy+ryqMhfcq
eHb13K4TWjD9CoDokOoRJUJ4iC9IoMwoG3nuZry7rdPeNcYzLHVD//ezYXxzgbjRXqnpfHJtfy7U
puQ2+F+DuDE7ktxykD+s+zZjHcTVWzY2mh4QdqbeDfGKpRbeFoO0lHjXm3lDpERYs26+3oQ4oaeL
kiH5aqYDJdPNVAP3QK9oiNxOn/YzHEbBqFkri+5XAyGJBZng3FDUWOVU9TQt31mwHIyodCmRdj/e
MB46+1iER4veVgdXxR0YSCvAWrzhBOUfBagyFB9KBcotD44V6YdMKg+BdNU3NhmfNCmDX7dWKG2+
ZMyqjsUEdNAJQKk9JM0Ta+LesQsKIhxzQ0eqvmRKxlMz3PqEh7IISv1T0fZv98u7qXYYJp6aJRrL
jixTkE9GmIqCspcth6CXaGnpBI/5QcXDK/NWC2ZKTrVleHq1KRtLUt7pBHs1iqOv1Tsf6mENB7lr
Y5Dg9L8IBa//JGC7z8wjPG9W3IhCXOdaHjf11JU9O0K0JDMwmakCEgsMgWExEdMTcrV3buisyuqa
MjwI0WsPagAJnUc3T8hBsJmhf2nzuUqyyVjbN55G7PBci2vduA7zu6iuURMLjBL5OZLcD9KiqzmC
ai85D1nPIEV5GCPS1PzNlvvF97kMZYJJCPav0Bk1ZMoT8g6hsT+H+h9/HJR4u8Q/gvXyw63rAlZW
e5FuWddHcdWiBqixD+XdOTtF2U30hvKu14JdDHHY93YmnNemiLM2RuvBoEiMoN6opk3jVk2OANYy
l/E6gmduoZwWCwF9nKFjsWTiEjn0OxKw9FYSruLHgexWXyMFKtXMB87cnQ1XQQhYMZSQX00xski3
6PrUJXgcGN5PbxxTPLa0P9xv/F9av17KbfJHYp3tVKKTu6eQhITIeao/mgYbeGGOq7O7OnX1dNDK
Ax8hqO6hiH/uje6/bxtWV2FN9IyZV/929hoS9vi2DYD/aViWYIwlqHQQP8Y5usMoYkC7SixHH0la
012AucduYIQqj346R2Ma5RBLdDAlX70auSGXutsiAs+9I2peSqs75Iln9vUOUgMsEtdr++BzYS/7
enyW37BdA4yD+Ek1H5wMukEvS2sQeb0txa8pG/pR7bOqE6AkEpSVBAIg1dHrxURKFDar4Oelp+Z2
M95wgF0DHxg5ijQ/V7YsVDvNS9JGiWxlm8vd+0tkDnV1i/HDUYDWsyd5OgsveofOgGIbBGhpqiPj
v1SwbN54rGTyFwCamazNhdxYMIiN//9TxQSNd2f/o6+leUc8EaGTS04VDsavA8fYtZCHVDuKaIPa
y4vHqjF7uttl43Mgjkg2R9VuN+pgaFFDt7zUWGlmRarnspDrUD49/GOFjyh+F/OD3DyxkozmnweM
lNHURjj/h0q4x7eK5mtauc6pfrGRV83WPjgUjbtw/Od2OlGgyYEp+u3E2KW67Vv77Cv2V3qRWId2
astxAW5NKG1Nd3j4Vb3PDTDmwKg687yRnLR5+BHb4+4RQ1bTbwkcpbYtCmY5cJam9VKXoGxBFx2Z
YK6HK2s8yZwoF9vfmQUweJLRyf/EyS/4IuMTdv+nbgEs30W1j6kZ7KCJFjdou9nfQN0R6JMAomKx
ui7MvBslNtvtQ/svNP05ETfxOF45yC/ycs2mln+OUHMgg5o7CydOiuJAkABxt7cladqkKwcAVT+K
768cXXO+N/U/w/+oLJTo70MOEH0ZHF3qKksCDvtkdxsu3DvDODUXbhHsw/7whXJttrXXRYPUMuBT
UFE8y1DsVz/J7RwSO9Kfrt6AHDaD3oBOu86AzflUOvPEMrkNqN3ojr9KILrNQbiD/AFu1rM9pNxa
Zsf+wWlAzHIBeo7WKdbeef8CozZ2B+smCTDPGya4IP5ptgw/jWdv3qu6+uhzTiHzyJJJP4ENgbx4
0jKj4thkYtWo9kGtjAD/nN8JsFZGzmLDjEYC8yd/U5DenXcq9sohNQSHNAlXcHIqKFw7TUsdi9y9
pdd/TkEfoMK4wa8RdmGyxsOscQ7XrrUXpwa049C/qNXDlqHIlUp6zkZNRNc84IYjNaxcJmjZ3IAk
UKVttsc1S/heotf+2ehW+jn/GqlOHABg/Yodi17ZHlrEAqvHdvoNXsPt9KMiZ1HjuSkr6jZ6P4SC
2mpT+xqtDzmz4iXsibajqLUnSdwMLzkUzLPvgGFTbQaGNQ9hwLoXus0ocWXkDkRkSCfAc4p3aGW4
xjAqr0/YYagfqEQm3IhUdFHAz/wIDZIHN/XEkjkUSLROG5ftY2OzTded+Xn4E1i8T5veZB7DLxiV
22mkRvdID+/vI9NPoENFs/R1a3iCc1a1myApHX/9AZ/+emygjgY9OB9c5goXYzMdHdOO6bDG40k/
WzeTLm9brqaeMfmC925Eh33jjjmHDYBlibgpacJMwcN7cF7sE4IyxV4GtZLOzCANh4w4LWmGsh+8
aUeSFY9mp1UQQ8cQOfGLmnZA4U6SAUo3QtW6oGcMXlWW7hzbZsRlrpDVbA9C/InIJPQ+S9KgXbfC
N8l4EIR4VXFxHMEj6PTEn9pRyt+xJsAT7nT5twsEX8n5DpKvfuDP1i1HRBc7NWvlQgln7bb/9/hD
UN3gGYF1bXDmtDfpbs7VwerRNq6g2FrbUQoFzJHVT+fzHd//mhiI2YXR5mEjQ70EAH95H4vTkydv
g12u5QapBD0NCJVaV3YCuzr/36sbg6zqUOWaV9erbBMjsuZHzeORoT9jgzpJDMGNj9RM+79WQIFS
inNXjt73b+P8USwykwS2otVrCVaV8A6l7YhpkaiV4w17FW2iTvqralfgWiIAo1RT09CSpSDnAWg+
XVee84PgAXuGArTeVgZ6vNMikZsAQM7v5Ac54zB8K53SBiOUdmd3vTLyLfSGVaMRC8AU22l79FIq
O9ePz6+rCnPWbUxedEMuySXEk1tELf+eyEeAtJlqPX3W3R4Y/2VcdjhowcefGnUQ09MlL3KzcxYQ
CXX6qppDpOe1Myxc5G5fiEtEUKYXcvgFUrvTnjwZ0qCEqNlKUAP19Td7DMUEp+aIY+DZsGk5+Wiw
1T2gc/oOOOIvOAf31GhUA0l0ZITVPnnZXIV9hHo5aYWcFfc28HlS/s0GpTVbNLi+KO9t1gDo7aTE
1+g41o4hzdP/30SFr3BxfY7tNZUE5HL4syDV/7NYPVMmGNblkLaETjjzlUONl4yc/BnbGe72ribb
6FhI9nODmZ+ZbezMv4Kec/u1Mij3YDKbsl96HRhMoh/wGEiE3u708479PHsBqq+YrUjq7pWF0357
YXWfVuht/+eiKcox6CYXsRVuSEqMavuQ53VBfivKIgplxBPW9Do+bLceRhBr2sPH6n+iljI+SPAX
0uaHTUYNg5ETrtioOdlZ+5MB5JfrAr3+N0w7yfLqK1kFK8sGlrKfGUyETpPWTUxCjOLRBLBKgsTo
+EEAsqYnqNDxeJiZgiaKdcOF4yRKjYZMq5tdS/9V60m1ghDtwO0zx+TVzSgaoK4crcmAUapzAdWZ
ebo3QtucvZW8t+DnTgmcWlk5MCBrytwyprO3mWu5jdURjxoSbp/EfH6/SPLiLKy+zdrNwLKzgsnm
nuL6aZHwZIYsEGwGtUYNEmHYsI3OYL89cKWMcMb5y1ePnKaWFkmDWT9ERpKCNAf9/a5yVFUbP4VD
FRbkTREHaIdOMfxNj7iL7tNCrxMIKlSLPIrvBeNTRefHgJiIShTiltrkmdJmmSAsNWxdU97RT79l
cCZ1WvbZKBmuNwH0iK46OLtUP95IYHrkuEFKHXF6lmUKin4j9lPRb2RAAFVugCIKh0zzNPVEg1+F
VVsTBVUrB+X8TP6cuk1n1U5dJ1+mhjPqQQULXPrIY+21ysgb4dcONE9TGN6kqzkkknj5Vwq/NRjn
Dd9hx08d4LsCDLIrYa6L7XiF4Nb0XWGnI6yEcrIyC57iZIAC9/w1heiGxp/GjfrxJg6YQym3tEdi
C/0IVITMij8jHi1hssPzt5+bELTdexZpdh7tJgZfuK8V4UF4WdzZ8m0oI1I+r2EYgcwuPKkBA0In
m070wrThgQ0k3MsZpGL+mKevxncVvGDW8iJE7cnjyWy3CB5mrvKeAklQzusbtzZiExE4tWm+PaN6
ps46AWQejE2+qKdVwq9PzZu/jXzj0lw8kmBVM1DG1zSx4CnAF0ywJigtAqVLy5DxauIgYm2g955u
eaoGFm9AW2VCXqZt6nw876KB/EHze94WGz7o4RPS7w+XbVBHjdcerkRqfJXGtpuFeRt4w2S5XjET
cHf3h+30ZfZpkuGAc+pRLmOF4vNAIq2ixsMW7Msn1OTVY6sB5VjRD5PMX4cqqtvLTqQwmH+LRH2W
HMN8d4j/ztkI8Ddks5MPYh2Dil/FSdtk+f9uWPbbk2/VFe+su+XXkCG4iigG9fypk7y87RPQwnLi
RP1dKwHDOYVOBWD/kbHdF5szzF+WmXx8LRLJcCYsweJv0TqUK/9bJgAamakP38lee53nHvu+quCp
N57KxAr+M4bQ2Khv4jrVbkZP4NzSaxXBgFtmwEzOkph0IVJlXxg28ZU2aCsYUSu5DmzcOWLuAdX9
Orao9F9iCod/Oc8B6uF9R34SI2f90ds2xTR6b2DWjpt2uWZb1Jdb99bwIibY51SpeBBBpnO9QE0r
1UqqrBqNlN6ZkxNBE+NbVX2o8UeMkZrLOJChhlKkUTcE+vhsWzA7Fz5WUUw1M51GHQNR9qxHim61
JbHtuvCYb6izfYkEj9gtuzwGpOi1T4AFvkrM+p/cNwQ9Mcui81AuQoJ9Yd/AjkQJYV/xlFTfJLDX
5PSEfkybqTSEty4CchCZ0pl7YwvGvzxtE6Z2LFJ5J94Ahp+BsedlikVGL38sFKmSe1M4GGIa1Mrg
2vQevzvdQirMcOKH3A1QO1uR1ZNBGlK7rOr5yYJlxL/+hEdJF8+FPrwAT5dWb10upsNPIeW05XAb
O9aeGZm4jGLES/NgU+QKwtwXmtCMR9Iw6DrnoMYv01aAzEFK4jOLWywulPV/Z14cl75Q4FC33YxN
dN1lDQx2yYJ40rPflyE0neYuyKevEaqKMIPBlk4CgcSD8Hv6OmrCrCS95fprtF2Uvk/51o6tBFsN
URdAakgONgGGpQnaCMcPr1oeGmiMcWuT3w7aCp3oyGkGsXNCvANbvUZY+lCFDs9usTuL6X5ei9L8
p+HQ8zSuy/BJTeUTb9m4XE9txGmsYjidFglBMPwNUtysntnqHXwZqkakDpomqJyqEzYNpUkYqQz6
lWHA4xvG1MEESsNka/FBQ5O8WhGiwnJxJtUrLx8QhhZharltqUa+LKfYmxmG7FPV+OjxYvt6jPwe
tl1Dvz3OoOATV3Dn3lelJ3GDe916og9l4X37VzZV+Joj5m8DWHpHryj+o+nJ4cBVmCxtLh/8OS5G
SqBngxKipBProduP8H1KN7nk6EcwtQ79Qj5xYW4Ukx3bL2FqhKSWCpTFWKrkRN7fpbLenwfC1K+O
yY9EDXOaEngEsHaVWLoZScRilzgn/8gqDtYQ5ihb+DG5sKgzGt2EMLK5JMlTfzmvGROID0oTL3Jl
NMzdJ+RPDGKv5o2JkiUGvMFugStTL+Zpm7fq8VeDv+kvqYNLPW7RUaqs6aFP+tp6ExkfVOLb2bfo
mRv0PkONcFDIl2ql4STrCH89sVN1Adb+nbI4sTXRWqb+DL2iZsF3+mnl8YWVy0HvnbOkHjRGhMBP
4w4so1t3ToMN4aPFz+quSRgMptBi6dIzp9CGzSd6wfAxv4k19Q5h1d274o4wg3plCNHb2tHFPIzF
vSrtazs6w67KnhEFajnP9V+AnReVu3ngKMvcZ/aaNYsOlN2/9menyiRa43wRH/LYWoTul42C36xx
ofkPumg+4TdsBJ7t6K9J3t8Rg7rxd5jsFZSwwDtv2AqH/kvapbnKIOsMwsFI1SyrK8mnjKD3dWdc
VQTefXPpp19zPwYAVVyj5aXUt3MfQZIN7qe6p1RM6IgdUJxJrDqP30Lflri2HwZZakItebe58deQ
/LMEoyA/6bDWEqbQYy1lFoftRD+eUS6KxIMiNCAWmvAj+qjO4Y022leir1EiBdEAjbEpuQpF9qnM
joK/pz0blm8JAf3txcMYc+rrXlo7b88z7HGfpphEVCYBxlpS50MgEXFEPH6xCRzwDlbfZrV1icOk
o8cAFJv945ddoKB7g/mLihe83o989YT3FMW0oYmtM5xwWv8hgCO5v3OuSQlSlxglrN7w1Wf9A9bD
mK0rENBwlRZiqvO8OPBVhIkjkScWRrnDiGHtPbMoIKU6iFycbEGdF/jX0GBexZlSz7wpVm1Gq7u9
vNG3eeI6Dfpc0XxeZKohppFXPyAMauK+t6DCseuVfxXCaTPzTmOLiNUDXXWRjCDCuEV1mnWG9/Vx
LpgXqvMVC4wLNEHuv13gwm6fdCHkqQvxWHgoicZ23wf4Yu8eyOZf4kYZSesbEZJreLbvp0Rq+5Cb
DDf6ubvAulK+3ztQj4rwFZGGOWo32AwjD+RClTddaKxeMHYheSP8gFK30tDftMe07fpDeQRdvRn6
bACUeUIwPDQSDV53TRu3cNB6xN79bSMM0hb6dYyY+ZBxRMfHcbbm+VsuV+d+yPMo7WATufgOJL+F
Jo7+SUDid5PWHx9pCtrgb4AzDXdJmgLL2dJ3pMy/rvrFl2EcqLgJ51Usv0l01ZUTpV5nNrXLGLMu
JUJI8ao7EYacWJoL+i45VyaQ5NQHWYQ7DeiZtLgRcpVMd+ReFpeCwCCiv33BsqKJqg49PYrQ+4K1
d1GW/FIMjTGGNx3bz7WIhxY0P7kDLzBTz/QCVv5CgvGZGJ53jBjE2W19v9tC/FE9zhStyDVBX8I5
u4smuqj+gIgguXW64FNa6Ucm4MHB3QqpxHjCtS6CwqTIzK7FHGtW2+AdF3S+1Uq7hn77Y/N8GK4U
p8uVAoU6+PMbX7NjnByjYy3sS3wvdbZeoXL5bAiBl15LqadD2x3w7U799PKeve8JK0zm0n19LNxa
yiuDY0f9bz8txq6ym1KNJHaO6j1s/61oSmSVy+4UDtshrm4jtZ6gNWq8IkGTuTdbIFbgiSOP+Dwi
1cQuLUyWLNYr97+fPrHwc0t/x5HT5lJQLUMD/RuOeC43P1eF6XfZFnoBp2crdhPte9XKSceYDM83
x4BrPt285aEjQBDDd9GPb5A9QeSsbBgXG8ff4Nvts/6YkwEviRyHQV0yZ3zgD+mF5+ka583wggKx
q+YuEe4lrJstsk2jbKoRYCG6752/eCmsAfx91n2UgRkKO/++1tMf5rVnscXgEGLcVC5ReN3lvAUE
rHhAlsOWftjqB3N+K1f/iddU+EIQN/pW9YGDaL/NYZYKrDNtDDYnwiHs9o1dNgy0kn9TjUTsr63X
zF4sOlF53cvuA1pUNJZEoRIIiwP40JT44w3l87GZN6EbvYfT5aKuofTACSAaMaP+BtYS5q+HS5WJ
WfN/nubIHQmTYtXF+o9Q6qIkDHh0xpeh6iSgboTYTiYO0SRh5wthHB4lweEFDw+Lrl/Uv5hVqW3D
5KzyuCOKnV/TyMslcH3psnMCGcBHtQwWVX4uPpKj0bFonTA4Rqk4sYm8J9DU/NwrBm1+Le2GMdWZ
pmYHNxiJfYGJt47P1wCZ3qNNGPEQXFPGNA+idHIJwjU7CPgkpN4BcT2ZAOV7iBUgTsx2dTQR6H7K
IG9xb+nNYFwadzuK3wCMjFe5PSyPwvCr4lPYLD/uYJ6oPw08KCJnhKMm1/ZhRA9FFe5/M+b2YAX8
IwdYVxQvk9m9ldw1M8w+nIZ/N4ZaXPfQE3sYcLwFtOpyPAX72Nwn5X+F3qZVfgG17/CYGRC4XYEf
LfJNxt7+KPQL0xyWs8oYNSjXovvWutKIZbHuvuso+vDvdeaZ5+JqRlBoe9UjfC1wF/1usPp0WpDn
5Pd5Jhp4EvPg6HDDbUAOODTbDnpbt3ucUPUk/VwYPWdxmU7QMEVHDI5MOVwIxlKAPTh9jrheOXmh
SfG53KefRhJu62G9ykYoR9qUIjcuSjxWWbDOpguofh1QT/iL3BK8GX22aLtOFs2U5NU98yB5Daz4
lDQO3MsvnKpZNQBA+L/e5TfE0hmLNRWq8hgCUqkcWR99Kr7PBlswl0uKJSBDGl/RS6hlrtCvTzUg
21EHujPMav8PRcw62700AOdA58Evm8/F6jARQ0uDUnNc6R65cnWxgAxOsIKMLLAxFOVYDd2NMqqp
w4CbS675AsD075/tTd05WwcPn/yukyf0+7xAyqGsEKcwM52UsQKcuarPburrH1ReVZRTFEQCBSCF
yUu9guT9+GdmFejdIrNVt53YQZO/bVxRB2fDoJaOWxvbeADzdLnJtBt4WK/P8s3EZ/u0SplSgW7G
B6yIucyzzYtGtFLj2LqCYDC3NcTnFKjFmuMcsjoksmRPxZyzaqG0fEPGC+TnOIaaVBjQUtznlRAD
N8Fg42YJ3SY7iw9CPdWsgE4pVweirK4V/qgyNnPyO04WkvqaTBcWhevwEgl854fLIMb7TKfZQ8lH
CL19c1DjY6DOtgwcv6fzMwJoIHRM4cYu+as19AiR3YS58JemCR4/VVnHxRIc15v0f3x3iCjNXw1U
z6gFIccYFzI1vaU9JPAsmDBQzCaQ5rGyvMb/M7E4EUVYg/DgxI+hqL8O3J90cx13Pdmj9fMiwdn9
FsXTHT8lwFch5KFl4TS+aWgJJvqvcFthyEtbtfHwEo1iCpMO0FSCOiO0FHcp5HVg1k8m7AiYsYqL
f1UdTjsD6wqgjeaFh1sFfbngdgmMh1xr8EQHRWH5yVS6zp6smjsR9z3pH0Eue5miArFQpqXIozgs
zWB8GriAS7f8cHZLbwMCD06F+2J57ObFUKSMy1cQNc+zDrU4K9ER1E5zxqyAP8GMMKOZGDSYLkEm
NNzAxcKRd4XFqAytWRlwu7vaHSVs+c0K0EDJIZ/7Wq5XL8NeanECEmOWtHzKeQQUcZzdCqxM8J/w
TrbY1jLia5RuPIkmmz9aacKjSaDMoqj0m5RUXFoPBPaDz2BPOKyX8tsqZ6BRuGy4XVfHcUQq1Mbz
WE2g6Mutw9vh+xlf4kJbnCE2xuYUPkFSTUELZutApmtu/OYb7x4muZ9kn31XfEU6QYv5raUqh/ZQ
kgVw5zuxWsJ0PCL4etRWxcAKNJ6Cu7MaSD3g1ZwqnMVAmC+1hQ7jozfFft/Zz05skRAqbK+CEHBc
qm2Tma9xb7w3PWGnLxhZaGwq3CNOojYNFmdkPuO7fn/S+ekOb5Xmz9nYEZ5qBcYj68OhlLVxz8wv
+ZY+PbpzpFGGO2tpkvsjYFmmWcB20oYbJszZM+DNI0bu+zR4aoj74uPpbF/Xk7ny8VTGW2Mc2j24
8lGSW1m9Rqls8EMDqFpplGl+25wzNyr4MvRrg/MK/pVJI34FzMRi7uVRzzwyHRt+y2Rerl24o8Vx
dlCv53JLg6iL2dFXrdRWVV4u9Ch00grqS3F4n6CizL9GjHfTX3aJgZuDmVEEfKC7YHqLbxm0QW/k
66khKS5cpbmP5DStylbQ9dX7dKwAkDXs1Nz6PybDL26KRlBKu0SkJtEFx5tjsD8XgkdUBWKBrGT9
6Hc8JLlvX1f4BP3eWCBz6AiDTtwdB13HtZbSqXpBWGh23IpzYp1OprSA/hpnnFwW0FhHENsrrTec
fJZepwCNK5sXxCPD1OnlpYFTWzXeguc5u9PcprY1GYOzcBi3jppE/D/JSDJ47kCXrjx4vS5C1vzr
vhUm20eAwmZyViJw+JwlJSa+sfQPsGVHGa+TeLMBe7xApXf0utoUy9FRYBmdlwz8r0ofnTojz2iN
zACuCXvxNcbWvz1b0Wx9Lepw4dSSvCyr91troUR7MrZGWcpPt1CdnDRJE7H69TiuV4GPKpwojVGV
Tci5ri5SH+YwZPrB5AZRgJaCCR/w2IJxOvwfH5fRty74V7imn4g92Uj6A7D0EB3z4k/0h+A+BP7R
zAJCTjOTSj4sUeFj4q81HtEwU3t6NaOAIDkUc2GcDb4LaXns+eObE0vT2mXKiT11spMNjZjYziUF
Hc41YQWVQ7saNfmV2U6JcHEPW/P95zxX27riPJ6z6x6dy54vbMk9Vgzhd0uyP1EEXg3s++vwTMeL
LfJHsHSjfuAqxD5NTsogGO9mIucJF/JDXuEpQsvmDP4/WorA520+Wi7nAzQZc8mob4tGX62zCFEQ
zqxW30WaBXCUtLRnuV17ZIsXFsgNdLdAILoRLY9d7tP3aqOvw7fL225RBFkc8DZrC36XLn+W60SR
2e4o3SEWkwo5KL4KIKhap9rOmDJPRqwupb8fyP3BgJIOsza6bLePsHB3km7KfcVU7LLpn4Zpy/yo
/vrIpWqCXZj9vqnRGmFWVBwmefFgc1plqKMAU+8hJUaRcKS3hhwYp0Pvj0f1dKHjsKwE1zWHd+3f
q22eTYMZVSLyd+cnunLVIoS6IBikLCeb2vH0nS4O4iXj9EtXuq2Dpr7/QY1r8SPrZBMAqlo+mqcW
dzCfcYDBMhr3Xolxv4JRJta/PXOp3x3mIzsBTKkZIJZvFdhz2HwAt2if0ETqWlX/Ucxh5RfT7LdY
b9qaaxLk+SfZetzN8tUD3UfVbiPU77Zs3i0I9EbBRbC57CuT+6YasTEM15kNTX5upXJsnrNhpYFn
U2S/TB6Ul1mwqagN2yKw8RY7GdGFseymw6d16WjmirXQMX9MkzeByTFs0x/d3iDwdm2AnS6dCAaC
9qSKavDRtB6XvCyXbSqTFEmhQAxnk2Jy7egH0xWnCaR336oruPnRdL0C93wu4K2oXJn6FZyrVz6L
Wdzm17zCC5uKCU/fkqLyaS8YQG5IZvB76HmdiSTnDgEqTYOfDlY7TgllExXlsrpx0xUfi7YmEbpY
+TeN519Mgye9KdE/0JJYtzbran7dCi6Z5L5FI38ZCr9n7QTg0JOHydz5JFaweW/IOmQKb/EhjkaW
4u5ZX62BlstrnJJTfCIaAIqgSI8Cw4fd7QFt+uGNXXKn6Z82WQQLaT+jpFniiVpqPoyDSNNVIi6w
CpkhH4B0YLZb8HAEFW56VuXMlMgXSDAsWcMq48Kgn7SmplUxi/gwiOEm/waaODUT8f53CKAdUJC7
q0cPdzL0EZM3deHrTNAsQZFi/UKfyyS1k6hVRq0HMVEVXIHQ9ZruUc1TaZatMmOVilxr4dusPQVU
56jTLpjYaRIw9dmhFFu6nM9+BljALvNZZQKoCEMH8SfTlsWbPrw8yRvT4bhGJwpW21p4iDpl4Td1
gkS1L3/zwoq7MmHEUOI0LwuxSAfPBu8Rr8AaRnS7hFMDrNH5ia9IaCfjjqfX77CqWjm/VZP8Aekd
ZfWUUVVDj+TIcxnpBHLmMquyE2GYF1HuM58BmVhNcc5nqWgvnbLLoBW5kndp3utIspkkrGEl3Qy4
OZ8cc+0rULu8khjI3NiHAJjX4vK8GHwifUukzRRbU1qHUCMlBX69u10MvI/FGBBqUMLUN6PNHOa0
D1AuG4VX1pN2QYRQrq7w2+iC4JXW4skSyNy6J4tXMUYtBxtHs8E2AWMazucQDKow8vdIegCQh5sF
5iMyBAo0XoRzBcf575+DPtkp77FLemdmhbQeZuatSrXRUlQG5OqY8u/M6na0Ed8A+Gj5iG6hPq4N
rzRvk5ZjFHGVeBHkSvR68/90uqBXSl5APioQaBjs5Tdgucz7oniM8cBWb/vlFmzBR1oMuTQqRuTe
R/gKp/yblPootxFMUI3bgYLpeojshu4hzXMJC0caFI5T/K+SP9bgQ5rT+DM8z65PYXJBcCDd4QiW
vJqx9/QYGg3J+E2ptVvkFrNcIclK9KikvZrFPT/3oGNvAdkMRZQhv2Uq4UHMjuoQksmhE2LSMAfd
pxDe4ZamQLb992xdsi9tjugPhlWTbeBXMVuN5GaJKLrhxkZpNPdcqDiYAJsYhSR/FjwKsljvmsYh
hqPtSVB3SOrFJmHG17fcBrAf2hh3Gv68AB3xuvDnQxbc8eb8ZRo3LxcIHMDOyiRBxi60CvPU9T7b
MFfeNmOC4u6+q+cefB93P6dIv6RooSaQWx26x9zyQkytUv4XVvLF0fd6QGUB0OHFWEgRziM2HoCm
XoiO4gNX4quIqFvC3C00XAnFVIps6mgOUs8OiwuKcwNvgivwmE0hP+iCUh9QKvY2qeWA4w952Zkz
JRIsmGLzWE3nYO23vAV84Pg2/T1hMg0sYnQPunEAYmi46x2zV1r64oVYsm+qD3L6l5l3Tue/No9q
CCY3NXA+ivxyNiBsncAd5KZxNjAZAkhMd1lcPT+OOvoqbXsLwyP/5F5kvu6zb9AMEhOoSr0iSRwJ
4q9H63Pa6kpaRDYF19fvawc9ImLxnn9IjZFgvEsVPPR/bxwhxScQMihC5v+JgnAn+i6WrQJ2xnXO
8svWx8C4tv7Q41FI3ECqtJUYbC3U93KpFWbh4WCmnWTGfyRv1MdhjxZIwtQG+fJ1vnQytNPIcmea
z0kPeOn0h7PcwFcpo4VYOKSmeU9uu19h0RnRCqERCOF+F8jGZeTL/HGjvfOl5Kel9DICPdPMu5fF
a88sz+TRN4ftBHMsX9DCn1NLBk90MrVta9JHDX33h9NXYeXi5OI8lXoUidTT2ytq2vhzrhX4OJtN
V5Ty/y1kdb3H8f1ttmNOzrb+aybo4kVxIca/N5nJoxyfJbx4TCExr9cgtxE3sJv1QLtbv+OsByiE
JRdVHkn4DQuTbAV2eKyuXxVp7YFqLSyoXJ4mYSNrwwN2pTcyYdtStvo9BX9d+aLW+sCLRDWFY+Mc
KQ5IxCHYMDTnd2CM3v30eGUCtZlaQ5OgmVbadnNVnpyJGfhWuCK5p3bo2tbX/UOfZIs7Go1iPIqL
pGdehrgrOKW1z2z7cPWXmV7czxZcZFW09gqLJWNkva1riAjaW4WO5teXwiJJNsHye07TGFaEiTUv
aPhI+owD2JS9JOwtZ2JCkYkDZgqhdgS1aNKcBnryOE8LiqF3NI+tQrzDhDPA4KikxadSxV7xFYAT
IkAMtmhdBkslse85Vqe3vycEWug1u4d0g+RX/I34ihyQ7hNT5Yuclq+boLBqxd0f0mLny6jnyTIA
QVdonsaHUZgRIDdR6FasOX7xgYT4hPHaI2T6XhW+HFHt9p0RzXgFVEgzM3RKmgUEpiydg76SBmsK
+h5ka8lr15hmUR+rXVEwDk/ffIS3h5IDSB2npggUc9eTV1CdDdpfYNdwVQQhvViFmMwLE/Ued+mu
04gtNAMUtJEIKpUVrfD7rNc9kUCzzgut79LbmPY7LPU65cQBxhdBf3rAk8RTWf0h2v8qzKkXetVf
qWMRFAbBr3QiDiLnBN5dL2/d+/rYsKSOakHOcyxboKr1UayZtoBfrIbvh2MNj/fFPX8Igtl0fyCX
kowS4Tyw2/dE9CBPQZufspQnbFvlekvwXdU7T/62PWLYmvZTrN7PfGLeQ80J+WcfRJ2Oynzk0goa
6W5nz1CMEAQz4tIXvZ4V6AMOLJdrh8PXYwxUCRM1Wo7scp4fpr4uTMWlTAW2gI39WCnM/ccQw0O1
YNhjlp7z6ctYWZwg89hdxmykIAVdMPdYomTyk0Pqsc+YGcCPdhfDRufON5Tz9Tn644IG8mCa0d2X
3H6KNjDuuOCQu20iPw5gNrPBNj4R29aMcS+TMQnCfpH6Ubpi+VyGy0YENLhxsMcohYW/R8cW5IOk
e8M7aW1BJxbUfXPg9G4o6fjGV4zr5geBElE4eDT59sh26nrXqeg1PsnibM04mMSFPhIt4hqQLub1
OkMV+162t6L+tANQA0c9O68XNFxlQwT90/cZ/OU7KeN+pWEYx/jREL/ZCR1QNG7ZWo1TMIPMUP12
LivTqsTMbx+DV3Jyutz0lPl8SDWOs4JaLb0qgG0pYbuvLifHZJjlkYtZDRCALTACUFqVmxgc8zox
CGdfOd31HhGfWUA1pxUMyv4ZjnE7HLsxMcdn8GlQHmUyEUjAFguXgHtjf2EgZXKW8pbJTtrXtOxs
yM6nB8geI/DFO1CJ1V7NJs8kOxByUWCpji0y5iXCgw829mwTD/1kiAlw3SXAoQEc74pxi9kmjfbU
wU47QZSl3STnekeULgrDKP1KZPf31pYfGWKRmDrxvpaFXdIaVe+dx7yobtWfBSz9WLx9m8BHKrmj
3+ef0YtPhfWzevwp4rGtAnhXE3eVcYQ2Jbh9QLe0mI1sqjXnPpfIs5hkSXHsCZcZbcxvb8b51fNh
/LzBrtqy+2R207MA88bcCNKAnAAJgW9QyABLDFSNBmS/9eLW17ge0do6toQhobKaVCFGxy1VgjAS
8IBovEsWHk7FpKTyP6jogtVPvrQiw5AN2wKDkIqx44ZehJoubvAPzzdiXY3qQZ6BLSYQKMfGhvib
oa0FPNZBlSLKZnfOaq/mAV4oaa8ar7PhY6MqHyNp+QWUBZicZaxIjewLNeyXeIWRgFBeoJv7H9Vd
NPC5Ttb6a9xvSn0hNBjM+P+xe2E2/ZSPHkrnQb6VaiMlZTCbjBu7yH9UqiUQ+k7NFOQnxVeY4W8A
qb0hv9CZDj6merP3rP+gBu3vIslhDQTSXRvDc8fHwTxLDmEUA/4dcM8EeLQxUhctn/2inUI+w77A
8NBwHo6fkMHrOGQwg9/5q+0WG0/+fUp2yJ0+iy5hnCDuz9e1XwYJSfJSuKeiv5t/l8avUoiDppdv
dAp+utU7OOIk6VvIYMCMRcfLgh4OzmkPrB+mU6Maq6+y7+HssbFgCfiaULb5gbXr88RN9L+tQClM
Ne7NMLbgy82xUKMgyKZCYF0UZq+eLfBTCbs/KlE6fMyAilx/VbN7rc7zxQTjH+Oyv23ARYCI0TAm
DtW/kW1pN97aDrd26cDB3hUC0o5nSgrpWKS8Jywq3j24qw1abvVdU/gkaAbu6IBT/ireCs2W/CJP
My0Y371gqh4akCBawm1QJp/wYQqwTPU/rusIocxUd/DsQDrRZEJiWh81LfH1ogCJDBdw383GPi5E
a1j6yQ8/pXGOQOJTMqzojMWGsaJZKGjb/vh4On3Yd0jev05QpD7p0n2Ek5qVzxn+dA6s2BuVWWAP
5hKzWcfMJU9/WWFDAs86wPgfOx+Z2FRLlYh7KxA8rS6+u3dSmMm5yeis7EkO/GnyU7u2J9HmQvKx
SntTWT/Ykpj+zgIYCqRUXhQYoWRYEGq2yTh9SfRTMn7QD4wjETbtE84RU596ioYS2t0FbSDc8pM6
EZvPOOewiboXj/hAOW9c5S7tcGfVzWTpUB45tNV/GU7qJZLSfMeq/scI/lB6raiUycHwcRdKsaIL
I5qkNuVkXzpXzwd7DmlponYFSpJOP4kRYNd+T1AnoagkqmATTIsWQqFR6ELctyPvTBM9yfYQeGVf
4Czz4DSEr5fNBl8MqdLyQSHnGzW5SHRh/2QzaKG528ixtHXJHnNNa9yCiTGfKlg9darhJWvIF1qQ
1xisrNeegl6VN8dbF3Udt+NaIU6E6KubJ5vr50YiWUgaqN84BZSta7tg9N0sztPaLBBY4brlU55Y
hZPvlFc199WiCOI8tU/JuqCQzOuqBnMO+OQd2a8QuqjJBaQ7khcfv5R00/OUiHlM0cHPrdTz2cr0
7JL23x6VnS1jR8veZs5NpKcPDRvb6m9vAWmMu9ZvctL5cSskhJTidWsPgsvzpDUDzyPzb5FKRKdA
OPYDHLrDhp7xXfLFxwyS/w4371TnJ5S2eSpBms2/LSl7lrBE2m7lvYpIH/g7vaShG6LfDayg/Hw4
1wqquGjVl92mOe5MhvEVTObnjnD0DhIzpVp+jbk9vBMDVoWLMr8KhylaU/ITmIv4kpwpMP+s+9hp
YVkwmipzkTBtL7xOFFNzL7/YmZ4i+Havc692/4aIutSRuec1+99trxSC05gpAcm4nJHcCKr6HXVa
RMxddkNtAPCvT3/+DWyph5nKABZEjCM8v55p5YNm2Br8BtC/ZUgTAxLV+1in9cu3KRZCW6nzBHG9
+qFHr0+fSlM2kVhnJLsA/kHq7hOYDSl6V6nIH2xQ8fJLH7TsEu7B+VuDkNf6CrGTkt+LKHUF78vn
LZDRqR84dc28PPWWqID1e0ucOAd7dvyB0AxRljiEXkajIRNxIr9rHG/IMDTmiWP9eTUcu5gOb8vZ
/J8AKQ7n21+VuuEEXfCP68gM9gYfIqRIMmihfXaMq/ckM9Zrf38AP+rEoMSYESs+y8xDzkJE5z4P
OWZQkBnIGDbhOV9igRkNyHbuLQHDtC/YeB7AY3rB6PikgZZ3K7igY1NNkhLIsfd5UJNcK8Bx8ljl
OgQoCiRSZNOf95IdypCtfXT5gR+PG237uZ+8VB0mMqjp3npLvPCZtuSZOY/xfwCzzIKFRV9EOPYl
Cvh6ntszp4bCRFkn2RdFs3CGPBmsDTkqD2upkFX5ZUg8tDWTdjsOfln0u4dnP63rtYI1O3n6nBMk
f5V2nS+MsSd+dMIs6FY4VOn4ou3YCN61ekMhiWVm920U4vXAtuCdP5Y+gagP62U1rZFIemhWMvq/
DXTyeMdoTO/257RvPXTmP6kMcUfdYr247V6omO1DI4wzYl0m6nXWXk2WVT/vhuuurpauvs5QmHkL
+Gw7LsoGPpj8q2LUZDrVdUh5b8PEwu7fWC72nhfKrU4km6x54iV5VYBgvm5pZqv299gVj2c6uJSP
mt9eV9R8O8bXqbJRU0RirzjOdkkM0kL8OAT+ropSuSkJZtXtRypD0zcV+urypcbqCEATmfth2GEg
UbrOwqTa3iLMw/rLCl+fRiPO8WdgBCptImWJsO6wwG1jReoNi0nyWoUcqtT9hqXPeJkoX26i1J0E
v/8ag2jcLUQoepRsoB3Xmul1oRrRLjoj+faCN+06R/pxxIFHy2xXbDNa8rVxUR7XARdfei0wqmFD
Oxcrb7Bi7gYvi4SXnjMcxWZy3JGfdcC3ofOyCa7Sw9Hs2khxHOJu7Cfus3Hqpee4S2dQwspibAue
0+p9XS73rWoZyKjeIEM+byKV56c6glyCWFymnKZ4Q+utY9vxaRXrcHOH9tN+U9SJ8C/NsznVHPDV
r9T27UksjA67wjoE/ctCO8GNIbJ/nSaeK/5odb4sy3EENKP2Xd8yO/gm2l21FwMIxI/zsWe+9zgu
mtVDLkmzOjNaghAKC4wgeGPYQIa+DfzOQpm17yMwOJTZcX83ba+lemKP67Xmow7xofzT/51pcBOv
m1NO2R5tWnmqOAEZVmuTMI9hs+camlvezD7sri7eI5S3mCRaM8zhsE+gtqQyIxBPdnlWWgE30RFV
21NlMq+AS29QpNr6PA0vQgcRQeQ3IusEmf5BgowjqYgVR1lugqIuS0we/YIfN9+9FShlFg6mrpno
G+MEgBE0rt10ZKWD5WjdsKADUsVo4h64QNWyy4yj9TrxvFynrV/FoJK3jwUJM+iEfKciZ+snPew1
efqCogj3eaMTKv95Q1cLHucKwNb/5FOYA7upgAghbzU1wYrCT6lmFz9ekq692n1QL7f+2mRGizLx
kyjhjMrsxTbJl4ywIqyR/K2MrvymlUiUoXvMtgDWtE+99dXD43dxmhKlfFhXFG6U8h8qWVJYwGLJ
Fr3PevwkCDZkW/+vSW8fLdUV1d0K84g8bnT06QUQCuwevc5PJvcndKCc9jRtmaWNHuVhxfMTZoC5
pt8oYjXieNtAjjQR+qU2j0O+aDTuFyUBmG+SJanSDtatlZ16JehpLqbmsLDWQZqcDcQWVfkK+VP0
NyUqaHE/qOlnyW+2/MMl5FZ51b6fsrhXwQ4JtJpkhi3S/A9gumG4zdHEAQZa8lsAIOCHhxfjxD5p
/v3SEE/2LerG6JpoBj/UC/6ap7P128U9fVw8xzMckRdbXaBk1SR8agE6WkmHXuRJqtUG77NURKBo
AfxJNni2QcIqk01hJ+kT+lMVxlVnq/LbO1l/XpccJDXWv7Qq+stQrDvZSYOyqJG4mNJK0+r2OcDs
yb+Ll4r4+seYWg+AK14MfhBP0WPdAi92QgCfL2KDWWS5s6lYOYA0WGiF1bZprIxkEAP/PstgZ+1r
p8y3JsSG+i+RQAezue1jJbMgYyfSU5ZWz3xYp6PmFqxRJ+WxNmaZ1VDqQ+GlbUfySQxF1FC+WvxT
p9gxsSjdKxAUvXaxeFkp7K99kl0F9+Mj8u21/MUuQivYH28DY1YThPXl21eFvuJeSc1bs4f49Qhj
X1gzRp67mMUje+DjgybUxH8MQDt2DCrU/eMSB8/oRMGqcZM8wDgSHQSLbVLHdvRT9vUOYqYcaLA4
euk8eRWXQ3oXvFx3ucRcDRz1yQD5gQ8ThYl5Q11uG1CuKEO67sWStiOxxpgeTZSAU2b6fhJjsxIP
S0nPguHk7niaItCzsMLEXd3SHUMk3eFo0OtyR6ca0QGTISm6Yti1kmDOLRDNNqIRKKKETQ49Qthz
3Z5xWOa3F9i5bG+QIEJf4A0sUvDs0zv3oV4dOwakioYpf0BFo9IegFQrII+p6kPWO3Zp4Psx7gPM
kQcimmMMo3rf/gxT0ijqlwekEPz6KmYNQlTEXHZrvjrTIp7BZCEFzF+3h0btPq4rengI/DsSpa0M
FmGTnJxQbwnmijQKTsp6K/e2ODpu2nhKrx/hX3k+qHYV41Gqnx7YCcpCZ2cSEi32t3LSPtBOCo/D
rFuTyLxY43hwplisN9CvS2U90jJmFAtds5xYRLgqZ+F9/eVPOZVEE/61kEOqLQ3HQQmOLGwDW04C
pM4hTxHMWUgbz43W8doo0SbgQIwl0y6Y6gVdHo0UsLN4OPl6DJnFQmOh0eER4A7o6Xv/6dvD0EB8
7buiiqwT7CGPG2EHsYp7a0yVlOXl05Gcoc3Y5k1ZXXjjOPR7pznT3ok5xUh7kjmWRv3gcVJIRJXG
Frc/ypPgRP3mG7NDpygz6OQuSPZCLoFOWQUKW8nnOVvDZXY3nuTkiY/7xBfpKn3S6mCtmbZj+shm
dHqCEi+/Ph3E3+tsyLJTawFlLxKpZJzlsddOQRybtF3gXhlPvw2i+I3R8NVs/cGf1hoQ0+8o0eir
7mpLUzOmwalQwdwnda1blBzAO0K7ySAOw7H9aCw86JiFzw3bqul7PeVfBlzlvVQXW8+LDvK1KQkA
wU/9m424UOFSzhdUd7b9voDcpnLQN+rjWdi0CdRz7vlPTUWHMFa3/X3dz8NsVRBXJpJWTPzICyvT
f60+XmMgMbOPYxqJrvpLKhLRI8vxPtwWHOzAXHU7CG0GlSBYTo62T1pxJwto98hQcKPXrFuqGMGP
HoLecAC6yDkNGBY2FuCt0XC485LkcxaoZcVwp7Id906kr1WWTqMjRo57iFfnkmXZZYfxVJGHtxld
kez1CmysHqpca5imnBxRsFlsu0IlfZpGCon8+FSC6t84zfkaxH21/S9hVewGk8KO6v2bNeVzRVyv
POq0nSDfc6UHdSEDZ23P1u/wWd2U44bLqJYzYbRM4ZooGjMUf0kprVzGHzJ8j8oDCka2E3s4vfv/
OXTlnjZlYBef/Efqz+xKxZg8NY9T0+Og7jwJPh7jhVFYh2ALUvvniohWeRMl6GJNVxMH0ZdERnj9
8VcAg67dJR45XwJyM9D7h6yUvCjXtFsjs7jnxuYguKaMq/PP6g5PhzQdwQUx4p5aeg22nnj8U4pE
tHKlrtibNA1SXnPZSo5ryFbinm9cCcT+HLnFY0Y1AyXANg7gI1v4GikgOQGl4gpNd7X/TCN5SIg6
ssokZdkdWVsUhltUirlKWnt9jvzrXWiCoIsulVOYl6dfmneN9JQYyXFWsIw7HvP56x6qYpnkNV67
aiuGVjITXl/mxc91YMQzwhH39LdWcXsEjRFaF0Ch3Gc2y4oeHAsjkYNZrw1wbwAaNg6DL1/1pXVI
8u+4NSfZAMfiEyrXRUjZ+A9hgnaaBLyKbUe8rochbPXp8vrPvYfwvXrZYCwavyZswnYBM9RIY6Ab
EF5sglYYhKY5BKH7bKOVytsJB5+l0YSYElfa90iZ4ZctIgZF120hLrRB6pOC0+WTdHjcGb0xusQI
By6SI63in6BAUIVYhSNmT7XY5BX2gXb14JpqtMnndXbh3uDhuX3BO20pmHUNmZiWGYHVK/z7MKi7
VdukhPs+hl4ERYCyqFNJPgf4E2bHWuABR+GsPR1vBB9tlE7Efk1TBhdgZzDs1BU61pYIjpotI20B
Od29aY7JXVLaVQMU+jLFbWZhiNOlV3RCFSW/B9qFIp7ysRyDto64FMKsgS64vJBhVbymxKLyxJTf
c1B6c2MThtOsGz2e8dMPzSB6W/bpNd7UASA42GcOQ+/a2aDN2C8jzbedtnFTaXWwYdWxyXM6T0Lr
B9KEHo7Ms7c7IRFSiVLEcXy4UfcikIua14DC3b3a+mTte7B3mJ76Q3mqkoUl55NAJ+yi/nNY60pq
hkgulGZ4+2D1r7Mnu0z1eVjpMGSIzLiMp8e2NvbZ32DTBrvdojfnYRBiCP49HtcjRvzdyJPttUdP
yf8rSrxsd0HoCfo2MQPJ5OoqNiFcj4iR9s/RCXG50hbBojs2sqOb7+3fgooQaYMLM1rbOsrimOmz
OhBqE8HANnqjnPxgARFRZbshcbVtcIMj6OdqnlQSG6rdtUM9nTNjB42FSqze/CJhRbflltbWRhRW
3Jx4h0sN9+KJmPP0Ikt5+Hd0UmPl5EZc0soqkDmbFlZOSDsYrbPCZoEaW5KQYN3PQAIaE18Oli+b
IZSVqiI5mPR9bdgTHNB9kg7JCL4/Jey9Hot+MFQXN9PoYMBSFGJ2igjWH20mgyj9ZgUDUE4bRD6x
pa7k+De0mQNBxpkn5uTQ1jo7xeCOk0Ez61VdVC1Qofbq9xEduio+FYjxFzW6lmUNcHQSDE732nlZ
U1zA46BxCpZr8MFH6V914vQFtjeK+CThHnasDBT61ult/+mp/QgVnw14X6E4ULfPfioRBAmkPLRV
YpAzLiEvgKRDcppr/SJ8dBe9imvxnY1LdowC42JLXppV0156JHXIImiGGXOZy/zzLCeEUZde3/FF
Rk3db4p3XBAlXYy+0G603D+QbX8M6TzhyIlW8k2uEBmdbNOZyYydrAKJdsjKOVXlY+WVVRKNKjGa
eyB6YrIEhshoFOzc6kxwt2vkAzqy4ydVs+6iKDcsUEe4ixv8y2XUbHUq4HI7CB35vau9hADAZL90
WTItzbLZpp1Lkb55WL0IJM57mhcBZPlyLrlSARusG0T74/2Y0WkxDF+MaTAkZzI6vofxmFcxGAqv
VNdAJRw3VDJ4MokZ2uRV3xntF4QWvNFSRGFakH7Sy4gs+LxWfis35H1dI93ieIHHKS/2KFvQsmf9
1RoHVmow95ynLqvTmJdrnI2JYJYQl4uZFHdbiJzczuDQCR9tIClGewa8HKHcJc+hfZbfd+4ZE1yK
LBfAguRBseOoZXy0RkYEHOycUO5dYoHXond0qYbt+owGLjYj3gx25f7+II4aBqhBel8KuPMCT0KW
vC4drqGg5fIyuUfAS/Kx+rUCs3KrnIUHprESX8B+i934uQ2E+vnaZodKyfFPFxs5qUDdYDYr0rsp
Inrh7/sDGu42sczXpLVzAfJmTsvl60tjT53QdmUnugrwBJtTX98+7c4QzlEay9jsFQtPv8afbX4i
hiiLa8ygJlyNi0g1d/n2WFOPb8RQil6AQZlPtMKU4FvRldqNe9dj/NNqy27BHu9+qpP4j91NHBjv
l+RZPJGvD6Wn05Nh6/bwjZMkpGtCKkx7FlYJQKMALGQyIdxMSpHstv4IlzIo3WWCxgG/AIq6OqsP
Ap3qOdcW/dbrs+GSMuk81qkuXiyuABrHoTgRbIYEYUZ7Fgfis7ZZ1nVTb9WngUc5yjJz/a3b6fag
xEBRi/MzYmZ7AagYqGXScKUq/j8JiarFeEoCsiiKtttFBnUNXpH0bN5PbWTXrpGBygAH9LGkTHX6
V8A7ujbwGmSwd5k23npuR4SuF4hdBUY4kGhWXJU9uU2Y7PM0joX54cPQAgdFQMwPhqlTEvsYVJ93
bzNBFy3Sqw+64u4LgDeMsU2oylf8pVc62+NfMYTKPsjHvlGqfd/ngpH1XujoilYu5qOYo5JHNP3k
HvrctI1KZLKM0qNVTuXEZa1A8uoUmjOKSMIOE/8dcvQQjiFjcDLYsaACrze1naGYnuHMwhM9r5Vc
nnCw+nmJA7w4161CKmlTJXuiD81EfohcBxsp3f11jm/J6UPvlJDpfrPPNJQFodC9QS1mvzxuyEiN
m4ewWv/IGRRs58W1DhOG6xleqZC+N9FGqcaPEtrDqcaNP1MyxlVW0B/Y4kuX72zUgJLJoBR6ODnv
JNvEL2CN0FvN6dsXQliBRt7vU+EkCiPxmyzoiyhvyfQYBjB4a5dRY+H+72YjsAROexC7ZGMcLQIm
LMGeFvCZV/Uh0cXy2AMfAt3PEMmlACbChBqvY7OGMDmiI/s9lhNXAOhjjKp5z2SR2DlQCvDdwV91
LFxvJrnBstNwURn/D8MjeE0oarv3gZwUpnOFWkuvIN/yGeDK6nzXUm6TIEdn+vTykqGaLJy3FzeD
a5X5J2tgt8KeBSxcdYrVOVwPr4QWXFEXAVs51JeGv3jern/4PIQPmqaqGRQi1KgipIV6kI7tL8UQ
CKNdi37vDqfW2DFRuXwsBrpjasDSNgka43vBGQ5AT8xNTlYVzOnjDWurrHIn77bXcI5dvS3Uyr/k
Rq6G2A9C4SCM4KucE6ImKqUsPOlMMWlIS9JnXw5JOd0pVyAdk4k8fRGMulQpQOu3BRQXFveJ+SLb
X0adscBEuRj9g+kGX5YwaBgYLyO49itt1LgK1dh5jGRkGvDvHgTOzRHYDRMqL11ZPxkmaKIYRq8H
WAFxFhTfJDYZmmNZywWMzdQmx0atdcDOae+9OaR2MxjhhqJA8d04cAxkZNfogiG9Vt7B0ldxfcMZ
LMsZuzSVFkDsUdvoZk//B28IFvT4Q2Y4u6vN/UR1ZX5hqu5vHRuUHWyI8MqEDx1vUJxTXHdE9Epx
D/WbX9WaKD4SlLo4chq8h0tnB/er05W/+hIoUcxAYIlCjKivNqVtQbrOSMjbCRRWguZJnAtEW5wE
qhGGB2KYyNvkX7bI/CK82EpYP+a6EkDObN+4kPcb9BPzkzGd8BIOSJ2gLGGHWYspwNk4Oi3a06yA
bLPQc+CSqtfYDWLoCpKbP+CUTwHwDD2AzSIPrLtpt0px89UD324z1sFmW04e/mVXBZxX0U0HXx+H
ULZ0crFTxuGn7ghQmO+bKdCCGSOG/4+/4SAqaDHi2o61VmUDxe5eH+g7eYYN9OQiMfkdWESriPNp
0SZo8NzPMFagylHrM0Ldr7O74Gw1uhHL7yikZWHuNmMHw17msjerIQ83xJJabaQI0bdcbRUOombs
Ueb78DY3UbZsZ2FEraoZpHCezu6CpI/vjzXlJqTgyBmDxqHzxg6XoSAW/VT/PrrhYy9MxwMttmcm
aMf0EIi910do9y53SlQKB51AAusDTKDvN1pnipiEFt5zBnKKVInJnP6MZ7MWEQ9oKzFH3IT16/GH
I7QXFQOgNZQDOOCKvp1iev0gfz6VPhoRmp3PBsm+lBf7pUlsVSbPM68z8O6K0HE7u5uU9k2tpB24
oGkJNyWEbefOFp8t+g2SRZC8g0b/nMXtcO0Ggah5F9sqgd6lJ2A0kKlBNTM6Q6MrnJ2BpUIZnMoL
czMX5kT9sVq/XsUhd4hndokVt7/WUYEIoriwl6yCWdRFdKIsvVS652oYeCfLopjUic8KM96CuJcp
yqFS7kkOm6zCgnDXqhgbg3f0IBLbJX/gGveWSM1MvoFoDChxFx8hKA+V6ZdvKz9BYM+cNNk76QYG
GkHspXusmMahAsr5jJ3jw/R9CNx2ciHJzdMuePvZgPsyKchkbN5TUBGUSUCB4ADn3vp/m5kJ4vdj
EOEq+XQyK2qw32KBImdQs3BFfZpyYvesQ2e68RrCZQOAh92TgfXeWuKjrF3g5v3fIkZAGr4xiFyi
4ij5OBtNVgjMks2QUPnJ0IkFEjsMaQsNkIu5EARQk7qpMAYVfmO46MSNaE9+x4tbsfK6RLC2ea2w
NDGfhRy8HsmyhSTD+o6f3SnzjGKM8kXhgv1l912mycjkzrDQ9196DNwLbwYOHRlf93d78r8SxwOU
CYZvrhXIX+QncQGdK9ipLKf5QSeEDfQ2OLrIbKs5y+yMt1dvyYSEywZ+WPWEMiJb9wThCVF4OBGk
1fdl0iLOe1iD/3nQPTvmnttKF/bwyYhtCeOQmsk+irEv3wCCw+1XjTmdAZHQSF+002jgkQKG/v0Q
8Hj0DL2kP5z7/8yeLux006rhdkMbx2N8jSqFzIaOClLkhJNqDm0jbhQ4ttOSklPtj9fSlldt74nH
+gjB44lrS+yk0vEn9aqD0NFe6ZRAp/seWJ4vHrBZ9pMX/prREakHJPXHUR6yAtiNz7BtEkA+lmux
Uu/xHhyKF0iFVCZkSGIm3NzVEW07YSoCsfX4O2TUbrJz/D/Ey9XjuxzH88y3OCeGvT8q5ZRkUcBa
mL+wWiuX7modtb4Kk9HcUV7Ma+aB8x4nnsKBlzEI0LRWeL45IZNrz2BWOAucSNPOfZkQ8CkWV5LH
91y6/oXd/pvRU+3GkPxl/qd4am5irZkxZjThGQ0K8kQF2x8whtgb8HqJ4ugWpOHaLSfKtPbcPFih
ScfdEh6ReI9oMR9O3RYk5z6vt59IgApqfPJPn0sxQ6iWYcMiHyv9sZJC8NUEN/DUx6R1WM1qdN8P
D1flCpuji7/ZkSIgNdPETwklCe4w+cOmcKw7I3Nav4pPgLfsu225lS+lFn8FKj5DZBSgFsXylfE6
S2y+1GnVog9NcNT//ju7BPK7rm9H82vQGCEqGHXb6Mpr7N3U4wrU7lQRVsNxOWG5odmtrLvXDRqy
6DJ4uKUkn+aNmNsXXr+7r8uQ1U5dR/+hPvOY29ER3mWQX53PF1bmnT4ttMIYUY8gzAlu7yOSb8cm
GFflA6KhxkygxFDDySZCm3jmq6EeXrJRk6Ov6hjXsCqz6U40GRp2WXGc4LXn1q3tebqVMnoW8RGJ
e4DN6MwQ6KhO5+Pydpf7w4u5OuySvJwiFHLs9APOyOnm6DpPWtBVly/J9UrSPR8l70wwpN4JImJv
e+hx4grKbJmm8oqIcITDLF+lRpx+GVncF5gx+jd2U82VK+fZzdhoiAd9QcBcsVXLE58aGIp9LdAY
O+k7zhIxckNv/s1rKuv8YBpU/EhAK/Ov5n+wwVamZT643MMr1tBDrpZ8aIuCDUCsIZKe+jZvCOy+
PZDt7jOsZPP2WLyEdjQNn4B6/icbVyNjrqJGgAE//pEQ6W02syZftT+1eAfoTl+vusOOqrMfte3p
5gUsACoC6Je5/2tS4tTiHywyrJzncqfBostzyXn4F0HUIekYwyILn43ZelKvlgZXA0ZNJlZixvXB
EDaOj4/LiGW90Wvs3rDFPbq0GSsBP60ylSRvfrWWymuxHODcQ4RBjA2Z1ueCMGFtUM6gQQkg86t9
Q91RCSsl+JtqG5t622dSihgHsZElnech5prXb8Hj7eiNbv6R2qC5+BLAjSSvpE1nXVZ9rojSOAYN
O9phS8DOPwhbbV0nG3m9qt046YfGGuCHDUN6lMLlBBmN7StMzJXN6zKKTcivYNUiCNXLhDEeL1LL
snTJNxRnBmAcZjAN9v+OY+gVZyFQUdQmwqimqVFAyvmAdEdJS/qb4vOrCNVfRoOz1qrdW3EbII3g
QVVuqT1prmW8T2+VV8TgR4i8wEpJXa9N43QV6g7IkTrObDYSbrR1FHAPOCJQ620RvlCUJShkxh6f
vXSfGqHdM1KtYwqxnbD1rU4ONGECzAL/57dnboNzK8hkFGTEj7NdI3IsqrzuWAEHCjumQD1BvwsV
VsNqOYe3YSALgDqvqnc3Hn3+sZeG0YJJ0gXhqxoVo/PzJ59U+5pXSovSNTUvBEVy5uocbgqGGGsr
i3LGyhv9wOStMbIENH7QAHrEMH6lUwu1sZmgHUr++IwpqAX8xjaIz2wE/1//HWIzxKK79hS8ojzV
/SP0+48J4XGyzGBrJfUyDCpQ6D1GvaXTdEibG8KLTfRrA5xYHrBsBiQTs/RmuOSIBc2n5lhrdFVk
38bSS91qMR/AHVMsZimjUIB0ipRHon9Zk89O28Xc5OeyVX6wLNJglxoYkmD3nmm08714NVeI6cuU
2KmBNT4VxsnrvQXiu7ntw+5x9yNBXzxX0W2BltRgqdbUhnpok7uDFhJSc43Yk71P59aqJQUwA3WR
OuDyR4nT6+tbJgP750Ik8NJQ8TqBhPa7JraVdapGbChBHhD6SoY+/PqQlvnZsnr/VW8MzCU4k4Gn
filNHgwvw3A/PIrymmv1ZCt/V1Wzs6MznWQ3f8xojIO48L7lNeVYSZ2fUvcTmT349xVwf0Bhlhtw
bWHMGejEP6oOCCDFm89OPnRE2eN+S7om7osGYNlgDRW7Dudr1gx248fUGeAB5dMX6D2TpvvMb1sC
Ij9RKkBuaEgDeb9ZPeh8hJh2AgMYEmEDT+ZGEImgd/uCwyVZCMh9/8y/bNr2IEkNiZ+OLe3Ca79t
JCbj3PoeYEmcy3eqGV4BClRNa98l8TDOFKBkWPm+jU4iFYJusgoI8woiDMRcKVbHHsNBupArEbEs
+XVnhPNUSCFaCvwx0P4WuNFCMzoMoMYSLHc+pVFBbSbXxN2Ne0jppXycR+upiC9X9+Mh9nT46oFi
bbw46L1g3xZycZaFfsVwsJmuxXFgWZqvFxeJ51/k9u0AYb7peqc51MxGaiGgZ0tSUyLEs3JVf2cv
+6qvcQnTyf2KQycLv+aABJS0oZRKtdD9PrU4LZS6QkkVJAt8Rpfy6XbS1Nj2+fD19wuhsmqnJS+r
RixYZ1TcR6jb4ZwgJOFlQX/kLUXWXJiOAiH6OSgyn3WwBCocEysopxhm95bKqhYGf25Hlg3b23Ca
0VQnykjlQX/smXt38T8Bj9b+NAjjqSfDcndxt2W8zetWG3P/evoEmi6XIwzRgC2fYkalifLnFEry
m/Ryq49cbAUxXQH+U9H65QSUWk9WnKXKpXm8BzBGrWJy4KdCurFUrx5qY1CcumMyqQqJrfS/neV3
R51Ve/G10gFprf2gORAdTxH9sTeOsuVqQX8FRxEbiiwmla3g9Tvmf1yggO9VBZO34aOXv+NmblbL
YN3f7/SY32vKUvAexzNH3MnUpZwSwqs5/AOz9P4PtIboUueP2wUo/JIAuxEJZt9HsjEqZGlMWPM/
+Yb+t1CHgFT+9vt+CtaYgys0IDuB1pCs+X2Ajglya7oGcyq+kC27Dp1g2r98ep+xZsjMsl4uWMTP
/CDz7UGrKwfGRP+TeR0pK2og+oOWTWIqZSF5CVcHd3HgMMSswSQkgTH/K+2M3x98LLvCcqYddke5
zoPeaMJcnnSkMyspXIqLrAqKQO8iteGkoLL+P+6Os7tFraT6H4lg1g+B05GUCaxl4xTOF4M3fPBv
wLsRCG8m1Lijv8adl/P0F+lsmycxEYQUqmLgYwr1solit7s2bUiUP01Ac1OB81gSpoN0xK/Qlb6Z
Sa84oKr2U9yAmd3IDSbvjuq7s/Of0t6T6FP0JVbGGbq3zNVU+wTrG6Hg+WAv7bmgSupqEm0sQaqM
WktSYLUpPWxZ+jOYJtQJJujk2K6zqqlLqmlEaSqtWY/AOS3vluzJ+7z4MI8F1Hc649gnCB+GDkQY
bGHd9ugUJHRt3NW1s92hxwdudWnoptamfTMULJttXImNTO7NO89ERnLb2UQw7JWkWHAFBahhzd29
WRX6tVqJAiUJHOA9aU5GQ0j68951gUuC2DdrIUwtuiiOwM/qtV8MVc2QV+Uo8eERpyETd5akwPNC
fV2PWirTp/6PesyVwYO+nvBQCmTbBdoeLnHkgBtJsOBcbhspOH6xiClFWfneakxRSriYyNtwJs7d
BwxgrkOyiMIWWU07T8yxFpLR5nxBdtdFMFZ93KfUW0Cmf5TfmpuwFoO4ZqO7GFyZbNDSPqz75io8
su06//7GLo7uRHNehss2OChg8fQNVCsGCDXcv0fZQx6vU92xvnPHuuu0O7I8pvowaEGso4vCYFmg
AWYRoza/MVHo/hpl+BjPpF+B0vrihfoBsS0jHV3oHDQe1qO51mJmzRniQqV1pTapCplzWFrVgWTT
wb2JkBZ7pF4oxlKUeN7ZIqLkj4IqBI+MUXkD8Lf/ggOf0QbentYvh+GQ+NVqFym7SbHVhA/szEbK
oIotfJs/Q2qGysIEB14l57FEa7BDzydOwups1ZmD/LPZ9eNUPpIYd107KdOwPpHAJYTI/lk9Hsfd
Qbdao8qkCKoxoILPkjFND9AHJKqNfoFBmD/nz7vVhWaZK9NRCTrjTZZE/7UU64qr90Uid7Dm6eE/
NwAz9csjNTOJD1j4M9CgAJPa1gToMexKkGVy4NFjdDMKgWVS11irUx71AYjr5body4MRKJtUULV4
GpaO7rtukRv9ATJh0K2GkZ7sF4m7HsMb2xJDhy4I8N0rsOF+FKne6eTktWtktffHoouTcJw2gdtw
suvuIZl/R9LIi2gRULLO1lyd2TwmAl44ko4aNzK/tho4vYtBEM07k22Whg9RX3bv6OmBJfmkQ8h1
Ba4KuRNPWUbBj4xqk3wNBSC7MVkYtSU0TwwGnzmju98LPeLlP/nWPnj36Bs2QAK0FcUn1wzYPiGW
SkgXKW1makVYOSjoya6+UlPIdgFCrS8vIHphQhRSYFy2fpiCV3cvXNxoTDderkkBNENBD+J6QRyt
JDdYvgm5j+fEInyiohOUMCHEj22hcDI3vRTkbuFsn7y8k+hf3ObWPc0VVp0YcA3gvbzqsVlmqGpO
D71K84oiJ3JkOvJAIf3ALr+/m+et+f8efK3pah3f4r2/C+CZXB+pdEjRs+i86y+W+yA9I7UUDROU
5FZuIhhVnmRjOR3o6Jp9RmbFcaFapPmMWFGwyjUGiI5wt/UIfEIQFNHLLZgCzGQIeGOjqbsMqJbl
TLHHwAfgg+l7kzHqBlu3ZN1WsOCto5HI3yB+8gMwnl2pjOlTNo5NiqHol/HHNpHFHdeEJTzRhVEq
/ABQKguUWWnJqYAx1PPFyAXBEv41tsaC6NlFu3+PpstQKdPHYIAAc0psFIZL356lCRDXl3VM7973
HLdIVJPmJ8Ap3dBmUst4Jsq8H8rtmgkelTMbmEe06zcjJg/rA41bihkBzaIfPY3EievD5ZEAwDrT
e2BtPi9drk4aEIonnRvPyrtHg8WA41sIr0KSKeVJTR/PwaDLJ1KsQO+DQDFBivSeHqcTFTvlBqk1
Anr7kojexwruD+L0ANfaJEbVD7M6RuiyfjG8znJosvLX4Zfhl2fZ76x4AjEVkajBmtWT+TPuISzU
tIJejBKI2rzy8yEvg28/wNu1cFQUJycNnixKYVJ3jg5rL89XhyJaFv7656vUvzV7ZLU7htKo5Qxy
8aoBcG3vg+Umtho2A5ouwzGBgHlibQP2hUT4O5FogBMMabO9KWHBhht9RVRrJT9rSOudZ+wnLxYS
5YwG48Fh4jH3DjB99ELVrxUdgGqdiayCjsmKJv3eSeORBJ+I26orUCw6ueRmUH6BEr/0vj5d2RQL
rUKP9nhRtix4eaoJdh55rTGQ3AijqX9KbKxRdEnBzFcotTnW4q7nSEA+92k9KqhtaIvMVIG/Jzrt
nGyFhLLBTaRdR804zhHMXHszQxLyLiX2qY7H8qOBFnPH+FsjklMTMwCNWd3cnOiAT6r0YizGmQZF
QTmjvJVgxbpfAKUFG+uN6NMCXcwdoN1URJcFgUvtrpyc+uUTAqsah79SRvq1GCglBn5DrMoXAxCo
XehWNaiRyy7T9AvlYN/kVW7yfBvgmb4yx6IM6WIz9Fjare7uClWKVXhecM2RCYSipf0vW6QYY/mf
SPE/TgvKdh9ZRZecF1DbNSv4mZzdZ7CBBcydzjLyZ8ZNfFDZ4aDSgX7ox/jZOatecMODHRKu6EIk
jloOhqFudEed/27PhRWuufjJiOkc5g4bdYOKiOmF9gAWmCIPk56fflHhCPgaM78u8jm6FmD5JS3z
tOLyg4MORno7g6Vb4EJN9g4/93ME0R6GXatntNJ7KJpOzKuaMq8rmbcwYuUTGb8vruum9mryFdRD
tNaUsOGgU/KHJpqiDwPxaUfRpb42d9R52U15/gzJML1d1OG+bRhltSe7xts2uNafHOK6koYCneOb
jxveudLD47jvME89CR05WtHeFaINANOTc739Jdx3m4bYFxmHRk0trDp0VhqEsKHGSdpvOKNjpRUm
P+lXdtWxNJm63BF4wieoTLZ8UBd5yyzhtJ75rRxTFLILclUxHlyGbFBNtUrZ+GsPv2RzQXEciwJQ
VkQpYQ+AG36wQAVEaS7rU8+43bpvC/LuZiR8NzvkvXdEDfZDv6DC7wd+WicSeCZCzqPte96b9YBh
/SkF5cZ/hENQCEvw2DgS6Z5lIGip1EaV5KroTClniabke1D7Ejbmq0JoC7QwNSAYhBfWE5/sdlUP
gBUDaN3kMop0LfWUClRFdiD/cn2aVooU2UjnfexC9IrSVrt7hPyfeFBMnjByRtNKhIKE5HRe4qVi
xFnoYanakMKCAYBkfxk0fflZsny+BurE4xM3eHAY4KjURK9fZDbBVH7qk4x+5+FJ/x6+KhGzjpod
HFnzMHGQ3cqgTgdGwAnJjJnbawcXlw3FL4lGpE8upIHURJ0rnlecnSNFOZMIiLsokaG61eZxwjRk
ZSfHVqvOyUs/yAJ90VK/poNrlJSr9ymTqu5p1VWGO9dDpg4xGrKpd2vmy0Ze0jWd7ltMSYWDiqSF
GnkvVCbE3k3VXiVQ6aVDsmMy1uz9BwTuHyL8Q2ZJBaAUbsTd2nSswY6J+Paaj+VxpU6tq33qJB7X
pFkxbcFWASdbxcEEv7mAr9B6VO5P0LBeDnSMfC+gnSbDq7E0msB9WEYfjL/33sBaiaghbm8QhI2V
eyynpBoirumEJyGDa3h//xJ0CGX1juhoCYvmycmBb9ix3wbwx4Qk99fpuUKdQmydaS0RIlTTeqyn
G8AjbtJzLnt+OoBs6AbWtBFX8eKxVDdwW+bIJtY8LovgZZpny0rdOSu9STlxvp6rQZ4YGjRCf93Z
14m3oyAwpsFYlyQR5e7l/szAJ350UH0tFBB0zSGlAlhtkK/06rneCl5G7B4TIcd0lFi2+63x29OR
IUOnUX8ggtxc0XMvn4RIoFtXctcwdfWFDyGmhuR6rlLyLSZJ9Ku7bNjQbYWjDJrUDZ2MixgfVPky
LaVIfVqcGuKZE6M/z79VnhQ059yBsv5dVwoH8LdgchiaW4lvv0UGMX0WYVwESeH/l2oE2aOklNOm
CTBO8VoAwGIreijIYu1B5LlzVNjggFHfPSr1MaFru/SxWpTlRYj8b7uE4U/v37Z7AxQRToVWZY2o
YU0XeslG7TvU5X7VL5ZXJMpr3lHUnztGj3FVBYsT22uECthA2LhMypQRyKirEhctBBtw4c/sPx5Z
4DvzsDJHQ6ndlLGzTg+LuXPH7kbegILpbOBynuS2cfcdOh/PpDB0VXwSxQDWsmVYBTS1nr5JS1So
YbapMsCE+0++sPH/l1rkRfCeb7UAS+rtSEmvs/c1qBrstw9/JRIkW7JUDU3q51zzvMy9Wol1NN0C
j+VRUxH5RjzkxgAGBUlwNVZYYbNterMZzeNV3uROp4XX3ilpsCHRnK34KsPkCwqmi0ljAZR7FfXI
GPGbTo5wphbmhqFOPG5X3NDrlK15wpYwb7zxd85rmpAmkjET8XmqqugGAAr2YZoRRAHbdMQGbuXU
OLwtdf/Ugkw/PnDm1d84Eb/BbOYvmT72qYpdtaG/YRjWAX5uaau+pRn9xXVGs0eOs1Z/IyG3v9Nh
+hh1JIoRFFTkvlwkyCRYEEFWnbDj0bqrGgUuMlspuOh/oaMZXLRd4eAEVv8EnmOAxbrZGd/wsnq1
V+Yta68OqcAluwvGamKmB3wX0Z3Hw3P5fDhMZgbsTweiw+mh3hgv4g/c2+RnkTLZ8yTb7htNsoDR
tngqvi6hZI++ka1DCMZm0REHCC50zItmQcymYFuQOypUFEC7onGzAmF3sXqGoAnUQto4OKe6yUbJ
T/0pxx3uzYwXei9qHB+vQx8NNQEVlugMojywPp+WCtl6b7rTX5JGQ/t8Wxa+p8UWyDaSpYm3Hyrl
IerRq+xfFIvIr3dQhCRZ++MBbdUk8cdamVqQ/1BlxSJKmKHxPVdg8LNGC3pfQwUem3JqcVA/HHH7
g3b6m9rSCxLIKfX2qqIbB7wdXTqOB90W95XDlzRBDNMKDGoUdePko6BgBjpIfJ8ltGaqBBrzHoW0
r/d6pM/JPX9uaMFSlGJDykESr1xUWD4nt2aFiGf7Y8nv/zykRR1P9ht9yaX7hCrWhv7Hk4Jx3ZFU
7SuTtoOv+M6teneU5XpqD0H0FV7x86UmFW0g62DzS6BCLBgbZU7q5agaga22I3aDx4w7eFYHGv7x
4KLSde5e0yxUr4vuZ/7jsEF8TJ0d8eKcXba8rhOtLK9j68jaSWtET9XPVEjSXVu1bA5qOBcKH+Tu
RhzBK6PvOxYtO6HA4S0NJ5UExLZhcTLnR2oq6AGZd3Kg63Q+CzPkZQXqVarLOTNG8I7LfOyzGBwi
Uv0BTfzPy1vjfKd2kYMPS47TgJdggvOzslLZYsCTMCeKUhFrYfrXjYiGm2Ax6hGfxBMJeOqO7Cce
QqSIRpZdJ/4tpib8oui0nUuAtMOCgH0h2ykNQr8wzSli05A+wxEg10b9HC9dAcWCuw2aMBS5pcA9
w6hXV1BswjlJD51zbSPfh10NXHlctIeHDwhDRRtWHGP6YB73WLBoM7dJ5wue/JX1jDYps/G5WPvQ
EhB+5s5vVo2QThuFfmwu1Nuu5nPaKJ2En5UNt35PKIuXerCdF7UNSejG1Qs096Z+IbIFYwxhmR4u
2/YDFm5bPddLIPb1W2Qd6J6lSV8aRv3Z9RuNDOSsEZgzag3ooSKh0N7fewXXQTlQ/C+SP4VrriBq
QK+hRx17OKOwgroKs7yAsfu6MrBRpA/J7Fs8LGt8VSTzFvKlMb3+boHz3iOyXWsJbCCPZw7dYPrJ
R1tU36fic8L9ZDq0MM75+wi0TkdXXup/7EcijmE+/YSQHl8RgPaOMDO3dZ8WJTeDFnEb/XYyCG1E
36fjlNuVRecD8p8rzU2cgAN4/QAhqNgq/Zb5TpGksFzxlGl4KFsUzgwiVPuMxDtWw2gTE0VlxkdL
f0LUl7avBBmcnyZZ1Fazpw3Oac4PyWQ/hjmzYxTvFAgTmA00oqczFNTd1XKznA0kW7nxr5fRkYQc
S4REUAmXfcWuj8+tWVbvJoSGwiNMuQw8pd6d6GbraM3LfjTjoYRxBkJWk4LbyttQk8kPwTJJQlla
8zpUptoEMUsMcZzYAhbT5Ahl6MuL4yKX/rDLptsgFA1HswFazBz1T6mvIjuCQs+2wVV6MbP5dAmh
SxHW36qoYM81ULn7aJlNIKctMNXg17GANoTVGZl2EfMiWgcYEhl0WDCYloSUL/CD4f7Jq7dpY3uR
1DaMNAKwRMGLaRDGwjsZELzuSUmdmzmvq7f46LkdQVV41POuxLcrTcKU1qx4rS7kel4KwN9+BJ+1
kNCTOZqFXkeytScXjbnRIcu/8uCR6EqzLNO7J3HEJUwm90N9+4uT4WKJ3jiIbe8s7lljLUw7O2sr
IRJqvYFMlLmkYVqsMUFkGBQkj/KsNSjkQyvMUW2lDzgkb4BhwjimNWK6QNwmkoXOk6xL0VDr5YPv
2QUwU2f2zVIrrvvS8/Izz9hFFSWyOlRU8ZmefUVhtbaQVIMdrZl3le3nGuuGb0FI5ETUxQeaBPwE
3u3w/b+B40ZpbPiIyXe0WA56pOemmP8LraHYR2L1kvq5M9q0dNYX9dfVj2DyI/OhLk8vwSxf/QrT
3P9I09kcTqqyXsh+0N42MrBAn7jFmv7qCCepcsUgKTIPkPqtWjwaohh4zm58tQJupZuWf3VK7bUN
6+vhhsIvXTAIEI9pZ4d0NgCdmvzlm/u5kMdazVU6n+O7cZalntiyKGFBomIB3BU6yM0C2YxVRyw6
UPUgYgaxNXVjUf6iErpS2OfEhE38yMyaG6gv9mvQwRBNWSuku9fCha6CuoZLhHxQJwSd+rNM/bLm
OpbuDM6PdG4TJX9VTdw9a2OhnKfKfR5QhC9q8BgeVquyicXhRFYN9bDMF/GWXOdl3ep5JF5D1uAR
t7n9dMyUjdwJJ+bk7q4cgTlNu1A7mtLpfmE6sJtwtlJLowK1rPVFiFBeBOpJcalaoMiLePr7LkQ8
1tryv/pat9Rur6i6Z9tp+t0d2hiFRWjoJrSBFE+lYxHFBolp+HitP763iZqS7yw5QlnXWKIIKCQs
fA+aYGxE617X5zYn5AGFGu2e2ngfxZ43FXYNufxupiUZ5iDvaq8NqTyy2HHULU173YAITyDSEWj6
mG0YWSzL1qp6nO9zhhjfSZqUcdBm7ITgU2pS5WC77UNUyh1moQHCY2BYg6j15QY6AYSrH2+2P1bM
9HZVhQyrXDJiYDRJx9vFAAY1pZQswvXHEGtQyxtMnnXGHlNvm6vWZAv6pNV0Nih5OqQWpSXIWaRM
8c1sFgc5OBYe4h2O3h/fD1P2kxK4PaIoiDOoKzF4ybgYurm7KFAu9B4w8K2dQclrZYyfKgLqjaUZ
LFbSpXUfU4YbzOKtUsq9vXm/U8S3dc/XODi/B4MYldGYYBsdtSmiQHnx965MFe0ABtCzDuLIVL8E
s6+Z433Vaut9igwEQIfIINEmkOiTmU6w4vVkBDqa4+W77lTCCt9MAW1xY48/aWihFGDs955WEysw
4jaw9iumCJKHo2yN5dP6ciV3KTCJVtADnUmxcwAaX8ghVmGbBgvqnsdY6p2u43sPy+VeBWOy//lo
46KHkt6oLD+Be7AcNDwo1R/BcEK8ryu8uYPTnl3uIR+N75hLaLMI7Lsp53b4liIgiDgHxQISe1Tr
fBzEuPIMQPUIR3jwPN+3431Lxeu42+2o9HMnCAK2pIKBWsWl/7p4laZA2Ahb3zAxZ/tSJDb7lOBc
LUeE3OBPoi8U2glXJHmo7v7H0Zs3dXVKPTP36MOM6NxGtrsRgsy6gMxQBHCykPGYs+hV9jFj6eQ7
remNRSxRbc2NnHWuQzFH51g5z41g/Z48tFhK9iqjbvaK8XGb+VWBOduhQcY5PcPrgErikjzs786h
y9ax9BYEJJ1oVAmIKZsYcNnsZy0RMa6dboPwR0ljvqWNHueiXawifGzNHTQUS18k2cuJE10XL4G0
m0oHX55A7hrVKvy/vh+bXUiCsz/gXTrp4vYXntcWNzGK0HtwjjFpQh4EJ+DHXYLbo/qcJpesMspS
6inONB/S+qeBUN8V1IlNbegVluw23/vPYVWzK1EJygJSVhVk48FPkD9EAlmh5eYfP+wNiYQlH9Xk
VXlkmkXngGDbrTlnj64hUKyod0WkdiXquz+sjYJKJeYdN813jFE3fFVlkaebAhplOkZ5ndvd7YWd
RvrRC0quy4xcgL76RusUJ7EFVk0xedE+0559qDQK71p7k72o0rhuYpf2EgCXoxavIj6RTpI7nlGn
bwwZouyQz5Dp6KIbM/ilYdRtRgYLNU132PQtYv5EvOUD+Et9vRHxnukyHH9vJ7jpdcUHexzXZ39p
6oFQYKcvi7N5yQpDZngye36+YuNC/qpP/zBreh9W8I8sfxj5nHNWwmLQY0HD4V75zj4hD4MdhE+/
TTQA2C5/Dd9lWtZ3wvEKzq0um6YZyAVq+2hAseQkIJcKZpi4K+Zw8DguiwF4aC3VB6LWDJXZHCSC
SGzI5ToqFHc+Jk4idjoy+G6EiGuQpK0ifkOvXP7n5Btp0kDn4oQZzxLYw47jytV3Nl05CZhTJIqN
pZblX0oqB/bR58VpctTDEIxx0c4RsA3x6qvDWceMveGBTNqt5GotKkBrLCP0e+K4ZoW2cOFehKQx
DcitPi6mujbQTqHjFdEmPoiqAJUbvis/sMGMm9zzhrkti+eX502rzksyChpjRwpSb/sxFwECi+YB
gmGFVSFEw9LXoTICF/MTInCUvvxl12SPa2hnwh0b3MysqUAN57AEED8ZHSPhG9YRCO+YghqIru89
WwEgrq/PolrVa2rTD+POWwknWFtyWce+Lf9m2K/PnkVeTvRi84IcnnF6kDcpyaOEmodPjhFPWBB8
F7Yvbt91C6mcfbPMagsz7sYm4euqHJUGYk0xnyS5+aqnnInu3QoWCoXNItjGW77ZsXaUinIwnAnB
ENawP9gfY3EnWEKqrwI5fYIQZOuTbMqvEAdA6a0NgJAa4VnNQ/1HQSF5n6xzlxFgo0U7AZmZUtAH
RDWSIsJ8WCA9lU0Xk2RyMCZAyiWtH2V4Ole7z9bdQBDsmCmwkehi7aDfaRUX2NUGf5fuHyzTT81C
vJwrz9YVa7DETwz2k1asolDnlpqpWM96QY1qe7n8NOxa19lC5grcX857dnWVLckOCzNKIS8ySero
OTcaMYribhYD3HE1MkGlf7PnO5hvBu6ISrCGSN8giC+N90BebNHbDW9bIF9YTuby2uHZPB8pK4ca
P2dkuYJNLwZom/DsbrdnEe7epUwvHH6qQ3rVm5zeXdkg62C97KwXrlimvegnfeP52JnN4/joPHim
8rkdeYULNbwThfWHkDldnhDOfSmgihLwul0FSlEe1Lf26KWeAGCHGcOCF5pH3UY14S46Tx0AAIcl
FaJb/RnzCCjbqouLrArYgxrFoDyQThYB26IvH/8H4WZXjIuMwmWKSscVoeSWDH260Kvvn23aQWI/
l6imzARuqBdsvLu0tS7DWf/jchNX8pN89xRFAhg90GEI2lrr1ykrOo46IahUKr+U5xnMS5fsFhKI
401WDnRTYlz3DilHOy+WRLHr0Il0/YdsT9/Si3u3Lz8QOPx5x4i/WVEyCdA6UhqUDmKxZhRc/tVr
fa6bauQSKcVgm1YnSToN8Np0kCbzpCNXEqJPTEBKE03Mcw6Kdrbvosc0lGhgbRGxn8jLMG3RY3J+
Sev/j694U50i7B8jqLM4+MMXWPM5jAcPmhWv/bsdL1j6jylgVWyOSEy91wBzOUTX512ZE8RyU7+G
TZOeGEfqSsQIsaMUWJ44dfGYTLu1p43HT66VtTTwFHXHBd5rKiQYDPzVQAyI9Lrxuu7TaQ/4cgdN
kD4aAm1CZ5blX+qaHp0NsQcjbLWsneizy/0G3s8bdSZBNglMCZ5ZT9RPU8YT2yqYBpaHy7BeowC1
8na140gZeH32GqiOzKjZuUfnwJ/4EurqwGg1ck9Noctn2UxK3RlrMlR3yTGXyQAMXTa0TXhGeWq3
rBoSb5uVyhvDPJw/3iFU9jUU5ceS1CCXeIq48qW9LPtHVHYZKO/KM5JixboO/Zy9SEHV7vysqeNP
r03jm61B48p//eIOjDPiyxWdpo71piPQNaaAfXvdf3EwBVT7gwrtDiAZVjrVrCVvfqTsEXko/CvA
rVESOyF/pCqqpzdWjklOIWw0VZMNMMTq88hvTaUap8xqckjvyDdDG/g9OP+7tBtG8JGacNtEnxS4
9oTrp8E0rBW06aaZk+n/jPZXClUNbNNaT6moMc5dWj13+pX2C4nXZHmnMWmQDNu1YArClFKZzMWX
Q5QbsR56yKFpDh6Ks4zCaq+ferm8UvF5nvqwPeDRj+lFoO06Q7wDXII3eGU27sP9PRyFS8NayxoV
V4Z2+n3gapkJY6hZFQYcO28Z9qIY8678nCqXanH4mvrupfUHvt73AkDlM8BoHCHyh+1gtopcC8B2
soU1sHJl5MmhBLH9ZqRM6AvJFVIsgx0N7st+zW8W72G/CFbY4S4qIqI+DYhsfao/8Mfwir4bOMU/
+mSJrdtU/JvM0qAYtKag6VYzJ/u4hjBJ5XHX0BmC+JcIMlGGRybFo2x9AkdwJ01F0sKyYeay9U/3
jcy48ecwJrHaSwrEkgRQ+DnK+BZlVdjrh9GhHgtRhNtUWreMsSbKjJT+uJiISQtlE1C3AAhxO/JW
A3rRCUP394Yr92A9oa4Wf083Uz5sr+bk3SDBLeskVDM4sKE7YQywxs2wTd25PvikGiqDdY+7iAxq
han7zGGjJf8UYrSPxfd6t7rCqh0qyQ0434e/d79tNZ3SkOl7PD8XaaWTo0S/XoaIEec1s8rIoa4q
RHyGyQMs9k2vtX7Y/fk3ab1SgusCVEKA/+9UFtY0lW/+MU22AbO82jOJiny48x4crakatl8x+FI+
Y9+2LDewFKGRXUAXjxgzyyJJq8mB3EdUWe+LaN6t1BZ6yApD3WEzC2/bwx5iw6knTyqD6x4dMd4O
h2g1f6eR41NXkgTYZBi0tWzAS4pnoHoIkIe9M+F/Sv8lGIY+U9RGfc85lYzTcG7GBPkWAd0thXdP
AliAfmE3Z9CZVSkGHmwfaMCpl+0tQiLPZyXLvyUed6uqhOUWEyQsO1oyWLwqBCqQw3xmXE90DPm2
6CgTIOkIPFCHlZxXyUFifcxjJnruS0IYNSz2gxYd6NIAG62k7fWgDAXKWXCRNYe08ZU2dLGNOtUL
HFc/FDwCfp2UzmA7nGxHxEo4f6HO3+L1dQIL6PQKEs8ZdGoQWU5yp9UVYUV/kySOg7Ie/LTnZv/3
Jh5jsBrGIJMLaivM7g+4eSouDxHCPDyzUPdN8KB/n5wGAo9xa+88TejxIbacyIturc9m0Ykyn+GS
evihkeW6WEkw/8xQeyRdcb43oMp/gQiyAjLHJmgQBlMapu5r1Wj643tE5PnLAIbAJx9Vx2h65D4J
FFjUlkIHLASLkVcZMTMjtBBI8deMQch43U9l1QSkjoYFZtQqS4fvqKwFkgbjF3cSwVLX0BDhqtOJ
H3lWnBrJzwGmK8h2RnsjCruRHFukUf0wIev8aRkyBFU9740DZTDSh+nC3s5Dsykg+HstZx2h0j69
c2WFtxPZoj76oCLlb50LisDP5G1/L2SvKUur3Y9FRtCvDazavI6XRnRkPSD1tzlsYsxA4aiH7Z29
N2dRIH2CwA6EHciYXIFAQHGn1OewMWXgwSXRtoCWOa30UW73W/5e+dzjftNgWr2TZlxI/21+NlXW
IYlz0kBbxjpBSh7WNhUPB4V04njA4VIimJVX4aDkhexR0C/nXIJW8ImoSDcU6GtJmVe6B1qh4P/h
DpZfX8kEqXl75LdoEqQTHVJCx5h9IK4q00j2xWOeQb9IiZ1QYdlNAKAunQfdr1+kuF2QNB2pci4A
KCkM0aWm35FE33JzwOlcDigqZl/CM4k2tW85MOsG07VSkasKKyduu232zMi99QBv7r8Z6efpzj2/
wPOUR4FTgDBKDYS+o6S3o2Zi9hw8PXdDAScpPNcsgpYqUvGdoMICoNE4B11Fy+B35UCWngoRJWHA
n595BMncsmEejb2jufY48BkcEwphEGKi3DAJUEVisD9ZvQGv7wgcekvCMbLkYRtCO4JSbLhOAggk
vxtxV8JRmLNSwM84YyRXXdAE45g2I6LZps4c083v8YD3DNjIVnsuGB6cXqLJ1tqbndkprm058tVj
qMJ3+0yfE4TxlCOzLYzk4cYix2SL71MZi4MCzmy2iNAYuOI4ZuO02E8cTxNQ0zVLfwLvApUOvW3c
emTiuQNbeQdz6kLOU2R1iSgyhPiteNP20LkXli77neUFchwFyyr3lP9xAN9LpcJW1eGBDmeLwO4f
YY8PmvNLio4VcEFwz3VrWg3cyL+6Bb7uE3IqBWkrd2Kwwa+CPaMJkrUV7CUl3rNu9Im9fz998iqT
2ywPTTcNX6uE3EUo3NeVYovi1WcNc0QtjxWJkrJ0pO+qH4jTz/Nvpv8Lkg7LWChav/yLxAgi4Vuq
DjB9OAkDAPZPUN3fV+szRm0uaclNgvyDhkr2JGQG9waak5Q8ENumP4OadMSCaYmG6hqXozgW4/ym
1RuXC/RC0gCcw4UQvq+J9RGwi+CgtEHwZb5OuQDzwjmNCAZaSbykg0QxTh8xjxw8y6gG4kP7B51N
dk5MwMItrvcmxmGcYFlX2FE8Ue0dPl021YfnWIm7pX85fI0fD+kVrApxW7P5cyCGVHB+6BjrMdky
6E0ZktxWF6A8WCIBY02DfqzA6kFcZq1Sjs8D0kZFH+zhrZLHZ94aVKz4j+3FMnytvdluSn2b8Bs2
sxGm5YkADEHm9SuIYHVF1DDC8150SWQ9TPcVA7vRW/aati2tTcl4Lny11+We0X2nRai6PW5HlfOR
xeYfOo6c0Pp3oninP43IGDNnD+bnJZTK9zkbmh4J5bDWkUu70Dkqv85PHAUVguHIPZSADZ3/4Dzw
/EHLu3u1AVrWvgV4L1+IyRErO70V2TVN07XNOuGtFceKZ1HkDhbp/OB01Eqq3hryuSVckkHgW05R
N4+MyPXLk3nkEIRKOhcP/s+mejLUhyArDKNjR3n4xa9W9rMA/9w9f/C2JMeyQ+R6BNp1moSISkEa
ZebcEV7a4a5PdrM8sS6j+DZoSEuW5a6p7pQgEiC/xwx8kliw03gUo/Y8Ck+iQvuu/K+06kp4rHYY
cN9WwjQa9zJzlu+2oAPE8MUkPCSte8fDF5INpLaMnr5UdPtR4QqA4zAEl4jZk1SrN6Vn62qfn1cw
E2xOdgX7X2hBQ6UIwvu0/5RycFqQ9ZQ7I2cl1k6bv+Q9X5iUrdfjdcZk3eN31af5b/JTDz5r4a1w
QofargIx7lnbhX+qCCTllCggTvJxpwHTLYj+eZYAYwi1dtOxRwO/M+mf28x4EpRvJCLHFdRpHGBR
SeuQrFbcMmrbaaMybcaUnUPDkEnqcjqVrfdUaBY3OyGVpArNMKKbaMiwNMxdisAASsxYeIv0qLqQ
axAEATYfqBNFghuhs8Et/MW2vm8gLKJrYT+lZHHSgc1gct9fm6IxqRBnAd7WuLJJOPacZKcVkdrD
2maFBjX7ihO4Tfr1qjWFN4A7agfMaqj9FkcVesXR+SIQOQdCVVkP/UKq+y4WqFZeDJKzHvWZgecC
H/yrVpcEpjf3HuLjMtpg/btULtRMIW3tRPvwt6AEyxs+0S6TNub0YIJdynJgsjzIFUMOr2qyf5GA
DikxQrm+o3/Puhw1I2S7Ecy48G6iYMYrw+mpJ3nc3gLa7LZy2rkasMzx5HXmyXwsTPWufFGaw7Ay
oqYrN5BHni9rgl9T8dqtFs95ipTsydyNeJlOecG2X/0qaNJ82yw+VEjVwOnmiZTm3BkXXCsCUodQ
RmCpO60Zjaph6rTRNLTHvR4G173FOyneywvrdiFr+31upCzmfN4KbkiDouiNUG7F0utDSJSqhQTA
L9bKm/KACwWaDVL3NfyuY6kd73psNQEvADcUP7XxtM4TWz9PNhPNUOQFDtNY6lTVmMFlU9MXtWpp
gwoudCfQSURePRDS44pPwRxdxHkirRWcpqNAdawyJHOzsRMvZPrWAllVLgGzwgaEHN2dOch7TRNp
YHkp19CDettOEV9Gr9igPXb3qoLqNZz6Hg/RvP9V/w0+BR6XNdsYR97Ip4YKcuzP34ZOHQeKfl+G
LDbDbmi+Fjk6VG2faF9Bm3qVXGzOCTz0gPKefLhgdHBip00L1fymX7mQ64Ch25307FKTZZb97Vmc
AJLUSL13371I3tYWlLoatVnT1abfmbFuM7UH2wIKHPJnIIZRehn7NdCCu2N5yVpQMb/uQC4w6PjI
1NsTlrx69RfFFLdtguKWXR/BImDP7UVrDVZO2e1z70bYa/L8euXw91vdo/ExRKrpFGGMg3fPJcmc
Qmz+90vF1LHoRnosVlZaN5qTpCWT04ZUbFMxvNAHjVLQDkCuRMtpToJRYJLWtQpluCxGmeNXQC8H
1lKuHAaBK3zqWCeE56vbrCdW8mScDwL0ze0/JueBomN0RY1oCGY7M32Fn+wg30u4dfmg8H1TADzO
MiFfvrn0ay5A4D/vuBe/oTiZLbOisVByTyRMBl+CodiXmlY26BwYuKg7VaDttu1HQ9JdGmKfOW3o
iJkaSz15nf7TjYEbWeZq4++JnT1lLwcElOC+ZcuCcKezLilM8GszYBK3JKgEdlXUs6KnEZQAKDT1
qU3XnVy7ukYh+ClFHdhvS53UnCFSzuoNarLj0MtIsQw/7vBRf7bOSzXVhq8dQQI1ir0Zk726HZ6T
HdpmzQP/kYrDijTysgYR1hYS2+8zg+OMXVJYupve7ZGEtL2y6U263s83mAGBuSJVqCDi2zdt4so8
rl3yK3H3gDa5DjjNHzIdCBGh4GH1Wbfl4yfoKgu0AdXIfgqY4uGHVQzEGCxBkQEKzYyTzJ1g6Fee
PdvBGPoFAynGUssd4PS1FQrJVw5QpRN4BgYVkrvmWfWW5E2152uSTebDJrDsyvajOfl81tSi2vUE
Lp4lahsobq+eBXRyjO0GOVqvDkuhp4gY3uBpWLMDyonyMfWURFTAYZXLBFIRHQNcIwe2UjoAvGo+
IVTV0kvaRW4xRIb3wTbWOV6dQrd6nKS8tVTe+SApYMDQKwbWQzoCKXIXBPk5UZsHqGegMZVDnRgK
MrUl5V3HynBtYXb2/EVFpGVXO+E+37W7AkkDMngqINFLIKfSNVLhtnPUwNVNfqYV/VDzl9yqNKiz
3gPBXeDq6RaQeA24y5TbjG4Ngv+Z2g6smvQixEldXON/LZ8Y4VirGvgb2D4p3eG0q/Jp9N18N/He
i1ytVVn9omqIjkf8+FdxMFm+5UH9OzVzXlMfJbCsegDNps1pdX04o5mQUefN4xOyuRpGsSW10kx9
bj3Z+iZAsMjgFv//IxNz1+2QfzUPzNlbB2pc5PdJC1jKp5tVzaIfMb1M/3iiqjsbe7701k8Ekn8A
DDk75jeKz2lNN4TuDBgI/QJ1YcfyHaZEn6llWV4XWA6ZPMs5VU7Zg1O3bUb39IVFV3P30DW8k6Gy
eKUbWxIQoVYXAAMtjzCgFzV9BEAMiOQEi5XZ6WMv+OYzvt+kCXBfVgna7kpCRUS4bicczgPGyT+9
pGnhR/xdhY/HPNdJ+ydT4a4JDkpqLP0+/3Z8jU6ai/wZCSNSI3pIo90JV4pRkMhIpoCt8HcuMUtL
n9CgpxQnZhvGhgVMh4JYuX2wm+h87pCs1ZdfSHTW5l4Z+J3tWsB+p9lIwgDxo7VWvJj19+YAmHni
nSEg4CCYb5ycM1WGr1agPJYJMSczZntrKLPyHHSkVoy1dFuM6VHjSyH+FAwmpG9CboP6canAo66+
K3HDHZLVtWsi3KdGeaMjRUHGAfm32ZsWugZEprpBbftvulW1OtJRM8iJxQgfzWchYPxWs6qiZJKU
ZqoF3kS71ZMjHv4ks5tvbm8EjhoMI0xzhou8N0Cu1d4FYC8eykRCGysHPSVQsB+8oxwwEK8fr6iu
CXPIPm0Q7b+7F0HAlDvnpcS3d8oc8zgCQb6KXfZ8ZQhZ2V9thWuJ70it+XiaZMnWX5YxFqgJgQQt
vmH79pkb9MOBLCUmmhjyZhEO9djUM/iGuqHT7+W2frWaeyrcFID8TuykMhgkx5Sk+vxHd2OFHQZt
CV7cqJCHWsnpI4oyzgS33H5kb8UXoMz36AKZULeC3PgXqnNWUgEp9F1oLXT0Zf3fJhiDQIlPtodZ
Pxun6yHUfvqL97R9bpAalZrejrpUSPz5pdppUbSAX/e0je5fFAqnQ+eC7uq35jd0fr/oZYKYWGIV
xACWwZma+HfMGE9Z5bg6OQyvoxVO7ZYf2X/yaLFSSkY739b69+l2LSnQws1DFgOTQCuqzFQYohOV
mXEiaQygglBVG/l4DHHZf8kv4D96XeiiGoQW+FkIZ/yExd5B+EROJJ/Nh7cNCxVvROVkPpSqau4n
S+Bru2wRWF6dfPRcqY6xPBG43c0szdsaYE0+zHuWuUEhNU/tPav+a60pTnPUe06u/57s97FWCogA
qtWfy447ZimNq7GBz3FVzfUqisBffdLwnRiAEttS6Aralmm5plk9pJuPBcxMcY6aDKd0J2QAgyN4
DBjTFaYOZR2WKw3YQ77g0IL/EWRob6MOxBpLEk5qk3QKbXU0D5vZET9C5g3JrkQTdwz6Y/VGA90F
j0fVFO7cVhzacUtUufw91O9k5sRqR2pp2NDIAnRQfTawkgCDmXr75PHYN2JJnvXWJM+YZD7RaOir
ZDitxqJyIacVKgFMKlBvgG6QK3bOXBbnTlmbP2Vol83tqxSetm03y6wq7weMSNy0eLw9/Rl0c4hf
Pcf/ePUOrULRfPvJiOwusW3KzwV8kOZCtFe1PDoS3YM9jbk+/dx8L3Wy+iKPviV2Hy65n5lJcNhv
ToX3Li0vXqPohKIB/kqx93nJI1NMW9Bw4J83CDJYOTL+Vo64YC3NdPtnFeyy08kIATHNoumowMIu
Mbb2pwCtbBTkeDKBVK1xJh7KHPGAQO4VyYD449IkzjXDIbDpc1hJVajfMjJ9H0tWtsG4BAOx3rHd
o8DEApHV8ROvU8D2ejgLCRNW/RTw+7UYwVhhyYvKA9ImbpIhq1Bc2xksB9kLeugn3OH8yXk5QZuy
G3Geo47cgF/UTVWp7y0GeOflqi0g8mpR0gG4RjW4nlwI5A8/R6HL4RhwMN6OTunlteEP/ZrXxO4W
6MGJj825KagaYgpVfZHWrE5ITmF0DdW8pEK1x6mD/mxey4KqxNlWrOAkN6tGPd62Gk9Dbl0Hi0Kx
AAOZX1q8/Ib6IGSibNvm4ndpInKrq3/tyXTO0J3K1dpiS3NuTBT5bNHjKRHYencCCKIen3GSgNPY
lB0MwhQgsLevUvMvaisnbO/+Rr7q0J9DZAqAuyu1KRcSOXi2PtNOpB5pLdZfFYEK2Rz/ouxiEWoa
0Lwwi+95L8HHFuQGRa/fitWI7TFsY3NIzwucvsUUSB2Rc6fTaM1w5nlERuQRR7r2gK6m9CR2giJn
Ex8iOMVGEu/hGK9Yqczrb6n1zi2nV7mwB+/Tqs4xrif9Ah0vg1oGH3YEIXeUvkWWhUknRt7HAHI2
624DacFkfIYYUEtLdGagsxXaiYyh+A7yoWA1CXGa2XqC6oLZOjPN8NyLg5M+qAR3YPdVnkBy6ltU
IhYKOC0uQnsUkh0XtIaRKEuONSdxNVPogY+oSPCdjP+m38jNWEpHW3D03ZTD8DLlufFVLHaA3hed
nj5o5LhHJXHtq6b77GG4y/c1OdoEta/+EfcEBnwycS9+y3CUyf55by794y66vWZYBYpCDr5yvRRl
Us71cpqInkT96lPxh19ft64j9KjPoO7bniUbv465sjK+dzKZVAOwBmcbUm1V6u7S4EAZWlWyectv
FwFCh7c0EIch09BOHJ7mITWruoDzlcNafMUEoZskUB747qpymfIZER4SNs8O5sGnfup2ETZ+hU8w
f10ciTn3PnJi/NTJb+HFgv+/TA9keFGhDedf9Zx63DkD7zmt3YURetWgegZzsxlfcp7ZsgwBwRLz
gEHlzh4jXUfwvBudZrdTJWvKi1cVQXcyNWNJKc279+jrk1bG2HA4/OyNIqlXvn4hfZXqqWq8U7Z5
tfD5pWtGrvQWykFAPDT+CnF4TsAvR5wbjT3FaUR03mmb4oOPsCVTiFD8IDbU+GhxVQKV5zMIflaS
3/anlThNLokSGwsJI7U063Pg3PjFtzj/Hfd6/gzz7mFMeGbn4sL9sEQ/DLCuIIXxivpyHl3RS0+d
wE3M90AEDjST8McRxuzdF/NFsISO2mKtvtLfpC6OrBZY4kU86jUtIS/7mpJFnxOWUAR4sTUBbVi7
aVrHBeCLpy+Ak84mENHwWoFOQqeO1VA5YsiWQ/qgdZs10CijNnVt2l9J9f+Y88qBTGkW2EUiRQk+
tOrzswZ8+gojml/xMpYiav6w00pmZnsT3NM0onZipA8MZ3QswuEp2rT+dnxp2gDbRHt4DCVrpzMw
1lIkBbJL0OCzzA2Zf+iuQqiuaKTU1QbovglWdqjUj/6h9FlDPU4o8pSFLf50GhGis1C0mwKnpYCz
gyLJOU0ho6/vWJ3kVUGAPQG2BXD2+0LZJqj+7Y+YQ+Z836X7k2EMf1zoR8y1ladqHxQe13d5kPy3
WFulOI+x4CCOX/Ii1t2bgki+Sk06zuw520EDOnm+M1+IRhQK7jmYm9o1R8ap+xvfW0fIOr157TEG
fLUYw1dDBzisAwmBoIGgEfBNLUYZXi2heg0Q5mOmqEfUxHDHM92zhhbQRE0tVRLBZs2sfOIl3Oze
gc1idLRoAz2ge5UBddOjH7zJ8+q6bQPz1XpDAtr9FOeilvrnLn1niV7GCTHe09FJ0+Li69pYXz86
wU/eCCakAFDC3jhNKPB00wG0BMHGq7G7ZoidaErO4678NQqcZz9+ikmFie/KrxDCVbDpYfwRTZAZ
WdRFxdgU7T3Wr+Gp/qiC346vl3+i97tYGg8W7wugfNHDbkNgMASxkqOPkYGjE7zXwmsI8mX7Dave
6YrpIXt1QIrqQW6KsHyy5ehmmT7eNsbiBbcl+GgyBnzzMyaYgaCx3MyznafdBvyTA/Eotsj0OgDg
GgDvJyIYZFyC067iybvaWV4VDOrrM+mA/DtRdUY7Y32Di1coPQs8jFs5b+hosvAb0IhoRD0YNBl3
kRt/qdS9K9NjlLEeyG3je1o9fTqhzQeq4xGPKMouE8yRW3OPYVLNIxcJGnET3cOFZKCDc9u1E0v8
o80PrYvliTMAUo8TDMqbNWAN9ePTLnAONh3+GsTM4+oT/3Ii1rSS6MXELNPSLw87Jj30Bvwz8+we
EvWytlYyO/pY3oCRdYoi7TDGwR1U2LBWrGMYzne7IJB1Mh1BRQrbw+X6o/7hxVzlDo39RQENd67a
u3ciTsDK6FejOnxL07WnIjNgfwMoXikz8T9xsqfbOdw88Czkbrh4NlwidoLBbRbdwfYDcktmEEri
mFh6T61AgmWs16aWqAu4G8dODgRbSQqh21wosjGFSlXcoD1W/hZKUGm6jChM6Yjl7AkBKYEA3+Bx
aaQAknsoDOfX4BlH5RhFTvNB7TBwDGNeG0tlKmsbLm4xnr7Kkb3xByAUgEF55hNHfbCsgQzj0gOL
ih88296YHZhUpP9uMihlwsOxnlPJEzUc8/Nz2eRKFur2NzPBQdN47Y+L405I1hva5gbF/rO6MCmx
8szqlX2OCemyprS8JTry4sGbJn3WvkwkuBnrzb7NM+A5303NKwRjjhzNQplmlhvZaM4w+v0PmYXt
aNsWhZ1RlRUeBXrjmjiwei4iWNABad606dtpUugLJd4CRKztgm9Vd5Vvc4hT/LauzmXt2qarjsgB
+suuzBqdmrAxXro05F9RI/8D3eVygiNu3eGcXgn0W1KjggB7wxxvEF9GnThwrjaEUF2Im4OuIxoF
vClL2RlPcpWbCznBWlvpuWbpgHhl2JN0bzen4vX/ufY90+yQFRv59m4Hc4ni2zKqCvZz7i9qcsVH
FUiJnE1caqa7IVv0r/VSlnpphFuNHET91WccMR6o2RtqTbekj5s6hj+2vAWhHVl/61FPtrl1idxK
zMtg8duImOQAfkXEyrZYSb5oUUFHa2n2F5K6Ba7QWowQxmEmbvCfC6h18507vdUWgUfE2j3CVhjC
w+7fRolJ3u9YDYQOLykengnUZ05tMeNiNOUudG23SLQHiBWHZRfeojbgHQ4KfkGaxf+L1ypPqHHz
HdjjUY97G6sxqmBo1b37B9bmjguIxrR5lNo41WGmC0sgVw2iGvEAwU2OLRer5SbZK5vNdcgEJTNG
kh3x8S75Ygn79e8hyy5hWuyAslCtmA0/J02qUqIY/s8RgFycs/Q2jiPghrXriSCnIjBpQ1/qucEA
HAShCgeqDh1mbxXr1CzqEZ078CVqqGrmt0fwBkjH06+t3jLJxj0H+Ks+hd83Yo9EaVjgrHuPUKPY
UuqnkwQpl2vY6C+ZywHT4ZgxUKISlnNk/Fr6qf/TxkRNn7l5Q1iVv63Q7jBiQiLQqIkXc7zyt/Ci
VnLg9z17kPampOadelYj3QIHEAYBjYLpO2vSogm700eNgXcQYv4aBrFZjxT330tMg9j8Ye8iWiJR
10uKZkKCHsQvTgzkwuAWXX241PYH3MgknyiFTS6VcY0+ShzzNp2YZNwT+Pzz1qXzEArZo+0xHhbN
XrUzYPkxTP5HhJMZ/+w2XQBAnNy5m8oI6vxfS+HkVMYmU1YH+Cchefn95UI/zkutgN5PGO+bxFgf
0kdsYEuPqUBQkVy7ijDp3sbCno8fn6397p08LxPzP6/WE0P/OrRmrwe6DQBhBHsqIK8mddud8+iX
QFDUKmKGb+JjeE52EzewPoLmQKMDj1Pvous42lXTX7Lrk/S4hTBN4PdRW9JyS4gWtq4LISxKxd6f
96DR/cONvz8XEd9VvowpaRWEabFQ9nURDCL1xgdBPVX2l43fYQ2YOXs+sNn3hubUbBq5S8bFlY/U
HgOeELjpX6scEZggmr3pWSriXUsbZQBDTz8v4Q+hayaQKBd4PDcVC7zHieKFtC+ykwYshyS/qtnI
nUBLSIh9/dqnITQIdgOVRR6Z5Y8bKzL+2gsGo76NnVUuYv/KX+h8WFHkCbrhkW5qBweeTVamJ6Fx
Bb/rywawwvASIkyOcUMyXaRfg07r74wUiw90seiR1GLG3T3rtfYJkohXFlDsaIqdO91JWH5QDh1/
Hbbu73rFxWH6V2uRrg9m1IekGfe7y15oI3hQ8TfMPXx/Fp1ZuaKFW8Vkouq7oQNVWgKc3l3W94Cn
N444S2r5rgFdJ6F2IjHoCZUi2ODl1EfyCJxEXYakU/MODdSKgh2cxi9L91vgkecFw2+swDbKSU74
yNe8EW35F+7NL+TLn2v8MwEF6+y/NopxEHYr6jPo/ZWDCOW1egxMpwWIphQxULokeXxOSRjv9G2E
Xy484a6MIfnDvSawpI+DGIen+urZw5EVKla2jx21ezehVwTBaG0YBNL5w6BlSMmjXQDs+nOjUZJD
pAfsrOwrKPAwjCUY2x1xC6bwHTSOIXg/YIx3yLu2CAtxHBkCjjCsWCW++XQJSEHy0XIhYiH/5HJr
7MXG8J+eHlA89Emiza9Q+s/IZhMgDUru44SWXAfKrQmg7t8u4jifn89l2u54jOVS0GXewE1QpPgB
MM8oFAoHxkSdTW54NlbyJHWA3OHob4+N2N6/4b6UbinbB7kTcrkqzbBMSqoQ5SasYKa8PCDvNohS
8raLqW3Bnwx63SaNAwtRKZaSrqPv0epWgAEp6pJKeuCS41ExvU37oDo8hY2KmCegjmRgfNWpTYZ1
tOHw0i0/efvJKcGn28bMeq36AX5UPQm9bGaWtWR4btvQiJU5Ucry+rbF9oc+auUhlj2bxxcOy0bz
NLXg1SYYjz/KqXha+SZjMja4KT+58XkfsyzD/4vbLMvDgRW9980m+OsfiovtUgNRDBwRfUveS0yM
RYxcqW/PniMjL19oD5kzL5PlYEV0CUCl+Uu0tAvxzv5e5nzBvAOBNeWyImO9HUbleV2fQmjSigyk
Ee3lfiYuA0eyaV2f6Mlvl+UjFO431CN3DpCemmOKehSlepQtftZwKcsI7K79MnCxBVuDJGw2fLG8
rMKig12Ie5PEUHHJkD8OKOmdTAryC81qzzsWUJqg2PUFNQ5TdEUSzm+Wb6h12JsBeVtknFmq33Ov
1ljxxQI4gkAmtqKjte90zgBXWuLlwyhwOKt/oL38JRQzk7HONEwbA0qk/x+oblOjRWrDk4aHF8On
ah7cLMX6UOVZFS5hux6+NeyNtKiEtCzssFejN3CJDp3wWSVSJV0lT3fY/k4VLA8vPtdM7S0twe3Q
UyaX2ZH4tEFBZZPaajCk4BTlZJezddcYdOEtTagm6LQ6SYMvhasLJcY9sSKzb/42cBC4eT+1katp
IJEMVj2bxi9g7eHtWbbZYF2xLiKvsBOjjDHxeoe7HZ34JVwRfRXmtrYGvALdcozTahCxfB7UfR/k
36r+bkrfEftfYXnZVRThM+jM2U7uUg+1xO/mXnnkcQDWUmYLyprYvdf12whSIhLO0jixOd7A7Nqj
PriCWc6+6nsDbQnC0i4WOvoiD5vm9dwDCeAOc4yTOkX6wzEn5NJKUYfO+sgrZwTG+lkZnWmmkpsM
UUpGz0pBLHoO3zF1l0lT1XuDvyGto3aI5zbqpD6Kd6JTyoaY2CFzSr6Whf7dDN9ojKlPpZr8p49e
hzXSeJMw5aMorrf6PzgQIhp0cnoTEdP8EoJ9jmMGtaTNHuSjl0f6bjqaG8VqdYru5xj3KL8wHB7q
+gyfGiVUfWuSKYkUIBveMEWbBJLNEhoUFrtoHuWk7qDFpyN7fiaRtvWL31418UcpO3NMpYY1L3rG
8rl8XEFMvOrY/z8L8b2pmQW9/aCZhd0Vw7SZ0k95N2X7yECWLlsEts/yS07qshOkCC/mrCtT8tTV
LLGemIOLWATnXZfxdhNnD/dN8VbTgSrxYmE1L6AUOlHnpyh9YEOLNsNOwmOD0XexvwjHIPLDQ7CE
nKed2z+K1urqhvz7wLNzJQAH9yWKZlqbfp1jt/Ass1z5R78EK1pi9Uexjqcs5FkNj0u8JHYTDSpr
OqTZPzxS+PwBIcC0GLRYj1prpFJPBhrKWsIZBOjlK8hNU15LX8Apg2lRuSg61FUxJaHtW3ptxlcA
iUBCo4B4Wutdg/Iv5vnog6LNsAGWQ6v+0QHDuCIjV6YJfJ1fLJfq9AYsgWfAlPt9pd4LLoun0BVO
aNtIM7K+kdmr8+6QQT8B8CuVEIlUlA0xzWAui/oZUAZOl8gIgMYi7f5GwSb/v9ShAtYrsLoHKCvu
OpvYBEyeoAxeTCR4U6wuleJjTEDIfBgQP96HJEf56i7PvX3ELfA/u+ZIXjZbSO3C3vT3LbduRu1h
QNEIBXcgobxNlRMIeAz+gr86SywDW2mI1F73xBI7IdjHYFa1LBvEhltByqNwNc9xJHzImvR3SBxo
sUQSSiEaqYHJ4BetbvPRWryumQAzZGYJ7r8PVlq9TQsmxp3rS5xzoB88MZJySm1MeU1kF844vOVY
5rO8EN9XFCEklIXHfcmif5Oc4iQD27fvXC4CKslarA/Z2ITCIFizt4oH9L6v2vZn2a6607SKKMQm
ZXglB4puYnRCJMuIKue3h8MGiE+pFdlVtNZHohsE72B3NBF26Ams6C6x6jmcH+UexGC6BxdH7PGF
KWMWXO/BIvOYeJjzEz7JooSiwE/HJqrCg/tdFT9rsaZtqiKTwSMVrwz4yi9hlKDWLVubBovROZw3
jUevQACHNPO2SKlm1K0fpRTzjBFbXtKqeCbG6Z4HqoKyor+ec+gUmscwZ89XKV6zWuTDXSIcYuSs
CY5gRQhYfUrHRJplxPnZJ07wulHHa+jYtU422eZIvOyw/AtxvtwFnr5nWI1oUMr39RqFfO+7Uhrp
bEQUOj0k+opjZ3nONnqvfnXXafRDEkcW52DEfO0L/c7yj2248FdUfa+6dfSnmiURxZBFZDbhLgBZ
qqpF5ntMHLjXFR+mXtnh7wCbUXwhCNZ2cvXFtOWLlhcD481UgjViTdk6Li+/cCPygET/Pp7PG7+O
d6meJdeafoXpkuJEAXzZLh77Q79RQkVB6nmh60Oz3YVNDT/MtDQhh0WfNP4pDMvs02W6mgc5FCN6
vT+eXn+JR92KktMAKKDk2pw+bYt52JJv5z184kTYSAE5Mrsp9d3Pxg82YltanxSkHb+huwEK/937
R9NoXp7XLoqDE81Nom4e/eFkTOge8M6ggT6MzIfkmSc3soplx/Ivqsgw2cEl9EIvuKWxl22URqaI
/fWUAyF2UKWXTvsTmnhhF0V6TBdo1H3UIe05ZfbzU3hxEy+pL/MU5DEDKW9ZTcGcutrrCxF5qYnw
6xrc3gVOpxGzulKZyladjOBfUe2iASldz9jBhNh7pqZMhvdO6Jd+FHsiSV1OPcBXgvf3N1fN1V8v
hBQloJDdFn0wFaLmvhG+ee2/JOinTYm0MP73YYrrHky0/0IhmBI1mtDXF6SoqkGvD3kNTChkpl7G
ktUSf+VwAR20Oy0pcGZOtjWKtPOYB8MC3Kk1o3aWuRglKKWPMdZ6e1TGdsKSSBdQbD0WQcM27ZYE
LE52ElVIMJexg8i73ssww/w+veJi2kPDB2u2JoPWVFfmoBK3BMVPh49w3u/+N5oUqzpqtyr4K6xM
v2cHBl4kmGNmEY/6u2h2nvXVxDAvHfkkLSfnQy4mceOCblmrUWWTW7wUkGMp5R/PyKfpSEcf4Rqh
foXEpO4SJCWnr9fcsT4HSzwZ1JbTrZ+4tV8+QNA5AIkdhxf9rU1ThAZCQcVeNSh6+C9mKZQ+mUCv
5/w5X4RLDyMMMELhdOQb38w8tZapq9DgqXoLwdovv1HzZclCtPd24u0PCJXDvyUxtN55+8ZHrugk
2feaxTAFNisylmfMb3LbjRnrCYMFmNst5cCAYrYQZS7PxifFl6ywo8U/g2wgcp/1KK1PYEsHIY68
W91aTvjj4dWQhFewzkoNj9Ox9IRAaMv/GxfmhSuv3GVy/zRX4XLaNc+zVjXrn7iJq2uvkDm8sGbv
gbP0zW464Mzj8DAguVDMRcfmbcXdu2pLAjokz7zeUhs1UsHX+lmHUOc7V531RLw+SAzmbiN6oY5+
mg99GS6yUaqQcO4BMAtK7+83iTVGSvu/RC8PGhDifJsLsknk8kbcNzz9jyEJfquJsTmd31VjM4P7
irsF+91kfcAid3wB1k+vae8qiHKh3VoM3sniptDkM2weeERpTL2B/nikSZzS718klQNIAB2Q3fgG
UVIWevBOClygXOWH+/l4KgNzvrr96mycGvkchwiRQl8CfhQmXmBB4DIDRQax36BfItaUrZXtsZPX
m6gb6R37iucDPeT1uogde7sp8WGKffu3CatM11PiZBIVJ+wGfVpep9yzwhu0mrrh+zhko4yTlvp3
L7ROJIZmoSrqyFxhCm/KrZSaYzkNk6tuBmiyrWXgfYu7DZfluB9ubgT3j5q79N1rm8Eg/Rb+gcTx
d2PbuLOie/CdbgKenOYAZAfGPju/gPNB8a16/P6+SJ36DE2o6jBbQF6stJoGwrIy/95vWK9BrzGE
BJURNDxIhEQKZylXhQPgHYC/9BSV+UxTUtW/Cr/f71CFWCNZQ/SfTT3sfE+YYWTlgL6I9zedxSHk
wb8Fq+HV2705fznGCD/PHSHdNT9ju5tGEGsviEuVtXieIE10WVzB14EWiSL/y+YWawDXni5Ojd25
kGVxindwDMMp8CCYgEoeWBVxlCbcBdY9idiyeU5grwnwphYSz/K7wViPw0M2P8Hp+woaVMYu9YEy
a19ldPU8+AzTA+Y4RWNvjjTgS/8eIYLvBO5+Sw5A2ZbX+C4RD9ah+iIHPQrb17VQqLrl4Asjh+lG
ZgXqyvMSlT4WK66zif88t3YHgMLvJ82AGYQwZY9RKMVT4sTjTCJhmJT0tyCoND01lsgXIINlYrXu
SsKLLLDyZnGBfU+mt9PpCjTy0joM9ZG9NtrPdefml+zfb26/Aha1l7ZaoNNkuF1Bj55LobeEWfF9
UQbmeQLrGqOYyRlHbB9CKQiBXkmhTJB2WgrUuPoHcBrpRUqAdLD1dLteWYDyg1fALc8dWkcf13nF
7MDzFoIoKFpOlUFgLUXz2L79Mc1FNRgqvl1JiZYRhVugTzEQ65/J0TqcvtOgnKsOqQfdYzasIDvA
V3hu/iZwk/Vn4UW8vUwKVL7Ieebf3dY3mvimwr1wANKlwo5pyf0tHbgTcj/GpVoYnoeAXMejqM1y
XdI1xmM2h23sJl/wLmFA6fAGHUXSmJiIA3NFZfomB/pReRBRIWot3my2zI4d17tdq8UmW81wrvDb
PBym4xfZtSvxfjxfNOacVJDuh/QQW6DMnk0L+suAGv4UGxLdjFe/FVP9ZaYxH4M3/cOLhhsSVtpm
mSMPlryTSb1PskdzUMK+lnRIMcDVADrue1PTorKf85okYQns7qz+c8T74JRN8zAFtS0fdxAjgsSl
ZZEXn6Dgforysg1cHA9w1T5JEI2wwwn3j4oc3S69FgD8VpmlJoKLXiKlwqziLMix+2cPioocuY6O
9TEbpvoJ2AjSQsWeS6ND38GQCbFExc2QC2/AhN5ySk4O32x6JWcJfaB0G8ZYBSyern5XqCqzLwiD
vbOQknBUbIorJcTfQvb9U9KFS26I4VE9SpD5dd5EMEaI4frs5Xb3JIGgwa7/Q8PFr1fu9xfsKxtL
gEo9KEBmEZTktT2UtIZdFznX7Orgf2FTfA0R/l7vbMjNCLMDHrK3a3p1w5IstwR06aLi7DxmBzEI
z3AyW6mJ3BBCPUPHd3ngLYSIMfd8Hdy86IxM0EH0HX/lDiXuJnlvMkp7N9bri5BSeifGn3R5SD89
h2KXewbyyiPQy3FTKWF+0p0u8SdDWBJ7R/OFRKuHhDUx9KgiJ6OD8RyHhIdRSLmb8uN5pKLyE+Dj
Poi1Dr3LMhKEPMtzdUMBxDNnTYjsorYISgXwSROlq2iOOTYTrf9evBuC+EMSGXUgvkh/YOx+tLNU
5Qz375BTOTfWK9nKEu5CiPZu8LThd4JnzX7HiGUI3xwS8I+RmENhWVZilO3LQbdTs4Hcr11SDedT
Rn3XwOKRAxAW/gm4E/jSEYLclk71QBlk/EwCJujVTtXLitAHMyxAK2A844JjBWGcepCuCP+EYUK0
08oIYGpi5POmAdrzMaHxdtzvOGV1bc6vdDH104GZ32NBfQDhZXDagPxOpMjSc4GAjcL9Bb6zHKoS
vFc8qWUQU3L5YRPKZI3t6m3k78FVJfmAll9pO4XCF2y2rogMobEzUTkf/vfhh96dSR8Bzb8UfuB6
NKKM7zw9GPaqXFvZSBoK5n/vdUxs4SLEWrpGoTPUrHL4Lp/dvFe6cERC3ekD1cbf8QHdKFxAjI8C
L61vLeXpnH5+fHlNa7GMbAjA1gkNxXCyp11uyyiVnRTDEfJSkgMyqBiA3UlL/N5jUZN3BD+gsLwG
/UFgIanRG0YxqWJi4tir2ab0Wu2cBTHUUie+pVp+Xw7+zU1ONYoa8ZwU4aTcnfkjK3igLH9TzA3T
MZ4RZBqxOseLUHiJp1XxW4XeTxFBMvNWZ8HQ+rXYNu4FQ4Yp4pu1xMLclWGhTI9gHBFjXunPkZ2b
ift1EiTuZCWPSu9WKDe361AUaCV7tZkZD1Xa0ojQiOoOXoXAYaoCNPEclhtYmQ5cgleKgqXwXFrM
f9KtUnMpIvNEpXEi3lLH7yAyjIt4vc5KtoVY3hoi2XtwGWuG0m0JoVmAaDFIo8sokXRGoAWY3zxi
Owip5lnHtMiSi0uV01DggkhhiZ9f2O7TpWO74kscu4NYIovRBub/1p9j9BPYCz02WqFViRjZiiJ5
eJPYC8tDRNDQxkWbYIBhr+YEiv3Huc0qMCrImtznW81RbsUqfH8aygKWIVIvZmk3ADp5vkDyZBWd
7Al2/d6HolXd/FGl2nTIDfO8WrUc3xZfoe60MFUCUv4yml+hxrpfKIqQmzntbUSCLIexPH14wHlS
chqM2avTeim4NsXB2QMdDrbt5Xm2uC/FTDpcOJ8xjGu+UsEZXeFLfrS5hj3O6FqrNEHR3tvbTkn+
EVUB6fx7QhgBlRpP0DUyTyii8+JgOPE9cqRQxISI7dRNAOrw6Qq+jLSG0Ux+sN3QTbTW+sWW5wS5
fn/Y5qppJj91+69lch7Bsq1ZFnygsbzCK+UaUcvXhYEvorKfLntB/DVSZtH1wi0qWMiXw/sQUoGH
l5i2rewt7TSc5xlHdDeJoZTQYskW82cVLDPWLtlQ7JWC7S9QLvXysiCjgCXSBUMkbavKjOOMAHGC
o8ysXGdQTvYi8kl+eyypsDRfI7nDwXHxzcofMztdhvP0QjcFKkqS5yYHEs6f5wdxSpOpnFi1rT5o
0GyWgFTI5bFL5es45qTdasC2zri3FwvV+QSAMs44Pjt9s2eeemJ7Rgatpk2xorxQEOwifMerbVMq
++ydBbHKXW6PMeBgyGlrUvNBVq9uxycGUXaZelaT1aCKOGfQPsbMNxcZZmc1E1d4Clg2sqtOV0Q3
CFzgeKhBlLGCeVwwwUqzRVTsAh4NcfjBsXqrW11mlT7hNxKxGQLJnWPKUsDoyh58Z/Iv62aNW7Pm
/V/I+bcGXuOmlN9bcGAdGNPq/X8LvsjvCRsoI8Du3F32Vy/x4lQryyZASiFNWggbir32OOZJ+Btg
6Tj7iIJ4DufusPqurS+Dboy9T1fyq6DA0muVoTNOkoLDYtbp85th7lwNXsj6D+4yIKdzAHei2TLp
smOeTGONca55o+S4Y377j3+In1qViYTtchUpbelloXx1zhfxURsQoZ7jqy4nn5EUhzVcYB5xoCim
1btNyHpRQNfwjwGzrYwKYe1hr+wtmegWvgw8T1URcj+0WPG9flekJEa6z1DMuwWZpgLlRzvvl9os
S7yq18kZZhRnoahC3CbSBJlIydF13HSws2pFLKfbCAZpiAjjUc0Q/RiINWFqD88VfeqbA4QoMqf6
ugrrorDmDfhcZHOGKNhNEGc30uOanedvb2zureyAOWoJGW0EbpfawxYRT9nA1rZJ9t09HktOHVwo
Qw0+jwpYleAqUEDvoMwtGa+rurzQCWJJK+pBC+tU6zrTcok2lX3vnwf8IOsFVk1AcK1iRK+U4aJE
VE2pcq+ytl4Bb4541oBgVvWLMVuFZpyD2uR1//ZkAsIEYmRJ/IkTWvKvwF9Fpnv3hEwekAf9jNw3
aiulYmYC34o0Xe6VYH/0yQeQL57ynYjg1Z5zCNmBF6kK8sdvibPYFqjCQ20vygyXKxKvgxu5MDZ3
+OygPfiXxFoNiSeZvBkHy5C7UycgV3WTDRPieQdX4Unwoo+jqOxQXeJe6e74gs4plYBQkfXqYhSh
ZjecTDaN+x5wxiD1O5RhE6ks3NqnehfnyHIfdYbVOt788JoqqqS+3cpbJrhB+w9jVGyE3c9QaOXs
9h2uQn+kI+VGJ0Hl/PuxSd4CiiN4GpmDwUpLuqNKJvbXDMLToDzunv9AOAD4QZE/LgdFAVOaBv5N
LlJHq6ftvZj1iarAAwNo2m7meVvdsxfVTtxgYolRg4ZSZmT4z4UrF8YKkgdJhY7+NypN8m8XOBlc
PfVa535qMuMgEJupFni2f6OM8asWKp6CQXXmld291530cy/a2kCf88qX9j97ILdq1VcDLL2GffCK
Y+CKGBG+cMYjl4PsHc6Zreg3ECyk5igfVencX3CDemSsBEVhveuvnbYKH9xnDrCCj/0vd3HdXYO9
Z3IJ1mapI121pghp1pjx5vlXT7fo8VntWLLPw444bMff+XwY1X0+4K7S2tOJG7wlWxnNS7nWbXNm
+KB5pMw0Pph37g3kyf30RIpt5nZ9lAGD2Iq76S9Sad0FpWBk8RAha8JMLpll1IFf5KYLdXp8FrDe
yw5SMlTJAUI0fdkSuHgMVIQKgZZi7VLwhQcHzL8cXzNFGgWXQCSAWWqY0YyVC+Eo+WBw//j2XDfR
8RpCcHxqtwL+vmdP6l1ojwR/1Bxg5clE44xQvJ5nihC1aZ50Pk5uhAxyi2dAPKl2EwPtPljFkvJX
8B53iALVozfhn8Dgr4nAk24I2amaqhq1/KZGFre3aryLUkbw+dW9Rg6wRc+tMv9gN1m0kl6H0stj
TqGi9qzeKUKST+gMohP5abEzusw0CJMEc2M/TgjKGUEZbF4NjnHbimtvLscl29zghcZEpMMj4P5a
qevWCQo6zOLAAywB/ZAkhLHJZ/gfyCvQcz8dAx/dzKEOVJeRwnIvMgICw8F18o0CdmeE8ZsaLsY6
Lm7z0CQpZYAEepWvtoU48RsPwxhYvC3rx3LbxMTqkw+t5c0Yzr84qa5JwTA8DjBRdD+C3QPnc+PT
Ydyeq5CNyBJI9rKZ97ojoIzKWWucx3XcREFUIRCCYInutuJiL6EhZYGbPYqlYpfc2u1A2xZuLt9D
uLAziuBf/sGa5nVg768bvu69tSihSmuQuMIS23gk/3rILCaBgCs41C53gCJC6xW0WscD7qWejWGn
aROJcaEno3GLOBanvwj3DmiTmN3ppGDepB1+cCygh1VXdyRXm/6jxNQNny2CmXnmHfqAAWKlogBF
C0cnixyqUgZaJcUOd7ZJMudux9FTKHHINWo3Yb2Fokyt8mp34xS1uMK9kMl7XnskLvO1N9RUPOE9
ByBOxvec/4URhV2umctqbaMP5BAiy0eE96CnkmVL3bhqCzbdDm/rg389XPZE4Fl/ffYa0KumGnBV
U0aMPS1KcL0b6a8Lj39RXD7G46KEIyeNyqg6qX8VTHz0LQv9HKvOk8HgojatBtkqieiZQIDE8sQ/
ThXjS/u55eSI1vwtkMTUsMe9Q0m8d5M1HzcYGAg9YZ466CT8qCXGPcjHnqQBiXFP3eTBbtwuWbcj
7QCpSgPTw2qVf3gllaGGwwdP/HO7E1X7AsjNThkVoibhuBaY0zOg17gtSCYOBPixxlWYKfXOGf0+
rK7fZiwHi/TjWSx7CinzIGAP1vMzT23YtGNJQwsMGqYFinfIyyxVDPXRnw6qw8v1vEW1pz3miiUf
kUv6GTqkYbIVmjQiMS4mS3N8BcqrQtY9sHlJuXVGFli02tok45unvMbeDZxlJ4lTeXdhQr7cHex4
gkCFAhp/Jnw+fnA9McPqZri/9r2GiIKERamXJQGQh3Z31CnfeTZm3lctpuap/vKs2PauNDsp3ZPt
3YW60ppMT9aVMus3q6fdixWxcqxBRrRb/T7+Bk+7LhCyVAc2BLcVAmW7PslOr5hFLFklLp2LRCrg
2cBJK+79RWs7JzxncQxzSJzKYB9CocDiT0Aay1ZOXc4JVLYi3DDDTnwLT1ZBpWkDK+rurFvxZ7ji
9EQlkq9wT2PT1XYigeFtj+K1/vNVrPSMiBuO4KbLEM9U5Q1/xX5OTX0bfs/H3aOZnOmR4EfiQeuO
KjCSmPnp0Ni7PLoAmEzlkYsuXKOcvI1KPbEJ/DOecotsFDo7ptHuL3Q4zQ5n6SblOuMECJPW7Rgb
W8nO1xk+VDVDjNpISjuQ0YRkPJ7f6mLuq/pOnj2X79e5bOrWL1k1Yj4bICw8wWuacch2DwST1Wbi
V/hzqub6ZRjYVtSnQ4g/UDYM8joxJPZvcRgAi5Cs/q+UlyhiHmNGD7h3Eunhay4mesRVJLuum1Hu
oOuq+D8NoJVbBNyANR507Z7IsBcRXy1ulaFQ09e9LuHtZWtaVPN3fOHOXlNRCrI3uH5KDQdriGYR
zjEhW4xd2QtL3qmtMQammPwKYJ2qT9q9j//7+Oean1dHzMDbuuEYecub2lKLDHjiqo108lv51VtD
lpyRpwdZXmNG5sKDevYsw9/vqd1D56TIekqxBZyI3GLNwnmu1AwSPpfGAKquTN42jWeHd/ukuV66
gj36KIvpitmhNVryFbZHKS3jCjHeIsrHxd4YgPgT+Jvnduep+vQt9z/+IXAIzlpKxol7SSonC85V
MLxt/jdqmGc4RA3SkEDmu9aIg9HzkwrgEI/hJmjl0IJm0mjl0qrDZC22gfFgTrVG/L7xMdCszdNj
n5hBb4DNwjPYqUidY7+hvlDVG1x2dbyopdndTmDvakLzYctDfq/CYJDHRW/qbxzc7TYq8ooXzQvB
5AlsJmI+lQJJnoTiotnL0FBjilXwqv2KkP9uuzLXhGQXaXZhAHpLI0Kpnv/AGmBVesvfqDb32LoW
mfs2rwOEI3ODBa9Pz3ydSAhn+VdWAlK7SpycHVhywLB9sx6xEtzVlusWJv7DLm+y9Ptr/UobDyXL
bQ3rPMCZu6fGmu9MoWc93wXpNG7/SIIvmwenBHDrSwY0WlxdZqAek/xVEzTSGTDUJ3nDkitPr+8c
iFMC/xkvOmRpPvn839kjEfiX9ykbhz/8S2KXqVCecHo2q0yR+7EJY9Du8KtNDsr2uBNVxccmk7co
x2NH8aJPIAot8wFo+aCwcemn695cRl76fQt7VJkI3PyA8b1tXYYKwx1qwc+EXnK5rK8wzxVAh06o
t6tH0f7DYixiP4G3ntKa2tpHCyTLwKwpIpuuDNwwx0ipwWK80xXMnnIhx/EUuqRBsLvYNshtJBZj
DpNVvVXRNjYPy7oo/vPlq8jsX+d4/YK/4XFVAjpPFyHkQOQcQGRusOTJKX0CXGRGd+Q7mbEKs5pT
a6Koichvsfmx+tsv9kRU0IpKtgiKYc1MSNe5zbVWzeXyv/uCqw3RJNMEZ6q3C6JOqM7mO2qOmlIW
thFcfnSIpXkLSF0SD4MxmeYnoT+ckd6XE/jRhmPVZpPPyw0Ps3DEf7EyZlk6RhyfgcKBY+9T84yt
g7TXHABC0hlD6XnuSpFZ6nVDWBwBk1ues9plFGguLuK8eYqpmXXrPg65nTltqMwE9RZWO7MArQv6
jT0Lq3eGXSgvCNK/0lN0g/G0GYPZht/vKXR7Iil5SSS0dnvb0jwfUzrdizDR8yzMe2mq3/7yUXio
Uf5DhDiWxxLT3tFg4qWzTHdud4EyD1i7uSVIP7sw6kJZQO7B8fTmI6ojSU+Gm+TUtLmrLQWSn4EH
rfCnVpW7jCbkVFsDeiFswN9rfRfLTMAEWgnuWpYiM0e4C4+3HE8b4KOlQuGDRFfrtqB386r49YMo
0qNPn6eedF+oVZMHQp+BQD7gd9SuCfJfSJRkZsAYVwEJMnmMX7JM+FhbnMAObI6HsDjiGafATJb5
tKiCM0TJRflDvFSzbMVzgZ5oWl8PjU644UXg5/zxpNsrc0Cabchcn3zhcIX7edc8Jv4EViJiRY/+
Gifsth0OkqFWgXdvLkgkQqnvEBEyPoMA4VkMUxhWtLej7l2gkzwPt5CP7F3x/45zmecxFWb4j3i0
lqNTRwgbgWR+/i+r9gbMVx0iko2YVdEHHPswMDU5rp2fj0pXhTwI3jC3LOB7izlK+4q9EFtGVdfN
XLEDJrC6p5Cad+my4TW3Y3qjmJf5KGPaUhJDF9bcchD4FeyWrNr55iAaJuqsSVyRmi8JYdc3nDn3
ONLFPQIPstx2MfYnN7hwCqYE/1HKImyBBXfQ+0dK9iRAk/+gRbndJFjLdiK3LgUjMkQt+INWY9Br
sku8Zm9WftxGd0saFDY29CqOd8gDTI995ycXoLTLjdO0IbCcERmg68swcgMN+VMj52lKz1h1rkfu
ewLe6YRPgMFvX6u+BU+407mNyCDDBDvpvHsfkf8zdmBSmzpLIHPRzqXhKnnUb/r/VDopXKXHZehd
suZdaoPhphIkpKq8jRg411DrywfUf9E95S45wjn7NCJ/57CwLCU94pWqWzU5o+46aqeZrTF9FzHp
/u446vyhBLioZa9QnCD31nL3H0MB7GVBMXucCX4fk3XumxeTfeM+drTdFnwbAFjUKhAmb3PhANI+
88J9solQ3A2BMPovgkGLuzUle7ww0nhR4PfcBn1XyhyjyGEvpv4SFh2+0oFTBp1+03MKRLqISDnD
dhsu+ytADE6xKnJWk4v6swv/td1vY+mEZAGoOrSG+N5JMgyOSPGLCJaQ/9486ygbjg9n5DXHBRhs
9ShRZd1QjP/I9mUDw0pVAovOxxVYig2zM2OIaRrzOhjTHQp7wd4TxiWgGU+WObhTfUw1cRvPurzp
yD28GbI05VYrAJa7J4O/JbKkRb3ZkTjmpH2WFBsSFlJ9BTpXyoDmrle+5LMey6AAexvQYNEZV2uk
ac8wMtACtUoEXdC7AE4K4kIrzodKtdhPgAjtPYi3MN3EuNSr2Jn3bPIqIPpWgTlevv6OW6u9WUS7
UH2ma4kihSH7o77GUkb9KgcCTE1gKV1hewi6PG4q265/fibRvi0WneAG6qnyWPF6D5OI2U+nu5iw
CO25LgAoQOFF4plATDbuExMn58SswEmSDOu9mDbhyc5vqvk5sNMMM8cdBGYM53DhnHgNwd1Y32pv
F5e+xqGS9ifXsN9YqwYWzaCknPvC+jJhizKNV36kvnymvf+gnRf3OHo6LBnya1e0i9MS0f+4KYIP
2Draim7N1Nc4m8Bbb14kVtd9ghVljz6+XB4T/OYXE09eUIaH+LNhlxzMCzwQDdV8UOh0OceOQhuV
1IO4RAjWDHwtiSdEZulcH1lpSApmC4Z/GTt9W+jAptfgWtFPzK49xp/SEWwUCPRV0qS6b3WwHZFB
UyFghAjIbHIagdI8uwovdOX14RFHuOpXck0H95z5uPVf7xD3UIrXZkfuCyWpSWVq4tTriLTgx3w7
3apgbCPTEQbXA4mF/GFfFqWKTYMVIPHdGa9tW82WX+UFYjeAbgVSCrBTSb4S2dMfIvrjqWsu/Nxg
7PmOKz1o3zmz73BfmHciPaAY4JFllM8msiS7/HU30bmWFtShKycAwS9cw3KLZTxhlv12MiWXjFle
Ro0bs2Fl7zAgSUfUovLk8cWM2ejFi22vxSvMPTeiNwOfYZU5H3UVZWBdyUiISrIxHQwCUah3ShYK
Jekd5XeSC0y2GJwDjvgNjnywfRqY6JYLE/c3iIMOwsEXe5VohjsrlJC93pSl/L6D7sCeK3r4zJ5m
vBcNrRNR5KoCW/Kq2RBAq10KZ2MkVsIM2jbiA4FQw/1OBd4ZpWUp0P8K9hPX9z60meFXU2180iSk
q1Sq4ODwcXe0KdQDxcCtaUrQFFgDRz9/z8lN6FEUkCsB5nDKVhXFK1O8movy1HbkBYH/RrQhfTjq
6lQN3JeY8APpn7dttKkptfR5UV4WjoTMDDyL5xJ45AT3JXzY0oHGfIz89fz2UbuC7aLVscSkamz8
HdSmKWqsIl4V9ueS/PMVAxZmKMJI5zgAs4L/ElDuPoiqSHIPaByoGJlFEUqkvYN87+vqqFdbSUun
rKqUbkiT80Nn8v9z+EzNFOeK3gqwPpcOTeD7K0dxbHiB0FxC/gFX4Q4lcw+h0FYdyteNgrbSmLQp
j9D0N4eFn6fCWLgKYXeuVcivne9qU51mFW4JTqh5IYO2ot00wteqzri47Db75T6OfzSPRkaipD/H
DgLV2YpXIqwnZtNBL3A1hK6xHm2a140f0lVMxmBLm8Sdh59YKF7hFZSBWIRbK1LUJqXvI/PisXpo
qcKcXAUj8TE3FTZA9WO4fzQgAM2WfppqYd7t/IX7giTdpkhUV+3I5oqVq2fVwhx3w/uQAl3Cg61w
E4bK1LNbXOnvIfSgu3iKFIkDX4Ktaac4o4k+ipVGZFSKBSB+bHmyqm8sgyf8vX7dTJ7Q8pK7psMq
NRO5VYJ0mmdOoF+W+tCoQdzyULK0Sqj8SL7FTYJ+31CHcx0pqt6nlkFVTPO+ci72ZEclbuUkSha0
gRnT9JDpjvi0aWZpj1dSkrE7SUXitzvhvMIOwhxub0d5exp1OUgypKiqnkpwJfXHYhnuwC4+oywR
uQ657s/GqkkI0pyOIvIHBloFj2nFV7fvO6cYBimeCwmZ/Xv6IvKPviZSjRGfwMrH1NQma77zqC/6
DKpkg+JpNyjTgyoXo2Mb0cfXpKpNEuZFQUzgBCh7F86S5oeP8JaKA5ym+WsjWZEikHH/iqXYRUZU
1haSCukOzBRA7CRpaCx4KA9KTwpgMMrWZhjRRjkLhZxVAh6fR0cnsIRfWn1y+XhqSYycgeo9zClp
6ex7eW46aDo66XUPb9fHJyOxXvUKRhlJ+tJGpPINZOTQu7f8xZECTHyFdErdGmGoPnaAHlKzz1nx
XVz28KmCumlFmCd8BaQhz79bS8Hc9ar2EyPn4If+y7BoNi9v37B+NyNY3GiZArM9z9Hevc4KNrSb
Wb1KmqpQJxAyOaCKhb9zGxOMng9BLJhO+jwpNkiyF9XOxf8+TB8ynxvJh+zUOwgxMwerg1Eba6TC
BUs7+tZVD1rEzGoG7OcqW9f8vzhOaqP9b6sxuPtgrbXmsa4yhyL+rPJHo3YHDCs4u0VD87lzGbFS
7IMWJXMIBhUCQmUkwie/v7dYsHr7U7IIOxMHV9QMpzfSDtimAGKlaC5t3vAq5bi2P/PwStJbyC4S
ROLZ96O/mlSi1BeypLT3RXzdxzGORXMmmKc9LsbY3rGBK/59NGuOm+sqmPUe/99ULRS5sk9t35o3
r04A14wXqyCGaGnvweEUtoTP8QngcA4vGmQ2u69ABMkKR0uzvn0wqxPVuv5y7ojZjcJAAFTdgFPw
NJz56myw1gp4KDWwaq1VYedqVy+nxJaVGxFrFwDefg6IA4l81EJSslfeHKiRRhqvWTevJAG3WW8G
bniMcH4xbsSIG6LMVoT0rhQ2lez/z6nx0m0xiwM/DD5ylywmaVez+qbYnsSrn3TQ5kFTVILxKw2w
sGBMswxvTbw3lv4wNf7GDcAIqfmX5dl97P+Pgsz3eig0Ps2gWpMsv95m3bKLd0hPowHgtdEESVJF
uZaZ9VAmsTa2uerqopc4yg6g3MknN/QZIzq56YShrakbTeica0qmeVVK+SYv9KBunsJ+lYHVQJMv
iDsQMXTWTXojy55n9851XqAuoLunRbPOstalpPLiolWWW1hQvUB0/w2GznSbYFlwueA6cjYV2mcm
lRqZSipZdHVnjw+FpAxeZwDT7hegoZrlwN9kINx5b8pmAo0J8KrYVIavvJnrZ9cYR7NB0d2kgZNI
gl56osWSRUDXeAI/DMNot1pXZy9aEV+TH7AvALjCjxUhhtO7YRmNAbppiZYXoCw3+eJqw9B8imc3
XsCaR0WOdu9gRoAYCNAsgIdahnQmQTW/rPHHrVIsbPLzAnu9P38iPP2wlFq10RmLspKEIZZmYWYd
kt/4iW+XBqqk/DVEdjzexC0/UF9WpfbVe4KYNe/jz9lza0UhvvyYNbWySVYJOfsgyaFpeg/2KL3L
tdsmvbSdrwm4dBTdUy7Pe6O7s1e9crwaKchcvRYjPVL/QKUYRZ+A9ozPO7/Bx8W6/US3apZoc2XE
jqG9Yb8QLJcJFTwsGyuZXSyBqCC0Z7y+wnpvMbz/FsELRXDdMlXoIp1qKN3wjwZOCAvrvcMKH7PJ
44lfywfIFMNPqk953VNV/WZHshNbYVZwwAfD+ofo+K06+F6SDRzz6hK+QW+v90UBbBQgI6VU9/KD
aInTuWw92NFFFWX1/IfO0Pm4aTPGhtLs0ZzOjvWl9+Pqbkr3QpC9VwC7z4jWjV4OZq/cLzpNBvn9
2MSInTXvg9Fjj5QtSdJLeNwBFKS4wChMGvwrMJ+36IbxnbFEHdd+h0vqSlGI19rgLAbP3sYX+Pi1
4P94HiYnrrpg2QQj93MXwD+vWg9meCWf5uQr1ExaKomKgsgwkeHrCe00AQIb48J/S22Pcvph8VH0
5dNjnc008ipx2H+OhOU563H67JxX1ib9CMAjPd3x7xM9N//jBE2+2kFZz3G/U8yTZ8W5Lf7NTIpu
oT/dUaTaX1czCHOewfZbSQ9ZEm5u9IWPxo4mpXs3A5uhReRMWvZU8gPyYtGM0VUW9lQspUSaCNJJ
kPUwuE5N3kgKgH206OSQMspX3uIvT5cIjoDIE5RQQfalAnoM7U+CuPFTofxVqZCQi6guy9DTXmC+
/eHWstcwbpfMIlpyDacJT9fC9jYRIz2qVhXslGyZiGMoMrnv1NS+wA2GSaAWOZjcN5RsWxg3J6JF
EunwFlTk9M+v5JsgMPxF7X07QXdly7+HHnS4ccgGwhxV5TYqrkXT8jeGBw59ursYty1X42Zt/UYt
mBOxBhYsQmzAeQg2QVDbQoaClDMeol8wua4DuWClGEIbzpLDBF5/f7DneFQ/RzatkVn9YX8/wafy
4GXJBFCHV+QTssRujPeLM+DSLKMGJtWRNP3ZIa9NnxC1bsyG2mBiJg+vY1TeaBE6/GrvjOdLW/KB
3wdMuZDMicjHP4NvV3MeI0xGm7F+kUrHyxj+ClUnw4R7EUM0OWJExCoFYi96YpQkIp7YCihNFqeW
APCi7QCe9e3lE3y5vbG+XWZu+kLhUj94+a8HcbFOLpqBDW39gv8fwDsESEJCqgYZjtECWeCcGABX
YaOzAcOiCJDZKxDAvygAONqAJ5KQc0HDAVpMFeFwvk1mtz6jg0Ymjf4s1g4dfFJ152tRWFgZ2Ffb
zKbPslGU6LBkizQWTvQd0r4FpOfkyeaPOFEd/+09KQW6neHb+raPZHXDPzpsO0yXUGI26w46qKVv
ZuoOjmzkJPIpHAhs9e0XjATzfqhjlnbt/GmrBJJJ8z0f0sgzYe4js16PnG1W1Pq9dHqXBx6aqXVH
HFsdjkCqT9m0DO91hGV9REzs5tDVsikRqjzqX5+9PrnLFLJRoEGLy8lizXtRZQYXcibIZAsq+JMT
Jw36MyuDNdOcUsNefWHilqKcn41YbU0obKFFUwk3cNABstu4jVAfpu9KIwwk1yrhKpZEZ5suFaW8
HVkGzMxuWmgYZH0RKWX7P9BwvoP2i63TiIQQARhEZLEC5TDOKNWRqrh25/F36fedKJPnN/hYM8xP
5DJCBPjpCnuDjs6sSIEoc3GilVN3dHNnO80V2aGfWDQJuMy2qsPn7q0uqBFMd9gAW3L53IsRLj6j
2i+e7URtGfLlMN4viVbma56ERvFuwzsQrKVopCLg4kazwxNDKhAKqhwlIX1pUI2DClAPsOa3cBoo
IGx4sPgawLM6m7xs1I4czJzRVBQdJvg4xLNxI5xc81JsmJVZe+S7W11NBwk6VZAQVt8hF0K68q3Z
STZ8ZZfeqBb14IkFlnbMWH2WJ65uFPuyzP8oN7Psz9xwM8PyOZ3FDeuMFI/e0JGcHRqQWLii4pLo
VRS2T00UedXvNtfx80uehb5APnyFuU9X8fEPKlWCV61Wpb2wTVCu39SndV9dQEFGqrm4FyQ9Q0Oh
ATU92HszJ+AUWc1DLPU3LbwhltC2P5YxEaT487NlEelomN7gyjJJ0rj+cBGLe7nn+NaeF134nc+9
N2Vh24hQs8De5w0RWIka9gXMDrxpJ5X+iAvpvbwsd6Qu4el2eAeHOqED1/vVnGCuI6CavIqiKGKR
vdMSPtlrqnbXc6i2F0Hg00xNJgAramzzQdwA9h/i6B1fvCPZ97xvf4rFjhfoTvyyny96Ma8rzPkn
As+flAbQpe2tXiwNAGriwUBzDGwYt5BM/appBOpXZve+0JKxnRwImXYnPiAAtYmt8XiAvFWTuabC
PHc9XBdPi3hJP2r3m7KzxhtFHwmIXISakELlVQXUdWV6JBFAOX27XYXd/QJFpvBP9d/lmhyVOWtv
99r0av8UAKFzIBlNwhf6J49VIlNSDyNL5Ii0vJPDqPGtqOmbIsI8I7nv+lPSbF8yig8Etbj/GWEb
bZUR9iL7fB/plDAuMibb04e6FjHpYFjjsfFesBExbhIKWIvKHWylhsyIp5sLroCSBmSeEGp8hyn7
v2T/dplwRIfwB6lVtLbnbVWRbKIFlfbnIhETYfXTvfb7wwN5XCFtt9n4/9Mm62+0IsBMMPKhAlCR
9fj1JpnEHv8GOOyYdQm7rvMBDx/9YnCNDPHcLNZB/YqS/fU5qyVPEVY2aagv0dro16kpIQuI9oBh
6fKhXYzu1u2kcJODtFUi1nXvsqA2CE40sFb9rAhIlJ5weNXG3aIdC8xSkq5cMAlyU+JSfEfs/fpC
bXAAhYpp7hLdKJpNQkS+zfISBRI4V3+eJz2sl18yCuy/x8j8fxoXp15v4MYXIRKEItKOfG70ml/z
3wDKk+L6M14kAK1Zai0tlJ7hKFYsJwZpiqPIniJ+NSyOXw603/4DNNj69MpLoOK7+5sDKio6Xnyg
8t/Ntj8M1qvYUuO5vS/NVqor+ARJVIBkD+vmOS/obYIrk8NW8TFvABUhCwiJ3rTorrDQethcILit
G1UgYUlcrXaaK/JTlcyQX7F7RulxUgV1azGGxU3tqsNSG1ZAiCTaChsrSPNScC77bDrE+B7E2axP
1b9AoT5kn/uTl43BjTdFy2jupLKwS6s1W1eiAws5bNwfvMI1+Vwy69BG1tTsgBezhQNUzfkmBs2z
dr/90N6jJNonPG1jnYz+P5SKUZCTt2BM2YeCAreZowtsdf1gh5avTUvxXEweM6/i2ES7oSSTM+nL
sjjFpg3bOuFzVZUOA+/WC47wZ2H3G2xBHEIKR8rhaqLJv8CVCgx1Qk1nyvvKFsDJJQr7Bf6XNQY8
QFvrbxzpWoWiI3l+A+TezxW3PmQUlXI+/BVDaxWumCDUCNAqKsJNj9YuHBC/zvZZsOawqTyHV2by
UZRR98CGpxV9aiwiqidZ3MY6HJvr5wthPyAVB8gBvVJMMq5U9+X0AvhPmi/oAiP0rmdLtHMWViCC
6sqv+JqBsF96DrtZA0k5PtZs/UjFGrFKQpzs0QO3SKrG3jmajvGCUawgRdnARanZQOLEdrSIPOxG
CNEcfXQQQDicuBeo3gY+hcH+rseIHtDaPlDCfmcvww1kb+afVQimqI7P4R6BQqa4iWx5pgUEr9sW
nWJfCVmWgON2rwj3hypk4ZT99nhqa0Ea2FsJHgUJE0d9T2hCcGRUxCR6rExnOJjyY6XbyIpobp+r
63gXX4gROAmjr+gpWoyXjJaLI4gYdt97NLuLAn1eyy1aGaXJGo2cq8nOXBreb369Bnbg+s278Qcy
9/2YGLHEbPzIB6JJNISf9L9+QgMBAmbMc50OqxSMAUDtwfhiyQgdD5LZWSDDyQMQcobP6NGfOxUz
jy5IZRQGz3oHSuHSffI9DKMVd7hO6wOa+NPQDrWAeGypXWRpc8Cm1rB+tOQZ0tt86d4zsWW+0gOX
DMYpVPGrltr77SebxPt8drZd99KN4a++AkS1LmbJYr8QHxHZdWiJsXXm5Q+Ywan9euhbXClZnYA0
xAEuKZXmsRyCGf45SyhEFMVarGVpTFnYxcuMSYNkTfqD0SKlGXyPr+phdcbc2/w2HuL/BJPKbSg8
CFQW9v2wC6LpWAlOXfbhWlDYHCQ9SRLpiKHs8AhvMHnRQivwCMF1sb97H9Ki+Q3DOzmUabOvLB6g
dNGqqg+rFffvqhOWjCFWgKDX4szeF1WWZiTXAZ5muieoNTDDF1lY30lEk1KeGb1UZ83rXEv9UXXd
s30DGS0Fh6LWUa2fCkPlpBfHMHJmA6WnqWQteE9mjUvIAHRBDu1+WToUeo/6M9g34tn7juwAXl1I
9pt3VKSu2Xi9Wpty1C4rEEEgLcpvXjfFhLOusTlgZ7oltXl75+QDDMODoiqjVwDlLj+UOQ3iWGhr
WfWwiM7QD1CejKvZ7gwBFwLKjiL3qD3O+uCJ0WOfEHwYQdCvjytWbs1RzmFLWiZfbbHQgTOF38+G
gGDzzsbp6ivJ6SZsGxuA+hHOw410+lxVBG504Tjsuu2aRig//Lci/UvJWDpReVTZPjP6wguRB8dS
bE8YI0xvYz8Wo9uCr91ffWXh69v3CLFgzSAMbNa9231RXy459S6XgSxDwnDfsHpbk00YVWxS+JVF
FjgLGdH9Q4+37kfkcCa9HI/ut8JSvtBXwnEgL247Fygr/T/SyFJ0FyYT7KEfaT48uKeKME8PHQ40
z3Lv9aRxu3oW0JJD2uj0RNFgEJ4XB/4rg2EcbkdOB21i6Gt7M1qTsQzgVhc0NNn5ApwSmH/jw7M5
qMGRXXh+cIFEYcTzuhx1JagStOibG9dT3ak327ucU6noOFzahwuueTrCifipOSytpyJxah31+cY8
o3qd1bdkp1k1GVGPibBvMhYgsTWJDNX8OW/S9n0I1CTe9CSNNzOMl7dhg1V2U9BCiruTN22zVqEQ
K/jWcRsJT9X8YF4dXGCVi3cT6E1lOwJ+d8H7KtnIZpPHOWyksqrrAqdvBOiYRWHCqCLdpVaVjblU
LsBUAjUHIXsWu3bYJ8Ga7fWXbvxg/lfu6Rwxxapm8FHo+KtPFZ8OwUiucqj9/hgwgX/22vAs0qPq
+N9ttpI+qCZr3G8MIIADJA0PWF4p21dacn7InAh2xgd644x3uENk/7WpofwEtrp0kOz0SigvMJdp
up1nRYwk3PJYAdTMsyA1x4vHvA9qv0DUMr3PEaNOxMvG5+d0jCgXyF2JfOH3bWu4X6pOsXAn9LON
yokkkdka1BxmgTKi22QCfGMvbUXVvbsmnamx1GiXNOYswDXHCWVBEQ+Q6pG+zg5OSvPEEn/hkc3+
/zbkRY60vVZ7Rawm4GAwX5RIml2keXkXad8kG6Foat2eG/AHdTuKg42E4N3JUSwHnhUVLiDVDx5N
G8NQKPZcY5RuhY/9QnM1/BvQ72/kUApUngwEH69aISFrKxhmb9i3SIJMogLw3hicgzGs0DwG8HRh
aSuVzzbf8BFY/KQKKmZZlyRtY86izQPy08IYwQHw5f3tp9oP9Gs0rdHXWqpzmdjaxGiT+b8ytInH
PxSg+c/mfXbV2z/BzePtdKVrL5MzMz/XXSjsDtlvJcSoZhJp5CC4pHtbyVVDzsWA6901rzlmzsid
cB2qxcx8vOhCx6oaQZQMPu8IsfPxqKTfZDfHmjoIx+YlyOIkt6lelJ6mHtmBmZ53vXYqbpFUVQCL
M3prXQAXzjIHleKLYo3zloLnU08uVJJVHZ/cfYB0G2v7JBjBo6PKhB0I9mKOUkpiltkr5vC2oWWh
iZJ08AJgwts4fgtbMTGtss2naxviwToQKm3MGMKBo796qSIthndwTaXOcB5JzAfw9H/kR48Hqd0m
Vdx6PYwuQ9aCcKgAU8YCU3DhD/bYS3iqNBzEReEm3vX8+hXcy4Mb1M5wYij3Uj0TpecBUvGAario
N+7sIdRGxy/DRdadKuVQOx6kbaorPl3vDawqxXDDT8bGmL9OhocD1x8J9r3v8xUDwzuV9PY4X5vN
zysNUo9jxCJ82hXk0dMW4s9psoraUooiLPMpnc6AdavajOHv2pbfA1jTW5zP2k5/4+nMUZ2KOkXP
2DuBaZuPK4mid9ZwodQFsBaNTS7kC0X8y16Hpmt9MtgvvDPo8KkwZuxVmvm7kOE5/qsgNU1cjmF+
Vu6f/XpU3MJn+gU2amTsEVBr9FL7DxFOPWLz3eoqVuqwhaBpBv2aqKm9FqzzfsdSmLxJ/4sF3wsw
5LG8sr2j9upYWVbeSp4hTn+krk6rtE2oeJQsuc3NtyvKXA5NveLVfHFCwBRc8q292FDjgqSyl1sg
johQ3J5XCuJlAbE6GOkI2MVcoh4oGuagR0nPbYypNGE5RPAP2oAyPBuEEqjk70n0VSod/n9euKfa
DXXGYaNsBZPXGiiwbNZPJP6YiwRNkfTB+iRpwzznAEXnCp/ZbkfjV45uJVHKiXEhp0aM4Bvb7LKw
zecwZmFcX0iyy+mZwVq3UA3WN+TyvDnjLLFIORISrMHAm6dtmeVgExjxwAv18t674+dchEuzQ/Vn
T4TmmdutycqSi4y+JysjVU2QjnOrc40ahDIIxfcZ3Z4a3EUw0rDJmgKhSNso9mSdE0n/hFuvpYt2
D4eVJGi5CfzG0DQ7BY/gcDBXevayTyBIr1MJHmmIu0nn86xt7mBbUzlQA1u6UEXXdTrnnWMCoJ9q
zveitT07gkU6xT/eZfuW8fmcyL0bj9+rbV/f/bH29nVo61DeRSRgzwSLszjNYd1ltEKCvgykPdx7
blB1/kXybw5JMOFtLDzYqLNdQDNrdWKwEzovVAJaw+2cObmmVhPbvzg2tyJaK2ebhV99engAMHsP
BHq62e5w3d/qXzOruR0+YT2JE2HYsz2N4U7d2EUPjo0Osej1JcUj02cQtjWbaTl4QrWPYSCZMfBs
cB5R+rB2cJqOi1o0/crpNySyvqCztJ2ws//mp8YP3SgLK6ZkWQ4f2YaeIOLxDytblp0g+nBbFyWc
oFmxAvgZIsh+iFeUB23dtVEdzq9qMm/0eFnXRXV19MBVcDtGlf9UTARW5Rwb2msJT3oIoCs3OJ1+
QOLSySayYnh6DdVr6j1U71ffS+vJZCexgisMxj/i4G4EweT4S6Zdl4xJ1i6jQisfXw4XvmOGu1Bu
hocLzLNsKviXjtbi1ElSoSrZZnv5RqfU54OzB4h3DoULcOGm9wDERXhMgT95zP6brq4Eb5xEjMLN
l6b8L3G5snivxZXS5ndv7t4aqZDoXpkDbFzNxWg6BVKtalthbqztwnW1v5bgua3EKFjbuoq1+7Ig
NqNDK1pxW1NQ3M7buO38gOMf+egLLDuFelLW2E4LQRxdPM1Ds9+WyD3QXk2OzN3wLBzZSmIHPhYS
Ttqh8r0lAapJt9Q1ehjJb0kLDJpFwP2nr36EA+p4Ooyvd5For/xrXXG3SXArXXC4czwFLJOHyt+p
q5AlUWueoSScA9ApHHP03KiMcYGY2hcC5T1FsqG6kEGM3e2gNW/bglxd8CD3+d5xai5jEvuqPwdT
PhJFg5wYC7h8lVS5UqElBMIuGnKBbDXYM16gC05GcVaMlP5yKqhYOEQDkclfS6Lkj6FOR0U4jLf6
IrEBpwZyoW/u8y6lpe1l1cmqYc9/WdLlzRjCgz6uo947sulFgA2FjilO7BUsdLvttfccxwpX2gbo
kL8VEOIxJCR4jFtVgiE8U99bPybjQV+Uf+mNL6QRxdTVu+aeFhnFeRlGBJmH93exjb+fwQ4P8ZbH
WBHcjQUsVQWc3wyU0xUyxAlObQI1jL4rwHrw6F5SrD6ESygBdyHt7i0nR9KNK/B60pUNP68qLvkB
3qNUVBOnj06CDJGfV4BHCJlzXU7MhdUtzqduOdkf4WPo2hBKc7qdVeeru+7YDWjN4VGxjudsFrtW
ykkOmKiD+qdTgoPNWNPMsoxbOPAtncSsVtbvY73HgKUYsG9YfJoxt470xC+mkz9AsDnctSGPaQyR
ygeLLTFhLRLhg0IHNyWKC2SokF0lxf/9Ta7mVNbroELhwT4ZhUbYIeAQ9GE4Tk9Ah/J0e+TQ3TWJ
ZqtPPJkknYhp7Hbir/x8dC5D6Zuq+N+sRAWmk8lIBj9FQ3BPkFMdErC6Vxwz5/TC0xfyCTL5rqCE
BSIqxtHzVD2XK4QqhUTgZl7W2Qag53qq+CYYip0XpXPka8kfB19djxuaukwA6mIwkJquNtLgOw1u
QRGBThpv2fgAxGurCFB/h4NsdY5UZZcXzB6eukK4+LoitOQaY27Lj0Isrsu+Zwi8FUGhxVvnZV7e
fPF+zqYlP7VRZa/sJ/XRQQ2PpOxSRCaWjyD5h02g6POZbkMCuT6e5nRowfSy58eGsaSHZIEMgqXy
z9vRyP7ZzjYj4JqVv7xJS81N7XkSL4Cn5JM2ZuxGBa6KJ0lum+cdimp+ojaX4L6/FQVg5TkzIx1K
SUSdGNGIHWqqRpx5pnQ2v9ryQPla/GA408TyIf7QeYltUf+e5NO13qYhxnnvLVAth0zPSINjrGaX
pygnQ/BXUqf2kr0RhkqGRHKylv7z73QWNu5daVUEsztXQ8a53KSJZEafRyTgERQq4tj5tIqFeHZ/
9eOqYGqb6IAySccznziMnJdoh2rDQ1TAup6nHewTq2TLH5npPqXnNgx4F9mtYNrxMwK99PmFi2h7
8mo54HNpkldSb9YyOau1I17uDK035GB0aLWm1hUWGv0MLKV6cx1VGtbn7oOBdjWIFaOlVMneCZIO
FEXdEpC08GUPq5SXOElxOYQsGGupMN99gM2QikHHfN15Vr+Tf1JcOwciQq2vgJCAt17YbX+d9d7x
LtChbWn2qn9rfqqC00wEajK6fDwFain8exX2PVEfLylAKjq9sLNmcs9Beyqj6J1WoQM8LzcsCj4u
r9Y40HG0/sx2i5kN3FbnouuPtByjjz04SIkuxxfahcIwbLIryKXevMOQqfaNL4r0IKUjMuMI1kde
dRX5DlTGqGSC2j85TURu6HUJYmuEGnWcGGJnq7ZK0RmptV2cjTX04NdJdNpv36fxlRVHv9NxgMFy
VsvyUtt9jlWlohhrHuLhH29J8zZIYaK4iOzt335WjGe/8pHUm9YQcbLElrxRWfBpEwSdRkOJFCTG
qJK0iNjqIO1S9wK39SMTEMcitJa7hxm999/SgJV/RYciNXbGIgPPQ64zad8VI2H24HowawtMFTsl
+4wD3X2sowYnwTJacTbkTzmUuhFvLBkDcKNk+q3MxluGtx2PR1+DpJKWVVS+bU8wF5EwZ0KNg3L/
QncrLBKYpeS3QO7g+axTZ5OB4VHMDZYIalh0W8LhVifEbuscOEJelC6IdQcHVUNfEez6OpP6gFA7
zSuLkckIlObX6bbQwwwG//YtdZwWSuK3BXBHMXXQuyNVqzj95ib4JOfF1aKJDY7WMkEZakj1A6hU
lYybnwD0h4x+J/GS51QVheg2y2PBBa1bwiKg9jAE6BW2aj+3Xu/G1Gw7t7tE0D5qU4/iU/7MoO0y
dnb47x4fuIgFLFoRPaLmYECIo9oojtTOi6Rzz28Nohh1Autoq5XklAa16YvFJfnD49xf7sotcoPI
qNvtGRd69wZ8R+pE/HmhNYMa/4twTvR0Ghwm4JyW7M54RmCosuwU92Z3syxenqjcHuGBib7mbgf7
jfFjSYbOuHfjhTLx9KDcX4LIS9kpwp/RDxHTL02riDLFXgZFXN8Yw/xtw6kN6nWJTrjbH7wYOh+v
TWMRDhAksv9G4Bdkaqct6J7QcvVxOYUaIYhevCNzSDkk7qeI2QtZArUA8OFltqPqcsmO+gCiwm9W
ZcYOLiQ2SRY/BLkw9fE9dcpM3l4/pE7Zb9zpbAiPwtFu5OCq6WntcuA5IeA3aJcgYujzwiFMdvRF
RcYhd7N1ieRX1MSC1dvBKpJu6lCiTB/+hLSUnbBSN/qgFqMfNhGfBJMDO7nbGyHi2O3tuW3uvXhU
y6ePHXr6ECCgo4c+gr9ZMNAygk8DhEEfLXqQ1VWpJYGlDTYvW1iYEYNWF+kNt2Ss+UrKAxD+Bm3B
tV3fh9XNk3jwFk1A2PHLDu9GE1xTZDXR7uXudDpFvFsbbDY7oD/2ZpLKlmcALkqZybdf9ptaLbdD
Hb8g8DpMi3m3mlGqHWVlZ7Xi4a7szzlwNZsRJU2HejFH+qaUYDnKY6qq0zf5AgsmOGBNqlgMiwIY
6XJVNqQ/nBQONW/SbmQ3um5BU3zjkm+MFsVJCYwIVw8qYPdorQ6MUbdTwv07rQfedl5NJ4Pv7I+V
YT39N45MqB0C8FdQ9dPF//rmonufZ5OB11wnsq9LCfL2lFCu1hI/ph75a8TrqrDgAr6TzMghUjfS
wDN0TvMI6nF6a2Bbn6AEdYzeAU86cifCfZmZe/3tIoQR/N77rmKOoTSsfQeTGgA/twyEy3tgKkS/
wgvr2DDe/+72D86bhARapc4BKx0MbBSrOkJD5DyLlTy6eTa0TtI2JPx8wfNcY95+M4hv3DJf3Imn
uf2cJfzPbErWubCoiv/CcbT7yh35V5hE1q4mXpJYrsmEK0eVwkyH6zOw/KQzqbLYBHbLYOjElURu
8FMkScXgNbw/wdXqOiOpK7HNmty3ayko6AH4RrD4DMk3ZFtPq7f/k8iE89TSoptjd2yNglY2ofXR
vLrGFHJs11f83g7I85qjurmWcNxGCMyrbOalEw2Dofme0/uOtL3wW5ig2llWcFZIgmvdHVvqHyAS
YMA0UUJtHtYU8Y3Tq5gKP8g5tGD0euoBH0pMAyfkRjil31kqOHD4rv5VlC5scpJLVGK1m1b8RvBg
/yfrGyfb4NYlDbQ8EL5HMi00ADvzuv6YEAhxa7sXYJM+zcZgZBL5R8b5smFMFUZWBtiLSoZjDYae
ae+ScxQpteSKfw5frHny3CZrwTnaTkugfw8l6tZ/veJOqByGS+juLKIe7KoStLfEg0GQoNlrqa9z
NPfD946FgX4lkqXxIw5ymleAlp8CjGvyo6tDEy/jNE1IU2aJz8mcpVZTdv9rgn/nfXruT+b9aY/M
MMl0nqaUiXvNHiglsFaO+OKtBD3UzjTT6A/jvz0tPZPubLQO+hGU5b9L7C803i/4FHcV+n9YQSej
c8U6kKr0SGTstCv8hnBAy+WCQu49h3W80xUrQL63xug40nyMVoAy30ScuIf333i1/7m6JYs43CJA
aPZiFoCTHJno0MkPj8PGJt/qFhv9qWkZjiPwzYpc/y5LgwHzXkNVJexD2FCpBhNtU46a4agfkMsP
RDVq5MEdxe/zIHyt/rq4YmcuUx7XBEnzFeoqrAlkucSvthMKRFqAZyVzzShJH2iHSGiyng7J8l1D
fvVdrwThdDz2VoAif+YVGozA7txgocwowLckCgMX/Tx1ph0t1sbt4pUuUEJ0miJwJq/g2SkK4vI2
eCLcL/a0CY3GuobuC/f3Rbur3fReJ+MVHK9SI1WPxTsrrj+pkOCHqLVYd25ALCWZfSzCF3jRjccR
qTMp5AR0vKJ67eFiBlWzgERvWEtrq0qZnbh03+wLxZsrxoyBNedPDo5CVtLgokhMi6hmTuvFQSVN
90L+un893b8XvWw7jlcsGxgWWYVuxCTXuCKav+8UYTT5mdLkGKmMICxOxysO14hYjBpt/43y7LWG
oRN5Kw0cAc0PX4CQzYhL3zRPQ5nwFLxKd2loWOUayfnHkyfLdB7TfWIyApBqzHGypdz+JRwloSXQ
qk31S8MLScG0y7hS+6WQyscxyW9xtSJfSistHch7xgQgG01l2DqbFYa5/Ruufa8RlL7kmEGfVGut
Bk47aYkx+7o1vfJAsgQpNREmjwdxTq/WirQvbcCMUazf71h5XOkzAg9s1yJy2OM1W2Y7x7coFgWU
HXWi8x8W0d23Mg52kGSfwkQ6fZmTWlixVgRRmaSRCzGWccr9zf8cvTXnEVB1h57YCwaRkXjwR8ms
ZTioTlewzZrgMXkZHNZVcuJ/caG7PN8zerKMO1MdrxrUHP9kYTHRqmUkI4g4hdFXDX1zzhcAEXzj
v5th4pD2L0SI+Kt9S1vXoct1UlbrziADHy1nXd2rHK3Nr/vVXUaNZg0qqlVnWyGtlTzzW21CY8q6
x1FnTIepMU55L0Qz7zJz+5Z5QYySLR7vMkR35NVV2pkoIJoqS+3aXFkiR8TXvffo9FN9CbdtZxR7
zDouBw5AD8ledHowgKxH5aguzOrNmJKdB0qdT9Fmzn+eq2xdiC7YCyM+mPanDQ6y2G6Qd0ozzmm1
QImJ7YyZuXaFkozGQGNJRk9Ra6ToTNJhk8L0y+em/CH8o+6IZprGouvzzV/SWv0/DRwGLBiYLdkj
TVIMMxX+uPrqmD9GmcWq/4hFO0vix5YI/zuYe7qT3/gcM7NEXsjKm8YD6Eb5xFj2/KN93jMlVNaB
q3SMely3o1Ma5I7E01tLP5X5Ocq6MCzoeBHz+p3R9slsQCp5eADJD2JAvRiClfFIjRRVQCx2qzpg
yKZt0R/SHmAqT4WpdDfKWYdxYlveMAFplSUNqM7Vkgip3vEll6VjmKpgpzgBXjq0ZNUvNBmEbX+w
lkDcEMGPpoQTP+6pjYSyZJxRUHrAJaV0bjwrABpFfo0MET2KvXm3Z5Dlt4yH4RrXtg8zmBiUysyp
N7cwFECdKLnCjLx12p4vuJIHWuiTI1+BMcNIEdeRGO2uHAM/vNdxmcXVISkSaDAAHD8m2NksbZcz
CpE07XHOYxEXR5TiIP0O11VPYGziwcu2FOJ8cKRmlGlZCwXiKhYhaLD3ZBmIgOVD55sky8sSCEQX
bPgIpMKj13QK+V6l1FSZENqyFh3A5Qkm8kWOAyBamrqyTQVzBhEPI35ZxNuiS++mqK5cMWHykSN2
wW1M/OQWP9pX3K+wKjs4fim9ED/TQQ01yRY4vJ2BKrf6VV4g+/po//jl0nS9DVlKvKP4UW6s4jK7
TlZjXFCBKyeMXT0tgxtVqZ81LDQaGCZCtdq1aJbEzq6n8Gh+Py3GlZEMYuQ6PHAChi8xygCgg5TD
kXglDe7i9fcZap5lzBDrQ9p1DFyt5cO3ebGq91vjY9bjaO9OFolGRR4PCpvGh7NvPKkQf4mVnvPA
OA999TkDt7CndP7XEehN6bsbqKAu+kEvS6zqLEyAaeVc+WhcsoaYbO5f9qc+wmPjSVqpbHejJSOY
m2BXowA4w7CF1cbbGpztOxrwfQGDDxKY8FT8zy7CirYHlgZ1qQuBOFDGJdMRiNR9Ouc3P36lovmk
7+jtOnAKI3Pk2g+tyjRbynTCpr6kSzuh1hTHuwz24nx2xhi+B2wttRpvvZTIFUtWnIi3rdMuCr9r
w7KbUIzHSw51GonIdFFw5h2LuzZL4NETokyZeY864FdbO2MJxEaOL8lf6ClWAqqYszI6OKAZaLMF
UIRKIUxiMZk0rDtC6KsOwaZj4jNE1ziDllbLVSMfUpjTe6zsU279EGvTBxX6bnvk1R0qD4cpM1R8
MgdzMs1Er2ztbHy8WtfzkCFz1T/Fhk93AbavkdEGdNwUOT5fnfJsAuIHhDtt8DV4k0ehXuhE1WRG
EUbtDLWc9VT9Vgj7LKrMwHgtqFia9uFeZ62RNcTlnWA262w0GJxbneYplKNRdn/01SbFh5uWX3W1
S+vMBaKbzACOgETLqla99MmGCZ/fLzS/WMXWmNaoA3pf14MI937aBtX3stnRVJGQaRkGb1QTAHPj
EbeF7OGMr4iso6RBpYto5kv+CMDM+zqee5j+ubk+7oWL7ORg2mhQkTNsII1pSAn5oyjdPF3PH6JT
0sVhQt+L5rxTfIh+6klHZClIzHD+CaxI4izt/+FHRlEAOm+Zt8Tp2+H7u93eRSi4+wGvnwh2gOBA
v3ZOnNws7V5Buggs58AEIXA9EUS+gB1Go3zTg0z+paVgy8RdSEvMvbiRacUEGCCQNaOn6QZdYlDc
pLlDqf4SzKeTnos1u7wpod43Iaxcbfse623hGoy7zcvRDMXiTxEJkk0RzzVd8FZ0G+VgdrAPkOTZ
6Lo13i6X5SXaTy+t6lrOkHqJOuCa2sUlLYMg5PHpNz3Sr9dU0YiEUzklF/KcIAsYFiJR6s2iQ85Y
hNBbhH0TSE+CLnjof066N8vPqxJCS7W3bt5z47YAIQkpsTfgjSjLQeg9DtY3CIW75XnL/pDQpRwA
6S/lpSSn8LrgrPr0nl6O3QYBAq6FsbyGSJQuM7ejZQ1mp7rjDFs8yJWgdMfWeTMbTrLUXgxuQpYn
D2qJ1yzrbD+TqKVAy7ty8YpUs44F/lVXIWgrl4ncaRph9oBhbonb53bBiwzzi2bgz1RdstXkoi7b
N2xuALza5umWerLz7fI3rZuN/Llhsl3S+ulmJr1pm/otCoI0cjW5SG1YQfnvqIHFQgqiV0Tb/gQH
46ue9IY8MYMv8P/Q2+3dvJkL6oUPKR6ybWu7Pt2lQJ/ynRUBd3a04ajrp0OH0+YG9RA/zu5e8XMW
Y94X/v9nmudyyAkp2HuW5M9crnFEi5YEFQQ4s5JV2ndrvUm2D9q288BH5SiFI+ZV9huHIjw1KQWN
/mFBxNoFCMXOvCDAijMG+lqVyCqNkeTbvmMC9qr3cXtnbN5p2/GDe9QuHNjCNePHZJ3Fv0iBSVwM
L16cz8+oq6cPpVwHgDdWbuCX8TgPHbLAjfFBG0hKPyeoW5z5v5gvmx02xUBlhgK2WXW9TzdSCuUY
tuX5h+G7TjM1j5BiacM2YvwaRvgBkJNFCAIWhuYaYqngVf8LSS4sIgNLWCXfDb/5G/knm+Cyw263
bJYKGaaxtvJp4SbPDI1yOlR1HsbLQw9TkZAwXuZQ5zbilokdF95comCSWttIgQZFpAnSyrCcxNf5
ZvpsgSrGIBqCqknB9kOUewjhogBPEFyBH58aNRKP2Xz/3r6iUlRuYh8VCAyz3wlE2zrcxB7D/XLB
02XYP/2jfVxqN4yaGJwNNW76zs2mHamamRR0K3BkuL04bRObA16+ijX52TsEexYcAyZmKY0A9/iF
V4ysZXhpKmrBGgRSaJEwVjIW6r5iYGF1BQ70VLGclvhczaT0dX2TcbEA4rf1qlo00N+PPLAo6I/r
0oSq24cADuFOfzhUS+KX4hPnUTU68/OVIpt/Gg6Fc3IXEF0RZyTdkbu4Z8aAg+6zRfzVSIizXi+G
zuIv3nTmBj9cfboN1OsXCChERCFzuFVUsVjuuyX/hp2ykstdJc21S0izdYhuh0jjJX8RgSB769mf
JoY2Jx36TfGLP6PfCjCkf2cjdZzJdziEGuFrrN2k92sY4TsbHrjzf2heyfGdyhW0D3QEhOgXDtP0
Tm0VkzZ5yQI6RrDDfPPjNpFnNRJJS2jw/qn7crFsk8Jou5w1aUxB/5w8+5CtOJQtB0oi6+3cnyCc
1dWsrFYscHT9ORkpPuKkBuTdolnZ6eIh5EnVrl2HKcLcfMX/uA83jIEe2onaxOoIyMv2Wkb8Ed6f
myd91bc8rauK39L1diJ3TadOvUrsxR1o5pc2qWhH0ZiCpTWLyCIwmXwubybPkinSlqDkRUyNxiEc
PmRuVSylqAcwZF2SGYTwKZBcSD7AgCxsxyPxmAZnsD6HQbf4fi5rVzgRaFA63KY6myvDEpYqGDe6
lRYg906/w6ml8zlDMyeGC3IUPNhb2LEroBHY95JSZb8PS/jwam9kbcQY03GJ1nsakJWVUKCXVb3E
A6/jvOBRtpU0s0C87ltqyXCeCtMvV6P4CNwCwqkbIZu5cLgSqwtWjHjRxQKSm3I4G30gZjEDQtIH
ct5/47Lben8mI50HTj54JbfuIihbWwMuhEmaCulY3HDU/qQqMnnbiypguzgTy+BaJDNBgq4vHsUN
kQyxVedwvSr+RSW92ysHQYIMGn0a/KpKRptGHw5cQ9pW5vB8OP7FPtAI477zyhS1Jv60FKBtpVDI
xJyF2UR1Pos8utsXrXB/q2U6g4yvtoGzG2kkArqORYScFsJu/5Y0GplrFNYV2NQtyC/o/UeaNODX
F5/TyWRGlTxtgH6fq3BobTz9r9U6XXbnBFqXj1sIByfY0TBQv17IMuCs0kZX9/ACVUYm4XA8/l13
YQXaOu0r83if0r+QTx/EneBIShj8W6+bbSb5nVK80Yg/BFm7LY0xpFZOPzR5dM7lxyvLysSbc4vO
R+I4GBvYqtG2zVKlBZKA9toMiF7utqI2AB3AqkS1ucq3gbcbKMEHHL2dECB2REn8bD9KtnpwTxl3
IcIPb7MLuDQrzIlIe4yG6jGKIFFK9W5bDnTpfM2gvq1zDQ5NqVRj3UR7kRhZwCakH89QOMPIa4eP
G+wcNjgzrqXSbJqEqEU90CrN/9yoxB6Mj25UUYe2s7lCrvDfVwYvBunEjb97QkckOZBD+rwUH6Ho
yDIv/JlCPfE7MrZz7Fr/vLTDpnpM/Z+SjhgBQ4QPCmBFHyDn8kXxyy31u4HQktZOOgF1yUjZ2QoG
wmpEQH2VDYhqqgETT3FBNCJSYtJ5+K3Xgovkfu6P6e77JkZLTaEOzIrnWkSLhfKMXeV7VI1fHhzX
oLR5B6qfpbD6CBMIN+5CHaq5iEwoJT+yqROTiKHLA+uzTPlxasZOHquRusa0vg/MFJN53eSGObpI
/SPq0cMYVGRFIrHLDyNZ7OrPahthbrWHLZl8HQ9WgFVW2PMIi5Rt0C8kR+G1mi68NfJsKJQMigWw
QyeaP2ow2wnGjwkISuopScJBilhVYdXGQr2DU1wjBZ4JZJF7jorW4QF8wxkNBu3dw+iHFQw1EQEd
PvufoilBv6gnPxIbnGarY8OVF93wdambVZ5ek8P4bMdcf9fUX3ach9fUooGPHdD2lJGvQU3a86GN
HTDWr096SQ8J456s6X35jzWwdfONJ+OAQcOtwbKRe4FNrg0bWaPX4EAQ4C/ePT3AxNKZag8Rjdh9
v8kZ2s4ESXIhgP/BpDgwpJudupmAjfEf5unAaTqaiAm+800YVzZ9YlLYLOJep9G+KaVvNTtz9t6r
TY6LSXz+yo72yRzTkJ1sMLVFRL99i1EObBVa6pLIhrrG7cLJ7WbcVUGTJLdNcgPtozxV6gBdSfJP
Afgh4TsQRXzMnmRMZ2t67rlITS1KXPjTDZY4/Trz2ZhcCMaKAJxkpJtRzzwaGc2a6ymlBQa+tOh0
8V8Heivk8TwAETZbuaIOqWp0YdtImjfimVwEaFT1T22DfBEzr24dV+T+XgoDbSwBmkwC3CbJklYp
UaaGHxscge1bKBTTIMEechhUJaTtP+QdT5+tSf6z+jiPQQEElP/oXw8xbUoLLEg4vtoWbtXxTliG
4fAhpWBGRl3HEbHuTZDaN2C4yY+Aba4SnusLwBdHqfE7tGzaxPJ13ARrVgID874tbH0X7xTJhRRS
il3OQLF7HgJ+JYGer1v1qxTmwkvXzyfnF/5mO9A0MITPJdePVL1OZMuAxVDudODCsrB+AYbiZ5/S
L8KjDAXJJ/15PgN8U6nQ+kZ3xoYaeO6fy/HJZj14UVQ1SiwNh9yRNSAyN6AdvYPk3X1xt4zwfZeS
0OBHh8n2jrRVDtQpSYzrhxXBSbtBE7cqTSZz1hFRzZHeOAeXYJMFYqOQ7UGuY2u/wsbs7Goh3/OM
pR/r9FXwhTkuuIikHZb4shMl/6fROvWOgkGlRtQC8bTsoCu8Wlt3MJS2h/sSfdJx4ZNG3zSxBj3c
0EGMoVOah3gK3mehQlkXRXEgAEiSThs8xN3FCBnDq8aNuu5rqKCyBK3VkfGtAYFEOQk5bWgcZfp5
fR/Zv9GhQ4rEwWWrvykZgBfEGePKjp1CeydaelfaBn++OotHijbmllTq6dzqVDFq+UAYTgJN2Cq3
DKQsK8E2EW70j8T2YR6Sctel2EAicLpBdF6vZd4dCpKz3/3q+p00X3qfD5AdgA1zXkzmT8Io8Tvs
yRwGN2aogSAcb7TLXxoeOqd+JNXpMukLF0qUUjcN2cdjOThOylNMK0rHDPtKhz15zwe8wNxHNd42
eHcNy8g5ChaBIjD64Rzvo38xsnt1dAPMU/OiuPEIO9weP5nQ3lLFjaYEQCXF+kSTFe5gJXLT5p+X
gldNgcAzs/VEEyQ0yDr6bGCUcs6Lvz/1xUX/QaP4GFSqLQVUp8wFjuaIwRBh1ybh5Yn/Gtk/WjD/
0Up/6LwegjuWi8j/gm+sF24azKBjZhnHgtS3IO0vcd34MH+jrZCX8bX0KGKtjuWDQbbwrHpKFgoa
KnyM12qmTYYcebkMNvVcer4MiJr9QhQ7n7Gp54dakySALyhHB2rxT66UVIVwL3goIwzz7JBelMpF
7xSST9iNohjcUBswlDllUiw+uYJAhUdE94FVnVto6bG8NO8xKqKjju6HpWiF3RkdSUNbTk3qI24n
8K2o+n1wX8myPnU2ww1S4FLXyvM7M8bs3LbBIYF+Q6ELAKZzYKT4EHe3EFgGD3LA8UOGcqSRlHhx
4tXvfLj2tSYYTuU/2GoZeC3gPLHJvGLM4posywelT/x7KUeoa3eylMxTq5sLkJlPxV/EMHBdTJKc
bXlWjmTbIauEQ/gUauUFpF2NH3eM+vj2J1BbKEqrp9x3ffyaBMuEpxJ62ldXmZddp+CCuFhA2/+6
SSuZ64u70NKdsKWuOYNFH8rwsOdilQpVJSQ3LxzDuyHfQ3Et/Df5avjsiwaHpMDqOcZ+WUvMZ4r7
pQGpBBDwYzz2sgZPvj5V/NtWkk2cEMpkXe8y/BmNhznH0gDIHhgtO46W8Ddbl3UfJTI8peSlhcGi
EeIH6ktrpxqmTEDlwQxuM0dRgNipQkYVT9xDIaYOkZTTqSdRiWV6803vtd/eVc9ypIBA1FW+6gT1
GvkzmJw+tfXqeERbNp6W3LQ0HaP7lZsb4YNE02SdPguKh7l2eJpgJSBcLAPyD1eF6wA74Sp6s6Ws
Y9oN/8qy7CTXcdUt/INyhEy92uRTkeiCY54XrOEIiKP8qrMyOkJ7iVm8reu09GpcrZHTb2/vQLai
EiyzygbjRRGcLs8S0K7NjrqBRi76vK7T+fKp1RVnL7FRy7afcjUwSWipKK4V/thSO00G3ZO8xa1D
GZAkw8vHKjXL8RISYLnAKKhSYzlBxbZ4iF3Peo9r5jRBUmGUnI1U2i4A4N+ZaCg73GI/kYMMF2kH
Qh6lm1Ka9A6XM7dOLmut4NTYTdU35bWFIs9DzmpUVBAGXtYuModu7vjzsl7W2Rm53Yf77uscYcb1
lQpKH5dGUwtBYrP2Nw3xXQv1Mbsiou6OSnpbUswAvqnJg33Dy2VH3G/1crc5T7WwRh1YxohOknfc
FrTJbcJ9FbegrLJ0+bdwj7ruY9Zut1xvpihBTu3nCHQ00BCUzVMXjZsMUlks0NHuJkHnqOqtA9tJ
3hLqrYjrtW4PkJpefXVdlQ/E1I70RTYhUE6Ey6FHlIVp33l1qTPIizbSIl2MPZnJjoxpALnfbdog
2ngd0RrFo5yurf7lNxhJIjlX1piMP5EC4NtCsE/1dlDt6hNfBLQjvfFYude/sxBgw1NBYXYQPNBv
bBUs0y1lolc3p31OjgbWAOdVmkiVVcNlfqubveLZGoTYxJauh9fQYEHMo398Ke0/jNhRPkP+8Sb7
tTTj+xT5zj/5P770Jy0B+eq376B8ZVT4dJESdZ8qc2tfKXm3dM+XN7iUmlhCwKNjwCLpQmkJuAOc
JzWNg/w0tjwRFAYAInSwobEMie8y8B++r89IJF0rvG3mZF6CMbaTX6ub+VluZFs7X3FwZ7CYZAYt
C96kdmTS0MEfPmA+5GFrcUKQKzXI84eZDafOZEIG2HudkniezYfN4Q4yfPSmbzxpY6KBgRhDgZjc
gwpevf9Ns+E6trIH/inAbr4azprGJ4yxcIy2O7Hnjz655KT8q8Gai8oDA2qAZj8CZEwglDvHCuHY
8McYRs7aC7asVxHcU8uRoJ6obsA1IjA+FDhGhQPkI13yLvj7FoUcupXScb5HeYTkvGEDj6Okoi2z
TYXP+t+oX7Z55BQE1ljVxU2kUNLGH4KSTlu2Xwc+RrDjZgFnFm/y8jCuY9B6cFO47Nt42qzXCfF9
C3e5Sbl14qrVRu8Bhjy7XMfF02BhdaDokWQECInzEKweQBtxCd8r7I/op6K4b1JgvhyC0G3PULr6
6JIJHE9M7fh4xV+mCtjb7urkOwHzygooi2E7UzMw4hHqGszLyirJUFk1ulggGCcJ2eswAAvbWdTt
5ntzWf9vOKczZaolTiqQYGhWJhNieAxt1foDgT1XjCZWhpDi6thoCOhAakofC/XYWEiG3e3KrsbE
XBig2ZKhcdA71UI8h1ZJpONCZ0HshXWWkLug5z2ZFaHsQK5B40M1tNixH5b4jEmAEBYsp9TSXo7+
pqDRlsuEaKfyi/h5nhJjOYhvnce19uoE3/VIu3KAVlsS7E6yfHYMTWgc8cmGpilNGdqLGZK6BeoW
ed2eR6HBy7dtkHjRi0sL4lpDy62OKuXWlczWt3zMzOsDpi21DB4Vn8uJG9JhNpScDQP8TfK/ekBO
Tu5XRbuK2voD3NtMm4qfQuH09oyyNygDy3c/VxH8bEtJ7P1bJu6lgc8hjTVGO8+H1D+qi5EGsvSU
ZlJnCQtdtX0coASlIp4M2TinMOeL+GA5VGEcnV+axa7EE+hF6GR+kjy4fOd+njdKuMFXYIrZHywM
u8/CPzMdFHg0Utt+NXOSai3nhC6vAYmFLzsYDpY/TZg+Stj4MaKzsMo6nWl0f719/jpdtHF4GJ6e
hqWqjCTyvcOwCgac8KWvL9vEHSXF1iMNQ15fJNQvJ9bg7zh/QeBxK5aNaaC63agK8Xr+YVZQWxtQ
0YOcM5SSZT8rL1x19v7OAZYKcO38s4n2wElaHAFdQw2ZehGcOiHxByNQr3tdSlGOgGIH+sCbLgfT
TRVHTFn/L4jgEF4T04uXtZ3/uSXL1SlEn8OcEWB8SLdLH/IgTbOAewiXhW8AUIPb6TGOXXiQhzGd
tqgZ7f5T1CG2ndE0aeqjEIrtskQO1qbdv8KdR0GtMcsPdOCBUKYL4nUV8L7kZksv/nh+kMllP3oB
IRkv51w3x2dwdhF0E4q5B0FZYCzVABY+ihgtFTEz4cyXiaPX1pzDtBkUe9VhBRkkwI2wIrDtTD36
7e1F5qafj6V2oINgdCvMcG7Elc11IpYJ4e4fjpZg+vkfZvkasCT/qjJY3wMLjAQOsuyr7+SFp0Bb
3n3Klb7obnGtAW8DU5KS24vCYQbObgCgkl/xDj7Hq59UUOMXId+B4q8yroX63HvhOLDL2tkWyzdj
88EdfPVvBpSnfKHtlraCVC32V8Cs3sYCY8dAF8vmUZXwE43V+C/b9Pc2rp7BTWt/Z9oX3O3V6b/S
QTXKalEovdnssnXmglSAtTv3OSzleZfKFCJNx/sbDWyvOAKKYQqsEvnBwn14IvEv5K6DKk/PqIRe
UAqtSIYxsDY9K/IHvIIlqHg5daVUa71tCpzltCi7iKsxDWQo7zuYT5jyph0EwF/WG1DzbFvl3iYk
YuXcHBle/b5JqOWOZv9STHBQHsK1iLWSKRsskshVaPVROjgOvqWUs2mnqnup4PjQf5RYdd4G0cqq
hSvk8AMvXA6WHypaw0NcpqXdfEjK7PSKJ9eQQ0A5veB4NWLzff2xjWZqonEbLj99jukBWPqIqXSf
SP7fKL+xSsoL1snB7Z3KlJvmIl3sWQRZySKQAe0ZGbbVUrG+VERVHqDW1ybu+UkfqTY7pQlDcYaG
byzeR/PpMeEl3wAV0OyD+M6Ok2OzEVDE4pUg+cE9kCMx6nKYBe+xQjZwr8AvDnP+VU9EGqwfdMkO
5FGNpP7eAst9llgBX1Q0i+6DojLXMZRNyGtX0WE7Iw+F8oZefO85JBo+4lmWDD6VlqDdtn/5ZLxj
di2q8pfbsJDmYtHZguEHApxNxbBEFyZHGlo+3zRdhXJElx0Iue2OiHkTW7aBrHKIS7tvhy1cOFmP
01Q04qk5kKbUqfkHpkHGmNWFLwRKaJ2fMRpNWjE/Ije6ogXULClEVs8TCk4T5ulM5VYIWfjtX1yP
4pHMTqvh3dTL1gtlRAmYEK+qFOiwD73rF5Geq0PvzrJZcUuYd9b3OkCmaygfAzqSVe2okiD7s+hi
TU4OGpCk9P1TwGiCiU9bJvJqdg2k4cIftvdICjQUaltrWmxDFOskpb/OR8gp9lbzDiaJTnn2RAb4
m6BtH5+pqnQ9YWLZavBK83t9NrXUSSu6wVeDpZ6mT523yt0XnocNcd1k130ZT2AQn7FBdnSumnq7
BpsS8L2EhjTZdQXGp/ub6qcR+dA5wWkt0t94YnFa77AfOf18cKje+yEBcuf8Mw/pkfTwQLI4sF4x
2jzGB38H2BrIr8qnK0jaMo4OcXKvveNHNAzIEDftW8T/eeD3yL/C3QfZ3hUpRL7+AY+6oEkX7k06
6cpW70MV+BjYiHz7yl04sLNVflNv2XGodQ3nnsvVlhnbNd7M41egn1JxvCNEzWsNdigrHdlCiwKw
WZr4gFaPK3WpeImFQ0RfgpehG+wUR4x8RsCN8HWpY+iTRvpu0ACpUoGraGsa03hrGfy7bo+2iy2J
SES8q3vm8xhbrWbmlqgChBkDwni7MqRuxlsh1B6H1IfgmnKL00oR8F6w11eOcFgj/Tta6y3fY+IB
Wm/bByJtL+Eus3leAzGFhqvzEqZKuh+q+HILicPte4bITsqfsRsCF8k6H4Z9f9F+dexYEsO2wqar
QMmSlhBKKJJFsvAjA8TkE3WD/e65seHO+CaM2zhP7yZttTxofKWXNO7uk8we7NU56s4WJvF2p2x1
hzRDMacZDcSIr9NNnwgKE8bcZf+Mk81kvl0lWTChUAMilsXV1ssmrsJU0HSj/3coi43Z9NB9wInI
0ezgSi5Lq8Y2Dy/f9+XMDCMaHc6zUBWTV9sdEpIcgm+fpixHGzo/C3reIFqnORijrM/U4WGUoFBW
bJTDJIZ5lpazpTnsGPQuFo5bA7QxnCYgaPiOknGubQVlHhP/rnCfFcJKAMZRyZSxNgOUTFKkJMSL
/Btstqyr+MT47qntpssYOve9GHBK+EkYFMxFk08JWGLNsjOxeCco43Ar9rE35ngIP5v/DmukzeyP
aXyNXay7bo04jV5JQNZjFs0nWKNn+bLw2ilgh7OH/fbC1My12/AM9H8oiE7lApUs4Llb1T3eiUGU
+sPkaNMD4JVul+fd+BD5dC9l2PLnlK6QDckTgQM2TCCgIyCmo0XB/XpPhiyC5qzmjGVjaVYAKwgj
qrIMOpWgNXcjg+aLBLmFowkB9AleesAp1Vg75Ce1+wCQIcF/NmfdwrIgPhK+TyBCzBt5OVWRF1Lf
Wf4J0K5Any85st+MCI9ZIXtqNWiTN4Yht45ezYXmbtsh+t+cbcZqSnZNmozkeRdsArQrBk2ee6cG
kYxsCIUq1DmTORmtqDGQAasGBa3IZQv5TyHd11WZfDsT0qVNZcycVB781IvPknxOI/si4CRT+i2b
v5JyR9aJCeVcTNNaThrLcgRgzcuNL0sVqUnBbRDC/XF5I6F/BYU1NGHjinO5c2RaeNCAtgipZDCv
fA+s5JOuxlmvFD09y2IczXjOWIOFxWUoWR7MdBCLzgC9fJaGuJhtF/oKL3FytF32g3wG+h5pMwxg
m2kZlN626+KdtMOwTlM/gwOsX/yOlBGOr/t2cATSqqwk9COD3QvYVsiMk2SSbL7P/ZHYoFHLQGc1
RPsx5e1rTZegYZ2C1eLYDTRz0cqPmqYw3nWSCrOVpV2udTeNYX0wvZrxzkno82QDmAmvqQzOdR7d
jxu2IKJa6TKT31ShvhcYp0CSoY+0nf0QfIFPTfPXsZESJcPc1FNzR/6s7WAFhxRMi/WEtdPWqbaX
PDffK2XnBQS/zdlhTq5jeP+te/dwELni+BudfAEmyMhkpzSuM3526P5nqlGq2vZ1/EinYwA3WlbO
+5+UebdC6EcSSuJUO3AA4gimwEeDp0y24V+Qi0J6D/1aLsu80C4ZlXW+YoW2Ii5befJDuO+UFujM
4SdHCxhTZrUFh1b2F7o5j+sgUvQz/6cctxXKaDbELSAifIxf27Mm2Keli+DzQKKeHNEZgv1LXAlj
TCl+pCkVnYQY3Pk/ecY/12X2QBzm2wckfcD9yATH6tc7QPmyQunXjZJm8QsqnI8Odv+q00ZH6mW+
IHWZxjLtJ1Vl+WrNKbV0MRko9eUQkl6QAS7XbsMUiIkzXwz2Y9oAfti6/psaGb8waoRxi+/m5Cx+
grxUfWa91gDgL47CFUp6EBsv8423BkB+g9AC2FfaKUuuzUh2dMZet81ljCnwSty62LCWU2NQH5YP
u7NYJr8vYg/35Mx8C40u0EbUoGVlQBTosFWBxoN/Oo6Yy11rqIZ47cDAJHvAUmnKoJNCixmGMTTd
5Xo68SJD9neST2ghjRkMgoq5AmiJHFI6Gi/Eeye8YbSRnyymEg+jIuyzdIfvAJh9L8GTKDtCf0D0
ej8RtBq4wRYskWofDuXCB9h2s9kDpK7WwJWiPeaSYA2bwgS4+0zsHv+xHn0t0MYZ4cR+NCV63gBP
4e4TnkVacLw3+TgWSUbyMFRnRy2ggbJIxYd7NW0hBb33Dau6MCilrMHjMEPf9oA73XCkx9/ELdji
nttEeCd8cb1HEyg8MsnkzdXrk3uKfCFL3/vUOX1qBkFe1k2HJmhJiMXjf19w+vijkPSfme+MQrUf
DDZNsttkfAL8jmwwASmAAjmcZlsKXzXSehMtnSEsmiZnsItP0FZeweC+2gYVSuSCOJdHvwUw4Zs1
tw5LJnPF91ktuFjBpTe84yT0gp8qjGm2GT+xWfhO4vZNugRQwDJYtc5JAdGwOcjLzFw3F0OpV0t/
xw5XFoIS4m/OAws/4nHq2YtSamOHN4tl3xkxyt3Nr7oLvBb3X0dc7hu+Bo4fUx4/sAWf8bBG1gZS
Q/GZOHJclu7e4psIgEzewEAyLTWh36L6wnsIlPJK9vpbnp4KqGQQhmlf04YrdycKblbWP07rRTvq
yVTqDw2Tk7z6YNAmH362AT1xnsrKLrduv1eoLH4GlUHKc/kv08GmG+BZC7tHOjlKrCNC3ZFq96yP
vswoZihP6maIwY8OO6gStikVUe6OMIl5/qotcWbpThcCb1V8g2E03akCnzj8sdzwyzh7IRu2zhNP
W7Q4M1VUkiuDDfbIBqMq5x2M+pi3uxsc/VCTxulpza2M7tF+2zcmg/tt3TZKoHTDPiIrl/PiaPgQ
K63OM2IYPDTGjc5bv+hStlXQMh+OLH/wGkcvWnbL7cLhDNp6mKj5e/xrE5s12j3gyqQdXzPikG7C
cJfnJniuGc4iaHlaJqtjQEuF5wuCLGdXtyCXFIkwYJFe54+UpAjbc4JK7hCRkKnTsSB1eS35OmDd
B6Xl4vUQRt4yIQQc6NvJ7xPVJsYbhv6s0Ob9IPalftoTNhABkClHOoOBY6MYEurhX4nPSPPDjLdY
+oxyHgu4oyXcITRutLsESz9XHZYRWxxTQM2HFrEZXL3x9jAUXuFpPY+lWySP288WxGOns5zZPk/Q
95Virmk6hQCPEVGJb0qFoqaXyoG954P+BHk2FFxE71pGdWIwex4vNdM2rtvbqWv2a1ufMPKbFwDB
u7QFiU2PkcYrYpx3lV7V/Nk8/vuU/6ugVquAUJNhYKtxzmNmWo//4CQV3wRJXMznAPhnG41I3yls
32GE57vEXqOVwwMvALnreNkZtLBVzkrtUBQqISJ8z+7+3rBR9CmB/roLCBinSt+6rM428hOoh2+E
kmLTXA3A4qp57mx5M3O0vpdrk2UiZ4MmAAha2OyhqXYjzI7XH557reWsupignzVqbSugBjI3yFtI
UNcWZG7y6rW2mLlDG1EJFKMgf3OOheSrPh6W9a+VbLGMN2cGm8fGKB3HsBpVBc5Cy188oqGC7z+3
uCdNp+Sxsliec5nH+oRNF7578aTQWyiS9Gm3lfG9dChJOTYOxge4ZP8EnscR/HuU9lCKxWbd5hYc
bMNDRFWRWPwTnm+K8Y+6HuQ8p2aeCYdyfSV3zDhV5p4b/T7HicNZQq59S+1arNd5gPg5XFr94uxG
9J4A/yK4Y62UBBUH6EbcHe4uT0xciMHjRpKs8wmqEV1Oixgd8Jv52EuB6LhvIC4OMRHc0rkP8eVb
T9GH9qlaANNKbzZvG9NPpdLYv3KbvWwWPFU1+hPTWk2Xhjk154AG3JO3zpBlmWmaRAO8jhND67P+
GfwpjMm+/ajp8mWz1yZJXxF3SP+u1bW7jahcww0pQ1ZIezUUWTm2VTPq7G0Hy74Ew5HrflEl8wS3
EZtETmm3ci3obkewH0JstC+p9p9GzGFDsYRjVLkzVR8nEiNYOLNtB3JfCo+gxcQgzILu9Nn7bIZV
9V0nEfldCmAJ1kklN4+cLzsQ5OY7nO8WaRerRo+VfzVwXgUgnoLEaAHJ3UxsbT+7laihXQwwgCNq
4e6Fxrt1Sf/d9gZI96lI9h3IjE7Xs5DLkynrKDDumgdwwqNgTlcY/2gEsThHnHFMfIOnFIuL/ir1
z/s1geIGwTwU8hTWGC7gdaFlBOxfkLIS9Xtv7yMNfwFZhhNtcjOeh738RaG9r9RJnGJew7iLokqw
MI0MLnXP7DOm9pwIFBGOVM5M2SembX2yGtLKwY9xzbkPaIagwTM2KpUSI80faaaF4YNZWXTjz5qS
8HYqsz11ogoxxOwOShclp0t2e/FLaE/gtC0iWQEc6Obxfawx4oZ5mgef3C+MbBwV787U+gFrNuHv
aFE9iH0R8nUqYcy/j9auJ4aqi40qDOzFY6tSKLx0VNZ2Vf4Zc879wfbq9WavOU/BxhQcMfbDN2rj
AEWx/De3UFRkDBwiH8Fu4i35fVl+MXrbTKT8R9Nrf13Gd+Qm9Fe+qYQlI1A5EPB6jPmQKAbD5jfc
4PbSAD163zHc+3cB/TLiiGjMZlAAQJrKWI/UiAj+Iw2ObA2tSwHVMCiAVdOBVFUyY+SWGVPsmMDy
cQZ/n7TgIbF/YyzBSEcFhkosoKys3wF3WaQ9RcpSgqR/h3KcZDQlgGvg27fQZyn/NMLSPq7JNsl/
F9tRez344326wi7e2NV7K6I0vdVDjs1EmozCYN638nEvF/qH7wvSsb1ErkKiT0CUFYgCSm+1aso5
2V4P55nv9zxnpT78+QEytru6P+xfE97fgygnt5wmhmra2uD8pBQYcmkPDalO69xRiqxsL9kw3BRI
b+5Je7baVeIqNLauWBTE6Z37Aj5kztQMjllM1yRljN7/s/WiQPPRIpqdppL/cv25E9CYNqsueOhh
ZMMTcfdiTGMqGAdEFlIGWfy8Pva3MU5f4RTJiK7vDrDcPJ2xta9Jn0EDpt5U/ooPuEmdeTBXY9mh
rSpEnOA+8hJMcP1U0eIkcCjeFftmxWwyrvH1tIomgG3sD0wsrLOAPBi9pPttwiJXOwVKhWx6hAKw
Jdlo+ksPYJQfgMGVvIgD7BYS5f/QkVfdy90w+++jEnyZCd3CbwiL4OEjADYzbZryyOYyEkgW+iuH
5ZdoPHGY9Z2orJDhU8gkOFkHb1YdfXHuUYB6D5scT1mIgTGBVO/uvT2Bq6iPb63YYrJ9M3f4eGHy
1JroYnnKXYawH+R11YcJEX2tL3x7j0bjf4XJHJBPag/6hF3rLWjcnGc9q77RjZRf+tBnCm4fEevL
A4omysiqaNsJPH56zXS7sNSt2sHTfA4YowD/xaHnAbmc8GVWbNkBEIdqRm8i/OuedPihP7mo/WN4
JtDT1jrcbPkd5JXTK6BL5Zi7CIBi+EROEcRHAEipUoA2WrHwe4uel7p6OqYN9Hom+rPW90Ce8uFW
+U2+c++0CYYHEwN2ZYiKoyQD2F9IwJFXUPSttphy+wWz1S9MTrDg2jwg6TBnJ9MNQ4BXVDWDMDiu
0cqebrHy32vwifQdTOS6A51FKD296IbbecqXkjlBFxqtd+iDuMDav23YSchEwpdMu2vNURrFsJoQ
G7nuDYBtT4PDYrTr8wLjRljvK890funLRDA7TVdmN8JOGYgLLOOttvpNZe2aqjArjFryDthScqly
Si7tPzDT6fkt6C27FPFOUJlTTi3r9ttZSV7y3U5ocfdU4mt7ZeU75m9GpmRkBnWgtHHzJ8MNX5lf
bA7+Zmrpzkgohuo4dKZAuHbmewSs1uBqjvXNP/4kP+Jc0L77ubPYCZnqF53as4RbX6Pn9ZqZ4XAv
00zMSaksUYpGYIT5djgq3uixa4ONr2ER0stuV8ktaaD+9Ur0WB26JcPb4SPfHKWyYZYaIp3r2t//
Ea0MumTH6D68OKHbRPX7iU11ZOBxxv3Oj8v6D9DwGmP6MswnqX5QSMhT267QZhwytdiQX+MFm0El
Ag0RIo4WyF/b+S1yr+H0FS0aZbh5y34NEWdGmLEBthPj+3X2lqOmPqKKVxScC2iFXKK53fdF4Nky
3uk0Www7tKYrZEu/1+PayYAxDcdcXzkCYweNWuV+Yhy5BUkGGfQ5tR7ZoMoJlxpuZpetPlczn8iW
D36ulxpQE+PN9hNx8gBJl9tabbu2h6/6gVaf9BlTbBFAyn0hgzdVko5DRzyEIPDeKH6ewngl3zhc
r+TFEtgWveRT/akfzMZWAjs9JrrQpEaWlMSrKjr4l5NK+6d8+ttaw0K1N155AaDyn+Sjhcakim1e
siCaRZgGOPHgwM5pw7sLo5n8Ef/uakSPNNQQGar+IjOVZcgzaB+j7o65iHBO2jUhC1P6HHGOZwl3
zbOwcmHaiX3hwTuPyuXMAwJrkcyB4YYaBseZUCU6LZyHkNCOwXPb8Io0PFRqdtIMHc681+BwwQ15
YU4bpTLZZzXTml2ItHq61eVWum2Yv1XEykQGrF81lSG3EW+IcZrmCh1hepmXbo3WxSc1aOx5KMcZ
AuZUJxL3qEqewM21JMJnxBaB5tZiEXkPEB3FDv/+vGGaE3ourfJhfYD7aGLxkWhmU68gc3sl8RJ3
KjgDaVHmalrUofaQdmZTWcOf8VOJw1cypv8sOhvmfGEIretfl9oLhDIhIa3bXfpROWwxILl75PhF
fN20cCQB6ZPWPTkudPDOxHlpaWyMVU3aCqlMa2uxsm9UX3gDwoU7GMWzKGtxqi91Xk1/avScFAgT
I4ciFldUG5j3gs8E7e06P6atMOH8oTDO+oR8l2a8Zq4vmEsdMrnrADftyuqiE57PVAR0GBaQM3S2
Do77hnwm4zYgkKpCmPEz+rhV0Z6T/8Qi/LrI0QuvphQsvrocasW6JTJQJrcVQNIA5e8/p2xtKx7Y
dp6KNV/4WYY9bkCnCm6jC5Zc+77oD5yKbkTlHI+fuOBe2RUK1CFTlVmGzCaFy0kjH/qINW4Pri0t
H9yWLEen6PUZtEtu3EzfS7cBH1A3q58ZtXlLfWez9P/yRhXXaM5TihicbptgH6C8XEQps9sZqnJB
MpSp3o9urxUJZ/Zr9CWBCViIx2FKXNA0FzCax0dSP1BlimzWNLYivkCBf+VXIZ6r/y0DX5YBrVp8
hxQlRWhOKvtDJQCVhE4KP25gBVnZMqhoWLG8oVaNPk8MldHvf66EApglvO9kjyjNIdfhd6ka9WQx
+T3fePC83fmITee+3EdOeYv7oBPHQn73+uYXPaLT5KUhpIZh0oW8x/kolz7Zq8+zPaCqbS4GVmcs
muDywwnC3H6m6pqCnPZTq49cw5THV7MfeVie3INqHY3/sOjDsdScNS/8qqVYe41G3fZveNFBbqPv
H5gRFZVUGGtwD/aeP0ElKQeHOJMSIV3OTuagf+RRLUpCSv6eiaW1S+ibE5/DpNrPBv+T4d4hmfK/
OM42iaGZoJogvwDokObpGYvuAHUT7lFAJRsxKhVB6xEnCwT/JUpKEis1zcqek7m8qapmtBavE/sG
y/2MmtAjEGKpruSAgMUEUko05y8xyaqHEhx73rcXpJo8eMpyj/tT0sgLEnDR27HjKGcLsL1VZsjE
o7PzTlBjiF7ziVXGN668S8RgzdRQgbe5knYy/ZbXXT3/iKetsVtCAcC3BZsrgnSBVNVJ9kcs6+dK
CFeJnmh0Bdi20g/MwMi9OMbv/qI1lwjj0XvNkQ/h52/rzkbfDb8f29kpTbV1AZ6G64jlFUNqKmGy
DpqSVAB4DrJ2SOh4WtX2ncjZlZ/ygN2pyc3Xu6mm30jbKk+EFYASp8kCTFWyRH2plHEljcyyXS5+
9VoFGXPx36n/FDvtO/WuPWbNLO6W/f6AkF8oC0CwHUftTvArJA/kZWyWp56FHD459R/dWje20iHR
jcYEyq1r67YON5HJK5Am8Cvi8E+OmULs83R6vzTmOcsgn8J38p596vt8EtwPZCXzINR1IQaX3ubD
PPROb3PoXzQn1iu/DUDXksVAIGHS0WFogTrMMOJ70BOCLhUsZTd1FSAkXb6SFm70PBToxXcC5Pu3
+8dqEqD1MWe952RHegeYd0vxudA13mjZn7a55+Z6U0a6ertV/U+FcJu+PtdTPoE1m1ydFie+x0+2
NvbaRdYDCfNE0Y9KTDNZz47eCXVm2uhEUT7KFPiCJ8XqqNu2BLMGBhioD6HIxL6kzM6q79gYpl1L
nc5jr7u2pqjvvueNzB17BjqhiGDsH/PUTdJ0qi7Iyt+kvJ9o+OCMaY6x9G1hh52+wYkAK86golM7
2KsR/yRgkSav90/Ld4vX9eScAGlFRghmuRCxnyH2sywlPuxiz7OgHRw5g9GZJxkn2jX+XY8A4r3m
OG3wTRhUVmXP+EcuQKRUCKsbH7QdhKZdtk5adztZhFhEOgW6yWdIoJTqJZWEnVrxs8wIXbV38wGw
Uc6ffNW0hjRyDg8HyIH2GjHckqcY/N3jYQcb9tOw7MYvJDdvHgQjCBb5lHC59J59pQzQh5iYfKod
0nQQNJorLghL1ztvgP61BK2dNNqB0Vu7PguBCzsOWSlRSKizuMU+kBI7HE24ZO4hSs1MspxDNL+9
sDTJvAtBTZIAofX3ZdRHFFaQdiMxG0D4cONhZLPRKIZ0bhKK6Ti+BP92TNFhhl9uSjxhkQNQW6+o
K3e9xJfIxw0dMWugG6YaZMoCaNVizJrtqNXopeG4lmFT4IRSoO8wpGtknFhGpXe0QDQn4a+XRZ3y
2gBfitiZXXymrBZsA9v5hcMq+L6SWj+y3RfhR6k9QmyR4TGetfUBNZ8tT8PVUCEiyv3AwsI/Ot43
8GXQlrA9Ld7GnkrSYZBCMXixcCQjp6xTUMk04cdmxkr3na0QOOizwLfr0MWQjBfdhitAlFTEkSZK
l80AityaHNe2FgjeBsGBuyTCobWbYYNjNgutOSDcej3UyH6sJpaSJT5iPJ43SERahx13buPn46n1
yEAcdWjqk8PuMMwXZn/lSv7qOAtaz7v9lZEqkjD9ypITYxyRH5rL+Y0S0uBA4H+G62rYLaWKtl+l
5tP87bxHTl2efk32RHe9I/jqcgm8c/0wRvDZD7aCFmeMOqhDLRxdFsATVDd6J+5nyGkk3b6FzBDT
7vinKcqh5b77d+H8MH8nvTVzhC/5VNGdfDbmNMzugm4hg1k6hv3zgLzuLVuUXc+yRkI+3t2jcRYU
47TpCullZVAzC6x/0qCJhooOy+ylgE7v8ffEcN7iOTSihP5xurduQjx94v2Y6f/m7cnuOZOZf9Xd
GY3GF/QJ9SR797sUtGCwTAzUlwAOuBZQWYzzuspPZDSRzgC1ixeVtTXbdcmLSNZV7cO6PJaMbbD4
sFz9y/iQHmdCk5/I/OOSYAn1IzppSvQRBpTFUqH6bo1CTBal/r6Rj03+eed8iP1LFl2uRHRON8bp
8WGmDH29YYpTj6xk4GTEul88CH3bvkwkWLNsEcUY7DgqmnClDX3sN3eGD50IKbgNUblsjXwKMuCf
FRIpV8s1qcaxDyf5dJ2htNGNevUPYMQaHpGHuYXExfFNVzx/Djt4XgJ9dRMRfQSL+OXjbdWvlFl7
KkhZqIspQjpExYU42ddYzT2anI8Re1oDibxTAgTAC2pJkaXtyu28ndxZgzi3ubQ8mbXChVfwctn9
T3MJtZd7LbksYqE97ik7Kb9zreGFH2s80IHQVziPSHdu7otRfAnCCjNbI8nexyPYvOr9U3uotMPc
ss10jx2SzwvIQ+ax9Sf65DeuT0m6jeYDaQ7mrFno8FM9/H510a0paY3MH3XkEhtfAcdZNifzUKtW
/GsLTTF8YyyX+IaXJknFv4eZvS6J6xlOU82mjm28KmEHXPQzO2IEPyUXBbY9J3TX06ZLJpmBlmvv
TZEk2b8uXQ4trfg78WaLwY1jgDoAKUXc7Ff/ltbmyP5gLen0bcsF0GC5Mmt5VXa+pwSqifrA1lLm
MR2GFcAEXfRabLcslKjlHXnss3rP55WCvAsYmc9GxSU5XPVcDyWeL/UUiA1/bV3+2PrsPXElH1GE
ClJUacBSt9IjKrZGOaDBnPP3tkDaGYnyVIfg3PZYICw5dbiFF7DENKqJdG0/mB0/pKpOwPyFGBm7
xXJvi+AAhXvcr1fY7vzgnco28k5nI6pfE8FqCf/1NOUstz4K0yU4t6w6Ci0WQIxlHnJFPAbF1urd
DN/fHyYyRwerReSMU3Hm2b9NZ+47+QcpQv0KrjRbUhLRuOcHJXRLjriYroS20sTR/4f9VCcVeaGM
RdO32uOYc/KZbMKiMLJPnwFy9qF0R+wZIqQIHP+Swt8SMRew3L9z5IYmK8/efslp2/Ka0e7t69Bx
kgw/hpN6nCgoGDcHWgWePPPWJgPuFNWlza3emWitREz/O2oZdrEeYIJxHTqAtHubprvjxuKfPvtq
l/Z6LBbsUtp9Tywp18aw1nzFjTlOtGW85aZ2ZXxAfULD6XwLlgBFRflSR/lfVSK9tGxr5U3cWh5v
LNGSU2/dxB7mHd1NdOtBUGnNC4dMpgJZsqmfUAxO1o+ME32RGTTyZ5mMcdnsrNSlhzYgmRDQ7Gfq
SdTumLKOEEn1aTneda58rgtonQYwE3sskuDs+QHBbCVzg+HY+mLffwbRGjxwnBUae/mBuzQzKPWU
wfTo7jWa+uC+EwYURYH6lMf/uHfZTOBxQslTdMlTmG37BSRis0i6WzTPYM08Qc81OTwvu4V7XsoK
h0vMZfesZTaylluB8aDb4DeecsmnnlKF40v7RcP8tx+BODoPYXjWXR+FvqROrSaORPjvCGTtUA7q
kXt+kgun044+Qaf1qJzLNqO/Zk/B70XSpg/YUAb2HGrNYaIobFdBhx1E5SSwxURVx+IBWiWj7mmV
rF6nQMB2MYrvkmVdh6UMEKgLJeI8X6IEUDAC4MG2pXkkdQMKv4UhY6Hg29X1wr0c7obE080/w+Iq
tr2hSwB8YTPCpBPAdmHBDi1NRWSFt4hrItcY9nDG04F+i3s5yrYZG1zCMI+n6AtvLzhKp4buL9LC
K8ShOri03nk5Oe6dnVQL/bQJTO10aV9kfxgoMNyizTbqPLOQYhogim+dAx/qpv20pPz80rOBPg7A
i501+pcuXpSuLvKfqbh7jn3kVycV+dgszhAeVSB4f7yn9iPm0ncO7IFpEdaQOxS/ax+bf0Ci3iBK
MUiWewhkRgVCV4bEdd0sFu0hQzMfkmxSlkqHgLiXknTKR/n8yZk0DAnvk/GdW4NQNkYyty4VOc3v
GdGRL14hYRABsKlOX14ck0XvH3hphQa7AsE5B2uKuYIfBqu3IHlZoQUxMQEUEioMuEsumZz8pxgw
akNPS/b2d1JL5frZaGC70nl/sWhEA+fA3aHPu2LQjAjvlL1PdnukCpoqqzRu4uqFJ8wjCltnIEHh
BniAoWhLvEvI/IZfDe8bJuz+DtBaouwk5C383EwOuu7poU7cPAXMsALbo1HE3drEcDaqCAAyylMr
ydFgWVXAwbWOa8cvTPjHxsbTsPaRbyLytBB9fZwQI3ZYAUVsSNB1t2A5EysX4Gs0KT149qNYh+nS
cGdEZD+dWsbInJN0YCDfdvtEBERZ150wkQpnD/aR4SqPJyLr52lPYwr1t6kzItm8QMgwapANRp0P
WxigZuEBMzPJFwr5GZCVSGdg5f5VJcw7PPALWqcdzsEKICzVMfsvoUCkP0IVRessG9wuoUxApfXY
a696blP8CbjhXL7zS6JartxwPjPnsO9KuCwGQag6xTdYGwHZvjfBTu0r8tBhChGQhOlWR/1xyZUJ
CRdkJe5mXqyM/IoOXANnmXM1G4802iJy5W12XSde/pBfUufVa9I71kfI9uQiJ4uvMVWLW1Xj2rBJ
ybA4RoxFBPPa03YATal7ojMVofFm99t7enftP68foo32oAksF1BpLEVyRG/KmLthPs0JEGDNOZs8
G2IPJNYrb+A/W9yANAhCOzwurhEhu0/kOleN2LrkVsh1iaqWMow92e1wWlJrpYvVaTuQBlopneUf
sBK0Xqb7o/cB0Gn5nrWDaaMEeNqlBeOv0VZZ9/GertrsB5GrSIT/T1inTFyhy7Ky+IQAV8FFYoMo
lzd5ekGF3mmwD1uH3f95NaDJ/RTGsXNRaSk9lly7spf750t++/0LscQ/UicdrqT0tiHz1r7N3zCY
zcuABu1y5OgRVctsmleD2mFAiHxK7+0HsT5f6oyh5U0YTY/3ESkk+qHhTLp8GQORKb7TEdg4yeZm
QZXfHc+0nxOY0cUND+Nj8TGJ8BIiCTNTbQnplqs3XFkDrkX8YLb1BlDy3KM/HXOowTd2qbM3/ZKi
aamHcUoOga7GWLRAbR7RjQZX0o/A+2S6QhsELtpPohSsE1bERrCk7wLLC/R0b23LL2NHZM4oAY9Y
phmjVUmGfgbG8/ggvGMzBys/3ATQ87/FsKSMyvm3ymuRYlYj6DDQP4oxw/ldGSCguN0j/EL5pXvD
g8TDnfTc2ALUlR+wM5cqpdRx9ZteDX+8+4Rye0X5CzyTFnNdCAxgHzP/9usV0r7FcdHoHRpdXPKr
wuk8QmasCyWFKHV4x+2dtxH0Tah9Q1xVYRqFe1bocuC1+Rg4HPTM1v281ND3OTdDewk4sXdwRtBU
WuOaXyrGKlXSKyb413THsFtBvK7Ysh0B+etVUinnc5rAjmk2HAed/1JtIpnrltkVJ1uXxr7dRh21
WBENbtsutAUXGD7DXZwliNBVp8/l4VUW1A7cD8k2yW2MMa3DDBLMR6clTz0ANGEU2aXeSZvBr7TF
mFy0ZZ4LfFHobgOjHzWUtuRlGihfu++yhWLi1l1WoniU6jrK2yhrpsjg/pDzJRGNpPJYHW2cjXB7
aKVKn/jpPNmxC5OzoyWsYCD6e4Wv3st48YKajOoV63X6EnF9Fn6Hv3c1IdhbMSFHH0E3rgDfK9ad
X+Wk+hMy7PAu4gaNLXTuuYX+v699mDYkj6wQ6V6CuwcDj42tM/7KeGX/gO6pwuEWlJL9ORVrVWKa
WHWMnk0N6yQPHbCBH54vEoacgrN6JJANa+LjGkyHjR/zh5V/cUHzEEyAtDWyHBBLDEFIklxTFldn
cqIsoIaZ0+DSNoofP6RHtp3ERVKPBfl/5udDDekCwr1uvFC54b3e+lgRa4aVwnge8Pjgu/WhT0t6
o/xii0mKIw07kegGon7vqLNQwLyFaJqOdCUo9WRsBm46lSlIIcoKBORpISR7QOo8QJ2310l3Ydru
5bq4fNNSV4M1Nsof3PSvpbLYaB7G3zmklkT0qIAr6Sfb50s/SeBeIDa9HlG+3FvsXrXKX8ttZAJq
8qmoBoFE7KZa16CLU1cmhpX8kmNDt4Jp3Lop1YyhY+rQHv12P3kGmiyGGirMie+l9hq6KXhGqPZm
bK2g2eYbBnmRgGiKawS1BrEfB35Toj/P886CN/OZ+ksQxdi8/3xse8NhhGNQzvwx3lDSvPeMEzpc
w5el3GyhgrU+TLhoxAMyKzg/l6TYuk28i9jthzWC4u7xPDV7n/kbA52yxkULhRUAKP1vcb7v22iK
Xu65MJZLyHZIPY6ccKQcPmKK6HapRv9RxLZfilt15Zl7zzbU8L+798Q0bJaNBeMSXHV/4D3QGkfN
W7gYC2OoYIE7aVKflao5j7GsvaMxVG7TVwczvchnpVjLvHG+ZJ+TXErN2rvZGZDm+uAPb1B3W3r5
NtSHIidI41xujxc+sMUEUtfX1pTKwxVcoIWuMD2F0YA2qFUBNhzSsMnjOzfHUW8Ofcu/OcdkBhTu
vCdp9R6MqIs8dhLZ3xRZwtKe5zdHumSV6b28sXCIuLmHaxjZaAbvPkgbMdt5rJXgshP2KRUFmv0r
FiXZFd0uXe1Bb57AnmWtrF8whxa4ZrK1m3btMOHh/vEcmPwau50ofH9N/zXjaoiSNRaC6YmTeukC
VVNzTOe7R2wjyPUlnu6quWltIcxKW1XMHM2J50N9UYBJYrtFvH94nMHWq3aoFzEB0NUxVP8MIw+C
GxtxUNswYqK6nZDUHK7BERDA2E9AhgbB4rPl4adzF5F8OdvzQ8qi7bCwz01x8XFX7GtNyYUd2EUX
HQEbcPLvG2l3G8OtJt9VErzmIvd1eohHLR7liqIyOK5ZFAu7UINoG47MgoHmxOUHMzjKP8mClRiF
jacxfiHt8OFKHHr4+2scTXMFsG2xZehnwHm8EUutR5FKtO6vznv1cZdQsaqsE8kNIYp37oE8aW7O
+8SqAwG33qFqUZnFeto01HVLMBjvDAa8bozWo4Lpbg3BVAh12gJh9U+uez2Ro6Xc/2AP9sfvB0K2
/e2U7t3TCgyFgsBQBKnbpyUctMftoqmhn3b1Vpt1l5RNFTGkn9AgPLTs1IiD6GVLEBMf6CrNU5ax
v5aQF91tsMou8KSIo5eCYRfJe+8KzpObFmST+X5ejRGwF5Y79WeH1+Q90SNitEgpaBVI+KlyCySG
VtKbYQwNkmXZNEmQo+RwLjMrSYU2rq/UVs0PPFY/6SCu9wFXW8FV5AI/LpwxwzOClHCVyDLWlIoj
4vfLJrOXQe4z+hC1sNpr5VJ23BSPCM7G/18CejHLCJuWtvWeJdb8QJEJ0pd2JjYp4syzEScobIaK
PJ0ib7HPUkX1+0eVjIN4d9TlV3ROoVPPxicsw1xFcftFHSiB1LCqbpMA0/umXwRL9OW+Bsl7IVSJ
gFwZSIfPYBptWrmn4sjXPxPKwkFLwOKaz7JC2mTvxKRJDGhB6JiLqEIzOFRnKwJQU5Jp2I3otkQx
sWPe3h+I5DQSIri7o+glFjJhWMAQmKtpdNV7VL59W+i8Alt6nsKGC870VF5GA3UvI0QpQohXP7pQ
pmQRAuiWeUjo5PTZoJ/WD8rsZy3cYyghBvUk1ZqEqkF92yTKpQGO+ZuYDy9EPH1Nvu1rwWkpDi1y
pdmVH8voa7ko39nUtD1cHBvCFTZ9czAeKv6jG3R+ecwGTQU96cNryIDCuJaO5RIAMp89AOa+8H7Y
wXeb+kBwF1tp2MKi0cjq6OlNzOb3pG4t6olrHbSCeiw4j7acIZu3s2hyS4S9Szqsz3Ac5tJv/l37
3xxTRulcd2nLMEtljokMqNV0Nik301m39JZQ0nUChOHa795z+1nRv/xwcQ6DUu9dZo+aNfbqplFd
hL9qtmQu7ZL10kh9ygBind5XcOrAdWewUl1fj7YRTLDurZbBg/pLJ0Ekd7Bd65lsuc/tbHrIYJLf
viTaPKnaq4O1L8Nds0GH0FCqRleAKmxmXxAt2SSIbdH076b1x5LAdnN1HQ7cxwQ9R7FyODC+luQH
p86myImvwx9Rnr3NHbQa/B8Ao7qJKX2tRRNkIvtkCLP1WDlE3a6z5HrYAy0zhyGqifkoMWNgJ7nR
ZIMQeram+QNNgSjImpBl+aJYJ/AnFmYR4GftXRxnlRPvNEW2YsJhCOJ3eh8x+kcID0IX63YIts+J
wJWI1RqbNt1w9qKeNbBOG2NVeDc8rkL7E5GzgpEPJcUMA7GE3elqi+eatl2nKXuEJLGS3fllgCfq
4neJUXlAkrD0BkXIxIVTAfVzZHhwEvrd/TMEI/Elr/0jS+VmAsOMkKhrMNXc8rWQxXsI2iRPCmwC
nizjSq208PzjXYOFfKow/RAkoCBsXILHC+l8xnMvaJac9yyC5JZoFNYxOWoLRBWMBNw2GcTEMWO+
I/uBBOXnRyHtKGZ3/8QgyGJAA7eTPgyncJG6HV8w8tDI1zZjycDuZQDsqYoZ1/qipB7ULTJSaDKi
zEcxXVf3m1b+tK0Z3faARvwTtmeikSOIFRqhs3YsAFVBWN3VITimleOKGw4UUY/qYV8pzoxmcMxx
fU5mjyEFZeWmWLAdxtFquxyOXzDNsMENy29OgSwkKRQpG8Z5B4FIgzZqmKRvEaGzmcw71w5c1D6f
+et97sJJWNy73n8d5MGagJ+BeFLPMVC5BfUgFDTDFZ57LXdkDjfGpvXyPbcfmXnDMqGohrZwSZDB
L7Q2Qcvn4YvBlptCsqe+dpVd6f+WSqLk2/sTvxo8yhD/k+t/YyHB5oYduCQTwnNXmXylcZvw2hGQ
Yku/Q3/QtnUx+IV10T4hSJ34KTT9wRZfG8RrWOhb2IiPqcFtW098uGGrClAyfOk9KiDOW6k1N+9f
c3c9FgZvjfiVRYxQkwJu7CHfRiM81tY51/p9WH2q/hewY2BemH6azbqGJDUcBXWV/Xbg6iUiMJfv
2YTlX9je+2yIBUN7l6T7lmJsgTYcjMGd9bwJXgNkLUfR+h3aAI7zOXh0M5M0yb0PG64TDbyrjZin
TIxmBRja454aPTXiT+b9nAv3A0L2gYQW1bxNIGRpxUkaXomMVdFU4LfNLK22SqY6BKJ8oyLpO7nt
mRlgVPPcP7HHBdG7peAVSuultVy9IkZ/2lehrRx5lSyt4DXIFPFB0gf3UdZku5tNFxwGbZJ6qL1q
4RJFlW0ZjcAg+Dxs/KXP5rpJXSbijNadqzOTC5VYDUl8/BBxLAXPTp/xplk5/B/M1N6h24DOxziF
ZYnNlFpAon5IbSQ0eyVMO2sMAes2+6LiY1V1PFRy26/jodfJs/4jTwlSLJalpeQxtwbgRvCqTn7t
KKA10ie76qNl3bqtnF6TJiksBBH9goRxwfhze8FUQgFf5NtAwZUD7exIFXaF1lneuId4UjRkmLrv
Bjea9ugisDEtPYhRV6M/JlfuTUCNLyoYNrqFcttqMS7aWunvCpofsfRkzJWlk7nNExap8Rpm0ROE
OobMRKE2EsEu/JIFQlnL9+zyVfeArOk2q/1TSETmFmrUCp3B06PqSjLYOX2f6+qhKjuGIco4hO4d
Oz/bkrLd0ay37Mt37eQpZ8qSU2bPzsFZoanTIqGMkpIUMEg0keC570eltP8QV7dRaBOqM1xu+loI
VRA0csokaqNzWgOk8BM+fHYMQpCCGzfacVZrXJlRbMav2ZoD21hFDJAxllCdoITRzzcSgCv0MzJv
K7bnNf34AGbUd/ABcWFL6yxlRpK0WxQcwFSONWEcgYg7K3OXhqzEzRfft/CZ6f/frypPFr2lfFhI
wwlqENpgS2UwAa+hH45WvW26IWih9k/tWyKOPT0G+AnVwhPGOocfGBv9lfg/Z8nThMwjeekur8PQ
3CcF+Nd+O4DJhxNpIsnBYmPEDS0cVcKQt7g+T7vW4tz4gPDuUFOWnguPRiSSncl6tbwe+IS+DdKv
z5qccjGlYFgxxzsPoa8AUAhks8tlrx3rxdE1+RXuAx039qdS1TQCsNzf6NeEZiBVy05ARSV4qsMg
Nm944IzBwfeQmUGyUnsvekjuIgIeuS8vE4yB+uxkScwFEPjWfWNtWhYPDWdXxPyykqp93mFAqpyj
TSjPlamyzgbIpmyoFq8/JhtIkKm39sq+bf6xzKbBLEWT3Asn5Vcms1/a5cYkCuRHywHOMxkrFt7u
y6X4DaKn/w0MwfTj3vLLQJnm8OshWAOBeznhy7GF+Z4eSu88oJdfYNpbONVBAyIdXTApC8W2VTCt
5LC0/pmsgZGlp7CpLFU42p7ukpxprPTlt/mxXxkMXij0obPf/FmyoHdAbxOhHelYVo5En+kCI78I
/dzc5do9Gy68xxHp+038SS2zHaJPsaTgL2IJBeGg+rkn6r7b3JaFoRsJg2Nj0gQrv+PcsAoA3Nm+
CF3fXnTfc1ijicul1ZXJPx/uMwE6KLc+VwNOeNetyJKyuucaDN3I17gpjPSoLCUX09B3uEKCc4FB
v+1VxM//K7rbEqB3GC6v6YIYeIEBeIu0T538xrHw7R8vCNH9rF89y1Z0CtpqV7KIMxp244qn7wy0
YgwgcnUxDKLb1twsZyvbNr6E3GEKwNUOgcAn5cc8f/ncluzcPV41wzOFcbvIqEIc2kBpGeEZ0YKo
hqwAlXA98AbzXsageCMRAYdQihm/3M6KtIy1kVvZmty/+2+wdqOtePNqmE9oDz1NRyDSF7vZcKdD
zhdWp3ktxpLjST0V9TJcuGTsGxghJsp63IDa0b0IslOVi5MLIHIBpC3Z2D1d0UFdgx4ueMNyi0KD
N3LusCsFzbmKZe182HfWO16tGGEHkD52i9FRdZhy2HUqzvF+Vdt9Z5MmL2nzkrq2rBjHbGFIkSyr
zW96LhLPmSmUVl0Z0buq1qa/nBnclmngmI1CztQmzv08bixLgcTrQaAUyjvbKS3yWo5FgAZoyhmZ
SfopkdESMlbCx/BiGWZoTjneQ9ajzUQGH46XWCsrADvOtK+ClK3McA27lYLThKc76NeNmvW1PaWE
EpAY5Cv5O0ESrqJYiWb1IWE6zcs2GEUek9AedkbBOX5EOdAUQmBXIs3X3FidcTm6EjZ7CAdpx9uf
JXycdvxpQ1z1lRj4QDrSuMOlFJfrAncTJ0JnoS3lW/ilkYlqb9WXkQf6164EVKC8817TuumJckSU
4YxnScjEtQUEKiSqoclGs2bMqoer6R37UU16jJUVyUQxD104OHMMLeRf9l9SI1OAWlXAzecCO8Ia
b6X0nRjap+WTUf0M7PngCqGd+rMf6Cwb9Gc4AAKgwL1fUqWL1H6gBqp5zYhkoG3qvmlbfwalXkz6
YMfGQn/qcEjfyuy3G1r23fLxHzpsT/Er67q25CBYwqW+3v/eN+5pz2zF/Q1YyGZH6M0G0inYz9HV
CY0dak9k0KzeqhyzASoz269JBWfwXkW0/sHceezPlQLtNVfBT94tOgqOhel4WoFXm6UV5zlMC5Eq
3AhPZ60/OwAv07IgW6SawRhdaYyOEjB1nltG6KADVjzrBd+YarqzDBs1iA4/XsvzYYmTwTn7TkU/
Am2hv8Vu61WNIhfWKe2aqK+eZ5rQEW98Y5LqH+CX4h6W3bM4mu9P0bFF+bNLNPWssQbcrnqh9hQL
BDJKdyH+OBYcuiFc/l8nhowaLj+p2LXIF1Fz562iblFf/Tox+6J6jUcdlzdqvNilgQ+24mpZe/V2
GmLl+CHVyFGHERFNnejYEIItExfzKkrUDewi7nosUVD5rIca2UgfcuuKWLOCJ5fMeiE9EVPd5C85
fvCo0bwCynf4Jl7yx/8RDXVDknlZX+gI/jZ8o/11eYQvrFgG+/vVMMOtDkczApWKPqgTlK5urMV6
dJmkSb43fp5xfKd5EV98zATLQadZTRPKL2rHT+PRXvE/5qMJeO9cpthDn0lumAozqY6KtZbhbcJT
uWp/bfOggr1bpx1BC/nQqR+xwuR0/BxB4/tWCeq860tiXe1Z7zrmjtWmTQftqYrL0LPdiy/QG7US
zvhYA5F39VzM6TgXNe2p0KgNOhTdNfTeu1HdsjU0kuPKEDNpPGMW/vIJeco6jWH33FX1tQVioojG
s/A4V777g0n792OFItzzLzzWnWeGAkoYigrRsYjfi3zjdVZRMNRsx3RFJE8nvLd9wJ3pANsTsLrf
rwvhkc+Fe9oFipCFwd1HKvhxZMDIuac9Vv1u/D0NphMi20qUN6DIOwtnG74dxW0liWasBqMSw+2c
sHHi+bRI7qkALmZt89YCn1kJ1zL5bXtDPhMJgG1EL0Zg3Uv6BcpfMgbW0zN8JLY5QoZQpeRwzBJe
qgCDXTXyXccOmaPKXbPeLWZttVMIN9PtNiTSvWt9RbUubfBoKF9Ro7CsxGn/Q7LNiXcrcyrZtu2l
OPT/Z9ngMdq3Z65af4dy3h1TA9jxXDU8s+lbwNZGEzQI9hEnZLPet0fz5p4uq9UlH8c7zvLnbyTh
hbJ6QtJ+4/eo75ZlF1odrCaWW1sq7Gdc8SDdZ6MjLyGfwhTruItiHTyLkciwfzPMIxb2zbqfc/0F
1mgzgUST52SfqU3KyX9+cjM8UTlD+a58V69IY5RsZ01crJofq4XXx+r9KXksIFEbBIOH4RnjNAFd
VgJOSx6K7cNis+aODEPJFP/vYTJ4mxXPp/typIWxxBO33dj0fK6IOJQo7sBOcKhI9N+57NnYLAV8
EqXGqnTLn6TaF+2u9HOlfVSc6xXscBXfpoE6dscnUXBUMb2vqWDqFa3Bh1g2UvZp2jiDCNEAxiXS
7z2PuLiVWSmc2QbTTJ/hg6djaw7umO4SNNqwCMNFEI1DDcKzy6r0KEKarXvft1aVY00HzE4AxA5c
I25F9U1Zjy59Kx2fyVG5fH25u7lxSjZK2wdASzA+lKNfsJKnaR5V58cLlavF9IAqBnsxksq0Gw5X
rMVQHjq9Y3pDoY3P82UzZRJIekI63SsAnacDHipedwAYRaQmYSQJlN1RXCMME1zZTw9+01wJQ2Zc
Br4p4nuFbIECD2rnl83fpMsmwE7fUkozYlvsVHsA1agF4VUXTh7INGXIgIPRkfKZDy+zK5VmqNnw
aYUm/BzIqEeAiWo/9baYHPooFfRHdKStvqBFdi46YPY12+6COa+gGLPgRP8BSDCm5eM3wlNfezF6
dJuJRVPNdOnAWi4gE9ycaf4ev3Sf2+pMaP1yCvqVFXrD43R6l36FmUNCE6t4aBlvPvSE3gnT6kyr
rzeXUUMYYF/fYu9Ec5oRD3I8W1uQrRtuCTLiXI6G3JvbA9FP4Mrqk2KbXzh+gJ2yXG0CGgGHp+rb
EEJ6pCJKqPePsTZDQsDGsNuug039fcDTI1O8M6COSaSxlMwQ3dzJIrTwm9fVuYEuR7Q/QDWJXFnk
0kRMWOar3sEZFihfIrJrJacnsVNxb6PpnJCETsoxAtbhqoslMOVuHjYVuTJdm3yzN5I69GOiNzRL
5dCNIJaWytxqUuCO16t0AGyZ32nM6MdVh2BBD4ha0szM1vABQ7WeOgEH6KAlX1JUba2RPeQFPn5A
XCGODW/FTI+jx/0TLpQKPK224f5nsj2cVp3Y3okoXEJ3L1327IhG5dDp/O8+HnSKAZM9EAXdk5DR
e9XOwXoma7jT52639rvTlBQJy0UZTUr1I3BumM2unJnJylRudzxQxcfXEUmOkKKWN8ivitJxRsdk
kl3BviS+gc9q9IdgmPOrP+McfxQ2yKLERSyfrnj7Y2JMJPp4RjoeFOsWsQO51VamNZMug5s1xBSB
x2RAgndmqQVeWOdjVCI4O/XUaJW8GPYQlCEai0hEnsnUnqLwNhsGO+Cqeo+TtVuPczbMn75ViEgq
uNYIKkOemcd8JOmfAb5zXDs7zt2Lke4+KOe+RHgmsAzMclUS9hLhBj7e7hRahboecItDXbHG75OP
u84/LaYbGZJfNSWln4ZXCnbTDrDXm8LwjqvkyMIC56ImNVfWs5vDN91sSAsXwgF/meANuN2dzVz7
VKXZiDnhRULfvGw5ok7IvjwQH9HPjrWcSdSO9VCTup5aCc2n9MAEeP990x06RRf8qSYUj8nmnWLl
Xv5txrLQV5o4T3tJcCYP4gW9GjlI2On+TZLa66cFz8Spi+gg/A3Mfvp/HZR7blj71o0mfG2Yrm0g
kF+RuQLaw7xO4Jt46ApT6x1YewRSwJhvedxxUNZi2sYYHcIzHW6peUecB4xb+wFDvRkE8O89Euz3
SJCMql7eHENbzCmJ7ZKi83efba1wInHbyAdSeKjMLpG6/eetJBfPcVIBL8AnsU0f5K7JXtqOjMfc
7jGpGZvOl0o0O3CHVEmP5KF+qABcHht4R9JDAphIN/mrO8X7dkvu0QKaDJlfKGjWbyctswPYAjGQ
eUZRpokcaZPzEJ/XTZ352Acj1EowiQEzyaE2lGzDShL0+ivIm3+zW1JBRfXMwVXF8Muw97RBrvnV
3Ej1GTHnGLDqh2CsXLz6iNKJLARWOiL2zhR8v1SuFbXiB+o6LOAnG5y6rq0Ag0wInSVC6s2dbFGx
ZTk0ljBR38VZM+XUQrXAUhdXVbEsBQtDKkC6ZfNA5CDq1Qa77qtO+8O2DWmDyKMaUuNZsl5SdBG0
dz61SRYyugkMlvfp+ZD1QEktt2BjhMMIy7+2wMzCuC2uWhqezFz2HRR+f4mctUkBK9vzqABT9Oq3
QKfLMvR0dZKq02KuQzUEaLdHmPtc96xNfmdNhLDtiXoubUaQCGRwIiqLObsv2Zen+Qbw6PH0kCzg
H7bV7NXiR+VJZ9gQUDVwSujAy+8xZzlWopps34XHsT0pYMKm5Co+z0Q59UJ8ivgrhcxW1jK748Q4
xqSXpD2UAr0bOIPnY2HR1SedYN/N1x8FV+eY2M5cwY1jMmqkjQdzBiX9OuqjIsDS46S0iuC0Kfay
u9JhRPtX9UfBDOtmbj+VCgdiYg4443DP2p+jeOQwUbwVbV1cBPu/fiCi/z+daTPYWlvcZOg8LvmC
NOqIn+xyPpzLJpZtduwZ8z7PwdqmSR+uL1vR89HXCQaCiYLxrrkf7m+uK6Cdpg7HzFwxi+1lbhpT
myI/WR3tXJ5FGs/ZO0MUnwcEOSr8DNeKQNDJaO23QX2ZPXZZtpCDu06aoX4BIG2NWnqXXGa9INO9
BA4+5RBLKu414Kbp1E6+NMa6jtjfg4PAxOP5WGaeoTpEXf9+/mxnu6Xh3TJ46itrU1FBZ1eoIK+a
DN2U1+6m7xLqPs9y0ztVAIsEYUj/X1IQaMAhuomItCx5q3Vz2+m7RQqHZSdy0PQCP5aIks0u4NIl
Zv7+kyVK8Y/ZHrVrG1bDWo5jj0N77JM62RBoA+FJ38ykbd+VCZWRxx3lCDeJk9ksI5zO1rSHwdIE
iJ90ptp0oKc9seaL9yGNhq5YpvAaDtTL5ehRaWejbAJOM5gZyFSJ/UIe6MhBTI2VlQIE9eZoXkOl
pVvSQ70AjYsA62Hq/o9/Idi0cld9929fyMt/g7RqGUJ1NpH/79pwJadhudsJsOe5IkiPifBweLz0
iyUrhnTHi0pQeJk9Jsw0OIZi6zYs8mFdGfg6Q5XnGW/jo8c8g1wREv4lKmhsnOuumCF1RfXTfZ0n
b2wPeQ1HWEdSXlGZPL7TSm4YXAJkQN+44UBDbCzIT2vrVdQVglPhSoI0fKilnDGDSRCFGZqFvC64
V1k102a9X7QVEm3cuiTfAmaKpEr/S+m4PSMrjoRLlX+7CnpidZmJHmK73PcmCDmY115qDTu7sFS0
BZVoaGJZZDS2u3oftgK/BQL4EOFc/zWFliEPdhyJmcODv7ddf5vTkbkkhCnTd5LDNxOFAyh50+YL
KEkjRPx5kw7lJBe+xFvZMoe2KfVR8YW0qx/ZMQkEUjUStxsBeG0IyJDq+6dysYp0Ufr2hxoLVW5C
Qcq+1d/SOf6nw7S/UPsPaOqX42KI6DKJDFYKNj+XsSn4tDHUwxeQ1FvvFj+8s+vwAZBu7uOwbI5G
VkPeTaKx0rjBPiCJiWJDFc6BRAT6fRDDyLr/BMMyE3h2c3tD4Lxcmw8sxl8wgP608HSKj9nnbiEj
zzrcTsyvFHPoOVRwcfToKfFwHZzTe0cOlrleTg1vvqWEJmHhQhRE2GnIZi3L59woUFNQ0opVZszE
pQ4piBpe88FG9KgoX/uGl5AhCHKfylYjFw2eJl+6gNi4cxr3x88588as80rtb8ZNreQPAcN+z3kO
X8Fvubm7bXbso3RRsAaxnKLLiXzFuwMQSYudj4xm9YUB1o81szHI4wzT+Lnosr2me9dFpnYbgFv4
BR/F5LMy6RaYYuoSByg8iEGiecBhwtWMCEVhIYfcMNOVapMwE4JA/gRMGb7Fev75YHaJ64iEn0pf
E0+kS3Vr8+yL8wfoakVePFnFWEynQwY6ywKcxWuP0Sj7FpXuHd6UsO2w8jAw4B+kYjelcUgfRpom
JNSiet6PYmENp3NXUbIE2/OXr6m84TXalwkhprocjMJm/uja5JGyXQTKd79zwHsa1Z4WHGMf47zL
twFThGG1H8MSmvuaWFUxLQVsAPYJeSJnBhCARz3tcdCg9jVwZM2Rs4e3qp6hOWCCeWxnT5YwFBIl
cetp3XdlHbh8b6fvAvrG1oPCWEBrXVLULTlILoHT6UJIiByjqoYdq4ggtbMQ6itDwEpqissDU8V+
6UYWPmuTGPjGOQVcCR4Y1hT8eNUwUHtVDrENvh9AsBBgEfb7f4zQZxvh3YSdJ7lQ3SWi5GReyd7e
CnqdjDUH+v/ARHHV1EoQoyX+NIX5160EYuJ7S1ym+3N401KKEvNejbTveiWDMNHO+Yl5OTa1NMvp
yb4RXLfFCP5RJovhx3BHZNFmOICdN8PyHsYeYxkdmkp91c+hgyCZyHivSj3z6pB9hLE/J9BVbjOI
ZlWOMRNTp+DBXPEnTX4JrbPq3/yK2SdpY/JZGRp4eU1UoobNmBxKtXV2sZHiD6MRit3D79ylA+Ad
qOrM2jYgdORB7RGgKzaN4ByjLnU5aHFSWa4R7alFoJCP8aV6O+bIPSyQHPuO6GPQSq1pGkH3sgBA
xinO24CV2u7n2Ozcj8WEOy5SqDSwNI7GEiChOebTbc2x/NEi3vEd8d/GMgHbN6iZWrJKeY9rjG96
8O19yoH/WY+K3lQQzYerH/TDJRoSZ69B7gDUHoRAl6wwpDk6nJCM3iB4eSs+Hb4Ckbcrk+oPBXGh
xAI8Yro2e3LkzNyyUt9x4kB1z0swBOnNXVN+F6lNRub3+AmAl3F9SO9Gp5gFb5EyTuFfMmdI5hxh
hdnMeBugN2x5gqoYhC9liqMBuVaoxeag9hzM/8VyCWtHOMW7yuZ9sparybMucDishEiAJRnriWAd
gxxl454qk0O2db1XKgMnIPAY6DiLGW9M7ZAgXagVIZsIYk3Doy1s/MHGhFif6V0K6C7Ss2PKMzPo
4Ubrs5Z3Kz23VHN6WYtwYwP9Q8oeEfQp121ecXWicMiPMz3fQldaOrYX6GqfNVxFyCEpebw7nVI6
ZPeNVUChLab6Og/dF3U2OAeCTLQU3UYt2tZOkC0bS/86iKSruQZuaod6Yo2uHBgGBFVA6K3VGgIh
eFM6C5fU44gXmV1nCFhYsrDXWsomzldGHSKAwBixOdUlnRn068Rzit9T9ta6fKq6rWNpY/QmLv2x
Zx0FLpFkFQ8KY7X3rg/Mn+c0heBeCNjfA1lEco1CpUjFFcBfNvV7Ckvwgm579IhROPZq7H+KJYAf
DVENJImrAKKhVCs0DE6FLOSNg1um5wi8d6oeVLSRDsVuiVZ3qXfq9JksvWFGDOPP4/O4XW/sUGFy
YnBC8Ixg0pzOkvtxAHhm6oe1XRFd1gxn+4nhpm9RhwzLWHeNsQWmiijT1gNwTbqgInkADQxqB5S4
UMKO2ePsJf/NO7BEnojsvqHd9YKOeCTfEG1E75bIzpZN7fef9WBPm2GamNfKaoMMqOL9nWc6hKD+
Fa4NSbtvT4c8D8JyVhNf9LzdCNk8apWycQGIDJH2vWPPm+K30qH4B4e1zMiO2SwcSZaSo9evxvZO
9yMaI5QSShzOk3B9Lf2mJmZjQaRJakTQYFhAhrcRkOwDmoKWepGAA40ze8KeAzaXckb0sAhHMifA
+Aj4u0uJivje9PPf+sKMVa91VyXbJjdBCvl/19e4OqFuS+r9lTSK13s9180zaip9/3NAFkDwsVX9
4TF5Qryj2o2vuV9Rvi1ESAW6rdlPBvtVcJOq1o2FTbhb+MBm8AKP3dkNjoIWpFWvXaxgRPga35+D
ecHIxcIVAdTS3L2SphKa0kHtrsvqskd/s2plZV9B9A8J8a+9FAhUWE8BREvT4yheGQdtZB+G1Set
WhNss9OT4Kef77scJsD1rRCYB8WgfhiNqXhtQdnP/lm0NNUdZJQbRhNkd/CoKSg9R7FB309cErmY
dnafqD+Qk5Pmn472Rnzt/ZbXSSz/58TJ+xDQyVtTqBxM8bIcKyiLoJ09gmrrrVUZ4qtedOzM0fOH
/RKIru1fTvXUrj4GmQeY5BIZ60gDMlm6N3VLZJfCmIzfKDLFkDbJH+JJwtitT5ugxQ4qKWBi0Ehg
ZWRS+eEJiFXbyhiL1WtuN+kWBzybAOON+yzFD28BmoxtqVBh9GGQGgTGFOE2pZbF8cHqM1KXcPOg
dvX4HtBHkmCqjQhElzll44+ee6JgsBsIhDMqF/kXxy+id6BhQYSAEdNNqTKf7rTro1jj5XAY7gtV
XEqt4coY5KoSgAN1qE4CvqlROqQSBH/TDaiRLwV+CVRlwSqL0YYZbuafa1rz9YsapZNuRSziNiWQ
P1lwe1GEYWJp6SKCGYGy4W7i3sGJzVLyk+h0Qy+FF4Z499O/KoXTFMwyImATtVh8h1g1pJLWEELr
U413beAyYaI212jbLM+Dn3ozkIedeGg0YpK5o1QmgAAcYUknYIJX6km9LhjJ/h3+7ao4WgLxp/jd
GKvEdm6KvxLDAuEOx4C/rV9OCryyHlOsaL0tI1VYwHAEcG6phr2kPHj0K7r6Ih//X00IV0oen3Hh
XT4TMVoD2+w9pxSb9rqanhk4z0Uc8IP97tlc3n6hebdRncMT/vT0+gBjeLBY4c22HJBV1srJYoSf
PlrH4zAiXTmvtA1PQ5iWCVj/xn6i4EsjEbadafttMrR/mtb/BlCvtSUE69gRfGYue6sm5VjS4ijm
4XZlEktnfzNBjB7i4GOgq1Uit6mj7RUBbNXifYnSVNgNMOw7nbh6GUgki9q07L43VPF9cp5vRJ6d
Gae109F1CnsWnN505HPRsdDNeH5nfmjmUarXSsP66vvYMRDvnslkB0KJwjDtNmP9vm1EHzDYrnEN
9i8rcKvCXVTnmMRA4k7D8DJ5uKyrg0ftOvtgugYFgbime6ezHCuJvYtjuc7bfpV1OLPHtb8PRPr1
4wT0jlCaqyUdLSbT8HINmdUK+EMI+wvomUcVsuepBVKmE9srZXo3Y34xhv/oeTNNF50ExCew8bVM
lnrL59cVRVZMmb5Goyeae0NcUrEch0sjl8xv9XwkR4LB7jfDN2BMDZteCJ1qyoU7b1fESLRk2dBb
miwjWcJPFm8EIm+ZHI0SNh9HRZaeLt43gR65o2qGrTg7/PrbGubqFWi6EEW8GbXHp3CGxXTUM5Lz
UC2ad88zqtXEd/9Vkom40NBrZGMZTROUlSrmb6AYFtSaAeTW1qTE/rO3M6nw8blz+YpuZRff6a9I
z2OeFOz1rkB56w0Df8BO3BHIY2V/xZN3ilIxx8MRO1Ka94Jmi/atlCQy0FReLfwh1bTtLO4wAwCQ
nZ1U7kWQ/Ts1TB+H6nMIXyi4eUS0cT5545Pd4S73bN4CEFgk/DV28JdSIsN923enblHaAx3yVRFO
5LcxRU6qzQP14OiHbreOEHY7vPdvgeOwyBsxpvr0YH7kpZaTIiIgl8WCF8FL9o7Hmbt0sJUKnsmN
CizAeaYVGU8PgOMTWdSVQNe5xSnF7iPnS8V9Nzgf/OsSMkKbMj5ed1vCa8TIlDIaqtabeoWpxn/a
1fjEVz/pep+nSXie9sdcOaTVtamjHSXS9bQhRJqZ96zz+F7XdHqYwGKp66aGyMr+lKqILpOLb2xq
ovrxDyR9bUAeP06Tt8znoqJXVLc6sC7pnuzoboE2x0SxWA5iWZllvnOE9lYBzZdVse5rfPrzLSYW
G1wILXi46+WLBbz1k+/Rd7Hj7gx+ok9aquljWPMxiLoiDFPo9Z0YNAbXOFl7sXR3N33HEi+avLTH
2GfEESfg3Z3g1sgLuUgBLKPq75SWYr77YUUO+x3Huu7U0PCTMQJEEEEYoQROolRAwVZls8ziSNPy
k8zYoevqE6T96NBmcjcjuVXAPFDrMeJ0aAZ0gN41m3dJcuE9UfwU+ZAgcAQhaWPukVTAl4X2X8FB
1bd5WLfaiArnYSRFxPwqm5X591Ucloh/f1F8i3d18O7GGwJKrjbQSR0/vRuliqR0Inztr/KkQ0Zk
Io0x1t+dlEdQUpP4urpjAG4jPWlINCasJNH8z3hZMeqe/pw9jWRiUgSJ+T1gQ1IkL82EQXDtV10O
fgfSa9Uus4NF6tO83s7Lde/SR1V7UO1VY/U8uCMBtQY4+uZkCVuBd0uC2gnSIu6gO0mmR4EyK+6z
6zD7aRtMEPZk7X+MPCp4Ezjy5phq9YvY6vpaDwRfQHcOB1KZBKY2w6CcBzh4H2MrPLUEuoBBzJeb
YhclnbTLsXfGnX7xOoWdvDg0Ez939LRviqlVfF6F0xcNY/Q3kdwQgA8k24f08GmzHU8Vt8xNocZo
4Fk03q8P/vyr9mjTJY9/tQy9IvPvN4iR942VgzU0tRXqpTGCKIjJFfNGU6kr8UCroxwF4xxHtTv1
km2Lyw8OVV2USSyVVPXQgVjnQPBrNATAfGyorCyyl0DRRA+I/ark8ZuRrJQrYmdo0yN8R3SDKgFk
mNIOYNmInc2FXItO5WF0hSntQMNETLo2j7WiuFxrw3QMetLaYJgvJfw75gM2JrTf9R7EyEjyq9kp
TDKZXiXBGS1Spu1RMbyMqr6BFgnzd+x2b9I1mTiu3n7vyIfoGhnI/OODpsdC4YvhzzA/kkegkvc6
WRw1QJXZALMg4rGk4tGpGXNgUThuYAoN9wTu7P8KrDnlK+IH4pSzfig+lrfUOEXT20KQGrycGt+E
A6yTSCFB8mW0RE1T74FgkvJB01eSy5mbe3rNF9Eeu69IkJe15nPAvdXqxY784IVPdA3lFATGEvHT
nxhj8Czp8lbnOnHAqdGCDyATCHhqSePh7g/Sij6nQduAPn1NOHRcIMRLU2ctjbrVKQ4OYeC39d4k
lZMOA9g55gZdDqy09GEOm4+AzN4BCy9p2U5iVq9Q84fhZOrV4bGDP00qqsi4MTBD0RlMCvbCIli+
6Bw3e6iqLg5WsOegaj5JaLLBIXxNf6lRDlr3pdoHyFGWUABQ0CQQrUEndP3WFlblsmDCrM6lx2rR
/x5tEdz2L+F8e+vq5vwaRpuqkBAjhOOg4E1vQ6qNrqP0F00cpf1jPiHAYPAdvIoRO0JTvcrnwmNM
heAh2/brnuoAxgY8QYi7Werb+bjDqe1FaVJ1Ujt9cIyXXlWeJd1bUoNZSgi16K12eakbNDoQN2vu
eGkRdsnnzgnN5JGr4wcMnJQ//2HBo1b7ViXBk/osd1MHLG5VREu8x57Z+mw+0A1majuIl4ajBFfj
LfTNNpNF4cS44WluMoyNlVfvjlkhgN0ztc4zb0YwCSYDyoQTPtR3xaUEVd58/KKJvOgrqj98GQOX
k4YwL0u4vSu0YQh8YD83Uyu/eVn0p1Do/+y0qWi3PZRnAHk6rm6g2/EurI+GeBLPTX4F3srHqQ1X
4fNEw1CmDmsBydNrFrynktnYItpXaPn1AhhyMSMPAhQ4XL48yH3rOdGTW/5G6EpEsKTl9JUqIqoU
aHq7AuCLfpfdOdoNjU8RMMp2v3DGDdbaED7PPLUD2ovpD6bchkbBLWaiAIc5PiAbleypVrne8oQY
nVD3Nioo3rfUjZpD0J+W5wTRgFPkbnx5dtb+zJczZgoSz4zboCUYvN1pzBRbjPb5UwyBQYYwL4JW
PMIWTUC+tQnQD/5I9z5mYDjk/q4WrTqCMHFMqDRTkpJhD52e1MuctkPyS+L6yt9pdUAWGfFhgjO2
Kth0VeO6fXV4l+T9i3cqzeCBUM850+nJ+kQAouZPXOr4s8UyvK6p/R/3E4dCj80p0jnjr3iv0LNH
zYHehSSDfdWFlIEQb5w48ElxS38JVXVzEL4ZRBqE9P4QCTnyiqviTS3kZl13br4dAOv7BjBPSRlL
vXIUyx/syiDg1kSVrgQEAQE0gtxI2PSL/iGJ8UJ48uNd3Pxg3sJYHkm8OB/WbugVE5g/0KpBAVxs
FHyps7Zqm5da5zY5Vl8YVVAzdvn4F0LjBBRnf8M4XW2Qvd8hriGzIjzgYiYB4Ll4+cuWXztos75r
ZutbblSDJpwGKAxVUL1mJCDTs0JiYDE/337WdIpRxLmPd7x0RyRta1tuespc7+C+4gkdviiJI8MW
OwXpr0t+McsbYRUoc6xEM6kJ0ak1o+t9m14oXRUXtLqKwFqA6U1/IrZZCGpbRem+vMaDpqOEB6dB
9a591wYlb3p8GIDhVPr5zCgQF/gPT4jp20ecTuIM0zsJczfCokokCLD6sDlS1mvsTms1ieme7Mz/
iDu6vUW5LRqQPoOpTwQf+yuG9GtiEI9vPOGYzQyZIY9nA9L6eZbcPPbS+WL1mILjLzEs46mADQ0y
MvyPilCEALfnHH/dA96GsOK1VUhmtJxm1eGDCPmLSY/ysJpBeU9CEPrJEMzexxb739mGLpDTvrZj
Vs3T4Vi+cii+MRjx6iTioccDysAKBS2jjZ6C26aP+TWk6DDKMrcUd0PA8HWNo+2BFhmuOPkDweiE
Yxj934V/pz0Jb2uuB5YY1nn0FqcKEN0BWJcmaftHuwpvlDZM7UBSZ3wJ7MF3Mco7wVmMs/fkHz/Q
d7M1FlwybKvwUMQLtxInhCh8X0ATy0DyRM3fEk9X5S8qOr9mjVJuc3ThuHfi471X9Jdy9wXMuiIs
R6HMACaSqDn2rDufD4K8VQlnBUy7DiJbWyUI4uIQ+RIz7BsD67LSopr32CDagH0coq5+R8VJ6rYb
/4n42BKi3/7s3lbPIWEZV7jxeS6SVv4tJdht3ocLNffEqpq1SQikskhQj+wjcLr+OH0zf++aGM3P
bsvP8Plvu4VgZLk3kBFIikv2srVlVyCCiuQaW2uKrSAl1FuZqesOB76DVrzcd0CkMHXpgadhkHm/
iPLChyA62Ai2Su4qnR4ThSYLbT7We67p9Gi5IVMkYy6S5l/UWgm9PnLN8KLHtpWPi6b48uf6s5o2
YfD/dLjViP1WOZaxvoaOz5BPKA12rEG7+0pSbxPBgZ1t+ALEqZNrr10YPVSXclMu/Wk07/anFAqe
gKYjCfqNtImeQ1vConpgJdEtWv6RisJrbUE3DVJr6gos9W1msHlUeLfSB2Zoeoltu2ZeJlFB7ROK
LF1xOvPJ3uvxGkauh86NZGPRD7vDCRmOqYJ5YL5T3P+D80RDmcilMrc0Jb3rrODjJoAOJzTbvwiv
E28kOPw3vWHbPtCIsNANI8z3+M6guUXP3T8Dl1/Rp/DpzDe+Bu+d/jk3pHoyGB57LRkljuI1i34X
i6FbL4F5SxgKdV4vCjztZ3vU5brGG8Bf+pDOfxozUGLF24OjSI4grbL/1gevS03hRiI33kPyKz0y
z8QMRk7PUMybf6DLYqMv5QACRSkT0wL9zCMS0FAVQS7lIqBWADGYf+gdNzUddzPbaz6JToetaqq/
PMHKq6Vjhc4ySy4HlisfC/EuG4Q3zGrBdvlRM1QPkTLYEsFMGKwCobVTGhbnG30IcEAp+jRzCRsu
63cdDahnQjbiNnmqQ8Iy/UE25tQ9MnyOKobJjoGA3igaqHozFfOh56CXCwBBqsGShfUu65dguDmc
8GgiPFlcqowK8fu/BPYRe20y0T4On58seTSoChwKNY4Oot7tckWeQkXJAvvUg4xgWiHipUJD57Yi
MlEwMyiPOftVPEekq1NFH+Bd0ukCJIabd3WkbxqwAk0wqfL5rXFnNKtzoGHU7S+NH9r/wXw7Hkit
kl9Q+PuR54tmJFcKcMCOeEI8wFIR8yWnLC9Jdc/re4Oqzl7B11XGpbiajWnQXgX37ygG9oN55SYX
jBdzlzXgp2RwOHIzrnihylV5+6FfMjE9dGyGUYmJH5soOKn2OUCw7PU1vrie4/nliU76DrYQ1cbI
qL/BeZTgIDzVGVlc2xpYuIfQdD37yW4Q33MfdoFDvAPiVVM7+CcsMBvh/g99i0EYh6OUuCV0Isg9
wlKi80En2Y+wuJ2dRlNCpybPresJSGlq2j1SJXVtFR3O5ulOWK0wwUivaQU4nKHrgdYEKzJ/KtUW
wR4GR0Ra/4ZZMZgD3H3zQrnHvvRPLzBCZ6h8dGw1kZFUOARNhBbVnGzJBui+eZNUoBXdtpMT4qcf
HwzbasYX7Wk5WtVoxaQeHpuESB9E/o3m/CjUkq9aGPzXFW0tSdZqzemO8bIldWyNLom9YkorgUyW
0nsm6IX3P9gZFGBA/DstMgfbOSNJVMUUsI5hvbL6IOpT42Y0TRq3OPtx3vNbISmwIi9hZsqHOcjk
oBoceMn5S2weO/zeZX/0n2/W70lFrRgWgQRk+dWGTcG+o6wAmYVGKlM0Ax46yiK6bNE80noiWhAx
MrDjvDvLieLdsqPBRTXU5y3CM8wz/REllGz9DcTrgb6xgO6iG08oicBoUDCRB0jK/bhYTFzUpBK9
iMw2u/NbgeIAfT0CrPNczf2uRQzdFZIJlAk+hRp7RrXwtI1HXr3EJFFJQdBxgixppKPszQZhraD2
eSap6hP69rfVgdAjhHMKG+5f1R6rmqIVVm6/+4gtfCOxao9E9FQwWCh21dLJd9rksNqk/gP4IpzO
xLidv0HmFZZtnbpgvTWdCvIr4gLF9KUVu1DWjqzGiNKJYOxI57LRbCdLc+ahKP+qLMOUunHhecv1
NNK9p8ZzMxVZ1t8tCtBUAtbKflat5mgXAFPahPOREM+q/xylmH1yczJC0RrC4ikzsrC+yhtx2WjC
ylvLvDM8EeFObv88aLQwYUGYTeAkf9w47iChojlEixEBbo2zgz/2XC28H8Bwc3p1v8J7tYbnRCkM
MFPmQbABvxqcvRfCGQf9ezW1QlaNky4Jx38gwm8enSe2N5oRuwTZMucK6x/EvSQ/XwtRP4rdTr/J
KnMD6urinRxfUsJxiQy0DghJ3Aj/AzaluhPNQJ/R8JYv+rCQ+jvUaEhDGljc/gPi+K93XyI+KJuj
9p7r314A4P+B8XgE6GWxIjX4rap2AqBYeTbx9RVmchi9sLnRBEmfNBlYjFJ4lo7V3ToxnHHbDcdX
IH2QqTL/auYNra6NQrx5s1M+dOaFFem62qhC11HP0clUOjrVrPuo5iYBmVfsJ8eE7W/QjjbwLMV1
5RtzqAaDvleNHRx1ICR0TcvIVhMN1ZqRgjTO6tx5WA7yvdq/RPnUnNnFTNOFSEe2trSUd+jF+TEv
MDixF/VdO+fKTQVRgr3Jo1NqKueXbfPZ0UF4zjpt/inXKSqHvB4pcsIiIEkVwcDlXYcb63g5sYi5
ajIal2sbmA1Sfhw1+v0gzVwcFJ7bVxiIXgh6SiDbQaND63IaoiByt/QnA6+l/D6sroSSGzzx95xC
e+Pzsm+7kZOwk2PD49q4LWrQtz0u3HLPOC8lKGzCskjcLewHSrBQjB9omw87Bj/Q3/8iNlkQtqMZ
uMjp4AW5GFMweCCS9NwZJmuBs96ACZ8Gcp0PLnJJTR4rXBypht1+cWKLGBqOuVGz61icw+MGZEWc
AYUQBL/QjHPG+kLhxSuHPExAfrBeaj/pk/X0Xj+FdDirzJL6CRw+IqU8ErJR8nj62X98N7XIXh1c
R1uO94rHpPDYNqR6SPMQ+MYC+WaxbkAi9JdSnP1EWtjUKI5eKaojExfFqHCrJ9dmtKSB3HDGA27e
hXa25/KgccXjghACvzDsEJuL+KDrxTkOzGvl+mYWqVH//xypD7jLrKe9hR7q1PKULq4OMOh3JKiY
acjQW8uascCH3MBWG9es+Eamf+phH0mBkvYQQdsKl8TfNRioj4QB2L4guzWhHFuBvha3dH+K6iFI
d9YOqJXlvoIxxkODctIo77O4oQBxxfnLerA26iJM6967ZD7sYB64BSkdQmjyRhGePKWoQpdm1nnP
u/lU5NgVeLVrAf/gUMV/4OFKQ8LIr87TUqtv0oug+0dpqT9tEKEkgeo1Vdmv7Uu7OPoZVx0iAfiH
WD0SAgMVGvkmWLhKd441QHfsj1qsGS7Zs56V8V91z3FYAGzDhGRZVJGxqhiqZH1w1wgO5NADurVM
QnoGWT2buwhhBVecegRekeiEU/VHWcBQJ62y+duMVKAcaQ/a2j3oDzB0nu+dTyj2Z1tBHn9wVUGf
x1Ocswmcj2zzVJO4/ivDSA2l59gfF7xyzRQFTDIbokx8Ej0Mpq7C8iG66E+kyqz3Hpn/djUUme57
ZEzzLm4grCMrC/jUz46vhfoLxO9/Rk3cBDQCFTuUGaMyhqt3GLkjvt4+0AckVdQKzJM/GlvngouU
kD1dZjW4p+EcO0+zJ04LGOWU3zOEKBTZXcaGAL+lXI+OVT397yDNcsxgco1JWpOCKAnBbAy5QxTz
LkS3tJ4dtPJEOk9JvS78RdNTXR3HusmdO9d75VL+ttsQH0HAuQxhs0ldaIgYR1pYSkwSW+ZyHQFv
MDVwITe/HJMEvNHF6SCB51RMen7b7VPFO98FVTrfmLontfer5liRSPsCCAancacqi3KkirwCMO1/
R0P8sqDI+WjtxR4DlfnW1lAzplIwwcK/JmTuZuR+a1/FDVAU3EZAsKA29GmeRaFl8dtcUqvEwEwD
+2zTE3mw7m5cB80FbmGPp9XURrxO44n+CD4S4N7KccAoGIhJjrj5Dfb7Oq9w74Mp1SJ/vNtAXTjs
3i8xPxq38VvxuPjWixeljmTkVi0UsgUy3QBFnFF3pi3ggnKAeXFmHzCVqP0G3LailWpmYpy2c+yB
BSHVszX/j54i6z4UBwdYPX+vS6HyJlvEbybmsLzAf4yobzqOJBtolFQMia/QOHuJsTKIQjRyKfOE
NUmb7/eqq6Vw9I8dBek+trYHtyBmZBDNE/KUd9U5tNdP0jNahFAdkXDimV0iWKCMKmKP+m4xSDXN
wP2OJYgIGYw2s8ofY7w1dfHDycJDJnjqRfR2gk3MPQiIRn4jMExUyDJ8vwhWd4/AiPJKWgdkxQu7
K5tEE/fh9jDPeouePfzXOqLr3QqvgVbEjkzcRlTLUPrYUMBCaC6aJGcl88zEw6UF4cnIPmHSZQ6F
OMxWXw4c8SG2nrSfQfZMsvPgU+A5Z1PioCnruFwSIKvkzMQveNclTlnuHesF8HKXCC0jHflXbXvo
j3f9b+9a/vJPxR2K9tXU+lbN6GgIcoZeKKmlIc/aaGZNgaFIsLpmrU95v26i/f3edAu5a7CPpqJO
SZNiSup4n9Cnu1Qcp6UhfJ7g7eZMJoBMvWOgObi5lcHWli1dFx5KfrKsoUBkp+K8u3ZJotG+6YBe
mjo2JoMFYxijiXO9F/8z8KkZz+HEsRWAOlN03ZGTua/AuMC9W6OL7Wehimg7sycrbissf0/Q6tUn
+dbfmczHPK4Cbvlh6KZ42wPIwVHE7IIUkzcnGRqhxUiDiY4ivoU14GiZaNj7UsRKRqDWuqIbpOte
E6MG57cV92swl0U/ayU98NQUvakEeEMGuii4Ok3feUmENnEr1PcAusGj+vWAa6C40sVOOfZcFS5y
zl45SDCb9oCcJDAyUI9FOqJxFpZiIo0gl7+FbFx65cUz7fe3Z65HlPX2PRj+NI5/8kjTJm241B/o
PqdlXBGj8fg8MzBac4DLyssTGrAb3P5pK/28iljcaKTtm9lmV50Ntnxx77/YQtzJnjJioZ8/WjRm
e+Vke4u8pOHczwUHpt3sDGta8DQIHnqMl7+h1WO07J/Hr+YNLqgrR4el8JkXABJUNHinXeyjIepj
TFulvePlTm8xlJ9qN7U5J3xueWicf+AzxNa8xjQeuDmVmJzvVQPi3S7yA0NzA+T3AbLD2Sp8jnYr
98feL3pArFOPw1CJMdEOWndwPdSpQXTJCtoHUfuTLd9G8uQAufk9+0MbQgdWUhLtPlbwyrcr9mSK
I2/E+hGajJP4vMWWsW2bXCBDJueArB7s+otbG4x6TDlN112f5Rp8Em8N+TYhrfQS4Vg+/Ku+UDA+
IWKZO4CIoBTvu7yYf62PlP0lztjhDYQKEfe+GW6BFr+DqV1wsQ1fzOBNlVlWvVYhGkREg+Ly22ne
f9bT1iVqEFzwN2DGZyESqK8S35mF9Fhdi6ZXeTD89hVNLr0TGc1TkaSQGMiuMs/Xi01OdMHHTMX3
/YvUvGPPLpTsDbQ61BSC5YAI/MZcIuZNY7axQzCIReFHLzypBry570xXGtEjwT3H2iY6ABWNWEuK
it2eLmiOZyo+aGc3VQep23uJKtfNXsXktTTUfXpduYhkH60CMrHNpyZfxqJaEUxA1DEBZXp3WYOH
G8Y5pIuj6GI12dRnwakREl09c1EcLxBHoJeb74ttaRRjWiNU8hGngKXPvbKRd7L+9+LSAXvJKAvz
D8fgebd+kearLSyj9ky1Y6SfrdnN9dFcthxttgcMo0i3P1X9vIkStDIR9C+Jm0V63gkys9fOi1Kv
uCCwOKv85xaTBFC3Rii84rvYjYx5qJ0APin2Ni2OXJhnARvh02fNMV1amVrElYwaSnbWNCfpVlTQ
7slF0Z4ty/H1QsNScADWMToXhThLU3+lNnqj1y9eQNoCHuxs6YY2GM4CfutqxDEZsSSrDv5vNyYk
nwq4YWV6+8HDeWC6mNmXOn9OpmeyQIBu9sI5dP2cipJfcW8aXGiIOFV/JpdGHFtck5ttWwjHtxgH
exC7p7n0OR42/Lwm0fQlPnIDEpr2OBarSMdkYl9HzV2D4YafG93lGxAQxcMeswgHJVGeZuyC8Z64
g9C+ikdBxiM3UYp0px62DlOZCMAqXe5J7YeAqOiW5/mOnRBCJ2+T9NPnq4PYXIfu81SgVLWn0omE
pz7IYKQ8It+AKmrLrTIdHNvCejzoH26x2P0dmUk4zt0S2vLhcEJNWk9hJCesX1i8nMTGZg38wr0s
+W7H3n1/6/cfKsKI7L50dY1b5zvnGPfrKoMVJBuEfJvndj/sRlcAO1gv1RzwaRJm38rNrx0TCkUk
p7z1zvYTnSj7NI0sujK/6kaXCCx7V+53CsJgKfpekVBU/l+/zElLOqmrX+uw26U0SJRIkYaIvH3V
fiNYjhxQQXKfkZx7G5X/LD2StMxYX3tVcMTfuuYg0zLA3W7xS3jSDmSnyca0YhZQ1vc0qyl+szJl
CjtMdt+npPZkFQVTWsiGcZeSXt/Egy9D5FEkGhxrZFaxzCqQxzzAifhiu2+w4qQQrI8DEKWcxUWp
nxj/cTc0trRfGFhxBfNnL/V9UYSq3SkNCU4WEw+rDRrPt8xB1jHOJ+r3MTv4POu5Q4C/TA/glibZ
OWM8+g/3MHtBFPTBp7Y3qqWBP/r6ocAGYq8Zoof6Lw4XQ6WzBYQRGtMDprBOIKVe7PHOKyHa4jqw
CyQZzufPek2mK+Fli2ODkQgLjPpRM07hCncYned3KSNCTvYQ1PSO62qax2NPOqsCI+M0krp0b2Qa
3zF6uWesFe6M20cDa5btFr/kooCzhP4QvoXDC5ni/Z59vM0joBd2BxyJ1RDxeqpi0BrIgeQKUyoj
m3jC1FTQQMHnownU5usVz+BGvT0S4jNwjHtArZrdU1tN6M02PCquXk/Uyor8rphQg/3D8FineYjS
8OtSjFH+VatdbBziH0DTBgd03o0UElUN3ZVvH4KhLmvSrXKg5Sc1/e7ZJGKdy75Q6hvJQ1LAwf/G
rhP3Uizu6M72zzPG6BSq/R3ZwSzMLBQ32MHXqk9UTsX2BnYRnNMkiePe8mEvH6VjTYM9XAlp2D2N
vb1x9ZPRfztk5ZsujxbSH/VpmOd5vg2luiUeFKh7dCZ6JHds8y/vhOA4QcI4rttrWXzDz6B7j5sH
TwE+S4rjoLHwCLXP+FM1GdUu7I3735Xv7mak+m543uXgIC2mKrp7YPaRTxJfDJVKULog4nyQT0Aw
31PfK2Su53cz/UUEZWujxzvVIA9qx1KJVd6r4XIxOMoLY/WnfQDPoDnSkztDiw8/4U4BHUMbcm3z
KDGFGlcpvgpzevob18qk0po74M0Gw/TV9lI13e4x5fmE1B+3kIt4MU/2ESHriyv2XZ8Cj+ZmmtbN
iE8GC4Azgej50qwOvgKU3x4EoVgNb6/RnAz7JwON5iNlJoLyWKE2eW9YdfR3EC1s7pz3nPItde8Q
4e+sOF4JfLJhxOOv44xtfCR2qmiCKBuHSStE3WC4mLRRMRNz3KwS92N/fi4nWKgx0/67GUFVlcPm
QCoEg7obpIl37JOF1R41dYrJN7UbCZXRFoVv0mpz+EMIkjs0l0m08BjIs4oVrqPNW3iJFOL8drJ6
9FUq5cxbyUjvRrLUqwVATQ3PvrLFJBzguvC4UhlO8dU9fRsVDNXAxRT09SBu8DsU+bA8z+NBZjVW
UAgTQfIKciYTm9Fpx3dmem+lgyHn7faeSQ67QcOmNLGodMJqTy3s5t5E6tZkwVMEzQhgI2sXd+2H
PyYctXH+tc0LJwKbN9hdMketGYCmzLFTKdILBsZhLzD9tvl4rVmuooV5QvM+yo8D6HF1lQn0pmSs
RHHFuZQ/OrLn8OmQpXzpRCw1rKWW3kR3BMrznWH05erMV1+SVv2q94lVNmHDGhtJ5gW5agLeV2lE
+CbUdtcJSQ74UYv6itwvtKQ79kC/Y0lKRRE4VL4EJK3nJ3JAQ09krmGAWq4ziN5P+KL6R9k/1UI8
e26DBpLAW17orhayav6C6mrNem5sPTcuU8mB+nE6ZzoPeWWW7AsIwmYRqPYm95JSI1TYNQqiv3E3
tgncsTAbEZZuYVY+vtw0uoEN9CiIf2lFLAaMS0GXRGwl/kgakUG3sy2nLls22Sbhk18ypEr3w8zm
qTreon+T/ZQn6/q+jrENY2GguZ83fA1eMb92mGVN7e5sjFw4toC0CMn9r/aBDp9VF5FA0n0Dcj/K
5bf7rxdmHB29NyKjYV45i8H0o1U65eyKsDOCoSdNyeVCwRAQmnSUrxjwEcQeAqSVn0ct8AjtrdQn
Yw9N+gf5Dy3NLjvACE0M0bCDGt04MWzHDtpE+AKIT9FwBZCBPhY9drj7N7ZvPyR7cZiDAx/ZJ5wx
tTb1jQlSjhuJtumRz63XwkBtyBj3226jfk6OpvNXxYobTq3Y4KRgIdT1j0UFoi/pbbq/ETtu6HfH
Is7EC6z0s16DjJLgYtmAGoFx8B4/mb6y/KFP5NAneqEJKCPBzx8OF6GRxrQvvnPi90uHStpXQxMK
HO2lV3lQl3LVIQTWva8OCHsno8ZGs3K52M23qeSF3uQprHhsxAj86XkU1aFsFheHpyg/IO91HEPD
wkQbHIIytw5E/TLAhIwKKXlUw99NaGKFNQktYmlxxZiND1FVG1lyzZ0mZSPNifhdvGKubN1qFf81
qOjZwlO7UUHSmnkcZaKOvY7UaPHBjNlh5oXbwvADp+e4UWiFmZdo1FSF9bsnsQvYSVq67HLMEsgF
kLyVgxIrgfiPO/kAoPVyX+4DW2p1E5CMJxL7VMoutUabXTLAbQriQPlI5CEQvkELSGo01W81iwn3
G/YB9ZiGKMgQbKDkyslyfCMo7r4t9TOIQo0YEdDxMJykZHKNM25eUNjoSw+QTwJCVXu+n/gbi6/f
oQV7YNPu5BWNC/EkjTJAE5Z1OukbHISKy80brDxtjFFRAlGi9WVIDcTYRwfS/kBfhoWL5C6di0zM
IRPr/p9mUJNvOIIk+pX0JYJiJUmQJ+hxttlOscP9K0o0dMxXe3rOZekvqhO3d3vZS93ev+CpvioB
4opJqLtYrpKSfogjOAIfSRCBhUzCFh/EH+Q3ni0+P95tgfO4w3miFCxUnfUWUewRXc2CqqvZ3tFJ
fo/Wlj/T6KB3MqDmQDqgvrc4dqz+D3ErkSY+w44oULMkXCPif42RZ0+Jie2LVtm5noyf1nJ/CFPb
O8CBRNNOJsu5ku5W/MsV354dQCxlg1cBK8HYoUsXoTioYS1k8kYgIjMFzejP/4HQWQtEZFuqY2hI
j9+GRnywqEEgJ8Bnmd+V7/yX9zG/Et8oTA1jyGC3X08FiSw1jpxaNTvmVoaM2HeGsWEIa8WV1XSm
naJ4au9MRoB2VHg+/HnIXD4zxGl2d8DSHy1MIeS9rOXeKa4pACQ38W0DyQPBwJZLaWJj1jEodpvG
JSmg3HmHReyKRAnhflT5auOslE+ULxpOjoUP0uOvY9z11TL6Xp0FAXA5zsrAdnwbkyhJ9K/DZuL7
7qIbc6Lbveyt1zxD/RkQbEzFabHtK0pCCGk1kJaw1sFPH8DsSquzIapytN+TUQJlUOcBI7AFKYg6
PFSY+HurrDGbpkihM6e4lcqzAjmtSso8YzmP/0vLdEZsdtH925b92ZMNUJ6YrRQ/LAK/mziSFN89
UFjXLi9gb4ttOCw1f1ImyieCjhm97gTev4PB5xncncDHjzeJN9C+lBesQq5N9vxJYRwNaerpD5d7
8f45wjkSimVEUCWHZ3YX56G8xNWQgrsc1/qE6ylNnx+tWM4/wOb6mJ42CQVYXq2GPmNnWzvumtFr
1/SSs9HHs/f9uvyaRH13AutVRKCX3hW9yE9Ai3geIgbUf2L++UAo2wMDinzPyvoZPpANZEIDdHvk
8Lnzn5q99pyndtlZJNUPY/KMn54BEHBzrd6tIv9Nkj3dX9ZDVGoT9K7Hp8drR4HGtyA1+dVyC9E/
N45EGwWx3pdhg5YjIz+Oe4imr8pD7FLo0TSqM9VdJl9etqGgS9ac0LCnSD82LmDik/0tikSQzGmw
JMadWcn24HNoIQjl+Cpg3RqlENkoock9hiGOhtUvrHmZofR3GirW7a7q3qqNZa84Fkr8ypltTbDL
uHJxOQ5Ky6Nnfo/Mruakp7DH1/7RaDMsNtR/qCcAJL6L4ivPOsmp1GIobn1kkNR6ZiO4R56tlnl+
sp4yag4LDYEueoE7Wxt0MvgSNVP6B2CklS56ja2uBUkBD43wW/AAwJI596HsgTSe1+XOuI1a6Smm
OKJc4FGIvpO8ZvPc2UhkziOmZnQJ6TQxNxa32kwpBoG4u58vq0qQ445tX2KaHd66XE6rOx469pSw
UHnRy5cQxk42plfGbXmyHDPxICAMLCuFg+SlqynFMRhx4N+LToM1mQnV3QlQ1JHUznSsEkkbw0LV
oq37eAAw8GT3uRVmdna/ti1Uj8BZoEWBPYT1772iebsjFlLmk72yvgMUpgIZbGMoY0DajCd3Pk/j
aMwcA9yrFnMQTiyPAxHX1eVMU1uqkIESYP9UBCmHd5iR6TxGQV0dKDMVYw8rkSiQpCeNrcoMN5ZQ
aaHdbps44VrWFVXRmMuSZxdIPyGDt/VsJVmtzoJ2ZhqvfJZUMrOaQzOn77LvNVN7IIZtN1aTouLx
EQHWce0yOnSPDjTU7TXoKpnWLF44b3oYn0nl8Mb75/Mb9CdsrEXRPN9ieFDn6NVtuylnrA1RJ18Q
ewd3+ws62KW1sdK6k89TVjI/OJA4Hvglr3mpxqVqbhmv6sKzGK9XHgStHbIEJ63bfbQAWD564Ltn
iv/aDO0cCkoD+aHlAkFFwmn074UDn7vI6Y1asxw3iXi43+xWHwOXjCmQLk6qJscNhcpFNGBdPrnp
oMxB1NNmmtWdlYoBUvHW7Nu2Vbx19377TFoRbZFbTdc2Yzh+fnmG7obB5qCSlbQ2PFFq1DRqZDZT
Sc8/N1Q///BZOJTsl1y8nv6q2o34n7SDHFvveqHn3tB2yhnCTuQ6eUCs79wcBgc81tzNavm9nt+C
ArqEpc8klhV/b5M90yBDZPqhwX433gFQ8u1R31MPqze08iD+AT+19ejPWvxdAhExE4wHYzxo9eNS
QEDxEWOZJL9vZ0Zl/M+OMN4/rXMLsxA4SNknm8NJ0CJBWRUDFDZ9kZ3xVe9ixRMI3DaalcYLLCOD
228Gw3u/6R+D9zbmjWloPjDsUjZYcTBxFjZpFRnaANMAWy8fpaCNn5kZBnvCPnKXY1ASq1GO21Ob
75+nmF/S2Z7bL7s8zN2CsmGxl6ysSLUuo4D83B4E+AvxYXOfAF0s32mP38hH1qJiPBk1itlZlgCl
KS5Tjolk1IB8fbbcaeFuXpyyaQS30VM/3Fxo1EIiqlvqdDlb4MGG9lDZ6+TU6Ca07ifWXMXfPH4G
ObvQn/IV71jXLLydFvjkgTSxhgK0L8A1hMndMH91tt5Yb9m/Ktx3ZtPRefPVzAusiYxRN6rJ8YbM
+Lmqu9Qvx6McA/T39jvqaUprG79lZcD3xE84nzEQ+J3Fqe4coDBpeVEgXpNu0kzn7Nhm4VLBI+B1
X5M1+3vJ1HcU4to1sQcvWm0b3GQ6/xxCs5JXTv9WKIiNPA4TXt/9yZbpZx9eg8G6wcg6LUHXI7Gf
h81WKUSPjDGuCpFQgw7aF7Vbgar6Zgp4z/8bdvQfKyzpn3c46Q6o+l1m39AQL0l1NHn6cLJpvkSv
r0EC9Joe+vWTGbg3a98kEm4kkNbKbYX/Vjyz/oUzaTz+bMURGYGt5kWzqc9zaZefsa2jWiO3mruY
VST/xpO+yk0N9PAOKE1HPMgg3k7qEAwo32iwh+4l4iywsvf9i71MngB4Jrw45fOd/8lkhHVDY5pG
l+xEhsNOoI1JjIzP190MEqH9RRPhvNT7pUAgfWO/a0CYbucdeRzAQyl0POSEW+M1q4k/UNHhcIAi
/L6xRiKVBkzXxIAU/El18Hqm3LOfSsds+zabGhCulTh6JKLGMBcUyL5Wtb6tZxM6vJWRlROQgrCY
ofjZumYBRP5z+Zrb9du5sxgmpkBIsOjn4GOahh8+Fb9GMKrpg569P074t/pk017+QHZZvyj09Kgg
pTsYFaoHEtWKQS47zJwVoLSEN6v8BhEyOGvHZ3Wa2Be8IS7BNwz841MM+U8tovRHG3vRxVnFqNXB
iG3QQJV8YxVPadYfQYZCmCNEyTRqD4uCkSZvq6PqMnbhBgs4tfRLTi4QuFLlwF5KUQqSc80ymE+j
Tc3DzmpAINzpD6a034thimXx1zCMxgNSGsE7RGbVxeudF9HTIWv6S/pQSKpGnPj3JD13EV56FQXk
z/8Zhh7vqalD1lewFEhNJXwMSdFLcPw6bhuLjPNu45dnqN69/raFk6PU9+U6qyHUrMfZ+5xYqnbu
DWVdRTWz6yBtfm52ZUrEBrwRcx1iIRnGpq4w90zIx3S6sTEYots5GpIGsyrfnSOGSVQQIEjQS1G1
J8DCVLp/YREqB8UIO7VS47ciQk/m4EOOOYZqqP1ZBF5wtsmtAUpWuRSg7v8lUCbnnesqpcYQtoTC
ftxjs/RNm9QQ9mtXbc2tyI0Drp6mwy7iU46AgAQe6+j9gOLY6dHPuEt9AFrKwjFHTgZ090rFvjyg
NhWFW4d3UqP1PpfsZlXvFnqSARtlvuteauLF6TFCTUWnl0iLclaczZWowMoJ2+yGisibdRIHkuiL
C0RNWNCeDlWGXaAbEmhJg3r+xXrY2L28GVdvrniTjXklNWWQBZO2K1pxExOesyREuqC9Ya7uJTtQ
SQOBTdysSUHN6mCNx0VQU82pDDWHXmbufzbun21DNHN2VeZXsrfyQNWmdRXdEoKYMSL5308nZGq5
7SMacoFR9kLMzVCqwqOepuqkZm6LJuZOiWA36MxND7Xx8/tKnsaPp1WlktpINTf2icC48mZu4Jhd
FIEJmRiU7m1+UuGOdNnP2FJ8QOCEbpkDaTzFxNWRUEAUh6N2NM0A5dgr+sfNaQ5TvEuymTpMTPv6
l6xQKKiyPu6JM0g3BxSPFxbJyM5l6pKA4yww0syBl8hH3t/DDHE7vmC5wxGjgs7kQVCejH/55h3q
mE8HqQ1dGYaNvVP+2LdjYvm7xP5fhiiRrTj4XfDGbLr46akS/vKyOU9t2Qj/52AN+CS0wT82dZt/
UC+z/85QsKOHDHO9DLXjtf0C9geQGz1O8lSmbw/KBaohwO+VEjgMxc2RCoALrYmcxnS2AbOO5kXA
G0DnBe8t2XaL23WJZf7eLgWlHEhF4QTWcrOH2h5Y9LrLE6SvZyT3Rp+2YVke7Hl5r1ovsZ/LO3GG
tv+yNWi3xj9c23Se22pf00hRcwajBQJa7cKQwXgYR34UacLlOCS9/SioVd8jnZb+NtBMSZqgdnJQ
JqpO/41/hmlc7OuB3oVmuLHOHLuguoBhyoMxoKbFXyl08qjCmFlToybaQdcrqe5wE4RS2G49pq1b
6V1oEVdUSTNRf/E4QYomk+RYsgkvjQODtknsSPlR0Pj3xbAvpcZ7l5HBxyxhilsDaWNjHxlrIYsT
CuOj+IotnwhNb5FJnND5hHZQqMkiI7yy6K/6rNstvmOdBh/XWWP0dbxWDjDoFIT7WubJfIKT10N5
SKvvgOcNHmFW4Ba68zZ85/YAXgz2xmwnRBm/5A8IlMgsXl+YBF6QAMUIgv/SlJ7h5K4e+2B4OhhJ
PDL1gxHJzpoI+z3l6UmjLmPJ+S2dKCgdw8Bo8jxOB2d92OeKqhAKYc2H4WX74s9t7rz9OqalVzlO
EO9H2MhTCIAEiuxO/gR6kWMXvKgpx7wo/Td7wsyuoLwIbo6MYGzR+or6EK1s50HbGaUR7SjSBOCO
VH4XBHPaGB7JQgGnAodSufYQMCKue8Ci4TI29WIdPL/ZXTObdqjSAEkzERON1YhnRK5mwVg2+u7T
c3RpKXJlIHkLyKSppJmCGol+D9eqnCZB3QseKSkaiSfyCxZZJ9DWTc0/epM9kCnIw2dSocmu8EmJ
lGu6FnXEMN5TKsjC5CSV9RleySb8KTdc9fjPy2QfLAp1qcUbd49l5rfUhzE9mSMF2nWGLTSaHvhZ
k34r1f8WR27p7d338glGHHMTOxxXodX0yajNkdE8FbeK0PGsSMNtT1xuIUyyIJsZVu8eQBOSZH5U
AUhK2lwkbnDYBYDHraYXROjv1Y+x4jHURIJ5+bcv8yxvpTyphtzThaGAS6I8urriAJcI5c85MIQg
R1iwz9KndrTG5Bbrad395h2lKL/YpFpnFud7n27Ph/YUl7IYjiCcwLL7E87LeREPeZh9lOFldK6q
uoKusp6O3IdDnSYCCX+LjdVoun0uqjmzrrVP0cX/dANcIM9PwTtoGIYiDKnBR9lwp/cCkfmWMO83
jqn+/4/k/qnLZ1NUjaOiVFhBICr2RJb1w6iEMSy7mX2D/30EEL2mT7pnRb0Ns6Nb/bVzsNrIhznx
CFcfZ6pxCX6bu50NUefWT71HleP44KL6qWWZ/7nCV0SzJX1kGU9vKpV1gXuIS0SnpHb2gFVdT61U
0c28EcMbBD9bkf/KJ/TwAer+I2CowX0mDg7mfgucDxRyVa8QefHKRIhRdTdef60T0DdGT3IBDBEk
31VNxLYTwH88rd43SArVpJtzMC2tm1DdYU8gOyUjhkKTNMVhnPj+NK9kGrokMX7M63gOZTE6dmug
npJorPDXq4Sxc6gCVr0UNvX9wmtvBUT72lAkeCz3ErQy/cMJ1sM2sUadkgT0ev1c3Vfes4yDO+Zn
11jVknYaGm0a8s+Vk7nITOFM4Wu5DrECkH1Fc/reuzHwUqklEZI6LH6CQJCR4o/y/lcS+ozYx9/I
UmzKuu2N+Ra1ef48QDHsPFwxyEe0PA+j/JERuHK4ZWKLYA42q5q3APfKirwCy37tuax9O3SqBasn
NoIHxKjqQSBqOXVk1Bv99DNbNSzvfdr9alYvDwX2U8cpmzfz3EFDfvI8y//9wbeN6WTmeEUQI2+o
A+FoUBbpOMnkzdIbw/2g65rdAOYWkyzZ14xP1571bMvr1+RMdIEJSXun8QRoWGZdNg3tHjU6SevO
HnPEuCNAOkmp97u05cZZQL9z0KROe4Zac6xKRq4F0oilDNDYNaJt+ZlsQv4t3hWfzlyBZAK9c3lo
JJo98C1U5Yx/q9UXcLnlXrBm/VOcD/HhMgcH8raBvY1YMa+E1LEg240DaHusBNB7j4IOMLLQL/Pw
QdRY94Ku4U5jYe5xNpw6p9dbd7KODACuYQFjC+XvNJNPZ1+I31tj8hKDzbNWU+W9S/BonplFkXrL
MZirLRx9WY75K4+IEbj5eP5o8l7R/89LT4OGj7hjIWJYStsql2q+cxD/i7C6CSAFC1qjZy/8Kf9R
TU6Ve3udUFrPhjvcfyXlorXQA85vVqj/8/WWemaUthhaPbm3n4pp6PVrRYBbfz2TcWz9us0ofv6i
utqjt2LhdVulSL56wsY5ACsxZQdpgkdXNxeTy3O5LoUB4kGBrOvuXNoLRRYF21PZqM3tn9hPXheJ
+PWDnpxjCGzXkmoC2zXnaknFy5NOC7TjsOWzUGv9V8+QCSYjcFGDhz+KzBf+27oXujkmMD79b/bl
uVHE1UozykCDWJDVrMt85QdgmYL2X2/6tsDZCVvQg/BX4+AdxvvmKPQc0t+GdyKsmZg9aynDRTlK
rRQKITmjbVi1VOtIva22sbt9wVjW39ltGyp6d7cEsX/50BjjFVyPuARkAb/JqRYLG3F6g6ciI4BL
8DMwal1iacEQ+7tGcuZLh8ufOTM7kZzc/F9uAAxYndwMHNEhiaqLSgc2+2H7qjKFYFcyMnJUHCg0
FAlerIUKVme/yo6ortOoveRdicgky+I/NnYgnHA1GgOg5Qfa76Rgflis/FdLTMWYJJp0C9oviYjC
rYCbIeIUqWH7eH9MQFDDUioVgP/itEQ+XPlcJ20OYO7dZOLKtLvSqdV/U0A6BtQiaB6TNfmLQoWl
YvAT69aAwCXLxXvempBfkxpb3Q/4rECaWXBINCYOwCblGGT/vMpCCpkRarJzztdMPgHskmjscRn0
Ph37ENvxJLa+ORTV5rItSp55VXtCQdlmjUuUHft4nMRNFYHQJzgFiNi/hdaNv8Zh1PqCfDnwRRpF
6BgqV4uF5KcXKSS2emzkOxY7e/cpkQM0Q/ogxxh0qgk/JQqTykpsQ+1gfvSwwjcodvZ7VHJDYViC
Wqyy88UViTCjrpgAiwG5akN8WJDp2PPnPJ1CEcIqJ2DTbM6aNHpsJSKqpbGPtN61pEotHihzEWbq
Y22qJ15IrTEetTvozM3eQVA7+3NaCZW+5yESPmAov5TCZwM5g/0/SMYROxOV9AM2+gmhWxXVymjc
KpWOQyhjJZ9JHcZM6/qv/U+a5Lg3u0noovVqk4xb6FrNd+wFyxeuV4p/ql4+Ce1cw1OURfENkHk+
QZUbK77MOrd3UoNJPG0Ew5eTI1COf4RiDGexZow/7aAi4WHVsjHAGMP2pdePndrn1V642vSsRHBz
OOgkOxPUTZPFEJU9zngyA1krUElvBfpBH0W/PEzcB6iApUvn7nRt9Hn3WSCBapQ/CUX0bs5aMLeY
YKvJ2fTBIq16z+nyHUbLK2RFtNpgUlbAvYWc8c2ZWU4wo91epRs1sGIdr4bgOEgxU1Fk3RXM9YxA
OTrMLdQQatpi9xlNpg/w+4FjADbXYZvJ3F1L/7yBufiWNgmmYNjx4b/6x/sGuWwtaITFgJvgNhdq
NCJdObuVe2yapBALTP9HCQIKuoVlIIAY/d7JlHjuAdWbLH0LG0EgsHNu4ukNY9pSSYxk1xc4m9tK
fzL0OByNf+XcRd/MM1hEDQ7aD9IKgPotd5sRXUaDBfimGz/U7J2j+mJC2JTSxmJrCC8VLx4/dhUF
7bo2FGRjbPhmUCHHvi6R+KtChsBWkWqrAdrWZOJm40IbC3In5mIIyy9Y4VlJaXF+8M+Zr7dhQIkl
QIFlGuGWONDEq/XJgrHTZdVyiEPgacazX1iI6Y3SsimZ+6cPKSmLCPduQ2pGEElimwg+a2QIDGJ/
LiGM/E2eukCNy6rom4i9z4VE0m2FL8oP/zXW5ygvXFv6ndjpwLjKYsaD5siq0t1g1NKDjSnpD8tQ
aN0rmmrFNYNtbkrN7OC6jjrNN0mq3pnL1hAevOU/MkamRA2u45i2FHfn07Te+ht5sKH+FG1FD8J4
xM8jM3chuDnK+aYgOoacfLCDaT0ao8VtUIfb01FPV+vuQxvrZdxq2eLrJayCm9z1faflAeTwb5nT
iGT61J0yd3UdMuSTrendKextB87A8qVhWHsLQp6HQoyoUTbt3riiqJhOnN9qtclZ6NBGOv2MjCTK
XKt7/ZCuY8woavKriuDztgxah2sVwc4YzcaJIYsztmusilJ690rkK/FJRVEu46TovFf/1Ay10BH9
nAz/Om/v2pawaztTxv25icFel0X5HErOVJOvHSy3dnrVouiaca8AzGnwfCv9CrG+0rxVrJC8O+o8
jy28GkT6YGLTbv1JXSX2qnYutthAVzmZsW3p4DiE0iWHaTT2AjewXSBx4MbusWGFIDUbfFdXOA4R
lAMZ6bQ1bS4vnqfGWA8ZblMEyt3FrzqtZgMT1vIMPU+X5IkOgcWpL6mRXKTm0xNKnBIN50zOXrnm
slEiK8B1IXLbJ/Y4lxbDqKx12i+NRClxyCcwz5p24QHwmOWXuM63NQ3PMpli0DEgRNykGDOD6hll
fjOQvNpS1BwIs1xD39hdRSq+P/jRV4Gb3mtpZuKmik7D6CKDgdloBAQpizZ72cdvPTKHg3xEuY0z
eSe5jyogPX12b/lpTBj310AOQt9JARHV4xd+oRnjKMyOyZk0EOgGBsggNnoPbHNQ4PDpc0AQOtkU
MAYqQDe9/pLBylH2CW76YEoeJW+EsXl6gFcpPJIeCeMe2BWBqCt2HhmTxIn1epkhCXuXbYGXA/Jx
3zO43NzONFT6CHhIWJ56qWxnKBsJfnEffZiplC5Ebl/fJcRxXk2lPfCwdzngP2HteXUeCAr+Dfmp
IEdoyCHwjQnqW6zGHxLCGPIjJTmzZ8o7ewTwIPg0RWx9b0alJ0G847v/ccqgGYUMGg3/hbKTxsIJ
68HIabmGdRGDZPqlPFIAiKQIkP14rzW3wgNCfecJM9c+v/BTLkvxQuI++XdQ0ET/lOzSsEq0e3hf
KU3Tz54NwQI8rOUzLcWUhpGOm/FT+Ha5k/bW04hM+dm9CrzoAzGBqyh/dhAasGq+iv1EB68dzw2z
soj2fR/2ngxnH6lnbAJm1S3QjUgk6YX00Fm9Q3tBICqWo96blBLgjp7ReVky6JKwaamN98lqR2Vb
h5UcogSsJLb2TQVBf+5XkhjEgsOt2rZUWnzsImNL8QavO8fnDxvXcKoeTap2cifmak4r2Innh14v
Q45At+0fWEK8qIGh55TBEXsqxbJIGDIdDs2a9AKtm7AITxArOE71UHGJYwDoBlxhRB1fv/xar536
x9Fycd5dJIbum/jt2ngaryvVDBIJ4hABxfXRLv3q/1fi4XXm8zbvYwlkW417HZLft1gZOuCgfDA9
VQM5tZ2bwrPKNpsbckuon9DfvA59XI++lM03rwO0QQaDb0Hn87r5GZk7F3fO5W+zTrVF3I1OJYI1
TLt0mUIcOCv3O52Dq1cdLEyZxA17ZvCBVeNszfkHcOSxiraYBFMMIB/VeLUQthhIF2I66XfNm3EF
5V1y44UnQ09DdgBBsWbi81uOT7nam83tBMqw+GNpwxBUDnnSrHLEblTRVQPWmfIVGQxMJkb7oqCZ
ZqVWpic80QV2ks/0EBhaBsRfY5CipfRInZLXfJHaSxDxGzw1GGQ1gaFhfuf9c8EQpkStUiMHl20Q
pomk7DzTaVj5oN19xY8c3z+cGMzAimLmaCQwvci1B7sa1OJFZ/2bOPyLmf3CHQ+Ewk7O5PuCC2Ej
OxcZ+376y6SkULUC035izkOVd41XYkrllGGILCgbSX1XbmBFnzO2rtMtwFLTjARbybzcqvFkvOOY
Xd5RXNx7vTmYF9wE6Zi+V1xjAImLJ5UDIdR7RsZHPgLow+rhqPfkntDDqkceJvyXt9RLTw46bWAi
EM1KDwPUTHpT7o3NdN75McKJUaez2J58oPVdXF/aUch91Z8O7sbLiQynWbToqcrLvopZMEi4W/sC
bClXcxxHEqybZNjsxfxV9tWFfLOK7byutLxK+DRHVR7jAoTCj4nVZf400Gf+O1iqB8HtHmPBJDZ2
7tI81ToWns8IbrqPzicFSF/SamJQarvn83JltiTWwFmY2xVEbelJHsp21nejl8yTd/4Tr36DtzSc
UDM8WftRM24Gtq4ALMl3p4SMEH7bP1ssTt2C9C7zYoMkjaWQ7sSVolJ8peQfOlNXqI8HTJYQiQUB
fyjoHTq9xrwJQ0Z1V3ft/wgsFkGiRXNKrIMZD6DNf+Ht7zA1eqgrd9nafgwnSzym+Ahelu7gTUN7
XdgkO/neb8YjMIkVRAYqEjKsekEucm6Kw83WUQgyHDfxeZ1R2T3IlE7PNgO5MGFo6iCT+GftDsCV
pm6LzF17DRWZlcnm98n+2GB4W8F5fJz3vat/lphyCXzJsJDk+Rz75PDN6efFp3aUTbIeAwB09cCn
v+WVgcjMM1xHmkxQzFbxBUuIOgj6XDJh/oqjctSz2mmy6Ui01tobdSlI2ypO4tHL33Qc+4h303x+
FMeMTNrvV1P2uPWJOLjHwjKtxZyDop4M1+pwPwIU7CuPG8P0BlKvCurlYx0hthw1c5pp0wvp6fnQ
GsB2PvDk/7fAjVzLLJ2zB13XyQG8vKVhgVberBZ6M2nJdCpc1PdDJajdvml7BEulIg4n/3Ry2dPH
7BfSXx4d0bHcaw3/bG7iQ7+6laYF2cUdz4Fb0aULd57hPuU/MbTlQ2F9zdBbsNykqeez3xq2lMq+
M7epI25xc5W5VdDvwtbR5fgvD2r8ji888dhCm5bQVSiMkXO0CYAwHqmqQqQLLEMKkT7ESpIXny2q
al9REHtPbmA0b9F80rBjtBAXDr2UfKbg0GVSTqg9RRU+RYjc78NjXlepfW29XxAMNbhcBZe94Lh5
+oSmCsdo11ErQ9cI+XqfZ6wmWunbw0Mh/Tt9/60zBcFpFzALuKxkUeTCQ2XeY6DuF6OUV5cJ4+hq
ShliG27z9g5uCAh0feWytnLFOBxoYZQZoSPdo2xInAKa90gl3Ea0v4RSqOOJmY47dm9CtSuP2ZhW
il4QtaA/pPmvOyCLaY0r6w2F8aG7rJc1vSgLaCS59pGmI7tSN7FcYWIwCwK9WG7q2pW7hxPEwB5r
eMFnb5caAaG6CeNi7OnGeGMBuxUzlMx3CGZp9NkJKiX7+Lhrzc/lTN0sOShRKPdz/dayEycNvdoj
/a4ZBLcT9clEol08XFRS2TNf/3OG0cGsF8HwteJHjQ0+ceUSgn29SNYMjehmbejSZTmW5VGfs3xA
Jrc1D/MDkO5JKLOEuaAByJa22n5851tTMVLzBHVBOWbtR07Ah1Ey5blHqnekU1/KIsh1VES/3yS/
h54izD3Tkt+nEYmAWKih17A5sIUF4jdQmlfs4je9+zx96xT36zfpImCdVrAhcH6jEy3LcH4mbesD
TRQlQDAkWz5AF/28j7FUOysoTQHgyL+2ht/lsCiXtdA0SwJjAXPZZx7xXt2rvVvM4/OPo1BU8lfK
4B3nopn15APQEK36JIAE+9QkgaS3LFx/uqgGhkVqoEbmGQUOK1ORL+Zv1cJbTXLv2520tF6XjMTy
NSZUrj4y2SbRJwqOdYDFn/TjyWnSkNwPqC1a4c0yJmVstKswLp0wZH3UYVoZquWbSNTvYsUulG32
5ouU++wtSdNZbrKNG8oxesfm7Y4XkpBzr6QN6HZ1xzaA3WxiDJ0RsvX5eIle4FumRsdiVF8dJxbJ
hmpW5Ry/4x5KBPEACL/1PlY4oew+BBt0GfX6nPaZyrnnovAy9t2xqqsLG0jmBOeHmrgef1JL90hP
u8Ke7pqc2WfLq4XHo3+L3K4B49Tk5vI4F07WZzlggGnFjVc494/JhWONS5UkTGZym+lL8DHTAXZy
NSY+xnfTLolaMPA0/cXLYXQnnqOX0QXyhNiEexIgc2nAtFBk0FkJjf/rx1z7w5sTuoKY69Q2JAV3
gf9/MX7hxs6wai6iGSv9dfm2H3fX+pynxkhJFYHlY61i/7bvSO0hgKcta2Jb2wP8WvLRvdQK5K5m
Ujb025g8c1F/XzCT7axwqItMCT3IjtnF7WNYGV5H8uqEHeJ9IX1dgHJFM1jZEFLytrtH4hhJ9G8h
NArA75DD/697b3UucZFDhl5W3XFBA/LGYyy0PR4K1Ylptj6866LZWwTO3XS9pVWVqPH+4r5HkcTV
hUHtOjx993PR7r0RZIZyRw2aihfXR8ZhsFq+UGzqCl5jCbVFF5fR37D6R9ZwomE6m41R2AYJlQPH
3odV0q5GI+9gI04DMbN7iSiUoiVkc5xiQESIqAnmC09OoTpdM/KwIY2TyMZmCMW9h1+NgoYVBl6G
Bx/JwIwzX4rYFyn7vr/j4S5rf2xthm/+dJn6lecbVjUF3ZfJ4MSaBbeo+L55GIxe35GlbAFyu96/
ozmJuLVP3vw+BfNnNuDhY1iiHC88qbSWjjDu632ihNfLKJq+QYrRQisa5sJ/wt2DZRz4dyT/NhRT
oGpWSYqIKF6cJh79ldrpHEVtNNQB5zb6noFm+i/KCfaFtFf5PUF3cqa4S9nJyiyGd8rMLlNTMbes
Oc7q28ru01GupHFxeMA7aJEcwTF1LsiCQvbOj415xaBR0mNOJ2GBZjEzeWQ3H/QykSi4zeBiEOBq
cU2sdtADlwfKUnEkLFA1A83nbsTNDMUgJKmDf36T6a00sMJsZXXJYghSTrZPlR9LVp33E176B9CT
LS6quRWmTJD4fY6ppuBXyzKR+UWw7gYa1BSSNeAjrDWu/Bv/yQErCwl02aQYNerVy1alabRuYYlB
ePy4MWchy/0s44f5+icxvAgeTuja8SEqSuA6IocJE1Kpwf7T28y6kXM4NoErJZAOcaxbEipRseWB
WVm6CTYKMhvqegdUyxhaYazDJej+htFIBd7/L9ykE8T3CN4OP4VI6LLPcfoAdT4EZj1/WJXLHLCg
3LgSx1e+X92tnwPM98fthBqiU+1SOHg0S/ut0AAbGhq3Wyam9qSPgLvYxmh5Y6ca2C2vtNqPB82e
FmbM4i5RLZzYHGVQY2WwLzP2FFUbaLGm3iNTgCEYpSk3UQMH+OEp8a5/5UYoE9K7H8r1/MHwJpAK
GRmp6P0pCSte2sAVUOccDMy+N1gNERMkMNOL6YcYDNxkxX5MLwHsEDtWoQsga/VlleE+o43TOCoo
KYzO4L3KmMg1l/Sj32LGhSV9h0ZicXoiSsDqQnPXpZ1fMwQSOrABHBOBWPGnb+y86mE9+F/QDxO7
+6EFRAwXFPoVyvdw7KRhLpuRIMVEKfXdk8GYVlhXwb8oywGncB0A2psubBHn61FcnUGAIKOw8/fz
TH0BggsHYpEYzTdSZEfuWVpNcNsULcXSUdKd17hE3REI72JeRFznPo9TmKocfXgXY5dqZsE5TB6Y
KMU4RfoePvU8vTicSKxD20qX7omwhUeZFDvrbODzpZKJ5BgKLoFuRCZKr+Mvl9bN5dS7HyT+++j0
dfMK2T2UoxprfDkv/RxwWwaFjUmraYrxmregpnXr1b2xYl7XDo+VCYAvBHCMBvt4Gx9AWmaQFG88
+xryjjDlvFWTbmEygzliLN8gtIQQFJmu5JfEx/nz9rWBmA4ivzaV9+1FcRHnHBdccTsy/pva4mmR
g+kQIdQsVoSAdquAz7BsSqsjihiqzELNRIdMo5oAdgeeS+nuCkIgYZ8nzVDWlFLGZZ/PP6CtWVTh
U5WT/j/8ZY3wfHIZnReAdKIeXGC6MLUmurpz7l8VRDgP1LNPkYqCDmdoCazt+GEed+MCBC/0H3MA
73atobOvYacKtHAKbYU4kjxEn76rUdTSeiGaesHRJV8NELDQ4Gbf25GhCrJkOWPT3xHFr0iwYZGD
Q2jX+Owc1BJWz/BEEnwC6NjfPLxQZRDIzXb254Hkh+Klh6l8q4t8bnIwp/YKvczKNDL0fuWQT0Mv
5OOZ/4YZDPb9p0/CexiPw+PQ5MILuT4mzd3RVkmiNvgAGgaCshDUiY7N05xqCtISglWywfInmUBU
QRNx3A+3W4i020BLtDWG0Md5SDh1MtZ3AKUpOK5GsT6TAvwsMwhEquQvRSkQTaI6xelBfFOMZfLg
Yhjk8RdijiAU8tAbdVEghyPGfpMJ8YO+V1Zs0qFLiPCR26lzpPko70sLo9DhUVCps/IKvRtYumAl
G0H1+ZWvWFgQlA+QSqIwMCu2nx/Yp/0xXB6BZPcnM4OPMIqldF/anZUwb3xLzM9sE5Vvmfylz5aq
Ajy4LIDxycVoQaW8be+KsFIU2zldk43eXumwTa/t6jvexcq4jTYskvFJtpNuvmS/alZeva3qqLW3
EXcE8wb9EEbJ8n816FiVS9/j9THUv2ULeZfoRn3E5ng7TgFaqapH1lF1KOocOTpwdKdwMJBqz7ti
FMIWAPBeCopfjR4mRVCj93ZE0WSUJsKoWAYaNgDELMZVac5UphJd9OFcC5RnFl2DrE0PPDuc72OQ
QGYyvA5/7lD0k0qIkvHAOf7VdJsvjisAOcf4vMzmQAWEViHKq7tK+AYHpHQtJiZ+oADkTqXFvw7c
CocxaojJNia9/UxQhbWWEfvgklBm/Bs2zrjVKmyVCwxirkW+qhAZyLfWPudciEElz6+bidv1PEIa
rLs6RsRAeMoj5EOdbaZ9buzrEdIJYjyngmCuG0vVizmcFtP1/QQ6QmOSRsskAvNmc019VIfF+M0K
EaGd0l4cvmzqDMt7JpqxnWCH3Ar9Wt2DzenSg7EPL36ZJ47wXRaNPqR0pN+wimy7v47MnR9cw/Cw
MzSxGIHT0eO034C8/UHSNoSBgSOuHvbe5dQs0e3VCQhTWI2d/dgqOPMAA6LK8extvOLSlR6uMfha
cUx0CPWQPi2W1lQWMhsPRn+gj2L9wElUBwtLIxcBGslrME4dwWeKSf5mW9RdFyBLWN5h7wn9Sfrp
X+L5Hrz6+zCrdEOWiL/Oyn/IxEpM6o0PHYj5we6mIEaA3SSeI1TBTkbj0ALTSY5ScR4MGfw3ciep
fjEpVVnGQZBuyrE3FnyFb+ufpAP5qKwiZZEKDPXOFSHOcBN81LXJiTjmbHZ/94ccFjSrLOzXnxIf
4VoZXEv+859xXwkfWY6YKhCrjjzKdJIDUtj66gOM2vwUUEtzp71rN14Ic2x+RpXF2ZDrd4K2QgxC
oXHvb4EpShkj46C5Sj2EYRFJZlAYsQY+rCBIsegMWxNroI5qfe8WcX1hJpmhihtFn/Y+YT+G8TsX
xIeO7wBFkTw1QRrA8lk7HPAz++mHizsGS5hxXNSaIKr9o4bkg7TqCtnXmqFCNSqPBfrqnT8WRpBj
n4vh3qw+rOcjWQsNK5YzdyNFeQ3I5uMBbMLntHJi2L1TcaVQv7dh+KmilBe6I6YM2/ulQ9Keh6WW
cS0rqWsJrB88Rm7teAdN+IRrAuo+FVTDOjdLipQHGs41RDrJKNWlPp/zijX7KjPn1qus+rQAu35I
8WPLYW6Bz80JwYGvWBKLR2qsfe9B3DsI/aUbaYfZRkV9qeEFZ5dDHlJOaqZXKE6e3qdobAkGXHAd
f147Y5kUd1qqxpQa/44mpjVngQQbBN6tYLZuUAXrK14UbHEsLuJTXj1rLPkTlrJlkCctjvJw6dBM
5R2Oyo0Il8MFBkPzEMbFu2RuAvwHX9lqbyjJH9kjrdhQufjHOiFXbVCR9VKoqFHi3eHBDoBlytVe
XCTLgiv0DCQD+dPfn1SH5Iy0zlLzFA5tDmgJyxjZHjPuv0EDZAfs8za02gpOW90DdY6KGDC8FO40
neSSojaSysXZYbJfN1JODUEaesafmKwK509IUmt0xJG2rbRdkJTgoAbcX+cHcVMix+BOcDgyhrbW
lGAlHCCWx0IagJj6OUcrETzqdB1LhZ7S5fNA5f0klMqXu46lAascvvfdnnEt0Fd8h/4CjGtHgmhj
NAm58/FsclYthAym8DRBOUs97/MeZ1pOwGxSoXhCmyNriUyk3zMU1r1vhaWJgqapcc+j3AqLdQaG
yA6P6AjUnJWDnZEufLxPtBx8XB2+0KFk35ydYTTudxE1n4v6I6pAk0djAP6XWx6yICcRuAbwvRjv
FP9Qdt2LGnSdajnwk9qYx+ckEnTTfG5mr2kbbYJyCtxSmhHdCl0J90rSRmhZNX7Lw0Tz8IF9XbcI
eEEE9qF8kfAEyw2KlgzuDdh0i/j1AftsM2pVkYo6WU3CMQBB4vCx47RvyoGraFkVA+QUs3qfY/N8
Cg3QVX7aNj2XNi1fLV9246n9UagMoLZqJZMscWPRoyPuHp216iCqkbEbPp92R7dXJOm8mLCWHeFi
OW+bRTvhRTcRJMCB1aiV4dD9NsLvwFBbFieAfT6wIQoLGTLt9JCyWwJX3uj+BMMAIeE+qBw5iA8V
REvE9YX5TDZMg27qlA6jQCAF3VuLziVUHclRkYGk3Ud2K0OCFmRvSMJHuElI7FKC+2I09i6ZdGh+
24lsejPDNjR0U6PL5XYkkRCD+bYArhoae4pFRyrG3wQuStM1quSu8MeTfWlCyh0M2MMkT2CONYMU
AHqIt3ZMEKgzShDZPz3uPe48SnN4I4HbZQeOxmpqLoKXAovPjM5bx3mtSp+PT7mhXAXY3FK9kuCo
GjplTWriDKNSaS4xptHu71HoTNQDaZmC15UEW/I7UkJDP8CfLCBN2tZcbtp3jSBAHKw3fhqgQS9u
qa8Nn7GEf2a9bWDW6SuNVjbd1jTLiTDi2OLT5lGtt7UqskhOwLrKrcblOj08HDJ2LHT5ZVEr+NnF
1j/g1xH6usTkARF4YhAKXomJDtVsvrBnkDZvUTFRpHwaKO9rLkWba25kSpgPTMoZSQqPM5QJWqee
CPtC7pHAOlVXKi5jbvWOOuLErqSuHuk1zgn8sCGmujVLjpuXx1A884MFSiaN+BmvtS4ii/+Kgvxb
w7DaG4lFQUfRa7ZPvyX60CPv85R4GcMceHnoPNgZkfuXcMQ8wT0oF94h2iTmU+kxIFWZn4vwJGv0
xDWzNZxp3eswGYw9W4n/bLXUJMXfSQPkPTZxgORsjM/sdeVo7w0cjZiGMYzsDTD3HZCn06DK8+Fd
eiFclkEZFT0W06V2xcCoBRULoWam+upUmWb+TBZhxj0eJ65i47Cge1uMoo2l7jqt46Ts431gTOxS
4WfpFjrHMFZdQTq4zbNRe59n9qEQqe8L1/j3+FmOsgqEMSuBHwz8qAr9P9tgQyGyPfHHm9yMsrqd
qFKm2zohz9D+eLTmn0061tOIInwQvLY2xYwphKZr8ix7QS+Akmav/RR5DRnbLVgupbXmFiErhux6
drdK7l5AVEjn5hDMgIXSA8uUQA0hNel3kZtv12aAPvcd9kIQmaCNXZ4Ij1W99ZT5OYOlvqfqbzUF
i8qqtxaZP97DwQ1i3/lylVdtCAwq/rR8UedQ44sZ8WUf9mf4iAl0lF8/zWFq4fDa3qf9LSivXiAS
B2yI9b+c3LimH7e0OnpJuYuOeb7giusRWsX9uzYtVqmW6Txx4UxVHS95dYqssNSl3kUcxAU8yG9Z
v0X516M7kNaZEkxvLmhV37mN+gdPCLQWQ+u82E+HgTu8TSZ5uoNvAL72nkovfQFdlj1xPVBbpz2x
lin6HM89l+sNg1PqZMOzeArdAcV+u9RKglC/NWAYS4myr70hB6WvmTB1R5avO8sIg5T8FM/4+CJp
F2Y17555H+CPNI6R+M89z/J5SuqJyrzUD7jsAX8/bka41lgm+MflgHtOAOz185JyRUtNhclFe6tn
Swcbg0BR+itsfQEfV3ayMiVxtuyODnXcfCtmGJ+LzpED9xATnKY76usgde+dlsjl4PS2tbsHLoGk
s16MFI3GyiOqrIhEGKbniUeI2uaW5REVI4kzWqf0F3dCML17HhsMzf07oB2noRP1JnUGDu/y+GJk
Tlct9Mr3wZOHHISFAriQYBWkNz2qKZcr2+22F1EV6me3fq3mEkyU/o5hpGYNdiOytpHJFH8tC1ed
zncPYMs1ViBhBav0+41KrunXtlakL3v1e7vzeRahhzhy7P576HUV2DqLEj8linGAoPFpMPVztrOK
hxP04iSbWtuUzQ+Ah6MiCeStqKv7zSb+vSAX5bVKzY/8EBmHR7V9OMiINyBVTufLJzfVDabRpJ58
U6/5uWNG6ZNn3u349sH1zuzD2YaBiXiN2cCxMhvvrkHPWlRed9ef2HJHx3vGHj/iVetvgtvGjQKU
mEMv8ijeKMl5b5K6bBfuZ7+i0dv6KGWweC6mfe3ylQmx9iBe1JfAfkMm/hgj4fdAfDQN43H4t+WK
Ob9JU1IMnhLOe8L6MNyXOjkV+ckEs3YDKubdh58OyaKQszb53IusVm+RUIq9ugTWr49DIKNpWtJX
j9s0Kqus+h8ijrxW7tDBsueLk+KxWMrfi7p5OPkROBX3jR14LREI2l9fH2Dj8M+xMyhJwCjUMUBh
gkUiOBJYSN1VIfdgO7kN5PfOg9qvA9Ut5p/wklf4Pb+yL38iGwd1DD0L9BJ2ZTIqpEsq8s1tPaqE
sclQqTVURD6ZpwSoaZe0XCpaVLnHZtKlYVsBJ1Zz+9V4UOKwNGqCTHnb8rtd74psyGradL7oKA6C
V18lk915JH3t4bujzu1AistsGaxoRa1yMozuZMLwj+i6ksteRB79byx4WUmJz8AthKyuVSOIfy95
LRcd/N8bXx+TF66M4ODM5CVWajPwOiiy6k6gLTYrtPeLE+aBR0EXqbfWzTbwzFBYUgewMuKj6MsZ
Bw5UXsPfS0CxepFDW+AxJqD3Va+frqiXrPJ8fToyjVSpL6FXmqmq17HjR/dIOiGowpu50/TUvTXE
XMrGPTA538j78cAnFujt/RiZ3xfSETMav3kXs5PKlvXTKV+lrthJ3/Xr6e5iRyiIkOD1d3s+Jb6h
+i0b2hyDMEA6omsKTlATAedpbNg8lUVOKq4qls96gTZ2Q2zNqMV+jmo+RL9O/TlH1d7yT4Y2BDNl
YmubWypM1bieuXjF+GjYwBTIyPrCzjFVr0fQEuu3SDbO/p/qhzY9JO0v1gt4jnM+xIYph29UYSbK
9+QdX+rDggJoQKHrmV4XFKvp70bLKba7A90B4t83KGeiVITlYMSbaszxiG5Fh06PHN+WjR9AHeLD
XoGf8MzGV4FzzWjqchYf/qiou8pVoqbcSZgtkn2QaXI1GsnJdOmN6jXqIG9hxY9ECkUuQjBDwaKd
7hWuGCiL5vryzyHUVgmVdDyK9EAmrpLgILm8/VYS/tBu0kkV8AToP4tH+Q3hl3aGRftoYKQsJW7u
JbZCFDiChShH9oYWgcIZ7PfUJ7Tz4TuEh8lmeWugnHUIxqg0DGz/XLk70KP0Wb+Z0W73y3QN8nl6
Ywq2V1/bCHjhdChJil7KfZCwNrOt3pu07xVUJFwk07SaGN7Zjmmt0zfF4QvZzeEjo30DJZBpHS7f
P+gpD+cLDvySe7xVtzXYYvP2zRd/HTnUELIyaCxeeH2DiK/ntCCFst4q8K2zacTUgIH5udO7F2TX
UIB+8SJAdKqTSd/T+qllIKQVTEamYiuw5CiL5c8jNNNGNu5IkBuTwEEIu1JU6YirWdXNo1qHIJyF
69EYpLN4eiaaztRCO2TA2l6ZMpcXEBd7t0EM6m2no6g700zCAlTJ9twPs2xr16D/6q54tg9MSiFw
ToEMcjKlEjY2km8V1/wpYiW56a926K3BIOD9VVim1oEsDt/8Z9StUiBtdaCzzEOQA31UVzusjLr9
kJtdyF6PsQFlVM05qsU0Ql3q3K9VKb+1TDz+xE/gdMwUb8Pav6XCC66tcurdXfjMRsz7Ky7evB92
2ctcaiqdM+/qAeGtXFfSxqj5f2lUuSU1fnf5vmk5X3Z3baujuzaKTDzt0YrYwj6tGxSavAGcSMxb
qr0Ty9bcmjHtRNy9PhwHhFWYNEgHCxLFij+UsSZoTUvfKr6XFtAaNqQUQ0Pi/btHFCDkdrfkW11J
mDI2qt94xa2vBrl6u4kOqeptTX9erPKQFG8xwkYpAcrowAprFeEVqBeXzfG4gLBdIN/xADj6xQe/
RVfQtuvlsMNVdR7aLMMlQdsf/h+ARTosqxVppg+IQX0U8z3xLMK9bKVzG5+kGqgyUbNGueZwzNAJ
BcpvrMMci+rMFYZuglS/yDgZhfeL1O904fk8r9ti/ZHoXKC+o5NYV74jngT1dH8HxAtDCMbJdamX
1VPxrqF3OPx03+/XvsiMWmE0FiJ+eL+JgtbcpG8qD2DWBaY/0dCiw2mPMlrS0wXeUFOsaL8chovN
feP5OR3O5wkzpN+DnwJlSS8JrV0R33GM4MuWNr9qMCxjDyJKNc4YvwwkAOTFcOByvGbC4+SYyYVb
DMgx8WwX5/1j1VLQD/Lk+Nq2zkgknruLmKWhoKz4B4BhjnJcyRHOr0yEUkfWh0IuSoATXJtlgSzW
YzFk3GrfCa806bVQqzwlunnOWKCsHHtCFBKX+MFNh/n7KpzD3QAyT4N85Nl6qyEnlxmrFAy63Jv3
TZAU9tO95OlPwhxE9r36T55RZG45rPXaMHWnuQulBZpG3Jwgdw7u4bRqpZnYI90GctYVAMq+V3BJ
jHhlEKvNOd28CR/H2fnEhz7Prwil/HL7+PtaQQhnuLczNYDukV+22mNrk+7risVg/i4KKJ0hbPHO
i1b3b/lYV8fuNNzUbN+13S1NkzPBZX8tYX+S7VnlHSSgT6bepeAuLHEbBe9AX05Pu41FcutvuMIM
W2KLmDM+TJ4rtFmHCmzerhjtOwPAGqAhEHwWblnGvOYHIMZ6RJFTSCwfB7HRnSzdJYLMZtuESlQB
t5zpjrf8szruwhHNSxtya3C2BhVvJVE8lrATzIym8guUkOVd8Bb2LdRBkP+jH0nwNqtff5veoJPL
vQfT4BzH4UzcwPECz/0Rh8zwKOa+Q6LzADJSUTKEUjZQyaL1W+OUHHoElq6aTvEGwxIrHT6OitBi
ycTCrjH6uO1JXbb/+2ZlYbiHgaZIkSjKAR6PcEeB7DywrbY3QsyUwv8FFckfUmTeddhl1Jft6LYY
S6RLjJzoG5LpQ4NK48bVjKHKUHBm/JbOKh5UuXl1w5eDjVXJJLyhk4oF4lCDv/+Sw6susGv2U8WJ
dx56h5tXfyKO6DSt8OG0cavr3VUz2HS8WOVG/2J24Si3jHfTG82inbMiAJtGCIPWXb2dDb++r7Zj
DoHF7O9OCBbxfekktH8LsiJWXhCnVvsD1Xng+cPrSDxhUBAQ/SQWpXpRq1B6kq5UIcxL9vprdxzL
D1DQwXZh0WDLjZnbU6RRSUBTqoipYbAThaHxiurpabftbaIJlByrFp+AVic/ldG487ZhaHUBfp5E
MEZAuaN2MII9SUsFDrVwvmIGnh6gRq2DD6OiLCUAiR66RrDcGBrkQbOsNEwYVZALWWI9su1vjTP4
KvpBoyRtsuMt/YVm8gb8dmwe1qmuSDQ+UrdlxwPuj1bEJSLHsPaRJs2CyPdlqE/ebooDf7AnwLwH
B8l0ZZWGA8iempmp9bcKBU/50OoDCVbxmJirdeJrJ/rit9AqUY15aUjm+SoLhAD7bOq5/zYtFb1Y
C/xtQx7My+5xzaLfPNd9mco5nLA7gIjBse6ZPsHfX1jzaaCF7USp7MzBRRCujJ6PHJTf21AD6RSY
dY1Wzpc/gPdFNd9BHNLN9adBrInyPsrAvPy0ba+B1aeaZwxgMtMuAgHGjgvY9XjJ733dGDU0evqA
YmgNWWkFg03vf7/T+Xds8BNAFviZhpRhqdL+gFpsmOHmil8jH5pF8o4BqoWyhgeaYYMH/dEzahvv
VSM0KzKLvKXcOfLif66lV7W9VXK/DxhPEpliOjBtS7ae92LNZKZENlJyuhd2cuKRgs/CSEne/SHa
I7lgKsjP6061Un5+Xbmz/EuuIaRnjCmtrnrwjDw8rQdt1owUxyJRuCVgaPNwqeMxaPDtoxwK+Aze
opBWWAKcLO9xpErBlwcKoXELy925yKW0+ZA5mPHvdIdmWgX7ZPqiIvCqFVtJT6ADbQTs+as6JJ7p
sbwMcjXeSSStl1pOhJRlhoeoZVbynoHLI8gGVRTSkcZCV7uJ3go3GCQKMx1qyXOHkxCW5QB/AQYm
St3BRawTrXECk/bir5zy/7KB/9YB784o6kvGmladvLyC3bQe01IG/ZIhp8w/yAQRAZ5R05RjDdzN
vFg/e1BVzLhdFMi4vRcEa2VMMAUpE3qcm4btvnEEKHuqNPkzQTxRPqjB34nrPZ0TC4TA3khCcU5Y
HfihkcLGk4kpxQ4G03okmm4kBapkGiWx1eh1ZBZV23VcfN+i4vcMhUK2xeKtGwIMlHPsBPo6op0B
T0OAe5c/22k0yoBL6MyjuFF/+V2ByPbvx4rgTFuy1Xl32/4cGBFD1d0UsJgpZvOFNZHt2yRF5loc
KCNOgeajmDWiirt6E5c7aqGcVavFA4NPyW9jZRqHSC4+v6JUenLS1X73rMQb47mBaHE8B9kP9znX
tFgIDdCJeNAP03s3gEzoPFUPae2333zHHscq5tEPOhzputAqztGXg8oT6ZZ0vJFmOOboJeztfCrb
gE1mNpojqY6SQJgFQFN7fY5HlG4gwPoKgLpCg64/pkyNKRn3XnUkqvvXKWmIYFqjeJmuzgxTR2RA
/jHjeFNHjvJWcjkHcoXt49/XXXfQjBVcbRfk3a8svnAPBsta9tSbqOVPjiSiR9a4rvCdJ9V+1yI8
LSKGlx5sOwr49hJrHAJIOKJ21uU/mMq21gZ6a3m1bG3GqjPiUm+1DaB9ruCzVQeMAlVNDqOWrjV+
aM9QyiwFs7kloBkeJ00npSFjzh0bMmhhNkEu6jraP6i8/2fu2QnZtOcV9Oryoa+n4vyxw0lra9YP
eUL8rayghH3EkF9jW0FQn0btj/lB0qKhd5NVu7KpkUXAyQW/B0v64gWahZjoq7cJrmV7Rgqae5rj
LMW9BwntS+vE8gT0QfGMUBUnHpq9Y/jHlC24hHQ4/TPWnYJGAJuBDGl177vU84yYhCEv+mSMMmFZ
OYMA5b/ftxrbWlpEgQzqyCdIF8mPFeZ3ZMPCB2VpHKnCPhZBjZr31PuOC/V4ENjNTMF2K2vTSyvB
LKZXpjZTXRDaFfcRIlvuUHTPQ4DhEbJ1RYdzB7f93COuLTHdOwesmEPKTK+zIyNzsituTVFtprmw
54m0GLSvGM+xdO1St7RWPRnpL+rqtHfeV0dU0vZ45JQ3FQIALYnPAgBgh5RFgEA0tYkWsNstInCh
jOnQrl7+kTgdfCMWu2gKei0/CCH3/cP5dO6B/zjrz3GTkZ5q4ew15u7GmqctRo+7V0qxeM19kCiR
qS6lFxX3oFRIfIZPuycS927kK/yX1sGOw1gDG0IJT4n79DPLAKujN9lON7uN2w9GI5I3G9bCwrfI
3ARgcn85k9Lkp9pC4PPRzCLmasZY6b0E4HnB1Uc5CaByGKQGfsZn9puFLy4adbmIGgw6ikSednqq
qMvom0MgqP1IYnsYPE9zhiVeP60x1oAxJlJJg8cdItk+g1r1Y8iiKRhwI5Z9lVFNeViDZZ1UPVT4
Gm7SvQT3BNsc81djzA6zsKdUVaii2aSH06ifkpvrdd53PCkjLYR1rsMtaS/+0mbvlAUBxNvUd5vj
kHCfY/D02t+F8I9x/1H80c6R6ymGWyVPeX/lYE7gMm+7Jp0Z0ctFVmvIhVKP+aMLVGeUWkIg9GAj
KnxWDCUqbJzUoVL5FBsPQ4sf2lvzxi+UH+QjGFmxiwGWWDURSQbyJo5hAfemf3rWKR7exyBM0pe0
AykAldjc5ma6Ve5GNc/Fp3vyqyZ/obHXcvfd9TRsRea74lB62MDh4Q9OpljUTA/aEjqHrkTKT+mT
B/IqqV0jqQ7HWM991ctauBG8UhQFS4A5NXuYSPKuEEBA/gyQ7S+0SHlginZADcO8qHmr00yEE/AN
KpcSiGr6IT4rRs2R/j27HMwmwrY73w7s96LmN1dsmEsA5ynF6lfdGg4VG6PdzrRMyKM9qjNiZIER
tvktEnPDVw2mL2zAeTDc7qFAcQ6AlL8hSxS7b3r1a48MBQyw0MzNwhISjXhiRTxwuJfq3u3HClgJ
w/6eNWqat6xcCrDjHBblkFtRMbLTwNZOEsq2B6gHFgaSWw6adtSVsuhOTHNWqgf+vLX0xbkomINC
U5gurYtOsRvBWB1Md4+P19abtSwQqGb7v3Q7mn5CVln5UdFQEKCov6fmLGxoESLePgWmypq1CGsk
v8FFy3MlmhTdllQxMFHFmrLoSHI4/dv+/bzactyaTXxWgq5wbuCqgXt2QnTHS5zLV2kW58FuB5au
i7E2hM+9s21sE55d2CAeXNCRrllmsAXUQXRwmBUzlQI8+8j4+aI4IubXB5bwokHtyc6nuwDuId2e
nBoOdT0tWk2ec+UJqKaSfIZPcmhmaIGAgs7lssNUUT6rZO2KeirMat8vRxNgEUk7xeduye8Sb5w8
KyEVHNwytEcgB7VdS+lr75orQUegxl3Zh+fjsXXAJX4F+P76KgEiExuBtvWuALFmYG3oQuxSmPW5
bBhL9bcHO98bk1qrTu76VhDkPw/2zhbcH6uLqVG33mqJ8SkR0JAIPupDvtN80rKKHmx3FBWNGZYz
tdtG0oe0QnJgtqF7XJkGQiq4CLsc3oy9OPX2/r6Uq8cjxhJK4kVgABu6apGf4rBIrNx753HiUym4
+gf/XyrH6x6AsInkyaXufzHPtv6wXTVRwZJRztQ65wlZtn3DNV/+HhiUR4zB+sAQJsJpEbv5sG0D
1/9PcT67CEBRN4fuNURtMB15Bfe0ZaVj2H80ZxpuBZmArZOspmKY12GAWdeT/XA/xpBta7kmFDxt
6KZT9DoGEZfpH60RGlarMJMpDMmZdS9Sp/tkG2n0EhB6I83KNRHswPcPfeoW7o1z61iGo/EIPhAR
cw7tbaLOif3KaxsUFn62LWI66NZ2ikMh2VHewItUNshqWZFeXenKkhIDIGEIkIqYWYUlq8pp0Kxa
aRK0lw1G8ct8O4yCfIbeNxW25sZ7C0SPs5D7jWFQcbM0bU4W8j5ZyA063qzHnWRJcPoIEH4r6wkL
Z4uMHkhvIB4lrZj76fsvKrLwNkXQJXFFk6xPyVTndZRkES+vZz2pAxK5rEtOKw601Oryq1O8Kj1T
z0n26v2cO65LgmMrbFRgsw0F1hRhvLIKulpCdVsCZS6wON2K9HYhfO9RPAnBcF0WcUlqBCH3GHPR
SZ86Tm6H8Itz9VtUGZBQnJpdi4bKdO+Iknn7CsCrPITgRFoulyeLeE/Alm111YsYq5nRc0TOKrWx
YSSh/1qey+sVauyoO4c135gmml1fieKwbqRoQ5L1Zc75AuqXa7RJMpPNvddYnyrmik74bxYcTiN9
j9w4rE9g7IZrtp1We9QSLhAc/DHFTGj+6Hzg+EJ5FqSDqJS0Dk7gJybm48td5kS/Hy0mlNa5fuHL
C50AW3DTBMj/AR7OZGp4lUyRw6sAd1dkjzNfHRULzhTrCWTyMZowS3ydRuaBISt/aSFVkyb+MoAr
gbX8H2Vh15WWOd7QUUVyNih3FmK1D0aFS11vwZZoJeVV7ndxvZmw9TkV4qM07If1KzQfcoDKzXxX
mO1ZPAHEwCtwbsYV8Jqyjf/UTsi+QF1RbvYGt9ycZYUfnbYTDcK0dZ4DH2oKF64W4aPxekxZe07I
aPklmoc+evZlC36SRXyFI1oU99YmxtD8JIW3H1i6qXDiWZBWhSvPjmwqjc+40rX7Sb5mBQCu40lc
uUt5rZ2FD1lFm7ZgnkAoQApu8h1pvdEi0YCpU7CrYJfcJXFhZOSrUhkHzudxOsuNfYboWCBWvjqV
6Z7xWUiXffUx0ceZZT4QCe+Pn99cw46XHxI2g4bZCk7tc+UKea7Q+cQy6VS7SUdqUSkJl3MLwzt0
Ruw1iFxuu0XI5NVCNLIe56NU5OuVhZ8/i2UihBBRk9EDNUbG4/i20ZklWqjULDfrW4S5HQsF9CQV
4iPQ35o9eTri3eXn7mG189QFJMKrIB7vR0GZU2G/rvDUBZxL6xXXaAL6zILu8cZEJ0nfSYSiikYF
mZ2xMiNAUEVrmGG2F0N6+qMgcjs+QEtr0u6zhCEFI2u/56Rer2/nWVOyyneRZPR59MOkmTHomRDA
BphF0PJlIQHM69ny9M3jtPxalay9SuHhSgJm3tsXNtQIJlbWS1naoyt+Nu49SuWQVwYP2Crj7eec
sDgH4Pj4h05L9W7p/R+v5U/cGBmutTuI9P+pVwxfL5v9h6tchdf8/IBsl8eMAq9P2xm16ucM8uVW
eC4Zi28Lt+xYkFEUJeiU/GQhhzexXVXH+6UnMmvRO0gzdi6MP8UjruWv1ryhptO8SiaKZH2lUXL3
ZyNA3ntXch+js6YpvdrPalx8t+PGU5i5mm/rbgyBx1l+Kd9JQuw0Hqvrkwvtmo88jbS/ns/NajLs
f/XZFQ7k92IgFoTeSRRyUWFQe/txMzSiwzgnweZrwY9SR82roMpVQ4ZSzeotYwwkw0AC1/h5sSjP
HkXaj0YXCFgOqKqac/3/v+OD34GnOmPxiCKyB6hEvboZ+dEM204YOwwRGprBLVZ5Q7+b2m4ZvDMu
h522wuSgWq6EUH6xIc/eizT+nnxpClamiy3ED3EBUBOlbrjaofx/p4vA4pE0p+a2mG9neJUE18nh
jZ1d2CqghskEgMEjiw1DDXKdI+EMpq/N3EY7LpbnfX7fo0nLEFfcrRfdy6s3Ocj6pAAH/Eddf8D1
tzCxShV2bSOQkOJdbuoBvobHLmy5bd7xP3IhEaZa/du8dEwhJbYEKXtpTnkUOme/J0gMSuYsm0oa
p4hezn5hA9LfWAe5fhgeMKjZH/6sNsog+1OJqjwvgBuqIQDmTiZCQ4auhURhvdIg5lxSY4vVqk9R
r5XXv2i4VdQhkS3gX59fmJHWyMEDK1wKwT+L0X1IXX7aLZTe6OSF2j2Fw5S1LJUBkLLbhcXPxgzY
PgFDAVOcAwrIPHaseMwoN05KjDrsXh2UidxJpo+W6GlIso5egRNOJmwraBDATBmVYhRzHaucOCub
KWt3p4XPCUmiavXYYdH8MyBBimAI7+2FrTqspWuClafZMegt0dRFK23w8F+5cBheItyP/M5EaCLS
WGAFbUowI4DdPiEp8ewyDkLgxgywXjISk5r5E4KjB9QcN6rm4WoVkK9C/IiVC2QcSkH2n9gjnUWj
vnGsMU4hqN1u6RKDU+3JXN4HgoLiSCRr+ltAWgEFxfViBcyfWbQnUOvZN+08GJsfsENiyDdmDSDk
pwUgat1QCRsXRgs8132Uy4tg/sIR9/5Fk9mrEVt/sWDcReNC6HNhNZSYS06HCcJ5JHk0JdbRyKAB
95/VGwKWJphKxRgBBOTqW6Ig9WDJPogoMG3F0X7EfuS1ikrRf84iScbm+suMn5l6RmzV4GbYArJu
ePhlr/8VY8sVaN1GCHimiJaMetPBdcHi4wTKO38ZbsM7gm+CZQl0z0fh33TWd7EGgUH1a3Pl7T5h
mb9+ikYpbOzxqkGGRMpPUgzWXPBdpGE1QkGrLJblHYQhCFE3KMl8SbEd+0Vdccwwo4CM2qaXFOSQ
wGtdaWGfumyc/UGmUe7P7yvWQK1ncsLW9JrNXTIh+jnx3/FaL8tN+3+a3lsMUTKVid8PPP3gPW2I
e96fVjj6wLwMf4AAzWX0EjFVCpfsvQsHu1vEXGm4w0z5p3gHNkANGvlkIwGm8kUcNzOSwqM6vFJ1
vunGh2D67bfyDWpnrBAbXDulSNEFJstKynVcwB1Fuxonn3b8mUZ3tvkrqWiH5nQ7KNPY69s0GA6J
LJ0bK0pyNGJBc/EtrWPOiC05XuGu65N5siYeExf92stZtHIdbKMW5yR3Sw/+Y0peOSMF+w7LXmif
TGUBGzvHnsoopM1/7/kQx/SbbHwR++i24ABQYKtL6BkkMfpDjsgkLbQ68qIm7HZwpHS9oowy4D7f
pHmu9ws6fyi051R1L76Xk5axSZMAZYtKiyaF22zgyxaBi2Eg+f4O6qhflR+6sVOxCQzbMhUrMoak
Mk0jOgMFCsu8BUqRpR3UfRcueuQ/moKaNkvYsfON0NxqhMPkxcoMaBRiSYmTUnH+s96MKKt68mxk
YBByfdDPMILgJzDhD5d5dDdQPvuA8tGR94Bx/wFGM/pHfOmPW0ROPGF+S16UIBYm/DK33F3ODZzw
44ARyuQSApzfzvR9QcnG6HP0RUUMvODA11ySTx+hxJLGUIR0UbLcCNChF/FShpHMV9I0LxZcU+va
7oo3nlRtAU8datSeEkpGD1Dnt4D+ROuTaJe11exME2nEbUmLQh+nLG4bwUy24AQvNT2y/12/RrFz
2JtR+jFUELt9UPMc5HQgALDQOoWc0Gf8ZYg24s+w6S8/dI96THlDHcpy7Ja44ZMfIxYqGozKJiwO
SRHsb2fbYvjMTn/l9ldfJgorq7ugzXVLwTP7IGu56vz7UzCK9U7+neOMGzUFrAWxE+m+Kvnzk7z8
nDGmoEZkVy3T360nDDzo40VIW/T5z7j3HSqzVFxSsW0sUxOkKdpqGNK95nNdRr4W9NVjTvyq7VFS
gJnbv037lGOTkJpR7Onm9/vyEVlayhArp75MaPb13kvzpeV+9zBR9aF0TQ0SmsgSJXNW04foefvq
zfZmmHzZDCrrz1eT9BbP/6qTafn9Vso5zip5rCZQ2lw2qS2GwTLbcBEYMxlRS/dp4hxbErhhljSQ
oHbNwq/ipnDyRmKksvNzXx8d3QH1rHvSghWLJmROG4ctn9xyE+EiRG1M6L8JlinsNlm3lQAMr4kE
plx/gq83Qzi14RAu0U3Y8e22qdeuOocHBKfDVya0+CuWDjAx14/o2UKFz/6mSWMrGKGRwAQapgku
FF0HA5cGLSD71q9dgSSM6lEfHTc1lInbPsT6HuHlobZwx/iLH8Y7jLhY9fE2yQR8hnnBSvfttq0/
RCFfayruvAqng2e+FYOfEuFxVeRC/kSwBqPV7LCczanODC6bVuBuB/efeEONqNI96NwDYknC/QGc
OCf7klauWPZjgRXZ1ICviS8B7+XhWVDlLUsXU8zWpXhxfDOEIBiIE5a3kB5uRJjw3tTqpSIhNpl5
08QH5aXY6Hej5bsZA2vgeOwJv15dw0cNPIlyOEI0oQ0LHHg7pMw1h54qBZtRPqG5kg4CKjS3MCwZ
A5Vm55ra3hguTCxJ91dlcfTkUxqlX+glGv/E+hLevtghIUon78aujZ9bGhuIg+vomh4VcHIqU1ej
vWAJHS0h/udi1jCjti+jh5l0yl2vpiwGRtevM/khdfjH2nhKP4TKQSGsSV4kTcq5HtnOzJ9JVV5W
AxXewMAKUPNGpGKMLVnNSaTmd1D00OlvnDZX+/YSDoTbwRLCgzPLoVqY06ftNip3uSInyfJFbHeQ
uZjh7D5DXUK+lytABHCClKtX1RSL5ANgAhwo5k0aeYmcZgyRCh0xmSf/OkGQSZU/EWYpI6KeO2NK
ARdQNOXNDfwGUXkVCEHL5x4lemtOXXn0FGhiCEDlUEFiXya0J2N5y6Rj/dcYutj8Ftyosd22ZR6C
r4i6JEh9thjtWwWV93RunQ9Oh3N0M07J3hG8lfY9+9hCxv2IEtJpFkR2D8pIKEEqdWNIe2XgpCjD
fohwFVwAfrZ0EtTgJ6A/GZ66rs81IIC2t15uC4JV5pfKgBNyWa9anYX1uK3wSg3wHrK4dfduyWAt
EfpyJpv3vw7vbm7cY1bYIjGoeReXFac1Oo8GQEXpJN+Mmk6Rub0ZHrjrbtWrT0MSdpdGOWpTG4EK
qTrhdtnO4arj2629OOcnCC+d79e9hgOQPpMW/CazmutIhsU0fzcY5TtPmYAgOYVH3xy8QyCMw20C
C+qw4z+OYe4FMadk4Rozcu5dJEvGwKYK0jhAI1jjJGIHMIYyu+HayHgvE6aaGjEM2D2H75e8fopi
762Xjbszv850upQZ5MVnMmGCmYRqjRXQnICebGRG/eld17byERJjg8v67oLqRcBioijNjtJvhlJl
994dQ/peiERj34Ae2xW0xFsbTtUeUgZnfpthh5DZr3/G9NK85vIoWMyaaMSEpljzpNomrEsTuCi3
phVh9STKpOvjH3rYEB9CKogytRuE5DD70JI3gHhfpAXvaLuFDvjc3f/h5bXf9qXpo2nS6wAmtdFs
KHEpRKrGvMdHPuPSyaQlCQZ2WwLn3pWtmB9H1MBv51gqUy3R7eb/wuldsHHI1Zs2O6u0tC1SwPqE
glXcYwPJF5PAR/iwxmVSEyEkQw0NF0fRhqjaMqdF2VFV0C/mEAelLgRPmiBO/8uux8zUSjWEbp+X
UFCoRL8kA1WDlbZX6XOHxbwyOmTdPhy36bGRUDaxgA5WpvFuGD/pSKipka1CKGEnVezzZLMzf0WM
sJsmF6MTun4NfOVIfiWiMr1AD9XobYRQat09eqJHtY+h9/7pWwKeeeLZf/T8DmU2k+nYFkHA9bAs
cPqVmW9qmc77JdV4G7rlrwOgmx5C2z1+0tXanMdkKqldOTBmCauDt5CeVddASD9D1t5dnB8nkCKh
LGLmMheiA5M6A1KGbRWiWUlwN5320GeRr/wK6i7DCBdYDJmEXefzRX5kb3RyNSkpFJWeJyGLTkfm
LVnMXmHjGV9cf2UV8k2QRB0KQCyN/Cj2Qra316bYMX41PB+wVQ6PBtUC0iVdLS5es9S/ppJdWEmN
ste1q8yCzz66urGRErGMB+zITAIRqFY2wW2QX68PqRi86yQzFQZ604Ar9foOkX8fDzslfRrXdcsq
Z/1/dC9/ef3qgfSbEAU+pFU7RiQlk7gsEnRtS3mqkV1BXupT46jJaAmQ0A6SZr2ysA5KcwVSI0Jk
BK9MkbA6qC/PH8n0wIM0nNDVlVd8eCTArNBkbn6CoaWePsUv9eqF4f5y9b6NbuYu6sbxzvOuNa9O
zeVGhXED5fqOypQtwKEYHVIgbbHPKPtJJHhH5tUz8K2SrAuCeEQRSCdlCMtBxGgg8wcOWATQNGwu
o4wCP/2E/ZFmtDJItXHVkMPoA1gW7RNHCd2SxgKA07RbvVwN38oZIueoqNoQzawdRqCtZ9CUB9QE
0XZq95nOmhC/JNvgszXRe3JG5gXZVaBHI18IigsBhO/063RAMZArvisOmaLi6pIEADFrZpOy9lHQ
X7WduKEqMWiT3WNdL7U5b5CbkibVe+B/Ogv2z+6guYlKJmGIikAMFfEXELZPVUCwcrQDuAmG2Q43
81cQ7kmSr9SANldDd/SOxylnZtAt07npmgjy6QeHVEvwDzKakfsM5lG9a9E68cIqTbEtNgo4QwXE
P4kqydYu7P2HLjyIpFDPwYoqeYK5+qByauVobG6aCE4RIG7SVGtZ5ENkbxcuRf/xR3/J2hLVZzQw
peeyheUwEdJvZHY+30HLCZ8RhTvqmZqHyNHDQ2U87+7N9qT2FeRjSqZjBbI4MQvsKE080SXuPHlO
0oZOAQIQRrC4Mtug8EKBtJl5SyVMDKhiER/+Kh90pQDOm1V/rMVBCN+hQogzmXQB60H1Ulhpl3Rv
mgZhg5hilWVi1pBZ9wB2KIPeP4svfe3b2rU3a8CqOsbun86pAszf1oyvYQ9NLGsT2/l7H/p0TtkH
kbLptXvs8St5+dkw+0xoZDF+gW8xw/mrknEXI4WcWFoJFllQ2Bpd1ReHCI2k32zwLhzjrKHmtWLj
DT/ALVxDcxsK0xLfETZ3hbiUaxmDAbk3SS0ZDa7760ai9f9TKK9jz/BA9afPnAad9uLtcw4A7RsA
1Z9DIPReEU6YQQk8HXykW2USmYmToIta7r6ZELU9zv+HtCHJMDdD0/M3gEc3VVfHiU3Su/zAc+t7
H4Hoe6VZBIVaLAkOJ5gs6AXiy4MAWlOVOYRoEsA8VvTEV9Bd9rY7/1sFxs2dKI/eKh6PSscEzxBC
wjR9uRlsF6NzWtl8e72Hcmqi+Nq1uzSuEgQpT0I1JJFY5z9a5uWVDj7xTly3PeCDDqCxr5j3M4Bn
CCcKZ4jDWP8N6kjq93BVCM3GM+w+Mbw5/jdNETXA6dOPJv0fIKOWebbdjqBhLgVxFkhlC5u1Ze7N
Fr7/ZHQbjdwPZKcHT0DPzV4r7YGGO+sTctdnjSbSKMPuaqTMXiGiQzT9LSzAVMiBZgGcWiCoEMur
pbTMxdAIjDg5PbD8XAGNx2sNkW3gHWNklHzDJJAjq/m6klCEsWUKuGIjUvEUd7hYMuTPNy+/gHSH
oYgRB4hmq/9Pev51btn9Tqn4Sg6zLmo38qWH4bnu3hWIw4GO7VMz3q95Wwt+MmXBa5zE3ZajZu4e
jCh24Wb20kjVnY8ZUifIoJ83bF27LIbAW1EpwjpsDNdu2rxVolTGrYrdNfHH5lwMBoqEkLeYdjqE
B1EKhYNd4dodwfvd+cZoH41g+O4XIVhBnRfQeKYwYQYH6utd6PnSP5ApMf9jvwb2siVpaQSmyN1f
luAMnibxoSg2WT+d2swDOiffZvnrYXODb9s9DdVZ+6imdLfV0U2Tc2ydo/xRvo8l0YHkmG6I3Gt/
CkE7R9Wywf2/5IMYwZCtvVeUPM0UJ8WhyUA1Do/ss5Vr6maZTdHvDhdJ5IK6CdfLPNUQh0AHicEU
6/JAFgjcMxoMPS2y57B6WumdKcBwjoXVWtpRZIqqHzL3frIW/dVt1rC6nFBN3vi3MPhaJ58Wct36
u2uGtYQXAUMg9nkydJAKrpM6eKtvmctNyLSK9fF5xQYDClhGrZw/r4CRPwk4W2HzTmddm4fPe6Jd
1BtLxHPc8nd6ergXO7N1Xzbx8aC5p56YMM4SiCe0eScJOH7YXIwwAIPUBh78Tu65huOUfk3RMXf/
o9bvXDZXpBRSANj7pYoaMwPMTazZBvxza6rSXQsRDcHt5Ytur1R5xxnfIzFi3ha5oa3cSz+hWmT6
iDxplNM9bS8LMBOlZEU0OrGvA+XxrYQYmLJPS+WU7ANiHXUyQVUy2ntf2ifyHHW6+tW428HCEsG3
R8uzdnqw1MGe86M72an1tiFVwc7uTkhxtMU9MzjFw/i+fVeroYAbl+j6/lZzg5HtZE4+nPkfW2Ns
bU6jBHUZbjVqMSaT2G6YF913mzHKsab7Qye7up2EN15jVnppD8qNRxb8o0rWsF4IqAle2D6A49xT
hZM2vHqGm63hi6Sde3h/XC5im7+P6LVzWbO10OHcpZTm5WoQTvcs8d63wc+0vs5ea96dek9z3OW9
DZi/n6UctuoW9+9eMVgwV0ncArXyZ4CR+Ldf/SFZOH3duOpqk98I0LS31jzcRvYd6XVPAx8WxjU2
O+S6LRaB0G/eJg1ZQZwgEO/PVlq1svFt2JJfLvQ25NDWmp8zz+dwFqWp9Tnop9jgPNUSru0PrgEq
gwf3U2OYTWLFrLx2vGLYfOn2uAqi2wxI3F6MggyYfuh9m5XQkb/s0bIygEaFEhFHtn40AjOuTsqH
RULGvD0R73fd3o6DyI3jkBJoyD7adVGJ+uz4Fu7/hBPQL8IvdQtb0eDGKVqnHrlHq1JNlBZd5iMK
o9toEdozgwy7xt4uWPTuah1SQXQbrfQvd9cXZWGuYXTs70b/sUlJ2mqBmGnDORUgW8d4z67TJXBE
UfXhLheHdO/JjRlN0FVTmgWCczCeB8rKY1z4f6NPEhEbXuR9Iteckj/7KD/L7TFh6a6gAuLwxf4H
bfryAW+811r5WTpdZHzN1dsC4XP/Umpl1T6eOdxjfyrL+HUWEW1Uou9Gl5xSBVGANIO7XC9qwaAE
Kh0gre8v/QMP3a6wfihkOvb9oWiiXtQKu2x2WgbDP6So5GTBxh9bpp5nZbegV8Qc6PQ+yW116JsL
cDr3mZ86rS3M9gbcV6rfuHQ+g0vPmgxttzrdfjOr2RCxQIcCcB4ylhogQBkKSLWl4beaomsTdD+R
FSt/W0TQxTWw+sQbtHBHwPnnj+dNUAU96W6d+FiFPlkoVEyNnEvnO7xbBafZUm4ZFMOfo3wABzsy
7f6RHDzWytivsrKdubgZ3XdxZfQAoTipVKEXd+o3svNHdS8Tk2UGXUIyzV8Sr3vz8G1Q8Zsruphk
LlNqTGWH5GbOm2ZR2lcjH60lJ3OGUGbNt0BM7T35op3p3sf06PiZEhldT+oqC/ztlFOob4nfBLnk
41l2EUEA3K5vLCJ+WGKMlHpmtsPvPDzkH00pZbFvLj3wU2isdSPSyCE8eGQ3ytXnJ4tQMMpl0U3u
8s3/gQCyBevIAGObySCGY+M36sNb+3ZVOnMUhP9gvKYHcIatnfuxImEQ2pLEc8LV0YxAv+Ng0XIK
rPujNP5uWaXWMiW5ekTuBOyx2XvTvAv7P0Cj5yLyWQhvctfYkniNgQCUsAwuFvCZg9hTDdgg88f5
PFruKUYmduzjQv2Fi65HfeRA58+QdojH10HJ7Rei9L2NICsInLY1XESe8+rF7TFbqIJDQlk8RJ6y
z9zKELGX+m+tOCYNxvjZF+r42oVuTFSllZ4U2QQaKiHTpR6kbbR8pn23WxYCi67GytRaX+YGPewh
k3z2aIGDAV2aHZsuBaXPz+LdwXVpqeWYiq/ErH6gPSmTLsTGO1qJd8Mye8ike1EKLhW1bbeuv85K
g7Xc8mPTj3swIibBbykfn5AUVuFbARPaJ7ib8fLm48rsAjL2QyLNcK8v7E0yTQ6VwushikC5H1Lm
+eXaI77UpUmkrLyScrlAumlI3BNspdFJimqBhQ7ZW/ZmmAo9j3Coxsrek5HyATuxiMLxwQiLsOKX
LFvRSJ8Vs/wvj0TmbHVxQ14J8ITN9WXZEMTyrO79+0H7nWZxcRJuAwJWgSW3kxaOdE7TrtciYA9V
l5qzlNnhcrRHPamT9I0E+6REF6fpHy2sU1UPbQfN6jrsBRbLaIrWw5g2mOj1N6zPCqiBMJ2jD3F7
sUCjquIcK7ADKMTINMKSmgrfErKbf+xlCHUKRM48lavKbvOzqm1kZ8v2wioi/saR+vM59rKwHAYH
pPhnmoOvqzpYBDMoxlSnCiQBVcS4SHrFGt2SDMI/z1XBbwVT9xckeNET9MOUjL7O3Mn24cI3Fm/x
PeffX2uO2cNnEPwGfs9qHmNNIzC1ZFuX+AGftv1rcEyroNvVd+ej3PX6T8bHqaPob1T3eSr5NxM7
866WrhMEoVc1UrDn7y2hBQmXQW1Z7hJZFeUM4XCfQnaD/pIrMWp2AcPHNuOrsWI5U3CsIt+SIA3m
ygUJ17crfALCcLoIFyMdOgXlVgTl1nVVD98uBbXpJ8YmkfAyhFnvah8ZWg+dNBt8jFz2UKWKY0m2
ey3vHneqmCxIhf57ofdVGYscQocpcb/RwUXah9Ou1KmUccVW2gcO8jtJXomXFjH2joymYi6TdL1p
mqaEg542RD9I1Cin1nVywfAx0pAGYrMu52PMtdUFqt7dCXvhsvrWUbsYwZSvvbBousNKg2Cw86nR
mJ61JRgEKvABXIpKktVa4J7bTR9bZkUa1SAIHNwR9jBFIekniiAeypKi0ddW4MCQ/snBJAPH6bE/
TfpkbQPRbFZ5mq5jOx0KZ375EhUlqMkwK9Z/vmILY8EroSLVcmpexFX0WEQgmfFKe0EyCVwZUtsT
M8MvXE0F0oudUFzcmssfT6p9PEHZ9oYxrlWPTdxczKybZeOy2el688LNN4jCmJj7ymF3QrZsjB+a
6t+h9DLoa0BItrgRoSLoxTBT3cx1f7DZ6gdkO8YHbYQkeWz4PmmWfjCvhcU2/LbekuDsbMisviWu
ue/vqkU7WFir/4+L+GFJBbRzPH5jqlyh8yfpH9Ti7Yb1VmMnH3SUX0SmrxTiubquf1NhN3roAtBi
9uXuyZGlWsHJI6oDfGzRcY2u3QSAegPs2xsMzkD7tSeFDYhkY0KZWQycFWeYje7jSb4SdKV7ePfV
l7Q+cvEvts0p48s1lDjp3T+qoUMU9UfgKaIIF7RNdV/cuxQFW5QSRkoTwxr+iKtDR8/BMZrn0PoA
fD+6SlId5p9ZOi63K3afTp2ppfqXi3+KjUH/t4PxM+mToL3vuKOXwjHwsOxG4npwqRutP4+JPJGI
5Tm7EwBrrxiTTbtRU2g6B3+Am2/yOH7VP8Ni38bcMlEPr25Qo3tvz7lBnYJ26edG8oVdhflag7tj
ULJIxDVEoOgL/Ch2uPIm3X6jvBhF4s8OXAtIN5hbzBL+MuABqDUnGnujw+E0M1OU71M9pbmjeHxs
aTDLlCP9XME2PeCdm3uVs+FD6wyUWrY+mp4hjhbyqEJPzPiNPkWvnhO94meg7z7Y54K0U1d4bBqV
kLLJ6+wwyjxNX6ytEcTd83Wia9V9Yr6sZJ4bIRsAza+PY3v4kQNK9LbBV0TQLoKOTsc4a4iTV/HM
f6SDqxJ+ZNr7etScebEDeTzxsEVk9s0I1ZPxWxROxyEnjy7SffOn+FrnAYfGtB2q41alrPBeIDKW
mHM5fvE8mEiVsQiqP2+NxZZPf7Fpr0Quvwu6d9M9uEN69deOlYl5XRG9So9kqOcnZFbgoyeZj1d3
jB2jxxKs2NCaOuf2K+W25yG71S7hfd0BwdSvOgsj/6rcqqR9dJ5JNjasfaqnE3MdKfr1aCwe/yrJ
7BjSwbHDFSBtAe47jO4iKoR3Oit9YaES5rg9I5c3FcDzJV/p85kz8Iv8l+XjsMpCGiYwdzjnThbW
WWSBI8A7adIc3vLUsGYdEYliGiu64IyeHkH7d6aNhaFG6M1s24W1D/rIZeWiJ8WNdVdZYnQ5VXGV
5v91PDop0SX8D8+kCwXASdMte14RPmUv+/E4YShuyzlT1NcA5skzCSbmXjd+E2RTljdHU+rea0rY
09bEblF2p7RE+7F7OwaA4jR2d3JxIjkred26A/ZKx7HaK/5blHNg9NAUARz1VdO5m6VSkFrUbsms
SZvZ6eXQQZgl8AlU9zqPcIFTESnMNMUgHN1tQcx82Vh3GJrASieQddO0VwA9K6DKaD9JZ17z95np
imlixs0h50QlIbkFBTa2ps2rfHENNvzcbUMF4M4ABk40uaJUbOeYGCZpxEtN9WhlCF7HPVjh4Mk/
s/nCc0yaddGn+XzYbWOQw7NNAnddwP7h6XxgFRfeu0ydzoQZlgOJ4J1I+xdNxBAY1+P4u3idkW95
LCJdVzqpFiEZcuwdSDxd3a3M/jCtQUlzT+Ans4PrE1+E/L9GQMCDcJHpAAiPf+LoMCGVd2wgCfgn
/5bKdyPlPfPPXv7/il/jiQ1UYog/z0So8XNr8H0rn5n2/IxTt/DBoh74JhQaNHS2Cx6jDrp86GZE
dX2fNG6ztyV+dwrcxZpC9VBjlug7ZlRU/E2BaoZg27q8hv0qGYhlQLhj/LygPRAig0nuw7NE/FEj
/4zL4JQssdQ1uaUUFUGOHKX9Gm85rm2McpNlANhb2yIDB8wT55oAi+sAZc3nHeqgS0x1c4EQxg9P
5YEQhV8mAL456wt6xN+50+Jl4HuL7TiG/5ac8iiD02EvfNgyTmzLhaC9TTjIY/7keUcpEuri6SK0
9byleX0q4pXkBz7t61jTB19NBNFIh76WCCCbLDtOZ80VbAzrUKdTUm6fT3kt5c7uikngKW3QQqHM
N2RaYmv2SCerymlPbp9KOuq/rz8YQ5Xa4p0dunC8K2SA1gbqXkfnGF0x/18Ygm/1ry0QpO/bsWJi
HBPn3njyxi294IOD8E7MXLn4EK7wSug9sSkW14fhgr2qGYAbjMifB+m0MpOzlX/leBnCDWalC09s
XkZy8sC+mfHLw3pksiynZrjNk4y/66V7mWo6M+uofNqJhoNq+F7uXQqJCVW4CXL5azpg4twjU3Nw
IFk+pW14LOJEyHPmR69GbpAGFXwgiq35LnkN5GF/Ph0jO9WZAtCIcy+BYZWKJdksCTp5pmAcgs0b
ZyBZNpWLNCPtxsJnDaBscfRK8iQqdX8mfC6nTGH0oahWvrK6qcG/smnLaMXz3EdZpZy0tCl/Zfj6
mkVJl6UaqoOTyiQMk6KSxNNpakz3JD+RFH27hMNoayT7SEPhvdfP6COPlZtJW4h3jsjRGaWkpFho
hO979Sx3636iWkTTqRHJ6k5M+msTlk9Nf65QSpo+yh9/Xd2me/HLiChGffMnJ0EbFtSf2CsUiUvx
aUpq8jTOhosQJ77E3YZ5YCcxu7J2khg+0gzkYtGBQSq9hjdUZfcrxlC8c1jIQ3+B5+HAUIfI0Enw
UPPCwSxbqm/9uguanMNmWVx16LtzuWfYkzczxzi3aS38TD4NCPQhc8h2Mlbg+qUswYRg1ucrBJQK
D8jRmebbdAQtf+QAzit8GNAsT78JDk78sE2wSlb/dB0OKXrXERGhz4KxwncgmFCK9eC4G2wanp2F
Xiko6Miupgs+tfQtdtI27Hvm2cnoaWsEiTXbCC6I2lqHKkU1PEMLSXNeWqIrFTrD6D1BQnOFqDeL
eRRFjI+ftEHYBaf8nM0xLWHsXQdGm056A8NWRGZh0+xic3tYe6EVzCFdtVbEdg7WFjUH5HCV/0Am
knwZqdKSc2RaoFC7hlzScGqvSyGbOHAaowvhqoWc6gktMYe1NcC4hpZI9NUxz94fH+RBhdZf1grs
nZJfMs1LR0mt78/M2ZwqFEKr5+hnacHiCpD6i7kkoNpFwRj8ctbEJTzXyXtlcedWU6uyTfxPdNP1
UILlBtulVGJJo9sHzUyjWiXbDfw8UABxJrA9aAs/pHo9Kx/6dUVKQ0yBbPijPJG7ey5UlNka7/8k
GSiW9hBJTB7YJKZVzX2mnaMoUlREmB575KjL2outyCuXf4R/BN6s0LAPCZZNsdBvVQmHlXSe9kLh
lV2/shgj3+PlHC2BGW7S7Y2HYKp73owNqrMH5mJYccFirVNM9Mnf0Y549Sna1swxGfkwexSkXzGc
DZUq+XEhFkFwlAXINEC0qfwgPDOy8n/A/J5MkXEfFZp3YNLLdbe9pl7V54H/g3GxB3d43HxvKgrb
faBt+hoym9eJv75YaE/t65oLUgFVupfvHN8/7qc4DV2L4btbU39ztwcCfXRNdelOGsjQJ0VqzbkL
cix3r8OzLXLEsaJyUbdQYtGYSfJD5gibXjpP2J8trEiEkiNbJG3q/lQwvII3hBSOn/Zs5a9qNEAj
7quv9iCPQ6bghuvc3ZBGkCZiCMzKIHv4qzXOK8zFu1cmThjg/ix5f9JDSZD0bhdf2VEb1B2DKwv6
moTY8mbhfR1XheGKuxpIwZO/kCizytCzfmrqPtmtj/BlZ80RVSa3qObaZ6wtaa4ZPJRVJhVwL+u1
+m7zeSj3lnYFnCqNBu3Vx+8Wt+mre93iHu2QYnkbksO5/pqkuVp2KP/n5nE4W8FlrMPZ2dTkvWw/
LZKP3asDPly5yKROYvI3BCZFineumI1gchmFVyhsOZg5itr3EIFTHDGS2w2vTYrm3s+lhLUuT+WI
R6/jEFlfaq7uDrzV+QjoXUqxpyXJb4EWxtvD0rGI+ZzjMYv9rCRis9gN6iI8GUcpp6vePL1DkWY+
NUkQNuQ/4txLm1IzJqG7H2nmufAYEqfO2kTZc/O1RtR01a62gh6hdgRICB92E0iXuCDVmeBEkdHW
5i6D9BFgvei+g8CQ9oJPr+RcgaA5wksS+Izwgj+RuRR3xEJQBNeyeAtrPC5jtZzf8Eb+8qqcxveM
gmA4MmCDagJpKJRkkPJyEOoQ/pv73mqH7EstGUipcYlP1fk1gBozUfj5YYhXnz9bbOHB+kdEurwK
LskSHfvNxMNt6I4d+k6VOdpWYt8W8XOGGR98S9O12fYiZq9BLN06l0R8dlahmThzpocxaVQEE1I7
XjRQGZJqDEwj4c9J32c5qSh77CVc8Tbv+dPwvwU/n2xuW0Rlq6IHEHnWfbpZyTaGiDbTE4yn+GvA
l9zyOT4ePUhx8MrpTLhhJo/3Ry5wPFiXS30btmCbNOUCHigaR6zUrel0DhJMsMbCrS/a2NAed9f3
skx07iQGQehdUw843B6KMACROd521nkZGl+TROIIoyZKqk0PkkL2Cj0vLP2Tn+ECdmJCydu648rM
GT83h2PNB299YuJvabh3Us0GGKZF9M5QpEa2W57EFyJnWT1pVe8BfhdNDU+7jstNwLsoAvhCgKsa
UtaCx3ggSBGi3d3l8Op8JUIpzuZxObGit/2mhsdw3xZccrKFO1xs5Ec5wsfr0KTQqI/0/02bqnNU
RcmmjBPNDGxST6Aflw0AKNrDFSWtHg8xk8JvAKvP1veP/UauJw9SBiz20iHE+9V8juj25DFwO8p2
9LAc8N9poVauArMAdRTVEkYAktKLo3Etq2QQmvbQTM8OIOTsgaUSwsmtJdFj4woMeGQq8XjziCzY
52ROtusDjV8whADd43CVKtwQnJdgNEI0qUyS9pLpDs3S5U1FgRcfT+08U+EDAacRFa5dOoC3eTu5
6BhF31CsXJ1CRQi6qFt+HRurXYRNRORplgOrBr0VWRlyPq1kTcKQLt1oMepVoN407cu4K5l6YDE6
x9dYXwlGTWvlYMiCh43YshPYsE3r6qosDuwE+Smcea0sHsCtKeCjjh8j6jlyyb8a2alaD4vM5lc4
geFCJVQPH9kv4bimEB0vcElWuHfmzt2hh24TYhBA8OT5hXmonyRGT/nai26pzu7qnmWa+YDUoj0t
OFBLGCIApAd5qZ1U2IwNxW1gb0yfGfFIhSj+jFnm3R3FCZQaVFdhNKzAZFaYINJMK+lV7pPDxvno
KXfym6mzA/UyP+PHzEbkh/1Av9uJONLoR7poVAQFbOBKUJ85rFOf63hQr9/dk7+iwjktbwsZ5PbS
iCTSs4uF1lrj39GiuuGQ7kVTIIZeEAddGeL+B9KinKb6FMW5pba2kDZKWbc63ML9b3lr3REvNJmc
YUfgtlK2fBgRWthmEDeF/XP+JEwLu7s8PvsRjqUJixxksY8obX9HCJ4OxRnNDJTUJ8tXuKnQU4cb
fQHs/n50nhUtjm1gXF94z0zTXodoz5IexXTJAm3PMvoMIUJraavo3p87WhhW7Xfn6xi9CEjGGbMY
lYgc2gQb7aoC2edwhfMlwwiDG8yTRQBfCb37TOXn2sDshbcPF0SeNPwuvLxcXSWQHDawJbVby+Xq
0xppgaj2qZv8zUEuQZ38ISTTXWmCAL0BT/PD3VdFMBiA4QVF6bZjMZpGzvZ9SY4VheDh5zuf43tI
1uOP2yvOFYPYYxvTp/cbI0h+RSA0RCxyxTzYRRu3HkO9NEkdZAwVSp/g/uIElEUEQi7xfcSrEEy9
WpOcxVXVcQlomM+VEi8AZ2ibl4Lru1jHAht7mojxnk0gFhsZvNYXHP+GaZw4hveKwqyqi2FqRCLX
gqS3mv36J7Ii3KRe6j8dszTnYbOO5+yOVlM3/TMBtinqbFNsV/IF0MgYapcsoe9sMQiGzhXBQ6Rw
/oX6CGv94LkwH9pgMVU82A2Sqgzopr1LtuaxQd+O53kldU9qgs0+f2WkL9R0VU2q68qMRD2anqGI
F4ZEElBnLi3fIslbm51uUgm22f1SniAJe3Lq6iM8L0jkd/4R+44blSda6HOGw8+bnejndQbrgSLe
HmFdOX74DcS257xft+Pze/h6rx/2JP1eLUsX7xUgH6mK6QdSpiyvxci05UUlH21NxrFCZUVmyP3N
3GjXgcoFDTSw2ppHqVcciXf1JXNxAMDJHnnw2SphlZQTZWoLUSByokrbgM8p1XH1D6WSJD2le7nZ
a0OTAY5Uiz/CffmCWp2zdwvEyjphkRRb/M1cLzJZpYjOwc+FyAgKYca4f4kugMJziD5bD0XCAv3n
22DercDmvVyvEUL9LTgrnuQPPve4ufNebku6u3Wstle5ir5nVsiXcBWr0WMEupja0Q7W8fXvfMi0
20rFGjS6vf4/hk7pSao95u4Oh3HyH8K/XGnBuUdJIb7xoEU0M8iQi+Deu2Iws9IgmC656kiBGWDj
fUnCpfxNlncMiQPx+5QLif05Ad6QQH5Ot4PEnaZ7lWIMuRqqJQXTib3W6kWbCbNLkwIZYPaSS+9e
7iYVWhXhVk3TbtITLmccFZWJdmPjQbBTFM8Y8e1m7uuMqnBMm5nFo79UV1TgwYEcFi3ne+xKsCAG
B7HgsTmZU9PQGYYdYtshHvNir173nkqupR652BeAkZiTAKv8KGEV2jsRcqIaKWZI4AAN13GJMUlI
xap5CKL1qXDzqTSCn1DcflyTJtsV+WaFkXm3lxpmVLDgPpbTpf15n55sb0I+as1FHtKFB0RaeyLs
KZpq5kLZPy+PpWuoFYrU8YcKZ1cGr+9Ed63GQRX/7GTUIhh0r7MlRJsISGDlBjgnpdQtAix7eC5j
Vp9w8gEimflFp4JNNCd8KJan2dAV+rFVWJ7i7nekE115UHkhqO+o3jZk0YeS7JL+lw2SGSjHUFml
1sr6uVrlwZyOwn6P78iVch75incbpOYLO7wf8Mkubryz93DciLskmoDqGXZYgMFfB3+X3tjIdkV3
4eGrYSw7SDS7X/ZImzzyXF2r5VATbdErNgAzgzX8IBoXvFvPbtm5D2O/Av94WoTw0OqztW0VLAsS
yQuOu+Uf8tmaqRCH0beD7fKwuSiHY7A56B0n/UznwJOodkazH6dv0tbcHTy+HSNqUECzQDXglhnm
9toqRFF3tzoiyiJkYTYW+ugp92Lc64I3CStv/BfjaUCj9ss3HHRQQT8K07IcqPO3KFfQb2+6VwKe
GEtybPSnyu/PXGXacxE5hXASdP5ZMTyFvZ8D8pxUawVUA5tMiiC1Yq8dKZ1rMeuMOZoQqeTJYym1
CDxTxJ/VzAkiqpLodAEAyvOHxHgk45DO7dwO8B669aFexaxDgvYmo1MlQnfmYNX04Ph/xNAbhhVs
FMsQvFQ4DHaSXtZUqxbGzLLeOVCwtugJ1z0AeHilETvYiQfYi054dVeY289e4KZ5yZIUYX1XG1vm
/MsZTGtZLqeqdAZsFJZ7npc7abkdsrKZIps2YxD+/LTPxLz+enRkp/eFUnDVTJai9JG9VrQUAuR0
rOklBInVHTeLyHrqnJhJR9IM7Y4ZmkTYlvQ5/Kp7p2EmhQphIEwOHHXmoYrtBl9K25h6STzTcAA0
+DrCMDZDK1ad5cVuWRZfdCMbOu/cT+kxL5OQ0WURZ2kY/tpFaSfmd8piC4gVcMlIw1tmx3BtG0HB
xbQiqAjWYrri6U+JlRAyPmCTBJ/TSv4VsCWU8fA+z6xMd1LUkOZEvxYQRqGB8Fy23yah9fTC5Xeo
YV38LekpZsDt356AHQ6Iszi61kPw1D3ccW6H4aB0HB+orcfkEbhx+2IPFDPgEUOp31XCciBun4M+
5m/93mZ+xHV09aLGEKsX7gz1LYtNXPQPW5pU0QFuOuL1HIBgil/bqwdXOmB9QvHGREYL00uSZkAw
HgEnZChWmL3e0//QO9D24Wd1ORWL6Xoa19txYxyjDscTN6iZ0vlfDtZs88Sr21UWQTqDR89kT403
UniIZtPtlKAc7i0vi74qSU9zyCVyM1mELHY4q5r0ulF1nAEv+winAeVPzcasP6WStmIjnncbiWxU
5xC2aU5T72saKRKxHLrXoX8Z8x+X3vTqG1bl53UELibeQHqcytXi7uhk8mB/9GEhEwNNfv7ZYFmI
c7kAmL6uYtqAAVw2eHOcFohJd24Ofmp2UQgtGQn0X2mfEzCuuwJrAffTVvsteWgA5bxaN337x44C
1LJQC+FQHjpPQCQRDSH3ldjEU2jE9vKidL4v/rxsnzuPpcb0AWsmY9IjWPhfC2aQZcYHNcDuzTFU
M92oOkBOs7mMv78j5jUg0H6gKL58ov0+/NniVOhMLLoCIvE8XzuEq/Z9w7yTTE/hDo3nONuTMsXp
sGJPq/OtvrFXH0EDakTshQ3h5JDWDqWLuYAT60j8c41TH95QASjnn7mR1zb7Q712h1lL1qBp8yzL
Q+h1AyEef6Q8y8EGPY04DTjFYZs2VDhMuWWnP6C9Uu+btYDdSbWno1PDHwVlROLT6KH6Gksm2Dj7
pRmflgfIl88ZbEDYGJp7AQJH8BQJm5HPirkCDUDQMVkls0vb2gOsPrG4RqWb9obxNVGUgX6pl1Rr
ZXjYOBWqLMtwoKZz73GuyjD3ZG+AxIfPtbyH+VGZuGkyNV85iyqi1AiLppw6zie27a6iDZlfVYOz
NtNo5Ocl0v37wmsNXMH9rs5amIW+KNcJV6CxLUkCeQsVCaYfygw9K23gRZSiqGC5x4PYMowqrVqp
fbwH/2Xf9KXFfcEH4f4qx9S/EoqHkVu5U4tWOZwPbWF/wWyayJEb3aMdC4WCa1KageyC5HHL8kBV
jpvIMitKzRmkCNNl/7iGtUdTGX4C98FT/+DMsUOz4x76oYp1gMcFs6dQsLvh/tq3LdqNwqe1zT3U
iJKHf3GBwsfNmplE+7kILsc7B14a5KcqHcfzHXz4cnMC2iWiCGaUE9DTtAM8GOaRHrkoWboar7pU
uRTNNKFNdoTXS6TjsVrlrjvk8C81hAy3y4+MX0LlfYXXQIoIgL2C0IHbsP0RRb423JpmR0Wr/L1C
kZWCLB+0q/YGOKBAR8OM8eAYcSFmBlTRu4CzsypE2vU81IUhI9ftckNcFJ65gcdfOCaaNaE+029s
nKXAQ+dfs736cDgY6394ENt8SqY4BOrmxqsHndlf4jtItZ2+h8boCJBeXfgyJo0eLDQh8DxfsdoM
OdRRNCfQ6RfBBwZiKfhboJgzp7rVB2/eGPhVNHx55153tIUbH3jkTJCjU5pqwP6jadvNNOfeg+WG
fj4rcqA8RYmTP/hpIbebmnCi0niyOIYgHmG3tZPPFymwLEICAZ5yEWyUyh2Cf7BiW5aBPY3L/obO
uIpLFMvrZwK7ELuftx8NkGwQ2HT6+l93Qi6+uOtYvJIApW2vqkD85Ve58ISP2yOA9RRmvr1VlXQM
yMAJrcqzYNPozYeKSrHm/fCYZUJhaJaJC4Pa6pEWG5sixj1irW04Cx1Erfkt7A/5+/ElHrlABJ92
fgZSjWyz2b1XLfkkmUX6ESHKf9yq4VTzPpv7dn2KLE1WR3dOpqXibKghTS7JW2bMP+Af7YZv1LMt
X1jc7kRYs24t5l7eL/4Niatn9v0GZ0SxI6niaaKiF6D6EOnCcpfAidLkKKQkRgSDM5hvFGEZrG6f
048AxN6jbj1DweIZRRPd90IPYfHgivcjLVo2bGA7NJSVRBpquaCnK6nl44aOt/7/GofQUOuO9D5s
nukIkIQRzqqQ8FsftvPnWGTQzpAEye+Vsl0lokozHZ1txQRqI0Rah0YBBu2UNJcR6YQmJ64A5Szq
LAukZ01GWPoqCQBUKSRLhI/mR2bRsoCOwqHviqxsA6U1xTW6WXCewVmRGNxDZgN81ted05BeuvO2
vm+zKGycM0H5QEjRsg5puBuWBZMR8Djvr3NBqca6bhjsrC5xUjBILteWcWcO1GZzszipEcNev5SL
fwVW8EHUmnthTfuTuwmAR8SkFMIWH64VwSyK7oNViSms00V6SlmwL6wT1jOA8S0RnwZs1s98L95U
w7p+uZcAFhVJSs1BlW2TofTDbyzKe/161+EaAPNDcK0/D1eMXsT+96I8f1ic+PKkyzCABqEdwAfx
6BfJubrRI0P67pRIqgzOGGhmO1qMOyKs6T1dWw8p9o8tk5324RgCUzCNhhw3rwhhSxd5QR+ImsLl
1ADBUjYruSmBSNhIZmmgGOBOa1ddsfLzNuInw+SSyfDbO8CD9NJ9V+4WEEwg5tOhZY6x/PPhpvQT
tcuCw2rFI68fAoaHj2UuyyDJ8+HFJE7CG9BXRlgJKBm6Hn676TUv/6Z3kmJ3rBd+V986xtwOEvCu
og+Y8pIOQHpFauWMpOp9Z4NjiqvtAZhuGWjI6VxfWdzsDaN/fHDQ5VXeF26mWy1c4k4lE0tSnwm6
KW9ldbtlsu5zGrRF/glQcqJKe84niGDHjSfyK085KeblMu2kZ9c785tEXWfy5AeTch+EILwWEdb8
qvKY+rFIfl0hmkBRSEAx4JTrRnMXpRj8g8BMMP+B/TjzTiNsZjnKN0ez4wKEcOCawSSHj3WgyufJ
wURPzhdY2yEXU1sj/4Bbjz4g1l68Gq1KJJ0mvDOsJWIrSv+zZ/AIsXAFLKOeTdGtACvtC25kovXw
FyTtJm8/PrMr+pw0YS8oea9McFFLARNLNYCO61QIjGa6Y7aWaScUXen5yBw9O28vjamK2d1c0Lo1
JP6L+Vyos5QYHgykQOx837RtxwFzyYd6wM5dgdm0yjHxcKGIBAETnCqtcR2dR74TUIct692m+F0i
vux84CBcTk3fdToq9oDhhsGR5QLcdeUDUVx480QyqVgTzxTo3AO9Hrndh9SCL11dmbr5LgTG/xG+
GfwihAL3yN9tS7CeOb52O2QUk8EWszPsRjBm7znF1rp7cOUQQtHI7Z/d/SfwjPU19i2Vg6OMjaQI
ni3PmZ+x5+EWj/309i1CNdQKFkym7iI5/xsVrynHQlRY1TSBmmejSFI8mxHMYHEPfxCXeAeLszjB
RtB8uZzLfteX/xUtljUMxllNrnSalsTm0twpOITl3WRDwRb1rDB3msfQUo6B2JAinAeTqtQQ6ADh
inODyuPcNGlG+5WbKuo/majqfw5iQxc9/dg/noVmYcs5AG312ojRKaC8FEi6jkUjcsMopITgXehQ
L/rAOS8FCdxRJEuXku0biE2IR2G/wQFxxUw3jUjPScosHpFLLF7qEDCgCS2AVa7AeU31N/reXMKD
IrAlxXxMxtdz168RNeJNONnUJeM+VfBAgYxnHeSlkKYOPeJALG/uA6+56TVW8/t2fbDoVqEkBF+U
UeK1L3DMOOEhjwgdq1E+sDGzdRI6ITSsEtCLrTMzO2xA52+cQKI0l4vy41Ry/EN2dSfMjySGkuXJ
6RXLCl5BTODdAEQkGl/UQ1RsTSkzJgbB0BPrKXYRqmmsGzOIIsahdPrAeQ6RMbAa2Iqm/G0uy+Ex
1NRPfWyJdI5LMPhby4uwQdY552VSi99zrxu77xrIKlXzEHBwEDWP3AXsp0sbhaX3JDdbn0ekdRss
qDmiIUO7fX0eg/PhlL6uUTK3xjsteo5pYsfA6ro+pwBXjAweGaBJzID7GI/JSm17EnkeL0mAJiAj
70kzbpgL748SnwQYIuDRFaT8ATGLZ5+i11ZXJWA8uB3xklzdpKAY9riJsFXtKBaveHsnWuRh+J+U
sdSsfFhNM5C3kCc9SN9aDygBXy6ROaSS4CzmxqfriLsUdUHiXTqAMWIKeRkN0O7FpfyOrhTCPQlV
LhLOQPeluyCqWqyNHCwHWbgGnYLZRN3RSGRlF7wYea5WWqTrnE0Qj0oGSzczV/W5sDFjP6BGe+PL
KYhjRgTNVWt6SYJbh1k7mK5gDckr5Ew+K8jrDSo5PE3E/shn3M1y5RTl9q/omqkKBKf/dhL4OGvG
QI83JpFSoW8zuc2WJqBVx3q8VphoZKCr/UnXbBSAn1zsrPY8Sl0aEqonpe8/tGVOsR6vviLq94ks
BcMdEqdP76PZ/uWD3ZDzYpcVi+3vLof44jCi7hn4fj5ejIGn5SPLHouWdYwJqcFaiwBAiFptId1l
aWQdPgbIVeom4kw1ut/7GIX+eU4sG/s+kWTz8jvouSeib1iLSnrCAboSfNPGzv8/q1AzFiPEzccY
50vPn8O1DTmS13wwoSFS8DQtrcqMPBShU1TRunY3c2UVa1ZvAyV4+e4oLemrXJMHHs3pSOEIW+wr
B0QrIu0aR1V0RBcg8B37SdfvU9taX+nQpiXETQ+oLvpQLij4CxSqKrJii4dKjPRjJxbo/Mwne9sg
nrLQiwKSrOCDJoAE0GvzpgFm0GlLzcm0AbmP0Q5TEk2P53NKYDAhs2Zg9BMXdXwoxYKmmi+wggjn
NIvtCGDgYWxZNSclN5HCyRFn2kCAZLqkh68HyFT2yWvvsbt1jMMIT23ZEI0tUrIW87Z1OYhCG4Li
22lDadIuN+QrkLoLNjxXlvXfP0FvLD3DLnZguFwBSpe3PSNO6F4q2Ky9DqxD1ns8O2d7kwQ7QEV8
/dpUfQvPxi1xNeXX9yW+XTpvVREQe9MMazvjfrTOlWaFtCMfoijihpYuYvyhEdKCE8plnpm7U4Rj
idP3EJF2tUcc+o0JKFUHtk8sibgw4MJhC45ZAw/Ms2SiMEXQr8TsfPutUwFXL+ayfKkE577D35Tx
lZC6pMXeHSSnvi3V4oBywN3DB1ZViQYYZWRd0NmuF652KCW3eOQz+iJLV2cRFVti3TJ7ak7/sruz
uOaj75pqhLCfFfgr3vPlzAuk0zcQmmWg27dgk8EU3EeZQhISWLItHsLJxscmXWUyj6Yh0xQBdwlU
xEU1HYFdhndg2QRe1SNtt15/9Maq9a0SHhZe2SHTmR8M+V9Rqey0ORTI2UHaqZLag2r+IK7EFtss
77gewLdekSVcd40U7rAGaCW1ORasdigCEZjClgD7bxkL7jcRQURH06sFlNTYOFtIa+qszC3JYEoJ
HuAYHWd14i/2N3Byymspb33dDKucZ8LvAcn5l1eEmxQjDcvWLr6pSSHkHj476wTNV9w6PJn+xgZU
/fddBu+WevIbewd0AgS11Pg8lKUutiH80hMQ2gcEMXgyaJo1EVOiOx117OIUYJieRa30X0w/LAaN
M9bea+HdJseOyj+xGTSW3j3hEtr59iEvBa/sdABxvX44uJngfUOdBuD16QfQZO0Mwg09AeRSDpoM
ZfJKSZqvluFE421yXmvwEg0Pj82yl3Ggd51g8HpHOUTexDLBfmqh76NZp+3nFaeXcaA5QW7T9Xhk
rr+fEU6vQYvAAqhX5GCRnue0TvB4XTKN6LVLu4hqQK6ADR5FG+gCMze/vYrimx0YxEiOiwFq93YS
bKlEy8zO7e34r78xwH1TIDwtRY34SyzSUXKYSCkpO7e1eclm3dzFttDwY1mCdxXoMD3EAOJK4ZF5
5rPwwUy7tWfmpHLqGP7cZx+NstUuZZI9NQcPINb2cBxxhgORCYTm/vqdpTM/+koODaVizFpDVGQb
6VxhmHJFr0IAz+kYpzlzjEe28dl+kLFI9fUThY0WVj1aMKZ2hWcnnRoCEJ5xmO0QQaFPsp9Cw7HF
F0vBH7xCyr1SI4p6HUeSFAc/id4MYoBWTBd1zVaNDYb01WsuI+NTGmY3w7p01bdGDl+SdfF1vtHM
GeQOEmztB0JevJ1b5FxaFx3ZQdP9Z8KXpMqhk6I1ulYti5htT+Rz5RXC/7v12WKa3VhBnePJ83J7
mQXGQHSMOg3afOHNG9JgVE3xqhQPzZ1RbSVHeSdyCklybOkA/0/QBn1UF1IaIyaNRT75GzACRH/5
G8OIm4ubXTrUBzNybUhYFr6LNi+JrS3JcCELhur8f6KxL/gmvvE8GwF9x/2JDyPNJIwURpfGm0iW
c62QRrolkoq8pX+RQInfRalDtAa1dPD4ZDwG/lBo9Vn/r1Mgz/Z/w34HsEuSeZYn0v/HZiLzpVkG
SYqjHYKeHW+NGFuRitARh2wBccYdPb7iRPws0hDnrjd1C1d09FhhwE+J2imEadUPF2iFdnz7qY+B
4c5pF4w69pSqF/Pg0NsQxJyGfueuKcMYchW3hAn9wyqM8jGBV9Y7Fjz6ZttqnbW7NMEJe9pfqI3T
xHmQ3eZfvIOF23jVX6ykmrDQHgEmEyEwxFn6hA+BHv6baWm283D9CmWxTzMkU+EvzLKEQeVCUmvw
zVlWRz6z4XUI04uGXNnP8y303QQyP6Qu0wfnuATMQbu7NOaCYP1xIGlByPPQQ8GpBoQZY6pILQTb
n6OQ32FHnOM9Gqdy5OD4SWN7LCtve8sexxJ9l+/3+snTIq/rh3QXx+YUyAG+UfnI50JnLslqnHNO
cG+rLva74IVNLUPKuunfpkS9PI2GQIkzLnWolNaFIK/erWVj1X7NvFGo5C8JfxCceEP8Jl0tzHPt
9vWKQtKLy1MhP64w726ms0pXQ4cdm9J2rhtNCmmjs/tOp48Ax4YV7z8v7Lq8XurXIv2qFsd2YHp0
1OUvfvDTV0b/TVNJk+7ZVwhe6bC8mswt3HRXKzY3txG7aj2FcLU0FwaAdGb7f/Jfhskg2PJeKs0z
dCkLqGuk9YLmi7jxwplmzkM+muFKJg0a3OR/oPVDCt2L6lkPPYCR6/P/xd3QyYLYYTsAivXNbQxC
AhPfju5cZRBnN2L3THU8muPm3DtmK3OeoLNfJYoBXDf19blj1F0/8Lv/Dn+XTPxySMviLc3Dn7aU
yxHvCcrsU5/ninbQ9ByhGqulaP73dSAwcXcG0NwJ2M7hxS7GHRWAjMeTA7m7pq4pi3BApbO8gAE/
hWEos9DURtMShzihvMOmBqr4fMAGpli6Jyafvu2TD0oOZkYBcdZzEK6SvCSHZG6iqgfy+JL3xpQv
ue8fOjU8eqEsD8Zzdu42NUrk4Wzjez8f0XhS3S+w4Sosj/OFX/wgKo4ySRByG7VN+KBXeTj9qbiT
/UVECF6imDqdKZJA3ys7MrIVK9q6ambO8rPQ3RI1QKFiWBdNN6yaDnq0nLw66uLJLPyhQsAGzzMk
TtXzBMAheCFfGcXRr2FW7ML8h+LC6B4K+QvlRcpAft4AzTfJVQFR/h8ZZ0zbsvGX4Du2Zhdc6QXY
ZF0ACUhvtdo4SuLQpabRW2cPEyS7NbcpGR+xY5X9ZYzAkpESYzwe9jGIMs/ggjKtlE3aUO2+bLrl
otMolY1h3aVn86UEVdcrAQeigPbVRPIXS/+eA/UvTPH3sKof8aLgpMd1QkrEoEEUxdi1I0aqnTuq
lxm7NEgK4bSuZpS9uvIAZdFPRHniZu2wRo9xzOSKFuxpTlC96PUtcYYiNAdA5Dc+YvJUl2RL4eoT
FteV0e0yrK92jlBzao3BJp2oxIOKtNnog600Y5rXsu9uD39YXTcU0Ab/v+4+6zF+ZfbKxp5cwD2e
GderuaSPC73It9Ghg7E9mKRXZ2kADSTLvbq60n509xwChznrVsY4YlVYwHHeS/7Rgsru9gUjuFKH
W3id7Hq7qziIc2wQHvb0bAyRz9idljDxzipU4ZF9KyW7O+hGd9JGwe4edV+2zswKOBrNF2LEx900
+J1mn6kpGi2KTikoSKRJbPMCQ7ZsNR9nTPQp0OMJ2Ve3AszLHCQTlJz2fb9CGN+CGdnTd4/gsUhm
pEK6Ditt5/BU/mv7XFWSMEa7lMzimXHgId+n9ziDzP8dmUe8HkdY2DuI+BlxbMF+PMHGlm8nUea8
bmSuzbiVTHRxNd42qdfxln9NYMOsv8qztc07KALM1/UNBv+Y70G7ycD5CMtb3ibxlp2Gjvb1lvxf
7/S6UZrDtXU4sv5QOmcTJLmDtbnHS3JUw+lCHX6mJ4qp9qPVR401+rNKlAHKHcePup0KIj0HTapg
9MkEXm/4uj+e24dQglMY7cWUlqsix9uqem/MBgndtffZCMtCvYXGkYJb3wI8v16IhhQFH+TCJ7+S
16qb0XfAeYTShdIYIFZDgk826VyM2hj91Wv7VwE5vxN8XLPdbqaFU4rTqO1t8YjFjYe9tLScrqu4
lb9lgAfwf9UBh0ixPP3sFuZBrTdrCnhX1eWo9MLZk+Z0YzdPB58hI42D/hsVgtzaQG00KPL59QVM
yPYWTT4AwFDVJlQqo8w+ppdng8xzieAThxktl94mnSe7vu1QYOLsgUK9bsRCenBd5ltmHt9JtfiN
X4tWJ/VMnfYKRZHBteicPNHloaFIlgck+PJTPZSUluuPCxMnKBQsGB0A6LMcwCI8YGFEpOo4ihTM
kEl58X18ra2FcsOivyp6vO0claHf0kO0W4ZdkmAtE9dKlkbi1IxPiPZ4QYz2lYEXu8VtUPeeIeYL
NqRF/b8Tkr4rTTSpvHG/EWSPWqf4HGUduj7UzbRdDTyi0QhzuqUoCWqi1AJmvfKthLpYMdU4o9HT
48/u4h99JIVvTyQYFkX3HjVquhRGjs4HZrDrnLYWLuiTNBgMmQD8Re90qzyeXQwO2bVI6a7qbcf1
3LriKYv9OWF4Te4wUwkbWUDPSLf/aL5ZFJQRepR9C1xMh4V/WGRr7sj2j2BpTukJtWY6T7H7BkMr
ZLi/QT5e61YFWTy9es1KOBvVqfnbnkxzbqWi2d3oa1yTTE33qdwh+vkisCb/fFaueVGbCDGO2N8T
iG2mUAlj9H2NY78FKBGemG6mVf5CoaQ6PJ2DJmQu2BCM6BwDzXVWXmFrBrYg6ELUvHtwDiEXqlfG
NfRhYj3zREBcKGPVjvf6Qf9oJd5Xeg5FPpAsOc7oGXbYzNwAG3WJWcnFefWyGkowuKnmMVR3JAma
AAehkbg5mVPKc/e4PdadaAu0sp24Nzhr+HCBf8mU+EeaYn89ysWOwqM9s1jctNSCs6XiOFt4PFOv
yt/s8zAe/YKSV+tmU7AdAO4LYzQLXlCgIPdW3YozukMzia9q3Raujfx2Z1aBih00gQC29DriDS5x
sGQbeYyD6BFDm879r/wCe7foHQtOqEwDBfIaK5Bm74Uuj/JsSkQYGJmIldHkhac8AQV50iSzg+5M
DmeKTLxWy4tQq25+12A6VbicdmGQDVIC7Li4FWgKgPGLs2cQ8zIF1jKPE9hxj6Urza0eSWo0MMYb
FmmciVubxGUGhb40OjdpvhqlmfoK2fIZwQn//zs4SEXXk9ZBvN1F0+SRg93MYSOiWYA6Tnuc+pqI
ItcQYCTW6VYYKKXg+wfcB9cM+vXtFaLrhlWq0Lsv74WqeQ2LEvQoIgcyoh0ioJ/wKks0ZKNcrVbh
bMe3w6iMQqGcSya41BZlnfWR51IJYousFHz0ezRcPMusxTNeb8i5fYlhuDmV+oe3InVkLczR1Pny
STeQjFHjvxK+gygHU/NHVNq3G49uIcVf7W3HSw5knF9zMQbQJy7GWfeN5EHjOlia8xy2aw9R3BNJ
XWqI7K3xTFXIytdKxeR94YdmIJI7aza+RFdnz7vxZiLwt3dkVQfUgvjC9J9ecL3z41wr79PvuadB
adm/A0WVZkkHG3hWhontZH5/UKeoWKcWgQhbZmZESLI8hdbEjYs95o1VjEaTz99wsWZu5zML49xm
bFbDQwT+B4R9je2khgnpYb98GVUoYs8CY19A1CVA49v8dLNmpxgAHudgrKYdxQZfFf2rGp5rK5NW
k0lnb1Sj9VENY0eEDnuc5mIFjDbynQNGOiBpzcvIrzgSx+wvu4bvhK/9NRj/F+BxkbOW6+RaHx7H
IGtcsR6JhANKwGlz8OsyZNdg8VWuLHXzQmFYsQSL2uJwbaaaWAq/UwQQGVXPN1Z6VcIXr9+McUry
TIyKxdNgQ1V09b1WOyaxLGNmDn9uzq9EMQE4Y3OvRl5JmI/gni8BfvZdXNzd60R9q0FPhx/8fCP6
i0nzsIvxpQl4FXvXSOzwvPaJ/n7bQBuXthzF49csUal/K5oxpPmjzpl4RbBFdcjAwUpghOQBZsHb
NH5sUFQxUC/3r0dtpzvyvX1VPuWw18M/w6i3qSTwKccG6bVLZX0Fxn87lzm+HquG+w4o1RerlSVK
BYcGma5AtQIyVodQr51SOPmE6MCgsHgs8UfKgRgAyd3uTA32PTk3yz2j5H04WxT+re4vlIORgB78
SefV2va9EQNNspHzJO5kvWxyyBvkBZyBvsg/hw7JHLpVBvT+JuAcK5zDxR7uzxbGO/yz4iWG0+NB
/G8XyISzDwVg3pLYnfMyLvcfZ9lwX6gIv33OIBUOHrIILmoKSD86MbhzUXiwlbaiyDFazm+kpYcK
x+y3i7CECgjMeG72jzMWrO6YxJJvCmlHw1YE8oS0mhECsucBLj21G//AGcTR2OZKs6tcEOuQo6Xf
h4sTRHtX4cpH7F/e8hT+gQhJES1EqDauBNhdAH8RcRWnmoV5ShHu7chyTxLxsTUAJAH+KNPef4ug
rqQQAP6MgiNqnFOfJARNPdWTPKMSi7epmp/4q1lRHoEzRlpv6e1RH+2GrQgY9i7FlT67CEtDSndI
RBFi4o8qcEZis8gW3n4IjiHV2/Sg75K3GFT6wSx4FG0AWb4IolZ2nCQRdmvaq43qhKTjk4uTXAFp
3zIZFebDGOio0ORyc8WWY/2EsHR1Ouw9hVoo5RLIsBMuWY8C52wM6HKqLkJQJ/+QDwxLz664+a1L
dGGpJJsZ+UpEepUdzrH8jjTouWUkRBQmMcgpWaEaBi5YYc0sAEYEBHf2NJ2mCQIEYduhLlgmtp+H
WDRcnbgSyf8G1byXGPZCyAuB0xXAcxn5n3nOjM58lckEoCxdeqgcKIQJarxST9ZYcJbavqxHeXhh
YQm6RvvK07dP6CagZ0OfBLUpD5ZQ5FSIeOTMxKtEtGfEGv3R+cYvK88ebBhjNhUclxd534RgiXlE
3S4tQBSLUNrZjcMg/WMWKefgN3T2T5xEj+4iK5a9O+6+ZQoRXyVz4bbmsiEk4kuEodhW2zQUzDuU
V/5k10YHs4BItB7PCS+1NTKHq9uDN9zpvKGcalq3Ooy604d6rPQg2ebV/3o111NfsPCBWqCCqA+q
GtcbM81Y+rtdXxDPPRUisSzOuMpAR/ATWf6uHme7NZ6/KsGTr9CHp2Ga1RZpnOfqhveKvQVzB37V
HPyCUST4d/rLbyFbeKwrAZNI0soVMLoWNyUwbu2ozP+4i+gbi66WuiHloct32vVOmAQOBHeA+70C
LnkCEz5W9yYvu6IQ3zYgZfX1y29mhTRFN1BKeP3h8LQRb5CyllqS+gZbjWXrB0wHt4/9SBMggqlN
hahsFkmNT9QMDoT1In0HwOuqC0bqDmE90zCe6fkyeDHgZAm1mUUc+6omQ4VEWW1ixjUGHFy01Za+
TucG0Put9oRuvEl02JzTblhqQJ2TpaNtxAD+C0F8M9AjmRz0s57Ig+hiufv1clbBa6mbIFXWEOz8
0eXj9z/PAZeaaBa9ekgTwITRm6eHI9VfVNBWP2trQStSZGVUTBtE5MeORqqfmtbDWX2+OfF19oDe
64C+siMTcUcTphW8bNtMOG1EXRb73jOd3NsIzpb2qdvea7loeoRzbK3aTY9zazsB6nOBrv/IyJj7
5ks3eMCsCLjs/DYRR8Gz382ftA0qEGdXLZNamOnIg3npVUw+ZLKUeucBWuHARPRPFKsS31jAFN5z
IOZQ8LxjAW+g9dpE+gkSx35Cf8T4wte6dHFIoLIEzIE8LhduzMzQ7aDBroaJM2hXOiNM40W59CtP
WXKN/ZcudX7k2y3W677iBst9cpe4txZ85lgO40+lagiXonELN0J/jtPx9Y2V5Khj3HTj+DbxAqsN
WhVv4juHlRa/h25EmvC2M7ovJ65zeQPecGcv82Dyq0oUYV/bZ5LRhUqZ8t/0u3XrbsJIdTqCZaHn
bf07i20ULjBd6RpD2EYP1qis1dpdU9HtiQkfP3SYSgE0Dqr9qHSxPg3ONnJj6lSXU+e/1y8HnDZ3
oCOFUDyd2Z1ijNNW9UsC62AdDHxa49ViQkUj0ZCoAGc7A96PF6vlk5hfvVXmuIKNh5Nxfm1jDg2B
IEgRLWtRevLJOqx3/o/DBh5ry7Fym+ytbOUoP1KgouJPA9tRrhd60UXnScIQosJ5tj4syqis7fD5
l4SaC8apAvlfQS2UxnQXkLz07Ts7/sqVzSjzBsNG9qppfPE7WytWjb+8kj4hkjFuBIn0WQBu/ZcD
A/KsvWdMXMJCFI2QMlwuSNYuUlHzDToaqRUDhuSqueJeDWK8uOPnZSIon3K2NHsczQ8uVZTJ57kP
48XiVlpkWqCc8wo/qDwsxHdtYeHMbC2P7X835d5c/dPDj5x05dDL6yYuYrfHPkhoG9h8/HvIcyOi
GjMGVNuH3whXQRT930ZYyosuZ0Y0zvDKbgI6XpUjoYKZ3pWTc/WZljqps0gy8DL90NGW9hLl/8ww
4jEdyI6sZ2YUfwqNpBiQGtEsvoaO1tUTfrS6H3e8qCLW9n27uTuCezvCZX/PNlNc1pS9nsegMCso
LVrl4eqUxb0mjQVNIA4BFfGaTbA62UNwkpem2bwu+37GQ60/UXC24erTxJVbhtgjcNYfFWY1XsVz
y17E5YsclfzMhnhzkVOuV516zM5bHoom3Q86hWgVPFSnSSiARkO8HUe/xV1K9w7Kobp/QsPaQDU8
VLtAuuJfLEybhsOWqwmSFqbZvi+tgEKMpMTZ9h8dvOsn7nkjwK5osvbVa5DKW4zwmDTQ4SBHRokj
hnYveDKRoMU69BG7Oc1iiXXjzF1VCoRNhF6IKySExLFghXHOj0i3juSR7NKrKNLt1uQOwtUjeTAn
rHcSD9+DWx69us5K7gUx/krqnYNgl0A5YNdjjwRSlg1oZBH8rFKCqw7OpAi38Xirh1s86J2HU0cz
fNRtmm0bTMqZg0gng6ozZpdJ9Mknpbo7op+XYA/QYxyLQczBWlIc1g2R26YBsbX6pDq25xULJsGo
03+eX8fNymUO4Y7tZlHF95Qs72639e6ZVNwnjzg7o+0p8dVt1ePb08uDOYcUOMCf8lbFXnudsbng
gnOspKfsVB5yfywjSuriPsguqaBqQFXZsLynA0+ngPlOm3VpdrwuQDrBbaUNNpHdxTYKeJ2GwbSM
ftsn2UzhlKWLeivyAyAnFhPlJrlTL9FRAt0Tg0IFsGa+tbg/ZdYC7l8Yuk88KSobo7oysEFFld8T
mxg1RTh5fmZDMXJdxt40bUvmD4lwAPlJNIIlzqkGYsck3+9756jkr/N4ClzFyXyHbUWpIo4OhrAw
kdnpLqT0bm9Tj4Ii3S3W1vAoB++SE10kcQO9Sz9B7cR+MadiRVCKA1d0wnJjcNnJtMlx7RucbEfK
ObS8bvh9uvhtnnuCyfmnVxwBYiynXh+Zes+Kguph3lgbvELqOYL+B6gcrnuljyw9aGcaRGGdNxUw
IGvaevPLmAXC1PkHJ7OP2dyYdjt78ThUyPBhxr3nPvtqxv/Zrfujcac6gMtoQuXVC2VuQGBDKMYb
AXJ2H6ylLrGxyLM9ZltU5Jj4zuooH4KkUDv10lMCc/7D0AUOiWsPX9MpPsWAqjeqNgnJakMk+62z
wf6SpfQb9IEDKHKzrY+I+jst4UxXo4J58IGBLmMe0k+WswBgUaPCrNa71vpEAZzZFPnUaUKffMuo
KCOuzoZwSCue/F/S4Vr+ItILmDj31Bi1kXF7XsNZ+93ZwYYpg3tLbhhnpgJa+27ZxPRpWO2usbSF
bQbuKHOQkoBO6iaMoaPYbbqmiuZStpKDeFUVgWsQgCa/UaSIeExwhn2nN1LnmqlKlio9k6fF+qPi
XYfqJNSnvQL/TRdk7g49m7FwLRl04VbxBnsk3zUSLrw2WMB2Ht6pxrpIUc0jrEJHCDMYW0Dy2Bye
RT8MWrj1K1aGq2CU0M5rwKvnRo+fy1cHxIPFj6dzNZ5FDLpJnDT0RFsV+kE0YMGPofJRbZMZfXlt
Q2Zr6bJTibuj/V4M3mwTPUHXhE51r/AyLoRvVLoe0QRBWF1hkG8Iqz6IVMBM+1Ze8O1yDaTOv4Kg
Fl2r8uqVKxUJbQqisrT+uKgbyP1RwsiLucpWkvCjqSU2zhV59ixYmWNoRhPi+KG83xEOm9Qwjkj3
s+DNgl863181SbC6CKtctKlvgYTvxa+yyvkmhUjkYsR7TETT6iHPPDdoCwOQIQBe4+8VhQ3UcrOT
NKNCbL32o3RURaLgjNYyYdcD+Fgr05LWFkEjMHA1tkpD9CSsJoTyFyTI3uScJ1WoQS2nQZIwIU/C
Vo/HsOZwL/XhferXlj5rXDdUrrar5TJI4XVUa1Wj4W3OGot/AHGRpXrxZVYKxP0oXJStPmsC/vNa
UcLvL25aAQIPD/N0UZUu67ltgepKNy2wEqLSJxysGcCEaThhvDWkA9JO/ufeln8s8ks08xJjVfFk
qZSRX+1HDyh0f3kjs0Pzcaese120d98swEOoQjJmUIBzrq/zsr7YcWsrkoRRLWlLGDZAWdUmDonC
CFkaBPJEAklLQap/5L7DBw5Pom/UZFAJRFdFMGVs1KKh5jlwd/41kFt3t/mFQ5Irlk3yZdVrDKt5
BeExXrRSpoqhkI2UaxS4rJ/0ThBkOgWY+WtH1uTnliWNNQBQKLMDQ6MUu9tYY6SecQWFSGYBbHB9
g5VNlXOI/9svVeWMdSCPAVBYOwUYOX+3D1um90Ko3wHCnR/2j9D7fbdHc6AlW8bL2x+lXGfksard
LAKnR+l5Sm5B7NejnbRmomABnLpfQI8pV6lfUcmKoPnOBEhy7wDlymCDxQm02Icq3fxu93qdTffr
3MwZ+QIL+Nb9JXRk014e0BPHCe/P0KSnLSLV5D4RK8hjuOMQVxvQgzE8eVRznoaD79KVM5OJ3hmM
12bASI8EKuroTN5TvRgRh56kpQ/mbmXF2AQoQnI26+Fw1KR0pqo6O4G+fZ1EBp8x97Fgv7qIhqT1
dmxxfHALGju5w97TnSvb58/xNtBqBwQPSkB5s7QCOIE/zp+5AjqlWQ9bWgAD3b3nNJe08IbxAUTD
B5zESqI/LUlUZhbaA1DBCawYVizbCd4LLNWqWvAxToS5k017Ql77vi4MBuZgl7NcqmB6lcbodSbp
a06Q0gS3rcS4oLAwT+78znnsOkDU0kX9aW6MOteAinzNuUB5QA8q8RGH3Y59WEr4j51BeEF8vHyK
fJ1/Ggz0NQKRHL781pSIhPLgi9w/gs+gasNQVbGD6X06yHrD6HEQrZfutwwwM+DPaNox8jvjfxFT
WHL7mbmmSzMDMkMMpnaf4ZIuTNYgxo9GrzYkm2h0Zdf91yUK1qCL7IAQXanOWETG2bizLhrBq+ml
4OhqS4MpFz7W1UPT11wj+fK2Fh1zR0k4ciH3mfumN0ErbnR4kOfjKrTDCqXveveZIFcB73fxjhh9
BJHoJHOIyUzlajgIvKIJG5D2XQPjr8L70UcTapCm7+P1y+WjrKwOJ/5VMuVnYWnXRIFKUeGnX/hz
cL9/E4Eak8dx9FA7HAR4YvjgrSPDMlezyuhfsC9Aih0nT937m6IKwtIWrWaA25w8+TZHSV5uDqvV
g23bI6wTUnCncecJSz2gkiWhqXBM050Hq8duKNJck7vMazL0bvAFsPezr6Ho7lwwyd3SZDmxVzu3
Cb7ISzgBnh+CsCn24JOJtTt5pNHZxbpSPSuFNu2vId00UgyET0aZAZMz7RQ29HaGGZHhM1I0HdvO
BCm9jnQXN+9JNMqUHp3aXS5e1HpWHFeUsqr5UFEKzdSQ55acxVdIBDY62Xw+piq4C5Sr1fIxb4Vl
KOfo5WO7gl+69mwOzeBenXk+GfhbC0x4ekjntkaHWK2X33o561AXZlkJPS9P3+jiQZ+U33itu8d9
uPj0sv8Gi3hRZC+BHe6zzecDilUuEhN+30JXWvCUq0OxksV8QucaS7A1GiTqp4YZwvVIPQQj0SG3
S4iUozvzIedILZazKi/VOIVfk9S/84L1Yuh94Okyo+7mVsOb/GEcpXR9Nq4ZAjn4NeUCtuvzwTdw
+KzWSdBdpz8Cioz/w8CZbf3YXzQ63FBq5fsy5eeXCmtdaD6NcgQyZeWmJQnQb4KNVTQYzdO5au5r
icqgIZ7nXmGmtCvxHDyLeBeuqL1iknuAeC6x+FfuFoX4WhfjoG7MW/dHISAIVrSWpEzQsJIw37qx
uXmGB+1mJSqEjbfWg2R3cDqkkEx+WGyc3KgvpLu8DusriQi7qWJ5rmf4F2007IrY+af+oRFYwWG/
UXOmOXcRyZDfpQE7HuwyqKnQkzoeu6cWOy6rc4gM2KEE501ppVL0gNDL15xuZeivmH0unXpKw868
TIUpsmVicDR4Gq3kL6TUYWKNp3OVyYeXcm0AzkJxKFSIcxRS8w2bfpQ22ZVOhIIp9S+OrVSVBySy
gQJwEgNQNYxY2HoM/KD5/jjDscfAL1y5m19sZNAl1he7oGlSxIR9kiOEJszEFiIL4GptK3hZwBpS
iWPqS5VgXS6uoYvhqcsJd9aH6hXdG0oj1/bZIubpOjgShA4Q/Ok+wjl0mm+AP0xtdb26FRTGl3ej
Q4U1e06nRcdfngqjgxGW2+HUan20t19Fig6rdIirfT1tyCk/8vPcFu9KGoqbN1KEXOWV10q1OfKd
i9PctNWKS/dQo2MriPIbiSyL4zRxk5lOGwGmtDwVl1laFBqrF8REz8UAXaGlZNG9cSu3N9eXvhui
SspKmyE2+J3yTTPmqkP+euqGzK6fdG4iLkZmF3Mo3ijkYy8PzEs3NjDcNTD/lHco7UZxoOw9K6oG
H3EB7UtcwjLgcW8x5kdwuLKLewdgxaQauBd/CODMpwcqhTrrYgqHN9/oHVsDkr4zeqWurnKlWVMr
1o6WKnvRd1pZKonkUXyFPyO6/iERvISjBDbzmygm8TP/mkQoXNgYnyV0RWhisXms9L4k+6lE0wzb
sZ3v0z1eJUPaWBOdsMqCpjnyTqcEmP7UqQv7rD29KPX8U3aLw37PDlq5KzPw49hOT+3OSNHhWnsH
xyVJZYc4Cq1PiUfztwvLOOG8ymbuhbz7Kny72NMHVVJuNoVnmdaWtHptI1ngPL5396fdae0Cxp5u
8HqjeC9+U5cU4d6SOnXJnv8mjO6dgoMa1kqsVk/yHyB6PXn+DescQ7FEGQaGovrIwR5SABSh2Ai/
ExmD5K9JDLtD2l7+FSrQhhqqaWpODGBg3SZiah4D+qi6+gAUvUYxfsubM5Ts/u3VQfyj3q1c+eCx
WplMk7lML2V2xx9YAZNLQnyMm/xQdei+vEzrOJnx/PWj74m5q0BGTUMFK943Pat2VeJKi/qTI/pW
bh6XJmmCgU6izAAVZ244Z+4zHfQPORxXrNXdu3GXT+oeVNeyTPXKbzl7RM1Zl18RufCJ5QvyfikC
NN6wyi7oIDIY3AKYS1tEVSPj2emFp8y/dg2xToTZPI1XpTrWPhXBjxLJJTpd1NbSGTirpfL5B2KU
6JIFW8yGNM+RyEJcpkys69iSoTd1e4t/nvANUvu4yAQP7j13ewIyoGkI0baRX0JgBKw40s5G32NI
Jw0RwnvHYueCUfMaN5jfwVq01wWT6ANiiQaXMkBD1vEp7gNik9I1VtghRpVD6g0ReMnpZCp1ahRG
nR5uj5ShaCnKGcnJgRRSguMwKWIHYze5EbTms/7PqpsOs/DYeQkNNqbf1NXZbZUrEDpqA6Akvq94
x+0iBgeicrIO+kb5cJRviqFKf+AxpNYdthEJY5VmPvOxdnoGdiGt/rNd7W+MdErnq0YowbWTVYvd
Zjl5/7hp6lf1GZ4vCY/1+zdFB6eJCyX6Fy7T/U7i7Uqh/vbmlrMJ4x50WKepzS0UGznXWuSTpC2k
aM+cU3LQp+TSL9cRFkpxhW/97P+Dpuh0y67C7ezBm7xHneLPM9dV6WMLwFlpsq2tbAaHVvDoMn6L
4GZhiamjHy5SXr1Dlme0O1SfnGWH8NlDluUq7gOi2/RYhS91FY+AOIcYrSO09X/Dm9ni0BGAYJS2
KX1Dz0CnMzj0SRr6YbgcvurwKh8MXM4HpguoHhS4wG/ekmeG09zCO/NwY+6YeV4Ks72dKh9Wdlh/
BbxHwNodeNEKl+R1AOnn0Em6uPxF+DntBdzauQOtOKG2z2oFPHdWMGy962TWnFTDOCdtqB/kQU2u
IEXKbPV7RL3VupWeWbwpTVyr7uwGR9AEwbYYvEOWiN/ZrWQcECg4TRH40Yykj9VMm83MEmX/701y
6dw/hlq7bAw8Xh4YXG+OT+65j8r7mhEoBO1FPQ6cUW3VWjqytxF0zFkLsoTzrm6FUp0py/hfLez1
GuO0OiK68+izfrtGj7e3RIpgno5Nzug3JG3eM9qEtwA9jVHbQREG7JlfYIjAKi2ty4X389lksSns
9RhqRopPZnayFOiKtowfsud6elDqoFk7KPw1k4NXucmeSR+Ne/8mUoY082uoJBbZwRVLrdDLri9v
iDku/hTkmyAm7iULm1wwyJeuqMk65xiYHtQKdsIyatGcmT9FmVYryO98Cw4qoZlm+4Thc7f0Uwh2
FKxi6GmzQcEveOzAnRxV5S1aghmkmBSburhgTzTuQE5rQwl0D2fS54sNs48L1rzn5a/a7cWu388d
EvPXWSLO9ZXDzl/5RjJHTmIQQ+ojoKIe6Z55edPe1GsKCap3X/SZ/pVBSOX2tyVHxqhkzO1f65Lh
1rNxaApwuboDOyTZe+JTPMX45x6l0yGqslxOEB92I6Jd9NlT7lvbqfip6T4c2RcdCzN6uoRRvCRV
bf8h+s39p8nsTnjVBH/U4e+ot1R+kmqQFqk09+vx+4p1onLb1rqAbUL2bnwz8Y1ZrOjDkQBGJ6JB
huxViEjGIjdA7EVAMD5MVdXCaULm9ociJCKU6Iu0tLtgRAKjt11Wl2/2MQ6AQeTGebHy/L5sGswO
tSaIiqIaM5SX9IMArwNHn7mCI7/v2iUs3L4mQXVVZtnTDcub9cRFLAoMkqnW4RWL9wd3DyBInEnd
G4CSTG9qe720BmmowMrxfnhjQjlxrdlJb77bUsmz79sOE95o2rlBQXEgAf6KKAM59VRkH9QBDNIr
qqLiwGPlyPEMuEHWA+X3QgmUxL6Bl4MZ8X5R3FGlbHX6VzNLqFikQ1Hv4psQ4OjGsiw+sanIUXDE
LI2hvcXOR9QXumFYO5p7L+84bSz/iFQ/m+R6NI7IiZOEGNETxoEuA5mtOeqwZxlu7ZE0wa5Byewg
VCeQUV/VQNIu87qw1HfSsSkAiln6FYKFPdXoVprn3OIRxUo9s2fUni5wIJOrdmWiarzEBM7xYLq4
p3ExWGP1cud/tgTDYj6CPPW1IBNRJZT02PvPnGikOkr/5Kvo5J7L31htZeI3y5nWlMs49Opgqeot
ba316U9anp+Mgi5qNUu+hbxJYFf+SsCwoSAz86JodXTWDJ013KiBSUKR6dGHcVXXMhxJbvgcxoYK
RoJCxgt0eFB0NQYuakOaf8S+GNBiMGMQ6swQ9Xo/GjDlTvH+F6aYk86GfCuhlm5BVjAfuRJg9/GX
hBvxeyeOay2jEYsrhGHYDwZVtrhVN5hfiEC/BL1y/6N1AIG9GsajskFNEWiTtYqy+5A2jfReyIYx
w5gsAGiM0/8IfIYK2xfGurAlEy+SRgvJZ2fVaVZvNcVpBMFJjS5RfpmkOJvpGFEvW91u7scy6kEr
XQ68tBAZm+oEK6d0TBFPLpXCCRWT/MKNf2M8bh5bH54I9n0dOZdq5RJUJiqNnUz1S/igY4MkcOkf
cDjS6JhwCJJr6GC8BX5rdJKVG9lLXmnng+yahpR/6C7rlOOMKaaIo5X+H/AM+8blFzAfFGBrp3Q3
eTN3OnR7vh7wfQb6kRwELKRH86WH45cALhgtMcfIk80/wfOBon/KnYbQo52I90LY1GVblPc2ZsRf
d0PXdYdGDuYt8tBw7V+qBrUsENQLcGPpTfiHg+svKKYQW85aWKrIv5kZ41DS7z0jnGoLIFDB5qDr
fPSotmglnTDyKNWIrUXr4vHwL2cteGlbeoHSGk+wHw5f+ARNE8DkL/+phveYhY0+bESXyUoqJ8WQ
G5vvveCVgbp3ec6j8es8JVyjoLcezop/sVfVjXB/hqXBkuatWY13dIFR/5er1RG5uKpTFWC6bImg
CagFc8tlw7olVUwNX0RbHF6DGpuybkTRqCIIGzkrJ1yoKDVTxwQYVkI3RKpK26vbMbYZfiRrRZcr
fKWco0PyiWc6LyL4NtEVH2xdp/JYopHzRKXskJK4ZSjnrfBrBHWGFWWTcDKbxSPzOsEVm8XabGrv
67eSkpzt+QkJupiDV9KVE7kffL7ZrDaQPAL2zn4kn3cRLr+PBshsK1t60nfdFV5ztbJQNNHpJ/zV
bxeMqV5TKvZGh+NZkJCNDhJp+tqaVwy0TsdIrL3UaC4yVkzxLsKBdDunsUnkEzK8F6bH+wdWW9iM
PR9aRdiTiE200Y7yrkwX68oq52sc52oxKCsj0HOrzAdJ909R2rFUbv5MpVTMwbllvy5O+dE4lnhE
c2LLtBXnxTonxXvEakAO38s0GjnZq/6k0dKU92Jq+VhKS9Dh58O9I5mVSCbI2i/0cUw3FInvA25u
F0XNaRTJ0v4Mb/tGErRdFHtJbN3HahLNz5wSYc4FU8lHUTJn5f8RTl4S3oU0bJRYInKngBGRJn2A
qymjH+J24f+p4d3LPiwLqQwbFFcxVwQ2hD2Bjf1Ww69fmAv8ZW/sYvGSCoNAKD+g4f8oDyrUD7H/
PE/W7WEMi3D3Y7rQPIrzLrR3E8K3UM9wmlaZ1ud/UwlTM1W0jPCbE35zumSR9mtsJI65J71NpeKE
eB+pI/biWCjmSpL+l85xpGyiddlCLnvYzCNPutUvgMjqeru4PFPW0obxcrA4JLfvz/t7YBS2q/cN
nUt+dchrB1uIcng2fC+ItZyHMCP8R4lZZ/UH/S+iq1Lcn/bdzzo0xuHnwG/01l9pxNUdrVbm+VAl
2FS8pWnM1LM1Sb84xMUBf6ficspT7Kxw2wDLMiSzgytJjJgRVTmSxdkzTopMpatrswoXY3ig5zF1
3Xr21zYkZc/uetJiM5UuUsaqvd+VtrvHHAUBzhl2dumVYM4JXYHoJ7u9R7nmGGsQRMWgqQtWWC92
1Ims0cMlqUv5WhjXgAh/bsRKCPIJzLNGu4KNOPCBf+ypeySetEfiwj0Nb11xnTCjnYzNAq2JqzhK
xY+0PFMGIy7vXGxuR1TYtSqpltj74dWlXLtu9DI3HRtcYBg0sJ1xtJ1x9n7fvSy+4vetZ7rJFV2r
4ryz3QtEiMNN/MIS9S41JLDfxexigtFMoRqS49cftq2MESvHzo+YVW6pELRdLZI8F2yNIMfFF9YR
I2TtmPleTdT86BduHjGp7mm8qRNAaRf2ytbs9XTOeTHZWV6RToSAktWu8qEopa3i1V4Rp6bwm5Qw
E4Wg/NWtuGeD1ptaV8eZMnqLJRpAqUel3XP+l9ngswLp2p2yBrcNlrxVpbsZH0rB+vMTYEO4cKoP
pG57cTDHq6l70fpuloS6On3HXgRT7hY/mPhGPo5Q+SpGuBzZFqyu9FEfwNbpcs1w44o6I5FZp6Rf
pt1N0+CDkqUGQ50nah4H7ARXq0xwKqD3fExIJHI1jKfoq9hplmhS7qtFLmc711YHJ/mZGqKLbH+1
yPPl8pe7clMtOmKVKL/sbyFJPlev7G7pODf4UEzJEZ4ipVCyCF8xachZzgI2MuZw1eON7iUX+UiG
MBjyO8f1ZsrzA6beV/mgx7bFeQyWden7On5dQ84mmBX8s77T2k8nNggzCF944X9IkrFpKklxTeSp
M6peDFTyoq4aI3OheHhzAdEU3NkdLZ3QiHqr3amCM5RwUzmZXZjal4ozrgBTDTvx46iRwQDPf4qW
T6IDLX+O4V98VAXEmUjpD8kFEY6skXTjjoxFMHT2Oe85cJ/hQtKQfSb908HVWSAooIC4jPWrIz4q
QiawFnsfJHh92kRpjE18DCcC2Fs9R/cdUIFSYwVAn8MhLCT3jWsIsyY9mXnC0oARE68wqr/l7Zpl
6z9M6WMGXm8Pq6UpBULGWUrkU9ecjdsl1zpbAFjCSNELDOYe6IEyKadd7CK8uWrc40J45dMvR+Tc
LDw59jjSoS5O5qfejSluI6hWGx9xXb+kssF7D3MTZSmecBDwoecOfqGFwbNhLEo/H25fxkrmr/Iy
S+tyvhaGmO+uEiJixxIyCBqf2OgC9GO+pSh8MPbI+lr+aBvGVAodn7tqCRY1Rcqt16g1hLglsVaf
Fcu6TP50amx8H86R637M8aoIvl93JyDUa3Qo1hmKJ4YRd3dLLE2vpXR9ZaGt65De2bj5rJqTj/gB
SXQR0SUvBMUqWe/SGweH//uOagXNun+Xugm998ar9nKH4Xsh+hS3TiMfKKyWsCXtWah+2O8w6fxm
weUkX3w0ClU+u3+ZXaIZJYMh3Hr5qNth/4WEpyLV5010UpkaaBDjmIC+Oe4+il3KY8L0papkpAiq
MREuKV7a6zxe2FZNNmJakugE7ou0o1kQG+T3EmKpIQg7zRDrUvneSTW+BLYCNl3JoDTctukn8o3C
BlI/RVHEDfC+PS/ZSPdFkMZwYtI1lIIwZgEmQ5IqIIyqWHupKaPWKpXyWJbhpo9F5c46RmwlQtjb
Zo2fM11zs/r8POuQzL4K6IoYGPV2gd/4c8B87DphQ1NUoVxm6EpBbmH34jKjO2v0nBq3TBj+7QJ9
DRDksX1m/eX3VFwhLxHT4Y9sgMzazaxnGu+XhwoMkvzmpSIo4Nd1A9vNCiVCr4Ozhmuq+846Wbbx
VhkUe92aJt57wJosQKACS4NpWpaQanogMunhWoi7haGcc0DyNRb1JlLizKh9Ep0mIFNnOg6tXUgn
sfHb27XWak/NCspM6hgXXG8+Q4Y9XbkV8qqZ+nhI2+ysPewJzEwlHNFck73nB3oa1YqGvm2zb0DT
eQdvDRalap2ahzQpyy13ECtWPHnpSAfWL1IeVTuOuk2cmCoLRCCQvrm8EQJFzIZyz8hnyOAI2bDW
en5SgvSHu2V3yultoM4HMUtumtOo+5Snj9wBtsJuPmLdpY25aScQ3sTz3hzThWduooDI3oF9dF/4
LsljfKPk3xIp3eUeCkPRhjAtMn6R+e2kV0ORSGh5HZ8mNfjlodNBXyneInDQW0HvVlHR4nu9eNbd
zF+nc2o0eQCP/BRMzOOTKtKSQqds/NGiZqkPA/Ox3ntJdTbTQks6Y28IIHTmTsh64wTcU75jBBlR
jt0DZJM9zZD6GhPcPOJhNmVWPQCAtjagACSWp/f1Dyd9vCdWK7DgMJm6oKKYQWLo0Z9f0M1BBRdQ
BUvvX3uR/XBnhEg79Cz9qke8djzIVpjrPY3Kd425QZ5wmm8PacOyi6+iS1j6a/f0YjyrpfIx0LGj
wATStH2MEDLFkIIZa6Xaya1hmDisNwWEdrb13B4EW8YdEr3t9gW3Uo0Qvz2oQi/HDzx7Bsc3H0UW
S9O6zPKGMhrJZs5wmiAxcuWThh2aEx12/mndkTJacJ3r/Cc259BJJwdPkUYI9Sx/cJuAYCtcZEsQ
JOrIvDz20BJByxh2uCy//IZgcmyDpAFKbk+7hX0CJc3yuP9M2Ss18CAJ5t2JtZVJXVNVlAMahdO9
aeUEHPs8geaGMl39snX5SE9dfP47Rgd1ZMSvWJxbtBZGsqsVF5t20md7oxR7O7rIsdasDebqS5/T
T7FOPTpp9NYZ/XyLvUbT1ko7E4iHwjLuGcKg1ENPDDIRfUhwhMuI+tBNj5j01E0ILVxQ4D9GWz1D
+bybtlWx8W/hTmmH2+WqhFxhoO985T+p2Q45aKjM52QglGR8NXmFMovyYN+25geR69MMACvEDVao
Upu1vm4GdOeQM6rxj2E0rX4NQ0q8KzC+wBizcNC0Wx0osfuaV0mxxHzObJ/2m4aQvHnFnnoTbdaX
P6hWEfV4rfrV6hXVIKEpCJ5sJy7OsYlCkjWZiPcxwCEtX8d5COdgB5/qZg33Z6yT3IqcucKqsy3/
VMnE6EjH9alL2BuKzXoFx3r4GdEZSgoR/CNWSXrBZipNoxpnY3Ezy03AV8TcJuPHbWAZWhx1adKo
eLvyY2aGzHAWNM6F7RtbNP6V4/baII4Z/BENbhJJCjw/sg6dzGTc/xv+H56bl+uOlDrJbmWYiMtI
XgFfatrtPsrOeCDORLI91LUES7QCr+lbi6l7OjbqZV3kbM/XYkoz85JauoCpFdoDdR7ORElsqrQT
SfoxjvdBg9/7p0gp5W3XT9mi+Z9CS83L+rpRhRgUQFqUNu+T2/HEDrSw7rqGaHf81GNRQIEuoA9J
O9gYdHpfftQ4K1I3N91vPEywDTnp6GIk+6FIkI5dow/ptDousx03lLmobakZzLEh29q401CGm0TJ
o3jw6FBf29FLfG3w8jnWeUBvCQ36ucdFBzRJPt9pzLf9u9EU1l1BdjVTzHm24UZyPteKQLl7GR/4
NJXqbhKo5hQNTEEWfEhQZ/VHpDKVyzJI/KYhifQOGwr4iZ0GMG/MHh1Rf52QrsLh02Z42Oh4TEvH
0NOHPMvsRPtGNTBXvtyYzgoMy1fIxzeb/cffsPd7JS7BEFeQWZZv5ngtRbGlacubhxKTBkcorcqG
XTukznpUrJetpaWw7o0E60KJjSFptdQb5J1c6cMIgvj1vT5j3d0gSKGDPkjtSQHSCOvKGHJkYf0H
xYiwM3tyZFMPeYU1+vt8U+iEJmsTn20ABPo6905055UdcNfU2DWzPY9w/ay3OPpFb5mp6lWncMXW
ZWUqXfqss9MQ/Ar9k9BV2KbvcRd6ZPdQgehiDKhXU3UXNIS9OjsUI8Arbv9Vj6ugrT4L+yQN3AUd
CRBk/kSjOB/zGKTrUPemHmfEdRsSq2O9MoM4mqDE42Sfk07klVKILv2S+3wyfmpUx23g1ttRGZ0u
0/Q9NsxD+Lt6WasixC5wI+tGUaNSQoIgVGhsu0l9xONnHagNL9EZYeGnRJoW7TN8yXjg+kHojMbV
EL5lmv1BsE0Suupw4IL68WuZg1eY3+Nowj/px/YyvWsdvbh11jt5girQQyJSEYcmQ7SkD7Cx8qoN
vpmngpma0fGSSKfePbATqd4Mc5aIhBfbHEoeoTOruu4aQgZU+akedIvzKUdCzMQRP/MqnqUi89in
bbqtO6GWZQd6VWzLaSgcFmg2ncJ68fwTJ02L55rJL3687ue9ri7Updc2U3S44SJwjD9CRvugq3LY
Dr+BpeEcEgMN+cmPiE47H3ptIzaeG0OVdjr5x1PnSBO6sBLwvsEOA97yswr5HH3X3v8f2QaixXI4
MHi8SddGoXT3MsOKqN1EYWw4TYPNUXVn8r9thu7Z3O/HnZnrbUnZz1zPpHXgi+hiZAyD571KI3vi
KtbBCq0c6oEPvxMzjGWHWUdx8GYJ5UMsAzanKkdE7UKyvclpkS0BNaFnbkHtEffX3Bs61GRs1DeI
1u3owvvp50dkGA23QvFHQdMr+ZiwZCoGrYjL/lGdgKWhmuQHkx6skTQdZf1vglTZvPBL+KkZNsp4
sOHZZYR3PVgvgxrRdNW+fgzHPCnOlz2KjY7RYl1Kjho3Hp7/sKEpjEcdOTthCeIJD3zNTMKSwlBf
W45LvL0KiiwlAb1Mkk8czYm86cJqUsgU9wlJaMj0Bnn7Ls2wWLPEDsU8D+XNcMUFtFTVjrYHrCZC
8QXhNFhtJ3Pq2sXqQdlv2HWZZK/mygti+3BBxYFSVtobQ0KipVJJtBuAFu65NGlxO95TIoNeuK7L
AL4GTLtUXtPyEfdujmLg6favQCPTCo08IUXpJ/DB+wq/S9oqGjJOtgP0jtHQ/68SnARlvPPYTXcT
qwMFhcImvsktzdNMwY88QJ0yK8WT3vsSF470Ot5wpzOOoVfkxJwELHz5/DC3KQqpxVnMp2SzmoeJ
E4pyv4DQtHw37tOKz4iPsvjaZ9Vj6qOTl12IfEWicQy/+eSIaqIFUzSyq2mVlXu2JPs/wcTQMajc
bDohoeCZ7jZBBdWtGJqwZxUM3o90huEJMKFgDOdfcknhZSqdEIfNuqDfZ5+DsBNkMEA+JJv/OrFh
RJIblt96SdLCATEWp+w/FXqhZ6TUL7VzQLz9ODB5vXWJl8Hmsn/0vN8CCSgyYfjbRRdLCrqmr1er
M32+jquYMPIjuyQRznWUUGXRrnmtj+5usyBvCZnzlCd0ziZUlqrz+2HkPqB/GwnT3IRJHkTB2E0P
1SkdvDQRs8cjxCjPMkvJJbIT5MsyDKgAzc+kCbG9Qan97mD3InxK2cZi4GH2b1dqEGKXc0O/i+Ej
Ma/XwR6G1lqBB1kUSC/SmKad3UpTOzdBuwIgY1++3FmUhIaCzFF/eEQNeoaH+u1ngqFFGmzL4tLn
mWLqX2pit9zV8ayiId3A2AEK1rAO+//Hlbv7flKY5M1sRoo6BfY7AgZDAeVqeCMT4tYu5s2CFZWI
utvCDnxICgZGZjSwxmBWX9Ac4bNNzwbWp1qJfPuYyT9xmw/f1nielV4KI/X3BYLGW+XePAzmKr0o
4mXrygxQpNmqy14AHcZEnM2W2k4EfWYIUINy0hcMXzyueR/ZpjLdH4QyqBH9ZKOEjgolExhtbYSY
AZXZmG9U+0hL2wC0GYby9GiSiu8JMcfk5c0UzBJzaMqCFCtnJk9C0tFm30Y44RqM50uH4Yrrxmmc
f4pix5QTKl3DIr5t9XycG7/39J3+JEE3gwy/45dX+l99VlD9/ZOepbggIdZknRcFZne5XUVU3tXU
wlMgFFYo69IQsv6VIYG8mmf4CooWhywn7Xqzu+JbY3L/0gL+kyCOOiL4sBKxdpKA2WtrOeqxadcI
lpNdozvcpzI2Ry+NkFGaqtz3Kj1qLG+TVOsVEN8HVkFLnu3b85SH72s3gBeUMCf6SfS5t81Qb+eC
TbZksqg03RpQgquJYkrWGXJF8j+jWZsAB8VqgUA1kKLQnY/2QapK89Dq9BFzx8Q3uzSS7IPIM2UP
TheqkBQn/RrFR/1ZXcq9t2xAA6cWFY+EMgCyqKUyXFNHa+V72gv51ZB85KHd+XHXmgcLkmWvWSyg
/wjfxetJv6sf61zmNom9BkMojxotXEMOKFj+4LXEqPPF7N5anYaWfyOMNbSebSuPJA7XuXCRPlGl
nWDQtIblnqGIp2CTAvXgibALZ9jqFkuJC6z5LRUaMjldgEfX0cbEUQOeekDvbRCEl5YJFw2YJe0p
ThlOpyEPzdhhIOc8C2ewENQH+Cgh1Tq6+OONTMFczi5OOv2MzSEBe6PCc5Z/s86mac+0IfzKtMBP
KbDVU1EVOlXciuRMIGIjdxs1LPXd3T1qAZp+LkqYsdMp2ZguQ8W658QolEFVUyZoEk8bJsh5XFWc
msSo0chUBKTN5j+Jv2L7IdAvN8TPv0oGVcV9h2v4lozV4I/8JyD7qunO8pfmQFqHR9O5wsEaOG2M
sUpMDSIJH8ItzKnDo7ae6Vb1uZvlXFJzD3+dvEx5zbKIn5YP3yW4SafpDfIf17oG86NpcwfrCT/h
YQ8PCE//DAHXLuKkxHbFEMWj9K7Iy3/RKjFxtJdh5iM3xqoKugFGUcvd/LTlOynwqWbknRsjFTsl
a5SSuUCByWsHqLUHOZdaSYRgcyQi78S25bohQFmACUwHRohYeqzY+QfmlB7aDj2U26jh76oJ+2qF
l355HGtf2SHzZXjNZlQ1RyOWggB4Mf9jklAQ7iu4FDNUhYmk7i2E0SlOqufM5+ucDMy6AyTU8nHT
buc0EHQedEnbT5YCka/jVAKxGMVG/e1AkOhLa9e0QB3A5VUPGDT3i6pktSb2hs+i+4Hzlu2fwP0Z
0lMJLoN8tzLbHMdjzLMEhrp5knyHVpCQE7KIwJL6qMya9YdNOpfeAPI4zCW3h29uz42+gu3tU1Ny
lkBlga9dTbGAhg6ldXft2FFwo3l/1fUb4h6lSypxHXljNk34JWhXQKoR7nyyZEyLJZiuAz21UNFk
2O0fDShQu5Xb4LFEOQ5zOTMWKTDIxQZAywTgl2DzCp+SEUzDXxLsS0DNteMCznblySUl+1HlX3xx
TdZHW4R+/t8NfZBgd1bDPU0O5dthWeXvc9u45J/m46U5yeLnhqkuPoqtgl0rgLMJ7V+843AtGjqE
dAc9vDy7HJ0zZ8uNXpEiyVQRXrU1qRGh89E4dzIruvFlE5DGPVBe1zFUfoGZirpqCkcZTRfGXBbl
TbRbu9iEEzXiuOkWYzs/DKxGEaUP76Qm2EmivPW7Td9aVUAN4KNqE5U8jrXnt9qF+t2pVIxK0gX4
nKmiIQj/yX5cby0idhiYezQJ1eizmeV/VW3zFpQU/L3G0hIxPF5ioAbwve8aEoFyaFujRVQ8VamR
Kf5MalfMNNPH4n2KpzNa9LTiZsb0wxGl3UqDfte8TRsz9rHZYABHte7/swi8JktxPfibjQJka36L
2G9JCNgRTNtfGhRS5NHUwvNfwSoNZGRo2weHtnBaEoaaXb9/Wh4ygMEAPOZzlkrpbXSI8HM6UMag
L+QK5Cd0SSjyAPsc3F3BZNpnpCjgyWfl4z9IYv6J4ckOuSvgPLF5q0mugXOjXdDYrasJoR2vLAgu
fsK/rUW22IFcZaUXaesC5sgbMEkncAolcKqVWJ/VLZfVXKYof2iDuk3fUO8fidxvizTzSiV463kq
7bi5li1cIh5xAsWZJrmdIO6eefaZjebQzJEiljytMc0INTTubQbbEDjmJJdQhp9Y/FeDDQ/S6vqU
JRIdCwVFdV4E3rergmGrZi46SQhXPO4hD5T8JNzzmUHo2BaLgcCNTaQZlI9tGJML7gSCxHdJizYD
sEmZS/HzQzyiEq2qb0biACYLawHb16DbepCvHApXkIDQ/vcgRZzUQ+6mFXQQHYpMaFuqJMPuStK2
STx2bZW6Kw2uwQMXhkzSG7jlb5TBUDXl9QiP5rz5JQ7STykU9+8S6xEvgLwT8x4/z8de2euEp6rH
pN/H5p28e4Uigg1DnETC4NcX0U8VlDXpOLN6fENYGTctIZK/Bx+iZ4/2rzc2MGBJn5Sz66sny3Ur
k3sWboJP8KRlugiDHRdUtgSr9DZo/ibwYq6FWJmAzGZT0XIGAWmZiqectlxNFqXL05FhaQTKhnR+
s27q3dSI77pDFS6FRAy0cWI6NAFt6QvPqAapLtzM0Jb26pqgLRe5EVrNVW95bFiaytbfnvzKvRa3
UkJK1Kv5w5uu8pzBaoghx0XQslvd19bJ2LAiVd7GFoMzVXvFSHerHZU1jBCoNyO8BZoTEBd4e6ZQ
n2Ac78uAL6H0zYzZ+quHhf/fVuwkWWhj2ZVzqfg43xKJ2QQxIG9Cq0clxz+YvYOrFmwaoxx6SzMY
SIMB3VfjcBjBj3LokL9QI9Czc5Nn6xfR8xB+/RU0yaqz/zmB4BQ5i+e4eW7SL1/WSlT4xs5IoeAv
QMujlZW7DpXwIvu2CHJ53eNDTaQ2KpjJf/fC/rRf2rtMC0upIFrN0Ro3YpqAs1J/YQAumXj4NtPE
g3TlT5yXdDAmPZZFkBjOoooDjrbtCEfI4A8FZy246tGWW8suDq91lrauAxX8Y/km8ERJ+hD7uqqi
9Z9T0f+Q7Nboy+vNND5pIoBUUoveWw6ahPcoCZYyvbyO3ik2IXNF4wwKpvogweIBUsOiwYxkmeI9
5LTjEHI+XVjy2fxplUlnqN5vqQ7P8KGGXUOBzU6A5Bzr7Dx/Qhg5UMyKmY8jYsW7SMCVd/2Van08
1V9bczraPH8u3IM3e8tc1URXNXSvaWJJ6a72lXkArJaWii35VLB3GSU2DsqycSUtFokMNPfMs+pP
e4PfgxhI3qtVQwpij0CtfCywoGdp9DBU0iupmnzdO2HiUvteBJ5oIPFsbJjhEHELvL8GE+QSVPLD
KJ587BaWdBFNlIUZQAT/jF/7EMy1GQ0UUKcKB6ZDmHEo11MbNXZOemt3ECgSQVc0szRNbQ+UjIpS
LNrHiHXLLZFJVf4B8nC2A9zvVvJdHP82UCrVWE9db9MYATH4HwmTk6365JaRfpARTmKDb+BZM01G
ZNYmKECpOybUTNRW++6gFaOrYrR+aK8mPaAHuG/D/9wxsSqngg89r7gWHXVSIsUvheAjN3ZiTaKl
KZuKBH4ie4Y+9xQtx55KhLmIJxkI6KwmeCI6f9//DdwDMKqJjyqH1UgBGq/LGZajBNVnWpFWR8JE
R0ncIxPwX7t7dcQEqzvqLtGGsPVAJ0OXdDRKVUSuNva4kuTHcJj/wO+KiVsn62LbEe7OXhnXRcth
C+zHfG3/x3zha/MonMHFhO0l1gkoEu2+cdLGUgerE/Nf1tn7uHsrbGg1zxjnWVNv/ZQDjP5mu9mJ
FgK+peUqoCELOdAsakzExeco9G6vj/LAC68Ep+D6ijImPex+M4/qEasTRZV0R02Gxyasa3HWnGZb
ys6kKS5JlafXaQOb26F5owxG7dqign5mbrP2vZaIzusoluEWkdpWCg4XZEkuId3ssgF28+MmzGkb
4Fti9i9L8O4o7jo0/Y143lC7Eke+NVFD8EesWPqBzyv9t9tJp1ay+WEomB2pdEvCM0lYzDVTgAaw
/UU8mHQ7cjl7HlSroQ9Bs542NTmBkYzOS2+a7YorJsSczJWSFOrWvsFeN614Q+rvOa7zMagCZtGi
EQ/Ux6+R0dB3KLAyOe+geFQHFFdfHYF64QH/xwYKWKPijlVI1EL35WXkn+A4nhdHexRTEdPCaHgW
tuZLxFMBCKpPsRPp4NgfrV29yycafx0KuK5B9XLlZYBuMlf+6PJjKmgHHM0jGKGM6Sn8dunTPEhu
rhMSGA6XATCEQdrSdzk2qlabEPh6WIN7Ush+MInavTBS9P9CH9UJW8R96LN0XIScEi6kt9S6l2iP
h7KSVffJvv2fuxJwZCDMSrxyvYTLGyqaO8oXWjNOVmlRrywv/i6kRFV+GTtqAFwdkMHs1Y1ms+d0
h6DlxLWNi+nIn0IeGvaopfmwBpR9a+mnn20sQ8737EMNmLjdZC8LDeoJl6Dx+QavNlA7Uh6Lt3Kv
H0QJ1y6jROgMP0DXgQiE8AeWALiIW1pxrbVI0csdqVmvXsMb7XYHaec582V5tLZkGMIViF9hWhqH
bkWzhXalsnFqFA5ZJ4DjWNslz0551CksvV3VsMRPFeC8/+hbf1vbS96zcYYFbQPlpACLgq2k76bX
rOvOxv9NUfJ/edr9/Lxpz++vkB28fLRHDRHNN/hmfUGmMKbNHbgwPF+SmYxV69dlhZow4rgMXPQ+
QASXlJbnzLKcpdibWZTBqQT2MQOVzxQyssmRCNHGeLZ2nab93gE4Q1W9yILXvXG/xHUakBCIjLU5
Uot4/aYXhPQ0CXIYkzyJMwoaRgEAMFVa2RLuY99RpDZs3gMdakOjWtxZ6comgXthlTs39BNhbiUS
LLkWjB7um6h1RsgusQg4S5leCAa6Ns5tUljIEc8FO7OvE4tUVlvpbqjd6U9C5/W46/gkHc9kJRJm
4S2QFal2BikhzeNg7+GweUWbQ221YQRWMlQoH0jLWswn+2VoWBnX1bjMyddXkmYcfXfDzQpEjp/B
9LQFQYFy1EWYWI7EMW2dSO5xUmhqikxzjvgdkU3xk+6bfo59LXuA/e6fYg+67xwXURi7tisegrQW
ik1HC/5JhT5fPY6NIQVed7r8Mu4GJmFCiQNjC+BSzYr/O0cFOg/MTYPKw1Wcea0E/W7u1pkeYzWh
LgGfibJ6kkYGkJXiJJflXNlSkl6ekPkczj+Uh1VCtjc0nxH2HsHFgVMWMICPBdBgkGS6xf8YszM6
B7fNYs6ZaWRqoBPP77pGZ/c+QMSgMLnyE3elouIomr4t9j4LcdxhcRfVy6raM4a0oTEXRlRtglYq
zTV2X6Yno8DWz/fe/Yt4CmIF6PsEcwaeEIHS/Qhu2U1VWVe628hXAYeAJ9xhppy33YNHobMhJIe/
wp7RT8A+6C8xbVSLvq07kXt+amALyfuPZWSBQKr7tCIT1OIJ0Xgo+a5Wzc0ImwyEiOIUcuTy+WlQ
bjWKtDvY3njnZ3yWp+T64feZO0QDP7dPpJpMZUF5y3LBzkKhVKBB4cfzAaiLI65bsncVYE+nygSi
FukQ7vI722hgGJ8AJCe+KaVmbjhxtf6PySZVewx6pde8sXa93weLaqTNzmfTBms3cDARxkG5sgTv
lgm08Xoo5+p2doNvHX7Azi5ZxY8FDg0Fxmb2L+jL2rcZQ56fYqpMzRlq0vVaA4D6q2MCzkBnLFl4
1tF4DQPMvplUL+rycxbXyGRaIOnUtKhvbCHOcu4nl/WdT0jLWseJ7aSpxLJTbooUgtKDgX+HzFpk
QEUXx0aOOGKe+qqreuTJJXc785+VOyalVUtHjB5L1qN1mCf5hZQuLBX/lxmqdt/9O1ntRJyMoNWD
+4W+WhhAiE1jn/lkeFePaPveDuOSuAMrtyUxod+GMUlXBxaOpDlP9Ckk+5Ys4S4bzQFtGSKUixhW
t08Zrd0fOACFb1bcWUcooT2OenKL+wkVDOkT1RzaVH9xC+X0JZsAyJWASlBikFMEZMfJwSuGHKvE
lLSwfDxLjreuZL94DIEBYDcW4V28fwg/+9JJWd/7xSOjh8M+iN+KkVEm2f49Di4DoNprGjUhee9P
jspmr8ZqF8MQif2AQp0ODvd8ovNKhn7KhPuq4K08QRMFpCP+kKjx9UlrDQRC7x9uX2t1zz0bewBt
KJBTSg1yRTXEAQXo9jQVM7UAe95CbGxp77j1wG0KVxUDb1t76sjCT3WaPMXC6CIsQDxvqPZQfPdH
K4GVJhFz9lGDK9RjrNqM84hm5Y3xmokgSgjaDxORhJ04kY2FHiWzboqjBfgTG/Szwco3MIJnGB0h
E7n+QqMvtT9kYUYWE644jTIY6tvjG0Vs0LkMfoGd1assksYk1Ng0hMO/fvcUZBxIAgzXkjOYtQCs
s1Z1axXvUE6Vr38IblPn+At6UjKQEwWoBwN0+uQ19iOnmkf6BRW4A8RDmA6RvvSN+IgEgKCOfwBs
vw8Oyet8IPRTeIwuq2/3Ppz1ZY3OhQBK5aX14rFiigZwFSvM1wpMx6fZtC+nefgICC/L9CPC3sp8
LtMh5Vy3A/fRglEHJNdbw342zfnWECziwgMwZN5LbRltzJ7XB0lnep1fSO/q1eVq2DK+C0T4YD8Z
Ybjkq747PT4MITpLY99Eo9/np90T9dC40RBYLGfyCkWsDWmGT1UkyEtrCE2VMHu3qmf5vEGffsF1
6Sjoi3/rPOdAit4KjCWK4SnGBeoLI8Up0iaVDYkvKnqVYhJJXa0ynPeQSKbJzoZ+v+uQlSmZRpkF
ySvNTU1lzsRs4Qfgv9yDT50GqNaZadz6kSGXZfO4p1SsVRPDwntHwSlrnuMeDQbHb/7FE6mwrFx+
xSdW+G/x8RUj+tN0gAl3x07bQNEEEIZ3QnWSLr7pH+HPeEGpa0h36GcHl5n6wl7gS2NVdiqWdnCg
6gDI7iHKUgQQAj3HQ472H8W/YBl9ptltOXod4GGqQLzshQl72sOvqhS23HM7JqFgoeDfSFu5iXTR
dADVI/kUxxNWmiOAwsTJrDT6xIe3SzvbWUo4kmCzaZX7r2UJSJWlIg8L5JeTCxVZWY0EBtlRTUc5
uyctBhB7D7rxRX69ZfEMITAw3/W8Pbv9jeZ6NummaxQa8nEOWSXolT6K5DrRhCSklCfjX3y4tUww
MsaLFd6tr01C8nR0P8vTWz4qnT6AMDJiVyZ/cO7eI18s80pxU+TCMWIcTg0HQgbNUtSG17RkjFA4
Za3ilylnPmn/cDFTMGh0AGUqQ+rI9scI6vj5fHLG2tWnnGrNuSDY0Mk8RrmebmpQQ7SPCpIqvsEX
tTuCUTQwiPwO9yLPJz9Fte+pOOC9LIsIRuWLQnZpnTzoW7UAZelH2Gz4jUxP82V0/8kyoBieOF3M
cJnmfbOmKZX7W+mLzPDHomU0CjHWLzd/49YasN6WyL9aOHpL0kFPCn0YpNLt3yvOSsVaXuv3i4pg
162Ww7/8TVRdCiYqXTQX/TsAUTRerev1L3P/PQCcFMRz3YLHT3iBvE2nc8oCSm06D7QBGB+aIP/3
uSdp4XSTemYZt1/9y99mKmeb+fdW1aeVZZvzCaOnrN4/fYTjiMekv44I+Mznz7I3MaMOPUi3zAP+
zUBzX/puQwlzt6ZJ6nY5SHQF9/60MnAke2YmAaTQAX6UJWsh00IwoZtvBt9pfH5U0ZDUPvEI9qiF
6dIR5XAWaMEtwdatU3Cl2ZlPPpWmVcIKYMCKwOOdw0PkDPwjHiR7euGRvqOXcVYEU4c+ChD9vrDt
3ceezo6LD5m5CC8vSc7/c3Gsg9T5yVH0bSOw0VrLJjpRB3156nAMeYo7xHIYFXpAK5Pbh2xcZ7O1
KvJ0yyv8KIRkvLAfIf6VfOVSTDNOCyKREkdgfBkQb8s68/UTOvyyRj34RK0MDdMClljLzuzEQFQJ
npXJev8xkbNicsSO3UysCKAqm3m7MYMuiE2kB5Jjdt0ZK+upbb44bdEhIArFTFA4SKMznMU3tU9d
9t/Yk0MEI4JhRYLjnLdQCHiFHCJ5+koCYqRSbRrJFgWsoGRCNMhZjhpgt8E6/VoHWY3v+FB1T0ke
x0L1S2DKb81MxQA3di0Ubc2xuTB8ZSZN/gBVXZQ6Lje+2l9T6coSNR+Au4s9IVpGlUOcQEYW0YcX
MKnz+oseuRKF68dIYnIS4X6MeLBha+bOvHJBNwx9PU4sWWflbeTQ068h9a6MZjwS/ZeCfQGGimEv
SzQxoT7Svm3FkqDlB4aEDKx+Fi16AMXAE6/PueYUvRGuZGG9z5ePThy2YTdIitL9NHVOXeTH6umL
pBJcZzfXR5b95QeVkxnpkxBDApz5lkngkQUr8/bbisoZqA8/DrKBBKGSbCTzpkx/8hjCpj4yOQRu
4So8d/l4KX4Frq8qvCFvsLEvdNwkbobktcfiqkuyWE0ojFaHX8zT9PnjN2U3UkcRrKMs2BIYnB7K
AflLhKN+YNkqGr6rOlgS58RQjwqjA56J56vIWPNKeTECkB7SVMOeGN08qy9SMRlzbwHvvIT20TDS
RmfFsn7ARX6QJH3gs5zLOzT30s/dt4QOuo6uC+90UqA5gOqjxCjNottJN+8qM0pkHhQJ5wzwU+IO
zbPehveH3IlDDNcKqFhQBKFPBmAfCP94ytcEAgzhO5MYdWtgHDlkdV7VOXo0toA0e0yaQBzFCzVs
8ztn1mQdzRmDeCIn0NYTh2JGqFYM+tmufxr6qeEXN5c8EbPfcL0+9IWb8VulttZpXk2Jugk1JO0c
egTJ+kNjb7TgClredQ5in1cwDbFS3A1xZ6pR8Lh22SWyuO8Ukben61cbsUFKy1F1CTPxHTISdX+6
bXqHe08TwK0T8tNWOhkN+Evdt7bVpfq6KrW70usmIPjUDVFwxFC2ZZBBgoL1x/I3GzVdMYKJztGI
Z9/vC0UqNuO8aHd7Hc+ok0tFlMQkbWvvyJuWfJhCyZoqUyBDdSUYB2L7TYpMKaYMLAv5zTRqmpx+
+IV7HcPH6BbEHEyGwcuu05DCnPMSEv+p/WMS+5MLBt3yGMwaXf6eTnT6tzDrlMfzD8sm/XKiS+LM
QHKnpE7OHp6wyY12A9v2iRHenrFU2dZtYh1bEDPhPvjVOJKGUmAWn7mD/BbY1ms2duIDKkTlMIgp
2838FP6+5mSJSQU+8gKBCkAoII8/PPuWBD0FbYsqY3UIfgF+H8Hzo4kpJpovZ2V+9vVN7xoZUjC8
9yPtF63l55P5qiysRdGS9Ch+Oj0G+80fhwaOYFTaH8NBTvF/gIDH7YEfpjzA9B02DwMwulblkXuN
WtnyxnZ8FsXcIX3oYXImflD06p7ReedgNM9zxmg1NFhS6HOylpKxCq55rDZylGurOmqY7n+QDXo8
dNuci5llVzBO6+qtutpSAPcEW4bgaLXNIRL/dF+TQ5pS2E7s4Ip6QPmKAgPTzs9Vy2izdMoADBcH
y34aJ/ds02SXsNH+9u+5dd934oWhJezszeOENXjc7SL7UxfCrvEvIiewksYtTPIBGZab/r83tl5z
RM01VN4sGzo645ul/yrPiID0epSQ7MQPWTHIAF15I1/5jvh9BHrUkLpQ5CrXL+Dbg1BFOAko/Abg
QgXJjbv54x/YE7hwUAkjFmuGk68wZwVg6cRlmFdrA8RE7V28QzoSu9Z9R+Wikr8zvcmwGfws0WDl
ogOPwTwWnClJnIinIpz5XnracRMlywLW2eixjEl932crgDsZAdccXSYHVSdVUZxvxDLdp0EtSo8I
YX8Vr90btsgN1tYy/fHhoyx6mlJOMXQsqTLVKrTfBd3hvliHorAH+qt9bB45UWc0AJrP/nrR+nC0
fR6FghgDNi3hrqlFLEhYXiyZCGY+BT5hYL0C/bwQLy+hpbCQvFWTKNW8hXCjJgJzanevFelWaMja
SIiTRbSi69V0pxT1nQMaHL/VdTkMSCITa0gFTJgCc+aW90UE7VJanoMwymvjmgsPeECIFQgJ6nHX
8A+NOC27doCT4ygnJlXUyPEqncngvRVPhxygRqClYJxRnv7Mn9qgt+jwBzSAKVNutrz6saX+fsgZ
pkCglcguwVr46RW7Wu4pRgTJM6CqV5gxKn9COfqJv8KUDDkm9DOwvtio+svRs1QjQV++QR1FP4FK
BMC2wSIhgZDE8WW6GDa3jxJuBWAmeEKQ6THb87jiIh1yuAb1+oIKB8DbJOlT8a49VrUJ29XsA102
l4DGwg8dLKeaCsa4DwaflcX2hm8w+l6XD46QC9iRfsxeLxSx3C1ki8DFmJZCNH7VFpb/nJogfSu5
R10sesoVJxE3QzCusGb+0JDLiGBgVr/T8pPd+WU8KEjPss2y+JNxP1e09+Uc7iRsI4LXXtbvff6N
XBGTvV/oPAkEyEou40bgYynoyCJ1whkFHfDVxGc7MeSli3n8UBb0iBC01cYM5hSWopsGAi3v+tbM
pGPARkYOLZWD+BMu6T8Of8BrWwCYq2v6y1eE6oAL1jxdTGmwHFYaepEfa93pJ0VqpDpKzFcQS9FG
hbZQGcARHDaS2jc8sNqb7ePTp941wX9YS4weV8QYu+Xo6rSBzep/XGfFuGGyl1YjARSz/W4dhtsM
lfuHimwpgrmZY5GAQBQolGuNgPuA+GIkz7xCVh8VbqBBxgZW6wSHbzFUlWxYoPglAGv4CpHJmwHw
P0ZTxlwwhcabPiWTFmtY0/hg/pG9AdeEOPhmLXB9Lgeqe/Kay5uHUjKR8ahCezc3clqBC8ZzooOZ
+6dl2veNJIyz5S2j6viQo30ZZUn0DuoRj8Cuz4JUPYhkDKHRoReYCqFE7IaQrjYyobpkgetB2UyR
cGcKbuwULQ/8el1Z72q6McU7m9e+ce4nalknTYdlYOL8GtDJT/XKElu8F9q9rDR8FvQmlHaXQM44
YuZZHL6AW5geP5jdmPtbJAQg9Shq1KGDwWrupJB/Vc20bXOy3/j469LS+DHw9km80KMOr5AphBGY
1ShabadhsxL4cnzoDknu4IuKSActPaVLneyPHBGPxneEiVeOEw8vA91+WhO+/1myvEHp19YqHw0i
Bwiea4nBXofgBNg9Up3O8EWvebmMUgnm8YMoQRTmys+I6iuxwsVN8/oiQwwltYV5Q0avVkd6Qcrk
Y9KrDO5gI8HOzJJa05JqCbefa5x1hfBMGPfAp92pdqV3hGvk3Dr06iOhTsovTwJkJV1/hlmPsHEw
ceUmgNZNM3qe7tDMYrCtx7PQL36NzxJSBpFRiNgG/KvpeGPnzTECnujVDJhYXwJAEsHh0YqPT1dX
k+F6aCrpbvJtTFlrzm2qYrfPolsidvtbnwArAkQx0O2eynBlUVZj6yoj3bmnB1FtmTl7p6rT06kW
pqh/47zcOWNx/czgHEciJCwH+ad/Gb3EoQTd6rtCmKFSxxZou+F8JgTDEBxyVWKgapPCVAFmOyGl
8Emss27K9POhGZ2oiuR/Wx5JNi5LmdkfAclTUjvpG2L8Yfnl9sP78nI0Ma7k0RUhHupaeIK1EErS
ydPIvtxeNVydrn89+uz3ePQpccwi0GHCqxv12CIno+pIcgO7E5in767DhX2oWGh+fzGYzRUN+/9m
Mq/AVhwMXvkShyrNCt/Cs9/hu4LD9C9hD2+oIQeuDZxyxiabHaDQ4uU+wxNwTSmJ9QXEqOoyOgl3
CJsFHAjJ7bJX5nAR17i4ApDWIwkA9NalkHhHr3ps23hGuPOmiN/21USFgDu9Gil7aWYeVKk3JdOs
HwXZJTkv7X+F2TxkyQMidxIB+vzfHHXHmNjw2E+wro1kOOqKM8aBB+k81ZT1cvnaERkmXFSXsFkR
W2HkZXDplHRWZZecQmKdEFz+iNvrXpZc4RLxhR3X44kNHFixWHNtn5bKwA2pPOxM/j7tqg5EamfF
wAaukN9Z27tsLvnKw+VW4ikzNRQhxuqqJe7b5kJxZHuZBznZkLwXkmECEHa2mxQuqeq5qWzHjCcY
FaChg2b+XR2Z+ThPbIdSet+qZ6ijCCKoUaD/PElWzojJkfwcDS40fMabonXwFxtzxreG5P1eTyL9
CNJLCB3wlRu8JJxao3sECOrseRBhGfK/k6YFU4FXC9dDw0J/cDrY7xSoligJcFeBdv9YcAfQ0/Eg
sE0D3nppA4EYRMoRibi4hMuSeRV8B/Jx5NnTcKFB6YX7j2yn87RDAMYNanWEjxtqr86KrQkCrO7h
bRKtj8JsDlrE+43TidEwZ9Rur6lMC5pHCAjLmlDJfp9CORVCDWjH8NRwBUmTK7iQ4prWySYfqRoz
m8ZuFLjdo3qnHkD6MJE5p6/Odx6Mj06RKJbZ7Iau+oVB5/hOeQFe9MNUghy7/1iOQmobjS8URtX6
tXvKDyYM5HsCAxMRTY8M2xBFX96f+V7ordWzjIW6HWFqD8Bi1A5PYh1PlS1XyIVSJ5SCw1ixvd1s
IDEEBUa29nis3mXgksSOS8gBqBEh9HrIs5smoiiDDW8z7XLpVrysoO3oaeBLHCONGEbRyPizOp0c
O64Sh4TwP7xlyupQJ9C3WGZV3jryN2p8cxo0YiA9Z9zCt3mlIA1gf+4Cb4GaI5SCP9OkRQIqzFdS
/ShPcC3yUcUODXHVUtOLVPsFTVumiB7/hn0eK638YsBbq+IlP3N8tM8ZYhC5+XCLff5ItyOPoPjX
/G1fWs5FQlYx9/9p07I5ODZS3a+IU/ymZCsjF1m51UtoVQEpNUZGZk+8GfXDTFxp9ajMZ1fYOO0i
45GwlerLxtLOLyca+l+YFiFEWm28PAQzc5Z6ojlEvhiBYqbuWWXSUR/xIKC5CrtBCGOOYAsGkRfm
ZiKtTetCY8YyniI7oLY3mB90BY7NxWx8VMGg/dccPgEuLCPGZeVH0MoDO2XgN8XXfLgfn9sXMWRm
QxxIP3kUd9O11e6MJi3kxGgxfTZ5Vc3Rp41tzOAPp9TGNfFbCVVwulr7DmQ9HpmIp+bu92dc403Y
mtBP9jQTVMdVOjySiuQzsSIiRB7IeQx9aCj2s1E4FWK8+dQFgCbdK7l4rFp5WkPX1NuMlGPdCtjR
l9vWidHjZ/YrN2YjppYZOg4035lEkp7JtwoB/Gv+iJ/RN8VPpbF7u8IZ5ztUIe7oEwBHZ6K8FeoZ
fiTYf+My+MMtIcPy+BV0qbDNwfaHEMFf83kPeY8Y8phbzM1yfXvBxtuuTcx6VhXvfbGmRzXaLv14
fwOiIZ+1qM3RVgXDfSa4Pu99yMhTwcrVpw8R+sanAAZbeRzojsAE9A4XTlyw1b2lAgrPedvQJQHr
s+/zee7F7uJH9woi8e4tGxMijCBZocN+PisBp1QCH1ecoM9FSPolwnCUniVAiRt6LNghlexcJIiO
xd8Uf7V6bz0dF3Go6SiFWOYCvZvy74LKG2ctze2DgqcuFj0kWXOOAFW9JX2cO7F/8lxmbgRnpS3X
xtnXGcNWk8pu6kwrdHeBDnpQ+ZA/itKqcv+tqToj5sr1Vfk69cacOeSZjkmHeJWkGgvMr/6/O2C+
lV3L01qpUK4LF2AYJ+eaPzAH+ONwXksc9G5vqmz2y4Do3rt6aJkTWWreKZCw48fJu6lhIc6TfUyJ
zlCakIDrBVeXLkdbSnUvlJKntKA75KOnAOv4NtFDkzaOJyzZisvRQRv4A7Ng3bG1+gx8YeyTN6j/
EJ6hUYD4xR9R4tzqLdMklFeZqKP4W43GvszsMSgQZI7+ofbqNtX6OlNwD1aoZvAYsnyE3g+1xyPO
3olxgFXYufMLfGwSVUZ3kkX3tCNnjL0yqGrt6apLdYj19zkGIaVuPlr68LY2492pr4DW2VdnA0kP
rSQuBpKGlokH3ZFzcJC3BCFkcqdi5uSlgmqSEwMPDM5GUzKKu+cei6KOKaOq6XERsXkCpZKHg7rq
/MTP2BKlWhHX7TCUTLS7CX97uw4P++obI0VD8lBOXackVUwuf2dQagleB3JEt7oQvLzVu+DrWZjZ
+ujma7h21Y0+GD/+e5q9V+YRyDc46QxQsEWhubsUxhE7I9jadq5Qhs3m9PJ96i+QOgV/APjySrW1
RCuh+n8Q0PWwRcTWNYWJLPhacO//svqU/K+avmZO3UYrvp4tr1vQnXYl5nyCJZaqD6EyCLZUZJdw
axaav3c1P3r5JVCZgyiWoqPomRxqVzb/CGsZj75GZaXhQ+xDdbakVIn5oXhuuS3CD6WFiZUQksy5
cqw9La1zCNN1L04uWrmdY1kX/dXWqXRjdpwZF0GMFefjFkFrboog+5RDmgSfrlM0LjhdDsCCW6Da
XSScCwtoYjuIaInAk6kv7iMx/AXALSeAzo1bmx3FS5HfLLGH+n63p2tHUiHFdGP9agYRwTZrpk54
IbwfJPzKaXJKSyRxdzNz5lPJDx9kFSN4aj0Zf1KYBtj5aJjRMFobbRatB2oObfuf4rWJ50Fwj2XR
HZB8fZFFjT5xvWLbV2BqaL62d6npXQ0UJi+ojpU/8Jo9Wtz7cP3GeluMSN+1GjHO2BJS4Xf/zN2W
6sYyRh/2/2SZW5lwB4blFBz//7zW4043Ot6XOJNLDHPk3TPzCs1szCMian17tonSJYq1VvwuaL9K
rdM0Pw/mHR61w0ACWPVVkA+Ww0HQQJWrCmUyHrglu1XXcLGxfKcUxDKBeVa9WJIDVDFcYmZPImMV
L77U22nliC8GgrFZbAUEg7fjaWuny2JFBt3ikZyIiiGAb2fslSAYS0XvAn4f1zhUvwVD8IW+ha2V
SQEvIGyZe0cOk9fHYyR/eKRXKa4OP54AQU+RvCZdfAmFwo2VHF2U+XtKrue0OZm7e2vO2v76zOiB
MS7Y3oJq/QWTabp3LXetm2Kum5z02goMthPR1VUh60llGGrtTPls+sYmHvSlz1dSmuMtcjtC/0wm
Q2hPHsU8HdFh86PQvHRnjmYjte18/A/zTABKiqr468PDIfdey2U19+gY8XYR3K6+yd891RBXR5as
iqIxFqWWdwwmlqzrB7nvOtP7RNUa6rGfca26qP8o14RVamvTnriJ9s5Y27xT51oW46ph52XCrrQd
e+BIP471H6gHViN977HBTRvrbly0jMEuKtoX8n0Gd56KlQQECuhI352zS6YzcboBmHU1bySPbKLY
4bQ9ytsL2Bo8lY26aOWguYD4qsQDEoP+runj75bd9gxctQfAQiZIlf+XsY403MhA3KGXq3Vq1tud
+rBKu08wM6v9ZXRxsfxRpNqx0z/mlBEB4gU2658kZR/uyyhYR+QLsS3UdnqP6GeHV/Zv3EoibLLm
79O44P/SluvkiSpzB1fCYaGRyCJzDgeRTnPk9Zb7zudxfxwqICN4kFW3jAghlj6P3kpHNcKIUi4z
xAKrOdX97eTOCj9TdTLdyNhsK07j/EItTNeRsPYC8x2nf0dncW5ymOGkKJkhxe6ewxgIFBXexFpU
hfwMv/1VulyR+/i6vq4jIqufVbVM6KvC+OA99Wc+Y+EzUiXYG/9Q4PyALrUBfI61I5KWGGRMjTaB
zISq2ALGNm+ytuopqnxsOk/sSlyUou5oqnRjhZhf1lAMEF7og/rhAqL1NnMn2x+J+BJ5JRCXB5ws
lfbfFr+rnyjunVoMeIdJ8Stwtucs7ldn9iKSXg/Sy3J/pVEStg1bPAjKsAIwKDhK8XVzrFidKRDN
O+hzGpB7/XsrCvJOAN9YUcPG8vxVU5gA5+IMNHQjy7Vho0R0872WtnAjnpxxvyqjCUR1rvzAGiAs
OafJP1MN/jdPZf3L+dhCTEe1hp0JLjFWKhYTqQxUrm0AcrsYW92fKv5vgIvxyipQtlxUDCwW97f0
vVYNTfLdq/Ds41ywPI+jsVoMh4nSURpGaWP84NgnL0bd+1wFbmLRlyLgx8M7LAScJxD/HYpxQ7SG
IeykQb0o5onpTwSk66H2e1wm5V+2S+SbROZwgnw8xiU3cVphVTQ8vfgITwzDW7SYjnGtfmwQ5EGl
/AUbitila6fBFDdALGzKxGxlB8VjhgtNWt7nlaMVdHewFS/1DFr/o3lO3NZNMSmEwZijL7iVShSt
LvNQgLC7BNsargDYLTLFSiq8P4xWxr1Vjy3WyyyEvhmKwT1t51qAtu/XR+BR/Saem1q0D4/BVWlD
Zm+mS3mUJ9zIUTMmKLCPzbf7wPUmKQm8NCwRdfgIByrkRrzSbfxaj1PVq3aQfpD5+4hevQ+qk6/3
aOmdQFvsY52wj2IPuo/mIZWKl/5SyhmBjAzXozxVc/y5s2rRxz3iD/FqysRoTAYGZUOeTwkGMYja
2EkldWE4yRf85TIHF82D/0MUG3LBTbpY6ZY3+CSZmFouOrI/uvH6ap+IlmIjpkZHYZXuKpILUcpv
VAHOsnBh71h6NwFj/gbUt1RAJpLfbQb0f5huh+Am2YrcY0M/Vyl4iYp+I/4v5Pyi06Zp5rxp7ujh
/j1ieqJ+ZEnyS3qtsmiDGLdBOU054TxFY3qMMHk1+MAKbS7X/rPrSBthaeXfnQ+Gxs0LtnniLaCr
rvndnxIaSgVRnMlmmNlN2qkPdNMTadsFbVN3NLWETw62+pvI8j9UFxo2p8Ec05SLDt0SuBq8TYSk
gNyMDMShJQs0nWqXkhPyQzK+OT4GlfIuxdc9LvByVAoWtJ5AKZT+Be3YjeAFfgajmCxCT8nnkaDF
Ul9wO2enEl6m7CWLRI8gC9bxpupyi6vKFnvNcaYasgsbJvpk52o4LHDpgEcwMAq4eaKCzJ72+L46
WQlHVX6KkrAdPXngCuGEw9DTBwWfH1bF/pTaTDtxkXbmmxBfxMz8p29v5UNdgxlNzOrxolH+Kms6
tbnHW+YmN8NZNUjCXb3+P2dKnSbCRlVbHf+9JGKphv2QM6YuditM5KqrVOXV89dK0ApYIyEIO2Zi
G+mmYV51HY42Sr6qjY0f3DCqwRk5K4wVUgkKc8n1AzKkXpdlBopP0l6M5KJmUcUsoL7hyKyLmY1K
KTZx7jfjpQpsoqcX7zSCP8VZjacyh58HMCINnbE8HQqED6ic3h3nNEIW290hNf2LKyfokclLfj7c
qOvaJPg8lGsRa8hOo26yBbjHpaaOZxC5SpCAPs/1PFWadrk+FZPkJ/9wKnUhVkVC13Z5EVlUafy3
hVYafodgw8EGi/LxCOZIkGmWVdJR4A2aVx9ulrs3k+pcPVAKlWO486Zl+IUKQuvGI8nPowXsoYK6
d3b/aIuKuaXPzySje+zPW3eBHRZi6bIdXLrBiBVDALJdl+uiROHQfmD2L87JwF187N0mEBXPLab5
rTKNHOaVjGuE3Qb558Rd3nnugY3BZTCmmLB7iIghaC6Vkakds1gEUgUVEBgtuAKadj6R/24MWR3r
tS6Ea366hqLkGTPf8PuFiJ/thn0YmXgwBsK/qhjFxXJu167K7vUPbluaDxS69mlyi6liSRgNS4Xv
Z+5tpAPi2sNDOSvB8ULXr3tG7Eo6Wk8b6TV9/OrzlW3zBxic69rOvxoAcJPf3gHQmgPucv9R878z
cAiVCPmKyCJnQJrqdwKQulsW9u165NkDe1ZPyEiRNhiPPk2VcuKL0ifpOGRqkdkzMSQczGZqB2lR
Snem5xSJ9iinvxqDwo4wS5MW5ihdNycJDjwYishSlfdhp4JQ/jsBSEP1/VB5gwleIIYOlo6dh1I2
pqh8nxQQQv2OuOu1jnOQgOSU+by+IdyYIIYZRQhDGSv/PBDBpfes9aLcHS6hiZVB05SBX7v2hiLb
MH5Tr+tnpXTnvUF55Z2eVOm3k4kGmo7QXYjprtBggRZfavO3PGevyLAm0fNoaFNqoz++bT5OZcm8
NVx4VdeTX7jp7nOIcNiesUbinkCXQHFH+djTdmM4f9jAHXpC3FcDSUJeSrmU6rgi4jfgRSlyoVvD
g6f7yG7iWer9ejrUdlNJ5nb+vi5EzYbyPDNDGfODiq3GqT/PkEcOqSF6GbdEu6SP/X/z/Z+sf5h/
JenoMPhn5oGiUCpW/yjVcucviTsDzb3SlA9Lvu8buGJkU4pdA3nAVFIAzGOatalf/XTXyOy7nrF3
9reCx3c+PQpJ/OKL5lXR5dVB8YK7hNShnpxFDyC2YsdPs6vScARDXqobLPxpBfkgBBxn8vjcVyw5
viUpqhF945WJiLkwevqPJJjMHB2DqxpxMWljX3wtYQIA99J9lbNoPAFWoYS0/PBNhkSQGbhNeTu0
qJ2wWfnnceMUKpa+sUjjbtQc5LixDAZfnu8HIaDLf8xK9ujFbeddaAEX64unGi90opqCpAcN0Dst
wQiVtgdi4Lc687lcJga3HN50nsUiN+wZ4OlRq22qIowx8NSr0plqPi7kRvBA2up5mNFPSv9xp8Ba
LtK+JXNpjUOBivpJ8rdCuwu8p81bNluTp1UfCmCMaYYV1Ic1X6YXV+XLkIPEnSDV3fRTIjMso5de
c6w1JRKUe1B1JeqDWeRP0X7/E7mjKRbcbKJsYyLqSRrbfdS1U+iK3sJAiPhM3emaVKbRaSunVb3k
osflmreXUSCUPaQrZAgptmf36iDFllD4sMDDptEbevbZ64+sdIETDDN1dU4d7kD+9CAIWdK4TBRn
e1dKAKGy7QfjgZuOAOU9Nk99+Yq19junaqQdBT89wbdRF8NLxJGrdZxUPhv6mF7mVCv62Tz7SLrT
cfc6/vX68XRa0YKFCwpl/820sj2WCrrC/t9+K2tfXg16sicJhR6nSt9Ey+IPZTJP/rJ0lde6/KHg
Xp5VN0Xwna/EPvQkTDw1gBQkXBWB05gqNlen/AGydO739AGXgo9HVLx30GRUb+UgjPQaZ2Icjklg
nSgfL7dAKb78YMMXKVHn51/3LFN/Rv3Zu4rrMjlG0YQH1BZd93yPBp+Hce3NZ8eLx+QI24f+0W3c
ikQTnaSPf0xE8jJoEKG/PW5kt4gUASmvoh61Xso2hsQOz3a3ZM0+N1hUp6PIDtqKT764voOsiAqT
G6thQhl7zoo/D9Bw+PS7Ho+/BKrZmpQte6/PlM6LKEMYKcBfImmeYX720R2K37a3xMcrXEyYjeng
pyQLWwRp6OoqKLXJcWtVJ6ImxLZEWPca2r4ygGRRhPvR4QWL7j+e5R/zWkqPG3zECasLF7UQj1tq
DyQQRyD6+9YCnSqU6YN53QfFKAU9cVDBj5bS0370qjYrlB/VUb9OPjqFXFmm3Kuq/1bfwdl1ZQOL
05AKDTFL9PU6Z32KEQ+VPbr+PJRi8zbqOKZrh3I+YOOEO7JxlJFM5kbH86IwWrZ0oX3/RSeGUr1w
QSCjedyDxaYV06TMi5Dj47EhHptL8YqF2Oni91FxBHyiBJw2T2Kj8RZYqaQk8QLgs9zbkUtUnmfv
9ZRXfpfOtee7NmTOnnJYsSnJd1q4cUgENC+r9ziDv3mHBlNam8F4ZdcHott7IQ7Wzf5rxJYufRWC
b5eJ/ROrwG8Cf5YKQ/M/H64lKkerM9wbVeakAm6blyuRzmRGxo0Fd00o020BNyJcU2apMfZCvSRF
J0xiYN9U6me0fClnoz2FNHjBkVdUbmzCFTDI5HMoKBPDwjnX78pZfiSKzwW/cqP9oq9qv2U8Cu8r
8eOBJ07+MHtDzQ1Z3QPLSNJ54VhBqaea+2/6QxsGKIAthyV09fRgYVxfFaTPSp/Qqn/z6yCYFSgY
rkWEwmRPYKKd55puB0a4R5ck4UzfSoNVz/enipRSHFqyKSjSsJTwAPxKV+/MyPWPEZNDAEOZuCU1
WzqZtD9Y1zjZQsbq8XhAUrk2ir00Fk65zBpn71QB9CvjfN/C4XcOouGE32Y2FAXZR2n7rhzAAc/g
h897Ql9yIlorBSTSRd03Ueh9Zx93oyTrNFxDHFP1eXerCY0T8VWKdOnLXkeRsyfOFotEICNx3aOW
h1MrKb9/JYfXcYVPG8UGJ20RJro71H8JG5Q5i0tvL2Rb+VMiIJrcxhj1z0/oesfH+daHunYsfFbe
gCXe7+cGmpmjzAcNnGMh/1TuDveQ5mJKfUl57ZvXa5M4LUhBAVDMked9xwjSy4RNpWiNVJqQXyeW
Z8wEHzM3sg0Y8OPDpFtBy9A+7SDY28r/R7HKKoLeIsM11PWItmyBCBHFcXEfWZNWRvuyPhtQCnUs
+LhJR+85Y/6VBd+2C3M7Q7C6zPbkODHgtYKUE4hHXNGJpKrGy/yuV7MOMO1sYxpsqPGoywirU33v
1DwvM4hZ+7AzTn1JU4vqd/w71zI95AJQnsgVdf25hvSyVVN0ANr3rGQuMm2ZFgOWfK3eOUuG3iU6
DbCaQa11h8l5GUqw/pCFQNLk7+AcsiJLWTFDNi58Y5iFg3HdF+jn370H7yfwL1Kk/9OppSaqh2x5
8ySQtrDIigfZRpWi7b9glveFHtzIZ0WIyJSrR5DgtTtF8ZcqbSa5XyukAAZPHa0bzJRIGRrBmerg
dyx/B3tQn9ntB5v9KJ+kWPahndvYU0Oav4XZl3aOjSTBjYlR4k9t1SvGLnZp8nLE1I9B+pOOGYnR
hs2/Wamj8zVaVyW0DABrmUhrfcQ/KWAF2fzTMAMw+6WXbvOUe3/irrw8nALyAJVkp415oyVxjvf1
Ll5MmOTdw9MKe0q3l3fwyd34Xs8AU2xdee22EJnlvY4Bm8MgRm/kkgmhjEF08f1iO6pydRMco4aE
A5iMbhC+8cy7PPcn95PRLLCI8eXO90YmhuscgLTGGvR2zokH3FwrNR6ih5/gNP7wLGVy1mphMkHF
z5Ksy9AFzHusc+ikMDtBu3db2ljlyt6ehemrb2XfLeaAL0fRgFMtF5OSYUP3rtMRwgyX/n59chNh
aHMy/hYnieXzjt08XTz97LZ3LKnd80Br00gq3SIJje2XB9fBZEF3U0HGtfAoIaWpVniAeJ9ynky+
m9zD8oo4tK67wH/lwO5ORVlQchkKEwEq7k2Q3NTX/kd5xLdUxaFX+/4X733Yfm+Ojt/lrWD4R9Fe
sZxKd/Guq1+skXU5wt09q4R2eZ1C7gBBbWTtZOHB7OuroBYgRMoSFIMYgmycKpC0AYR+fhGE+mb7
pjJtsUHViwyfwMO6fOpIRB5FxmtnkufNEV+ZEcBWEETG2u5JvJuSXdXEQT1pWfm+m4SiE3sZDxyD
6fiGE9W7aAcFbNzxflOiiYPPt6AZ+7eAhqOMGqDYgcXcE1Ac3+tFvlhlPQoWuzp+uu6XU9kw32tB
I1+MztHUsYtBUmEQ5tRTphflSSI6Vi/veT1+WIhC89GQdZnagnxOP8gBPsiNhN2OmvgSQJi5KfCt
ZCxY0pPAfNKIvs+naDxcQOe4Jm/2eXJ2ttdX8J6MB7M15nOlppB2Z+c9JYjRoXl4BUzwz1oNqFge
ZsRcTjbhWor3oGgHT20fY3kTy3xHjtCFp+6+LzmKzAhH00RLsJ235wrSF4rsrxCTqJuyT4PG32PT
zs277vYgHaFtzi/dYk0DbLPiZcZKj75+3OwLV/9/NJv9CSVXB8Q1ZzCS+Eh/SeM7CPvepTltNBa4
VbbCzZtOGVVWDFdHjJeQYr+xmz8PQKxC3B2uaG7l2+rzvqXFwGLnFZSwfganTyo10xakwUiWP8s0
KyR7Ov4vbqfHOMbCNQtdvfj1iZhnHEXIg90YhGc15zxHKwzaWpN+xhgYBYmIbgEzVhy19CFL5lU0
DXSIU0q+j0O02Dk2svO3rTt+8MIz/Q9PGMMjbC/GKoLq3mDYBuvGjB13yCqdJXe/pc1uxJNOU6O8
2Wq1sOw1OTyh8zk+IXTqxPDiHf/0mNYbxnmHLxZ9iAyYJPPxeYZdb7HqexcpRhMDB9MEYCa/NZdM
8oWETfzqljCh3vobXr2nJTN8mARCosh9iIGkSU/Uw4X/C8CoVtVKXEj6HTBV+DlBWaKYFnUoPFI7
UM4EFxITM9oNUZIE39eb1P0C0sGXeG8+Nv8iQeiHe50vh5LD1efeXCn2YY6pIQoRkAETxYheMq7h
w7QY6QC1n516oL+XlCEYBmoU7CWLnLMWhYwl/TZhkw6Dg9c+MAMNrX3Gb6RL1dcodkXcac5nnHQP
STIps6/mfbTsQR6mNa6rqhWq/fQyhyfDyVzp9craOm27GnqTI3R/Qla2STvIm3rX2w38hDuixTtD
iATvI8McrHbFSTFcr1xNcDmHHpp9Wd1rdv6VWfR3Z34xsqOK/oxOVusgzXOFvPoH80KP7DLKTJx0
kK2Ov2zTVk6Zto6PKw11RZe26hPI0i1cPzNViPzi2oWCls80Ma17YVgyeFSNuVcjXXOo4A4280zT
T66J6eAgRYM69ffJ8PZx/ZbrAcroD22rK/U3QDQc3Ls/wvM1H7x7a3yE9j6bubp9kpABg+D40mtJ
FqO10NACn7MnrYjnjOS8OkIunDGdKq6vY5aHc2s/L0RXoHm1MuFniFA8e6+n4tjv0QqEfjAetB6h
y07XOZy1X7vpR60SMOtreJv2xG6ZKW23GpE9Dh3WMn5GXycDbLDsufPNmlEGGN/QYH8ey1y6oQKw
0/hvEqbGApTis99yPlR/g17xvREzXu0r1DdXA7Qq6/PSvzyZ2P67CTtRCmoNxhLjh7lUIeRMfgW2
A0Ct8tWIFuQPS8MHSct1l+fwZun+YRe49ilg1OKT1f3mKPQpRfJz0F4qe9Z4pPJdYB7I3gPM1GYa
6UNk0jCKOtqNHUoWtXtjVQqIjAKrbuKNBA10T8pQkZ7WMy2a9JZqD9dEvHhGpYNX0/1Zl14l7e5O
JdMK+JdgpSJ+W3kQZ7rTUbVi2hOPAZC89XtoUqTFv0MHm3429yvcnFx96XDOJ1UU/oxTXEmxD6Va
4HtKeU3f8LyX9MmItpureBdlitx19jyOruROcjN6bC+yK3pb2YQDxp1Nfv2Fc721/cEiLLhmd8UZ
xKF1KRhU2Q8UzBVr2hlBPHN9DYham/CfaslfJxWpo0AoEUY36FAAWVk+r2zYNRGsFcNjoA3ieVdo
S5cHeMpjQF551ydVnyDeicA1SOfroGjE8dwO13XIuYMa5pCxjrMcPe0coTIj2UoDCtWgWoWPMYXr
9sge//Cd1KqYUXOl23Vh0DFAlfaZIIIRBi78tflDcb+d4nhkjXe/aEKHUcyDxVwBA27qA0biXOBv
XFNlujRrD6z7WOknZXdsfkRmkE354aozmBHMG+yd04lefx0L+9EiYFOtcq6uIEwe8LjRs/NsqRDV
khlVcGoqNF49XzB32iXylotVUgr9m8FbOeKeBtvR7rd5x3wBIfuk07zuVoChi5LWKsunna7z+gzR
zzKFSzN5tv03nrUUH2Du9bTnICi6/9ZA7pYLfWUdeEbVjWcFxVvhM9evAx5bHUT8gi3x4VyJFTKO
rCTqlYH6gCy1NcoOVMFBPS8FtYpNbKO1flwCkv/mRufulkgl8Vn8sguRib/jt/2rwmrD4HwAlTDi
Db86Bql7ZlwOZD1x0BFVtyhReNk+52Fzt6uQsSRXvZPo+uca09tHC/eB4qGtiJZlLsi0A/zT0D/v
lio0fIzkW5R9zh9SoRArsu+X/bo4LpDAk4poXxncIRbO+j7DfDLnm9XH/7FEAL3HMQyEYb5PpB3B
06VSZN/iPP8DC8V7bS9OlWpoIhtu8m9Id+D50MwdlPVUi9a8UC6eJMxFFFP22Wx8YMhXmHwmm3m9
iNAxlaAWwXMXatFatzzOhsQlpidjruAgXUnF9vJe6GpCqsmsQ1jzMi1skPl2qiUiKBls6cxPLgw3
YyFPcTtWU0H9TOzi09wbRmq9aIkh4puwvddSmjZHHHY9kvputMA9cZg6wWAf3ERnjaDJQxlZaSo6
RlPg1WTv6A6X0X3RCFEak1waTDnZVo0BVo9eXjjBSx2zQPROLDc8vt7T2o7gNlqtpDBB5gqnealy
L9UcvfiGcEY/TIFeYbEOkSxPPmbeKPLJIL5zxHAGYQP4urpKnxZaguJlA7TJZaaYdqO4jAMAhNw4
LLwOWcXcs8QwGiDms88n3EAF6+ZcPoEBuawKnPJdc8RDOVp6AsWIvjLYTNDEkcDLiGR+3K1qjeKM
Z8+0an7xtbXunEzCLuX2QvMZ6irckFprnl2SurgUk5ntPz0FCLGVfKQFz8f9ix1jLN1zRnuG1tx8
xJziuPUUkXXT8+Jrq2U4PqzzLro9wAQ1D5eyRJgPZGpwSkwiD4HQb77nhtdrRutMTD/ic5v/ijnX
LhV2pYa1Eiob0B+4f0uR1TAPQA12/yoqi4Zq5ZxTe3qxRL5+0BBp79IJvHmTw1DimLDz0yLiuM8b
rDjkCNKsr/F6MjUNq5iDPcwqt4GxkHOuxChZE3zcBxmQGrP5SIZibim8KMh3Bi/yKYfVwqp9T8e3
V0OS8bEclUDcT1bRFXTms1B8erfH8hZleTUNOC6ZoDKhmH1L1d7U5jV1AvABXvprVFyNDfVVozc3
SAy98HI2yM+SwwAZrVODugi1IINCXYkgUh7eupohV33iTRN/+8JIgtNww0sNueejPyfGSgLxYqmP
LXP65utWb19lIV4fVKD6aD+pE5rVn7k1Puza+80NOpDgw/v44x9sEqdFn2JwHSBU1MrTIfjnEXtO
aWsICq7PJZZ2KaPoH8oR2/Nddp0/F0Jtdy8QgWQ3YsnSsJbewrdJIjedK6bu52KWAG26phNLCSKR
UTxnkItt09qJmN6v6WNnR2LvK3MfahOxitjIZF1lAUjzLUKW0I1sMqqNiqDuUAXIz3b+rtg4tURh
Ldcg7kyLRe7R9lmU6izEDCpdXCHhWnThY4uNaPfA+6ualY/2yIw4RBlT6UqMSF5iZLiLiwGNFRSa
fYTUQt8zTIKKhNaVR41KD9aGGoXBGnsiyUzDmx8ZYYno3gNksrUbq/wnEn0CfdyicugP2wRwcmD9
8vt6icrwbLiV/AW0FCf/BPapZr0DzGIItRGZlfbi+Ga/NHVp95iFUP9/rO0F0qBIZFR4zTliPCNu
TpSj2+OUqR4Zv+Jjdltoin5XaZHte2iLT5L+QGPlX0Num8uhAAEPH72oQk9Kvq+I+5uDuS59KVJH
6xkwS7qSiPC/m0Ft0Abi0NYaadh1Tu/lLjuyRVicZLO+Oy7DQQTbK6Aa+0SKjrHxw7zIul3FeOET
mI1XuLaandYdV8pu4hJAJOzWmtpCXnxwv/16qN0hMUzEq0JE/tLcOwO8RF7zRGuw9CQecA2khRTQ
6SxPDb2ssBTYD+KY4kRH83PH10Dloe9zpSEqUKCxNJxux6aJzLRG1P6qesu88GnW/VUWeDLzDfD0
gtR/04U6EHNC77fNBMZTdXN7Uxu2us82GzP39kWSJvuYJLEkUPZvGFJTevKHiT62byVzK5QgyM/C
cty+mQSsEOjTh+YWR8IEqBZ++6WZ/3Nbkn49EKpf1OmWKj1jaHITK8PQdlEBKNxO6f8ZfGtpXP6v
zgV3Ka6uHOtmofJNXHxUxeofhjoPhNQkzUbgVCS6nOFaDiJfNe/CJWwHXEs354GxUj64VYiE5r+v
6eo7rNC/13N0ldX93ZTz76dVvL8hc+a6lW5ODOC1Nm9kLfuJAk8fvjNP3OInzvppNXY2su0NxC0O
7uqa7p4Gwl/wL2gqSkrlimlJGKCOI1CK2KAhejiGceO58VKCieh3tFXq3QYBrkHtzpQ6s0MLVrFr
gWSJhSkr63eKYDnN7kS13Hht6FZKMBcpMaEx4fXymHwx6tNNq4nNAxcVrG93K3X5CQxWbyZelljj
irJj3xIgkH9zWZ9xFqbmTRNl4GFKUEE3p4n8O/Bom9ITY45cv/vM0Ov3ZT5T1bf5q3DqJiCoX46W
Juy3znVaAILGeGcfXdQJ7HlCMOtxFB+/DnMeaWzZjT8YgW9P5Xy2+5sMWbDUoi5bpPXUuzDIDsBh
+buVftevSgvWIGlGFmQIITt1dZniRevwv29y388IkjPa23N+jivuZDuHDIVY+QemX0RVMaX7SURP
xM8d8QT4HJ1lQqDXZLR+9i7uja3vmx6PoPYH1rk22ske4Hzdh6xpcBRqLe1CcN9kyZloujYLzg8P
YegFQyTvNgspD8mLrFhVBZnZyJJ+oK4RNVDkf2MHGTxnWSy/qMhAncUQsa7HoRDdYRNGSSN6XfJJ
JghNjHH25rLHPdjVWr0Mnbkha17HYC/KCkZf0gUwKsmsMUJlcdgKHhqDT8n11LsGSOidEvhuZgbh
9sBPrfoBGyp/C6A1Ro6/OCcFxlIrxegwS8ApDkKgnjMFGSezzpve1CiUC1ZJuQcBYPaHKfjLqL6d
lGv7uHPtCkgPiKSs6coIDIrKUG4FDHdstirwf1niujIBc/2E5zpcXN7N+isHmq+Wcn6xT4Zu1S03
2gMIp+hI6Yw+A6zCue5rybA3n79veKuxBP7sVxwcBhv073L1kNXkXOspJZpXG2VbKH/Mer1WynFP
lWxLlV/oEjh9WLTgSS8yyUZlQaaQmzYtDG/NQOreDD2PB4B0hWRmF7OIB4MXoCZLvxqhuuwHQ+13
ou6fiSy1qbKyYsY+eDBDIGeuaKg3aPrI1lBzYA8YEuXcYg/np+wbOUqMec/FUIVoqtbv+pMDx+/0
pnJ6kVaW1oe0aqA7zL4us4tGzfyhnNdhQ/OfCRYpeGv6rh/2qOPE9BEDS1imtAXpb4m1wnqwLjIM
JXv+ljb2CJURjZhPOJIrBo5tQtRCSEPeZo0G+amyEPIoCBHdjRk925hCRaAJDUHKjIBBfmxn33ba
Brmsa46Rs1xMyCfr5B5PYIBr8nil5/jO0yr3JxAtayxOZJ+5zmGEbOmi4knwuUkKUBp2n3LnxH9Y
yCaK85WttosfIxQRwFwIj1O+iIjyh8YNuXvlE5xhHYk6x2DVtlMVmGvoDySQX78fMlWxU37088jQ
/XnTmBt8skkT/5zsOqdQxxRxPgVJFWiLb9pkrozMcJoB6pisryd+gMUyMwq9UlGq3iXQlhd+bmUl
ifDes6u5R5m2Jq9fVURZTJ9mE0nBCw1FGu1PehNdaO+NZEif5t0/eURYFfPmGV+gKAc5bV/sCj4y
BAyxo4TORVtsBK1RerEvXC7wckxAwOeZf6dWwdbkff/SkOdw1609j9+UFmh2dFuAmCq/CHZEOsC6
PGPyZ+xaIBlWPz9/hmVFkcmBd5DLAlFcb1peHB1DWm++YP/o1aVbKw38kmy8epYAHcQDW78LocVt
ctJ5KpdG069s7k8MOQcFhNBr3ze2Oq+aG7YalCuDdM1jpdoPe3WQbxdxo6td6Sq70BMCix0s3ypQ
9AuBMIWiNtL9cynSD5PdzY2RKf8MXy+QpTFGMruwcLH+UxhwDSc28USI6775CUgGZpUFAhXc6IQs
k4WVr+A7xgYWs7tgrMBtdYIrm8V9iUpjN0OLHlrmnEpEu/4vEv9Y5KV2MqOUJauTJ9TxemsjzyXd
s5Cszl16laZWGXA1cd/uZLyajBRcUvgV89RXcaRsb/qRr8+VFKsLg5zE+DDrtI5FKdcdDbq2c53h
LU8nmUlKmPIYyE7xjdd37MqInQx8i8tKK8eC6ga8QxMHrpEsm1LjX2d0RkkopoHLcbDznEdn5HdF
/qX4NRuYcI8pGDFTzlK7AzbmU2kZZmvIKz+X2IPPHCXiRGyGLp48R/sEU+ChJxLDmwbsu/Hde0jm
3pHuO+UNSe2aiRK569fzduzAdP5RpQx8m95fATzqKuP1XTG4lLnJhnbQUgWYEnU/8OBWNtOmJOqY
/e9aMsLVpC+1qHFe88oZ4U3WTtYMBcwv7KRIZz37k7aq20QRRxo5+bhgTbuyoZ9Y2AROyZirfRPj
iip8dPHVdxsk1wLqrHWvAl17Gjf5ySOaHUfbX6B0SXtRwVMWucWmwDbeM/5k2zOSG8naHIzpqMl7
IrA5uRfxCyngdFWjDVOyyB3zLOxuKnC9e7oAGoCDYEcaiEtaYoUNz1FIrAz7dHoXgl5577JvlXRT
oamtrcxxJKfMeH+14ibT8sh7qyVpD75y+k8cGUjYxXHpNK3VWxfsM/FTcKQeNINznZYDRz/LYhS7
Nm6HSvp9Dx8GjJMnr4NNrD7zfQQmI6ns6a1qs+Wh1Xx/DRpx8Vix+MbYGVR9wgKciwXWHMFSu3ul
U4AKwvoRBEI2k2n+fxsdqUoaSWfmZQFO+tKMLvRbujnpMt2/tzMnlX3Y6itFkv5ja/am1aRfzg2J
PlN+bWJbkIc20jrS8yUwd5XpuHOXDKWGqyKcfjyFkhwRZESd5Cpnr2ya9Cs8PJIY9IKj/BNT/oSP
0644tCBRXRB1lu4sEhDrk9R5DGyqeLptGwxP4K67fm7lkvGgFweIKX+oUIVHqQB19MSSKXNHWY/y
wGq9HTUTTmDmO89kvdgIRN1fpp2WDKQQgSNEiU3M5mV5QFJoYLPkdMWrlzjdzTMeKHk5tF6JyIFf
suFJddQW6EPOR0b9UxWNbxyEd1RTZJG9iFs5ANTCP4OYBs7iO40PdDo1nag5GGF3QSANlA9ZGowM
AVG3VdvH5mLVNqWx6pKDSm+7iaX7qK+Z7F7As18odgLNM68E9dy+sL/65eH77nHtikvyLrmFIgGl
0rPqV0zi5xF7RrvORpada+mHRGexHA7keC/ofLE0iZvCpbp0deILc8Fm9g2D/cxIEQ13XP5AYjRV
fiMMQ8Dtmqtk+735e9CCCZHvR/ncp1jLS6s5b52Mw9FmoRo3lf5ljvXm+ghy0/CZPfBY/ko4SsdM
V4lME0uyl7ToQnQgE2auJRBmEdRSKq9fMyj+TVTbL7jMe/TQQmo2Jzk1v/pFYFI11r2vztfw/dyN
ysgAfK3F7DgyjdQAOrZCF+RV35QGUwtq7dLfzsSStleUUmXGK0ENXrIAXRnB2v3V2Wkx46e6wme+
S5ALOr0ZQP8PnJ7RthFqgyBxCSaEltPAM+TYARjoZoQG7tiYoeM5byoiD2WjE9rYiLEFhcY6zeZX
2c/Lwg2mZtiihh/nBrBjjlJk5LN945/EDnlqMIRHj+pxZzvpEO2gytgkbZBUvRdNRDVehGiVHL4J
TyhpNLn1uRnamAHu2Igb1WGlmtn86T5Feh/w6cClEXgEJI5Vv78VVRKNvcQoEbWODm+aWSqt5eI/
sDFkjQI2Dc3zmnM5cSHny1D3PSFjfH/sQBEkx7/dElJdDpA1C849ZXeQiR7W6OjD23MuGUwLWAj4
TXgI6N90oNDL4XmOs/hglfOcbwTpf9t1VT9luHGY8ACxD9JBDxSR2SYjShaYVQJ+4nmVY0HY3M0B
LfdQIneBa1VgRa1ggWFRZ1i7+asrXfNFnYKRqQfEBDt/PeAy/S8VH44RpmgMTK7QNvjCaH9u22ft
3O0caRMZhFyyoa8iFNEvhF15P5Hw6wKlLmKsytf5Vwc96n71iPmnX5hrC0UXTe4g+l3HkhY8cHNb
Eu2/tL6GiYybMrhtU/QWbUUcZ2ByQsIMYZoFc0yD1AWEFiY/dA3XkffSqeB2OPUoBs4jbLqDYAwi
v3rPN+Bsh2RkJxk0qqQPMA2WtoqazMB2gIpKSKYl7kCFSsT7jZdWWFiz+kIccmusnYl/BWmkCzz2
427lf2EW27ojIO8cl7CCFpTME5FUy657Eord1qDVv4dP6Wl6lAYqbIGjHIE8AEZ8ylCKDrDCpGsg
kdX8wgvLY2VfIQWMYP3ieqUE035C7D0fs+PibdcxJqSQvwAgUR9iuAAuDmSGAEdeVvtSIJVW1QU5
2bfZ9xduuuD8Oy5RzRG7szx7GzKpNzfpAg5/dOHRyjWSfJXn+Yhj2tIMxIyM4EQ46z8nZmSAcPKw
ZvCiY928pdyNTnypm4yIowQ9GDbyc+YmxW+reooU/IwBdZjwrRf4BTLyh6jPOvKZOLH20JVRy4n4
OMjQsZlEE8YlkjbJ5wIRW5IgQMRSSxu5oPW5TKbs7QmSoZWDrxwjjo+ZYuoGWRne5OnNN22Rtxcf
/1YOjqctIT5ROlA8wIrNDUNMRlh+8Hy/8AZV+nNx8sBbZaMV5SNpPIeaiQDBAGT2DpYzrMmnbICG
LAsMj9QhVt1FOgcjjOmpoVa7bf9ILj7C3XVAQ4aXMiF+DTzeVkFEdbbIkiUMcR4WPgLVhAzleLLg
Z0uyWTT8zIHl5PAsjgUcZ7poZcB1bkim18Bs5qe1mk+VTTIBsuQv9mq9SinMrSZg3d8LCOpUpncZ
6SrFcIqTv8WItjiKQOvTMF4sQPhJF2Yd0D8M0udroXDVszQEKE5YrQu5W/PSqOlMHoEKXo+meMui
H1Qy2mgEQ4uQXb38o6FlCFmbX0724DFwcopj4X/7vrghqUi/0mL6odsNXjywqHNtsVU9xd8mLat1
4cAMwt5X1TXr+U7uPfIEGGq6gTvHRR7Ax1fbioB7kzzwcxIR+ctsyKvaKf+kj83n7Cx6KPqGJjrw
vmlxRglQNjoOMaKg0Q5cfvix+uN2YMzfC3kMthW8bclpKkuB1ybfByfS+AbQEbQ1K9SGLege4IfJ
OCSs5HkgH/Usq5xgUab6F0eC35/qPNQmYG8ao1uFykztYqJgGNVYOpKJZmEqHuW4KYD5AIIpKeik
NIp2g/DOu1qfPjheBnLBXDETJ0vlKaqBFaqCjSHkfKX/v1OduY5mjcdXoNxejS59iXygsJtKK7dd
6UAnYfmUHpJw3xzevzzFWYPScPZATzPLHwdkyWqTGbU2cRS+oMS7rsG9cRepqWoNfgGBgchjoCat
/DVGvoRkMml+eV5DZaBAotqPjaDM/tnI/C601sKkAVY4A0xvE4gLWUe4U4/hNCHFAEhaFFkIbq65
kpV/PPGdFintxX+GuR6kYOW2v0ez2hFHBNlwnOTmSiRuAO8nmrF6fbXDm4DiEUMhfkzG7A6ZJHJk
lPYNgkGuNVXcXQ+OaA9/8+Nam+0oT7FqV2QNMSI0y9aP+3/NE5bIvJhAV1pamWwl5p8rVUkdILZq
rDoLdENhyZtyI6ZabiX0BWvFGXm67MfhVytlbHtvHbFFJbrM86ZX7aBptUqpf42SB3iCZjnoP+3D
hMVHnx06B8DRKOv8LBDB13bAASuKgSL45ZW4s8NxV5mJhY4hfGCbReAIKassy0cX0mYdQZzH9lgq
0QzkEkIeN1qNqTn5vm/4ddcd83COhTypHH4TYheS3yvKS0/hvduDa1IdyHVQT9/Y28iAso7l/kOi
LFrBvbRaxFVk6YcdUECi5aM836onZn5bZc6P0QgkPmHI100DkS1oskVIW9N3ONdT4x3glmDROTB9
EOksJWdItmtDEcO+eNta1SKLJabwrOdUwHLpe1Tuo0eLcYezfEmpmRTMG3JxPZLf6KWGvOwfs/rp
bnm/ZmWpMJIPTUnlfEZFadB3DBq1SAzv2Tqj6Z2Iiv693pb+N7+KGJbNwXFbybVpNlzPBvzsKAGW
52y+L5fkI2A5esW01Xc1Tqi8BMNz/pgIn1rDpQMgXwLleehbvFu+UcV4HQBTj+dlGfwk/CCjn0LZ
FxWkMLj/ABlbA5XuF6ntTiMYmfdXI5wElNiIsnUue8+09Spnppfl4lkZA/pdtYqb82iCvAxphnr0
JG4sTdMIthYuQRwC6z1LoV24x+FGC+yYWTZZmQMuN/DG81tfqB6XIHjrKDPd73u3h3rDqogzCnBv
Y017ltx38KHTQXltVW5vbUjiS0I9WLEG9rBGfWGBJnfBpzbRqu+xd5tztzHUbD772IChY41yr9eW
RFSzpsYflsbN31JZOj15DXltVeS+PAqvT7R82fKHTNTvemcfTXiuIXJoruP8JFoavP9xyIGN5AVC
F4gbBg+z28VW00bwQXLtUQPtYA/bAZbyKjiVG8fLTfSDwcSXzwziNW6nCzx4bzrY1bpxPA7F/HMw
cKR9KYA6E6w5BhlemI7t2iPGlEpnJwJOonCi5ayapIF0GmLOxq9X3Y0Ih+lQyxxeTrVWzjXh152i
TDFJMYp+o/5LNHq2emhPlb9nS0HjI/Jaw9VgH4yo47Uu4nsiAk87NzsZOaCZuD5fIPYkNFOsdngQ
DYkNMnuV6JN50YiDpP8VbAyveQU3RTpBeGR4lHWsLoetgkRISjYcx0266A77iPDC60N+/74I7b00
2blWShK0LJeMCQ2wmEKkY7xYSSJ2crcZm9wzGj6OdUgtiY01PjXSdFhtComiJIY/GtoIET5dQjwT
zc4dcrLCLsKoNcP25PEDY1fFEWj4q9nxf6csDzJZeLa30qPRiRL0imhAswEs3CLzgbpG/dMU078d
g7l5D4aF3euf90gtjBkb9ReeTWJzNxfpKoDGCmY39aLdoDXVpWisKWGqYnrLv/oL7lHD2yd/iLF/
RNs9O4pKdOVELMgLO7zFe+k/pLg/85hczQykaeczD1bNc6iCcroWpDAENqXHr/s3LEbSd1tcBk6B
oWJKz1UpGpPsBxofAtaWe7GFdOyUI3duCNJpSxq+Yduz4RyQR37uSUrJ1C0JFU4QUDR886x9EFJA
kej+tvH7zkYOTHDuR1zwvSU3iw+eU80rMaOKbqUbjdZ7pGZj3Af4HR9MdgtwtzUAir6AfdWcqWbJ
nkpkeqpCNOs4+nN1g8eWvM8Tq8QQS7vj5gsxTnZFUYALyXxznsaT1Np0Y9ANkG09625JE7RYlnpA
Lz6crJmb93WQDn78k/DB/2y4rlWqkZIvFoRcYiIlnnDRuXmnEfcI93QleA219ijHwhNS4szTq8u9
LAjqNZEVEngoiWGHNsDU/35FYfOAjXxIKDXj3qBBxmSenMVAiwKsN74nVD14U6xleKx344B3mqUQ
ORK3Y8t9qiibOZxYSnKAIoalzuIHPhwfUwFfJigw4LZUGUjzXpP93gJngs/DhPB2Q8kBFZ59mvzN
tHNig49SJoDB09vRsZrULXD3uyCSwnVkLbHW8+/Hs1JuBs4Mvn1NDFkU5f2ytevDw+Bvr3jvHUs7
nKUyc+p3FYt+HO3b+jgzs0EW+/bQRNSocN3uNHI5ek3MZNuzETVAf0WxbVxTuiaBfziZu56xEIgP
vaGoyv+hkwlm6saxNJW5Vvsn5oEIC2ZKw3cIPSYXDmPge5scJ/JAziNUEBlo9hklcLAvzOjM2K6i
/MjwfZPv1i0A0r2z22qK+QMvCc2FYq9fXNxUk3UykHY0DHqMZkXYjm7aAdfyURw0PdNLwKEO7Qeu
gvxX9SOybCTyIkh+vg8Doa+an8nmHF0i3HEOMDXW9RLLpJ23UfYtCSNinhYizpH+cLxilENsGQVl
U6yaY3nr2ldSamgCk9ysAQQ+BZlgeEKaHdcvDMw37NWZFtAOvjvBDMzpenWlxkmPqkIm3nCmwHjr
U0pq1nM1H8bYLFJKZdo45TRW6iuVg4nGZDYMTRQBW3GVTDVUkj+CNF/mRDl7rBv3+xMvOI8cX8pg
0g8NToeLPZU3uSAlR/8y+QlPLxi4Gq9EOW5WS5kvpwzYx3K994Ufwb8XrpbfZyZJBMsE3Lr3Qj2n
JcEXwAw9pgO2p5tZvJmhdKHEk5hYMetzrqMstIR/9sgvE158CsxajJGf/vYXFrE0dhNc7ICrvvar
SIHOwxAnY85OTJv/O6FJghFU1RWBrEMUIhoT18J+iaqc2z6sWh2YThl/w5HC9CnkoBRunXJyySlh
Usq0okq9/DAZANP3HGFvPlO2zl/2bdN/5Pf30IpTR4GDUOEUMZowC9xcof8aq4VRlfENZyRWRDKL
E5XzMSbzT3TBOwAf+VRYz7roYk9eGWuXOHrFSO7I0qIUVKoLZGRNg1u0ZyIDoV27Qxl3pEf7OaL7
q1/jITw/zSxD8KYp/vcy1jTb2I9sk+baZ2yMDIq2Dvczftt2IPm/OJkFiFgverc49BbEp4o/NUn+
RcoX7MY+gweBmNzMvRuwV35Lx25HzRCIc7tiYj5rMOf08IEqoboGKWrmWHSrLqKKBhU8w9c8xPPL
IzqLcUV5x4zQ8J1JJVDKV1OHXKbzTeg1Ju5WIdtseYe9GKPgX+OPZqX+rHFWAv87pkl9cpTanogT
UDGDHeM7Q44b5BWs+jzu04H+l6IWnfvdDZgJGxmynvmDC+nyDBRyEup2bDVon8+UoiTK9FaUk4GF
JY8SVGR9u3cJgeBCvPNFITpo1eN1yliZDsFIzX5a4ROiEWcxs9NuST18DSpNPKvO263dSvjMbxPq
ltKGhK5P6WcMFrrMEl1o0G3fZfXdUXHbJ9EB7FppPt6w3OkI4VIA8I/KqcyLbsQ51bjnFkGG8Be7
R6D7AmvQIhdABJbyca7If/DYMGPNCHOFtGmpzXQletpei2wU3vlO2lI1hYByZm1n3//8HLpl6JUm
E1kFOaEUQaO60VXg42IT5ZFgaxWPIIsU8lvsO3pXMXuEd/Ub1hoDgEJHGoLjnsaz/LNnhf9Y8MlX
0zNBMuE/V9iYFGlHQQgh5o7VDP+joZ4BMmBwzu+O6JMSMQMx69plMM5JnrZfsGvs5Sk0nd5X+jXv
S/5ENdkxmicBRmzGbzah6KGapSRIyOOJXnFInh9tenrwRkYwXM5TNDgNT7sZgPs8tfZk7NJdWT/y
wANPqvALj9cKiYITvsHCUtpnY22+cmPs9bqOkd1X5/ESy/PwMKAJyR4Fkcp5wIQjW+He4riR1hCq
cO8XOVkQWwP99CsxOqNeoOnoO1VNNjLI9hSK21+VaJMITuv9y8WZqNQjlpJnlK19ovWRkXibpW/l
/x4IilAibzFzSeeI67mJrczuO/ILPrxi+xjikOqRI9i5rB8eJZAd1rTtgmVy60jI6GWrh1wpsSTn
vKIwwUbwJ0/7Xo1DBCDGlbzGRFoyHfOb1KJwQCSXShX0gWNxLAcpxNVM8OMv8iL6wf94y5lOeAMC
AFo86QOomsBmMVxe5yLZsWuVdkAmtPbm1iN4m+qSdY8tY5KDDcq1/SBRrv4pPz2dvnUn7QsUxSl2
kIK8Z0QChmTulkdIxA0agGu1YeNAtBAAOvEHovN2kljoxnPh0jr7nF+1Bu5hSmZVYNtDX2reKdGR
mkQixe7zmD6vqLy6ZgIn/kdycQcrkAZpo4FSOpDBtqStoEiA5xYbZNFxOHGs6Gp5wMsKTKo7CNRx
tVNAOXL+1/b3uEu2TzZw5gx2exT+3t9RuuYJo6/546a01Q5ry8oSqa7uFY1ORBz+j+yO7q9M4rG2
Bkhw317j0pWyh6f6QKj18m9O7k/jb2nmdAxarE2gnbi909cRrDywobbZ2/uwyGPHeSJRzxR1pE78
j0nD7GJ5QT5l1XP4YcH7MvfQLbzPM9yxlCTiXiMVzWYfP0UVwDgeoh1oxXU/bxhSmcPGtHWuvXLi
Kgto2yarL4Tm0VWpL6bocAFj0F2gnbh+RzToSwFjP0j+W/mDMxDRq4johGeygZGnKyuhJij907hV
nwyWIF+ZPyCF0rscv37i2yfaHpsgilrjIbbCB8ga/o24GvmSpDQZbBxfFT+0LFJP3jEM+b8tq748
zy9/GKXz0zrfuCs5Einj48iz9OlgHLbpMfpCwgefmst3Sb1dEL/60O4Wj7F7lqYxZpMq2D/3aZ1d
KxnPC9dawA3r2GZHeNc0ruh1EwfEvOSSBmDkgK4xzaY9zGJ630h8SYAEIKWoQQV/NVkXy/T/wP2v
z6y6zxuJI9FXuU4EgePEDVitYk8vIKO14kVR+791DBuw4NtECedB+u812MXT44sdl2woWo2QaBFA
9HSEgtCMw0Kwte7m7jH4BvvqqwA5iWprsg5prdBhlEN8K5ZQ/tmbzLkN6XakXNvc0VxQI/l0G3hE
HaRObMdBmIcrBLgRuEE0YgIZjXLNkjEZoni0H8mEF+G7zJ8p2Ub1uInGqlilbq7pavHIZqdXIeHq
YYjyfPf2lmwXPr0tjXX0X+Yl+uQjxUTbH2e5mpyDmfYObirCUj4vWEFB6m5Hd1tr/X0yiJk+lDgY
NPxKU14YxPTmK5tODtthldR+QO8g7PHcXNTu9916wANWE0vRBc8yu3dxDnYStxFTBIIRF7eSCYyT
PMZ0XabxaiChmG7mLvdd74iSGrVprYMP0HA2Prs6lA84LuuU4+K8Ga5irrlgLzIKhIyWM6KR5Abw
wtFK7ehXQXBs+IajcgZnWHW5JvloRNlllUL7Jt1dVnF2usPJtAfJQsQ3ptVC4uTVrJttcspl6YV6
iLBJ4r+cDgX0Wri7Y8WmyqFFlpYJwBBlrZo/yJOe975foVEr4gUoy08Uxc2Cv9w+KbvnVqgmco/s
59ZeuOsnX0nLLBNzDAsveDU+KfNgFIaTl0kNwxnOzJENxI0BLrXEnCg1awU1LGmG8dBGBLaR1Uu2
zXbtoRB88CgGO8qkmnOV2gKYXa4Zc2nq0QwCjmRfOObQo4wdLjh0gm0t3asVsTefcPMkrTEtO1Vz
VyD0BCjQAUaJZjtrAUbPcrr0AE0rK0CSM/7fcpngRdbXMqguFsDDDxrmYBk654XgSBzcRyOXrlmh
DEgwob6XC60Z19eCihRssefa0/J7bxqCVYPoc67gMZV7ClWe7iTePN0xNYYXD1oeN4XWJjzbx58f
4Ews9miHfJpRVeylhkPkZFzBpehjIeoLh++s/eM/Yy9E/1oCmNdBCBAU3Z2rEyhJJVtt3YJKAF4O
Vhcfi614XDFsqDaMjXzLXf0nhNCZ5lbogwVWgHNyGltsarYVitPZz98d6z53sOAd1jyfhC9aqVk0
JFoSvMKhFhlFts2gYdnPwZCK4ttCssk4Kt+sfO+H1eXKiepMsju0HWZ/OhRZEGZudRLZwEygjaKQ
V7Z1CdyFPHMU5J8T8SmXGQCX28h/1Fr12zpdjdhKnUGaFgk71VehyL/WdNZgzt8R+xII+NMhg6jN
Hjcfv7amkrQjx8zgz8/VnyCrVsuZLPwuuFh61ktf+8/tFs0n4sJlzVn6j2/he7JjAj7Ay5noEZLE
xtBXOtepH+I8TJrcHLmjKJZib3jCNRo0vTONJE3aFxDz76HIo58p+KD7rE5q6/3CJxlr1JhpBmme
hF8xExMFyYNZFhsqzmdol3PLwpSZTcX9Cfs1K5izuRjX8Zq/jzhEAk930qLxzEbzPKh4ND/a4QT1
wfPgJWteWa1+gSY/CVRNbwveJclkReDDOGNMgLEQ1S5Fk96Oms6msmpeE9lHry+1Nk/Of3UBA1Kj
HpptZsGYGHf7b/R0dnJTLubM2iuOcSglpVB8p6RCZunjYiFS8Qs+YLAxtjyelO72NQtWmyW4vvNQ
D8Kuo8whdc2X/6T48v6+L1r+h8VGVqCSnEcMB+BtIHAutlO61GPlhYC+vB0Rl6S6u/oUx9Mq9drG
ch+vvBwH2hkmBnNRswADtwn3sb5iqynJEqTydM9vHHXY/vsqtmbZdF3xWkED+SZq3uf3ffKs+N4z
fUdqAgBhJ1X1cfUBR232G86Pk/YETie05VKY/Hr5GBQAb1ZYYGeZw4k4wWbC3ITCLX8H7RxVnWm6
MHURv020pQRd4aKpo7A0V+LoMXYZ4BDMhpbfRHRIjb1vMXdN9+GkA68qMGFg/yxZf0twFSmu2Wtj
U2w50YPwqK+V8HqCWlPBvcsOKoK1yb9TWmZbo6A0/DPV7i0vXK335bZGybNCkZIzDzA6hXpZb14q
0En8OMnco6T4SDVf+kwRxVOnRiAMUkZ++TYt8p3a2tGmlmxRAviB3nI9sqpvyoqnSdAGQuy/ITUB
wdlmtioM5YWefQ8C2XmNUfE7TkU4sdSJbkubZFu3XRgziZ8yrUtosSgTBSarGP/rtPhdWwdSrHKN
RwH1GgvVZMfdLqyTm21moFRw7mXo7niLhcHRvCnSovA/WIk+Z8OAdxb7RnI9oEljHTIy0Exnel0+
fwQsgWjhF7xbpACyYwZL+zn3XVoXgL6i3bxhLMX8tyux5UFC6Ue+MAPvxTL/PSIE8x5pvBbVP9l2
ThQHMHruRSVF8zMC4LQr4DLtIxxsH/zMW2+iotQYOmkLvnvsmrbbzNMdkmVNZdrWuow8nRaEtxXK
NRg0C8AZR2Vm9lzr4gBZWR+4kjC4nDqtJL0tSK+pnOo3q3Q7prz0o1kCVm8uRw3OItyH6WtnMLot
JGr5gaT4W4qeIUwQ1YUBE3N9zWXq5GfAr1+XdhmjbG0bjwpuWnSFl69ce+2mCCA9yXRqWFXnayR4
9h7FDbrG3CraE18BXoBNWB6LNJtFlwmNNmkhvwCEsi3oQb4BwPSKysGnansuoD9igZmm7wXwhIG6
LNAj5SXm8IJ9CfrpU01CfoUbhXSgOXzJx4+IBKlZ5VoVieqhD1f2jgnKnEpG4td8xThahlk2yPDG
xzfXeSx00Gi8le/dOEF66cwqJamOgS4ufUaZfJXJK1AYiniKlqy5p4mIuDk5UB7zRCIGZftuzz81
EpvGPl/sL43q5as8VddZLXkSvCNRpR7k2gDtHHCPnoAd6rw7OzEtNth8rtj/bRTDOrLpnYzbV6Tp
gA0MoFEDdwJIsdWFAokLtw+y9RHiJRJOIHemzEXk+WdDvGHRopD2XvUeJGDL2H/bFwP2MCdzzTXo
ldRUqySBBFUr1CHRrgrnIBL96YUD5Kn7rv0/kQLGklOCMbGEorw5BTH6F/7jEwji2143d2hdzIvU
G0maJ+2k4kRYRH4igcfKcnAo7+AzPT+VmwkVAXapkpJSwSIwdmVZLWlfxxdRyOgrhdOAVChPAib+
hno2VTr4H1HiKUeVmUlSlN4MT7Mqv5q00+a4YqIBUKJnQKrFPS5fWoPW3xyp1bb9r5wrtCUlqKsx
B3XIPZWand9JGSUEYYg4ToFRgM8ugiNZMZykc55R9frD9ZWYjgnSAQhxkLI2+QwkwsSDsD6n403+
yyCK/j0b29zrMmlgcaS/XB3//c6Nu1VDSCV5yNZwxulSH9PE+8VZOU9uWoBpmuOFtTgW9+2U9b4m
apWyQ5/SAUE8cbnWrl/Wh8cmN+eb1Vnesx2sNwgT17uQlQSeyaY4X4ywOgNQiqYvkBzlxSkEnKlK
Dj2HgjO84x46tenDtwPb2v0uXevFAEmr6HAPhntXBxa9gANJRdrr//h0Cnec5hjFzp+Ykx5Dkqui
vH5cdCkg1GlxaAF2926EDyFP1tdck2Ux584d6qx9Dkyh5YZm14hTHFHFXO2JbtM8WYXpnChFRRMz
OgkMlUdwQVi0ONNpjyFo8bKr3rp0VcqdJTDP0Ff9BiP91/Zy/1d3FEa0EnzOiKXRVhY36Au8OX3x
3cOlCjcAq9RMP1Afy55mnUQVC+KD/PadytFNy/ceu0ELHaBzvUU4BTLa2iLV0sOOCoatYTRabjvx
47s816O6rWTjh6FStaIQt6YvX7TFCMebCEve/FfnmVh2VVygiUneCxB/JlPRECeVacUC5SvXUBIl
B4z07wFJRAHqAWypMqyx54Wj/diDBJB02r+67HrXLL6+Qbt6vv9rTtHEzjHxEz1pprB6eIVre45D
Xr1smnu34SF2rMnGk7jt/Ee/jXutJQDNx5H8pcZhzLl8zR+wZ2VAM/ywi7uv3Gm2m4fvhwqQDJBS
z25Y0ekii281N2VeLz9Xw9Jpr+Fw8I9d0AeY//n9/p7262LyWIPkxEfHI3LhC2MbFRZW0Hz1ukrC
fXx+rT3+l5qbKu6RRP8pn7OHPaJhmgFvclBK1LnJ57CC5fBk+sEdL1LXLuiL8u4PWLcVZ9Ue2Vh/
1eoIfx+Izxbqp604evcN+aybVtDRJikMvvRoHBPRAlsH5LwnHrZq0AzKZJ5mN9X1x3aRTXV26fBY
AOamcSPrPlxjqAKfaNyracXRNSo3tmvb4ciBAegsj/0c7hTKfUIcI55dAxZ8a3w7H+mQXl80pVwl
yuZy8h6bNvMnBeJfY2WDKqcZRWq7+94lBNIaaV4VVVZEe1i49iLdJWz8P/H4tcb7SPOnDAcxtMtI
hBtlaO6zSg7JXOsEyP4/FsUv8fkX7r5MVlCkWwn4u62SmY+9Way85pngXP793ZMHz+NL5EFhH2KK
CME1wNSvZyJlPgwcMevkXyviina0OY/MFe7cYH2rFk5M+/xDLQRTo4+7kt3FEaRIp0s5rlWBUFhm
LT2gL4VDftHNIeLh/ucZc3/SJdWBS9WZSRGY/g738KjHyVNo9GxDpokXJStNLzY5HbB1UTsOBYpc
+9iawUJhKOH4Z2UmJ2znxDmTBSHk/qj+eoGxVEdYg5G/IHYEPvqTm97oFgQiX51VR3VpXRFpTLMy
p6yTeHgWWc/c6MiBFxxn+IlS4AQzSIfmGc1fNdabXrv8aZSvYie6pjRt2hU//KkB0Dd8U0664QsR
h1JECIhAPAkJbV58MvxQHrd78+kY761VbDEF/7x56KevqryLqAhS8pfvOYybKAVqJRuqwtlNGKF0
WpeWrLiBlPQOWoP099YJjmVj9SvK4+b7sVJjmSK6WhdjeFu6chJCCwyUr+6FdmswJrgwHuCne9IF
DsHEm/J4n8h455wPoiWtYityZMtHtEhWGxylVzdnhOjpYGSLeno0FJqI67xEdrWfJuFbuPPGKwEs
dqmcuZ+emeIY6CRZEZ8JbSrs1GD7e03lAQtZwna5FMMY8zzUDk9/hKKQWR5pwIDurnqs9J7tFopq
c6Rr/1N6eD781Cyfv5ODGpq3wDI06kBObg8KHRKrlHjfa0gxk5kWuSLZMna83709UCpcsIXPR92v
R9y62jvEiLKfUlfZRyNLvungxpzWtFm1vsZcNoJV0XJAZiX/cYxDB6APoKGZuCp1j3KWM8fNjx3H
aQ6o8Pilf/VEWPu/yCITuAk9awIsewtu8n/Ii53iz7JzwR99vvAni8S0/l/3kPh473Dr3KbroQA5
CJ6qiKvbRvohazXgEaGrhELyH1bq28XQt/ZteBOP5y8c0zsVqS4m1XmTWX0USkpJEcKEzs+mjJyI
uOD8nSBGG0dzVrAP74kanmZylgviczQ1ud+uxiqMrS2UDFLA/Nc3Deq5Ymu/8vhMFvZuCRMgPzUs
dyV4TcLl7qyAtR8kXqSXnAhx+xmtQrgaCe+Iy5+IL2kY/UIDlnY2+/8ertNNixqBGOcTuTzhNRtg
6JShyFD0NnioACE72Bb8a4uSlxtdgu7EavuM9AVtTR0i/mOxOSsJPybmpW1B278rv4LfIXup/56d
vjOMHwkjIhg2QGBoq4I9heuLJhXUpN/pXMoHXXZe5WwjNZo/pV5KIrfraDfP1ceZ6txCKkz203px
PmAr/n7IxTxSC3ol7w2MpNDlgAcqH9EuXf2URlAsCzqaGQqpJYkb9+lQrNapBDkX24IX+CDNdW8d
QGThe9Qe1eE6I0BIMEAY9XTqdDH9XhvmVQeSHRM247Mgdfw6ZwQH3fr3ejVNhFmBy5XjPWVO46HT
qHj5+Ww0q1he7LdKUHcCIvjwTumVGjRtlKLmf3yqhqskg6EVSHO8SmvxYDbNpgiPJL5LfzcPHW8u
PaNah3gmyTmEO8kfNf1EENB71zE2QseDtKhX8gya8+DArGd43SkyQMe9JXqNfpM+clNrjnlUs94e
8rkVSriblzP4W+OoHfuHigivWRT74o4vZHHQxgNWZAC1e+Cp/3GY9eWio/ujl7LnI2BPhoZUD5kz
0oz7/FYzfce4etVqtpF44xawqtHi5HvNdh8PpjGysic32OsbO46Xh9IGses70FDJHpXdjOr5FpyQ
SGgvspcNGiXPpZVnT+kKAxgoZbYnBHJNkHmnRK5k3VqDLfP9asnKgoAuK8Q2G53edd4JOS7DyEvz
dNxNTiAq0/YuX9kT4zj7vRTjfLKTiC/YIbasS08i3ybchYh6JUqDm97vnsRZrb5MB7Iwhb8muisF
rUdqGRtI3xl7ggmvB1mBJeiFiqtJSvQUEFnXRSj/Sk5pEqBudd+8PakCd/KlFBypJ+9kNNzwcskc
PW2WqOp808KzHshst5aou5KVzMJMGM03rCa9K/Q6WDYy2/UqxszNdChx7Yb26+1nMGdWevyVYw8Q
h8QCoUaj4y63HhOu2LC7z1Mhp9YqARNFmDLosUH+K8+sWaZouX8Edzzz07bwXb6k1xxuNkeroVKY
V/f6wlFYgC0tus7e/Uet/jSQLID1latHMRNvpvAIoY+55KoXA5BUsArKiB+Roso7+L8yQaUyU6rW
6gmipVK6pTt7FLRMMibrH69rvMg9xGJawfPgq4RwUhIUJesFJbYxu890BvyNRWnrezAc9y2WIzdD
joEB2RjV5sjKlP5LnupapH0qDy0zo8tbZ8qArk+Bsg6CDDpTgIKm+4qTrxJXe8740mTtT9UY+0PP
rc6I/9lTte6ftXNsjKo2RPZ044xadZoLEcG6MMndwNodq/6/mpqWHnZBIHsOISSbGQxErY/f5cTo
Bbq+JXN5DdkqgZuYVP6FyK49iEBHmyP36Tf+Q0rMFNuvr76JKJ6C3f6KjN9K2XEzNf4eRjX5/A1h
lTfZE7ZKLLsbDLPiWf2YlJEOEEG0O7MGBz6iRgcPllqY42IlvJYWx9sdfaByXc7PiU+zzsz139rm
zaVoNoSSObdJ3LJKMx9wmtFl4E0vcBosBf+FmpYbCKJhIRtHk2AkJ5ClT/rW+nCmb0zvoSM8Cbll
iH95CkAi1HzickDako4YmjvynI1SFGm1HNTb+aYDYty0CFO1F1bJ1lb4SUtrj8xEYarLV4ilzXLZ
cKer61M5BwxHBoM9o19CkvrN53FIFVo25mXeXRJXvEOqYXrC2tJ/qUox8QxyuwyU8ncpCg7uty27
YUkXnCAifaOAFshtyRiAaWzQJPptncOcvvSIzAkaGNY59j7PeEq89jedw6aWc9SWnmoE1OYr8Rjp
KBIYYCimlarwsNoN26z+ijGeYmKVeRKT7/ZSV1cMV4phSKA8pl/kVsdLAWWMRuZIWhUHYdYkTzEP
5FO+s4FkosX61xfsEEBJ/doKs/avMOmXPc+KL0mhfD4kbCV6ZSfmhmxz9R+ppbDl6Ue9b61lfP3M
hVceQg9jGdG7/GW/VdlgOS61RNFyPBAilgExh2exXbetTQJjG4XkQhR8iZti7e+qx7BY1YE09zSx
lDLCNvu6mdg7CTzhZq+DbLpWzq7o77iwEbC+TRPCCVc1NRbL8QXa6W0dP+/MvlGiusVlif+xpIof
eRBVHbXjDQX6qXd7JlMwBjG0HEErZtNWCbNkEkvPHu83J8660BShXEJ9bgPm2uqKV1+5F67opSGX
tfA72qp9JgdgzB5/tfkvYf6GzYfCHd2OmTGRoBp6xAYiGbOqkh69A4NVGUNNsRtY7Guifui2HJ/q
255Dtp+KKXqr44+Pe0MFTiGU6Sww/fnuph+pDiJwSBV9BnJImcLfMiOuvfZwOjc6zVUQkkEjIVWK
Yu78EvlV/JyFc1u4iM4LfDabeqUw6+Bj1lWsYlnWbfIrqUPlK57Qlp+BbCu11gYAAoM1+kWfq7dD
BPiWY7hQ870nhFBOm+ODdHM9CZv77HruF/MUb9zIbPHkKvJ/Nv0Lo5M8Pp2j+1c+HUPrldcLDg7x
FuPlo1rAQ9bw7SgCMkO0PTeEd7v99DzD5Q/T0WABOvfuJYxmsW6XNMMhVK8i1lhk3Ij/eQh2FdFt
CN2H5xURYbGcFHOXT2EoCUGuFtAOI35mTHRnABtHSbhW0e5E6SlZwKjh4lCUOaT6MHSsnBl6xXvP
cav1zbGfT5tWuawl5YGHJy6veIEfd2FC4CbBmCbcDRUxUU9logIah5UgOd6ul2KGlCFyldj0bU9K
zxbWsvavfMHCSPheNBoqtQXz8fMoxiFMGUiWXYV3WIlhGnAovwsqh+aKeYpNEEuqeGDvN2Go/KeW
Gu3r4BQKSuQ8d+YOrEDoBPB/+EBk2Z4fFPzgGT0QIsxFhvL68sDwDNQ+cl5ZzMp+H2IKBgqhOhmI
dk14n+j/lk4XTB8XFOmPSlnyaBn0Z1WrCyl4JE6chQg+1CUau7w0xUzuu+SpSfyldXo9ko2rluz0
z73ndsWBhyukqSykAiWhihJ9nJLjKuJkSUWvCVYI4ZhNJ9EPbk+VNeocJsGlXpcngv0eWECLVAno
snOF5qZjtnOanY6fCph6ws8nnh9hPMmBXm2p08i3lsOlIkrUMDYC4n04IkhXRQvJEl99eRzPEapL
ey+ZQ97yyWWhQlN+NVEEEqhb25hFHAMgydFad9QE6b979FsOOFHTcgAAmaG79abRmbJqs1IRELQx
6n9I1I/4avv1Sf/nB/3+9o/wKEJ6UWgeT6fem8no5uuaAPL7YTuJeEhldLxNB/anYd92pYmZ0Bqc
nXO2lWwAm9oFa57BhtYHpiBAmNQ113IgLRaem7SDPJzVZKenFTaUMQXwmJ0NL3V5gT1aeoE/ybVp
TE+cW7IoGdxBOlRtvJ/3y15oPskiVzGXajCkZSR8mXerRaYm/baJvh1/gYeiihfn2VHxWV9lQtps
9FFG1T5MvbxJ1/dlVOF2w26mVNdM61wxYVpYRUKAflaa7RYg8Inx61cWa/PZjIJZTD7Mo8LCLrU1
T0IkWNGfPpgao4wobMZQRx64eHbEfuOfB7w+7xoIf+0K6m3s2gnzFeKJZrZWDIdkvonstGWISKrv
ajZM1rpcVd7VXLt2BJFOsY4OvofevH3Ew5hZ1zQaxVsC/uY7+ljsOiZLhLrEbDnX240uxw7DhewH
R0JajeiccYxnBmPUiFDOW/rzJI5zjB8IGGCl4UfSfMr9UfLk2X7uWnZqNpJhKrw0YD1dN7jH35Z3
sjhnoUr5ipvjzV9ayOdnOymAAnnLIJ+ASHT6txyZFmUTX494ISbUDqr0Y7msc8hqK978NLckZTsD
A6/kGnjNDa6q6R2xfQlqn8Cb4raQCCFZ/T9xQR/V3gIIQx9jz3c0kSjg0emSDfEplTZEiQSPNs1r
6nONQvI2y91ufsikOSyWiu7EY+NCOvWgZkPJ2frXS8qiIjQ+xPNaVCiQoPo8IZmix0tIXIvjDIO4
cvt1Skof/0v1kdM2lsatuQjj+2PiKR4caqvid3KMaxvT9ZIUWmpcZTEHLHBmA8G42pdJPPMsyOJt
zw0GCxxVJa3bFcYqNrrYns/o2CD+ELtVNx6xQdygmwMlg2JQcsSGZt1zndW7XpR6jBUoPgdQWugE
RQxcx/kLXloQhHUey/LrSseVChX/v38ULVkU4Fo66nsTZ1CQpUdwLR4+MOZF9Y+NM0rKoh8k6x8x
2kSRRCeRRa9JmzVKjx7ilFrWdeKeAFuBEPxK6JHLUlWv3kHI/1YKBWbCgdDvlskrPxp+VOqxuX7X
PMdKw0nRdhntxFJ2YriJIZn04cT3dL5S+jCAs6tqfXAajaw2k7HPYOkwmIcrsXzhlLaAAKEw2EIM
pvriICeauuNo75ohIvWJyiX48Vm25H2SFcmCVAQXVFGGfsUnjkcFvkh9RZDWNEpoHDL4/zkOQjA3
FK1zMfjwTdDAnhRTolddqyA0xJobexZTsGpE8vDPL2dx4AelzRtTJFnx61f1iqdOe7VwPzHqAPX6
SrsH2lfZ4LaXLZ1iVi779cX1fBOVmFPKzJ47wQziWkrdkYpF/wINsZxCAccRoTCK9E+u2iyErXu+
X/HLiC6L+hZQBDlGfdo1hNZ9mVl/TKUxd15QMTcG7hjxomoUPMyE5W1iko43gE1+R0sYgJzGsA2x
gHs3hZsF1njLU/lYcT7bU1cp/otl1L2m68mRceii/RyYZ+99ywVUBuHtswV7tTmJUWvNb+e/ws2T
obrrXT+ESzHq/gsAgAYOVB+QnasBNRBlu7Ouxoy7O/b3EkzwZLDlxFquEOJNVkSV23H4cTzoD+Ds
yDkuc8kBxQAX/N//niDwqqkt7+3QB3YHTlYE4kkXI2WrZG4MuSC8EI2YkQIthyNtTtucKD71qJAr
Prbnk9XfxznnGL72M0tGjX1x0KEEFpQ01NvehHX6o0x/xekI4EYZLtC7jDTjMPG56L4AIl4gLuv/
ZxB7tSPETuCt35/EDwK21KuWSzWLWmM87nT6+GSGMTsSSYsX9gBXVxemBRBNd8UrXif3pvMJxcm2
1CTcDkpG+USQg9fPIzictGQv7MqRwrDJF8ZRcqVMOvPTWJPjUW9Vl8eGUtIHBD7+uYniHsye3nNX
1rF8fh/tN+atBJ1e9tpWtL+J/iFN2NtGLasH1G4lXD1HSs94Es+iCNnB9Sb3cGoqAOgXo1zaGjza
jO0YpvuUAcJhAGO42EnDNSKK/4BnrgGp+yZnwdDtMWzobsyMwVfFpfUAfcbOVV3Y8kdu8cdvSXQY
qIyA3OGgO6pbEgNrK1K/dnK9v4TCEo2/AyUO3A1OIqUzqZlt7htZ8qlUkdiR8zQ41SlTMoWuj4Rh
i42SXSCpsa7IPqnDOdxXDl6Vu1G3YK9S9r0d7DlYyQbqYUa6e8+VJeCfnoqAb4fvROBJJ38/aYcJ
AxnTEPk/zZNCkiwStPE60JZ0F+bHUQ3O3BnKmghr/yrabmypM/EqVlHE280BiAMXOozQj7QQEWkm
r/qHnjZwrT5DviJrpFosPCXzZJOgKUZcZCMdblhCsIGFH0HVYFmnKQG9c29qNLfwP6tb1xhcVYoi
wsKiEJMVzRNgAOxBm3e/U79Jbz7r54GfGQG4F//+b6+l1OuFIPFvRl7kOLZL6KBo6d7XJsoijK0n
oyKefJBxso4OFcRt9R2z/rA3DjZpiskjFEyJPH8D/YodUHmDIg7N201cUdCGzBCNfYByDxEx4/T6
HuHBTIYbjzybEcUUW/kYOBLYIaudA7/TD+7jPlg1VTpGr1KqpyDBBsuWeF9HAwJzKhVeOQ9gPR6M
tVTtzY6+EkMb2Jj6xs1FHoznN4dyztCUrN0I2YmL45mjxNH9JifFEs+Jbjm6ojx/vx5/4p6uR0Uc
01ZrilFtH+TEjWuaLZhCwQ+li2yvfDuxYCLWKSc9/rqjyluhk2QX3vpkOzLA/LbhKNOvVcOURRhA
TlwnsqXLRfo0TFbHPz+BHpvuq0Irpm+soMAoWlxOaHUqALbU4fnOioq3Nx9ZWsTI+gJTfLCP+1s8
L8QAClg0LUaKOUAVwC5hKpxbAXCh91KtiK/UudwK8ZvX0rLLR+1pX9UYpnPRGvU7uUld9eOD62UJ
J5PERT79j9X8ZvbhavejBSQFURWHx79987zYPqVnTL7AKUmYbr0tp9m9t0On5rM5RLyPhKtNvWyv
cPdIJduz/TkSzxyw7+sdCq0x7GsnwXw6MpkfSu4u+jbIXBta+WvoNQqBicKglN88N0XZGPi+rIc1
6FtlmWLwCmA++nSjVbik+IWt0cZW2HIGYlFKSA/NRU7wCp0/Cd5LyerZNjHiL7os1Kr9xk7g+f56
VDLHy+B8JlNwwCg4cLzsCXiuWCRE3JZU6PNGcCofoj/TJWEb9pnZPiOZ+aAMf/gm/J7DTRoH0PAK
ySnc6gu3lpUY5MKmK5dsL0G6lb6xdtvhByzw4KN4wyyHvaslh7L/0pJXw6JHAGG/f5zaJ0Z/gNEY
6vWhsgXxPvsUZY7lVZnMCopehVXr05Q4Y1qFqcEGYHVHuG87cS8xLoSWwLcZhAHvZB5KtOApJEFz
4zztDERzQYSmNRwWG04+QitHH2uUIa2WTrplydVTNZQUccm2/R5RnfPRuONz4dcdu2m4p3wkSwC4
mcidXXuUorOakU8I1ZR+DwZUbN8Jdli7eUwRmKuRjMFUReyCClQbhxVUy/LwxkF5ob7Mz5pVzSPc
tOXXezymAhpGGYiOovGNhp9tLkjlKnLet1zFWUi/Yx70kbrlgJXS6cXf5VolLjyvpuM3exAIw4+m
bJyHmyR4k8hyZgl100F4fcYLm8uHn/kFjvlvO/S6TGDKSUGtKa078E1Dsqr3t0lrZ3SSQDXQty7s
Ponk3XR31saPo2fY1aUhtH9KaUIIs7Mb77wnSrgfHKEpk/APNE1rDUDt21Y6TgMKzJ9brTEr24ou
suhVyUFhK204gNLzOpOMj3i4LRZ8JzlMqNzbpNth4dPGVP2lDy/RXNKkV46Gx1oKlWo6jEI5F/hH
RcsTX6Xep7kw00jB8FMXkLFSkEGWNLxERPlbC6EFR8FZBeRoBtLYh24QMqn+gk2d0M1Ks2R/QiXt
vUyAGxjijcqtqBQxwN58BZ+3PmfIPZqWfi/TjhxsO/oDINy4iH5cwrC6huu2BOEImBd5L5uWhWlo
kht4mBJoKoKQgtl9Ybr6zaAUpVbi9eOmZyp3DiqNkmWrKrjlOOLznq6+yp86ReRBhnHSScCvBcGS
dDbH+Ypz1OPgUVxatxoG4Q/QcVxt0Ug3JeI8MgE8/XgWWD4uWvEx3deEh6JanEOan75DJ4EaSSeG
UkZTZ6y9ng81oEQBdAzKHGPKuLD84ujaIuzHrGtgFDt3/AB0warpaZv5sIJ2eswgWRp+EDG/O6x5
dm9op6oyyK5gIBDZDqfFL79XJOX/x+/doIt3oGhbYFrTURBFIoJj/3GEAwnYbV7DUIqHJ7sgRro9
YnWNcvgNmEBaDUL40Eb5E+s6lfNbe5w60f1iTXgaRGGDFIcnZeRhEZxqNBTdb9mvJ+HfcD3U3iOa
U9yDVukpwYGdtuuyxHbi66bmWCozayflFqEtW7QcnaW9CqlmBqI/84z4BS5sugS1ihPcJNdjZJXp
fGDcg7Bmxo80RXFvF8ZTR/vnDT5I1W2rlEhrv/uFRAK50bBJQBatbmRJkq+pcnlQPO6O6vcvHM5Y
w3SSGOfMzsR2cZFOa7W+fmPlTg1YZV9+vbDb4XMpFJ6Jwk7Z6i8g7WZbXgm/sd89GLCRtS5TmpPD
e5VZgCP5eSdOSr6ttlFydpGbC6kVf12zK10DaQ2S8JUzo8fT+Lomodn2qlBlLPnMcmglSDE9V+CK
W68mz9Aeg6eDgjj2XjPaQFShWfs/kH+5Y9NLC6yCHROvZWdSJAv5BklMmCrCQKEfPkZhIIjd+l2U
bhYU2t99WBSf3rB6tQV4CvADGWZUPs0zaM7o4Fjoi/nMaQ84Suhg6+1UliW8E9EGb8tbx3g5DGQf
kHgTWvvsPl8L+IYiLX1LGd+hY+ufq6zk2/Zt/xzBF4+L5SColAEVGdsyR8JZJovSxm50nZTQaeZU
iHA0JSHhPxiFrCm7x/N8L0Y4S+WBvX1q+rRAAMewR9Io1vm7NUoHBHNpGJyA7ESiDrn2ErefN7lp
PSxPR8sBsVtRpwSSffYxmLlpJVMzzPngLzHxxvNe3DHQRTemfrS3XfKdMce1dUpcbtr0TrocCspd
NoNXrrT0qZmyCujyjaN6O/bPcx6/Xlw6PA6hlKIVQ83osC6PrRSw8b/ymFD9cLDZC05gfe1txldF
ABln+Y+eP3sA08ERy+L5QmIR7Zh9OC0XKlnoRe2uJYHoQpN/ndwdtUODEdekA7jsLrHtGI97hquD
etvBtoaGgvkMWfY9KMxfIQ6P+FgKVHA53POmQFKU7p53eKeWK7BmHn+q+QLJ3Ob56NbAdFdABm9v
yT8Evc9pgH9FJ1AYjKcWsTIKkT5C2TR4EUeoUYLm7pOdvXNKw3BQFi49B8yo1UDMWK1suMec9jaP
IwL/9wjAWCvOjK94LC/ArnBgwmNu5OJOYdhdlAINJAHGkEs0mJ/ggFRZklNdeeUA8QTA+gcKtKL0
+c/kMKtNaDBKYhwwjLuZ/QZGszzaOaSFdvrlpSO2NC1zfz5V8RlhLq58zXCOUWnpEyluNFHGsoGN
Zy9jpGXnUa105LOdvWpcRqjoPoCpiChgrLq4ExEC+vEvHRg+YSbqQcYA0wbYq24Wyk8lhDRsjAp5
fs3ckmsG3Cts3Dbe4tIT6EaLHWbsmw+mZBhp/CUsVNvkFT7n0cWQbHNmDJ+dBwVoX9uMW1WEJdgl
ZIILJuyZnxYdvUkRtjqTJYrDBK4jayO0D3zR7p9KTGsMNZqfC53b/G/gbagCTKPh0HyST1LSGfcp
mTygpzTjfN/DAjgD3KK7EWH7COwl7XyM7faiisBge4D25FqWN9Wj3frOvffs9ASsZDONzr/JJVSe
7lU6r6t/QTMKiFhZ7JO2mltn5oUbJ4TeBLG389WlNMxZz+NPsUk3iLd6ZejrfYPrbbFMK56Ae11O
X2HCw2Bg40hOxqHkrHGC+nrr+Z10G1ooKGKOvlqZUWZhH1zNcX//0MitAL3adrTcN2IIViVYugBY
IjfgITrx2H41wv1Cejh93bBEze8ywDUZ//1NpdH1F4jKTO2xVSQgM88JT7dqixJkYljnvXmZu+Pn
2qEQb1ioj7NYp+esz6MeT6nai4DVJm2ZRxttSEXWvUSwt+A4PJgB35J93pjErERLWrWRMNv6Ludu
6gmowNBhNJm8OGTZq+bngaR+Nl/XYl/YniRf1WMp+EhaDgM0UJgC3DbM9pkNKxqmZNQV7+qaSHBN
gJf6ZMfl567qOyARp4iN2TS+eebJoCy+2whFxK9B9PYicR0/Ndh/N7ih04S7OjpxnfqRE8hdl0BM
sZAT1LDh1aYm4X6WlGbzSoKauq51TLxNbAQnfmFxbR+dyYSvl94W3sMo0XiU62a7bDDHOW0m5L7B
uaLmTEsf7qIosdAspb8n1+7jXefqj7wIh8mj/VvJM+djXqL8VGKdUM4ZnmYU1nqvMsV5VCvJ6vDH
RyvPJTH5mlQYmeSYtWvDDklooy381y0dgAxFtFAY699O905+9qutzGClYp36HerKmkpXECmKwe+Z
kOuZ1hXbENYfNx2V6A2RLoC9PAIQBwPIlane5r4KMvVA/JF7vfhOOfxbOhC1pvWrlcshuN0SrqGT
Xd62576mPiJbfvUHKP5xDkF7A1GCUVxMyG/c/UBJZZ6341Vy4hJ7ELf4uwLDO+RnjbjSiIcYjHIx
/x9bQ5FCkvndwrAGoNbZS9Rw+LMNMIdj4ccgvMI8dWV3LiiIgGkuDr4T/oLe6NocKfzG8jo8ugyS
p+I1b9acRcoLwUZV4ybxB1/dcOkchKQzuMTA6G3+LcWSAc+x5z8pxHi++MB5AyUuyKH6mOfyMDS+
IAfTnB08PE5y50AsnDD4JF2f3KxUnADOE7Mh4iCszghLMLHwl5g8R/iTEejNNKlwckuwlofaqCQX
H//6brAJ0UG8+QmPMWoga7LSQ5TiU88RabooAsIlQbG1tVctbCvueCyH/5Y8Kfkb5SdU22KATSoC
gAa9WVzPm2/pqikrRTSB1VPANTCOU2+RJ3S08Duju8XK5jO0mNYGb8krOoJX1d+QAPbPYwKx6vQy
rsEQx2dJ1uD1MyDUIEc20BiPIlF/3Tr0vWyneWnBngRGvCqJQITQbsneXlSGbhdaazNZYaOJDIG8
GtIXsVRII7+GEs2j9CeNeJKBdDOc0E0s2Auw70yiHBiE1DSUi0MDosxkXQ+iDI7xofDe2NV6+LBR
a5K9zDYH+3uqd/CtKnhrjuyPvArNLqlSN8fw+ZfRM1f50C/2pc9vg8iKrG0uNvwVx5qmSaQdca1b
Zfkfks9OCF1ko2Qv3UPHtUTgzklBaDwkz0Gj3jVwct2AmRCJs0n1GcJaj+zcxuWEv+8LeJdEnQ+D
v5KJRDaTfN6AiNWavM5slwcADgFD+CSLMlNg49g7YJMkro1sRtQpLmQlE4qSiX1CBjPlKqCHuCe7
vxO6i3jSsCKZN1Z8ace2o9mcWFgZL/6YPUeDkbqJTqRDXD0r7JM0hX3n52Nd0vi2R/gaHAZPpJ+B
UFAUuReflpA+eBtkYGooHO6Q7GjJozehwMiKhaY/ucPHEUjHDfu+RS1+kAdwaPy2a4ZiBm2XAv89
vUurxfY9ibCUMr9YMKr98ehmpVCQt6GMTMs8Vbamv9y2LaFi1rwgm0Ckpq1lsZsXAi0eJHefgwWt
zRwtFMhPDYii+YoyO3pbQqhAWK4/SCHBOGIXr6yn3l8YOFBZ4ztbY6yLunyEDUC60nVATKkkLiR5
8XBvHND3U9ZynVvbjd2kUUbEDuIurKz9rdcCC0XNGKDZ47mn1zJmXuhTKOwXAo4mIV74Zyty9tvy
6cTG7CBT4bR38rUXhsKULNHFlfLgHHSCyv41l6uNG9mtvN5VWYDBfqsSDVHsL429yF2SLGyayIk+
GyVCdVJ0lOwmSeOKg6pV1BaIoifnjgJYFRMwj1n/bRJ+pHfJjciAoBbwKuXP38cW80uw3E4mijgT
mbLvUf0VzeGRARDhSiNERbxHKJrzeG/nVu/qog2D8Rsq7VYbvwXlu9N6ggoGl9YCz4a4D8m+ovET
3F6xgZFb4CbswO1xxNRuzc7D40v9l96R2RNAoBGGpcsKsiJgOUaBvHtbQShhUqBLKgJiyHZGmhJ7
aPD5VST8U5MCna/knzOdncaOtoel78fvtBsQWI9C+y7ncuM7V+KiFaPl0iy3ZSgtNLc+lj4BD3za
Wq8RNmJS1wS7VjyP9mNykP1+uo2imlXDaAyivJU/PhqyVmdnlRAaUCVsPRWhu4OKTu999DGRYbTj
MntLQVc2YGLh4Honi46lN0MUGmoWGR7ii2b/jU1akIW2yFY9MqUXqesQ0P1xKwZRFTH7J3FQt9fr
L23szzDLxE8NiTF0mxnG+qm9NxZsLN1WZb+fzkMko3YDQKdr/WuGdygXbVgEaoasfyL3lvJh/Bev
BqZzPvlR+k0m/bj4r+N73o7NQ6P9kK9Rxy2kvgiTFS3d30XOylqvaEWg2UrG1sB+wKqW8Ci/Xh5E
z227hQncIBUWMNv30SrZe0UjcVPNJPdmvs6ulQz7L4LoJITPAZGbjloP9oOkj1QTSJTr85JmJNU2
ubjKQtcd/9CGbaJKx4omS2Lvu1ShMBBSMyIYmCZj1hjqRnKBm8Gu3vW7H6U7lGTic5J/aFBBUTub
4bnakBMIcnDrgvQXQIQYYr/ifmPykexxQcMaMYI9//ybR/6zugvqIS+k7NqGaGvj8T1qAVfo0PqN
mtFzJ5OX0mmiH1xkOrGBOFAymqBBqLdyd8HS8Z76kgB2t6aZW16FbUNYCPOmf9poDlQlIxfegWC4
9nTl1eFObH/ER5oVRlflnG+QGbTyUJeE6ZsdmuSgsfrHBe0EUx0KSmJvLkio30+SeJku4IkURGix
ev6knzrndqde8LW3xxyyHFx/Ga5PzncepClz4LToUQyOn1ay+rst7Wd+AAGfIeY9mwrobijHj/oI
MmnEPvxTSEIXsaJEculwAbgf0BLJC65kACKsP6TOveFMAV4GX9ICYArmumkqtsN2tKpY6OqvuGJN
gjwupdiJMlNuu+zq53Qwoi1pYfW8Aii3mWDVhf7YSXY5YfEXlf/+dBWUflnvypHhTpU3ufdBg9uC
ehhOwpMQS0HS5J48Jik8uo/7OjC/6QcpGFg88BAhzTQ0dfw89kaaCbj7Jkdggm3JWwAJqtGvUN45
8Kf8vBtZihLc+3z8bW0mwf8OxTN659wdf/ThPwbi6htHBqsJFvXX8eZKAppCWs8aY9cac9Ebagrb
mGf9oLHjbZiHcIZp8rG7IBeI/NXf4HO0FjrQ1aq2BvuY/tS8o+jbg37ujWDRXOnXjUioqxpya0Ky
9c5iI38y8McCB+Ugaitt/gpFFCTKHqsI5Jv3WYPQoI2WJrdwcC86V/OWHkMi/HH47dBDWAUEaphp
EBtgWXK9LRapd61Z1sl15d3GcrpDSH4bjRTyS2f5Y28LH/QvtN9xKqcm9UedzdY3JciHgxWSR9ab
/3iqse1dToavXm8XWouj4eFaCPse4rNZy3sOoDaC10jT2ntpIiWuJz+pObHdG/aLs9/uNkYEempI
bUOFq52yUkyd/wd3z6QENCIYUnpFDHkTH6S2zhQv/XJzhTYt1IOrqQfbWRemdIB+h8KHpWFmlZdU
E3QhJPYwo/GprGF0YY9eqSLCQ9ALXD1XS3nIFwqInBseHYsz+27ZKj1gCUcfC1y0Z+SOdtCXumzq
xQPfQR6o8UmSRZqYFgN+lVes7wYngnnyBVWgzPwwt96V8jluyqilFS4Glud7/zSv8B0cIjlxmF2h
yvnJvgZRmgXhn93L1+7XQHWWJYnsYyO1kZmiwNth0uktqvlR0b19YXQPZeYJ3my8+FYh6Cvjv/G6
qILAAkNVuLv37eCjTBthBPW7mtYPlTp7R0FG5bX1ZFl1qNReWPOr56ZU+WW/8+mhleaUhD1sgb4p
4EhZpwFm+cIZuj1QxRePcccY4lSoxOW3vZRuRLiyO9KICdnpW1VC8JGyHFNo6ejoNoqjxjC48nO+
osFz0CrCoy+GBEhi1h9sgvRjWzepsnaUeXsljDy12xLGfh+intAIoRSq+KdNiUUFj9M+iIqMjAgq
2I5nrCnfttIH+tO0oLta6Z3ZLzOitY9btA0rPqIQWUC53L1QcRd6bImgN+V/WAHm+WPf6REniJAO
G+25H/q/xD5Lg7VV21g8Nkd6RCVTxL9n12gHiLQ/3lkqZ1zu5wxa/238Xho+H75XZprfUpHdu5r1
BNeKEvIQtVPNJFmoj7Cd7v+J5Igqf3DJEnqlmQ+1XHXmBYDOKa22HelpV7jjwnnnQqPqKy9boWRp
EM346Hco3PzClD+ao1w2cjaBNgkqeL6Q3twsi884Z/csgeoIE/1NR/PkSTXoJDClxZv7ganVAe30
ttLPgWz0z0SECb8C072Z37h1tlJO8Mg5lpqj0SEKHRFKKAt5bo1XoAZqiLPzkBojiF8fG1yoNtvN
pVPAmI8kHpVQzZCjXqWDzRwcTEOO6JyZvCWOKvY4/hppuG+Z2kpi32woUSxcxpi84+jji7n2qwGB
Uvm6YXt87ucqCSAwJSYKqoqS2RCX4U8p2BiZA4JVdOy5806MSCXVO/cC2YLCh+0b8U2NHSCyg0I5
RUy7e7BOUR1rge6VhjgQbc1+lblK9+wj4aay1Xt0b2hBElyJF2qhu8Jj+9VPwKVTxbUMX2Fh8kUU
AXmai6q1VoTVCJWsnaejOaNYCX03Ulerw5qjEJGborfxwRUpAxRHqIS8119uR3VgjUwQkayQL861
6XouMrAzd8EQSVnOnWVycPIbQ6FHn9aIL0j5qjOsSR+5M9q7mMO1GSgfcQV6KD9KYQGjUPMvLJ2U
4AqDnNSvQ36mmCe7WG4RvGKVbfsESKXhF7ngPbFwBBSyOeecKr1c32fliGiO7stdr3UPeaHwEtot
Qgyr9EgLHzJLjOECTyb4A3uTz0NDziy9NsB0QhGuWj63qG64d/q2RQ5GuRwylsKjSc4z+yYKS3X7
kNJz2QhxKj+6ENFcAMHnzjua4buhpB/f7FpSGdm3F2QAyJtjSVPyS+jE7leFpoy2bvamRWpL0pQD
JaAflxJw5fqTsZi5Etokg+PO92/8spsT05oz0CM72FG+KWR8LogBmYFoS2v/CTo0ohakrJ91L0dJ
riMj8xo9C1oMRhbWlhGB4wkAR4Ex2SorGxyEulRcT23WVl+NTYOg8iyOckru/I4SfieayN4j6KTW
dUqb5YafMAOeosvYTFn9efZnSTaT1Fp2mrA/sxwTI/3bibCVfyajgUqhZyOI40ongzZOT0Qd+/yq
V+tr9v9M3hboAkJKzLNzjDMWYFvBj1PEvv7E+O2UJQU0A574uLFPLlkiLalejV/mdQLUOYr9N5/K
JU5srwX84lOeVla51V+7VS/mOGXC8PLkYt+FMR3ylhr32S59gIgg9+pu7/bJy3z8kuqd2r9XVJhB
iwo8oZLoYcz9abgYDP8ld/GXqW1Os/HwEZKP/GTuWKAUuI4nSfOby0RzPEbum5P9QwQjwqFv69Fu
X9EP3XICjPEXGdW3KFuWuaVCaVuSHPUXtC0asU/5bOz7LMOy0raIV+688QDQyQcWkw2DeQQJAjHA
nNzyEPeQIHE1pcrhcV30YN1nUkrELPfAmxtyjqDXigrkJVRq1Q+DKyekmiqMHkkogD4UAU+/ryEt
zTLl+DMv1prFRtrbaMqR4LsA0/zbB8+FSt7jm97AhxuvAr8y0K4oxbby5jzeyK/pds0FcxCANnV2
WWK0cpnVyBMefyRiP36dUJdJRWITAaRfgg4zPx4G6WZDJ+ZmeNyDi+mxxsp4wsscrxWmS+uxMFHA
9niwnF35ZAA+Yu3TgCG+55DaOxetRg+97+VpLfMOCm3ZHxoyytz2kSBNv+unvj55TL2sE/gyq3aj
oD+T1YyPB8Ll8R9t1kaubZ9Knz+WbCjLrKV3HybLMSIRIGEZUuYj93wEUvapDMqWPV1YQ3OdAn5H
cZnJwBaYv0T9dxD26zqhTJxl7fuc5Q32qrfFI7nkTlKAFMTcFP6U1TMOxN7jfuj+ec90z8s9L4CI
sGJhsLYYGwBntjirBG8R1E4RNo9b1TADP0B326+ueVaMOC8vmjc+KJHtuPgayJletbtkMq19VbMR
eMNfDpA0hqBVXxBygzPf1puzcq6yUHJLm9pySObNn11moAt+9tpyvchf/uhs/4iXybIaMZJW0cPL
aaD7ymSUtWFdnGZbO/IWQky4RFbKup0EdyYCsBmgKGalvSFuVo1cBibwvgW3WZQzSfHbWnJGQEbK
R0VLxhddtFPtNXpfjDdxq7bXlymgB3Xgmv3/nxEyyrgea+r/8/jPBzdvtGOmsM4wv/8bpxNdncpw
O5+419ErcO8OPZAqclQp5QtMxe4GDHB740k1GvFXxXpR6tG1lG0SWQ1RazUySta+7fQ8+MrFpzrb
6WjXD7YvmvPYLmZPgsX8dtd5FCuAqnMXenlbRyu+Hc0oi2OBRR20N5c7sH44lGBEEfl/eoipLEaN
rg9nFKisqCVQaBXy5F22rC4qeK07Fg8S0fWBSqL3L2vOEW0IC7m+W5Ow+QazhvaE8yeT/M622g0K
d0wJ8yqOWBuBA8KtdfNwEbEl7hyqlE5TDw0sCnCYa6bEEuP68AimwjqAIKud+iD5xhV7ea76RNRr
/eH42Nzc5YnVMugGzcBVyhY/YRJtlkRYWlnUhLsdzgVUDmvA33CJoaA4ZjrAdDBM87A8KNi8Q37X
VXrB5JN+Ekj4TwlvDdfEvm1R5AyXUvyH+orKoKfk0fDb9i+VieVrlW4T46JavVGBW1uM+GUIuY9F
QQjvBp2hp6UTTDEn+RSi0sDU0Yb5erUfthVS55jhgpaDjSyDZNADppb+Iou4SyK+Qp1AGor2iVMI
rf9W4rjHH2XkB7BG/cBBhAoBSrIAtP8PYeNOmYFPwRmVQSwOZYGNJ3Mjhzdv6vyd5QuhzsW4rzpo
0ZsI2/qciMjKACbuFCVkNFdK9HMU7cKli2DUiEpUjkIPjTbYZJIAVqj/rGBAZxFrDGU1X18ltdEG
ZYkCSfrqXSReNZmALrDbeEw91EZXSotCGvvU4Gbb5Z8PQGGu6gBKrR+HLUCwokjKW0tTj3P6KmpB
2zbgGEO2R6B6uuwG5TzolAaKhNSEO09xo09SUJPlmnpPIhz1cy3upclomkvxp6l6oVRVLgA2awW8
c4Ufy0nSHRmkgwag/ssSR6gcLKGm+RpN2CxyjavjZSbDkf7M889JJmEcHBzVpo9H6+8m7290Pn/O
UIpqlczaL1ucZ7rCGsnYpXmzZ07FXJaSV0bKNRM8M9cKDDlJEUlfAZY5YkJLh2qcieN9J20b1PYM
yiYCjkrukmInnDyzmGrzDeF9o6bdly5lcaZd1ZYTvlgTddBpBTD0GJKMSzjbH2l7ayIl6V9sqc+8
p0fFlDyiaZrc6nAiNaoVHQl51JY5gF/kwkAxJ8k5Cmb4ED7LcZgOyRuhSGn3PDNABliA90SatiWF
qTKhARqqGJ7PNSFbcD2gIxjQbC1Sm+PLA1ZmTQ1LP5TIRg1WbRsXTwjaJxFBznltCLGsu9+dou/S
Avw86Uc6hb/hoKeWPd7755Dm6YtiKZVx5fjnC9hKtjJkDBJCn/l5MCRHrld0hb2fK6+zQUQERlpm
zaIykZpyxCJQdw8uhSjwVpPRPaqRkFrfuELZyIFlWRlam1g20tUCOFDrzhKJJy9Jb6hqQZf9uASz
JBBWZYN6sVOMzK9GlFqp3G5ONpKd1urLTjsgARQ6Gx1qk/hj7RmHCoqm4bSK+O4q0X5SIC5uyzrH
Ire++pshjnIyUkoSfat/Sy5Nfj4uUj037XaUjmjW3duOQ3Cuo3H16mrhTjO8IKSqqsVv41RTQMIE
/9xZe8e2Py/YWpCBzWbqr0Q0ae6wKkTsbqWUYoMSIjRCCq45IJkwN97ysCKnWAlOTWMyvgYoHl7X
UGBTdZyQUwQOBIeQpKDJ/nwFnhShSJvuz0exBtbSg2+1KCvda7HMt0a0xejlvbqn6ldThVbRX94n
9zCHLTSXFCZnHQell3cLsVU30z+BTGxlzSlXS6gqa8Ag3JmqI5jFuzilWLOwCwdTe/Wepp1N/QlX
NtKg1aZlNzsmgCYeUCAXmuaarDlaNrW79FDJ7JbNXU7SHBdQyMLFKWmZ3d7zM5HE8z3LYXYx2wZ+
sbVSD9tPwi/E+G5jrLVU5ysFkzleZsixt3PyL05cCw9skMQbYT33X21u/3xKVR3JA9coQVtpPkeQ
saTfkCXzpyFJ4Tx/k3gqP1+vKaFCGRXQ/EbhVsJIMV9woVWCIgKeWxqo5jClgoFuvDd5ccxtVIE2
IF+qoHCEQfyxPlFl5/w0+oqisGh67H7sF7lERZ+ayrEa/0TvZinLDXy4BfQak1LnqlAwTvYKt1N3
Jd5po3j4JSRDd/BFKFUbdfWg+plhYj6LKXvF1jgu1XJ4drR9Jh0dDT5srYCdjZRlnqEEwPPTpK8S
jSiItGIBPCtr2Z9O+YL/vmOrlNGj/TgeuRx3AejhmL4APdE1iFKqR9XeBkqkFugOiOA72MVTX6Bb
g8pR7/qoKo/Dk1YnwIcQqmWRsjix49K5BcRVsXoARqocNKu6pSe1mzTG0Mgv4gWx4FiNlO61j5f/
TYEG3v4paD0jWmLY3wf5dE8YZgWmwJM9q2S7rqgTeG2DaEZDeSL/OYZXgb520/as8XJNh+jJzvwC
UzJAFOM8APWRO1xubCjZPU2JmXqZdyOuP3XnZppvFLotPytAGHU1NTl3Vi5U9T7uwJJGTZqh6Ot7
G894iz34DL3o0cn5tcvOGJH4gYwBg0o+NcCZJmG+1KnrrXdOIrHvzty6N58mZGTodQLxtl7g7b9i
PqoillaDSFA7avKSY0Qtk0IjpEbHW9+hzNM0Ht/WcDuNG6qXUkNTZld/En8QXkBdBmFnCZF5HJJ0
qSUKM3PsbYBndC6dJeMX/PnDaiBDVi5ubZm3DNzhK24T87uqF1bodG4asNhagz3NMdyf+aCxshax
wGpt0zQFNuW5ceMH68dH9xFnF7qk2D6xwxX5fyw+lTvLNCbI1tvuu5vxDX0OiYeImNPHrc22YgRD
BtlF/EydMpq2fd2Xn2XEpK7KuYQT79fns5vpw05wk5tTKRP0h+STJP0njN0CGsD4RZNK1+BRiQRm
Dq+a+0c0dpOR+cfJwMx9TywY5Ui35Oq9IcfkL/p7C/kQcAVWXWDY44mrHan7jQHwU6GpBeoEH1ra
AZ9JjFytivR2gAQqDS1pD6WrPPd/vKrMFhrHl2NK+MXETpPEABu+iuNZ4jmKp55cRWB5B97vBktt
rnDohi7r/OqUlSAZ4ALpYhUXyh6SUJsszNBMDSvj6rWPS2kSXZuwTnLUh4ZCQQJ5150xkvQyRU/+
Y3vrfZQ7wZPVRP12y15sASye5czgz6I4D6uFuoLcfz1Pby/8CBokAc0aHuJBmFCet12Gwr9N21AQ
KQyUAnoTPujEbmGMyh1AzbPcdiAGhw+O4m6lAXomb+ehFUa1FGv6RTZiM1lHWAKO6SHtDTfpsMaJ
G/5lhyw4JmCcn9pcrH5q7fYBv3/M+V2lx3KncWMrUuCEee6O2R5lShQ/trACCgByu78aM12Xfhox
em0g1fLL4Un17VuyjAycOJAj/J8bI/VUJYL16ftnp2fRBZqHLPJpP4ovfr+rCtxYugEFcq2ODQoL
Wy6lB5qE1YrPhG6GehUGM8QVHw9Nmxmb6oKdCfWaPN5bVka+jcPh/puWmV7+Jv/elzcsrXjkf/yE
nvwfobkw9uiYxxgZUDKPGKXTMedmd9rVCYpnoFaCqGl+z5exb4V4Pksjrl94BP1KOdOd46t/Bna7
g5ULCGnSkOfNPPdgL+wgZoAkKVSYVC62Ae7glt+kjHUyFoRPSy7oN2uaWTqGBKOla+jy6R1XSSP7
DAPH8wwwwH9c8GtxpEIq/uB/j6ME8HMKf4DquaccBHAqYkE9xrskpbPoe7TivlWeXt4AAvSc5R49
lvVbhWaJePbThVuJTvvpN/GSljLeDeGbRbx291FtHU3Jgl9KOV9dUt1GttSFzaliJ9LgeWo5i08Y
pOIv3qO72ymI6zyDNK/NiSnwK6rxU36/0Vc4DEJ1D6GQRNtBRt1c5OdCcWd5v24AqsGdrsEECKbE
1gFVGAZDX0gvyP/9xtQhQZh2KY4pi69iPvLbQewYKp5+3eBQv2CRzAjOxtX2aCZNm6vLMW2yhilg
1ns34E7C28Jbyhx17dsc4DMKn4T/Ig6Ry23GDZRS2QGTwziS/msbMKJyY0eCtKUOBWaIIlF0LVOr
kM65dGcA4EHPkefGJzDKkhtIRFB/hQsoN6/m7t1XrJpsb5zZEMWLRGUNB58Gjynrt8K6E72NunG+
orVwe8J0xWglO9YKtD571lgQgWBhJvrsFTdtVzR4e65hexKhTQEobmbq8IV2oqc5MYcPA0D3vfsq
sXa5SdwUroisxToqhuh8s/7YxgI8wsnwUL283IXt2cCwZyarpPMpqMwrf8Pu4ugJwfaiqX8gsROP
7FB0Ou+Qd0/EKx2E/Pz2Cuzgt22EXkAgNbguon6AJV9bBAvlvbfa+3OA0J5trTr26CjPkBGe6Uo7
h1Z2r/X2tpsiXN+ahVJSmyX+5auDrXj2kujY5QctP2KtpnlNIK81WlJXQ4iPHGOUsd3g+iDU6oq0
rGQTakSGw4AtoBo4/3ozw0rYEl6bPMmBjL0OTt9ZPEszNwIH04+12Kz8/oAai2mtKw0Bmu8DixDG
DOsJzYI0be2QyHf6yX3fP5Xvj6mtrHX0Hawlp1Ka10Q7uc7BahQAEaNI1fXq4y7CyKcDHsHL9LW+
Mh/nQ3xqpow25EdQk2vszso3017shydcz5bmUqe7pBmP0PkQY+YT3p6N4lpJtEpv5V4m3Avd8Hz2
6NhTvX9P0AcLo4cXuU9JLs5HK+hPBhA59JQYQygMPdnXbew1uL95UyAsZiuddWQYufggFHNt/nx8
tJDFlnDMPih1ic5uAsYCqXtZAom6HmZtLJ0D7oc6T6U9RA+nrxQuIjhwXES8H8OMedr3J0iiE3Uw
x+4kRsmkLZF6jenBfr+HKdjLxiPwVpR5W5audMgPi0Xx2LTYfbeAhd8UepcS5TjewQIlF/qX690o
csz0b4kIksLr3M7/+HgcA2zP1x65nIUM2VKTgKXZLnsey3+R5Zko0mYZz0HZmgU2j3tjcwnp5DX5
OuGUYp/sNuCMvcJ1dasojheT434pWOxQyfIdMDg7OXmgVtEXeIJnPj3tCf9/7pHWJeWlqiCPO+Hh
QPUC6k8vCDHmDM99Hybpiy7eQtpTrNTQ9dTcF6unhoWMdxymcBAT/jie3pN34OCavXmL7eaUSDqo
gwNtlLKzbM2cScSAg+xRI1hucSxaU8Xs8qYPzsm24xssLsYtz2eiofl5KIR0zzhjhsCFL9SBiucR
B4vr744pvFk7NZ/99WLdo8wEldT2tEy3FecpMHeLeEGUODMRegjsXV/jZ6LTEfFdHzsORlkOY5S8
YMrwkX0s/R4e7xCflZZnG0RljhONQ7IPmmPWFlt1r4fBZEiIK2DKdLNNqCY6PcMqWTjxuEljTCMM
bCxGVq9TqPqJfx0VUXZ2mxZhrD7ncx25T+8akB5CEH2UbPmph0TkdcqRURKCkTkHorwCOte7Sh6q
rN/jt2MWZMsKi4Q149fuHdiOpUD7j9qFJqQmzcz50SOxV1kEWXcRzN6eFoyOEArzPUGF816USkL/
ByJzXEC0LfvbTxQyu+EKmxkY+K+qtHRCcHSnodMmrBw6kk7Vw1A2gF0caJrwxHs8Jp6Ri7qHVqh0
HKeaeZjYstE/yrH4UfwaPvKU5tfTfC6YepIXpQADAUSdJn1wELvXlJ9zsxZIo1pW2bJR3XhQnBcQ
JG69oe8mY3wS/zOtWWuGbXM7NfCikA4YBlBmC/GrPw1GcH8bvK3JcJltKCOo+Rfaax3KB/Vwd2dU
rFIeFlljGssscRlEeVb/YkQSc9sfxBZl8nZRuQ0WZ4gAT28i/xc1PQb3vRijwVXe/OkWxXP8XsQK
uronkRC3wrG+M6M+aoARpZ8iivBAG5rWUf7CxrCJN1Qvov6QUpmtA+2K9azAc1JjFdk4pm+e7x8r
CRM9SCmyg5Xjqqdt6Uoa9g5FNk/EPi7EPCaVtsPFu8IHt5kjkRHfB+yYE//Vx/bYncA1Z+TjEg0b
awSG2FWO1QlPvU9o/YjDJkuPtpzL+AHW3CSCtc6h0RYtdUYUSQVWizwpH7qmjwnfNCfzeuOFt1Ay
467JVgCc+T3KY7y3hcAY7ExCWUu7VYy41Uu6YbDppOj+C9lrTHAhWLw3eopQArWECy2NkFjDNtq8
NVAHwe50SxFMPNXolfHJ7niAXEA42WDKRvzppcgn4pzPiBgZsUxtzNMNVrfYE5ALKCRYjcIeTN5E
z/0Z2lhtTbDZq5DOsVPf6gvb3MIjOfVMqsVuqGrQLLfkql5xE2f0R8AHmUn1a/wrWYAbxp+N/c4L
NrhxvcrsCZeDD/uRSUfHlei74r6bfDh/JinTShcEfws+6VvMhWto1gOkvUEoMfBrcJtOiabxAQaB
4udmW88/BpwkQ5yI2YZpBBVW1UW74pQIASrIARUFxVzB8e+bOzX18QHbz1RCYv41fwmaE5z/3I2l
zJEG9GuLkaaMl8gEPIX1iVV/0gNtv5nPlHXQQXIFaotJQWs2x1ynvVK0sK/GpPhUb4vw4qXjmIGV
x99EgngtKY+RtoW8w6HB4IW0lrbopD9rojTTldWHaiLQG2zdkGnWN9iBnajksEgdECPkhJ1Cmqdu
nvds0/SGTRfSdFZFCzkGMgHJZnZzCbR98OMGl3OvMPArri2bsWCAUYhseEfA6URaTf3WNDRAgJPy
srxaX5W1uv5LjGya9FO452Ek3GSZOQddYyGW5/RV9idK3U68BOerVbQRm1JKDNxlwUm7nx6MH+or
kfHH9fVQQdy/wk/NWTJmGTBI9gqdAQMIieZS/IITznXS7/tnpXQTLX+W5fB/XVCehfYQe//XkvNq
F+p/lQNrvxJJkPOyHPCNjT5zVhQXCfoNYoaSCtg4cw+Oj61AGWIAJZoPGXL8N2INcJDi6dSH+Tw/
9U2lsoYW4amSZnfb2SbHrBCA06jrVWG7QPdgvC37AlvevyErAcHdnqJI/PMni+gJ0KDiuIBtuJgN
f1qgDzqqoum1D9tc3NT/bgth7rYDTVR3wW2iAAZycuVKsie6naCJquP9Wr/y/l4RH3+KjqpZpIXT
rWcxDsGMJ532vbNZ/82std+v56u9wkFE6jxySpcs2cpxb2qcFeOFbkgktVhyM91HI5VL9SXgrKNw
Dvlls3iR6n4nE8suLdSxI3izOndPPGM3DDyuhxG+rs6OhRnZGmj3fka+kZLv6ren5D4MDVCGvDfq
w6CapkvmY2IHUltODUVucDZs4oRwq66e+YEs6GLES7J7JjPdYncpPZsBF/gLSyDGOx9pi/GonVME
koDZe3/h0HkKxGIrPDFdQWeEGmEJtGSneCURuqwxhiVvUlhzLcUQZRudzEd+BfFiDdMdmHV6ZK3U
PbqtMr0xXHCSJbP4KIsMdL9DY49+585Wo6ibEaiehhyVm0XvwkqC02TxmXkiOL/SUOsuCSccGwd1
KfKyKtwh5FPEbr87maZKvXm1vtRVFBYGw3Q/Hn4ptP+yidWPyLNxM/638IT5KmjqIsu4F2l/zo1q
dji0QnZe9qSPnQNxhxo55rYfjyGKrSvC3HvCxRI+FWaR3/t5WRHflDQy8dxrb5T1o/EKkUSWw5Y7
2NpT5OwG65yF2YR2nYXNTCeNvyyLS/6sw2BZqB9qQiPTP+dDqgzZmhOMiONw/fYmRnexwRBGb+/K
JksfXnjIk7UzvgrWlfQ1GthtOADahWydQUuhGNk5xu7zGyyzdP90B12P14V2G31vzEWu35le+UW2
fZYo/xMlIWWTgV+hDLSDR5+VyM6lP6KwEknoWUr8/uS4qn10yZdjSCip5vPRoVpP54EUMJR78j5+
ZvgKb+cNOrljrsFiOM0R6Ypa/99y/HluUxX79pBe+TGkp1BABc2fkFMK/55eF7gyDTc4pC6s4RdR
s4/tqpXMcqkQer8ENpuGS/I3hbEV2WbMwWgRfeUEBA5W3uTlKMIbwGnsEcfMY8TipNesjQkusBaB
/ndr7cUnNa4zvOeg84RTXrtKnD1Aif0IsV0T4klLyFFD26tWwjaQEhzMYG/4T3tsViLDtXYUydXK
OrWXCcWY681xF6fZfMvE+xR874OqkwaLnVMConwGMnLATW57J53KPMRquRtjMFbJr+79bvAin8TB
lddIy0dsXUMYBSH6Zwz6sa1HubF8nWc+AbdI/Tto2QmS4eCM9k0LaZ75ZAxB8BEZuRiSeeuICuJn
ei3HMlJcqdsyrPwu7nu+sWKYg0M/McNeGhjuq02oMOI89taiCgQOFSo9xgsu3zmQZDpH/i6Vbu6/
R84yHTg5Qe0dtoLBAQ+jJZHQshsoHepQxlAwoMaSEIl86kmjl7QR7kWRJKjRq55msp8pXqwKdeGr
RAzG2vS5wuCnMa77gHYNHl7fX0RgGEoHD+x+nURurGYFiEuKZJHQLY94GRuQi7xkzNFBXPExj00K
wzsqRze5lYsoX6Ph8J9/wOnxILt4NZj17b1LYiIyw1AAt2P6RDkuEJbFGnZVkUqiXW1NFz0yIb4F
b8Tea7bBZi8PN7zkMiWPvawHSuHlmy9CBNfsKHJ641owTP539GGg18XBIf2ySVAEbkVbJwZxjb6m
NYrrdR7/BwVTc5zPgrgnbw+KLjKi39zQGIH4iPFNwU46Sphcpsa1u2OzmNHYIXQ51wvnUtSj7/wp
ecTUEBrls3HW0NdvGv4nwXpdWQODOBLdvLkAo7IDuQ5ofdYc7fKhF3US9K5IHPNierU6enq8nRN8
TOiSt+/K6kfh2h2xOQjKi8GEk7UMYYaCukXvlywM0Z0l7ZTEXpnfAlvcDiAXG6aQ6M4vC5xIov3e
d7LRfXTj7HegqsD0vOH5u+KBzJPov838J6OmhQIqBEyVqWknenD788UNV+jFrheEwdcXDV/iisOI
G13x3X9kOqIx6szomApn3SbEKY3F2FR7UqYkD/3f4fL95Wr4DxnhAcES/s6No4Kb8dqFGwWsGze9
V5QM/GmdHlt24CzU6/ubeNpCk9oQLaCtYX8oN4ESFxhalYJ+xsdj3tFHYmGWshCenMdVkxEoqVz1
iGkvPMHvlQRzD4sMAEN8Ptabg/ZgWJ+F8b9Sigy2GJM6PT1ctmE0fGvyY6HK1NQSPBIvep1jFV8/
fkLQ7BI6pBWftKWVUmkKyuO1TOcaov/63NZziScx2sn6oEYcJIDoFMZyBUfpeVETb6jr1dPt0AyG
PzX92hDF3uAnTmAwvrCwoOadrof0UJYcl7KNIXdeaBN0QJyPdWuIkRc8rSZ0BLiUkkBDPekSUd1b
+8xjlLHOSLun1XAJiHVN7LTkgCdU9Vlcs8/RKekWHWqHeaZRod8gmgK++9ma+ujomJsGBfSQkbvp
HYtC1s/N5/LnmkLGCKeSsYcgL5w6ozvVqSMJRChPrDp2qUKkQzTrzZ72IoqrioHRfL9s3xbNuTSd
AuVaIu9Qg6M8ETajWHqjDD5xe1qKvfmyvnwe6PugnZTz8WWCztzRLj3rQcU7AS6tDKliLGfJDqDg
luR7mFwLb8i+3UjFnRzVAu47kQVpn9uuvNUd6tbqM+umsxs2qZ49deoxOsa/i7W1Aai4/fWjDxyE
t0X97i4/8QgtMVMwr3cD9ZHHnhe4m4SLvJrtDQWfCXJ6SmCoPGKiXxllfsPhN5xHjkL6HZIeRP7g
arVQhSUjnvzimbKDloI2MDB1AHbwcI8/pn7C3KEhtXnnbwI/0HK3WTrxymT3ege+ipM8svfYobki
5LDoMRFfnk8imcwgV7HV0uytvKLa6HIhHkLRm1hfzDCyaWLgcEkbkaW9UmeG698yLW7ykPGtLn6B
Lvp49AH5n9/MsQf+0nlDpzgOXvEQvUvXckp+xl2JRT+rmy8Cwuo1ax+mSSlC8LLgK5XRic7TCpBv
n7QE4bBSkfiGUKBpodXjhhLxqBo8xsPhqYtkxNT7ZOOH1gsHqzeMfMrUzN84sE2LG0iyxt9EImI8
kLy710w5loX03p2+8u5aU3N7hjyakrmoJMoO12SVvw2UgjBse4SBd4/N0EWD+bBmG5wnVZ8rFhHj
A2r9GOg1cN6wz6ieTFQMUWok54c53MbhhObb/VC+XyMwlYj1JxlSIGiB7VMJCPtSMR5I2LQIwObM
h4lLj9mGKdJjDU54DPr79ZKygcmyFQccsRppGFFh0XWaygqgww8zvGmWJ4nB3Nn6I5JWP5aEOZSh
FiC0VI9VxCbETfFFUUrDIOO5Qd0LYsmenawaYlwNhKBHTTZNa6HqjINgkm9h1bMT7fv4fFnBzx/p
osNSLPkaF7Eb37TByLSebZ2wVycV1PiZ/KihgPocKzRo2M+Glkp+3FoD4N0Wdnvx9dgL8RMKXz85
MIUUswoYSrIlug6U+fsixEKtP7Z5vfvpCdbXWSvVFUra3Af0ORZ+MqzSHohxLseTZjMIIN93o/71
ErFSr51TfeXcQmb+hr0ZyfCjvU4byFLdNfSuqvnWOp4t96Xnucc/3O/ZcrjaSrjxFBcWjOyk+DMx
0TY6wbLQta2HQLZufhXZANMT3H/SIUtXcCKWkn9JBHaBTFuYMadqF3Z/EqTSsVMAw6DlOg2jDiXa
lveaiUSjXnrNnQWBvhTYfmOc/sJf5jFus6TtTbugbvKXW9rdJPQuPtjpSPMTszRst9CoLhGATlF0
5rET+WZZW9UII+Bx1MLoGS7XSPWGc5JMYwPHpTxuHBDIhubkZ11QJs6V7ZkeQQSyBPRA+nFGLBqI
NVIs41enqWe4wQsooPycAoScy8SRd+FXirmfsrkOtFc72K67uau+Yh1ht7DZuxpmiR5Pkg5MKDQj
/JQ36CNzF0L1vN03XvB6rvpMDMgBfijor2gw8bZRzrpfTqPhFHqJp6/BNtGCp/hFXya3EmNrOkWP
MZOfvjGSK8kp2/MIw316m6BJ3V4BO5hvPWjWiofBEq4OqOVH0eG5YUSvhL6RwAS3eROxEEp+beEO
9tCd4vHtQ2O9shWJRhDS+HlrVKM5iagjRIBv2kClrhfJNFVXPlU8qj+k8vmK8jlxLd3P+Yqq7H33
SqVQ7OY9W9DFginqtIPMeyXlj9Jw8ovL2+7ULA7KoXZWruq3rY6w/yIk/Mc7kmmmD2YnUV0ltfBN
SV6sKgmLbiNV1S9TKnSLFBh/FjcHOtw7SmfdG2YWyGhQkzCy1FevVY6XpEvX2AIxeg32OQkvBPWm
ynQI1nf83vHAh8Gp+fhu8VNsDIiM+7lKcTMlYSLhxUNFXDrfxzPm/iYdIw1INw0JJHuzDRMB3nwo
plNKlytHzS9sf4Vg0g3lb60xxMEPAXLEg//79mglsvvH+0rx/L55g3s7yvLHYPvPclJqauYTlyAH
5REeMd6BjznM+Fu5Xa5Qvy4b/qzG3J4VMygcFk2gnF5JycujbjbXMRm+xIPdmBsVmF7uSxkMerp8
RwFesYkE86EAdLvuGYjdgbOob+lgyHO3tA86nGtxMtqp1tudjgOfKj6N49uYDrr7pnSTJKsv6IeX
vCw5k1RmedVqoHJhfnxViw5fmPBAWUpqlQIQ7e5oV7lyxr66nnao8Dq3BAqtZgyc5KyG7+aGhe92
aHXVXjS5ZNHTF/vIbmu5uZjJcXVOI3kjROV41mOrU98wTEE4raa3/wamHTNlZveBmUp5aayOEm3x
ERaNtFhkp6G+YThbe34qWyu9ek8sy8ZL4a9H8HrCbayceG4dwsfnaFK+hesudTKtf4EAM2/dPy5h
KE+3ekaDfrRw6J5H9GQWm3utWsbJkeleJ4iNzOGyZhCSEbf2BPTt6+p0MHO0aRNqW3+iPzj0KgV7
4P4ALs7YAFtDdE17CpfcZ48jQGwLOskwHbhXsjk8g4QcB2CA4aF2re/fW3ezR/CDLpWjytAYkpBa
+W2cpHTiZXwk8vGUOaZITyNnBjZ/DoU409qJgtNVrPqvlJ1a3lniWYWzoCFVHgL8cU+gBlvLIh2n
/i4WJXGfcErt+bGgRC6iut5Qpaprk0EDEjhyR96FSNGR/YXKBi42a8euWOOT+PXAWdt/vtvDQt0e
wo2Vthk0TFVuUT4s6vg0UkDqCb9nUSObb8NkXqmV9HYlhMq00rN2B5Ghs97SqhrrajBQZ2APQpOY
m9u0mR0+ADHMiicXek5F5tTHEqt85nEyY6kqZYyxBWOxygPPDkSu0ts8YkNSgoUAOocGwMZ1YJxu
JwupY3HZcrsPN/y01ZHdm7Vibi3NooJJTDrOi9LGDSkyLClBEdPReqBOw87252Kaj8gLA2nRzEBe
fZcxGBUMqSOrcT9pt5xH4wl/YeBwvCFOVEvH1GUh1VExLkmofdkzhgn+nvySzYbPv168qazsHX0E
btEUl0hKe75UagPj2yq5d0Xv7uiQDS548V7wY0HtIIRvf2FXlAiG7YwifKSehYsWDIwD/VM7W0A2
MnEPli/xUWsag6UtT+tOwyAqopCfuOnkdfSk4gwgZhbddA7I4wTzvw4ADDg+3Cv+S99G3KC2pqYu
ZVTX1Y7BowDWoNn9EjdFZkpWcCA7izvymMarR/UL1rqZawGWfEbYtbLWmvrSAzqsZ4OumoRFylOl
QU9ixqNJUe0q7p/yJYZ1/WfehpPGRRJHpzQmR0nUOE+1Xam3VWCtDO2jhQMEo4I6jRf9EJE7AJj6
ScAboUWurDEkdxfeia6e12dzcTtyU1UXT4cxlkJ/q50Ba4963j63ezobsXHgCW7c8O4BBwYWbmN2
WZH+uYnfjf0j4FMRe12tcrOL4MkoZNEaQSDvbuhIoxv12h5Uc6l9DJgq1MtZNpebWubAlzBXI3M5
R2ipASfjPx4y31vh0Rp0XxlSSOil3FuppQQGg3yci8ZA6kPvC7QiE39DkifUaLS+S8qCQ29zcyit
i58n0/JcVhFEHLa1qhKotKm81OnxKwQovKgot/dvGaQVvlOCsW/9HTKlSSrBzJYHJtiJd0w1wLt7
+CosV6tXU3v6y08UJWl/UoRGIos6Cts8CHRdOucUDAWFS4+MLspRtJIq/jI4S7wgEgOsc+NSNZW9
6C8H5NGmO/PiAtuHA03vqpw1/qEXnk0XfWFMoKhoziPrkyf4zcMy2Ipk25gKoYDgd0SDDCOd6hYM
mCcXkhz+kOf9J4TkgP5v1wQBmPsPbC9QbP7i23ERXbH/k5JVB2A3rrvO3JeeyX90GgJgiE+byxSe
qyP7CXj4zPEHmGL0OwpgkcPqe5QNzc5EHwcT67WT0E52jHD5nA7eZOtqly65xIseB60S71SeFPL3
93kb1M74rDMVjUfsr7tjQGBTwBQCjfajr7Ep9HxgVdCqGyZI+DWhmVjd6tVnyN3E92YyWJh1Os6I
KnjBQO0ZhgCnWKdOJrNv16NZubM6rAojnlAKxLSuWsaC5LeFJLWxmlQfLLZV2uie1XLJLOEGWrq9
4g/Cb6tcCxyv83PoxdogLk3njfnX4DCjmKNNIPoBOQ2NzV4fpyGjg7fcxvDPngYKK0aIKcd4UPZh
5qyvvnDbtjHW92w0Vrbft35iv4s6KG29e/Yvhz1IyG5Mha4IfpriB/lwaAjd8bolspfoB8BQ8BNE
eNXUmuXAxC3TCd44NqbwAwA/DI7b1iP4NoXTnjY/iQaiqxM7BHPQloVx/wK2tdaCOEXUfygbcI5s
OOaqXfCyLXgWmu+eEnYU/0cOxMVN396k/lrUZD88rGrLkRB/Uvn/F7KS68ub2T4fjN2xmHqNa1wy
KgR3LzcZ5767b9mN8g4sFfJRBCov6OcjQC3CVNJU/S9sxy2W2wrvYb+UILgd5E6hQFDRTx9BusBU
GHMyaWezm/3M+cutN10u7YVcjDffUgLHHClxz5CPkfy6bbmBFRg9SUlEbWAusik/yzEDCNHGO5Fl
ZLnM8RM1I4bCMhqZ6eVgw5k7unuN18DniPBCcavDLtnHbAJjV1Dk/R/rz2KWdGr4grN0IAH5I73x
HAf3F6zrX7ZSbD2UpjouuVdnuTUtM4lrTx46Ia0vwmgl/aSRI52B1NbIY8QIx8leXkhjtBesytIQ
OA5Pb58w1SAUW4EowQDluJ7HMyt/ST3G6mZc2vnTYNug1RT6cajv6GHUtAgTuaEVMt3wgh0r/3s1
aLQEn3M07lq064khAqJPNSIaFtgl2Bg5jQs6ahBAUdR+KnUKTfDXDgcgEowZ7BYLM4QHnTu7OBAG
GMP9ygQpQgldbYwaCy71LkFUdjrongEENtuTsh21k1Ul6wiYH14DWMhLXxQ8IbHQfb6cWfVZromb
g0nrJxqwHT7Tdla6PjAlSRoII4KQ9MDCOoaisC5iIR1mBymdQnmRtHzENVqkOP76oMaaHnXMlVVh
GpTDTeQimnf2LMWqHNcdi36Y9kbLZVDkV4O3pn56/v8I7YxhdDb6MvwW3EpIUkbthPC/HF3PXk9I
Oa7Il05mVrDOO3oCm/yB3eMk6DEmU1hZk+1Z2v+cm9o8s71rgkjY+dLh0+BbsQkuZrctaXgKSHIU
osvxoQufKZkwJ7BrarVBYRqm8qpgZ56CLGVV3sHO5q+pbR1V8ek2tX8dk38vOjpPwRf9EDfZPCYQ
JNEDLcGICGvvHxFnX48Z/B0oy+eLH0nR3BIA0VMRUpD6OeTFup5ALsU/N46OmHC9aWXMx4ppKMGF
TpPLdQVAUWZJf7yAsMlj9+fi7S2ADiUJ7EQIc9StX/b9RzHTdlRjGlKQ312sAF/1SjuRACVJcyvH
9rUlqNNr/MugSse22wMcQ7VF20hvROBTi8zV1O/1UNMHPOLxPx3mEzfOmXyjiAGcz7HNybCc4LJ3
dKrHNvay6dNFVP3AFsbmyaBcyynfM1UPtW/x+n3vdNb1ybx/Dr1AwFT7xj6dF7qfqGeQWtR2m60M
dN7Enfm3esJnRhHRUTmhFfQ6sWTcZ5mNjYlsEN/MbxupZgvbeW2ksPZ61umJFBemOc/xP9l3wfWa
Dv8bx9G89ykkShRu8S6H6jqZ0aBToXTwrt6EyiBnuHP6z+Gdc+Buf5ZXWLCrKFPN4wj8xiq/gw2L
eTSz4qrNw4kLOS2Aua6/U+Ft7nOOjeCw+eGXG9/XMa8MRin1a37Tc7DTTuRV8HALdw7NQdRtXhAv
0tyfqgad5lUeSgukKWZwQen5bXYvmUOM0vTTI8PhA7pxbKSENFjEqnyPnA9FOQWEMyzcOJr+dDg8
BpA2XCScR7AcbRpicE6bYz2Xr26fDEGr5H7XQM6X3kE/vaH0/ej8P5gOSS70OMHyI3gt95ghx2bu
PLFmPZPpYanUAF9jSUEeQne9TpMZ2vPgWw7m+fBY0QCZerjPtmRaVBdnSpgs7xiM/PRGVsw1bOCP
IvKhdgg1diZp3SCIcf6ifGpqVdyUtWSdNzD2piOUA+vKkrnK3b6mz46AOPPXAn7O1ryWgRN6cf8u
hsOt+JfVHIAunBxSHYCoAiTw0Tn9U9KQpSXMpzbTmwjwvFef1sAw2titCKXCeK7TALPMr3A4brpO
Zeuxnl8X4grkoesF3m9VBcPyYranLbpgcJJ4MrsMShjSdiHSW3wNFArxtxLV9doD/CGGoRmjzNQ6
EhAjHK26hsU3IERUOXWLw5u5nMW+2FrvhCeQZbHWv2YFR9eyU3URs8Y+0LCeXxd06ZQabEET6UXE
E0SeBQoNZb2UWTwn5bo1fQZBrbsDwXmjiWQFAucm+7vvesyyOWty+zgzZ3I3su+Tgz+Hk8gM0B0Q
5wv6okddA5JMdnZTyI8ypIQBLXN0tL1SMyxNWO9m3Tp1VAtXV6sPJ5A2sIhJEA+nnJzf08b6gUoO
ZsRMQO9qS/T5brXs+RrFFKnvCbOyRxAIOd5iwIfjex+oy/If+bVdlTLb9CDkPJIrvzr9yAaXk42c
Wt3PYpuasK02F8yjNu5QuPJ7M119Sb7hgLqfRn3yFJ0YlMJeQn102+EEMeufYoj3by9m4/xANmDU
axEu+dj++J0Jq9/a72up+AFBrMDJEriRqU9G+eaJwzORoPd/js5HgAKAe7/STrem4ewXDIdcptc/
eJNs2RLwNnooGcJPAWOB79VQsHzdVJjEwW7Rm0ANiLNCpS8RDvnDepBodj/AGg5cat7BLWYnTHSr
E5qkjZdxnqXyPnjQpgR0+FefymjmekxWD60HgEntob9UX1+7EWbbGegfNySFtIgCBUlJf3+Exbwb
Fkj/+N337vO6jeEPXY0vVIGVpkLA/MwJP0YtT8Q/RxXV3uxzJItFXqR83KBxhs+jWw5VSbjZzCht
wXRzCvi/hVmzo8tExolVIIiNtYJuJ+X50rKhcglFLM82DfpoP+p6p03QORTfXvfZkz6uLYF8HvEo
vm17lFziDHAh724jZOy2MG5BMQyG5ei0K2mO3rCfO8omFS1PWUVIyFmKFyuEwoI4YuzPGA5xLFI8
UmcYdNLWpK3wGIHmTJffrtYqylQMA2qcahNVZrcDbr4atxRMeBUWtOJPEP6dbk/ZcM++Hq/oQ26Q
3wK3MWvkh1vpWiiT0xbQKOaZUCAMhHeDaDZQvTE65BPHTc81hZlymwcXTuVZkyZS+4uRtTMGfmDd
JiFL2RlJF1Z+Xkp6ukpvYPMgI+VRZDVmcxasVFE/9tMnchtnI29JHmyALkPydYnAMNyvITUzrpHu
356jYs6IMnbwdHGhzStp32zbpJb1KD4HEglzFfVhFTW8CzD4q7h56qQNStRW8iVoPsyMlCp2OkOH
HIwByHDCQZ/5B5TwgaIJVtk3dX7x/ZUFK1+S6wvN/fpZmGCBSDMztK3Jw/YvdqE96N9A+Ur7F4SA
olV38xrkTKGHeKhEZ26kW9u4ePphAeV/+2jF3afgiGThtsSlYZxjpPPNQsRr2mo2pDkEGlQbSExm
PIgKCqrYqD5bWNYCSfotSlY+Yrh/D/bPksTzc8LcRb1WB92hf9qWp9+H+OHEeU7sPZjtZlfsuzO3
dLAPCz3vqPIm311PpogqALPGuhqCwu9VF0HvZWtdJtJ5LsIiMDnQyg7LdHwDeVCw78WnPmOjaWFi
3ryds6cT8MWPldSadTR3Or7ePycI6Oa6yPR7a1uvu9cWY9qphLfQ9k/AJOTagAy4Kpok1XqTbYWh
n/arBD5nnxhJYnyUlgAeirkRkEM1UdlWOuQgD3rkZijMCV/09k4M/eHajxAb5DrCkE/YXMaqIJOR
hu1hQTePcahczeNkk91En7BHXT6PPQlqxsAG36tzAYCNbvxVLLPP1inH5d7cGyEpW63J9ImlLtRU
efsmsGvXWD3bvk0DtmP/qtKYBt/2zOaaCfJ1SuyMxQicEgwMg5mXoLN9ezv1zNR5x50SsxpVRN45
0QjkXWCzlwQ6o3jjZMIuCk6qXFzChpZJ9TtOyuTtX0R3CfQf+jAMDUslDrCnWvQF8uRF74REOv3M
j3i5HJHmnwGpHuizRHLguHcPYdbPebUK318OyTSV4E5O/B3qT5h7cXIiTQbZBiQAymiHXgrxCoxt
/S6A14jal9Xn1U9+dbtZlaWTWWgAhXtwlF1rTHSDYOhQqZMIMZVwuMh7DivCVyDULGNeAf4qiLm6
BhFVN2lgpLR753tSO5az5Rl/+8urypZIHMy7SXqllRYkuPwVxckMOIv4NK8AcBhVZNVgKeJv7KyM
RDjcMjGk4TjAkhSdseYG5Jn1b4NOajQpvKykCfSrlGNnIQ3Fgh/rikldLwSDn84QI35cxsXIec18
eKjn5QllZBIlEb6xgXp7Nf26IjC9dCQXFbdF1Ke9Y/7ubXKZL+xGv684ai5FEdkDGwI0gCuIubB5
4HxkIEegOJV4t5aoiNaPUu9+hDPQ0UbCBPiTtJ0yY+aNmfGf72z9zrYTaR9i00ME5eDmZpHt/Bs/
J26/b97nOPfVEiy8myzdPUXvH3VC5u5W6YmtcbdNvgASFPSM4RtmDTG/JCp6pXmoJepkXpR2cyHh
Y+NINOqIDl4OiaOCGt2zqZheK7TrRzdDx+aNphKM6QfqUOTqtSUqdAygfzPwHV1oZ/IKy0caUoYR
RcofM5Y6jjUpmnsszCmgIcE/r3awJGX50FkSYuG673EEvSucgm/8bAwjOkT828slOjGYqezt5Jo+
+Zn54aqnCFpMQ1LRlIaHsA8HABP9sQ+DQtIczsyWc+OOQr40OgSutsixq6+fP8W8pALklFm3AfW9
tlSUZdxCmwz/IsC+isO9LkUzuOMMb9639pke8nB9jQVmGDtWBKCcGrrcsOw50dUDNqvUNhh4supN
nMH5KbqCWnaQmH1FK89zV94sIB3E24rO9dscfu17KsQbvp1CBcy/RmBYBO6Y17jkwOQB9LFzQs9Y
rPxcZXDHl32Jpza9ACzWjxiOWJWGuPW19VBSb7wNGPYkIN3+gB9dOqgAUou1e9r38Dver6Umsrk0
YNLCr4+X8kM+fBrvqODppOrrMB9Vle4TS3HP/wM7PEtM1sPyjeLH4cm2b4WOeVevoVBUZnHWwL/i
vxlLp1i0Hru7EWL2PPRrbQb36y81+YOr2Z8cpE6p1SRKP8/ABdE4AX5I+iFbLsHpfcvPgyRJERGR
XGf3NEBUgCq3zhqZ5xsLyroa9lYE9TvdcVSGwBCj6db1xMQ8yUoeklupiPzDV1wCQjeS10iVrPsS
43tM7t4by+ZucQtnPj3YNR4qEvis+8drTA8sMglPRDTmpDBFTnzfM6bZonQfqQSIlNiKbIpu2Q/r
g2HhHvFecSzbxQVkqeyrM7XzHAf8g5cXPPou2qZZie1PpChnLcstup2UkAyoXk9RL1/NGHgZ0+yb
ZME2NLVGcrs4ed/qeyYt9zUuxFFngj1tvoW1jvJzS28RZaYxRsf7ewFaigk1Daq9ZmK4efICLt4b
CS/h5YBRsRjSBaOb06fdQ93LwBrlEe281Z2+OOlTxIs/BeJwCZabF62JN6W+eYJHtFC4sTtb+YuW
KYgFraVEj6r4ym2GpWhKDVF8M32bDqPbMBDtC/+7unyZEdCivVPTMqZZeOPGR1n+2JeLnzW6YuTR
W2AfmXnU2EksRFaXw/MCeaYTaF/kFrW4ak3VK1CmJD59llGGLqdDwJs1bT5Sb98KWHlEZOqivA/q
CmvhocD3N5E3Iwz8spnB9WXi3UI3BT/byaWMo/64N35XVqoeejt3dritWQb5ppRzMG249Jj0nWV1
4GfpSnHSAbmZkwziCX6F+yMPZGH3W+WrLwTwzda7HAmJ/YrnjrTimjluKBORSItZuAdLf5+pOFbv
ShWl0fKO/TxwGTOzKMiy0YQyS2heNV25PbTCa6HBT7YQNOrA6WILNesBvXTNf132/XBb8wexa7ac
nAcifD+d+7+bft++nvuCZO1elv8nujbJ8Ka3Pk7IhbxCcK2CkG9NB4g7kvSVYdqOPnqT79YpzpFp
txjHcM+upkLQOhkgxKLGFSSptcwQ3B7kDsxPOyTNe4/St1cirSyOOK91mOKSCUpi2hp4odTRccNi
CqIcFr7JRj8xdL8rL6Aujle5RBgic/1r5TLmeNUJ3UGMXNMqxE51W7wD4ZTjxp89PRZABR4p/M3b
gE6ZrFIYC+oDqQNJRBZpr2ee30/ifBBBuLWj0cEbpk979ifiovrw+ls+siRSZrZETrUAJfY+rowH
UZ/VbD3FHGsj9xof6uyc00psI27Ftm7QMIB27nIMx5zDroepCRpJTlLph0f+ht6DLx03ZM66Dfkl
NxoTQgC+HqcIXgvGIMLpnS2NseScOxd/N5iTozmI1yVSo4znkknxXTVhr+jbHoMBt1x6ap6Y6tyN
fKPADJhWWrS9qrV2PlI68mStxyoubwVOcdIEbxUqpiaVG4DTKb3Alpz1VFSmbSaV/PimETYOABEO
Qb8SyUrLOCn7TsumdOZgFwoIKfXRTo692IbJO+AZGVmXDl11UIK0LWbug2kLwKwBlAXaEBi04v+9
RfPl+Sw6uCkGOPz6aYACDc8q1IpRQuw8aeqCZGQCs3m4wWb3jPg7BKw9zQGv+Z5EEh1SdBD/pgEX
KZwx9sl/8laV+ZabBWI33Twkt14S8ShPUBz+BpVVP0kyza3nstqrYqPsEXzz5b9inLGAYtEoh9aK
R+DLh8ViwkLSUYyoJuPGfw4LaZy1CwCZtzWZeeudQHxF22AIV1RiZujQbOVQl5GCG0UbPT1uauZ7
Jr7u+uwA1xSVWn81AfR8PEFCCDrQHe0aeGD+n0FEm9PAQBUMOm+uQaaR6N7R0zF7dl7fWxvcMIpB
ZXILdWMkL46X3QvzHIPesMoAPK3MbQ+TCnap5ULnAYWpUg1SRHn1BYR9L9tg/6nkP7z0UNKLK+QN
x5dtIJBdLoI3KDYeBzcbBPb/e90sPh8qa2FnSq3XcNWH4HzxMHw/EK+fDVSOq5IkMrA17VLyuKkD
33DbW//QL3Kp3GZ8b9Pl0YDY7daYn2RDiHiFz7sSKFmO3O+55+r5E4Uh+by5t8YQK64fwvVTkwZO
JpLvPNjBVtFkcaNclDSxbQ0gnMenDqUGZAY372eFiR3GUwnDJhjrNi7xjFQns/6H711kZeYXVilQ
v43AcgQVV80w2xo3TGXNrDQHDRajPIc50U3YTOIXCA170JEMXZFjQrzYNpHTm8qbNhScFXPg2DR3
ynq6X5lCcs4ntbtOqApvQikMUtMwDeLtwqNYxUe9bD8crDElx53ILHCPKSVY2pvS09dw5D1mO972
mwh+ivXCrrp2xS93nBOc7bLaeLYWFTQBB6FLHeh+bz3PFez3DsH3GTTFB4oJJVbjsgUeADGQ8/Dp
rllYYmFKiOhJ8DCsI4GQpnVRD1WL8E2Vwqb+q8VQ3UMU1fu2rlePf4DTMLIUm8ANwDShbVcP05Am
OiFtDwgNzvqH4ZctM/uelKk/yPbdsd/8PWOsyOOH+L88wNz6sJ677GQJKTFPHyJ+AFpTorMxnajh
25F/St4IvPeW019oIp2pAjCQS5H26l/TvYf00XM2ujfVJoHhwpECHAIf8jx8/ywBImIfyYPtGfLE
XOyd8V8l86903Z8y2qe5jfhdlc9vwceOs1c8ERRYCl+/u8xroZ9REuDKJ92RhP9dD6xk8bec7Bb/
EeQgx3OdJAqQM3yAgEoTnkOEW8sTPJrqrN/kHU4ru8altdry1Pe3zmNoRDJyg/d0rI+CfGp6m2WC
44P3cjl90pOH3AYRYiEfgikhITP+Mj4zibiwxcHoznFvImilh1hHKkSlx+vMG8B26ok83w3dTqRu
8b7Sj9nXEQve4NFb2cHiSswlin3ESPNIhh/AGf5sI9twGoO9h4Tp8GO9q0nWPhXxfyHeJGBSTX3a
qfmS1i/LahXcNOegb5Y8HTYQdOxD3L7OMrhgaxf9puSyPvwZnxhOm80ljgxXAXdZCZKlg2BQW9t4
WOlGjep215Nqpk09bhYzmkJgSG7OJXx1cunSNSVtb07JE3U9yQ8ufQcAYOjx9EpK5DDNFFdKbVqe
zehRDVgaHnvIuhZ81TJko134rnl6fTIYT+l1M4fYNT58BkT6ILE7jS0s8pJPZ3/PxcdsLovHbs1g
W3PrKCZdoXF6gV8/0Ol3fr77AMi2wRtL0acEcBs5SBHnrLwpTz/mSfapYMsMPWy58B6LPSHcIJFZ
CTAVijj/7O+voVmKreW6n+vqG/O1LiW60syq8+CAVeuU+Xv+h0OTbGd+G0jL6rAifR575EXYvBUa
t4D1KDTfRsuo+scbH2a0jRUCaRqwbNCQbbSJv5H5O2kivrxJt8+Hu/oxtTEwFP7TWdZGs78U5ZQX
cpRqaYgeFlwP96ZMOzTNsW09Mh1ceL32tDZ9YGJMzQ/6Vi48jL7/BMoL4cJ96QQ3sWASoVCR9Piz
W4ioJbu6g2K/2/pg8/wRJf00ipO0rWaUdzYTsVE0l80lI/0SJXqgqi4Q7wPMW+7ZRdQk1f6vQOJ9
yUlAcmibndvriDlNbcFim169jebFNfpCN+OAQi+HKdLPhIaaAgCDmM7vD9S1xtCEJtCDXOsRrd+y
ODAWCiHnfJVjeqXM0pNJ9Qj4b42UGK1eHY9nqTWVSjq1cInM5WB6dCglbLxWrpRwiAC9HRK/sC+2
G9Zgtt1MA/VRGNlR/ZolZvXo350v6pChdC1Ra9iFYFeLt613n+gYH6yPwBBjLLQtLpgIO3cK5CSS
l8u3y3vg7ZmbAlqOsrvC/cfqs5GNkh1imiqNpeW5sXitu5W8S1Z9LefR+zNqj3XpjuFI7RrcFmsU
7gL+ZRoSYh+p5xtSnphiW8+4nPUIyN8eZnbfPJRKMVogB5OYTomTbVfQng83zk75TIue2iWi29TN
0kmc+23LrlxkQTPO0p7h94dBTUhmF2F69lCBkNWCngDA1XRckFqI+P5v2OdN0mZ4QLVk7mjm4mx6
pcbd8sL4y8+bskww8R/x2TaXNYnX7Rh5u2pR9RZjUd6q4Fxtwi4uLDuJL6kFja3f59KOKmHHdjiT
Z6iifmiALRKMMtb2hIPfl5O+9K9LsyW7LEL968ZQKLc1ZtvnHSoLgF0uxL1oyjVm2xi0w8N7pKso
UKxtR/htirRaA6Fahu5ZEiC6VK+z44T2+Xwv/Ngj2uqQRdqUu/1FEbfVoaD00TDoEjyyETNePD7i
k3nv0CxDIKfDJ8ay1nKqiSiKcDNuonwSuBYCWP0Ldl+tZiaJaQTXF3XthPOVd/WymWcS6Xsd+O3v
ynurzgZt+IktGguwUsNp3tm5E6eV+i0QWkPSTrRzHDi3zHE9xxOKIqWL9uB8A6f9qA2lNZqydh/i
YukwY5D884BSrIrYk3K9dslfNaQYxSqtkKTf5ZT6oK7sny+4gl5treZvfm7xUlg7sD5ZQFAMSOYI
3j+si4zjyl6KusJzBeONLDne4ZYZtSjuKvt8r8ivnh7i3Zr8Y8qbRD45M21pEuJUBlxuIYAdkqDy
Oq5O+YlC4orkbuqvLhbH+qkVxwawlG9pbRm5BlsarfCqfXG/cmbtP25aHG44Cso3fkrif8OaCKYT
WxqSWLKIpvi1GWjLjPTjJVxd/I0k9LFF3z14l1etVs7YxthE8WG+4Xqbav7DtHGD6M6zbIdisUoN
SBgaSA/9iYd2EDjHUrtoddXTFIYEpkxSBxmcil+YRsOaFYc2Vfgi7xQtRzaDPw0jWLpDwWDzh30n
iRb0b8LlwV4ky6zdrfmELMuseU923tjIxscEhLrzDUBDZreuSBnlAOSnYgtXu0h5V4zAxUXIdbWH
BNZ/Amcn6e0HK4vEyS8nFhRfe2HPcM9gbXVkhmDf2/Elt0Qmx7QssARQaMrfLJhefE4PDzBSitSZ
nEgN3SI8ZvauVD7nbOgsN2/arPcuTZKWIYJGLVFDIEKuTXLS2gr4u7zDW3OqfOfq0Td0v6xH7mOt
zEKot0rA7tebqTUFCtHNNCWx0xAq/ISYbcLT28EVp1K1h6sTYyQgb1icom9tYERpdq4wnxAbfEj9
UsZRBHpGvwW3vRAhdh6BYV+CRgFLCm2nmsXlmO3WB4l3HFdXrS7UH4vDzb+Fshsp1AbMRYf3VVFx
c6PO/Z6pmulZt4AhB09/3Od0LDKBqORK82I973lA7Me/G+mg8YP4NlKgp2lYGYxJj/QuVuY9Mr9d
8ro+rGnBTR4DiVSfmdmzFbUv5H0MZx7nCo2f6GJNWw/rIuuZ/0S/bli5xGN+Ral1c8COWns0xwpi
N+DeQuPu8rXeL8zVXFhCQO/D2m7tn+3JH9MEkGD0xnDOGS/zfnaiwUaMfIi0CRkFM9yMj+g6it4/
49vNgKZfTMcKdhF1U2U7AM5PZHaNCLZJPEVlMOMgsGJvzS0qM1GlLWEWSM4Skn3KWPY0gVUYhbs6
cyIvsv8yn3RRcw92nMwH+PLBUWXogwFulhiojdxmfKGQdNWq6qbzZTESQwC0FdS2c5BrPKmjIP0q
Zra34i7ufmHLrFfPvJrF7K/3JvUmjk1N5rRkLvIwbxXJrEsVOqFCmCP3Rs0f6+gMS/LR+gakU7Lu
rr015Pa35WCwFbiB2uw/U0hNQB0rnUXI8XlS7LPUv2xx8zP3MI3bNDJaF6wtMKP9pJ1m8AB1S3jX
8sqyq4uS6gx969sQPTv+S4xUjqnMyoGmlUVlP0kakz2y9jdUYyFEfYTL3JLzv5sghDZyX0onYM/r
hZF42ZJ7bNqUbqUPPLvhpL+mnG1S9Kdc63Znd04Vv79BJqt8fZQolVf9F+sg0qIqMxMAUajla9vZ
pSEasNFny+ggKG5CsAFcOSF6KJypePO20R+pFwWtI+bY5s0CK1LPuo30oA60f0ZiY78zIPESerKG
U05P3ul1bEiaObna4iCLQgMmwBJT1RZwqJhHuYErLlKRqrMfUtQSVU2uRMtB+xAj77BFnFJhtVUq
BjJyiYpX8SoLS+7bNDDBhIxylVluQREoV0rGzU1UjKzXOUhqYqzZrN3GiaOQDZBCRA14cdsuy4ND
Qt73DJ1ubJYVQCnW/E+txdaFzMl+QARz/4Fga69JxHv7jRY5Af/IxeWR1qiwpBIz0t61p1ol6iZm
cqi3U57jqLRCfi8znxcRaetI7Y4W600YYQ4MvA6/XGteFCdnSAz7eehR9+Ch5vCNegje9XiDWak0
Z5qxgiDA4yUugVl7+Ckq6eFE/8cmhDHVtIFj09TsTgzv8D2dFCTqysemYxlLb9P52zhD7xcha9HF
oIK+2jtmLFPuxu7BnLoAQJyypqcQqI7lQl4D40sIdgCDW8roQ7ju/XIBDhjKjgGd1AwaXt8V4Hpg
fgxZ4sEa/xTO8HcDvIvpZWqBGgoTqnEnQvLlMNMnxVLKSMKOzYXMPTYWxLp46qWNZyN6uWoLys0k
Xxs7zlCNIjkl4iaNe76Zd0aSoTAP2rN55slhbGjY3tTdn1TA2aTsG8gt+QxB1oT/O6QYhN2Ll/ba
Bk9i4f3utM5lcjd/ykRFzgOu7Yz7fwCXnVHHXE1MSI300rIbqx8JXKdF3o5mGAH4laopyNXKG1NU
TXDuSqEGxUH8+S2erquTmsI549haa79zAx2cZZryFQDoX18/kykEuzQwsTeO+OZK+NK33lVYO0WV
IuLC6IKAFJV4Dv/5sa9pD48cfDX/vg390+td2tGtT8xwtPAsgxZVq8iqpsxGh36fuTyY/wq3kLaw
XxmllanZoWFI0PrPEXQNPyHCzo+mf3Opu5kp9lfNXcWIm4K0K/gaJx6Pm+9VS6stvQFmp9MSyHpi
5+HaicU4Y7i1EPkB1Ln48eMaZ/36TOtM0c/wSMrzvknROuRV1hxGl8Q3qW9ts7ocb6MJXV2/3CT3
k3czRNSIhPbj+ebjVL7eVrnKZFP0yhkt+ZovQdgOHAytlUKEXvJkhio2YUN1UQM4ir5bp/FiKdA6
nxkGJs6ycnGHKQoY9/JsHVlMVTdlZ6X/HRdrdtffTCakMHvlUxUkEpW2UDrc+/uyCuQ6ltPtFpHq
IUNE6dxQgcYTjkFES5BG3rFGcOgAIHbQkQYcAoOMCOHyJKmafleEZnuyAGIW/1uzBBjx7QlrpPq4
XVfMKxouTTdLawsdWpRp43uBepOu03TbOoVJx5u5/ZjDDWUymflZ550trot4RPrB3HOMP8Otj03e
lEQZM80qq/kRBIeAKokNJ5Mhv4Rjlsi58MajZg4pldyItLeOK6UrtlIiAQALXKuU9nI/+l4RTCTx
xQKxV7sgi6CpPVxVPvwWCRK/Sz2/ZDxyVi+xH0zG9vkXYrqiavAjTbxmioIVMDNIkI88LDWAfDeE
ZtPwevZoe7/njQNsmP944oc25kSbO+sV0RDt4aapvNje1T9mPgR91LlYwdnJzO8BPeEQ81aSMVDq
qn8Y2WUnoIaiEQIsRb0oSaOmqaVzTrID/feVYyzJecVm3EIvOEntGnxuw7wbj2EbyZ4scAekFmce
0ey63xGjUJKeH+YiWVXoflPvxBr+1AFefJT+xihm7oh+iOWyzoe4UJvAtc21sl3+yFEQlkRqwzHC
rSntWm3H01SbPk99oBDovOKrg9WAtpRErpQ6y5MZt6Y7gzEWOv18+GG5saCIcswBLqEM2Cu6GobV
sOcAeXXk65H+YmyHBsXYsSiw9dn0KH+5cVnKZynEuqWzNZHGxS42s/UBTnF21UaoUo5sNPr+SGvg
glkljdELaE6UVTHo3CU1ndnsviLArGoauyXHhUq+E5KlIF6Lon8m63JiFhCf/b4Y6RzHA603Tl+N
KzJfVodVBqBsbr2mVejLRtwHipB3tPcoDZcwg9cc4amEppYeZTjMzVhwn17fPwX2mfdZM9Qr/AmA
2pJpsNP7UOXGrApZargZ8SkPwyh9UKFd850C2BmXnrm6LwT6Utl3TPvEgFxvEr1Ekv0TqzNnCv86
mAaINqdHd7/VdmxmTxebXWu81yoOo6Misv19ymDYQEZpoZc+nORY+17a1uvvy64RAwc6fSOCtUWE
lGeINswQiR1duWOKFhppNPZ0urp+QTVMxv6j6FlQ5/UYk71R9ifdIWdCIeh7s5mgvPB2cUaQ62D0
JL+SgY2UnPRMuanjjbEfQc+Gog6CLpQ1yMBv3SmwThq0jzukJjnqV4IYLb5hh43aYATxBjg8LPN5
ehGpA9xQy62+877whL1ALZ5VQt3q6HBRTaAExdA/YYlw/NqXPEzFovpHEcLn6uLbcXU2nZQZT5pf
0SiT+2NtWspu/aofDC24huj0JEjKHAr3VEtALVbVv7fbMaxYahtPl3sz0cT3LaFqlXpgX/iCzfBj
C5+29gSMIPYB2EPn9FaxPXFjazf4aK9PooFUqCegTCwveDsh0ng7k2bkGS/dmmdMsBX6ck8Hzhg/
SHAIUXGUx2Z3mTXAzpQkjrHSGxxO623yrSi711PMb83aonMpPJv9rOT+mAJ6RZ2LC/iGaLVY/kXT
g/Lh38r5ok4AtDE2ivSjsdNR21a4ojkeMnkBzTVf9f3+RemRf1TTU/cgFVt3nC85H08fIL+lHuIq
GGyio38xo4kCIwCEzIzpS/Z12qA55Fzj8S9Slsukn0FwM1+hWAPeT6POVtvVh2QfCt5IkkpjG7xK
eiiGelbUk9S0r23AK/CaaMBoyIKapqNITjVycLMthIasRgwvlBF6d0XNo3P2bcUEB5/b+6qwyE35
z01FW1j71ED4nAORmEDEziILjIkN0iFAbaC3ZUgwAfqhWNO5HAWRoZVOnACOkv8uqN1XOmuXVNtM
x3uJCfPoTTr756wRwobHoLcDbQzJiW1Bi1E9WdR339n1npVGMl2hhybcYgucWUtYZ74Cl0O9g4lL
EMCk6RzRz6E7mdi69SWtSPCyoMyYS0FMo3jNc5b5Uub7UKDW7i9Z8TE0nZNp9r94GEueYl9JL5xN
2t8buW2CemJVgxNBpBJIkRN+/EuUBsMeVxVn3svQq/euw3ojL78p5dC5L5whPm7Q+/gbFDlB6uh0
I2TdswYPEbAVdSa2H92jDtAD2GnQWc6UyrbTJXSE2rkqnmXl1SXCCgA6C4cka2g6A0geWcm/kzQX
Q4VKKobDfUjhu42ful6VvETAKX1Y1pjL/2UiBz4ayLt0Xuc4vzTsEgMr01qOk68a6w3iECP/JsTE
oJHynBB73bi8IXOj87WMg/JyX8RueX7NzSqZB0AHqvP49G6YXxJ32FlTf3LVwze/7E6c9f3UAfLS
jm9Kb9APn0ss5rDlU+dzqZ5RdKvUxXJxkJNlaap/CkHO1EwUMOe1/aVmH1t4WrGVN1QW4SYSmIMg
0cngRDNui/dvDVDTBxga1Nekop/vtyHVjQs2vwPzcCMGIxwlL8kVdRsEx/OFq4B1CBJbUm5jD+UI
8De6LdtCjtyamzfM31v593mlaRu6V695TRceQsCoI8ZVgjunc566ymqZeZVFwLjIC3hlrmwdZM6u
ZfDaQnxwZRrrj6t1rx3UB5jEnOIYrmjDAcYTWqanIv9Ja2hGKEoNINJOAcwUMQGrbfE8hGbsmaYw
7of0KcuYvW1hxeoXjR57oVNp8teiQxPqZ32NihmvCTe063Rvv6OEiS0uj4zi4tOJBRhqH2HpISgo
aZUD7X8FHK1dU/2T8gQJ9nLuLloduhpIHkzIt6+aGJvq11RF7Df1e6Byqmnuq09yanqIdIPzmp6s
pMVdQWGRmNglMMequUKlMWpqb/hJSe0uP+YihLQPzZIpkvUqD05hnuPaCXLEmyyyz3tqSDs12v3X
x0Ke9UHhYz27XiCLNu6wI4+Gxhd/J9pnjzmHDtYZuZm780zFWuaqPCYOsVWFT1uIJLraZndEtcH2
g1t1yIi8HZ2M8ADeqqStqQyoxD/QjL4b2fffjqj0X/jvJ/flgeL+LNHDKsQjHtuWTIxc9p0tNDzP
IjPQhcCUvC12QV/iCi75StWz6Ludbh/zdzklghO5dNZo42RHORkw8rzRZLXO612nnUeNwvKY5nFf
du75baj74duuhp5Bg6NMHKMkxlK55wgOy1ffPDfaw+RlFvmW88+871jzqCWbQKC0Gzb8EsJNiwNH
NghgaKlG/kyH8BzGpv7gAiLDRE6wPE9F0phKC8qPzzf1nuw9OIdJybECxDeShnxIHkfx2usMfwQ+
yR7UMULdoxdFZNO3MpUhbHCfFunoD/zj+LC+A8sBjdO83Xo5qLyqRtsBCassI6OPJO1KP0f+F039
5ZR5Mgaj/1HwRinse89y/lt4W5LBJ1UyIqB9HtveSFGvlUidm2Poh+Qr0PnN8qWJ6Ew19+egDmRu
U3/qIrfpPy4X5jCDnCgOkBVfvn1QgE7UPJ8pSWdkb29YcJuQgADYQkletFcglaTnquuT/MhM1Pyj
wi4+bf1OCDfwCNZ91ZvTSgAVYRQasWc4UWYJNBaU3qR6GTxY2QgctUff1heMDhltrBCWIqQqMHX+
MC2iU5DGxOVwHmnTr80ACTPqj8pjSWlMpktzdnPeLM4iqUAHo3TJ2qsx0rzr/94ryedmP3v1P1Pw
9oXVrMDnI3V8KxLmUhKbf1ZekwDIbKUmhKLi53S4Ug3w+urJjD6Pj+m6b6rb5IPJ8h8X45DMisj8
Eh/EjHl3NZUHs3XkvebUtOasYDHXqPguxfewjmbaFksgHGNHf+yAQqjn05nHdJWB5EtNLNCE6t3V
qe7fljyDmxb7SumUfxY17USvNXdo1n+nmfNq2VShMHAZlfJ33oEBVhJztYPhWtXmC8P/Dq3eOrRp
Ik53GK6Yn2aJLqlY6alD3e+jCL+FeHQX+ELsZSuBj6O3WQ5yjQ/BJRAhgbZVdF0l5V4V1i9Xq/+s
Sp13dit6EDCLGBW9oYwbjgzUhwaUNu0qUAz/AXIGV9Ht8S1te0lGf4TBSLBkAbL2zq/kLXu9qZ1e
mAsmp9Q2fjmlGaJfjraS8RcXq7fQH+ehVPwbEkVeZlUdXt++HDZafCGvoFP/CfoMVLJojTJNrFy2
SN2OyWsNNYBV7I8sUmBs173cOUQDywFku6+Pm4ziYxDGGDbAahrweRVjuXAUVEZgIykK1jadOuYP
+YroYaYH+0Ii3+7iIecDzxRvtoMxmc1IgOR6SCCeDSO1eAqYk07D3s7y8dngvkD1iBy7PsgR3U8l
tj6Gspy/Gl0Sh2p7WZ9xu4h/iJl/2yONV42Uvm/4UJQc9H3FE175ziC8WQPFrP/jtKWoyduKxFbO
Fog2UyD3r5cbCCLqwxkYEoeBtuCDhdHTKVGJZV9mGumeFdDE8QsGscoRoiWhGeDN1XefkBBj0SYq
J23mahDYr4zZf6HkRgfEtHvWqE4//eM2hcniVLi1wDaZ/ae49cHZD3t9YEoRgUfwhwOSw3FLu5cL
zNNBxYcLahbs7aRC4P6UpJD384E5CtN1Od1c9KMq8/hO6rqgRAmrSTtoq+rl3Bw1qeUzD4H9GEOQ
GxI+uctd5vNGcMFio+0xS3nNWwsLyUyZiJbItT0us7AYzI171GlNF+WCpDE6PfJPFbv66VKdMpSJ
lPLUpxjaGO8uubr75EkEYJBCj/rK1RgRIflJfNLEm4ohI+nLLnUsmKir/GyCWpX5rY2T+adyUUCA
aSILYqFSuMuB8CNSsg6PfMc5f2R3FTutYDCxWC2iSfRnZLymaRC3HriDaTOW/ldDOIILY7OUbfwM
OldUZyrBqQjAUO0ppxOMaZz4aPK8/OAnbr2snhME066VIPY2qsbX7XvOyjc97CNuQsxPTfaZ2OVd
dkNf44OhUL/wsuHcbc3Uqs0I8Qeivh2udDxMVQhGzk7V0HisDigEGSKSL5h3q7KFcpUHB0rQl9hM
HwL3nx4W2VDLc0ee6rOWZyMyibMIIpuyfrIiHcagBbIqDsbMYNK4H++CUUMBiswPZHl9n6fOl3UY
qnfrT5gsSsOR8MH+pezGh3TBJwI4nudLN8eyH1mCFrg/ejq47xDj3+7RsUgwxwl5EZfvp9lj9rf7
ONjAYaXXSgf1o7Bqzy1dc8yu4p/oZhZnsXQBZOj5zZyEEEPMZJ+Tqf/fJntyXlGnP3W9KdV8VeNI
TQVkCb6kTxnj8iqZhDuJabG4f+LpHgMQikDiD6EUfBSRVsuARo+7wW3VTkfWcnoHIA7ud6T2OR0J
i5nNfsDslL/lNnNT2KaLBMCMjgzPSfsFuXaYMmbJ1g62cGdlTpogomLy5gS2/fJEqILNGjDnMu//
Wtslj3b7aV23SkoLasDr1JWKrHq+UnwmSrUO7/HccWj2fmk+nXxchr5+TcuW/1ptNf9TU+bXwRT5
jQhVOKvJ2w4+spvx4iQc2kcyce9impO98hiIfRjN1L6eP3dgltkNGfKN6k8o370+dHw0bDd3MOI4
/nVfSOItHa2XOPWvFSowvPWoy5bEB61S18HvVVz+3hBewiBHyjR/v+R3TstlSuVG5w0FfYCytqeO
a5PPaSo9ISH31UE0GVW1pndrYqRW4VkhUZUj/5YrPp8OOi99gGaj82/mgJma9cm5R1Vc8oB+/MZ4
PKng/kbZBTFY6NOm7p1dsTLYN0JWQlejYDUMZH9A1Pdcr+eY+ytgNTeV/pYA+Rp1PvG0E6fb/fmE
LZSA/boHyJiHWJx10Aa1FVzWn+Gg9ndqXH656hEgW0x73FOzenfy5Au8wmfkqr+jKmACIGqvp30w
nvgYuNsrsB0djUa29cR8zU4QldWGj2N+gxvYgnSMuFHmnI2o4hYMPodR1NhbfL+REVWweYzvW2nP
ljGsANQ3ADmZZ8pJu+nHaTFsDNrQwGri5hDKPUTiAohMUK6ti5rLaaCEUeLVe9HGf+ouSpU8dQD5
Ot7ZBoNvTk6hjQcjwCae0CNcTfo+MRi3cfJiAJhNrhjXaFzOORyBfvQW6N4zphqPVeJvasHpCiYX
GJzkfYMT95vBpCk719i3rEIQ+M63cBBFI738LN/Db2eIekJNWqESfkaIOtxKY/maU42dNeRzt0lT
VLPFJBCen2tgJ+0wEdUKNIlB+5SzOnaiGN+0nXXn0cr7Adz7yenWXMks4h1vaM0zSvJ6bb4o7r6/
SVy5dgICnp3h0lDor4llyW9NurFyqutXF3m9AHm1m2dx9pD7o5gl4jEin7YICYHG2NmH0ZU4tUt8
vYYKxXRoTTGoWU0eTNpXPFbI+c9Uypc0qYwPRFHq2On0eRvobQ3Jwi4nCGml0gjsQO7I5vlXNh9U
UAUsV+PCbmvyD1yVBLl8FDxylSY64HKyj3JHbGR1X2iMcStSTX2llnKk0XgQukCjes3aOCiE4Dqe
djmAFsaRIHScpt1vrTuNUIaTySbOM4PwL9ngkg2UhRcnsP6ZKXkhqMSVGwwG2nX9cnjxOBV7fJKQ
qni2sEoXZ2GpkkjWqs8mGumflyN3hUSM9OIH7PEmTm5a7PG5rpR9Kw6KXpeqIRpcKt+yjCtG2bKL
mLwTclQEIpzkCkEzMzThUZcBVZBF+qHPmE5JaIr1QPAu28V776nH8vGHvr80spFuogRAWOkL9/C8
g9rR2+VoF6Wiw/UkvebUks0NQr2iErLVqWLSFAZ8ikQ14OQjEtO7R+tsBJx3n50PlUsofDv3u4+8
cMuukPZUw+GDyD7Iyi1CUJ6ujegB5mQKiGo59MKoTc3Ta5tFf3BoXyb59dd62Y/Ln2sifvw4K14o
5Xm7QhagNYTXdGECpH0eocJQbOn0Yv6mW5VI9DeBDi8gDtb+cf8kiQme+tIqxkftxHVXbjC9+k0y
gjlfqF/Tf30L84z68tZjDdQZjhLvo4Ykb+pnWLbXwIvS3V0AZijqydaIVJZ69ZGlpDyJ0uefYBDc
0PrJNqxPqhIZp+YI/p7nxfiKjLOEO0qLADqeno6AWtpkmS1MJz7I0t0Xbp8Lnc4Ha0jXd5JBXYtH
O7fBAGYKQHT0I2AKPAraKzbTE69TzddBgAP/DSndjaRSM6PwGAs6pHyP4ZnOmzqi6MNXiiMmUM+p
n6J7XBpzQnb8zCmHddGLFOLzw8vyHt6kD+1QomU6m25lM0iHL7Xyndlroc6ex/6XcPGsJ+4yoao/
U4QeFdw7401TAtXCAv9S7tKRSJJlrpMvRsdnb/ea/jwM1ezePpls/dILp4fPxP+jheE5M6VauyCw
k4pmgTm4dDvKCnP5pH3Xzzg3f7P3Znuu8+bZC8gT9748dXjzVtN0G/VF7sz1hwlMFKxUsI7XqRQ+
q+EB1xXNeVFzNHG8W38loujyoWV3Rih+t545L3t3SvEPVvYLqG/xUjly7w+nPa09yoMw7cOoXUhL
CwljBn/dxiy/YqZfCIBfT2DN/Ts6V8p+AVLsumkVI555Mh3TldSk66vdz5ciDcnK9zsW8XqYjgig
YzH7OquHNkFpZHCOQWChVIVQoQXhD43Do2XXYPWMIMlzwapbNL8XCMdRYLbem7e35/GWFFfyG4jj
0s4v1jl6RthiKOR4NBI9T2t5VcxTtMCUWf/74/UX+Qsyu19+jwSNUP1OOP4AeduR/GJbBHmDu6Fl
Km1tu4NuYfPmQ03guvVqwBDC0kQzr+QCb+oAe+V+8eAgEgpsoUI2LxxqSgMY8XaCQ3FYYSWUMZiq
HP/BzrqMlb4EaVO7JPbYhDUBO0MqEB9WotiL8L5/pOiFNgE1+fDCbBGk4/RoPkyl2XoJYgxiHqmL
genpf16bcsSBdjnFDYWeWrUuUOuQKmv9BB6oZGW7VJNeH7OydB2g5LvhZpj4Pzmx+gGM4JKzRo2n
94KncL3TrP9hGX4GF+BqMfq9EqfJIzyWNedZXEgZOAqg3/CzPOdV7mFcDNT351iNxHpoC8q51Vk3
PKybnu/oomYVWuUoJegsj5zkwwfXo8ukdP/nwW8GOEI4hIp0YriJtVUjvOMGo0cqAgl4gGWdbjne
a4BhMScASsXEaEoMCrn3fnJkSoR2skMsG95g1PwEDyBKwZXJuR1VXdaAkV9jkycSmaKLokt40rUz
YL+m8vaxL353sD/Yq9K81B7lcLE17xfvgvM1stErA6FYMLXAmq50f++HiOOUDh3IIoOuRls/R8RI
DWL+7+nMrKh9vBp1zjLksV10GumtsEg8i1w7TWUF6A2z2IAjRWIdEC3A6rOtBatUoqtukQ3rVWjp
KaiDwuyt4SmvrMkW5ZrDkNj58IyewH1c0ivangZAJUbcsRXrjytI/A0K2PZZJrEScBZkBS4mT4Ac
p3il9IGJvXGW942Ps5A6LXN0OyIHN1QflKGGOVY/XO6nWvk/KAxOV0OTtO/0k2vdmRQbU1axbMWA
NfsfTdop6QJlVHQQDDCam3MgqKyTFsoD+Q/J07P5BZnbIA+TqaX7lOY03k/ZoiLM4nuxbCWz9WMd
1sipLJ3zMKFQqTdBCAzY54IqjC6JW6nM5w4MWu6pDMhU3WPiPg8QUJkyaNo/3TYPA/REDo+yiG6h
DtJDH1GUosyq38AY9T0kCoxT/wySjYAcc0ElNwf3E1YhgruUuse87mujafrDTxExF8H8XHNya9WV
j9VY6vtmCPRUT1LgFgO3+ibNE1XQ/lNht+cSiS+chlSJLml9eGC+ZVQu420qGa+t7pRck/MdKfiV
pLamHdz7FNNB3W+5SFJis8VS/yBApVT3CLx1YlFcA0D7yeusruGudLWzvMxtmMElouWyFLQw7iRL
dNN43JBnL9pR/dGXVBXS4FMlEbFAGs7oNfzPYR+VnYBn2/7FCxNHD8upAU4QXk3xtQq2Qdg9iTPW
pcSuNGCfvYad7POm7jiRjaMfwz08Nlq3w9czGTUAbp6kt0Q3m1BFALsFttgXUxBrQmulhNYMU6Ld
oEuY092Ww9In0HCpXxamHq6EwBUIswOF8BMN+F8tB3EcZJAltSeB015G9uAREYY56PThOoT66nvz
aQ7dfStwoL+UsTVDSbYdPi5HH2t6nNc9i4ox+G7ja4sZdbOXZMDgY42Sbdpc3x0/b43e0N+Au3Lo
obnAayDE73xsYiVAPjp9bh67flc3b3E2oj9/St/lJS5kSoX4Hrn2JGxsbAW2J5Kochc+lVyhjHXb
cbqd+EqqFWPtYrviksSOIFHMQuZuLeframpOgWlYo0vw+T1blr5dfcJPqfUlxG21zudRyBDqJTSh
Q6mmgG07p+YAW1Y9NVUbdGBIv1/zWzzGTi8pQXSX0xdjedCt5LPsfee0DtTsHeelVajzxfu5cGSy
dUMU4iq7i5Yy+mp7dJeJ1dImJhISxCzQmTEYRncTAk7blcxxH2zvgEYo48q7UhopS5QDlf+Acldd
zqj+lMJAvq6n2V9LWmer+QyaFY6pCrqGC/yJnbfjc+TQX/cHQH1ZKukCZ0rA2QPNKVZsiTzUKl3B
A11DvKdY7JLFd582CSPOBO1pcHMKRZZsEd/DtjK21gOajj44qdJuixfcjh1gOb9/QbQDdFkUukJJ
hTIhB9lg3H3JtXPTxmCQgIUua7sS5gx8L8jX/+2/Q8JgFO6QnJlbjb53Z2AgzwjF4i8sod3nsigw
nauk9Xy4ayWnMsOK3QtQdyN4Gug93uaurJb2TOj2xdDDrCe42syTMpyUGYOtlDEydAfN6PLTD/Ak
poTLn6dT6qT1LMVIS5FVDd2hNZzG4pvFOJMO1rZObNlIqO4DelxPKVLaZKTk0Eom+01UTwj7Pdfc
gc8U6jWDZpgmqUK6scBiOiBcFmmL55170E1bWH5gK8J7wx3XES4qn/xTqFO6Ged0Yb/sKQEO+flP
PGTGs9bW+Hy79dQrtMp7I+Q6zg5jksGOuUaaiZpFFp0bW+REGFeD8Dq2rdDN0MVGCDQBaXUjt5i2
MQ8nVL43kQF8Pp5ncX11+fvGLpmSyrWWAku8O/ixUiT7BNeE/LNOWVX1//mg15cvpBQdJWzT5dQh
IdU2ycwYHgm0+th3v6Y7dosgp3WcKNSAFSohnpAu3PT/6EKsTxwuP5sf1UPnA2UWPY2ZFsZG363v
HRJOhCvaHqurK07x/KZLbtgcnDU3Fhg8ywVECLfPsT5+G5RyI5Nu6r/K8cmwKEqmij8+udPkW4My
zoov6vWWeaGBPXTHv+8Mr1Z5rQ8u+g/21aMcnnM60N846H6fyPRkYJ+chssYvSHhopBC3DMpU3Iu
KlwiesJbAXZxj9ojOhIvD3oFCKdaiYBgtZ1qOdo54CP9I10EIwkl4Dj0CY3HG8Qm15KyhXZbJ1/b
vKfs/IAY+3ZeFl3fpN3ceTLj3j/zskfjeNn+UfghIhyra3QRv7N+5EfMeDdYCo7xejZ/IQLx9IhU
j2/IgCaiw9E/KxvYyokn4ZnwjL0sU5u79vIsK/SkXmUFPeRevXT6DpfvvsshXfkxy5eSx0cxLmki
t4IH3UOsV8Jk++sBmzUDjvVLxsZQAHxTfFWuMF6feahyM0aEfptQQQnpJ5iyDmLaY3dGfw41UZWw
AVHaLR/VFitP460qyDCID8yjOVPY3eitbBcyrQquIcJShn47KGEKGmobRQdA9G6EGL84iOsCavaH
DNCM5vk1zOh20NhLPnOR3N3Ggv1v8UjyDlmk+rGcKkMRyvCL4eiAILXUpjPO/RjpQOU69LbuCJJg
yjPqKp9xJgOJbKYIMD+EmnpNIRDN4B1GZkdE+m1K62ESxVAO+1A5gRWRyBtHh1Lo9uuIbHPLhQrM
kl3UTB55RTDUUnwk2uh6ky3Sc4zgfiZuvzL7SVBT1FIidnuwtpQ8bBj0s0K2p+6xJH5kwxz6tKnT
pjMnB2cw/ZUsbm2d5w5s3+/JDdIZjYcJxbnE0UjSiAmiY0bHxVIkYJZvf41R1e3f6VW+7oC051O8
w25UnWu91TszEvq/HjMaBg59HiM1JIdavDOm6ovpl6hn819/mrw3DDv4qIvVkdFIuOX39iKpUcPt
Q39e1IT0GkKlcpDRuN/isGq0GnVVmR32D3Vnb4wNGlt+ifXGJuHbYJfXp/ZUfDojUwCqjmv6vcG2
QD7ekXUVMNVp04ECW1RprR20pgSVz1GNLyZJEx90EU+Ho4GRVknqOQ9GpKWUQn0zhQz3HBMuw09+
DNs4/VP8CW47LbqvuYPUugbZd9IkQjVQoKcAoITqRYJaKlQxOUweU6TT74tJ6yaudx/fDbOTjKww
ChQDMN1EC6VaYaXNENEYemIePUCRIN5zTYSK9KaQMyRtwXHmYKxn9ISMckfp3Q9jeyX696nhk+us
qJuwgMeBBIEQSg+iKBnc0O5DbFs/Rph1sriMSbGLHkZ6j8k1TzUvERdeowj95p6wzS6dXhWp7ihy
YH8HYzpIIjUD+suRir29dfcZJk9Bpx+vvctqBz0fTqXkoo2q57jvqm8EZGaW4S6KiT7kIJVtbCys
AZm749OwCqkAZ2sfrHY2X5zGF7Y71DdT2IpJcQAaJbymkYaGR5DgR1XJ09DitlSRsX5xk1Qb3HSD
mYMQzE+DTO8pAJ/WWkPE2jwL0ZKkf+57RRxiNpAbazX+p6/2dwMojyM8F+ajoOYywXPugkqMhIHz
J5yIPHsG7yHixo+EWo5DESIKC1q8GMNgKtNYc/+JLXXPwz/mMsoyM3IjlE2fhdSfKe7cxMSjN92j
Mi4Oqs95WKYFr3j5g5v/N71XpynHu5VEu75zpR7bU+9jeAvHsUA6Z61Gck7Q8sQnII9eAaDrr8d7
9wdg2a735202FE5CbetSVKqVFnygIqt2VyxdHMkn1YHQkm6+lyToImwvXb7sXCUNsGoIGLLAOlq4
ZoAmQ/JhuuHicma7Kr3MjD6HrqmcNJ7JmFWXauY6NhovXH7ZVNtBLw+GeIZHcJ0pMuBbBu8GbBjD
/QiRJEtiRALcb7e8SiaBHpOpKMREQ02ShU1kl6SwKFY3Np/dDlNgiY5DibW/f/lDBjlJYZbnQ6IP
8dbXwOJmaBWOxWsp4iKJ5bafE6TLewXxBHTU7XLHJwuake6xfkUEg4QKuHCt/iVn7TsTfqRR1amo
tK2CR40xaIm1ZjECtI70ekzsD39qHjOhdVbmmHV3pk/cLbRY1i8txrZv1qBqoyraNLNhD3H3Fx0M
PXxrvAVeURTDamU4LWdKndFqrFJm9qfNmR1fv2Sr3op3FQp7OrzKdys2U/PrlJ6h8IDnJcGkKSrL
aUvAbffxEBp1jDWql+qT1HxrHhxvfr7CpnEx1/nVuyx+HifV0RniFQhZgUP2E1DUVY0T5EPW/Q7B
hWKx5MdyJ7okPXDfmOyFxdnfrgCECWJb4vL7lflt+8UsaJKtJZNyZ9CaLeZ9ZT5vErQ+TpzpZyhg
tPn75ZDkqz9IGap/YOKbO55AXKqYXZD18a6T/IQDyVZ5y+AQqEDPJYY1JAa8z1NEmfh1oh6aMpcE
9tlzoN5ce8xNbgagmHJ4rLTyVqlX3I4bEq4R1ObdCV2GNTa13RYir5m2+7m2E2iECFuQpX0K5fcW
gkomSowVjzIQtCzoOlTt6giqg/2tU3nDqOStQMIisRsNeh8sawKl0nby4QsdDWy8LSXM9pUmDdWo
T+0t8OZzxhM4m0ottpbNzcncszTSUTdmkmeyf3JRXvwesY9yt4oYEt60EhKchH9p7EQ5TvWuBNb6
5rEhL9I0HIA8X1Avypc0yUa7eeVKiuBhN1GG8tmlHYGLKvRXAKwHf/viO2EHfG3Z8lJHjL+zU6O7
Un5LS/5j5+dM4TBAHJQvGDpukodiatzrzBGJbq3HPgBPheRubDAtIP2WhDigQr1MllR0YdGDXcfS
3kFptY+8+UT/Gd7/xtr3cCT1ajq8YH/EGK6ROjzw5e0dMYxBx7yPUxioMo7+xhQ7l2i3FzNqKkFm
n3kBYTyENVsqyvwP7kltLUvQTJ7ArjsHPelJ2FRbVbYiYrfuQ5nLBd0lbU7sBVVRPVNy+Tv3SiIC
Ig5LuPkJYMo8pKWEWxb49Fgvq1u3dX3tYs0IRw9DktHJYNMEbTGlpNmY8wQoGTSlMUHVI2aBnUGd
FAPd//7bjCMHsxwnAmY7hCa08DyUJTS8nRmO92yaDU4/RQQ7RFvncMtx4YjqsNvpFcqrUfK8SSmE
RBVFgGlesgm1zyiFmgz0JSUT7o/UzYx4UYUBD5Um6Akk648TmLO6cbUIKt6FJSXHXiAmovtyTFgo
JQj+1EnBaXh90hqEPWVUMWZDBdeUmL7FB73DbQqBIv3xTyK7tkLIPq4AWZ9d9duG9W4hVbKhMoTI
Kkm/O/fGSS8oWJuUs9PhcB1hZOu5E0vj2RvLrKB33uSHBIb5qweiw3gAqbGOBvZPPncpSCFkll6I
beGO8G7P0IlV3kGEhwXt/ZDlD//WLrU23m2KSEzasy+LLAcc12rdfzX4Nc75EEtP7dtRy/EI5NRr
nrtG7LuxCD4fqQddAa9/QFX90P4fZOWZFf7Gfvdg6o3bsKWW6TLg0Y0tOJc3QVPhIZ5X+e1OSBZC
5MTYzeqaavTdhmE64ghYo5uyJ/hg2xpz1ckEA9aR466ryfPQEPREOUm33k6g0ghMAQ4/xaFANlYD
o2eUygSav4YBMBBQpGr7yt76RK+85Spbe5yTybZQuF1ElqzHNuevjLIz92t9OT641xrAlB1PXMpO
RHL3o2lNhpJHn49WethmtnyfgR03loaB5MjuAuc05v8EN5VAOc7+eNHhfhWR9ASv6Gxx1M0tWdga
+D/8kxeE+rzZfywIxr5XiPj5IC+SqaiiBI0BkGYp+eKtXEjHzDA8CkyQyZvVEBRjN3qQV1YUlBty
vV8ipfG8pNZn1dHSKkP7l69RUEOT0qgLruXlzDLv/6twGVb1ERHuFH3E1Q1AFz2ExK+OqeVmIgLR
PuhOvDPfPRoyh8knWBd5dUjAFULtDBe4pvOJtxAGhKNuk3OTHhDBLVZ1KS5m0jdXc49mCYTlB7bR
uqCRXCvM82vVn5WBmoAaYAXPoglXw5LuJHzOzAiw2RbNqjJd7JA+5XBvZD+3nxEi3zs6Nfx5sy1M
MtgrvvnXMxRwBWXn62+piuiXgE4yQJ1JZ6r2MgEL8xOqxCnZvmN47ju6ZT3XnGrJYfKVqIJdyzbs
tFWkq1wd0GumtELb4wJ/0xlMseLVYvEpZ90OFroSRKLKLMtHySN8dVG+ezs8JTMHnqbHiCG4+b43
aiYOY8wdJRb+ly02itqyycaa0YizOuXbkTF43WauuzgZ9mrm2Wu6oPpErnaAwSoph+wcoxQWO9Y4
NFNarGq7t9tkbQ7Ky+fWeXkuBWhrlLX1ClpwCAvp92s8BnIlmcd7bdAMVTObH1Egi/O7Pb0+Pn31
a/ZkNLCytQTsJdxDX/fiJhvA0nqwP0cwmJmgXcgx7Zt4UMpOId5mD1gGWAEc8w2NwTlo1N8jNUr0
sPu6ebkDxTRl9AgK/76OBWG28q92QVhHRzHLfBn79V6rFZn4LlQ1vx5tatEBD0jRAspx6sgxvZgM
5ktGZsumliTUeb+6++zuo2fMJxKKu6kbi1d9UqNyzESwYS6Eob1RYUBfX80iUxuaddENHc5wK4jA
IQ20541RrWb8d+D8IZzCDEP9xFwSVXfI4TTUCXaOIWaBeZz9lYG0+tMwY7b03WobV9vH73a3BckX
VLrH8ETQfQZkS0MxrZHAShZOmg99o1HGXCQtErrk9C51S5zZDT5/SlQT84pQ/eHvTwCyP64GS1OT
ftmTJWST3sinG7bkimtSO1dKIz+bSKIQLAn24bUZHwI3lP5tVb3qz7Pl0xOxpjbm3ixTo2O233+F
OAAlvnp1rkIPZuTgmj35qSZ1ylFn/AYyD33/YIvBoXOQIAhlay0/E9v4GE8oEhPbVg3vKyqdyIiB
JgmWAjCLdOmkdeSXlIHMJD4XLfqZz7DE1KmuzMfSAnJ1qmVSjnpsD+2AbozZ0ldQ2c/LZ9qsZAAA
EYPLlaeO77zeLxQds6AlIF5z4yMWS6oN9y96PvAWftwpmNI+GfzwXR6ZYdwe2U/I31ExzYGFmmK5
fEHB2emTYKCA+6Gd9QewAf/iDS2h3ta8xY1nBYk6tiVm5VG//KIc/oScae2mme/4joNfn9gtG8/m
PYwWVqjvzdxBjPycuIz9wOO2rFDiTIR1EGfHc9QypzjLPICLaq9JFb/LJqi/J4iFpy0l+yiNvMUw
iVOBgMPeih5OAHuGk3gMeuBqFM4PI+YzauoJi+OqFCjYMKymhYj//9/MdFhvB7+vN0xEPaemrtoX
wuxKLIqt51yEzaxv4dUCE37RNsB/A0qJisdlaoaZyZdh+WWzqrQbiH7s48deza8/HeX33OysnzJE
NtTGbY6PHRy7uwbbRQPNecm+ggZMajLiqHwtEoe/1/SBdUjFYRi4YsxKTwOkGU/+iOu6t1Yvs6Iu
H2/k7eoW/PMrsdf5DrBoPEHPUEOv0HLYR5gMCCNFIV2YOyIRESKpa16bk7WDgraOnktirzWBCgN4
6dMwvnhFCrHAmGFIEcwAknN212Bhta521MgT7j2i7+EriKc1ZEWSiX9n6GyDJs3amXDjrF0fAOjB
PGNbW70P1v5+V5T0K8Cq4QwbB3C/DUtgbotYMC4wK0r3tzKbpVzB9z8drVez3CIC4A/GdVZJpH9i
70sdXy0plA8iXeiARZ/mKjffn2z2hMGDok320VxhzsimJl+CcFmEIuvt/EZk3ieKMDE+4hVS/X7k
VyPWb5iuF9g1yxqsTLy6p75pgYR0LlgCsxthHkjOxv9XnGsEoHlq9urQqpf+aeLtxuxYqnzuZiAj
rIjqCDnjiBeRrafd8nDoriT6G8dH9wtyD14eEa3Y5tB+0CWuvrCNRd5dJb2BR3E7UIqJD07bLOvV
ftWvrD8QigxY/Hmh9yaG+CyexXp6uCp44zNV9kciCcnbEplyk2RbmebolsK4qMeKcCo1kTmZBTpE
ZjCWIwQD2MXMlKYKRHm7spwZyzsGjGGZHvs9b8imsXnqRxRB3+7OukVpOxGCsLc4Dlt7+XqiIJbZ
u3d7VHiwOHJCWIyok/QDMz0RGDl7DHEgCp0yDIOrJJUEg2Yl2Z/wmR1wQrJPdBdPultzjqswbnJt
IZy1iM7YsKjeve5rTZ5sHCsjE0NzIU77otJ+iCI1V1IyXxzihYbJW7nWR8gFrRV/BtirvKR9qOs2
OZiU+gcX/PfLMcINNaWdFAu861AYbQbQOBHzj2Bl1jkIH8pM+wMmabAUW2+O0BlaFz4sWUzhSjF6
lCwXwdn4xxYXNfoshRvKA1CU9XvdKoaJyXuvHOlk5ItE0KlqP+32fxdCnw/gYJpwcboDwAUfbobX
G5doU1fEqlhEDvOURfu6rmyBtzM83V2Q0gmJejAmyf8o+yW5oM2TkQa96AwA49cmw4OdEKk1BXEO
1wSTI091MT6UsVUoJFLpj/umkQavQYVf5BFtg6VOjtJjCndqgN0GXcLtTYGCCy1UqZfdQsdVNA7S
/2RU2otQrTUaSmCg2PC3KF8SLj12yBrdwIz1jECnYwlag2T46E4rmRH6fMTC0fgV9rIwHVX6B4AD
BDWGNI1X+QGlZ8TK/kfGaifWkzd+ZolKtlQW0AD5knxruIC5ypkj7uh3pFbbc6r/d70q7APWx30R
ZUgK5GmYn4a2GWia/1hYfC7gbVva1btCMv/jVTdnijx7QJTcr3tp0DbiwyAD8ylmYJNt6/FKyo71
22r3OzacBd+JgQNkHyGDR4dEtUqjEEjehaAscT3y632EPhGElgCbF/FpDKEZ5opc8hq6YSSUptr3
S4auvCNEzfwI52LMlNGXIiNmFCM6KvT+lpxgka0208pMInWYt1bzm8mpqqY0PQq/SP86O2hNsqKF
TlSosVYdg68qZhdLAQ30IAWaCl9VcNWkxrTuAQhxVUGzEU8+fKPbHLu0XDajkNmOF0lGUhyEdS5V
hciGgkUiGSdna+fRfvR6E8Bey0yZlzUpiK+5zgXojlfgD1CKSkU0Hw1S1tdRlwcerR/iAljMB5k8
bdxUwKoHztxiKpxTnuI8XW+L+xvghEURwtO5zRx4uUrwSLF99rRTASE3pA5O3uywb5GUAzig1qiu
9TmfcFHoqFlAWOAWBlJJPkY3/xj8mtSzYD/A+3bgTfHM25TpklK4+DpQFd8nNHIyNXXpsFy19mLS
oEK0OBgvm8P+ZD7bWxnA6G0PxA/Rm9JacpUfY/RC5JERZg2vpjl4PV4CM7OO637QS7AtPLCp/gHR
+X4BedHbiVCUUJNMw+k/eQUhnfUgtgdp1EdhxtEAFjhRWVQg3ulo/1pCTmrbgGyadD4rDGTuC/Yg
Awe8mgLNTVmxNlrhm1m5g+Qf5vJ1fli7D3iyc1s9aiRNDvJlbn5y1voyg90m7hAJrr6UL3n5vSts
qbLFaPnj1Ok1utR1K4qWpD5ona2tWt9z6BP0BJI2Q84KyyumEZ7OUU5b2qV6hgc80+ZybKjyrUxe
AlnZF3s5JHYqc4XKN2IgT7mwAhFIOE9nNsQHrfYEib0r0jJwH5OViUTThc+jVV4nIEWXo7t8OmX1
F5Ud0zp+KUKHwG738X2/Q/XepgqUaMvd0bbCVuMq6WWdeScApb53Xu+QvJopj8vhl8WHl4Q9v0/9
/AA/Emjgf0L5OWseu6tOaudxn0MO9Utsk8QDdiPW15rhpQG32UDcxrVtCxiMyBMV1ovwWOqN2L+T
kuLXGtHG0UJf9YzWOV3EKmqD6jdcMm348LbDN3MU5vub2mx4TlJc92W6KJdT1XaV/Ow9D7ud4/uZ
5kXG0E0uznEp4vVs+xzr1KxiyK7KiL+3YUXH2/1o1VfrG4CbE8wPiizTte5H+A0Be8BLO28EDHsG
IuDzruWyn9Mwpe+k7hY6XGzrfrCMopstF3G0dZ6/M8lKEQub9bbcm0+rfNoMLfxO1vi3Mphyw/bP
qdLWuTJ2S20V2QQSOo+qnJVKN2VloGBjwTISBd3+XiOuObp9hRr4CAbVD3xzQqj14DmZgB4zd4ln
l6Kib9aWx/d4VB7clJuoEVdoYnc9VQZ0HicAG96pPYZ7arB+86Brtt+V/eDBL7OrpcxvkqXFCFFT
/G3crdIW8IPsmaBbHfe1+Vv/tEIv8iTQRjlKHrx8TIhvhYTPYofnogCaaszjbUGhx7xLYAseh638
PgwGi0HgBO8VceOST3/BIdYRac/sBM9ZkJ+aGSxE8Q4qtvOZpEUvbgDMMs1W7UZld2U2ajrbPEgK
mo046c+LBhFyK7KLc+G+HDPGVOhOtSDDHJt1sLZNx+5Bz8lLumZdWODeslABi4h47JT3F36Vmzps
1igDuFYpvNi/Yzzqc6tW6ToVbnlbQYDmTjVazmFM+OZiJk36bxhSuylC7c83iPKSAIdd3hAbZ0S9
6qDrvSxtkX8TQCw3sol5oOyPSE4SN0i1DULpeTC1SLbgf0EYJ7PRMtdGGx36sVECpOxoGbDIbdHB
7rQ/izsZeRjWwza4QiGaC9w6zOXSaMCh1JvYy4EOdl2ZqLra97bdaDdEqu1ntg4EXxppkSbyxmrV
Fxssmdy5UeYzipc3biX4uAieMt0uD7zJj0urVpY8Y3bNh6TSdw8/9jj7BCw5oSts3LB3UCHJhuNT
TUhnu5iOtGi2ZjjIpur30vQp9OynZs6r4lo2Asf5jyofZ7V3SkIjOyQAwpjtmWyxv5sRS96/uOaB
y/16M+Lb5Ys3O7ygMqYzxHWSfLjtlr7Oqh1MMEmwvtDFX+3v9Z+wWurCggPhCtIE+UQoCkBXwr4U
ZwXVICZXTJVN1mhYThYbKvCUxN3WqGt9a8IXIpjrGPLoFSHug+RDC+M8rsAfJJXF1060WcbMc6S4
poaZ6hC1W7HBKQhdQ6MUWZZWp+O+ZGhAYTnXyou+qqzYdErECbH1IcX3CpX6Cxa4yrXBj6OtHhbs
UWGR8I894ihd4iRCypIOvmds2uL6UUJ0gq9AL5ejNMfDOIXytbbgz6gmyzHX5LicIKb6iYVc435h
99Ec99Nzynde9pAIBN1HEPGofeofeuhzhXmbY91H7+RgMLGJVbW9SWuabftVZhEF5tQcga9pmo0J
0Y6DuNHIRbnKNtQ9fUNzw4qtz4LXhCzINdP4Sjwfvw144eWcV8FSnefpXB8eLGdKOHQqWE7Uxy0w
6BDcNSsukkIOiL12Dbr4VSyDMAOTTfB1kkQUz2y/cHrvS9nikxtoXy0kHe5JnN+QMSNN3jgsBnt2
ETRz3OMjgHbbcuT5SLpgWhNN3nBd/hXsOLG5InjPoy0Abx+o3ShLiJJEcvW5neFfshOMXqJqaSoV
FZmLeI/aJMv/yLM/w+u+XyBa7eWJB+eDVHg8vu8BdAB0Z/FTVZaQzT2lJJna6iMlQ3qfWIHsyQBl
fnDSRmoEkl4CKPXts264FheYX5wjB7q8GVsw0LQFHdJU9PK7AupFZ/c4zpKA+JdfZ8b5RGyop2h1
jLlt8e7UzRjfF9F32gAyPPhw+T/NKUHpCTsoIo/bMu7roKni6+tVPRWkYsn5HSVAhDG6EnwudeDO
3rlIVuoysGKTYRwHKOnYKckJUpM8cdvaFoUW3nNeFAexPaVS2SmajRk+kjRo0pfwDj7TdBILPY4Q
unlmUAb7aoNzih3bSaHkzNDuntzF5l/xoWg7m1ZEVtzmTDp5Zb/aqrXXl5l+fDFisuPBoGmdDiAi
H++WfR/dfWKb7ifZ4X0yjMfyjGrPdWIVkuR2eS6mdC8IAICoWhO563wf5pJ0f7cHnmPxc70Lapwo
xfjCMwXI5wpHH019XyKfMsP99xRyUREBj1FK+0kHiPJ+5bRWAO49SARjuX3WZnyz2fOWnnstCb1w
kAFKa8jyB2NM6oCcYnHdgf3HL7gKjZJvKLnU7Y6G6ZUYZoEtb8QO+ul+VnHbjzlpKuzSKPPDTJig
ffCU98aiTjOI+diU0WEHV9Hi0zoCLOYQVQt3FPU0XT02fNUnTlVSmh9t/0Sbp1Ihqfgz/VwZvofY
hxDwO/Z+h4BisNW+y2SiL7DTD+L1zsZJPhFknw40AbxQiqehORBXN69ahJ/FPGvJ0Hfjc7S4+T2s
rhaXspzhPyFWLMqhpkVkgYhTgKH26pXm9k441pinRKC/oVKpxxwgzBEQSwzak9Jb82IDIbO+4oBt
dOdJm5g6+eHWv2GJMDoIhWvd7/5NsXMiFWi3Q1TQrvGpS84YtrvzuUpudnkNqYyop9idnpLMlzQQ
s7rPy6NeY7KODg5bKBnPnnypNGbo+UYB6Kqk+jPVLom7O3JahEl1po03miM7mQctcHALLkzTxzR4
kAotNttcBaczUN3j/Bs2/xZoxGSa0eUXvd+DxqZ8pWmxUjl6ZsHhFGlixZ36EKzQ5eC2GI5pVSsQ
B8E6R+AxaMqbmys5ICT7x+258IfxSvdxmAC4jymFIGtIiZZHUgAa4ajJUkOcX1ec7BpeJNlSGCSL
qZl43WdhBKCPLY41JlZMLB2aw4rl3ZZ9BzA0IhrMcW0pi2fsLVlbDrJb/KTvTRYM97KR1ZamHFoH
VN8Dkp3v5idoyBt1o77/6wqXNlNz6IwiHu3axi5LIgza95HBiEIV8jnQJ6avWAwOxcTL13CvAEDR
FaOBvXU6F9egxoZVjZJGUyODV9n8RZQ0Yahw4as/bagJVXqav/VUHTS2gpjJL+Mv8dgE2s+EW7/J
PKTzE5PGpZYrmWOBeXvd5bJL33uTW5fX0duF/asLzCj5OwhcxOXoT2rxeKVrxL6qtxHGJUlAUnC6
XDvVha7Mq58Wn7dw6OMJncvZCj9s5N+vld+K+NesDmbPNVescWHppu6GkmUH5GQtDeala3FIu3ck
Tfvs69JogM3WDc5BkpRuCI8svL5m5TSlkQg0uj3rbkAFHFpicpzBr01zbTSsVyd90QwQaJFCbrKy
mSpu4ppe+rB3Ygkel9ijelZWZj+YnvH/7cwwKQAo2IcNdmS+c24syk29zjU8MWHnTdTtK3IQF65R
bTO1rqw1rqKesncw8XwMnJD2Gq8nj5dGPEP9rM2wFEbjWGObGvs4kXeXSL1Uq/cjjayZIDv4t8IR
8x4sjWz06DJ13jmksR2H+3yLKd8Ryop3GoSfX6oJ0ozaOIbnu8wNvFxj/om7pd8CUaQBfWrjfjeF
1QBtTv492XQPs9Hl2HkCIoO9JoJSfR4ac4thaD3MElljkEpYjDT19cAHEU61L8hSklIOiO9dxH8M
DL1TYiwL0/dEaUvL/eJfpqsZQnq7GgJDYqIPcxt4rtkNwPATRYWWjLl9r3GIkYfHmezM7s2+sFhc
vKm+t5t35cMT4x7NzZ4XCotpCJPtpAfTkmmWflptGiDIsYCzwhveAM6N3ff4y8IuAWx/9/4MlJeP
D6UDaA4cL7uShUDT7KpNUfcTZt5Fn/YdpEaphDn5OJxmPZOkcUbz7RwMnhGxNJ+c7XPU/6jVs+3h
ZrY/ap0oIZbiTB2Dg8442aZlzOGqi1uRsLLTBUh2NPPYdipmkfkTQnsjxjFIzhsVF+UIVEVyGl0Y
b+hO3VrT/l7qKU+3af/feQCyKOp83YE88l4mLKu1CjBJnZBbKq8kSYYZlnAXlr6KOjUvM/MhQjP/
meeo6WrUZUN6wD0Tp4dpdiM3+CNg6JGFIdEeKrBLZ3DKnn34K+3vwhgFJbH/cMNnj2x+cCzpLGyj
1v1w6xDafbHpYT2oAC98537jKCur1zSmNcYTXZcKQNsWBDjbH4jJ3MSNhhQ2PGMTxu7pTOQVb+Mv
CYie2gPQP7JVcBVG90uXvNHffOK7M9J0UUYcamZvOE1v4khSSgmkOBjWWzdJkFGGWjxCY5e0ia43
cZ+fjXyDynrNMsrvUVwpDc5ABiOUW5vE+BG9+MtSLCbf/yFRWH2OeWCHz6pASZcyEJ7vlBLpPCwJ
A3f/DQvz1uFGN8b6HmBQhiBH6HBWqDi6BA3n60PguSnUq6ei3WSHf+JeeUn1C6lMLHuiN/g0xFu2
/Dx1myd1lPsv31a9xYcPTCa0WH6/HizGXJhcJ4iBOva2rA2aU3/0AzKDPiHmO43a62Db/k+cXKGv
ySpFl4Y/iCXw4J3erhO00afbD3QiY7UvViBZ+S+hoAWVDZgQQSJPaSq7UTZWcWdqQn+wMd1o3s8v
P6QzNLpViY/g0AVPmgYMjQAxz7I8RqeUb4RMfUZ/kn4DD6dbiNQajL5wcOfeU0SCGAlU+i9mtuL4
LBbwquNnm9K2CUr4GNqES0E/piPuyZBzegmhs9LGNUhDWA3hyyZ/oWXmAwebX5R0lhuUJ5HdlOlJ
UmEvMw+pbMBJCV72n3HeC7aK/KyfcYJ1jm1Aa2j4flK+EiRaEnCaHc5ZhkoZTpqDHjyC/m9dWY+S
d3WrT4hJEGa1idJY2ZmD+3N92sxtKAxzH7I44ItXHONSvVaX/PmG6AvRwsNatV2Q0XV+UHyLStTc
An1FEkAltpXgbchBpKxOWeMS9ZU1huNZQ8xTbH/FTBE3YyCGUFN+oVXRUF+VPN8fZoxDX9WG3voc
TXMoiiQlt8fhLh6HX2vdcF1jh82XltAzTdO5voqopKxrQ+UiOy+TpkqLTCBSG8RIqiChmBq5QyYU
RcuDGJ5W8X7iiCi06xUfOu/Tny89PKkjN7tFAJCNMy9+YA9by/66miVnWKwOQSyuIl6yVHTm1Rs8
fPFADw9Yd7hgQ5gHyezsib6VBFIOpZqisWHxcjO4yoCcIELXuGo+P6S4BuKDRiMXQezZFvmArr3z
Z7QPzBWs+Qaqkkv1M7ONrSx3lBQVX6BDTOikwz6oH3d/HOBkxCv21rIBJIBGs2Zqgs28LpwH+NvU
5sVZsi5Yy8LKcYcr2bQo4hqVCPAhUu9GQU7fje2cVw+2NNYs9YVr/3Ma0CuHESZMSsKGa5eRaMnn
7qKtjcWP2CagkvZMirPwCgSqkqul7qC/wLJ1cHZqoW6No7LAvu/DU8YEo0beR2qUkXP/FW0COQBh
D2HIc08sY96uFZxmeBBQYcINOfX735w0gumIjp4jGPHZ/TJ0E8dEMRkVqa5LjTJ0Q/Rf8Z8/O9k9
k6RdaMYfxTdlPeRMn9/3DqYph4S8T8Cl9phcrbs8EkuTxDhLuFbrlHbeQOhhOEbbAxhz6DlBuori
kc9K+QlLjScjnOB2kL+kk1Cbg3nNtQC/T48FJx9x/fNce+hSAF6Okh3qp0zKjUFbOCN6K0HVBrT3
ZJJs4WApsO9VhSuvbbPYjymtgQokpouU6boFUGy4+QVShe+P78roPA248F0qjMg6kPaTIPEGl6Sm
I4GNt77uY3wpC+ij84Rd+aNeQ220LByJWkR1rEyP+YjvYodrY71/jYXRCQpU6XU0pJ3J4qpyd0zO
2Eyq/CYt3TTViFC6Sln1xIMD0qCWOgrT9g7Sja5lz5sixSHgn5Phr7QT7JGjqVQ04IhP+64ypZnF
sHhUA+0KJDmMEm8ZC3N+eIs/mqpiYLYGXgGP7XgavVgfufOjMaOxGgklUdgqBGoDO1Jva5WQ4vw+
G3xHeRg45WpkT2+USrX99jbZ0KKeK+CeTcVRv3ENEu/qoI7x4nVcvstqvhmhs9GPBaT/Gwu/ANvF
0awKphK2+0m354jdmkudDsG/R2TVZFHBFdNE8YdkyTS8KODnOId3w1MsxQ1uQj9+9s/2GLYUFUdn
5nYQgpmlhDZJYGjxKARNq+SvRQ1NUPP5CkgRHNlv1dLIp2jA4XtytwQgrjVHQ85cs/7yhIbmBiyU
Cu3+RMaHJBSRi6GrUXY/ILSZ/H7A7icM2enGmJrIXlECeHfsAI+Mad0EgTUxi/nF1iNHdoMDXhle
nQmRel3yY2CsevtoRy85CvrCY6oxlVmF99HmHv/hA8ctptHcwAwPARdq5/xpvAd9Nsh9A8+fbeaL
9YVfJyIzWog+5NbtJ+PTa3YyH18LWhjhoJgLnFQAunRIfhocaca6WHt1z9cdaj7Tv0Pg9OfUcBMQ
Ps26hYYLrOO8sfIvsFPZxdzkdQvj0n5NQlPtd1li0QODTUm2GDNIXRFKtmh8n8Ea0/1rLCr50M8L
ogvGsavB4CDXBDNR2IYYx55UWSKgyf8fi7VXY24Z/E6d8KTHviRht8U64uDZjEMN608rHs730bDL
iiiAPHOVNvFp6BQLgUcaDZ6mMXisBFrPk/v3JCWmyzMsbKuqCsg9Ufbdm/RUA3QFpnc+XVQTFmFZ
lSozPMJVhoqWwacQ4L7gLxaUI2t8ECr7FWjFTTlZJVSxYBEySYiFSig3HWRrny51wrnvIBgT5CIx
LgtyUfDDJtISBxoISDwvoQ1A5xxkQGSj4iasdeDQA5Qe9pAZ23YsEyX9itISK1iSgKT/mLAToHyI
H5/BfIfHUZf/6M/4TXwgmLtzITkgbS2ytKnXdnBiPWYNOBK4urMHg7yNDAjRBL/prI2caD8E+zPH
VZ/N9HTpCRFMUacwNJzgEba/WnBc/TCAsFr0UcncPOR1ZzZDmAbmqBM0DCWGNu/06MQAbdxXkEwq
psbmKlLFv9lnL8AT9s84X5jzfMlXdvT6cdhRhtIm8kr7qQWek3VolKvaoMDUOOcR8UAKM9LVYscB
pB/MmZvzE82N7Bnd2vCT8SEqdE/FxdCyFhrkktgBDxz5TUyZuPq0vJcXrpnMeYGn16QsIDI4zrZs
HyCJ95WZkKUa9OADh7PQuRBOGYlu2TGP7bi5ci1yP2XoiozbD9G1BCmyq5Mgh1pTNmdwAnOoTm5N
FY1+e6BE6mtB3hetbGBvSdmews15M3LW47zeA4YRzGL+ijPy1CgXSs6dDHwa0YnMp3ok76FNI3Uh
N9C6s/ocqxzqQ2HjAdBjCpMOIdZK4X+Vcz/6wkIZ3umQCEbyhSiX+kqgWpd4GOuf+URFpGDnk/mX
rCCDedmsZqY03X4f8D4/gPHBG1AyCFsquXj7lXldfWfWeff6omdZ9MEc1O4bI8fHjBjFMyvBEVTW
S1+zgGO5pQU/rzBx1XItfYQfpv5hAUL+uz302ks7xfYPaLNY3LQzqGbTKhVsun6PQNUs/PorhVO8
g9iau0YqCTHmyCgs5gFBnbaoy2BVtXOVfenwlb3Gt+jEo6Dui+JvE61khNWR7mVgMW11nyg6wcki
xvgrSJqgIJ5rHCZOeYQZzN8VSYzzIA5P5+SQpQ/sSvFoKYLf+KiYISSX5JMytqVrfWIjCcM8z4zf
J0Lp67BJwxkF+K4HYQhVmx/3DGl4a4XJH7zV2Zz4yMVi9wZsQlzAxXhYRTbAGiS8t+5uGGGLTRjq
lrvH1OEEIotFjl95gykJDaHYF2gOZb9Czr+d0e4D6IYojK8TYmLqblINnvGrP8MCY/RZ+FAiR5fp
WS+tk6AuudyFBDhXk5ouxtD4XrbVnJObDBxi6CLRDXd6YMPmMHKqru77593FHNseEZEH07XpbPcE
9gUvmZMJ0CUqI2nigmAyawHPXtMQbEdbjcHajDG10pC4i7qax7kVqWZwZFjR2AM9xm7QUtSrD8an
/h8bT3B7u3dp+WZas+6N/68jD8N+Enz+UsMxZatOx8Ffk6l+sNtK4iQyQQIDkpKwPqu6TjAwnmtv
TvqpiqzYXQ1tf9crwmMhi1iCnd5EEfsgZW+4eGwI5+qV60AMy1h5d6q4ZBd3gEztGvfjzW8NZGam
+Em736HyJS50Xvx9TgsdEZbAIXq0gc8gzSWih5XxwGUvma3Pm3BqlCuxhcEQyGTpTjScfvfitHFs
m8s4u4DAVeq0rKYBEFBcTYn+wOml8pjudPPQDy6IabsjgO7offxeP8IowRO6iIyBG8i8TjDxX1jL
v+8lDfOBJtu8r2MxbvI2dhbwEoArefSG53j4FafesqV1R5zrU98cOsUu/r6GB57UDNvX7CWJm/AZ
XSouu63883v2azWrG6YH912SIuY9oFW6Qq3yxcjxdUAnH74M1n46Ur53pQQ6D0J2wpXKRjmzlibu
FyIV23OWQvayUhNFexTWX6aUnTb2HeuF0UxslEcJRKFgIjIytGtOMKtmFcEt4VNpBaNO85yOe0eu
GDWepYw3ci1SHQL9pND3w6XlgPIKlJ27tfj1I4E/dZr+MO5uuB20gzTSqbi+k8FAWtaQzei8kDJ2
S69nRqHtF8CHwO2NtexxA/TsRIKnKSzV5eXsAEVPQ9+Ib9L6lufUhVl3u+/gqz2RQmrt6H+PJHhh
zEjSCbQA2AO1Rr5xhmV1AWn4Q8zJzY86ELuoFntSNZJZZ8mAlAOYO3OEDMIJo7C7jr9LN9QlUDNq
6So+MWEYmgVdkatZJEYd+eZqm+z1HpgoIsWAuGlPCEhA6SMXTbsLEgIX8LW6RGoj7AxMKgect5gC
RxYlscLTLEFXK4lBALlXJfBiAy4R3RKTPv7QLxPmhRlKcdmZlUCQ7gkmEkD6Lufp4qMHsaL617c7
m2Dke2O7FsopX/PYR9Z1sdjgUr5qVskVqCcVNGbqE2Y3LWz/e+50GgIN4UI9fazfb3cSuKcXljFw
SXFRdjJchmQ//0JklhT9y4tNzqic3o4jpzlNhhrM4aykUJkh5k/Jezx2qIjAVmmegTIGjFlWke+t
FMy28KtIsXXNOeEH7OGRdw9Wo1tmdC0t5Rt6b0oU4XmtZKFzEUgQoQd8DMAino7IZiF+3HJZ5sNm
PsQL39/QW95QHrwJBSOOSsjuRH5BLOsGH3Yc3XZIiqMOhjQ6AEuXKFpJWQwRXFTexRmZHd+L+9ml
tOXr9IN17iY9WllEF73tpmbqj+h5N1Wwy/biw12OyT/DnT2i9qSiIeiP7mO/k+1hqFg9SGjv6yMF
d899RBZSaDX6upAcIBv5DcryyaxRIDtdu7VEc2cPtnqSwqhdPGQm1eyvn89HVJLNKO+OncCDHftJ
4Yw2yoR0bQ1jbCEFKHZ58U/slPk4ZznFYR8CHJyiYAzaaTpmJJS3AmPzFfnvzME2Iv1NCaNwQb7n
YN0PtxH6kNKJo4PzM/sbtHyjsccKVIiacZ0jJbbgePTKydRDUshOks13AL6XKbCyuXvYZ14ruVn6
VEIRtavsQ9AP2ThyV6u2J7sPGkwGOgpURLSiXNyMQnDNzdadfX4ri44O/dW3TlP/aCvuSGwm6Neh
+Bbv7Ms8laTV6TWYUA616MpohVEom4osJjcMD8kPPEzTgs7nDt6mZcFeHlMwGqpRgDWSmaJoAqgC
3PT22VNFtRBKcJQpMBJ94+Qwc/DDE+irGpIDv4ex+vZyuqFaNZ8cAHfBeDmm31TSsydG35Z0beRF
yGk9rcyc0p08t9AP8FuWjoBa9eedS9hsZokKcwvm9B19PCxGXUjU1p06byA/HIM/0mv+wbotU15S
Py2OhcH2dzoJwRpvE5HyyLDMpYEVnYaydNlsTfitPDA6JrH2NXZIBaVScBsxamMZxWNEdkPIyCDS
npd2Krxagmf6CoIESEV/Dg5OVF9Ig4YUYhkvLqTVHuEhT4L3Q7wRWqFf1UeUmBGFVpKbqIFze2wG
KutogQCz+B7oEDy+EVPbYcY/0CWfvUsHMXn6b+/o1LYQxz9ZXtLNGoQ0OfVGRSt8wVaZtxGTCrfM
wtzsiS9D3pinaXgXx0IG8kiQo04dAvtQjugrPjtoW29iqL8ZVMFALV0Zzh2Y6Nsq47jAnfKaoXGI
PnOBHgcb9xDxiXtyeMxznk9wLq4GABv5uXA9QsIePOTbegtckzd2IlB94wFsS7goyekrFudch0fp
SQ1zSpMz9mvkJTlLPpRArq/GCklpDOjGZ2i3jTd7RVlwtdcuMj4uOWn7J90wSp+mSsli2zeM5zYZ
6ok33c4WPCH9s17V2qA3ork84JYey9zc2Feu/MvG3oQ+YV/u18LXZ986iwv3z0hMEY2ztngW74v7
9GPwLT2Rrj+pFZ+e7mIeYlP6PbJvs/nGUTlqYwCsM6wQvMKPJOZViKnadFASp7Ki7O304Oz0hvZO
Xv4DF76PMqLGRBFGB/bqLo35h+XKAFrVlBwNCCvbcCIWiTS2TofBD38CF/GPAIX+LMxG3kTv0sVC
LgKg6GhF27B3hpAPwAbnQzE9sRwe5qb4KOExQX9OzRoFV+kBoUtFLNRDlht3YNhuLwfftE9lN1hJ
Cl5+xsJ15zfJoz7CbFQYoIBnv1bF62NvAJU82dOssPsONCRw9iJGU3zJsjsFT2lMHMxTGyb+cG5m
63pvwF0V9aZsePAX/7cb+7NdZ/g+9+TYx8/4+O0NgIgPQfMcYttfw+PmUj0ZVL765DCwGQQYlvoY
SeXhWHkDh07NjwIaC2mi0rF5V5M9thfOghdN9QcTpL9eEd4hJiSR3an/0SB5qmLD+9RGrsAS0wOf
7oAISMmCdEVTVxcRj5MzFTqjN8XShVo9uIKyZJhAQN685/xY0R7GSw4LzsMlKpa/6bZKSLF2gf0G
6fu7rUpFdzx57qJciSFN7FYufCkjIS9V7y50H9sBWn1FsTjea52MQK8EEvEdKeMQQ4cafh7IQXXa
ub8IPe4HqM5KjRi4Uz24XYlGIHariPgZSXSohBdPx8osfFR1liwVRAGfZYurVkUlcHd+yMODdCF0
OoYTAUt91R2Ufh3ndaTv9kvqVWxafsogeFvEl//3QtagoqPomElIInEDbWasH36XfS4iFseH+Lfj
ZaYCy1FFain+XmdkWK6TChdwfSP/FfmcT41lh24aBgO6DxKZEMTpQzB3FaT1z8ZYerxZqgRTQgpO
mqipnbyhq4ueHR8ybYBl1vkCUo2S3OxGpxJPDGWuq7dczFyPV/meFlw2h49aA4rbOIf4g8pt0oXY
Y2YbZTV0usrhVv+KVsDb+9aqbVtJDYNHewjWp7NzFBbdrD8RW0h8Lo6XmM/CAMTAlAv47scDG8Vh
MtaAm68QydO6FUtnZOJwoB9ceR/6gtMOd3unNskmw8md3nj0lzZjoRQr31cJMWxF/FXxnwyw7N6v
WZPta4tyeykoZrEFs1mEAhz8KknthpxhHGbquf8oZanR40aV2k+wSr/RXQk0pPPNhqL11iI2qx/u
Y7i9v+YQUPRCRlVqgwJaOr0ZB1+S8pu+cjAWwX2FVW9ifi+VNYY1sxXvCmTGzp0Izg91chCDfmGt
C2D/a0t18zoZbmCOC8mhWVPdDrzOyfqiKoqkL4HFivxPwAW891g303l2Ub4lMkU2G6+pUEGUO2fx
gRjr4GxWO1dnuQOTAQUkyjyP5lud+456+ieZ0uxWGwq7uLSM9fjDRaw9FUN3Gm0Kw2DgWFujnEq0
x4Kl+NU+Vds2VllLEQoy2ttFelLEX/4YIGwnn/OU8kTv3H5P6DMoPEtDJuU8tC6V2QmwDSTHMqGY
fL6Lv6xaVenN0Jh/9HPZCbmn9aDXiZAOjDncDRSGJoTiyFbf0P/c5Qxbjtgu+4QXSOfpUgcgA3/t
jqXf2pVPfMop/DFcjPVTAFSbixnMfkkrw4I+rKJicw9PkE6+propn+LH50fx3jlJV25hDSWlc6P8
3BsYy/gLkioIRdCdShvBU6Y9K0wP3pzcfUPZAI6oV0VGgFFJIhQcK2vUlaUeIMqhtsAce0xtyyd+
moeL+0cS4e1Ilj/bpgpRJ382rlSIE83RxivFRcNHx2wXZD0IifKga0REgOmVL8qZk+n5yA7kRadD
SHrRSHWBeLlESvjITGRLTaEDD4XBtQMqceQyimeIaJhy3H1wAih7MAzWFW/6TqcbqeKrXhp0mZGk
P7FUdbU9ASlwb/TLatu8JQxUsk4vS4eV7OLfvHMwvdlzJU/ozGy2ffF6YU7s91TWNfcOhxXuPCYX
NtrXgdAuVuL63BJpJSQT7+mpyM/h0HkgbpX5I1WLacmmKwF6QqTeZfXHnguIpuFu6oEZS0GwKLqD
q2PNwrOgJNqPBiNWhKaMwcsoS/2htmKJWofIuGDDJ7xk7PWg2aSAlIDcs731y4WNYtzQKtF6fd0y
m1WF9IGOW3y3Ca++XOi0Huasgv0+ZhfjfjLTRoeh8A/rGI9LgIa5CHDD/tDDnFodeftJwMFSZmvJ
6+yx2yVyITI/ntcpyO3JTVbnCybv8WM6x9jZTaFGshYgDQaqDukf0W2fInzGIY9yTUAN1ZWwD2PQ
RHYIhjtfAwyXnsrIRtvbTnw/aQDgZ3nK6lICMnWH6pQ///VtRHLC0oqu4OrtL6MMGidXOaDiTdQ5
zDQd3uuJOZ64BCYb/jnrVVX2ikJ7arcGC06aJRzfhlHm/foMET+4IzcELgo/RrOnhRD0GUWHAzmS
pbAs6O44gTQlsZ2o0OAVCB2FodTfdWRTtgNfhbYZ4nd26i68EvD2wL+6/IafuAKoSPa+x+ZAYpYH
5z2uGFjx0zJ5AJXQYnCLHzlZkzKghavQHr8z2jVagcz2uVCsuE9uqwImaDHry+DeQFT0plgFzDmZ
dNVhtj11WkxRKYYDf9racwLtE86Vo4glWgu+cg+FrukM3d6xejpnv7Q0+yTuT1xij7mNdp77kzQL
5GJaKHNRojyV07MOFYY2oIxlICTkrF0VykPQ6Fi4PPfUPy3bcl6smRPIQIB9Whx9S8hWearnXZNO
1dtDPU9HipzLnEoXJMgBcwwqMCIzW4J1lVvTiHQnoUA1uzdg7sZKrWYTqe1uNVFECfuE/3tXmacD
mKLN4rd+O3a2cifmUra6POygxcGqRxgcDMZSY83sav+K6Z7WWu06/9q28L3551yTAwKQv2GsfYvp
0QvkST94oV+rlXNty0DJ9ZxE4EVqwkUacMQL4qFCreQ4QV/n6k/j8CqrRWrHTyNF8ZDFHtwuTVnP
WvFFA3h+6ZQb+th/9E1a931dDeXh7E5Nt6LzKadp73w5JcPxbo2f1lHznk+GRy3uVseK/OcQdz2G
W2pO3od8FsflkOTUEPdFqx5CS++Bg1QnC5rmS44Fp9N4s6+CE6styFWHDNwx/+EgSjYD9q6qK4MU
xDEg8yHTKLE2uvDOZ8htn5/4jBqWLl1Hn0TrSJf718ofAiehofQl75dZUhuJlq92npcrB83q6kac
g2gTK70MnYTnnMUN5gc7vfGhTLbzo50WrOH/713eNcDfWxejwlu9c90yagAQKWvBYheYdqR7Ao/a
DCAMwi0SMMwfQyFYwFMU2Rtkm6cxwLtfSXPGQUwNi6rpGSGLMtOGOWE6s9Jk7vN7MgdC714ZnXx9
3Im1GQrbShQmRlydFKAclFAeSS1Ty5Npe23cuchbctudzn+k9yJES6o9VvgQwmSC8WCkUzgLqkC8
p+lDFsJAnr05T0hPuryYZ6tU+tvj2YCGFTvubh7dDRBrJ8vR3BMohsnMGp+Eg56+lTmS5vTH9nYX
U+VlR4/K8dguI9m33wWmBvfhEJkAVI7sfkbGlYX8cDsQZgUhKdcsc7715tzNUiRbKlq9mQUsR4K7
5vgaZOtyfF4r94is4Rol+fk2e2M1lQd9RbMU6but/M+3B+w7/KimXjMe9uhdbSBwfF3ktKaKFquY
FqF841QVclX3vtrGJFBLpJsajHbg0ucfRfnvFTCeF7uK+TqJMfKV/QlJNkL4RtK6Z91XNxYwzgUv
u8iKeKhXFh6c2eqPnb72wUdjKXO498owKvQyEXQZyk6QeehoPQJt/lh6pHHgrFsQXZk/A5CgfwRM
T8oF+RO9Dplho9S9CuGWJirftLChpLZC8nEiXi2kyZJofYdey2aOOoBJV6ndaPBBQeWbhlyryaKD
cFUhYGfK8fKVlrvuiTcDJ8E80VhSmt+Gjd/EVe1eAQvAvKMZ9Ca5hzu5DtqxYA59BVnF0qha5dm9
+VtOfwe3BFQjfob56Mx0xQDOI6G3oI26TzsrswxXy9Kz+zd1pruYraqYjj7uBJNeu9CfD5gfDOrJ
UELV8Fps3ZAK7UXyEWsDez36kZbOkmi91kNEgXoNM6tmZ4YoPcmnNqAyOvByl2L25XOPxLGeQv61
dwPG6g5RHYWM1m82mFlME229wLrFP8sS13cnmDaqfvdMY9O9HtmLGAD17J5lkAUc+p+L1IUjZR09
KUfG/aeLcvU4Qj/okSMp8UKdJxEt1BcWn01QCKWegZvOHYeWA+FvZDuyjshu2Xu8qCJzEild3F+m
hEL4V+bGpGC7k4e2o4nYOhxReg73zOvCfosnPPD3ZPdcYHxd5P/aEIgvBVntcFVo0rGqnjVNl184
t9sk0QjBZTGbkppevJDvaeQJhAjoMJ4UsXZ01cDEYwKlYWYQdYshrCvZOppJJyLScdZssPYsHqyV
1btA4BREwFvNr9GE9SuvpWbrQHnLqrmCO7FE8PjiuCMfeN4XZu8M5A95Yoc6NF5IPXT/VEX7T9ki
yJb9rfC1XRvsTikXMXR7UJMyM/v/ib9fo01bGtR8StfONC6jwKXxHxZ6DmpG/N30zCViQDgFm9vY
lQOsRqRtHr1J+HMw1f3/ONvgkhOo996/bc3A2XlZ9X+Elxwzn0VGVTznxLqvHrjmfYOBIk0i7EFt
/pl6GixbxCDxoWPIYafmLSjfy08JZy7cASKa77LNJqvvFKPGKMDnCRoayz5if61nXnerMzh/fSzj
lFBxglk7JhDyrECHPRqk657XdZUGYRFgGy8cKw/SJKVUTk6bnVAPR9NWriLAAGzCPeLqDlD1ja8g
7DrXU4j+Y2zFmtIg/zbPlJLjMfbS20KD+2uV3JN+po5nF+X7YaEVLDQ5ZWqOyk5AuNX8jXgzFut/
7vBRzBuNbfmAanaGZExI750v0sz+TxPgHwJQ06LHxLoZXcIGDfEgAvlJ1Wq84l1wpLiYDz0lMWP7
L7OoHFkXEe3CNQfGj5U86fuPs7ctNEad4k7dJJiwhj1bmGMC83MBPOirsZuh8hptSVI//lHYMR/Q
2SdLC2KAd/cTOn1ffyaDP471QTPmRwQ7e9VPvT9FOLNXtawdT47GkuGDQ0s0zdIzvRsqfPxdchrl
nkvgpPlczJ1tsOshZLGu3vuEYkGBzPKeSBN4guWD6qhU9fqFc14FwaIvPp/AxZ+Ad3xOKWA9qjD3
JD2Hg0gDmCV0nK8Lzk3ETIPkd64DHEO5vhpT6uWuGhdVeWGx4H5LwdaRUygZnkpyqYEWmAqa1qN7
yYIjlqQQLiP/fCdN5+bPP3YzXPn0BC3VD89HKiGFjRlECBWP7pOY7Xr09EzyOgPR3QI3ntJJOhlG
KYIoM8FxnVstTptpXMfzy1Ivwz40t5+cS4yokzLZHzDIxC7LasSpB5JwIHkCYIVsyR+1gDVS2c2L
4nx1jylUPTIruDoVfqrdrofC2rkixDYvQFNZNf/r5ZvZLz5MMXnW513sli6qrZwAj4MpbZQYefMH
RLYTuAzn7u6TfT34IJxDPayxzX6syL9a/fYSqhsYj09Ad+05xIMneZbwxMQFAhtTOlL2+DpvFxH3
br5q+Q1sWBZEs4rbmYdRyR89WJTgR+dIBHwuG+TNxmfsUg67Sr63i5cRQpj7mqDF1AkSi2MOPS8a
zBTEkZ4p4xZp0acoQXLDE2tFCP8zznDklKURwWjslk0GWkpiYn3wYB2nVBn1DvuTDRZFRUHsl03G
uUDck2w27E4d1VizJiULudwVexpdGZyllJTfCW5kBjLtBOfIbZgpGfi/VJzVxjzsqCDtCvSEqsqd
Kayp7w0GgCbr7CZuki92o6zOF2ALJJxvB1lERFoIEjLoA2ZeKEUl9/Ry843flPLlJdsct+uFLpEd
Ujo+O22A8HQyOiQC4HkTyRzJNf6ewv7gahMihPPHChvyhXCDCpHm/UCLXxHCf1t2g1aM5OvxcxoM
JpQxfZtHqCP4Yzrp1ouONhmTJZ+ZJQnd+drnqzjZ/caSgDAaciTQu8MAMFb+n8j/bLGRBFbflhf9
GYIDFHg7nN/1c5WfMWt36XBTPPEDAVNqcWgT5xsFROaq8bqVAJgVrGP78dJlmJjohPtSe8OGway1
NLY5BcgJjhb1uQaQOb6Yf1WPn5GoQMNW/R1s3HzBDvQ2WOe0mdpn43BxK3/gODOm7UNCK07Sfya5
8PVE/syVv2GeFQK3pfZCXm115RGaGzcA++AkAjiYL39r35waLuG0sqZxMdSEO8DJZJYkXywYttVD
zRBhXgPIS/VlnDchOkfUeccHXIh4zG72aJpaiDQpUHIuR8t9Mi6z5JVWTkt1Z2XlUjbTBc3fjSNl
daa/vmFEgRmCRbdvLY6rtBHL2Lw7ixRm2HSmh2e/TimsxCVN5C2Vey88PUjPV05GX7yJsejLaQKr
GsU1j2egIx4tpDsZESGCJUB+QT+BJN5YrYW74J87Z0dreQNBqMiQz1D2sQINBaZqKfeO92cKpVNM
OzGwmEkw5bFmZJ6bM7Zc1QgTCgtsvTX8dD8WQuS+LqjPMAA2h0MbF4rVL7R3K68oxr0pzmKXHXaS
Un7byUL7hIwIWwN0z/LWFKvBcr8EAFYcmgPAmd1fq3cZ6ivkmp0D6FizZ0yggR1No5ql+RNYabCO
qyqI1PAnHd8yLzg47Q6eM+wGZ5VK8s9zXsi6wMRLs9o/KDOSYGzyVV1Xf9ZNWeAYknXmeyJqKIZN
nUYvn1cliTg73SF+r2J1C9qUvoiXRHSfMlKKTGoaEkH52aNOlxG98T5EIwAekyQLuWyHJntj4Epp
7sZ5k5Ur6W/4Gy4vFDPOc0cm2KbpnCtV8eI6m284EZwg8qJwC++bl0GtILpi9OlM4GOp6Qd0HuvJ
Me+ArCT5UKy/lHZG1sqBdZIPBclIz8w8IVsS6oG1KB+2mTV8JLnPW2iB6P2XoYfPEEcTTLkp16Gk
JiyzSBVX5Phdzhcgi5ShONbJafRxmac8EdPlusFB3WG1Lzhe7g8XFWroMin1gTM/zxkE2wb/Zm00
f4yKTIClkS9C9tr95yWnZs4zw/jhJCFExxsMf+60qfhGbWFTMrNawlYgI0jIeU4FFeO62cnLlTEQ
7ae98OBEr+ua78pikvkxJKkanMLpXF1rdrsv5VyBnaER8eqWF/TR453RzEuzr93qQ6WtYgIBpLL3
YQjTyRvICNKPTa0xX+BRN/C1USl7SeQGQhDcRNxNPCVb1v+g1pzZ511b2w35mrXSKMtE9n9Oj0Fy
wVx9hEVgf3KMGatNP4IyqtBvYZn4GP/uqX+JdIQhGCgOExPvc8BGfzPCgm9RFB8uypjEJaCf0wCy
tx5Ox6DdM5yoKrjdFNkpPiDvuIHrPyJcA2Vdtoz0hgBzXIY4drBbK6jtsEWo9hJ+GSC1ZFR6SF6X
9zlDIFk5OJv5v4usvmwPgXlCE/yi8lOEWStzwt9zbXt+dhnqSdwlnERXd+i3v5Q5bWB+iJyLtlvb
DOo+4SIPyZRCdElq1Hjol1YTMM3TDN8tIcFSBgLB7zgloX3OWPIlrajGQQvc/0awVZ65CZCYLAQ0
TU5ARz7H5Ua76xPTE2s9ve4cCKFB7Yfzhr049H87umv2l530HpgA8rZUIVEswzLcTipi51+A836N
pWbFp20tjSC+VcU4gACIvj7B8cS8i/U01+X56vpsUljx1skFtQsftDefJ+ETbXslnqfxkZKgXljc
3hCIC1GRvbyYxxIGWO79dh0d6DJ9XjZw+paRoUZqF5d5ClZ2xxNKANDBJhd9nNGm81lyOSk5OP75
xfhvo/dwmeXNlHY4ouLUtv6Fm1TD3yKw60NXZC6dYav3w5Wd4T3QLw3oEfaHhcJzzfNHpRJaElKb
6JNZ4DQVJuWn+ChZjPBJdVB7MfRAJXLJuJgM/YHbC+jOxCAgylOFKZ85QUhKlHqX6hVmRUBmkYsa
+z27tX1LSUzyy8at+s6wUAsdWtyfNB5Nzo8rFa8FB0DVDU5yzMQVSDVrPC9rrhZlWAepd3SuydcY
LQzziXciAXjf2CSertTOK0IYAUhdPKSWo1v2aY2RZgDw7hPOnZdKOn250PIHyzm654jZQzZLJLOV
btNTRmTXZZPAnQbulxwbtAbZ5taaLUSMBG3UxwEHkGErGq08l+R8CqD/Xm1q8X0u6ny6jmExrn7d
+vqImLlUKtOWT3mn4Vl4aDVs58gXhh6/U1Ea4JCFWI9C6+2tE/RnOBDoEQdwe4VDWmCTL0Yls6o5
ysLC92cQ9PLIpdHTIt5iFZpgxbfO62kqKdbx6UrMpCPoe5nPppcJN7JbWNB+g/Vtxviy+hcrLtWE
TNHrIO2L9GoPRP6U1DkKYnipuIcM0Lo82SmWrrBRPn0Utq6VyswZA4lYYvQ5NA0nfwKmCiN9MeCV
L7Dur1/OG7cwGYt0lNCRIwIzmcE+6M4s33/xKqL82+BL2k7DDGLsFwPpXPQyHsPmV9XzHuxTu5Ft
adhpBjS6sK8RGMw/44Chnmw0OPUSkI1cQ4PNDG2AiaeloU4863AuWCt240U9HOdCNEqKOUKVbE34
CPNkWZfmYKBaT75RTq7B9LzcOuuv7wWmZRAEPEduHG3HWYfX1I/G+Gy44I9nk97yHLbelvd1ZmkY
lqvfhTHahlePRcaRcKwC9d73B8odYPERiAc8EgoshftY/wewgWSkbfW/QdZ4Y1RK8jfOjylBCkNr
7hTiUGXB+NmDurBg6d4CAH6JzFPc0Ok26heuY3W6xs5mL2X5Ctzpl4LTK8ZOIOfLfst8/FsN7Vvx
Wk0nD9fV9rw+MNaE4YgeD80wV2rcYHGH/hvRPaeaMXI4Wf5+RpqAfuhHcNGYIWOm62KQopEspZzg
k3shrNhnoxvgPgg4Vdd0vsyYFay8mK64MvLUd0W6mZUAtu9WJJ3RHqf3rnS7+D5FTuYHiwZjTyzY
DlhQVP0NxoIQcmIlnqstCR6OQFmf7HhHrALQOxRq3ZCo6G6pZOnhQ0MjWm/JYvTjL4yYqsbDjNCm
+rEL5ZHo4EtfBqQtGnjg1dANpUxLLWw+WU3ehSxylNDOu9dlQIr0Sk0ZCrIphQaXMZHLbOR1krit
8y9oZ1ITgjuxAg9kL2tUewWM6kB/74Y/Rf1IyIebTTW2/lvm4PBDqNqLkI/IvVITBceuqP799Npd
xwhFMZyWa2ELz8xHyQzUFDceStNMKaN1gVKk6dHh3AYWpYlbyXjYJXiqtx85GE04FQ1920KNKUsj
wLH9EziEBjbS7ZV+AtEdOwU6nZEAkuJMmwT/ecBxXIQZQ+EVrM6yvSTMIENtjb6AfVxNJE5ccvZ9
9RJXABaNWhNwM7G0EQ7R6mBwxbDsr2A1jAvGL/5mCa6IJ6JI4l1NAxewdeUOIJV8cY/G+oJHDNMN
eBHfQ9wibh88w17OEoD1JlstwKQcY9yPBevSj6SlN7NEJjmlPQuIwOG1jKKY6ecKfLMjBhHeEGpZ
/J04Q+uPxJ0zNQK3sSXyHOcx37w4TU3v7tJDyvV1VgwXCkBAS+L0Vm+m5RzN740pHrEnL2ShUWzw
ewBEFCE4kywrvG5d5Z/NFr1a3uifdhG8ilc2MnuVTjpDSwbvyAms1I0eX8kSEZggrp09cHWWaM10
/boQymzuxfZDF/hmEMqPz7uQZ2CmFBnzWVU1yUdc13iDiWezflpQF5krGHN0p1WIBk884OFNCzYk
Z1bXUZLjpzbDOJy1TgkK5feTpNB0YY7xTd16w8RlozmDJ+czLSLyzux+7uBFD1oJh3ctTr0D4CMj
3TS+u6RKKHPmk1TmIQmwAhzSyXcWqhUd2X8Hrn2OWnRqrElORRBWnKAwBMJYgBIwNjRScxSniapj
yF6UZEyiJTLjh+OrOGk7ZvTR0fOe6CEr9Nsk4kyykV7ddYFQCXRZJlxojT1c18Su/x+ngEqUgli8
F/iDPrHl0yBf0POeUQ57FKLThV9WR8smzm7XjhOQ53l0hT4nuQLbsmsp3LJQzeND4rpl3e0lLD0+
Sf/loW30om0CZsIblgkh2mc9reboX6b2/vI6RUjfA9GsPcnE6Op5qeYffhxP1+fLqntaoPBw3dWI
t/tRc6oD1DlHuE9sJpCHTfoj1Zu6WFjLTBh8OOZZU2RW1ibQQSlJt8G/12lULZSTBG1MwFZxN/ts
8bfsZP2dRLoMpvKmTNxr8PNfEnP5alNLfoFP5WCoKmlz/yQJy/606UeGuWS49lXl8P3b0YBXXhKd
1EYfJjz8D0cr2MkXwtjC080NbCPp5fQwmE8Om3Nzo1mqdHGhdXpywxtVlukzcI0YDWvkPm9iLxrX
MU1S8+0ZhhuBE2XXnwnJXJN0vfYeOSgQ5MHkPx+4B5IuMI2BYcs3dI3IX6FYnHBGDwAeGov6OtJF
0GCM7hBZ0Mbp7mJq7yTkeJcussQ1mYekRQ0jVtjX8I4HQjzWtGDDyiDuKF0f4Ioj7z2pk1QiZFsm
Xmw+NZM5Q5TlDHbPsMOEKTIoPUM+wp4CjiofQ8G5+Ocb0ydlRcz5myzA8PGPTojt1IPid9PsauGG
njQxRIgoDkvPju7liBqFgJXU2danxQEEWa4rKxFlqUBVwGgx6tCTr9Dn+nlZPeXHllYIMerUVbHW
9i8hYfrY7ujyM8NfxKzyhmK66Nd1g/UtXxlr1dBGf9Z7oqfshoMpGsEETHmBbAgyeh2wJh2E54nO
q0ZbiNm/DNajMuaarH57BqSK59PnwXsnT9ft0oWADSghnhGMiN5AztgwWwOLzghvtuThX2vYCh6a
JgwTCJOGyHgFb0fxsHBUuLt69i1b45ZXMZS73N0GI0617aRNeUQHvnlPsuN3lq/MktJFmqoUO5Cu
vPCQHLo4NtEHc+0Owxoxwnyxk29G4f/Dx7u/Kw/sD2fUQVycuURWIKc3lt7L70IWG2q99a6xbPU9
1UgCD2Y/Pk+tU352FnaK47lr0tSm7BjJPAfVFdVLLVlwNkwtZMHTjGB0Sz6r2FMhCu9QP0JwdGUr
ujdZvad+YqhIPNSmliosp3XYg6YsILFVh4z0xrA49scmcSclipiSDg8Q7BinrdahQGF1WFDE1Yli
XfdxP6EDj/dy1tyydgqftScNtNRtmfEXdAYI9kTdb/Ti0F/AANxahjaSmkTNO4hGEt8chFT9C5Bt
nVe1ASH3Uxokhx/gTxb0cBwgYjF3euKCGbuiuLkeTu2X7sZyN1+RqG/HcI3fwIaK23xSQj0/3Uny
T0/vJ9ypTarzuo4U6Au8NhhHbGhPhx9D3TzTLw3bjtWWa2omNZ1uVJYoD2lmLHIlfkfUprAbTW1T
vxIk16Zueo3RsqVZYWLflKqcVsl5A4lzdYtf517mSa9ixffAZv3l+swri886Khuc0KYgQHRHRaqb
REzBwm2mh2+py09ZukQRzBq6bcIFyI86BMtNkAPcMx+GOwsQNAPCp6UzXolnCzhvWEnzkabeLTQ1
+BxR26T364qJZs0Sn2XiDGDUKyg1TYX5oVn6Mlqc5Wk1W7y5VqxKKbsQ2CEYU51i1tK08KtfPsHZ
ZeyPcNrrQeyPGcUExeb84CtgCowXg41SCaeQCqqLcPxAyq+TG8FlOTnMSw3BmcYP7MSJmpRHuzCY
a4bjHL95EZ2omSFpn8tisgyhvXlUJF26yLIuyci3Kr3jGoyzLgZ1LihvOBJXy/QLwh+MXr85kafK
q+5Skfxcg856tXsATIMtkpMJgmWORwHmFlcpNEzM72LD25e5E/BdIsiWfaC3mqvOgHVcutoAVv1M
BHvzuXNMFHp6gX0xYzBM8bIN2mY62zWGHTu436uir3FeZfdjFEI/cMdCDmLQSALd7WENJTEEghbg
lXXiCoyHUDsspHinXlsr/l2A6VPApebMI1UZyRBVs1PhuF+IVHyv3J7YIJqOBJ/zgEWEKPAk64j2
FHjhMgiw98yXNw56hTidbf18aE5RoXLEKaHKjlWPcYaNIcnw37VYK4CqJsjEeFAB6BifTNnssaSp
yCC0NXg9Vqg8zzlhmmZUAADyKFicFed2VOt3t6DeXlJyfkZ46cS3kv3K+jXzVSaPH0Xb6bD2POyw
/VWxC+oJ8XbQNKXRlgIycbKXoWYH50s0LpxOTDYhbR11i4Vfa73oIdtj7Ppb2UOnkKNSbeoGJEoJ
yThhOZBWC3EUSQJ5yDmYso9GUDnq8aOIpMH0/bf9vIq9pA9wy5kfBp31h2tHsXNeRBROwqKkvOHo
f6WZTzT1H3NVeqwgRvlmAGFiMoats+izCfhbCqKNaHdkTCopMLMRompyjsjeUBik5yBOj3sT8s/7
jphGUMaGNBdXPIgFlS/f7J4jHdgvhIuFX6Ryou/GKOfgF5s+sD/pnqrBkLHTRo2PrfZyHMug0tbz
F+YPbfVlMYooNEvQzUlmdyo35i265hGyBhk17TilKqt/42V8B0svrdnmH5LvzmXZOcmIk0NgPOYS
Cwe+4gTr6t38mgyKEjF9dLCUm1jSvgx1lrABV88Ig8mz7+AeYLicWf59mq7bqndpn1rJUJ7+GohP
iPQla40ZfH4nb5savPxA/LUT4glv7HKs3xjfhmft4QKvfa8AOc0EeB7ikFPP8U5SsC9iCOrieOtI
IcQiYtszesl2ocK5TC2ek2Opl8ngCs9Reqc9LZ89q9xTj3qlmbV2hMUK9CdCd+wUsozQ97TJ88vI
V6WhCSp4vpDO9xs2m51Ziw+Zu8726GW+Pde3E0p9iVvOqzt10TkkFOWfJe26hSl0Wxm3qshuUTlt
Ny+GiJuvtPjiHJ2ZfvOUvOxLY41IW4LHF7pvOk6l4rctL8eGIFuYgTR/jfl0xZcB0S/CS4s5hj7n
6xJCTUzLMHAVWQCAPyIopP4/KfcBpCTUN1Y1ue3wS2fr02dp8Wh7V7qZAHN4MsdoxIEn964MvjWV
SEGCMZ7pbnwbvkwOrfwOHpXVHY6+2knqh+ZXWmyz2++YQofbCQf125Ylkfxy+g7wBWZbvppXMzfj
3/Tezc06o75P/LIfAhZblUm4LKYfwZg8tq0RSNEFOZ1azW5e6jquFP3mUGI50OY21CS4NcYklUDa
jXEIQvugxf+pgDiSQsWZO7TBfK/ULvB/Y9u9dAY5tfRs97j/AsPz5qob44y3Iq4tICpaUYb8onNq
gfm5Ta3+uoSRxapw/gNKC6CLCnuiwA5JjgoEUOMShYxLG6Ti6VO2M8uxjEpvJW8pqlRY8p3a3rxU
bcovJQHCx07N8seIcFU3uuM9SLytstjha9rROsyFQ9A5x1cob2Arlxf2PFLe5dRGbX5ppk99Bdkl
S1hXoXOR3Hg/7YWlljOAp2CPdmaNEstM2pO7JU8BdbRgzMTFdUHemMU6IYqDoCBkg0rCff6HHote
OPeAmDXROCS4xXwHzIje7X67CZCZ42fLSDKWkiVVMWh8zpKgyBfyjSZ5K18yd+hakTINpeBkKNvG
4/A35GSiD+yIhlZDTMuXmkPIzdIWVx8eBKli1e71iKoQ6XRo/9oGFZhNMAjBQwMiEUxRgbc24Uy0
9UGp+RJ/fW05dBaRcOR98PCpqirvpWIIpx9ijF/S494PuUXPrkWr3M2K4A2mmKv4C5GzRQEwHeqL
XUGSVkcGThzhn04K9DlzlgBzfj5mr1iJdlP92NWkVkzaCDyi5y3xyTNqAsK0X4W0JMY9iPTz3lau
Attvpila5ITBnxy4JtqgX/2EubAdbTpUAtpGFsBNyHCjsOKvvjRRcLIVfDmYPaLzNLrXqx5THK+S
ddQl32Eftv3w9z4uG8jsYCEoxHh5MDT1dUl4yMknJrpPglBJiEYIJCAtwb1Ng2FpyV919t/JLze0
7oHDSvaSXcvTcjb8WQNNxK+pMmdxGfLu/4iBHxYKtBntIPyGOCh611eD7TTHKo/c4HY4RU5cUXB3
a42oZJdqV43Oaay5+QtDz3kb8OnCkGaO1FvjLBuVNnk8SwpCJTM46sHU0+peeCpAs+BLrBYAqTg9
k1D0JcJA40DtctH6UXpSzN0VQ4iip5gIwM6oB95LOFivcXe5ls9KrXtW1ciG/An22uWoaW1+ugKS
cQUZoUR045SzV4fV1xgd7I/4TjCFi5kHCJgcRRijFW1UEMl/KPr22ZMnnWz42mpeycnfvnSeAa/q
R+lpxloj2ejEEq5yg4lRe/ETnZA7cNN9fgj7qNh3VnkloEiFQ+sP4skFCWMhhD/e+fORANBHrG+V
CU1Drqm3//9p6IcYmQ0lbwSrzc0lTHp+pKddFEFXVamyCPryXM+63umF4o1ijDBIeAFImPSUmgoM
pe+RxcuEB6j8BjlA7XmpLHzUD8ya/wwemSmnzG62aBmh1F3ahVjYysFulVpNvkOUscqYHeYGTbNI
S56l+Kuj/GSXE+NEj3XoGRXFfKcQsaaZadvYa3b3UbmLfqqnf7ZLzNWNP6BRrgcwV73kxlCcgq9F
X4SMumvV+lJCS+baT5II9INbz6FI/Ku73VvUEs/eeUw3PsE2ALd9b5VlmsYyypDyZQ94Pmd2I8qm
YShaTOxrMl+UXOmPaf+45iTXSv+A23JLiNkS/krsSGiMJ2StBHXCG/dwKXujzTVUsaWvpRownvhP
CrKnQjwJIiOE9qtLqEHyx8gTdyb2qqpE7iAHfDjXIWHLZYxB+K/tXnFRNu5Gi+42GqfXYm/4Q00M
cqq1Rd4rVkZgDmlmfaWpP9gt32hbRY4/d1JAyvoedMOjn7v4+sBt6Sa/NhpeJy3q4slALBadni8h
t0kkj6D5LSQv/e9RtG1DTMs546+mk29e5ZbWjsncTRyEJzQZ/ZY346oDsYAW1xj4eBOEqLnoX7Mn
coPDuZ/cnz4nWl/nv6l3e5dvE2KwZ8YPOEgT282jlvSCmx+/gA0cqX10jFOejyeneBpUlNkVUFUs
DGSfaNCNIL15WW5bOK0rGF4hRmfMCAM9znRBB20fYFnlXtnYbsVmnCWYz4FEsDsDR+oOxD+Pl5mf
o99Z1Zxowei4K7EEnp3sTE0ylGIIUcsQJaVeIvhgEF6oQwSlefMTDaBqNNV8TCfjcTNUpXIjAudV
kKdHXmWfKfXPM3BFHvW19SBOVeBIQoLLoOoz/4gSRO5zDEJ5BuSv06kYGt4T5cgvr/XFkv5+SS4x
w7KMvc5g2PFR219hBM6XQdZzMLvKxxTHeOSh9B0sLAM1xpgq6yC4tk/98VSzOFv2ZJjoKjb5Z3o/
Aw2Dvgf9CMR6itMJTYcdghFzZ6YvUPXApOTEsr8sIPHpGl5QU1ZAr2RHMIjy3uVuJ0brE8vkkNuU
V2p/zXakrz9VvaHoGAax8/fO8aA/VquNK4FRRuWZwquA48JhmR1vZzQTK4HVa48Ck3UAk0jrb8Jf
viypqveGyOYgWNCzhJjqBvYLlFjdDpqGmvKgY8LuxAaFJJQp9G4USPYwyA92UvRs+Ny+AdaCg82D
xdm66K58esjILi0+S2Glf7pNRuGBKcchFtV76+7lM6xQwC2Vt24IwX2RlEs9LV2PYSdhPbYF3q4y
L6WmYR5AZiAYS16HCYWEzSFJ+RnjAnfxUxre5oU0PYVlIEQf8wYZhzQsSB+GoNr1FlUSGnGkXbxK
y3sSWRl0pwk6vM4aKwLTkXB9vv+qpsGbmcd+SAeBN3YnHUYdGou0int/qmdZLkNb4Jkcy7Su1EZb
EOrdYPb9h7BhvboGHmZ9uWeqRSx5eKWH0krY8A+b9VoAgHSp70WZQZF0iodD4kF1ET4mG9/6x/66
+xoen07YhehaaSQwxCim1SQerNJUdeM0WbdXe2OFSIx/7Ug6I1ZVO0P/l1CNVTCNlcvTaoo1HRal
CuMGH6iz0UsB0JYcuT6nCBJI45MTwBZ0jG/ZzNNQzm0Tkx+WDf0TbVEvtofKAugWFoNIhKImJDlF
3Zn3WqCYTQvq1SCafYfIcWGJHw+J6mQ/SaaPkjqVtobk+R9QrvypxtE/Y4BPf4aSvOdq5zhu3/gM
FKp5RPh9asgMaRS6nm2TB3jQ6Z0awQWEwuhJ9hw97lgAfQ8HM7UryNuGtNBuhn4YELl0062U+GbG
BnEeLXgGP45gtRoqz/rxXFnzZJp58A+Z5Y+o7gnJAKsjyVa8QiBCex9DzFw+TAgB+X+aV99Ong18
5jDA78e5MoP8is/8myI8KWQLr+AmCWehTweQ1B30ZAJYvxw70oGoZWsfHVocd7aED1iuhbnFK6nb
wjUhQKtjOnJ6JP8MgZyXc89I3yBfDftzeB+/kJFMxu09tHRMimwoWoWXCy8GvW79fHib3CYwK0ID
sZqYwWhh1mxht16tLYQM9K2PaiEgCRCwAZMAJn3r4+/E4JarkL2chwPowL0yNzMBFicbwOjjolBJ
TyfQ0S5Thx0tl8od27aCyAPpLta8LNcEsjADASxYgeZ03w1HncoR26Vu9VMwSQ0jDUAec9Tt5Zsi
h99f9WXY74xaQc/jFI8zA4GHcF3sccYAqyVAXnBcMbD8mtIBnReP18hNn1Lao4c0/IsEAIOBlBS3
FP10RuMNZrEROKNBgC0Jn8hLN129cY13C4JFvOk7tj15zo4qunEiFmAZEW8BR6PwOxWBIouJPscD
wUbaRx8QAf6wuyzNZ6O+d1wOxAb6RdZ9+LqOSh/XRTbomF9xEU9VeJdxbMvwniWFEPOGSjbaRg3Z
gfEfn0fP9AOeVUskfWDI34OGv+EziQMot0gozhJ5pyDRRd9ohJom/eFzkyrNpwfBe7d332NY9QrW
cxS1W7cuEeyOPi2byGyQsj7u+Q4VtoVntSJZ66C3rVVrzGE0PLSGDivCmYy7Pchoo2+/BLX18GSH
HVbKcAt0eaUxAkNsoixdGvoP8VCpCTewq602I4/ZQk73RGYejradm4ptqH1m743XRB8zhHBTwF5u
CAUnsA8z9t6RKoHx8c1cue5J31UZ+ULOoH9D+LkSt0oUFAVHGbTBu6N48lxSfAnSQGQBnpzqcgwm
bNssT1Yc4p+dgh9d84nd0E0eex8StZH++fimsgEZPz1f8ZxEeAKq1zBKov5fZ7ROK+G7eTvvjf4N
i+3RO1I+D1DgE5D7XacXToTrUIoN1B5psgQ3M96zBysNRQxV25vnbGusX9moTJDtGsTb+SGCI82y
PFUf2L5/8ea0cMPP5P5LFBgtbXYVLEaquvU7YRwlAUzRoJeBEJeeWgaWC2hI7mr8w4o1QRm6VANp
7RLzrhJBLawG1uZJWGxsk7Smt7MIXj5N0TY3uuu72QH2ALAxz37XeH2SqFkSVWkGruMKzIlYWsXo
92nqv8mvzNGseymEscXfnf9xNf9w9CCEq6n+JW23P0HRPJH6eMih1RLcmiIyd+qHuM9I58Omv8qb
r87ev4+MBzBy6UVSuYJ+5LC9M9+S/RUAC0cUrC3DT0mQmGmEX394Stpdu8o9fMepm2NzyZdllo0W
iZTfP8VUO5HwwBxGS1VaE1gAAlekCifDeBUc5LkUySjP98kpulw4c+i+1hp3B7MKpjOdQ4oIC9rb
igId8vaFnLyexp5S+DoXYaD1xe9O9NyP2IaorDroBgzMzADsDlRC4bLddbVRZDU1mWw2AADoW61W
rkeUeAr1GrZAO4uCE1YMLxFMtbJ7jlxcMCVRp7xX4NWA1Rc9fdajYdwoqb19AlS79gX/TRY0uXt+
7/BkvO1JHTRUCRXZWg1CxNe6DpwRxw5xTDKTSWt5GjvggDLRU09luJgzziwv0Kv0EVWQ4B2Sk4Ej
feXOQLZE3TPnKuoWa5+E1DjM+vxv3itv339NUOfjYK2/jWILYYQwoImhzeQIQU/V0Yc+FyT5zMot
QhOfRFjPBBHGoy2pWotf/Jj38LQsn+9nHHchROYwfb1cZghUD15NPXR1hz2EU2/i5yLaRF9gI8S6
w71O+CKDAIWlyGfUxOCFJYecpP37+UA3GLC0WaKrovSWfzXVnmVA8Q3XGx33yOJQU6ZLzxAXgid9
SQqMgLySMrZgiTlkpMgrqLoWFUM40EYkaZy8GjhM4X/vsO4GJMg8uLTPQvYOtRTYP+CiswtaX3I8
lmjQ2kC+5xHQ2LZal+5eQASsi0fRKSvBkldVOWtlVVSNGcJagYuLx3eCEc8fp1Dn09vOXG4C4Bjr
1FCF/DLEAEveln+IoC+XJe++YieulVJu30hG2iToZylHvrAxk05Sh9NqxRH6AbU9WkHy8MYQuI0A
oHQ4XLuG3gXFw+uIjnAdmHYBiXFJdK3QMZosCJmFuvNcJx2kvdUhpsplU8xIoLReIQCUVlBEcC15
hpljyteeP9Vm5GJ78Rs5r+hbZrPxqV5e0kwRnW6FN+bDZ7FSwCT7Vvf8UDxI6l9acF7P2fb4hokN
s92pyGwqa8f21CqC5I83n/r3TaAfPrJK6TsGiGHPXKZ+P77IUcmeVO0E2otBwsec5bxggDqvloFS
PI1I4/0wKdhzvnYLo0DEJVv7ojJyzuHmzp/R3xNHCEJfT6Nc2B1d906sP/9iFXunU0qLnglqBorh
WeOBDqXVrwiOjE+lUIYlmocFBdoPlv+gUNqCcdePF5vN6Kiwrsgn3ez9H3weCLwOCVzvs6WUvy8d
v2clAG3C63MeOSXxUiwjDGlW5NJHUZ0panFYTDFO+ywNZzt1/C5bg0lC+5flpbpDXR4vKgzBnX2+
pkadghNjrmbNszQPsK9OwPtbggf6W8zfeIVayYWm5otGIpMKisxguj5XQ7AUd31iao5X9Fq5XsdR
2FRrXhbgij7H6yl46KtLa0HRehp8e78OM7mUvNM7HzVyNQ8tg8t1h5ITAdoUf4jPPy42wDRKaNQu
ZzTb+2JLPX1xnNnLAelD+P06Uyhf2FXbfTi3Qd8yIl0OoAFVynVLgJ6fXE87BO/tOEW3Y5XP4cuv
pVDXOi5ij2UbMEe1zIu7L5oeBu6uOLKOeC38ASN+jKumVBKXk33vQpIVe2kBx+ABY5771+uucA9d
6ar0uL+UMDKNgtiGgodjmJaFtQlrF2+sab5bOPy2bWeo6YdwXQZh7giEeAOv4XmNzp0v/DtndQL7
h1Wh6e6ALueKCAEYRIFxo7U2v11ORORlT6EKcKEKe5UAuT6sVs2EAUgKJGJrZ0gLmP3Ej/BfbDB0
tsQo21YdhPA1eTFquu5jn7kCwZePDeSAm1mlT1fTS0ckU3fUYVzmPGB9x8bG/GVQpgEfCIpZBvdM
UfgYKACeWQ3vb5dX52sqfEiQ4cg1BtQwHfAUUIN4i1qNOBm4Rd69/D07uCXW4PupXJ8I5HCoJvCu
EyZhBeSUAm1nFaPbVz8scsxZ0jt/L/+HPxd/QCOJg99/ao0zWiJvnwI5iSGrXYVrC0jYldMcyO5u
cNukHMu/l4gW/XsSxdR9MKaSGP9BcFv+uciBih2pKhooOQFxAuQmD1uRsJajh8/kHXsZd4Ck8/VD
Y5uNN/oc8FPyBt5n8PUBO6dCduhYQjVDgb0C6yArl5Vpwxn3rG/S9cJDPBTPo8HF1EstbxKuwDPT
TVyxhme97SQmBx1BzcXe+Wbvy0b4vdmwHj6EL08Y3KZd2lf0P9AHNDIR/JR3PGSoQ13cGhcA4drd
+U98vX9JTQ4nI4jYbuht9fdHUMlE6udulWqBRoz8AgH4qEFvpF1JkEKBkXrhB2hLTPVTNv9L2oMf
S2q27oHqFkPmCoUkNrdTUXeD54Q5dTwuaN+RqrhU9hV658hbOHh58geCRFw/wmGp/zOTZ4FpyD0l
+e3LXgxxtMD6ucWkz+ATZ11vEBjOOOFu1pVymTMA7r6GcJZZolRoweUp7Fd70taU1mfb6Q22uTFh
UrSA5AP2wSptci4uGn12/LnZSk8hh20TMt+bnxwS3u64C6Fx0tIOyBfmrDSHrd8g1HPavNWcxXhN
w3HLxvkcarK5LFjKLCf09f77mPo5W3qEbJ9eqt/xXdEEvfZK9+KxfFxiUfo/m5PPQ6+v0RZPyuaD
nITokaGiCYpsyEBYg11x2DXf5tE8j3jwxUiXeDK49jY8SQ6nA+DJ8+LBDUENVyqoSFo4HiYtxByD
/i6G4YQpWORTAXcuEHfgDXuOL96tXSJtIfmI0TEppCT9ejHEicFldsL/Tkqu3vTvuYNi9PiThX7I
6KIsEAL/fjHdFAutHqwrPdMipyMezxt2WbTGHyYvzgbTFanODkBMPD97M7GfXgG9vXwlEOEulwb2
DpnPCoJUmOc3K5ebx1tg3ij8BNF+mpBcRpF8mH/hMq9dSmpZrFJ7WhwaBhcIDWCkIPeVE+Fu+13v
+EAUUeiJqis5VrK0UtDKGLnadVOpsr31QK5ia7h4vkiLC09ROZB247wWbMWtm1AHPOT5cxoG7QQY
W+ZnNqxkYjmI/YEeZP5THIVacw4VNNwYZMDcKf50V9RPDEpBAfTaoqPSfczSNR70wMaU0JTl+bph
q0cWR96OBYY2xppRsG9+qfKzQqEuNwCtHKjL1dMab+WjrEG9u+5bbGtmug+4UpoP8lFklZ3pcZUy
xs/tObMWXBwpfBdQsIBS+ifCydbuc+jEFfu7hj0uCI3Ibgpitd4YX8/QO/B4gH/uKzIE7JLsQumV
MUXTDwlkcKgs+aJhZ5flz2CuPwvVxhiqKoPgZsFS1Qg19A7B1DV3WHU6fuNWSw28LzfsnuZ54to2
lgjf8r9PonA2ZH7+Xoa00k6zYQliwR79v4ClwN2ISNARrNCobZLTKJaeIddkNA5nqo7B7wNwsY53
kiyxS8B/aD5L8AlwSoBFPs9SId+pIwvm8y1TRXMZOkConxOSY4Edmx3wBaslBvKEuCKCJiLY2n+n
dkMtiswD/5NFxhOatEuQX+GvSMzntOsK75Em3B09CEGki3twhF5DMRT9AaHc3Pa2seOtoKK076VR
3iThDeWHY/JiBZ6QKEYBRzOf5XLMrl2m+tD5GGyC2j02oOyYRbmvcrfqqEfBHF2G6uLGSxT06PdK
UCZipQAEIuMZ2esyjYAFARsUP+3UFGln+TsHzafPoD9gwu1z7xkjXbE6dllZ0ydg5PSVemuB+GbN
6y6L6ktx2Q14WywXC1MSA6AkdjYAUIDmU+rp9W7Qf0kmwRe+qzT0AO8gNojkoKAAJ5Kov9fY0ZRn
Nq3lO34vSatidw7s2lqQNtpoqEwYoBfkfO0xyjiYQb/twA6Xh85X/ir4O6uVj4u5c1583BEW7BBQ
En5RAICgZ8DxnMytabQPNycp3LSFJPovD7sgHNqJzuZZ0HnkwHX+7/QvIEgIapAwB3asXsZvBua9
5+EP4czPOzd9Z+wBPPZC8BCRVQOtfcnWveZcY97zSyO/vpx21G3uTTTeCEKgFff6kaUZvWapjdiV
CAJYFFeW6A5q/WgA8lVXallv263+ZV/8qzZclWvyhnTMUf9Chq8jvEY1YSnilT9a123kz4XOq7GJ
M9oZooaBTXeuneW4YOGqcAPSSOAVnXdeX29gxp1RdVQ1mtDuJuUbp88495qtUJEXDdCt2I2YKdHe
6txDq4htQd/VddMQzAeNYrVAxPC+JpktmNZfbn8WdAlFWeC6DbkyX4XpoI+h5fhsUrtvltZHkU8O
mlRIuaZv3Mm5MNq9aiKPcFNmvm1YvAAG5mln/G8t6Rwy/IOA56HkOefRZ+OtJgWc4PHbF28TECxB
Mlr+GeQ7WfpvrB59vDAjjIkbLg3RP9oOq/AiLy3UK7/DDB6oxee83G8s39mk8mfBoBay3iYMRHEv
T8GcPxyHmzmiol1U7cUVwGL14UD1x0QandcTIL9mKwYkeTPHkUYrAfGsqqRhL8NbB3phT+ZblYmf
scCrRrlJrtIpkM5HcWi6OBNyrsqZTAsv1bn0yrFLlAZhH0EF0TCDcynCNxu/Yi4QBC7Yk+V/gYkD
Yy8yuDA1JqRBzfnNACQkmTxTRQOr4sv5p95VoLnrcrOjGjxp7tFrCABew9r33rxtMhgSssP/nFsG
/669BtT0RwNPyERz4K/8dbkYlpKXR1g/0M/hNh5psqBmBzLdcV1nrSDQ2AWL0bWHOgJA5reEq4yJ
LPaOYTJGwss8bJYXrRRRaYa2lTle2YFJzE5NhJ+ptgJA2lMe5kNf8wQT6XcKbIK+FlpHbI8eX/qR
im2cLDVH75uRlgBOrJSuZrsOFa4748B5TYbtTSvmdY/nsJT9RaVVgqyJEDLt4y56HdUOv8uJNEjG
ufsb1fqLeiKBwrGDJLQW3fovqPxec4OPOPP1ORlQN3u7yMuUYiYWTqznPFunZfmDX5/haoLAIxzY
hzfBz7+2MtwTySN4s1L0hG2AZO8UWuErG1trt5qcCv6tg/U30p8uE3mLKeNUeoKjc/J/TbXBqzft
FlK7IqIvmO0BwB1zBsJWtFD/Q012IiUT0CquyeoB+xYW9+Qs2nTwN1P2/jgEyEeoEBZOXWVnIDCB
ltO8zJzFYgHZm86+2yyV2nzzwKmZ8OgqiwHl4nGUHaQDlhBPmcWgEdAWkUDYnU5eNCoC0SkJHVYQ
xbzCGd0jChQln0RtscUmHoqCUtxVlcyAZSWwtlvGsnyvWRW0+faDcp1FYmi1gEsGAy8+L2wJ89cX
2q2gFV1X6bBSGF/FS2shXCHtiaeiobriNwcFzxJ6JmZT5ZYeI97aLX8U+aj5vsABQEYMg3hY0FW7
7142SONW+wrhKR8IYvUqSnJb8RK8jinz+QuBebAu3btRITHS2KFqDmhfNROflkKYky5bYsrtul0b
SDCyC0nIwpSF3Iy50abNYX+6bTec7sNiyCa6JlKacvpi3SH8n9F6APaOZnIgF+Qi0gWaendveT1q
SfvdLu0JB4jO+Nxgj4nNGyNqhrEbFBBWx5k8br0xsZJ+7CPkSSPrIcni7Cl0zm12tjLRBlqcQ1SL
ImNnCSSuSb0DHzkr9H2f53GbUU7+Vce3NRdzXfC9Eu4DYvPkc507H/7U2QxIILflPx78Su32rAbm
tk5TJW3QCWIPnJx1RyQ1syTUUMiOYVpF2K27uKI48AsvYfPHoRbTXy9NDUjXk/NrbXKoyHCO+sfF
qeFgCxkmIFpcz4yDh943bHPZ95ADjMG8ycSgoGyQFu1n7gIhHeOSkUAQjdTI7o2EAgrkpCIsH/vE
v/uNRXMvVjKEho6TzkVu7BbPxNJ2QgXG+E6JPNoCZkqLOLfcM5HQ6rnF8jjn0Aa9CxzbstGqRmwB
M1prbopOFqmN9ar6lzd01BdQe0mwIXRb3ejDxcSxXeVx+G+EjXWEgC8b+O5onv0B8LzuhlHAUleg
FHX+r5D1NZX/2FgYnJ8CZQjoSrQY87aVdXqmMMgCmMpXtmNJGPaTQe74dQdeQbIiD9fqnXJN7sSO
UCeKr/q0hfiR+fszaZyzSDa1/4BG5qytBrYk5/qSLrrxgf01dzn6LJBU0WPI5nQIF1AsMzt4fKDl
HsyvDAqiTo5An8mm/dk3IhhFVgm5UH/L91xMWNYstb8Y2yPHenxtAiQ0biMTnbStfNmzWesj6Mew
6Gw3ZcfpDd5TdLjW7H99oT437FaCdXCAfrqHbQ2DkmH/O4zXc1np/6yAGoDsfRWfhqyC9bOkIKzp
U2nuJrBOXyI0f8JAjUGGH5dOAXZwwBo5kkGX44U8Np/EqSPw4UzRirvw/vOJMOj2jMaY0b6PPj05
8wrOBVF+vPqmwCNTQXemrSwXLXzJqsrYXZ2hVK/wUQrvVyreSuyyVkYaHVvg0lzrD2EbajYAvzsY
GivThVeo9mkdlXsoE2lDxB7lMAZj7UU0YtTkzb8fiPGRo9AtSWUb6sIGkyza6IPSw1BvBrRcersJ
spp3nYYt9Vj4N/MyOmGnnfYLPLkm656x8Qe9S2BHbgqgxzIAvarFicjTot7B3CpNq7FxKKV+JsSv
o6pu74em5nx79IEC6rNZ0Dxl4HtxrXGnF8skwDFc6tSykPJNNkZUfRqXmeeWY7kZ8FDPUbQrs5u0
2u7Cl0fuO+k4nXrUr6d3i0ftwh84ncb6OeC1nFKb/v27G3luMeoKExXMXoI5FIVGhSSf0bpTYjoW
lhlnQlhMVVE7b0lytuk9CfnHM+Mkc6hH+SVT3yfmITq7kkNL7eIPgmRMd2PbrkgB3HceGam15ZAX
IpPOQWcMIrlI5FreJeMIjMfPatXf2EKVjMpHSvTviM5ylr117mQFC8kno4sta9qjS2xV24WFB+x4
1QlcdiLSjDSZw6qbrRAAxAEPWxWoLKIn3x2h06AXUf09UA4f+yeMwsjMAO+7xh2EmRpdhqKjFxxt
aFtcLMsWNdUF/mWavBQeqt0AH4wzOYo5lnavuKYbF0AvhPTX+51AKz8TGEAEEx0px1CE7krTk5rh
SiIE4A5m6rru29EU4ytb0MoikLZjjKgd7pjO2aYHG9vK0UPC5RNn8m/aRvLSIWV6s7+WC2FZiuri
QSoxDuZVKDcFW0Tel05AW/2XeftSztcE8YIqjt+6tH04S2Fa0gHGQGeypxoHZR2xo6UTJH/2l4lq
E3RhIpaUam5f+dboeaVeKbOEOYNJQ8QGNfMJr2zF2YmlwF5zY295R4gIsgNjbRbMJi1UyB3mCA+s
2SpQdsfZEvsNM5MUfe7iFQFxr4ZM8eYPEYkVfT6P6MAL22UNldRJmOU/DpHTrF4rCo/+kPW2k2ze
5f3LbLw10vKZ7tHZkTv0/g7ImHRvIbWeY/D2WXGJtIxvvD3e7CDYTffZpeoa9RFrlEAGXiE+nd9S
OaGgXZiNxgM9X6gdtjX/i4hwa6wDgvRNiUbio7iojWGpn53qAeAYgGewYYh86T/bpu9LbsbcpvAu
0ZrZEe0gQOOLf34A8ZMM+yhWINfb45XyJxHvkLeR048lyPU0TQm+Zy3Mb5wQFwD8446nnVabX3DT
dELegn7BgFvho7F39QJF4fFZYDCBMvkDHxIsiuUMtnYPyjA/JWKkTC+8M4TteKKjtuueoCo/CLRL
UIxR0B3XB1EZ0vG+AA+sM0USSRmEkTAfGfXir4mcxeUUXMrEoghHb12TqX9bAtSJ3KOflxpBWhcU
7w9vtBkgt4U7M3YucVWXAZRTgaLRQdV6B839qgZEFItOKLjx9LrO3vyheNIcdDYj6Xg+Uo2gnEcI
hXl7VR01oPIzBhU/B57ynGgwykCUV+YMoEUkkUnKZZU+e/khC5yClkavHC07ttYNhYBmTiVsV64E
LLufvGnE2sVTkl2jXvVdbltb7ucFHy12RGcF63/pwi/hE856wCSVBqFDj2eHQ9zaTiPqZkevNOys
l8yEuJmHapFrNYfY7Qo9MuP6zCzGeYiNBGIAbCyjTFiVeqEW5e6rt9bv3ZQR+Cp0NPUWBSjTID9O
nnohAIJJ/KAimaipxhwZeiMZp5H3Vg8RgpQFSQfvNxS7nm7zTTlPBlQWn+wHJvMfZwHUI+UuQQAy
TGo2tzPfjy1r5113MI/tZf7/rlQVrdgH6IzR7aSIRNMkINir/PuSElfYUZzngAUOsd+FApqIDPAq
zXl/UHzDGZgmdT7K4ldRtE8s5SG4nJZzcSCuy5UTQ3cYPAu7psqIjRumh8C974suwymGFmZ3QXj7
UHimviaV//x6cgUzGv3HxiTZhJ12RftYRn4T7QggcykJYEw/Uv2fO5peWv7NyROg3zu6jptuEkud
SfaYUFbBBeRXAjBuDsvV5aqweAXA7Y/T1ABlRm43w8vMW7i6uURgfOKQc2GdsqjGdMKUNr8OxDmw
M3YLq67UGoXaZbMhhPZrxSPu/T0mvCfZHspwU9XZqbm2EiZDU+geaWeMMwnUpysqilB4kxi49zVu
/4hE874VSgktivl7+aKGleqmiL39zIoc/L0AHcgKet0vk5aSDZC4UbOcxcy8jN4TpNa+fhR8Z3MB
fe+r2HEsan0ZuyNwimMNZ7eqrO0ub/mH3Y1sr9f5kMHmt4vNgFE9MNhTNuXoRJdbW2isNIb4+Qw/
ZAybfXkmGHzUZG6ctzGV7YB6Nv64er6CgePAGg+5k4ljQs81C+nFcON9HUFe8h15d799dpfgAexv
QkR50fHi1QR0ff7Uqj0gM1DxIFGzOAgtwH294+lJPHDF7b9fETq3KKJa4oVM40seWp47REdhLt3l
emliNc+5AVxP9cVhURbXklHW9vVmgvkjdDlPayDhmFrVJH6Pgr+39WKFJK+BSzYvEMhniXrgnbaV
p3IJ/GZxrvYwVorb0CKCU5Ji5fSXICqDZ4py54IjPz2kvIjItj6y+4Vpg1HlQG1/3oEOk/qkjX9y
0+WFLFhDvFaK72xHrXihMqXtCJ9e4FaGq/i+r5VD7zOwx/Z99z+Du7/RqjcD83olsuKlwyx+stD/
H19ETLubuOOf2LC+GlWKbz5oKEOSufCJ32O0c9U/Qrkt4lTIAuo3Q7Ksur37pEedeg9TE+1OgpYY
tXiCZE9l+55b/+y/545wkv5vlBxnCGtxwEiJQgylNxI0D86zB3Wl/1gBFj1g7z/Y8/zerVjG0ahp
gQ1ISKMp4bo9eWceI9b5WtqRncYiTlXrupXGHLuop0seHa26f+sohv3b3/ct1ek9dkMI13tbOMf3
rdu1vaAQ9YMWDmKPKumgdxV4tcPXanwtuDLpE4sTNkDnTBXqrXS9eaUhVzuaDR1JSCrD8pxbIynC
YTpc/zOHCbr3v67iqKYVgRl1B1Ere0EPXe/U9jT9CinczD4IVPgdGqc29snWqTNEM8wSmLkIPatF
OHMH4CzJ04o9A+2wKTumurUXwQQgemFHTZzmLsDapTeN8sBfW4AWlTtptn6NX3GIP9Vxn47H6mku
bhCrP2uIunHRhcjKKxZva0H1+qN2MxH3Zfn5wSQ5gwATnpqlFETrVjV5yydstDDTyWDgB+V4f65V
geGEkl5v4M0Y+KT0IxatwtZpbPKtf7lr8T5aakrGh+W4kUpgqZFT2yZTEoo8M5gOTXHFN6HzCKGK
LDGcWAYGLxBiPdRXtvhOO7bJwc6OwJKvMww210wl9DgEE8sc6QJW7Z2icEwIUocGGEzqqwXpTj/H
yRjEccSAEJdP4Q+3cXeB1jDPLZM/lasdH08VqUsRtwIXB9Khr3kXS4su1w0sJCS2M5JvG7eTSYky
Z8lDFW72uV6M0fDygOQVuQStzMgVZlwGWa0a11kQLANXG0x+kvOGT7eCDHMChlyO0CJ/3OFOOpG1
avTsR467pnfy9GGEg3f9ZHYV66RXynSrYC55ZoTe7SSQIxYKN1dAqk87DkdqNqXpHAT4365sBWYb
ZzLyUueWYmJx5GZW5MHIn8M/kbx6Su8UIXtyawqlaT6UMsLgaW2QJYmWElI7J3dr9B3/cHIPWIl+
HVnDCIv42QTnjzY7mNt9U9K+Jfqd47hbPc8m1QAZJiYsuGiL6x+xk5CbHBRZzBvVmbSCBNH6eRv1
x5T4o8KhgpUkokdTP7Z3q8Fm4RXkUoLG5r2xA1+bjCrh7ZsGvBV/+cOo/CqQbJW1HJyfp/TTDOmh
F879JN9Q4JMDP3DaghM2IsvJd9OWfEf8AgsxF+w1875vk0wVEAjEVaFz4HCdEfHCVSDFsMgKHeqP
kiLpzEdXAMG9MonqPNqTuUgzCDRMsLJz377kMhQYnf8x9kW0apMh0CtcvoL7UJyrHwv09T/zYVJZ
lxAMT1NaX/qGrHZlHmGrN235dWYlvvaG/qDETcE5Mz/0/tlWSOS6AmLytr2fYNh31vVKJ+kDKPNt
Z4+vV3/HTFWkR4y85fZ2qCGsMelRruiycaVlOCRAdyksjSH/BdHO94RyBdG0gaPMt//Gbzyo8oAi
hn6snrpqaghVjbtcYhyJGCke8WtxX9LYs5KUP+tL61ZF+V+94qv9y2cjjh4IJRkFnHhmQ+R8vxc9
fbFTEBA4h0hGjHA2mgfCt/8h6KzG5x5K4FxWw3MlzXALHGMexf6CgtGIfaYyFDGqotljM4pw8Euz
nvdi7ys0bgxqeogM3qTE2T1uucPgmNTe27suMRDDXLHeYVr9RzPU+7kW11g6oE5fNcGqje8ZG7gJ
ZBsxnYOrIg2K1IeXNiGAO7CBvBp1TSXe4MXVJHLHf6QR0Ju03P39hCxobQSsfLScqnZuX4c+3/1c
UWWxJZfEFlCmro//Zod6fj88mJxFO5H7v3llUEmZgRbmY02/FtF90J31ddgQxZOjNXdsxwn97hc0
cKnhYN1rD59NsTFItDjHdtGvYXqN9n85t3S4gzeluIzXAOcyIKJQpeYu4IkE2wZtyBec+Z5yOEqh
FdFPd/AsJlczhjBXfNYo+mekNT09W0bLQHVNYYMui5fTVgAMH7YWbe44oUiu4jfXYOOSXlWotsxb
SQHPb6tfHAvh/BKrTsYHENcqQIoYiEJ6npJsR2RUbAsMn4fbh9H7oV9yTeGrXb8LvI+ep9Op2Gyc
3OZYWyunLYW/to5NKWlqgNiWSwo/a0EED9/Ktaz5ZaNOIJG/EzVreRNmk8sCJNCimXwgMGQQEFOB
8Rw/NyqekbaDg7bNDc7zc3dCNMDNhS1ZpvmIflKiMRFAfEHf4PoShC9ODVTdCfx2d9Qxt4x9gBRl
eRj4B1XF5LQSmSi/Yf/SrH3ndirBw55oUtIkQAwMycyXPos4M85xImgXlJB9HRxxZhvgVr3sMIHg
3vvTGkI356jWQ9iYwP7GsHrhhsQn2cK7nxDhHM+qHmpyTDBqcjlDrxu5vmc7fEq6j7VjXOE5Pn97
PRSDW8ePPNqQndwiSqkWPNs4xn4jyYC+JE2xSD2xpJezTo4Zp2BuYbFd2ytPqQLzjJRnrW8tNjO4
5hoISNvfUkYBOyzr7aC3C9gC8rZbby8u/fVtgL83bXstcDMlQugw9+bgqwtdH0PQUFj35BAW9UpO
4E/dvZoDvRNsDIPsQDovQ0Hg90JVMoWIz0CLvVEHIeb0GqFsYXPAihdkLTyoxtJJLyy+ckaVar/y
XK/G5zbm7veP1k4F3QmQyt62EWxOTYAGIrmkXg4JeFBptTAW3BreQ+zGlPK9hhP0KLbI48mm5PJy
PGc3GQ6F4Wux/QXIdrofF0S8mP2/dezVDxh9bdS7g1T9LpWfX8AK71RAP//ioul2gXFJKmk2dwV1
S8oYhwYBK5OSOMROPFUcVI1Whtdh+o+2o4SJBFZH2R5iuxJK5m+qCx1E0dC8Ma3YuJWTeNUdVbLm
mXkbXo/LG7U5PBqm+mD1l+ww2m/WIHi/ImQureEDrppREmSXnmSvntQ0VeYzJt/dUpGD9oIatBG8
RoCawoylU9UNRIDA9H1raNJf6G0fGe9KHfFTY43c21skIvl0iPPKpxpmreVybsM12Ok8A45cOCsT
IrujYjyZTaUO7Z0mxxiAjYILxj08IwDPa7b8689FZ664fukB/vW5/HvS8gUcoadoWAdKYLLipata
r9J+WTGHcbThQ1AiOLA+IUu9LguT+RWm0Yr6moJTiWCZ4vEHsJITVun3eZPcdF6F+CLinX8Q+n8q
uYnx7CrNx9mnI2bc4C3IMTgIC7o7oNO2veESfFta0v4bVfi1gU5PHWKxe2bWbLSHOJ4dLa4TJXJx
4UqqMx+ZUXQbiJ/RkgptSMhIrF6QZcz1loXyUkRWeMuj3pJbP1msTcktAQiFHvwjio+qI9NpsPv/
TUjkV0a05CxjcRsEnopXvDTJXhrfafEhHRNFqhqJkkgwZad9mRzWuwVoVcZv5+e67srwUELKkkjV
BSZftGYw6dyfWCgAPeTtHd7dkrsnSRHEz6tOa/fEkwMQddQ9sOAmKL78Mh2BFyGyM9W0yR4MT4Gs
Hkj0QjkfnK/t57UedW162I6CoeXMb8oojRWLfzKDvjPOU+NVMmjxNpOd6tU6R3jhZ6jRKT0BOVbi
eC6/M7ffRUBOKoDHuvkYXaZujZFe6j05VCYjRELGA4KhrqaZLa0pUtQJ1kZogzbnebxLX4MXsQiu
OrSJ+i7971p0eGi6QxegcjdPnzqsxXXXONlvtvMPFYMCPqdpmAxFg8rWgpDtysjSn3O0MscK7OMk
nofdxWRhWMfwFhQYoZQUenqKw0F71HTc5edbgmJrJalTOqz3qtq1YecK2JR3DOL9kq0IjB4+egks
nxNayJ5pDYPR+deLQAe86XHjBnPlXhF9JObFdOJOeRL/0NAF7BFzNCTknzOdhQ4+HaRrtP5w5w5z
QWDjzQ02vw5pk5gnh12gFu8uezmKPs0vmwqQJGfDhB0Zl0oky2bKzFdMR9Q2RCIv0pBZ1t9ILHcQ
jbbaiXg7wj46kaeBqACKf9gVk2wBuRUMBfF305rilPKlcwC5DpxjbYvHg1RNi8PQxpttVvXoWiPa
9gidh/ldZO6rM6zProJkhLG0dVj+EBG2nprROung5YzNpizEulSE12HJdAanKuBYl1MZ6U/nyF5s
E4gP3N2Tu1FUEUcPEPO0v74CrZjZCxAgMArmdKZah/qG4J+c6dvq+Yqc2y725SfsNYP4OFYIzS/g
NRrOAHOVwFPPSv9X+8JRSqiwynvwF8x/K1Db1ZdMQhzGu5SFsoNOoYLHr7NiQFZMGxURGFzxlGBR
bS99T32NPAQTKr9Qi1q241qywdjnDJoNFzjSTceeFw4GOCLiGGlGHujvc2ThQ3nQ/VsrGtf6J53j
IjDF1l8BUxX532jM/26KRfWpWzMSxQ7WgeA5LSVpV28lmAGrGyCMi8HyTjItPCgMtfTYNiV/jF4M
KYKSNxVU7r7ri6SI+Nnxhv+yBHucc6R9RoDM6TSEInPvrKaGCUuOMyISJC0/2AUSq96WZ7JlLVqO
Mv2Be319AFv1h15mlTG/056gFdE1/1MSGiEVkSNe+VJxDjj1zKfAx1nAbcRQyNsGlzNWNIqEoo2O
RkfXUG8Zf4vwqRz4xUX4glbl1/iksppYFkYcb/gJJW6+SxHn4ga/kVaR87ZJ2cpDrYvbAMzIXdPe
Gr86BmfqhV86nPd4Qlkbp8hhlJ1/ZGXk/G6ZVZw5iLsHJy4Z2/pw0MHt/VhaiFay/LBCZdTZEB/Q
C0kCB9b/eTud9xrZMyJGZDUaFU3zuM5+5I2sJffwsQcKBjPMr5DCak1MPBOsFu2Ae3oJeIl7FIGQ
n4RsT+Lzja5Wsr05cUO3lIgRYqHkVddqnwsy7GJTcDI9cZD+258zN5zOPIp/EQ6TcNPRfCGXERc+
I+F8WgwJ7LYXKia4uNOaYer214IlqRLoucDGZ1BIWo24nG5Yhsj5xvNcusO5zYjRuliVIKU8/FRr
BWshqX1O36cW46jKlx7MkJ224OKJTZdCW0y/xgmk44wrcs4lqFZPaGFLaVbl8x3sUet2oZG7j9U8
Jbing+cTDTep4e5jg3naO2cTS9WmFSidhcTLX4cpqXPhux9XpZDDHiR2bPbBsDQ3reJxo/qutdAp
/MGMp3foPcmoZtXcna9nvsr2GlUOPhsjTWT7nYY3sXZ2Z5lJx159pu9DlQu6ddBcPsSpV9ea626Y
LszvMNey0PdSw/GkP4phoXxdgb5KHWqP6LhLy02ls9bFMzgYg/qlTdSnmjtXfa8XkHFiJBT+emgz
mO8Em+i1YaNrI7nrmjF9dPrburXKj0Sv/alcmj8wzIsEutfpgSkkWIluq1+a7yxnBM/Y+2N7Bmqy
LHGicmRzL7/jFBgCOjjyKIESol5/1qUm6f7N5ePT/Ale4frDnDrmT8/jwcH49MRIiYKAfG8DDV/f
wEMVpWVlRaBzxSSupmNofMASbpASBHV91SPPVisXZqp7W77ur32vWvt0CB/a6zVh//0DfKz0ITdH
Kplqllin0cwAALdbb4NY9j0qWv870P+a10Ia6JQ+zSJcvCtKFm2Ke0I1yNESVXctf0QGFADsW6B0
U1KbE/r+tKIT0JtynTsbnSxk1D+oPYeHvHWPYnPncLitOD0vkQ4JPhOIX0iempIiD8c3lCv25H0F
iVDrrAsqu0f9YNihqN+iODT8+uvtbvIj6M77nO9ltMDvI7PZatpXOzLX+OVjg+3gcevSoVvO1AEl
P1f176CBsXeKEDj7d0agyZHeU33OhMy8r7LeVQao887NvfWQp1+lCdEt1gtlPeiPhZFcHc9vu/GN
8oIbt4s/F8TiSEShLprv7M9d0iSJ+rscpJwJ3acFnJYHTh6HfS7PewiteO9jHrh2tMor9gsjZBUz
mq/5GBIasifnO8E+KE3q3ozJGMKoiDP18b9chAm+Flow32pmPQsHTDl4lmoY2sBc3OulElQ1HS13
LfdEBNVBKkfhGvUe7I5OIiRh1VpxA2TBDBjNKWltLFTioJM31lJpjfAVv1AtfH9p4WjUj4xRJvtB
QVH9cYqLpVCtEU58sllEZ0Az6X2kB/sn8ADR04p1APoyp7FnbeLo81YegZdyQczG8yOuTX85IDtb
S5H2JwiY2Gi/N1IltudBVC6VtBOttRtQcbWwqtW30PDoeJTP/OnIzjsBmgXr9fubsgmFb2ql7qJ1
fNr83SzWae8eSYizojdRQWr8gc5fTr4ycSZEeVbu0pnKDGjiADvD6YnONeMEn1HzEH4JCy3LZqAH
5jLTDwR4cX5lcOzQN5KGNaxy6+lWo+9gRyiPFdKlV9l9Nl9tBPYkvAG0VqnUCD0Z8QP2NQJpIv9B
yUS7SoUejuIpDl6QRAG6NIq769LGgrCeKVreh5an8NjghXKecQxZ06tHDmmfx7l7acbW5sk7ZJiX
Xj73Xw42HUDZkgGxytGiIbJxn4k97NBDEi+AnjOGoTtIAQ2tWz92p/aWlWC4TRnM5ksjs7XtrYQ3
DqtOGEXyVgr8aQnl/JzMgRWUet/gXB7WkDAvllxLNviaK/ZDgBM236rlnSvUJ7uV3+aE1A6K79ix
YSgfcJ6syeCK1UrQWgT/sZPdY8imUwloFVz5aP/drADArV9r8p/rY+4FXbRzBFv6PkSHWBq38g+I
mQzVeLBoZ8Pmc0Gb4uA/QYosW6uJFcbBq+sKn61+vdMSJSa2FwFaPUcr6YEYq/895+rvGaCc7z0U
8tgWMVwL7D0GztFKue9Rp9tL9EvdZFFcgsNhzRGT8n5JPy/SmEDGhPAl8/Bq4Vu7HxwZzmjYXDBW
8p/BlMrM8H0qz9FVC1PLM57uf3BdZw53TW0yYGWrUjFvMqct8mx5YH8NstgjqtquHVYS4pTPuqhi
M7YhipIUJv1JaaZvAtrwSPoJ6MNsus6WQpsA9cMMF3pIBGfXiO1CKQP1EMq1Od51n1RjAiRkxx2r
S1IWwDONLTOiNzCOeY5gAHYA7VmiPsNjkhq2eQ1Sixwyw4F457/8XU8u4HCJ9k6mbOL4nrIJBvvN
KVh/dg6x/IdwrEaUr9Rg0iH1eUdC5/2uYMKF7Ilg314/Zh6QP03LARPmhyu3SoM07bb+G0OVLKLt
kyIdnBim+Z8yOLVb6QrB0j242Ev0+29IDdwSU5n2E4BDcMU75KsbDZKQa8nUDTbcAO9uAccWpGeX
ZKQaE/EaW3OU1ovQRwl40TxwmOrCwh+iV+0eeJVgiII3gPtZLPKb+DKvm6JUmNkEiXnhTFzKseOK
FkUC2floa4f26PLyXuDWskP3Y+ExyuSdjHcFgH9poQHWlpr8vsioJ+/KSA3N3tdcijQiLnIK3oXU
tj12nFwDdDfEIYi3euNecjMeOSzhb/kkpdoCxC0ox62nl0Hqx8EXEhDfoUO02mmEFAIHhfpyFwXp
4BUFkZPmL9/fSvBySQW6RxKeXWWViZGmqvmJjUXRQlmnDZbCkIODAVXylymIjm5hK3IC2PQM5OV/
a+gmX+z6SF4NiYDF9FwAsyqpAIANERS5+nu7euNlFd2nSWuU7EAErCr5bjC2IQM0s5YrSHp1UEtZ
otSf4OB8Tsn6EpWY9CeOe1c4Ln/Z/4jfoZW7u0HEjx+2K5LL//sx7ofmZv432nXhajeQqxppHoJZ
74xBg7JDG+0fgU7P4wPzLhMruBYnbB0HqATowq0TNbqu7Lix/4CCunwFMuHJktgMN2En2uDBJMbh
tJLUfS78otE2XPuziv0ORo2+oF1jIkCwYRPhnb6qBlCKgwvuPl8prMuK33zwONZkGItClQvUiAsw
vuuRErjrRWg2W8EtwigO3nHZV1GwoT314OnvSk5Ft5wZON7ADwbOws4HQCm0HjfCa0yu0cX3idt9
iN/PVAHFWF/PoJXKivOogxGy+ZYSo825sMiu0t87SL56xjyGnDW8H9T+HOS6mRhJ/dr87QreZPCR
QHMQLFlMrZXqEm9CGbRmNzBdM8V7cLLlxwySnAoN8kNrT6D7sdiJ1cM7xvxNMtcT/n83ulJAfS5L
k6t4IHJspZ0vyIddGYIaoc2d3xWO9vyirM2QW+f91Vst4yuhWqdsmF/2e8/TVw5xrIpkgDxCazd6
FRzvueoITgwqe/nHXYjsJqFNxVuyPdKYhVPv1nkMYHXZMR3slaw48tUGNNx4TRlNXcFV5vO4y1pv
3a+Gbpu+idxWY79jL89WM/A99fNyx6qpzg1YPWPKtqVBG29mBOO9w0JZz2P3jwp/fEk2b559qJJ5
PZZdMurTKKuIFMBy9e1w/8MDiVhJlp0+oHA+kUwAzy0iGakrzOpVYPYpI93Kn+/7I4CLMrxTCKbv
3egCQ+oqdE072Qqv+jP8E8P57rRcMMmk2eikYH46NQ95t7Kw4EyfPl7JeWW6ApdbAS9Sw8bAS7d7
4foxuAeLkbMt4TRHXwGVIdxkcBfHcEy3LQLeBN58dq6GTwbhe4j/nex/3ewhG0H3emwN8Ukou1AZ
R6BsBIk/u6k7sbOuQssHk9z4lpAdV4NiqZdTBp2qshI0Qmml5rBoXeWCfpL3CAxvsNAAHUTny/cV
U+td5tmP87rZ44YgFrz3O336zLmAUnbvDm3GwZNY9oYdWVY7DeEVAriwYEGEDbwjIvooLUfIDlg8
PXjzkNKDgEdGNKHmBwg/L/zjHsZe7zvUpqcm46aKC+3MxE3/cX6MZ6pJUcDyy3bN/Ug9nN34Kpx4
8nmRz7VOtZNC1QWbYKbgLc3GAii2PmNWsTJoryO92Kg+Hmj8mCE80IViAtmTYIXS0MsSjc+tmLjv
cbXLZ5b16ZQsSHB6T/HSTLbw+5xpzzhl6dLZWj9EMmtm6pgvR4+YedHT47CAUQ5QWzDcYF3nIG+e
OS/W+kwYlmgOXVJ0IDgS9CPlXECagWe82Ihyt7UOaSolSvhvPwQyFUMIdJA/mfXAyoxNcNpd24JQ
IfNHZ+a7e5/GSuo6P8I4g5oPUSNGbptjyvYRmkVciWX21QtkiAxebKOOJq2TnNjW4mN0YtYJZXOq
wZRm5ku0ZYsL9MlqEgNgpIYgBpv4L5sVODkOQyor6UMKzJqUeTna1BIS6Lzz57jeT7dfzc/C4Voi
OhD3zkNf/VodOsVEXD+k/CVrlfgpjOhSboyb6/fYeTX7p8vAJ8zcLTVekju/yYUOaFmvZe6FSp7h
5fu8aDgYIULgjMuP0HwFizKH1PMvkTTWiapXNfDfGL5/SLksrdAlrxuW1cUIyHUSBRsMNcn1kyr8
tPNcQaS1/Z9weoANukMFZ90+4sKsYt+NrrWaxpl0RLFZadEiD59wMkyBnVagZFtN1I+ufb9HjhSg
jDRikUlbcCktMQQB15Hlc1txjlUN6BouzYm9OJnCrJQyCg/XQn4fWvZfBu1d7p+HI4PEW28V188M
WntKcQF6n2kAfUiIPznCVYh8zCUmpe0BZw+gDR4iNRhbg/wlMxEXqaO0ZCEo3fIogWjrOe5uTF3E
A0XECFJZdIA/+0sGLblsGm8fRCYHfub6BXO6R5nf9fmqwndmcvB0HZoRmJL9urXlgH76YBMKnWFi
3hpNXeXaIdwz/Qj0ltTIKEp+pbj4XIyyl3jzFW4JbWCsdv6Cqhl1XLX9/GOM+37Ej/Ai/c09lnub
qTMx1vGI3hG5qZpo9a/REnRpSnzRTC/EfD+EK0pZEWpSmkd3/mCvPDSYGjOB2GhdYbbcBnZN5KY9
DLQhAIitvwaVDVOhj8dowuuIaBHMGYzz1VO5p8Ls0qhr70uNbsvT7l+NJQyR15EaBdMsSWtXXrzA
vHNEKUhm/MZnX4LJwFyDmiwXqrCd1NEI6PxuUSVHiZdIEJeKHSTBDYQmHPHMVgovHoauRlgirIkk
iN/dgWYb5AAAYVcnnsep6gS5AP3JbiI2SwmaYs/TDQWBh/NWD4Rp/Lpc4wzHikOQGtqNyDq/xnLg
jrDgIB2JElmd4X7chOAFoehUEZtrXfnxX/MO4qOoapTxWA+aRhafIYWCFTlpexGcfFT4dRW5XRql
fTR0G8DYM/1ZLCBCzzbk4/RmHOENisnydsBECfCcsH+Q8QKCKFswNgXBwRHayhp3VW0tFSsjGMV1
cP246ke7URu3hNw0of1VzAlZe/9at7oqElVXjA5SxAO7af9IdKhE8MKr9jm4Nzzw9QTpuXIznTp1
rZUlvBMJC8EDJO+Ca8A5kj+MRN4fNJg/nByv7a9OjdTVo3sUgr7jF1WJ2cQeSMjCHhVEFzpfjL4V
srXNCWh4+MP4mcBEcrW55zHr7+FLtNQKJ8xgH8vRLB2/s6g3qg1/15c990uAfCd3yk1oVvGNmoNY
qd5pN8Ip8v4k+XhuWzvG/NH4JlKR+ycUdkg1qe07WGAU5c498nYQGBVdyxhdx7a8VG1oy6ZNO8vQ
dVvyEVG0UmzM5qsSh6W/jKrpDFuCWAA67Tt3DOHDd/t4NZdBnDUGfBfytpsPSbFVSr8uyTymIGH0
B008BASaixUaCUsQ6VNJpvWLkhWtYTsldBjJsjRHLdTQce80R0aRhuEUxT2PBfWbmG9nSQJ9AG+t
Gh7qJ/BuoA+uUTbFqIHYMwIkl+dKhtRWEmdLh9a2Wy51zZ/Fwg66UalbZIcvb00rJS5uQ9PcFEHV
CG6aIrNOP2bZuwIENhGzSWqN0FjIoXOtNgptc3AOQ5fr2hyUdKjezeV9n4Tlo7AESwVgsmm0ZQf+
eGJ1rgqeEQWfBZiqFt6JbK6Mz3GTDhvEMTpjPo5V3IPGLnrmihmIpjY8OrFAvVjA7dybhjinHd0R
A0bA/gvF75zpBVQFsjn1f5fFYTlU8xBXybDMoKtmRac4H3HnlwptlWc1a2BfaGkdkuhshzgDvWq+
K7enamtqM035hQhdV6Lady45G8KY9CUzG1Yd0i0SDMuvU5d9ldejW2mlBwyRaUJENzvP1xMKJYIK
9qfuXlhNlulCpWdtEl1XlrtyJeN+h+nfyEKrozssWtCW+BGNh7jzhcR8paux9ud0/YoNa+BedcA3
S2L4+gXFzBDUvJs3o+drk4cAO/tNBbyl/3NMc2jf6kcOHycF5iP3W1p7YGyt4DAd7f5c9Iv3UtYE
89eQLn1LJ5967jSRCPIsxBhu7YDMaZZNT9hVJGdzaNJ+gf7bWS++ZR8QUA6xIe/G3jfYTNFJ3bhP
kRPgx7ANrpXY7XFGrXEvtR2Hct25N5moLoBE9Hl/suoljbGON7sTWTUpUJGwx03No9RheVevwlJT
5mqlMXw8tFmpimStFEedJU8kWBevMf/6cTPSv3k9DAXtI1HoX3GacHGs5LfpTDTETBH4WkOZK1Df
i59LwdZWydb4Z4IBFcZ8Iegtncm+dTtQr+TRKGCAidLwCia8KWPXVwLmLj1QwBhb9I76LiE7rznD
8J4alHyHMBCKWwd0bxGm6Jp8zkzeDDXP1/pTn/rFhPmxyysQETXd/UO2oUvqOWYjuwwmeIAi/xP8
8LzyesTu3CcT9Ntv/0O6w25PjJznfRW7nRe20//Y/THskesRJ5Gc/N73JnBLyIRLPoQ7zIO05R5P
hFJNNTR8LDiagLR9CXkcgmRQQfmWlcPs5oh/IxoAXrqthtGv45SgW36laNOarukOGdjOPOTMGCBK
mBuAdC8C4jHGU03+D03/O8dSBjvuLJG7/EEXgr83OuhxoM4UBYXnUtZmS4yP3plcp9sPBASGTWjG
KVU21z+dCzTgLET/y3MHxqZYx6hOf1Rt4v5K9TtqcOsB1ruZGbwMDlomHOyFGlqIJizlBtLiOFv8
WDEgJ5dX/MWruLyrWk0P/wYxTZWaLhhUrSmdjsQL88qT+AOmT5okcBFwRj6fsDy00xDn0T1pEd82
ngbdAgEF1XeGSGwq7W7VhRFKl5ePLoxVNRIopoYXULhpD4f1xb7tXc2jgtJbtWcliVlYj9dhRxlW
InLAHQ4/kk6il2nOUbAfbgRrtKwBWu7wdw/TkxiDuAM/026jM17TLEWfxd4GhqFqjHPB58QJ6IGk
MxfoCkALKNpSSjeUSMbQPz+kllJZRnqE6d1HGt0AchjfXYG0vtyPOsGumtVs8+hz5mB8Ow+wTzz8
eREo2pz5B7RG8tTvq1YnsRaS8HU/s58xrenwFBxD0tbZBvf+9Jdv8+gbSynRSYrFU2Q9RmtdtClP
0EtU969pAjAGdS8k9As/J6cUSEmr8n4Xv1oE1yN18OVlIc8rmeXylM7xgC/zGWX5fWdldzbNuAwu
97OhsCm6lJvvq/bEREMuhC5ehfs2NWn7q6m8yjmxzg9Sr6NO9hkFXw68LeVSpu4F4xa57UGge4cF
aHnt7ZZzCNGgL88aCLv6GNM1+OERk3M5fRZLQD9DqTvRFteGxMZ88dGFa7Kn2dBxjto+gJDKrmIk
GRqulrMJIAFX5ZdwcCbr3VTph9aU8TJb/ATwTQ+C5RROXKOaQuDjzkh76wAY3pnU2okXXxJaOp8m
TuGAfglyGsQvbJaL++2ljBmk6BZX8yR/fX5JoFqY8XL/wZFInni3wINZ061Mvt/dFqbaHACnAMZ2
yRKRU6qejy8ZFR6lo2EixbF0H7ITYi5oGV5D/8OXk7102A3vj/x+nv3cQ+hGkU0JDoSQTzSWAprx
VJW/kCaQTjfSG2p+SpDk8KJlOkK2l0EdN0X8sUhj3Bm/emzL55hWQotQy2RDuqJ/WjJmO//unrnl
Oc/+rbDZ0OqQP/IW1bqvNc1L6Bdl4vXOfPQvIwCn1NCsF3k2r7kF88+LzDIRtowFTj4yHfsMkDAE
uzD6AYKHEK/Yl3VXdi21hlZsVJM7C5pYSB19xerjo/F8A+S241f27aeFTma9c7GEHNzxB3FU/JAe
z+JJ7/syFNjwSVdJCLWpak+O8iBSpzC8oH2OEvhOrYBXhQi2tWjiWjuo6EIqVj6XC5CtwxpZrKrc
BLJd11zo7ssUMLCTxl8pZrRSL9luxRh8YDDKzRTDQcCAOQAdb7QAj4LRyGbcfRN+7tchln3BHiv/
+HNeFPCbKmWwx2VqeI1dpVzQpoOXnsfIfjw2qRiA42T4CBItns2ypsO0KBVkuVhTo1+rkhzdFRSy
hcOLv22IZW5djOKt/5yPO3EdRLUN8eKlnqfa1tmpqZoZsyjZPZlziaImzGp/HZyoTCz4cTXwdJ2x
t18EpoJEe/XcOEbglXDs5J2Lc8tt6GxwkeEFsr7Lhpn5jbiFEmH5geJAO9oL0PNyQTFKmQUFRRW/
ksW+bgWYLvk9i1RZB67jOmwCW+w7ivkr9LAFAJyxuqj5YGwGqX9tS1it5tPnLAWk0itciQldas8S
swlJrjAtF+q5fL8P+n0vMy8o9RO/YlubRPdgdRz7z6vS2yV/gYLZRYjszlr53AupWLEEeYuKOQ/M
hktXeem5CMp5x6lOfPE4fnk7E8vSmIn9uHdaZFVv0XVrU8Me6OF0xQm/kG0LCMeD9MXfDiIRRaNp
CVCvvMu3cyK6A9T73rHHZ4sR9aQDBm1tdujaCAup54G42CeNFllOW+UEV6xi+ShpUpe2MGImIM7V
lrOK4UjQtJr0Eh3wiDTgGY1tD3gQjUjM0q9Huyi27Xbx5aeqFHCPQSNjkPE6a1XZsm6CZcwgUFGg
19KuVRceOw0ZMyLAlwz6AKJK8OTf5COcydcPBen3Tt4L1y9du1nbYEFahUarsMm8gkgQoS22mRX3
Qb0OLVjxsibWbZjXt0APxQa33LKuts3RwaFgRKbp9E0gzdPvtN87cRrt+A5XB87F2ON4PGub1lga
/nQdGQXqplld7s/XsYpEeIOIrxw1HPWcv3O6oO8zFDo6TnvmFori5avYZ5BnmamHvr3rtAiv+YQJ
QIjO92VPP3K+p/76grD0WUQwY5tHWNFBlCKXixeNJ3KuMdPMhfjfS+vFC8q5CzWpUT3eh1AVhCo/
V6uf/91Awj2K7gn7BIlxLoog9lm01ux0Of39xoXJbe4OPjLWgAroOP8lg8H48uUV/mMf0jdUXAiB
tUnoSEJH0Ae2Itzbc7x+07hXZM8RxEpxa/ddIFtQVTkL0C7ztnPs2J0DOW5Hk1I5qpgJBNL6NJcq
XtZpCWzg73Gf64hxvJQH2ixdVuLFMnartEiCXLNvEcvTWl71ivTLDnKIOvdmRtCWsunNSNKZwUUR
pSBBqq5YlFnILI+kSTjkqt6rHO/ehSZmCUHELMFCfzHa01TsvdAO+Nb/TpwgIHb4JQbqMgR19aWq
AH00pRZJbbXT7pDLQNqXblt3Ej/4jw1kvWN3n8FU0ziMyIKMtC54yGGcyH237lZALNPY/h5N/ZuO
yzNYseUTqs63xWjtdsydyAy62rFL5IlIk7YpWG5EJmvAAPtL3ezns9fvAY2JQaX+VmWux0QlXPPd
+KOdDR8ZBB5Iv6WYea+6Ia4FcSmgmUOp5Xudr+VYWGhSeaTbWHdks0egoEXI+f63ToJQdJmvuz4b
QVnBD0WJ1umG3kKVQwuXPq93HVsHr8E0x7cuJcTMVarp0JiRBEGVi4VyC/pP/4eMi26EuPoP191n
WuyniOjuFXvqJGdO8R9BFOYPCLaHr4KGtHdICMUrglJsxytDII2pvR/t6dpT6/6JX/jYdq9b50Lz
i2c5al6FWrx6vZ7SffIt0V/3qnyjD5FdtqBFspBAh1HY+nS++AnpSXmIxbFHfIM+H4ZPbMzIz4yz
f3StPbW4YGF/JUQgLQT+k5mNd9HveCftt1wevz/v4WwxMk5dbEiowAii1jPEjE3JbIqIzMRwIANt
dUiBu4HZdF7hwZnYvv93xMoAH9Wn+07/Xq5264PPce7LHGS4whb5UFBmlTJwYLZy2gYciJ0mWTgS
fnzg6kVN0os9AA/3jN0Jh3R29g4Y0adAswR8S6bYnqY3Stnz1K0Llw/YWg+oZqDNwjHTCEzg2Up8
Y/FvkLwDedYmW3+Ywp3y64CDBTVrDLvLyneJQyCFo006orKe1oLCvVSH/aqHzCr1j/BtE6/kAjcV
YfHgT9YAtBAt5jnB7xD7X1iN5TVepM41gADYVPgxcScu6UbaIee29fb1ajGhHo3q6dKnQri8wu7I
XZm5hvtW1b5xqRUOPOFQThdq+Bu0fz0p0mO7avGz7Fv7/7ReBsd3x0jGsJUrATyptJh429mb0sGg
gtt2uX4NQnGX9YM5Eg5ociKs165EU2MY4eZyTeb9KsS7qe8y7ZpJoq3pEYkWp7ex3dgkvKb3fXIy
p5uBbqP/BlnaUTO0iydlRIu5fm7DD2nmBFMvYUtXHud4Wp+6+goPAcueXm+cS0VZNVLziAq7aus+
OvJoHTe4iTfE6tK2ycj9QrCxT9BDaAz77e8U8KE1Q3DO0U7xCcwI6BqVpyL5z/bqSjmRour8FHhx
Jlsapoz+BziBacyRWpQnjffds88A26rXO6wGPHlaBdJEHk+9MIzPcai568qyjBY9vBr0Xx8lpbXP
xvglJQPC1iFJb/wKmz1eeJr1Z6nK8lz74e47xwtrERbfn9+kT0UrCYZ33tjPn3lHXOLNkIRcIJfZ
d4SEecRaheOTH7af4YeNWGZuZlBLGNzQi+cg3G7tK7tZRp3qG1fkG7sBlyEyVQm2F1sZzkPySq4f
wqTjjcUjqUHoMHQgax+wcvyHPbr/q7WnA7oJ3jlwTxJIS76uEQ5/M/FfQUzdDgCMG7a8AS7x+b1g
IuGqeUspKjKhAR9OfdbIsQ8gfdtPrbLzqEwi0OQykwCR02e6OKZ4VmCkFyZ3qoYf53uJjSH8BRLy
23Gn74f5uQxXNFkm7u5KdiGfbzgk4plak4BpBYlE4OGvP6g0nSOjekT4mMGA3JKlYDk/kIkDrY2x
B18y2slLUbymDmfYj8ovZ0eECEORECzDwXF5XPon0nY2oUqjoKf8zft2lNWoz179Ve4IpryUTlGO
o/TPSOCRR6wmNLQPy6vxMZOKRkWG/Sm8pTTMMN6oxvzrP17CrAVZXwYuLr7CyEWwiyFGP+36sjJ+
/9v5DPWFWSnPNEN6SGfO7XWWQlvlAR54DnsMitTpM05f9jvaXgM647mDiUx/dj5TjXhvfIsvhRGS
iViUmDbaSe4FTpZ1kVkfBcONffiPEZCujR1mprDshwqCC5OoqDqjLrauUKq7azikLbc2GIxfxUDo
JIiYZf8R/seYV8WYIJ7iQ6EmfS5AwxJZqfn8wRqdmemTgsv84fwoSOm6HXlk7doIJaZhtOXLzt7R
IcOotNJC87eDlnHboiH6feA/Ik37niT8SyEGhtdczrxTS10bEMEzZou98vpoQiksiHXqvFZcZlXm
YxdZ6ohlDsqGPCH1NlXbb1y5DPlpDmFix4GRGbiGeyi9+Pn6otJxR8dTXDrkSGfpiv+0EUUglsof
ActFqsLE0+pymtpMThfRAtOGh07VIzWXIrg6RQeTqpnpoGht2NmtNbcjAlvQRUnqgbXr07SzSoWr
842RZsQz6Xue//chMV2g3X2ga9yZjD6nft6p2PFb/4ea4xMnNRmUEEquoijUJMKZR8+xICEonn0J
pAi2o+zWaxFo+WWjKWdzSlmlo0T/9leI/h3jaY2JyhldeUh6mc8aXi2syP5v2nxCO6XPul2i/ycL
ald/Ul1CNaLB41ea/ZxyP71KZUGbrLXnMICLjMRzDB08fsEFCFoHeJAG5hP0IlcxdZnqvBUWtsam
tn843vtnGhmZCGVrIRMsajWWSisxKb0KQ78KuwD7AUOLUafNe5u27ky/QvWFfy3NvsWGC6A+GQsR
WSmD5XI9TEdtdTbs6pfoUAXs9a6795EGa3MLzj7SHda/902jgCtvp1fy7QPcfa/WmmuI8mEveMUS
9i8BnJWg/MEXqwlQ2adNkdXVZdVhQSc2HLibAyXHDCH9j/o+l11G9tqL2m2FEH8O8T1fYMMsNg0R
YBfDTPL6BdjAUJSIYL9oPEQIx8kmsH8SR8CfThOfMFWN8ADcu1dBrcFdtqu/qnZaPdDYh531cmsq
IbEJ/jt8rfWgy7UUKBMi9HXtGCRJoMWtzOsDSeNh2VS01hkID8ZYYHDc8e/t32A2TxJIYfkON8KP
pt4J5dPJfjQLdPXf21p7jWxgVGO/GklQuLrAntWJzDPJUFM0m7nXVlyW+57rmwCD+footKj5vy7O
cWh7J9VFehE92s0b2P+CBmbXc2nV43DbUWOvsSegUrI5ikcdDgZNNFmCKdfeu21+cou7WeJFXQSr
HhjbDIMikgP6oIkLwhML6RNEgcLDEerqxqlrpX+d6VQlXCePvGdYuWdzBy3b8UESNiHmYJVOJ6KI
r6HeFABx1pWke7PLMWm5D0BidEf/TFk6ARM9jYBHqpMWlwc6y6W1tNRumQpmsaWjS7xW/IEAphCT
IkFe+IfgCLuH+cx+NlK4QSKu6uf3ZgML6RpoIRquaCMUU3H4k75sV/SMFvMkXsVSd4r1rHzxJ4gW
e0mDJtCFgYzjh/3AUZBc4yqVqpzvnSWvaSgaCzTn6efijpj9CrqAvSHxba+B+c4dS4E6NDDT10Gk
jNyqxWzZnHUNYesRb5LBpIMZZ9JbxIddfCKWyVhT+wq2Ua4WI6txrY5WnRcUMg4NnQ7lk/xyNVxX
rZcthJS3PVHirprN1IGAjiG8OxRh079c6MHrUizSxOVnB2K5ToGyf93n09PoUmLBphAbBn22KcQH
EQihoyct04x0BhUNp7ZpiSWMwwviVsZQzuCDy5VOiJcUo2MclYAI3cfPRpkxXJ9wUYXZSHxUSgwU
Z9WX4ttycMtNSTlu7D1GCQZW8AMhi2ymq+tQGEpQB78XK+Rs+6G/rR5OZMW6y25v3iR4Ct5YgoXX
MdHwd4bwdgwK1NkCNJ6KyeZF5IocoblbcRO/RmGvupS9BlJO/UpprHUK14foXUedghjsJRK8M0X7
70cVe/ZDEiJXyg16LdSRx26l38skGgmzH5kiFOAttswbnd7OrTWTRq2xoiti6zoCIBBM2jW4almm
ayBGv2oql8AX0L3zZlJy3rF2C40pVAETXFviLf2GQ7wrY4XLsckLI6+60qfvlUUIFjvBVD10E9mw
tcgQD+o3uYFU4cyyH5mqzXSOGAtAhG/kPBonlnOXcj8kUMJUHRsFGXuJ9Wx8p1nXAQFbmpxG+Nc+
LWm/w3iXqLFmAbsvMePmxbMZbt8ZDgXqTT6zhiNxAJsFzlnq1ozxyEmzl1qIEb/+vH5yFuunF86t
k3EygPUXtJ1987+ytEI2VergNiMGBJqKt2S1gLdVQaVV1S/RPAs6jny6gPeEYGr1otnTFIizVZzi
kFA9ZTa9V/7G4YtZEXhr/hSIUNB9YF9L6ZitIlimLexcqnnFogMuHkqktKtpyH1J7RwzEZV+qzrW
x7tq1S0ZcL2ZUBiALs4IUy5ga7Wg7etW3gau+XY2tEx0fXiHI/aIHKbsO+J7j1JMcAnGupIOxMg/
ABrsBUCvwb2gS8VcBdsTzDA/9aa3SZiREIjpvi9mG/XQsMFmjqS4sdfJxOhwr+ToGDEuhOWruD3n
4VY3Y6YcgxVcZKFUve36BfZxBphtRziphbWHfw0dha2Wf50IYXAkBVQHbB8l3IMj5TnTH2bv3+Ud
nkYbBUFPmHEVhWfK/LpSGN0ZtF+1EakfWgRPhBRLu3DeqPZ/7XER+NJHVzMChaD8CJOi7xo8crsS
kYxcx2+CTgRW0GBeIKaa0NURsotKysu58v5SbUdNy8OpP1GXZuv/T3FCSBqOjqq/XwLyDO3yeUWI
TFNWT1KxpSb7swuctNmCSqfP9gFIQ6coe0UxISnWifzno5xVSX8Qqmiu67+gjGHYGhKSpbYUnVvt
p4h66cva+6nKqg7n1YAxLr/US8FO89aYC8hUmXlg5TfXSfnJh7k9cjaWNaMpFmR2P0T6gDA1BelO
Np6bCN1YS2ZZ5Mf6nbchuK/8bgEWo8ImPVtJ9FDge6++Wmo9BMxLZbTjiVhnpBB2pol+jXXjyqtI
k/zoCnz6TboDHJWkFPrMBybxeH6UPDSfSIr0UB94lGnlbWbDNPONB+ss1LEKbRLzOMkjAdfBVDtC
10U56Qn3jBIWgZRX1pLpFezj6LKvDSBegL2kGltf6ln67fCiPHPuSnZv/U4zzunPlT4vES8u7l8V
s3HR5YxvkBNRqyvtAoWKqEabHo8DSjVFdaOgwZyebERvJDU/Hd9FANn/5Xb+hsIW98/U346EhLgL
onR7tQ3qqb3VYpxasUSUBtUStbB5aP/spGDwKrnNGV9lcL8fhypYr9jygzI+MNx5wa6xFI1r68+p
0oNLPtlKNbzY1tXdCMtMBYk5018bHCzFwS9o4Nu9EpUZJG4qIeaOErQ/tz5EqjdMszKE8XFVw92H
nDtt9sZQ0GkHGGZCbh5wHNlv+5fnaA0i2dZjoZ+QSU1LknLuxGrxTB1W+3WYFVD2Fa57jUewzYA/
Vb39VEsWVc7B7v9EtNgu3kLLo0Vd4gZNe6KUgm/lmjlq0c2LJ7Y5Bl4RYTcmxW5TKvNDoF5f2fxf
HDjRsRkr8Y1UMIc4jIf7re1APW9PTiP21w8sLoFzMB3G6GM3T61OGxJliko4EPRF/oyFrxL2VbCl
rjp/R0kq4yXhrx4B996E+pNfrHmg0LeTdy29W8mxV2A54+z2rDogX1Z1M7prEpaFBcQogMg75poX
HtRrecY56+NrZla2fu0xuZ3bMPChOr6G4AV6eK9pgfA2kloOH/zJavb0Y74uGw2GcP6iy6phDFO1
7A11oN/3m9sos3aEHY8jst/p84GyWrxdPX9xDeYjnHSGeOT5XpQQnoyX742RgXWEJ+JYP99Q05e7
ASannSdw72MMEWAEzcOgfN9P2bd0uM17knLTDlk9RMFJNOjpPIV3FBPTaQEFVFpk+PtYu8T5Ai3g
dCP9ABCmC0hXncCLjT/+6wPAvFFbNUYyOPdkaEtDgYzyT9mGBvkh1JVcZn6Y41AOfx8j5HHebD0f
QF5BXlPqaBRZUzE0R/15/Eb6/g938PIbPrmfVDScyQ4MScYpxSCWRlIhJFjJC9frRf2ZHEpdCumD
Rv8ah70JzNsjS5+AdgVrSqr8/3+1S4LFzDT9EvFKpmCwVS1UWNn4StNCTfXveJGxonm3U6gNkfjb
9bwDJFySwCIX6cDCs+GLgXlYR4pafiknrArgvnV+ToP6VEzFXoaMF3shLxSMOVoZZzw2awx63ogG
Za9pMqrOJzMn1iL9n31tzUEgfu/3254Cq/cNQaXrZeB5GLleqqADoRGLArNwiqNVsWxGyadbCpek
S/9nqK8K/vbrJQgPMwZU4q5RX1p7DIrN711Ert8is5VrsJlprN1Eaq+8vPBG/qoNG8xeDwMHLl6r
g6klEYHF1ilUiPNRZ4t2bGJHLgN3/1Xtp3DzAsIjYz0bm5nt4vQNIHtvOkmge2oBmK7Jsy+MIwv6
+Z0sCjUpmfB4kWOwSmAS11Sff2Mdz++AeZaticVmeBuWT3nX71l0qRy/rnM+FudqREgJ5VEzfuPi
SJJyKZY59wDS32W4obLPRPXEvbgaFzEhybHR8KMDZqlaLrB7qPuBEPwU+thAtXJlym1PupjqzsRn
mey5IC3stG6/foZ4bdw2A3tHa/aF8rL2x36gOvgQLimGBg30JYFKAEyc23m3CnOGfogi/3P9cNJV
e9NkqHP9GKImC5qZD1S2n7jGRJPYl9RE+ixJVj+nk9xKfCILyXNs/4JQRKYd9pMwuTY9Sa+zmvWL
VMmyd9wpDGh+e3jLUW93DDPQAxP4kLKuyUpvgMs9rR0vQ9pi7akEW7Wr7IP7k0eKLfzsWrcuRLlD
qqNheGUgwflY8oCjp+Y6ZI1FVISwSdJ2EFKnZvA8xLqUF9YNcJi/vEdPniFO7WL1BK9eAVxOu/Yy
SipKf0bT+NwIBOGt//+9PPcawOgUpsIftXZF2rHno2pG4NuH3nPEnb2k10EtcITtgi1LqcwgIpr8
OLKwAnDLbtUoghHVGtoJjapgs0lEeXgJi9Dz3RBLB7tFzdlxTI50ZowbvVJTNNu4+wNyzCAVTKpZ
KSMaN/OHUT949BedybWM9J4+dOmFnv7FYSkQHgx/A7O1uE4tRz6vpWKNRs2n4DKx+NstFX0qq1n9
WG0VNdPaAqwZZA+G8Ik1SwZKV0Oa/pA8SoDqBQ4NNQs/1i5/yvh3x+tB5ivK9ZWJ9YIsDGxQBCxm
7JJtE8ge0b/Rs5JzelQ5Qxpu8Sus3WQe48Uyq/EQSJlOsM0XxtFD/tjV3/EHhw1eC6iU72lt0H3y
3KNH06n0dwBz6xiwh/P4+dXsAIDXWXTgCiiZN0upkoqmWNUJOhkf9LBfqovE/E2kIffHDhAjL2lE
OVCDlBMc5x8QEm5ZxYcyglhuj9mgmeTgkn01bFeoyhfl3p2MeKWKvqIuBHekHbSRO45bmdiiwQgc
bhr1yM2lmvK9D4xn3M7UVkFgOt5dZ6cP4XcOR6veHy0/rN48v2/ZRNEhNJXju763CgHtklU0HtYV
6Su5IkrRRTyLpuW0lvVfJDX+Z0ZT6KoUfMKW+rscdAah7kHcyc3VlJ4uzq2sWR8j7hmsBkR+XJ1y
qVZWsuL0AEkcsteWaAQQHHbvrtkEvbTVGH//o6gIP5BmWQRDCX+B64ujm1ReCpsufT4xLZVGMqep
1+EacLzzrkDGCrSZcRFfgR89phpgAl6QZMYBvsxHdBNTXMYAA2pdy1My/Ai8N2xPJaXdoX2qIuvN
ao4/4F0vo9DUxl4Tm5G7KLQ5o+lpSPLxaPjWKZx55nHbeN7ysMA+Dij76vgw/TevpBwIWwrd/7rf
6rZLBktMoAspeKeLvJYMUcrw/NBuQX4CUvROoonkVfr9hJ62h1Sqx6tEP7J7O6EL5huH9nH5nIMY
WnVFk9iK7wfwZO7WEkFSnfRyMkzQV7mbpKHkLrV/4jB78tSPdeOXyzTYTz+A+mqT1o1GVxK235e7
4Gx0v2Z58z5Uql4y+uz0n0zfYyMXtLWCNOrPipmXIN3cis9JCakS6KVQhr+ionGAtTag2zGhKjkc
0PrjnnoUJZfD7FhFA872IwppeNVbnh4wH0vg5dtp9DMxY8zrTMyHuEHnOEq3ijRtLEfTEeWsm1Bh
mVi8r/eH9/ab9iHBbwu2dCT3OJbYkVyqX7u0XCbN5UgsEchZCzSUQpjfFG9q68rPihdWbjBigCUC
TQ4FxYMQYOBfiJZGU8flyJJx2W5HEBFAqguS/YuX5zYR3bm1kpaMpwTkVlDitLLcpmV3tzJ5rCmY
17byEVGIcyf+oITdeyJZ/EkdWLpfcjvyL8vWwbpyo9/RoWtoFyi1Xpuy4Ib3FhNPNbuuS8uo+GRe
VTT8xAd7CyCo+GbFrjQnjMYKyXwQgSb+U5/IzPZAgcid2qXSDkeZS30u7tB3W5C24TvI+0lRglD2
rdGypzQK6L3HM+iGvxfc0EbA9EPWFQTNIeF65Cj2vWcPX8m+28yDuo7J1Oo2zE2AWU1A0Zr35xgA
QbisP7PfeZZ4FHlNFi79NYT/Xh9qFa13hJ3chDS2mn6dAJIOVxSpLbpUJ4pRDidO8zYe5C+KIh8J
Ble6aNyvpRSjjadGf2cGFr/HG9pVTS2RRVVOrsH0lYgH5PRtu3QVb+CsmK1xNfeVmGuAn/7KoBIL
8ABkYjAYi62d3UPm9E37BxEt3KHLQq2BA7wTrJVfYZxKc5KWLwalbQGM+QtbFE6RgPLETnNlC4gh
QTPbHHRHtpTENpjuIvtl6E3W/djVs/x286kAR9m4IQDj5LD8LrfgG2CseJ1EMDeOq+Jvfk0UIiZp
2T0wbkm1HCXlyftY/n2VMB0ZgkQD3lZ9dw/MsbjmmzQLS/qc48va5E/53nSS4/IU4HUcpYNZUnT9
R4tL4luPXY9O2eKj9V2qBxxW/l/xkLb2ntFmd+ZOLUO26CabtUiJhz9iDC1S1Ktr2WgT4a987L+f
gP2Xk1DTFO9KxJRC4c8G8IxHhkh4oJVAdnhK7YNIkc5kRZP2RDGs2XqgoVXL40I4Sa9y4PaHtHpE
SncviepzxsigMH8WwBJM+7Rp8DRHY0z5uVmVEszKbbABEba51OhZbxMtx3umf0gSlfU/qiIWg5b6
mmXv/+H5gHxgW/bJRUq3Q8nL0B0NszYczRm8BFizg8s2ID5srnmgLYTlzVFa6h2BC6gaIFsPYfXJ
lrPUw/EZM+E+1tZadthnrnjg1r78CMNbdagba+5Z7vtuv6VE7JCWF1GVadYri8XKvS4PHeEoW0lr
/lpbzQHgOHqT5h+FsGlEUu9W8F7jgjB4x2s7jWhC2r2FIeZrxs7k4MxH2CiK2nAyfNc417Bvd54F
wdNUqlIXCdyma6dZJfhALCDaSernW9QUohrkZgOvj0fA9FJUdiB5iP8vuPh0Ph/AXDNhF92ulAr/
L56pyKYdW7GIDhLymCFxlPS+OYoW9IjU2cvZpuhUS32QOpukhvxsjDUhudIcxVlboz/Qp1WNuZBW
0PmIC9Hr5vmjJjRFzI+0yvsURt1pte2XtJ3xjKPPq0B1Kri1oyu+Lshqp4H7AnCitMKJLZoSaUoY
llma/fp8Jho59sG/ZOzQstJAOrOyvrFgkffO924fir8gZSJsc+XlJ4HLSH/d+Nvrh8VlrytdrMSw
l9cvJw19cScutReAVnZlzfSKpLrmcsFwb+1Lwccc27+14tEpCfTHgBJwrR6VS6m5L35SkYhSEnbv
ODLj60aYnzx+BuTBF770rEQbzTtxOpftMddvl8ThTM+kqejMWIZDEfy4UIbbTYmb7l4YQb6mUJkX
BayjxSlJtA8VefKf6RpBUrjDw+TR8N+1IwX0BFtcK/QXZK4VQ+hvYn1vgf3drbFTOMOBL/p4hsXp
tDYblJcUMSewY8wiu187uOpbAQcSX7PXwitq5jfmcqYl8PoozkvN2bK0lupGgNCzIQ86Scc9JBps
kJYKH6+dXFtJepGNQEJPznktIs8xdzhW2MIML0z3n3B7lCj+/hS4HOFhC7BLX6as/4nlixqloDY6
mzR6HJKt8ItMNc9jHbtEuGI4c0SpV183zj0BwKzwP2fx1+Ezxq3rwYZDu19Dhz8TEYFBac1NnRC1
aOv57G44jv+1HWuCZDQLIAvfeoc59aEYiMKct11v6UEN5zorCKO4nRzmEAU5vrDPHTujiAgnvi58
a2X3sDPOY+g+85/pyKDE3X/LGFHquZ5ZjYa6G0uJxKgRFnULmH061ueS4/aGVo2F34aIvsnrDvOX
4Iw7KjYTJKEtqvIQ8nj0Un18zy+Mz36lVWFSxvOL4rVMP85KPJsW1r3r7O3TsQutRnw4EKMMqbKU
GkrdLkmOX19cB/FksqcfSnXANG/X0YNE17iCDhfDduOuOFlq/mqk4YUA5WRRfU0JtUaXuOdgVMlU
juwdLGvSQsa16x3r0mT2o0ptucCuVMUR7/zgIhRvqsouZxHXRYNSM67EPecK47xul96zX2yid6FU
7Pmr6G0CbE3m7abBv1SW/QpkPKyZVOYQb03msN6x3JWXai5D3Rg8yU0ljqMgtHun1/p7Vl1Anw1/
BMV+7DRrOfV8R+zVq82AJJtOSJLmV387dTripQGNRBwxGiV+94hXcXRCOlPsEmJqHYYRJLSTaIT2
e+1UXe78Y9QbZ6hcgi20mlUuxyRH+6QFCxoihnBnaS+6st1x6mJ1rZYe3cbNKEFFAF2fkQKXv38Y
BP8dzB65BMJQslmiQhCzorIb0vKZW5g4PizAXBZTohvmUz8VJPG0FfspHslOWYvHugPZn6TPcNkR
4/oVFjwm4kn/YGolPn+gmLTrrjBrBcLl8vfi8ddZlRrAlfdd3LOgPXjZ8sEWmO2zBj7iHfLuOgFv
HV1QHWp6IfS4Xq0NpGK4rGgSSqgULPpofz15Ar2IYi8n94xr2om/WzI/hDSIsNxYd4xLqa+F/bMp
UqMC1BeMozCQdLt8Ta61cijagOyt/X3wGxORZZjRyvzzm5HvarwS1KBsjWBbGmb84ZpeajPEhMd/
X0M2FSe0ElWUtWJI29sKaOWU6B2ODEhUbKS4s19GDUftYmhiw9do2B9kUNTPTKBds8XYu8omTqle
Z579hIoiYtzggP1jydGvqhk+LM4UMtVFVKefRBB3TUr0oZsdDmIRioTP6PLkOVl5Dmoon+7FNFWD
RVDZjos9fFLXfotPREOheqiCOkdZyuv+AWAklx9sfiaYNJclx8+5vOcPhsVgmdIInLoqfIxU+mlZ
XCurh4C7hsgv7N+I9kA7RhkRtPSzUeQ8HA/+Pe/QbdAPHJY8VVQGzVGdJsssO8bTfeN4jsB2287R
kRmn23UND50SjkCWYtNUNNXW6xW/uHAy2AO5oy7FaHS8VDpYAdlPgCXtoE4uyOsyPGlEFVYERcSG
ULbmyRC+0KGi/ug0n6ptDWCymKS0Dl2sMoFv7Lf7kMY53LfwHNQgcayPhsarcE/hgs/NbMiz5Ekx
op6TapdKf4EZj3kpQL3eN9EVtZTm5V93WWy1Cxj+jVvpbdIXBEqIlmpgMD1y2KhkP7Q++8/s+OAT
vmrJSUXlN+BrHuQ+b1A/+b2/4VW8UijdCS+vO3huDda43Lo2LZACqmblhS1mTT3sD9cLHBK19Fji
DkmEGnzxUsOOQA1Z4SHXChKA9tPoPLjRJXr6c83ZRGGBd2fcAeDKwM07zFLWQD74sRu2EHdY6/I4
DhY2oMJkH5F0ns+bzNJVgryyXrSJfnLdmz1Zl5v2IV4IK+yUArsnvkhieaJZrBmRBAORlqK15+Ok
qvojsz7iBRzYr/KIHAwSlyK6JcK3GUslBZZQcosZaKCMPulxBf10OHRkpKxV56FirxCbhcJ5R7EW
pGt6uEuXJcJ5BLJe05Q1I0cFFYcyP/WEvv4X9JVho4ITVgVJKD+kngsHV+i7hnhHOC0KsPeUa8aG
J40TOYAhEF5ZUS64xiFn7RadbroeVDXtvSGYzkDVxQ+gEV5UxsimaQUtgrh3QSLSntJqKGhkQqKU
wIIFHtY4TPxwWEcED9VSDVNTyRMb4dQ0+3r5QSGeJIrAZBbSlLa0pyj1pkogWM/WO+WKHCHSe7cE
k+RfFOKrFft5tgqLaelFGlxTLNPcl6JBrhSOUb49kdzifKl6yFmRTXt0reIkDAczB7r/EfGFCtWY
OlS6OrexnZh1bT313bxgkxDEd4o/XRwSzcWydbXL/Xpey7UmW/2VyiInDScQuYHglgkzX0uyS/cU
Ej+gjTpjdKjHySzt4ORy6LCWwhPj3ZwoYucFUQZq1Ym1xvqZweWr7tVwrxqit+tz6yPan7wlbc0m
w/V/5ImOVK3zj0og/4eYPGW9l/AK+NTOWM1ffm6bee7Ue9oOJchYyXI/fW1mmLF0zLz7FSIRw2J/
uLHlJJbfG9Fy14qTuLZasDFh4ir0qJGNtJb0kE9TXaDPESYUzUEHKz5kq6dFPJlyMpV984AuDi6b
VxgiYTE6tdY96KJ/KIPHQMYeBhY4xXY0Tkf35DzGeJEHaaYfQ+zgc3uo9byf7FoYxYCZVugbLp3P
5ZKBg3SWX/OLVpQ0+fDbEk3KTYUwVdjJXvFW/QroVDCTupOgO1A6w7R8gkER22EChPhXTRO3tKP4
NxujjtWi78cf/S28AMER6kfv4y5d7f2MI06sP2uTSGrHSBZJhfI+ptjJceCreOwp6ue8IK3SuLD3
vsQRawx90eLfzO+jMDDDJr4JN7KyugN87SflT7YNMrwI5C3gLrl1As8CoKjVTaGHb5U0xBLbFkxC
KauB9KM+afxXmJ3R6jlQ8bmyZGRc2sDi1Ft54QNRqVDLq4hghcOdJNr5MbswpkXVoDDElr2Gdbms
2q+sj6rkZLry8MIcn1a/vnNAA8PzmbTRyMK1+4tA0/SwDM6Z+W+Rg+bQtst3mHIvWrPJoi+L/oD2
ORSn6g1bDyVL4xiWWR5sCSXEqZjnTvcJBeICdXK0qqHDHuHO06uEKXa3jFRHbQzSFNmzZh7bxgMD
44xGOJe/B0dL65s7pc9p1f/Q8p4BVBujhRkAvMYwD6ZQnYLvCYutXsQjopWewbRBgLyKM/sJ99gR
lyp48snF1P3UF1jgIWwJ/+08vLjBY9MMdVVt4ZfcUOb2iVLpK2EURxZeDYddysvGGUvkOt69sOxi
IYzepy7QHkEghN+e1InR+CMl6fJfeow4RJQZCWMYjQlcfUSh18M3J7PhTncZMU5qWF5TCAo6QkHU
GoTaodchR6P6nhn07yItPSRsr6UhFCLtHLZWPfsC/y4lLvA5UmjYQV5BROSrM6MLq5t19Ki3WwoM
NKy54H73E/IJeYLTbMwvm/KiTDMa42c3Cu/+FIv6Y0nMMLKuvs3iExuJNVtt0Vb23AuFe0svbtm6
x9dgv99jv5Vb+lJPnS6sUMkRJR/Pb/plvC6z6pv6Fns/x5btlkgUAMSBsOfW9pPxfRgqrTemBVzM
7qZWM7ynyoH3FJIh2J811SO4UHsskIn5+ugbH1piqtmanPiy4DolGqhzxPhcPIVGH8panlnS5A2F
4srpR1sETR2tYGbJ3EBhYfWHxMuoBIc+nmASovucfphMiDuqxZVPgD1CAXUhpYlNls3wmahclrAG
c+HiaOjoUWBkhyRNe0BLQhc657agLbNejgwk5Pm7o/SVKywjS5JS3OnarvvWir8uTwaNc81MB8V2
j0FrC912OKjAbPaIk4CUbNCye4AkRbyGTSqzTMXpORdCthneWsak+Qr3zgpwAN5JcXuS7zbjjsk4
bEvXpJmZRfOkyHrzUig0JYpZTnxQqvkgmMpKHoJI7UipicZBqW0CZn5eFhitRUtpuAD8Qns4UakO
pKSbtE/WDJRaV3nvFeSm4Rmu1EVrpwxSeVql9Tw5BY1GtP8QbWMudtsUskiDjYGlUVYGLynxpsWx
owSkZf9VMiyg2n1fee4SfSF3yqUxqTcnt+EPPW/ABSCFP0XhBCtWoSs5Xe7uULEsoccpgzANalfh
N4IHz0ecP95JAuMkqo9Z90KsBs/lPV//pxubHXLu0Qwh255fbu0cRyegTeie/nnZMJ5txo3CQh/j
GPXLlyhG//xSm8+sch8oui12poLBIA++fUxilbXDFXMkKO3jvgxbfW4cg8cjWTPlqkIdvL4L6qJN
lAYSwtWzl66j4hOUnynv6iNKuvNqArUgDsjXJ/06BlGwxhP54UiI5cJFnF6K6B8QGQMzB3lWfGAU
0wgX+khxY86VqK7PTz55vRPKqb1vxCqZff+B9dsdW0nhfCGNN/GFBeDwzK1rfvkd/W8kADeb3GXV
c7fj5/MwH59vLHad0SKwIyb2LTNV830qeNAJbuKTfsIpYBqezKgNJat7Bn5lfJRyYm8P6wyKI+Rr
UnNehFQb4GK0lPXZw+PJnb3G7G1j4bsUAoC51Y+86W1re0rcLpwqDF1T7vefulqCHkgaKttZR7zR
llawLuWJEoFG3wG97eVm3hSLHDfu698BQRug/7fxtPDuhu9vYL2qjTG3X9tPOpfYezhHT0M6rUA7
UAoW3xVDPpEp8rzrQBDCMJ4vB8/iNtwYc7spRt/NRHdkRRTclYoZIlXIxNcUEUfS/upMf3dYNgvy
9O3Sd3FZFa/TIUgh0MZfLCg49OYINnGtvv6M5AQx2ewRgVyTDKKO9b7BIbBmjk+kfyekVST+bGQs
Gb3eH9p2HusymqYFPM+dQcekBatxcQBYOq7oYMTtaS3C/NUj/TF8ZSPFkgcZNDyF0WSAAqKlzxT6
IRhn4ba1tMe80hAW/6wEw7P/xn2kgJoHG69HUkqsj6TW285c5GQWG4g4fnkEV6RXpH9+tB0vxBAk
WgMsPkQ2KU2GcgF95Q151baj1jcXOkfmxITyKM2POVDE7qqHRY/s/J1gxTuS7kBwpZF+QMGztJan
DHzXfwf3Km2dIRc27SJu96KHU/IYKF95m91yH6FBT7fygxXUaNzS666uP3UP/i884D41zeocGRbo
CZkr29bWndjV8qUSDcN2/7ZZsMQ78gyvY8p3appjx7kACbTdMSAgHYAfmO3LvsnUn+GRMXrKSs0/
smonMzhaSmT6AMK609PLfpfA0fd4IkTTYnN9M2h4zs8wkMnSHlqkyu+7qwS1tfXNDlU5WGxcTAQc
IcdSdcGcRBa0W3RaoCkj1onKMeN7Ha+XiglQDEDWFv0PAxN4Iba763akjel0km/0ZIX+Cjan8v4+
OA1enuso7n0n1vCW5Fw+r+SwVDZTo2+S0YbK1OWXdNTNIq1aaXUqofvt3vsGrEzaqKc/ONA2gc1H
fcYRtRAJZlNBOydgjvZvfeZdR1lx/q9wHt4OJvtYPK2RpKXSfZFf6gnHzNSHa10qnw3mJvgsrqAB
73rKvqbVlezTMupN+OROTFg2kNdB34bfMHyPImhpIxdjJihoSTPbOg/eXNNoh0PfKG/Zom47dzst
KzBOSA0dLcjOAri51p/1WCP3AlfFC/K770cgmK28D4k/uHN/kO1m2KCdnRxAUYEmSrUDAIPgMhqE
/rsl71g1Cqd5dZLjdk+SkxMgojJ0j8s4VYAyVZWlDbvI5OxpkO4QjNcQo1OT33U6bwpEzgQJM7eY
a65lIykRUeaikHMmq5rXbpowGsthVeAcvLrvzR7D9jhufyQZSl72a6f2BrKxs7laXEQcTyMfGmqW
dAxYWaey7UGnreZoPM8V8HMdQXRPq+7LAp8m7LUwUicGTUhosQ2HcHfw16s/vHHBRLJ9PzOtqW50
caVegmwsfHHRDgkb5ZcGe6eEXMb94ZS3X7dwZ4uHYto0JGFcjnNDsWKl0CVnreA9U/Tb8bbfshmT
KJDxgvc6Lyw0Uch0rm85kky4tpHsWrmVsKJFHIOE75AlougYx8arPdLO7nR0bpe2J70ruQD7Wwht
fATHDtc0+85DhywtOP+d/FnraHOuCnOggQg7rAry6egQMCW1JhQrSNlOvscjwKvOjJaVN9wVuncn
ZULMWT3LPg3s7cii7orU7gUu4ZlDDWRQWdNke8opMvWTUfYeDOSDpg2LxfRU5S+Y1fA8Cl/zsaXG
AMbD0BCD0Jg7bprtk20vwxy4I+jehdBDOudcw8B1zvp6VhiMsYSBRwsAuwrapp6kh4DpyoaIQy+C
jmhZknvuV6/overIwHWre/PNQzt4l3onO0KAsbauZpfwr2y6iyCGSTZYY1k3i9qvHt7+Ce/eRpVD
iv3U1mlITpl77GNpkNdrDr82yEuVk/nbM7hcbwS9qurINSKKkvufU4ltwdiDrsnTqEsjGK5k1Qbn
QQz1BWwAmqZ5ZK6dTsZk3TTG2gAAJ4xMJ8BHzFmAMD0DuoZna3lfLHPAIzV45Hori7utY7S9zpf0
+UcpI47+ZzmzdCCIvS5coR7nwUMZNywqc5qbIAKH2kHglpyD/Yje2Aj/apRHTmWDYKHx6V5Puyew
oM5Y4TBpyfm9N1/jB6XGDxgIRXrO4Sku/om68Ike/vTs+10lyieNLGAazY4mgS9BABUJUYCXSsY8
qqHP7qTmVdz/4wFpf63aUUAeSmdBIrxgCLZ7OHhIjXAYQ1qExwjpIwFW5h8obdCc0B3C8+042W+K
MkTXw9z2GOBpr5t7BCTS/xNof8+piuW4f1J+NlX+Jci40dUAxGBUM1y9v1BPFlo6axVgLJKYgaIc
Hu+dNj9QookWUCom74NxCtHRl7D22hJOh+uYmBNeOJBnPa80D0JXtknljpkFcUGMaA9lXCYv2kl4
V6Z6TcaWu/khMlaeOm5AZBsx0Vtj+EuH1Wl40qCrA76n54aqYbFyvFtZzHUC34/txMOyblp5CuPh
KxXhVXSzwvJYBUHaoGJdojv55pWWVOykvSXVLYxHBLx+Tg9j3sYMXicBZZnwrTqzbDD2EwZwz0aJ
HHfgH+fomrFkXmwnu3J/4Zvu2wpom3LyJoQgR6bjtLV4xBYbHq6fz/vDrX131998ifSbacw2vxPp
Y+BZE2usgxTT0NlEZPMaSKkaQXI+f5JDzjZXCLROSl3KqE5fFuLKW1A9fMnQqt3monf4lhD/dEi0
4apksC2D7hBDmC/5sEOBlmoIyTpTrWe4JBJzRWQFgTh/Rc7gn1EjVznf5FVUMLjSNf3Fj10EumS4
aVCJnz6Kid+/C0awZC78f64VoEziX+F8nZ+MLCfjL2zP8zv2D6cuF+3K5Yw6Oc7xJ17swCBF/qFo
buHa4QsB8LWpLNDGavQnz2K2qMmNR5+I1JKho9x2KPogXrogI1ZEZWIoE/pUPvkREDu6JYQia74f
W01ZiSYPqhQr0tqH6ckWr7pAQGCCRFocSqDB9oYxc1jy8H7w3u4pZOYGAzAQ127v+52RmyOKdVCS
clZ8zrzRhpSwqaVzF4LdffUCtTHJ5I5SoCYuOkEtB2HELWbGoEFyeTxJUQwUp2r+xsZxQml9gA29
JtNUyH7sMuYRCNzV1I8RhyFPNYgplW5gc9eoZYJ9fWM/2C/0saUzUWD3HbbeqBiIeoUK87ZHVDGh
SDLZfpywGAHpeFo6ka/T+mg1u5BNaf+1vvZ1EfSPVkrsDXE+1ye7ewUbY60XvxAcIq6v7eRQ6vZi
9fN9y2OpKVHeslIiZlgEfu3kSX2wD3rbEnpN1F+dAn6/YZqwTUblFHnEUM6gBZqy40d28+ztazWT
OIz/bdHU0yqsqPiGlr4U/YgnYMDbNcI6bxoBK5EpAg4Em11GUb6mxWJdo9WfQylXYBk1yoa891fi
BI3Vn5YcUHXPcKJHj9ddZAcX6D17UyzY6WohFqZrj13W/3++c63NNJMmIi5XYoBZ+nGx4T/SGRbT
FQovL5hUX2ghQfcZTnM4JL6wdOA76oSLYATdt628gJcFRsmyG1ngAZ/3N3EFG4r6DD3l2la5zSQq
t1rCHDrdNKy8LBEOZOjJRbcE9gVI3D+xsFGEKG7V6xqDXhOLNIsksI4ODwKsqtK5VhRYd8vbbRqc
6eGfet0xKbNkfr8RSK+/G9Vgv7UTy6YweHT2tKUQKT9kflB/NkOPJ1U4WFB/Luzfh4cfbqrMShBv
MYunsEWIdE9hsw3uginirHLP4C2g6tlh0lz6yQ4rUyv4D0jOg1CtG+i4p/hP73ifGCxhtsP+Xcan
zweGsfygJdt7GSr0J1G8dOHW7ah/OFsFR/gJVYz3dkdIrZfsybxWXL6QbGpKG061KuiUHtcoICt2
K4/m0DcgBDxv4g8koUhwBnOBuNSbL0kkciR0HyjI6wwL44MWj7rnr0nXBnBtHIfPu+VWsYnsv5Ec
9qAEyCmEQHrxhMUZVbtDWGayo/o02MRoqSElHK99DPXXxyyN7ARljfDW8mW4BEXIvhLE+lr3Xnyk
/gBkLWhc71xWNlC555IER7sQ44d6lUd2ZXEBq5dKJ5VtT6ehdpbAZ94xcYp6GJb1jOWZ9uD8AlAe
TgY6j9EuOfFXOuSyCRvuBvIgelVj4VbAfH6Z2ay+g72Pi5ACHTGcYgG3ms789drqr2xa2CpqBiqS
XXwelFwrlGX1FJFk6FPRkXXUf16xUVxnyk94+8ZHZQ8e1+8LGno7LoSgaOVjD+HjDJBdBhM/xcw4
VEiKCOCiHUEUDYpHNb8ORV+bEc7ZyYgOttZGgt4E1KS2sn9nfq/UaqdfZDENkYUwC2Osj9gvMegb
e4nk4PVLhR5mBB4ukW93n4730UYqrVAlMo0VRCBkam1Vc5acwuxVljvwu413fgrTvIqYw1tvbG4Z
PySGjAivnaFCZIzyvs9UUiTYIp69I1U5f5RMEBmL5Q5Ywo3nUOzEpfQqwbTQI/GEM7xmLqIrabpE
ETLRFgbInEo/yH0dNLdI3HSPcF9YL97eQnGIvj9W8od3c4YX3uXa+ClBgRefNhFtqonlhI0r7r6O
o2VA4c1gxdtAvVJO/x9/d+SK59Zkh/p7Cz3YtNL/Bjk0wxjuGPQx+x0CfqUbzyGjDMoTy7+TaBXj
zhleEr0VFkTImgaxTX+81m8hcpC880wz6EJ7b02OAh3JJ6g2AYD5Br+I0GyILkLEzpTlTK6A8EIt
ApBQcd2SVfy0lgkbxT2difAmhAkpMkcf0/mtf6aiveMNsDBfVsJYdtY0ZcwAJzWvR4j64gfViPqG
LtGCuUr6wkB5HW3Hw2V5VwVv64Xi6Z0b1JnmjL32ufh9jCtFXSs+XPr0+qLrZhkCPCrzAaO7pYg6
9NCLKKocqeLk/2N867kLDWC/eWKg//GABTy5ip2ICRZIGVL1JKKAdcEWH0CfUKOMLwFgpk4r/xCO
dDSUP+bXxcpw+Uaal+9ByYvxJnEAjpi84gJqdR2Xrrju38dWR9R8T0Vmyw2vqOmMC6KEi/anWObz
inGWqJaeQbbEPDto8BRGQRxtsFAKGJKGqe3Lvb2YxLZT2NQFY34yhaEjaTvNiIII2rNzPrP3hKcS
j3RTH8m27zugj1PF0AURhv8qQ7xXwScS6aKnV9hXVXdIPA6yDTFT12jH4Z5TNQwQJypqcEOkWf2p
KRQBj9DrfZN7tLTm80ZmQ5BMiOQrnFS9vbdni41bDtAZbYsYTexNP8uovyoQ3Mwl9fLn7tYoivIO
7X7p6Zpp+GwQAY9rpxwOcLrWLjleHgXktGXQ8UH0ijE1l/UTlK7kSHN2fyPKaCo0oq+rjYfJdfFz
XXBN3jB0731bpQmqUnTzGDnMrqu6QFSBYSLYgyt3C3+EnwJNc5kKZi06yvPUeTYI15+zxe0PCH5a
u35b+1dSHUwwoPsM20eHHSmF3ySnl5gJA7dn79FroAtK5xxUlzoJyyge7aBU3UJOt3Y1Oo4u5nol
ZFFZYLdrtQm9LUhNQNm7rfH7f16CQG5/hGhBNo+VXVEQviAIA+DYYdHiWVBYNBO9l0cbsxWjlq0H
2fumnB8rKGEtycYx/MLw3GHKo1nniRSzMlu41DICZo/U0S7r0uYw6IAMi8/MutnQoXcA2EZyO53Y
Y85Hn3QSW5E244oEnxYlIzuKAAojw8JoOAj0V8y7dVnoGtVA3gX4gktm+tlGDERkMcbU9CoDGARF
8VhvjoBYGy+HDOtOPCiXzP65FfuFjtNwmqz3eLCQQ9KbVcjNu4A+y7wWsBUkcwkj3WOc1Kop59sq
rbrhTuyeHeU7mfy4lr6XfsejnUyAwZL2K5gfw05+tjj3Xfiro3uCn2BLEdQATnYFMFmEQqsPBZ1Z
FzPr9/EQXBYH78lAWcg617UyiOcNfz0Uvh+oXjAaKzuhsTyCLkHYGWGUzk2UbRLrGVxE0nbxcodG
EPxIAy+xwR57Fam9pLPVbZVlY8ZozHEvwX3sNgo5/niJz06a+Cv3MTtdGV+uB2OT3iLtVXrwuYzB
hT7PxLjdFMVwK7I2Hom/71WiqUJFdubYvVU4A/ZBRivoFenMpZUkWUe+ndevjMmMJ/G3c9UZU/Nl
chVdp73MPGzTCbe/RpGsDGVPUKGPEfir97OYPNoc4ZQxsKTCPHrwngUrpGuelswbnxhvJM49Bhdr
FpMBUFSxxjzM80WiBnZ5ZNeIidxqcO/9oVPF9WvVMX/lXGB/d+sgqhwwCG3T329/7hT/9OqFoy07
UFRdrk3RPXfxBsvS0+v9OZ/Ugba/VZ5/9Y6idy8S8odprhJ+ZSEkY1EFCwxqTrFntaMJ3EXwoNm+
UV4LUxpwS77vAG7kcZ7ngnOS4+T+fUbDfw435fnvCfbUfIbofzr0WFZNn3QUZpxVOJbbuFuIyq9u
ztkVDinFlCaurD+JGN0HJHY5RJ4hTKuWEWZNdfmweDZmrEZFGJCynRyettQkN79nMjoEXpUWxoIX
7webFYxR0hf1R1j37C165fX7EUrxBQvChBbXYrEQGYHbY0P/EoET5D5HLdEG9L2pTkm0DVZyXiYb
id44ayTEySdRRd5MRPAwIXlUcjjASOVxDKaWaFD5NK+GiGXeuSIXeP3bPAttUpRdZLWqdEW7i7CU
Pysa///IwLfxj76oWkmbGTILb2rZjrWww2V2h91t3RcDmgOX+xlYmCzwQ9fYbqx4nf+8u9B0e/Y9
lRZg6LfpePnEkoUFysJoGqfLDCU7SSCcBcOg5zeFhsUl5uxvnUeCA2Rf6KmKLQy7Jk1Upivo3aS7
UiPFQgqdDBfneuAgoFbjOzuYF6mnioqhudSDjV/+LmqA1w8y4GApuOQ/DtFUiNb1RF+gBGHtHYhF
3HtsnBgeJJ8q+tClZqvwqdQ2V19pJBs+min2c2b2eSyS5XcaEaR8H1GkdNslDSWv3wq300d333Xj
8LCDEdQilH4Jk2sctrrhyD45m4ObL4dWNzAG0Ka3bZa8aHdqe7Tt6gZJxqVa/ogyCU7CHmosNlhh
3AYzhRenKWLa3CLrg3bVNq8Q7tcQ6DqDoS3KaBJZvLsfrj1BKAnZs0smwVi/d+kLPwewTRvruH2r
K69hRT1c0gS+wsEEpZLr/Jzu70ceByCYf7U+m9yd2NeJqC3q1TALenEMRMrQBuiD5CMWo1ruh0yp
W7mm/0Kidur5b/bhjNaBn3EPk1RNEI8jbnW2v7UNKuNCfnQITDnp0/GFoohKXHM67qXnnef3uk2R
52GH6TY3bJQ+/qMP/G9o2sMTy4B5gL6ys9gokvpm/DRwuQIDfgRdkaZ6O1BF0aiDgey8z3YO1BnS
2Fe3vZtQp8y7vTC5mDjjmX60ezdd+v4ldqD1nzUJKmUjdm4HCPW3i+9eI2LTRVuOs2Ae/w1xu/lm
XM/kfodqQ9K+zHiYifpieieLFquxR7ZeY1jPM9hg2icYUtN/ypvg0gCa1NiyV6Ow0yxaBVAfZPDw
ZrYNCHPwgMV2IETaXtqXwRh7oV2caND/ruKYmR5ZIOTj7etzKIcuJpV79hK7ky1PBDItrNMPDeJR
MaYad6yQcIxXaeQar6uQEiOCW7aBjkLEiDMeQ7jVWXyfa8CRoAZUyxkGX191GYlu5ekdbpnTk39R
qVdNrXqFfzO64gS9NX813jEyYP0OCN36CcKDCSowhhh6eahcK38jrYprh6U42iv5bwvJ5TXxyVtH
nGRQ6I69kkFYT+LvE4wNu0+rXJ6pcf0g/S4V3TkTmLZsN0YKevhF75MWNXigXfIfyQ+sQ5vkv17x
Wg/Hd+KNUIlhp2g43Z/by0tqdIW9dUCCV/eJY6FynYaA/1/ENk0R5nwU6KgoV/u7tptcQnEG0cfS
fEhBp/KlZAc3bfsCNpA9fOEK0zF4qWvIAIxmey9/criOs13toleg/bKJfvhc+N9PnFsgqGsoC8dD
H7yKpRC3gM/OHndK3kAm6wmRgxzfT04jajEYkKXotLqUQWkWUlKrawZ8uQeX67iTsaeC2gwwwXbe
dYRh7ieoMn1E2E6r3DZU08rbGwc84UZZ48oU/FT3QrK43NQG5061kxOk97jRF1HAOQkoPUF0sKy2
sFp95MTizuSicnhQtT4jOaARdoc/rfm74sXsqiofssuZv2d4d5sB7XyaFc8iwsgtAfqxYTl2bHwn
N9Hub3Eue9STQZWaqO8h/qJitpwIe6+8q28W31IYKjnN3/yYv7wCopACnz3hRpQadq3v7ESTSl3m
EtyLFzYgLb70Qsz3r4VVZGDqTCQQcEbttFiDbJ0De4nIg4BMizvriLgX3b9Npq1zLZE0NTjSHHKv
RK1epjyRumoV4HSZWweqLR6jBWTipSVABmR4WI6CIxalLBhebkmQhoL++bUR2G4FQrl08CydqpXs
FIIIKC/KzXkYaaLmChCGlHhhHWEDEKH/8JqggVgYFk53aqvea/a33trx+Sm1PCuINJOUj+jHEVBd
D0w/lWsh6I5DFsw4X6wHuEDsiXHqNCyXKU81zbIjXipmkVznYSzDg3DZUtnftcxxwLkMhN9kVPTV
lAiAB88yzrMtuB6pVge2qtm7WWOa1QcWbLEvyGOLU0tXms/rYVJgKRxbHmqg81gY5Cigaiy2cNjh
7N74wbAUL+fvQtNBx7z5RaC5x0SHT4U6x0mG1946GxSgAriGjGnW58YifLCT6a6AC9dCgAZoEt4c
9dTewiARtePCDRPE3aZB8hQ5A3XTVw87mqomRKhvF1KH35DgxfKOKNo7YQ9m2NNBvrZrm0O21c90
Aje8IqBi9ZiGd4K+8DJ/h3jfaUR5jfdCF8fc8mYqmcIjTANeyITZjBT/cbdRMTt29JGJsj01M9S9
OqP74ZX8P4/UpXI1B18bPiV9cFguQ3bVQ/zFNhH4DntjjDUWeIwNXvaiNXN/lhqiRTzhur6fdbIB
ecV1sjXuQufYC8Ce7AMmTVzPlNUKcdt4ydidbbWtau2Hw11V1HUG2FzAbQ1z7LaY1wCZEDv1Fy0H
230qLijObuB+aDnUOEq/41uup7791H/ytinUJDTf3nQtGYMJnAVgItXoQEXxmy3ZXGHZ80iEfPw8
Fzdy8EVS3kmJbcXTWywEm2aPrVYBdOvQrWTTuXlok0ysI89mCGUUinrIHm0ZR4JSjjpM8LxhpMBo
67mYu5bunkVEqozb0prSLx1Pq0hD8xJL4WOUJR/aS3eeyrEdIsg/p7Nfp99LyQhP4SFCNWeyMkEh
Pj0YAm2wzprXSoUotMqZxX8+MfXM8Gmta2P1IML8va203qyslLuI2t85roM6GKrcon5m/ACmbgok
mqsiPj0v2QrB3xBrWpJ3p7cbvtEy/ftpA2rySCBwahAldURW9U9HToQCBw8PAKAU5Ua4yWAmvmUG
0hZtzeqJy5UCbqzfaOfkhPAL+UZon0pR/Vzybop879tORy2+TltN41dQZYfgEro+9NvPC1ERjDzf
kkrBmQsvN4jWfAo0fvA+ApYBfO3jjc49fFLWkNKuUANSK7RFFSJPWLh1WA0PdW7eZslAtrMePST3
FteMekMWagNSC3+7rRDfhO2qDxgDtDiQ9xl6g2g4uK7yBW9WqTjGaBcQA3HMqMlrSfjCM+MLDDCd
ebHmj/rJyr5KwILwod5UFT8GPoHbrcSURBPP8y2tv0iAKX4jy/1o8Xhhdatb8FBIr8dgWkSxodjf
UdxPsxKkv5MF/k6huu+xJBFIMwx0kbw8918u9TUETlPZvDdoIpA7FfJyWzz4KFoVeCZ76CRDK8Rh
cl9/xmz0hU7qLfC6Vb2TX3aGomdn07VKQnKmVppIJRmvV8x02/GZNht80Bc5G16oXkwOK457iCvW
QcHKpyo+IZupvSiovY1o8m4kNeoz8UIo1BYF0hnUxex4LaakLhllDqvN2z+CEW2TdL5LcwN/hkGI
bN/pSzSi/xNh4SYRl8B36eNfHL/ljjbzridW3wCeACwGWhWW4Q+HdQyI0KyFTFW/hpT3B+mxaXWf
U2qaO4JLHPztlrq0MkcKyMxgRxiE+j0SMMX3bHGJNcvg5ZF3kodfw/b0WIiTbuYXi6GOFOo9yIEx
uaokNV3JvT+Tr4sMg1rmLswmNUZkNKHt38b5arR54JOiA8mCh8vX5Fgcd8pDHI6l6FIg17uPxG7h
LXPrRtbVa6G6+CdHmWRHJOpW/D+oBxkLxq6uQ7BZA3MZ0WYjWXocoYytMNtOkv6DMfxtwCV9EWO0
qIZNx2W1SNeqFmzLHtQ4o1q3oSxv81Vebou/PT0xeAvEPMVUE3jpe2ELt8uukjba0TGS9UqZZqgR
W/68xpuUl9qlvwL0y0IUOWF/fPGFgr7nOYu3W90AzBVsEB5nV4AJSuPa6b3uIiSQuXPq8qfclK02
aXJ9fJizNxVzNT5ZLFZI2g8DefU3OcQFv6v7ZsDiVgAqzT/b+l3yxOXWBCGbajfKUr5yxlpDNgDv
z01747ufbnIf9/W0j+LU5eKrM8t33I1anArJHAo4e4uij5qAc2Is1ju2AwfXfxyAMVXOGC0hH/Us
GOV9q6zg35WKWHGRNA/kw34d2wbyadLFR8bfpo6PGkyH/IECBw13MLvS33MUzI/lLJYLdcE+frbV
8ty0W7xrw2qw7vHa7TPvAwPI2m1HNe4k3B2BwPnm9mpuorwfZd/IRwIubbQcBwYy7r5x0+pbbKcC
lpFxW7U9yc/3Ef0jq0VRqnzu92tGoQMV/i1ZULyCb0ozbA/zPTRV+uws6q8ZXg/1C/+NZ/h16JJf
XXDXpRMJheu15WPzCwFr+zgV/v0DSyaLi7O4NtdIAM6z033ynb4uQdKmfbMQR/hAKUQaDfFMaPwb
uW0XFTBsh/1zpdBu9pALKxmTnP0FbYvA+JWHris3wfcg3gnmOBhT68PlsD5QOpXtKOqc4hjoAzqx
raVgsra3YUrWsLUIv2lZiFJCu3at7E1JUJX1I6e0FGbNVkjggHdIw9UdL6PlJ1zl3uLCZ4ZKkujN
sl0J1NKGMfduyyFa5fC6L/2fFEIaiMoIIJV6VO79/qnv1rRYaJy18I21f8t26eYWzKFUvPAJ3X0i
nIKN3UsR11HyilDWkAbMdHfJEzQ9QuDYss4L5jsalqCFMR+k6TQrfSxZf009SGwm/df/+Y21pGr5
5wk4gFHOVjDYukSYfF85EWEEKYKlJEVtIpmxaX0VAwlyBSnkTLkgaXw4MgSunaK0+fAbi2t/ttAD
a3ZYwj+7y30ySELxpEStC31EKp8ysX4V0EIK0YU1MRgBsMHViSgeaoOaUnYJOk2uqkR9cGZ7pyim
NgJpqBjsDEOfrshxYE17V5dRK8C5Ieae/AKH+n6QDrw3aHE3ILiXRBJEYljZjghfDpsGb0OWR77C
9CmWldbyfveeb4R1xKoufkELHV6ThW31giD6TGju2Gsy/hkLKz4JTdaEEeSycoW99+yiP/7sI3CH
ev5AKJyOLUT6EF3jzWIGilK7X60OrWzu2xUOWtkpmkN2u2vvEzQk1k912kFUr/Llmf4WP/AN1fwR
zElRRus/X/bYxSaZBMVBMrEv3BOwP10Xm7UjAlnP5GYvMa0hn/hkMjQdUoUve0d17Q7mwUoemH9L
pu2XpfP0t94BrS7y6k0ti1f6lIOJYfpypFX6wZvkgNN+C4wetOyWI03RdsoTFdQ8kRlhdSAPpCV1
9de6PxoQjq+aIXdrZ3Sanfn0FKm/VRgL8Z4pqkcYf1T2CPvmKjmncn3efgVoW1U72AAarROmsTMh
iDRR4+rVsdm9+A3QWb1ncF4P4WU5u3yIXOjq8I55BLxxbS18iaS49dPVlfAX2S4XS670CGQTk7pQ
2w9jIpak0ezN6SgE3ewxo4/WgEIAvxR/PlqnqIyQPvWyfH+TOUAM/hG8O0Fzm/WKjaNd8ahF4ZC7
LgM5fc7kAra+ayU4eeY03q8N8e5tJW+CcraL/za3E8mupDW/ypW2QGioMJdSGNABUzkA4ST9uqPQ
y8CBDsiRZD5DmMe6KpZbuP9vmtFnAXiJDVQ6TX2Y1Xe4VliFEqewUXlXjjYYufXO3DiZxUA8rkFH
u/fTTfu0vYxWnFx+m+0CQKob/6hURJXpiW5elEEh3QqGwEVJRvqIBDZTxpKQdehxcVhoRHHtkSAA
xe4tZf/v0c3t4cZTrDaLnZRjTjFIV3h1KpQ5a7dlRr0Q71l8x2bU0+gpBbq7f/Zovaf2QRtoJjPx
yHgJyJkVe8Oi0BnFWB5d7IwiQizveDet5zrUCV0tdDRWYHW4/IChBlmUqGzv8BB0pi40ESSjz8EJ
0E/QlOGt0AgKgTBL2WPQdSA/jjw5UwiNWp8JQNotOCi+s5+otArZoavqG0zEF99yXod9t4jsZo6k
2jxyuZouUUn2rMgRn1IXiBI+MgyaN/aMDWQYx3E1ihRueq3lYCycMLhuNIrRtlKkG0H/wLWLqRTj
NrDx6T6oKXQ+OxrMKe33R0p75hW+X6H6Bxasyxlfd95JFdZhWmvdXFqAF91d1Pf/Jl1HD1e7KLN6
mcLXh/SST3lbEpPUqatUVOvVgy+mSDjgrOFAkaaV5mYD87FTh1jlSwIgmi0kPFcHbhNNBTQz+C94
CmisLl+JD9GY4bc3IzJjJwQskpRQMW7H4Xfq/ZQsTRh747cCsOxF3O8yaV1Kpto7AjcnfzQdr19c
+3oQ2B4nXmU0vn/o6ZoXSWdNc5UtJtwodExLxHr9o4I7nnjB376/nelS/2c62lfVG4YWA89rGab7
dg4L8CMr9KS2eHOgU2znr5IVTRBfotkOFKvGleCI6pQmXfLE/I4Dhg8+0KgU9G2HT3Y46Yge+FLG
u0BfBzXGItWbTi6r5o3TSnFAZaRQ81LUAaai8NUfXsmpQ7r6Tv4CPi7gkQNj0Cc6eRsGyyIgbWP3
1G9xMOXcX2XUSrf1H3zbfBOq819dQH0a7Csfh27Bdeohew7pkKM6bWoKNe3hxJJfqktakv/mXs8k
SOr9U9g+yAhsLsmVO6EM8969qKPHSQNqfgpkkQd7xBh72cQDd3ThYbQ3fV/mlxOL2wn+8kR4M6vd
YogBO/PhuiJuq2DlQXa2nU5+ILGwXs1L1PADXiGrP3QiuExprGbQzecAW0QQv9czZ3iVlN7rvH/x
zmXraIuf6BjiM0bIGxi/E2sfcgHIfmz5+VMnXq5ohnEGIYl0TydZGGF36E2QcYO7DKqzwqYKREss
xhnzDYVCV/mGyLPzsl6kfORJYNOL4EhQEQeQeyTxHfWrAdXJOhkmhvbyRILik6dGWvOP8VOQC5DJ
Q7wiA3LKkgQ+whuLthBmCYDpGixcO+ZwtVwryHlP+N13XWp8EOotUiAKCAZaZK39vxK2f3eS6sTU
dKCETW2VKyMg7IOQhLSkPm269WpAwTkYy0M55FPpfUFdhjUh/ocuNd/82ajoonIb8I5benRF44kX
isXiW5UZWwzY+MoZTk+JE+i5FLh+QqFfhUgLQMc4VuOwjX3K3ALt/9139RYdXMsJr2gD8Edm1koC
6n+9f7nIhkLS93/OtfgqkihLz3cmYtPFm0x/TO1mwMwF6vkOKY4wEX7lR2VbuNZzXBZs1fvupX7O
anGvISFx6tR+xr86quB43AJwmYKH1h7vqHQlesZ2EHtcQFGppVyE34gujvgwXxqZqlSQP0VVHMA6
FIIlZUzLNLO2LTMe6PvJ4w5Q7FWjfOmK9QwLu/J0XxpptT5fw8ETBnTabXCIrY+L4sPbYtleWM47
qeCy2zrG4naYvyY+sHTiJ7MyK1ifLMwh1rzSWeuotxySafT8DFo00zvuwi9jFwhUiF2XK82vUAfn
wQRkv2vC11YUFKlyuylVvDQXZSFXBHWL0t5bGJH5cLvIl4hxRw3NKioeI4V2hXoFXQnXWQoJtizi
GyCEozw82uNHcvjWf92gLonJDrm00VA5K+Kjnyvi6fj7WolWnukl7bRF9dLQuz+qUxPEsl69F0vE
z2785o5tHtrQF3mF+TPObfrtIPU5CF4z9GNd7aHJa0bA5lCZdwc+5rAAfjwDjN0IaOqThVRL/s8B
8TtJEN33q5GU6LfHKhSAPx0jLVgUQ2++ilPJbi80ntTFAsgahJkJCyeFILqYwpcj0R6rVtpz6l9b
G6V733Z3/nKHkLtoSnrJcz7AFs+xoyOt85CJrin0g5IYQ1I4pOmVHBzYNGbHf2gIZ+TzLeCGDUdI
AlW2srd2YLbyx9/2PofZR6Nbq2yFGIP92qcvSacBqcusRpOyAn7JeQwDG0Qlocf7gh5RpbdXKqcv
55L58sn1Md1RMK+7sip/LnFdqz+FM3GXDxJeK7M3NuXGQIbcNunEyom+KYUcnZkLKP66/mP9OBpW
T1yXEVaAX8ntN7naEXYM0Z4p4C2FYXXkLAu1/0lwJtVkVXNdIL+V9h0jMSMEkX80qa+miypyX6RJ
yku+twonJp1liMh7/5kcsNGEYYaFy2Dt8r+nV2UhdjQ5lu/v00c8/7QcO0RCAHWaUebco/3DT743
jvWPIVoVKVU1eZNGMXSw31mXOfB55Lf/6Od8t46LtKSLD/P2q7rStBSjGUdpHV+LoEuCIw7JRvDQ
hyJRETuYh83V+d4DoYuAbNmae2ceTRdB2JMS/eXOemcEwOFHnfRAV4b5AZmfz0BPj6fas+5LL0QD
+JpSX0VRa6T+c67fbjXJVJaHboq+LW4IKFtUm0cS1kNzNtgdNa836c2o63193ydv0VUJ21Nn5jvV
uj6+mKDfcIMEZRXnsMoFbGowFqWR4/5uiwf4ZRO3KewBnqCp3fLfj79/x91Ixx3l/7pebEk/RIDQ
I+8Go/QW8x/ET4+kGrgqhGAR4jPwd5mzL76gE9VHHoo0mcf8NwlGwxwmRyr8NPE/HoJp6n9SoM39
nClBZ64qlDZ6ISs48kHjqfRl8G7uN5xTjm7lIygBoauZv/ycw+xjC/qASZ9GDpFDAmXejYG/niGa
w7qzvH82zdwYT2J62W2zjmwTXLmCFXEodvWBJkMCu+1nk0CFIYOeI4RfxWuic3ULJ3AmPGOPU7+3
hD6I4OMRmYLaealLqyOwGvByTYp9dMedrhk+c/pIM7z4LC8+x4BcWjhaMJxuWRbj98JoAp2vGA3z
paRrEhdiVVpkC+PPgvbc6ZPzNzJFC1HTeDZAjSk9vClJmDx4bIxXb6XezTRPNWlVMaG8bKhj2oAw
QMVDgL27WemAGLePnZZfxS2DaEUE8syIyRLIVMGXB1iuVSWgKdokvaXmfMvx8S9uf+vJCgAdOh3l
MBH9I9v4+5FkgqXrpF4DkmHEQL/nCvryFetel8UXVyhawtDxb8FP2oVHjXt3B+xxDW3qs71+insl
dnH4j+D1Lvv9CPPfdyymvgn8RAPXxk5U/qoMPLG2QgZqKE1dRcwAstOZGam8YfvFFvB2IAzdh6rI
bC1qaA6TJuRxJlChCq5HQBI44aLB9+wOS2HTrrpz0yzY73jx2aNSQYuUvGR9jaf4eNWFFdbNs+Io
tk3unYnIeRJFV8MCP8uNm1tCVQ9OXMCtSGn8QmK5gTVlio+oP675looPoTSAeC1n5qWX0+dd8EHr
h+QRl6rvT9Pjhp8v1tupUyVvyfAUV39oFNr/Z+4aCu9kKb5++2Aud0Nhr6+8COh5ZEc9nw/5L9Wi
IgPFkdq0r2fe5eyhSPRVBATdALg2EJZQ/nxwLA1xw/MdtsFOgF+cnoaq7bU+1Hn/WHwGHfx/iNWo
OGc3fBjviq6/NlbFzixvLc6+4NN/lDsgiqt0cJdEOs0ugJW+XzDuBDKYvOZeE4SuhMxYGh484KFq
GBNVpGq/SZy3x2DSKGo6DxUxsEbwdRDfz+1yeQe2NT+wwdUIc2z/h3CWz+q6zKTCodTqapVTIw7R
UyV3aBKO42WeaO3ZcYlh97CbuX7y/CfRvYkDbD2B+hILxK6LGctZN/GcfLFGSYe30bzjyYGJ+glh
KZ/7dxAnDl8OwKdMKPObBLBh8EUOg3sYd7ZIn3VMytF5Hikvz5tfw2/1JioWLmUBsXdYBrdeDSKU
P5CL8meJSGSAVtdIKexykPSmSIMMgWX5zEUSQ+eC6PmD56PRtVAwbzqTTUoBkYlR7T+qw4Yk0fjY
PpteYql0C4gau2X6BFXaLZC2gG0Fpg3ZNbxnD3HMkXWIx9kYaXyJ8NCpeh1kK0aOeE1ptHdPElxF
O08lkdheR935yOG64Ktig9KFT8YObTj8Jfm1w8VKLydK/SopXGD+K0mK1g+pxBS+/PKCiiauv++w
q15ot+kC49GWZ8tLaj30U87j69gd+tes4uP+hn/wGGdRZ8JSgtyR+q2K2j0TmmgaU1x6Dnh4CI2B
0Pxa765WU5iUzmi5LHBidoprjdJF5pVv4H74q8ok9gJYoSDPLpW2hwaXb+aO1nTBvtlStLjDh81A
zEjLkGbDCuJ3EvYoGZ54yFp3d/mRTE5q6UsS9+d8rlEuoOnqA2IMiDNUrhh4MCvQoimJ1ihTURwq
AK4TEjNgM/CAoyKx5kc+/H16S/gndx/TCbt/BEJmEembR9THeUaCAbW0QuVg9qOJUHpWPtLdrI6Q
rLKQIDKdhaGM9U6MSCm+lM+mWdyOONbktxfoJQds8uy+PGuvdUmP+rzJqqdHC2rVZhSGHqHhoUvy
SHvx507B6B1RDYXNFd6WqIzYGZe1xECgForoQze2yxfwri616Qe6Rs6U0uDIHkCucX5jQ1i3SoBD
NyftitSda8L7Po6a9rUgDNSfOpBx0TjbXCiBLuHqwSvix6G4/kkdIp+AkqjqBSsk7EENnsdIH2pY
b0Fh5z0FgdhiBWGyzKZ5N/RhCoC+L562y29eQvEbZcKF6FqtrHXEke/THMPyxL7PRKtvFArcP8eL
uK8LJcQhElCaGcZK+Q84evAEyj4NdWvyoViCf5AumFEedx5DmklEbHpFMvNf4NBqaQIdCjACEyWj
MQzIy6ysiL7XBMjRLsCNg8dOL0SbS5QnuTlJkluMfH/jsSiCVDISGkfIb98N+C8w1xKiOMneCPgi
1Wpb2FJlggK+Evwkx0qur70sNIDlBpxccZVEQKm/Wq85GkDG8PCYnCPM9oHIvoZ/8olvHHDs3gLW
rrU2Vynv0d3BTHAK8nezD0uyzy862TowsQLyXAVGC2KZewYFnd3cFrPvxbtMofGU2fwKdsa7EAUm
dmKydzxGD/qYD9+m1L/fBDrYoPr7QqnMnUWu3yQ4N3u9Pb0EpjoIa5R1NpGFZWLF4ndoEXPLOHt5
yOhUIDfiiWR8756GO0Rd39e1UhJCUiuRGnKkDF6OFijBrXoHa9cpcbmFJlNM4rZy7wIjWMCkGHL3
aAuaio96hj61g0bdLLgxGIuW87GHOcGZJmb/kcUZW6jd+3SUF6sXKZXQs1eZgK1OWeux0IptDmRs
aVoDpblmhwI4KZ4gaLGf5GHRYXiB0oQkE+1Ksjc796oBX75bHsjmpF1OWvf6bZiWdNiRRDastSyf
U/2AyROOJgajxU8GVZU1YkvdnSROdZLXvI7JokxfRFuTGvIJL+Ci9Su/oabeKz1G4+PA9BKvdY/D
E0Qer/v1iB0tRzybayS76qyloX0Ou6E+PyJQfmkes29J4wmmkPYZj9EsGTfCHlMv9JWCibAmAvmQ
akUgkCbcJZg5t89Q1Hl8k8ZVAVW6HHY9MyWIrgx7Wc1vTycErOQThymbwvEuKMMLyBnDvay3PTJU
9qsgsJJUHOfAR9xE7x3PUXZwM2SqaEJz8XsMi3ddiG/ddLHLDuSHy6b0QiygjnfUkvx/gHCaUiQq
8nPPE6bD5JTXEHE8Q6F96vGRA9GoqfnG+3bjcWw3xDqTzIwhtiZGmcmIHNSyLdCi/ehP2mKpCHv9
V9Xblyz/znbZa7saFES9VSghBedT3FGMaQG5pQU7vZJn090PT7V+awEQJ2+jkHs8ArIwxxPVM/wH
DyrTIiqy+5LAIsdrhf/RAQXkFTQhj3VZ2qFCAuRmKq/SHBO8SRF6ux/Z8xcDAXx4wW+Dv6ZEQRKv
lOGdNQkW9T1KZUf8QOMM5u+f+4Eh0SeapZj4+bfSFjslHhhdFiDmlTZtCiHdvs1lff4QtWa425YK
YgMww26lOr08WWgBxslrga/+ly4CWKNWSLXE1tJyzw8IQmmnfYFqzODMPkki+HrTWco5zqkGkv2M
6VmYqUeuvb1Alf8XSqIYdGQRc89oobM/7fOG1+/Cx4/95qRoq7gLERJfbhQ12yda1HoJxRYpiBsA
Big23wkn+DAc1vOAMgCvhx19CCXD1JAZdb2p3Yk57ozT1vbzc7NK8/XbLdCJ/IPHmiOd2pvu9lDO
mjLGVPnOX+N5Ex6RCO5IlR7R2Z+dC7oQTA3iCgRd4Zg24uE1FxXj90avI4Wka4jXMO812O6/VZJ5
z5/1gKILohgfuc9Deq6CYzb3MLIPld5Nkq16nMYy/PENleEkL5RH+TX6CzxlnmVnnKC797GAzy6U
eKZrB6rxUgrO2Nrb+ODa1KufvAFQ+uOKfDXDE6+NUCEnFn6uS0534B5cz/jG//hFtLp/FQsR4eXg
wXU1I2IvEU3r8Zh13tCGWJc4lkG2zj59XIvYeqqf5O/vyVJ6l01pz01DT47nFZEOMDJAZc7z6IFi
iuGbRMNNluSgEsnlt955ohBfI3Il1pbjkPGNL9bl4Wu0hSsP3Kxu6+12j1J4EqcCV7LUqT+CtAn+
EstOmBKe2V4HE2p7t9wPqiFdy+VPpIPabeA0/Aml+T1Rr1toVKBGCA3Pt+BTaaefzFK16Vny4TUD
3rksns+sn/ufVYEe7G4/IOpHQ9TIo03YpQ9QhJV9X/KGfAvnGJj1BOATswC6yYuDSCz+9yAz9pYS
PSS0Yn3ZrIUu9SzGKRS9j1mcB5L53TTT/Bk6MEk+dGlgY3+SrDrx/Ru0MxgSvOn5Qi0BsbcNDEzV
nlQ5KsPwDrxK9ybSJYYlWJRB6YKOHzffRyyZ5O/KUApJnEyUCkaxuLip3bzeyQ9wYqvPmzNt0b2P
Xnx5nNyWjtDSPWwgb4oc9SYCcQ2jASt2iNch0PDt8Z+NHbhLKDt/LTUVv3b9epa85zZ1RL+saSCs
Mq0ac0EC4ws/JghYABALnSKSe3LQXwfeopB9xdG4UcDy3GMA5NfiKJLueq3BA7NuAa/5oHN3+Dc1
UCTP5hr9VsrYbPS9nr2g6Mt0RSk+6YFXdm/eQPDSIxZ91zIXXbNpXlWcYFtjm8Dxd6CvA/pIdWT3
ttiXQNxWRSAhbDXilFx/WoLgsVxaYz8NjMNsYUZ/HDE83fnwGNtzHHqNUHSuoL9N4XXhvXEDN3Cu
cphbnoFbpzNhpmMon1JruXj2ke4lNxggDKUTgh0XTWvxQZlqATyECKZR1q/tsr2DtzLDozknaY5J
JgAeS1Alke37G2VPtzt/hddR+xOTnoiiLtoUZHCfExnm3WAo0iHu2LvFckTM2UV/9rBDqTJhNqzG
BjgxvhXMESunQkPXQGjc9AILHMcXIgwQnvUZcD49XZnuC+9nDn6oJNKaXB0+ywfmEpn4FnnUrTnL
G9QQBPLYBH61orTp0OjgLXOsiV+Jpp0KeNT663JfdYfxYETM5tI6L3G7XAa29uJKCt9PZIwN1tFI
LXgHdoa4RNtZqbyx6YNgNnEz4UdUnvDbIqnRG1xjPJDlL4+EyXr2FDgkqPnXJ+21KpXd8HpnhAl/
UshSbnVY+dmuSlmrpnk6DQibbxrvVILRc0LUN2PS6ZxGjT/GNkm20RAmcVMoapDLM2jxSR+y4gdS
XCYEKFpvx2OYiXe5bPs75Y319Haojxlp2GyVy9t3Zk7cHkB/xODqqvbT5I09dSjts3L4/8p7mBVi
fvwZOaCEBPcGXZJh5iGdQwA6XZjwZYq4HW38DVXPgv19eO8EGeLBkaNgeqnet5bdWslzL/xWn2i7
mLhY4xCwVGS3bTXXkDu/SfDniyw6XMV2kolJX3xXy45VVUwmVYgWNbRk1kiS2ccrnsIZI8kgmh/A
5DFiameWYC5rxqx0pAndeRJ24JxYiOhDDv9V1C73JmLM5LjjV22HZ+E2MZPjsYdy4h6AJ3pGZTF6
qkn4zDbNSDSYfuQ5USQw/Sry+PBm10/Uw0igeE1PzrwjXdhzOwkWkgzAmXGghd8y7fLCXrVMbJjd
r8rOCj8r47nwxpOam24aG1lGHtNinETqW8hRWa15vgZEWhZZnRtfl0w5N9gSrYoJCzdHdlKehvmG
nJozLhWF8M96bHN0hnYWXI7VDp3yCz5u/rViivgo97hKvw4Hf6PoqVe7KAhyuICT01bH0zIxk8/U
xJld/yLbvG7fE0A0tlsKSjAEfwrkYRAUsjSJuzqCSdsc4vDmQBOFoRKHzKheBBwQ+0wpkA824FT/
6GzZIN0U12fdl56gguSNWOL7Tb6kDywpr+t/oHRslTG3y3Km4FM0NTNqyvA29pIlJGV0Ja9ORoCk
Cg2xYt+WJLVhGMOTyVJlzWD/UqdOQuV98ReDTvdptOiV0mSiijXqXjGa9x3ToFE4jZAC0PkBYT0E
iGeOM8cMP6qaBvklYd2qHwWe6f623nzN+U2m+U/p+H+x39YLsqmOT+S2iZaGtN+jz/QfhDezknZK
4pssA10UuwkDGWVlbiPTZsyLJtMrmo4gEAaGxL3E7SIBIRgZ+IbbXlCnanzrzs12CVEpV+eHbooc
CUMr0JDw7f6mdQDlSeFrlSy1XwoJDXcqE2OhlhPDMm0wHQ7rrOiwt/Bp12tpX2qbSlb7UPvzitMe
FNjCSpDA+xTzN++rRu8uniMCPyZt6jGKV7kQ9s3FdIGgwyEGIzIYvEa8dLm3DBj0lDvt7mekwZX9
u/+mTHp8Ikb1heQGqZ1d9rNAGvNjEQzAs4Kss2cl3dLWT1+ry6ei2q5GC1xPAc7JTkrgiWxW49+E
RqERwV4YnQrvw+WxNTTVWUW3FWVsXGcIHAVpFYKyu/AMuuXRNnmhm49O+bB780PXLOGmv+b+bmfP
0NIv0POmNOeWqEeLfG1BH28NZnOD/PIChOejP2vp+lJhRfXFBch6cGHSTLNMm39Jwuxsfb2NLLsN
VKQyH3VgvhaExtbjW7cP7FnHsnOiQy9FMkZcbzIBqjar+yuu33KPFmdS4mWbrEydg7vybKDcTW0J
udkYbyMqf/LUVcItv2p6sLH1c7Ur0bRKK7Cj97d6aqoZ1NqE6rwfGhtyEdaKziAbUu3is4/UqLvW
ODWwao5tXcJBj6r9CdmXfQiTicIz7UB2zJ9YjHsnrnrOY6/euLoDyIRNoBE+UmH+HpoNO3bvmElN
8g0E+ZYLZ9v3X+2dzIi07NkSnEYZTsxDuuxWlCqodVepIs7JT3eufSWWrfsa0qqcJiag4/FgePLD
wY3CpV4ZUYtrpUMrWhSxMPER5Ir2hXVi5HTNv+Dqvyv+ZXcWzGW2/nqMsHrOXyVfquusRqBP82Lh
fa43rRkXyFMdHC27Z6VaJRUWVXxDLvrfN8GW/j5LQF7uZNRW/JBVxfBAYZTn2LrnR5zO1kqXDmX5
Q9QK5JZOjsIziKk+iuCxxXFdNer+KIrYyZ3XnnTMB0jJv9s2Bf9b33MkuWID0i3QQgDAFSt7moXv
3h2pDDFUUd0ZkJRaxyUJWqxpZNZCGXrU7gbKSMuI+f7yUWAP3f6yaI2ymQRpS+Yr2RPXCQvnjQyB
oDIOK5PK2Pqd89OR4PtMPtd0mcmispHdMBzN57U9bquPvtEveujn+qGM7PT5bz+8PvRSaOkVCZgW
9g6dwC6DAt/FIjckrD2XOf4fXwX+cC7n6h6WtoqvvKLH/ysuc7xgwy0WlakINrn+uulm92c2Dlhg
El5Wf/UKbnmNA5M07bCM7LS0kaV9rpdQtzxCnqcYRfnqiCwgrSyO1g5Fs3GNuulAUWG5m0HOEvyk
kbsjFZIS/mVtwjYU6YYCc98hElkEYnHzeDklrLVe3POAbw8eIvp/O/ZEFftC/nEBDE/7i450Vder
oEa1SV2CoMugm2X085LMc0rr+7gn1jWXxoQvkfXkUlQNWHX7mqGbfVLCjF0co/n/VvQLu3i+dyZX
KgEn24CxPg7lHF1Kti1ULeq7IhSCj94nrypesU/+CYPBMw8GGeiZVFL7yelY4x/zBReyqxi+dTRr
/rKMus40dtCL1CNXAeJj2pDBOfyDeYomTVWrzO8AQoQOaVOVinWljZZP84v5WoL565EYN0ARFOu0
uBFqFd1rVSC7bbZQ6jmqomers9Gnvx1A77g34KNglf92jomeQoh/MZ/yNeIC8lokPRcysDl7SvI9
Sw5sYNCld/2Qe6BpiCn8fmhnTavjAqLo7pl9D9e/MtAVp/olrWeA3Rh3MNe2OHn1utu8egU3Ah4b
NUH36o1LVsIfsV1xMElPuGwtwZoQGmz7a3Oy8vTq34ydFnizWKiK0rrxvBUjVOoa/8WWed9RKBUJ
KMFqfuZMjaHHPPED4BeMrO3VbZdC67C9dtINAa/Sc1C4Pgo8PkAZA+sZFvrz/LuAaDPQhIQaiDNY
jnMr/fMZIA/6wFe1fdfLyP4/QERd+5WXBylxAMYJLZHzOevQwPLJqosjW5EWiBXvdbL5hCC3imbH
Zrb+RwlGXn870DacGtQZxSjmYBX30hPjRI+JFZqPSX9imNXNtL6O+jbQ+6trlhPGe7k+VKgkL2oL
uZ6tSSoaDsOw2FikBbLhFExTRlostc9vOCdd7CAisdxUyrPFUXWxYtIcA8+osirL7YgU9oKHTyeO
N7w4RI6l/bLF1mYXmIVk9BRePoxnyvijW+rGWDqQ/MQWZJUpU7bAPPL4Dk2NkJq/uMPuaEuIF7ji
pfcWBWXEkPWmOOI70mwm8b4rX3PwF0vXoLFtSXjnxJtPQakDApB9YaZCiqLJtDenouJiXAUstmgA
PAFD0XICJE9gl8xV2kk6FG6lYWX28GFQ5+bB70WA+W9adn07XLsosPz/3GvJetGarbP7pHfsTEeg
0yuwHEZOQfCsdn/hFA37E5FSqo9mKL5c0M4KV7s1rnLtSPxYwX0FQjKGlPRlUmUhZKzYqLpu9fIc
xPksR+ZOe5EYIZ+nAgbUrqwbUdtXEx+JYU0POHs61Ybde2HSx4UlsC0zgDULIi99CaQbIX+mzky2
MJkY/rfeQT7SxVI8uclpGqz5kgCXUbR1O2usvnoU+zOO073RsIcYC8HwebzeJ6q0HOOnByecX+rq
XaXu80fOi8y6HIomuOT/GD1qxphSb/tsh1awJMDjUFY0WD/aKrc+aCqQgufxxHcYyGm1ToZODpof
i78O9+VaJGA5of80GtUn8M4lrEfcWMimkOP6iNkHXIsKniNcXQ5GSWBqLSSce1F5XuIlo/alKzBy
1wSDZo7tTmRBKnIcVEoDJHxCmT9wQPh4KSSIWGlF1it/7sUDMTnOJYGit9aXjCwxo6OJNtfSOQ/Y
emg9uhm3GpXjfA7ixX6h6+TcrvcJ232jXDL2wOfx8SdbEPamlCwkLbSJ2x+u/pKbeEvATLNnJEkY
RjgktASpoyVJ+mwVGF+2OEPwWp1jgLuh2X3HngAPmlFQ6Rk27H+LeJMjA1qPf5apHYCrVN2/dnvL
vjlowbXTq8vKr8VzQYOTEVXv8kKYzyR44NSYz7aA+N0rWchG7h7SSgxWP2LezToS4j9HiUJbCiqx
UIZvMC9isQK7DtjOVjIa+gPdsE4lJiV+ijWZmh3GgoA+qWlWuu0Q8bdz5s2Vu5ZEg6RgBywNEOxt
LavAqMXdCCPZN7429oylTbZjEfMEuMuKlzUN2dON0R2kLAwEUUNez8EwE3QzcDRorXfHbPVYsmUK
/Z0nYOsd0yLL2HXZeFqhxAmo5f1bhG1+9HHDQSYowapVX7vCBasxwIQxwjnUl5Vnb4Cl28tz8ivH
rds0Zqe5Tp52EjDPE2qDNy3Inp+Sh+EGv/NdwBI3ID8QwZDi0bZWB1evu9Vxic14XW5mZSmfphSc
ud0y1n9x+FASmCxVuvCUYHUb+nkYFvdzuSuSedV6rUYVLTgaGm40PjN/BTpIM0rDFxo82yX2ljYs
smfBornDTwNo5rPeYntYQ4VQAhreG4027n5KEymNrkSxGWS2jlJf8mZTIsQFT1FpbueCunhikYcf
gUrOypQXbrl5/x7jKE+aG9EYWLlVoLGhdtZy28X1EV7VgVc3klEVN5PsbTbGtFiWrpegqTeGRNUL
uaEGGQs/URXxDlei7d1o4WHIC1kQz/QvLnSl7454xEfp8EPKYwxHsrFsopF5hImd9Rx9B1iHnI7g
TgYMqaMucIKwYrecIE7I8qTj5W7az+6PNNKizWx6B7uGCwc+vzDinxxsP7PreX6WDHCQQAY4k7iW
WdfsfgZH/jp7PiyJAIEOX14fKq2b5o3Mt1RTNOPPaSr0a3RAolF91I6o07PuDaUMCbOkjsyIJu79
TzST9rIo6RsyhWoJD9TffFQpJ9qwbFY0l04x4KDySoCUn+VRZ3quThvZDIfvpCeR6JquEhBjq8Gd
CGU20GLIA181+cw5g3fE8AwZhshBakr85amSpbpnT8/h1IopeuUqnxoUZdhMioztZ3A2l1hes0Vj
J8LtzBHsPNUH0SX+yNxU76iWI5Ma1I34LvOvMN5JxRMW2BLxT1g12DPA5M6zr2owz5Az1m8u8Ui3
LSiKSgV9l7ZKTiypIH/OE1ktEWSln0Vj8xLWyi9jMRqQ7SRd6R1vf+FBqB72xPDmtGajUK6CoSwX
AIMtPIj0t4ugEVChsVBHlIkWnmvy5RejN6HgTCIzigIiizPid0MjUy5ojdLnVVnQDMwTpUqZG1vK
UNyXtdYr4nKcQaHF6Uajs3jfupO/nphhlPbl10O48Sv//aflphNDSbsWkF5fYdLZC9u/MPANIHEO
1pK2GFOiVCQTEKJWmRfoXiFNATxHmirXBN0K8I2GEIuFAR7ZTiuujpoXBgmx1UAO2Qkh9mTvYRoB
LwJuWDXmRjJXjfuMCqRdhvXI6K3ElSqEZhdq3hA9ACHDSSx9AJZoBK9uCdRqI7mxCQ/0aF6sX5FM
h1KQj9aU/7EZv/aJIzbF3ENBd0JFwuDcKTy2uGEf0cxVflBf4IYdHUBTHYy9s3tGIFVfQZacVSYd
3VucpqvN3rSFarHY7kgpL0vAQ7xHjn77/RYcl5nJlBeJldQyk6Uubc/3lQX+qIhAQAjCP1xYqMxW
TLhGd+ChtH5T9n2AqtD+yXobJHCQ46A16VkNvyvfdFWBu84BkaCZtCeOtft6XJFAugWTHtAB0oRs
YzHnOCWtdGWN9LzYPCZ8dUhs212PEZuu3ZplIUDNtcwNgYzKo64Mqw7RxYG4MPwNwJnirNyUuXvN
1VZ9aMoI11LEUzf6p1xtZcCJl+1b1L6JyybV7f66ZrFJ9bug0pWVNifrhT2KhHx095ii3H8qvcKx
MINSK4HiByH/IqlaOJLRnAZyHmVCBOhJp89XwXHXOjZH85xBRrlar4a7ggS97JFqZxl0/sE8GLFS
4HduoU6S9vll8dgXpWhX9WczRFYCtqr20GNV8AquyRCfnds5qWGoddCHBppWad4XaZYYNAuShkPq
D6MpGgqLqmTIzd0ZR2033zxveLCFlv9WGl5Z0QfOK2M0xNg3EThDaYKcVNQiSc/WTriz6Yrc03Y1
NRG34dLDug7yrYYL6PJC4UOCpL+N3/Z/SdClPumm5j2UrRNHc6rqlmpB28/l3HrfEHPV8NBF5v2z
5O3UB35jQMa6HmCXVvmyaw7Q6RoAFMQ9NVgiWlNlCPeM49IvQfb9Hm822k4d3SCQOs39LSf+F1Ff
z5OhBk/lOfi5UKFkTohuzPfdulRI3w6iZsFee2orKdxkLijhgUgEyHkMQZ12u8LQA/J4r3ZzHvPR
LnTyWf7sSmJLeUANgtbkOAeYcQLsqzIcN6X96qu4qKY00/e22BqqxLYn7RsPQ4d1K3y2W1RJOLJ7
AP5VQLaCX4LihCv8gR/99ac783iGA16CisqNNw3xXHTkIMLQ8Cvf4Mdmj6aj6VdJeQyQTJP3kp/2
iRT7Iw5J2GxCBYh5pg6Yw0scCVFltRXtybLI++nrN6Jv0rcvPvvaqTGwPcGiIJkaaK2U+BKBTPq7
jsT60Dc288S/84RwSHblx/0ZJdj6nJwS05vl2XDhmFtj5cc6q0KNF7TmaF2jdf1ZmDuvAeMUMVeT
VQFHNnpsYHSN4l6nlsdzvCm6PEbv0RZDjTS1O8lJ6QoQ/OaELt9Agpj+V0OYKz9ddX1F6mLzfle5
Hv8Aqck3uR2v4o4xz8EyvHCxr7hQhZrAY6ipssAs+u5BAlTJVnhT/SOxKrCEb1abq6lmdPs6bHh8
fpNzkSDohHKj9p80a0yLZJx/FrP6yQ4q6+vIpFqhoFYSVTrUeIuOyspBzV4jIj3Y0TjBw9YPo4G4
wZq1YxWWvuzypnYeYzGMGRI6trJ0kjOefcaSAqMvDkRSrrE8Dh/teIRWboynY+R9hIz3C/s6cmnn
UEVaekKMzOdRR4rmOojhoruBMmFjhqzAiLKVw/wTgxBpmVMFCFsH0RCz+boG2DgZcjSVdivqf5Tu
Z+PEUimSNLF959tF6ozLIRtITdwrli+UJOHpJGf69v8p/WO6ev3AnLuuhuf5jOdZf6m21IL2ry9o
eXZj1FygfNDiaYOERFKedcOY/5TnZpNgKXzi/UNTcloL4XZDjthPFBf5OhDrbcypbGLxqrR7yU0H
QA+PH99Hkb0jWlR1y7bfg6A/ITnK6GjNW2pjg91Ot05xrVn8v+X8vcmu61qgc8fRlEbyCxCq86o/
G2rG3TnuuKWyW4rgjl+ot6xIuY4uLifkmjZY86aWG0SA2y+MsGeyB6cuwtYSbRgiDU4MEDoA44Y3
cy/63a61UkF0olwhly0ElRXlqA7X32lBAHlWTm2JB/vDbgMgqvFDME3paHakUhqD57CYBZlxh6Qz
nxz4G+l0mqetLjEWWYN20VEXO7DLLQQhKszyUTzggqKws/SL4R8YWDO1q5bq6Mdod++dasdsyBwh
dwZfea2e53jNpov6qVh96ViaiRD9LqXbEmi416YsZMBkaf2MK1Qs+4TwAhe0LhLaGSIaF7ObWdja
o0K9wgf3fCvcogqCxCZJEaCc/Cs/1fuL+GB2uGZaXCOIgJpYpfZnhin3jF3AAw38kPLdf9knLVFP
fCACQlxcbWik5uRLeASCbhLpj+ZVRnKVjsfxByddogN6H7oTVqSfibLiD0aQrdSdVvEl3+5VcfgD
lYRT6Z6lnwGPGhapOvsx3hl/l706Zuyc/YUU8HJ+LSLAeqFUKnN+GdT7ByfxPBybqU48idnpCSgk
fHMGAHoI/mzh9TbTzuP9C5VOToKreWcPfotFHVzwlVClyo6uE6c3at5h4p/hGTywYWc41UKOAKek
Hnlu/72B7QEUoYGFFHeS7ZBuLi8I49pQ0nFlUND4qc8fjo4OyF3/F5by15rGTfBFu2wqKmqnW5Zr
GanPKn72aozvo0w64337/c4psP1uo/EGX+93csyrIE00iFplNZH8kZ8OaqY7ompGb5dXWYnAtzEm
BMPgWaFOIcoxV79cTXQbd1kJ7l1tTw5LI8N/VzBSr7/14cPnC70E8Uz1FgbKIKPVAqi8tSNgGnPD
lMY4jgy4qUaQd9g0WEVHc2C/B05mR4RXjBYo5Ctbe0qkTkXjGmmMNa+DUk+NZX691cT9McuELYk4
chj4RBUem9s1RqcyuYeB09B/cPw5YzNC1j1GEWPCXlyEVIYYvU4nUEebjYUYFSC0RbVW5qbWufcc
WjnoPrPqwOYw82RINqIO7zRKqVolPulEZaH0T6eylFAya05AkgfFuVBdxgezVJIDIwoJ+93v29mX
pBPA9mlo3me174xT+SDNGlSmTxE/eZxAgBLo8jgGGUNSLKk2JcRxY/sxM85JpfmN1fvfk0gRpCdt
h9ScmhbznZ16k++dL8v428w5iGh/61uijlo7An1xyDZJS7TA2AMeVsmBB7E9KEmWWM86oMpOO2UL
j/3xnkmE3PWKYey2ipIWXPKPd7ecUlPW/+IFdhfNrDkafUFsJH5f6tBhyRXag4sJYLrgNFjGMBS5
g7+iVngSSmTQKlpzaAffWBrfhT/vfwyInSw2vl3vWHbSyamjrxAgsEkVzt+mU/UbEtGVgUGuz04T
D3HWD0hgUiINcDYkoKd942XmBGMPtGC6NqiwXER3C1rgEocSgJegFFdYo7wrz8byIxiY+opzusTd
tyrRfTfMVgHqrc+JMS3v/e1MKdMxnZwTcgaaT32dSVwnWTvHWTqoqcdXoWW9QUj0DDY8YvAH2yHf
GmcXp/OXWCKMKKg903tuyatgW0WmvYh3V1KX9ENTpuCNx1ekhrV5/XL60VBCujhY5ntf7w1iBMtm
3uw9GzTMaPphbux8bqViAQmGhmi0t1KcVc0y2b/jyUrUI/6xjZYX9Kex7t76J3o+xbs6ESpITE9U
anLQsMUVdKOESm7KcjEAD3dTsb27ZA3VG0aCDhvKvu5nyACB60DyxjWSxmM3SJUU+Hdm5qYgKzep
G+9QKrQftp7h3RsczoWltDbZSd/bEFWpLgtQrrCW+69+43zGhyfPPdt3iWAI4ZR/yga/PHmQoPxc
G01DqAS2vqmFQDEzjl83D6bbNkdjt0QVgdq0BFBzcr7YpF8IxwUF/+osdJhSNg5+uTpUPBqM7sT2
9WtNyf73COLoIKitIjJWUnp5gnTnSz/IWvUIjMucIAhPmjKZdyAngiXPvv/q40vaM/wMkFls3C7Y
4dF0CBodeSWjvWmi6kc79b8lQXx1XsyJPSrrqq2p39ELMNPBTcDcXwfeSiGt8J8g13CdVOns1rjW
dDLE7sfYpb3EV3GnOaSfDha8XbOiLltZ9jlLnMispvT8G2B4Rp9YcsQlQsHkaTn8my5pXRBXsQv8
rzzr4XNRZmYp2fJww1OSN9bnt78IoHlMrCty9/mCJU7rXhA1jlrmlU7E2TD1MuZxSI0xm03fwzpc
GNj3I6T81tlAs+uYyD29+0asIp8gsUvxDR6yxdjhiQFyBTUwDlt2/h3k128x9sSNuvCrdPFtwO7J
t8LAEEUcxO/in/MBv92MkXshfdSYNxj1k1eYYoMiOy9J1WIbQuaUitz5akwKxdBHuob+nVvrRL14
mjyYtcY8URfmO9FWvlNeZkdj1zWaVCXjhKOq//6jURx8yfqXyeVdPoWH5dDzpw8XdJe+gXk7heh7
MlJ29ci/mEbzdyh2d9D5EsZTRPrfDEQm9/Iw4KGVL9M0n/ciDQwI8rpwPy2Vfnula/m+Jf0Suif0
sDzLktTL+PZOk2DqvBCCEsiUMfxP5atkCB9bFA4pSsgk7VlFc2W7NM9iKO2IvzFlphnHwDiY8djY
D1kRz0jsl19+lZFhZH0ciSKFenb7d6gQbJxa2w4Sa8mPEAdTwydGjF0PEcuDjKjLHZN/KNGp8toz
maYqbnl8erlp35equ0n+eFmRBd+/zTrpUd0N+AdCGIYZQxKmzMhTEkVvDF/UXlPTaCBmEdAzLyNG
Iu5kQkRZTNr+2CzNJy+JOvpxydlwAtPL+u7KBUsEvtADtdQts5w3MYphbo7XaJVnUC+MRLgmPhZi
V6bJYpieut2BjP6bB/sb7IbSePkqYN1Jtcbj/G4EfVrJvd2xDH3Wpk6MabJfIbgQ4FaeVPF8JwsI
zG79wHIDhRd36dWuYgjmGwYSkjLZZcQnc0Xoia/YfCMXtqAzNyZuGDCIKDxvJB7ObVuzIJIDiynN
ejSXC7RtjQcX4lTZyk5XyV2/8oLAk63FsZbILCgYGYGdhtwFPeTeHwQOmnwZP2oFVIi5zNtJBzgm
NVfojdkwoANzIqraE+JNWEy+FFJINyqa8Y+KfMLxmUsfFr1JDN7AX5CJcaAfiY5cNPG/ZUFuzY2X
pjHRvDEsDcRzLgQvTdsYgGXIJOcnEpGOcnG1Lwd0u0yMEVqY4zsImvvALgJniT9xAShplLN+ftv5
Baulj4cqXLBeHJl0qwTSqHpGbqmqnSNs6HXaRUARBEsRjyAZzcPLQ79N70GX31fgTrsxqmztt0l0
RRtgLrRIFMwu4wICIrZn5YEERwjquG4G8796X15Dxx2zZUu9/3qsr7yfnBqr18Et/9VQqijNkhPa
VYCpmsB8g0aQGgmcRBGWk7SvI6rLeRgSOltfpcD/PjQ9BDOqtjy+W8IZ4Tsgll1q2Aar9SCCf0Co
2Yyj9TXwMShK2BWWviNYYtQxogRsGg5q4eB92ywK9KDPH6dXxp6fgqwHLyx5moYNhzbnA5HCn5ZT
N+gK06AH6anWiuBSrmX/TX5g99hbff/iMQTYVb874J9LvcFSYkP9UJxMyKGsEEYgS3ezuNxT/M9W
OUTfUE7IdAIOzQLV8ykPtq1p9cF4G1KZzmv9+nMBGwydV/ot9RsNDZEKRc3Cj/dvU5d6zpmKr/FJ
O6bPn13+n7EsEhddgAEPjUt6ebCub/y2uajwNF355oXhzliaNrkCO7Te7GP72rHM2iUTLSKymBam
J6z2Yn+CVrgc/YApP5fjUS3MFfFHaafoFPdRJZ4afu6gn12AFJesSnbQkTks4ehqhx7FR8xnLgmf
B2xSFPOKvCLYsqXhIjF1t+BS/PDba5Uw+VseeC8Bsz886hh7IU/jP9LWSviJKdgWGpO7VVsI6+SW
2c5J9XUWoutCCJ8e+bAe8MR4R1NnizsTm0PBA59qr+7wVybhC0zgfOtn4COjJT88efGwmCHY3V1k
NZcy3as8tohz2bOaqDOyjJgtoNsoellS7tS1QN1Yu5M0gEpmSmB0f8SaznnrVZFt7s90d7kBTxlD
ZjcQO1gZnlHVg1yNpBATOQfIib7WVKRcV0nYflVslbWGIGFHRAh89kc1LRZBu0LzntdqcCwH/cku
5THWAF+05h/Ti/W7sY6pJ/UlaHlkqWtYRb2IvK7eBlzV4+EoFDFq2RH8yu0V90eP+ojQ/6zKMNNs
08UJ4JWbdtLdGI2S0vPX0unl9pOTSZDdXyyLBYGCPC4uJ/tc99qPaKK5Nb+1I0bW03XiIeZev3Aw
a0GDIMNcqYxYagM/jG0DROuIL3YD16sSStnMuX8xbu/w6B6rDp9X+xWk+Yqh/mRQ4rAMxrVQ1pxQ
3Yzae9AHc9D89ROR8KjHJJkdSQlBsR1La9YYoRf5yrQ9B10h6hF1KTlu7D0jq57aF/5db+bt2Jnp
2EeMv7X240Iep0g4VFaK+8k7JcMlwKl+RHMiilnGoLuF06YUfGGQDH/h+Mtdz86d7OEnYrVKlZOA
Vyim1CEoLSe2uhxH7idy1LpmQ+oE71IRcUqFyCXEZPGy+prJbUuu4PncmSDhA5A8cYGeT8QWm6BT
NM+tlcBUR6MP2Gassj8iEVh4VF1WDROKFgVlsnMhSILFCltU2A+xqU5PHbuLLESX4PwvYX5O93Yx
ITmOkMOxSAhy9W/7AMf64K9QX0zvqfiX+Yfyc7uBZl4l7MwzaUxkxOhTPe2Afkt0HOBjXrtKZrvA
8vGloN0CWWtkqjaClMMuhY6gCJrIKnP6OnPVMyZIh72Xf84W/2VQcbOm82UxJ5Npv9c3bvZLR8XB
R5BjhmtT1yY/MeeJVX/m8fgxtOZPu+hcL8keL3qGzYwYaBIVPH/JnOLIUWTu4Qqhzk+6XhpcKuFu
gx0rRTH89k1OMeJAV7rLQ+a8bKqepwMGWxwdnEr3AqBDBsquARxmSZTnuMZPWMWGiFxc8JyQuetH
4uJF7hrHTmvCy5AEPjztaMCoTCZfHnReQwljs3N/o/Cm/iptBi+behU50gXmLRDhcm+K3Fr6dalJ
r39K/m2oJ0YpkzNINbkB01PD8QBspOnsyUjAOk/d12aMfcpfdW3w/ZQkh36a6qR1LQldXdZlmlUQ
YXadRe1eJIbvLCMsLPPvFtTwgVl+1MQg3vFd6Jjmiiio5zy7+6GFtLxsMIyL62s6wZEMDxejGN3H
G5ERksqdLT2rrvt/yQ5PRycOdkb29yQH0SrhdEaeiHwRuhZaQYKht6bSD2ibrzjjulW06huGj2U/
L5LXmwGC6l2mvnuFe++J4V8URAuq/oHR26FgFWM1fnXqf1tVO+BGnei3CC+3H+5IlCFZNMDoP/JT
E4xOj195vA08EffpMuyjoD9zWA+eZQ8hLv03BH+WuXsK8gGUv7z4kFa/0tnEAUD43tDcvmEzsKPi
CuNa94TvXexF22se2q1AxgPZ+KS2DS6hyvTnQX1+mGb87ODHWA0h6k3gyE4cATmpaaGEvO7/xpZ0
YWf7CZ6gsrspeCfhWEWr31iF7KFeNDov7J5cGyzTT5PBs1zKl8k+MfaDY4Pyp7BzHPHimEuSVhYM
J6gP8WnqA7QAkjObYsGbwB/Y/v4hbfNxWXRnJUMRIM+g2XxJr8dWkGu0DiAqjU8y5YBrVJOj04YA
OGm1pcPBm9DMJ4UNd0siR0xo5Nu3RnN94PtxjVjfdXdH1ORt0ZQ1gTrrSsmLdVOCerGWURX8hshD
xCfz+Z04JJe0VUPMD8bze6xPgNehxlrINowpMXlA7Gq1jGk4/yf8RH7cO0SfqIfVIuMAR3hD5979
weLZ5b3uchimgEOqdDro4eiXF3AMYQ39nVIXLJHG58aKZRU2DZccS6SEpPuimUjxTYuBfYvquZ54
StRz0babSO0A6UY+CX5AE2ulQObSveL3kfatD31I1Afi1xwP4F9BVneo++1NhykS6p4h3FWj1Lzq
ntFJ70Y1uX7hI4ZA4gxnEmE3SvbKQFgTuI8OlUMYfisMS/Gza28WsK8rp9gnccv5ccdra/MG4O6K
s1YQ2u11DJUd5yjI2EToOtG5RABfXU86q+/whnrl2BbUm260c60RS5u6Sy+NdruukRoFTyUKiIvS
cXBebpNEqybV+G9UsUU3U6i82xev94Z7IS8hGyZQwQ3MHljdMDbqh6oz6Ic1mpKM0fnsajZBfxFV
g2Ntt+isiiII6d/ZHSaiYWf0lJV3Wfv7QiPwT2yks30gdf7s1JS8IW7AonMEAkpHqNUbEF+Z7uFd
YBMoPuaOrwfBF5lb/SnZHqNIKHBY1HU+Zbd4CvWND+diTiAMls7GiiTvqfmONnXJRPyzbPbK+XRp
oopQfvJtPVHfe64XdmqD47VkJPuY6QwfyQ4azBIyP/frTkwqOJAs3/nXCt7xgMNeaQxQ2KCTFyDM
XnnC1TAADmy7UxqGUGmEifokshkf6r474AxgU50jFEF8ofwze68QOvE0GWrTuDV9s92JOWFelf0T
4w7TJC+RhJ5pkTxBAdkNz3lv23qAruP3iIuWYzGzvhmcdY5Vp1Xj7OChNUNuOskIt2X3w1SXWF9v
+ienSvw/+XTDZspUgfqh0nQ/lmTkFwyBCbFwrzdmN8p2Ayp99kKYkNjjb/qwi7qK8f25a5i4lgQC
e2WOeXL0lPiYRKKllwaVPAacORoPnpQtPN6C4GXyAJQQh09JjbGO7opVbNOe85yciFOBSl+kVk24
PDFt/CuZw4VEG8nwOodnUjkJx+ly2XwWg9CpJwyxNKVxFX3HTD3Tzm58A872hXL4ziSFBTrsRZkk
mLAixl2XlxWTv5Rq9Nf/D3ckeGHazm7CO4OJW6JP2Bp7fYcDlKs8GULUkE3Fmx2SWgzcsqud57Mc
CoSD+neSsutl7fiyOY9X5yZkJvK+LFraTXJ6GoIDYk8Q07QPLwnSOZomvDlLWziibFK1zTZXThMn
nTRusyRWSi+qmXDbjcULPqx2+3TqlnNxAxQsfepFw5KYpBUIhqspjZo2r6MMdLXZ6cQaW8EfE/1T
29bROBU/5zJkpArSIDVwaf1n7kAtnebYxdAMVH1YzGDQ45Q1a7cN/bY0mEoqzWNXpRr5T5AP1jbc
xUi/w0nsIsfFwUXQmV6TrGElwRIXQdhWG7Br/G5TQ72v0aXmhBapjdGB5OR/YTujMQlYknxMuEK8
ExJeYdlwRc6Hn0xiIo80CjIS2oF2xzC90+0FyrzmUmimwewJA2kLeGrXZnavM29EMrZFZkbTFGCN
cL6YQZEITTcSOR3ziUIdj86xDneFV5c50OYsNQ32phJrLPLetPMCbN51asRgpTq1wPgZ5nmoT8ln
1Y4T7fFLPRK2UiJdiwAtiQDanllTqX5JB0UQwytEnoNhn8/6ZNTbH7gsoezh6Ldh2PmqNWfbw0qp
vW99aJSpGCElnjao+KsRPUPiawvx+pICB3ybdpshxqVu7oIu/WBpfEFAy4y4w2WkAUXC3ab6CpXS
69jMHPyZSgn7he0xwZkb7adxwlYvpYjO2suFRqlU9xQujjYgI7qITjN/yJ5hNcZa9SHmgQODXx94
nMz0gOZbz+f60kqNSzPsbXLPTirvr232/l4Z9UQtON3kTzVRbZejTWBoO2sF0zLM1t24dqDPdXFx
9nxled+Hz2C2KD0gjW6Y19zWcifDduWLl+lDBU4kx7R8tBzcVBmlvi9FysCiugPRnHhKXqV9NqVz
x7VgRoYzZ/j+tx26drX1PzgtKqh/QptVN+0QYKgtNCoHhOPWSLxtFqnWURlt6n5OpynUgUtnruwN
m01TGuvpvWpmmZxVCVapABCCCkYuLkVE1zWSQ56jOWsjfpsqB24bU1hDlNYLb6/gvRwbZdhJAaEq
1dh8PfiAF1wqVqZ31WSMCUZLXtvYjo0puM8w+8mkMB/FMSz/t3Ke7SPyW2r1p/Rwocl+RkK5yKgE
ZtUVL3fM1BS4BPeVNNEa5FXCXgQDlSd/mJvpG2qFYQ7wb2gRXhyEG4xNL0FBj8ANE1UmG351C3TA
3Ij6AFRdctBzNXv924AAthK3Td/XYfLiIxiaoX+MrtdZbtaZ0D1HlB2xZFgEDzXFMs+xbDFsB/x4
g2Kt11KcQKLnVd1wo4hX1j2AxpFfQWjYi68LFNVM7khCUgO5WZ7tpswG5basDdBbm8Xqn2WPYUlu
VujHGJNvjdTaOd4n7JYC9mFGEab/g00vmfX8xOb23yB/MgtkGrcxCakwCyOmMTC81v8poEJBGplG
xSQqUN1W6Oj90vcQN4Qy42t6tJVjomWoEDE5/JnrHmOqoeFf+12DlbYKONCxomrK/purHq7L/okB
0ZIWfsBUYoOjGdGHbos76cyJuG5+I/HJ/NQ4erMWkKvWksyjb9CE63aYTiZITRPuJlVdXgWUK8jl
zHsI1jv7c6iE/86amorBNlyBPlE4I6qr3xX9fGfiq8FqUziSjQJZWabMNqvnhMkaFEW0syJEjKIM
CJyYh54z/Nw88JNgar1daQsTwxYbCxyojxgaNLeF7tsWK1l65xY1JnsLDWP2aKdX9T4gdLxnOaUQ
jZPF9So0mIQ0jeLu7zwdcEUgwKVRGKSZixvYaJUZHZuj2AId5E4tYltJ/4EHS8SnQTKRGGoNAHe5
xNO5sFDTqzCHnmkC2iNIz4C/7rWqws3SiV25oo+LRH8fxQzjvWR9DM5kb+L3O+fRc8IW0EPfDtoD
Cvr3RDHcXaBwKZAOLjuSOJ11GIACvvTGj04a99ahHw7kG7h9tg1KBeVU6JARxHZ+FJ96jRr16db3
RmrdNBAgfi9mngS7liSVAU1pjdSFhbfeo7Yl9KER1RQVxs9ECX5jiivu7Kqbnn1mMffkb+iRihLR
pFyT/l2dprgxvBNx/TK1xRs5FjpCcDB/V2jEPSWzpmtcfFK1x8PCak9aY+kjpB6wjwNXmRjsKm4b
nBOXm/FgpFZKvN7KtLGGYyK/S3owrNu1QzX5JWPpNG6/tH04SK4FNm5izFJ7h8UlmbA2a882AhXp
sVA6LfmtiSOMSGNbAbuE3RU79cSL/eVwazA8m0lAMhgXOcDx7BFIpVfW3LILM2tyCmagYj84nvZP
lz4GZMXDbR/wxIL6KU9RsFxPkHUPm3c4QnagteXaSVInw7NaJIDd4PiCmrzZGd71nGmD9ycIe42a
NJxqTI3MnjvSlIoTDm0bLkfxf4ZHFdSd35xwPD2coNIJ4V9urbtvezfAZ5XLxpvu/n1wOHvMZmMY
cXHFFYqJAu8gbcm0nQiM5dOBWm3kBSSiyy+CuYlQHosHbNkDER50wD6ZSl5y7QXL1D3aS3+fAzyz
GCST13E7g4SssQ4ALecg5Vc87irdxj5Mhtq+g/XCZawYFcnC6z3FubyZ5K24oBHazD/hfDTwWwL0
k+rXuU5G68ZuC9c4OYJZXCF8GKzByrax8HQHkFpy/+5nFR/581IRLIs5SggPy6ptVf0u+An1/7MT
s1kO4Xq+7GA/F8P1iNNLTJo5zugs1Kp/KmYLKBa2l0bwjCoQEjmaROP7lvKJwg6XPLZMK7VSlPUH
cvqpBIBwG4LZQ1xoDI0mPuc3agmIlrZBWHHwSxE+f8NdESNyv+xvdlADG7UKeLj2wtvT0YxkkmX2
Inv+qJc9Gp5MoYjlU6og0R4prpq0WLlEqp9jtpiAKFgIYIeG8c7Eek1pcm0C02XLUtFjCj77qh5f
TqpuPLJUG1FwDM6C3N62zOYReYdpKlNgK9mAdPRVaxZSPupnDOC7N99MUA6U1idqs0TVHsQd3X9D
X9EglOZs5ZSyAnUobtLe2lxxcA3FsSXI2Pw/9F0LmqnYnfMQdamfAjIV2Z+3Mq07FvXwj35ByyWX
5rDKUXHRTNTfSGeCZLikVcdZNRV8uXI7UCYGqsnlG0kVPLfrcijsnS7462cGkNRimkkwV94NbNVA
lPyEfTKBPEv3rILEXQ0NgZHuVDZhiCg7As1bS7ZHnK34k6S1MDzVjZAtv+4wiBjB+DOUXaB7+htZ
9eyRmREzOpp1lddLYu1kVtZ8rNeQ7S9crZ3wagIUF5UcZrdpTbsv/7lqch3cj1n2QHM62eL3Y3K+
YTDqhwsh2usFe+4c7Gg1Cqt0xR4Cz7vjJyfQOOMr/ya8HUKE7mbkWNYZ6zarjinVer3iAKdL16Oe
e4z0pnHLn8WlIJJQ1alTiPT86WBrYzIK+IGY3KyqCAO08K2M80j1gWUGGSQUg2m7+gh2LEHLCXp6
nUPCmof2q/aY/s1UVwNoa9muKJU0OihpO9hUUhfcJG79HwIXOgbpmKwNg1kWLeXGdIIwqg534lHf
cHXjn05zu9ar2WmkCkBHfOsNVTAqhTTOzWk5hMaSnqcP59VAkIkJjK0+L2Lp0Vb5WpeAmIcjVSqs
VQAEmLzOkXsf5zmXW6w5axdX0k7tYrZMsibyDcC9iAPwW0d3LvmBgOd0Lw/a6M1A4loHrBVKUAbJ
NPTkaKmle0lLkhAdvm5nYaz+zL8rASohlxnniLQPDtWWCAgUhLSG3jc2wSqM30Gq4/IiZJ2/RrqA
yzuyQyANmXCkb1Et9R0ncoVUi5e3JnQ/5u4naHEdKpyOoSfjfoAbWuhA6jxHQDSbeXzbjvfS2bOD
QdVUn5Bu6NwhZI9lcDBvbR/FBP8Etdj9WkvNUF6ab3ychDniczURjsK0D1y6LfKpRcq39zegteps
yi5+ji8xEuv3ai7Z/NTgKlfL5TgqjuSs9+pRU+rGPq0O9lNGQp9TdwX7jrsgdYRfIPWEJzJurKzh
BwiOzQKOBjFyRlSK2JhvETtlS5nnKPn8s2mChqWnCG/aCqVxViEQozjX1pETj9sgM/iowkRQSTKO
3D62aSSKY23kNscqTO/9aK0cChxYCqpNj4udFoSFAbacMgHs7Ine7Ns54WN0pk6oA0ZrCDMsK+9w
A7Lhd96Y96DKEnRmAbQ5jZV4gKnnlOn7dXqmyfbxlRD71Z2sB3wOZUnGKiZyvBRIDZUIdmMr/8lg
mRw1OywYvsNoh/zzKrqIghUERGKwFmE1AXGyk0nQGUvbfigbhfP2HSncRyyBvW0j4A/PxWgQTMsU
V0cqGL5yKssxL4Rx45HyjoFMYSj2KvNEXINfp3QoPLBb9Z9p+sGfbleyQgo9O0FBrWMOLLIxXxI9
HBJOrLVOuyB5Tzz/9GJBq5zn1KZlULfwAq5rQuMqzlfdrOj8+FeQoYFbM3l/Z5a9ejhytmwrhol+
x7aRVu7vrmBj5ssIZpAYb6sWz7cR5AxscUbZS+HIDs7MxzwqbqtnROFNM6dzeV4cGr4iWZfPWZaU
utYV+Vaf4NsYQ6srAJCjwzlHrktw1lMR1D892i5XfNkJNMCulP6YzvH5TwvtzJjtkDUC0t+umZci
te6l50ZnhzErPDwvjWdLyVr8BTXTG6YYniKGUXVMannKjUxPgcZYYIDP9FCG4YP5GVJL8hd5QvSS
VE/gJosWRTB6MKO2Bz4h+inc2CmTue5Y1xWsL2OG3FS1oh/VH73L0a8tNRsiYmXcr6FuAwz0hOPh
9loCGzE270tFRCcSLXpo5srAEfZ2wxXI07xo3mAA+VbXU+Vp49m4yZOnwXOBDovcG0+xB/Rg6nAP
UhejMW8+DxqTmGrYQa3l1zDsZNmmKbt9Bcq1GmljjexI2hJBN4CcJx7XvztrtSM6AyqtCjcheQ+Q
89FjRnsJli21dgN7Nd5727wG2AxSmeB19J6ydpZdOKAIYZg4L5B9USJh/k1wyf7c63c1/fYJqwNx
vQVU/yYxfCaSyvSdFSNP6cclw6zxFzb1kz6rSOs0yQvKXLEFKwWkdQkp0XwJcF0J5Xcd8zJKGOD9
cB95j9HO7mZ1LaSmmTVvpBYKafvD33crH3myOyx1iaMuvWtdd468SkciQ2x7YiQ4FBKfNxRTb3qJ
W8R9ARpROeJWkhYPN8ZuTa895p6wBt6thHKngrFKEJR7pak1i2h+UMvvLbsYdRZKr4dXlRds0HhH
k4xMcKJbIpXoejp5CCw7+djXOxuadtKtoJ/gTU5E7fPkt4epQ4iMAR5EgkpGuA07IHOFsMpTHs07
b/bu88KpadHVWvmgwG/JNO5mU4NT9t8eI2C8qeqREEOkjk7180njqGWK3b7HcclH0DBM+vWEjNdR
PrMzB92Wnpz+6ViZOEsVpbfRGnkSrbRY7eepEyYLMB2VzFp/qAoMEPRt5WQFToeUzzLMNsDthb2m
bPPNByE8eyyQBbrqtNvB6AL8IhPtlQ2ICJ/AfYWMuGRbkdxRt/gfQOvgRMFTjq9OVphSFwLVLvZK
qWSRLlsQKp3TPsAuIi+YcsNZdOaQogV1mgV49IdCOgDuDOJVud9oQkxMqzcO8iYlJoKDVoiFSE2Q
oJsH8KjD1Tmpnmzoo45H4LB05cIHUk0pzljk/A1NJFcPxVTdPW+sCzLGTBCuZUw+y58O8spHosJS
YWgssrjxp9tFElTPHFC30XjFK5ut6YRyHGul+74B+q7GVndjaZZufYkViqHBI/s1IIjHicjbGD1S
nmVDaoWglEfl7wyYchBiIfsO4lo4XJ7pXpzhxHkIKuC7PWvl1TLZd1X7Yz7KRCN+08ZiJxcb6uur
zI0QJhmDs86V9OKhQEBYO6KnTX5ua8pWdxXflrfGnH6aLjNVNXQAxXyo2o1pIhnDf/SNQlKRNMmh
S7b/X+21uXFr4k92KvInhPgWOoYKsyu34nSlAxaC8RsMS8CegmJPYQgsAcoMaL93bKjbLXddh+KO
tA7HLisJm7CokQPD/+0X/ofWr6UqUuOTTnsJux/ff50sOZczjgV469m38kdkS6ryKEK7vjLN/shj
acCsPJKej1jgwIj1dZ/e8a+RUHIukAhGI2OJQvbbFlBFgdaEmFReOx//YdByKqSB59cRoQbRAQbG
G5fj+A52AI//DtKUYglF3bbVriR/q7AiikvevSGe8Ww9plyxZ1f5gc2v2MjWNZDv8vowqI/DfbkE
loQQQF7eGyMSmTV/KIGGvfJ6I6A0S45wb/1b+arm3FSLF9EZ/FA89jXt3rRbeUlikUiQw5OA0DlY
yL9Ro5pbvX+iXlCmZmH5eatH3Lf/GkIb0Fc94EifAzrQaCZ+e4jvbzbSa9HlPRca+NDINo2Rbbfk
l1gOCNJIMJxl4x8QA4Hi4ZiDlit9HJGlF8Q/Hp7FmonqCr0p84EDE2czDpEW1p3q3FXQGjbwLAhW
88ionmDVkWQaSJTgx8G5mtVFg9bHFYWe4g9z9kIvFxLZNIgwardQekbOSkkTc+mRh1MpQmTlDtD5
p9MWthR0b9nj8HS0rY/uY9JxkyOAi5KAmVNCO1Vw+xqc05ecvmWMppFim2tBXWAS7Ux5r0uiZljR
CQyXe3FYdsXx7QNzffLf1CNWWv/e53kKuKkCVT2SIikbUMnKPSDVcE24NMo/x140S6ug4YaYPyWD
OJlNkPgep7RoU2gVAVAewVCrV4bdRZd+ng7UGP32Om9NUmdn3dKHPmGSFEz6Rcathn3iBCNL4uUw
4xMvYhvVT9gydt9M6vMZa4RLmlM5/U5GSl1WCv59a9ONsKvav4GxO9m0lTOqPZWYzuuXTdAwvB2t
hZjJjktEULfvaxRGpUQb5JdrL2YcghhsC2CKMp8u+E21N4FciwzLfe08CHCp7IJ0umwssHQpuqxJ
Ci7QvYtTJHCbKS4LX1OqVP+UVbzlPfi8HQLHddu7Mb/mZFKzA8hfz84ob+AoVBx7K/Pt3iOhxr3c
NEP/x9qZl/NOXeTunMOWtzgL5ETxHWD1niJU0f8Gq/HMrCoyVbuwwD2Ah7MChpkPDUfDkB5rgyEB
OZtKA+FegSTeXTSpQeeRkAcNAYtqva90NUio0v39bubRUZg2+7ZiWv9IvduNU11kjT/AWAdl9GyV
5WLQ7kZ1r4hO8ourXyzYJoYIBWiMJwf5MOWyZxH54kC+uJDPG5knWK+85oD1ltDc6a1TvWG3N0W9
3Up2LH0lb5yrbcbfTBNrB9KgNk3fO1ZpwLtq+DEp9OPfXbY0Rgfr8OvwhlZnzafQynlPKt5gOhxT
fly8yBUSV90ORwIJ6v+Fsdg2pMrlcy0NBC5uJJXSocIA0ZLd5ZtMGbeULwN4wZ/mNF2jUCbpc8To
PNbdue8sV4aV6UNOJlvQhpnXmDJR4iRune3KToW8QEB6rUKHVUKZ3kMxa3Dt+iBi0YNjL6ppdNp3
hxzGKzBAuF8wXip81lHGYsec3sj0+EDndDEPYOALp8s9PFGfFYpLXXuimrzXGMNkXz0LoIn4fLpX
AHEHRCcLnBTjC+Mq7xKwlK4JjJ3qYRn/EYtSnCNjIKBdgWEKwIfG8tT8XlH8CJk+D10bifYktat2
uYpTIHQff3CaBEEEFkOWn5QUEShWQUrSnODDreu4DZQSK88xX7oOMDWRusC5VsZTKNdzjEz0+fj9
C+7ScoD5UYbYjgbhNYEK7lMbJgMB5fV2OClFX7Wi9Q6A6SfP+GrwsqIyR33sLOlox8gnKABe1IlA
EjSkx7SX4Twypc2rH6kTx8CdrQ28albSnyM3XElFnugulHxktphm003r7uvczAlqnncoafizWUnM
u0ArUFCpU5249QuWnj7k2hmahj+uYzLxyKM/wWlketcG4XS/ao7fVSCyVch5vHakCE4pW6G318Rz
JqcUiA+/oO4hFC03YzwkabpSKbRkwS+g29vuXrs18CHjqkMmjNcKau/dccmGy3m3/zxV3j8+UTuN
05hUY4GXzYEo17a4PrZY5U7RBbdBj2z8isXqxxlSRWSAceKkB4U6xm/U78tpm051/FbVX2ddUzgT
NpFO8oM/4OeWZie0a+Qt2o6qvviesS/UJN0dXj8qyrP9Ks/niTaWSlELZFnni0SoAoLdqWEJJOVP
k8UqXL4nCy/yWykxD/mkz0jwgv2nCKEj2LCORKh+PfGm21f0nFixhkpfM+cprB2wiNBX7TNk++0B
m3xrIzwaCLG2GNSjNUBTHdw0noOrom/sr/7BVj86e0vpgbYQ/K3HbMJ86nIe8W9fipRc+0prVxdb
POkCh/N0AY7ulbG3iVkZjXUwZyO3Nu3SueMYmeub/+Ic+v9SkazsZWGWCWv2F344p+ghwqCU8OBw
R1cWLmZqobBduVdE1/2gvKiBvq/oGsW5J/dLtmeBWzTqDWbfEhxnnT7G+Pg0kAAt/XfjDuXSSGIN
xAblt501SR6PrXux1Gv9ANRBvoHPfRqyh73IjKLKapAhrtclbUMNmQ0H1R2u3bqDrjBA1DV/r3qy
ye7XAO2toGD6fEA29tibFf/8rghJLwDs6dJrkT9jKLRyPz6MibPUma4n6o7KFXjYngO2dVQguj3S
/aB1aTz3OyB42YT7PFcNZrkz0vyNpLo7alb0DPNuhSBJNzP7JZKpeKBVXksq9kMcdFTyglPK8/E1
2Blo6GcRF8zDZnHhJ3sGqtVwvua7OOoZOCq+BPpmMlSYPE+iQ3O9VOy2ohIv0uNU+PWD4ZSGAKhG
s1el0K+/vmKCwXz9am/mSAORWd5tngE0ee/Cf5DBoudZCdd/WuhuQEiIgWOSGmOHSyrirw+MSIk5
t39SNniF5gLAXDkbUfUgpS/4C1zLxwuVXnbQMtJrs+dCWHMi/xTz4IQGicygTaJcCtMb+RPLIrrH
wYwh59m7AgT/E10E1QS4uGUjwWtkP6HVCTpzn8tsg9rTBEICMOeDhagpIgg023y6sJs5pElph6LA
N3eUOG4iJgrJRPerULUDCBS1cqr+STnbbuPs7duZUyT43ePZ2sXv8Lledx8TMpI3jXJdyJp9tH7Y
DzCw+0X5w5bDLG9MNzPlJcKtrzoyK5qsFtSAs1Er1k0rWD/5d3UNBCK/t6qKTxnKfXkHZNYaMaG2
bhh6Jb4lhd/Xm3rfKk1dA5RNnjDP/D+wuCmvysF6oXa5pGSH4e+u+66n79qGVaze7X7TEEg7BuzT
eqsTDxrRkvX0wr2OgG2ujqq7OccJAZjHLOlfHbYZqVZIOPyd/v/j9t/FkvipkcCjjDTJlimClGXs
f7yDc758xw/HgdJhgzkMzXW3Axx8ry3xSiAedgKD3Bs2RKKevDSNahXz0+C2snqHLZAxPYwGCE9R
jHoiRHJO7CQof8LO8e1wJ5uHhrLg85Ezxu8KJXNh83NVn9RE6WJHBbu85HOiI+VoElCX+Q0z3iqI
Ji3cHou86Pd6xxB2pHFgSYwxpyB0CG/3eirKNlljZjZfWrgLb3ujVW4dg6uNAahWP4LCExHpABfx
d8tYfXItpzrUwEXqiQcwYsf7x8rNhMT8cG3zPjMdD619AkjQ87AHG/CYElbZLioMu2LzPe2QuLKX
o9OsmTy5aVxYOwVAmPywLOBkwBZ3V5ci/fPuXL7ZfsEngFvhRNah2UxTS0RG5ElOBAX1CmG1PGyi
vksYmqKXbk5oUon7FkJvdATokF8uZYK9/ubb1THQVO3PBf5AgIDXCWdNin1cYuTJcDw5jMHTtHxp
/fx0CSK4xsTGD1T8M7APMTbC1Y2AMQk6KCjpbA8mVnsYNOBk3xpllc3BGD/LXulf0iYQJXdmP1AO
hVIWSM7ayvi9nvPsYLI8L6fwx1+bKOWEBksbOrtVzLdasEyTpczVuvKZvXfdJ+Dx9OoEL/n2qigG
4SMb0I19sAz5NYaDt+nYZbW9BwuaYjdszWtad00W7/1Pj10ZrmYv8ZHEpQA3ucGCAFYYa2AmMI0/
zwkGeq9HSIHZPv4UZA75RmWcDmEPqyCFyQgG+GPIcOnNOCGm+1gg9fPFvVNeR+Sn+jdDkyrQYurF
z6YGRt8s6REig1ZlGFk/ua8JD5Zf3opS5uH/JFX0w+jdbvrImmvPq7LBfBcM00bA5Q6+uW6mmBoS
yHjtyTALoO31yrA+iPBOQkcJ0g3SMzKHXSR60Dn+GLwucaKtZY3r675rIIqGxt7TzSRJvyRyTmax
OVpqo4tPA0ar22ggYl35mq/MDjSJ6r3VvUPdBwzJ6s5CzxLmJX9entsOVcerNk8f0ELQPzlOB5HW
rEHyWZIekQgjyIQ19JT0p5tc3VUiPAulfQFrw2zDTGXxcjuHoJmNLUS48+ys32oZRj2Q1Md7d6aw
KHIaThACCOp3eGV7v/JXgMfU2yGnOUtp5SXD4jqefs79ZbpAUxX3Uoi2cqkVoRerjBqcolVqT4h5
hJgEqYyhte2iIx2Mp3l3cbQPUSC6rovIY3C/tQxlbHzLC4kG6nD6twQZpEZ0C61L9+KyKXw2xCEN
okqTEFSM3KGXi/XAiU06rrpdY7iJQd7Gjdg3mqSuHAr9Nz/8gc2U1RnRLLfz5aWZMjKYxoI9wvBg
mn6R5HgTd/5c5sSqt7zvy4IooxyO3xZCakfQ9S9kAoF9q6QSEjuXLTNOXRZxWK4WYBrVAm8Xvlz6
FXknegSV+PuiikqbhZ+/CTood0Vyxw4kyJLjXX4ZIJyzsaoZa61rwM+kx++g37/15JBVUV9usIT0
3p4omFCv6eQKbbCZ3Hdh+WCOoD/xT6kgZ/b9x+y+Ln/vuJJns3YxCrWs0uNw/t/zpjJQaoAjhmz9
g3iqjB3M2VFXUpWQyw+Gwt+L4o5xdzyLRhL9EpQvY7JW4OtcJcFupFBHb2IF0Ed0lClqE1kQYHQS
A2tLqJR97C+wviX4LeZqZ6lTNyMrxE9MO13Zr75SG/BWiO5vxTbWKtYQhcFaPQA4NW7nq2yysMkw
xRB2ezQrnr49WvNCAXVeVgWoP4NGaCXtz2pnaUCweMj+Z1aVwhaqVcellAsZWtZW21ZJsPBJ5a6Q
zK4E4t3JM4F6yLWMXp/ENXGvbQ1ZU3mkHXR9UdudgwDAIHSCTgFNjhAVRbH80Wc1C4AfXI643DJg
mPaScwiVnVQmCAWD5QCbO62YCrJcfYh+VxeWel8W3h++2fbYL+jHoOWTiAOlvO2JAUhS9LV3KAWV
xXFod+zWuANFU3V4n8aYeFWiqQ1eWIV6bN+VgzzOhbDmxAEDGdxhPTOXv/wtmLyPOCz54+rBVqEL
rtzfLRlpGuxZF9/wzCHRTJ2lr1e17sQTcg/VbEpZYZz5eOp5cb3+uUuhnbPnYr68qkI/UC5CMIv0
tjTtDNdVgfgqrKERPzcBXb3VY+M1d2xAG2jAqikJ59b1EcP5GsEnnVUte9jgupy/tSB/FtEkRy6D
hXEiWcpDazSJwUxTwu9rz9xJ6+70VrE+WufbvZCzUsAl8SXOMfcj1FvENqcuNKZvfQXNeV18VAAo
/H//cp2aAOu9bn4uRljltixPPH+Xsw6VRXNYcUT3ed202mKpPiViblyEdO0CtC64ytFNE6KBy3nR
laio2N/GUk3pJdbgJaTFRmf/gkvhZ8YcJL7b82sJ6CXDk0dNyPftL4qAk8HnD8wwQz6NamteeuMu
3GqEGhwIlDAB1oyRJh8VzAL6FKOVZ3/bYWIjHD7cJPCAbEw07ogQZazPt8KpVV3bOp/zUVPi0Bzd
jXSm4/D/pxL0+MWBiSwOlcLFo4ZDKEK9b6hYQC7Hoz0WQJK4TBeQj+7ijkW2yI3c8ihuBz66sewP
So1ZFxEFxjAx3nr98xa/9QEohYDurlJ7eV0evbOoHQfY4C1t9SuyZ2lTFs15R79xc1sMxHMFGzPF
VdL/zA0HcB8U8sybnAN1w+82tujwlNOUF1kH5n64Sl3IRkTtXEKKWW7VQYOapQu8Q6yJZ949+pR7
0YZWt+2dWorEOLc7Iuyejh4b4IFN7hWJnnz+pkfpNf0ARc41RRNhRVuo+Yzae6YqHBtwzkXhEPic
IYNLMjTuveLaxKeAKm+8xZD9gXOo6UxQ/JPZ/vlp4arq7IPwjvEyYdVO3rKuPRUKb46pC5F60+UR
G4gEIDL+xHOso2WZNBusjzSHBeVDOmU6OrGwlBMCwqm0Hk7E+v4fcFcAo0rWeUhJ72yJOyZZrX+/
pcLxdCyEJ4e3nk/Llp1/mBfmnHdd5gcCUaZS65Ef+uMQOpDmUhRIbUwOHiKCTnIZGsbNR9mOgCp8
DgWnEdCnPqigvrlNm3ja6R9zcwQf+lJy82RTvFzkrfjtI3JqH9jb92faqISorn3lqvpsV8Xb3P3/
PMJm6CJh+73QdIATZsXzo+hQZBAPy4mmREZt+aOD6k9bIaD/glnkAEsp9f+tC3TRsPr8VhW1dcpj
0muDedwOIOnVY79KQxv+3XNrBpDCxBZfbwOS25C2xZXqfsoe2477o9gA4x/CFy1N+yK1P5hEPC+/
VEuZGFcbj41Ad1HrzsxR1zaG63M0qzgAq1XOPh8CM9CP0FBtu4E1mW9vTSfgKQ84IIw+sUAmnwDY
vR1hJtYyCnx36i38IFzdosxnLIDG2adZiGrewcFbp4iSAcQmEQb7jTJeCVaLq9wSv+tq/DfGJlBv
HASBqAu051ZZ8mnmyKPE19tlDeUXo76Oc2lRI1FQn9f65bHSqdT0PYd9yqMw0JZ844UVSRraYgG3
qB5t3Pa6DjPP6Aja36d3Yy0JKkZQVT1EHmXThSY3uV1qCGCXR3EDjBKVlndYNmBOiF73H1VQd99Y
dmZW1rfOPgMgRS5x205qoH/i3wOtsEIjOlktaIiI8JV9zcKDTXT/HNUVc8T20iC5ij/pskIxnqzF
S4+UVNp8pwTUlulqbKkrE85xYlVSdT5GG4d7q+LTQyfohw+r64mVNHT+RV2r+21ik55VqC/vuizD
kqrhGP5O4tGJMmNQk71ZLQdEM/T1mK6KLl4KrhjzBA9C9D8HNdTTz25hYbwscx7UnSVuu30W7A2Y
BFtq8AI0VQi0ueRUHMqGYdnEnUrYoxkcJpUiXJrxAl3nKo1oPKwkrimQ1CeY2XKAFae/jJW1D9da
p2EKqrGifpmtNxOacLB1aZv0TfRwcMXRMY3RtVanrutf/XO5WoeKLDYCHEiIaJUmpc2SUqgBIkc+
IWxgxkp9sXfdUr37PF1eAQASNBOzL4yPW+Ful/M9ler1hZcMcf5SAquYCT2acx2OZW57BZO5eh/i
XcKcobPPHhKZV1XjhTvfvW4G/ucDyg8Fy6A/raf61Xih1lF/iF/Xa79P1UbzvQU3kGS4u1HeeOkm
W04jor0M4vI/I825dgn7u5PQN/DwbiClZPtemxNFUW+yT217ix3k4E51PdEi4I85gRpdUHBDAI36
CpOYAygDSANh+6wNzLuT4tiGwD3UEoY0/7qvILjlYn7hAKaS5CuV/E43WRF2/vITPmY885xHy1jO
vfHN/2gUvluQayJTlzX0WI2354LUPTPfTsv9l36BMjP6DTA+uxVN847qb5jOGBT8CC8vF+Kzr7Cd
/oaFmttb5Afq750QBIicO1+DlE60HpirTyytQLFbiwh8ig2ncBky6Q7TAfBVwRJHcfXKFiEgySdb
cgQ5A+7UrD2tDlsmL9gcpEVnIY+UjviCB3kgp7KsLp28PMbGfsxK/6v84C5Om/ag21mISYnV/8m+
iSHI+t5iCIgcBrCu16KGq2mrLrhWI1DV44wBT38ZWV5UHij6ONTf4Px1MXDvV65njqvTMuCxsXLv
Z3y0Tz/twra8rso8mxZa/nGniOCVr6XKyMfqyzf5RheKNJlZLCcz5aZJKyxbhkDpGoCAgDYRxsZP
LHVCJHmuLlNMfFGC5mqdgeVlMQuO3tirGnyAaOJSneUAOIPsg1Bz6dDSD5RwMpW4/Yg4id/cHgFy
hLWwAybkvBXSvsZ+B7EoctxNXaSHTihEt3kzvVwtLz4eNTBBgUB9/q2BlZz2+RQ7/W+2BPZhvZOf
1z/KEWInlooQPHcL7P1WwmyNRFAqjOEHDqs3KaMdgUO+9ZIh5tVaJw8fnjFS6SYyPE/k6FSQ1xAj
DbCFfdH/C0PuSyDnb0FqHQmCzgXZVben7hHT224cWYcGBlrLjlgbqVaP2amaMJVheYrink3Xco52
xzHWpLIPQUALNPbRUy1YxBsG84OvU43jn9q1ilHgBiPxVSEb43CdWz2JRDx6S2AKAJ4A/mkqr5MN
jNVfcH7v7LKU9cohTTMgv6r8eBzNLih9mOtbOgZeCaxiM6Bhs2ozOoOS8czjFpUaUjdjamMp3LYh
evVIBIf/Ofln7OhMjnRn0Cz27+OPU8JIhu0vJeG9FCQRRot8utgUssGtDP4q7/a7NTBIEolPLpSo
Pan1enm+iz/ZBkTeCgE4JmelyYI8bENCMDxQWeo5nibsUbH54h6Slv2J5UlxwuBYQ3DuxCRQIb5M
76UJkH5mqOfJL+aYx8kuGZXulGBIFIFZKLvgRP6daTgPvD+oHchTI9nZBnWK2s9wexnq/+bpOAfN
qtl/dbQ/Kezw1mC3rGJer88V/7IUpUSyjOD7GfasxVmRtAnal414eGK8e0ocTUgvOpCDqfOymxJJ
ZjAq0FTdDInn0MTTQsDa22BpPnH4zXxhV6MQk539yPbITE3shZ1WAz5crMGaESnGyAHWzPRIQGMy
cjE0vu74ZL/dcjgbXsSBPJj4AAURFzf3CrfxrRzpLK/8gld2Y2iIizU1BPb6OnkmooateVtfwRtR
b80yrQlRFb9dGk2AzsKRgXJD6B2FjyA6ogzlZX5vu9Mqe2ClGSJvyEtljSjqna0lcUF39CYhBVXb
UxRJ7g5DmXmhHM2IT9fGBr5lz7dUSGKkMN64n74hk0Vcy6dPfbWtklfadrRyRSt8GFgeoSdN+Dwu
4zJYENiOMAvKb6lH+uxpJrgVq5oYSQm44KZcDnE5JnT499TVvTMiRq8XhaYfSACU6qauzdKy/u3d
ap9K410+uI6/n2zTgUWYAd2oJNd0JOIfDJPBhhhqvJ0/CFb0VDiwSqdj6ua3I1v6sohCs+C8ybzG
XuczVbxN3W8nTjKneK9taKApgIoYYOKySk5lw5U8zee2YzllIbY577rBNc0Z3coDxaR7LK3bZt+/
JQuKo6lDHBJP4d5G7WYc36WGe1uv+jB5Uv6gCtHv1+1V68eSqW0l4rCVXCZGI5+ylScv66qxI5yf
8eC68/IAkM9jELGzng4ohl8YDkSwjjJOTx1S5GuJGm2U9AAGATg0SDZTZzTZhyxB3SSsmoaWz5v2
xmnaH9Dadf4GvnYa/35DKZeRDcvcOh5lrVPiGRUXQ1Y4inSJhjRmUhuHds74snxgRP3wIGmVJxcU
mSTVRDei8gKrZx9HGJixECffGuQpQEA4yZZi9QQhYwO7qHRjbrfb2YIhcJwbQh30TX2wTD6KRfYe
illELAtmw4rgRtC+/9wO67Ut7JxYMe/bJlp7Ey9NxHETMxBjZsEnHzba67DOAlvu+QRKkJYQe0qF
4ENhGg5Xmt67zVG6y02OfHgDrsPhk6BUZK7SDQ+tbwlCiesVfhC/+kZchbLyDuUzkjzGeIw1xwcb
7tHMi5hSJQUazxSIzgm9PwGtI+mOH3LlIEsXVHe8HaX+2ypn+YEjPe8Vb5QPcXhmkZNfH+28goJF
hogAAaG3+ZXSB2jKSL/3CpZnivVttiYFX3GLya7+9GG1Osmqqz/t7fcNYFCoJUBw6EbMlE225Sgt
v+i2vnaSwDTxzzXY7ZYRgwY/SwL7gqdS/aPyWIBOwrEB8f1Y5nwhN2KhfH3yPe76mQNgVnloGxX4
a2I18qTo8rOfxkJgF9UR5BqibMpG/8Nax7CjLk+i4OOEhaHldo4SYLlFGk12QkCwntOoFqnzFGHj
FUbwUh/Cavk+qs9AFX36G/H0b+d+74zFKa440rtvCPQD2Fls4RE2Z3uDrf24D2U2GFvQfMOhqZQQ
lJ63KB2fCn/bwk5EpPV/5ZbQv6Zva1jmkTbDFi6AqedoMjzmifdhjYf5/WZ5wb8Lpft6z5A4Ge9b
7dTsg+Bl2mUMq4gI5vEGS8hftQmu5xiyFYUrPkwKKYRHYouTWkXDwLip1T2/Ee6wpjtqAHEp9BC4
I3zehe1dMALSKjoCqqccJvXsM2F1pQqasJqGyCkpdX5blykppA2cl7ohG7tGD3nHPa5tt2rYEq0t
Sr7zAS2puKAEtkvliW0n+cXh9XEVamX52k96M6RsLE1QVLy3d2Gl13LQSVVrAGnJVUZ8LNRgWEZ9
698x8VLONHmEfaOEvwCoGhXxkGp68o9Avor4KLpjyCh9JFkpkPrK5CVUrQIQvPwtLczqrX0cQheM
0Dw+zVMZy047QIKnfJdnWbgABPNRg9P/KIaR4QVmpP1dqg8t9Hv4/p3SA08D/BX8f2+gAr2K0F4d
Fds2QOb+sVQKvYHHznjJHlew1ZZNCNQR+TMFrFOjA0H4Wyo5qbZDd7THD4fqMb8mmtpVhcip8UW/
ErpgTDetdQomt+8TXitvtE/zDDkXgiqjWOd1DtpgqEtVaoRf7TX9yvbqUZ/rkgg27fykcjhbR8+P
SWBI5efITccLbKhl1a2QA9vD48WQW3AvgXac20vfOiwsSDGIrhC3wRUnH/2wzhKak5u84IeZiWFA
6F/VXaA9RZX6HBxi9lsx97AvLLbce4IyJQE2TAZx3cJtlAyacelOBxuTpaSs6KQBJHUQ5iAnHuZK
4w8i0fMBejIb9lXZv2V6h30pG+X/I7UClGzRIzDIvkirRAGauAAo+bAb4nz9pUc2e5RpNStItQsA
wR0VrByj8DbFDOOUn0coz51mLhZ2zdKAWXxif+QQqzyTebYLKY9bC6tQMnfKeWWinZ05qwhHX/Ge
nCKNHpbeo8FSa6grkjn14oVqcCDaKe/2ZiHDAjO/6QsyZrXix4eQ/152ULBVFGFqB+ZOfoFdTJGl
quE6LjDHt6VHBsgtkSVMUV3jlUUQRxP4uEa89Q3ZTiXYycpWpEYTKXtBFhRiAvckbt5YAWUuEA11
Nalsei8OcWixeJSQkfmpCTJgIgDn+a+KbRi6lKDAkBFZT5QY/wdwy0GNC/x85dZsTwR7frzaWgtU
UdfdHvwQ/Sw74+mBeAaBQeg6IeD4qV7gwBjLOctbmhO5PJ9SH51vattxj1n4RozhG6TbrYWRqz2A
HFT/dQg/p5/ym/t8++a8+Liox8yFH0+ABwttHCsBTyL6+XNES+YwNhPrDqwhACgDbfU40EyK62Xz
i/DlJkPhGocVPFd1sgyiiuTHvSQd+tsxrU1tkFGH8uu/Jx4U3kk+hG+RL/YnkhIWcma2It6T+6xS
bTwv9MP1GW/Wk1WU40N1In82nQnWEFGE2reYXc5k9FUqRcCgBKlS7Di4ApTMZ3C9OXbsLn86MWll
PYJIp04fPpYt691QFTFgD4a/4a5A0KnNMeV/avl4oBMaD8DvjsuNgCgssPGQg6Pbcw/Vv5qFyMDY
KSLxMmEH1pcHZJafZGpc4Jdm4Qz+8WvedxYBUFAc1JfIvEzlo/DM6SiTd8K6v4Iv3UWRqv5IIxtg
ONQK5eFDdXzYqUrTYOhTnza/Ey4BdciN4T/wmuf1g6Hn9jGBxznm+Xvgr/3yxcX9RReEhPqdGOxw
V7Ub0IBy4KZ5KrBfHIbpub/0CYtHs7/RmIMsV6IeB0V5NyBKQPUhLSA9oiYRxrUyBLFC2hWJ0fQe
MD27MkqOCnrGD42Pq2gWz+2Xy503AjJadsvoDdUT5N5EAJC21GYv3zkn9bZz3+mSj0Jze8fLIM9a
mwGnFPF2vOCDgPesfZEs91e5PLNU86FenhjI4t+qgComaSExRl8JPdAwhrY8Gvf2aAusYV7vV1Lz
D24kUVPVOfD0bIXDcFBGuJDkOizeHFDHSXyRYtpQ1EFSqvHKCPai6ZNVicXdCApI4k5+vAh2hAS/
f3/3D8PXMckBIl+5Kc07a6YhQCKW6/XRVRPnsj+0N5pY3siZBI80BFmX4pV+dZrq9AQdcIgquJFP
xYlPuHM8qzH1EEGc3PBySz2ZfKCzQg4JLC10lMfzY8QpvVwtFgz1gq11lTvXoTIV1NObi09gRuPn
dn6KN/Kw6lCoDZeMNsCYqtqk1s5L9+Ya8lysZICXFaAflERbJYo5shmGrwlwtO8uXpmG12MeVxEF
8oCgeDqgncnJ1FR6MKowbX/gSlcS4sCcYXrKyQw4OhM4jafWrKssI8e95aRrKQt+H6dgyAvcCChu
cBj4FAD7cFfom4+p7Zp/CwLx23SE95p8JV4hm9dZmZDlx72Jw/Ppi+rE23G3zLbRdH7VsvexGGuR
BfRBefjyEp4HHQ3/l4l+aDlYEb5RE04y08umf0rvfN/ISDyovmiO4bNJnPN9wk7aSvMRcwwYdmhm
E2G55HjZMl6UAsIQ9bIdnu4T1oz7KsJZw8kXwYhQEL6vfKfsDwCOSmadao8iF//22CyYZNbCazqX
0JZdkevb1ELYp6llaB0oAdZ8uVuJG/MteCsiED0Jgt6wvk7NAkSlGwpYP5M8yIvPKHz223GsumW9
Pv8VnV13jfVmCxvNJTX+pSCBguR7f/DuhwE2LoFWs7UZgVvuMyv72oVNgDv/pRYYDQt/fd1Lp3IF
ccB/PT5mMvGfAuPlrufvTtru+eO7GOYBfds1Nar0+38x+fqVyyOLXPSgd8780Tohb9CXh7ukwkm+
dRrhyiBRjrF0uB/bXR1zg6/HAA5H3+MzBUlDI5QWVG/PJicbVwyLyID5s+2ERBD+PxcqReEBgo+r
K4mtDPmDxZfjk5c8Iu87WyQO2Os1cR0V2YdRD3E0EOUwU1PTy7PF22C7I0p5gjsjA2CYAS7eHYMs
8svUPJXLi57WymSbxQJPXJNV8aQIRYFZCNNKRnOoj7exJSr/gF25KtFIO5hDehPOMhFZEfRLyxYg
O3iVadnCEQw2MYb4mmJe+h3BAXTVS0fKwYZxUg5rVBphz5yv6PrPQNRVZ/tTnp4qII8xWLOlMPMP
kt8td4fURSCTgWXMHLlnHfRlBHcHw3FDduaTzpdn6zeQAmpqfUZA81E0wNiprP7XHmfVe338YTOJ
gJuctLAEm8iliRBJFlb8UN9up+WCrscuHAhx902bXTCEE77sR5SnX22TQFVp1gT6AlC46+h6+Nld
mfgcATZ5aOHUcveLXSneJSSbdRPEga2w9ii5WZ4R7Jn6FV4f1SO3rIecMVSFNxX5vrrqN1dHl4Or
G6Q03CV2uZWqUq9pDBLxR5GshBBYieoV5e7ImsHpyRlxv0KU7sa8yc5vq3Nmahxc75aRViNH1X9K
FIvpLQcg0TLprIqUq/kysuG2uVrcIuScVHiQcV1LzRLttcYmMJ/SWS24m2tiUmRwYoXKT84qj2O7
gU/h/A16X+N4AfaYlCr7TqM2YNIU0EVoJ2PKl/nOiRvVny7DziwVcNU3YWsx4Q4y+7ck8aIlr/X4
RDce0zM211bwEnZh0hJDSJT1Jrd0WlwJGMVpXnMYYmcvimQ/Cz3xM3x+6vSjX5OZQC4say4kBRz9
0rtl5nCFbHwU9v03PYe/cBwkXsCOmTp2TKClXHz68suy541qVSRyRjZ7w1ECkiY42fyTd3PfymNB
TiiGfdxNpN6uxf+z3hoSNYCNNh6QzrehJtH7mMG7C1djPJX9KtyQK9ePnwNaXmRG6WLB7jJucUhf
KKHhg1GJSBQcV4lcmFYuPD67N6b6LelnhtUdgwPNY0A3c29UQknHn2WXqE2Pk4c8hRuCmrPm1TNf
bHEyqGBvH2ANN6QA10jrvfDk8Ac6i1lS0nyNYUkWb53DSedtrX3lg7gOtxaotKs86tLp3Cz2asqL
LqyEokHaaYOq6ksz4WalytxOHrTV55d2jkdw6O1IcG7omqO0VuRF+UniinzvCjdvODGvnhAgVOwB
yZDlVGjoz5J8sqjvuNwdMovWjIyuW0rs/3mxPrsoXRVgHwGDsBXA8OHm2/0IzigUWGAa2RAAUKog
EnKk+3QWdlHPwLcVERCyR48kuntzujdPi1OP/UYD3MmbFkPxQsqvRonJOtBxhS6u2xcp3GkeUyRx
u/4PWxGVzhj41HtEeqyYSDD/geUwTnspQx2p5a1z/WZkC0Bnx5sNKgxa0/wRjvgij7wrVRRppmkV
ZP48mlGn5GH7NgeT/yDXAkwslwUzjQUp8yPDNat4pk84ugvB9I72DoPEDv02aBX/gSONMon50w1M
yrjuVD9H8us4LKr8QLl+klVOy3FK4G2IyhSXOXxLzOs3SJtSfwOMrjrm566OT13VVtHVlNC3l606
P95cUcb34KjUvpXRrpJXcIyRuPlr7JYgCKevlRUxlbs45YsSX3J9LTqhgM8nU4gAO962JwsK6hQD
d+n//RIcZ/QPiSGbyGssV+V47v4coZROnnxcnk/PE9n//1s7vhfO5qmLgEUv3OthTZYTlYfZMaL5
8Ye8pGcc9J7c6140A6vbYLewGiGXG7vo5o7aPP4tUwXPN4t+obVXN2EMP4WhoA55nuLog0TZelhq
CirD8JpJ3P9Hrx1i0ZzUOiQSVzVhIrtfgurf/BBy7X1RLip1aKt94Skx6NuA4pE6iTjFaQCG4iyq
r1NltezXzJrvq8SvaEv1KYRRiDarWuKhs4DAHiqssXFLwZEwS/KZdZqhmeotJhAXc/hZnxwVT+Xf
kOyYgOuyjZNME8nOs4Boo7uZmyla8GHoyQjI1Q4J/uu7NN40Ff0Vnqt71ovpnEo7U7cnFI53+YV5
WwNHuuxNvFCdjvIvXPNUso1Ll6YsnfEMKO6Uh2OJoLbmyVGX1Wrm93WCMdMp6kue1I72T8cBndGe
QQ0+4EPrgB46YdrvCK05FKS+jt8KCsrtmzWRy9NFGsoPBO97KBqXIx5sQHB+9dC370R509+NRItR
GPddFp3xvYSOzP4Q6Obp7b7fcegXdlH87IEo9gzpnSsVpdZCyIwf3BCpiWCgi0FUJN7+NujO215S
ZBBPaf6j5TtFz3L9zFqY0R97w4AX5P3ouoE8Cb/5xCDmSvgKNhpG2EB3q+IDFN2KUTgmFXjcTNi4
+hnyBMJAsVSCeOtsht80mxOyMu70CnnEYmg78M7hDvUNfNdchro6lcgzwMUGJkGNecIUC/zYRo72
+cyDtPwRsqG3glwAbCDp1aiCOTqo4rMUO0E1ETy5Wx/1hp2EF0P/hdSP1QjDysviCPp0KCnHeBVs
tYr11v90/4kZXKPFnpbOWiBiUSggCrOFpu1RKKrYTvg+AOVu1/646bA7H7X6/uU8CdJXDGJxqp4a
0mAD32zU0QwzxSrWQD2vxshak32S0p51ADXeXcgwoVZOTGVi3cFQnI0tFEr23MYEs0vuOh6+0CMF
Uz4rTC16H9fPaq2EberPhuRquyZwULq6+CjzdmI98lVEwLY/hF5d7GIi9SnqLAiihk3Gro1kQ/WW
CG6Cp2/cD75SpjWKHJWc4wY4lLDWN6gIbt8ZKeOQOEzELczdSxygKatNJ+45fyXu3L3EAL3jj5B5
FzqXEY4OCjgFdzCogkYPxkFrgSf3OyzYJao3UJtCYIGLykSdtYGR2eOoz/N+aEhwfQDA7rOSArj6
rlaIWkhbpuiLNWlbpJmbrBb7ezt9acQQS715Jqb4pkZssdUUV2MQYKQBWFt6kQp7TLGxl71gzkbF
y+dhbhI9rVJNpnaFYofVYsoNP//aWdKvFhNxck0AlOaLMp/gQD254m2F8CQh5ZaCFqG/0r1NjB/U
YVkjsmd54KWYmVqYekS1y0LwFbEzvMW9+Cq2MShTYuPO51yIRr9xcVtkTi0TPxeVLFCHOhXmRxYn
JJLkM4raF+dIlEKea0WBluQ45Zf0cRdHqpNYJ4mXYrp7VQ+s/dUWBy2GtUlnL0LmdMt19o+axOPM
uZjflhNHkyoR8cBn/CaqHofr1/RcmVlIy+PxvwVV2N6LHX0l7NaAiehEYPdppnRoDz1rJdeXbGwY
K3WNm7ytxtsQ6kfqOG9Ha4V0g00xaTr/jMSRIkLs5zdVS6jpcLPAhdW2JWpJYiZKRecylg1U0jCP
BUHtRL7OQImb9H+0WR081FaDkrx5pb9KsfnoMlmPLvgbzyNFHt9M1pbv0iNWqNJNVqw4Vq8ugbeh
Fx5RS+dY+Q8aTZh3snUIojRwMKtMvcJHuUB1mnxz6ANw9a6S7cefLQJ36YI9zMhKbP6i8kaTc63T
nmSYcYScsuitSGz6N9lmCLcIy2uGNVs0U0VlJ74VeM8x+ONBJO9BDS+3H2WDaO7bh+pG2fJCoxzG
ThazPjstlewZ2LD78gfgvwAKpCSN8PMsliw47R7yQYRYX0stZHbmToT6Ed6zujC816p8cyM+J5Oy
LVSNgKVa0d7T3fZ+hQBvvA1HaeBdM8TWf7vGbsFPNgUCiA/zE4/ImEDfZTVnAGIhc19L5dFlEYqm
iKbuRMQat6Aal18+mRl2sOVHwYhqjHDsnh3rqftDvq42X9ACYXuRDqvw7IfS1f7Pemi4cKfCIdE1
+7qvTr/mkuD0v9d7XJnw2fWgVP5AzwrajPWfbd60/fNr2+Ozo98WhZ2l+AVcIpMmnFtR/Rgw88jq
imhm2c+UDTstPqcSrv7Wu1FE5wWOkEWNf/e/PXMYmpix6v/2AKJuNLuP6Q4LEGHmBwUgqR/pH9Uy
LLVmfgmWWR+tizd+R5nxInRjiTwWV5C+qxbimmDEAVqQyX5b8dmRZpU+0rgQK6v4jXfKtAwW4Pte
e5T0rEocofSOfbBAVP4EkfqTtr7odHbm3vCm1di71GW1lOnWcIPIKMi2zoEJz0S7DebHoryYi3u/
XNTA17P0dOm6ZUzQ4mwrq7P8vKO6VOgTvHXGirl6w7DhBBcF/xG9p5aGum7vYJY3TRs4gc2yiQWF
2ncp80ce8Xdvw5IJpEsujDaAvKLya0cFCEzErFCzU5Q3RBfedeFViHdjGhaxxHQbCLBXUNnUgdLt
yrh3X6jYdPHHCbS1S6lawpe9NkPcWj3AKIwLSxkt7KDRL0zf8KLJwdwFac2Gd1IkRLXK4zqbM84L
RGU50Nksjc4WDVVW2kehXbf5NlD8VtktF7+CiW7dHLycndsRGd++TgthygM9uSxmIizuO42iRMy8
D9axUR7ajTGcgmi7tiWG6wxk3UiQx9xzN9lhS9T0Hu8NI0GEDaiys4rfD3t2ROiXxBOy7/sxQlpK
jcPQhY27yR39ghviiwByAw1H6olDngkI1RZ3RqVwJrUMT0xseLBPobN3fNXna+16oqH0v+t87N1u
4eozcPB7CkueDkKqFXC18TrBkT1geNlrv0b+jB0G9lSVe8Q+q0DR9FHGA2hr4eRsBtaLbB+LWQfW
qCTgIDBfSB/PgHQOts9+jc8CSUQslVc3UL2KSXrTDvlJCEpYfFNGDGWc4XGjkgV/VLjmOqqlmGkx
L8oKmvzgFIzOnOgOIFMBgXWKMevXcLcwANC70yrz1VVCqtXPqftb6SD6F4CxoZGm5L3hjpnJqfvK
1PE7QrWs3Be8XWI5hPkUG7CcwCpPsJiRYaqhLuU3NtO2VC+MzARIQiOzVo3pn0mXP5SghcAhVBpG
Wgf6cjqbvJWG4ABTAt9n0d3xuKFdTazd0O1XfLzveVM6QhDJ5y+kmqij6YlVIZ7j57rNLz/w0Mar
erFnzLUDTU3RQdVaPj5xjQ04Ww1YX7dWPOh0quQkf+gg9gnSiqGBkjniowY40Zb/hitdXfo8eEum
lt+D0ocoStMTNvhrj3MqPzxxeC3bvwqWfnKiqPldFjrE17GOCggEmu30pG3UGp5uijpBbk9ppR5E
JBMLMewa1501jic+x2JIUpozxUWVRo1/MuYf5l7BbLGnA6f1nGzXYqh9++kze7oREjQ5FvKVnUM9
aRRlQmXgq0/gUyqJsFLCg8NSy3QsMnM9aVZanFCHlueRtKIq9U92nYC/cv7JQroaPobMi6rnwiGx
Wo/yLX4ofAu+Z9GXPCrzEmqa8kiJrxHCoqt7eK4S+Ap44zS4djGeCKtW4wD+EVIvLlzG/6XdFAQN
jy32ju+bgi5Uh+1XEU8O51BbazHYPA/Dqk61OjWZFC5HPa56omGOPr6HNEIUD0ERXJ7vNvLVzKjR
VzHd9sp/yBGaBgFS74wExd4cpJC3Nf8OxgjGHxp/5XUxFPI2uF841DWV7QZjh1+3KEWqnBj3vsqp
pXAklwrQxIqvSC64Wbp7lnyANTqEJqi0d8uCxzi1oOG+UWHWkI6l9hs76zPgBbwoYB7Ncx/nmSrW
kLoRCHwWsEhczIr5nbLrgZFcW9nPPYRYnqu16agL5bCjBq05pogA1OwN+muJh7ytT0eRObEtMgkW
+UuucyyKElOP5HWAq/YGmZTMTUQCMFPejbvkHE9gfVHQoOJuB5e+g8pxh3zYtOJn6P0KGWrOKvxd
rctyARbXOEMeYhQW0mt0Q2G6cYAzLUzR7fE5mIgFoJyAkJh7CFF/LxfdOhUteeJtS22nygH3zAm7
J89L/ms71iw6mm+ToSBjR98Uzl4LTmC87Pfqm8fCiCbnc7vF6VDk9NcrJxrEIEZqJsvY7JF6HlOv
1wqDFqYKzbQQ1vJQbN+Dxj5x7ufHFggIV5aGDKRKwkxJP7ogZFPGiFCmqBeRVewkXTnam35PbcCQ
2c8XDFzwA6X/11lUJG28vVyNQZVduGI51zY2HU/bMlQ3Qu7cQkPDOecgs14fNqC9nJLWhxpB/eGM
k/Ye5R/3C5D2lWJivmK/ZqsZVRmGwZFHlekgWAPvcWDd1frSumTaT6v8/asx7aYM5ExhmsWSZJ6x
gb+0C5wTNos9BhBLfOirY8Vbx7si6HC9bdueE2ZWF9YBXtX81wrTSAP0/pAnwfSuIj1KWbVuGYwn
LsgOIMLuKcpFrQQM8FK3XOlmL76wyIFaVXMVldDQWxVU7et3x8rbhY21Y4SboajONd8X99Qlpap2
SoZItTUucI8840/WGsC8PQ4Mh9Rx4x/DmlcbpdCm3hNcPVCrP/cuzcJ8klYKMpCWhc7F5mS+nZtT
XAa9lzcYf/7iSLmdN+qaBD/2OfiY7zXfIJ0RlJO8iwyT4300yfAl6oCh+e1jrFlAkPMMuXSkofm+
2KmGBCz7/s6RJR19YgTkAgHkoag8X71mfrskNSYXYsWv/OxFXNpDFJzo3cDrcWyj9KYRKDyBV1p5
48cgUmULZO791xruCuBc1kDISdgrkrr3ASjTJ6t5Z4CEOhwPEOBXEwZUVyDcWoJgcT8vBV1M3NDR
LHxX2mN4CMMT0QvMwbKSTWyZSWmfKbJscRI6A5jHIR0aNX8CLdt/T8SiguTxT3QrNeYW6t8meJry
S5Q8jsejlGUjQE0iCFWxNjLSDbagpiPHWWU1ARLirFxRh0wyEqWq94d3/HhX4DjMTGS9TkPguK9Y
dCbf1u9GQ9zqFy68tVFQzNjPwpNrDH+luD4CXw/IO+TpBla1vR9XTxxm9voSiT10KtIbBvKBbQxg
QJfh1UAOT/4o3O3AH+sbrswwWdsQMXzzGNbHPXHCeWK//hsaWBrGfJIJWy8VlSfOim6eKPQbo1aa
4hAiENCLHOCawxK5rsM5Y7hPvKMOnKHi3PGED88E9/idTUCNPmI6imlp++IFSVyGavVpt67XZx3L
NISqNAse/ekk25nBbpvAaucO2SWcWgqvKlv4l8E+w9hmYhN/dTMXyjxqq2F8xlVfScZUkzVrGWdF
wDvBGEM8MnZBWhxBbphFS5dctErYHmCTOFhGCvk3WRrdmXxSXRQxCxeeTMQ61H4Bv/p+5BVyiS/M
vvtmcd7CTS1Gt3THYzcbykdF86oyofV1khcn6AInMMSzvZeuyN3+XVa3+1DwipdQg1sRTktrlNOc
3Lo/W5k43MmwkHcaZ9tSlG+u+vn5zZFGBPkwm9AOYBDJP0eqDjhRoEDdSLSkI6a7te3OSCt+njw6
8/DPWqNjeIeO+U+uZ6P6OBPEOX2TZKXjxKDMI1UT9la7pkrpj5B90tlG6EskLI2HjM1IU2nyfVTR
a8JliL8go7AmptyHVb7DFZqrrZsqPVC1/OT71q+quWnV0RE+mQj0FBaI4jSJX2yaF+hNBFHWr/g5
sns6P5W9sUOHyG2tHgwXhWDOvGfAezLE0AI9yGBdBVdcnMkNeI75XK0/s1Z42NyAdWh7qopDV35R
vp+Pj06tSMkGnK89msUVK2wddnUpQCeJijtvW0GsZ8eTm3ZmmtpbgjFG/Xlk9Lmnc30KfbIlIzZo
A54ALuYtvDO8pn9c4pFWRelwg7F0lEVCDO7FV431aXa8UQnB0rsDsNLsj/zonKzT0rchYqI+dDPD
OH3HyqoVEkgWtjGRh8FZX3Vmu8Auq2dWYT68On5Cxr7R6ewrHxZX1ofE//cDJFm94CXhdMffZ8xI
sYT3H/mWuGmv6lrzBXOUFTJ2opNeYMKIy/UqUQKGTnbXe3sVM4u71GKgTP6yrWvICzSRao2VTv3O
sWnTTQTNfOC5zCUKKk2nnPE4FKpHD7ywymtOXZkEui2bU65nY1SzuTL2zvI32fCaacC7yA6KkWzs
j2WzCFRCrehHhplFdnJVOI69gTKD7aCW+y1UBZtPuIe9i9KD+SzIxGFGpllW8K4hMeYuzqh1KdpK
0I88IQ83R427FQkYJY4vYcIr4suoCPQCrfEk7id0CldW58r6+7uAcBxiQfIcqGxTPGX77F59wm88
Iy1r7ibaHnKrxbew6jWgdKiR10TJmGe92EPsGFxNxjWVpO888CRfdgaWVI+r9Vdjah/5bcdaU/k/
dILP4YYfDsqsWm1rwyhcFfjR7U1VyXclnI5/aWEH3KDxc0yCBh2vS9o1CC4Lgw7m8vPSdurfxe8A
zS6+VA/7OaFTugT8iV8xew4IqzocCfq1a8mSIvxgRlWN57iOe6wApuh2inbtjGKWcD3YLkQ9sak2
YH/HXizAQESvpK2wzsJzMsYEMqD2s4MosyOK/ExwEJg1dnoEeTMeFADQt3CLK6MmNuzyoh5mklDe
mSfjrDgpafuDq2oXSiIX1fYKimqkz2gcEG8nUnGM6R/5nSKhOyinv37gW/7VqpPzx1zC4Y4Tq5v5
C3l2gLtsBRp3sM70MrmaV5wSQWfWpDQVCkwmV6Ho0vOOoglD4cqnmScyB7pqLwndlo3+3TbDseq6
A+IGvcg+kFPSzAxTMXarE4mowMFgkIZ6sjczFEa1vHWCX7+HYebEqQfcskXP429gHhGHl/2kA99a
ciIjks1byIVckwn5iB97BHbRjUUqM40Rke8Q5qnT5wf8GQ5EoZ5MsiohmXbeg72Vw8GZrveAAGk2
/26dzsH5CRflL/bqlUdDonhsfak6OvhLEbkHDRZacbR5ldZflvZfbovqahSE2bNYklzLUfKfHRwI
ISXSLJUT4vTcQQmxnsE9lL7btbXKl2BTvPKzDkyCKGrJZXMu7GI2LwXvtiZocUpney/S3MgVAjXd
S+QhM+JTflWdDyRx2oofu/8BvPxAbHmxyttaAiumw7HgpIEMGdtm4ybJ2Tlsu1XteVvTYk0KRO8O
8r8FDmK3An6qClRH7SxICJMY+cnjPFGKqaE6VhblwFXvB9vYMbq8BQt+/j1Dp2Y8eSvqoQdjLx5k
26UljN4jpQZD6/TX2Vrbw68Um3ZU7WmglF7EgEm1HjE+7A94KMLxVKoOD9d5Q+7M5MuersopMNOz
8iIDbQWkQmQz72H2utjEVOUtlacsEha9MZ35cmA494/CHttXk84omLfVdNStQD9ydKB6povTo46V
jS7sFUCMfyxOw8S4YBkp5c9d9/YL0rrCcxORNMbq0sssC4iaJS/1+RoTshvpxp1Yt+zMM/6sIja2
wlxrRV2jWs6JmlcdAjB6tcGStuQPpLZJw4OOQHB8lC5tAlJReU966Zhpr0P6ZNftJ/1wrfe20tJ1
USyfVtX7HFDqJ6PXKlnbuxv4F8qqTTWYz+FPbLv6gZYri8gz8gdYNWUGjF5M9PkofVgEpsTXGnW0
baJAQMEoRDXgiBJU9irnZ99yu1GEPCDmvB4dr9gV+LayOIfnWkKON+cD6HyPH7g5UHfAWvRA3Pdx
iumXl674pYtq5FYjTKEqH0x3QrgzV598vupmtw+1SbAd8jdOCqSpemGkCW6zgXasPsuKjcKmTEha
t3bhrEp0bOWs2Kshm0e4fncE7PMqUUq4w3LHEqcvfJzeX66Vjg93yIZHag0wrSytqPcn/ZDka97D
UaU3eb1ZROiHSNXjXSU6OqBxB2qTr2pz9nM0GSvG1ZSUxB/rtYvKebJM9LMoKqDNXtoLuFp37LGt
0OnGlS87arfhnhzrCZjz3MXTohUetWRvOw0g4zewCbsQOkWMBUYnAagycF4jnL6iL9KH7qCuGakx
DxiBTcRL1dnMXnMepsCPDHBVgo6qJxPGW+DLbPAkDN+5bKPIzmIiKpQuLR//Ij5at5k2mDBRfEv7
18w7PxYbUhKkJ6sCuEMDywncsuCVCVocQh+92Fm+5C3qamfz9srS9Ab91enqFl3hoI5WdD+nNOno
QyJDA/36yD8N0Wv6bBlTtlyjtS3x9MZ/Ci2ujB7fXGtfylrMtNo+d2URMBlEft8sPCaXwTTu8DTn
MzvALDQTO4q8IXA2mvlhrob9cCIv5Yz/CGOHELPndYdhQrmFwdtMEvJwLMA5lXx6Iy/3BGXYRYUP
zcDj/6OSo3mfzGlieCNly+35z5WFqpcNLMMyudNKaw9RYiX6PWrw2sylDjzDPjsJ7Gtcs4+KTmXj
4aY7Bl5QXJ8DdWv1eEkec1JkusG1xrYgtZCmVqsyo18z7c/EA0gawedCavPQ2kD8HNqZum8GT4fX
lSdqFvCSTu2cWBTRCXVSScjTSorg+1PaDKqORLC/winIX8sakNvUeqCtI2iR/rrAsK89TbzdbUBG
4z12LMtSOLEOsOeZJRxgk3bm8a6yTFKb2gc26s3VlWhIPnlabn9uM3mE7WeErzb38rvneVICWNbU
9FfZy6Ha0YD/JQyhFnrYpj+tPp0idRwvsnVMoA2ZBEhEEMfSaELTjdN18v6k1h/ZBsVam86DuOhr
ADl+6x1XY7HLf4tCl/JN/Ty8J1VwLf+vqMC2yogueK7UDhlUypcrHyRs/puONcxU2WFGYuJ5fhRx
DRQOYFunhmcRK8VXiq7zcs+m1nAnjlZ5ataNzjC/68LxgAq1mRoSAYv9/W6/9JNBiFx+Xu5W/6Z1
bGUgLxxARN4uRajxiUqd9En1+oK6fC+uf2WoaAod+zIlMmAYRD4Rso/ogANPsb4HO5NHx751E+VX
bJ/UO9ABDcYIXEQz6yPvfycRhCSPp8dceiS8nuGYEfh7UVHjQkWTr2+HDEEmnOgUxLCChuedf839
lgL91k93yw5OSKu8Rnf2m2i+DbPOi1+uZKmkyXu/8ILpDkVyY39VmrjXgoDUkD9ntAI49aGC7yxN
xWLYN3a+fOCGzQ2R+AydwYQH9+/MO+2kQTSPGiZmewTBL1JlszAFF/ZWTqf3Teip7ZBoJxz7LjP5
Em4a8lHZ9YkkwrAZL0LrUJt1AscuFrN+tOYxzXETx3Fx6FxftohLanxcW/GmpRaYtNsX+MYLLVrH
0nihjtNSq7ISExW3nYZC1ZQdfd+3EtPJjxoyQnjOWKzJTX9qRR0PBEDjJEM2DW2lhSnGI/g1a4au
7qPo/kHB47oN9eh8lf3b5Y6UtYLyW+iMv9LQMLJj4P9Q8jSZ5qowOyHEjIfeS4p+qWl6uiosLG8U
CZhlE/XPQWnT2QhTZ6cVy1vDE6g+uc+4kIAc+ZI3iaYcHdZ9YNRKqpIUgFrVGWse6AQUHw/Dp43H
EQX7RDWX061gis5sG/TRAWSk9nLtYBcBNLQgl2747gUYt1B1DLOdQhwOnHXQirJBdsYanDKgh1cF
/atwFEKEd7chJMJPIxWrlMRnMjOV5Qo0rmvZsRc9A+KtXhwCFsNF3KuR6OzZTpmrX6oG0/W0qEK7
5Ndm8LNOTUKjD586YLqF+Fwo1xFid3R3dnMT0FeG9qNCXOWeCgI3QLc5uwRfpLExxIxGTnaOPU+w
LZiCeElcrvMhKD7i+Dj4X3j/GwQWIr7Wo5784wHozhKfzquph903nwi8vPWmwHi97jl/OVLfdRwE
sVI5KuACBK9iOA/7bsQTdF400BuzUsPYqOVRDB9iMwMEHNWEOlDvm2aBT2qN2Kbjy3XTRoH9+O66
Y4oOFpCHFZMxIjVfixnbLDzpJsVILURIxqfq48JtBoLEtv64MabOfNStvEQPUldsIjeQczbrbbvt
jhKZtmnyzMAuzAVBHNtNlxA4AnJg6lJoGhR5scCsZm2S6AtN/a7lmcTwqlJ8pTTvggQmGfG9KL8y
6bF0eqvKEEtlEPcdhHAjshR7gqNlZCOoVHT6bcCakqEb0RlCMPxu8XJ1oi9QZN79BAUrm1ZQw4if
oZEaew+CnR/gZA7aN6GqmP3k6RPj6zw3phgE7FYYyYDa+rwogZOZSch0rBW/WknUVnzl8Ru1unUK
UD3eY7wwfkChGmR7NSVpEUXX50mBo1IW/mCRrWl9uQu/W/Go4ZpbcWk32U1n+ctabF2OO+F2mYSO
dL6Y4f23QBRqIxx2cI5tpox1gFs97VcVtN61ek9WMHJTTQetgmplO1geMWL2XQBF1zid/fQhu4Qw
FG2fqRAfK63j05Cx3cKSlI92xl+PwziCYgut22pLpI7PsM8LdvMoO7PwkaticJBrz5MlM/ecjTD3
k6cJyMjL4+nTAn4m/eIBPJlMb3vftqrCSpS9j/qfwxrao89UlZWjMbNKYBPWflXOQ8dHodMKGo3E
E9eolVp9fXb4H6nNYT1HdtBLm1uSVGJ6uXeQQEkAIGAer26xOxoiyzMKKzoUFTdcNf+ZgO/L+0Oq
hV3S0fAoROBNKsRuR95l0DotakUB7C7f2yBmUEbmbA1ggsorhWmI0nGlZgCDJFavr/lumi16DZMm
MyhuNbM52bxvD2s9c+5p8ohWyk//z9CpE0QhJ+E8xdIXIUdodbyrpjQ/fmEuZB15zlz/FVgFS7TO
IoG2m8Pnw4jxwEf/nJOu2q4jL7LSl+hFHj6RyYXCld//v0f6hifgmWdsrGcbtvojyO7bSlme1tyg
BBT1JwjWw+4mhbUSQRBhtpJJ8hYB2D1a2AFUAyMG6VIUa/X9W++Mn53IsvpCM1/IUebcOoTlMZXX
2jp0muiY3GCHwRRId10fy9aHTS5XFPuhK7icdQ5ESMuJuqnofuTwd6y6Dm++2yIpe/1HJ6aBpx8E
oPpRWcUhwp5TaMukFlWYmlzRSTxe7lp6pPQUH9prTfTsV+RUnhnJiOIj07PeTX2yahpyQJYfxv6M
qPRKoueDqWFzD3B/mSj//Mxk6/S3ewJ9kZ2+3Ig4iUAfOluzDzrRXmcq0ShYKiBfLhIpMpdg+qXa
aj/rT3XoFnBRwqoZvsYLC8S/WIE83SeYJ8XlPrazdX658dfezedYyRtdBKGHZcNVhzhdhnznQkFc
lcOHUoEKlinyvjjpWZxF7LMqz6pcf97mmwwk6gL6dkPOo13EvBN55v6BPNyJGYNdINOKca63GQeF
F1NTekPx1uc67rSO8b9kA/LPSTMm15xD7mgx8v7uEO5PDkkSp1/rfjrQe9dVfH06WByHHEXPYzN9
YPPcSkNSAsRvuXUQa4VzNsLU5E4YWubN0lStI2SM6tvxB5R32xbyFSlWt7nY6jDExSVh+oCd3zkm
0togmsPpnGu6XI3QDE1l2magkbMHPMJy7Qo4BqN/8CVipMOadJuNiH2SqEYSgEsaNCvadbn83WJD
QIWVqGVla6lJBYvIWrbmckKuOHbfBRNNDCOg1DVLxWL30y3m9QDF5N5d9rltjBOKliKjDygRk+Hr
O9Hwv9/YoGfb4xe39oPm+UEwKHhXh9f8h3lfPOv81rW5a3nRiccPx51ZLHT9hLQe3G5KYTokGqk2
wxZxb6WQXgfJwhio9Cklat0GJTXin3Vuqxc0Leh4erhPwWuzrqhmQGDAHZ/9M9viRCyHwCTWm/tV
6onEB5BvMSODGD5odSGetHZeUxkW70mrzrGt4IM+EbqxFNt+ejDwpYrHj3uRqtDi9MiQs9kc9KI8
+uG5K9vT+VD/8UUMHvVRnusAHvuko8lufmtWsQ5ryjuAFmHJsQVNRNdWMWLNjaHh231x5NjcySvt
Ruf0LmU+/oZGdSN1UZPFqqpQQKgXjdJ23NRzhcgLhXICshp13uELnw2/xN8RT2dJXGRhzPT9jqbg
KciqGa7+SvmWW7/IDQBBsxacJq1lqsu6ewIc6wrKz161sIqJ0m1h56v6ytCMqSi1SDGMoDqLxlWL
u4aaj76DqI48/iGjUeH+hPqyR5GpvO8v2vSBZNGYPm39aBBsqjoTTGsyJbl4znLDIKaHEQ6wXh5o
iMm6Nf4CpTRof7KaaGjHR60GjkEKVSLvON2a+NK5e6wRhPSUaFEuC6cY88DrrLbPwqGhDFh05GDp
t2TLZ2pXYuoVe0C4GuuqYLNZUhe4G+GzmQcL1tvfWphCXrGU89PsS9koaOZzsDxwO3r/d39Vdcyk
Y7BNlAVKDNdw8zxJrDsvCDls6OnioqMLmnD7oFPHN5p7pgpjLDvLaDrv25E8lAIyKCobT+Aq4KCB
CEQLCcx3zr7u5QVRi7SOALT3atQQhvqR+bRHpTdYwEj8KuhdnCiFvsEkZwpvwLWXTyiNwqADVpn9
OA93ngN6eFKb0qkh6lueekFJGF4e0Qd9rLCQoBuKNY0zhhS/rqvTa1Gl6hhlefVwdP8JTnYe/1hg
YaHRE/hHBOpYBnNFWyVVwfrWiW1X9O6EGX+XTlXec0tE5VU6iafw934HurAr3SMxUT0O1iAXJ4nB
qMGsQc2pRvPAR0PC+ZNZ56YKTeIbx94NxNBBOmli4ajfv93HuzDdM2cYwRFfrXXOo/xkzDbdhZqE
cwIHHbPopph5JjAXer5Mlg9DhZOm99A/oikf98XgCZ6RTUSTzYr6HyPRbYz+XhOCin3cXU8ZCARK
h7DodV2AJgrB00pucIerZbwcGFVucedNG+tgNs/5tjAerd+QvyXQfFdv/ZVNxweAGmb6GKwjKqI6
u8sx1chF0wss4Lx0t07CGquw3ipo+NSeh9sx7ney5EmsjvcP4jZwG3HzuLwoWWMbQwVaN0txepcu
kgEBRzAFBheMVWhWDmWB368oHgy7ym3/x5GioQFPOwFzbBedlzQj/wpmqO1N1+5k+Jq7der6tE4+
ojcYd1uuWWRiPYwSVfcYmx2y2uVIf+22ephQEVL3gxjgWdl10W/4293zN0DrYxhn63ycxvsUoBP3
NXZOW+JLbQNz+YaByr+kQCQyH5FOL1HV1feMmAed8JQdBzU3zHBaO5udEzEpaZfiHk7dgwmjJKvZ
AJqewpA3UzFrH9u134NBn/q0Wt8j5I2MaLJxOP9U0lrtvCiTnmhfh1+Ykbk1hyKdoq0QnrQYvlGR
sjnDpxgmpJCsX8Mx9Wd99BATxVusSvHC6nSxL7vfZNgwgzAWFFuxrOnhlEyONbnEpaqva3nBQrwP
u7Df33xbzhiAQXRiEmmbSexgI+JJPU3KdNBTPLWIoSRnVVVo9g2Hf+ci+xY5pq+5YksynLZe82fp
X7f98F0GA2P4fexBuLndgIH7/RXyeE0xP2jZf4uNigBewBeIpkbwl3qtCy1HDLQTq+msLq/Ha2PK
ZQfVIsCF2fJ8SrMsVRFF0TKRXeKBiRULxR3s4YqTfHI9lfaGkVubWJBW4hgIvxHCmN9QI24rc6tS
a/PJzalcHUhOdOpTdXXrRhJF1XfiKEpcytxSocvPsXjAwCF8W4gfCJb+otQPcKGvoCnnzrn/UycW
8WvYzINrJ83JBSg7hoSGiPcmcv51l4BNN2ZUFm/MZQeckfDa2j8GDdh+eZy+Pa9qzqmpGaRbrIb1
ia9ZfCp8kXZjyUh8tnlhNN6qGgsiSWVHj/8eOLd/DG8u1MYGurcnP27dW7fj4M4eNFVb8KQaa1A+
3jsvXia7rE9NSFKejDJmWbaiVzLXx5ZvTnGQSHlrGlSdoSPAPJ+K1ggNZ3OiKrcEFDfUxM4A4Ad3
n9c6Crj5Wm20b+ezh8fzF0j3dDqFfQZw2IBXThg1/15XrmC/Hk8uz0nTGKNL/ql2xf+O9fku8LrL
JNGq2jUN7cRude6nqUgCrhS7wqJO8OePeWYZ4td+e1bICbEw4xotu+GMNfGjcGahC6sWWkMc7q8f
IrOek84o++s4KGf+s7XE5mhD9MldnHpKSW1EB1jbLlYySN1+lsYv5WBRstVaIp27edSHnt1nQ8kF
o/6tF4RmNou0PrC7ygJydF3A48WkQ2Eg2ft/446o+3zocw9mhpWqI+QJ9mCXollf+gs0qYyOFlIt
+hexht7Q1fYxpB9GCQJQQQUtsAx6YqB5Z5zDZmIjV4xfWZ42pR4WGDrugozmeduE0CyZ5MnMoAKI
kkTSpvuQEAXEvFACTYCA/bcMr907FBCqRMIx4KxaSg5n2dXEcxbWjmYnl/6cnC2oBk+6SSkSbXOx
SJE7mFnsrvXq/ff/qM6m9/IuZ7TCpzaAAG919735kJWiQIJQx98yqwEo6deNlZVqPuhv8brXbjTn
qqWi4WxNQbo1lVL2DjdJ/5zjdMNE5EdaOEg0j5AIuE6Y8OVEVLPnDbvPujM7+d+yBKZ2IVaW2AY5
pvYRv3Sv4H+Qu7K149P4o+p9Ns3DV8c8sZL9t2QxqKeVgUsELROvE0WXeDF901lN9WXCIxnSILHg
qjgsUqc71TpesczD8xjBn3S7jF3Z4Ma81Kb+tbxZdtvYFH24nhBHjnAW14CJ1jGPh2B/uuyg5QFI
pe9V+qkeq9p4NkgoO+1uchXvQIJvCH7CNcBijYNcopnVh/z14UzbFg6GvcaS7Ww7/R0uWOiItF25
ya/bZ1xSjzi614ee9RgCxk59ZBnZ1lWM7QRT/zEkD+O4/600TRSAAYJ43pSmzjnr83mLfGOengoN
2IiUmAAJlPt+yrMrIzDxsqjmsNYxHUQn9pwJv4dwCNttb2CGf3LGQICU8fEL2K7/1uOvMOxEaGtJ
gN0UqScuaH7nJhO6YOSnddKZKJ0OCC5tMeOlX0Hd720Eo5H/PoPVxWf01xyDdNDU5+ptV0bVu3RT
YVfPuasXTVOz2/klGMOmdWewgj3rikiZYQgEIIf2nRp7QF6HGbOk2aXTYXtsD2KeWcKleQ5EoXAB
vvsDRPUrn2h1zGdqVpjyWKN6TgBYrYv1otz+7YG0xoiFaCU26OrEWAFrmJ4DMsYyNm2jPXGwFzoz
eOXWC+owclRuhuub6CTZimcKUwu4kmLgRF2yLkcHMaEkijI1vP5DBU8xPQg1ECBUpR9aOl0p3MKo
VJk9oB2R2Jmz3zQWqTU5YvRiPS7hUKsBUbERSnZklnH+qqXUO+qHPqtvQOMD+FAdg0Nz4KgrNzlN
WBw22gUTw3bXq7oVFGi3j5K5nKWru48gtLOB4NhN4sIQwaknpqbDz8n2DnqZqjPEzdSSIEDFB8OL
1+czBvPABSnMGRam6HHcxGUO2pJOwksJnaGa4gxKQzr9nUS3L4zjyihMBUtqnctBmw8OLeI/y61x
NecvSQfuTpjzpIc0Mxup/Oqpmt5G1I4kIjElg9mnvRO0/uXLVQG1VIuvmV5pc3gfa8p/h1sJcYGk
FP13CQPUIli0gXZEoA14Iaax654m6c6doDk0R+BtCFqNOXvsuxaerkOwmMKgyVDJg3ZiNmjIMGy0
14yd/xfBZny0oYuIhcxonkgpcQDrCU+I/+xMUm5gn5iucs9OM4HfNRwtmGCjSKZKGXiafrhBIRll
65J08CwfHzjWv1bPqVTHIznf4+52cRXJBYNZx3yWXYf68hTproOwLNcmHorw4pWOx1C2cuBr2Lhf
oO0gBLNoYXanuEbHcD70EYSrhr8m5op/bOykD2pIjqyY0BZClXOuxG60drhYpMepKSc7EelvVcYU
faaXBfKg8ZrRN7yyLBCq1PeCFdQu6mtBlgfTe+F6Sau58r6Faih+C92PJQkIVBhXNLzAqKbjKdGM
O6is6ECUe0UCvlaxZ2Gc4YaLHguckX6LWNRBlb2WI9pYYaMUs1pDiROCjFUtNT8QLDzLW0b8PDTH
HLx/wLFY8EfuEHt3sMT4PMOjwxLXTqUdOl3oYJ+BO64w5v6m53j0GOWT56a6ltqU0vHo6Mlc2Zii
C0bslZngXC6HAgB5Yys5ZkXG3UItrDbd8ObgB/xB8curZcjIcD39tyjO5XfPJl8noBxZsffXC2oZ
ii1VkZELk0Wd0c6Dhjba7uwn0Wr867vOYuUeZC9UdZZRwcA/XAQgfYFsYjXwEvx0ANqORdfCtvTR
ujdTf5wBoblkycUTFllPdeVminPAEJKyIowyKp3ovUS2VMzqOwEeX2zPEVwseFYKM/P7k/mQdmAk
u2VSuKWFimO/b5NAHSKyBGLJ6lne7Af5A4iomWd5RWvtd9NsLqe86FcLEe82O6VOP8+7w8u74ylP
ak/umtVeT+lKsD5m3ffFPpE+G0zQe22yhIZKeC24holAnpuVUZaBPBO7S0N0xT//0u5Dgqq0gfkj
wbqskGBdn6Ku4nZC1vOn9f6Gz/ZBdaLeZdVrrmJ7Iek9rfwhaKDhnIkXY/3FUBXwXdXqyI8/nW4b
QofIK8NIHNPSUgj95chihI2gwoLH+QXFtKV2nIiUyQX+0epndAsfdgMGzWE9ph6A+OpAawPW/XVg
hixRirWAatThveWTDRlqIMZrF8yKiUwtP4cTWsNvM8Gm/+5XGrctlgPffzs95HhLJHlPhDd4GouA
KHpMN4DZvU5xm6B7UBbVQDjpXB3+mpvs1b9Em7h9tyaA1Zpt3p9SD6EgKRwF4gtw9bFC7r1MXGN2
H7PQFIu2pOLeeKMDCIvazpNfzCHdNsFaZrkkZSa8xuav4ldod92zXKS3aAcs8elFVP9wMJP7Dc25
W4WuJ9Nrbb6chmzDmryU0dVKk2ZWVZu/WGk5oizy8jtYW7YKyAKt3ZrjGq9cPI8xNTJR+ixfPsnE
TLMbfLHi/fjOlxGCf+ialV9N0a+2YpP++TKQvdJMWRk41OVYXwnqgX9PdB4+GeVCEKnputCWQsYA
cFGFy7ehWlwz99oHLppDj63YS42DhxCiX3q9SNVXSR+X65kiOnq+SezUtQyVjz5/9hZ/FZqadZLm
lzithvtxA6XmBc75ioyaGU6tEUuSUO3roKA23EDY697KTnJMim5RroL30Z83eTtdp6h22tWwk4B5
Xx/TjuYDetdvlSstAN4c60NpU42f73zRg0sCWx8KzVsXH1vc+zLkT468QmwSRWUSov8jh+Ra92RT
8PObVN/xWccZRtH4BnP659TNNIa1DWrDlrLmsdhJtDTcTEy1p2xaNcX7PIjwKykqKFrYO4qup3c8
QO6sk4sV8EJxL1wHXZz/CMvCCP5jDn6T5oIVUNBUQ3gbOjnXQ7WanDAWfJ8+MVwdAB6wMvlwjS1g
VPcHP9riw5KbfikfNt7x+/tdM34Obab1lRN80hE/MF/3WrlzugvXzdIG1T8Xz9OeQfSQ0L735+v6
yFomHKEdUWJF6Rqudt0LoHGTzPStjcHQqtltWSlSDWw+vLdWwYPDBqNolLARyd6WCCswyx/83Csr
MlVylUrtABCnBnCCIAX52H/IgqoL5uBXTgl/km2DsZaq9VzAt4d6FD60GZIHJeGKjJ9p0gWkq47X
EbY6ugKggliD2oE6ul6Qziif1uen9qL9HEK0Hy5lpAvEE56oTYJ5xNext1dso8dMyD3c8tq4JUv+
lthmr816EbMX+8YAMZJS89Mn9klBF77B3xaXPbLy85eGK1dw1QvWoGI8q0J7oG6c43M5kluszEgV
PGtc+fQgTGB1X8lYbMXcOp9+Z8eX7fH31HLSdiup1DOLQlNU7Fn5LTl/AE1HlFS32MknDwCDFg5G
tYDunYgfKRDOFhNX1ut7RBAlaQdhQrn1rKRLqEErS2P8vbMd6BERBzVHgE8D6XtGuKXRnRLXYoHd
f7XiqT/4lZizEQWU7ea1fxt73v+zQcTeTBZlWUl8wLDe4++uOilZyJHKS+EQtU30RLmxOfGW+F0U
1mcdtFFylhcLczXuzXXXPFe1H+MtrEWgTo+Y7A/7fIYBaOAjkKhw5vgah92LVgu57qRJetQyjTEJ
OWDQ6vrthFOz0v5qfL3N93YT1n1AydT7qm6uGQztEFNu2QHq5qQ/PbhThO1DPlO4svCUxKDVZ2OA
RwkcVMMNDSGGFkfpC0BGjkQ4N10rvxNiWpYIkRNXnmaL8XQYCl6xs8xkKJjAI5dUwjLv9gOxtO1L
e6Kt7kU45KUk3wEAr1zIDs1v2YUQQ3PNPOYjHLd/fbQlbXtGoQnUyDRgmgbQpqPElEs3bMtw0Fql
3nwJrC+HHOSW16jjThUwXdBdJSitST7ph6N+0lnJku25CHZwgvSsn3AUFBq84GFkrDnOqJz/j3C2
OyZh1Zg4VjEb4kiFYw9yurfe4LAbjgIsFNFyZ6vhNDKr4ySeixvAZMMDJ0xmE82FxP81F3EcHg8D
hFWfkErQLOus7Wj5BsjcFtvrvYayil0P6NVHU5m1XIMUM9/F3LybrfwP1xw91pELFl7wAFFHy66w
/fZTMTg8CRyeKP4u75QuTG4FHYWOqDsgzDe4lc7DkT8YxRxoaH+I/Tlart1HILNG2cdBwXjd1qQ8
0VdTyKVa2U47Alc3UR0wrSakmJrqTX5arNK0uD3rjespXIIOkpkt4HvkG+QTlVLsFQq/eLrGwomn
3Dr3pRnlJsiAxFSLndt7WrmHYvsJ+gnQQYvO/Yi9/7NGvof0DD93f+wxe2+Pai46R8itnkFKz5AF
pDbHteJzHHxJFYNY7cUfVo20bJPFd7yjfxqrhuuL3hhpe3KqJkTTTHyVgAjRME6KjpjJaBI/TaFe
uSYtLHQUVsN0h5Affe+HZHZFnMOeiGOV8RLaQK6qkeuinIG3yMPOKMYM08kYAgCzNNjQNzIP8SPo
OmymJaA94o/5Mgp3AGaGtg/XbiY10wH2VKF0/BaOLu8Vt6FVq3fV9Y66vafansiCKJCzDXrE28kI
GF5lgU0J27Y9Ykd16KuZkoWkaBmJkDpzVJmHJ11H+ftWezykI91zlkZUue/juAi1U87dLCwOXPeb
bf0/4E2KC3sNgJiIkVfYwAaHQg94gg+9jlcYT837OcrXtG16xnmAFWwMg5rEfuZ8mTOO7PinXakx
iwvEshaGVXQF6hOTwSQoyUrparCvWGYiW/yHfouWi5zqnoKFMXukmm8JXRguEV59v0fLcPuR9mLl
qZJK/rgDAPGn9iHcsSnfN2wUMCzg4QEIem0edlZRqOyvMR0mELExf0B5Ib3q/K+1te+gh9TtR9aY
yxERIo3JdrJJe4KCsH0jWWbv5PhKB1ZND01SLwS+LYNdlvX+pjZ6+lhmPDb7cUN9CtRYPhGgH9Fj
+2Oc8ldlOPFnvm8Io6e8sGDBjRvkgXVCFB4vIGVOoEU6SAH6D0+sjPd1nCZF0HBjJacSxPKOeCWh
pTB0RkhzG9le4yXoQ7XFPaKIGoCbVKFmHTC8HzJAAfJQ4n+JGcYDAQtTSo9r9UkVgCUKgE7xu7+a
HH68qpqc6eRaAUMfsLO4X95+0Rnw6Dq3EjnvQhs6ObmZtpCmBFfrwVjYM/xhNhQ5bhl/QwU/IA//
pwoattExVT/Il1ecYhccVTdcnJUHWRol64bDzCAD8W04vfntOtG8zRVhr0sO40QZX3YJFvyoh3f+
sFbpOJjCbiFnx3Qgic7x6I+Hsi7CU2tbA3d6AZsnu/awLnN96AHzF8WFTY3bFjrThsqY7eLk4wKU
WfXXRj7lEj24wjPwuyrPMV9G2AsiAMs+fLBa/gRP/cpF68akiw2AbeiZlDIL8X7x/wos8EGSzW/8
sCD5Mf1OBnuhiS0p3g6ssTisC6xNQs+GPO1ksz1Ir7LQO6whUlNhfW+ySYfU5cIf2ZVE4547h3u+
KJgYWqsbfIQzFzBSrgjGdi6RQhJmzR3IozKdbYnkUGLqBmJaJr62Hcqw2R/28E2GtQuYwjdwUqhN
u25DYHeuxTK06UEh1gh5JvsoXi5vcpUwC6PxKLKc1vbY5Y7TTSTM88eCAHdL9aVXl9HmHi0Nw6Q3
yf9MVNOQr7/FLeVv8p43CwfuuZr6r7ZUzEbiF93cccOE7rxGfhypAaatrZd3MA2eCMFD/IVkdbeE
6g5S99dM7whiB171Pd59CgKd3VpW4Ct/tQrRCvK7A6qK3T2aHzh/KDLNnY/KpstaM4yd3SDej+1d
mKifTY5L6aIDawk4g+cLKFsRGDm+XUdp/CQG+3vJUbdg6Vm6MpNhYQ+Qib7KDmdy+kw6HS0Sp8iM
u2vyYSLYlPCyPVoA4gosgpKhAXlMTCerWPfoNAWUxbR5koa4aZctyJP+zHQ/Qm8b1J2BmavRu5Tn
gY/F/0EUyDWL15hHOCuVuenysyaUM8oYfaAivukr11Jj2XUombbhZVxEamGBUFKTPVkVjixtCpiq
sjOzOr/oHQY/JigKoqeHRRhxf3zDOJCOknYQ6z+5iNkyR4tWz26s/u4ToFkF3DzDl+Hybq8fv+3U
AKPoXK+KvQF3yrcaJVIm/o2/2QPo+EIkTR273mT2pTBidViErDQHaHAhJz/qi7RSPWY3RLS7eMa9
lGIXsBD10/yksiYjOFHZdVuOemzayhoTT485TesJSquS8eMO0sXH5audc7E5bVtziT3Ig/Svs+a5
pYBw2qVOFjovwUZ69lcIDNeuM2w1bqCKWH/s+pobzjcxRqCw6dbEk7AOFRnkG3rTNCjDHi8PANe2
Izx2A2EGuh0NxcangXmL0oCRPJHTn6Gkef2mZCQvdY9ntZQQC0BkHJ7NoVouDfNzYRYy6DdiQbRW
pDOzHBCXVyku2/l1HpmGq+zKWI9Kgp6heWVRmbvZESG8gu/WI4kyJdwhsow7COmpmoGq5jeDrBHz
uLvZynKR1hpu147XAPzMMXDf1AWQGSNSk2UqwxZZ8yCRlJ/Ta8LYiYU4uqlLX7hMtal/YHC4d0N7
HZ5wYkbDCP5EJ27xZW12I0keV41y+DKVY6Z/a/fkXt2uJZX0j17BKbkNzkell5s97tgyA856vWSd
zH6WLu7lQ2vbgM2DzsJeDz6AJMQlg92NiiotkjbjVBKxF1uKhNX2qWUhgl2MoEKLwtyb8wCnngcv
Yau1omQDkBMvzXrMKPH/GiISCigItrz/qtbHhk8+Nf/USOj+jALPKzsHrpYc6n171MhzxDIFopsq
7I+fKc/iCJSiEt2HSRiCRAIvzPZ4qi3eJzZQgZ4UGlWLSYyFtvhiXJPVkULsrVV+jm4aaQWrLm0x
+x4IZLQxFSaDSAIkvRxENXVa2GiwIPZXe0X/97Uq5aZF90D8Q9gSv6vCtrC/mtWaIFO97swW3r38
OyaKLOYPabA23RwiDDvIzYbxZp9DtrvVOzA4CitfXxdJsfgbNPIA1b+/CeSk75vuUG4OHU3JbcTb
X4hnygtDS5Reha/UcMiJtTh9vA3ifknkRNBTkdoFIFRb+v2CQt4wF46Sj82qkJiLjPPPGA0ukHJE
DBlpGcsxwKKa4YNIcsV+hTIHPTh7lyDz6HsLJXj1d3Pc/Pli6+a85H0Z1WY0eLiMbS2uRzwLartF
cVXGU2tO7lehzI6oWKS8F8X5Kozpz9giimbrfOS7Hs/wGwZ0LDcyFrCcqLAmA5ZVvN6+rbt6lYH4
sefAB0rH9ZBjBFxLNM0RnE7fZIv+w3MC1On1Ea+ajpE6T3ap4mUpGqMs5/Luac5Lyx75mg4fuaSd
wm3O+1OTNZ6Jxutf/KklUTvyo3BUPGG7InIjh2dA8vQgulmLwsZ36iio7+e5Z+Xs9F3fSQJBsGDh
ZLp5IZmzhUEBnoNLXa2eFQRj0vksk93Y8vaSRHILSHe6dTcaDNd9gl3Ht+gHw2Ji4gP/2ZrWO0mB
a/T0oQMTIum6umrAkN424rY6b7+n3c6jhdjl8yxoLPrlC3FPy5G1NHL404puTMht93GCmpvWwxJs
acgFApBuSAVqWosuwKDQrHWLyLtO9tAQ1gq6SA72uJfvntoAW9qPmZEn1jN1rtY06JTGyjORr6Pn
pTAQaaR7+VLuzoOmQ8suWC5Fji0jsuElzVnwwOTD4jnl1uqK3K3RTstARtCXFtu5zssOVbFSirLE
cqIgQkKS5sZ6yr11GLOMBjTryAC/iUAgqo9gT8ebBqgUgfEzfDxkEjdj8X7+NYj+FKqBTBLScpko
DNpCDdFK5538DYYTn3A2/6brtVHp+sG/bO+PaxPU8bMWByIOvU9uEIz05c4iJxps/ci/NhloHUVR
aI+Dl/0O7HD72GbaRBK+Ys8sViBwvThgQUfzjqcVTtPe9PmPLRdAqq+x/PolDpc7fzAk8ncT7KR6
eCrptrfGyPdZVhZy0IrlkT6iWFHvwxY2ItxFI5w9R25q39WU8iVaSYdZzhEw3KVarJfHEvhCGNuq
qre5NfRao8TUd5nk8d3eN1KTY3bmVuD0SqN53btqiiJxCJDnPxAil4ZbeSE6YS6JfGyfQ20tRMUk
Zop9TjYTZ0WH+uqzvyy0/RC7STjbvYb9jp9F4r/uNdeHSzyDqsfAD/QQ7o7HLkSGZ0c8Mob1p0/n
dD7RySO5xaPc8oiY/5gqJxFza1S13x2SkmT3Ygr+f6a2wU9lJPSlzIO+fIyLmruZSd/ujIuhl2J9
nJZJoiay1m5kw/3SG0D0jZ3uE7lFv0aZqGsDFvHblzEIY2p8N7l6TYU7/0uSFCBz28oqBV/xLW9A
OOt+mkFEDpyYn2uiISRbtEbSp3fNVFItRNOmFZ5kXBBPdpdgq8klWRAZxEas/EMAlJhmrMQEdWY9
y73kt9Suktuz+IRjZXh4khFcixg2VzhASb3tmgQJn1zg2mlmFC7iIgFB2IYycX0IIE8cJebvPFci
ruzWf3LDmZ+A5td7qx6/OtXmgjM563ZnOTGw6VdCDu9QrYPVs0lBfS8mk+nlQKQ0qSt5fanSncvj
aiR88V8hpjSdGxO+Q9HkOPtG02ekM63+Pmb64ynHT2doPWKCvNrg9Mvk8VojE6ZKT44HF1UQjB+H
4OykUEuj0cHfWlPjV4BRQ4fRapopt+I7J5iyXNjVP/5OKr4LwZ+KBRSBdukcXLxSMjQ4fKtBpfP1
g6RLS7tVKBRdB0l/aAE0S2Ifvq//CApipPvNRitCbeYCKs2FnZ67tRhooc+GAvfBep/Ha0cUsvth
0tfb6swqFGCxpBrALBwYzZqzbGHAkTtTImblFpbP32V/2CauZo0d+AjflOkHnz/CUZwQ0jBvrhUp
HnKo01mAdPXiXImj9Gaj/3qqtN8A0puy1qemhIbNY6LC/EXCKizs/cUr/rsfDhZc7fen7/rOSsHU
6EemxAkzJGxwxXxSZViTw7HGUOJ3aG0VRLGCkFACvDHI6js8w6N7xH7/isWke6Zz+8O+vPpSURdj
2ZLfteVeYh31ehv3XvvwUqL/86yqTWEh6U9yoHdNuTblGdfoCYWa1Y7ZUq17vNDtRKb7CkudvPyo
pZ2z3nG6zMGA0SHWQfxsUVxKVDcrhiiaTF6yBdHhYBQrmE6E8J3QE+K9vKgVBedIgNVLLiBiYr7c
62wR5MiEHMntf9DgJeoC/vGMsFhVg2xqjzhC1cqmucVAuovfcPK2Y3U/ijoPSJg66182D7SZHQqP
iSsO+HAH824BsHlovpArRgw7gVv2XdUssNOg7Ky0ycxgJ1WRc3DWRFizyzLGlQtMyCu8MJ2/fOui
d+XwAXI6f6LFWlyGtllg66pi1HDwautNBZoHYgH7DY7KcDKpdntnxjMXisjXrGjj8zsWAJ5jiBse
cBBVb6zJdsh7qrwN8KETCcdPYYD9gjk4/AnmdyFwCn26MVzaAIxZToFH5kK3vgt6ENncP/jj5f72
CS8TFjIEf3Ls5UIn+MyPHzILIy7QxgkTqSs/fWk0I4uJwlufSWmo5WCa3nVBKGjLL3KVW9yP/7dx
fVqwUhLy6hOTV0tKTAiaGvBD4ULxQOcqkTQninHEvL386/Aeh9T7Du5aTr8OkyAkw3R7zJhIWhq7
u37AEO0GVwTYfI5iF+Rtgx6j/4vPv9qbKkzxoQR9HZD6Oa1zCLInyT4N4X0/h/LBn/dAYwpLoa6D
MHol6dKehsBYdGBHSYcWhx8zul8rVDxUS674SBmWcNaBfW7hbRpZHT3+RLIvhu+KNQ6q67WkSBYs
PxAqEB80i8rmq/oqa0aJKmae1kwR+9ZYOw5jGUktACdwsTdZY1XE+sIgfCo+HfNEVmFtJUdK7jny
b89yFeMN4aJPYToMomuqTiCiPDI0/y3IhD24TwnTrnq/mUrapIYl6zFIkLc4OskrEEh0cJ98OOtf
EHU7+SAahYG8YBqgVoc9Fs0C1yeDLTfYVFwxOBF9fIyF75G/x489BftYe/CO2yrKdSvwZeNTOKzV
z08TCyRo1NrtwzYPXG5PFNyC57nKCRgtaTeWXdLIUeNV0dv4P+EzU+UTJ/j4hjwGXUrIu4FoKtYY
IQPCuma34feAhTSJJAmIZNJ2xXza/WjYppdPDcEy+eBpBOSLTTZMVRYFC0Dh9nxePk0Z7fruJSuP
mRBjg6g1A1RD/HPv0x4Arvfbm2wJ6Ta6Cjk+bl5OkXht4L7W+cgmBaYWi4vEbSAFJ3z2cAMH4KDd
AmlJ+YB/tO2AyNTKtZMo4xB28V5v140kqB6rQ4p5YyzE0n8e4wo5qZtt3+l9BZL72SUyKiPCaO5Q
13rT5DmQx7hLfnUY5yA6mL0zhEyN3Y/cJdqYKbgaiiVzi3VaCpMwOzSiczQKIC6ilHSlpL69NIr6
OnPcsxzWn5hd4HDWSDtw5vEeu2rCJiEuCkjxIOHrPgfkcE7EDyDl183Bv4OfF6YG+EWwjUwE/UT5
yGJqE+gtYAAK0/wIoyCLKoYYl26+J77zWpCM0T/95nEU9gP9baR6lcLKl8/THYDArzof0Q6m4EHP
ujfQ9iAaigUyDY2PWquVTykr1AvzmwkEe4uFNJA1DYuARxRmIIWIPXCuvCZO2QhykeC0HEsxqQur
q0fCvv1rnIL8cFT0iu5hBKeT2/9BP9XZqMTAnsH88ouYqIjEg1nyycVvnuUZO8EIfLOTq9RtK9gD
p9lbcwg1PqDVpyDOsyuirgtBM8DuiAS1vWvaht4FA/Ykq6Urh8VK4pGWK7Y4pvyjsCXEUM3sSZBI
T8/0uCZ0uq7FZBpwP9CgQgSwqFzqMnFkY3t9GeW4X6kgF7sd8mW0j/6Vh1aMzA7RMVBGB88K3Ita
fxNzKlNfgyXxy4tIE1rXb216YW44FKoqKOKHCTFZMYz92AtVHGAFA+2Oo18mNQWEZRdVeKqA+i1q
fDOELyGxXYUHZJBkkEP1v1z6YraTuIvzbQIVi158hrXtcaXiaUlYDoqd79HUEixcaLCZXCY1+Jzz
yjR+KKiseHV3MufKR7UDZIcmyoWFQz6NuUwgnURvKDAw02rPzhCm3dyvb0+RPgX99pT6fTv7IRXZ
kI31SIvhce2vZ2R5dnytRxLNBS43nMUyPwGbghjkdthzixZsgopGunYgM7NddUnKhQAWh69Qu65s
jVGkKlXuTvWyBSGIdlV4pYbhGDxfnmDPk6KOLHpNsagD07rh68X7Xk7AhMKvlhboguzUmFARs8eQ
9DuV7cCGkBMaTehei4QbkgM5yVxH/apbHXVYxxnfXCUHDUBjGq6vP05fIfYmpqUbqZMwiZ8m5ln2
SHfY+O74C6OzkJtSQYnUGqSLR5iek5W5jxzEjZkuxsBQ/5paKmUzeSTY4YD3KhgooXfxl/mwgts/
IwfAf7TdKYLSNREZv9sgR8/D+0NnKsmUKMGNqK1zQ+geCspXMD619RwDDOpvfDLHT3UkSlU3yVSH
pOVlPcuzQ+an07OEnB1siVbUTLqO00ukiRNlf160xDnAEtXmc6uYcEXBPMZHUPL2LmZUQ7NjGVJJ
eEi69BC1Ar56zg8DJ+43xsiZNADdGgfRsz1SUVRoVTgxCzpyPufcCOOugnPSliRnUCb0ctZoiQHD
ypzvj4oieYsowukcQ5/kA8GQ9D/vdbqoVXjALrpckqzvzkSdHfIYuyY0ExHhBHUGj+gvXGE4LEKO
hVuQYsXs0kiOEFEX5c382Wb3yCy4ooOBFHcKmZwnLy6f55CNfFihGWneFJcJhawKkq61dN6H0x2v
USI4RrNVHvF9v4vOHQKc1V/OV43XR5gNeflkWeJlfPliiO0+q6GiNxUkinPOz53uMAEccSwcoHu+
slnA/t2vp5PAsDiBnpuoUx7TuYFNPyoVSSaz+IhH2ViPDG9Zx6NZGFc3XZPl/JjHq2McPeAJwhP1
ekdK63fjhZ3WQOU1KY31dGyiy1XHX6MDXBAZV266csx2igR6hLQAZVstOlJP3c+v/betzN2LPAY9
kvT8qzpKNjl6uht8bTce8szBqqH8ZRhSOCADYLsmUIk5bS2okgZbmy2dUmmLdzy+T5xrtM3jHUK4
tZOXIFJ2eh2KQzGdTMtfU1NXBdhhyb4HPLwf5bl+FvljjOlTjzQX42bPGoSUr0ZKJHSu63xfg95N
yVqKvqMlhVTt25XsZMd4wlnDpr9nlUR3crW8J0depSxDGKuVFxyo6HEeuXS+e1XNkI23f+ShAH59
kzMJ5ByCuqKuQaDO+MMBeo7ktiXKF8p3xieRg5cnmh8sJ3CJDk9EFQ0OdtVwzt63wAa9Ods1W0JN
v+jL9aByAF8PW++FAHLaIdvmiXoSr8ghsBoQr+wuCqSB6T9wM1wjMv/eDIyiGaFyD0eIdimtn3Ap
U2/6ait7+HWgGIvsd5DHDBhdBY1Asmz7rQgCwMCA1jow2ZinrqPSCtjZLkkgnK5+wuZyl0x/6X11
Ef25fEFaCEtFv5AU4NFAetNXJMuy1m/6R9Wjx4elqft7lFlBnS6s60HV2+Td+Fln/TonEqscR/TY
RM/eeOLBbbj4bq+QZRwaA3+of0/LejqOVG5Z3N4DeB3CcOAEQRMl/1QHYZhZetnyxbchaFKCI4CE
CSUDLKdotZxDGOp9BxpG6ufiMYY+0zSCunuL+JHjjKFZEVnMHt451ggG5E0qqisNhRoOxJNagnek
JlI2h1vFWVjk9he9ztzYThehhq0yKeASstZScWM7WoozBne3REN1JvtH8HonmH3DMqbLROVYpnej
6L41Ldk4Ae0w5vKbwSHVAp3LSDGuk17J1Voc+uWvFMiTVDEhwhL6W9+bbXsf9G9dxcttbdrAUsWI
XsCwR2QA4EtlC2SORFGpZlddauqQlX2DR4lDLK5/9xyyarxIwmTA81+fi+NRZB7Q/SpL5Qsik5uT
CzsEKIRbKZ3zRSzWAvkRBUurfc8aqi4yNxH4mfEVqFzdo+pTTn1+3c721rICfHbfGANdeCX6cjh0
QGSCD4A+wYlerDbwzdh/0nZE2kdd8L7c93U5MOOv7awROCbRDXb4J/f4nvpZ+E4oa7FEOnMrDXDC
2QLnT4zLX9EYacNMK86xj3KwjTT8SdahdhHr5gnfAV+dz/rxLqspFJz82+cCLdgOQNZCi3vLlRha
OKasBf2thNRU6jDOtcCc9c/6ooYikc5X1ywfIc3ZlWRsvZWdqdq0cYVuuF9BVD00ZJb4Q4bjAcf8
0mkG4H3PB7R0mKo4HoYcstIHqIGNuTLJilBbq1uKcBrU1YHmUNttNVg6aEB8uiuoq17THOu5S2eC
Ac444h/WQQwPS32+AmJIStaC1+rgoCZ6TH+693Z2WQt6TqQ9RBbqUbh6beCMQea62b55tAy0h6Ry
4cqELtkBh0TvTKZSdCEp/MwBgD71O0Le3xDwWW/CYyHTgl1WIttZ4d+B0to4eS3zhc7uf7VxH/l9
dPARmnvvKSsAG/RoarGu8T348HOQ7lNRLnMfuOhUkepBZX5cHVzop2mlcnLK/Jh6vW/fgAPNszsP
igqb3rWylgpG4SwE0GCfafq6WrXvdjXJshBmG0qGvZMW2ZO46wv0OLx+TwvW5q1LrHfwGWYnEgnz
6GroTABsPrFJbiLDuXGiH4IxOXuT7WQvDK8gVmCVixCnmOg0zzx7LLtJJxWDiKPvMb9U8uBofXYV
zfUX+IuM4pqZmVwUSUj093wW3aiOv12s+W2LYgNJr0hYMlUUxqJhXDne2ujR6qSAeNFqCJs6QfJY
Ec6csu29GXImBLNs9z37jIJeENUIGtxg55GzITXQ7VGmwCIYbrYbgoXID+IBuR1taYhTWikwQFH7
lHnuTdF6CRxyRR+q5CPNvcSutCxbCHFy5frdqIq5JP2oDSjiLTdxMNI0K9qhmhdWHDsrlBB8nnH2
Ff2ltkesEdVGarj1FB+WOLcloZSpuTKq9DZjY11XC+XgCjkhnTefMtmHLFRiU9d2fpBUAixl1X/M
nt9zSRPGW60C+zLNdFSmJgBs1vF+fS4ULPmJ9CNobeBqrgCW60PmxkHQQfmX2NbaQIrXX4IaWwnF
ATQPS9xVSTwEje1Dzioj+EO2NS9o5QMIAuv+7v+Dgrs1ekTBO2+xyuYQYg6DWA7ZUJ0h+2kxaEln
qPYP40z/BZa2Ue8N9wJhaj8LCykRWL2vkz1O0g9Vwxoqvx7QxI/PorVHsIkBol7Sozw6rkkoBh/Z
ywcwtQSaZYcYVSkySbOz5l6pa7VkjqRI9eX0j+u9gfrDShp6gRMven7N3zsnkVJGAgbJ3d+lqqkr
haNHSi7vFESWr/AljEjKVW9jqY5dsbCad8oV8Fi3jnPIa9mwWtHrk+5LyRCOAPLttiq15qWAnbJ6
Oj4ZTUeBdpO+GT57iINOOlQuFwjuf4lA3MX6rKKUBW4rutLenLH/iNH19SGZm0Z5mSFlc2mQ2REA
CBOlg2ji/vpjHuEQ66NFgpqztrjnKUJGIRZMn9DLkhA3kc/BOd1tWizrsa1j/X7l+T/vhiyfgILm
HCgmJj3m1dJltXKw0XaFty58ckxZOqWogxZADZovgkvQfM4Ph+C2GBjtiRPu37AplngXEyhvnWb4
YmfMGAvNOp0fu4EPvq8lSyfkGNi/Xr5QKgJZHl+8miih9Ut6ybuMVaV8RVZpy7Z0xcZlgeibYtik
FAncag4TLYA+8TZrVrGkyJlGLWaSOK7HggM9tkZ6LYpj1M7YEcPlYFBxcAcp8B+HQ/FE3Xop3XA2
ACQ/mCesC6owq7sQpT8VICGY3JNppAX41YYWsOOwmn4LpdJ+9yPsc2fomca5j8L7YMjv42A+/Lhz
SY7ZRTHk6Ha0Un7wDoLQ3V5JUwZF2/3cusNFjiyjn99bGzrHAL4IVbUpTonyGrQ7eMC6J+5f/yKC
xCdkwbDQJZiXLNO+DKCPzaVs3f7ADi8d2hI7lt/Qoalk8gBqTq9oW3LlJKgJuEcP0ksR1w7xe8Dj
b3c2rAC4dzwr7FJMdEYHAWmc2oALjDvj73oYpWuuak6WWB1xerbZY2BbJV/z9fqfidmXTJrc19h4
1XANu3OOrnw3AFVANZffNg4tw+QupqHGd83ptCiftxGbehjVemHTD7qSy+Wq3q7a8ECixZJLuZL6
Zi9FvebUjvusnLB1roeB19QP3N7/W27N2/q2o+qEeFDkDvdC5diMerXzvGUbaqehvoZzKQgqOwsv
vdEsvOnKW3t6eoF0WGYSMGIQgeIeMoQLH4E/DI8H5ydUtEtl269exddfCXaz+e1mrnAmMJVC6HcI
moiYSk/ctNCYFMS3QM2gSIy+KufX5gEt9DrYeQlSTnYYza4K/7rCQf4W+bPM/Rs/hOLgPw3jpkGK
9EdF7UlamblHMyqKNI9BEynGHnKFTwWuudN5epx3Gmru3wqQDHFjDihBCE3Aih2u2CyThr80KEZ9
whpe9jRLMhnKRmknE14kdJ9YVI06BPty+zBQvAVd4vSuojyzgC1NF95lwnPV4Ag1FXCs9HFA14BR
ARkoJVg6uNiXFizze3J4RPD3VMrYKzZQ60xAus/OVD2Y16sI5UyIwmFdiRipzKtCl1FU13x6bBUl
7fviz9M9VUXGyG+E9VbsOeFibCrIEFpO1F89kpaI48YSoIygWH75NbkVg26ZBgouxzDRWjM8A5Ey
z33lufb2iqlWlmWk2M8eFBwcMLGE8QMS5znoP1gRkdhmEF+bCGE94mkSpU02USQMo5rLP4wnloHu
y9sekSPaoLC0E9cGT/wC7ltvMF50ZP5pHknhaaneDfUu8JSya0RVuapeZlvsywGnZh+A0Jo+sVPj
BFrDY9RZimbfoHmOqmQ1CEJCqU74lsy5R3drACZCYmpZf2+i5DbX2salmRrhUVwvoIg6Ynpap/Oc
wgWZUTP/wZHdijgX1p4M1BTnfhrp52RZSMIf0fNWl97MDdALTelzlE4IkVLi1Ldzrli0W9B17iug
lAZ7R65KBdvnLfUfo9lsVTK0LHdzbH2Wmf8d+dHsr9iVolNVeGEl1PVWeIrh2cerVBzoonGjadVS
k7vn7mg/igED/GY+gJkYq4VWfvpvdg6LBTwVFtUIr6XTt8WzWPmh6gNeXSt4OGPUSCqDWGvnkDw5
W2u7tR9UH3dSkdGLne9a4RbtNfcgL/K5J+mHZISjksLFA5wHv7Hz2RVTF04qujw2CbFjzEuM9sQ2
rj6d3dlNGR37QDosInnODSfnZxZbLh88sKfpDq7nOi87IS+LmpMCgliWjx6Ac31CMSxPUj3nn0TC
jgUE946LOLC6e2+aOwAygSenQK+mBC6UALpyQXcZIyBKQKreI/Dh41IffjLKOLuWWrKjhTEL+yI6
r9PY6sSxfJZ1uM7H9mON0X2f7Y8g2FvOSM6TA/w4afEk10jOvrgOeC8fejcU/ubc8k+FLt+G/w8o
j4BjvXejWbaFsWCcY/NmJAKGJWAoz3AMxmr7PbJ2Y+0uR5J+Qh1ZOFGtMrjCOrNZbpntAsqn709w
n52Y2dUu+5YBBJb+CwthaJdF9UJq5uEYrxj7oRDati5oqMMhQiqobp5Ghz94sxvP5YZ7IeMP16TG
4Emm6GG9+MBZOnVyU+uLP6UiO6DUSu7yIHszwKzDZpToXPt1E0kBWnQ5tCG1Dq4H2pmEmnIIVSX8
dp9xiNdG1JzrE5ngF1dHII3bZGMrTrSAUcXE/9VPoj6lcTVhoZ2CMXDmOJCgUwAqimiVJ1XQ548F
aqQ4CDNoHL7KbnOZrWH9Awx/1SFW1QXYJuI5jejtaKO9EdqZHcbY+fW/LDW2gsK+UpVijSLEHF6D
QR8XQl3EB9b6uEahHCn/FezNzFS48zS5mU3XcCEcXjcDtIvbzVeewu+LEyFUDmIZvqEgXYQKsR91
QoiGq/7iBDv8EjEr6zCAYkjDTWpmumYvyrzy7vEWnZwNRhCUVrcEgXJzyLhIZnnRz5+dcDzM4rQV
hsQUGrEFWoQ+4Ejwq9EkK6V8XQhQGAKvJzJD+VHaQQyrY+IyAxDS0bBn7JwpJenZn6UHlFB9yetl
7FGRqmulRFm2bYj1Q56RVI++ujjQNpL627CqjeeAUByD1IppLvoGhs9LNEghzpenBbm4R7buWK7b
cjRWsEDj8MWx1JeYliTvQWepffCQ0F0hlVqW1DH2YZb+d81FnaG1tXYuT1VxOsca/j0Rmcz4fv2/
B+RZnklqDlkhJT81+MKYpTlAyX+hNX5noRFMDikBeVPwtlNe4QmgvbmZ3Jw1kAOkS17zVb8ywRVD
EQ1auLqiy0ggHQmtOvTBuGNk9KqZWb+TESiYuEEshoq5XWYlDWCE5FiKGSCJI5z9NX70nRevlsAJ
gmYFYw6EmICtgm43Gg65haEvPEWv7gIn0lCALlgrJRgVEqOunDNA5di6hgPLXEkglVdatUGtZ8aw
Ic4G97tfYKs1whXG0o/Sq1mWA9v96FH5k4DQaFcFYNoZHQ1+81zOE+CD01Ni4nkjgdD8PHnhqtCR
bXNiNrvKyVfb+Yh5RoR34dqRaBBnsqX2RddkrSaLF5yZtV/T/p4vdzyOMsiPYCOzK1KXqIHPw6i1
53ODWQ8qN6x6HooMg+f0oMe+seJbA2fEbKta6dqBg/AKKgkeO2rR9dpGY/rcriYqHW978YRvmUcD
rx+QcmerjyGYw+RL+GbX4QeKxDmTvKD9iig/ElpRm9OpyQ1Wi29TIgQ7Vo5eRNcAJHymDVkcTo06
s1EsShcDVTSSAYZEIRGsabZxKIc2shAPbbUMR3Fo/bUbK2ssTqcSjXRQNu0Yw7Ce1Bbkr81gir60
XnA6dnh2g4+VGah+V/WvP4rezmV/6o+RlVDbLoAUqpd11dSgOyfFN5Jh48JVz2Sj9qzJr7DVmt2/
j1EmNuCGs6UhnbAp5DRMlwYHamECcS7iDd6P4pF0yoXsEmDdR6cQjo/sTHEdFAicgALGFm1GiArB
F+j89uv5ymqMqveNsSQUTOEoajmEIQWVaiRHs/quyHF0AdQiufNsq13DekSnujqYFzNybWFfKW1P
+P7fGPi/0asqW4Lgv/EwlagpLZM9bwiT45BXZcQVYHqCAmIdHl/WY1uSxZac8tS3tDTf2QObhniW
EjRvVetkk28NhOkl9wNRoYELOMEf4eQFb3fBr3nuoBhifzGOXI7JdEdFGoYq+zqT3YNx1cell23v
o4m6qJSYL7l3aqdfKPLhY6VxwnNM341UNWpP27/mQJ4kvkLn1cBBfEiRWQnH6q4x2f5Y2yVuUdop
yDWKsjX1srThhB//N/lu3N3GD3k+BEUr3WengfFMuNTGOad0m9a69LinvjhDA56dVAsJCQ8lOksL
9Ihain32upGOkSemB2gSj1cSkeJh7O85ijzcizQEhpjHhpoLM/0rwUfhK5nRnX9dgNTerPh9qXsi
6vW2y+pErVSEwd1g0ZEoU/7Q4Rn0RVDZ3sK3bvcdW4KhwJNhWcEUSdxNuBwlL/F38ZqMtZnabhuJ
Zkzz3RVOE4vDR6IaV6Uj+LBQa8fzKE2j6ZxJhNdW/QvnkU3rbTj8UwmZD0mngDYTf0uMgLwspM0s
hr7A/m90EqSwmjoNv1lulkkHa0UrSCko5SyfN83W8ac5+AtaSCOjwfW/54kQYiC3CK8LnmHVqbv2
dxTLJjWSunYMZ8lRFf44isRI6sbyMU0zpSn43sScbGkAVVDQqbU7N0Csi/Q0VJldv30RcMspQAMv
vk6py9y2QOEbOlQ6ZkWFYQnYaeEAr4bGCVfi/nTjslaZz32noR+vzKquEXQMjZbiCdrD5qZeJvaQ
yBZ7Twr4MKOj9VjIunGG+tb0hw8bPREHwRyH/MJxvgi3W/0kB2VtKvIWe8IuR7DWUgx7WjSNOYGv
U0Mw3Yvqyv3d+dU2hsFm5XItxUSfQNY0qhXp8/CO0ZK3/6S+8aeuKBSdieADBPyRSDDR0ZkSQ8oi
7Rhukj1yCNKcmc4qiu9I7Mr54ZVlTIz+bpHSUN/JpfIe1rVC4cW0N+6KWJ/Q9yfnrnaXL2u9oHnD
/KbACZvWeK+gHzJKq6DP+OyQTsNr1qNE3VZ8kMmIJr4uNhHt6MSnKGd0C2Fb31XhmCQXlbyo1Lm2
9IJjmV20ov/f4kby2BClxNfwolKcPw6ulTm+f77+ebj0nqeVaVKe0gIPfLp+hSXanzyO5SbhrLe0
V6nlKSOytOWykBmhztkifz3bw+Ivy9vZXGNhURPSr6WqFRdN6OJQaKvCp9Kg/PuG/B6q9dvyj6JG
47FY0pQzTQd+PuzF4ffCLYuL3OvTPhS9+yMC2bsUhk9e0VmfFgyjmuGnWVmMd5PObcF/UpYtKbod
U7vnJCFvia3f5XxK5DhmB869Hn7F3PlU1IY5dtqGrS+X6gK0/xq3GrqBDDMAxlP8H/+gSKF0OR36
yXjw1UF39/4Sy68cCEhw2vj6fQ76FFNokh1Rf1oZknSRM+wjkY9tJNWfffE+1O1csPb9umFrvbC1
wZH/WK/X5aRe9we8QsFIYYHKVQ5VlHeWOzLfBTKF6XTMx/n9P+dL0ioWX5BlHmiJt0bg3HdkDLoT
0dNxehggikGwNoOQoa3YtVwRj0jtn60QST+S9inaubwSBgHtjIfq8AOeuCzkQ6IOwI1qR4pkoRZi
WlF5dlXz3C9lA/UDpE5RohIZrMNm4uPldd88+9uS4YrvjAKlKRUD/30p/DoKPiBn8xK/EtEfMHBK
t3qzdrt8Hlr8yRl2RRQMCoDTVOOCjRrSxEaN59g30fbq2pkxoLfGjYrtZbv7Mw8NZ7WrBGHn4CLc
PoFmPJwsTOOSepiftnd/qm//6q9upRgV2sz24SDqAb1GbliD5UjA0klHEcnt6XhosCWwh74BfWod
Gw+HCsGXyqbhxh6xIN96KzgvAkvpDSeeaYIfqxmNS9XWh1Zkm5+NpO8fUAl9B1rucbr9qRpFPLTl
ZPT0nwK6jsVis3c+cyw9Dj/en4TanZvWaU8YScaYieyD3/bXGgRSyUp7yA48tcuT00z0bhjIG+bg
dNQpZTGpvQwsuNOr7wHAAmuQfYgfacSrVm5/XkOvIHOWYHDc9HFk+Fh/0q3pbOwl6sFOFoERAvjm
i6rjBBxqlUsmAKkcV4eNGuqtLeMPx+htxowE5ZPX7ut5spsJkBea/+dl6pPbzBNZLzuW/vrRvQYb
jSoxYix2bUS+7vnRGIOhcjHDoo4RGlqvy6xRZz7R18EtW0L3Rd4VyzidE5ur22w0+IyEf5wA7ByX
7v9HdFenbvksGv3mohdv5JgZgMKkFdKqaTptJPJkUbY72BaIopTZ7DDffJzLrrEc7hXGGSLJF89x
RALLZJHZF3xM7sjYJ8a+NGVBUTZ8QALDrnmi8PbJR+7CfCadq24o8olQ7iLeNjjZqn27ZhbV0ovz
nrcO+dFDBIc8MdzNhj5gTx4RsafIIvwtLFx6UKSxH4TyUUAbM3AbqFYTwjE5QFuwBfPfwKt+Zd7c
qJ1XDIKM6qBRgYj+vAhss/5BBKHpSatlIWqtmzErU+gcrzjuvZrMrksbjYlQ6PhyMapAsTOMtmTm
HuaxhgDuq2tWw0gQcJpl7/DTrPz1CInL/cHf1P5gAVNr8++XUfsdBnxWvEMWDADZPBWX4D/khIg6
ghObgNE+p9Lx4H9n08iWAG6yUHBmSFovjcb/QotxiWLcshUmbdYBauhzXsqaurbfYPPwXHF1w1MF
kT49dxHefC14k68fHXfGAZ290LCXayhjRzqlivr0ANnFNZSRy0dsQeiCe6uWhbDIgtbTi/RrnR83
7FjpxK0Go9prgGRlvZjq79DqsU5OOjpF0ss7BasDn7q8gMUvp1EfmahnyW0IBoi8tiGqxXxgNLQ2
U0cm86tOiFl3SrkAHLZ+9A5vs3tlTVMDe3cuqVsECXdi7DOEHV8oQauMu35WA4CpBjETSra9SFne
tTyyXvaSShlYgWc3LjNdDNdrfkmxGbKNoLWxXCnluOoDSlc5iDwKWbuR/P2BLXcMmeI5dGYoN7Jh
ar61Q/ckY2qlugydcpXBIdOsH6jx0F44DDnD7ePX4Fv/MaAjci47yoYXZGJMvCaxJSFN0OicLlTq
bJpa19LxsM/g5rkVrRgweWMENsUq2LvuHzhiGiX5W/sm7rrrbF5+0qj0FVNc+02Yknw461pesLGk
YqlQ1OLZt9DW/XIROkRpb725djL5HCHTPgiinqIcUfJTf/FIXt6ActXx5cX/c0p/ii/DcfCXN0jJ
cnxyYm1pIoVTnBG+i4QjJBjtyPtKSa/B4kXPHM3JzTiXroJrPTbeGst1qSlg1ZHZUOByoh2LS1gI
V6BNqB91Wvnn+252ulGcPYphLTlaiB9GTyE9pScjg+wZxc5fENrpFhqbaS/DK+pQrCqc9siPNZ0R
QIWAD4kKa8zq9KCexXk5brGlble3RgiuamPIb7heZJMC+PSEFuxEEy/wUxIWopZwtweL3GaezkML
vzDI1nTykOlAUYrMNFQYFa57f5X4vRUePAhJlEral12NPHUnppkwTAesktFN5IhtqM5qlt4TopZe
Z3dMttlNPCNwo/5Sqb6Cd8BXLyuWRFWPeBAewu/48h6mwuz5TLC3PTgE5bkTT8XBbJ2yFEprNoYv
qHCWTy9TMmKXw4AYP2VwfO4XZXlsVt0Ek1TUiQXIdJpWBd1OgcXQGg0MW1BkiVlUIliVSYIkNhpg
J0l6wcJCOk36ETGVi552ibHLQwaluYth2AbSDAJxGyg4B89hww+V5M8A0WkUcuh5OWUFoz8U29+w
a3wQp3jdPetyLoQk8feVgNl5ZjDAOA4cFolM037FMVCEZIybbBAFyrnnCqU//x1RE/s0888BKIYD
9BVF1rqDpgWNRjWud9RuEoISsCTAcCFl0pGnzxphtnc0/HA/piXIk52lASAVLDcATgC0o5Zw2JH5
Nb29NEldPTiuwY9pMwco/yXRyubVsgjoEoAftcB/gYDQ6iPAWhafra3H4csus5TsrgSW7iUthcSi
WoELcebJ3ewTBmFZrdwtX4lO18SV6N5SBG3C8pm62i3krZbHvOg0JV8B4Nl7DzF5VZoBTO1p3xDc
HqSTgXQoMp1k+rGOlkZbjPEpX4cMop2kmW0LHx19Rckogp9tzH2cJeJwzBZjLta4DTIRKYVwvGEW
7E+33q1qiOIQT7nSfwQRFRkUexOEDZMh97TdK7N1qheZ5FtEMqkrc1ZFq9KW4LtKlBw7yoHWDt1e
3xDKf9QCd/3XRsKuQUHyWrA2s/zxxgYW61O7F5ZY1JvsMFQGAO4ynsmyvrRQMVvmXmz+RCeM5mk9
gaVTkLGKpaY5srXo0z54TQ+r9kG3mVWk6T2bVKHU0mFPjuE7WezRivCcWPh4FqyrXQTYyMVFh2KL
o/lK1DiMJPjsQcebtRy7vBcVaP5BiRSiUxEH+7R0XNzFjyNEScg37KWJ+wDwLDofLj730PqPXpMt
Nmga/PrST1ghMu7J8YApssTxsBJAm7cezXWu+uiMUY156Ai+HIURKU9WJ9u5hktR0MLC79LCqzUG
nHypHcp2mlKgGM0fEmsZ9Q0UfIE+LxyVARsf5eyVoHdsQbntjVDPJW6Z4kKmYMnP/08vGC8mWfBM
KbNd/IEfMjdwREkHGAw9rTcvnBPVMIPqDU4gU/vwcgPFP4+b4koPScrx8nbPvZqhuGOI93Y8Hsed
B3XJnbnlw7TSucXLRYoX5Q8O+1kv5mxf1GQf+98gkf1nkV3GzH7ym4s+83Yr01vooS4bNsSji5Dz
GzH++c4mgmlJi6GuvCaPhC5FDJW1eK8IQAS/D8aWVsN0msAaNQabgVdxgJ2KHT+gZTDJ+nOCN2Jk
DeUTLX8brRViAF9m1Vc0FjQI/znArw+iunfomgfnVlWUwBlwNgAZ9ItNw0W6vZeYU6SJ5WthQZJ5
0gPG6mgTeXpGZEzPVcFdtAQ9wt7COlc1se4O5ah3cKAk5Qw+o43YsSb547ztY4FWaj6DDM9+Fj86
OOk94VF0Zia6i2ysvTNKKhNvkzgTJ5evTR7EqHZ3BJgyEeilg66w3ZaNaCkIRSd5IW9JqMg84GKz
4S1Rl9BDKF/kBGadWISg131DHwOLmVkfXw9vLhCdqCvG2A1PpIBJK61gbt1prB4FvnpDJt3/tyWt
nKOy0BbULzLa98YCxjTLQ2rKeKy+wjFwKIqOmAMG7JRngKTNXExXiJxRM562uEhvTAAPAgHneDVk
t6x4znMfxIaLVKTOYiE87/qnyrRhmIR7Lc8+GilG1ROefdI2JCyQfrZAeaHaePBYBvhwoUupFCdC
dJSfldIRO8tqvNnT2d1tDXF1/vXb02V4jEab+VS6/TEqYX1ycOB/PMzrh3MP5jRtz62N3ouRQq/x
fbUL0yNwDhKa6Z4wWHQCxA9L7Qx2SISbHytKHe48Q8ABLoTOGcjF3SBgOxgNJpE5QD21TSetwKxZ
aiXKPwgUYwn2ES5c5UEsV582ggk2GaK/bZn6A//trsAUPhhZadwp5PbJzGKnT9oTX2tkdFcaX1uA
R3M80pCxZnw1iseEGMpyKAiCUVmcjSprtJyYZUrGtLfFOg2+yEfZb9nB5R0wiTF3QpuXFP173QlR
mHZiOxx9FodIV3G8ARDG8+ULs0lQ0JVLzmGClSYTHca6fsO7lbpZgZ0ZrvDC816dzQneqjU6bJXl
wm/TOb1z8t22okO5NF3L/W0E3X8BwtfLkECVJFBL//CL9oFvd4BnsuUecamFWDgP0eqQLZzOjj2H
WjWl1Qy5l4c+qmHZBhsEqnDLX1vZl+q7WLAQauutY3DafzFUCHOY3GJNhHEjJIMwXnOGZJ6UAL7o
g5naAIaMgHWSYbgtqmBDVAW5MAqaclg7xe3kypoxB4ImaeC0IXJFW+Oo+QU1TLc/eltq/vE8xpQU
4qO/ej5JgyxKVfYZPBJeOpkVbQN7lGyzj0Y0rOZfBaI6Hj+30JSYnSQ2Acwp0OTedm6S64hrLnOZ
nYeVDA9ws/cmhl6+KrVrq4Yh5cGklHbt20zuWWaKPQpWbOH+57QIABmuuLN9Meb7BUiD14OL8Z9k
GHL1Ey4WFwOtAj1up8WVGgfpu42WjzM8aXMeyYF6cJxgzS5eXpCUmfpdxKKdYdeOEJMvBolzLNbx
1MKB80Qv0iKJmeWFnmjB85AmZpcWsRgzl9IIC47cQfHSqxtgjKAH90ZRTi1Sk6FO4FHWYYKKB42A
fCUp0U1aKSF59BK06INnJSD98KI0Cv6nLpPfxSd/ssdinV4fzXkwYuLHNu2UBFDiAzD51XrJBVul
egENtlPjXk+8Sga03I0gWW2XUudsj8VeeeCnI5ENSrXs1D0McjbiDVt43pGPCKrkwuaHlwnHPgXS
8MAqiHUsxxuaXWP410aswaLGH03+09i3Eyl0lv2T7TYwQc1PySjsypfpNRAc7KSgJQ+HHoKm7Y1i
j77eVywxECigIh238bK2cghty+RpZrij1mB9dpCbSf1bTj+bPoco1fk6gGIAYvuIqjHBKnG5hRfQ
a7/Y6vFJaJPa2TzDYg1zlOy4fHfAdO0338njs47o0nI++IMWuYXopmmkYYuIKRdQjIO1zUGhmGVS
9q2PwijmxAUjl4LB75TgLtNOFtc4wdxX5rXBGL7BWbU9oQ2n6v0s491BcpJd+IbYXyGU52ySSD6I
sjvDdSluPChFnxBDy3zoJDl2evUbVjSEYWQwtIQRcrI4nlZTU1UeOI24eriDiDCS2Tk6u0fNszf2
UeeetKCXwGKm7Zfrrwt57zce0JbPJL22C0mzyESDlEi+RJyLAoBX9awf8AzA4SOjEnMyTZJ/3tgj
Jzj18FU4P/FKo/XQnpkvJpeUtb15E5hhFaUiRYJEa2oCQpVkxNsAw6RVaARajUuHLioCBeAEerxH
TmqJDV2HaMUzbYgt4EQ9SGMuixvqVK0q0y2coWVnO2dlal+XPWW3TnfoTEFPcGvvH84ugbKFge9T
IQgd4My2btZq1Ntw1/9V+Tr5Q5Lb4O5EOrd0qNHf6HpakvksfwcVH394Qe23vRMobhYphesVBjfw
dLuE/uL9vrLwpNBV/0KUiNGpy+fPRYjseMoeHHn5+FMZXv/lxgPJFwEEDNQAyimv2YhUDjUPr9b6
66N+J31hc/ROYI+PeCrnIWez/+DOq1jPAJO4hjE+Q1xWcyNWihEZI/3ZMAw1S5nmhAxCXAe3DwFP
1czjZ7ieidC1Q5QV3K+PWhY2vJD0l+LprTNdak3kTupfn3yUkK1x9dFup+WFFkzfkSyWSohYTxFs
1THH5HKhqil492gOjNZa4ceLmL55wKdf+qhCmD1Bn4r7POc0AfkTwu420iBhJu9ef+QcQheU5GVp
LYMWb6CvwJpMWbmp6R+TM2pRhSdBzMATf3YavPT4Iu06LK+DvPqTKADOhsUMJuXA0T1YvqqP/YFW
MPnm4xz3J8lT6XzskGx8VZp2tabEHMIWD+/3kAskqxlCPZiBwGhx/teYp+JHKA9nhuo3eQRIf/Mj
+nM9XIuu9+v4tVwNP0zJQCqqGE3DTSuJrdcbH+M+2SkTSAYvV5xnr8vyJiqCtUTxalLFtQaaIzUx
yxQ0VKUVrTVpwQwD8uL8BQN2x7VwYu6KRbCp+FOalsVZlW4RUbvEjqhkUV+KaKI1AGA1t1zXWXcG
TkHGn8fF+jV+tG6cmSE7wKWxzwV2KhUPQQlZp0j4MY72wLui/JLdw1o/cgWXU/81yldOZlJ8fQps
3Fmih1kfsvj4B4QBn9LhatXxL6KzWv9PGudYDnFBz99nqE4b9ha3MNhPfTW/z6kzzdNF1DETJhuf
3zW3rhjlhXqTrYgIVcgYns7RUBhkEYwbfjp9uQC5ePKBFnca4CfzLt0uEXZ3dgfRVgofi1yz19hX
06w33P/853sR4yyUr8kGYbPasm45tO253/slK3z/F3yppqQlZ7MnYsBrJqZi7uNTFEpIp1iJXIwE
4jH7/9WkY6d8KgnazWlHKxrOAXW983gzii3LJ+RtXDFNnkGPKdsDn/se1vZfnuv7lKS4ANxDpfP+
0CJGFBfDn+xTDbKj3QVCX1TwMGZbhDBcBHhE9AcVQ8f7dkxfLoBagbflmilsp963kGL1n3qC4F5q
Mt9nACfc+yagkr1uIWIJtQnuNIff4cuJWk9DkdyQg6rFN3RBjigSe8YMm4smKJjo8dSKBMle13B+
L+UjlSHDjuv5iDen8gyv6vinkL+Cm/nEVUBOSgJJZeo8XXJH+zh814E/gHP+15++CA7v9wAGfRL2
WV7bEMwHfKu8lMbHT5uBQvbIJUMFKwIS3qrMv3dDf6PEOl+TbMXBAIzZVaURGcCR8GaKwnTpkxYM
9hD2JBuVBHX0oSnAeljrHFYUi7NWqw9IwJ8IkTLxHkUKKmUvDUZJsAnDtShallJHeINxYSolkFK2
XsPi59EUi/R3NoWZOL9drn2KpB3CLy1E3WK46AcTSbznYAw/d4QEaCWe17EgIbf3TOQR1VMW/NUL
3Ipqx4LSPgWv0VqyOB/TrXQCJsELiZvEkaNPovX7izerCQ2t3lee52tDFWlnXNw9jzf0o0wRmD88
xA89eRTjY45uJfAYSZmsGvgZdvBcuUEAp1r0g93WmchE5WRmYzwDp4puYzyDPl4UvVbp0wWVWdcP
u/B+S0+E45HpHX9jU4nUAt4gKdAeq11sX02flqhEyNysmWnXjF1zcMl4h/nluApihZcxHbV0/AWs
GL0IqDSFxa5vodOG3lw300cyPxgJb4kvld+vnN9tt97Jr5qa572i7rvkAX4+xmrV3lbrimXsglPw
JlyNV8nhJDUalM2vr+1DTpEUNOguW8JdLFv9OcSrA832zO6KP4WWBRBliT6QHBMwr2kjel+qnwaV
Zj1IRzMbm9nnSrRQW2r+5yJbCBA6aE9e8NUbWj8Q85zANcbfYV9SXBzKdyPQLL1gP5mjFkwOsrWs
LcD77JoQiWtFB/TJNdrnmXl36QN3qwyoiNHOdb9DPDsCzKI9yIxR4gwbY4bAIHv66tZ2qD08HoQ6
3fuWYdj6lqJ93Cd9Ig6a554b2VZCoGZMxiSH2wVLBlXiY5QlAYXG6uLFN+eHZThDgBt7/kW+AgTh
tnd8NifS5EOK/q71KyIGGEcOaaCA/BR/nCLcBv4N70gy0ysfP6a3vd4QECk/27IcUW2i/Jffw2aL
MUb7p+hW5KwvTns37+81QsCt07H2oEanHvL8FzspB90LF6k7RZRbsmKw0gg9oWWCcc2qcQ721Jlm
ZF1HMe2M/1EUzUvZSNhCEmZ1x7Nu5luZ6sIWY3+dVJ7KQD33pYd7BwvHg3ezZNa0Te0SE+/xpP+q
joLI/jfgnnsh2bakQ6amMxImkhdYzSzQkZzBAWXF3Ol3DNbthkol1bBusZEid/auC6qWShficAiO
4EMyKVSaRoUvo68x/Hw11ZJYyEbLZznqBPh2UuanXKjLjhHMztEO3dXqbf0Ci4SB/BarODhdy4NH
1myrjJlfcPs9ln4pFW6wDsBOBgDTPbQQzqmrI5DPzPPoQjszBl/o0rcPAxu8siSnreugp8pKFTlF
CqHow7ptmqjFh148cII82CAb8DJa8subynCifosiczI2S2cs2A7Vh9OpB87eIQfmwu0BOEWqoGRx
r1GA7OWUGwZ7K2wOcS4bZWQh61sgFZD/8feEzqJ4MYRIjHi2rJRyWvzdu79ufYQoCj2DEqZKya71
NYsTWrb8rpzEmcIADoJWxZCbFBWdDmqy3/fxj7tfJAbLntLHVPCZoQBQEOiboLtx6aCRpf7ZkOpe
OSFmzN2LecL0alq3/ZpXLUNoP2IGigb4ntjj0H4SCI+UgL8d+CkFCaRJyv4rMyxr7aoqyHfmAjHy
jqUv3xmgDjHHI5zNxT6Nhkb5qrajsJMf7vFGxPLIZFqItt7N6DcSrkwlaen11NSIUVFpc6c9JtXd
gWd9ID+vkg+xetCJemGMFz9qXYveFJHlJPUa47rpQRM6epDKQdZExef4+0A3LgNiK4i7O2cBSg2m
34Mcl1cZaIu4aMA4qsizOaEwzQAv/e8QpOzNxsT7d8MR1zwrIrVt/0dypag8oHyML/rgTOr280AA
5qZW2pC+kkssxbkeOejq67BH3E2DXsuaMr9097+f4EOFmvZxMhbplGdHFJfvxZrfnlxVApwur6oO
xv/vMeUJcchjTudm0QL8TzLT3M34uCTrDjsc81RdpOM/qUnqal9Dx7ddMIWrV9LN5XF1kNLoX/N1
k6QIdh/CG6IznZS1FGjm8XhEkj65/CuDxMz3kbAw0eKlzM/i4s4w8brJ47nT+9AwGvemYV3M0u0r
yFV9NNAa/kyXWqJCjNjxSurn9XqIFBWcVhlC2+6STF9dOepVvxlTSP/vairp3rS6ThVNXMjd1teM
e4pLwmk1IryUUXDHiNzu3MydAvq8QMF6aKnkISo8cFjNYmm9HPxjQPbj5lYE61LcdSt6Tc+pqHxl
g92J/t3COH2/sZQqkC/67ZZlyLBDRK38J5zWKHYAiyRu+XPEvcpbHeWhBAZVirMJWRulzlvJh0wW
ku+mWsWqETxaNUWm0j0YJ5P6hlrT4VQ3winAEsc9TKnMYpramRxXAuJhbWtCZ5zfYwnXZjvhSBFh
75qjnhoyfOoTztALW/ugelh9FZCKd9BLOHerXhxbeE8HnW6bxZvSBpbhNrC9ungUgIV8mnKMxi8i
wXs1a7/Y1hkwjL579J+yJQ+D8+SH86k8YLIP/6jxNfI/uTegaylvAZ85flk3HJOF6QHto/iFihX5
q8j942h5GYsdjAnUJLdIn8XXnFHOixhfAQApTcOcnPS7KQsJ96EPBDFy8Zp7LEsy5mo23KwDD7wN
EbWWPgO0Jlro+7+nRUNHMwdJUX1YAlqe+xWTsVYCkzMd7lMPISCZ+f2x1pEpevB/fBE7HDoXFNED
izKevnkShcatP5nmNQ7jvk6iRWiJ5NrTTa+VFh6EaYQ3ULHLgQ+kTBISzGGcQxgFrtn55xHMzFPJ
2LVz/tQbIM2fZfZrqILK6DGsFbO7Dtnn9Z3Eh77NeqPnfyuNHvgAukjZLbqJgclvAZDbP99VRsit
cNb9ZZp0R/dt+H8Jb98GJ06JICh/Z34vwf3A8hRROoPvQiqVT3ynKPbZEXc20+zPrBB9shvOnvxz
ttC7kuW8SoJfYAhqhipJV5kACxJsQjdGXzk0seF/mp87Kyn0Zb0YM6zd+nsoFCBg+sD3OmRejXIt
QXLOQ9c//vQX31jAQzpqIp1SxvdizA/QNqrVlfDTnTgEOoqIlg3VpwwgQZywZi6qJEX39Oy1nE01
1TlxBqb4FOdj6/TsgLd+ecKZbgSYBkAhkvjy8F09tWA3Ajt8JLvu5X/pxSDsSAhvm2Sv0yiCBEzB
IRubS2NKSrclVDiQxdS/nbi8zfML2xhSFqrFUvyJ507AtIx1c8+DVi2E4251kn6B7RWuei4Kxqyn
Dsg7VXHZ2yR+sC4aldpWmRWsiVi8EtVgdY4jN5hJgXcIn2RR5UrLKVvCqEUlxhH45Ts8waGo6242
xwtlDWbp+KmKNSephdFHoZEw4Kc2QA3oDTmRJYUByNWAvzEimVMVv06uXxsQEYPabHy2RvPyddil
w1PnvrhCteVMh0rLWXM8QlQxnCH1sbtvaNEcSAWN+cTCEwunCzO7TpbpZgIWkE5zDQu7yTVn6EIr
0bFL4wUds1LQV69XmJGF8TlSiSneKbc4uDkn+cVbsLzrVWJ873+PxR7Wq9WITbj+J+NYnBZgLrww
G/JYdh6OjZ/Pv+RmvIXcGe9RzHUXjxsZ/e/DpoPv2N1PW5csdyhvoHAGdcHFqXE0mhQVQ9bfJMcI
oQnbV6p+VSTmFUs592XiygDp1YOrIssvhji8w4NuIA38eAXrwvc3S7FuZ+eIBcgGcSFwIZf7XJhv
fLVWy14DJXv4EWUFldsz3Qh/puUOFpW0rPHGw7Lbx0b92P+Cr+QNWpKhTd3QJycyfHss55YoqY2e
H9j41rL5MjFS7LxC9Lo2aDaoImFd9baDakc9RP5lYcFRLWHPjDYOug42OHKJ83L1R4/fq/DjLFjM
nF5SVy2Wf4ugLnrzozAuGAwZ9PQTHZf4w7L7AA2qJG7tt9Kx9xI/fM2s/CaKHc3fwE7Q0fJeLMFK
jom5H5m4mqto8MNVpUhwUiOHNSsUq1y49NLNEkUsk0KOs0ILnB/EC4xwiv60TyX31kS66XI7pJKQ
OQmj13nsjP8puvJ68O6Itt+HS2JokeJE44dFcdJIC1SeANhIcOlwVk9MuezrR9ySIhpxowikqnBJ
UU5N8ZpPPezF/whXrBLwray6ZdoDZ/cSl10EPPHwEgsnR1TjEBHJlVuEPQUXdzJNOTur0gXwdcgF
1vZXP0rlfXmOsRotymTk8dH5Lq31+zENs/PRBNdDu1rpUhrlyXzu1X9gkwmnt9QYYm0fPjs41iA6
9d494iKm/49pOWzybF8NB04I6D8XVjootjJKTPX52tGfeb+Y+3hh2w0HbqxRQsUC1NomO9c9d2ln
RBaCVhCXm1BsWrr+YALzFeSWlVo8lXK8zgUtcCn6SekLtC6fccutVLJ0W3bubysjCjkFNSCSsLSL
niKGzEXhymfYbea6AKuXyrbrlYn367CugPCqKAjo+ur2+pHiMUVITm+pUIVG4E/Rub55EX5NHB4R
/nShYm5Lr5ZMB6TbqxoOPeOvlAjDnwwcOmg1Ok6abOmb2dfqNj40gqx1gGPXwZjvrDBjj7VgJMPZ
bEX3s2uP7pm6v09o9pnYui+dCKODO8bOKzfa5h2vGVrPGHw9of0TOlfq2wAF75gQW7ed0RWjDBub
fjhbKwaEtEbtDnUVEux2KPfbSg9i+YlFTLRfs7hykjLKQ/KVLmQ3v/UXB83noKxzHLZeoazy3yAU
RmVOVzkeO6i9HyuCC4NHPqtk+bFfvpJ4YeZe/kgbuOP9CKuCTtopC0RJMtI5plrTqx/k+KKYnSA+
JGKTZfxmLLK04Tw3mm4MXVrZUfD1SCMbx0w0y6Rw5yF/xUSRzfKjlZD217mJpNSBpNMWgMXU7efq
PmxQ36VHIJACoNYK5VqDIQsir2fpqnkL3iJLO76/CST4a6kxhgjaC5wu7TIDx/qylZCpXzN1KEOo
+YbNgIsZ8bH4TxpwtfQN0AWFbTafP+3F6zu8UoAL6ljA2WOVXZPLYKT+OiI0BxkMcyDZRzGF/AJW
03O+EbPp6lG9PwN0jGp71D0cV0UaE/tMjOdxQ9KMqDjddcAmwckRcvGBGaiG9ywIB2+F8TmDwEd4
zcZlnaf6oLv0+8pZJQHu3hKzux0O3eocQhhiYwHeN/T/3nPJ/da0Cwy/3O46PQ8dXm0fozn4qjRx
e/YJIjoWqMau8bHfd8bI2xou+4udiQjkyTBJ6mAOWhocF0Q04kIcINeAUj9B/fKV9RMSPzfcituc
LgRl8lJ8+S0kCi5JxRoinFqWRHlDJSb5lSEbQa4PxjDoaiLUhMVcBu8SslizlTGYgg6oIdphwXiy
ASo6xiZJLWgKxsYaf6N98hU/yxFBfjoL4Xi6lheQ4BqJLu9ImWpfMRHUXFIzpPcouCWc2sxH8FBm
3sEci9cCiqIB9qzeaAmnP9b+7LQ3KHoe8kGaleqPo5Y3g3H0KQV9jWa9q3AomEGtnpZByUByrc3+
UVj9RGcuNtei8jrERlKn7YHP6x5VDsMRfOyIRkO6liCN0c3TQ7Sc4q4qP7QyaZOavqdfy/A1h2I7
cL1WNcgLzPAi82F8VrbGA3QSqY3q64aXgv/8wvIe6VDPIW2XakAtXwVNVFRbe4sbeZtdEtBZbel3
93ebe7ozJ/LNqxuwzgbKVJLla0VxAwH0RaCcV9dKNxFtpfU1f2lm89QpjfwBGJpK/w29eJpTj5um
84to8Q4fZ5TpSERLQq5UyHodkO6U0eoVPOj4mWOJdUSYbljpSCSA7Lsq0tpD9EgO3ZUOMA76D5zX
2Et/Z4iSVy//7uV10Z1DL6D/bcHb6/DZKHwSSgrNfgNfmFj+tYKi2YQVLmf9svpd4wfpPwtZX1la
sgNe0XX92u3unmMMV1hAHYtoMppLaxZWsQjdidWfI2pDRY80sntJQAJ5K+xIn2wDlAAJ93IwWyzX
zMlOBkeF9ut4669aBXljKOgjSJjCvYVY3QNoAUD551VX3fDUsboO31isnzYZT5005ZPSYF48VlPq
YXyjrJ7ruWWE9PHmozNOkSTWsAdkeR3tqDz6mWSo4VANAMbiTZchjA8Qq/hzW+hKhc0iM/XdMMAK
1vOj4epDvaXDfp1ydSLhvw8I1Rj9ERX6LYzgBdq26RCnexoo2XCRnGEco6QdMAqCCCsgQk3ZP1SZ
QwvtpwKJqIzDK87J915EGsFbTo0yVjxJ4BLGDYjuNrxtKG1r+TcXJtJH0XX83Sj/2KLU4yHhY4bd
a3in0fULsV5RSguFDX4OH0SRrbTPtk0psn4WsON3ytNSwhb7Zr9QyH1y1FvdEfwg9dxBsIjGoCfm
37EFsK7Bl47sxnlqvpuVDj6dSs5sihk/GCG1dnNowLSYrTykngR+YVoa6Ludqp5XyrkK7Vq7IYTi
AMLRdYwdvqLVagrO//UWb5bJeVMXry2DUL6XT/j631DXyC7TwC6tVimL94djPWb/wPXdgH4RsNFm
ShHkOdTcW0TGJr8DAA7zZGPyQKEArZpvfDlnvTRxflLUz/F289+GWnSkn4kJKp33VhyyyWDHMOfc
HBwhfR6P6PGZDpGi/+dWA1MOxJtCK+Q6BWorLijfQFIsGNb8zdRgzFhwAui2Tta4uwTIvbBnn+FT
5DgQIKaTxavUzrPwwvq8+VNqnJUctKbemGBP4yURsqtCvmvf8GpqHSwbnoOTgdGoNYmHAKbrEYhx
TwdvEwoapnb+2rgIYk2L8811MgefP9OHb09qVEPm25WfDKT+dDlt0DKuhEwtg7GbCA4ELSeKfegw
mT9A8yQBhIj5+QXwIZnLXIXV77e/NQ4U9Wll0rddDF97U3UwRQTqtd5NHuvWrfTne4zmLcQDkYiU
t9aW7Hgk77Hld6qwihfwUWxDTAK+2TjOKo1ws8Bag8Jt2sJKoWWzXCIJwwwxe2DNg6AxqkGYmxd5
2iVH1YYjoNAHegyhAN6qbqzMugpFncsGdhcjjPnuTrL1KsVQ0VtzwsqPC2K6C0nPRqZ510wiwZaS
7guH26hSkuerzT0N3JSoDVj4F7Bl1/PoGfdqgj0HQ2RiDX1DXboe+9eK3051IxGkbxoj3CPrd/kW
C9A3Y3JXrJIn/SFyPhgRe4RS0a0pWiLmk3Z9lOQc8N5FY2Rhst1kkxeybKFqQKe/fmFDCu56zT+v
OxZI8UGYAtRy+7w7ou68ML2UF8soOUfXErqiAdPA1NyYcm5QeiiIcVncImxPwA+avShgJFitj3ou
hwEaf3iVZ0/vDqpx28orKdBcxIgce7Nr1EuH8EwMVklTxqQVDePsl+LfUUzBpS4bkwhGtW+krifT
J5du3kHB4ipkqozOcHadvseEqEl7RF/2gxTP6c5SdrFrMGKrXA2VdJO4h6Fadqm/BihY8TdcBD+X
CWrqJkLmhx1zMprRL8nOAT0SgGk+N5EEWxD6kNVbDXVqWIe0VwSDGWP3aJbgZf2syVDgUnSvp0qS
d7gOBCA0YLE+wZ6xGf3CfqRw9MZ5sKvq28YbI1DQQq1Yay+hJfHxO4iey4jfCA2GtCRnybzaPULs
5w072djhKwPWVokBhUGh2r/r4Tpy5r3YGBZBICebksMfgM/tQa9+JmhfdjcpYe9qwGGQ7q4UOmiD
s7hiuYdR0KagnF3AA7OcM7UZGDIreB9JH3REtpzX2cjqkuutJ9KUv0go5+C0D2zkaw/Ey8eH1qHO
L3VWeJ05BgLxvQINda2Ye3DFqmgB/zawLh6pZPkMPbaepk4d3obqzIyR4PNmc+RC6/hIh07AGMRp
q9F40xbM4PM5vl7t9imiFz0AcS5aS2fuv9BRwpS+431AN1QX3cvhdDVzOZw2oCvY2HoJAbFKGz2m
lLkJYCGDmq1pV6zu+UAqutJjQU4EMjCPaNxM0LN/dudszY3pJpVBJ6E6tWWIEqiY+R/PwmqhE/sX
4nvTQG68j/ztFSwuMqxnC4xxlzGm0z4iSA5BdOtkVsyx9o2c/TnQklRZMtRjPOtQ0sFTViCxAhM5
qS2nchTm5PBmR6GAuqr73ZMF3P9hAwMKv9EpOE9OfC/eO9cHTqPZkFQrJKZY8YKmqhM+gTra2lqq
JDGIN/r3GxNddAHW8XkeZm+IRFXooYSPsjAl19F04VWIQziViWU7p+OKzrqV0tDxcXlcr91FskQF
Pdd4/kdLO2RFJVTiGDkdZPNTpRF4k+DD8wLGMhPQvMY4UQ1XyLbWnmDWgX02Gzz/QfGnYQI3/Dnb
8vZqFfypKGxqghqvRKQzvz7N0obV3eog+SXd4LdRUo7F19/QHN690LmFxVbcEEoeGGiPPfcrhBW7
eQlSETZng5FIGNrULxdJoA07vLp3O4HhKyg15PvbNPfok72koDEopK32/8utoo5wVRIpPmakIfu3
XzKREGkCMvFRPRgfZj8PpjYWfwWpJJr72RI+deIPovzr+G60+UM4vNnZrtTYXMVKVIU4GRismT9r
7PzwRbrK6LLRZc9QANS4/TJwpkfC7wGZGIQNVtX30PoG4ScvcVooXJm/0WNs7cPTS6vBqKeha7Sa
PRqBM1lgZZct5UUWSKZk88L59bzezVLVmNqv/1rhk+NPFCr1n32HPABl8HJjEjxo6KhamUBCS/RN
4Z67OduT9b7fvXaixL+APm/d/bzu3qu+m9mTMkMk1gjqvNanXGLJIPYvvybQDJ/FyaVmBv2CBR2i
kMhTEjkD0hfQ9ycRgPZH7G+RXNaAR56peSCJQPBi7MQ7O3sOZj0hyPfIBSCfOEJFoI0lMIAuY/mK
x/gmIkFSXaM7CfdbkBNyr9MhWexydRiGJBIWsjayD15+lq4MJ1XeTYcBWEs+e+tp/5iY89DYpK3v
YJBPXZ97/FuPSd2npOz3a0llM7+u+aOwqZQoWR6zCLILvQv0STV5rS45kY74Jke5B59PMcD12D3Z
z/lvU6fZMFt9/KU8B0hDY7taImSiNs09zR2IAP4S+Nhd5x+LEGpMC28YgMK0n6H655pRWee50EvP
mxpGWRFxUPYvC3HWgg6CeRAmu8cHWkcm6S2su/Yi9BT6bgXAvlNi1KFGIaIy/t5adflKm3pCmym/
IAUTKPg9x0pJhyvxUAkmtkRHfR57d+t+YM/c3cbcWrtwnC0yO4ErOdnCQKc3ZoRnDBrJKTfk/q7h
zBWXGs2DVNiSPx99nika3T9d4ACGZUPr+zv2jUEMtFMwwlYRlbqRD9iZNAXCzMyyC8veeINUYkQ+
hMxLYLcx5gjv9IIlRwJ91AAT7/E0UrYI4MzVvIbP7GMEzD3Ug2Hm9vuHzjaPYv3WRrVKU936C4q8
qp4eNffnnqhBnHSdrLT0SPpPwNhOUCnyjKc1ZVsIb71wFYLr4kRGXc/JJokfOqC4jp6EpeCRTbMY
YukoGOlMSLXOL4fo8wtrpxK4w2D3lsFxFHTKps87tM+DOv16QhDhEhPLrAKABDE18cpQPsgfn8Nq
YIZ5JaybbN0z0Hz6WHjYIH3JXcOjfDdU4Wmp5dQoVvKqhILU98MuXmMb88MwSAIQb9GqfXhfLXCw
cjn5RGNmelEbnVtHz3mdkLtP2eedUX5jEQXhCLX3zkxOsSw8MK0M35KHLe/jDgm6+4783OIYh0D2
x45mi3a1xWZEHvpK/joy/xhsTB73cxljaLBXFhy+o1C1giM0zhUDKO30yK/EpK9OsZKh+jvh3Tsj
sPPbLGf6t22r1qIsLsdzEf7ervCiHdkbiluS/lCmMhjc1ZOFx99t3Yqe/OA8ek/BYmxPX5AiNwQ+
qA18vvsrs0gJOkLDfne6WKY3/vzPUQUjwKZjmHJi59/Le4qb20JcTXGFGRN8TYoAukUb5SkWKkkW
JOu+04ZR0i8DFFKRejLT8dncyHEv/3We9xIS7kng9CWM3AfTPI/FA0sq410EmzcxXxCngwRC4Wbl
jJsOXSLc7ru7Zy6uhfxTFG0c8LFQ64kAy48zB4tMrFYeqiYIfvKYz/3UhbUEF2ra3gd5VAfF4Kd4
FBrkXz1EdJ4nl5lm/0WXtg9G8pTPrtJCCIuTHqAzQXK38ww/IVyOgBD3J3kFyalR8frO0TfuegEu
LI3db+64aRvJQzRPiKm3wdjkr0QhzA2W3gB7M+dllbgUAa2517//SjQEitu9MHEKm4i++LFP+ptJ
3j+gS8Brcg4rs5puTj/8LXvmNQIJwASouDtRGS16c6hBy9n3Z9R4provS4eZpFSonIt7u1qL7/n3
E95HtDlrOv652TAKIhyMVN/7YJR65u8BcihmlVQSV7RlTsOoJmRUEz7kSFqF1rMuFy2fsC8hFjb0
tXJMd2QbHyjXzKk1PnWMe6DfRphCIIcrbdZki45Ruezar8veHvgzMDBKoVXKkhGW/hInuC865FS1
/iDaNxtZZBM7K1UX9ZtDiW9jETqYNb87nKgs/2Sg70lAOYfS27kfXbwpyMRuJpa4U5cBzGXZUpe3
9Fq4rRz0qUvfm+pU/UE/yfbeAJ13n+U6+40c7sbJEZJhruWS1CMHRKOAnqS1tLb8FL9IkgsHpNGd
ZiZlaP6shCo1f+49YbKLB0ItkGgdZARtU/TcRBGFe1+nywgNzIMxkeRX9lDWyXnnfq2EYeVwX8ds
WFywRU76VIBaQxo9TyY+tHPpZH+zgeCSCmyy0TKDKVHDEpjjynPEcFdYc3RTb//VnJTDjTEXaJC7
DU5EK7xL5pwtS+j8pKHC8lYYhxuSlV5LxJkvQsWqOjbiBFH8zC6zMTchA8ar1fUzFUjufK3+YBVu
Bk8djQXB6JFeZmNLmmqj0m5dJCDnNP2FOvPqSlwwkt9DbYrMX+2zL8NuQjt1xAPtMXaNuWjtZFK7
ZRJeUZN5meZgvNTnLgswPmHrn4ObZaLaX80UHLH1zm+tCVwB2v5vWR+33dkajcLWXJ6Tzu24mKY0
uXbYInfimWiIq/Xv8QW8DafMfLeKNLahNcbB/kY4r+ftGeYmGt8pdvDZJlKRYyIYdZP/P69e/SFl
dpH1wdlqNdiV6AFczf5MsbzocT+H5CfnvEZvE6BtIq6bLtHbZaHdlg3Ksjv+SPZ38SsoraqREjkr
okeN26d1yNhR/Rmqg7/dx6OI1xlrRoHakCSyFccg12J9wSFj6eRPHj8MUa1wdbQOtHTO40ASGS/H
EZVh5EGBqbC0aIr2hxgycSC4B9V+SX+3gjd4De+g1zpq8d0Sc0UxWFENuFyBfwxUPhbO0o9zUqET
y96pkqfjbRXazCbS9SPUBw4pe4GX2hQbt1hlYSMVWr+2t3Uc9R258THxabZe/qRZT7j0FRpT1KIQ
xMJtI3SGZg59HEbbojZgYD4EfzUeE/ggFXT4rrrF1PNQ9/HEZT0eIr4Z3DGJBLmkCEWqFHsGhuF1
hGLnF5Mlp9Kaj+a4S4PWYwwdlx9hj1ZE444RZyNYzXotJE3ssAImlQlz6aJEqGclLOJb9fujMOHy
kebHSf0SB/MQ2AXriZpYWe+ZPxguU5A+WuTJ2eGHJQM+rovGkiSTd0mGh6909VaQmZmU72MvsdCf
/nUsGCJV2+uWTP9UCqLM9LU8fhOxyTGOpewvLhn+DUxfeqGnM1yX50lIh5UNi1zE+YCUoLbrq9+o
PTgn1wmiaoNNhloOX9mMpWd/eaz17D4Qdoadb0t3sPHPNUziZAfJ3EcdYuvenPpqKS23mM5E3dL1
S0+KvzfnVKfBXsH5lwrfaltDCNLky1b19T0ow4OM8SPniS8MkEH2pklfw8PggWNZNFbz78F0qoOR
SCFnlewJSzHlnE5DaNkdFJJn8kqIhyprBRl6TPPqJRLHNBKFH4omYgWgtfYde/hVU7OHfBLaE1Bg
fKkIFo5o+9C3iq4jRu8Kjf+T84Wn3JWttgWhDWBMLIrzYI/IdSJ+NaUuJ8hx1OdxKc5XZm89i4YH
/feMQRMBXgutUINdf2MXQPpNz8BF2G6mqXO4Xi56m8PRJ8F7cF1ycow4PonePlJq2nr19fM/PgN0
ybRQgYSr0g7kJoWcMBHJHyPBwJjy8leTpd4XuryLKgoba7FLhDzx0O9mdug8g5KC93/NhLOu6+Zq
gQHkQJe5408OXaSvAU3cEH7oU0QpqPtEN2HUiAbakRtpc8pkOffBcLHKM6SSYXSVHl4vXSnMrlw3
AOaQ9uSPya8LMk7g3CuoasK7JvqHAmrxXM/H2U02VOIReqTZRWW+XdjH14DzW0bCrdYDSZ3seGSZ
izBtv+h3UIam3UOxKZ+6wg18zap5bDErCV1l+TfRvOI6b7VeIFP0Or+nY/QnOZIh5FXWLNXcjR8S
bDakm55KPKWMElrUPkXmsz7uNThy0MHQ9lDOEtqumMlnwnKYCZk8wciRD6ure3SyMmpJhwEkhwc/
rjmA7jNKEFV39qtPBgt3R9F04uB82kWOsqzFxtBXZEcrd+wtpzjDbk0oD/4+kC7Xct4sAR75BZt7
7vk/C/rP9pDz05G9DWn6bfDcR44K0+UwCprGqIildjqfpDGzPiqrZtOJ360EOgCvh3bgYDbSwutT
Lp/C/uA5S+xuEkiMlVqYbKkuMerExdVGxpAaBeXSdpW7vqflT7xiWwCBDNx2YE56/DzdFw1ysQ1v
qMnGlquEInDfKNGa/OfOetGpv1phLobFOFT2sGuZZTgQKzVaYV0S/rNR3Hv2JNFkit1D7VNGkaY1
pWyAKQQ+4QEXvB46RY13SYhSclsrViic6HyDvTDzQbFNT53I1InvQ8v5gfaYFlagyUqlSKpLiSg7
Q7/bsG7J3St5V/AoH239w0y7q1NaMSDrFQs8pivj+2QJy+A/NItiFwtjQ4oWTKCrWh9Tzu+ARxuL
qjnCbN+f/350dwma87SstLis34W3FYstf1x7O/avk0y1kMpsa+hQmLwpKjChp+w2WBnAIe6A22Kf
eEd3nhvyzN5l9+iztsvx/Y5nILQRkfGIit5QbjXz7tUb+Hksdmg+hgXWdi9BBnhwj4cxwWRnJQdh
23ex2G0NausNxstz8zbtHWfZFYW36BsQMxoM7lqXdyIlQte3JR8VuEx1CBrur5JBFC2bGr+4Nl7e
rf98QQbSOVg7fnn+DvsuBS/y45K27tPgCGCWBlhZLEqgOaMXbjhteeOwhpZ/aDj9LEg6SaV2W6Em
kmwtLqOTW/7+seo6lxCunD+Zrvh6QTOsvPmyz9PYEV0B8XQIHQTB7WkBKM7U4hMa+As0sZ3p+FHo
Clst4cALCwAJPYGz6KvCNTqJlHGOJqyVM6u0aoDqnohGMoBjxmrl5vaxnPeafL9q+mT+CcMe45Kj
UUSCzHsT1GRGmGIzP5JR90GhvZQUtuQyPOkoocZ/8yPJ9zBMWecSZERXitIEs1BqaPzf/KVGeok2
T4XDJhHcQ9+Kbw8zkDDyTdvy7SLbvN2hDO0T+zaorO+l5zuDop0yr6l74/8u2vH8X5ij1q1QTzzM
5CKbn49fChgLlqrgxQBYs9X3VGvgmRy2F6bztg56xqObPrayM0TC5jr5yDaJ4ly02V/9kOaeEZZD
TcqSgM4EI8rvd9H1tXPnwIJp6uxnvwHP1z4TYwMp/zQsozcIjd5h2VnIm/iedN1txs+6Cdrb9oFs
71KP04PtF3GNy2dQeH3p0Z+d7peqdpO00iSOPIMuQhYW40qcpV5QXBA2DVJYJSIlVsH9LLwb4iwA
vxz1aOlH7p+0viJkHMrVVBa/GSlXY9bbvMh6vB+HwbZpNiOLPVnO+pr3bt7JNzupwFsOZtJr7uMn
vHTd6zNwRHSsIbzDVRXoHpjgxCBFjwws/a3bBBFXbJ3HN3mDq+7D5YWdomAR08ra8/3z7+Q6qFJN
bc3uG5LGyIcwinBtZs5ZKPImUPdLZ2DvqOoGXalajTxLfKnVHbgkJT46cB192g9V2DpaVHJd41e3
ae2KmKh+k30IK4SWB2pvTcX7xM4Sq+06BEL+q0sagLq/cHaT82XTWiUN+S4puqFoJqkFaN5eOmCW
MyPHA0OSjoBSdVEo63RrDnlZL8TEr7F/AUTEvv0vxbrlowQMwv0T6lct0TbmpvGnPa1fBgvV9b1d
Uc+ltgEJ0lWecn09dEud9n+bJLsVkWDxvG35u+hhKFRj3Uslq8d5KKcmf6VEvx2QOUlnjczDTSsC
peLb71U9zoN7bAUan7vNi13Mww7EpTNUv1XSwKBDDkjT5X50FuAnGIAdxOo7k0izYh5mLe8SmIEP
AU65E2eePfwaFpA67seGsU2dLvGG1l1vxy4XZ3Z2rTQnhuz5k6YnDqJUUZR9V71knDWhaoc9tEjt
6s5/lDCq1DVcGSIMfIe0ditXjHr1YhoyAH9LRlW5T+SItFru1+WoQIXv0J4p8PfRsq6HlLyDcNi/
Nu/HZp4Y408Q6ZgfG2jB5UUR/ceujiLkRPouvy6obFGawpgmilnj23Gad3Z4ZUEaCWSE/C7yvdRu
1bhM3gc/AGijcUSRpH71FaZOU2+eNeH/9M03XwFPFmJRQbq4Q7Dl3DBgvu7+EIxbW+RGR3EyYP8I
Amxg+0PUs0bX3G6H0VGnfM/UTEiMF/Te9Slg9h4M3hib5Ab7lWIVqACSqK+GjgctisAdJISUYAbg
FheCqni3KlmJTMhfnG85rReNlSV8CXdNGiQ1R6EfNydQ0weLFSj/10rJ7XW+DQFojDiWjncwudQH
ZxYTty8iD/vHGkDfdlxqPLe/bW0aFYMqTWPmB+Gnfg41ezkRa91wUqhCRxhgVyCuVREofyOfKbPJ
7y5BKr1eRd/MZFlI7dSatC2PGxVs9/lby5Z1LtwIapy9pZEUetvb3bJOYhKEOhlVpS8OAOSxFbPa
faxKLINDJ6WH61GdvSxucgEVLtHT8YbFfsnRT03Nq0F0ZEHYu/HgFeZ4INIB1ZUsrVy4gPiaSjfe
VCuUDkvdYPZNDRC9xqc9JBDuzhPyzWm7Tn2dGn7hFcbql01+7TkDL5vYbiWCBXz0Xvi+ui1FdbMY
M1LTs8tQR5yycNrgCKNTiJ80U14Gik+PGQS3lkESgwm5S36fVTbrqzTML5BFS6arVHO45Rqz1BX/
9TYLIGAoVKf80xWe45yl1tkOEb32rSl/arGro7+Oc1URi0MdSKyyy4OGQ0rGCtrX3RivEe6gr6tx
R0cV7rRDXTjKKiTOV90bwvaKEPCct85yJbJwHbxE5UExM74APYPfwc0mLpgDoX4I/v76hZDoYNUr
fNKwruMRu2skqtnon5ZT4VKV7jypcpFOgdr7GmP/3SLH41+m1FhWtg+iQiXKZKNzVGW7J6bGANrG
wHN1YVkrRsLwH3XVnmYx3n1KqzydP8mo8Uz78ymswS4LL+DzErJS5C0OB5Wx3fana52+s0x0NGPE
O237i9saVD2RInjzTXKlfJ4dCub5ZKBBp108xh7544twYnzN/hdFUzhcxOQQrmbcnIOYjNpkK7c/
6nDn1VvdIl8B2azg4mok2amMBUJ/fMNnnFEigGiV+SXK4Q5VCteAGj5cuceS9BKpVhoMWE9MGcg1
5BK2tyzJE86g093d6bRwfoyFGUUbxGqEDS0Rg0qTg2MuZ9AmXGAUY7TQ7Zcc0TLIGyuZZBAkf3mU
wiDSHTz5HqKbTLMTChVb9v7wNK9me3BscJW8PFtesX3b39m6xqvMdyagzY83cF4/STevasiPbnRd
xqGxc6m1EdQeUt/FFhNuxjdP8DcheNJFMsNmM2TKryc3PJwHJzszmHWHHaHv+jOlhOc9jaMmkKFf
elw18GegstTUZu4IHQaYj9ZJBC4Jw6355x77egtJ8hexcdCNRklwew/UzEsOli85yGEkYUengcmq
AVb5FyiFd8DHG6FoOCG04TvsxHTmjWQZPQSFKvqOj9xFSMlD2H502OdfTP3jiNFCvHMzSELw5yuC
nnNWn+xHCaIu0rmEcKSv8tZDVBhq9cSeTrJxU3qtAZoLLNwNoiWi+NWzQ6hinEQZl45wHdEkYKl4
NRnJZKvA2riy7QoOECVKAcyCPtyzvED8de6Z4I/u83TiGn8gglphNzvdfuMdrMIW9M5QMcyNGfHm
SxE3P4H+fy4/+lq/T/46Hb9Gu7WghDbtXgNa5lZc4ZZgMUMzxEMuqKMCrFvNHH3EdW7Bv/nUkSLU
cjuLDm709PfpIAh4PzeTGMrCoPYm73D7VLVHVLD9lbjB6YSg9j6SQN6Fi8IgkmkJMQ6U6gKyWyCK
/rdhSlq69ijtd4e1DqpnTaCDu6tXsgdN2Ld7+LL0H1MqFEioK+Dp9eVVxxNNZP6KeKmXTfatumj6
HG5Kcv15II8oK/Al2UkaACzjCA4mttjsGmPpeJ+qRnOqqT+nb7nz8UAKpwa2KhEXF0+/mSiAV2rX
8riVZXrmsQ5W1Hh0rjq6GjbjCqYlRrXYiy43uDpWgcRAwAvQo2vMlXae2jQeF1aFy+uhGqIq3MF9
QIKIsho+aY3vGuD29epfpjTRlWBJRXXvqa1FlhjMmab4iCNSMTOHQUsfS/allL2Hl7L8q3gQ6MJs
CCforFS3Bz9Q0kk3SXfKAkc5Um3X9McU8HobtVm84fwRsrMjUxadIYb6z7fdpnFReTHUMfT9vy16
BhqtUyCOr3enfQ7iFDKQAlP1zjJKp+J5U0sKWdcu7BoK7fm814BLX5YHayz22XkKBu0wc6tbNLAz
YvLy9e/D8Pj3M+c/vsUXrSprqoiEZU4Zs/inBPpheG6eoGwilulg2zrGsXMnrdUaMGJsNJaisl3q
tlUwHlGM9XNxvP1wprxT1KhlPnzxuvv2LszyxG269WaXWMt4fWO4he5z0EGgWtRKzPbfUjrWJ6YW
XgfOxNmtx6BDKraq9RK028ge6lAGzv5454XGovSBDiHDK8+xMXu8FlRpgErt9YSF4nqTcRJyUq1Y
dKJ1bmQ5Yxlx1I4OjXrGB4OwfTA2qrbHDo2efPSIAMUBajOGJP/vbqR82PlqW9wwtOLU52Ib/6IQ
Zr5pOhPBFE+iOjHNW/S9RSclQlQxMgYvuj8wCwC5/fcZ4uqHdygOkmt2qlQdMNI20ueD+q/BJGi5
Vg9eC0+LrIZ/ftWt+GQY5C1OrEMhVmD+aUaQMFeaoo+1MoypGdsYWH8/N6EuwAvFgwuE8nmDfQqW
570sPBuk266nUyInPK2Lnd0rH5Oz7iZj4o23HyozW8oghBqGfO4Rx2IFIfjp8phIzH0EwvWNsOIj
t8tUvG4PL0qZu9EISnDSyXw6O9uuLDa/WOQy9pHrh6pq0eMxFNuJRgP3Yk6Z9Mrg6yjyRA99Bolm
riLKMUzPQyv4jFYI0rBKE6sRqdDufA0ldK6B5sAWqxp/2yeT38xsinmTRSVm0xdir+SZzJ2i2AW+
iMZ29JVR+Rf1DdSFQe5m8cb//T4ZYSu4956EZy1Ys9zp/YkYvSzTVAfmeXDitCb/8JeVmYMHc3dv
JIY5XwzIhJHesgfmjFCo20EWy7RKw2uY61qLRuNAihr90gYlQkBS/T37o3GK6/hujmaNigwARkk+
JIXmJc66tB4PuDepJCiVA0WirdJoRGsKl8fULMgS75GOi8AHz/6YETVczIBp8X7U/bHPH0BGJlbp
dR3IuI0vHJi0IyqLoayQNCVt4wudfH6Oab9R7vU46Wgg2or76idO+vmJ3ga3tCe0wWYqCibyydbP
N95NySBEuVORaYtx0K7fXl8VgjL4Yh9WHOxbaVSChmcz6MrUr48gwBJ1nrRJWOuQEYH3qfsw/hap
zTKNCuvZKuQ7ZNlzuI1u2MggmD9WDEXyLwkK3KP8AiyibpVplCaJySZUn+84atGVk+c4ZnQsVePJ
Wv9U0OL/bYDRUg6NwVhx+O4fXRsKwG0QSHcNR0ginR1b19Zf4T0nJozTQVCRg1dMYefWnWW1SuxD
SEEmPZWPWCXCEH6esf7tfgKszC1VECZkE6Rwb1ivubKSK+ac3VoRYqImWQOw/J6eqjGJR3wk9m4C
47E2QPAOVzkWDk3P00qrA+zEtq3/eUt09hUD/n0ZsThVq869lUnTJcdil3SnSUa0rKcyky6bt0qw
wu6dYvIJKBqubd2BH7Y4YOPDGpmOMNDQT3PTsm1eX/KrvIfDTu0Bd/gVYOqxzoBvdyTmTK0CETvX
jDy4XOF8+cgA/jlXOd7AtEa6f2XcDV1m/wtwD+j2OIovKMiUvT24Q3lvtH129e+3M3xqWbY+lCc0
V01zG8H00uoi0cruz4zQjayP/1s0zhzji1XNZEBs9grpVCRbu9lz8jsWKzzz4axDCXm5pUpgVldf
ydudoGipPRzoLIwfcLTB0bmB/abcm9XfT4qFfqZ1urkQnhons7NKzudadsWH4DhWu851sZOurWb2
DjAA0GaK12V3s/UCMFLdFASp7Mn/ayrCXhPmvt4n2BnhxL0k1cGtVO9XRqGLVnFmfhKlVpr6DeY6
9WiBewnNhF+5G2B/m8xukpjyAyA62Lz5Xd2wjsn65pttYOb17DMuExT2kBL2UunEnGd9NqWix1UQ
KC0YBpFnBesgbgRPIQ+2Ja31ArG8HcgPSdKoLKdxc7h/EEnBpEN72Ld3h+/9m7q6oCgsn+p1ZLvC
sNy6op9D5DZ5WL/jG2IXrJzQXIGoTSZms7gMgYpk1sV+vW1g9cffMey/Wgu+K0As4jBGtfZZImWA
g/EPBH+jXyre+80cut4jU2TJD5gILvfvkU7MCHXV5Dw9gzeao5AYsIynggnYJiegHcs79AZxP8pT
ZRzOoSV3D2LQTS7igl2f+ZXjF6TIIcJYlcX9Ou0A8RTco0HjPAnhvjrzK+sFjjRzUmBH/lZe1M/j
PoGXRbVRxAVWdLylhrCwfUA8RLaExGopF8OJNQyrBZK+ybhOI31nhYWsEsz0y0lgtcgfhxctA8TH
DXib0PdKEl3JbHxPAm7UfWwCePw/5NAo8WJNlUVzhHQ8rUA3h4f/lSDkuICqvyq/EcvHFZHs3uko
/pqboTzunhnOg7ZqsPwiSLtrKG9EM6kSDGBt6yoAxGJOAmn+c+8ixHUk8PqPe8uEIbYhIrSAMwdY
jFbrQAZboLFrbgC7cUF9RzOLFwu0gM2K8pI3UrG+ZUK2tnVMHQQrH54tqcLENtWVcyycSnJGHoZq
Zipuweo/U6UBPLCqS2BFlnQ06wlmfqrj5ntBmIsbBM/7PYvcOc0e3hAtOU0VhoRtMBa9K2f6aMOH
Yla6q313z7lOs/Wwp1r55a/fIM/hC0s4qryM1ImuqVhLzQI6qivSHpFMEqExOSlAaBKqKGYMOmIo
dYb3SMyJoMEtODta/djdQlMz1fga14Zt2DrwqzJGWCrWKFRuwKEfxFPh7QSIXbo29sS1YmS4Ds7Y
xgpX/FNxWePikyuJhHScKhkhwfIgKBgHiYfIupQ5A+o3xbafYAE0UWCahh8S+hRWLgO+PfRvNiCw
xmF6j0CNhGOQg3rpEPbLguSCj2IjqNG8xi+JosN46wZ+hi6+ORsa0g1dUzfI8FPfcalIMWKGSYBu
WmzP6H18vN4r2uBEKZARfU21lMOhFhAt/kypKEiLceT5GWVPja8IfuNsExmwpIjZyNMHVuZmfb7M
AeuBcyR665WF7KZTrvKPTX7lH6x7GE5du6zjzOq3oLainj61mfPKXIdrxu6uFakwOz5GaBm1ccDJ
6UGTghsPhN8fj4apq/YPS5jm2NPkOhljLelHdSEyfgUOLJD9wwHyyCcb1P60brAj/R6aI9ZjnW5J
NwHAPTPpBlWON0meuFAUbJuXFNCbZwhfbv0xXmuXgD+uI1WRsst+06Roqp9FlXDRIRKhzyCAgAEO
I3SiosAEslhzl4cSKk2BD85k46ky2+WEOqajT0TPoTQMjIxq31v+52EbzQ1uaF/XhxchcVzIP7F7
ibmYVA7YOBbmU16pb4yUrjoV9rX2Qpk+icq++c9/fsiM8yrvq+3AHnZR4sdLN/3E0VvP9gwgNOI5
ZilStKWmaGGg4WGZFdDr2QzkPsuGetylqx0BkM0G89aL6uCSJXQfX3bdqLIIAWrjYGQf0mz9oHCy
zwS0sKYtiNvYgpN36XWweJezAU2WbdFHnygiRY5CspJchnzEqD6KGl2LTKG+fgicOhe8nf+FdFKL
5hu/mUEZa05C1kKxXMJjbMLSTpQGgk2pUfxKcNUOGNnvj+tNiGRb8VYV3k4ibRN99nWQfb0PY8Ls
y34X+9tm4RVjXwz6WEq3tpyLTTm0mtrPcNQe80kP5FmxYpkF9MzkAmr94AHoIIAGyC1msOZvIxlr
LRI5bXhiwkEWVQT13QWMBSpSYFbnVBTm7IRc98heB19/+/kbNGJ4Qa/Xbd1TaoiflHvhTKdjqWbh
p5iDVEp2o67jx9hZxDCeW611zcWMMC3y/iWuiLO/YuztkqraEaCFB0M2vdPo/kmyQYWowqkI5mAn
AIVrbzpRt3o57x4Qdgi6cIkpkRa8RYiP30ixlni9o/JG4Q74lBofX8MbkQlep/I4n111Bz8iZ4OI
uRC2Xt/lZalinTmk234vnS5ZZGcMRU/JA8z8Dz7o5v086euvLPzGBfl5O1pgSZaW9W1US+9apeNt
6/BGNkC0FQVsprxCp42fgt8VhoX93i91wYjquv5nBkczsdEv6iuYu+3dijKF/SjHOuFsasc5XhcQ
mOEQf+v0pqH4Vc4ne1/0BITQVQl0PZhM6faSH7mQatw1eKhor01J5aoTWI6by3T1OKc6MQj3VVyi
MBiNx2FSyApYv0C6S4gUL5w+qYWqtMmHJQDzk9dNt4+zf8oi+tnZQm+Hh8nZ/9ej5xKaaG15YBpi
+dm6U6oKuY1gNWYe8w9VyqmEjqRngz52IQ97NSN4O0ijhOUw5vh2y0qyW/BkkEPjp0mhvjuuTV3C
9FPkNK5gL+GmVIZZOQovEMQcu8xCK839spyLYafGi/RtWGjAjtZ29B6KqFjOwM6lPhfCKCIZf36r
QE302xS1SgKXWrYb8ztt1KMwSbRdQrKBuNgOQf+3TO1AccVmIxg3RHBtdArUzNRh7rE3ArXd6YMy
/dbPkQMMvGF/zcp4yr/8weC1rqp/GemrIXHsImagUPK8YzgEC/h53qqJHJSR71du8C7gTf0jXMIb
h/JPfkALDBaA84fBQPvvIa/mM5av+s9McbVwo15Sh39qwZgWFipTl/i0cgB9q4/AZCa52jh4+KuJ
7L8QxB4oDO8dkEoC80wh34NV2JUL0R+cSzXcbOfsYqmtNINmiUFHknbjQOed8RbeP6pW91hH0oTl
Q/GBaQQBOnAHLvTWAmI22OQT7hiszoOCTFA0R9ZTMHSRodppZWRzUjSQ+pNOAq2hho/EYFZVozE8
x5IyVXhs7uTOmcEyo0+ETn3TgKx2s8fp7GREmfC/bal3oXrWLT2VMaGbEIQECEUGhlwBKSz4bt72
UcmzqGsxrfmzNDrCXhhh0Npf9Yv0W1Su+lQH0dHZWN7fysQH11grGWi9g51IV9zVT+c54azAl9/8
GOf5I1nIpy73Z7DZHWAsEWTrdWpJLYrssakw7UKm7h7wm5jQfsj9bP6DF2ESyH3LAcRr/8t5DYUX
yN+9TfKL4M00RfIcWZfUpeme7bAvOulvZJggcD8RbwNFpOomhNDM5W6qUN0d6tKbk81kVfZLdj9X
afUP0SjhkE2rBOmqRoRZ/a/wWe0ogHNHvKu0ieaLtufYzHOlKbWKMeD/XvB4ztXUwAetd3tgAivx
LNCoGmQQM8c7O2/ZkwAZI+xbqb3w000e40MqxfJ5QY2ZIhDozF+WNjrsSdqO98PlAYpR6HEjIU7W
HLb+Viu7DJYPuPvNvRwonXotXySFWPFy/rA/QqPh7sbK9Ktj523k0FKonjAuQnOnUI0rBnx1Ekrc
luosGLGWSWahgQsGCnUW1lFAWpqZT0LY/auInLvhFkj8uCugePY25V3R/qZkpQmj9pNmvl3hkiGb
/+n35vnpNnhTmuugBUDHXdCWwZNLUCLwPwbMgOOESoIUJzr1X87L3tzwDvS4Xa0WjfROAMNbeEyU
SJfWFhVcndbm/4wdi3IeHdtiEQBKD+Jz+F97OJQPsiqbjbVrP0VhNwCPz+k9wk86CUU1YSpEKfUH
MwAANCB2iD46nlWxsBNQWhqVVfDAE6y0X451lcWQNXOYL2hLmSvCf7uMIdfQyxspajtyrlM/mOM+
6+6scSlRTPelKRFKhCwd60gYEQOwnNlhavSlK/h7HlO8TOkdx3Nv3b9zQCCBQz3KBn7cVT9YICDT
6L8wEyQv9mkWvFYnmeyoWwfo2p9YBr/ZmDkwzLUiSj62aJ4OSqy8hTfYDXfOIxahSsBpeIWVfy4D
ZP2Vxclc/WnYOwswtNG7uvHaKzPpjVaKuyVdXxWWD+AprmEqC0LGOUJkNTWypjWFTUH5pHO7LzgH
jfvo43KOz4Moo0kCqFGO9Dl+SKJ3j5fkC+zpvXZ7ukG1BcrksUu1AEop8thmkb/yaH9tkoo4x9uu
vSIlRUHF4rDvYx31/Y6tkz7yuD9oimHSqeD2MR+blrLbUKKLNkxt0pgu2G6lp6pobVUD/V6dlCTN
qCFIFtF/uerrMeC+6pLJY6Xgg5sswG4ceS0vX7uDSG3a1CruS0MeiFcDAHbYvVRlp1VGJqU2gFWI
odonex/luGQKu5UzPxQp/iT7XVUa8Yfr3MLRjozjMtEVJ7FppTkzc7l1juH+gF+ecoZ867txFAvb
T9vvnbO3QIdd4egtsHHwEQ8PNDX5uUcHoXGYnhYTLjDxLAHjzoGId4KAVddRNw4SZu/rKw1BJoY3
Th9AR+OWCXUp0ww3fpm1/lrBhE/ly13eAmx+qENcatnBPE4Y8lbPjZQ2Ol5YNlqnJJwODGmhCs9p
mxMtIQ3WveOE1KbkXaiF3U0wIoiBM7I0XudhnI/j+8U2AGBlZADkOg2MpGLmduSimjb4Lxt9SDD7
TEQkxZE84atZF49g7VfbpdddSi3Sls5Sl4WBhnI5GB5zbPwi2inmSV5BhDwG89TuXZ5lI1KO6wTu
suXcwK/xQV2dgrAj72i2Hg/NWO/7KHfUYDmn9rCzKjn+mWLD2Jy3sUbuMy1uLpXZ4oAtXWNfYU5j
RCysL0ezX7t32Kz9Ti8+5ongX6MxrIEuhVlfvitg5KCnXps6Ne3txxDlOyZAZX7Jgx6q9UfTNdOP
YG/yvrd+dKNM125nWUbUrI8GFuBxF2UNu+edgR9jSTyp9g+j9RvA7x7PyAUBQWcU5MVzFNTYROma
gOkbt3OgGr4iSlO4LRVMrBEF/sRXMTUv6scqMI689yxoNACIjXyHmL05eVsdGl3uaUOkgewHgNCl
Bta4r+ujRh0mC50O/5y6ARVlRV7ZXpK93rw0EM8KUr0j+WxvvgvFfbIaqtDL3/Q6gHYMGl58GUKN
RZmYvbbnujos3T9VhjeVc0dxuARPOLik/yp2C5f8l5eRBN8XVBJNcEeFqWQuR7lYi+rUZ8jrKehB
HZBQ6DlA675/hkPUomoOE405j647AUveQu7wVgsfSftA8MGgR9/3nbLOkNrIbxJxmdcYN4aQ7FTC
7X01u1ciSSJ2GksvRkF2rBp1mIhATuTRdGW4RYQT2hPWBCtCdb+fzOta8j3d3nz+A3hcOtkQwcLF
zmppYtnRCuCsi1NGp0fPWvz2+4KjocCEerahY20+6WfTgDTmz11VobGWTrAGG6KvfxSZzbvBtrz8
nhWuDYvoV4J1mIBT+vBLaNiIN2GwMh1zLVfQBcFr00Rb8C1WukSuedh8P8BhIX/7kV7kLsU4QJCL
s/q9sisjBdDrgtuLBFgbc0YCh5dphLfmP/rppVYLo8/qlty/n77BgF59FnUwZtIhhEg3Z/mix6iP
uXXiijMr6tJUc/ZaMi/0KZK9DyIvr5zUNKtIkT2XOHD2I0Ajf213kd74aKKBf852w9fe6ts4Hjor
AsGFUVtRlmjruKoeD/p/W3o2T0jjEzpj/Mkg2WpBrAzPXe3Ygvl3U+6Pm35T8YuW2EIGf8HBZOcc
/zQfa8OBqC8WJ4AqDexdO9cmIMJuaoU6gwV32X7prNcqj16n+EwN//2+p1quOrnLO1ZqqGN3fTrd
6/NDeqaYPZ1PO8IHULmWmOUr+xKCKP671sJ0bMIDMnquqBCM0AtAjJdAkxtELspEincF0Hl9Rcur
seM8nzcGWxaNtcsmzHJ9lHoSpSU0tFzwxCEjt4GMDDRlfjem9y2BTMihHY2t3frMTi4iTgCdTiN+
K9mVHIKq5UMKfWWyQ82cYrXMz7TFYACuIxW14OPXN/4ZoPYH7GKCZ+MvpawN0aF9pyLI0uNboSsY
ABL7OB4zrC0tUm0Oc7I40DNtYSVMfZ+DuQ9zeDeQoIPdNs7rRpJebtkPm/zXAzRmuus/PnPgLfMt
iH/bNRMdpTDRSjy8hwvbbdwOGE3Eq/odkkCzbokHWUkF+Uc5qwNJ1q56vY7btH7AHL6eRP1B6Z9Y
A57LhieqsXx7XnbpvIlALWzaQjKV+3q8QxJhKAakf2Cw5UQQgA7Ga1GzXGq5+PpgT2LUkix6qdnU
WXIjI0f3XERXkQmQgODzvG1UTIH+GQfaC5DASGKuuVjFxZxUFz2pidgQsso4whFcrtmBkafoXnhm
T/EUEl0LvfdBsRaLNszu6oeljmoX9L5VJjvz4h/D0FyNVs2Y1XvhsTZsLWoD7WMbufi/V8HNgxEO
28M2XJN/eQ0aOEKFtH82rtc9U9YajLjVovgcvwGHYbvZPmfljqvevrkMFA6yNS/x2CGW14zQYsAP
Prwju9cf1UmU3BYjWaRxCrWskFbXdA3GnJ5rXMFsRHLVw8H/Yxmvu2/d4LzcYxr5Hghlqm1puMHZ
j56e0WK+wEXk50l+ZaCqXzJhfbmdYP++pjyts00cETz4Kc4HXW7S6dOxVlqmJdzuprCOj+KL6Ygv
FiX75UZTSYGNT5Z4A5bXkMd7gfqgo9YocRAVWs/VlMGEyA87KkGaVFUDjerggCHHSlsAb0AAJoA1
PC2+GFxxvHFVR7E3nKKkWYxiw/gI0z9wfUkDblKiWQXDyA/iG4/hDSDpO7PykzD+gNsXFtSVuz+s
tth3tucBzLfS9AcKR/Ozp8o3mtXux429Ce5KSDVkEMccjm/jzA3fWeiN4EqgGoPjx/GRGcOBR+aT
0jnVn32KgDG2xD1rH/i3NsM6e29zpnAkuiZ5rZ5J5pe9rIdn/EYKkovnMrgfjYslNRlHypdGvn3e
XxDvxarO47MAuQEFP49whtqNk9Ctzqlnc58TdOIftSvTSPcygsKscNVPzy/H85ScStJeJPbWYaQ2
Ki/E+8q0UDatJQ++yMofuFu/mCEvNJMe3xnklsjY3/97N25SckyP5aPL5whNjSavA5wVgjH5e4NU
b2zqN68doevkeO8ERS7zPaB881++3+WEO/3GLKdxN1rBJBwx5Al6Y556RWs63yCXyOAP6gW9S30E
npVwUVwIGpvYeCc9yHsN/2dXD1KgDE6b6h7dE3vialYHSiCH35/GSYSXYVTU+PlcQxFyRfzXjROZ
nQ2Azu8W1elhzkQ9qdxIuSgVSOZx+MjgrVrWt1oae1eC4IkNQri1naLj5H5GV5h5a68A1eotXHT0
1vucIemJ7+EFfZEWTS99vbKqiKY5TJiJCf62Unbwh4RDqk9Mngby5534xI/YNWfMUk/88LCj6/Jz
zuo1lLAtDKiJPB27GFxDO6XcXTk+09TcHgI94/q8M1JS7m9TlR/3DJWmqgLPmy9dfRQfmOeNpXtI
YmfozOKyLfGm6kt7wXfsFRFH7CYRS56Ayfiz8kBK1N2TE0C/v+s9uF6NwAanLFViNuUJmzgsT+KD
zryGTo5zwsTdxM9lPbFEYZTO2VBOjrNNsuNfZfXQjpRkOYgO/p74ObU2SzYunhT/21XlAj3+hW2X
9FmHfytjTW4ltTTu3uu/tMQ7ud1cALt/E8AElGZ0ruukAI3S+PWYdkDaGCCi/0cMbutRlbtUBdrU
NyiQXfpNxjJilanJ3tVRY2n6zViRSS1BNmkQZyqFXmy6Q48rZ4gzNgjy1iAm8A0GFitSCCgBR40W
CSoF78i9UUiZCoyLk7iG6sbq7OmX3XNNEjNIqlKkD22hQX+fhMEPrjmDyBiHj8zRpLl8irWJkISQ
zRVWwtNSZZdOt+m4P1cwsODbJvjJJZu//2rD2VrqLziMbe0H1ejHNGaspmm/Z5Lp/Pfi2+2gk41Z
PdgU6I61k1xXQs8gmEDpX3WChZ6veapwgOLxNqxvXwZt46Z/osWe9XQFhw0vheRUXEwaVmnsUmSv
w5LVX3HQXHcUR0wgzAfAMX45FQ2nWGGe+aRoRdvinnsvVcr6zgM4EbhT4vnMruQaiplp6+QoyeU5
/skyBYrlXHtOPWu6zECrf+2V4bk+Q47YnKJuLw8QDXwEOfuISpu9mG8QwmjxqrivE9hUgTNHYHS0
c/3TjmFY0nZQiXwCaKQqVtOQ7tldGyF+xLHPHk3iLbun3/qWq4K3KZ2/b/cqTBXJhlsQ2vM+dVVM
vMMN3QQT5GIqY+hZIP0hDB1xnUoUeIZsYiAkJZmvdWst/hrW7rEfMpDnmQk/yDqWLnmxW2BvsYdT
XZ/lZ8ZR52lKgcXFHl6TtTvX0WYXas7B9w3u/tFlquDi6lKJJklUrCalBf+XR5+Ci7Bpft2GFRQt
GPLH3HOj9GetxuxIHn35Qpcq7p6dpc9T9AQeG/rYiBUE0Iz/YH6ScDXHjTLlFcoR0+5p4sm9y7+L
oAbQdeLd8Lj3qESGBzE+b8GotakOSSwOmwCgF9ehPeMaQ7oe5iA/P7xXrU9YJXy2co/CBlVyGEJ+
VWXFULzF0yT1Bua2VzP6j7cOaX9Zh8UfVMrn3SV+PvhYEaI6Nfk21HbFDejcK+Q8Ylk6SKrDm6ok
ruBf3RYCTQT7wiMHycB1OWl7HcaHzq5njDOXasoodm68N6rKhLC5re/jPmf21WiolMGircWKh5mf
X46vmc4iDouy4/RMHpkpuFiSqy90thTnKXNYvZ8bTN/xZqh6xtJ3944SqILK6VNClt5kuO5I0Pha
42cHWB6lO2aFOhSyxIbdC1M6/lwcFJfTCKKG0zHLTl1uEmRtU5Z5vurUwxrWxAcDWHA4EEKb1R2R
ZIfMEd9DiEAGansICpI+fU15heaRRDKuE6etheueJGwTYBYHlaM/Ho/ZfaFJKsIFMvIIuYOJDwJp
mlbFPMpy7QCRk4/S6ogQ+4BGn/JaQaf/hwr8GsJzvc2tKgWEyo1mJB+sYa6iyHh/taGWQXhl9ddx
BTac5vMu/JYlEGiyY7af1DJPzsEw1Pe01PGm8xqYcRhUe4GmiRwhnXE0JooPfMuHTlgPez8DU29w
B5a+0uQS1WztG5yoy7e3fyI2Asxpku31zS6mW6ydtbo/ubODd3mBTCzVGBlDPo6RfelE4I1ty6uo
Fg/CP2H/dqCyNw/bBgV+oM9bl0WBYv3OoLxm8YlLIQp6oi20zjOIZbrlC3MeiyRKjPouiDIM5mHT
lyK488EBsjkj0zheywHToBh85gKR+FVp0YMQdW1DLRTJHT9+3MeaY3Wy/RgQxH7GLOhXrF+jO6Hf
8NsQQDNXEX0IXA6/a1IAYgBSrc/vf6hnw1MtiB+j/gfQ8luT1fACgUxhMEi00gmqKErrAwOnqsvq
XWpJXZSU35LxDB+HLcj9xOALsDy8UqnO7BoJiK4MIcbVLOKPUNJ5YeaL2XrPc77uBv/dptqpvB0u
BJlmgCVkzBC9O5XH77q+beXC7DOonEK8sQLNec1RdoLpH3PW3oX6LxQ539Wi+TFz1SSqFyK/iX1g
+KMK5m6AYXBhRppetEwaEdoFQGwKWK0u1Vd2SZllld6czubqhRiH8lytSa/PEuPhHyzQZPbPMBEL
K805l4R3CptKMKCZvNyNSsHEBOH+0gCHc0LhInXoVCXicmtGjXF8t2HyAnpKxfPw5/+1I8zCTd+s
bwPkbA9RORvxvkZS+CNoImzDf4G69UTmIT68R9rdbLk7U92Bs2jEEmE1FloRnwtRAyjochVj3LhT
XtEX6lkIpJj3ipVRJsUSNss3OtR1fvnq9MKGVNgScXrlUvcxoxoMtwkBn7GTDo7lkHb5P6ctp2yD
GLjEG36Z5/yc9p4l2+/0Az0+yxdI5BlMTCxoK2UQ/FmHJ7NpIjqUk+xhYZtDdxLQ6p5wLwJHw7h1
nWqRV6IpuIoMeLSFmE0JnEGQF6hAu3LL1wrcCdx62xYecckJZvcjF6IGrL0OGw7PX8w6E/D8nsC9
g9Rs3cWZ+f0l19fuM/trKOIsUOPoc/IjQr1IGeoMSXNA2tqb7qfnsJETjuN4jTFvkDdg3qCn1pgL
LfKocdtRypbTJVJP4eD/2die/zYY8Cd/kA1UCTYtSuf3uob2y+yx62Mwk1RsQOc++RcGmwuIw0tS
SYrSIDAb433O4TmxSqZAz2D2xPvhAgPuYwDCIQC4SDVIKcMF7HxR6Vmhu4pjDJVEKnrniJLne6Zr
k15dRA+nojxWWQZBZ1sjFRX+LMSeUKot02JZ1MbY/iPX3Tg9VIkwFsAiFLUyqUQfBB/HX+wCphBP
9X5EGoZXuvE4aQv/v8l9W9CyhEsI7+GFGl24p59dsaWFD1KV+1IrySiJTZsPXHhgwSDEPai28gd3
BZIVyaFqS/E8G1EK7OiQ9m1DG30ES1w2kfNIxHXHAroKE7oAbJUCZY+OzEE/7ofHmUWqnTYnbNjs
ItoxOJVyWbicvPXIXdDLc70JXhoe3lOgQ2h0PNQM5W+WRCg7BELMWFfgCU47M+ksVKt2zoJQ83iz
H9dtnqN9pHBPMypTtW/Oq947wSDwI8B/p7/++SVHh8TqqCDiDBqDkaidLCs0KiNRQThVlegnKj52
Mz2qNprqZc92v1yPCW9fRjW4ZaCaU0fULr+jcrZ5Tkteu1lh7JJy7pE3EnE9S4kVr+iLIX9Sr0br
a2xXTS+YJV5MvcfvUe8V0TV24vksBTb6cz6wOCVfQtGs4XcrC9B0Znug0f/FuNWKLNQc946jqoew
DWlpk5FrcS0KgVCrKmjjMQymqRSUIAg2sao2e/SupqVLdF0QvgdkPi4Vc+Q9tdB7BpKQTrf/r47M
sAmjXz3UvGlDqfJluuXbmUxoXlYszZYnkclrE24BfggxgZsKknB7x860+qoSNoOlK87GN52TMLS1
t0ltCu/BuK+NILL55Rl5zsYbOjsMoxu+JBchcefWdXCW61AMsdTTOo19HCd4+r3rqS8hwwAGl+Fr
FLTZjRlFX2PR2RbXV3JyPpltdiCg1+fsh5hFuMFmTkfMQe2o1GzPwtlhn4S0TWrE66Z6h2xCvR7S
kAT+o3P19Np9rW+4It+XNEtZHXuTmnGCIefoKnJCTLVnpeiINEu3C0BKdGP1RsO+O8LVwdCm0RDL
KdhNikXESL4ajhwmjBBV3n0kc6EscyyCbV+ngZaKjXBHcZzqkhqXzpBKqnjr40ZzCuTFWyDn8TRr
niTsoP4TQ5O2kc75CaWY2UVPxyw3K+CDq0mYVQhId7Eh0a0F1SkpEXMb5Yoxjw3vZSQL/n33oaS4
m4Hlw0bDY6tB8KavVMomFN0eBgDOtw9DUxBSaUxVKf8Jzo+GOCi4TQbV17/7uRNrXm4R3sFhili3
TpJhdpiQCAHBRn9+CVhvf8u28zC5S0Y+77dlpDWTdH4uBmDKBveQzj+D0fsRDdEd0GrTy0ADCwQd
2wis+z0+agXDKlcdf6ibhe+ZgefExzPQJAKqRizpLvBhJI1HssHJ33M1TlrBuClxw7HRHE1lBeDn
c0uCkJjUH5oEJ1At2CpIdT0df/Iz7ahaX7By2iUeuvfUCXKHeWlW1IvL6WIu23ALiY4DegeOaXhM
XYegcdmMdUgr3Rs0YFwe/jAMIPtVSd9G6wrkg4L6GIz3suePMMTAgMGyap1pnM/Iwm5niGwFrPZM
wi5+dWAoI+qoLcBhBOYVxdBDUhcJFloKJXcs9U+vB4zIonIRBMPFe2re7kV9dbP/ykhU5HWNhBfy
+tKD8HGICbve5GSV0zqPi1zexVoU8G25poHTm+KhIRPdFFiN8inXHl8i3LxgDVgxjPdJ8qFZxW0n
/eM2FerOegVAZB9PAmVM21STIp+ob0W60NmCOnIKhChMFjuUaqafEl+a+nO4L/n+5avUyZfmC8u6
NRmRtS/KdsDgojgo/STdX74IgmiTvaRIi7Rsag8IkQxkxuTDHwnSBT0GVk4OuUpFWtJiejkTnyuD
lrtI2ZnxszsDLTpA51T12CjzJUG4y0tbfaHcao4++wFUcMz7zg5F9kqMEBn0APwIVVR74T9G6Dia
LWIj00SvKJi95zBr8FJqF3fVd1sfgUrMcETN4u6NQVbKxkCvYQJGz6uvzyIzUpyzt354qsykqzMs
laBdqmDNhENl1gvwE9utkd2KDTVEAHNOaI/LYh6sGhzLSFAjw5YDvXLdQmJJKfgwBU0iBRT5B7fg
rWZQ24q9QsMA3awkryiIWGv9DAQVpC+BZPQsePylVnsMqCzV4mu1bhC3nImB1xUJzjW1MDze8/sa
Ta0TA9st/w1AF8dTjO32yiPsh/3HHWGVtm9c0VGSdyZLoVqaDn+sQ2f9Gc6EI+LT5/csVYNh0u0O
b0zSmT7Mk+ldIQ3pZl7Y9wGbssCTKmmKnTpjBakqdEflT8CKIr1td94Dtq7CaPvyY/xqEbKOnrn9
0XDb7sVzYUpZxrxABACEIWz0pNKdUAHdDckZq/Bx0b4aZHTrHIFmPro4kLimAgdU7LuTvUzr9rLU
tB6TvHBqQCZGF4gCuOZF5HfDF6YDVT1+CuNmkgeE7xej9Wt9p86gcjDVv0djk/CA+ZtQzKdSpNS1
aksqUss7MGm2jppSNvfGm0CFIC6+D+N9MTdg3E8vi/ErlCCLpYm3FiVvp1s2FoQ9xxvV4vbivguN
GEQ2zYybx+Lsm9GTCPGicFQ2n0O1Ana1xvwGCrduz6IcZV34bZnbqFCB+b0ZlBxvF8oypZTZopPN
iRY8TNsLaXGeeyckqApDuNMzHynS7uSGyyauh0UZCDGkOldyghn7bJfPuTjTPflHrNq/DuwM+48V
7mkoDyArPdaQU5Ed8M4YJRYfAk6AiXLVjbdHcDNBQZjpdmpdUYea4mJ7Vtr2PDaXrQdO+6B6Lcor
Bt6Cpoa4OYUqKKvX65D6+Ehb3RVYsBbKrFLqOTAwWWncaW25LDU4XDg3fC8CElOPmqck3+vHCZX6
rtYVHUT1qLBhcKHhnProqd8O7Nmx6+piF6wftCrEfp5ZsNyHh3Qp78YkeNP9NA90q6VzUHQAUoMg
EsJCzuQ85xdgkkONV832WrTWccGR6rNYHfA618rWcvQXXj0vkYZFhfUU8SMWQDXjCxmiOOxCCO4Q
AnBZErByJfTScfzPKud9+RAp1bcCB1lUvt5WwqOvuhJMjLYyXPhL0RSMLHpPXpE8npuNF1P+vouB
hfjMvUJPtmsrvN7NVQ6rEKIjr7+WJa8n9sSQUy9Rta3kNGdNpU/ypSZeKrUokuySkzisO9qglY7G
Q5hjlF/wtly7hXQnICPY1O2XS2g+HBH4vR/RPsjMhTAZMHaC8LPjvWFZkMbWg9fRJ4KUG4UoUut2
tY1Ai0kQdxnD/ZK9U4/elFzfnTdH1nQEwreqt3o02czyinjh2o4nVxn0ARVOuQq86mf1xhV65E/D
y4onOYOuy9deyiZZ4prjxUHb1f/G3z1i4uWfDcoi1LSrTgpHE18Jb3V64dLHPuXJKOHnkGVdpzFx
e3ZF2b/ngvP9FVl0U+0Cs4QAqbaguyeAfvoOAizExLzFADiXWFUCiUooEXDQwtbR6DN0y+Qo1oMF
QmoENjcNXS7vQfM2SWcusHMUZBiJZB34PbjuLqO7eH9hCvtb285IMQKexZTfgZNZyWX9qaf9V6PT
BAW410OZ57dmr36YuwuGBlybL2VwRsZMJbNahdMhDWGObtux+kK4VEY8uEaLQXe6yrz94wHylvS+
nGakJc1XJ6fGa2Vzg4hPpdsqLOQ8O7nt9lQInX/mLg1stnCkqLbq/Wu/rswubcsfOvyir8HXYEuR
m+PhuKjsaGh8MX0dJSxyyUYv7/ke/I+yzx8Q0rg5Z4vNcOvfrSfnnXnEuMKPSxsMN7fWGQ/S9xG2
Zsxeo/CkJq2nmqqTrw20hQDCthfReuJcu2ZeJuuBEggwVvbLM0PDfU5j9cw8Vu8mMn1StKFlnxgt
1Hc5BZ0l/1B/Ky2XCB+umFRQI244Cl75q3zDt35agIKwM99jnvqpl51vhf9xbU725oVIty/Sbhfs
EyzMGfxcp1jA9GRIKCyV9j89G7CgW9AwE7JLEqS5S+4kuF9zmF7TK7rLu8ry8nMdW57dCJQ+JwAV
i6kSpah+B6UFlE8/3cJj4q+XyME9XiUxou9Ih3+nZxRBxd6UzZzrPM/nHjynAxg8q0Q+lgIEA7mt
xfPpaNjtllsA3lHUn65/Drt1LhQpFYXqHVFY5CVY8FWHWranLC8RViO4wPBX783Z5NWcn96B7mHB
G1xw5j/4Sp5reTPEg6I2HNHvML45LwV+32Pwq1gmqfZR1zJqDcljQrj/hKQwThHuenMRjYI4Hi6C
qGGy1x1sCrB7caDXEa8SJt8D5D0hLigsUdUfhAELAzamc5EHa3DkiaYWQLK1TShByz302Ih2MIHh
+SUmIxp8gBjxFFJoxLnja+Hzh85ZPLW0+58l0hKYMi9OWJCvh0Ae7e79t2O2Cd5TPRWt5EYCGL8r
xAZfVSoybBzlU+WLyGvRxoWb9Z5/0egq4IIGNOuDZzCE7mKrfQy+JJr2BAfnsT2Bu04wc/hOQRKc
MEpV7BEfbpai9gnHKJrOG/SuuH1NDKcJR46yY6ig3cWNi8Carv4t7FNfGUR8I6rO63WHRjN+cVrx
xeczsKZ6X+bo5p28gg9EYDV6lfKJ0mjfARdn8IiciQhvgV4czIVtoxOXIdC5REhELT0+VIHGjWJj
D/e+4kXD3C85hXfAhoYXEXsdO3NOBsvGgG4mBBwii4DAqXDukXKPpHkPDuax8L8TYObFCrfoarUu
yE1JGbqMSuQAxSoSqAC+iq3NMiXyfrCfb7ADn09B4e05BPe2bp3KkqayYjvFyruOwl2PjSEmb+V9
kL8HmM7SUemcnIZhEkZ4y8ECkmrpVJ7goowlr6M2/ljphqhCxKdFmbSnbmC5nmGxKkjdxL06dV9B
ZJeYlb1UeXAzqTSiF44+NcwK96GNmvjE/s00FnJlzUp+3azcb1jpv0Ac0etFexAXKUfafmNbsYxQ
jZfxRrz7BCN4oxHNJOkN5BjpsJf2TSw5rMupK5Nb7Gj7gQ8gcAKIj9oEsFLifCyAq+J0Q0gkmaQD
Cx8RQv0sk7E0YZG4Mv8Uwo6WIC9KiyEldVq9jrk3SRA/55uxT4I9HSCZptBjOY2/H/R0oSCkUhsa
HwneSJMnKHaOVTyjC3VkP/ZxvKxYiqEMFxhYg8rJjCUrCMPVr3yzrjlQGgnciQ05Ee50OmoM+By5
qP7jMHRGDJEpkZq40kYJYnSxiYwRysCeTrxq9ccZZ/edIB165lJFxUGuGphl7/NvcUlRQ7s0w5Cg
VdC+q5c6oT/0UTLzr997JVtuZvqLjS5NR5P9ud46SW9ey7pRGU4D5tGdh9HEXXFK5jycmp2p/fcb
mGyDq9/OheiKYU+aVrGh+HWkDttgUMmgnIFZ/xddo7pg1Q7rXOE7Rn/17fqs+r7dbEmesQLLSrEX
rl6QVWgB13MqvmUzeFq5cxG7ZeG2Yv75pOddlAPvF7rjPs6Y6xXI9bAXqtgoz7M0lT4CBjpRyzgT
kE5pvkIE/yYdE0VyJpwzRPp3xtN+EO8B5S/HbqZBJCwud6twgqK/NGWOv6gYvNU7tcgkdOTLRLsu
aUj3TdFrb6OMC5a6H6TjqpVT+wnDQvqO/HgIv7LyeqZK0Uww45xKdeG87h1TxTipcBy+RAvtkOi8
9NYw44be5u6HZoO3SwrQkNek3BXSD+7eabIlxqpHQ8at32v104tb4jAkQIn21KwA8BLaVBM4iNhU
f9olCTBNEOw3Hq+sHxLP5GccID7tOaeaK5Nq+jx/mIRHJ7BcvozfJgRVTA7BfBysxI7tLQ0RwgqO
q+/eOhhQpU2M+h9b6kUcaoar+QYDWJUzrO2Fs06mGf3iuK8yRY/ZZT/pF8sCxc5LRvAc6AlONSgQ
1ke/4MwJigwF5l00j8DGkUqUnmYXUx1EZnwEO/lFGIq+nxpXJXr/8C4MNntz2XIP9DlmyXCywwT+
/rJcXwZVgw6Y/dzow3ZbZRsbgoPdqZwQ0GeZ7SpoKThZm7KCM8hwpCmtOt6ffiF9xy0HXQ5cGZQE
YTUtKfT5OAvEx3BQNvTd3JNMwHnl9T4bupcZ8BsJ9yp5zxfg1leG1Lc1P+sjDDABwbBnxsI9Nj2y
xqNWLVi42vlfi/1Q+tQaOgJU4kPRwa23RzN0Xlss/omRxpTmx6CdAX7UCj6ptp3mCkU1UVPqK9Sv
KTCsCf3h1myRASjlkqyjZjpwAsEByXHckRO0HWHo6dZJSFiCqfhUscC2iUh5inTywPdFUUqgHq6o
Fjr473XaxCmnwyABSdwGevB5qGtMd72K/lXHyUnUOd515P6vF+zDe51jFmsxGmOV/QGmtZDGFl0v
NnrXxKdR4prsTYv1o9yZ2UeRQfiWWPuq+/KFr/reWfrIjPxKYismXRXOSw3Wd3N9p0+8j/MNqv5m
W7L9mRmx7PTOf3hgG+/hAIzcxWbrUH6BkpD3mP2Cyq/xTnq3XnX/ECrcSJxTMHc1Lp8nZ/0CZExy
IArymxm3fxb++LQgZcEFx76xUZM9156qY4kuL0T79KuXmdBzBsPKpNpkvHMnShc+tZ+yCXA9HvXi
BXlFGrXd6we1y0MGaw8SXSXwd0vYfk5eudQHfRiWhtdzRsUzRjpnpd8zCO2gb5OpwwNH6Fzy9KTa
AgExYqfvLsJTR3iLdH4nFflSo2WgS4L5HWY+Hv8oCe35201Y+aKg9cU6/695KkPgJBTo9MXqhw8W
RJQEqB7txTSblrc7zd2x0oDrtv+0XCYpo4Wmh4/rx4Xsepk/ptwoflIA9+wOcSpx7P+n2bDCrGDU
C40kgF+zY0wqa6qPrZx/nDzDv4Xb1UntFBkJY4EUj1z1F5wf5F2HBMmQkS9+cy9d1N8FEtDpDCDg
weueWEOVuo0oJ7s8Me7W3ysJpJFyHO2UMNNMsvRrmUSo0vCcQrmrXx1JiVriDdJ1F4nJIPV0VFQF
1ReAMGC8Bezwood7a0AaYoMm0JKPjJf/cpdgp/1ULsHXgvQOZS6AOQ+Y9ikEdcFfZhAKFwED6BJu
n9j8uNlI9mT2YrjYB7Kv0+WQuV4hsvYPZs8ZNKiH+TR7NKQQ5wZbbecIE2QgxK1ptvmKSm/Hw7bz
/CuezWz0OfmGzziZHbSMDrUmt5zgTRN2erukdGFH7Li1GBHbtzauyPHOqNJcEOZYnxhr5lQGufym
pysZ+vSIIoO0OAujYEFYk8HETqReaajdWfWjHcSGuIzl2R5vGh4feR3GDo+51DbccUSY1xF0HU94
p2Ps6WtkGlRyt4KQH/CH9tY29bhnwu6ePO+5RYFoeSjf65kIYclrbBRZCtASHhxES+X567riY/N9
mE0tj/8nIDqnzrYUIEXtc9UQmha2AgO2qPNZvbycB6pB3e2mdp8PjxY6kWNrwRYa2/x0mRSdi+qn
if613lXTAPy4KHmfB0EpeM2z6FHPUmlwr1hOU+kCUoBdGKnYZqLc53ESTU2arChMzQpkRitGcRhY
jJ0ksP3DPE4z43mHLiDWF/1xoukRGKk4DAmxURYDdCNRw2dwO4vOHdO02Z05sVwcakr0qHwqUQ4J
gUBvRO1bmtrcZdjE9EOWnUhq+tl/DC8T2h/EaHuUw0uzj5Zm3Xblc3dTgm/C2D5kifKLbwYmoxB7
lyvSscnWcC6QW97W0Rut5yBjHkS3wkV2qB+b2PRcZ+FYAkb+ZWTPyE4I+oP27czYOHmt/C+GgEP+
VLl5NomolxchAGM/fvY6+qGiDooRMdj/cBUB/3XFGhrUOjLpdfYnX5tF8PSjqMbE1B1iHREAKgQl
zrjBR8Tet2ad1siKdwIYMZkB8xrb6DOV3smB1SL2d6mzS2j0vtdDl4kLmIC04btzEJxySHnRhbga
WYE3YYA9LdPR3xDcvr5dcNpEIL/1BrPIgT7mYfTwFXb09IfGI1at7Wnzb4tIJC9HbdO6YvJ7z0hb
oi3lGh6PHjT2lMeOk7MZTiaiEWrtvfbkadZsWsQAMMWafXKeeYg8p2r4ejQ1SmO5q/Pvalmm3Dob
V7B8hu8XvGDHNUbbPIbFM6a2CYrZ0+X11l9Nz9c1gxQF1qvrNxWUr+S6qJsP43EokNVx6yoXR0Wn
HD1hkV15NJZx5na3uZnUeqK7yFpTU4bv+rUL7zFyWM5/J/+C32XHo3rYGO3Uec1BBQZbgCYLe6Hf
JSvvz8t6dngwAdGGJL7A099qoBpv0+0MiAcvYJm2JLu773LlliCRZr7PDrvUJzauVP1TYKxhHyeO
14gbQClXpRwWNSygT8lWpXgxg5yLSBslaBdS3/dxRfxPn1wXQNwo8ZilYdfJaUkSuLPii23N+PPU
BefCZSNpM5dqqdVzxryXPS8jTsLJXljRQdzB3pXlbxzxtmLnyVzKRsVNXDyht4tIT5smFU+834pF
7ZfkxoAz1dYSqr47dRPZobjD47VlWyT6NI2IcNjTltAIZ6aHUg8EXjf3NvH3n5xxlAIip/81iGhv
9wkAo8O7OJm6WByODLztUAu0yNt/93dC14igQFbsWbRCGf5scedqmejwNI+ysJbzRzjhFfpa5Mqn
FV4JLCTZh3GXUT7agUJ0d0wr5xoDpuCpGSnazWNduGue/Ve/IQ59kI9I9oCdeOejP2rBohtA2nKQ
+ZL2U9dJrGbQEKKeQjaP1mzxV+Cp6mvROE/K4bEXAOqUipkTYp3MrX8DZHODX2RzQ/g0L2kz+Eyh
Gn+nYAufVnplJg0bRRn37AV+dimDChTcQ2Q4aTtaSv89BtyadMuwVYae9l876wz7OFAJ7mIHxXOD
oi/XEtepdYybjuk2gmYPK4C30S6+mTle0u6j86CjHWT2eeFX+reDfz64vdbQEOJyDzAd1B3vtduU
GsTtzkUjteMOHi+EiLjrjXb0chMgrDppu9x14h2aH0Uw0rzp4Q9FdLF/WcC97aQxvkLiMOxy1e+D
Y6LrvGjjGWu8usUe/AZzjLFFYSM/fP9/G7ScMArYF3HA5xFaWZaRoJS0N1WqveNoqDXkC8le57TQ
R15lG7/OAQUgFtZguUc8nJA8Kr/h/QkG3GmsRchg9wppkRXj+nBeamUc/3120RKj3Z20NlaR4Fi3
aJam85BqeE8vI9GpK8RSeMwYS9imVyYK4Yf3578dQG4RW2AafU1J1URSkLv7/TxW6iuZSHIW+TrT
5c/Ip824jMx0Dt4QK9dymYAfegZdsqvRwuvQ2rhBw+f7CKOjYkkBqxPtorcM92iJPk5SBbktwZAf
jE6ZqymEorHqU27KJz8hMCY5Xbzs9PCZcwj8uC48ZMHe0P9kgmUkqh9+1TPhOByWsyqJMvORth+g
d0slHWC7JwEBwmFPl548egrOMtgQbfbcaw3PFJDekMwPspkXbjZ9RErjTPx1hIDEkcObyd8FKq0v
fHU3CM9l/45uSApc1H1MaTIKrAs1Eo2bmrm2JROvoMqUvFw21J40PBXQHiVGMM03s9UPIZCL0neq
3SZ8cln704sUXBIiWHNy7rOQOfePlazVnrLZFGAHtQqFkwCshwmBibjfcKcZDIhcuKwa6D3n+5r/
TJxIvjPSF8QxJlqVLA6+H9Kiikamx1lfJhRrMKwjUx6KL81OKOK16NiyehtV5pzAkdLUbKKiaMem
LDkU+HiF+u0KjDSQCvMHJvIfOVgI0I1umdI5eyrwb/rEh9Ar/LxLnwJZoSPN0QSKKkzcpjJwpgLB
5BysHVeh/RjvwINZAFlr0XN7gb8y0ELlHpoLsAI6nrQt2ASCqxK8nmsOQewb4RSicbqChOQaoufH
aNOoa5GBxrnSO6w/Obo46IrQoa1uk2wP3FjufSd2ytNhAkTHlQ8v09iQ5Fh7UOAYxvdTHrceUVZB
65+gwFuBAPpUWyb/ng8eBUOIAaal1r6+fIjE2bB30OmXGZM2rJ9Xr154Gu20lJua6+vS2yajrT1F
dRql/YZSGy7rWI/sZo45xbUJxSAPK0wToTWmSc6MwDKBcIho07ZIxH+E97HG3g0mZtG/LuslkvVT
NLKjHLQeIxFvAf3/KVLY1wlTQn/pRbXLhMSfQp5i1IopWSP8oNqMOMgr1ytVTsaYd+xOoYa7Pcs9
8f1jbaE4h7aydBueMkeGetVqrwJ67KwSAIaQGepiCZr/5baenM4yVXq0p1QOcOuJnNTWbIJwFqiF
KV+RX7rn7ZIYi0NyabJbIpRPqHRRW5uN+PjpC0lJt0Mbo9buFMt8zKKdQH0y6nR7fugNrFFkJ19d
ZS57r1Oz0mn/aJcwlIuw91BsMloCLBdYMXyI02tQJrtRoraVoW6yBgcU+Bw2ENeQO2r/7luhWVRx
KIKBViWKcizg3afMW/HDofaDVh3HzQe/ouHrq/kKCdGs0f1quzcdWdbsyRod6qCkSmQW5AF8OLYK
GmTOFjGskQOrHVGtd4F9O9vreRDKW4qpatiy/ReO+Hc4ymauvXyXCZKND6it3V7YG7Hu0IB41BGr
ETzlt/ZBy63OTzHWVuAhTUCs8BrKutv2Yj6UQmOPT++SIra5k4NB8FP9u/CjUIhuYCFsXRwOF4aV
QIkn+BWZ2Ferg4ntbDdOTVva9ivC/X46vXLzP4sVsXauMLCRUMey7rt6QoNcwGhQaubOTAzN4Zid
yVwF6C221BlIz0kUZcdSWJTnUOASQSXF3kEOnLM7zJC3IeWghT729KX1e4P/jUqO4oVMJ8ewKAQO
5C1Wa/HhcX2I0gOCr8EK7/wbuKyEbpyNii2xZAZYIuICoVckgI+bo7F1HBLBxaBM3FgYC5U4O5Qc
5Kk4jtltUmYsMSx7ciOIS36da088YJZElKabehTBpJh2wiwOm8xAYoYOVkS4ceBvOyHsyJGmnOaf
Qfo+cpTAslP0TbeerjK0ImdM7dghf0CrKyxssbP+ZSjZAE8cbnxbjD4tQDED2AXZg2wmto4zk2Ku
V60X/vr5EWz5IZLoDzL2aAlZcozEqYom6scsP8UuiGczqFJ0eGzptEDsOnYf4SzCyGwnXxTZdJRR
DwAV0xcGbzxfuNJJ3MTNqaAiVYJfWwmCuXQpR0+xHQOWbdtjYquANG6vYnrQH3iVtGUQLifn6gLD
mHON4grfy8pLdEFWwVJHdLRP85jUHRJh5GPuhSZohWlKsgE823MM8M9jKlrqSWGkUcegLCV3hly8
MgfUvj/PSeTkz4oIpSJmqGHe5TsRLA4mu+jiqMpcx2KqqE1Hh/0LvSLOFW7b27XC+V20Q+DBY3qY
iT8lanmKLEMeRcL0QaZIUXeqo3+MYY1kc7YSzO8mbO2b2SnW/a4kyz4ryyFwv7Jua2UYh84yotDR
sKITHBo7eUyaYDn7BvSDYHwl9jxwU0tDDKefVKLRewwS5ILdHqjjb2QdF4Q6aUygnNtyUnjOEqae
T56pQE9aBn0r5kwR7BclKrBge6QIYt7SFm5GOCiilfWPEDyCX1l++kxwY5IhIuv8WpRjwEOPxpqg
/LwC5gELWahspKooqHK9vZIB3eYOByIU5fHWMGR5TchqlLVMefuEiO3wYiWysdIS6A/ANkaHp5pe
vf/3T+K9nyi1ImQ2jODgV77Z93mUsXpyre2PPVVCCDPdb0z9uhYByqRIwYOKOJNqGkqeN1i8Uo7k
wyDcADvct7jk74U9YEhA/9EgpB07395wpWgPkuZ/KgW4gFEyPUn0pVsECwzsDjIEVbIJAuD5rN0c
ZAyTKfrqaiVGrU/gyYQ48xpksbUaB9D62SOQGsVTKzmBbFhmdXFdBef56k2XpaDjRIwWIK5S3kxT
Q1GSif5Pge9gzJ+YJLhcFlb+nrADHMSCfl6/XPePpQcexmTRLytJuvG6O7OY/KOrOZQwtO4CDOcT
djcOu+0rZYqzVhm0P8wL5Fei0wysamQNH8jiq/BjWBF4s9gm/h5EscDNajfeyPLm0bY0CzeYEXIC
4kT+oY5IxTBmbEA6Ui/5d/sZx+JTAQmFrs2QJ07gO8hjFnTtcMa+lNaGzkyED7Vkb1Baxn5NioJE
cXGRv06PDXyEnzFTO7Yyju9eTBsBbbV1Sh9oDyXdj+cKJI+m03CHiAWr19lRdxIDhUCknHfNgkHN
VmpJalvrRAzgnZnT5Q99h52eUMSODL7gDnYPVCKpYhy9aFUg5yWYa4VRFRsh8uaEU0m5CNa6htck
Wm84/jplB44EnPU00B++Paf90+Hm06bbOvMHrFg/KOf58FNBzeLkzqG10YW+1jfBmsRK3zCWwiwr
c5Dx65xYyNIZV4KQlOGoPbLEcp2khrCZRDqnJyG81hqhPv6UsijqEeqM1xpGNVhkIXHcxmaGgqxv
WKtn9O7clQyFxfjamkcopr/UWya+w/W/OGIP2ZrrPs0EjwOHIOGrdyoxdC4GGT+WP/knr463aMa6
7JdvThTroS/WEp7sgrmYQ9BWM4nuqUhMxFodPUwGLG/NGxaXYyFvWci5VKsMuLWkyIf2JEySPX3P
YFBmOxBRK8GJhx6IJrQdc/97696GfZyfp/Gqei1uihVrVUZCPVR9Jry6lW6Px+NjgAum+50ZiJGh
NWvgzkMIaPyLDfbWBs5aRRoVthECpRJ5qvHflwJTzqYC4ia8peLP6J1kew56kUaKJrylqxcfq6pI
hjZQJheJ6+yNvea+SfqUxbNzYUiIFdWRx0T7Ocgu9N7/Qs3Iplm4+lHwNXMwK0eu/nwKJmJGw4HN
UV0frZal9ZnweGi+rZS6LZsxEAEQzLSbYXQIP92dX0JwZOdipUba+2JlcVPtROg5acanuH1FCERL
gvqBPzEFFBkLuKA8CQm1FwUHLUhGFeevC7KHmOgw4u8aQ0OFNftZgtZSlfsl/UkXLU1QwhF6PAgZ
Qb8vCI0J+NiVbXKdKng12y51BXD7d9vtwVDXPeK+EGBS5lbr9a+WaYtf/7ZTVNSSurKjTTmYOcTE
MsahgsFgOc9QatcItCsZ6h/kkWGbbfij+UyGXptGuMPqz1rOowAA3XSqTGar+z4dnbcPia0btmbo
r+9o6CcdeWXNfJsb82qIDXIF6flpaqylmGmTOrqxEFa0gN2nU8WeJzvL7EtVtY+vJeB4MUhtPrEc
BsJ7HTH6N9n3nT7z4txy7yJ/k3wgtGFLyArotrIgQ24sshcN8dDiQhGeE7kRyFvvHhQsSA5Cbm8T
mwyAfYMjNKcE7VUdJmreasvSjoABeHezq4gwzws1M4sOXIKT3WRBkFPTIMYmBfuUJlUY764soeGP
taS9AgWI9ulOSBmrpW331P8CTC8eClo0NKNdsEJq27kuUW7OXtyaMnK0W6bL/TYvf4/8Vjk8auLp
fTzRBWHBzpkXAAlHf+4e/UotRtTQDOyUjjQJkHD0mlhUnPMXTxlca2hd4zjd+lVI+zm2VE+41vne
9g8BScR1a2oAu62yhK4Lk9Xa8JTNHlpUT8EOTbIcFW2UkqPnGTv+n7NXrN9CZboM+GuOiBg9X671
M4onUhx9cgipwz8tnCpsrVM+ZHwRO17DYJLwgiagDyaaqj1GtEmgc3x+7Cy08oSqFdywRohKQOCg
tYh6mj1UIzhpZbgAVbvNsSIECVTLTmlrvZLSrq+JOybTNyk3AnhJ3BhunqiDT/VBc3WNLNn1IYfC
CUwbuDCY8umJsIS7F7FGMtaYyJhXkdL4DcoypN7lZE7ePChUM74Br41gKMGK07bbTgFb9NwwjHDT
MWBHDoLxiDAZgQKCNSH6IlWzeFuMyhwPcHNzSxFzh8i06LQV5uR0JY+bib6quiqUh1Log1bl+GS6
VLi9JAYH6XO4wmLz4XqUXjPhZcz9plzSlVClb+uU9aZGd3pQANYBw91EqrPSFptcPW+k20q7DkEs
cDrON4a01CF3uJl2tRq1fSNdJ8B9RErPOVJnyWVoLOlahXVdm8/oiL4JfgDR9BLfpcRIHL9bftXM
NRleOB2SjgTG8VTyaUNu9jhtUyWLUQhyTGXs99yWNJ1gHDDz4g4JXSULDnAde4jo+z+gi0rZZ2Pq
jQWcqofJeJ5Wo2vZwWN3NcGwFh4cPcT+b7mo9F4AkcyCmnr4lDMSwEhwgm4jeEupu4/pcWqlnsOS
+MSxG9MWnXpz6GgFIoX1TlPEN2yGCwdRAHhVX3kFmxcGJUcLwHi3JNpCKX7HIeU3NZcdS70mzNlK
Deec+yVFSRnsBWj8mdy/s2pkn1ULKGvYTTfxIUrxIoSi+h1uGTsp7LDCOVrrhwCu4hJLb0JS7/kY
6/mnoFwmLe1pQRtdQ6fBFz9EK54uRWYjmCR0kH36Wp+jWVgYSvnSfZfakF9ZZsS3Xc0m6pr6War8
pG8PeODrwCbz278Dz+e/JNDO29AliNId3LaxpkTSF3ER4VtqLGce1UdjNBnYl6sXYx/irAyzrJod
qTH0IJ3ElPA6BRK1u8xNij1OKaBb1fL5F1Fx3swBzW5bjNXwJP5uj0ItCeyfj8+uDpzTh9PJnDmG
uW9lVSRKMwKEMIuHBJNxYIPYTnOCIztAkuw69B/BtytierBl9WaJJexlkm5JvABxnpeAjQMCIVJZ
eR8tYM/WIOkxDlgbqqE/MKptA8KIu7TW1CugKCG9iQ2CmKAoXWbUz2QcvoC9oiZXccHTFk5IHYiD
DnyLJOiTazH4tadlcOlLp5ei+1+1QuGGMsNIHTQZ1g+9kgjduC8YxBUHWynxBPs8uSSWGS2n41Cl
RqBsjmM/kRRmV4ezb3cvZNgSu4UjjMF7DSZdDDtzKkUZ/3A0J3jNrVMuKdfEiRY1jHYStx3pPgRa
iLzwBJd9hG9nEXla95itmh6O3Ep/O/vWGhe1BcUAOs8tj/yO1xlCdcXbdKVAjGeYucuTDraIll9f
ymnH+DlU7l9IUR12QD9nkmxZzZP9ftFPliqvVt2vDpwTgdkB7NPz9U7EP+VwmiOtv8wudmuEKFLq
0MTlvTBGr/a0P/f8TBeEmhYn+5iZFcOjep92Qu48G1E4s6Q0EgOENIJ+cdAZJxD575DNj6vf9iS4
r2AhyikwohNl9XwJOaA+VNhxUYoTWm3grBOmtSQ+b2KCjbxk/Lp9fp0twfmjATVwDtU1bZwW8dzk
UkI/9YoxzR97VyOlOHQLknaGQkQ0jBPxwY7IaeI/XME+3G17S6kVbCWFgSjcgw+3MKDQhfGecjB0
B+aRrMf4ixgBJCag0k2me536Uxe63yhvoZw6QM9YJv3p+ltimPHnLJ+qsevsBvZ4MiSVRXou81uM
Nr/9EYd95K07iwrEisqiqFdAJWmq3IOBD8FGdMnEaSNH58ub2FJx9kWgqqBkeWsaK9qAM9J/I4Eb
vsal4tU50nePlfVbH2p4QEntcsnKUCnJMEg+9BgqkQ2HGXqivaHzgTwSowCpJVl8yad5hdsk3Dou
vzPfmWSzKYzmK/FgM47maK2DhXQJVurptUkyDLamTPxGYWRvLMAwOyPHqM+yYDdn1dTsmOli9Hsx
199go+Hzd9l+99C3ip1CApzYs+8kBMlLH40dMzI1MLWIi1Eq7l36GXur0rHhSaA2hyh4MfYgJhws
lHSU2z1T5qLciTYbukGKoocbRiryBP1sN9vn81EGEkYTv0Mw6CwY1RCYYT0+RvxFXFrs7nuKTJzv
GOi/R0HIZYim6rOUPjX8o2Y0E5JuT8WETGtc6dtgY7MeEy9AqzglH+WI57PgzIL9XFzvzDQLOKnX
jARdMGLB/PfWWQysTpX0TWJe7Z63/+PRTASt36rhhUCkleV72JP3jAekDZBwajCU55ZRm+Wdj+lX
/SPYnebnNpKMleQqEvvP/C8cq0/O8Ql5OI8vYhFvh9KNLNQKSwdVD6N01hga2aoQr5XvPzn2aidd
2eu3geqrm1txslmjThhgnsnhELefDRKDA6VM6RuvucFDyAvc1ncQEx3K8n91xbDNdvUj4oyc3V4y
pterira4ixeH61ilm7apG8Jnh0fI2XZcOaSxiSzASPs/b11LEIK7wZckf87XALM0NpTLmce9bRBF
/Tfz65ILmujykGXcO5pMiuRjuV0+eHnfb1c8+pZRFMpyA94XvqyysqQc12JZKul3WM6FQF1xE3Ym
T/xnGvjNC13qN3cHwH6ql9tic0DDHxKG0xdVBwQr/5kWI9PzCD7iVXnqEo+Q6Gu3R0ps3X9bXRp7
3CxPcamB37rBOg33Jr2ScvzdTsqPFMXoSeowq1gqW7xZitCosa1CbDRfBD3JDWB3hTRF8qVje7wd
PVeZY9UWkGtCGOMyhXB5BQmnwbmhaWgTkDzo4E70ag0pP5Fih8uXKupZffEUFvn/9YpdQtorPfWa
jED3umHaDSrci6mKhnW9CSLZPvWjyi5/YPUNv0KeMUujvjlk/P0je7YLtDQ7eeAJsSJDpMjB547o
BNmCeYaryB7+JeNNbdw8Md9pzTvz0z1/lnxqPNBEpyXi6Z1j0Jw5sZ2AujwAutBjR1SzFHhKXlqu
P2UOEdU/H9paMmJCU1+TiP4nYDB7eiq4BV3ufDa3KEQXAkrec0GsM8s8cM1EYRx/KihVIEBsIZa2
Ca0oBi3KNrQJMZOW2FzynyKjtsncqq2jX94E1Tc9q15yx5wZyz5hXAXeV+NrradeL7KS46GjJcuI
2x/xWcFcf/MaOWGekkKLYP7x4VpiI0dYfk63K+zH7l6aNg9XU9ubkZwXIWV+W70j8j8a9bIIdzPp
Zm2y6uPms9XnA4hE+oegU4dZQbO3jyQ0BMBkptSdJI3EORnA7UkQtuFugNQSXvK6KNPkAEEZoGA8
1bFS5sSHZMTqMxZTeL3LXGdZsSD27UK+8CH6SGKDHNuOo4C2o26EehZK2GE71qAn3MiwJA79MFhG
LaBXa9YGbEiNjnuLjgUsJg6Jb28GC6amloUlHFcMxjJV3tjK5NnKn8Jv5+k1qx7rjZmxDTysyQM4
AE4O+r/g5OBZfHCfG/68akGnuo7D8Yom3TpC0V4ZHLoQv/WeZMxbQECx1eH+fhdWEE4aR2P6Zhp5
cKScVxmAIex3RdovPLci+f0tYqr46PxJh4pHot5HG8NIOoGjwbPNHgzAzydC6i9zKQeuZ2e3V+rD
KbpMTCKr5EpPVCEQIv8U7IPrGVufbCGXUM8W6xN90CGAmm0gCB3aYJN14Cd+oYkr6sgv5OpUouPQ
wX1YOzTx0+iV4bGiEYIFzaVxHTPwVXRLS4rPv5DvE5h2qivY5Q2Sc6R65hDuUexAFO+lUlgRTunq
QeWZfCaVvmN+3oppKvJ3dhl6RDkEVExU3d4i5pI8XeKkkJ/3YcN+/DeZun8H1R1UzLsNHcX10jgH
Xo1bDKCYu69lqifCWnt5m6aqQtadC+0bArhERkItYVV5nfrWVAxtq9hw9Alr3+Nau09czaNqgLEH
v+PN4oJLvGlZl76EAmefSu60blmAiajSeQOUcNZELzD9ckYKiz9DC2rgALafgrD7ingwCorg0KoS
f0CmhTZGo2NforK1acQjMYFSKf+olej4Wj7yvIZ3oaZ2dNuCE76pdThyVlTfXcqCsvlSRxCTgWmx
GaRvkF9WfWvhYy1PI0GRjvagqAnAIO0HMde/M7jPWD+1h+lk0m2p2tvD/UflnKKm7TzOzIe3vg0N
VKF0CAiz8KmvdUCMasyxWt/TipdU1A03Y41B/I4DzSEOpCnSe40ujM0Q2UDd264PDhxPxSoPjPJs
O9M85VDXGvtU3t96T6hYw3VAWEcKz2jfIdoq3n7ntPpDIyP9ZkdemtMsXf/BeIXkx5bmk1F4RcaI
yTmCkCb+R9qmELeubkX5buxkXsvjNk3vMinAYBoOfmA5P6ohRHw/dxP6FnjqIjx6CfTkHzEqAgAf
z/jrinkR67rJ51y7/NRb5BGFEn/BPMvurHq9gXU7S7fZQpTvXdh8paOF/sEjIu1brXAUK1v0OC87
Sl8f0gtkSFgbCTifAWf2KjbFWVTdi4294+0uAvc+0wNHIEyaYxUbkhVJIzDBn+bGgvhZccRxTu3u
UrBOoBspJeDQNjtN6fMmOx9vQ0tXoQ+9iGQKsTe4tNHmBv8E9bxgtQfh2oCa0tpYZlnvGs6/6SaS
V3hYa2yLLZwPdgvrbLc9QBqLgfvRi6fovkuR0aJEDsLQ7veHcc1NG3N0JzumFVnGrDaKeU7gZj+I
XmZzWtH92ete9BZiumYX3nC/7NRhKeY7NgYNIRzeDU47iQmMKQSkaDXv69qZw+/y06KRE6KC6uGJ
IpW2G0hGW/H41tME/r6N3tmSt58ElpDh/5XrLShGJwSwVXjYdU6b7DpVWq25Pcd8fj1C9P8n5SMY
ayG++wSnwR16pmVJNOVTXwBYZkgUJa4WM723THgnq+Q20fJiWz1RKe+IFHOAeigjwJsbAHZqvTT/
XsEXZzs+Ukivuw4Q6JsxKNvjcz2elilT3hR5QBs0bxhSDdiL2tkSzNeQW7/Ln1HwxbgfnONWLzIF
S4cZyki43C6JEhyMHnP17ib5bh8EWKPt+7N0P244nx0T0LKStDZ7nbTqri7Yq4ywLM8t6UEsn4/f
Dzk/UzEhqTfMnNIfoUq/Zc+zp3qGDbMGGFPcYD3g7ASFooPICMUJdCg8vEi9YVC6L/wsI1XF3kH5
U/ZIdrac0iFLtcO+2GeldLfigAJp2bbIgRMjYjBZ8cO2X2QKoEELfvM7rnKzXEAVKxiMhdbb02rl
/6Wv8krcE7V/h8Wu5mImuqIi4U/Tjilarev6V+c3qOSv6isdoFgg53bAZh1/SOrk/6eUwdyybAXV
5MlT0RWeVmWSKiUH+ZkhyQGq50DUz0mTNxw2/bmpgAtWVFW6xd4kHtCAA3W3oyZNVJWnC8K56aAc
EoKf6/5D0L4YuiNpJ/zwA7rlM3KwkN+K/1mo3jRNN4wjTvIcSZks7UywYI1VAQjOlhodP2T9B+dG
luuOqiO28yunTHbbuVhz4VPdkHya7TTA2PYEbUfpoh/v31bHjcV4lZjy+AdcyjQwN6uDqnlGz9m1
GmlByTxw7qQr9mbNxrhai9Llv9iIVO0I9AurmF7HQJMiJr0l9NGXoF7hi9Ot0KY3sirzBGxC8RE2
XBdXJgqOpe+uCaoJ59k0t155tqE2HcE75foqGos+iznyvjRuocK3i1sQnpNUdP6cwFfreJbCSvpO
+McJmmzj66AHvSlwtsEE+gkv6CYKV/3mkRRj5YyjPU9Omh5lkVJHZUVg1l4Y8JTN+R/WMkDMM7k0
qbSQvnUs4oQJ7b/EElMgUmPVvIoLJutkafaPM26H7hUpIf4J/A+HEcTv/LvItl14x5iLeOLwpgG7
e87NxU+jAasO2ad5tJHhJBogb8cKYcCBQnJi+J/O3hNgBCDXEh5YEjurCM0wECesAX6zGlpLkQ7g
/IxUKzaQJkd/Uk5NX6GjOgTViTpS8I9pszCX05CFDFFxv/k0k1moBS9D5yemOxitwW43oM1E9ySf
WZakQpizxtxiPRsnhD88T+8uClowZSsoYmhC4vMaRXTFN4ND8XfpsLFIoWApJOE81/dYWBmPh4Ke
rkTVpgGmV1iWtqPEpIf0SQ9lUc+MwSHveLT/JfktAyJfbk5fc136P+46x2GdvY++1PSC5X+nilxU
QB/EvFaJjv+cDkXO6sehfCDvc79WeoM2JCZGWkO0IwvwvK79JUNMlGsL2URtKCbTR+Zpruys5/WK
t1XZciT7ldpe+BOd9/mRIaR+AotWCpURyaMvNI99UyB1bQZ5cxuR8yYfV84rFOU5kk+b7WXvk5Dc
uxqAuNO1PfIEVwUicUmnMPGXzxrMqZkRoLwe9xd2J3bpJNrm2JDj6YhGgab3hMfIpdiVFZ1dLRHH
m1VL0VOYzSYAFs2rzQqyZNdcKA/rs8MW7/RoLvNwSYx5n/bHv5AcWEORj6uMHZx9p7v5D7mLfpd7
guoXwzEMZ8gWtQx/ZGT3lv8L8bkAFIpGJqeH+NQ1MoUZGiiSeFJEn2bczms9icGTvwgoQ1DOA1qO
6QBDJevb+sPuSCis4CCFQ11S055Yvphb8khgRskFYgBUM6qFFZMzeVccOZmdZUfYlx13Lyd81fep
RUmBvobMU5tN70ZMUAnUK+rx5tOwo6VEdlmtU1ssEFeOkpstrBFLXi1Q+1H28WGVgasBh+1BnAWv
FKofSAuLZuDObbtH4D5Ss5HkOrtCBP34bNJxBNAtLQM0IUvXVcseva0T5qq72pbjT/NZy7dX7QGE
77wsLzC2n7kkQrfrba10Dj3mDcwf01ogz1nEjdY8Qjj70r7L3oMUvoPvTpsjyKiqzo4w4iHe0Kqu
AmmWCi3GzNU+Dp/fsje7GQGduB2ojL7wFeAuZorutrHe/g7zVDM3YNHT+SjdRmS2nlSUc8d270lT
TeQASMtxu7EMTkNSUX2A0QMFmL75irEfdoGQBG4ekb8FJ/9OQi2KTlPPYmYxfmBTqcbUs4yZWbPs
nOOKvdjVnkMkKFJjFHbIMoRFZdeHNLHJEWe5ViJ7npQYjQIhFBefb/VBRuVvGq/bv0ZGzjqqS+ZH
tp6byIw9dToXUvvaLPh3DvIsnyt4+pI1G9tN8MQIZefAbbZqMgMnCzTBjezDUyFGsDetiEpgK0cn
0Vk8StZqIe52UKKaZIcQTFRTIgyey+i7isEYiLbU96CeNm5Wh19xfv3TTM9W0X3aXLBgzaTR15g0
kDdoi5Gir8V8bevF+BnwfIcZm9x5hYxPd4DNi2p6y3rN5j//RKkqJ64c+d4bN1G4rxXTr0cBwjdH
nAK3PL9MA0FIgmQvDbJrxeDdvsmKGjUzBb1bIhsXeZuxt0NtqbEWxS7SaJrQEsLBf+zefCx05vKQ
GNB0L8ulUqkoJOYU3oJCW/SbM6j6Z9xPH8WDrHYhciAs4cNIH6W9uRUBPzIe7xWBod6kVhcXTs2T
RcJSJrJ9e2kD/W16+7Ivd5OvcBnMPBmyCJd7yK9gCY1k1OLikLwlJJR3Z3jwfMMJMY/8N0ioA2Bd
v9RwYPLf1Tj+PdgvoEzW4nMJxsYZ0HxTGsKQQJ9ssxJej7t4KoVTdtnTOLlfArWnob2Vn4OLFwJk
n9jklFkzoMer4CQ2gXDMuJIVJB1wtQEU1eACZ5oGFF9OfsGXI+jJBYerCAP9yx/JfVz41bEm5osu
0sUUUere2jTGi6hhqt/HZChccNHyPu8qrQ1xnyREAAMp8o/GZFKPpCkeqpV+ANWcQw0maaB9seIV
r6Ap/T+18cYGTdERb8RXQXpmFz+o8kQ4kyZnWzchmOlA57wmLL918gv3f3rvmmVCSKOX/sSgeKW0
fJAybbYM5RQWsrKeHYoqA4zuClTU5yBD6k3YDqCRko+DW7C/Ity0AB8jqgngGmImY71Z+gRG5bzs
3B6RSdpoF5VnGYs9xl9BTWYB0pa1A/+ctSOkrf+PmY7fTdMEtd5QvRV0xxnhJDPUc8y00XV2yeLQ
e1Co+az2Z75/RW7zUIA0paLDxvgF87Ajl0y57xzEG9j+LdHzrWFPLWITL8dL1zoeR68VFLbUeWdE
z0vxIA9A/38lV6VF4+JlwD2TKqyPZCzUh8o5F7Bszb9IGTKq99WQqfi/k75Y8i2uw8uRlE58GecY
JE4NAwcnPAU4xbL3jkMGW1ty+GsJbJidWNaoBVqjoGh16tlPwwOyHZ9XxWSOB4rr6bAQuH4YexL6
XzAq1qHhM0OSyQHhJZ1Tp8QBdIPnfm2tdLz74SqM8n+GOkm2FVgAF8McGjTLmgfHZt4zVXGpreWh
NDA/PLE3LJR3T2nHOgNYK8wVG1+wDexp/9E8FGv+/29mieRzEvJ9L21ws+7gz2adOWbO3RFSvOSI
qVTwH2LJgl9hFUxEVwROAegdpiwQSHcD295R4dyboa5Hkb5MRlDEgvWH2cJk3zkIT740+SYPxSDa
UgO23FSnN8G9XOGLO5qeE8/gp/Zq4PEB+Z1xXTRtvOwa5fWOYFa+fDBmyCGuM47sP5EPryiFrP6C
JzAOgwRFyzcxHtP2eca2i9TlWC8lCuJSvrSLkTm5hvFS8YqeqJvGRLcfOgjSsoqPh9/AvXQC9kAE
KU+unyygpEx7+zYkwPqV58T7SdErAR/PaEJ2xUguszHoBXr+2weZbChVZULEQRIW6umSdvhaM1JJ
qqz426ysLsdoCDjhwx1ihuj80ueu/XJt6Mzn/QPP6+d5uP3QjYgV6ZDxDPXTNqXcT8h9LsiRS6tR
36jpZeQtl0Q4m2SKwRAF37DMjjnAE0XDhfHdpIgPlDCwtqWrDBmvG8zU63FqdcqCk+ST2MdKXzAD
cnSdj4ICrEEInQ3wnwqDSPoyy32mUbPkXIjvR4t1zeZyKWPcQebCF9KPDe0eUFJ62N5rpF/g23B/
zhg4TEtgt3pFj4GnNQcbDlYfLFLbnQ7M+Qh1JfYe9zt1OIpagxIHvc5RH7goW+6V9YImZMh7/re6
zUaNeEtugnlcR1Z3NcAAtrGVSkSHHmPQIbPG5iG4KHMLrmulhWU2xZOjvqIxfHQ9MCF5T3r0EXtV
wPdCf7JJi00QQK9XB1u4tYTaKhVaS1JLs8pmjWRRD+k0yAGv6sJEPN7CB9FlvGPhSlrnUADJG+Gl
HcuFBKBNbPaayABvb5I2hZMkD4twlGoDIm9MDoF53O25zRVYn0tllzi89r/GhY+DPZwEan7wDghS
Y704P3ICqFRIE/AZo4mvwyAUMrXffXxlrBdbii3b1cctZ39+2L6mSTwNyRYwRH2YwE83PurJxABZ
NBEe3XUdTd7BMCSiTmu7zC4NQ1aJ+ZVsZ7GKTDvgwcuB8/1BDqplD+m4+lr20iLsPMY0fMLwuvVU
iiyeEJp+pZZDtAxTSgCFMphhh2IndZIvCZe7AuKAAc6hLyk/J2FTkwCUPt/nKhirKJ4jVmNTPGPx
mBlRLk0sZKxg4f5Z2XhzuTBqSxBB4hDB0aiL+480ZNRboR9kQZAudvkCgkJs/GHCsfRrU1Ak2uMC
I+Y7GK+gg16IrhzNUVHFeuXZVh/V0QsMEr9khdiD4xl8xM9635JrzeQglR9AzwgOaQpuY8hN2814
+FMKB3v9XcnTvdtm1NjVDJHHkI9lBNUdtl5yP5Ut+sS4skxWEy9oTYv8oPVWF02Y8K1P3/oV7k4L
XFa1Y715YOs3oGMaGcyaz10OwT9Xt8Keq1VyMHPjMkC9fHhAs8UO9s2qdeGjs31LTVToTzXcQCoj
aPhcYFJ4jkNPAKri3C+ZOuYs7BWuH3UfqwqM3G2qdxm/Zb83fVRLLDWn2QqYfJ4dDR9eOS4pARts
hdFSOcFLo7iV3gudu/txH6DauM51BQg8NIB8iWt6wXs/HGX7vmIjk7kvcLpnOj/HXkJx/KVfICkW
14lX9lu+ZS8IjuBoAWJdHBdN1poBEYY+46kcm++oK/joMjcQZ86pLPO6I79siWVdy3WedK2lnCgw
BKc9JI8GxETxIQPGaeJVxPeduOGN3A2ADV2H1dFspFaxqpHn9YF2TlfhFYvNRCbsg5cLrBzJKKsa
6Q+sZcG50SyoQkNgCHoN86waVobwceq4dULhr8+J0Vh74EDKjj18F1gkN9pkh6TAQQbwYxdEFpIU
M6/idMP/eRrtz2Y8ls77ewSI/7onXLN+1V9l35eQYX1lh05LPNqqMZR3tmLrBp58eRqh7XsBX1Pg
i8UZWFWdhV22a3KQ/X4dqpC0VX1QpCLDwyM+fO0RWlqrJfHqYHbTl97wFP2Y9NR7MqWPXo2kKXmR
h0Wv0dKdMvxlbXUQGeZmRIQQmap95fXod/o1w7v0yVK0x4Sgwawk9B09w1ifNs5AluGlN1uUj3E5
nii6uY/Cz3HaG5voULO+bIY/TPsbCFcf7RN2akUBqLH3x01LqP2IFM76KsT56nwdE4svXpslyGUs
9BvMOmKuQ0uKzkpFuFeKwFWy/laVdBwNMO7XopE0vUvpqLXl+yhYd7IoF0EcLYUMt9brzZVMsdNa
DRIW6+B0pF3/FFSbXMsPTOPPpIWFEbbJVBfQk3LjUqSOt2WGM4fnluMKPHuG9+5U8f4FE5ZRsPey
f9Ml64ZOr0DBg+W5nTpV3OhkgZ62TypkeXR/NdFP2xOLwtVaNDX3GaGyOwJ2cHFK8O7wKBtHrlyK
ZtlvSpxC78XKYumlwspqcpEGsGaqVMWJ1tESA0iUsoiftbzg/wDYl4Cu8WkZ0B9f7qZt1FKCpTaJ
9R3p1o+eQbA4ny7RE5rYdryENPYzHrmWjhMSC//Qv3sGLctbvkZUqvzQO608h7pejXY4myh01An9
zI6WGhYsNQwU7r0RUBzhwnYPJQq/qvZ2tqKc5fNZGaxfx26UL/a2SUZHzclEhCNHiZR062GFrgNT
TH2qaVppKEFtn1wc/oHaintRFe2HAWoK2b7FyqlXitvkDhzM0qTf0CGwpNoHyYFg23Wmp0f7EJEI
qaxuXCSUm+VliUTc3yLp8/sZ7nY77UoCcgl4M+AOI1WwG/dlQ6Pz2Apu+jRegR38k3KHAWyBsLn+
Qh4/eRagSQPqwkBlLH2JJB81k0uX4bDeeKI2Km4xRCtA6zohwMicTC5KV8505gSSm8B85Th2b0kQ
publ/qSU+YSgsfPjcKlCFXVDzWL6Dfh4SV77fpF8PAwuG2FOlIKNUFTnk6913CDC2xIHw9Qdapvb
mJS1T3LLCSHx+GAmwaK8tPkUFOoKE1lI7cPpQUxWq1uiz/Fi9ZT5gocmIaGZPIHOrYOWBboOdRZ1
afkKwht/rAWHqT82yAXiIOm4Qvjia3bYbgoEa6YyvF8OX8A8/3afGBhe/DyTK2UECxFpZ0rNjpE1
MDSzgfe6lMC0jlawq3/4hzA6I2w74R6CMywqFOYb4lfVUcttKDbVCSpv/Nd8uAdxtHiZG3tkeluM
vtBFmz9O+T+qSsP/hNVEQScEZn53BvBZLLjezyQwTdI2FHMV0l7a+fN2iID0An89vkOijqUrMVM4
XoFCgIoLSJDYyRAX4ETSy9kOAogj5PAD0aq0MUI3HluVd58skZXGKGNhXeel8y7eeaRaiXw7Etey
Xtb3LU5UXZiAwLYC4+j3z0ay8DQdMaALpwihxH81zy/mXpJLj2oqjPKeW51gRfiqo6Zant/4KOUt
bR4FKv3DgqkY/pp6K3ha6ig3G6pZNgyiFOaPo/8Ke1F7Xxfd0iS1pS3dL29iGiAz9HZL5YLcX8MN
vTTmOyoGrph3gNWf3Mgpk5GN+tAGMj+VDvOUyq434g85Ll5PF8XbK5eKYVrcTfmIGeBCXnCQ58mT
qupjj8PFU8DrA61TUY5qJaRYT7XroZ8tNHD6tiUy9nHZ4F+ibMc44GwtbZPaaJcdVmr+I7idXXQk
cAAnrXhHo8yKlAlw0oSXz23dNcQTGoUVW/cBcl2A0uivBYrL376ArROvC8+uZvtLT0qpcdhwKIRE
7xqPuYZeyxUNRZDwPwHOtOSb7v1x3J3+Yo59RtIjtplxcL0HiVCpRYIFlmR67BVFriZtSbzesDXE
bTpYXTIHLndMdugOQwvgFek3EPPigRQHl+C9/Jrpj76N/VDY8o2qkdnAJ+q3GMxnOyJrZkmXZWcP
GWXjRNu3VI7PUzelWe0zgG+RIFZMR7sdnDlk77DKOKBrqJgeAkPkmhK+BoGEeRRPXNlWenkW13Qh
b4leMekFivouFr7HncsWZGjqb3pPKeVXUQlRFxCR0eUWV6uh0Vu1t6aTsfVpi9wgv/kdqYgeZ3W7
/qOKTDmPdMb7kljxu9EAs4SsUqKnk7HdFR8CdhGNyNjI2TmpEV6ixlQqezTlErUsbI8SKCgjv5qL
W1OP1nM5XhRB8lwwZq1ftEftDCNt3J4YC75AtTtTyAedA3SuAR8LUefMBi5vYK4hBuqk0OxD0yhX
gRPH8u0hD5se5w8uCF58SskCE28rdQ3Z6C6UVj+bVWhumXXeyN5BMLwCGtQFbnj8RLlf63o45BHg
7V+FlsC/HHFKpv6XGuIg5AiZs5GRiFKDKq7RWKChQRpq5ne9gvB5LayE1exWvlcvDNIAjW7rZU0Y
0wq50htvXbo3utueMAXm3If8vh2lGtnqR2Sb7CM6mwI5Tw1Uo4ThAEkm/j4xrYwYLmgJhVyJ43Rh
+05T/lFdZJuYfhugRu61eQq2ZYDdh0fICk74bM0vlbo3N0MXN+AzdotuV3bjgh1/iG7IzglnlHGv
3KDqoXKyaaq2fRB6//N+ajf327sR5j0gjBsQrnhkwRaurKpUcrqLgGdikYEVGNxPGgrWW6qRCKXW
mY6itoYnx/+AL+REpXZPoHvHP8x7lr5NtUAwLyltXmJMZU9LCNtQd6q7h34p4U5K4eva9hT8aJpq
nM/RosBhCgFuY2sQdX4372M8HeJYGsgqZfB4onjtX7HPgGkcDUxYZ0nqV9jiQsMq5PbHpewfllf6
tmY3rdDJjXcMqi4vM1xh6+OoJ9P+vQkH6MjrVBPLetE7XZ4BWxRYatT7JWq1R80Qzttvflb9jZgR
P/o6x56oBNFYrEsigE1gHbTuf1e30iRBR6iu2d6Z67bUMfAPseBw/o1I5DOEhKgAyb7sfEajyuLO
FxaQhpllTX/Y5Z+aK5Bvv82CM4ryKOcW5eaW8iyMgJ8a/KdW8u4jpB0284xpkdsEW4JfbpTBugYf
qmb+a6vvEkjulzL7vnJ6XB3Q01pdX5uusavyFv8nLAXhn4M8kWajF4TSOFwcjWvfnwniEp0boRad
tUqZoFbeyma39B64kx5XnPErZ/Shh9640cq7RmsJVwricgwJcJMhi3HV1TZFTK5DMSnkSIqE03/j
AVETS4wrcnErAp56Sba09pSLH2nCNShU7sL9O6my+aJPXJ2NXDA+8EfJwZwzNCnhrkEXVGW5QyWN
2ScDhrCZlSbctjWmqAlNw8aRjwQ4ulxByZvLfdUusciK3aRtOMpCM3uQuLu5aBb+mzAHrw7e0Dox
/KoOyGafvDbrcPIeGyPIW+kgfyHLHafbWuFQDu/RhlfdMOLNKTPlAE6dmQ8iyNGWRj2a+extsuos
8iVjRxlxLYlsNaxZskErvE9UHRqeIDV8nJXroOVS9sMjBvk2LPMpDMYBYxtGOKCM2AT1YI88NGQd
z8uRptJU1eQYrFWcx6801IQhQaBwi5wAlOQDuwHPKJkPsuw2vDlM6N0zwCaphmXPjxuQsJR9kkl0
uccgSqJA6acPCyuWr+fITNsxSUUYzeFce7rqVlhV2zD76rZ7NkN3VY1/5nWAi+Ddc1nnesdubOYf
8VcjT77EyR3qkKrmh6dDXgP3lw+CTDXu6tmt+BadK16NCenXy8zqqWdYH+AmylSVPzgfxFx3m9z4
VGeAIrPZKmuREh4mR7OAD9I6m+xm1+g9N4GPD03/c4C/l5Hvf73U7CNHn492a/84MW9QzNw9m+XI
94s66cP9nnPLS7TTgHdD0REReZ8HTOHyrDYkRE9VGeEB0ehw/C7Of4jNW9AThKr761a07kIkyYZS
RDc24JHTq8sQJqxuYVtOKtxzPYraD1T15iuPmNw3GMTMet7nYcm96I+et2CbiKtZY5AxOz93ACVV
+LRLK9/afyL4ZdCoiriz6AABFVyL8bi08XSM89pBECEzjrMOALF5AygVtie38En4OkaKciFeobfn
SBd+4GEohrz6Oan7ahSFkNXMvykoIbzlMi3D+ou3ykfOkVyedBq93X5Fk5YoXtd7U2TuqlBgGxbc
gEZGHN79we1BqmxtwCO/AYvH9mJPb3BJwq0dzpQwjg9LeYnx7HHjoyg6hfBZn0DMEGMdlBIvQvVS
mpvZTsHplcRZX/bX+m1NHIPGyFMPrMr97nyIWmx11a2OJEAR3lvwFR7n1HAutKxLpGxfjIbN6Hzm
L0ryJ9mHTdmCd8ZvcktrHc3ZHr9u1aOFMir2cBBmAr2y7SoLp76Id7J8MGODDWcHyEIoXE7yKSWx
W7EckZnDaCvr2N0nnhcUF3FicpfnzK/a6jtQGVYWpnJ3H2JUIedOTtmDuDTsQglMFAgWAus9XGWl
k5i8cbqXdw5NovQnmR1KZ5/ux7GsyKh787H387Spv6ZFK5uKRfUA8YWDnEt2SLP9bgwdrSeo7jaj
Ba9HcbBWrgboO8gHd8QLvHLCe89xw2sTp6qMVD3AZ0tDMf5MjukSBaN5t5DVdxhFn7gJZu2Ymtlq
+PAaxCJGIQ+XomaTlkR5ymBt6+yOxQgx+WpOKJapcEZJmCw5lZ2NPZSIwg93vCyThYyGZhKo57Mm
kH+9CAuVlH7Ogs4IEFuBZbt/wIjbGzX4pF5H8s3+kjayXqEJ5nlDd7qD6Z7vdi2BIgF3qORyOhPR
3gYcegGaZn1p0w2QoBS+88j9sICeQjeqLicLiQeJXwjR9xqRllTaOe8fVCYFjQAY1FrXdEfsFGEq
yt3oorMHvc7Xk9ZoDMUtKajCj1vY6PFa1158eoDZa4ynprfYl9PVFv4mtJfwzaqEP2y/HmypUUyc
/dZ+gdEwjfddks/w5LGc6n07ENV//jfGjbY7pmRGRajlODqJATk5DdJGCN/pYGsfOTv7L68G3Fz2
zfm+3bCNeyl7DVWKRhiS0t7ToU2v7L9Glntuwkd8vQenkHMY5eUt1uT6hsf6hE0Xt2262uAG5o6f
Z9UD7lt8T4SAEpkkTIjfeeGLdxBr/W8iQzaPTW8Ua9HzvSFQ7sgVudOe5euhktwyNF6zpRgQPp9s
ezP7yXiTsNaaBp7VCbMPUxBpt9kO9FvwAaICXC6EthWIyW8Wb4fcbtcnE/MgHsPTvrUFcGF5Yrs1
geE+QbOcm8taM0+PRaW9yzCH2DTENMSF7bdSOIzyakBaBQ6gRnrXzuUKoGAwS4YV+CxB57n7N2P6
RqbPoayVk7XavU4T2papXNmm3GdQQeKuCetRPWmslc1085sYYUn2ipka4JT6G+EaSygCew4wq1PD
/qDWnB6cYKinbeSSJMLCLBWRcwBegDWN24XiqHKlzTEQiDg3q+d5mXbct1m3cOgaHwCqn5fX5rwm
9IyuqVWkkTgQHXLLuU9sv6nklo1ug9OMsg8tWCo22C2FdVtoicQDpnr6boWdSIkUraDRe9yIbu/H
CqSo5aAE7toPB+XyR30tCMLlslC3MtdQ4jhvql93zAfJU060XZmSmqgpYpOd+YC65gSlSum8azYG
4+sEcl+MuIfbjo5DHfyR3ca0TGzwT9SUNu+4E5L1c1mkBouZePwzOhVT5JnO7M7kTiix+Qzi2+8y
cj9mZ6KeOCeNTFFhn9SDwnjecI1qML3doczddGCwZ1/yz5E3FVNbqVotk/1ibEzJOjXiNbTMixUC
eKedA+aa6LHuwV5+Xfu1HX6Ftf2Dt0+7CvHgNAj1fr4UZXM7LnvrzfHbXN/xgP2dKipdpFbNK1jn
beP024mfUEoij+7SuKZTmgNma5vj2rgXVAEcL/FC3zwD2rQTTPxSxFAmd0Ermm/K+xStSSAarVCm
iuBnuWyeW/rYulIan5uCspqCNXoYWUB4fSnTZOiYUtgj4H680LA63nIiK2GZoSPToyESnJ6SAeKj
VhPriLtDJocjlpC1jkM55Ep9BVcW1xuON2Qj1SCYkxsxXvqgLz2tC1+J34BnfmtYRTyyHLFeMSq0
UeCSt2ZC00742YOEQ+2GMAoSsiPdC2SacWpkaavznJiNb1KPSSnBOKq/vkbASzAtzc8=

`protect end_protected

