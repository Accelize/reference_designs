------------------------------------------------------------------------
----
---- This file has been generated the 2021/11/22 - 15:46:18.
---- This file can be used with xilinx_sim tools.
---- This file is not synthesizable and does not target any FPGAs.
---- DRM HDK VERSION 7.0.0.0.
---- DRM VERSION 7.0.0.
----
------------------------------------------------------------------------

`protect begin_protected
`protect version=1
`protect encrypt_agent="Synplify encryptP1735.pl"
`protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinxt_2017_05", key_method="rsa"
`protect key_block
LweKQPoQX1cws2X66icOU2qX0t1yiMUqwFMhyEaZpjcS+yGZd0eG+904THRykHL6kFj6JBzmGn5z
ZSz6OodBeFpwRiRsUdz6o/s6Pr1JlXNwJpwJv/5eGrbHzy41qJ7PMQcgM2iI6uIjSBU32gVKRH7a
vipmdcmisF48bqhWGhdwtISBXO4s0h5LgF9oe3sPlqr2nOoB66ucWPpL02lNC5hyteATU/ba6Gpr
MRV+WCKsX4lriHLoBCd/g0vgzTdrmol5zx1S5pizLPThjArALHc5+sqXC+Mg4inhPpNU9xexMoKt
Ra90kZ58q4fiibV6DSf5qrTdVymTabYnJBtcwQ==

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinxt_2019_02", key_method="rsa"
`protect key_block
gOCBii9jpJal2hiUMZTpP41t/kHv6j0B0O+wYWsSJtdG3DNZfscHK6/V1wXq8vpl6SO15RUCP/yf
Dd6aelJuhtUMrl+4zmkEEiI1Fuar9SL6mACP1+WbOunO4UZItsU1xqwsjd8YspiRKnq9JbouPWX+
WLudC1ojVS84HaV7rOnL96iEM2/hwVXS9YM07qzHC3UWyz2CMYwP5cJ4fS6G4xEXHZin2nEkDjNX
WvMMFcTYhGTno/xdwYu/DU6XyAm5agc/xWbbFVos18ZqeFHVjrHWCWb3bIH8m1wEso2IoX8ftOR8
mYMUuxtTUybG2fIv9EdFI17H70LXZVjpttcb0w==

`protect encoding=(enctype="base64", line_length=76, bytes=877488)
`protect data_method="aes128-cbc"
`protect data_block
vn0tTxeXroYRXAcnK7XRzlh9xE4gRjag3b0EIxe6wPqIp0gdkmTm3z+0q0Nd0RtGVLaQeH6cCHWv
ogCVyoAijW5h/NT3WiZfbewr254x/jF7y4AjwuvwzfcpX0eED0GWThh4HAuODVYIt2GEcEtRHrFD
VZpEbLynbR5pdlp7iVX4+LKc5fIw8WnIOMAnRuAVza5McaivlcmQigyZUOUl1aAUi1iIR2XOAZ9O
2aNBl+Ma9IXAY2/gPfuDeEXEXcf8E6xz+pgnN1fddTESPPBk/jcDj76BK9rmPJWwlxLKSpd9X5d3
k6EdVE0QfZnZqvhF37NH3bIoThUThfVN4HgWTgKQFeqYsjvpwkm4TSZtDigZwG73bEZ+K26XCygm
G8fyqjkvTm5cXj+KrqJz1eFUx+u8iDEpKhV5tpaE58hUd3UB6BtyWGABWDgqgg44bdBjtTPAcuSe
5bjlniiT648j9wa7Bitdf0gFylGquwqDtb9i3a1/D0VnkMDhOWzrNThMAYP51/PVStQgw+8JO+nN
QEtP28X9UkHEvoTBpBtwfOwugPX/XKWZJvE7fve0aAhVbsb9cCU+Z2L1pWnOkoj8IxV3zRctAkvY
c/7CjAuCVsHEHLmdgxidQ2wIJV/Ha4zLotqPwpHnhaRSgbu60jftX2R6xWPFT/26ILkYXOSGMUpm
vlKdOfWhK8VDr53VsZCFyXDHIQvzStGlTOOWBJ0qAw7S3jA48gFPBVz83Mpr+ZZw/ZdchWFstS7Y
75fxqJSXFXQIO2b0YAbaPlIGfTsg+jXIV+AwmSXRHXYhrTzS8MjAVTSa8fHKPaWou3MaaKZ6qVWM
4WOIe2mwCH8tRw+TDT5yoDLgt2Tc/j+ISRMh6J3PQtPFdTNgXCiali/UxbqnTJaA7zBBM/zpqI6O
Iib/du+/23JOi4BEq5p6ioJLrtAiKbcWO4KECV/4euheWEY/ixGLLFNgk/9JBPRSVOEggmpENUZG
ObiXu7Qg8pErw8vqkDRt55DCaGb/0wFvtTuc8dWbTatl3eAXXkzLxUZ+uElV5jFsS19nqFO/jgII
EKIAlyJw0K1zAPzn81xz/4jo1sidIr9MEsF3WeVH967qRs//RNqAdosqxLUaWeWXQJn0S8zCNbK2
AUUI/UFZ69atgqUIK+TdFSsTMEYhZH7hleHJ+hQQKtUxhAyTnQNqzx8Ib9XnAuRv4GoQY2Nydvbe
niu89JWlvBIe1NEVI/g12fMxVtm7jl9MIbkXGsYxP7/U1vBA9sEhX3H8SlRF0AYw1KoAjEACmD3A
jlqeocCnsoEQbNEXK+TgSc/A8hvul3oGed0HHR9E5+hpWkjdwlle9liLlITJ/qTy2jkOaU9nMEoy
S6y8s3NhH68GF/FuubYH35XOQ/v72EG04qIBdIo3W7UbQg5ugRwmgTF9XYV/We0ZE5g29S14h4J+
Nem+FX4J7z2V5rRISV8XMFtLMGjmSG1yoQ0GcvfsAO04cZ4i29xee6T4OguqvLb15QugdM8oWfwg
mwVZQYfhT48mK+zOaA/5pBeKDBTahZoTnqnhlzas6hVoW/GibCUTiokYSevoC+xGk6v4iFPYPd+k
KaUIISYbmi8MJHqFDteD+ZlCyC9XKIlHBHr4A9p9Ug00qMwfa0Eu9NPYMDYt41tcgUg3TGS2Fvhc
QM5os7Su4rOGSF4MuKw16uWM45i/jDuBMGRMU4UXrJFatkUPraAF7OZ2RYfM4mkbvKoFXmwxciTr
zFFZ3B3d+/dN3mPTuzS7NGNQjddCfZru2YVXhhNaYmAKAP6i3uY6A3L+7C6zwMVtICow0DRfOFUz
omE6550lUdhvnPFPz25d6zCQ5+s8joH/48ZL1hQhPTGYqy39s0+VBlQe3SXZy36tvVO1/ex4QBMW
N+qDNNpODFnAyHcrIOP8ipzZ/1g53dHyQgO+R1/4AG/Duik2/wcFy5h/3xwkRD9idew2CKANk2C/
VhXYyfvAiyuXjZ0+9haqLD8MXIrzdrPod8z+tpw2fRUgfaO5B70ax50GnzJ6QwBn7kcH2V92q1+L
QrNfOZVFkgBSTHT/yzv5SRXNSNSrJENsmBPqcRZCYyYLbOLAIGYPYpug8/s63BnDXo/T9Ha3w5Ns
zlAt7Uo5ZAIQ4HQbpVWYL6ukwuhKkWX9r0+HYCl+jXRNColfHr2liHJXhmGUhjRQwaDPI2jKJCY2
IgHiP28MNIRn8rkQ30e7mM+YfyOlH0yzmMeVUeOZg96Q/PhnRypnSWPlKVaaYz9d1/V3qqMSHt6L
4AqoVrhBdlVb5eiKXlyxT6wK9I7csE6iPCoaCtBnTQKKWCcgJxELd0f6cvi9aI+O86/zYI7ej135
esUrWpvzCO2l+KYYyH3ygfEVnlavZgAvt8pp/iSF6CO1jMzEsB6ACwu2gYvPGVFz9xxh183kHcvX
A5mMF3QXygnlpUQb697j/p9Ew02Xzwdg3JQEROUflqH6x+vC9AFg78SorW5UbyN7jrUkfGDgwE/j
fV+1VTdQ+/eKxAAVwg2JGBXY6FTrVgzK6wVagsQUMR20h3xswr9AdsIFsBB56/IT0lbDCt9PtPME
/jVBD4GB6AdakGxnY2da8VUSiw4YTqF0C9N9UNrIukXiNL6fiElU/gz3p9YraMFFgrOEOJxn/9BI
ZBO3kAiYmVr7ZmBCYs5dpavN9/H7KFUtZT9BLM7trtFxAGE/CvMD1Mbq46gfT0Zx3jYaBv1Amq19
7z2Dr1A8HbAeogYYjO794GRIQCuMw7fZd3EEOJRFRJTT2v0ht/J+zh71igtdffmJFMDjhpMHxsfm
F0iikq9s1Y/45R4pYZLniYo8i8SGleH08hGNSuW5G5ZBsMbjMxqImE4ggRs67CbMd387TRUsdQN7
Ezq/YvR91jXkbx933CWmkWiKab95jWHXGDduC1IA5+oef5lQZu4YItDjGZUVGVO1BSIGh1ZVdc9Z
rF9NoFZ2IcpzHse2Grpcqusv7Wpiif4hEW7jGeErJX9MdDtmhlhf4keeD7Z06PXzQm6aiweGZJ4x
PZP80r/ixxAZlpG+sL2yhakOSdPbqenbGUtMgqkcbFbh4k79q06rNx17NXSPClYqQyg1YucDIn5X
6UZIqqxoerhGLblZT1B2gM8cq0gcN6uCaWFkqGDgsT2urdE1brgUL/yGtVN4sfoZxb3y6vsb5LRF
LSM551nBeATG2CMDPfa8u+iRiPx7tHAJ+adJPisa4cZFFgIOW5APTOt24bati2RQtzF8isR4Uj3v
d2DO8+MVob85plAi2Cd/DF+gmjO9YfXTq5E6G8J+TN43U0t/peXqErKU8EblATLsjhDn4/Z/Dwv8
hL0bfPPe/Lg61VaYRJGuHqzTbtbfyIgf6ZM35GjaEF4+yjJGDWLgkdSyoT60uUck9Ixrpnl05yuz
q7NSoH8CjmbfxSqs++yYofMCGMh96YmvYizm4RhGuM57RrJ4DYrKcR5DXdT2Dc4O2eEaWsyAG/A+
VhmV4HI2X9Yb0OYFKRxxow79IKaTBoF/sxN76JHu4EWQtJkG7Cgf0eajfzuirn+3qlvDjPYjeznw
fTEWFrQfwxgHqNiHFaa5LKeLgYfwa61HivTiOKbIHNfWx1IGrEm5aGxa4uO2ys39KW9UUZksP6x9
deNz/XtHy4KmIo69PH0ZqSW9p4ciXv6SLP4q9+C/30n07gAzxm42xLvtRAGg7NxEDdkR+k+1+HMh
TjCcllqL0oFrZZ1x8ulsILJcZlCIGy3r+mzkYOh/MLOTDWtB8hxEZjYpl6qputkXRQ6CgWl9KWXN
/Us0FdVmHYgiByb/JasE3Z9djG+xUV5EN6P/tOthTMAZTYDSezxnge5mVQdrjMFeJLwdNAe0Q/m0
NIi6GhOaAAhCJC65UXi0boDFNewTf/08uHf5qv23ggFXVjKnNRHIpNcY/YqoZQj2x/jkg9/NcAXR
UQ6uPtGsJ//P92RVFVsZET+KIRnvuzGxAKi679eT7yYXYutXeOCR0HQeAKjJm6vO0ZnShipD8km8
52yEHEs+Cb89P2N2cPslswLuv0E6+kyPiYfm8k6I/nkQJthkgLt32kz26O3Yno7PnZSUPJ3W0I66
0Y0C0sblLw1OnOgBlXOQu4BfVef7VTQz7CTWMqwWNuS2dBNAibk58mq5eMt70aVax/zy68TRP497
I0QOLZEvDwXOZXWhSfquUPjQ1AzDQI3qFM9SoWdBEyO5+Qmo8egCsoGyAaa4hIhU+hFWi05zhM4O
Y+lPmh28UMXFvAnD/O89x8uvNxXHUI5FI/NxbXJqRxQWS+afb1DtNgE8qqv0qHdnrJHTf+MClzP/
SMYwbSalJJV76HxF0AZyZZAPvtZsgv3milG28AkC184/KCD9p+aTFxAcmc49gDxLTHREF+aGN/3b
bQ+ROn2y71gafkfcpwF9DobI1u48uJ/WOQ97POM7i73vhTYhDxZAT2hPXBf3Hls4dEjewyFOtF06
ABP5b2JaapIcoQVwncvO5trLh9yhrWZ10zKDYk/pR3vUsJavN/27W4kLa0l5D7Q5CeKXjYqDE3j9
QRH5N3oXqLXeDCwC3hJdNIhnPD9Fsa5K+RmhDyv9BqNGFnvSRsXG2hf4DzDlHOz6QEWdc9j3oeiu
UMTtv1Qoi1oSueOhZCzR6ZKn3+pO8TgPkdta5rKpmICtFQG3ozVRk9AS8P+dDVmmZEfIIYBccBWp
1MsUdEFOsjl4PWVAZHnNDQhex/Uji//AXa6V97mYjEUOxKNvMGgEEAIp7qpecnNN46tvoANAj9mh
9R0I1fp1x/Cn6FQ6S/Gp+FJFqsbtX+5RLnOy2xwF2/4Pp25VtC9eMfujszuCtDtMZyft0ehBukkK
HcZVA/38MrYBjD1sxB8cuikCJHhK47sro3LjYJ4fv8ji0m1s0uNz5RzFgEeMx67WAiHbuc2TBzv6
nP1RqclBKOD6NAmdAbXX3+wsT+1nb8PvOdS10EAaixaFmjwv5UzjaCKW6MLnoFOPrL/shjPfphGe
YgSAeh1dCYcLyZAqeieFAiCzGBFLwPuz3qIRvYMK5Dz6i9ehBRD+IihPtDxzvMnwDnAs2nI0LCvW
TD/YKVfYqQ5boWrEUbkF1Iclmjhr5wuR+cbToSrYFLBczIX2tpsJ7/KdirxDEAv7OWuTdI0K88nC
v3qZ8GWvdAVE4GaxIPdUaKcH5oQpR0CL6A8/EJyAmV5xn6s+hY8AVJjg028zEyd+Is6FQE0zevjd
dDafO/+UIB9nRWmlQZVUBD2j/sjzs2Pbw0ENpxczLG/MlF9dkfjnxqMdjPZvD9UyM/cYOOOaPTYz
0B6R590H/JrlvnnHfmvRTiZJzcawlBeaP4RBbno55uUnjemT/ltt68RvPnTMI6BIY8eV0H7PkAJw
sQV8pGoERngtYoxUJy3+Hhs6BH63zyx29F3v219NmZ+Iafgc4gHeGp3VDHlW7BPncjNaWbnjEQxi
jMHf91xz53h/eTlqyRM8dQJ5eunlTk2drKlN1WGTtS3zMQGEIKe24O+Yx9ncgS34zaZA0/2V5ttQ
OGDyPz7HPem9tu4/2nsGE6mMspAdFIiz1X2+uXA9K3HKhmT5NVUX8a0IgwASug691JF1XnPoofz7
nBsnVh6dS0k4Fr+CTWM9JsFDTpivJIg+12e0UMilA4qVHXEP09Tj1kGKHJhZQC8Bdx3eEQiDfKZM
tl9j0o/Uq6ouVT7rMmrO4Gw4j5kRwYQJ/nChOpG7ZWGfgQ8I1HJ3IyZhtnLnzVPl7a9ntmiOswQH
zsEuf++e0u4x7TMrmEelhE14FJbDe6GKpRnTbo+U6aBIfjoYd8yiO5N68kRSYDS+PMj8Ljdfh0ti
kZ4BazBsakEYoNsl2vt1GPVd5oU810oxX4F1AOpgn3Jq9JkjMmv58oDlKR3YzOMgGiTogbZnfYUQ
xWVIcS8RjGFAV4ygnZPBuZf/KLIu3SCD1ElgFlOcyesAdHI7JuNM05mzZCZwSIsXs+zm/MPnsxKq
s6wR71b73W8oxu89lESF7TK/ak3MYzsA91Wti5SCZC3AaiqH5dJO1mZ5MSGXvWophtvi7owaGGnr
8NKaGWBkMyi6RrCU6mlLD/7O641hg0WC4Kswr5cXOjCgfzlxjhNqN/82AG9q8P3Ljgs1WJcwBGSc
kVHic2UahppYmGBAi8XKeYlSrcNI8y+niu/fYk1xjH189Urj0y3N4D1XPLNmmgEyqj3O2vLn9gLQ
8x8iaz7I8+2OsSm3Sp+v3d4t6H7HLWMQFnWOcXxsTq7sVwRTqj2wbq5bao3iBKIR9rnjkX23F4RI
oDcpzKpuTHbP4rBMb7qjyjbBj/prWxctWhC3RRlFsfObjX5rNEn4OqRyw9QRIIrFXV13umR/n8bz
eaqtun2wUU0kMliJvHVTKz6611RheqleZHRvV0x8dXfIlKI8C9pMhezvBYdV6DpXh4GL2qKTWCIX
R030J1ClU1Mk2+uBm414HP5qWOV3zjfXIhV1kvvq6bS0RTzP0bSrBVyA3cM78f10FhE3vioZh+pg
KzYCLOVHHqN+g0M4gJnHFkoiqclyv8WT9GYn9SlhgcVGJWDigTxFV+Kp/71WhaiabVFTpt8fFVBy
L+IDWJSqg/w9hfYsGFNtPUn/xqimDVzG/cTGCJmemRNaCLmI+FhfDKblYIhUZUBbqvy+9IvPREpe
XAZJgPttHO3yecwjAsQqD8pQ9ud9OP/sWFNx+D5dtSAEVClnM5M+pxSWl0Q50J90kd9N7/iu3XCa
EEj/37Aj09OIHH8DNCj/XV/wEIoXlNPcfrw/Vl+GLVUoz2PY1CQzcTJJD/xT/+mQXoGaqbFaW6qr
/Gl7QpV2KmHNMr5u92tZnN/a74OBDtkzjP3XaBoQgm/0m0IyagwpqJRYpamZtcXbedW5IO+STmhs
XrbVgyxI2wOfeWdkMtU0Mz5CLzL5KScwdx/ZiA23jP78UoYjyVai0T66qTb2c7cSjPiVk2/9usGm
1ikYsYa+ofqPTEFc2T25gMBqEyZI6ohwyxrTvjnD8t2nr9/szNZ1vWNQqzRpMM1dIE9wfFnM2DW/
IYDNWGVdJ4fnGHDn71x6ravgrCpWUT9mRhh4D1A6bOYgVPjCR2niV8hCPZ6F7lncOC5aX7cXLa0l
gEaSaakAJmhwPecTjK6nCOM98s/+bgr4uNoi+BQS0P2/Jx9ADqyMY1R3m6Z8RXP0MYFyLdfPFrTm
cj5qoZIoswpHF6Lw/YajowdSQzVeIYkv8RatOBfK6LOmf+Gr47+KczBNHh8/WFjPx58WriQxPvrB
NqRSoKU3cFFqbCIrmkMqVQKaR5Hmws6ZrtPs0ulkgmKTQUuQ+hzenmPB0Idy++gNQGI5Knydr44l
u7TIgKeCknjCAufPOJI38K4/Xl3eLG9D8XSzQ8G8hxA2MkYeagDVJ/L6c+/IaZDyjXivmq1mICPg
Opl0RwHQVIcGhLK9JreLdh5TTCOsZ8IqjJlpb4Bla1bFhYf8av0Qp8KbMNGhlT5ywNTQsp4V/an1
hY9ic0jOnbkzQV1mTZAXWWjlVgAKSY+JqlzcoF4Gfigd0JsOeJ8TbVOiIDM9diTHBNy8v4D8aGpc
ew51PzK8n7oYfLXvYorQrsY83YHA4yo/pByeqXkhOXvt97y9d2mXIEPsjoHOLirdauQlt3bk78z6
eKY2U5HAWwy8KePJMUSH/DRt9aaw66gcsSiqd0bmrzPOlAfX4zTdQsYkNlbeVeaYF/v1V/lgRvmG
2Un7NuSST90Qc5df2dG6XsB5i5XYwpNVU8t97kQ0CJUyDgqMPnNx32Z0Tcx3ULqKpCddFnj8YMQx
4sdOPUKNXH4sTzLNbLvbYnXIQhhDF7eZguxxpmC4tAkqDoMKlxL/TmPr5yrz//YDj9W0XGFApnyJ
CUGiolUA1yTfbS/v7twUrA3ngnO4QL6320u0DtHPtTXvIfIRHZ3vRhU4BHRTZCatHCG6mhIq9ZiC
FcZuDMtqUYggtWgiA2734llhEt7/zbkl9HJedXmBwKmyLjwO0EomgiGqvswjTrCZkMJQr/tQFWP5
8q4d5BiUtlOZNwTeKGlGg+QX5+dQQ5GQXH/457JvMbeM0CHSasY7W7lKowCLnd7WE8yQWy5J+UxX
Md2VXvTBpyfsCvH5TTwdqhs3oKa1dsETPdgkX/sEg5fPf0ZEyzeK0cBpGWKXVXggnIjCY07vK2wj
IdS2ZMehGQpnkkcT7dlV4tCR4qHq7wj7/VeIqFngV+8p9qanwsY2eJJWrrEcdLOrL9VwL2flMvE3
LqMW4dFJeM05DEZTQK8+aIng7rI6gjFOm90u9EKgBTo2TTsZ+LiDIM2Zk1qFYRU4bnNuztuBIUMs
gyvk3qau7sgf+jw5xugbcrkW6oEMR3CqqV0RqK1crWtBJ9mORq1xya/ptyKfPasWEOtAhJ1loUBj
GYgTh4U3NlecpZFda11ava1roWxPikSzXvA8QsAgtN0/z/HTI6QgLwfuv35FtYZxoWwIskm0KmRA
9ahvjldSa7gEeLiCB1eKNTTD5pWEQgqNkWHznR243dVQXKb4ZeMf46PF3ofiZnQGw30u41pCWZyz
HS7VW8MXDW0SvDH1/+UQDJVQOPAR+8bHt2SrTzEK4YDXOA4gfUgTZs8ssVmQOEw6YgLXkWflDpsn
vSC8gPd9ish3PffRGlqINiUqDC/fRf2JVPJ8Z5CgYcYKtulVD+O+xqm3UWSe3zTgA3mWre12g/oV
IxNdWRXBNlh1BYUCGnFvAM7amBxhBGZwgT7xTnrwtg8aTxh4j/YwJOG2sCzRdE03VFDfqcvlgvhc
BedWyStC6GjL5pypjbFGJWaVkbdj83f70/vonc7t39K6u6lzZaMncCBAgUcwqNxuOjd1KQjbpUL4
wUIaGDndyvsCZCX/VxNKXx49KqPMcgIQQoQ6D3TVmCgGQVKIhGYa5d4rIVmbWxaBXqJGfQ4Wo9PY
PAzaCxGwmc/8Duu6HOSR5VXWy8rA5DQk4CA9uBwTZ5//1QLlumvMhbjSVteTOXbQXg7ISwS8m2HJ
T+HWkuj7OQVCkCJEr5hoWaLQCcRaI/KFqmy3vDQWJpMRcHi2waG+RJ4Eln7/tzcp90oxVdBSYP+1
kDSx/FbSNSPcTiaXkerxo+I/T6q5iZ8+oBBCUW4HFiAes3eIC8n9E0bhOHYQDFDXE68cCQgKScy1
gpkZ9NVlT5qaPLPODeFH6hevUw56v1T+9oiGGRIX8gOSPu45PKbsf1ZFybp18dICsJ6TqdxoUxKf
0xr78qfLmD9mRMXymHJQs+Tku1ibm0QzdvChaxsGGTm7dxgczUlW4hSv12+VtcDlot+0j8qSNbuJ
IXRlOZbkniVJiJOx1F6ptNKpZqqsbU2Fa2qXXwyeUnCXZub7ZuzXBOlJLsyMfZgmNfmhGjIzaV/a
XzOKPAXr4e/VIPoZXW6JWOQ2XK7tMWLZqUDRM7YpSiDPzcKU49bvuR2X5lTqpXN5Hhe4F0LyVCgt
HELUAdVzStckWFViPgxlimYZmF4hmk4v8juk5jQ8LDDVOzmP83clXphtunyCqjWJ8+CzWl1tffQd
C5Jkt/aCoY7i7SVznWXeqHtYrsMt6YPFPTPzrv6nRMKKDD/13qi4YOutxhIJ0aLlRj5j71gf4E64
FOsGE5LWtx7qfFUXzYLxQjRwj3TZlEPL/Pqp2a7Q3ZK7AwdLcGwgeCJKPxPVagFDtbFjC/Gr899Z
/k/l1+o6J0UWcYKmC4akjZdSaxYN/991REFmKZ6fOFP2qNbgSjQ74NGjCVlm6Zq47bV9clkD+1iO
8qDJyi5Fe3ptf8cKfYJ+XKRbHHD3yND2DteGhBETVriTpClIsn6CdHE9qcRAL8zX3S4nwEPq48MO
CanI2C60fqzXrT+Iz7llGEgCVmRnFCOECkseTmRRDaWvVFsgfDqHzlh1upVmMXQF68yO6jfMt/pV
SVRtOi1K+LPvVJqnMUpWO+WM8gZmGjZCG0eVm8/amf9OyFLdj3zaLsclO5vyZgDsISJOb5qkNXZs
tSmXUbqqqFG+g/3X3w+ojRxjmOBeBDAAFjpAxaZ4g1r9CSsKh0LD9LzTvXyq1LXOnOn+5g7kCsyu
1TBifYSJSTynBRBdZ1neKKth/fzEXKcJDhr9yg6oR3cG/cfMX6JjU1szlDwdC5u7t30VPY/xdHL8
kDxLWcoJKWQZi3KnHUkmUWrdxKOp4edGEVtggp+//A2zbZ+S5XgXOxiGd3IuCuGPMh2x5UaMwE1F
XjHEfUOsOqwaGRIwOnj2Pyyere1AOAQT4K+7dkki11Zfo957eLAymqRMoluZbMF4xMwsU89MvAMg
pEliwyeNWjAM0830FvmdoFbNfeT51B4PZvc0Q0FPhwncZfs8CzHX9ErBLFE/BMUTonworJRmzMe6
a0UsnEbXKDroeF51KDa7yLbXKKaqDYKWobyeOWStDFgKaqLmD9QeSrlxq1zx/937fB2UkAG0ihon
GHNnW/ZgaPg1M9WbYJ8P+OXsW3GTwixTnqkJz4Rz45UfFm91A+lCcuSvjsD2Q0y8XLene504EXgs
mUTv8MJBH4Lbzm+JEJO0pNYYhWh/ihocSPY45HX8jJIcG31guEHUPEoFDyeXtE7g00bemNXV/HVJ
wgmNwYeBhKaGsftZPiaT5P+HVNt3GaCgsy8W2Qi4dQ0rEOYcTuEpUIyGqLH2pH2stNd58xu5KPmx
QUOO75lD+oatAiIIJ7yzX5vqoD0u593wgn+MFBy4bWfCAJRn1iyQdWm04NM8ERRwlBVIav1Kd3gg
38tXbKF/QQvPzKkO1rchscEht3NEEbEZvaawbaDthueW0XOHIOpeRdF2085SzRKB01RDj05xZK90
KJ+eUe5+eRJE69nmA5z0BLQUZg7iDsw/ySh1xugCl1zNBe8lJdOBP9k7Z/GQLOt8BUtzISoiZhu9
0Mpe/WA44jJnNj66kJgyWOVAsgc1Z9KxZhQV3c+az7vJJb0xgGOQ5eypHLO2LWI94HT9mOW6Pg2+
jsZEtQZ1pHI0zGlOBqQ8Q0Hh2cKyuPEUlSSwKDnTpI2a+B9kOEj+cMtkEGQnUafV72Ty33v+mRl2
tByjNFghC2DsKjojrKL29t8uPxV7+tr6foSICNOmzZN+oMUUiiWChmL8Wm6PoMzNm2enKfPLyh0K
DAPYH6UfL3ynLEI7FUeBjtG/bODnzIVdnSq7iLJaCR1Nzbd7UmLBbnKIFfJ6R91KR1wJUS+guD1S
gE1PhhYmkuf7CbRiWsRJVhdtkZApvgiVPN2NTQ61veK4AN2/9nDqKUPZddTo3z1gDaRc1DmJTks9
f0JYn8FMdTKRL1/LrvmGicAh3ZX9p7dWsPVdcnHo3zfarmH5iV5O3itDOrP00eoDdkF7ortIxzZg
BEpDaSrtD24VhNDwazgjGkY+Rzud53hFQum+hogUCPmGQs+fuxPlANupSNRAzdoB4MH19uXeMXr6
oSSgONde2H2ZhGonjqs0uda75guTT70cEuyCUrSqHTNnfC1ZEom6+Qwgrysl5tWK6TZOaiRx71DG
897pxJvxzwpGqtYhekqR1eSsw9D5I8RkMXhP7ukeNNrvUG5hwQAS0gVkYYnaZl3DeAKWYhfQ0w1r
pwgZc3AD+KYRbrsLged7rmG7M0zHQxPgqNaTmfrigbqLdgx3ZdjMg/PbzGXt9+UIDOSRUV5GNe5X
xBYXpIvGsmifkZL3/RVs3ZJI5jA5XlttCDjdyJrnIdgQcGgakr7qP/XNCBSShDCnVlicMyRd3/KL
F/hcYPAGluApyulaF8Py4WZYdSoVF2vwrsj4nqB9/efRskEAXMyiIHbEQiYtwb9fjoaflRri1LWL
6PnkSHYpJiZKgXLpFxFHai/dxu/8qmFsp6I82/AEQbfvOsTxSpars+akzgYtweB31B8ULe1M06cu
MrlNMAHuOMlXmKIKUig05neAJ353XIVcNL8yWvbJHcEAhugwiLQZqvGjxJwyk6zZ9RoflBzW3F1C
yYYr/OxUrT90c9DkquNVav915CWC+E81XsyDsCVocnIFnP8T7e3FLPc+IfpZ7Qornt98JlSkSgyi
Ih9FtB7hj1Fct9c2U0BZSlsNMBcEU4gQ5JBbptGbb22HYl4LkoEnz3m+bQKEFwDl9Ipwe2qQ7tGZ
nUvzr/M8Op+5xVggwjZy9E5ZRZj7IlWabYssU6qKflo5EYifV4OCBvNBMPWpRuOZDv/RbV2nMX6v
SNCxDtx6ZOn6DjB3t+7dQmyyFaFYjCBsffYqXzauiAo2O+gPBxlmp9SO9rB/eER2IRbYAv28I+6D
6QMbyYEh7wNGtWWdRSiMrWaJsxIxnobbQKzutV6QUeXw1aWoqv9KDal65AD4mI3nIOeb8dS1M+Uk
29UGcxiVl7LEqsB2yWddHIDdzFQePUe9uydelhsQUrS78hBqy8WiYROQ7hkAe20OwCQiJujtucwl
aszcWLbWz8R7hfQhnTZW2oKcXyN9YpDz+niev97FEWJFxlO0bdwrtiWmeJh9usYxjo4cQgdz0rCY
2JpWPUOWTha/qExWbOCDVAM/q4kiWXDGJmacumM1zP6B+994PVqUT+Lx9w2/HdyoI1RRHB5CG8Mz
E8XiPxxbV0Eh+9qOusycH5zaM3bXferWuUV8wgt0jkP+9bhz7Q16IwzYLr9P+z+byfqdPb3mqKXr
40YlihcyqpcTX/IgZV+F1jJlzTXBnXfQ4K66bIKb2JCl+ieStbf4hHZHoXFDmCjzhHHXDo4HCrea
606Q083ZlZo9m9RFKfbZqLS585XOenl4avQnNgEoIyA4dCEsAVZRneI6+bUeONKZnuCuSROErP6N
S7rsFCge1r/BWGcr40FllW47RyhIIL7H3uKiKK55AHcmZVrIUqGt2OWaTJoQHnDMtewMCb83y7WS
LpcOUwtxFNT03CGpvGK6E8cuT9Rq7Ff/M6g1AyqKuujvTZsNhHwIWZRLeOH1+fg0dWYmgBzqiUTe
vtlomAoYKEJ4hWhNtFgvmC8cEWcP7IZ9yaVw3ZMqTv4W7ehZAgPG93IeUgyYpaYP3yooxOsrylcC
iBmftVz8HPX4bDRn7ViuEp4AZ5GesXuJ1F4MDBn4AbWTw9y90qJFwlNPzPUuLZxG+/gvqf25e3su
RYVdQT0obsusj7c8cVAqnnEnpDkjACKRsKor9bvEpwLdmvwkDt6JEtbMJD6Oqkz2VkrC2oCdmaZH
BEjeuC3jY596+fDYNyTHIDuD9pbYxgiLCu9hxGlgWfYoB1xN9BBtgOKJFs+QhL1tNQR3u+wundaI
VnFr+SWUsZQw5M7D5w4v60W71RLHtZNGAuqy99HlDTH6zk45WdTa7TKKvaCu8wQ1Eo5jB3G8Rsmo
Z+iDo//r/szCOq0FxmyCZI0PIf+lsNzUAdcNy+dsgdoMbHXSg5IF1O+639NURab9S3DUGaoG/cbL
L5D8WosConjnzrMcXx7ET2n93Mx61ACqAE91s9aZVKhkLOGm1+zKtaqp3evCy715FCeFyY1l4aVQ
aelk6aVb0aVl/06Z+muDFgW6rNsB7gr+gHUoBlscrJMibZpvIFDD2UDOC7mlOS2lalbLaCXKmyD7
aYH6Dhkn035H4PLfg2d+aXXeX9xSN/N2jdDy6c9sew6ZOV6m/ro9aCcs7UPVks850uzC3nQi0ojG
v3asaNgv1qcO4LWqV//oUaSQmc1Xvvz0lqwrxQYTpP9zOu8yU0aMVuYYIsP4E3oA6O69smT+gFme
dXo62BP8LJ4SimqOs09dcXQLwuuHbeYEwQK3t3sIbk1ImpD2Dqtqwe2zdGpQQgptQ7IlYF0/Yn0e
PUmhDCneWXJwl1iwn3m0JjYfFoo32vOBJ9qTy3ABtJZFvGmFY3CfaoyMgE9/VDzw0wLmVxfVG2CS
qxeWJ8ZTFEtYLAoZdT8dU8YNHEuTvwwJmuGLFv6DUlRfCc9uyrxzlk7ioAoqw132+vH7Yqpln1Ju
H+ZhrWnWXJOtn9h7lolsD+q2RVjFl5Ydwzj8y3GZvgJWhm30U1K3Ji03xvtceKTuiOfM/v56HSNl
omF0TgloTPXiB1N6ArGhV7g/K8iwyjArYTW2lcSwzMS/FlKCy5RS1EgUwsFzfHHO/mLRDdsf3WHh
tmlDEocxKfuW/Mx1pSXngVW90FBe7J+hvfD2rwoutmsxogq5iCUUmcwOyxto5w+A8zvdJ0CYw2dH
nvHFIkPz6Pdtu059Fo6MOvP/ZmJW1V3ZnsF4aT/a/dzstHUaVB3J2fpEDHDXKclyAh+qqdOZrmzO
2+o3ild8/zHNkODtHCbfqkXBzVUqevRXt47d8YL5dIVmoVGvnME8DJsYzedSYHQ6+IKmav1x+rbI
QQ7JqM0UKHkWTXKm1LjSqDT5UY+0B/n3QgxpbUF+XAPkiyrotFsDch0Qkpl/JxncfS6Db+AErWRf
y0o2JLtdkatb23jMJwcsBEl2+/I+YvF8PYP7GBPwyHLdNlx9NIZkkAyuHLTTVmqs2pGLjrVWkmtM
bwsvTcD3tSK1jUkkC/wH1ZGy7vbnL+RzpeMPY3EWQ+Y16NlHha3zGJNmmsXYM9PxUQ9sBCFESrQI
BW4uoe9suybqXwMmFBL8blY2qrN80XzYTIun995Pm9RrOIKd5m5IgtZb9NKe8OdRBeDvfwZl0MW9
ql7q2MDih8O8c0wem2l3WQ61uCSsNjvgnY4q7lHAJgP0ixyNP5He+oJeKstSKs61277994zFGwhO
JKX13LSOhukGjLWserB3pV3iKY5jwgXQgg6t9szhF3kzP6gCtEF7HcmRXukDcgetFdiPi3dMrtRl
MnKHMvxtRNCPhoCn/5C3QTICTC75La6hrpLgg2S0g1LqzFcKZhuoMEw6xcBzpY5SGbf63jujeI4D
zY89UMJPlnqHX6p4QPD1+ZgOLye6qtRzxEc2pkuhCkMLJVG00rU4U8BKkt6kplKIB/nEDoqvo5RL
4bXrI/E0DzPzxGOhyNqP5kKBBPgysTLml3NiSPVGqgXqEgTPbAd1j1KL5sy9EAEQnNF1MGATQyCu
0v8cQi3ysDpqjCUqme4BQN3sPyMDVEhbnig7f/1jgHAIlpviJP6AD4SzxNPHZXGbDUZvkktAvbPo
UNkC1Rx3SxD5Q6cJbeYDd1OVSbmo/xu0HtjgLKo3JpWzY8KVogD86Yl8rR2U9o/5nDP2PFB4Y3e7
KrYmfveDhgzohr7sgq7gfY8ed/ZYAqqdQ3Xtrq2YGCl5Dl3lzLQ8GIr+pcFmFQoNnbm5J8My3GA7
BxWWraU8KKrCzNBIurhTPI7u6JF+Nkys/eSBNo3s7W3T8BnGMA6QJzeNOvFN4ouL2pYqBFQPdlhT
AAFAJP+c1GfTIh3Sn7SsXZru7oOGiB2I5at8pxw+tzc0b3jvijA/ErsV7cDVz3p5C9JMUzO3Rj8i
w45QkkPDxSTwNgdXcI3m0XBy/DrGcc6dB6+9eIbroZEB3SIGzaT0a6367vEYSu1ytZR5oxoPcNn2
qarPaxQ0QRWOatbhBV1TyymlvdzXIiMJeocObciXuUdPveJ2+hoX+qAFOkt12+/0TxxiVtuX1RMO
hcEai64u/3WKGMlaB038L3eIUmJ1S+cGjvKJVrRTdsDGeugTVVM364lmTNi0R+cTpUZvfTMNTFuW
FEEHM1XGOLzQdcTzxgDYehWUGnvM0diVhN+XvezJrDjW7aDGrqfwsoJsSR+B69anNMfhjxE8FJD2
MJXEJlDSazRDB2nfupKyu21GWdbkiM0Fk//KDrU5mzR2Mqw+SeXmNEDKokIvKwCjT7i0SVr9VjPf
A1EvdHS1xLei1WHMKGVBSba2RXS1q+T3FXZnZ1Q0R05PiiDVivWVc+VvqRd+pyHgjEDvCzWh28M9
oPS7362RSeCeMhEPqk70Pw02nSmv6DRb8faXL3uFPotbDauKPdpnC11vBUOaj7oeiWMMV3n37HMD
ewwa95WTV6ZpJPhhQpR0Vr3Dc7nVUW4530zIBPJ4dG3TCvXqewLUd0F9M4wEIA3rKYHQgFTdh79s
3lBgtdDXc+yKF0IXw7++2tTtxX5g/uTQwYYNw22Jcsm82I8XvtBeJg7akPPJRMEDX1QKj+dSClYa
t1b4Ma0jxCaehQZCstv2OHancI/nD0agFdNoBc6KFttOXyD/HzJteokcvoPaf0wCeYQtTdyHM9Zf
7y/ScsyC2xSSbPPwLjkpTIbpJsL1XW9wgwk19aDeVXbU4QLj4BYK2rF3vnU7Tiqu7ZRiqFZgoPbW
P5gAcQON29Xt8qcQt6PRrS8WVuSuCspd1xFpB50I6cT5DFj10QEquV0FPCFqlA1RXU9/jJIeAQT/
NDiiERqg9FebVN7ADvmEnGX56uaNl7IgO03F0L4qv7thwWdCxoIdiYMetwfkH/TVKv44cXSJ3rfl
79K/wMEPtBaKTukvsQDUFcflxEiab+MqSTdwRvjnZ6fXs7fNUCKptgX75lm+vFeocSCOtpQbfR4N
9hP+eKRJa0hbEJkoLX8JtnGttX4DZtuqnylr+kGmtLWAi9Gp5A+fsvBl5BSWxUfU6RykeVAExx3/
78qqFNvD8DUJac8tO4Xerbw6I18Z+rCyJfd9dA/l5cNqxOdwrri1K6haaV00MI2lOKD7wX/u+bwX
E1lEH6Cc79OuLU0fil6JhuZF5bgMBCJcM84oVVzJHpmqW8IU9j5YKU0qEV62M7aRx9FylnDi2x4P
uY+QHusNeuFQ0EcJiumAhiB4ACB6u8eFBSIXV5jA0prQSlXrg2EJFo3XdRy7+uqB2hwcSqnz+qeA
SvHs2y0pXsWxhYA/GLZ0aKcoeMuZDNMag9vGGmg4Hd/MGHi0jhiuumpR5kQWC+7a35krkbKohmpc
Cg2VtKa19YkbNLVnuAz3uVk+8jxqlPL29EF2kTk59Rb63TU/3aZvmVXm5dRASnwMhi+fu5n7hoD3
HJ7a+W6uW1AUojK/YdW/YgQeHeR6XdvQ5e2GKVbZq4OJBcN5JX2EW9iwfj9wlNNgws6G+sKf2QFF
nbJUpI+x7C+bMUjOaLgNGKa+MLZpazhmpPLrz3flq3qi999u9Neuz5FjvpVFGpkz3EApMVk0arGL
G42/Qjz/+GJUJnZ0t7R8jsUmMy+A6m7tN/s2+ll/heDoTSHZtpKPMzNaazYbLJKGn2Aju0N7Tuse
73ELfjlJRKEbbnaJsqtjiEt1/WI6RjCh9sCvjs6vCAmLuSV9weJVc7frideE1XcFO62uShk8MhIE
eMKNs2jaHF7MArv2vXDu0c33N2umGERTjRaFOpRxeueCkExLJpllZKoVLUyb5flQxn7uYfh5ekG2
xgye5sAbJAMj+suirkH/nCfgIeHxuCUotfHuC/euOJXVJ366UTVxQyNLUSjzE0DLnLKQ32enHBFS
DPofIpriVBw2nVVuoRJSpsFVsWuP1WDKxvs9At9D2VSegEHATlPUWSSMJ/meTT0bDV+arI7tWhdx
8jS/qQOnmhsCM/ZaJX5MULX2H/HAO1SvCXu2DmlCG+yfTvxPKkVP3bqJk9DgZGSEciCfF9S7RFkW
v9CURUxQFPXMElhhRjXldSk+007m4i/+UjWnGkp2Gw/eL6jDhoMmxAwX0clBGBDsMWTO686UyVAu
EkxN/KVsX+qCrRqlpTyE2w3YFcCC9qTdB2X/UUKmF+2MIr2MxHm0HVmPAm/sYPon3J2qT6VLeq0l
l5JmRGKwCu+vb5IWEeHQwqjui5kfrkkhnaJyfRa94M/QBt+FPJk6IT88lrUA+eIwN6xw4/sJhYry
DIVuUQ9TVeQsjmzchutpsZF+h4G/uawnL1n7Q5rBX5UJYjNSAFNw4f4+f5hcxfFu971BDThw65EP
SaSa1x2DKX3K+T/tFW6FEwFmrEJ+Q9Nt/WwCQmFggDZFKWfIgDUrawnQI9HIu/FtXn9pZP/66nEi
4AP7X57LiVAIIbjPUb8vuRaczWW4r8OJ+T0E02gOkdOq4puPmNMfMMN4mkDJFtZmhF63Iihs/08K
4/DgKhQTW4Xy/j/DkHt9bsmzZnH1+qiNxnB1UTIdpwaCQjyHhpCPk1SV0c5afsyZKtHOucSRxEIN
mgc7ZY1VLkvdj2pitNIo36lUfsAlQwBfk+QZr5CJyU+SsdnIB7X261s+kL/nYyu4v3z5KoWeZmZt
A+1guNOCWLnx5phIxPslmtFB8fpIZhKxYu4khl2Yc2tBikU9qLP4AuzFvj7Le7afKoOw3IzC0iec
9BS8yNmsqYbvDYcuGsDYSr+kSuYHC+63/DWIdewVztNBdJuD+ng9VylG4L4psVsFY/k7wC9J0GrF
jyJ5D41S7TfkvLQJ68btluBPvi4m+xQUW5OMw4EUQHjZXcNTWPvCisdlRwX3OyZ4b6pNZaSa3GE/
+81d5pmrQ2kPDdj+BCHr9/YcuaxNP7RPIjva2cisx1HEo72KqDNrvaumw0X4y76fOXP/ySjmy7o8
Qxktcfh/k6ZRU8bwrD4prmQ0FmQz7c9R+YLbRYf4KqnMugb6bwohb0ta2w5BZHpZAqmTyEYnxpfv
6lrr6+3iVjVMtT96euho415qVRBw7pOxThBHwcpEpVrHdh6SdvXMXk8G65sSx5KOV2DByBI5TJJC
9o0zcGbFXE6GXOuEYiLEANkOxwG9rFI5jRoBOzrBPQBUm9zY3b26zwrm0jzAjdO1yosoF36LiSqx
bNLGC4rSAZ9tzP0YXE5AVq3T6wTOnn0cw2crU74kSIJV0IiY3HojsScX5tjNhSWOOibm98QY/xM5
BKkUoKzLTXeWPUmJX+iV/2w+23cuP4/6ZbJLIL8SNNEA2MG0sfOyGYhaNwtS795qU/P2SmQTnq1b
K+2EOCpPkInk2kEA4yWu7RNAt+rkmeAfvDpRmJWGtpD6c8yOoHgMzoqnkJjXfAHEDWmad3WRB24W
14jqoIC3joxZ8N+DK97S5TrNCoiENek2Nm0YK5bueReBBcWKefTbekUxIIhGyOGejL0Fg5A//DDC
IDqWpxRuPTqVfod9acsT5yDERTK9XOIOokoQkkXbtKTgJd/OcA1df317FHXsCJn+6n+3ZhVoioyX
+o/BsD65Uvrkn1D9dPsr4iNrvS3OzEFBUXN1iZ5dYTS9OBgODXHUrfck/gbP+Zo0tEPgVHlT1VUY
NJgwtqk90fa3e5OVjHETdTQR4z6gOd9EknzKNVwJVUsqXXLl29mfYdl8Z7W82/akheod3h3/0BqY
Vyruk7VRCq5Kv8Zqh6znvPrLwa1lKc83SynVy0fQ9boj9OGyt6jsXaGqwk9s3yxRIu/gtPbiQSpM
yoAaeqJbBL3hONV/3e5VA9tTI5CsWihHWlC1/4iKth4Ul0WSa0YDMoEJtAJdiRuVIZyaThvunhXp
5PbprbpJcGhHnC4PZTTA7l8AZLvnDct0ZH6W1wRqwdpcJ64hZnP22ds7GstqLAxupZmUOCmn3Ub6
yCNUnEM4atYioltJQtbM0uOmJtCbSvIwNJMXWnkFJLS+tWr+DAbptrZDMG3GnVr+JlrPhmdG5xwC
gmtvC+IRBzknCeKwc6bRuqJ/Yx7GaKKsxIFkx82OC7lJzwlLKfTMR3MGfcy31/hHuxZYWKZC9CEo
pXXTLEbtDRHyDeZ/dpDiyfZdtdZtxaRqdgtjfqVrFQQBc2DCU/y0smQL2Ya4MfSVpBu7/nqFQHLX
sZWK1ZiGs3FZ0bfg5ld4qPK8rH7ydvejDBeB3bdEQq0c9d/RCgHpd82I4IGZf8Sn1+2NcCB1E83Y
KSC05w4t+p4o70ViuC9i5QF7XwWwem+23hyDqa4B2CG+BnqDHy3vnjq7KS6yzNa4SaLjYd9oebbc
BsMTSzs0mV3g6Q0KH8AXWhQ2+J3KALC3Z61GTCu6pTqbsSurtSnX3xQ3x1FTPkhhlFORvcaF1kqb
zrr0ZQbALnm75EGb+szH9NRk0uOjKgmkXoQbnsf/Fb1/3L2V98JpKaOU3m3yJ9vnwitUfKakr5Xe
X36yKdOqp0PJ9vSNXlveM3a9px+P9bg7V9NKR2DQ1wOY5PywKLZj27/OArsqyHdo+fc+G1UpUvMo
EBUud3YlLSGxLrp8Nkvn8k2mb6CvA2SaMH9HusPVextFLP7Pl8gwjZo3Q6PmeHofbuKN1LH/W6+h
Gyj2gr5NdXK62dZ2YNZiYZahjRs1JTwmAE9I1DNz8oZsuI8m9iY+tkMgHbsh66Y+81e0y1WxxofJ
395KgSAsH8xXFgGXpluBgvH2qUAKcYzFgxd3hwhqYfuWIYpUZT1szRRD8u/6QZXMmdLsu9agJyRK
AodjuZcBtnvOxYRHMKmCvS/NR68QQ2HDFwwLW2J51ICAgDppNavC0uy+bTGUxxq6icwcwHmS8eay
1UC0LHVII0/p7IRP6zQMnvmZvOEBNJvo+Wpz3w9z5B5KtNOQcXdigF1osZYGFW5Ckleff+uCJdQu
cajbx1SFdtRJShrWmKQV8aHmAGGg73vSbmVCilcWb39cMC2IoS9qg47QvFqF9tFKYPlfi+oR5q3i
AT3TJSlnl++krsFwqbV6/XYBamVoIFke7CFW2UVwhdhkxMHlOv8nyvJwpjjIT7IGXUjU3hziOq2l
jIalSGmkYpGQo6AGdurHYdC4lGRCi15ejEGuVFRDrY1NW7ZLlSdtpjc+3Lq9W5bPzC+2L4d5e+0O
n3TasX5db9Jg3l+O1C99Y0Twg+v9V5JOoYXVoQ/fk4FToB4mWswsNM9U4fdxlxM681j6gvRE+F3E
d+SLSIvBvVWYFrhhZpPwIiIMOGKc7Zjqu7SSiXRZ9Jb56U4NCTJGyoyvYtoMCSsY8l87wUlxzf5a
VCiqpspDcPpnSGc9OZ45KlYCY6SL1HDzuo8hizolVGXscA4nPo5Qtf0G4IMQuphUWf/ZwISFu2QC
tEGoDoCk6ac+MdniSXKedgRja2eLSVRU6nrFcW4QZMV7GLechozDXSLvHU30cKKQN7QhpvHSzCI0
PYNh2Ju89GnutpCMOGxKafJx4ghGa9ttEwsW+gwZ4EUNc35AId5DhjAUcTYxwxmmuvy+7J++3DUH
DBrISqz2FW5U1Vzdlfqt2PFV5lko/ONtuHKqrESDx2gGV3giV6r5LW5LkxtTTqfDdYcT8nAAH+wB
dg8Z681KKy3eHwBjPepECs5tVcEKco86HleLznlWANb0WzAHvsJhy0lz4JNz+YEvUdQMFf84QCaJ
J+VCWXxwvWN5NRvJQ/+aoZqLqRMVjvwaWbmCYxMRmsW3JH5fDATC62J/5XgbSj6FbVJ1QdhSwKrS
sRZL9nHCtaKiySZEQM8wi8OmBeTMA/nLYi9KVm9Hwx+J0xp0dRV04HOa3QYuYIwK2/RyApUrKBJJ
r/tpe4dZJ9MSxN5jo082aIM2gwCyuPvlHcHdyRj666WP5DVUgH59bF1YIXMwO6La6na6w8eWSKw8
16VLJsplEhbR4cu7rvN1/ASEB8TC40ejr9YKyn2v3ftObyMYIQL0t3l3M+2aFQFtBGix+2NCPQF4
6rKjoNlaJa401zAvSWgzTtaNaof27sSRe2HYGZQVnwpeVRqWlM8brYAsGuHaemIko/l3+ta7/eML
WH55f8eAYdhOAEVJ/9l3BkjBtTb3fXRzYjTSFi4sx7Po12xMTcPaE0O1fJXwddPZHkqsAhlRxDzF
TZuukHXZ/QOoMmHVl0ZxlY26WvcbZVGW3LTGFaLuDxYBWNKsUekq/bTuzdLGj2+zwOBFx/dfQ0fk
W5xCkX7ImmaY0kdwy46DBBEFohSeaMi6lkK3/NiPif88dCcpVyO+aScfxQ3ngyBhEYin+JrZZEyX
o+tAWIQku5MCWI0rTt/qWRAXcfyvRzqmB8s+hrToSEARb8ft2hBZKUCb3FCDfXXjmxp8/RHF/Uwc
CUvx+bIuWOvfrLYqS9ldV3niN3oyT9yAfAEasTmKfEMGrwNdiUytn6Fa65SB8bhOadgB3e8gF9vo
N3oBLEkvY1+RGPhMwYcFLtJt/jw1dCU1Azn1iVp8PjcjHdidJsQUuByFvCS5qPQrwNX5LM3sk7Tf
/AdiLWURX/NwKLWbZ1okIOcCWRgFWOiqzRT4urSkgP0/zJ3ev5XJdG0z/x9WmXGv3Kg5NkvV4K7C
VYsA2BskaWz9P0+BtxKNqeeONVJ3ef20nStut2VJX8m2yyD7RfSZrxb/41kupEdVHlUoiaKDEsSu
d4OAR9Efplifxip1WN6e9/VYgeylsRrkaPldvyq9Y2qRXACYdb71uEPem3C3za9/tm/I5Dp0Iok4
Z4fWwAkrz5mPSoWHrfR/7e1B1fU/asAJrYjzQEn7m1mJdfl6vRBAhUPA93JM8TtTiV3edseOvqV9
Cd7J93qPsCejbH7O9LrqnAXRXfkNQtRbLpqm7Nq4oe3prZWA9wbGTJ7C/N0Mm/U9bIVCHXd+noRZ
1gLyZOshtivRLDjbs0nCQMRSV2rOrbqHIQuuy5FAalZr464A7Y6BM5cM8LpUY0xSBfeZEpcuhsp4
QZdDqSXtkql5m0WaPhTiqKaDLbc6Sm6+IAs/Q0l9ADDg2YcNscf+e5LpTlmLdScxlKlj915l67sm
0CSLcfB0zqW1BmzjkQA3P3hmZK2DjZ1awFqKYIIDOp/BrXmW8lqn0xNG6NIRV2UPxn4TSebMaJb9
K1GhzYgWyYZeGjaoPkRVOQLiFUppmiqTjeF8GzqiiBLdyGb1xu5BYW26XHABa5OuIfAaYziYlGtV
UVindqq/qxqhotQMeDaGC6Y8z6pwfBX2KjjcHG1RsZr49qVGaiMX/zhiwOlDRMpfCMNgbngUSMNG
FTCyd967DGUkrG3EIVGwW/upmwsMEcrHvj7NygbyWEqu3N0/6hd/mljR8/sZk3SLWFjMXBNQBNN+
FhZlCF8NzRzKXi2EUwmVSCiJHPNzOhJyZcWszg3fAwbbYajLCpinQtlwdaQ/WtkZP5F5TZkcCLHt
7zP45WmmWf39+PCDqcZi2UrMQ2jXG35EiXXPIR/Di4NT9o+D5y6GhXNKfdy6ys95FOEVMFPI/34h
oYlVlR9AwmAxUt36PA5qhi9zsU0aLP9+4qp9YZhVPyXMK3VA2/BVIpYKjHuUdvOMxQDxmEpn38/q
Vs517JLH8ARBHsuXbeiWBpc/r93UGCF9NiDBajsC/QigcbJ++KSDwugogWvUxg2RJvOI1HkOMcgZ
xTQ+NKrEn9IZoptUjPQOvXR+Jkkuq0V17CWjiE0U4LCeXX81yt+e/UHgPfdsgg84CGwNyDDhYISW
qIj+62vXwt/XWFEYQRgigduv8/xb+kgfOg2HDxBupkD9VyIod5pRODpgRUcr/skeL/gV+6QDUhYG
43WebxZG1Nm+ZZQ0CUiQo71unM1okhIdFTimcQmcCJaaQ/GjKyG8TFCBjCWb/GFI40ys9GcD0s0l
4l5V3uLhNxK7r+cks5Zvk6G5DMBWlU94JMAvgrjpjcgzMAGXt2wYWw+viwWQ393BXO1h6UGF83F8
TyBSK6Wes2QBlXEtTTYkTvBl03vNUvQPoxYLY87By+T7BltcIXtnuY2hDKRH3Zu/9E501lPPuCaK
l222seU6H66N49tNRxf5fw8NX0iOROmneNt7TnccS5oc6OS/KugUaQJnKTTJPW7WhQcc1f5ZhPAi
aCnALdw6k8QQ10nqsdBu7k1hgLU8llSmCzNXRYREe9U0sn2gTN6eg1+i4iq8hndd/TFgxoJu8h/m
4uJYEmFdPsEyysxPB2gkAq65NQn+bsXJ84F/0AGWd0qCSkksGGUJ61Z0rmF3aQvbbr0LGn010Hy9
jNRwTwRmjLIfnwiohCZm5TiHWLrXfPZS4eUzSCqkUILfrUW7PPLU5EHx7ibDWC75LYMP+qLZXJNe
DlV73JfP8Ru8HFUShFPEsv2Hcw/VbczB15CTaYOQM8BfEJkHaBBVO11RuCgP2cDB0svFGto9QEPB
h6xGRK1qCyVaGNHo6kMQ/2FgsNKoEbbbsEGmBEid9m0C6nhB75Gd9WSyciZHxwbqap+M7viPhSV8
mqAS4/JKv7q1fS6vKYHXDeTYW26PhuvfS/bDWbeMat3N7ucDIrkk4zSjV9xtXvGJkovWhIgypJWH
DwbngEfbKE6P87KhF9ZzZyqJ2CS/884xjw8LetenCMZmKIq/29XTsTnGOzrQVEidyiBiorLrJAV0
bjpqrA8g6v6VfsbsYnZ9VioTLG0tdH2SvW8Z3ycLcAzbZrQbNYt3KkofGs/89Li0noT1pb+UdmPd
39/UlT1r9hhtsxEDO+hooNKAc2Btd7HiwNGDirKs9yWOrV9iCh+DvfMaW2nZeUvVj0dK0+3DtsPV
nN12sNLCjdKeC6AY9D3B8hnq4hTjZAvC9Rdm4yw+PzBaq7uPBYIorMGYCxlXyNHVZ1D3yJp50UhG
iE6u7q+7M/N5ncqkdN6hnhdETHUDIMisuy/fvXcoWJu4eNUDzrPVGtLy2fXMiompjaorNegLBe/L
s3I+aJCsQqHnS58/v98/VrvPcgcnUB+y4X/T79tFJ56aaJP9UtKNTVvwq5RtMq6pkDKsE2u57g/D
474/RwOBQdmSEYIf1eAvXUg8IJGDIrR60VpOwi2BHxmMeWs+6IYGMGHwbWK32QFp2BdEnP8SnmNS
tvtbTOfdXxZQtLHQKs0PZnTy07HcUtK6NX2nZxJgn6ogypcs6o1qt17+30At+HYvNkOR7EDYcGGk
3luEFS4lmrUWJG9Lbfw3QmOGqJfyd2ioXQJWKivTRnlnWxDm0XNA0HzEjDce5E4f2gEHkN+SHn3R
w1+Lcx6NTWXGzuJ7wg69JlBvTYZ9PEPzjH3YATTT1BxG45nSpmfZNO3n/UOx/vZMJLoHnRv8MGBe
TzB1Pr8iCsVIs8sGMRdzKwVR/c1NKdI0ds0dbXSnj9SlT6XGs/vB8OSKyHI7iNLTaiD587ZAb4Sl
t1x/K2wg93T9frLaQSs+TDxXX1QxL7op/REr6FTbKoMxjcgAc7xgSumBocEDCL56r2d1oy6pq9T6
VxjWun4+BpcWyc+U9zcMwj5axpb8wS38EMbUsYzRYuW0WKvzcrt4W4F+ahMO0esIqw2njY5MATmI
9H4XyCEt6qpYYTG+Ilz+J6op5x2U9sMAz3c2ZX3WxHgoFMhmYbhVLrznsgWFORuGyoYZiq+iZ65e
Llb+mKPeluJ1rwLyb+DNfC+963CBqEIgOeJS44MCL4EN2YSzl55sTtZ9EIardrwbYEd1e8aPtJLy
7TTeJsjekhZ86Wp5wJngMWVqWHA4ZR7D1azAPyNUh4EWwV6DoULg/BQzi90WKq7sWpVIcOOBw+h/
NBTofHdbLJ13yEVh0BR2F1owO73WeBRQ3ANChfpHPsurOGuXvGpH/IbsxjR2ZILekXZ1iFOoL2dh
lr+iRoGhqr9wKHtdxnkXEtAB+Z9gg5fXsdkdpGZVoNo2FpTy9m6VyYdZhMwhopyrjYlYvVA6tqc8
l3sI3KeXNrgLpZ30A9S96HJVnaef83OnbhlP8dzaaq/Ytcc7EXkhkfuIaLgAMggTjujOlwCTa4rA
NKJ5CuLySzIwNEwBpVjyEaO3O9Y9cQcPJWW54+XvZXUvDF8Mrg3qWUoxmvnpqW1be7Ei7QKnViht
I5M79Jsh10JXke0vwUrUjowL2+4ZU34pkZfjd8dF/QJ6lt1g73cYNQU27IvnpODJWqUnjiPDJPUF
nmvOlitad8wyrrHydQd3V1vKAXEWQt3KvGL3FuAt7P+BezVUFBBeiFdLhALQiguzFOWkfv2qboHM
oGiGOmufXSHidOrrEbQlHlna84yUZrDPjjHKQmOBO/l7pkJs1tZEnUGOmSln9AbpAE7FzUwP1wa7
BqG/+PEOBICqLEy1odrN0fU09CpyHLGw2NCDsfQVTa263Cmzw6mWJMKOgEN0Kx7OMMFnIC4EyeEL
dQno3vjJRdW6fF73Az9YDhbxZXARZT5AIhYv1EOyuJV2lj8uMatRVWo9M6nFxg/fodbSzRNZoUVJ
Xw2bR0g9WKUBj9lebqjdyhh+z9YmZX31imxCBbruF12nvX3X9SryMyKSY03UobYtwJDp5Hr3kr/S
E6tsDt3k7vYL/YU3FUSsCl8QPB1us0IMIc9hTn0kaB/sNolATzyb22NWhvJ49jfQQSVPDaXTsRvG
olKZ+vBbKnUvCKcdShzL2ndVhi1uTxbxJ5VfuATA8qRJijDToKIKlXzura1IAWGoUyyUxv2IRHCJ
iz1uZev0zO7SBp9r3kvQCa0VoyDmzmaFerVc0rXPEHKo+B8ZiVhfbNl3eBUwYTZIhuGoTa+vf3Sk
lkgx0tRe1T059xrUUrymWDC3TUV/2XqI0IYtcPb1L1Bve5SY+mjqX6ZGZCDucLCX3HBqow1mTOge
cnhbJ0SovcqLhKZcvyf7Fk9z6NVNbcplyKcK7izcYNsM5cG5Ek+9g9wWVGqzxV2Se8D+xIvvwbjE
/UdcgOVczZsA8kkhZFke6vtyXvirmYQR9BGCIFfxiW7NWmifoiWvDMaho6nlbcZ5YvxVXXQCzvj0
xBgWKa+xDh0ZwdY8y9z9+qWTRqsWW2oaaUEqVP+BJtqsgG83siI3HtWquaHcOKS5h1rDpOf+u6s5
N0uq+o3DNDdmmitgAkHLVxih7AJxRPh3m4GcnTjElAeMibEEtCVG5BlzKo4UXKwJmfc5rNL5wx0I
6GZ68Y9ZNPaPSWuIeJsLBNwjelqv4hxUqGkP2D7yeq8Is6eClTf20EBX4fK46YT8RAkJtMDdbp7A
y0jzE1JpDI5QQiMmBtdVKQWbNoaEE7JPwM0pVF0V2JAE//xpXNkdlqP1Rl6UOxCOadNcl1ljxdi2
Kt2yjc22TFBhj9CB+kDlcGYAk02cwoaXsnSL3SF1gWLTrFgRSYCLzSo66kGtLr+5kQOrYWerzaX8
eeKj1cT9R7Bh2yWlcUzF6wFEGmW1UMb2Fv7EVlXyBfotdFXICLe+55dXXqd/sQEAZPBG1TJlwkkh
9gyCxtHqGUzw6DiXvYnNmO2KJe3Nino0SfInUpvM0LbmNlKQEJGXCxzW0c48KLuqhnuz71Un0ksd
gVDkiTIcpc2iR+WJgToVOM6ycRI2tdGpmH7Yu8bMS8l1R1Zdp8BpVTaxrZmMdLgbHKzonI6wje50
NWqVXez6h3IFgE47uq4dYfY2U+ex8UmbgGCQyK69HZGNq2xGmlHBJxDnBhv8+M9TfLLCISuUgySZ
t4HyfyMdGNFUZ82rc8DaORJ3D6tz/fx6sCS7DJF13AyPfQkVENJpESFTTsZeODPh7eDAu0czNZgo
JdhYwTwOkmL3zDAl2JJSHzxmZe52Bu0xBzlvnD6eJSlswqU5hIKF3QE/uJ+1P1YQ6zTRszcXTCA1
xkOOx/b0hdochrZKmj0OOHzGERdY8YAlf3lyEWkwh1/rtfL6kBb1pa1F7vueFRv6oZhfplZ68Oss
6ECT2TQNzEEnh7cV4XXZWM858f3l8xaIWFqT3JG3TPeZHddE4UWFgNhlExGPZjVrpjZA0Z1/rx61
Pgvscek+JLBq3gJQywWwnBMTWXd655rMBzgT8si0x/+tRtPcxB0DIo8VEB9k/61YHw41hFtCUxjM
uIilNRuixZ/hx3VNK8/BTRCZtwvVfqzZ7HQqPrt6XStJ4jMKGwWVrKMSrqRKcQjF/CISTusKlFIh
LrLWjk02ood8r0jF4F3GqQt37fYGPqAH9UN+BoS+FdSu7pveWcCEsfO3iABu11HE/9rMpGpyeQ2D
ZAfhnE1wv67v5WvbTIuzL8vjcfuMrYYiiu8MHjh+8wI+G6FNukP4wjIqB4Hg4GAOtcIDNu9hUzkx
Hr8fhHIn9pmWgG9PEyWwvPypwhv2GOd/kgqBsM2e6t69qzVBQlDqje++Do471gN3FXVsnx11E0i5
MOuHm1qOjNyLKUZtxf//cghy1/beD1TSka8M5fbJWDyApKb6P3WAAzem8FsIEmHyjy8K9H941fOC
lpsBNqaLfonrk4vJwU5vO4Ay3eUTSOiTos8CVQwIdDbfP32BOCoH5VRL4EFsSwSN0TmsOhVVHD1J
l2ff4xzTrqcUztlSmvb6xSflVdzxY5zcJcTxVJSqv4gz5B4munfyEZOC4sjEV0nXMS2VQQLX+6Xi
1s/EEe/AEfeJ5raHeqZ15K7HMlvxrMKpPu62/6v9BKyQh8/sTO7wnzbWxRHYKpyJoKwdXrwVUSkq
Z3kklz1VE5wApw8CzzG+Cpwe/fuBM3FbnTbROjsjFFyTtjvKdFOp/lnxQR4m+vAFPdlWA6W3ZDYt
weCLqKtl8ly0uRGk3zl7u5/COmudwepQeCwFdK66l5Yy+HKICu9FeRD2BzcDgCw8LcfwnTkq907i
8rDof6o5uxwqofX/YLYg//rdHEoPdQQpYsEppcwSqru8ja/8Ib5sAw3OwDlW3D4rv+erxUEFw87H
1LlNiLc61LOIVIK3poxTN+A+mEcIaNWusWYhv4hWHNqcfuM6ZGXgDT+slLS72f6FCBNxyIjxQl2r
YSDKc0/mEjtvkSmTAtGjIAypC9+Qd/6JvoVjucgZdxWUaX8Gitxht//09hnhlv1Vc1nEA3nDi5i8
R/rgd5el+WFV1fHtsjGI8bNWiuXKTXhzDXlYUjmCPsfsbelCABdVizh6tSrZOczfiHTTnIGdDB86
YQzUhG3ZbhPLoZHKnc5ZGm0n6g9SXqleNbPtiy/3dCcKxcneeNZzpVbp1kD0UYhb7i4HWJxVtxse
C8MQcBrVAWqc+pbhloyhlxlovLy72XUFZmEJU8DGwg77mrtrCLxm1evpdp0kQHZ/FDLP14Tvh0dO
5dTMhepToE0fxgmtaJidQyNNzvm1/2ammdt+cO8qJCPluQJlfPVKkaz8BKY0kZlGokIuQeqWVHXN
baKX5fVM6qFfXgBj1IXrBJs4cKYJOnBAVvvpo4X7Q9rpxnGQuLBlkGFzG54r8HQEiYoFNYsEyBfd
sVYXCgsY2Pa8YGnZeJ5OpYvSg4ewBG8EdOAxH9kjB5eu6uuGi+xbY5rLDJMJzK/L6pCcZKdyQsRp
VRHn8mgYntLv5nXjciGw/Y58KjWWE8sWfU0ByONw81DtuD9L30RVlZqIcedUVGh9zOORmcfQP+bn
qXwBemlpyOg+gQVFreZ7g+zafBdRKhZ9/v/PHrzh6Ida+gBDssEFtCZrYTbw3Ol3mt3IlcQWcyOC
TXCau88xtPFPOUdXWbnzossH4qCFg70TpqS8cfotRtRl8SNICeGfjf5U/0RZS83jI36N/Cu8lerx
+L02indLcsFY3x2Ma7rtFnwW6QLUcAm4aUEnENMwMpyarhDPPZHNNCQ6AVsGGbjsX94cK/owwKhR
JRVydpw6/fHUf1jQxbZ+rg1oZcZcqSWqYNNMBcuuGuD4VNGEjEoXuWHTB5Yh9M0ge3c5PZZhgqoO
LUP5WP9DchfXv47CfYMOXHg+B2RadLQmN4wua5rJZ2ZgqZB5Ve5wjpP0kqJ8sUBNW9cgRQoB88BG
7+S70JyOber6VDFM5lNOlTRV4cs0e/Y7g3qemlRpcNTd68yxgZmVwd7YpxhXt0CKXPogMvNOk22y
mWT/TfCYzkb5HhB090bfJ6FKDaafGODi1BOBBZqbgTLRcwNz2dQdj+4m+SRYWY2tI0EaijGjCUCi
RXbjlDTD0K15IqqxYgeHAlNZMlrE0Uye3OWv2ipxjhFrgHoDDfSH4ORd5vEe/l0tqCAQyvdKmOZ1
wve0S7ER1Ha7v3UZ1MBKeItmHo2JshvR/qKYq/mktuvMbIiAYHIa5Qh8FCNfMMe8azcO8PK8eajz
Lxq2jtw3teruk43nnnudSvzU/tZ37PRr++k0XTqONyVcfFAEqNpRz9gAeqMa1qVqIL0sSseja4TK
iuR7nTQYRToGf37R51yvFeDH7xF+Nc2muQOtwls5TGKasWNwZa6SIVNLiVwzKXMWLRO11hIEgf2K
c9zMhvwVEF8ROYus0d4QVe+3qoHHKAZLeHjArB0EX1p7WLsplK4RPOm4tsay+h+Rd3pmncvgnGAv
0KeN3UKyp7g+B8ldc0ACvglSlYQVkSIcQfckiaAkamnc9u++5IxgAudl9C9iEC+fj2cQqDIPn+Wb
ejEHYhPY5yEm3q1lE4dywUadWeEWaXoyNS6hnKAF5w0sKOpZtHFiK1qKvfu5KjE8o7p/h3+w5W2n
epBCZwiwXA7YUyPHtZIycvjtRQsS9RP2zeiIwgLm2KFfMiSnO+ROcXAT2KXMgtCkViIjRRO7PNtd
uZvb4DUdLHwmvZX6C6cn4qrjx6LB/vfie9rnQSa+e+CuHXxKfKC3w3Hd3MzqlNKx3Ls0FZ6SrcLc
MWf5OO3exCFp//bAqHRO7fHPnt0m10A9QQgobX5of7yatFl4l/p51HaBFa9wQ2VWytBlWv+wGeaL
ohilMuJ6elJ2yohbMvtSqigfSqpkeFxLWd2Fu9BzUIsMsJAhbZiFVQrx7+jp2Lz+aebyIXF81Wc9
J6eZYcJ5YPn5+kmSURbSsASh2D0N2I7nUhWMKHpvVjgh67PclTOFB+33GBLvzONorhnhb7lABPfO
HjCInS6xXq18z3CWs7KNrQ2OgVVbQx6OyFFZ7qRnvAnXqbVVSbqnBQsQxypZyo3Ki5oYLn9tRIAQ
mOHx+WL0x4mBXvdBeAhrzKAr8/2HtFceprOHcFPbeckiirbHFJufkB2pkRA7MqUH1eO9OQL+Fjeh
EyZJp289bwvc9DDcAQlCv2MkBYJpYNvmssB1j9KBPhkvDK5K/IuXlo3WZamvwebFRiCYa3M1mIfv
fUTgXn2aL5boGmbCq02Q6N77J1VjBrQiL1RU74arWq/j71+cH/IB1P216GsCNIuI/bEQSrXglgFN
axcCTDTv1lBSC9xbsDyp32tjgSPaWKDp60z7CH5YbCzwcacIl01LZebdE6bN2uPVjCkcejuZDI/S
9yzwb0bT6dYnM3PsdbgGjIibNz0jMy/N5rGWz1fu9ZBvzb3dtgtsG/a0sZP+v3i2qLbF31ANvYXc
tdjUr78A9yLeUXTXWzkTPDON04bRXIUwWdmW+PLY82hBn5N7/7FZnGa7Q+WlY5FfQuSoK7bzR6jf
oFc590SOzI169hFwdTPfkKsGMc01A7Ofx1s1nI2OLO7JgaAxLwGSbqWZ1VPTQPm9x6L5jBKS52aQ
k/bBHaubUNtylqlUZfgqy8PpcWIIuadIWqFGAgBCeFt9JiSyjgURtTUVMOj/LVDCXXTITzgez60u
wmgSDtGeNoNP0HlWfTkGBYMEor5bcFzDrP210qntZxQP69zN1Rr+KFln5+5k/0C8U4Za4TD6xEpg
bcWygyWIsD60rRn60/HnZkiH0QiRn+hUREUeT0PdcqrM79omyZ5EGNiRlcIow+/g2auoXrxOfUmb
0T+xpW9AeQob6Zu9Wf4aKsurb0w0sIvG2LHJoF6q9FGNHk0+5CBFGL8V66WMG9N2JlWpQs0CluA0
Et+PqhEp3fIOykowXfY4/Wdz7S/hd62MsnugPQBwFbbXFOKr1OtmdDiwxX6Ai2Nn9d7hfWI3qaD3
DKa1fcERVh9Go1pmZP8/QdbkeB+DGNpniykjoiJYx0u+nMr3BowOWOFjFUgk8KyuxNC9bJ/MBti9
+zm9s4t2XLIR26PLm4dgt0VZwoYTitIabe1MvyFAzVtzIwAAEgokOZ7Q1TCpshW7ljIiSDJhnQ+A
QpS063Z16GVlyduO532we4wpiqLmRJixPY4jD4a4twMQDsbhnVlSiF6O/me4NlFW73zeKt+qq/it
39zUkBHsXoMPbELhFBQfiX4qWt1PV5QX8ipNcpvPOZMepj1Rj/AvUSJaP6f3LA1GKwjAsmvKG9AY
CAin/RFIWZVvqYt80z2WuFKxFOpKrW+zGvSkwxwgc+OqKafCOR4LQ0gmJdoHMzigliIwJyTMJQCg
E5k33zscIpwPfl278qRQlItKTpEUMzH4sIOiccNrFwSwynMf3+hBhIVieChuq7fmsAgCaJJMcmrv
TVzx/8jnKCUoHXA6dATL/m7V3zhmy/oiIQc0MrTfiW71Grhj9iNREqsMCJHY8tCKhYuHz8ZEIkya
YyCnbdMLeKSDwNGkcQdN1VjclhWOhDPcqUD3qztBPQ0XznR9f++9otJRbqxQevtJsCf3TG1W5rTo
BMgu1H0NPic6hLeYU9pD7a5UzN7YIPCVEYpLRRekQuKE6EafI31sFvtLOoIsruVqS13k+/ItsXuZ
320jICrGqlJrqKSIab/4l58EbEm10uhpk0d+e4ZtL4ggPlFHYMCGw9EKogfPI8pmr49dhneINf5r
w4mAyvAWY/XsAxnvpS20n4PQo7J2cofAG0sEqXpTXhpgam4tfKVJWGyvbqWTOii/ykNnDBmM78BK
rC5utaYuN5Sc7iwsxZEKgTh0E6t6AKLaqnLgUXX1zC8dQnjaOCAt63+VXwY9J2WiANQBBNyP7yJa
whqEHQZah3Xaow5Kq67PmmHnUhfvCThsAwbypDMremekYMmGGJ3ha9bcNL2qr8oHTLFWD1qrFDHP
x76/CpAnJ9GroKxssbVHwBj/Gv8A7aibURIjoFP2Rr1emAs5vt3l4SZX6bYTgRSI/X1yKW5V5KAE
w/inLV7b/b6tDjAkCf4O8s6o+VArSCAwlQTAqrz/UWtiikgCSHqbEBbpTAJdaT1PCI6Dr8WjK1LZ
Q47GOimB9gHRJC3wFnlSSH+sv/HX7rseHkx2acQ8MFmuIEXgXLYcJS3Dyp5jc4WDgIUz0hbQCFqj
DDbrXtTKrMpewlSb0pn3QwxKjqNzZRYYweWPdBJinS+XB4jsxZWTdfJRUXvKjpWZhjFFqGiy7v4E
xmmuXnKwjt2cIpTq2PaqZknivqrlZfSwP9y2IhGnbyFFoii05+FLM0EaTV8z6RQbyEtjyAqkDqoT
Kpts2TKtaJzyfXe3cA4yyqicqiUbYZcIkt676FNLaKUd/UhAuSRolEfEpYHVkbLRsnq2DhFa+SpY
UDOJULJRe/YqguTnHSN38fs1R9cpD91+6tonDs17K5Oj6ZQnP2WeTCDkWRyE000x0eLByDVadjI4
RilRjYcUKOb5mdQp8IFRhx27WUeMl2TSUPeIR1dSZm0bZmTipqQtU7EUDzcuO7t+HXcpLObuDB0h
D49V/tVk8uPtXXn4phovFzwOmBT5AjS338svn9mvpGr7pGlkaZ7O0uojc/gGDYScZFCX1/mRxIwC
wYLgLqU+Z5cBWBm1IvcnF+9kjybQ0mCtPOYeQ2cgXmEZfoQHCXTapegFlO7DnswTChV29ADFF+d/
axwb7ywWBL6moIIk/zI/nXa7t67FaNLLj4Z0teZbc8LhWpJ792n0LvV/yRCB4/UsHyl8WNNSqfuX
exYwWLEy8tvIJAr7epD/OiLZuJWmlylR6zXqi/bUQvrZqngnnuuaNqaS2+LMHDtTPCH6shTEEbcp
tFcWf/KRmaYYAB+6FTHW10F+th4j95DfpRsbwIfPD/ZtfqfUYGc7Jb+sqeMZGAkjgLRIhIEQ7orO
gX7jCtN95yfEVNW+b5+FcFCVJEm7Djcgxcc4cAJWJoC4b9QG9xngSlgyq0aiJ16iXirnujbQ5qc3
ne2Sl4GE9qNNKsbLb+6xQTJ4/Ogf8utkXxhWX/RoTuy9b67e+sXaiodnf8oEZ/GnpEzGwrkOjzwz
kFogkVcpHx3xw82EtrBkvsSwl+yUZv76pQ+mWYOwfzI1ZH39L4DlF14ABDF4ied9Vmz4gH4SZ9Fx
/WJ1/O8GUCxViMKyzjuH+GaVRhpd8q9Aqd/QlHISXM5IOd0oypqfQsHMoyz7gMqjkqiBgCo/zfKA
uEfkIFA4w0bWUt0AqhK7SVWenlSqDNPOKmxJc4YnDPvB56U+/6oJ/9G6JjBSFs7dm2m3yqLcUGy8
G3yl4Sqwy5w3D32BKZ5Qp3v6F5nX00H2q6JGBRLlas+QJFT1U53F2F6Dg+DrBWVr/tRqgR8rq9KR
IlPoJP73iHtUxv9nCGHn7qPcgduZ4FpOl5MFU1JHQJerUobApzYc38/4xh3+USLSYjyj5ObktQBa
qoAVS0Zgm1hCf4RNcUbFhl1lmD+iVPHVb0cKNBSz+P6bUH8AVNYLHUlnzsE/TyBzl87zMiTzBUnz
rmyLtT3g3nslOLlXxb3ckgj1WfFJ/u2Oew/OtEa+cHra+YHWjlUbYY+3tIJJgfRlhGCug3pLXmzb
+RzjjPm4ndhEd8D548g/vM5RzvAK2wlYk+3pP1tBF6QQ9xX1as/sdjZ2ixj3m0DW95J7vH6SAePG
EF8TxHNc2M9Wqj8O3o4zJfhh7AUqSdjSaGh4cG7Xs+N+s6oezkxzE43enLi5NfmRTy7yCB60m195
ZWlteh8EGlwNacZqBDmX/pzWJhmNLH75Az+uXuZ2VaNNmPCqxXcyHeu0ay7HQqbrOfFbwTPqACe0
V57+EjKyFiDlFg5UM0XiwUfOAlZF9L3TRZL6yz3k/EA3xnOFMlQgGrtnP5FjmbpmhjC2NVl56HPd
fq5eMTeR7NlyBs+boGagriIndEFsowykGHUoWr0c7w845XIMwuiMLhRGEnZnMY8obDI+7ExsekmA
8qSsVkYlfxPNdL4SCEM3EJPVt7t6mIRheMjjsg27sG1c2o4yayoC+EXBC5oVWW6HrPhWynlxPtUf
qjw4pSAx76F8kfk8hSKYTwMwaRwZ9HNtySMDWW4tcHgNXZi3pwsAcNIlPPXgyPp2367Je5CxJn2j
TrwP+6Y5B37dyooqFnPqRYJGjJ+G53sopPsKpH8u31Dj4KB7AD3Y81nxyf3jTpE8BpGggSbVOQNh
7pCl4ez5Uqq75GmkMXKCE/MT3A+JACb29JMa8tWFS1ES//LJ0SUFKD1iqRpX0ju4PTS8aBsORY/C
HLTCbVG04vxat8nbK/isagZdHVPVEoAXUX8wvhcSx/8lYXJkUsAT5XaTN1xJRwIEDQfoLtdQQZNx
xpmSLFXd2lDdTPL8a8unymn+leS2FXPHizDJs0pUrFBMhdJK7GFyVHxheKTTcbBOhSEKs9k4W1D1
B69BTF4GEQ9vZDVf5W8cKs+BtC5fhjRiR3IBgCc83pBT24JsChvLf49LMIQ3lPCmKRmzz0VLWu7e
02WUJLlsH9O6iuc3AAEpE9uoLeN95vn3fz9z70aIFz8RZvkWAJLvlgLKGQ4VmuJ62aJPbKwJUNgJ
l8iO3RiITw8NPhT33cdq8LraP6pAsZ8Q3TdW06ltCEC5kl0xCD0C1qeQTcxrVIpvrd1qL0gCm+lA
u2Wk64e6/Whdvul+0qF542QzHSWpznpQ1nrYLxIVfx1wwffJIroBZy1sUP532+fUG90ny2yMqdpM
PV8TYISOBxc/H8N7tmfHb01avsaYb+Yy8fp/ds8YNqh6jdStIMJBApuCZOP4p+dxk3YVmWpUcI5p
f5VR1+0zfiAPs8ZhgtiSMb/P/tq6dtlnvG645MK87BdmxCdrGI/ykMSp+1vB02Rf8kw2Rnm9KdbO
uPN8tWdUX7kQ+4Ja2jSVh/3K5QuD0q3IMXj6yE+xbSYtqhcApBbyHd7KLY/NKTL75pmYS6MjW1yK
uEV/4OGlyW39qHkJhJBbb++iASrRF6TSX365VIUAwlpqaL17bjDtBsD0WkztOHjES9PM0TpDUDRY
cZO6h9v+c2SXJPAHZPAGPnA3QTbxkg1ynIo5CmSfXpJLZL2DBCEp8L5tAz6kWzbZOMKF5bC42Xdi
iekTolwWWpiX6649Ft/uAl9EwCk/hXqOyK6panj+LtuQCHJaoHsYfaip5RrobOdSUOvInJ2Yu1HE
4fxm2HlY3jzlFQF1N62+RpVaaD2gjgTRO7iyWh93Er/Zvj+0C1ZoaZB8uCUdq4Zwwtg7FWttmJzu
q/G5Zbv/y2AncjJpj+sAXWV7Zv77D+ieX3XYejAZQNemGm7rz7L5KcCL53PFckuXRmlkX9vnFe70
JDZh0ujxrWBihINALhLrsbxKovmV9+n8kHuA2kpBQdB0NC8PhViAiReThAp6TGWTp75W8JHqfdc4
dAmgVM7un8kNTfuOWncSoFWwTYV7mJFZnyfa6b3D5+cfR47gAdrftuZJov6ZeACSJYynmkihUAky
kl8gNCg9/Cd2SryKcMLZfz/goawZejgXPBGwJhesr+BERAR7HLcJVF0L+KSqyhg57Tp06oqoA8px
CrwY8uvnUytIPcvRKDNfcZTBUJD7suCPTuQXJsj4YbiWoZKv+6nwonVHCLszuPWnWBvn3ImcVFfk
bXwFwwAYwhjPlkiDsgqBuwXlPhx2nH5YSi3GG5Y/3qxM7KQDO87m9fznk4thUq10m0X50Q0rMiAo
GjI6HNjgqgjz3gVLs1NbPpjsIDUg6Nlzh6ViL/Ro42r+d5L3XDECRUfAjPIwCAs6uBoVXF3OEIUy
e7moXD8POBqV1HFLMZgVj5yk10lvzwePbFCtzf1BOONcsg77J3zaPMjD58gzNokh7orqmY4bsTkz
3RoORFF5lFcfa4fCq/JXKyZQbksF3dpAzANmKPCHusjvAOFdNg2xZ6bqQhj5J+epeB1OMuy5V/+h
a3PUh815j+8pYCWHrZJu/6OvRwykYGNRy0BArdUWg2iI37sGOaRtBE6whsYLNIVEIds4Z0SNnYUi
8JGwaI37YCAH4mMEx0C5b4iyvBT/tVTmj0yEXa1QeMHv30LRlBdJm7HjfUVHgo1qzUnA+kUekaCi
7RHG09FqR0sQuCS3Uq+bvANv+bixr4R/36YK/Ph1fbNmn4tlLKEGh9Z6oOyaCKMscJYaES4PPrKx
mSNGsrcmeerbijxPC0cSnm6ksicDzaJiH91+Bh8hML+AvUX+QkPb4sMIc2qBmBP0WwRj92xy7sSh
DfybEgKRyB1+0XkCKetQ7YUm5mIxhq0weAV5fkZXbUQPOFY52Xb3asEINkQsaV4te2zwVO8BES+X
DaPWTdAYo14sRRyvCBvMxAjcnbE/FTm5ezegia8EWRrv4SWcFevgzWjgeIUu8Bu4/KtuGXDy0nsO
33aVMrkGOq7AVL2vCvkHwa5KkXGkXx9Q5AfKI5HJwskwhqKf7qx21qmp5+prl5IZ0calEu6UwnX9
89a7tX0/6bzwRH2ym8KYJuFUW587jxk9na++t4vKvsYLBTkm9itjdJdAFHznELrw0Rh1vKEESRy1
qQo8VZdyFHdnOHgQXHVRGw9YDUQP97RSW5V10Do+BflR688tF6kF7TGSgsKO4tgwPIKYP9b1IHcV
qRQu1HIaW9jE8r3e6V/KQqzdX1c81L1AcqTAdAVHSAt2x47sw8SfLqe0aISIRt6mVFTB/3EDIE0d
qs+G1tAGUSp34a2hHViIVYinudMqHyX0hjbSZcvTwoEzFm6wt/aLKhuiLYqWA/Xe6uNUCK2ACn66
MtEv5jnh/yg2j4iuUAV6kfbx7LjWn/KrSBI7OyPHbhp7hWtO4LQ+PC0lE9C306PIYeYoXWzwtekw
bhWfKPfP9hjk6xw4bHM8GSFRzFhTQD89DYy6PJ9bwxkdftvVRRL9xDFrDKDD0A0QotF6B/mwlh1d
H48M2j0YV74VDYQDqSpJ/dZsLZ8d8ZnPbM8CwddewbiyOFDRU2UBefampmTsph4ENPYMUAGKD1c4
erEPXLWLohxa1EvVgvtmMbsM3yK+PQfSciaMUaQusnu1SxmsqlJH9uG8p42MolpZK2nvvPjsZZng
Qrr9qqB/ymzXTgXy+p6QBm14PLjV2GYOImhh7xOxq/tjlvSF2gKc44N8Em7yIdRsQxnYPFl1dhCk
9++iD5rluoWTXUudRo6wuiyI3gEqsnKPorLHQAY6qhmfv8qBRC7u7hQCwRkF10ViENBbaQO2p9Cl
GDU37ZoJEfCxnobZ4TgKjLpFgIaiGQQREFPQb+hoGKhfdDrysJksdre/EH1vl3uqW6v4/tg8sK9h
Xyfn9ey9wO/SEbaM2OA5jvp3dbqYE3MZ5LHcNq3FUdYY9m6460amwDCbILVGbvGV0r473AveNYHc
/29xe+b3G9qTtkKrEJBZpCCK1OdOMH+FWyUaEeh08tXn85BmOBDx+77DUaIxIZPOHLiH4VdCP2vX
sdJX/N1RUhvJixUurHERIphmOXSqwwhG2u9aE2O6y70iSGk5dDzelLQK2VH3U4iT4qFXluSlouT5
80xI6vFMupJkNHZvb5S6b+JON22JrLxPMPh8dcDU0rbr8pcbVWQoAokmozTOVCEHrmYCKafTRG4f
N77PlMLfsIJAPcmCn6BPIZ8Q0xkoq9fLLoTa0AiB9XmOgdfUXCn5cASpyfN8pYEMivWbLYsdmos9
q3CilcyNVdcxGuoh8Wvr67wYZZS7BouWWuObHva+5E6MEKsXamlXAag1msSa6LejwijO8CNX/xXR
IPohviupHM4cBhNRnqej6THuGtHSZJYEkIY3oRbTGnsHDNuq97Ena3RLijnjRB/A65vy8isEIpGd
wG4JzDq9lGsxYMmEOPGlutbBUVgTSRB0if3N0AGLbiGBM614r7ZVZkxOIMyIiY4tyIQKFmNZsDXQ
rq/ZmVYzH2cyXpdhq+/AM1a5qzRpdiYljFdixGWcYcAy3ybV9mRSO3Yr8coYpHNVoWzhqXxymOaD
mNMF1NIew6ST7F6LUgTTG7aTtRKipXnH3CMXehQ27f9eTO8C+pn6Dvq1XFdrgI5IThKLaW89HD0P
0wKkBDElU22CS3FnpyWE5rAHG+7ESdRltkGAsorlUhHNKkr3/E4pA92Rlg8ZAk3O8f7ep5MWk87m
EqnZUCq+Usu4NW/PtIdm/6uc59mw63qC8xSvQADoNFq6Y8+NMNyZ3XLeNOOlr/m0VCxYhLLPlv3n
eow/ouN3tR8xy4B24/82VPB/pySzE634+2gmuUkWpn/0lg+ziDAgoLvgAGZXNB3xjgTcCiEUuJOP
7+dFPugAXFEq1MQOQp4ZmNQT6bARjvw0TnFP9rXEDK0/C0+N6P4KwQlIJ0KenY4FUF11Gear4Kzv
+5cgOQU4uhE4YjduGxY9RPZSJmXUpmDYFN0LZdWCjHABN/iP4a+HHmbrE/HrWf8blQjBHv+UbVe1
oDEBDCm03YqlFvSheR/pQ6UPV4uNGD0GneU1CqwTrCsHst4M9FJoxeUASqJWl/azK07EDZFwAoWm
P4CO4elHnsI6hKZy+NtwikGrqh6PKbIhrdcb6tirRACLChYTkJdYJJVW3srtCOd0ukZnawnC9/Qb
ZiMaRU7FSVdPMuca2Hh32YtsxMsLqBhnz2R5gu/dnYTCKyREZzWfCOGMkFZkzPeaAuFPolYLxMQ/
vg3oKYStTLSZmEDS25QE00lPwTMg2F3qPfi77cIADbkMvnUe/+mPAZ4R6Se0ZYkErf8eY4Q1ZR+F
H84duj2G6nPFOovMamPvyCb7KZWgemQHpgwUwDqKciwpoEPzUQnWV7GlDaHYCayuM3SAPmdI4/qC
FlWuIc/MiT3GyAzeCE/h0R1tXqOThYMeNjPye4puYSSf6fbMp+KVOfpamwF/A8Mre9AT+dtKlgDT
whtRZgkWV2SmMC38RkNTFksTgJ6EQyqD7bJrua7sVj6+l0e7YxTJGwFV8sijjUj3iZRoB8yOycCb
mDRhWXuCRH796ZmO9hKCB8bINGlAvzdwnrrbJVJZR/H3LZ47j6sYyUlTPnozlZ+sWm08Hkp2PfiR
O2ofXbWbbqGX/gcI8NGwZPAhgp1HDthYE8GMpseDBbMkqa3YVXuFv0v7N0iLvF4jwKfxz7z8crn9
Yv4CdKvxFSGpAiY8ir2iRfTGAbj0thMOKLNkxSVwdjFnWMnlpGJb5NW3KvRt8atUdVoU4uTcGlVi
bo2FPCaPUeobbTDmbf5DNTM6H4trw1JVjaAk3fOb1+EgzPm+85Joog/Uskfcfu7F7j7XVhhTgrR3
n1lX7zEztmI5oY4j4X6ZRjJjujyw3MLD+dWM52e9zdeEzW38tb2e/k6dOFtFX6GLBCy/4G1Z+3NP
DLOeXschtBXRktRC+J9vgoAfx+7RgFFHolz5HbxclSByDMBLxAq4FSuXJyCm+8TsQLKdpvvqMJSs
+AWAmHvyhWv/uRoI4pzYsbKGIwXADqGuLIKrT6VOggPirAwIj6AylS/A2jg5KoZOnX6//mBIoq9S
vDgnNEu+UH2UE/zDgKvEow5g1SnQPMpWgJHNHud3YdpBxkrbR8etzi6woj/BazN1VS9mydFDau8s
N702ulbTDFNXSvZqpdYcMj4lz4WfPFvRpgFloeeAC5W3KMyLpWQd2xzpBkATVYqWGqY/DeV02nx7
vn2eI2knlhIntb2xXNLLtJgkHjlwSWss5dx/n0aaD8DHiZzfj7hn58fHkL39gOLCcrzV9Jl8/sFu
0eCT5r11DLhrMtdACETAsRfTXYizcr38LQTGAyvWjs8BEwcZ0SP6koqND6JoJrnrtaYW0CKS34tu
46qbessFCBtnvGj9WBzyYoCkU6xoiNy1AeX5aiRfPfgDh+K9TiOMuMDpSDJj5sHPEs2Zcw4wsi5a
lu+R2NcgWyjgIMgWSOYWcJ8CNEJzIs9ETBOaYUX6WfqiKiaxD2qZ0nWA3uI81uv+jITKPTlaBYa3
KXWx3eX3JtgTQfkpaA1mzv95ne4IY30IxJ6kXq6M/cbtPw4KOaFGECgw7bme+jm0idMYtQVuJGt7
l94dAqtorJGyA/PhqW5M7JFsihOz5O0/QILKlwttcpIYpu9RD9lKOrgAdiSe2xz/DOJaVbw56790
JmNnfzdgiZzhg0OWnXkR1L/TsXRvfbKQ+xW5GDzY6j6/fA5GR7RPB6h7+EGArV9SvVL/L5ac4Cax
IyUiXEeY0ZnTFknvCsHGVdCOYuva4+WlQ/nyVaPOREJegvWmZE5PWsiz72HGoNNV6pjkyB10cwro
RNg/QkTshePVK0dsZzssWNyR+MUHGoGpE+fOomFQO07mpIfFKKc3x6FuIz5PsGxVmi0Kub2FnT6m
b3tVqKHM/AtOl0h6tm9FNXuIDr11jfkS3aZV07+Rk6u45WE4M4AfxzSVqMinslSo9FreVBrqxmGG
9O9JoanVMLSlhIMPIVfIWlMB97BS/Ad5l9R3TFGLDeXbf1zXP9d9L3TIU2Fsm/Ogh1cvJwVjwPoF
KbhYBvJA7J+WG0LeCl3T/2Syf3DFWSoeN7E8+HFkSTdHxWRfp//lSavxjVETwktzN2TNOddCvsJw
kLASqyaB4qqfvPhr6BYTYbkcybAcyKa0kAXO8op7/5TBZdFmKt58tj4OtwfJtfjmT9K/QO340Fcb
i7vuNRBzeWVpwK39AuA3ELHtert0s0oMf1tJzF73214Z1Z3KUymZ2iwfZVkgkhX/i6i2y+jxovrF
kcw6UEOHYMfTGMMHpFuC6cQWOhUrqj9S2yHa0JX+jGrfO/kCd9PDGgUQc1IIGPr67lerGsTIWlwt
9JXt8xKqM3J6099bUnD9KZjFbw+7umwt7n00Z3SSuGXq6ZeTazZZXhkgOtLYPzatMgaTVE1lrkmP
OVWU6fuweMMePuc2qQTmOsTcwcklrMtjuuY+gzbURiaxaAilvQJqmM//7kD7gfu4DUs6EwYZR3Bm
VSHvCxOy5vAdX5WWd9kO7OMix64mJd7ydYMuA9vdVNd2etVQe85jq0LmODea/5O7+W5RI816Lhoh
svxKQleOTUOH8AKFkNB0fLBqK7LMoGzxcfm6MvYLWN+EP5AxNJDNXHntq+yMHToOKs41XQ/QJV09
RGUS5zRR0P7DePmnCmIYWSrWTIVwy5i9U39UYO7DuvoNPY1jZEimZHN+SlSs+sIH6Nzg6fM3XtqY
cdsiY7sT5YSZ3ub1QeaAvl5KFmtt0XP8XnomqgfwAxftJbQewWTvnuYMqpjyI3P3vXzbkQkiECKp
rTDnGTVK4Qwqfb59zDPT1mCDqeJ4vbV9WVnK1EKMfZ/n6XbdfhgclhxN0yCxL+c+f1cyq/mqdC0k
BbsZyHWVQ25/MoYp7t/qss2DWrY2n/VHgj9s1V20hyMC+Z6wLzdCIXxzgB615s3oTqW06UQ3XhMq
XI6WSWo1TpcbNwScQlfcCDRymVwp0g5X7sofwyvY5JqaZ+o+PtkLf159ToryQ9dgvWEOHkx0RH90
SI3YC9O8JD0tzI8P36QRLfv0XSv9fs8B+abnm7ovEAfiHJsyExmsbevj+TH4ZHj0AI121AFwJoJJ
1IAgfmf3QrNaBNzPAU7Q5nYTYJvKiime3dshMhSadGGdgBWk02u6AosDLqz2IAR+xSSrFCdSfXZG
bVOJo1/g/osPBY1sjF5uqy4bOXXdjkqgapIRRiEg0N3wvXkWjSKWuM20U/Yg7FcpqegI39Cv2zdf
ETEaJa0kiDpQ6L4+9YNadWxkgLlV/Ajk28roeFvRRLYpO18SgifK51NaZh0307G9M9d2OY6ShpOz
EvMxsI98OYcd6RAEYrowbClFgqBbrZX/jhlQIcB5DPSfc/UllNEmS7gmWA3ILkol9FJ3b1XmwyIE
/a9cygENYPjVwUk8ZJVsk0PPG9PgjMlU9sJnMelI2fWepk/qAx7erkRmNCn+1YGFSfT1xCotqRoW
BX/B4Cu02NI+g6VJdP4u7qgNs4fNXN4GHyVys+6xF44YaLt/7LR2Ia9YCCk7gbpJv2wiToIZq6uu
r7THviiOCP4y7a6xoaUfCLjg9BgA8+YKw0h0PKd2VG0HSojxa6FTx8T7mhBuK7dVdY2UOGqozrS1
OLQycrMyG05nqRFkBxnO7t1bgM4mBW/mMYc8lIblOnNVBz319l6GCRuR+NJ+FTLRcK/ENitoRV6e
Ats1oA9lC+HHXMvMJCBpOk7h3VbgqBtQZsMssz8pzcdnSHd4LSMwSrv6PyBkSjxd43/d828ToJ6F
T51obdwgyA+YBW1NYA5l8C0PO9c6qSICd0mbN82S0l41CX9HLR3Boj83WsB3QVb9pe1qjU+T5qBV
Tq9Rx/qP8gHHU4J9FTybsmoTqrpBjtBUmoHnEYdAuPFFAH30ETnR8BKJOQ97bD2HE796Bt3u95bQ
/0Mo8MeK4AW64P/pZIhvKfMZunGPf6DlAT80CJi+PORFrDqB31mFYPNOK69rDt+g1m4jbS3bkoOn
ZQwQkmWHFhWj4BpnVzDVJp4yL814VvAmCbcm9a3bSeuSG9YGgSUYM1w2X/Ji6Z2iwc6hnteltn72
pgAw79DvG16q457RYR8/+fZspIPxXYwlHQqXvBageWexBSNz4mgSPjVwhD2V2TVzP9XM0DLgdO93
XbEwGLAZ5atOSfjZ7Z96k3kg9a8RgnkhjX1BPQIy9+Wc2efJFMRQGxaMJ/EFTk3/j4M8Fm5tkHlV
SoJB4iXUk+7q9NZWpsVAd4DB9SkLIWh3LBfnT8xJOeMbri+rkwxNXPOmWl/P3213/iadPAj91V+y
d+KZDnXvfWSv3p7zvwM0VqP7LdqdD6rXyStcqGLOsI4LaCLI8t3EOZKy8/2hpSNgal0pdcgEdrZS
IoQQ1WSL2sidvYMIa9sdw49MfyzH7mWs1DIF1fR6KJ9rYK/0tkKTNSlDUopxHWKjvP+LprdUt5gc
tCMWpjokFceFod/O3PtFcioBi1m+3U99H32GJV2Dqkzqh1OSA5PF7SgcUMcFRibWScs/G4mvzjL+
uRy180eMSQhS+Iw5zRSrTIaAR6UXjXZyq/jVst8P6/Bv6u3mKqHikC5fcGIuwmIizTu0jDbk+P2k
gV6+vmnZtmKTignzuosQ5zNackzBpPLbY0W+OM8UyOQDaxvytDOMTvcL56H2DuR4gPiZWeZxvpe6
vdFpz5ugNVIIlk9cx+GgbopBjd/sK0iVY+5LCDAB0mgB5lDW7HbuKLSzbKORvkfIL1ff9DTtxqqu
tc0HOnm4KklYOIm9KqH2VmYj8J9wps0jEyDq/dje5R3jzsV6hBIe6UCf+h5aWGsc2GYyrDil4LCj
AgtKe4HGW0mgKIp/kvRo2GKXsWo+TT/Q9n2mcUGYV+elI+E/nOM1vycl0Tu2ZNMLeqiZ3HbWye7i
qbI8qj8y+TicFKBd+vkuErJJk4ZgyDubN+m4oba5ax+LKVSYMmwR5w2R9ChhQ9w23pfcSqGtyh18
wi+lI/uVRh4/V5NcNE3N3IRxiVlEQFgdrB8L/hweAXVfkE+6KRcgBa0iUnlitVf9V4r9h/LjdEee
1KJDNBStEVBaENRXcJjjjEswXli6c0Rnsyz/XPyV1oqHuORa7qp/JxEHR9R7uLCetjO8LdQJ7MZw
0xAiVlyK7RU33G09RPi6Q6Hr9Hh4KgxPCrYRzEORIOfSRxdNymgFG2ZFanzNvxzXeXarvog/q/3P
J67I0+YRtzVwOzsVIPJ4cV8WJe6hXUHryPdlY9NT4I/Zm3r/0tadDjPUCj+rBf0pYmTctOwQsjXf
aEeCj4rgxUeAHzIgEMcdZqq/66o2qXGwwrR7+bSODeOpjHpSBHGe1248rq2sy15SIU+ezfyVp5P4
7IivBJmedIkibebI5JviRYgfl5RZ/XPi3OPUjpJp9yS3v650d5ECrOucx5z82x8K8GwuoRB36/pc
uc9ihB4aJah7jwN78fRTEvy8Ik9SXTBuB46TQ77i/0HLF22S2CphZ5Fd6a0HkEgzc2BaIy1wHYht
xoatfVmMF4p7OQTwuw7sFV7h4gLgwpUiaLLF9SH08DgTwUkvwuJIa89UpdwWTgWUcqXyEz5KsLZP
x17BRt1cMtzTkOfQ0mGzzrQ1TZ/BwkoLREa9jwHPP7l3hEo1QkqDJTJA0PUtfukgXwz1vvYWXdg0
qcYDAMGrcSjgEw+wM0HKlbELwNFLQgs0QonD5kItNUKsrr3Ff59+9XhJlDXnaHlJoLsxfzMo2Pjx
DAHwhxoA0x1fZe4G8wOpwD1VjYgA7+UVIdGcHbGkDYgiwII1fICPS2yDWT+dMle7CPrf+XeBKrkl
LzjAmmamIIPZNmAFc16lZHuhi2PIjRqlVXRXaNlTbTFd4L9Kpf5o6nRIMI1cV8DlWgA4P6mHKNLa
cxh6ujIjHzLtJGJX5OKTNs9tbwsOE1ZE5XgF7FWCaLoBA2sHSlz38agwkxG07pqJ0lYPUEIOVgR8
wCcnwq75bG7lC9cXJ+SaRjGR/KKsF0FXUl1m7+gbUeeMuPePcM931HDX1FcN3J6lTLAwMDgDCPer
h2zNQ99foCffO066RjuVhp5ToKXMW71RYIQlg0pJAM40Z+lLT21sJjAPyizOVJ/xQ9/tGI8BeFFj
ViEFRZxolK9ikqZYO0Z4x961H5RQUWUCf8QKy09NdY3XbiSYojdss8+aRIpH9B1Tze400cDAklKj
ap/oLGiIh32TT3dNt3JHKioZP79vTgt45kHe73+PlWjmpbBGJsryMfYD4EdrFInFSIg96Fo6Pf8x
++2BNX5FxADnxhDGQ30ypqo40a71eVflH5kXuOM6oEUcAbDkZiiPtFRhM4rL5QFuZYy9B7joeNiX
JwJ/AB9ICEuZ+U5rutCU2kTlaGm3fD2yK5EzJzL/8zFIDlFSivGHY4EzgDj0sd7CyWcjbS0YmLWP
usZR1588JmF+9jzxm7iElFoqQ3C376O7QBfyMII80HRjZjrndOIZHja7k381L2QW148QgvDXgHOW
AQXA4YaD4YBeuHF5XiWLvRbvz9cJt78Q7tyWTHU3SAYUwRvAeejxRuOktbcx2oaSLExvEfmLIcrI
K06vUXG0JpTNSHRVl9A18Ybjq8+9W/Jo5lxUNQ0dHRVxvXOWUrhyD/SA+vdOeHExwgCpf1TJ3qXE
QL4y28qwlXbwF6GmWbOQ4svDiYlfDiiweuegzVsnkLy2IfRbvw/kFCJH8RNK2wgTBI51CADLNNFJ
RLg5JbfsNarOoORAL88ikCe7lIY4tjlvq5MS83Rnf+fj96U+LS9i2PFqGrXSGbksGUif4PhUwee2
AvEMo/W1bxl928m28VyZoaumxN82HxcT/VtIkswQusp1To+4HWvq+HTMHVF0lkZqprJjq4WEYdaq
Z60ab2WO3UBPHyGqVrRZv73DhkgFTEDUBFWWs5Jkw47CuS2A5omhgsYd6JVdql7WhFhbDB2q53Gp
olTJHB9Ofiuum25/GOArLomveHb9qph+QpiCOR/61iBLz047sdrPUUtvL3loamjCsnYGlHGZS7za
lG3wPaYwEfNAdVbicVQWB4uxWP4ouJura+bAwwM1EPP6hKx34y7O+0bmYUX2ywyyCaL29ClrBbAv
tyFlKTB3xfpgK0a2oTlOHDTep1CmToKXH++hMsCM/AAnots0ghPbaCB47N2R1uC0y+h9Rq10tklF
8VIv136p5j1E1j4EGaDte0RQN4PKbGArOG5frybgMXu2c9G7f2kby2koTclvge/fpQbFvoGgAH2k
hWSkZDL6qwbW6vnXIXO54EXNoT+daIv9c89m4S6NGufGMiIbIym2gRFxWus4dDTweQ6dX6bj2YQs
IBPJclbtPQcCn/VOufF32cYsUosDd7JVncERDp3mJK5UWMpEfrnKO8DQnEwshkZKG2K/kKzYa8bB
ibLwZe+YI+yTRHW91fEI4pQHZkNRJvCQw27b+QIVN9h/Kf6iBmBYHg71Nm88ix3W5mtTYd7Mxo+5
4zTOuVrDul6QnoFVtODeIqNYZp/XshaMQfFbh++nI5LNbNgSnJePt66pquJi2hXyztD8OMpSHuUu
BirhMdoVeKAfNHdjyqAulebn8lYz1kyX3+cFOe2bDGmUHA8lcRfTu/XJ1iXLFCQUlEwoTF3KYIGg
mi3uADufZwz/12/oX25nczi/tC1VeAHRcwQAQGsdf4Q4VxX8et96ODa4SS9tBhzyoI4zuAWqMeDE
pHdwiTf8YRZJASMBTh1hyS72kTKD0zmJpcQUjSp2uttBvS93XvBuZ+e78EAAS8ugtCYe+LBRVoAC
s7ys9bPZd97VzE+p8N1vVn9SQ8fhC2OK0gKNUuRS4Eta8NbFAEnN9aRjzKapZRGpteh/yg+/vtBK
+9vMnhHXnU8eeSGWfu6ACXv+t+Cl+ZKj8BDf/wREeZmLDQCxXQ1c0HYv7z1D4ZKJtWWoVX4UmN1e
Xr3gGU6QbMy4YNfODs2YHVRYMSZDBK4m6uZov9BWXvHkbMo2dBcij2RrI5icptmgg3F9EaaHgvr7
SvLv+iPaA73WCRW0Ys3jDy5tOp3GMsdVAXdCyeTqTYAU7YXXkCFIp40JvORQnbrb7/RGvtGxhqkg
O00igf0MqDogkzFE7vE8ymO4YAHOG9Ug1js7V6Y4mU/Mmzdl4mlXGIVZEfKSJEhL1QFYMWif2whO
1iLwbHovtg4wVZ4xCOWKkwELJOKbtR6b6ow6NKtF76yXt3VFkDEkoCI89XTsZVsTlxINUe+mpdwq
8PBUVmYez/zI00xX2XFQnbHh/rK/PBAZeipw5JyHlbib4dtUNc6fj58QmrwPojIFfQs8wEizX6C/
rbzduk8kerWc+zuJaFHremF+RSLbgEff2haVZKLjYScfCL+uF85pCJmFAibKLt6tuirvllf2xtUF
5rM20lWyeUdw5S0PQQThs6K6FKRzj4JNgBJlrWC9Y5Dm3WAyOPvafLICsS/jT8S9zlW+EXOvPFXn
gFnSqZE/WSEkav82E1xUA2OG172optm+NnMfe2IUSkEmn4wNjgIfy4A0/ZWbDxJNao8xKgsdZVVr
jhy6P+yGojuNKP6rrJL+0e4bvsD6vKNL1WIZTOuy+uvqFY15tejznXqYbJoDTDTuhvVp4qWAyMU8
zYko4tcr+0eFN69gxBfqXmNHP6haUz6RuVqN+LZWROgAM8dFHZleHD+Ejhs7Wutv/guH0OjH7351
4R2DVcZIkIB7i++kYDADgcMZFYrEy9NnNYkELuUDVy63pkg6wbe3Ajb772VOVuLbzk66lhioWvvy
d5VIYgFDO1f9t7NVlgzDvp2Ra4JHl8zH+X3X5kdD9JhuR2JbI/KnC8wzVww2v8iX3LXye/HBvzXX
cTIlmUk1ygvWqI9zNpXG4qokiuZvzvsAF9U/7UR/bctvKAdL/pi6I1xtanfHGTySjDSlaJXM3f5g
LgC66yD2jBkmUB3axewu8WOPNyu9UhNVk5zrCBmX3rWNPWcW2abz9ZF78SvZV7jD1gSp/bhUQaHb
KScj5IgO54aUIQS25+MtmEsu/NVem81gjVyG2BIeTBI4x3EL3M1ztP1GptHXqXy5hMR/tPGkiUF2
A1QIX720HgwYLWM/I1kb/64z12b3skTlch4kpByXPTsl+rY0MbgL00AFlDYSvoz08LydFdHRCnFa
JeVALvjI3qhdSU38FH+8hDBqxPKnGnvqnbUjtTDEkmj2d2h+aaLFoIyKlAJ51kVfXfeKKNPW1mbg
V5JyYyvQ+iiBUlxjakRowg3LXLzTRGZ9JSXkUZzUlQz1JwKbkMcFdq/Y5DjUuD8JRh0USMnTIrPT
x2mdyjaie1QKD+jO7F9G2RQWOoxU4ZYyV8UMHpxsfwLwizjxRF9lA03tmTSjA3wmi0kPvFtaKSTu
QB09e58h2EaezF8a0utva/Le3NI+lALugTqRNAkyInVB0s8YaVLMl+Oc0EFSxPvft9d1Alc3HgU5
n3I+dN/s6VujatzUp4AkVKIIrL8e0EjwmyP3oQghHUt6d6iH7zzFsHhGDCHyizUsoWRjIPURxTTI
YHbn9pNXQrwlubGFO9OY0GphSk7xDj/oSC1XPQNw/Xa9SvV/sQ54Sf6sL0hs1ojsX1e1GqBFFDh1
sMd3fQkLtVCcL69hP3m8e1Vej4AMF6vNeYFDu4A4TFyXhOR5RLl21Vo1YfKQV0Q1MdCgn+bXjIK9
JF7U/OqXFkYsAZVWqh24RYEN72coqwNkr9XqfX8MmiokHMxYYk36tr0ll42nb3+4HKQp3fpCLz2Q
cUrv13DjmjQm8LW4azuQ96RyH5d+dvnuZ3L2q5u8pd+xonVBAToDDmWA1R5pzw3T/+K8JPNo4wr6
w7cNlnAGMpPQPvLLOpIDHj8inXXzvN9E7lc+s57g9IPQq2l7eZhJRnlqdg6HP7WGK3Hxro+524o8
dB+9ShxRI5fHET2xuzFfm8In7GIUmcM9clhWqx/u/QxtEhw/OPgtRU6e/611optIfA3WfumZemog
9AMvGROVrqtuqmqiLlE1CJJW5DVCLOiPFWLtjhHnfCatU0E46nQUevuC83DGhJE9Y78jnXYyiYVT
MDooTzR+5BCF1Diin0JcQST6zpNPhq/DAoKumkoW7P8jcNsqfxPj9fqIesWVpOE5T2qVm/jLb6zq
ONpAi65yVbYSOaPVxPKsvrEQsPUB5ijQWQ2AUMchBhiNG7ZewqzE2d1jRN5yUVxnzNay8vAzw8C2
sROsHcBSU6sjZ+zc7Zk1F45zz5pzWJQ+Z6Ensm0pjwz0AZKlKbxPLZTv41uigIGnCDqWecrcgYeJ
dFruJbNYRGyi4k/+obtvP7ZShk0SToTttgnvvlyCelVqd5NQt7xmkcvgrinBt1y9QExrRaI7RpYq
V3XTpfN1qFqZY+YoFuz/E8Ze0N88/LssBVcyJIQeDJ3Q+24NnY0qPCVHkO6uV2E0j70IIFJ8AXtG
V127ZM5Z53orvjZ36D/OPAq3xUgWOegq0GHXPpYOBYP+dR5cCArVCGEOtQeJmtXCZ/FPbxPCRy+M
jiU0gjJ4FDey7X2VJyG296MvXQ2nQAw8jTK/VMqjNbKYn+CSKLY4EBASh+bPpAwz3vkb3jpGr0oI
il/8R6FGuOZF9nIjJHX1GU9pOA+xYmHS09THsznAII+3I47eh6Sji1gXA2XAa7hgFg5xRfkw05B+
J/hHI87GrWzLhdUt4KYmpx20fgzWiWOd8TM2G/2Dmn4u8K1hUoAUjwDEQ9aAGUUg92jIZYcpqMRg
shicRBgjQmIovO0aI+3QukKF668dgIWe8TdsPg35LbeUSXTVR4+srzrgtbIl5fr2ZUzw3Yfe4ksV
YD80Ky/ug1+7FvjgX1foid2uUh7KELNUlkiPc03X5jx56WU1P3Co7mXCXPFHK2ngrlMPFpSLo1Ml
qGzUlHATyqKAFUVgDwS7bPzi5lyabZ+PkU4IJVJFGDbL7B3mU90f+87KGIybCs4XKAJGdRgMkl5W
r7BAwRRc1ZgDPJ0qW51iIkCOp5ARU8dWot0l3JxG20hZB26NS9giyhT9eirzUcF7IQkyBZrHk4sh
5K0Fkh0WPUs7PAyVkdQRev54ghkr5p3UvSAqvwvIK7BznmZsaXuKhDFZ7kCpzlI26IUsTTqP62cs
nejguKHusmoutnoHr4YuezRTjWSl6xJmks9qmtz6f+p8rRVTGAD9ctmGYNbnMeSV5I+hS4STOqWF
tBxhfiBYhonGslOEvk6aMM95btQcixkwcjDuSAtTV+aSOU0wn6b7PF30A5IlMchZjOJ83RHlceVY
0W8tEL3LlJvs5bPv440zlkl0a+5ctTeGV6GqB1cMLSmwYKjhYJlydz4SIEAe618p8NAxfCVn3E4a
Pf/c38oI9pCb2rbuUg+/TseTmCb119Bz8jpTl95F9Rrx+4K39Jvz/H8bLjAgMdOTh5Iachpvzk44
x5YmA3feH7BxmSQInVDpjstKXVWWKtbnb3eCMA0v85L59BJnU8EiBJTHrFtWC2xDP0DrWYvX/zDy
nmvK3Is/Jr2Z5+xLsIxWYrVTEWNT85xq+G/dM+PVTHsB7fhKLZ5xVKuN4obodtn+WJXIidBFoFFe
ZUpbwVqvB61aptoG3BbcwHFmnsiFp/2O5SlSw3prP+4EhhTyNlgRbR0u3TCAexzHDcdsN8AGAAIh
1KmJfR07+EuGvTm+Y6Q4acRjtfHE2BIT0817PuNQw2/IUK98NFAoQ7JDwVA6rF29uKeR0wTQWGdb
QK2iox7Fj+82igcR7+/vQdwGNgZKYBAtkiNgZiV5WJPl+wPjL1o44vBuMU1Aq6UBTgRirM4bMl98
a93xvOK1OnT98Sq+Htie/MLzsfr5k/3Vyc0eGanbRRHw03PaSwKTo8nc1hkEgoj3yldtyvcMzA7n
gtVPagv+Rq/AIsWsu5LOm4NATBXLJoXJWZ+qeQBJb5eAQZPJzJeapWpihRNEWBA87fGPpadz9a/B
1rPlwOuwKvlIbrdKgKDEHGvgXHvq47ttdnzqVKwcZKypVSHHDBBoOr3xZkmvp10r1bQbj7dOjJ0e
cSqDJUhyrXmemSN7U0obcZcV85/O7OVZ3kvhwit+Slsn9myeV+0Ki65F6W/XPLBVxS4MaXULSBT7
xmcZLlDOvHgwNQzM//qfdH7qV9EsdveVapvDqo6rULBh8DrypFTvxjdetE9G/RreGebyw+QyYFlF
uE/k356aShYGv5qUkTzZV1tbQXp4dL34QX7epX/WlGEWWZySlIbjKTcXn145UtL0Mhp38pFBmdAG
FicalT+mA75+vohjpqaQ0sHH0/YVsd3SKzID3lWo442DnQ/EPJxjFrqsWd5XkAADCHVS6ypxzjMO
MwbN8VHHnakoy+zi4uUJNwGi+SdeSWj0FpRAtnMfiXBiAfl58fTCjqnw3DC1TSXdBJGYR9ByDPVf
ChWYDsSDX90506B2wIjnJ6aFgpLPiLivt4zF0r+iwAXOeWgO7PyPjLjBlaPyZVdrMC0J5UoZvvSj
aSQEqwAHzjh9uKg3RY0mF8clfUYvhudvWme/VCujTAxKrBYfK34Qd4Zz4m9L9AoG40bLVbKD/I6I
f7oE/MgIoENbk+Tc6g27dzejfdTXBr9SVECcrEUJ/4mDX1e1z54Y/whDeWZkY8wkEsXtrBqowtEV
L2bCZOKiYaPmsnLBjoTcQkPEcKfSfanGrV/5NqZB/UoDYmukCLjDhjCIYwYV4LvErjhJBefuH25p
ApR+dMwZjyygdr8/VrN3JDi3e7MF132wgw3rIDpiGm6rqWsrzKJmL560H7fQDQ/Dmawn+0pXoLAz
h1z/Tsnj3eKAupM28FASJ6QVQJComVZkQMee7qLNvrY+l8kQ9pqTqDs0Tnj8pbWng8aJhkEVurkh
hH+vZGwcgCwnL/wHDB+0e2Y/e9Li0lRpIcnszgwo6IDCUnJ9E4JUH0Q/z+xc5Ae4hepQkWiT/drX
LW84SBn8D8jK7QFWe4U9R7uQW7YGBuCE0h4zabWw8QmLUmOsDSQCSWhQH5xx2j8tP7/eBsXkw+5K
yBRfuyIyL9TPdcS7LIIHKb0JpEmaRNz2C5WIWahzIyl44BJCJuM/3g+24UrPDSi7uRnITfICYdn0
YbjuwXcf/Fre3cHYn2oxA2kfAJZFU9Qu28I4REqVYOSFL4jeUMdcANh74ZZ4inRtjUDiL9C2OoQ7
KIr9K+81jQrFMXNOk/DzcHU0Sqpab7+IQHE0Uz8Lr3Eq6wApUXwghWRbJbM3XORfPFRrwzy5N4ym
gAWjTaDLjpOxv/VKwertJiwJi/r7vnC4CUgqINBndeKDuEq10mLqBXg42K26v0aU/9HxaixBMzxW
3RhH/gKwyztRfW7FBH0PKK3A5Ry/HE6+e8ylRCpakdRFlmBoVTrqDedLYjCvw9TvRuYQuibRc5db
N2GAqx7bF923NyN4ENEaEFpSK7jvFVyjy+r9tbpQQUx8eqAqRT22lAvvsk13TrKe5bZqmpLD2sng
0I9K/ctdHs1HiUcQd+nQDDQnTjRCwJAuHkR2OKzhxZatGx4/JraSWGKUjfmfX4qcppfn8Av3FaJj
jOQagvP9KmCeSXv5ZVxCbnAUKK9Sy4ZJLPvSuB4J6qgOfuPWdK+Y6PmaGNyhYkYWd1Hzt1DZzIwV
lbtJmTzqR3uLc1UnrGnLbLzBYWdxV9ajGPmKAlmfypvh03ilnTTyhmp0phgWrZFkdUjSFJlCBQJI
HaOuRYEUqeV9gKqo/RgZAu8SY9T2O3tl+9oTfawQ6pBOa6/I3D17cuhVR2Ky1WTQBxxOIZewGfKV
C5mwl/q23L1AjI7xPFL9wV2jZ6QPnDg82H83Tn+A66a2X/uSTuNiyjBCBTrTnqzYrv6Dy/3Cavuv
t6DVtRv14g3++Do/1HMVSf5ycQM7xgpMDJ/7hedzku7lv5AFEA5V2sFwSgmVXg7bcGWuc6mzl3Ln
aV3kP7NglPShqawSUfIyh2p7PxQ2xAa2RMi7HrcxO3u8FvD61V5c8CEPaY7yACXpR0H2TQ7s6rYg
4AMoZ3YaR9PDHWEtG4yJcscyHpoCtjekaBbpucARGxeQZGNWxo8ceMKWhSgCRNe1pgLnnSlzRyjt
2tooTbRK6TxKK6L8u3X9hs9xhBrEayXQzdUbiwxrbsz+DxovEV36pFa4Wxd8QrC5D/HoRLOEjpXF
1RYQYo29nkI1TrdMw8iZBH5OtFRdA8cotZwqu+nRXHo6RH2rZvjR8Qb/IMDbeEOtY9BrJq/pGl/0
qo0BTUcok/Ueoy4ZSer0JfQwZGGXafb7KfIMmpcH3jRXQ+h14a1eO1+iLUbZYVoNxMvRNlloWk2j
h4Llx8Oxhy2BTVqZpOgH5d7qH0oU329UwChsRlJO5NgHzgVVfvdNxfWsrYeMHhhz8ZBxnzvtZP8z
fa7BpbDSLiNsOO/ltNFKh46ms4ANZHQ89wHhJpjV7ddy4ahBrSCqQyKZZ1JIaZR4a3nq0Ldo84pc
Vw9UEm1Dbz4tsoy11R+XzxoKjUD7h3tUKtf6YKpjULFZH3MnbUjtJyWNjWfwvjf4zGaDXu+HqZzb
3HAbA/okptyrko5cv61SkeqtufdC6B89goa4hA+XQ6hJQW9UjWCXGt1+HsxCXB56YAoc7Jw38Ti3
aCyB73e+48oc7+zSVJS35nFvH3nRUAsH3md7CBiTJGF5glYIvpazR+m37JKo8WjxBTHY/vqpLDg+
6GlKfCxYx1cgf/5nHTSYQmzujox0+MizL0mnZlUhzLQIO//x9d2SXBnC+L4/QKlN3PB5kgS+Px7I
q4BH/3VGR3AIlKjSYjburXBNJnzROZ9/skLVeiyAugN61ownOUqFDYCuXPJqqZT5ltH1FpSot2OD
uvvegtLiCK8MEKMABT6id6HWSyqglGbKXMAbKvqOdjkkY/YHfpAxSu0xW1ObMVO4wRgm0PvtqKy6
FHIQMuMmLf0YEL2EGZgyyPOL47dp68FqeduUNXeDBaoj1LeVnlZaO2gXKnHxclGXAbcUZ1m6zRz2
iXOPkOaKCosOjAWmLHmzAzTDbosTV+8MCG7CgnIPdbA5sueHB9VhII7jsKVw3XZCdSxInkKkN4LR
E53rktxtzfv5Vd4Ge/LanzU72zABfPZkxQbqX5V2OIJFWYBCukydHvtrUsqZWPCUwv1OOrEF57zq
93xRL1z8U0YjwfjCFLqtBqDiyYwPwEhdpofsESNk9wrWKut8SmM93irFgzvO2S73I9ZnvkorQvTd
hdL3uuGlkc7FqGw3EjfifHcH9InqhhqpUoCFbxAuXhP4+2tj3YDpYR0TveDJy/RWWoO89B+b2zWB
XykDyW6HtxRKgc7vKxF7HfSVyhth5W1qjTvG+4uxpWmE+6or0EEd4uLL0R+95fVDuszP/A+lM0/d
1RusPleAkYCSyHj8fV4QNzET6savmwU70chLCob3W8ztKvnmkDEnTUNzZBR0IuLrRxnogL7E4wjF
6uT43gO/kAVG2nQUuPJfcqrxQH8+14j9MZZbDIle6aT2Bk0zOXeXUu2Blb6i9+9IvbWqnMsUjNLt
IGvBkzOcGzkV0XfVnOLYoqt6rSWPTaWr2EVARyU/zQKw1XOF/D5tLRyfbBwqINALYwEnmlZV3bHg
Lp2d8foqN7TzIHcfDFyJjAlZ766NvZypo/IKhr4KjHw4dkTg3dcc4RXpIIyAY7HYC0WQHKOH0jFh
2Zmi2Cy/aNxcqBzKP3yqU79ItGJ2JCwmq3774myEaTBaijyq+og3OUps6/QZHVOHE09rV116OLAQ
XSFUj5nqQtPXbatF7W7bE4pDo7U+0VrELzIKC3tGjUkD06bQ5FB4BEeSPBSN8idZgvIl4HINlw6Q
nCH3xmfpi//m37j1Wb/f7BvRIeSgU6tUcIHqJr8DjbXhLMy+J92XYhUj4Daob7bFDJvaawUJletl
Das1eB8NqT3VcvKre7yf/NNOlRmw3UOWQAlP8pBLfgBB4Uwp4+vC/XDbUItIMojdDeN1kvDBVYOl
pVL7b0QyJwb1ixm9O+WtldrmIe84ceyYfHA4D3KgqVH+H7jSr1ix6RxMgMN3SyDUgh7FnO39J5hO
40fMPHVRwKqh3LWZppqV4idzhrKaJNmSt5g2QE9hFq4ecjFSI74OO67awfmCpdBbUut6ByYIdao/
mASHjgafXPYWJf/stXdYezYTATM4SW1LdX9RJYtk1K5KGge4+fawdhNaeGCuUx7uhwIs0BF072Se
y+8+ZctD+thwPeYcBNQU9V+qyBgZFaeMsEyP9RK7UTNH4u4XIxVliqeZvvQn9vUZSLi2j1L+DJ0Q
Yv/LdwN14VIyvhZQuM2WaWAAu2Ifa9SM2Ktl8g41myvKALQWHztqZcgYioa8uRPiRYFP9wll291e
BzyQ5YVMn0MNOlrZKmu2DOS3b88V+f5W6TNalDNl+c70m2BOb44q9DC+KJOuwIgHf9AA5csdX2MX
l+0bLP5f6zjVQWOZZC1ahiW/imS9ayYPibx8R7i4FymOV1bfeIyqK2UAGRY4EWdVbAFEsZOnrp+E
QsdHjWq0KJiUN1YuQ7uBQ6qnsV3DM3YWeFaA4fqC2BwtmjuV0VX0Kyyc18DLScfN4Le3b4QiT1Fc
vyMffOhAB0waDjO93zFyA58g0DvqdJbbfAEw1EV6zWA+DtCXiRdUtZIfo+PxjR1Gqrp6uC30LLmP
Lr9fzjtnzqP3VXnZ/DG5xAJ6I6pJaYMsLthZZ9i79cm6tEaXVevG6yU/C5R1zJzzR990jx3PG7Z7
3myIXAP+vs8AHvYQ7TbSw4H3WpyDSa3ezI7RYIxjlWnVmku7N71Lr1qf2a++AnHa6OVhkwURyBu4
ol0eOh5NLZPCUheOdl4fPd3i3JamVL6MFGNdS69WkIE3NzKv7/4W3VNoxpf+cpSVhWGPjPYiJ7Aj
1VFmh0RjEoGbEmRlObc78mUj09B7sKSJhlg0vTE7XpcDePsDUwcQ3ZoqpdFPI9GItDJBlnpc2tQA
5BJF0Mc2nxaFeJaMR9C+gCTE+wSCQnl+00eiT2tGyz+G9eylRwrKLXh6THlgGPnOwM67ZHA3qUXC
UoxshGQp5ye9fst09sjDKrQqcTWCgAyvBL5m3UxfdjLPBN5jJnYkOMI6qNmubfhpHMQZqEKh/yuO
mmjaN7iYhdV0a265xiPoKwdar6opcDavW7guVOfacesZ1+tJGzD2W0W5nTz318AwJpo7N58FLDoM
rq5YVvOUkRwd0HBMTcBHEHVSnXnFSEH7fPwv5tYk5kB0nUnILiAArgBUP04fPc1mflOaFMkc8p0i
B0hSoEhEWQQnbvq9bBwVSgdOGebFhjDR4wOqFvPeFN5V43ZNm4Xcx6BJJuRvWA6I99m1febCo+fi
eox3944mO/GmbiLfo7vHIi0cbi4vHphBXfJ9A14jJdc3Ahx+rRAl+vV9dsQkU0h1m/Rhqpd8aM65
JbIgGfAXbnq28QAKo0sdxHl0QHhak+C4jG58B/HmDPYqyKW4XL7M0oK9I22Mev5cMj/7G1HD/Z8r
gpkTHboNrnpIzydpbEQMu36lxI7C//wx9FqYygPMnPIcY2vrtepnz0rL+wsiyOztvuGHNp7mpFX0
Rf/zoK+yoQ0GsG6YOqB7Pp3V51rm2YU6Vf57tj4DB5JSZ6IB/GMJIRPl3EZzaidoW2i0tSZ/Q1Kz
Otfy5DnfScwIhmiboMwcLWhYirscBSri4CDpY7Ni9z9Vgt1Gtd9WUvQkQ/1LDd6wlDL80VwvY+ew
Y1GmUmCWFNoxDHAVkWxuRYXFGmxwGRZllzkPmXOP4VcUCDS9LVoj6uapAv/E7w3gK6/n97NKaRWr
yxkJfHEq4KoET2Ul+5c7fnYwcCUSMiFfJlFXPh3iOoxxwz1HbLVa8eJCfcf6Vbnd78dxQP5YckcN
KrKtRxfEDVP8CQqu9OwITSJ8qRENoi6xLiBXQMh55VxC/5jpNgLjipTnt/jGVl1OqKyd4T1gkIoO
Psxuuc2i7a/FR3bcq7sXyz5IVgpTuR3+z3R7xafRYI3b9Vp2wGao/UsxjziBEuOABSeZnQ52di1t
OV18lxqrt3WK57wBRalXI1gTZpM6CdwWDv3kOmx1RHvnAyxX/BrwSwaelC+RudXe4aR51/zT9TdA
KGSDGZl8P1C08b/kAUdCb7yKDvk01pbpP12UzvG3J+jzXGmActXP4Mo+22ueCwXoWw65SERgbi0+
31YXaAar5ZpXEtPQ9I9S/e9A2+80KGhSgWe5+sEehLd5l7gvrIp4/D/azUZ00t3yStFOsCmfCaJP
egciDTyqPKaCgeWa8kx4k6OoQFuov3bANBsuyRszZSes4ZZ9E0N6RymgpnTxvhpop/0ag1A1LoT+
lxJlf5epVv4vGF0TXPSYfsfrlMLjmZzBKHPguz8uQfAU7URuN/2Zrzi5fm9UjfRySeA9PxTf32su
hjx5X43yATC5tge62e+uAnLSaegzeiQcXDpvLhQ084+Hwc4KwzW5pMupekvwC2hJXw6cbA7OoyRs
XPnGHS1hRxztm/KqRb36hKyrchvvjxJM5AT/kUL4EHC/+ckGp50mAl5jppr3/2SciliDPnZ0IRc6
yJhKfeHGf1HBmW76P+IsdibrWknn/avapz3UlOlaQV1iSTlck4MfUhRQt1VKU8JU1oRO8hlPQEqd
/U5DvoCR4h8MCLTFQ+xyO4S1WId+d9rgnavr1RHSeCO3tsjQv8uDN1/31GpNnKl9djVSr5uT/Jah
nMx4avJJriPYhYROhO46zHPvsVN7DZ9O8vnwmKGHWqmmj5DeNWZPdreVi2qOo1MFHaTWE6Qk9p1l
bNUBmk3GzpFJQq1/i5ij+tweeKnymP6C4mH5bLe1Gu+jDBenlu8S3iP5N9W1/6OTCttVp9kBBp3r
8RbkRf3oQZ/sBxQqwge2dSPnFKv6LY5xvodOxBlL0Rzo0EAuiXTN0bbEY3krtFtUv6Yp/z1wmzgC
thT4tKKAt5OGKUgt2bFkxnuuwe4t4gyUq8xyu3zFE8EjyHOgDlY2DOig62zhmecIEP01BRx5o6EU
WviG0MuiUcW5+gn/mbylwyQwke5OiA7ZuolbHRJow5V2LpkLWJ/ZyHTv6wuntrdLMr8fWgfpDLbT
VNAlLXKdQmUkUNaHAJ1DxCcQo01z+PnLOcad3tmumK+k3PR/C/wTc8WaCtrioE2EgUGeDPyNJ3FN
wSK1bC9DSOK4fyrx3BROCESOnhh39f9Mn1Nj2fghaf0vanUtJjw2deWZxKeL1xAdLwH/yE/8uXNF
VivNFd99gQ+y17geDFfkpaN1DfNbsF/X/h0ayKc1UyYTaFdg3RaDaXNXg2gQk2aOtjFF989vVwOL
ytiGCvwepo/o6qDJ8jBDK6uN+rc+6HuU0bvDw77XEJ+1k75J9x1NSFE9x5D45tJMwa+Elg67R2x2
GfeoO7AVYNm5k7DVfWdQ/KUmVu82vFIYOv7RoMbyI4dw3naDdmBYvaAdJYpkXr+4QHtx06DZNVGj
cNUbkN8bYGqwhgYSfq03UmWC1aS661GlleOb6MitBYSeohkhz2GUOCdftysMeg9dDb2JVbxn6rQW
U9mvryDSXqe+3DYvh3GQqHSmCTEQy3mWN+vO/c0VZQvp6hmwYe6pf+6LOPOv7XA7pSW90fRdB6qL
LkeGcvAoNiHd8GY1oQCsAUpZGh3YBIhNb/ejHedesh99H6PWE6ut5xVhWjfsk/rFIa1moOgMOUj8
GNsRsAUi1Y6D2lgYCCSGvLgTJWhsTpMQeJgEvFb/4tVU5YviySEkY055q9UxtbF8w030L3MV3KmN
mGQrtMvHdecN6iOYngGSB5CGYMD/t6s1wnP/AQeQuKg4upVOPLrGrnl2pWz60s/02wnyB+Nizl4k
Sk0aEw8ITlH/dLnjCMslUSnGOk1WkBuQvRwwLbDiz+BT4XWMUxTAzW4EAMDdH/gbPkSUli5/73GH
0ghoDdHpt1VyMNZWep2chsEKrU/7UOVTb56AckKHuDOYZlcC9J05ixdMrK8+U+kxnpIP0buQuOID
kSqJbslRR5PKd2iy6m0am4caCw3blwYn1bhtEXLAK6TWdXZKiJu6G4g3gxHfx4K6PPjL21HOXof+
IU0D2+i9oWNU2QLjj2uzRJOZ2Lw6Xn9MEA1w23xS/ue7daBJdFVmq4zi8FI574EHUR7Nyy1zJjcu
Z+fFlE/gb20H7ED0GkFoQpqh9VWivWJ4xqLT2zJ4fPYgSBJGaOVtYFljGdMYjQA64uNJPKDmpQ14
Pwv3pFMgTO+T4/w5WAc5fzOsIoNQGZVjI0w1ndhdBnKvjrLkpZW5GK1CHgGTPCPLwgVf8mw/AaaB
32Jm17oKqhKSBWRMqPo7BugBb8veDDRpyEwhIVeMoB5SLYUIk3dNyxMVwXGHA1PnzW4z99mAGW8h
2ObfCTRMIQs8WJfunsJGcsZfmtueEfDXTNZFvPzjhjIoW8etNpnJIxQ2oMN7ZGYoxIV6nJkHbrAU
2v9x0EBTpaZu28HFYoCCJhLHc/pQKJ+Kx6ERTOgC9Ab7KDnE4UeJqivdc5uxVbAWujJtRSMWumje
A/3EaQTosDJDqQSdYzcYG41ATLOCehbGe+bG9s/qI39j+xs68EeLoGxdAI35BQG5sq2+OdOLQZS2
4/hTquqCvhWKvSBpM1jzKUFyk1JCipWJejDR8a4H7qw+Wt+ds8TdLTx5eEQlLAfc9oVUOzEj7BBZ
j43mtpEe5On44rJLA/+oQC1+mFqqQteewOc8fym0M8ua4K+PYHpNTllKykf/ENJUFDy0FEXgcGQx
Qq1mTEKVid6dCAwRHknKak2mZdNDdqH/2z9Il9morfBAIe9wsGYRxp9B1AN++mwXTu7T+e1vFvvn
jc6nAsq7j8wlY/MlGuQay1k/Zt5ZPJ/4eDrEK7fBXV162qrHEQGdDSdjjvMxi4X2H+FvctJ7Sfbh
amtwhz71o+9pN1oDSSneVKUksp7lw6LnPGcTFbzh2e7nS17flrboIvERGLfyP/Lh/oJi8cTUOJec
jBC1w0sbR1Y+bC/phi9/QPi22GNoIB5010zEoyJa1N7QufLeJAfMmmgSR14cRBuoxPj8wazylam0
WfSvqwJtFcZ0RchRCNYUBlNNgidbUWM3BQ7asanNdeiIZFRByuZsH/LY8vhGql3W/vVvhNLwWoFd
OEqu/f8MSjJNGOUu+NNPsmdcEsVlgh7EVU9wQnm4aPU0V1qGmhPHOnBVX6ar8lG0LxsOPU9PsoLF
2UEII/reh28FWP2U8q2ugHmkyqZvEANLTj3x+goyFJhMocRGWX1/Jut895DWU7Km/e3e646RcV5L
wo1+ccFTLbHC6LrxEXg1M1JpleiSHUhiAsZCBa7JtOdauymwlDGvKn2Ddl0Q8aJp2u+VEYBCVKzI
9GtAUAClz4wIEArfAfO+ufMbcRJPMu+cfoKwUrcAXg7G2HBXwPzGdkp+99WBcbPbnv1to0GXVn/E
xFqjEW1uQToARkUBgoreuXrhjudkMrXSp640kHBR5qpw4lx8gw1hiIZ8I1Mv0aC2dekJzuqtB8ZZ
2/2kJCD/N0dpzyDseirh/XzLhShVIwtryrDG3+FcxVz/t0RiV3yYSYiomCQicqe5OtzJAeklMxT+
/u0dleckcKC9GUe5lpi8mvx5v11eE2aGKCaqDSmV3DvlY0NvlixFgFr7PhM00wdwl17uZNCH9Ens
6G86qZhM4H95TfLdStqe6q2JpRO9J2KcpkjQkUwu9SOktlXUHpEqIVJa6fDBThcAJ6xxCsbWCoFV
T4Rplo2B3dDS+YGOeATyzwA5ONgqkVd2iIc/9WwS46Iz6tFH2hd3z7jLgNzZJkoFq+25wO+gzTsE
+4evsq8WMlYqOu2o4gQPqU/trCk3C/qO/G6v6TZoUtIpYFlAdnzLz3/8ohEyNwb0nByYLLbs2R03
CaqjUvIZaP+UeJPFIyJuHEiRmaPg5dae4kpfnouQQQ5HW0RkVQQ7V7VhzAg00XNpdTRPHKK5DgVu
FInLRG5/Gy1SqcSu6ExsivOahXX5qzVaWJI4jXkShFGh4gQlhWLMe4y28W/Fuh1XJdXGDecm/Blz
mpgWFPNlQl0txLuCScF1S1jpFfdnuCEfGeoSSZptd7MepjQPMvMzE2VUfYn9eTt2xSJLsj8IzNVe
RHnoDhW83ZLDbg1izkl2xfOS+kTTw2oGAPVxGcLjA8Ad/oyw26YiU+vgfJ+ZNbxagKYp2oqw5mBx
mkrVuERhI2zF3Xw1iMWbazSDGFHs80TROgwMg7kRVyc4OKSIBnBRsMf9D4TFDuJsRkvkTFM8ODf3
cPYsmhOimzRur2wYz0dzKuyUap+g54BB/mevvYwPzcGL9enI67LxHqLi627+Qf9xHvKlIvzGM9MY
zTNLkUEZdsdBOSvdB+8+Nws1UPgmhH3CS9duGCf5W7YHlPwEO44NTvieD3m95TzqZsrytU41vfuA
tAlKMp9ozRWq1ofaPmKgCET9/0HsXVCO08HXoje2Q2zz8vsBEszROCc8qgPMqOMNu3XWMpYuseHg
1FZq15qBxvOS2t9s6qzT7qj9x/C7pMCeT1T+JVh5zYzcy3DRsGRRaLhwMcXDW78r/SosYdLnU0BH
QyAdf3OmvVKodIXI5Ksf2KaY8Tm03lMc8E4rgFtWjehWgQAoyHU+XhLAJlo6NWvlNWODucgILn9/
jm6eHzCJEjro57pSkGyfyq7FbbDDrc6nMj1oHQcHRz7Xlr0HaubLH2BEYyFc5fIjyJYyYfdrUJLO
6gAn0pi8nsM+v5JXAirL3iP/UuJKd0Er0RZZ1P1HQp03hfx+O5ZUlsYKccL2GrUxiam20CCceJ3j
fBgg1pd12R7esveCBoy/QwASJNbM59pUi5jwVWwSgMNj6x4WS+wNbFZxcbbxOsng0ERQjr6hx0kt
NkqDk224q9x2Y0GRrm7ymOe8ubIFwFET6mf6EJJ/YjkFneGxDls7qUYOGM1ZhiO5h1Ef+SlhXAhX
v4JdBJuw5rZae5SWjlsGE2+XpfRWcR3nWom2Vs7Enjwhtvj3a+CjKUOBeA35S/PDVtnPcdvN9HCS
2qQbqMpEUkR6D0wfVJaOQ/zJBru4rNIpHS3CPhfh7XN6QRIIrskdLWmou2+B3TcM1kM8ZAn8uuKp
/BQeKL+zbjmcMaPbBTPQHkJ9sj6sKYyyrAkBfOHYB2TPmUDl0TDNOz8GjjYwu8epV1Px+mer+51E
+/OhraEHiAAc61I6823P6g7NZNhag918tN0ektdHIBflgz3g8lDY7OkuJwpJcNHEEpe+cgl5tTg8
yImDZuce2g2YYd02xYlLPuy3cV/tXHLm52cCMmAlp4oS5JLdmltxPetteXogcgze35E/Bt3Uu5Dd
jKXftP5Ns9e6UXZAOu15SOI8UM+87f92jiMF5ngoZJHTVpfXpF4Ju6lvZgpT8QDe5VPfjvMOzddn
hnUQa6bZKi8qLhl6z8tsxVOWeAe86QSDLkLKRtL5VGLMPeIAdNQpUNn/7cN299lgKXmA3u1UkmWN
/TXxEuq+wGQsWXvf0DZqd6/4f/XZwbOfk8NZcjjU7RLMMdnsb75raNCmdHOAfHomhIPxDHDh8NzY
yFCAJx4wcsU+uEsKJf2Lf9q3sXl2jTd5R6sazKnUPTpc1/1dDF95ukEIDB9NsthdVBWDz5ucG3o3
WAXwWpK3kvDc7ZoazZsVcLxhSQ/i42aLkFgkds37i0d6mpu+SkDc3Wff6Mztzj2nP67al/ZcRDbk
UkwvdZ6NmBWSlX7Yhl9tzNNPuYBBalHehqKhLRUXStGjgj4anFKEewexA0o2FlRpcjH4nWLYcn+0
H1AG3hBGlmwl12Uttjkc25wvz8gOQepnkMN6YQZFwhTpFg2h0NuGlotaZa7JiCHe6fZRHy3Cwxxe
peECFdWNK3y22fl4JYuWmNBkkftAZMY1izONOt2f1HubtPG7zRTRq3pTbp/B/FaL0qaGyi7w/vn8
ZBgtJV7yGae28SJnFP82TFA4uo3Ec8nMcniQErmRHR/63DFJN/M57DprFMaiVZKAan9j3eCIg46F
l8Fjsvb7mpjeflbYDAQWjTa4oh+kNOo8CP/rpNpsAmMK5Q9z0JbsMYZGaRRxB3WkMzUoXrSix6SI
mqCxIQS4GT20y4Ja7+6NYhu4zNfFvhYo6j3RwW5s2CKZ1pHwWaDXG9KbVU09/zQeR1eyMO5LdRKY
0qZStpsFM8RY1NODNNmjXaheF93WtDwJck3WWW4c9zz7eF7fswDAjCfe0xG+az1ZOV1pFJvcJ5vh
axLQz2nrcPwAJh5y8vuV+3lxCwvU8dHiEf2d7SIOE/eBpnnHlz9P1NFpLzgFDqdUK2PaS7wRoNf+
Frvvgtoi2kzV18bRHN7FXFPzjJdosTKY/H+XMv5pJ77Umq7zlMBBT+twiDehu/uNsJI1aiI/G6hs
P3gdglgf127pAytOitrlBmPSmcIuh2y9jMDwxGd18AE7JAUyOdG2ImqzAp/Z3XihN/+Bd+fa3RO4
dLepMwdD1FHyQVZU+1kIAzoeBddq6Wb1gm7oujEzNzwgoyD8fdUHyYFc8vIaltQprktrI8iX5tXH
3Osl5WNqaPFfQaCwX1avbqEnTIr8n4tATevLMjZVqylkiVajWztrdOo8YBixSBd7FLEygpdgePII
EkHfwpcAq6SMdrZOYdRh+JY6hCuaTfb0yNrqbWcJKFXSRePDQIspbU5I4VEVjBL9DnQW0zaIB8pR
+LpOKaG7M06tRF1nO/cYffzVcdyA2C/rI1BPD8IdWxzeo+qM7+C7F53AGWMdovBfAY5zc8A2xia3
0gMR7hl+JXdP9JaiYmplRUS2jMQ+TOQB2k+fRA8k3NpMrACyKcJ8csuf9VHhY+vK3BB3IxS+yfbl
rH5g6kTU57ZZBF5nXvIGD/5unaZ6XSj2v+8km9B/JOTglRhenFho0ON63kRvuTI8ngp3xKtPHiDf
2GwH+EJzivjfg0Sj+yLYFj0jQzKGrJdEuneEsht8byZ2c0MDG+8IRFQ7+mZfuyELxFTrmlB+yZ8J
2OLSisp2VNLIAfEIgTbAAF1qobTsn+lpWtibfT+bbin1PpgRRbkIkmq/kFB0U2UodICSgmsNfw1n
nz218v9JxqoqsXkXyPwRfvDGFS0T0n541j0kyLmhZfZOFJz0IuXGccIbknbvZSp4VG76Hd4LQ6Cb
CFfs8c1PIYoVOQ4z4m2e7S6b9l5auU8J+fRDb54tK3bu7QdNKFi5Ld6NlDEFC1lXREMfF5EwciqI
MrqXymOcIBR23pcrfO+HyECGanuLifcRe4ivuPCL7JUZ5sIumY7i3Do0ZjgspLdKt8sUqTpzAq0n
OXbG8h5EiioN8eCNxK5OITDr2KCL0Xa1uJgBnVSMS5trS2qm6/ww3utwAIOk59ZSfgGoTAVmul2F
PgqC4TNdw7j16f4AcQZTdczPlaNgIT2dg2HYZ6vDX29uNz4iZ5uVetFfRBs+mWqwV42egAfWigpQ
Md3PDnb//+1BnfE1tmv3J2lD+phZgAWqy4Kn7BjPkH2M4DBI0kuPlQLXnqaSKe2vt3nmoJSiHnyq
ZW83wHsqUwUJHHP2zzKvgdlhyWpt5pevLFKWyhO2+jWmIZ/6Iy6i4yLFhUjFpeDskkJF1QBg1SI1
UEnJEgRB8AxRpEJFFFZhfxWBKAATqiOQeT4b9MMI3apVzBaLAnDD3dth2t6bZKKyvduv/f9jv5EZ
9e0Mzlajf3gGAz48xk8PwvPUMzr1boaPomoi0b7auQJ6oQdCHveJjQSpn+PZgcmVbJhr+/ou0KqI
SMloas1MxqiCSqB0eF2T9b8rZDKbYqaJfDB78e5Wlmy8u0K7uJlpCkddqT9mtocU3HKwU+AOZfsT
jVrcv+OMedV+5BkeARJOzrJofhv0kFbIRveTw3HvIcAV8yC3z4pZH6T86YE9O4/UovhY98Xaf1w/
4pxRY1qg3MHxcapGDOwwloGUpp3C8nHWDN+wvHupQbcfwBgA6sIsAqaF08perEDDn3ZvKmxMBhEo
GvMpj0/LxMuSkUxN3CL8isKxvsaRyai6jDNSewRLzNUxiJTl9+VUDmiNvigJQNkjX5USp7TIvdLw
evpsfDlh2IV0/EokEeMab4vx0EHvz/HMieQ3C46tklEBM8J50ZSoF6xwGgAdoDIBvbe1lAJDr0qM
b1bKTYpLaNgp1uAA79KAZwf5/RCXLZVQh8xnE3UoUizJSoFBIhgVX37zyh4pE2p0tZSsMz4Sm6pF
41XzE4f7DGscjE6nIkYsAwYaOTRAo8XodO5j+PnXoL8Os2dveTwaq1DOXjFUN5c9Uej9PkREfeYr
rKsVM7UAm6Ktv/qnn3wCNi23ULjdFvpEZonA9ZKm+GZkD33NapFsnYTmUbXMml077sqsRp7wdjXz
R3srUAu6FWZlF2vivke71/AbDCZkTbw2nnAQzyK6kYIEGv0LbENS8LS3Jv8hvm9xzO/ieOkMdmmp
Xf7E6dNCbIEXW/IjvlG7A1kvuNkoDzP/7kO/Chc87cz/3uAxZ3RH/1n1xKGRUHH48G9hOjkMkl/s
roWHH9yMS4UeHJRGcSjEuns+MXoeKuV5i51hvIIKPjIinJnKz9TAK9PdDSH2bSUUARNk0PhNUjTS
aQJzRcq79N00BHyej0qWcfT7MpvtlPO/+mDJqKIjKzb1pgiiZaiZ+/2X2gdBGVknX01Up4oLajPO
crv2ZRD+B+A29lQB8atZ9/RtDRn+afmVPgF22T6FBwRx+48xb5PfM4Lbqd45RveYGMlSW8FmrdjO
cXKHtNFWYbGFQY1vQi39Bc7fh0DLkRwovMZ/WDgaRFMycfp93Na3BRYKkOoK55LzoJaW0h44E3Oy
zqqysWoLm17fg9SmVdC6Ku1To8/tG1byPL4z3htIcyjtXp9K6VRn3QxVn9LOyqvr3WjZQmBXISOX
UlpJDMeBXwWaDXhrPbw3aPHiTlkujH03bek1s9JLFcV3IJ/TBDkB+ShndPpaiXweRYXlzqbWAh4r
+WztRNN6Pf12OD3hoxjF99edUEPql9jNCyAuoI0j1JpLmJ9KWUW3rGWIqxZvPPmMoFBDuIopCiIz
l3j/VBNjKUAGBL1RE/HW8w4X1JHh0GXvxWKcAViGBopOSrLopnj0FgNrGnUswO7afAXozbdqECLU
cc+aNo0niJyDWW5HcQgba4JmQptSdk/vgJeuYlEBwe+y6sSArEq5yLSqHCwATfkMPNJ7QExEUtTp
hxxxjMT0ZsNEt10jH8TCNgjbRy1K369MN86Kvq1eTt9QlzOJO00ZHmzGlleP6MMcs5oIqN3EShiY
d0cns6yT3NxuM7Ctimak7dI04CTToNjTRDfyC228mfe/FyoqUZUzHS3zcNDZeQPT5Y442MSNjlnQ
/eMZgwiM/dvXkwDpFZcN+25K/lSZchSiiHfjwvEeHexVrKGXEOFVL2slw8PfLQvkyMaSSZrptY/R
VXdnQURRyg/YCYUNkXR2jw/gAuXUBRv9SB8p6GkN5GlwGbXcdXlSrnlAhTX5jL8m58uE9dBbReK1
FhKUCWtVE1VYcXWnN852n5GAi9pQYxPlmKQNJAJyMuDlfAPzshi0Z8sqtwO75C1oOwGBIU9Qcyvn
N6Fya+nqAKQEdMt9tFS16DC5vhthsoGRS8TUrLNNvOciZ1ULAWpHdPcQMO8IyYlU6K9z5h+Piwkb
FP/2zje/TqFcFMeN60wbR99jPkVYohnHr8S3l0LUfl6KKunSyf4LYNUxr2zveTnWb7ek0n9rHKdz
ZiyO8hj4oAEysBAeukIcJOCWmLxNKZ34os+bXX+ilpeFSjETBGWt0YmxgN2mNNSj73W5PaFFcz7/
ynP6AHqtyRJuZ03hQVZKegzhaswORKqCBs2pzut90+f4JfBMD9jxMAYiC1HhFAF5Xa+yqMamut78
uIniCK2KY4L01xw35DS4qBfDYIEC0Obi7ECVgxD6mcX/i1cgCpoZOZ8j90fBuaMa8SQwIOl1dkVm
xRePrSmyDtJnxI1/IyXE2ZTy3PSreiIGnjwE3n81Qfk8goDenKABam4dSJIkDLitmp1rNMtXd2dd
ckAGeF05GsJSZ5ojlxNzqdCRlIlJ+tKMOb9i9nzf6wSPknNHaar9Xj6qGxSinRJsGpFtP6rEOFl9
bBDIaZ65P7qcmmlcBsdWqYei9C4hgoMldVOQPjmxab9l9DmhW8TofSCboZQ+qhmDSh735kVa+6/U
z5glsFY9OH0tcEfvBVCaQEYf2uAKPs52Y2idgqyDqAfjWEtzuAPX651H9CMboxrsqoga+KrT9TBp
klV9b6Ud2CK8niurIofXd1TEqbHrOIQpsBp8bT/in1TkimlB0npUIgPejXHoI5qPzx7XlDmYHw0T
PH1tzspKV2ncqkcyjePInrRAlXggbnPBL5oUCtiYQelxlBlEkD+Va9juVMMW8nyWrw+INjQ2tKcN
l+33q2W3sdClyC0yRp064DUOhJ5g4dEaEtyQuJUUMhW9AFc2iBCuJ9vqvKQgSTKgwC19o110yy3v
cUy8Zoc16JVaI3w1gVbohfe67OoreaOcvgDubK/QO8gVEXmth8lsT/Dc7kA/xznE3zSFE0o1R+xd
GKD/hcL679Io3SQGfaav9dQwBiZ/HSh1rbCuEMLeDR2h8YkeRS51kJttw4uPK9t/hBMyrQUyo9FQ
mcbNDzQ54+1zl2bF3ShCv91YFB9k5MgM+fxG/X4lTB8oNOuHhn35mWwOASledIASEoyvJi5PzP15
W8A76V5XHm5dBNaY68JB8rpDIMPN9MYIki7vqLYDcWGA99sKIxjmujWe6wMCTSO8OreDpc1FhBLt
1PLnyGUeC61/h20TuGor1vr9ZEPT/dGnmPWumxkRoplmstmWlzG6PunkQxDVB8TplEzN/QK1hVYY
ZgxXnWjlHJvT1FRdBPQA/fhApmewSNNMMQplXlEUiY7mT6aW84c2H0/jlQ29SPber2WwSgbej7oT
DhqoMlBqV+MeqPOPW0qHhZDbjcamgIGfq1p3qY4VrtjKhaJ7BwtbZeLWNyvsZWwDIMD/7Hn2hztu
vQ0F02i0X2DrEeGdkDQTKEJiCZrnVpGs6TqKGL3lsUQ+o3LOHo6YjE3InZzR2zqbbAWY6Tlb9RNV
es5w/UrmpzU/Pl3v6tqmCJU0KS6e1ihOkRitJna4qgMAEGyxNrWy6DUMruI/UjtGO/EfWyxAkCXK
yc8vQfQNjEpQ6Uj1vb5muS9SK3P7fAiB4BuZg5cX6jut+gX3HNZFXmG8p0pUQkiU3JFtE5TOLOUj
Vt6TFm77lweVpWzvmML1zhXcPup++Vrj5zjtBa1+qnMIVChdH5LrClXJ2AElSW3kUT3T+xjDdwM8
wbN85De/k6kOLOsewVrQTyVEwInv1UzISw0tjgvNirnVJszqWmQql+6k0Lnu0MzSdubU9V6MXB8a
0sqm+pnCHvovIjG7y9AhZ9MIyc3qVUx2YQiVQGiJLTz56wP41Bg6lfQzQGT3PfTAIuMfc1Jplc2m
incCh1qsK+PKmUbtTr4zmDmY97ZaXt1q7Pi26fic373m81ZexPPYyvoIyFLx3atzZgXVNidRagtg
8md+5E1enZV7FLiKkvMGy/O/b8E1mXjvyEUxqQTh6BVOGka73fbTXf3EKUjyCnpNEBZoMidtt+u/
aa56CShoU6h+0BtfGOO+9WQmWghSztEnqhLdAK4CY5USkvjp+Sbv+SmD5IYC6+v0/wQ60PzOvy6m
0zZsKIhIcdFKVMMeiBQOasICQ9jGrx1a6TA27b/hJxxsf0w2y+R43QOtg3xz40Oryi3o11Cx21wz
ar8HIloAp/mVeqFl+vU0CHHtkaqFnU8R6DD5WgKHmAqTrlg422s0zwczDFoOJHDrePKb5NZwpDFH
/zUmsVkhguKUZ8xHcOINBZmBKc4fTo5z/vWZePFYPA86ZqtAzLKU09LWxe1COu8uK5sePUKgkwwI
NEqFfNu8Zy99I8IG4yqfpfzQNWUugMeMAtmO6vtSRB965//VjQ/eBJ2zcGaoqh9mlLmcjqMHb9Qp
9AiV9kLxpP4svHNjckmw3ZL0wOCj44QALHDD4SJ7ERvFSn0a/taoWp2QNGURVEuK9wSPhISZckpF
68iderUo3CshWGnRLeSsrviT9YQL/Q+kioas5RkUBE7XToDZr1qm1bGiUpUqNx8WT2kNKdP9CjYL
UiauYpXynBCORlzJmNPhrGOA3M+HcBY6pTN97QWwQPZPenzhM6z55/I9VYda/WBASa9qx4RbzW96
BJGknvud/bGoMcrRZ1dqO/ti48VB3AJFtte0AeJxxdO6YhuuHkHBULh8C4c/gyDOdxR1TthduHIk
syXGhbll7r1iIArd9h0p85zgWR0cCmENKQFm8m4QSHS8sMKnbVZ0Rqf/wO6R1rhB6fI62NEu9+K+
gw+muquCbfnEfxqEWeRcvCTrxOBReeFrjjMMYeRlsmrVM7AExsBVhrYNAxq+kxqL6xMVsMBzk4sC
O/L7QbFpvY1Py0DmyMhnGk1upJrKiRXkt0d6NTITCNsxM/R0rpTt4vQ292dzJSpCdQOV1lVKR3qC
Izb170jr0arjiHQoI9RvgJB4mPPnc+Hj//u80FkyVpBKOdye3FE6uO7uQFEsSwqmXh4Aq+ZrZkJr
fA43CTCxsAuYb53W9dAyzbz5r5s9t2e8HQCGoNxrt7MRCi8y1re93TusYGx3E9KJBKijrYx7NFRt
rnQtPUKtdJ0ycTDUX4asVkMbMbECm2Ogyx430SW1JDoqpYYoTR1866Pg66wprlgKJSw3sDwozxHA
Z+wxwEbVn37SYSkmZuC2ZXpFiK9vIM2uudt0WrBgS/M3lgZ0N3Qu5eH9JeORx9ZjqBslCRMkur4I
2SrjtaRKgP5YoTIw+cRmVCIzTioYojX3f50JCqsqQCZpioHbwtNtOI4UdNttXgXndk7Fcnwvozs9
JhhROsOGma6+avgsQAUgmqvmPTkVJn0JgnKC7u+2xkh0RBwGsp4YMFbp1g9KRWQVYd2q1/hFMLdg
lqMXrWWrLPUsKgo8d62raJPT+IuM8BYOw3LItdlBzwuA9yosEKjzT/b1AhbY5pEmIa0d/X7+7Eax
vEpm7oectf1gkK+6ZDfbrIWBOyemQwu4jzZcwUCwE5olRy4n+dNl6YUqjeZ/NXBWRcvRLWqw6QEV
coecHnK+iYlkqd/VA/ds7GgFU0g4KktPcxUylsodMsBWdV6uR34bP3wWaoDp8kQUBHZoHU1au+Fo
BU7t13+IzY3TRa/llNH1V2FROkD0CfUosuuhyMLakLyATDzGoQx671dU4Rj7r8t+ZLFNVCPn1Y0w
NOCFr9FK2GQ1syKRZH9AVSEEarSDk7ylycItDiwz6XUc+KWZN2jzKui6q8eWerjvPgcyWvnmeDEQ
2FLjrUaVoS3u7JnYdEzFUECLaUUm/wMux9mtGU/haeQ5Z+BCLGfQ6c0gA1QVwYFDLhFgvsU6RGjU
LQqtPQbc8kRSllRJCIl09OdFdD1JGLmLycTCXUQXF3GgBz80oPfQu7gHigz4t/b0RWXFDclMMbaE
z09VdcDmKqsDWlIvY+ZKLvKVE+YRyGr5hyNHb042EOg5LJfOpF1qCZYfsvDgJ9SLi30JgRpfFlVZ
XOiS7pbARMytIHNPFiyjYKfzHefq+rCEYmZCDkkexFfahsh6JfYhdBDS/zrfJAg97QSM+4JDwIaj
hb6g8vbQUvVEkbwmrI+9Nnaqj5TtT8HK/9FvZmc5a/aIkRnsNbrqC2enwlIzc2yahXInZnwWJfyN
1Rf5P0GDVARfRgQQGDUdU5/ViWiYhNdNG4nTITPFOrYGICccy9d04kyvzk91Ug0/5buOuCOeZqhU
ujm4fHHnZS7xjaK6b1QJ70hMIA1HEiVldsjyosLwcrHdPJHvpDQZJeKfN6lho3eAdp84MtrGS8Gx
8wv4CeGkMookgOadfPn94lwXBijKQjMn9i4p8V7K9didB6O9zJLmPxsyu1rmnN0CuXen/3SAmK88
MQNoOUC5fgZGEGhw8NbWwzRPw4HIslVpzlqgpy7jAWGnaIg4DNkrG7LlWWROo/uFam5LBtUoX57V
B48llquCHq4/2Y5pJNrjL0flxdU6EwS2s25zmaFJFiZx6oQi9Br4eCptqkee62/esLh176lkZ3S9
fqzFFN0H8SZgQVAKnO7Ut7qZsRNji0YZXJtLUPQeV7S/f98rJV6AaZIwWGvVUjYamWYTP/m+7dSr
EdWD+INtflV9F9hjaXmQX4J9JvYIMIYT/1CRIHXVjSxmFiLdMgG7pxlbpb9LGL8LHymbEoMVV37t
1+SDBo4T1abWtDGYbZ7af/g8RatXdowMR0gGkIvRgYOU807gpKsigi+X1WTnSBqPFSLdReuFYEqH
bNicFe+bAZoBoXum6Nzxdbtwg1zKOo4/wXdOY+xZpLGQYq+aKT9mJFh4QJ9P60vnwL98isQfaw6k
+ViH0ZJINzkW1JRtJHMoz5bGoHYi6N7mzMMOIeT2mJtZ5rVx11uUwns+AUrhUWTn1nRN7dbgR6o8
ulDuSW7eUqtvGQo5UkbmAemQQn0sOVCsKAykV4tDkAxpDSVgnSnFOA36c20/dU9MX4REX24iDVN0
wL9DrBfvAYphOpckWSzQh0LTrC5EJefe3IbXorRlyRa7bIM2J6Uefz7S0mNh5usQjG4Eu3IDPT3j
IoHTkC1YFFfBx9xoJ+LMg8zzMnFq7+KL4A+V6S1cjH/hCGkbFIWalvlS9gZhGoCotSEbW6R8bIz2
iVWGExiDWv/mv5JETzZkMJNB015T8cFD95YXP7BPINAxuKDCxynCzDCg21khPh4pC1m35jBzoINN
eFE2gI8uI0S7la2E34QBbFwpsAFpdqiLY+XXRZvOUgvha15UOVlT5QSgK2S0k0Kpp4sM+G+VO4Ga
7aI/83luLT5zarIC2ZYNsQTd710XQINatxq/a5TvrcvopD3qAjea1sAVnjEeVQYY6NbYhkSaVMnH
mnUSapPm1vVbe3Ifx2LaRpHB9vGUDctgEWUmTh++pLbBOHFrQw2guDNBdrCtIuqctfX19xfn/Dv6
QAGyPDW+b2crARamfH0j1JWFxNwD57SmFy9A2Qx4QAtllLsfuw2rRYFnyF1HN0Wbrv4qiSxLyqrg
vbLcYrZv8EFe0EnBe3j7MzShJb76MnOdJ3O1UYF1dEWQObTiw/T2bCR67ihubkws6SdXjv9RcxAt
llPCrcCIQRi2lGAH3Eye070EiUepQcs5D70qdTXFnMtOeYRFpZkMR5VBqLvfaMIdX9Zfb9EdAVGH
loyYOnRXITTZ2aRUolMjqVvb3iue/J7YsI5KlZXOg2ro+J8IwaopxHio0y8uZ+FGDa9QtVVTaqlS
/ihpD78WqGxaXbkPfPjDS9ANjxdJBxXah+ddMq1yyk4JjqGkqZTBGIWBMS+Q6FyB2Pm8saRpugVa
sxIUcOQv2Y9h1ny0T7sroFwGtbD9/Dz/8txcJfxSocy8f52QZfeRGrQKgyTXNNh9H4Yup7Xnd4u3
V/qXb+jup5FyauwG2UvJYGnWIU++/XIO1TB0SmMyXSp/oXvmdVnMSitqkMhcCZcsT1OFTUMPwlan
sQ5IxWRqJy8422ltT8doU4Jj8AMtEszc5MhYQAjGpWIEu6MtVkiMfiBZ36vS3yNFdXsqsxj9rIRU
2YOwGAIVVZ/wcUc4ngZhZzl6CTjFGPuyXvjPSdnvFUFnnbrQksTXX6OgSRMu/WZs8clWXxgyWJ0i
Zz0yercYXOEneMbEizZ+sZul2n5jMdADFnQdLAInOD6cbvAjjEIlI1M5knmcoK3TWw92LXpy2rBt
378KNZtcHJK5KnJHLLbvQqZJoHzyLBPsmmNcUZHbUae3LKI/h944LmpeBT1L26yAfqIOBMpUbAa7
z2fo1InBkomqSp9y2qd+ZU/VhPiQtVgTDbDtdB4fb8imwE2RiPA5KAzgBOJEND9Opdb/9fGcOpaa
oeyy9BiCnxPyYGdBKsW4UHCpmSvX88T2C33ctw6CMpO6VAhz8NCahx0AOF2IlSs9fo+YeJjbqSTY
HRSFaNf9oPzMABU+rLHPMBrrKGX3rTVy6d5e8emTUc2EvthA6DKJA8rSGPRnjW5QtWbGwbE0VyfL
P6tZD4g9RJS3cagReUN/RNXmMrcK8yM9uW/TcY/VHpX6ZUaNqh4qEA+jL5H+V7+FEGwnij0GArvu
JDfa4LBbWpBNUiu+8CiFdzpqctyszuGUhGfQ8KRbliQKICFvFSvhJ4pwjt1zL+ddFxA0aI5P7CT3
hm5qE8WLNd8nnVerSHMZMcC9k09ACPYrCZG65eS0MwRUo/6IMANARvqk8UMvyLbrob1jwetid44R
NjTcAhMatZMBrntukLIJZ7jMdYo8Nags5dS0usCUUljbM4qMzsiyG/rXYHplnera3G0bII4xjaT0
DWbh2NId84WDZia9zsRc3r/7bqr2XyAynzLUZOCL6xj2EoD1oZaTaARQnAZNrqvU6UZYtZ5Nilea
TRMEVBBKEkWL2rTob3w6FWup8NcfN6NWCFrWOZQCNg9ia3Gv4RNucjRtWQaiZ9ma6SdGHnlD7Xoj
VVsZjnHk1AevnTu6heOk0W4BCUBIFEOC8OTVQwjTfxLk1Zx9HkQe5MRqL7V10Rgga4rQyIIfrP02
GVa4Xqj8smawzXT2oCbnye56ehNWASvGLjzWPaxhRYda1/lzOk1jXuNgyA0bX/U7WU83pvKFeEwo
GcDHELK1fRkIgztCBrPxB2o0SR/crrCZjiaTkr/1RbI7L2M8NLN2J6Hk15zThPK4t+s7W6bBWFev
Aa4geNqSg105lzeWdONtrxdfMz7YUyjNNiXl61R1ZU2OtAlRWApnE3EEQX4agS5DqCFg59aSTRtl
XdDbjl6d4q7aXjL7/IwBr4CDA/lY7FJLe0N6fdQzUfho+eATMSqx08JFs0yM/8iroAwxuBFTJvuM
SOdVnadVJZzb0ibPFAK2BadY7AQ6kPCF/Wgup9GGDvkfHriJGto5Im7bGYlYD0ZsPWxtvO/A8LfD
dmatNEYrH8O7plJ6gCMZ1MQo9MbpCUIDvghv+G5TFwz80ctNWJVTTeaFl1ZVR8mME2QAvmyeHTOM
88iDk1YijEqwyTPKnfjyisQ64RyWT6Nro0MbeyWWmaPedYRTcstwErRJ0ECtdiLrrw0wxz4OlSdT
sYz1fyEmkBi8TreWEUFH6iuRF3FbnemVHlTvVvQNQfDLQOQgKe4YmWeCon+KVhZfSEQi2zDbsE6f
xAcUXFrjghBAzRddLSg1mDrVuGXgoBd1bfQW/WEA04dgMr6XRUrIm03EL7m1maA/oxc4HmAVSLH8
RdGAbuhmP8M64N8MJZSyw2L/XG45MetSpzt/SAYk/Y0uxoq5vaAI7cdNh+bm3vDwyF2+DT3mB3pf
SE/1WCoIq2TxQd+xTGfLqHNALqy02QDLVN5mOq7TcD+cGe+pvPXCsYp+CAPxe2CHYSXpV7bvW+XY
qypbPETCIAhFkdGxkL71cfYf//VwCXjyF+DMa0PASaMO86L/J+0NArbMYV5N42A0mgyTExP6KQnc
odvsQR9ZLMimF3q8EMCqI06/QBnXYgOxERXHz53OxoUueYK2due9LNjLblw3TrsAGQtWTjWQRlBd
XyvfrQzjkwpKGE7l29FF4oC/B9cj6i/iASH/FVk4ccQrmmGU9K8Wcfp7bsOrn8EHpm20F7c60uon
lcfstQuETwUnW1YQ8gRU5zPjBkk55f5pcKb/uhaFQYcAlN/hsFUFpCK2yzaL3y8IuZk7nZSquPB+
UEeaWIxJjf/sDE8fMe+8+qATKzIlA1qj4JTzWWOLhT/NrI6q42rG502qo1luCvdoYaB16AyMpqxb
eiH4fng86bGg/6KYJS/OQOwn9Jd61ZBT9WOZR8Ilr5kztHw83k/AMb6zUyMemRiudhMmZxgct4IZ
PbJG3ozYpK93Zu5eGVUR55POvTH89rgvtWJS9vt5i3KqRavleXXL/c8wYn/jLPQ2iNFeSODLX0hU
VahC5xEDxDLgcUCK3KFUFXjukEm5d/mTN3Ls3mhuSAdlEq4qzIRnwLl7fRuSaEs7nMrF3PsWmgQy
wMPoXJcossQ/eAOKNyIYSphwgj9EU/ut5eNlmpH1WhtpMDPzfmHrX3xYfh26k0AOxVYqSitgSQG6
QNHohtzw96cXUR3JTXeNfsf5DfLObgpHmfauuCf0IOBrjUcr2mfOzIlvaSzMj+Qpdpdd//ZlhRji
VAOQ+ry9YG941To81P/8GX9/bVaw6mdgcO45QTzaFGFzcABLA8w34yJBcbroieZRMCk3YTleZWsq
cWT8+/n/XZsubhm4NdQ93N89J1s44JZiJre+ublKeQsgc1r4nA7Q0ge/g9F62fpmkuFqcU58Hdhw
Ig0BJqCadmGFoYh9Ft8udP5EZqg19vzxBl8lqR0el1dX+u7T6KC3wkMcY34+tbL8Jn7Z8pJWvOIV
FZ5cTI6sdtIOtU1Rcj4Nvv29EmXHJLZBxS7KiU0FGk2gNHwivdHov8CeSK4APEmWSm0koy0t2NjT
unDS3T0fEKqJlI5EuyR5KR5UhxQTix5ZUnblKc7CuWf6Q++AF7580ihY7PMDkWPRHDuO9YMFPGd2
mxIy5sN3hN8+vfSzxZSHcC0hOCVJb96ZlWPBDgcTp+YBmqkKnjgoyI0AomUqJ6eWdW3lLol1S1SW
YMVW55/Am97vnEjsMvFQScTNSVUb7EUwQVBPys1hC0N/i6ySluA0SXbyMIEysjZkgL+pbCH53XeB
Xqaq3ZIIt+td4/U+i+6MUaIWqNR7E9fYJPVDMZ4dphIcyXjwHaQxaHjo46MAMOyuvH2SfnSfNAkX
D6xrAHel7b1o0mDl0RKNa8Ubhk5NdgjGMEUonPEsVTF8AMwkbJvtX2m3PDeNMzYwp3Z4EFRoF8nF
fBG1Kh5aSFMAk2lllmOV7H3Wb0yCYVAwiPeB+LGoOBrDW0DXs4XzZAq8tBct+XpD82qCuq2ffHvz
nitI5cWR/vY+dJhNfeVgXD0PjDiimblNnvy7O2tAb7p0xAGbgCMQJNuS24dO2vCMEZCU4UAdIufF
L4qacdsRSzHKLpKqvF9KZvDN6w8aXnFGto7AURrVqL/12ghKwexRIECGK4xrYYlU5+SRmSWAPZ3+
ihjGwvTT3F3ithNO+lTdsOPwqmt62YAKyPLGJH7hnzA9Ln9B3ZqVMuOBBurbAE23D0lKLeZkzlGX
111CPOQBh2LzXT1EJUnrUat11tS+XwRkKjdxSIkYv3Gih/PheYA4VHLJng17wF3EeH2VDgavGehq
ObNlzgen9Nz6RizoXT0JmD0AqVQZv8Kv49xseahMBwFiD/TEIMmW0HqLdn+exRlwEftzWZob7huv
fjsBEvDqCvsqmV5yG367HUHg74eyparmY9g0816mY6/3Or7wM5jLKb4QjPGADmInQzzJ4Z2FdBAC
HPyWg7Gi/jkWplYMnX2b77ydPCck1cxjXxovoDaCACWbO2j+CN/IHJIY1/j/BhHh+/TJh5Wjfn6n
q61Ndg+PFPinKX/233PV8Q8yQlyb3RcKrSCYajT86mEBMabvrSzZHCuP6c2pHpahiQa/BwRRrav9
Ljis8qe9XfLak6Ocs7n9Ie/bb/qpG3w7/ozUn5D3DxItGflFtS7ye7L/hNMOD56ne3ciH3jxHtuo
zoz8kHzgF81bBRDlOSEbF/+yEdcSFVJgdjkw9X8ZouOtQa0KFDJtTnDA4juZtLd3EF8N2NYMOR61
jNuNFmJnaU5EMvUC6/saAM6Q+tOnE8FBjGzck0hrtTTp4cupAbWG+ttFVhq1r3wL5MzHxwDqw+4y
0uR9egej7pmw83zsOuPMD/h5XveP3KTQVqVH0iAQFBm5xDlkugwqayh2tGb0Sl/+v0FVjf7mxkMh
lw0VKIk5w+LjCGgygUZhFGb5iLbZt6z+4Kea+6tbNj+GR6yMnRSGS3cSAvXI/1TYL+z+ZpdKReF+
q2kToGqZZoio68Sj11fN4kh1xmrQgcDiItoFIkjLM0OYlpNolU77EufXr/+fqhTIJaZDVQRzdqf9
sBPPKOZX7m8YurGBRGp5tmFQ2Ekon2fPd1/VXC5xJOf+r/mM5+g4R7N5IBWnkxLmcSKa2kwVhsuW
0WYNWqW53e4BQ23YcAgtLSoJk64mA0hYH4L5mJjsRuPqzcPgwDS0JLapvKCfv9kZtuiXQJq7yOPX
0JADo9xNVq2f4mhaMeYBPQ+ejMz48IdvwPVEjbnW4nqGwj4+dLTn5RrxUKhe6tLhkIxRtvuoY2sL
gz4IfCVg3BFumRDDGK7fn+5sS63prOeAOwMhD+Q8e2zssPhge5Yh5ULMLE8gWKnFxO4mZodnuGnt
zExxCsa+IDwY9RKgPccvDYHM8RPAmsUdAGCZJh8j3dlWZPcyb6Imo9Yq4CsnA6LIZOgiYif/32hO
+E5QoDjdjhk8wa4SNnrkN1AwOSIDK8211hdf8OHs7zZwVO9LFMSc9fAZdT2niDa61GuONzZSXKPb
1xXKNzMT/I9af4CBoZF5dNQbzXA8v/5zf3W3mDKG7GR4BRA4/6GV5TLQs+jGM/wIGn85vxkFZmw6
e6Ho/FwBPoBs6ej5MHS2gaXGvE0hIk7EvmdyxEkuOXlVJuizZtwFrftJCd2szGdXz4Ljgqd7I0Yc
Mq9h+D56h2mV8xO8NQpvCaHvqsaZkIje/XDhW+HaROHGR3R2qsdsy9TA9M2a9nMN3Kmh+iIUGxiq
AB00GU57Puh5cUcKdWsP9TPLW70TSzkMalD4GkqWN34ltkrPehTPulj8+pKqSbUCp9+wS3ielDW4
oHo5ncwSNVNcyF6lW5oUy763fGGdP1MozzmeaOLLmy/LaLSnvR+9E5y3cVB0kxa0mdwwx2hJNqcq
T5oB8fS54x91q6Xyu3hjMBe+ZVeB3bYiyYvtk4KG3iH4fiiLgpU7jX/hlVwqxDsfaNiGAYDKOD9g
vhHAZmOhc8yTLHrTmcyPJRQqCq+3qCqw0mXwnEkxVXEK3AfL8Adh0v65YSUjo9bvmSKlYBdcdbwx
PM3Ri1GlW6/CYW9ZyRvWRqnnFj5LKmr+qp9zkpWQOk74OC/MW+x/nfGIoK7vWiBJ5gqzihXpf1d1
dhGTeXJaVY6sSz3gIHzGWX5U+SlAc512mWNita9QWNUSli04F8emOzwN0+WYW83FEKt9J8naxSAM
NTIQcyBg/6+FLGDG1cFwGYFWzL827W75wdItP7rH+GCS6zeoKsg9E7YFOVk9puRGl247vOtC+wQV
iaWhtCan1NZzhdwG6AzeGhpjV/51ldsBZaKr1sq2YtyHW1kXq7/N5tYatfBRDzeHex0VP+BnJvBC
2BSM+skPyOlqyHZRQ5MfhGVAZw38ko27GmLTchfDCg/C/CC6bbe2Nx/c77mlm54XY4ycs2dE2bTE
gQ3hpS8FliEt0/4teggwcbyAhUFsjr/m/r1nrVskj+nawcQKgsqYQ7mSqPoLFeQPmAesoH5/5VBT
gG6K/nREN90oy9mvJ7QVhoiZijmoCCHP2IiG4ddqFWVj94w5akUU87cBqu6tMEjREpX+TkuHhGGf
7aPk0MrqOdxDSwQHjhOOz5aynaiFgZNrs74jFlFmdwIZ1grlq8ORz1iFQ5YiF+TwxAJ2wb7vYYBb
8mfpmtLCN0P9AfKksvDaC4Gkwh0XtkqA7eZaX7dzirtTxpGJ7QPpTeDFQxEZdgx/op/nLczr3TsN
bhvexMJ5usd8yRAab8ZcD/I4VkDZKrgDSRYM5n2/hO0ZED1Iri/8ClXRAJohg+0YvHJ2xkH3oxrm
GbZ0XUZOndrsbIJX9yo6Pu0v/s3AaNaaNdX27XE9eulUAoGSCDSwmRbcsZ1x92FvCPIa0+7far9n
GZkAu5r/dwW1Q//343ROKxqu2yYZC9WU3cRCTPqNrcPDDdAM6C5DO3VK0y1Y0sD7MpQC2csIClyE
4QsY8Y9pr2Cg/uSy7kbVJgSKf/Vw4fC7WiLhcphyQV0UcqjFmAEyhXec2sZnCYtGkn74znyztvgN
PCZ8WeykV+JFqia/m98AFe8Vic2D/lRB7+cav0EZta+xeF5P9U6/FmzQJpEKxwQLsypWtlT/8X8t
O+tYf1DCyS0rkhQyej9qz2WMtAqxOWid9Jijr7517bRB8sJHdG2Ajj0th40CJ79rRbT8E9rVUXai
+flhw/WQmjlIxJ71xTMAK/KiEiiwd+HRxeUgC941tK7EpO7P02sham8JflejsIhtsZIhnunJh1+I
N5/JqN20/urCPQo5HFo5eH0OL1bOfyRQqWfSFGpTj2xRPXqXjjteUhJUQN9/9Jj7vz+iJSiRdkNU
bxWtXL2F2F/yBvQVkyppjuHPcgkR+CJIjIbvCBOP/3DfduRyTwTiBTyZA/hy8364JZub7qiIitHy
j6+bgW7majOqKj+Gmq08j7WmxP2MNRto1n4TCtlhzV0GjONSer3SmkBEsznGYz8ED60x7fcUksez
kVhfXm9xAuhcu48IqvH+6Tv5BSRxnzy1itLT1hL8g1YyX3tgcWKX8A37p/QaO5KCIWDSh50xv62S
hNqYQfeGzRxEu3F783P1UwMb8iyskvpOHczlkcVAtgoANOuLsq91maWd5I2LppFa06KdFF+Q1QTL
lGX1fH88QnJE0Lo9kzUIz/gYDx+h2nBJ81nVg6VQqA80Oy95T0yIzevr8RELWkP5qEp4zuJ03AIq
3ts7V4jXtAT0a2Nr5e1YBFuc4s6GeUuHXbeMLTgcS/aA/AxVgwuAiStttkbCAXcjHfDxFFr5dzXa
p2m1FbqD5WIWTvqw0LU/s4kf6SMjBestqFbvYVHNZGIJT6iN/ci7p1QJobZPGtgNIgyakw133g7Q
yWG9W/qWM8QapCSldrfWxtIpZZFvt0d0WzlUoK/z4LnKQDUro7RMH1MzLmlAV5Qvx8ijDhTsdBBS
+fewA70zAZTNdPhAfZEIKzOakoBGXcWmMr9eMJAqlZuTJnOjQ6mD8P4muY2vf5QqpCkdHKlLWQhU
Hsgwq5w3iAhXAhTc/A8K2dNrNFZ+LPujOcJ7lsxaCGnhbiBdSrZq9JvsLQeQwPXbk/2Pk2X2Cm7i
QCMJlaRlX/i4CBE6X9NN778rNoiRtmqmIF5TqvXBE9OpQ1qbR8Iw+g6DGbCnZPhBHe4SqGjBdhhc
f8/wq2nP3UXTDx/ZMqG7Z0Lz/jyx2AgOk2600MEYpmW5qvEIuMJAaHz1JPYqP3p/rQQI075t6ERq
w+KLUmtpgjyhXxMfP07URMlSe9jZTh3hzXToNoBBO+szBpmU+g4HpfwrlC5UmADVOQgTOnqWXmwv
fOMi3CAcjB5AYBkTnOO5hHsdLtPLKhsRtJtnWa5L2+1CJMmSy+9Pf02WhgSBLBtGkiJEEIuERBh1
0eZ5LiSJK21NJyDoyzvQcuy4qpHCDcRa8YGHHAU7iiCrwlOaPdg4lp5JukFe6KqDTTx+bdMpzip2
jjFUvGYZbFn19x08cpt5lB8Qpt97HHlfXw2dmIVvZF7sePe71HIPyU1wusos2mYkcFjioiQoitde
BvDZr5sY7sb3aOyTtd8YtV7U0CV44TERkalutHyxTKyWEwulLixK7OcJOmZ0TSLEPzILV1raZaqF
CxuPgOWIXwplzVqXaq5MRzlmYNYK5hPOgtXkdSmlOCafNd/hPi1yqQBT3wrc7CFTa5MYKOzL7QTX
juVaG3AOMuC5hDRJ5XPhKbCTFA5YFyZOhiWkD35w5df7tOLet44mAgnJpzkz+/+fm/vAbNQJckod
QnzT5xl3S+j3HJiVEH6ZB1VhRzTyFuwGkLt2hVXQBUNVgLFMlkzEBVkfwcaUONcQVM5uiS07+DxM
DBhzG69uFc25fXBZCi79K369m5HoYQSEpYA634qbUPWLpHq9t2GLhy+UxwylwQ9y/wOgmp+7MRuj
p4KYl5rxeV36hdu+7y/r9EyMBRgYnKQxV3AK88BwTPxYXh4Z1jpqfqQCXByajkm4lc76ZvZmnJsD
+c4knDvFnXayjk0Ve+eqhEa4SV85NvK6pSo0FnGaTSGVxSSTbD50R9at+A6DtiTD0zZGRtEvq5wz
DVVIjjprKFzEK7ei+7DA1uD9MWP0pmJ7wzolQL9h1dGJzxwfp8fUZI+bQVtH7BBdGkUR9+xBrua0
k6S2ylcehRXPze//ak1aGzCUkVjtfQOrjv+PEYBvrdi2uBF+NK2JDXCykTqMW7K3JLXB97mZ6qnR
td3vbVZzLari6Yf3RtydvWPjkw3E67wbBbDYrS9i7204vKNCOmzFrwDig+oUUua5JastIVxQli7Q
HV8ZnMGIDbcj7dpGk90PSvL/UMK+Tqcz9wC6EAZ8qJClvweKCLpiexW0ILLfZCxYNOHBZzP9qwYS
E55fE0JRgIOAajBd19b1pRTxqhQ2rOE0xRbMhbGq4Se5NL11kwpsZLgBCRpSEH+ruAzB7wqjlsaG
+MK/tQWYqotnP4Qqt7YK304Db2eMvEJfT5Ugi0fqW49WQKSfsCQr6Kyb6vNPNTzIFCW47WxEXPtj
gTlQ2gI26dnYTVb55VK856YylRBrI4HmzqjH9lLZYxczokrUJq7LonueXbAZ9G7kSyKdJWaCOVT8
2e2DG1885F/v0+TzvUaiJ/zMZ17BAgAHR6Vnr1DL4XEO1SOF2tk1BFnpVs64ujw7rNIZ0GDtdsHZ
TC9NhV/pOKEg5rH4dpuW/nWW34i6Xf/vcIPFLnvjdrvR47soaJd1n+cttXU9sLFCfLRwvBT6KSMz
J5vMhGQ6KJm/6qtqk3xmKhn7Jwv8Xw23WbqwdT6O8nEITUtw3xq27b2jVsDP+7e6iMDSWY1CqRa3
0HJcFsPGxdILJY8SmPvynMWeSBQ6tT4MyYbNTAxExPxeCuZKp3d5En2NtkGFoEStMQDgeLETq3Jk
T35+GW8dYJLHb5Q38pNcvqrnf7nSxTFKCNhfgJSTpmhFG1IeOdcZbP29jR6JEdLI99DyMfKsPegH
AE6WiiNu5b6T3kWMK1oxBRy1rRxIGYQL5vy9LGdIsUikmlYKFit4aBs3h5GooIxHa1bwzEnYbU4o
oFrVkp2fEpW1N5utW+Pno7bjxqjuByL7Tl6yTmbiu3uvgeRtNxCVhEYZYWp8Bz0O8/Eeham8+ec7
PzCHx5nwpq1822q+ZPl2EcpUU5N+ucuSOK9c7Qtoci+IjURlg/d5AGWpfESveab+MywLp+1dfi7H
8rffkh+y4olg34EQ1tv1fHPsxyIXy37MfQ2qo1xTLc+8BdFwBbEZdeFmN2b6ox15OWzgQGSd/xqr
yH5603C7IsJC7/l5/ofz4BSfQ1DAEhL2q0USX4swq/PNHJeVaQu/RhOgHm51cLTWKzYCHHY5RDjX
TdA1igUnD3RY11JRH+gWOD5XL5wd2CdSBkooqH2w6At++wKu1/jLEUW2XqofJ7W2Qi1RszOQPTdU
0pWmOpxUHj1Sk+nz13Y0dInNy9K2guKy9HD/oOQzJKku8J6xChUzbQ2p8IL+x24oarasp6JoXWmt
0Wyhw75mOnFjO48AspuDUZC9833MVHqZrk74h6wiayt0cxcsUlDZUYRe9ycFWyAl9/2dJs2/QRxW
x5xz0LESk/D1hDQi5/LlMjFME4eblSNWfUezdWHie76S+ChJaliOPXCUGzYGncWkWPNh/2b0P5lw
xeqs6u/rXhw4i7OhoiYcpdL0Nj/kT/+iFUTZJsEb+9Y2krKtZHLnK0pZQ6A9/nteDrG/WK0DnEdU
7GtInG4ltWGRABUbWqzGPtWY/r2Zb+CC/PF+S5Y+Lo1Wkx8QIuZ+YYlKcW2tzz2UaOTy3/ege9As
yztyhP/y0LWltpcXz8jMIbOPQZHpP0BXZ6SyRmQ3QUoyNaBgmudWpfdOQCE7w83zIN2gI0Wusrgf
+mZDubqbcbxuPcwZIpmamfiAlQKzxvGg+3pdkwVYnehRzmjtaB8gMUPLXq6DVImBMOHziwWBewOw
WK3yoYdxawlywYphDViLz1nQEz6YT+5kULQUFBNSEUEWf0Y+wYbKmv8zMbWdhvtfsAPdPzzzm+8q
kfeMbds5ZoGDvaconqUUZl5iRu7m6W8QQG2SSdOMwfV5jrQqI0izFoCog0D/RpmNPsPydv0pD+GV
A+aMJCYOajntyzqEahIaqsXBo6NvxG3hTYX0XBXlgduUD3FsjblbfJ1jW+KMsXHUFirAUaYyxEb7
3Lz0y2N2n+dgq4pbSvFGi9VJjF+wGcquRBxLthXKnLeiqhtu2Yqmej+jLGZUC8FFmEvhx9rJ2c/M
BL0K6QCNGKj9hDVfM5oMNmoNrMW+WuPApjnxtnoscx3onLhYDlzXLG+6vtHcBC1T463MgUfw0vLF
QizWTg+UaECmVQfAjMrs1pOlO0jFxaqB4K1sjm1SG+2Fr6tUZKg96Ny9+T8fIBWK1MrbhvepOpVU
tyc0oO3EuCJ5scL8lK//JDKTI4ZF5KAR4S9WkejY8CM4QdekspdLXOZQqkMcPvateZecKn/Z4RT/
1eRs/dJV6z+xjrTCY+w+vqxctg640ORzCBpe+UA6SqK8qhoVqk2pCB0q4NgIXL3xzAvxJSbaTJ+Q
YbFLPTJ2O7KfpSkf2IyXaXp0BtdtrAtS0wbFLCdbT0cpk9j6AhqzP6w5SWPBV6arXgx++b3WrdaG
YGo3rV2dsvB0apeXzTGbIC61EwnAeHVdsmkcZqbOc1CZalf3UPCVo0JOZXPpkLhn3AtbvBdwonbK
pj0ZXwPEiYxopqmQ+htxwlNgY+9YCP1pS2RLZT4RBQYwTPnNYqCqg56dFQz5WiUE2UACh8Wswkj8
K6uM8eUC98YL4GjhC+g1HackB5OE23nMIPsPDRzjy9hyQBqDYOr3PE188fOxiitCm5zHDNfz8in0
K1D83QDiSVz2TC+XRkLsxwo9GeWffsRAVoulAxNByrrRjkQWT4fKG+8vQk51Q77H+pwd5n2vTDgi
OXnwOMkgBRvJvSpcGPXtv378KIpqQPYkV/HyOUrxVPrkTYVefpcJb3D46SYH3BUbMqYaFgC4WZW9
+jjj+Ic0fMnmCqQiIOXCrwbURGVNgPl7CY4GsF+eUMvzDy4eVIc/SCo0cdq6XOG1Q67iPReu3V1b
rMTKkBwG0fgcMh/oQjoi8r7FIvidiAZU1tVYciIEvHJZQi2Eyg0Ie3P0/gXricDgOPnQmv5VbDg6
ohq2EhGRWiAujEp8HQV8B2VOepEuZ/oUnZBscu2A2yr6J/wXs6iV+nR5n7PpSjVjpYhTvCyIsSMX
3In/GMAQCYPedms2UYDGWJJT+Co5bPy6Um+rzdLuraou6UxE+BQfurRuT0syGcV1f5K9Sw5sSHRB
jDYGjQEZ+iAaAoNHQDQseDRm7Xvz1COt2KM/UoNGadHRr+kR/wb4qonsyI+VEzKSNv5XQh+jQ4RX
TFQKJ20XcN/jnVB/M8K2eegfxQNGL2kVPes9n3YhOvob2QBUiAnOQA6qpPOLFgPU4oMxTmaI8qMl
9fXlu4DQm76YqB2/IwDyQmmnmbchsJJmVJ9Oc0JYvX158B/kiHDu7Xo68I9xy5uDWBmDHeWX5jqC
YUHeCUOB7iiEfXslDyl7RTky4+2Y99dUiHtWyeXN9W26iUWi2xZ4G/ECJ2g3aJk60vii2w0nUkvq
1+0ANQN6gmuwZZER0xEEhcq0r7u17SKwsI8yFWyIbgp/raIgelNZz3c5rsFoopcOXgZjcrAGG+/a
seLISXP8C1mvmu6o3aXNVGCAUhjKhhkJfT/EpnoNQ7fU8SM+AbPWROll6E1/re/iSkn7HJLgExBG
XJ36c+i9p+nA5X81u+N4aqAqpy8oNGImyblSpSK7hlzkey60+JuMuXXZ9svlKygsYDbXhDXoj75u
N5uM10vVuonCImvxK7NhU8zwkl2y3TbRUZUFaPOj+BNFUyaRObb6v7AXXRizN7GWtgjWTFbLLWp7
cE5/cRUX9wNYfs1Pt3HJyz0dETXiG05aUZO4EgaiMPi8/JTfFy3FP/zSVjxFBzq50NnN7eHPf2/c
CEvFWIXnHm+aqm2QxLChsrxcGM6Qs+15ckd6sE1QEe5I1N5DujpprDLoGHfAXFJ5y5Vu0akeDyZh
JwHWYc+dWA3H6cci47s1IQhXS0F+5HjGL6cDyhBWwqyz7ty2T+Ny+yFGv4d2RlPYuotMq0lCJCY5
fInwmZVtcIEHJVsl+RRfhKZGoMFs8rAZ1qf9+fUxEtJ3uE83cXzleJOWjvTtuvpI7IMSzdZNlInK
naNscSzNsef4C2gvilRAEEBMemoXuaYiYZABxZbQwJUBPrCzGuWLM45kF1XvRin/CBlClWyo645d
jRHlPd4AZVJ9FRo7GGfISvYZEvckidGxliwo5X1wVA5DRqXbtpz02KOLpiL3XnFI5paxokptV5T9
ZxvZZGDqx88thytqoRZGJwUx4MIVQG/Fo9tesSUrQoST8oOOozBpQZbpTZL2FLSGhMDXnsEz952K
zAaVC3DbjDcDJ0ZWVgtI21ZeOtQn0M45QwjP2uI5W9ad/a2wyZX9sw1xEvXgOyH2p9uLjJ0xzYZ/
n8Ia8QyohozKsUMhgXXiWFYr6k1nPAfN9Yc5IeUZg0qruPyEZ8VHl5pDbZGJFfjNjdFzuedYnjJC
2SXODWwi+sbm9jP2sKuwxiDr/vU7CWeh0pJndsuGGyWHgO5+1OWHP89Vc2/BZyNb92W2N5kYHwpE
xp0wMrbciYJmCgJZ1HDAd9wfpW5Kvcr3Y/V90WUZpMbIGAIong09M95admN25M4UZo2rqcqJDNYs
vbdMPkvu3GcUdoLC4YioqkOzH/eP37h2+u7gsICB4Be1S83FQ2emCzwTUgnRe+8SBVA5xSWB8wgq
Lhd46BIKTBpLPrhzHTOkEoDm6PFMhNIBA2o+ViZxLq8Kz6h3xR8r4qDaelWtmeOBMxClvcqgf1d8
Dra6XXb+/7bb0KnD71rP7+Ymc5zA3g1hgGwf5wgQLSTBJ2rTrROQSOR5/7nDWUJntgrkJAH6oP3s
U41G9q4IE1nn+bIScADM2Zfd6aOJahf1X+6eXQqxe3r/7mzX8ivrsyYMXGW2LMjozTSH+o+ut2kY
HgbnZil61whW+Hfrnu7UECMlmDobkfzzq11A6i+RaQb4cv8NFfBzhriVU4qFVak1Z3NjphsKYtlk
x41ws+xcbXDh/7sFlk/2HB8Jya7V8380KaM1f6MfOueMxVeEVxoxuaceT+Rb25tNWHFEvvx6Eaai
moX4BtXOfYo//HpV0SdPfBMJ/4KwWkNNnhtOcJkJ3ToW6EdEF3kSG+KuZqnmBPJcpZwq0v2Up1tM
EGD0c2uWy+dcNSAzTzx4idzoX91efhO+PVkOfDUbeE0cu/FzQBvKb0+uiRHhOsGAn1qrQiA7q5hm
VEl9akoHVa6ceQ9P7NSiWDsZL4scrPHY77mtnUC2fY/9exjA88yJsWxs2BfmyUxtObtjQTFlBbA3
orKqTETMCc8JwGBEDatrmMj2J2uiAqhE4AFi+szU6VRClkp163AtK31u8BvczDRNhqlh2EDdz3Rx
qsPHqak7bWTf+auGaLoBf2KWDOSYKB+1hArJmdsnsUIIcWoGkGDSllWOSjzQeHoo0lawp38d5k7a
DzUHlg9ZhC5SVHwZRfRyC7PBFUIsLSyRiCONjgnmSIj6kAo4SMTo5ElbnxJRXCUaCzBhBVS3NVwl
YsBm5jyKeeWSKk8ayat6TyJPBlW/UGtkHGdjsexd7mHu1fpJGy2n3ecNbTHyZ9RmEvwBoCbHTYWx
gTE6Y0C2x16MnUMPV899SvSaNfnxbt5dQ046gkmOU2SyED52nkTLGRkvl+SsnkU3q2ucCm98JoIA
scf9Ku9wtL4YPfIEN/a7yecVMN58LQ5fZ7arjLG2QYbwm080E90EbQYwGkIX3SSwb7J4n6jKtOgA
pCHMWRn6nXyAhiv02H3RIeEo2K1q5OemvVX/LY6vbPsCj8nSZV41y7kFwIEAo0ilapHkcwQhG21U
2+u9fDMKslW2Mw2AnYJM+ATr6lCQPPNJle1Dea/5+nyx5F0DdG4+uV1+iPraxaf2JX9a40jgR78o
wdg25TLgPfaWNyDlbpM9Al32sd3/rFmjl6/buo3dvPzzDXeaa0mRuJd7LxruWkWgQ5DyKLDODTCw
yzE8GppmIzIhTTwBprkMmEkjJfM2wPlt79sLQQkPh+5UZ6DwLEcSI6YZzQX5niXF7oDJdL4/H4t3
oH8NHluxhDviIOSH3y/gnFzbj/xKCsZsqLEU5qNnScpcOcI4TEiHp3PMOA1khQqhTltep+l8+r1y
9ehi+ZKZ2saYRTtHaBWuVlSXkEk9w9KDmx+j+5NXeHvp7H1BMIg4W6w8+WrmQYng15wasUhrahEP
4Gzk3TALvtUwDRsZfp4lDYyu+JpyFHGCjIdfQEqkNAqfJkhigjkYlsOSZBK0cyz7Rs0SLjBQNnvP
lljSUQwBUdtuDFALU0Me9280lxqgzQVf8sFelISYG9QnoFfrfi9gMGHp9PcDblt+EXl+QMbBq4hk
hwabikTKX+qOE6iEDrb85V2SrhldH/q1RHUH2oL7UQ35liPUDMUYai2uSMAPnQZ9Ng5yAwxS6+MY
oLJSR+M4/N2BnU6y3o1RqhyloRuljgmQZ05rI2mh0sZ4yI+J/Tc/M3CVgWRCvHheZPfnNyEOwcVg
GTAZZlxD4ZaDNc8FE2STVUR9g1GtaPRVNkBIH32K8mMRz1fYAfpUD/0/qzOBX6Fni1sHchQUN4LL
OEBOYEQJOU/hLJtrab4yudn5fS16flZyLC5DDVaec6sLvHnstSiomZlI/M/Z9lmNJkeNAlP7Y8Sy
l7X6bqnxyPquP7Lqk7r93inP8Zg3JX0oZ7X55nwxAaqRIL9EezvFb8rjZPKTGl+/lOhqc7Dz2TOF
NjikOhZosPF09y1+53jykKLIjQ+PtHW7wXeU64whmQbSR6OdyzdGVBWjsA7CelWtAnFQ6NuxoiVj
eINpln4jxTDHS5m0qKJhnnNNN2JyERZ3U4T9BGUxaIo1U4G5flAnspH6vhGjNuRW3p29A4VVaWvm
CTJAXUlv6VOpSkF/uKfwE2jk4eMruG5wKe1r4D7ih8UIeVVw01vZUS/N9pMlqYLzoCTVWMLS4GTd
6YVbGtZtVoXk/Dw78OyqHokqaAG038icVdjtVAIvqKBusH0Oh0qxhM/SxihDMA2/vthD0kMqBuOE
nvhDCfyBf2TF1I6DG0Bjot7OtBe7Jms16DDrOPJyLMZxGCoNxvD9h5lbAveNMXlT5nN2csOAXYVt
c+bPY4qtMZHJmYiY7dMzJ4xLMVJrHWImAnmPLb+zRAb7udx4LsSDyyelvn1iMmIso2qHW1ni4vtC
7qzDQXCcY6eW6Kq33RNnQS0rMJXkuMzhCsLHbovr0NFuLcQvxqeXmypjYjaiGsYGEOb3Z2x6KR9I
QB2fsSELHNABLKPulcZgOJeZKXyJhZNiTBxyxBge5iqfeYDIfQa3c+b9ZMDzAMIzb5t3RvEFUby4
u4PJ6H93xubHtmdLZyc45Gt5BsVLJcDN+029rQ15Zij7VHc1qi2jLUxtCl89ZXzQE+KNz9kj+Olg
wHPSZNjfNsw3l6MhPw8hMUZJgNSjB3EGohgd6CLpApOKwzx2yIo3AHnjuiuCIv3cooFyavOZ8GlQ
vipFVy4DITDtpWnYaX6yf14bqmLA2YMrglo8/1ION94TzURyURZwjKn7khZUOv8omr3ICwGdDY30
uGEiGP19Y93Am1o9PA47L8U4F39Wdv6CTvnA+u8FjihAIs1tJFhs0UW1Bh9/+F8VnwTQOVA/kQAJ
gLQuwrz+VrSpwEIqrUSvIhteY00GwatyIAmbEPbF+kB01bTTdbXLaIBP1etcAm1W7rbWj7b0NhEK
6FpUtqXpaCn1Gc/uD+hdSS4ClDS+Tu+ONLyq/a4TBLACkG3sH6fmfBjFlYTsQhYIacIxmfzYSYub
X885izHhz8u0r8tq1gjKIjYMDusNyEyQ351q9kF4VzWAvl7aQalr4vq4jSFG6dPh7881V8s2T7Ko
TSSGz4fbzx0DF8DOEWuu6ti2Eq0rgw8dyoEFjXSmmMDkGynfDfJ20G4twkQPb/kRtYmu1q8QH0X5
YDlsh+VAqyeMnuSXY3vD+7M1JbrnVAnnoZYrA2TbjwRnb4sjBuFVo1qTrw2QH9ClMtbTU+zrQcKZ
TS7COzqe05cKVkVVy5+p7BS60mQ/dS/qCpyh95spbI36Cs8HVHUriDcAauAjiTO3AyyJtQS8ywPl
nsYuF7Xma4Uz4lSxKX4qItt3d61zMpFUZMke04cjPrJ+7y3LQ2oGWmTkyYNH4aTvmEWA41gUp0bB
SSs8g7y2Qx/A1li0DxoIcRNPJNh4EoV8enn0VUMjqRwSUrF89rFD57eosGi2bP8j4T27+ZlWC8OT
i7aohS8+8DjivXMQFwaWOFuKi4T4dEgW1QwSwrSzaTpgxO2Uyj+iDjR45NGKKiVGnmhCX7jUyp6k
coP4szqc/hgFa9ImP73oqiQmvtm9SVGkitXVtJ3kWb/pHj8skYT1vZQoUZT2I1YdES7FEGq1WsIu
OWHv8f0YbA0F9hpfcnMrK3kPLCtqhR8QIcTxXkIQghNxFQ5X7SRIk7HhpB2QBXivjvxB/77p9v/i
W7yZssMob1amZRqwnNXwOH11bEi7Jt3PCfrBSRL+nBeip7CAXaw/nCnccm4mVmWAdiPkVxhZu8/u
c6P3/7UGtjfKhxy97aqemJKLGuNXo7sR+7S9NFxatENxKs8snSL99G/plzKRqK0evJT8YQw+Ispt
NzgU15soy1486EMf8dBZmtMA+TwWk3zBhutsXVea0YwZ0YrwE12koEf3W1c0psz4UkA5PG+cu+La
FzjW1N3lZREFxTHbHcmF1+eIl6Qg75t2ZgIgsK9AZJJDt9WJh/HVddK70XSa1nyjQhrL3O/Ue2b0
8oH7de5DPpwkqriL1eruBgOcOxIwA7M72JM8mtDE9nWa8mW8McGIuc8aH468KGSxhuNDJgkY4gQ+
3RD8IfpUyoVkOOJDPfm7q5SD8E6gi+tjTZXroItfLpXjKVtn3Bma9xWVLmkYBVE5mAPD9YHV+AMd
i7XF8/F84jJvV7iBUYa8JMGRAQXiwmnzwkvL8F1X2CS4TvedS3F0jBfeIAZhi2nFEOioABPIE3vN
wfP+IWxlusn9rfGhp/nA6n7XJQqnL9zcssVEvlvI2CEbM0Qz00jInzBdOYZc0D5ufnw2yUrJuZwl
qYYyYOUnjyCj9MC8y4lienl7Uzz1MpLFQli1ndo0+XghiJ/DiuNwb0MlaLUwV659XhcKlY+yz9ql
hFScQY0E9tte9igi7r23N0jQ2bGY9atUyeelpVch1i+XeOpoJKz12700OagTJbFgyDxcKuKRNeOZ
lCwu9cB3SE/a1E/P35ApnfwPJmZ/ICngRCTgxO6R21VjW6n15G5Lr76mqkqM8cf2BOTpNz9YEh1k
PZGpft9wEBFLxKOn7KjgktNp525cDa+0psgzEIDOInr4STjmHK/xBpaY5g8eOSmT0CUeeB059Av8
WLJg9NBfCDhZ0UJ/h8XL+uX8CUUNgy+Y9MoaGvITgKhMhsKjeWlXmVUXlN/I5X//BrHyU5WZrfKn
Qf1g0QEHr2nIkjb2ztYF/fn4rLtwLI8TPzV337CbBCQap9Yl4yEvtqVUdEPbxJKoL5FiKD92U/7j
xe232KF2n8AGWAfjS9axAlU2fUcRCyevHf/gxuYtPO63V8Oejips8gs2+nIh5B7XFEPfJASv1K+4
WxI1wRQbgu1mN3wxWf1Xpk1mXtfCIng7tPEo6Q5pRB4UaJmxf6Enp/s9R7hOKh0VXj9FVcAw1aT0
iivncv2lnU5JpSwUOoYuUuHc0a9eHYhsZxjrPgI6QE4PxIh2fRst9vGGY4GS2XsqBTFjZNyTkwfy
QFXEEsxF47L+tfVPwKhiQ2hvFSSq+061oKcKmKOn+2jLg7/n9FZT6dkdfcFv7sdW1VhHzUOYzYzk
yEBi79bDbOs4xzVEddzCJkiNacTttyPKuF1U1FlYTn/cod4uMfdKhFaHr1qsOU5z6sF+MH/WEEeF
bT4vpwZH+RvXDaTNXTjAmFHsIORhatRqU0+cNUJ2EPApbnHXtpqo6lkZd2yRPtuPL6vgEEmKTOY9
Qk7rTQAUfZ68kiaRNML3tLrH0H09SVHJXbRPn8tGwJ8ebEzKe0qVmz44dyYK5pA4ZDeksw+3eXCo
ZSt8fj9wzoHJP1M8T3m3aJOM6L4gdTsKuT0OpdZhm4RboC7/faLeRQ1Wt3L6lJF8WQb2oPzYcvyr
eHPtr6AUjaxJr6gi7j99QLdWU+CjA2Vakn/MP65DYbmIlulPazblWvWm4ofULlUNrHse0b0Zpl+1
nHvbRzxjDO3ORbgJMVRJ+/cjbCb3YvkgkHcE1Y0oqQmxBoDTIpUoN8glVssXsUfaoLNeYh2qotZp
3w/DWMEA2n44pE5aJ1ZaHKy7ceJRias7jKQU0fK4y2PRubuLXtARr02RMWdxPX5TPJZBtdgq19ZD
y0eQtp3vtwd73HvIYR1yBf2yGoCdgJF8aVsS4ZkZJ1b/LFtxZA8/Z3Ak5TEW4BxaNivkJbd+IIDB
oJg4+/O/comjiJ3jcawUvxt9OMGlS7Qd5Abut+5W3U/AzQ7ViH3T1ULhbN8i5ycVr0qGcsPx2T1t
u+A2HtwBYcwyMj3tEC9lBfu1sUZ3LAlbTdfiFCM1cUPvsns5hgxxUlm5hUh4OEvyFLPhOTS6UlyG
5ZVwkMLgdB4gnWUYhL6lFsxTw3rzajbNKpbZbs4Lno6hVfjOwty4XRfkGjuDfyVWzLHK+Dx2SvdW
hnnHd6bALl/8S9kKLjJFjXcvvLZYEs1HyUXt/ziCHw4OZs5hJJZPJ3ee+MtKvrToABSnL2wq2zyB
d50d0XtH+VqOgaBAD9m58s4d6ja419ILncCzxVz6Jl2Qee504H9XqYDnfxecPWX9mPVUDFmDsuaD
EMLeBUvIwuLLHszxns5Ab0mK73uYPsvWrfrq462VNBrAwseLTgWd+m6qz0au4/HWyDhWiSRiqEas
Za6SOEqKDBhJ8VlVgwpJn23MGok7UUZLfRHoYiSvGcWxTRwIPRZTMIO1tUxBHjAiVmJJvPrLGrVO
ZRvLHstP3nMQKSW/jjZ9vBhxgUgdmCskFn6k/5krSZFqPkgohrc/sNyLcGm6gp5p6BFqMTM1MpHs
LK2Tu25kH3kiYwQxc6+vM+n9BSL6awmqZzlDDadAnPIiQXHZsoAnLtayWw80b46cPl5/HBZE4Ckh
KpEnW4WGiA8gXCuYjhrkV5dLxho7RChK1VcbyLxWEVjQshE/y7kkZuI1XkGwvC6OVy4cEHq75Zox
GpO+BvBkiRbxnyXIyQ8JGEzv9i+nc50crpoNJJm8u39GlLxCYVapo/KphTlReK6lbUJuJv4FXtWH
ArajDyONetg7seRgmvn2/mTPumCubVSJi33+fGRcmMdd0IMSLhHU0jIoxFzyQ2re+pb9Ni6kAVn0
49f0BM4H7ezNdhtnctU6QDrmPWATSDLDrzM3xRVdgrCDLn2tPfz/JJhf9VG+UOdtXdIDWoFWwbgp
yFvpw4CFc8oyhf+qmww8Ahk5sd6eZYorrWazHcGTeKysQPPZtQnq8MN4LqzD/PD9XF+GSXrBaY05
EXkE/ExXdhjilpwMZfwPFoWAXW46XLl5T1eYKt2L+uVNmD0uRfDVkUMCS6U1i1b6bNkre//VhAH+
Zyyy51WYzjKQ/sf4ODGXWd00Kyi8fYv0LNN+8P+hL3bbtUamEhtALh8wk9Zr5GffNWg3ERgoW7k9
kjbYvLFvR8adbtjR4GK2Rq2BqeG6tniAwj5bGmFwyQFag4/M5q/xnsIuzW1fKk3OtqQUooBrNthk
0ZSxZ8jGAgmdrvLr/kg+YJS3EPj2Xs7jR+DSheU79Mv/YtirhZR1/94w0mVFDtQIXKvANOwxHNlc
BKcTyRmD+0R37h6ik8gQIgetNdIEeH6ZPunQMU80HXNiNxSTaSgH3TmTrbvaL0Jh66CBAQi0Tvjm
vgDTYSHjCqgJX1lGZiEodgGuN8Q9LxXcyxpHhfaAMVLrazqytsdJCpjigWA3uvwF3U4ZeX9cVd7e
PFUjwgcTqFXdHSjuEvTkSnsLrhxAVA1S1KY4M++/RV1lMT2sUiTyxpP/Q2wia8mc1wayhHz26KyX
UAIhAeqp52Y5cs6E5wAt+XEnXyKWpvfYJZfjHSVOmlZoNZX198MBfOtc3+qO2voFK/aYL+V3eA/z
2honUrjD5A/UoqE/djYRZlozIPhIDxV3HFPNQBCwovocZS0rYUYcmuP3bbQ6DeTuL0CQdVuETAJU
l6cZtSeqsK1SruM50tb7dkD583fDX6Byfn+HgVRA4uu3U34Y7zWthSN1xpYEXW12SRo7tdEBlkq/
ULJo1eSPTTbRWPi41/bxUKMCWvUe8ZQHxfrcSbwSA03XNQuNsRSQZ6BfXZGb4eV69g3ytxrl3nQT
bRYYWVcR4pWhe6IuhrHBlo6/bWylrJ2bTvDq/Fy0bjMlRx6poxiS0awViInMxKC/hvnoc7q45ASc
zZRLXRmZYp0Bl0SvRViNBK+mgpg/29Yh33FTY7MZwWBdZcXJ1iUFX0Aw/loEgO9RufyT8/3wOuXt
8ebWVRZw/+QnNUPR1WTWuOoR8ahAeTyn4lt22h846cyctlCw/FuDEQeY4IutI1hWaKtxnLcSsc8+
Qo24iNI/O4anOq/zlW3mkIsLmEtzvEo3dvxG7d6QdOovoOZsKWW/MwLS85UEMP9a7OTh0c20BOIw
JZlzAYRE59yDtoajI4yopc6tuYLW2LxdIGMbyCPEnNB3On9QQnfk70zfl7zEOqw6cHlMKIOhb57e
pyysQW2QQJP0RTxVU9bXp0NUMvtZFqeosXfaxNF39R8PtfqDMmSm/j0G3R1C4X/TVk1aEpSQmtza
6RktV2dS++2yOPDabK5y0MgLyqG1s0g9XgSwLlNufk6CNEoONvSGxbiYhZob78uP/ArzODkwbppU
ArgoDKkYfwfXlsP9uNf4KoPymJlWKRifgSGgfsRmTu1ZYmdMDmrm1ZnTRpwBHlmii4HQ2ez3E+Cf
UP1N5N407UUt32suDxHOIj6WzNAZMKrviuVAVgtSqrV0DGvpY3Yhjjs1EwxH5LlOaV7Dhn6Yxqiz
mte5Vqk5XwkqVWkS3srkcvBv/hs5T45h4yzvTXnoeEx+w0WPRa+fNFQjtu2ZWIPvIPOZjM29HrhY
03Dk5fO/cQT+jyyL0AjM4K6g35WUWjflihvG6+OAkKuFLD45tCYSqn9HzqVl96vUCg1VoTHos9Ie
hiHSqMMOwqloCripBrdDO3fwNjJMmWizGNBtVAYRc9Ry/PcOiqMn+CFOlB9K+mu0a5c1/E1EGqX9
XnIIADjVxaR0dHQL7RdJu2QeSAsG/1PcL3b9lS7nxPAutH657/BwnYB/GSzxqQtx8BY5ExfLaQGV
8CWChccjF1nWqC5btE7wS+b+Knq7SqUCFiC/7j9Peur7dnDcR4XchAoHCgU3aewVVpkjdSIXvtjO
Z2uduBJMCmXCmEkIiQOxilx8Q5+iyxtLrapI49pFNOTiCXgmtPj3dql8ir0udHCVyCmJK+/z9MU1
3OL9Zl6DHWnq+VJcPo0MipJMokk5C1JlouOeDNGGA73P/JLquN+euFmkL7Z9hv6yJJleac2YjBXV
OZsMAgi/jxpvLAztpjz2lG1sFyfOEYRSTy2VlKkg20PzwE/55j3ilIHz9W0uEB/m2jrEIi11T1rR
SNVT+NN+t8mkyOE5OaEUOjj1rMOwUbUbRRnwolyUtbiulKbmAYp8sQuM0rIkxht0tO50ZpU/q6M6
I/vFHlpu0DkbSp+Rp5HUVPtYpVjiLx9txT4LOSHqcpRoGa0CH861bTe5NVANH9+mWQFIg9NfJQx3
3Fd3gR6TkOkhfiWZ5Gnu0d11pl2FcgAc8diULNucHQoH1Toszl/29UvqGY5R4csfZU6FFC6QnDnc
q2jTHGJFJ21ug0UmgTJK5U9SuA3m702V6oeKgg3Mlk7woh2NS47vme6Avhj88HLTKoJZOgWFDeHO
FO/KOmvsAabXzRttNlQXWD7QYZ5OXaTZ7zvM32d+zLpIR/TXjMkyDT1Wzz01mpaxZoORk343Xt20
y8fDYlqkQxM3V2GBPHUC/f2D1TNI3jx87UsD3W7+zbkBQBOZ8JAqb5t91rWdh7dN5kCkRnGjTj00
K8E3GYzV3lQAAL72BS9S0FfiWY0TDHOLQqbPPPUtQWvBVZRsow0A34KFOS7M2sY+sG11rsbgqkwf
fkpV4E0nEJXrrkOXAFVj3Gn+fXYYXdkNQC1FBrxe8RgpAB3dv0XLIU39rN06ZXjCxwKcBdwz+wxl
L7AjGw/UVEm6BqnqPBae2t6j5PEhPIK3bx/yDc8hiiPWEfVS4FHvHNLm7RLA1/+YrFcVgChtQmic
+mAZLOHrph6Cna3NVNW7u/yMyCKFU9Snh0scExgQE+xQq3fNYgCDcm5fVufWfYBB464B33LWozA/
1UWxkPmkE9Ehk03xhHccyJ4p8LVqVZFoaqn5zvxUGq+YhGy9jzJaVdtQdqTJPu304pIJpqJ4ETqZ
QG8AdN3JhwaiVf5c75BtlSnd25MZLHyLXzDw0PPXRWzE0Iykf63Ccn1EEtdWg6bIIw2C4xuHVIMd
/XlsFqJCIc6aV6hbbW7wkuEo/r6aQfYtZSZPwlu/tYw64HTx8gk0uYkvh4cG9rTDsua9KK/gZ94s
m9TAsR+biMk4ps/W5S0vkABC94KEDvT1aejZC2o0GEHqr+dfmtwd3ZwvlZuRU67JKja8kDVw96za
U4rqtmZcwfBdulJ4Fa1FdowChqDgS1iMYK2dT9+GdONo/i19TLutOntt5m4/YPzK8MDlglG4Ce3l
6kpQFLhuyR8Nu7AROe5gLCe2+SzAmykPvoElpBeh7mj0xCga5Yvrl6MESZCFyOTSCIZAD5+Qm3Bm
Chp7gIVXaOoI7EzWgxCeocSGVP/wniXqvQnFzxh1ZwyaG3OOInLLmRpyz2iZjiJCxxqlaaEStDeC
NSeczLml4v7T3c1O74RlRVJkR2maP6M1KxnRSTXU4Te+Ud7AjZD67wCok/MOPqE6+JYkl26Zizho
TMm4g0/1Sg6Y70j+2OPxi11k7szdqvfjzA3NsWPbCjFZ57BtCchJLj6V2Y5/L/0uLaYJm8iRy4K4
ZzVr6jyRBY9aSS7tg6TOXixvSTQ3L0G0dDLxj13LAg8B1IcXYMsd2+ddD159Ax8c5gMm14ni1jnW
kZrJRrlDymBtARmAEGvBnxGcYX5Sf9w0dZJrC+HkGPIr1LOeyCRAIBVxeiwSj+zfwSVqyBQu5+06
zNtFt6NAm4i5rA03tal5pQ9PJ4plOKPQ7JJHfLXkHAT29FLL5JVH9o5R5GoBrEeHWYKeDZ2tg5Yv
LcGmKl8vqGhL5++ZmxinB+2itJRxkHadWAZaqOno/TkDAjvpLGHmSpPF9DVlQAp0NYm3TT/1+vZ1
7Y8dYxk07I9vkwrpQlz5zjv39RDkOoJiQv4MbIkFqvo3JI+TCWGQW4CsVPIuOrUK4EaqoPdMXlep
RaQrwjMVbIy4dlK3KKHvZ+r5iyjjyimBXKSGF17ajzDV/ERxxWV9xR6saqr9oDBUUm/iGEwzQZS4
NwzrwvYCvuYkUPf71WGmKUFRGGdOsT8dsDyGaqhbMoQDZZgaUWVwWA2MPDc8oznFwEp2gcEGgK5V
aUSYbWA0O4enjzco7GkZdB8F73K45OMfwt8rBlZ8es8+zvh8ErJb+MRzM5bgmIjYleynelFYl4WM
r2pglVjSvMfby9BC36MRWhxUwymC1e/HR36tSyXYLQ5sLK3ce1qQKls405Yfx8i39S/Bws0t7q9M
pHFzNeHOSBIU5s5F5ko9cp/7ie0MUPGQutLmIv2fZLTO3o95nho0aLdV8rH80lkggA3GJbS7CbnC
M6CGFGOu5W4dTvBu2yS2mgIVLnACaenOap/umXpkIs7zriw/o4gwtL9x1qT08uagZ9bJ1Z6fvLzR
TeIhkoni4U8FwpCTPIv+miTO6gK4IzH7iu/2Now/FXumXXTgJz+4qGDoJcZ87/4YHaCP+DkuWl2j
DZV7vYQGMzUClWakWMmm08eNowzgeOdAsQUgMZT0bUwfLwFhZBCmZgKrJ+Gp0DbLNg6bDMVw0gym
FOEKC8lGhbmWPg+SvIraFsP977os4+MBP+4Liufum6qa6cyQSyzuhR+hhJS+VQo0yFlohL6Ma+E2
4qyVdluEEDCTdJTbmyj0xSQjZoZKKaUg1wQg7zOOy5k9yClAYwO2r8OGEk1lD9Tt90PLnGpJY0qj
KhbGeoRknrDLraDD08uSCdPgZTHOHImoJFOjp4ryZjy1MujyJWvW59W7WKXZ7c2hde8QdKqrSyZ3
vnYBo/cvuOIzXSEWFS7/GWFrAPTFXHAoCMQhd9ALH8Mv9jCv8CCKpPsJQtU8ZRREx7mgFOZuB+fR
rUl1uZXVHUEkv63Rzla3dOkPUwLKf7lw3Ns47uIQCP1P/JgUux//Fu4jKWBrBwy0TsJsQH1fMUhM
xcAGQMyQz2VVLYU52a9ORguCAwapjNs5h49zHTJ47WzpDZTjprM+qs/M/cCYkU77k0trkTV995Vr
S0+92Da9oOo03Ko9/GxvJ9C4FHd+0uRdk+w9cX+qJyFd6PLKjK7hg4LAU3y/rFRfQr51Zwy3ZKYJ
iMrccM1Qy9WSCJzzHZ+vc29M2DHnEvfw4NtXioxprc5q/vxwcvQag5h5cuUPq2B1N5pj+QTumTF0
pkumvMzjlbLWimro1LxUcc0qJGM2zhWstD+DzAj1qaxvBbZeDbIelJ22CFF/rxydlwiWy52LZNzd
1X4FKnpmUphCPMXGCHrZur5MeVXYFEjDlUCDZwPCnp3cdJNJopr8vM6mbngo5EqP8OCkmCxC+lNl
3K44biWo8A7CVpj5bx4/tJTVQISGEhmfrAXpIIU31Ejjg5eCrjE1t2Ef707tuJv0DvTMOHZNfJyO
tcChbCqTQqkjDGMz6y1sPuTB0nqbOKGQr9Ory59dboj6uWFiEYibCgxAvm4fF0ontoUrx8QeOXBj
YIfHuW1TtKFuSmxZ9Z5Y1U5rHB9E7c9+OqFaZay46/EXiDHv5V0ya1CEDQaEqKxFzLAYTmxjBB3X
h9YJrQWwPyC2ebwDNDUm7w5iZt3LH+n/30a/X8e7IQLENdFl65uXQ/OEbhnWgoFH1gme9RJ+sMde
Sa26qdKcdVAGgs5Wd0asaGTufn1r86KzPkkEX+S62agf+5mahfBlvuvXr46bxQuFdZ6qpPGPpC0s
I290COhGtXJJdMUKf6sqLEDC1lbpfiEt39cw4rBs/IUef9P5Ab0eZW8cCtRQ9yEy0RP7gtAxGUHy
jmeGn9LrThY9Gi8G5zoXvo45qEO28QQwGOHsrzp+bvY4w1hDHE8kFAT3qbZ5eQfh0UDITjy2EoA6
nO65QqpQdoRxXeVUhI3ibZzx79CNBETtOSJs6yr0cALUXb7gI0ZaFWgudK68WNFEPpmz706P/UJj
YHS1A/XPrThYF0yww4mbCweBZVLDcxCKYUI/ymYOaIgIPs7/3bO18Q0bYMHX0dRK5mFroR753Bni
oscMcCjstWpaxtZkFDgeMKD+pQmDOaf6mONgCDe/YQed7aomSqglVfbYlog6Dad7c/OVMI+xYKrn
dB64/qvMo3STV4tvl8IXcgW6D3ZsBqRbfhFEIIqfPr6OrL5XM6p2vC6l80veSEGT0FKx6CNRVSI6
O0mOd3z2JegBIefobUnTqZGOJm6HyHDIIZWrqolI3Xuf+hO3XdQ1O1XGfKdT3jBizEUXeggyj4f6
ow2r9gAyM+kxv0N77goQ2lkV5EWvfQtAhZKCsQO233FIKm/k1UNzYcdBq9KwlSGB6gIazfdM5Aph
GKULsSFq4MIzL8W9idYOL719BCrvtO45KZXKThv5mrH3AevZQOF1jZ0rr3QDVLTxHppcuXWxNC7C
RAk5qxxLew21YTdLGyLspVvMwQ6TuDaeP8ucnk2JI28sD6vQOaN7GDnehVfgRswg1WlUZ71x+vOh
a94r30nstWZULQoAZydwHn/hO4UGHjuy/ym+/88TCUrgZMnOvWiR7tfq2SdF9w6Vkjukja02kCQa
1LKp8O7a6atUPqoI1baLnx1RbmJVYHkjL2EtWVA4lqvPR+Cy4qU1qJn8wwvYgg2QFO+BPyrJwJWN
U4Ldf/8xvH0FLwWAVl+54DXVdbSFWooBcl8lzfi+caU6VAFO/j1/8r9fjuzprFNBB0tLYuzZNJ3r
dGqGZxb1jVu5qWABT5KrjV0k5SbXJBZQ6yez5wso7UrBqOYHCH4b6NTV/j4m33EOsKI6lV2nZpdd
8qTL5idhqTmf0j/RHZ50h3rtGq/ovVi8aLE2Jvav7y11821doBh6ob3EMC56FO4bqdS1gXywUv1A
Swcn5vVMJwr7wV4VFNlf6nTYlbwr3rkfZkhwtifwfJCIXKqUmo23uI5iMQ1bjS18Kkp/j45etiaj
+8V92iVRmduh7ouA0aoRp4+64Yz3cUB47pd3Lowi/e/Tj4d9uT9+uNPLEF/7tHPI4yM+kzDmXYNh
x5dgGoUmzM0oY5YnodNYwoeBsKBSEfPrFvCn5t3KYoubKDA/WnKOvif63wRkKDsWVdFc87PInv2x
WoOAeRU5uPgviRTsD8Da0uckc1xXcFYN3xwfXIjQtSceGC7pzFOnRiTPrUpzZpi4lTBtsGmWZvLs
pslXukUVvrd1ZtLcjsHKmvt1FZSjf+6OlTWMbhUlN4jEpEVemugsOxsxPAfBSuFfD+jBLZPylhL7
Ayv5AeUN8GYxDvqEC1LFMOOBgWxbvEYOwg/FSZgPfGWfxhhUmqh8ClvAB6PsVeupQnMX1dsF9Iwj
Xq1N5cLLdWcFP6fqNR8s/JSTRuQlDK8l9buwwkhvkS4Y4kLNNBUa7ZgmkKXPRPOnZVkNfh7geSH0
sHIKTPH9aOvQ/wPBP0LhJ7Rvo1EiSqwzWXgot80YD2ajsVcWgKMMMamJLmPptfOhUu8spotZpUrO
hwV3FjNaWOK2SLVCh8uCTGHmrnVdabUxAtRnVkKCLfiJboSKTRM6jtAdcVjTfJBUGk45XMo01G4B
Zsj6XEMf1WHCnjgkA+b6jpWjG3nCxcryEXp2f5Bd8LwNdLkKr1RS6VncZdN0FKJCSRdDuK4uKmVV
xgvGRZqdxpucdpcWi7P5ypR+K/Lk0NNSSjVMF8Zh7T7MrM3Wr+l93lmxm0MmFAfiBr8JSzZjfA9k
ylNu+3dQNps8rwRpYOlkqUNFsx5lqgaIgWev1qPjsFmAoYib8HzGHa+FvSfLMj/LFIy/jQIz1jKF
MgQwjf/2HjhK0CBrUi9EP9EwhJ943XNasxHdfp9iT0caDtQk9/iT6FiOq9UAqwMMIJgYTTb3j6bR
t9XGa8V0RHcWFqyXtqyM6dOh/FjFxbEbAA6sixs98nvQELDmD2tk5MAUrr8xPp5VlM4RiMBW7K6l
jXp5G6wlMwaUWuhfpzz1WtZVw478MnO5WjItRQWPtMZw1mxWx0xGF61rt99mxUOEXdjtnX+Z5BGZ
j+BSh/cMqVMd9Y6P1ChjWs+7/cWJCBYUtTqCQq236EP/pss9e388DA0dMjKTABjjoXvwaLSgUMXl
tuhzgGTO/8Ym0FcucUrBW4WIE4miALWd4VTqVON5q/sifynJbbTLvIMtEcyWkXujLWMolphhXPlf
ysZAZ8rzokdzqFoAEce44jhb6rkJMu3BHF+gJfUfJMWmzXzDI30sMOK3Zesz5N3MEdEwfZpr9aeg
mdhhrBr6eKub0YQ5bNwwMjbu5BGyLv0yAwPPr6srpqk2MwqqPF0sseUN3z+ifJ1KcTBU4mNDNZWE
DLwlZcKeqV/JHq9wAGw+Vm5KhHPWnfmRllnH6mDPFeHdOv4oxuDD5uzKuWd/SrmDF1eK6iuPf9hB
3Sr7fxqv5lM/6+litoceGTdNJYqLtcU6L+S0nqtGHu0mKrTKOddM0cDnLc39cY1Gx5ebO0kYZ9ou
0IztTf4aJ1VeE8j2/GLqeUD/kgkY2TgF5b+9bOUUZuip5HPllt4QKzUhXOA47edfKmNkYNMWEt1Y
sQ66ATPMpCgOXEJpELyem03uHFK3HQksLAqchzyvhL1JyLLApCRe1SWqbD3O5A7FOEiTuogiSc+p
q1VRQ4acGKhRuMd/35VnJveclY3RmeJJxT/8jTTAsVvcX6aYzUHY2mtC6bFRblaUGk2Py5d4rSkJ
yrBpud13+ahX8wQe+KkW/x1uo+yjevg0IJXOgjuh3KDBPOd1IaeaVJp3dRiYAWGPNkkuirYXGFQg
55PoCxk753LqAlOspr2Tu/Rw/evZyHi1OX4jezCvb7Xt88ysGBqIzEcCjlNAfFrGFDm7Vcyz0sc+
UJe4YgeeeOm/bEajgUw3skwqdgvxnHKBG4K286ERtpcH6UE+BPIVMVgDK5gzMwdSxI5wHsP7Zem2
KMvCwDhI9uoho/oo6gJhxZTuznWdWX8w4VawX6vQR80EtbRMvZPHMwzZKpS/yC1ggtM23BwGriLQ
LckaD4Kjaz0LRaRZs+SNuso7xeX1Bn9Q/MS6x8/r9kJ/VJ2H+N2SdbqeDBn+xwJB9kHwU7J1KKSm
C2gXV73zIAtUTRSn2sYnZ0AGFVTLTIxw+ezJqF03oWT31WPoROLEL1JBheDKz+/w82hPJ8D1k2Uc
0YWiydZVNJ7Dm7d83ziasLs3rGpebqIOQoPaukgbwnXrYui0L8T5CIMPNjJC0RNxN8Jneg+O847S
s99PCJ+7UH+khS9HhkrdgCO8SYMwlDsqnmfk3GxPWXYP8Cz/qBP5MTbS0UBNRxxty+4OKWYNQjqt
9XOZ3b4NyZImh/2TEPkY8YzvoxeOOJF5ePFgBNTuanmL6WkA3bdTpwNVV+jfOcm8JyFONZn0gJyP
MZsOPzGDmoNh9vuqBr7ilbdu7o3oEemGHm2w0SsXK9OB0BphGnixupzR2G2peX2splyG3WU5Fznc
yXkNHDlWTR51DVtSNmLP2I81BT3+hPdxScEXpnVqCOYZG0u+14ZX/jFq6f2LyuQvMMrAjY2wKwbb
J5+kdXDQjiD/zQBfZlya8u3E4/UBnzUWmUxCHHfI5IAE2MIMpothT9/HlcW2T8KRxp3Q47MbPhCf
phSyz8O7tvjX/GNUZczVRP5Fc96A5SPN76hy3vT+dU9npvxQbqFUUa8W/Lu+ohvS0c9G/jVzJNEJ
1gVoeoFwqm6b5L2i8DAYJO7QjvGpt6lneyCJe3luD6YLXYpwe/Gq6oBlVFT8oq+/iOCtr0F3G7lD
tPwvmjHeIHjouMvXZZh0ROrG4y9douOYJBk6c6zk1ltRO282xwmZ5/NdL9r8KOxkMC1QJ1h+kf33
BuytrkugsFKdCgjQX2ACwr7N3BNolxeH1Xhoj/QsW6JeCJpYoY/8L90IbPoRUp6imYOrAQj+1gNw
8KfmrvrjQbwzDf1pnmAATHLBXFm7V4c10V7NUDCXTMNljWUM1FuxXIH7RNvIeHSbTyxj4549+ibg
qYpJuRMhmqJGEpgQ8kKdTPgkl9GvAjhlK354DQMRq+vSH6j/D0huSvVpqbqovF0WAPpVYas1NDmB
vzmr5xWNzgeaTWQuTIFVc+6YBCjw+Y96u/sJt68V2Joyu4Mm4kBmI1UTDMUqJUGeHiH5G9MSk3Ft
vLbtvpjKGDLga4MfMViw6/IEARBhfyUeCsekVjsO+7vWX4DXhG2E8cve7YZiMj2Kb7bzO+T39Efn
OCEalkR23oGS0jTaDc0o7UiqRwLDuCEKEkSWS6k5iSHPNCSa3H3HVOLRoA2nZOs5RVrBqBRv/dli
tndz66u+DG7gytCEWTglnvb9aHyL6Daq0/0VJzmaZlscSBE7dOqY94sf8pFozLPx90LdNyId+20V
wZxuIeI77m/g49PTvIWEb3wDrXlq7zO5+11Z6Z4ZOsPUZ2VnFMQ+YEM/KxA9yn6KaJlzncHax2vF
g0QACnzRUfqan47pmc9pKZG/dsCiRAWdNYpXv5VEppRkTjabu9pvs5oJgZr8plDjLuHupAig33Nc
gpgFz55YOPgRjgClJqSmKHc8XNr2Whzb2XMv/pmiIk19Dwfrt4ftvLxnaf1ZVkZp93ZCpWmwl4O2
rY8mj/c6NCso+cx0nGO0egeIMEyNb4Br3dTR7zoMzFDoCUTCzIq5SDOj/H9/AE2zxBLnFCrdHfCa
TwBn39ZNQV03T17Dv+wDtlfBLCyJ15TJgCPSEdG6i0t6rQKJDWQGTEjJbpLpGhuiVRCruKeBkk6K
dZ8xlV943qI1yHSTIrPYClL73XwuJKFrl707u3ASwykvio+V5UJ5pUg+QUL67PKm1fADeTQVrZTk
dhvxiUDU7nncm4qKgecop1Qr0EmrUXBXUor0Y/OwSGJibnJOqOMDniM8RvDK4gSO2TTVrOXUUeX3
5JyGyoI9glZii3ITkCtvccjg5XK6VN6HOpe1HWUwvRac5BJl8ynpvfOQPnfkRVSkxH7Mw8/oTNva
x4IM8ie+GDvFanG7/PSghlUFnHgkwpQHy+zrtrc3hGAZqqjsdh/f/P3zzSmuvItV2eEz9doUJOYG
5UjWrUC/k3nZQ/ctToOpiyR2yI1drjOZ/mHUjI9zadtBJgHV2gCDBY0Obuj4vdlcO0eZh77BSI6E
E3V8CBwY7zuGVuGrcG9CjArlUiQgoeYwT4m/VB8qCeJzvSz68Q7HJ6t33U3cJ4eXWSc+hIHpVl6N
0fHiddMqqmCSfgr11kcQLYtL/7nbRHqMqhR8KR69ekBPs03oL7RSFuMbFGJhAN1PFaDcddVM1/M/
MOiN7HESKiDdYsvEO3YSHUy1QzzeZY2iDsHJvgkCrFdBf6FzYQ1hUSfRb01YvFmf/fRpcthER4sg
NHFHZhFbiVi6KEgSvA6cepz0Grsq9p7uXeH2dWF5wh/x/p3kRaWezJ5SQl82WHJaCK1Agogamlpf
NpB2HLOL3LoFgP/qzO2OSU8/+TjfGp4wiRgOuDTiFVBeT+UzgK8XuCGunO3kpOPupaBzlsQE+h5B
NAT6Qwj/8/teBdyXD6aT0zqW0mDTmuioLVc8inIWXfbTIgX4dwwuB6cHj8vXGCFUn/RWsLbDpEG1
ynAcWn5LupYVPlsxYFxrbxIDZ5lB7Mw9UL2VJRJ+BB/3UXWvq1bl5qTaChoLAnOzqBNJHuwE9vhZ
uI58sbqJGvcXbDqdMPz6zsuTbXlpDZpNB7uI9NpDV5e0SNnlKdTh3LItAJbcKCvgq7ECHKV2LAzO
n0iPJ0H1FWpOm7/QTz1OsnBmkR3i8EjaFqYtjWzY7SIFf/cd3U7J9rME3B/kWkn4k8F5pv6blV7H
Y0tiaNpD5Zp7SbND4xIf6D5y+SoqAYkOQz2QKrxYn0crS9S+aXQjeialfMfPGsRSzegcJbkqv3t3
rrIL6QTUtprkEgnesuO4ECjEpTF5AIpjJNlWpve0QJyh214L/1s/s02fdY1lq3K8d0g3tlQqnZFe
DVOH3HZ5fH1onN7uq3pumJHJMWeXwIAprepcN2J7Rw71Mikm/lxt7P+8eajU8nC5fSqinxTSNv5r
wUPlmxT0jmyOOMaUC2t4Y4dvzz1DSFEILG+m72kos2ozP/EwHs5hWiDr/abAnpzu8OlYF1nl2SMg
foCyfIT8XH+T8rMGJ+njAuJCFb+3X4oh27Ji1SVgflBu/0yqMmW0JmrDHD2E+drcRo2IM+0ZXdn/
x6C1IhPL5d9BZjZTCXT1j6LT/RO3/PVgOcz/FjPXxlK5u10fSZdq7+pK7b6D+riR0t35ZT7wcQc0
Uu6QPCqZ41ynlVOCKSRQUgNzkgXerqy5yUgS6QV2jeI2SYmeZHBZ1Pm1shVHtTRiNgwpJrTfFxMC
GjnAm+12lidl3Vfk9gJ+IQXLF9QQLZmJHjKHKWCD3QI4S4ZDsoSIPu9TlXVS1Z0xv26MLlH+qKcT
IxXgQ6RRG6EMhF2bdq9KCw0xSrGn7ejVAY2tY0gcMvN+BkePlMR0NMW7tpk0d9xnGKkNlDwF4zK/
MjNrZL0TF+V61AhaVRxsop0fFvk8bceLxNZO6VW2Ps6ShVsQw8fUcys5nZTbjoMVouQhP4E9iz7C
rK+jU5Cs6tntzcXKLoPI93XJFcKGpf6/OpWm4uwDvUrn+W+Nr6YjHNONNGL7hYH3UN1VcmteeN0l
QqJeDvi8XA5tNbXlLY+8IJHBA8hW1uIoEZvPp7kAeRikFA4kIuGgzFtMmra3o0go/dcK+8hKys0Z
+f9PAGitOoOAGGIuJy92e2QxPdRSR9h7eT2y8Gybdb8/dkqiuhPbDStb0VUQ3weod+kQY1U/wWz0
Pnsx/Mt+TKfyXAQ/LbNMy5vhg+7MoYuprD7CEcV9KrUuHf7Nf/XCFAmQByTYI51NZZtsSXdU8xh4
rJQXbF1jbT63bVkZPe0s1gQ9FLubzA2wml45gMejxgYL6y/k0xVdV701eCJkqufuuXiwezHukmwp
fQOCrSCKGfAAz3PYcW+hp2BVzbjkH3sx41252lS7DFsLm1+v4jRro64c32WsJ1C4Yx3UDz1jUAyR
PDmSTyXlxf+DT5MfEhLuPwj8V04OAOIfe5KKSlG2iSHSxFs8H+T1Cgm9aSZCWPx79ZTnBvkcUFtY
k4QJU52ZJt/2V9u2i/13ySNDz+uiHic99pq474RJ70WfMfrMAHMOmrwKrAcbdqFgdoefaIefpl2A
leFW1rYfRK0zSVyP7RuEAahPyi7arxrFP7mqHTymrWOF9LZ0svK52qwiB7fXS1ck1yla4LQXiVao
PJkl8JZ0FHvoqJyLwAeKiG3KmbeTryMXsTxKRAxz/sxu5w+XeSPb7mAzgU+zFyZg+aLQ5IXzqxc3
KCE7FIX1lE3IqH5vDjXuO/kOi3BVVWBdeveZ8evp+aMSnaU0rRISHQmRvoeysCoMEhBElz/cK1K8
coXO+lEXP+OVrS3CG7/fIQigeKlHDHXc56tFQRT3ZBhToprahppL/IertKiQa7oIwz2x24jiDJY9
TmdnD12uqGxruBXEGUYagd2d9hifLnv7U0jrR+/Xlu5La4GyfaPfAVOTAA8dTxCfRGz8NjPwfaz/
NSXoOQ+ZZo6hPMiEfgXNXSKiF0d3JaMbnF0RFp3ONg224/D0UZHaf/97dgqUfeAVL5NxpvJT2XLU
t5PBDpIA8NM7oe3AUiU8qZ0+TeAZzuqAV8VEWP7+qf7J0qdaGzOWLtGo4OJfzYqmCwO46fb2ctqd
dT7m15k7JK7C1Gk6Nv+EmYlD9k+YxBZphCMKl/dE5dfyg1XkGbMqJB8YTJrcF4lvtR4lVlfoLney
8PJwvA0SON2u5H3XtECwiEMs7cTLp456KdnQFsXRi5fcvafDkNBkwHdlaTTEMp33wbRm4cWpVcUf
83qBbSbPgL2/+k3vy2VNIDR7PFBCgu6kKJPdNg6t4z0CN3LdwFvuF1DzX/uQpK4628mLbF00eiVZ
gPZSVBjCDiuK1KAuufMMfcnUzAr0lKMGIio95PHynqUJRck8kNwNGU5w0azl8fwBGWwEYz+5fCZF
KoMVHWlOIg0XbxZ+iaBhfaZAwhQxsZqjZjJmzLkWy3vNzFeXvkMHN+zvmZZW5LKjjc8QwUNp1KIJ
vEbcUNHwZk7RTnkIWcfq2bG+i8gd/92iqyh8dKkmD51kmoTqW37UKeXm0GRymaul3a9v8/KRUkdj
Y0Hsy0C5hgXIRYs/rpIalMTSe+0SBpXm5mU9T4ybuPYFc35m+CkMVY/AVD2pdNg3BWs5vMW7jsVz
XOL7rLTi0i2Th+Qv6XExSo6v/zrHy//ss82e7o6Xvz5A7YLqk9qscG+EZpE/43aYw1jvNqkrhFT0
BJNO5Q7apY9IvEjFbo8vbqBDYioig7SH2HGd4NEciS7ln1suC4GOjYA8t8aax/jSXxzWbrH0hTOE
JehO/R0iBJveXg+Bqn8eXpyzqoWt4Q8evUSrfsczgOG5neqf2tD78KrQ5L2FkFi8QbWKGK3S0Dv7
c/jBl8NGw3wOXhLIPKg19ytGdA6YXI9qGGq3iQIgZVpZuwmq25v5pO14M++cVFEKMKN4GHbzen+r
RHurDC96K2g/cE/ccYVj4I6dMHAteFoOpIFf6aZ/U7nU2741j8gxIsoJDR2rNDm/C6DWUpUX+HSL
suDS1/I3y2hvtgFKzGF7nZYgOFTDRqWsGo+ReERpJ3/+3GZw/+C9C2J432LiKTLvdlDUGxvk+ZaE
mT0PScxg9ZuIZ3aXRhPova8CFLAKz2YbLhwDPpJc2mcrqHRW6eCLLr+TCJeDslkezmpOU7Ir55US
wsJZzlonrCWuCAW8cRoSQKeE2N58JVvD2uocqmslYyUoBzoKe96EgM+yeYy+QTPSUo0IBIbCtw+U
TvXgfj3PYcOh73rW0tLpunYMzQbvLaWvB5+kRtWUBP2UCPrYfedvfCAAw7QrneO4v8sMzNtq2lFY
OnfnaGQeqDk+H6sshaGweDtLj0mkVUrEDJ+ZmAush0UnIkJvfk9K8OXGg+8oP7IkcX+ThurrMBXU
AxdmlWavnQyFO1dKaBIAjtC89BZpo9Ep+/89Y1wtJpX7nlZjVq/orYc4F/xegLnhrqyf2TXA/x35
n0am/vhujA0FJAz8Pon1LGv8DxzVi2ftzqbrHumV4WJ3blYn8YmfrKAkkofIdP9BsJcCUZxGz/mY
w05uPVGk1xZkfHG/+uq69o+1ojyCRisEcoexEukl1BG1OFRrhNp/gZykwO7LxTgcp0mW2t1tkr9r
uQYVtA6P3u03S5xQh04Q0scL0ipz3cQxxeUSsic+SBLmbwuJdKZaNejf95PzLgd5YqlpN+aUJDNs
z9dkHVwPbJyKefwaUxREN8M6oZps04n0kLOyNHVnG7cf3XZo16IRxrfSvb55agzK8gC8rKK3qrq3
UBnx9NjrP1JV6+iYdmQt/n/Ge6FjC2D7eP3cSHKpWJWlnW/lkPdkoeab5cLiA4gdd6Jb9tIiYxVo
x4g4sjGYmAfNNJWRxHqiceH6brlyw1/L6PdbH+Tg3gWDycYutlzVyUmr1uueun1lfIZ2Vi9cdWDd
sRK+hdcjhQccusx8FAnE7U6vclcfOV24RmaJHKCevIdsZzosrw7iTyjxAkj+sof/fZDJ5afmt6D/
jwws2+emvJbYyu651WWdO10t07YElrF/jMWMnRZ8soUxVu2xt6Y+CRx1w/+d7L9Gz3rJssFo2Y4F
3frCDcKeuvOR2MwT6FlNXiNFo3GmEZ3IvhpA3wPu5TYER0lJEil0fQl4kZf+qq+bKbjZKSysgq81
OIuWr3mVoCrQtzGa6//294XT2cCJk8OtoXB+2nbDPvYzaAdX6RJO+0t2vsW/NsC2/qpeUJCJXGyg
etgBJjqWZLblkmEVpRNylswzRy62vqPkGAVcVQvuTTdXJX7xL3oQEj9Ut9OeAWe8gEynr3hMaW0Y
TolDssQedWPn1uVlxFa2Arfe9+7cFy+NliZoSNQ4rxo95Dlm9fR7ZlivmLF3M2i29pNZ9+0mvEvc
utC2X0eec6crldFenVnwb+x7cyoPOMuDLiAc+DGTCfDbFeOrynB9DBxw6KgFtaharrAwxzlp56c0
VlR0NMHJA2vkW9AgdFR32Ddls4fmrLBjW7jZyM2uBNwz/aiGLhHt8KrylyyFbk7RthfO0sOo3Sh0
7b/MZYnyInrrzV9z+tVk2j6PTke2pc75DUzTAykKqy/zu4Ey4GVblxEgj0yARvX7YC85hXfXnJma
m0U0AMkjIB/oZrZMoGxEYxkeP2OoT6cLJtLcicbiH7n4YQoZh81oTQrkp25BRCoyRiJIqyT058Y+
ZT17WlPgmVU6UQT9NbXHglm35GrQYfo/N0DCc/vI43EKVmInCaHnzrR7h9k/p38nbckb2HmkoF/w
0soOG7NOwq1fFqXTguCe8ioDh/3gnVHFZHvBzc+yC0q7BxH2kgk6mVGjBgc3jBmNEJikpCm7d11h
BHz3yFawDXbEoxCeRTdZRQxAXqO3+EYKFCLRjGzgYKArwAxKw+k20E8Y+hfIen8HUkN0Muv/Sx0V
fwYqYLBGq60aMGmCCDWOkfT67k1ttNofaUb8x1LlUM4+sPEOKAXuDQYvDmpxUWuIAAhdaeT2kT6F
EWgZOwUNL+W2U08rJwu2K5SouUflqp9X6vyl2O6jiLZgzjEEHQd5PyclqCxb1u8dCczKtAh8iIWZ
PuhRG/Z8LkLw5c5zulx+DZ5Jy+02bp7l3N/5VGzWURRq0iZHifzPX0paBERZLdaGkwPzaNEPvlYN
PNcHoPp6x/hyUdDp08LA8Zqx5WFXFcX5AEMXZdMoyfB18bMVNkItf1kdmGJBtNGJYfV1qTDXvomb
ADezmj+KHpdYUm3Inhq+CAZM1WptFtgIh2f5SeXWO61dN0g9froR4xYhjERpqLEnrysPAnZugYMT
GAt5bU3875hL4V6FlWblDhXT0mKp+82cnct4hnlMXWmQOkkVceZww0yREAs7iUGSCuriH0q0GRwC
YnoowvI0ULFTkiU9BDjsj1WXavc4Kb5dVOIVqe+uF3xPzv8mTJxqNUHw4EzIngLi/eturfwrmuR/
57yiCvZVMsdOojMfzwgd9S9tfkNG6PQXJhTWVA6dye0B5Q7GcQchy4iQuCNJZGxHbs4dN1KzoHlI
ssa/tBIU4ImVgoYdBlyqVVGKbvt14Vy+ik1zg613b5z6KQB19j/x+AjeyicM1x7GmfYy7VK5FEXX
JUE6+iG4TF4XIDZQEpDota1A8p+v4M9AXA3Ti4iFttDZFoY1dStghdm1RpKMRCXrcodqwUADlKxR
rDONjbQ6Li5GcK9LjVXQs0C5X4kMMu2aETndWKitlYXFu6+LhBighOLpyHuFEFR/aQqowThlBUtc
FIvoCqQDAss9ZeeeGC0mr+NwndyD6qDAgUovYBvrg/6RCcoxIyctHW8AdmIz9qNtvSOkOHZTudPv
sDi+1qXzvfLr1qGnWSoH0+M1ntLq1CexGVCgQmAiCwh1qkGfJcpl9ETPc0WxJkfnfaV+FFt14Hmt
GIqywTlqoicbYyGd8HV+QTMbqfltKaXDNUAyzcP1x/0wbTf7rJbj0ga+SwQmhKa8jfM3m5sBx28t
Nq9X3ALNYSfd+rKRzgLa/OsJCZeqD6+V0VeI5L/LOswCGjTFQTgSsutQNZ8GA6lz876YX78BWO8Z
fueizGrHZcHruu/v/eFJntSKbBZ+hoznOIzbjBqf3U+iCYJmmGYU5J2bbMCZhACZp35nDQXkkoBq
xOoMd5PLOyWHQa9Vt6XHBkuJZD4nei7jNwCwey5DIy3Mwuklr9v9EsJXml8AuWUhxxIMhgHk1lZA
IeLXTkcx0Yh07OVwNeSiT8r894EcAI8iP7Wrr5kdzsPlklz4rq3wF1gWjRSmHlID6soTCLpqGb+b
VkADzZHKEISkA3JDOgbot0P6D8/lekzYP6S5xde001QJ3R4ZU3QkpAeR0rXNjEBVqTbs92oQ9mRo
nFZ41pcAV77AqV+03mcmLRn+Pbbib/njRo59kXFTRvDfi8jZsahKKri/KQosvh+XbVBwUYJyRQ8C
yuZ8oPu7bT6H7bHQB3lEaJy8+WRM4zB2G83PzupwHcw0rASSyL73VgU5D7l43LgXhwO2CQBPqdU/
vbwdSHgrGop7NjMKsUBRf6VfKpEV1qd+y2ZkClf1dfToJ84B1l1mEPIro1dsR+sw8QUd2fmw7lWb
nzvfF7GJUfyY9wBYJKJWu+uQ4N87ceihroQFC8e/ZVw8RovvzrExWOhrk5tHZamb5GGVn7skUjxK
JybaT9P8UNZrnGc9WSewztHT2nRgTJL2jRACnokOs49qnyHG2gfoZo/nQ95FAx06Q15btCLfG0Kh
Pq59dvc5hmAvCuCTit5JjF5qGMwKOU3AnjJrSi9f4x81E9QTJkiojS3oSPtRLb0KAu2jwwQwygZP
Ukw0tEs31dF3CmqAKBuexq2+9u1xrI1/hlJhJnZsamS1MillsNvFc4nJxjc+jgxMIKRua8nmnIl4
Mvv06YNZ9tG4+EpbXYexET5X4N47Gwln8DJcpm+vffcX6ntW3T42IRv51Q9/bmVSw56rxcKMIgrg
vf82z9QpEBf8s0strp0Jlc9gVs4/0ogsBKdoOrgjRJL19VnBEmb3jXT9GoLxdFZI9fBGe1VElVFg
nqRsLIQjkFOvr+oSVVCFakYCWXR4iUIyCtLRskPNtBXkBgo35lPp5ErCQKtouNllkXEUkXfbLWNB
VEgSa5BflSUz+9Sm+bFhlq/5KWAImGotDibCBIZfH1kY7gx1hwRHYL7u+whkniIglTyqtBlz8kAu
cscHZkRQMSv+RMMWF12FofWZ9rgUn3VIVua69IHg0Hgk5wycamYN5KLWM8hE0T50szZNgCwCSp+a
2SkSDa17AGAOdf19sYnclv+fO5X1Fkgt5OFd9ZsWKuNWXdnWdqmeyeUde9NumiGSf0Cxy15J/9ph
4dE7r8G717qvFwkqToGj9VmF0NUXh6N2fqJm0H5IBbbbU31cRmc7h5blHm5tRAbqQ07X+yEEqk7v
uXxRr2d7M+E2i+ztFzXrHa8ZK8AkHv5CSWOBKjPU6a1DxLPhA+2E2J6MdwpF2oBrcZ3EZcf2pBWS
bIQJeQ5ny23qVQQUJapj/O7wz2PhUz79TSlqwGUrTA1BLwazLVnnGGS8LEuBDnmkXBhsO+ryFwqJ
8JZz41wcAlEXEj6aIwi0EsWfonDsf4evmR/pl46Kht97fAKG9Pl+d28/stjCdFvW2FWHM0fRXSS1
a8+Db+Gdk8Nv8B/eEDrIHBxAoy17YawYL+K3JUr/EgffGitXYOnoQEPxSpxG0kZ9bHqTQO9rASZX
Lqi2NU7ODjlmMLpnUSfkg2OsJagqNTeOJkiBFCruVdlaaqtJzwWt1qG3vdn1+HDZ1e8lnoxJW5Rd
TczdufYizGFCXUAYsiRNgiZC4aUwIU3tbGRip7mN5fUJyPrZUTH7+4frRowOI9V5DPD/tu4NB8yu
fztu5BH49A5B20V6dj81c73T9M/vx7ziQgn2S5VQKAR+CahD5Rl47jRSwoSAqSn/M8BnsgWCSgNP
2zkHsI+feJnnivuHEAf2LZWqmXqfSc/iDOgXqRs4lcwr1JNSTjDPmL9taiYoEApaLdIy+dQkGZmx
yoiTxSAnAUDzlbeHUu/Dz6+a1xLukJcTSWKqRd4hYQuC9yfkqvPIlP5YPcQ81KcMNH6jNT3Bm3Zb
f27RhlVRKMacOUNke+XT2w9F64jBM60ew39g66vmYUC+x/hj6xJiFf0xG5bivTngDW0n/xa8l9xj
kNKY8E6wDnGPPcR3J45rn7fNBIq3ThKMVB2MeIfLsF54s0CfDCDnk3VY5m81MdbQ0Nvm7XfEGGJt
Pe2BXzRZyBfuY8aehsXCC2Q8Qm1+dTlPOpThU2fWTTsu4Yd6+WZSwSZeDLrSqHeW8X+EO3Jg3wOg
347bCPXUaak1MLGuJg+UhX0B0sl84JaTahAWxijU0eqqBQoAVFaXYYop47ylkQwlmy7IU97RMMAW
dsNVgSLW2WcPMWBjDTgsxsLhvME5pMV2vHTkJ8r/BSAm8VUW9N3s3femANbiMAXBSmEZuBHeLrJ9
4n4EinAI30hlDu5nFIopqcJ9ZxrwDqB/NswOExH+HJ414F2+CXle7Yeb6PgH6UGHTddhg1OJsMZh
cTg50m02BY6MF+vyi2MBGzt4HbqDuQ6ziTL7S/23+My53WeuWGbp2icB39qe8u9XykLKqky1BGSP
/oXg2hQ9ZR4b3kOg9ZB0IbgkFZnJ5j4+4zCPC0ncGmhoauBvteFAepQlTDodzmb0zzJZi8ERedUE
Ij5HCsFs+NfDt6ha4168Ysd4JfxP6m9OnyyRPmJSeG/niHY+5TKaM4CZ4syy0EdDe6DW5joaBlso
CUdk2JwG/JW5gJBzjn01TV89/qrJv3/yLBhDLrvQM2diDE/PDuAex966dnRipsopzQyo1AguU2Dr
XEpMn1K2VKJqBEJMqxvYMxR/raXvuoqXsfj3ay6Tc1jPKMlRC/tPFT+EJAiTvd4S44cHyu7lFggb
ehnZ2EkV215itLXSg7xGqtQfcCf+O9tVw57goHp8YHK2ktZ3t69T9P2ff7iOmjSWp/ImzqWdoYwr
JwHyR1LV9HjNeAxl1O5uJ9SEj1nTnmSt6JFg4g+A7pe9QN8PTOMkq4HPK+0BBYm9RwOZrrKLf1si
HZxI/RUXZbNJ23Y6FUaw68z0kKdMxXqQQwBAVemD6PW+D1MyqiI48Lo7Ue1i3xw7G5CpU7j2MG7f
uN6F08xUU6PyyDQP9IL2jv9Kvpr1XVy3ck9Hz4BaCQTUZfbLiz180OaoEJNTnGqRZx1vNfVHLLdz
UyQ9ovZXf4TXJs3LZq/BIdD1JYCNm5sEw9PTI1vkLL0ME1Y8bY2VEfkqBJ9FiuxkFQxDxKXYqvLV
Ju9YpD2oO6pzHoJg3UEl8G7za9YF+rsQlmeTnXnTkxxN9fPJglXDj/hX4LdQYHUi9YFF9PIaTUxa
/Ue+AIOm1YddMIDTGKJZsG/b55+VpTQGlrezdTGODdxkfXoRAB5fHX1zuYCvutZwEqt+W52IC0Il
9P6b9YFB0WP/zLAzIcpdrCRPfjV2xlLi9x5UBmXLfBnd+7xUhYX+Zr48Zr5xbNlxysY9KBpN2ELQ
B4Cojg3w1LDYoeuqAueSWGPA5mcaUBOn/aHKf7g2bOs2k8c56anz47rZ0sqq+bfhj0HZvyOJOLAE
yTTSrTAFaEKPZwg+rcV9EPnuTVJaBX4cGtltNcd6Wn02aHAxlSquAmT0JUYyz7Xer01fRzWjkrSd
dpUEQ7JsjvETAMIXCqbKL8Qkt56NzgXqM50ijatZAsD/IP7TMLjJQfdIaccuO/FswSE7YZtOmPNO
KFc7m7VPRLxYdl4G4msIC6jTT5TqDVQqXtGwo//UThDK0FOw66VmaTpsoTv3h+F8sdOnPb6hPZa1
yDGJri1t/AtEPZR8lPtLjzVPh9jqL8AX/jJG1FZacM1uJ6I7uM32e3yneWLOMPWqhMsN0EJEb/U5
H9xQilwHVlDjBNMM/hGtWvsBu29U+vtXrUMYJn2An0tZ2sIMEVwSVZ8o4FIpiQVib59YJHl5NhDO
VZJZwXFw6HMKl1+EDH62YhNce+a2yQN4T/+t3+5l25bfEtDqXaX6D9LrixvvAygmktWDoFFSBJM8
Y3ipVhRZOp7ByeFZt698b3+WyWoYg13MTxvG/TPvHng+esNSY6bqv0lg+V0ca0Zhxw7a6f5Ad75n
Fvg6SrrB4ogdf2eQshl6fIYUH1f+Z+YIxhN4+zM/CdRHQx41fMp8CK28/UHGMwMUxL7TcslNqQFX
IIYms4NTsIkZkE2gtHX56iGySiZ3pm7qLteBPQM185QxuddF/XeRSs4DdbwHyqSVnC3ZAqqIZE1T
PfoFRjLiD4vtl0U6niTdWvelFwoT3ATpOsrGvWJZhOqs3dFHWJU6jkNPoFrXPMrl1kHI4er/vk+N
L/3CboBIEZ5OAZGRxKsGVXUEPHiwzJI7ngV+LEbTiNXNqSHgtIUAg/SJ1DNkA4SWGF+JtuIvwwNS
8qQ4ZWDbWpjFXg9vP9n7mPIBuPFfH58Mcv4lUUK3YAPr6x0lxo/Vhk/NjPXyDGUskh2TY4FBu8DP
6GQJT/G4bOzMNu3YCUZi9Sggdpd3Bh1cKYzxD4IWayWHbaz7alFwuqZNBsdXEyoFh520MqOZyJVf
oPf/0PG+biGV85/1frCJsgJyHzn0iYejJGSngwP6iePsa366P0qHMwOi5BHrlbrCOQttN0KqJ8Sp
Sj/DwmQ5sHNMtPrM2YokPXfN/uj600LLEAkVmNzsIr34M5PMOKNIhoa4p8RrNQWxkavSr0sh/5F7
BCWla69vy8Aj8igwFiOanlPDRbjZZYsa1Nmwx1NyhRMB6wqsiAUuNRnmYumwR6I/QuktC6z8Q+z0
6pnttOS0dTQEH82quDLNX46XPq9zb5CetlTJmo6beyilYEbTfUmbL6ePPnAL8wuuSd8m6lY9xGq6
QIIsq7t2vxJBfSnR7hHUc6cb5xylutNVWyg40m5mZSJIhPlM4VcAOusO5UJp1DA7gs99rkydpQfY
O9ABm5ZlvTtnTZUKAlc1A+fTKsmV3+K6qyZZIyi1kfYuJB4KM73tjwUGzO6guibr099QQNpn8XA/
8r2k6RMJWKDvijDjv5PlCjghHq677Or5wTbtLuTOGe/7nrxItQSoGjK3DBXY+Gelix9AVGRMcMKl
f4ChDLhbswO+n19+QJ32BDyvnnO/tWVbqC49CvPpbqVrZc9H3zEek1tPjJLakXGA8uk9cHnYzIPa
+tGTvhCvbaHOzOHE8Mai2RMx9Ptpxq/7Fqn+IGOxHL2e3YqTAOs7YUFJw5NAJa2YsHQ6GiAsPCW6
Drwmid1BuHmYYVwQE1KvX7LwPzU8MJEHCuXWIb6Xs4lexbnFehi+kKqHjXu8dnRmP82SRCwy4kse
9lpCAWrMhbgwE6Sbt1CpoEHtzQUlGp+lOeIM1U8AWNj949kYZyP5pKQh90lpBVT66woQgC7O9ioB
c2Cgsm4qwYOxKPp0Qw1LX9RDN1NOKp//pllUBndHXxbKqeuKSQsdY9ZnoshBMuQClSQy96Yhc6cz
XiQYIIPkF2aqJ7VUOyTjNGqpj1vH7Ih8WDdvsTY6E9CcGRTVxJXgVlDxz9P9TDgTykZolU9a8l3N
UyWzobURKpwFSN8thHbqlAyetdlZHafNRCaEgChpWl7vhIUQ04ET6biGwurjMKav+icSwvnD2Oi6
2Dyg3GoAGQIYUASZtYJVHyK7US/IGRfyCDgkQjwjTutRgWVRlq2Tw6IkxEWlaZvFhC2nLUxXecEc
1QOnZx0kXA9ExVLC10NyrpnRgGZnpMf0Wg+a5989mJqhxQ5LaC3MkvRQ6SeGa3JT6okPaXPDDrok
FrCKuNPhDMmcdYihgPMEcTiafHFfm7Umoq/y4nCDX32YBKUcLNv4iss1OSNCY2FAi/uaIn4nbR+j
ulkUiU+gvZ8dwHp9phUhVzuFcjyq9ypIjMhkKSslYq+eF+EEdtylCitAwoKn6DRNjy0ZzsOm7tA3
KGkD0l+cbTtp79x8yAEauR5YV2jRDcxl2swzThu5SLFDTgKnttLdBHcl3krey01T3vNpKwCR3xaI
C6kNinGt4/giHuXvJEw2yCGWYp67MkLjX+S4dsZwKiGZLsKrIn3ToBGssTBKSTn9O9ykj+MQdVtG
o4cDeEg40uNyvEYibWKWpsR7U1AZORgUNan8h3UO1KGfjUp43KfeiEcJRJpKFA0hfoEUNocTLaGS
CaUIhv0fjKTpHPgc4DOyqDlATxfymxCQArrIU+TYCXq9Y9x7WVe9UivRD+T1M40Jf9xZyQuICU7f
opMU/3C4gmztqb5i58WoyQJymK1I/6zJJoUz5d0/rzA6AalM8pv4MpWt2+J8NmZ54XTQPOu5GbRX
EVAWeh+7JY4phjncRWja4mOlcR2tz66LB2Hi/E0TCh6nYzAT6TEQYA8KFbV3sk8Mgta2/EewKSWS
9G6OwC+mdgH0m+GvoRh2CtEmuDNQ0+a+AHojowad/NhQuw7j53oZvLq457Kwj0PfBIXs0r5NSyAy
Ppfyb5LIz3RhyKKnHkjSLc3kAkkXE62hXY4JfRug0QqgqLhpGxBLKVNmnfyFFwdh/RzLtOQy2Hlq
QP+sVwfwStU1sjVtphyJq9Mn2h3LJvYy2ECEefn3OpPT/VZ934aw6O6gc4uKob+so9FOcCRZsu6/
v8+cVUyWo4Z3pHUzf1GtfjLlzH7RVo9y8dHZn/SaUDP5lKBjJAlmWqtBC6y4ZPQg6aqwagdWpJiV
HPv0EUjenj50qkcroOu6QbumfaiaYZWB/kSirJEkNOo2dCpbhclvUwW94N1ynNMA5zOLRakZ7dm1
h9CYEO1YiqgzjePwWkhnepojsr4W3lQpivzSQsiwP9a1Iz3oBfFtv+4NshZqbeHpinz7G64MzWKk
OUinMl+elrxG1ULMEqERt9zUwuts+OWP8XagQXIIqpI3SEBq8YF3Fw3svSEqSZAT/XIm2LiaGE9Z
x3pl9c3x06CIWL2r1J6vk9fePRcDnWXVDhjAT+LE2sQM15BpQipbZSkgh/lGl91/0L3oYLrmcrfm
eQa2q+Q+unsJaiouZ2O/pva69CdHRbGZvroprgDkXyJW2Ww5YRxHE9jPiRSmCvNiWdcarWpqxVJT
6LBd4Swbd/6xda8PPYMuxbDTmduDnMG/n72bYrlNqpuDjQW1ZdK/6vI9DbMmRtpuiLURvsTJxYix
zFPo+QGvS3UNRZQrlnNaKdZ7/HzqjjTpoog9IG51a6FHl5Ff6Jk1JJdaVHAcNltYVIT4OBK34ANi
Wf3GaKL6ybEyyZzLrqjeR07j1AtGdDtCs+yFcDAmEKwmvOBA4wvSjCRSjIid1AWa2K0/n6vinE1Z
CBuHn0DsIZBKw4fL/zHyzZjt4F7sXacIotCGc/opaizBa499Xc6XZZKS4AaHYurg8nmfbuF/izS6
4iDu0Xnqna8+4rhKNCFbjbmtGCjeYFgkJUrbaId7MqSGcAgyxdJFHsqnvqWo5hIMmOzDDcjkJ1nT
8+skReDAyyNbDgOCovlqLkuoKUB8UH8rTnFmxIUQBLFVFHDu+fyXPRNJrdONUhK5i+QLDWLe3bfK
f9ldShoU5YfRKm4Y7qNBsDE9p5tg8fzBHMle2y5XOkpqpZkxKx0f+Te18gllHch4122p8AJ/9Tuh
a6hogW/hIyFjwxo2oZrmac2QG4gfESzkp0WcNED9FiSd3SNPQoi2RnhGwQ437qcs38AKGyWFnVcC
qN2oxGxOTY3oym2qNIR3FZSSccUv3oc5Od0E9geFXCnWP+NOlMvAjzkwOHSjMGCFx7r3OWQXXR62
1VZNnDC7tZSo5wxWOpC96f4MBf1o21aQ1H6cLsYa03ivjr37fRUWbg92BCJmm4Q7DLyNt4oIQ9QM
xe9ZRodillmzn+GT01Ks0kkuCchnUx+FfbEJH5hLqc3UAmOs8Y+TmqBgwjzoZfFOpZkN2tyQIVIu
a/QDqLGy4kkB/zx24Ke3tjgN4OJcNTfItylfcyJgageY2rrm0Y+JRz8fVjr3wpr+1Q+0cpYfuMpa
0JlYWxlQesgWOh2Ln8GvL3rgY9AAXgfr1Vp0LWIkGlWOag9yUYFiBXkLkUQazoy3xmNbaYc96+Jt
8uEXG4cTMD4NUBFT//oU13hMTLsQijz2qzwBVd3Avu/M6AfW87V7U7FmYwkpHeDbXFfxvz4VGJEM
rFpta/yBB5krDsDXm4jEcg6Hy7sJf7XnIEnXR426A42enaQUDek24mC79hyPSiZzam0sy5Oimrsw
yR+1FlSLjkOwrzKb4+pJdzAE4prM3FEmnw3lfnM8dkRJfMC3cYum91OmFsJk2JIVH+A5f6ZDhOyp
c6IpTkdCXeBmW26bPqB6H+1LBPG5VUa1f4OoCGSYzVzCpl9YDCLu7rXw2T0CQVnZdLC+6uvnWen5
2Pz9cgwsx1di8UbajzWupwPvPHEeAy5AzAHSmUoxnv7kKaYD5YI2nbI+t1bHt+fGgOX14vPPf/no
2lXcxHfjUYOeALtqrukxVtUDS9u4THk3N9fbqXp7xzLtpusE4zqJqo8is+A49RbHsOiRhKozQlZB
PRuVcWtCOIilJpexK+1eR3JoM0oT6lGqwq7c5hXT9dghNsD/Amx5akBB1p350yv251HhfkFvp5JR
1F48LzydJZ7oXNFvYQLZT2eI/Gnwz/rbtrTARbb5xLJdrXMH2a1moK/wmOBh3rKw2cSKKF8eJ0OR
kGKpC5BnHo2YD6gYs1Y7CVHBjXGGDJq/L7D2ZuJlEkIPA0sQ9cW7HXL7pqDWjxOjnumh1P0naHB2
zeQMWoIx7ncekEjOH7myn7q0V3/sIsZSJ4NelYiEibUaH0yjud8MD5BZhdOnm/mg7qivS1qGGCbc
vGKV7/ctWgjELZM7NWrxkXQVTyRyCy1ewWFW2z75rMUIu0Gz/ty7ke2QpIpW6CdBhBVPeqhIO9LO
1NLCbiRxD1iioLTBZb1Avup973dSsu1foqIwrEmnYQRkwxk76te8SIqJkmigHIU4UgM81Ek6eVNL
5oKdOufDhBxzfdz8d6s/k1BtfFyv9m4TrZsNJwbK0wainsvUrDnjVB8MKYcwC6JmrDN8OGXYjIRB
AHyRFtIV7VtGRfqrnqna42wlY8TSxw10ePY+UwHAIK3Mvmq4r425yZtpoJw+YBbihNQ4VRCNVGLl
e275eJG0rjfGzewEY1iWD0JnoVs3OwmIZfq6UK37+NC2O+7rsLUi+lz+BVLZN5tpHaiVztUpxY06
91lcYXrNWskYdepplrcx/FgVDUxFDmHfNjxdKTdZZCz4HlaDu4w6FaE04uZFt7OIm0I7B17JuFYB
hODA50Y7bxUOUFufHY1bs4N+Fk6W9BEXSWoUnSOznrrTNHfRcjmb/+V04B4jEhVjCNQA+Qdogljw
kCBRjPAV8lzs9FTo8rZw/hIRiPuaJ9ADKMbaNkpFU1hLgV9OBjf3ArDbf7NEeuee6rYGBfDNyepF
IQuJHtNMcwRADcjwEptSBwoJGPVGD+imuIFYAgc2EueHPt6KN2wUJ8EX5dvCfL5bfTL9tMOkcK1M
diHysMvHMzknRxL8/VGdl+AFIjMBI01Xe0k5Hrqc5OSNHTIeRn2uJnuoEzyRsksFa43dFfEnHPPZ
NYvl9sGjEoo2Qz7q+bhy5SkD/dkPrqtRkt3P763v6DzfUtY1gHZOSPSqWWeJWqeYucon2/PYoF1d
0++X1XwwYTSYuWtLYT19uEAOeHoF3r9tHYW+sz7qlKSisBSXu37hqu/eQreudk9fCOU0kM/wRGJN
vc0NTcFnmMGUV4NvQeoGrNXEel+yaS/AH19LlFJIBM/e00eTh+Bgzral8s9JiNVAAELVjmfb/RT2
F+Fci4kEUM5PpQWoArioA9d8CUMRnv/e3Qnj/FhjeNPhTuUwwSe+aBghh4mVeGJ9Jb4QzD0VSVFO
+USrD2ZrMVsZoidqAf7WrHGK1kCqz+uLRFqAglyT5C8r8T/zaIYRVLAkASEj0Y+V1zPloDThdNvm
mYtJ4/XyWz/K5Z15cHPrxEaIFf4DPn2CzSodw1724F9zTDICwMyK6WUmME+OVPgXqqvGWWC7NSfp
9jatpSZKfCfMoOU3T4SqqZe1nd77bEqsZ7nv6wG1iJUWPWTkACg/K0dlEvbtdFIQ8iFN+DLtLuAB
KROV2Gk1Ck0sa3PV/fVp+Bn0PO34Zc3CoNy0buTXlEW0Ja8BW3mUktZkA4HSJLIPKtoJB0NJusj8
OeIMy8chXnRzYd56mroz+WBxV9lHLi5g/90fvKRGIWOYZWTtS2uhAPvO/DyFra/z4iwx0UbI/Hzf
q3AzONGlPMoIDP21vAae19CGKO9xqYUgHY3wsX3U8q4ThclnUQM6rqlpNM67ivoXPFLpV+OHjS1i
pOWSasqqulQkRYa1obABl6q4k9FKIdYJH3rUiohAypEJMWFJhp9+I55aqoONPGZVMDV+SWPqRjur
P9LoSywG0dukYYUKKJi7swEbWAW0jgJFm7PGuHxf/lkuHcKeeDNCGlNiD4BiguALRkRY7sqC8UAX
a7FVZzxDjm3j77db3UIfH2l8wy0e5FzGgJr4wUA7TZKjuHySxXMdYTsQ9ILBB/wBwwkKhdESC5IJ
CZ9cV2mGq+lS2FxLMKGBNMM42MQIBGQkCSs6kTLkNF2sozginuK8AiLMBqkrbWKi3gvjTMl7ppNr
tEEhZ8w6NfGmTzjD+FdLvLFoaCHhtsoAizaKAhCLH/MirBI1TyC+asT+bdT6DJ36Co8JTSjKX28H
alZ/eyuKNYUTZDa2iaFIuZB1r5pd6renrBnLmcfw6+U+8sWO6FNUNLK5nRnavE8pm4AaEUHWLm+8
ZuZEc4bOuGDcsi05j7LE5woxB6W3tYf6ufglb9zTD/YUDtyeyF0b8W8Tomez3bGOX1YFbG7UuR9F
NAHTU1FY3zIkkX5g31UEzIUVpd3nqq4VH017G3dz7wIaA7gG88+LNN7K171MgpdAdKWRNhGtVMaa
ELsdgCN7DoHBEthpXNg8xdCHJPPVijveDdH+s1ac9ZZIChSnKd8ZahfoM7sGxO9anb0J4iiY6XC7
1yuMzA3tlmEuwbQfy4LUzUc5vynWaRCaDgwuVe2FauBbkbkUoV+xkxwTT/Q59mqDWE/o4j7XhYQZ
k8FZ1p0FmglGCZe27s5INmJslaaxkVyn4nTTloTCUnzhSX8BVYYnhGhMmpvEVrFED8a3Kxm5zyQg
f3jOMbjCzVTrsaR4YhxZxYCBKVMjT2XS4jBm3S2R9fZJEaSAxUT3d17XL8JGWJ5mzAmlMClH0/b3
ZgE7j6d0DCoWj6c0SaGVm3TyWdR3qdSBDRCqq+CxjKtr0E1JXmBMrpfr8RjwsAHEMjOfTZqsg1AU
jPj5GqX3sTT/aj5so4k/yqJAFQUR4pBBJONEawM9lFQ1Bsnqz9rESFKvpT1OiaNLl+HDbxDayB5I
I08f/6NXywGaUPbnoyLY4WOELZmTlzc8sz320N0cQsM1T0lODIasWHJ5eNe1bAvUxiq5UhTNvoyC
sYjoZOoswIHnCbMwCOa02qqk06VB7saceB0Z1Vnq8cZTGoJtI8/3SEmlrmyM/robo8oPaVMdbrtW
LQWTLsEliJqZ9pn5IpjsKBLe5m0zMg/pUzq42Enbl24PSr81zQpwHzUw4FMFzVWBLjBZQ2L2eKYs
yUsqJdDXSfDeFm6j17iaLmQWA3GxonXBFApLIj+5+MOwmX03urvD4Ax+UEu9s4DWQnjSn49IEJ1t
3no95jgJI+POzsXAQKgCjmSw3KtZOLPEjJfsJWwj/fEd6fbr3SWjf/cxfa30iTla2/AZyxhuKlh0
nKZ2NGDnU2nx3tYfmgW92vpCMCDkq1wUVYCN8LM6rMdXOHQ9GOXvVY7u0nLNmAXimrzQ5wow6KXA
V6GAuLaxO2G0WF6QhPIcCz+IDyD+1hNEWe7Nz//C79lFDSp/sho0rKv0jpEEmZHBC1MfGWFuTugO
9HX/t07S9/MNmdYiC2dSrJ6mUrJSMfXnSGhM8OUZSLE7VZqnpVx510kbP2lEXL+flpgWyHUOWs9b
kw07IuWxogvHB6lqD+FtFmBQVQGf+YLDIuA/XkJbwD3hwdHo1vHEtUzuchmWx03EKHZvlIip1ibv
X87vGt16ELc1JEb0JVWnrw+XN+LE3JGV2od5WQMhIxtFXE6Q4XNyJmO9ac6MTcp+qDdH1GmXn2oj
DWsQeWCg8R4b/Gwm5qpfATBXE4ZORw1rfwCXIVAbjMC9SY+lFqv2cD3ierwuxItAUwpxmIwMj79H
9XdmdLmh/jXnPt+q5KYqf/AicfufgbEb2ejcVR96nWRyJIzlmPpsBNBHh/t7OBbtx8LiIJYFj7/u
IXed7P/zrnXwt6UhTX+c+5DYGgFG4Q/ph2iy43W8PaKLTCDUfO9cai8FrqPea2fDaJXmfJWswNVT
fgxSYy4PP8T5GJCGNUNrJRHW3AoE4iqImX57up69BQPvUzeCTJ7Ubp+pv4SVan7rcIHOxb6nzDRa
oI6UTFNy6RgKR9thIGOkfX1y2dVyZV1vhQpaKpCAC4DP9/htDdbcTj1bIW4B025x8UXv5SipYmg4
tgW0+zENgb08YJaW+ob9xygo+eVY4e9w4TSt7nAOhwkZ0CTsY5XrI/pM0lElir5yEMIiQNNfUkql
5jw5od6nlKiKEO+OTjrJhaXZqwRMWNPIiefccbPAUimiC3LoGzoFiR0ukU9Oh0dGPMVDQankSnAw
bFisAy5OYPogddndw8ZocmdOSP7sBQaRaTTJOF/tysOJr/1e93uW/44BZ6N2dc1tGFwQvZSHcU0W
qrBXbOyxO8JCBj1RYB0GUh3UkoWFl8oA9AO/kuQqoDdHhBykE4RQDyFMgYa1/HcOtv/Xo8O2KDfr
vpl1JFhjQRlMpAKtA0XenppqUaQnHJ1fXnToKVyExrvxPa3ZqbZiEENL7v/wuVSkb/5kAFvCOmTX
hWOuKRuTSlQCDrCHKcQvLAIqCes9xqOioJX/kz9oQQPNfNjG9lhT15uHg1KNc3dh/1cFA3ZvtRVd
ddquGfUzC83SUQXKKJFbJHHnPi8tyUJNVE6zRQ7vjSoIRd5qMUqStoaGlw+/7IAMqnrfLC+4JouQ
h6VvlZUTaRH8A8SEGUljZzbMRB9/TnXPqigyStcfuHMATkt7vmBdGqbmLIbvulTGCdGMu0XSbDzz
nzLTal9vzfoyJmnTmN+2qUpigoOpKPzB8tZLMkmqAzZWnZLuL+S9ylgqY1R8XhvmuqAdGTg41rPG
1+rJBbxWbNok6gpM+g/bt8JVbz7DUiGm1MnnYJsk56nkngoiTVKeZHSFVrMRgvPgrhvFWlhwbtmX
ko76jWo+Cdz1RlhwSiCj3jxAvnk3AcbPZmPO3aOlASn++CGUJVkR232GGrpl0eAKXJfn1L4TBoG0
7PojQA/rAPiPGWunaEwniRYDD94g8BgU6hmTkZkTQ4bRJ6OBZOQYXiBVRaEbTDDkkuziKGYAjWR+
xGGxcm+ewFRPYppfkXhWXU78v56DhF3/6jUgTAtpY1377Ne2FJIhy1pKDjhz2iAap5dyRt+ObRNz
sSNKYhbPKM6Tiq2mSt3kRX2FJXtne1F+DtrPXH94yF2JlXNl5/X/1Ta21JPyHFXXh8sAMI+2PAvp
31bo8j2RjvjN35CS6I3nkJdDztjbux2bX4pt/s07e0Sd4AVhQi20KXhcCeRyd2fBHojwZ6R09so6
9EFwezRoRVyyO/6QKVl3JMBSsFWiClAjHRV8UVxWuKT4MyVVJwoAiXfiV6hYj95Ui3OlrF3rtvuV
qIxTi/y21hiYwYEmU40i/3aXT/VYcySNmxg+yj0w1o8xHQQLyZtZnkvVTt5j+uj8iicjbZTUYQzp
ngfoBghfgVtcWErwUj89LZ666vYYDXeNtjMJJxNTwGpK9sXNzvIHuH7qcGektuDgl7k5x1Nn3B9y
+8yQKv2I0ZkYcLHfHN4vplIysbfCieSFrJRYCuDITv37PKb9Zq4KjLzvrR3LMvgOzHCTJzJ8Y3IR
Vw+xPmJEnCKLtgYKxqHY91oAx/l8VQEgxJWezJ097kyiiuZcK17LLtrfM4rdj9aBum/WtL5fwuNp
yUbYBuXWMWCgcVgwhhSOH2qtsCmUhrcysHAfencCbt9npMDP00XSLfVLDfC2q0JFYG+W86FvYSh0
ieDRj0nPrAxL3Z5ZCmGzIcQejuK2KDBsJ/vPQsJ7etz19hXXYkFrPijugwnBJE0W8PQPaBdkA5Sq
vKI5e293T4VI8zc8UN5UNEAB4nZCaNufj260o/JvVFwQjTelkRHaNp4AsvEMsY9Gx5gC1TqOnppL
mJrlajxRfLNMoSzDe19dGY3Fep0QTkS6HE8XOH7K0oY56wQTdQypUctez/TszlUelFUpnJB5U5sZ
mElA7GLVvQlbL2ABoUvzOscdFqgBbFeQuoQAxaFAIzb0cdUvYnN2keuAxkPBSCdht7KV4YrHUmqH
myiYr5czHo6FtbzH8E6C6Hox8rbx/lToIjqzFkNnJFRTSW4d/HKwvdGW8OXPSAbGaQneBUGNd/WD
DxaF/CcVJYrJHBvuWYi3ELyiWSbOKSlhRwlZnZwggayG7odnkb5Ax6Hv7/tGvfNlxUfqD0KIeY+4
jLkVnZG3W0Wa1NKcbGemdQsBz8sstZol4i7WRP72QeFReia3LMklj9FFRJH48RvbV+ZnXZaT+0nJ
CFLcKPPJ6644ZXW1kg1i5EIFpwhT97Df86r5AK9b79Xd+n/Ji780ROJ0iPeOltjlOnxy3R9ecqM4
09I4UKpxaKea5Mc6dt9rfvwLgATFyIfUqLtQre6unEeGIxj63cc10jt0YGqsDjUaGqDXu23jg5IR
NJCPvtRDtfNO57Lq18SBNlTy9YKAxUAexHChsBCw5iHZTusOq73urlfA1gDnJV187iAdw5Vu0tq2
nfvrMC4CQ08ysXF9C09iGl8W/5KYg1qV0hPmRNlJxTm3k+b5m1h4rB0pO6aggCNIzvPMC9xcn7dU
IMX/y42A8bST7eY3I4MXlA0qDQDSUfesCQUhKAqd5HMCSS40GshD1+51VHn2kojUCayyrViJgg7m
lWnLlaQWW5VF9ltXmq5tMbmuug6ocreEW6wYUy01FZHbsLNqGBlicbVMRayi+u79uo88hB2FxkGl
dojOrOSWhXJ8bMl4djMUFh4hM0zV/SRQ6crc8raV8n1/dCHfqvEBgSJ6z7GnSdwjgimKlC3+986u
2u5RHFeh4APbV1eYJ8I6FqE0mJF/HO8Oll/DxZdDk4gWUwLWF6Cin52zCr8htKiqmB2G3ttoym/Y
tJS3i95YYbPh4F8E7IgTzw0aDG5X3HRxpSyjASk4JSoM2/PYRiB6T5g6SfBQxpEkIwrdw4qzE51o
KdQ83Nm8/ujkaxSJWxpRHxVBP26+xayRDDjyK1XuFnE54aNm1NGXx3bMFKcIGCpxaiBILPFddl3D
WUtv5d9zwMq6y/7C0xb4BxTlJ4hxdLnJezxxCsqq3n+Wq0hPb2gAZlOQz+O0c88spdWgfh2s5KUP
VPydE8yNMXVenqFWPZaAC9GVzUcMphhJnabP7HAKYfGb65Q2RUCgsBBjHz801SEQ5Fu6BhBqFr/M
BDqY+B4jYMk+hKzNQEiad1KcYLhvogh9n5zKXWxnJZJmidvpAuQwGeFNC32DWW0biqqdLo0wbU18
SrNSFRWIoxKuyvn8rfg7ncX6C3eRPaN4DqrwC9McL79QxUHyyLmNSMupyHNsJOy6jnLFz9P6ssSE
LMPokCYGJ5sa5e5wziOPwpCM+v7T2/+b1bNwhEfuHepgqGYPQqYEszhLf3oyMYXnEkHFHtgpDSL7
+NkdRCpsGkiLQSUv6K07DIqkLqKND4fOrx63ZDM5Aa5diKLWhwvzrMoQqEO645UGWvYHr4PqXdvM
nG1gCU1Khgw3kpcEbcB47aIHjNWjLcNxAwT1GxmYoh/UNgzs+zJvay+vtpd/BRmQWdzO3UUfdRJB
JavqWmnaUt7wIyevLOPcCYF7jtErmKYjjbBTthxQD6qbQD6H9YLf3+zk8yZ5XQTm+NWFdJdJVYOo
eX715U/1N9yx6TBGLmfzsybRlIxUvzVrz8G3oUI15uEw0ykw5PWocu6qYstwpTWBAEM7NRQLI4+p
+JmuTw/AsBNiRjNOEmBYBdqcX1MPiWWgGgAmQyZGycGt2Qyc5d3q8p8fvQqWnpkrRN+cmAtkUXCK
abCgYb7P6rq8Adyojd10VK50aWH6wrjANUpI4ThpPWrzrLtiDbKZveAU3c4iLyTBoUJ+TVL4OOBJ
TwPEX5/EBSCibgVQWdAXp5pVf1kmiOZnAFEKzEN9jjLxUKP5/R7UyEAs7WsjHv87ImhMy2/fwtkZ
GgP3LSmsMDbm5oLA2trklVNopTea+5hI7x201g8K7rfoemuEgqcHpXP5O2cqXDLZCrpArI2p4LnJ
3web/C2hyUBE6y6pFXGPUA996uN6MGY3nCqw1t/4xSW2dTySEgL6+ho5KaXYFFcSG+a7d9hNAqxC
QlEHjhAZ/j8OtIMPUNR0PST26Kb4LqE9PnXFfAJNyQVmf8OAGTxyoxXe8DoEy9QBDje1JiMMs2b8
3WEmQC9+7CXc77fHYo/DadfduqKfoYtjrr4ih3rmmj+tmNxEfe3E8HTi73FszIxDrAEGmTHRvIKM
M9Va+gU39LBdLaZ3d7C2Si7QkbFv2hQViTpCJMJrSiqZ1q5aMHhanffbmO28Bxb7kWLDA7NKHy9R
tpBbrUZzy8QPpx53qMUjBmiuF0quAYrZa/Y52Lnh4sXzph2GYKUz2Kl3hh/jbgZpw2POp5Fcs7bQ
VlBXsIlmiPO2xmj18YndA2pMBfTv8gXDNu9MWw2CRujQ/Je+jsvl4kpKs6w7Bkirt59ewwY5eUoX
jJwYz9r2TW1DiTbLnvur3wDY1+uMaikCrdY1sGrt8oneYH9T/e7uZYhAOmtFZtBt6haIah3CsNX1
XPgiDjQn8Gt9gVJ0Qw6zCBZSf4Fv3Lhp4em+EVqD3NIKJO7oPdRQV522WPVQJUC8PwZcqup1A9on
HcZIQR6v5tCyM8aGhTk9LZwLz4QGaIMxdeQK58BWcKEFp05XZKlm5sRYIozNQ7J+HoeEvxfFGYqM
7vuwhU0zhexvQn5w4ZEN5OQ4cqSYYxBwPs6JDXyWnTUE6yfCbJ0K7tlkfclnrk3rPpDqTA9a3fv+
mOaoHOm+YiSaJABUN6e7VaLf3EOvXx7oTCATMm+n8N6XvxlAywIZnS1IGFPcDKwMQ0JpdBx1we3g
LkMWYcKGnhQGHLMC/iPyfE+oG7CLFDZGrHZv1/qrKTmC/m5yHJIKjmSePDAx8y9E9uqaK+INz+JS
3xBeqz8OA0CqSSqQeUP8Vr62JMqtMRhWZGM9bPofxt8vdVEYrGOeF4sE++BVTKB+xF3bqY226UBa
7kWUmnOyGni3VH3/cSWOGAOg2oCswVhePBTB1qVp/WTd9VyOAtRVpTNUHdeBYDmyv13HDPc9zQot
3k0htdsSI0jCReuosQtSmQ6XFYncTT/8ICftwfgojkktfmu/N7GvqMYMLuOVgYZ+YzX7a+knHxIH
k/fNhrMNB+qBTkZx7avvU9zE678pizCaxT6IolBcbLzdyQuSn+MjFpzaCTGcsIy3lBK3I5SpM9Am
zHJ82MZYHael2GXosH/cwY4tHSUzFX8LmZ7vPM79bGiaf6mkgbfjwpTc9belVwSwwBTBF8AH4Zgg
aibx96BlR4B5oWi1GooYuf3GSpGOLxDYHiMyLo/Yy9ZRCVCuyBstlw0p9P9qFVhXueF63ExW8cWc
fSyaPPphyQ371hOf6DtqUgNQ03mEsyrToBffILlf1hZFice5xhHLSUyDgphyBXJ9nHg9hpy6Q6Ps
LN1QX7dAdcZo2AmdE9/weNMWE/qq+T0oq7oBO9Ns9nIcu12ON9tl5U54zz2mAZxvlABmvTwe5gOi
zARJTUYJwUM6sEDsw35e2fg2KelJkTSdimRy0jlrQ0wKRKyev8RiXmUqp58IfJE88eCsk09UU651
cDflxKA7fQ1ONJ10FEVENTYxcXvJnnMfV1oaT9IRn2u4G7OAnY5nRwRgdWTVR2e341dwUfkVM/WN
f9ZIwaD5owrfc7GCkhryJZFl1yxRALZ1y1UV9atoTNZwHj41gGMgrGM909epjRddUR7gEeeD+Irb
caShyKiaz+fJ9sNWrbTZejtZm0qSLCX3DZ7fHGWM5iyRPNA4EkM74ufGCLN1D2rPyAXWTWt/mHWs
Le/1aV7gyoRdLXUS3ik64bPhciZpMAoRTu0mIwmJXqpVzY4la1rZKcst5/ChsSUF2s/vyfEgKSp+
4dhgpV+QvqrfXP8hyeUiDS8fDeQT37FCaByjZaRegdtGJM9XUlYcZvaGTy+LDd72lwZ6NPuZDU9l
JmoiKxCNT4oxL0jJKAfNUkq2OIzne4G/UQe9xsI4c3oylVO7Kh+rdk2GMTMRcriTRoKedmX0HO8a
7ikRKp42wsGua9TfPbE9GlC7Z5uLo0RRy5z7ETlH7IBIH3pF+rJOq4ZQn5AMkKpVqRIQ2GQQdBdd
grdRwWivfc9IPDHONNizPBe9YZUFemJdrclZPYdf2XgdlF67V1tfKK4mEaEqXudga3yUklc25VI9
P08pIhJP/J8hFhT1Wuwof0Vh8ravYw1LT89o52tDriBDP2FCi5qp9hDQUpP5vJRdDGBKGIFRjhap
qCsWumb5pxg2o9Q7/uNEtITjj7hP1xVKeJWDaD0pzsjKJKqyqg/FbcF/7c429+8reF2spcfZkmTr
ertv48oxEyu0igc1DomM0SAv+ALBeM+NyawqVI6SZn1sIp7zJjAGNUGq6huYr+Ti+Pn12T+qR+T6
0jpbDDnhsuVWW89WLB8GILQM4BnGvYQaBziYeXLeC1J/jdJMkZt7ShfyJxLR2XDhsrmempfvLmtf
zOrJyCHvu62ZVFx8okV80qgbiDwEljV5mBGRn2LkBGjQj9TKYUP6cBzy6VA4TLMVFF1KaZGZ2vEC
HcWM3l1QiLoAqcb6ERXZzgrC/YttsBmF5k2SSvgAAjtrUPimVf8Cc6dURJZL7eR/5J7bMCXuf2R6
NJz/ZupqdithxtnorlYI63Hy/J/IqHNheSMOg87Uk458mX7gGyRuHwSURGAcj24nGATWo44s8Mpa
I3/Y4IMOK0y/aLq2u3vz9FtYhy89EXI36nUgfij6CKjPm9e17A6M3/wWoDbE+sXOJLZa5X/epuKX
a0igJwdLBvh0llyWmbfTUvH915inmZFGG1YdvPfkA0C1VZmpHm08qldrK8yNGtmA1PhsjFUGPegW
uewgREgeAQ8SOnt75ZzT6XLZqst5qDRQsteEvV6o7fYPx64wflAtfAYVjtJ5xsCC8yw/J+lSHqbK
zDkb1MKWg7AzD5UbbQKxLVKWtqWV/r6jmOgW/KAxcE0ObFBJP4kn4+RRQJYrX9ncH3YxTOo+SNeW
YXErCdQiMzn6M5Y9NmfT5ralsTcKqtP6adQUvllZ/5NSZpZjddHY31lIip3c65fm6fdr/voMfUzS
XgpjVvlVtRfqmOm1EN0I07Mvo9d1cPDVUgrCJ16M4I3q+Kxy2VMnQaJfZgmswJpzIIKCFMVemrct
LLiaCvaBD4uv0jVwjLsqK2zf9ZJ6uZfdMLTGwDbXgGXIQoudQNdLk2vbaK7eLUUFBT0JX3INyYDY
mKikGYjHjRF+/lS21h3jduXfGnNVwbkS0gZsgSpBIuKNjx5WGYllHgIZPGuaw7Vr0F1mfkj3YftE
dsNj4P1PJgma5lwhAaa1Vk1S9Sa0zdp4vDHt1uf8Wcylvd7Dsw5/owll8P2x1Ilx2t2Xf/hy3IMw
bUmsoPzuK/uL8EsLj2nEm10cIyS3nJKGPK+DErlvVVP+ushSrIpIcfwx32zC4bQs/BTgpPOZSCa6
tTONbt97vxqlVYkyhTHXMax0gWyqsAhpa0qryR9dJZNug83oUFY0+bK3DOnd++6KkRYkldCyMjJx
/z+ei445GHlkuL7wS5HMmh5+6B4WYTzrwa/i6ir4kJQnCE8EtAOeKOIoPRckbvjE6k1zcPEOuBuy
NaPie4uMlI+Beshque2Wbw07BqCNDzQcWL7ADcGV1Q7SmyP6vNrg+Ar2q1d9aKp7LelvhPQtLKKc
he8bUjz0cqyrR+/EpTekBPqwW9bPoz9llHoBg1aj6FxdPOrhG+6urAjMt4K/C5gp1ResUiJZ5oBT
7I8xj26zYtMDRxMjx/9XcTZrdvKBKeBVasyWmLoIXLM/ldplT4V34A3Qg8MWbFcf+9+KaFV5SyEd
uD7+ZSVx+YUpj8RvsiHeK22f4tbMnlBv5Kh8c44uzh+HcnyGuTxj8MrksyEj+mj9gK1oe95w9SsH
NKFdOEwjlMp82ANed9snhibHUjw2n6FYI9Pq+/drydZtn+jfv5EsFJR0M2WN20ZJkhxSrLKvksHO
PagDStJv08c1P0htKAz8XJLTK8nBk5rCSkNpZPre3cQaKvptgnugs13Iy8JUPSw7kKBqp0KdcnX5
cBgoDqDACxcr/5jJfhzjQIBs8rK9zSXOGGi8WmypXlKONTxb10RK4FB20sV2EgCC+JnLN5VAAKVN
YnRzcIWyZKv+NymG/QoVglsTcz2l6yWRH7Sgci59hXY1GjM4zB9UnP19DRZTc+bZfa3d61Su+Oai
WehhuOEuyWI/ZfdgTH7O555TggqKDsOLqQqnzhIYJyJDXrTGH2Aosj1urEnoxi3o/31IKkTpGexS
CfBW+Cq6qM3re8ypo5olq3JlaBeJgh/G/Vzw6e2Y63VEmgwAmw97pjWcaSx2NSzRNfYXQhYmoVzB
Gx1II6nqiHahIoxogk7XZhZtfD1gZOfeSC9VLJ19WsCUAjLWZWaPcEqubH8ofdh2dA5svHcn0X/l
hUu/6I8XwuwyKBVJ5K0HfKMCr0o5HOz/OEJF5TAa4qE4wZHx2lgoGVXZ6Tw6EfoKiI4GMRQjgm7Y
TN+/mnNT0BoSFu242fuTG+02FHSezgcbv1Q71o7pt4ffoWhVouAHgL75OCikOUeXiBIMUSrId2xK
Fgacy3MfFZs0RoqNTVHxzt5f3AkPdoCDSboRb/2WWy46EYqMYYcaltFCqq99BTFS7KgnT8ZvtqEB
0QeMOCPDprDZ/na5YkWh1PcLcm1tgusSuDHD4DJXjgShIrMo4SQ1uLLHM6eKWtgQDgeEuVsJPcT7
9QS1O8uJcQ+4Tw/VxQElk9bvFsaat+cju80yZLqjqG4L56YADfDMNY+8mQBhxu/pva19QiQtBGv6
n9agDYQbUAzGfQJzs7dRfxPQA1sslCDHrmzBbmxJQwc0EwWC0J27A+fT58K574R9j3zMJstb+JYg
qjkkKiszDaFw2gfzy1Izfl51+qsm/9v8larELNhwsJs9yZOnrKpmp3giGBt8nn5nabYAPxrKmg76
0zRy+rF2ByebKu3vuokzOcLhRu5fFYL3Noxm/Svq0uRZvsFeGwzfw+Haqe38oQ3RZ3oIrCtBMf8f
7aVRjsYwwAlXmqFNwYuQDvOURI4xNSlhf11BHXQcZWdwiBFUs7rNdYslAgH/sN8y4WadvTkgsSeL
HW+e4wVdsofmTPCQ2gEnlkL07NScUApgKx7jnFjhLqHmkSzQuLd7+cAz5oZcHZVvz1m0WPKWaNw5
HpVyxbJbapNRAm4Sci9vke1osfq0G3ib1RLa9Tf9/mB80SEy4FVuvA3lQdIQKvHc8/cVoqcp17n1
y2b6YdYtrKm0e53Xp2Xwo0YRwIP97qP3/85X/0KgXZZkR0DAJNVomLHCWZAwkrQwEiFUrYrXwe2U
PLk6YNM8AGYl/pKcxUY8kD84A98HqdaoJybMjO4U9qqj1vwIODxddCXj8ycbxwf1zQ/lb4WlRk/D
HTG6tkmM2wZPia6MDcHTIiJGi9TO08sPLNo92zyycXO8qKhx0/613xHH4Cfcud6I2dkg5+hxOnaD
gveYmXCqf1NfBONUR5mdg0/EHeqrbUaOFnNyIdBULi21lQslwna8xgF0ByDQLsemx2EZU063ET9W
rWjoPHUdLJjilErZyyYNTgE7kxOjbrQ2Jan5xeFTtfgpNF2iRjVW9niNmrs2IicnLtF0GBSYSw6c
6yaAAcdIUvqzUtGEBb2SnhfHUlLVrg/PrijO3ipuPT0FhVaM9qSbdGZ5UIBWy9Y7D99Avp/AX+Xh
T9KV0YiDSFdIb20BaH1wlQnE/QrLHd+AqZSluNV7JMCHvk5A/SLe5YC+0a+ZXBqiv7EFewyeaqG9
cHQW8fnbGZ5sgoHVZ3uZ6DvMGP1oCQ5j3CdyXKKg9cLL20x+WIrLI7qoqA2NSWwXuAEAcqFjgSAY
aFaNKHNcmeQ/x81xRoxLL8yzU6sBC3Sf29Lg4fkK316/KlXT5r79oSBLoP0MEw82STe8m6b5BKDX
FqQ+4YPyEWSWHUELpP7chee52G115h/9pxd7OgVIWl/CnpmTb5w10pbD+/g8krxLWbDpBWf1auo9
NMpHGXKY1iRVb6Ec85pBUU48yuJYDQOhnjcF1z7lioUEp4jg8GB/vFsoZKseDX+Rn1aLcmTjnwXd
f1LzaOUyzWTLaSsBX7PtKq9yumPMvlO2uM8z4AEwUvGjFL1O2sXRtXlGrctMPqmtpLOHwgtIXhuJ
YP2UvAJvw58DiklK6mSXw0KDA5qGKb+7acqpCxfRNXQu6+rpjEv+YlqRVe6yGUimz3MOHPks7V3I
bp+e6q5yTcRvAvNLoiE3SJYipElr9H+m1HBeWA931KZ3i2FhzMfrdRpaXnLusDr+avx0Xzf7RO71
wtuhFYEU7r5olX5ncUfbjly5qk/lTx3ErEY5BwmfPUWemZyh8ZBMYhWF8ldYhZFyMiAX9uPupbQh
S0KghNqBj151y1ON+yqnnthZXig5sR7MQMZa+cBiAe08ty81ekfa8n4AjcWfwOP78V8GQKWwqfDn
Tx56x83gV9nPcCCTKsLCzDfKpw/NiWGxPz6LXJNmpGv53rCgDWjoTXHvl69+kLjIQfY1rN9MJrnT
DIEgxAA2Fi8vQzzvWTE4+B0PX+JkJygBVcGPoSE6xbLi5APRRN/W/NCse/89hZ6P4nTm1YEnrqDC
cRUQ7i0ajiRqFUeXafsXhk9kTNMcTejOUlZ1DqHKcGhUKeughO4XJXWfhJZELdzIHd4ohLll16Ao
a6YqYuu7xTkYhKOfG4mCqtP9s1hoik7u1y8pqvPs7rCAlK6bMEuQ4fVtmEZipbv5dqy3cOkiC5AM
YViXJGIolIJRW+y8JSTZdKbWotCBEiZ6sb7uw5G4FVZRj1K13k1raXszfG98MqMNeLLY5unkFk+P
8spKwVr3ig6KmoexWIeydQfdDrQppPhozWkTUnoPPBb1qBZigFNTLG7y9+TgnevZNgOSrfLz/lRR
StiviOHgJFTwQcwsq99D/VC2AZtG5tlSE2bJZD82lCZ2JnqB0rhRbk5M0RdrQkVmXIU4xcUG6ahf
fPJvqAE8HrJRtOMwdmkl3TzeavI4dSRuCiVShC2ia0ncAGZ/zCZIF2pOk6ZiijRCOmIuSwjNFV9q
nJiiVgi4B76eXXXCNX3dJS6PGltVtvjY6ezYEEy6pRKDyYckCMed9I6VVSvtvkc4Z/wxOH977rVi
aCJU9ukI+wFu4eynveZf/4JSDnZ+z3BOwUpTerNZiemOGMpdVE1gZuNiyJLquCxJEa0ui17eK3fe
a2MP3/LtVxvtlxdy67/L9jdZp89Y7lwa0Jf+tJSO2fKy/wbXsa8HHhoe+F6SbGr5vL/ddE91OSrE
MSyhUNzEMQOEiLyPLvK8C0/vcNBC5/b+onofrO+/BMSLJywCVFYGlOhYuWGwafQteozO6x8DzsRT
Jm9gV30D008yZRNU5WVt2ku5i/ES2MrhhtExi7msEmhQNo4VTFwY4K/uNX+Kb4iDp8mJumgtSrCl
5tVEe+buxUzZn3Tgc7MzU/dOBbBvDwqqPr/9IViXP90j6BFnPyONZFRzeyePfWV1KukGvJGWJo0p
KYH7vmKF7nFa5KSEbj7jWyUKdXxWhtHUe1W9j5uyC0II97cCw7VTT8q+/6gKaEcWY6lI2RcsYjmN
B8SRmoCkTGGek4BIhJe+r0dbQUFD5lOM/S0JDvYXZUOYrtwAfXmdFSEUTR4qWkJaj007VvLjRjfe
tKZHafhAZwsLCBC7M9QhAMluCwleW4SKnQ+tfec/l3g3TYaOGRwZO2rpV/m7bLonJJW50obOYNJV
MxrDTk+lrqTsYMGYeqYGxyPnZy4n/WRwz/P07MIpymZYJcQySWNhTQ/eXIkbyWDPZKyGHUSiaw4c
T1DHSuX1l6AzpInJReWJgCDcQgf/lFzM/8sNDGDHCLJDQcV2cdHw/MYhm3SUwCKPjeL9bPsgup8j
4uwqx8eor1dNibNWnw0iBlMzQW1ODWuQoIVEkFiQ4KB2gr0AZqiT9TG6bmMxTizLFmYCsIclUfoH
cbLccDWZ22oBV2F+Nio92xLvgyNcoKN3qATau4DHUShuX28LSEt1FhxCMOxTFuQ774ig+rb+LuRY
bGz/eDlWnfx2d/i2rvHJzkppNvyMw5UZjQryunn3JgZSY3Mjhb0/nnuw6+eBanjBS7Npg25Q26Do
H6EM7X3pLtLr2VufKYmnhEQpzplk05bCDBVsqpL4GQsIL+UlnGgdtilYOL8SaxKplSAFftgOrTV7
ZKZJuXXlSeMb8jNUZ0ULa6mpwxYWWSzSgZvE/adYRAOGB5U+P65M+uUtaEaOGPJRL3zrgagDAJdE
d9O/gDe10l44i/GE91CwHhJ39LFbxWtc8rykkKWxE7vN00o4kEfSv27/r86WmyUI9j2yTD91lFLJ
SjimjGxWJVnPqKAT8uRhXa6rfJVZXvx/si95lJ9cWdOZ6Rd6fuN22ViOFNkWBjwUNJiQ3xk3T4ZA
1lMLfX8OB8V1qXBus/oQbWsfCG0aScYFe0aPrcMoA37ix6pGBfvFLeCZkVb9mRzW28EIGTmtmB17
7m1TVy0gfSZkFqhnJqcy+UTGEvSc1Y8IGn7wAZzlKVWrfS+ahombmCyu4PLyrRkxCzpQDLyooVb4
EeuKF+NEyDCF0m0yoseLEN2aEiA5jiQnMBvR2HFgl+pJNkBSX3gI43Vs6wfFOUS307+qEvDjq+gC
E2G+88i5K5wdJfn7jSol4d+jJlxk1GSq+wBLWvhNtAmmLRfl15W7fTkFlZimbQSvBxoXQBP58oRA
LKDUtxO01o4700xCfKwcMC1QbQR0Ljsu1hnfZOak2t7TR02L2tRRYnEAdFK3O51Dk425TYMjK+ZY
A+2MUVx0bkwDCunJbW3nNjx5wDv4F6OEAYiMImERCBOPtna4pKD4Zx3u1pUD/aPnZIIRgfdOoepq
ZyZXUt3C8tB//QMrABQ8n4W/cvCs11Im3ovQqzQIxyHaAmp7wtym3SuzoP/T3JPcHxJ3bSvD4UI6
SJ4lhqCM/yh2JohDFPvCjIdYELms/GqMnQf48cKBdnbN3OfruZTSkKaZ4CIIgO7Jdp5CyV30XEUh
amt5UmTretTgBZB+kQOltdprukpjcO2DZonnG5ahT3K1cpBKN4oK2qePlcgGelae0sXzl+ksWIrE
ohSJv4H6oNO04Ev4VL1b/o+2iDONJkvAxOmhHKKjXFbPf2T8wAbzl0Q6mdvOzeqoMowlF/moGY6j
gFencgkllLLwBqObHtGtfJ5XBDXWC0uhGMm85ZvQiZb7S21fJlSuJ1msyGTzxB8Zl2k3Cbh6K8PK
jw38r8OGRAE7l/evBKH+ZM1Dm8EGcdVNH4se+/WLnsTsyCjLcx6jUBdDwLijLi+FWT9qhrgsTUBD
zx4Lq+jcN1DW1HLfjPtJCBRlY/f3U6lt/xTHp6EStByHD8LnPq05PfPh1TNCgWuD4yPzalOXMthd
4ZKel+uLxgDAimPtPa69bgpgGw58cqCSEYQ6Fbwh2JI0hFANlC6EAdoIdkzPOXTDBVuGZ7/fpNVa
MnvItpaDItbZHEO2I7kPsxVF0ObCS8Gy1JJOKHAVraQZuLQ6a7F/UbTsffNRBJWXWFE1W7LStYun
9a/1+nJ0S7NWMBtRDdjEEmmhm+qIi6+8BFrVbajIVZH3J9dymn9eBJEY4B+L2DJ96UOh7FlyZ/EA
bD4I5ER+S2pQca/TA950ZR5onCGCuN3yt7A49+X74jq7SFlFD8W4mk6+wOFpYmsgO+6uGpvSwFrr
8QgRD3DX3X31DFlRrEMuwgpv+NggyAJKu1cvHT7JdUDGKvNVu24KhAsJ5E28pCPWibEK3y9UGNf3
vwmKNpU8jSti08A9bixyyuX4ldd8eHD3KoKzVwXuQn/pduuPW2cHOTbvN6LYcRnSN7ohMeJIyHL+
IGSKud6CJPQIz2XCxorVfpzj8mga3jbQJEnVYNUd7EuCEie/qINjM8hvxtNODGjZ+B8bT3C+XR4H
tQ1+1083a03KHEN9MXnhsZgJj2bC0aiDTRvviaEkHTuAQctsLwUuraIuAoDtTYcD8ONUmLCZHYaa
0K06wZ8TzsfkbWYzJ6stgXsTHVU0mQqty6iX7XsbiqZk2K2qjVHUxuXnc4jbZRxAPvTDfkzQuie1
PItAn+FzsFoKRJyhB6+/hReM4YZG7OxzFb/QlU/Zb+e2Au2AwFlYrkAHyQNURXPNfeTWyt28eB3c
e0DaA8wzj5lnIJKkARr0EDKiBmJhB0vjkq88tVNoHzMvlxKFh3OGfepNRJgUf8iXUq4zxe/OscKe
AMTMxrBskx6abT5xqsy7kLpAAjSX53UmPxQrKIbr8Rbcpuih/VKxyNym52dVrbl+kWSprLfN5z7v
9vZkYpdY1DMxMFRh9q0HfgDGFPmupxpo/A2Mk2BzjR7WkUyG5Gnk0c9GfSnKH4Yh3oli9GHEfsWD
5kjuZrZEzYyNM0f5fLuSb1k6rrJbiMmPQrS1Dbqwwv9HZTiLpTFQJTtoCuOGOgTeMnvAZZDIuuXK
RQGewVwWQm01ljDO5DV0O/gAg+TPC9ZDWvA6lDH3hM4fD+NawFaMCeT9KSFLyn+B1jLqGbRjDvBP
FsXO17B6qIfbkrbxgIFCBoB4FNL/6HtHdD/ZfFfZE6LvGi+qbz9XNa6smYjpI3OdoQpr7sw2YOwE
Kr72SLh4OWGdvlwSSSSpbWlQkzYPfuhx/zHQwqDI1NtTvXxFXQeYqw1B22/ityLBwAnU/4nA9M3X
HoHDHnvqsGJ6FWmQOjmjVLyPg4d6nK2TH24rw1Qg2q5i/FnsdCz0G2aox7/vvLuknskWQ5AwjFy5
Wvpj84B18GjCGMDLOGl/lUf5J2VirqvmUiEJK6iq817TgBPH1ILh+Ub9UXB/qd0Ep08wfb2tNpfy
n0xlBNXchXFF67RQYL9uN7blRdAKe8Fq8qnKWybdFhq6R6Ms7E86rzv801/Wj3/EInfXVZnycMMm
REkRgUmT3WoI7ZYbSz3IvBGRkvGplUy5udqJOc75/EBsCWytVamaPEP1IqAiIXye9ZTneIrkdYjF
8E/Z/1klbL/1ye9l0rabmbPH8mWQnTAslsXRDEKTgzV8I/nxD/yX4wpmJimWNOK1nLtCVylKRC4+
qdK0MBxBDLkixwJgpwqi/UDiWTKcmO2ekdb+c7g/efuR+goW94jEaZM5xN+jOMa2jeX4AtHwWGCB
U9Efhe1JsQYyegI+hefO/0mwPnRxgSYXTDSkUbSj6SjTndtpFNF7igVuQNmzAm8+UTyTz5aHg/Wb
MuudiMpzrn/XJ8rUYHqa4VnTV+2rZr26/17Ty5Q2C2OMMhFBSM6KdscqcwcvbIoRV+Gqhe9T/R49
63EQqy+M1Z0UJzWchbZHMMuSSKj/Ax5rxhgcEoXALPed1wwU8DP2ZMhItjlh/6HUDcg+2pwxGgZZ
pngnn36E7rZWLWMJh9J7cBkhVJjMq6rOyEBZgIyXUAsWIumter3R5mwafDCmZYays9gtLXJny8Z2
XTjvcijZK2PKmKoWk7SJZGmlqXtNaXCumYdXEWkUpc5K2U+kx3rQ2VzsnqiQGAen7Ucv2VTHt2UZ
4OPg++12k+eBFsRYuZOi69x7+XUhIDQGNcn5XtrLcoK04KlPeQStoGHa7g4ELFyzAc8hiytX6cda
oOlOb2559Phf/B4hW9Q9mj6eEPlEyApsmBDcC10owx2YiQyTV2ZTDtwnnJRRbvsvjScwN4Jx0AjH
fawNEbhjLapAxQh2+uXATZ0IOT0bup9Hz/q853YiSxBoWJHDa/RbL+/JKj2bp8Che/iotyeiWL+O
Br4emHRaWnY61/GLC1tSx4jxhDwSPDMM6x9aXUROajPsFbp31w5t6jKtiTubd3QhFZTzTV4ATN1x
pRwVgWQ1BXn52166WnoPnBCTwLjCpc8c7djXDgUk5cXT38bW8J7j9JkL1BPIHUT+Mlugtn0qS5su
ebOP5kn1rkpN0Wb8zn+iJP74idu83He8mm1PW8CiOsDW/Ka0X1/FYksS+2s6S1NbuuGO1Sa3U2t2
4G4yVvI1RSGLAwPYNRtoOpI40bgvF9nNw4NEVX7DWieCKoTIgG7JWtAnXEhmd99PT8HsBvvoMcAr
Yoa84fB64YeNNIjCT46Smrp3tSOpk8Q+JMwabrg1wV4lUTLNlGK8102B3A+A0Fdh/m1AvHijYf3A
TXP7sC6E5nLpl9A6HuLNwEIXWBXP16Absm6iHLhaUpkV3KBNRtTMYEXnFj3XbhmszRbMoXwVkN+z
M2hEAt9BXn8mt+/LyXGNlkbp68jAEgtjkl0TLm1rbwCifDd4qGbVxF0Vdbe3DOKFp/25RBdvFnBX
BCclgs3krW7LMAdchb4FS3bTg70KIrRf9j9kx2Oyybdu7fnZSWhKIIXTmzFwfLOoan6mu3jG+lVg
BJyavKOGusY7lps4REwDT8Hm7G1QEwSKXJQSXZrV2gDZfsWDJq39a6J6b8st4O3WU2OPR65faQw/
4XywFM6iTDvRv2yjgYH/KcVx+Ldkp7aNtXT+AXkx1GxpePDGz9Nw3Umlz34es/3qci33jHOeAirw
iXgwvsTVmVnZnLQpQFNGr8mfLreWZfSA5GLr8dRmiJ31M5XrJF88vHJwUPMdrusIzbirUA1wjii9
sH76aq4objXC1WZBFUWWm00t2oBYxF0w3gSZ1NQYxLCoOPlg+JbxR9IQ0S881GoWdvUjK+1Peb/X
kHUARZ/jL/zOKyDzk4A8R010wbZPVg/bti2rnn/3+5lwhKRHPzoYFMXcLre1SYb+To9v25wk8iEV
iI2fYaFfERAneeTMpsxNxkcPGw6F0yZiSnItD6P9lH/MBykflZoTWEjs4b50oO9F3bBVDiTegtFr
WARDiQQC+qfysLUppS61B0lYYg2eyBJwlKKokvCic+BPKONxz9AG4QR7g0afuqPjk0tj1STAnf3J
cZZpoW6kAvM+bgTkONQzvv27rAzkWfugfgrWW/Rn2mrDHEz34D+vg4QNIJH+Qxj//epsOmr+fEVT
i0MEfyJHxU/CZqMAaBh31JD7smXHR8gg618CUwvAOaetdj+ScgAADyUa0k00zXgIsio/0Y/Db43p
dcX0lL3iyWq0X0erCQbxVNKd3ZtWtY8mYuEV+rqe9tFMzZmDk2sSvEY+38GTQdT3P7Hurp4Io4eQ
ERWLrsPuL/8owi1DSZxJxmo7/cY+rh3sFaDGEAEb0yCLEZZjn+JodM6z1ke2ImVXTQuIJSQZJTJb
IjjR/Q4i9Ze8Amn7PtFentVjyEDsFIonRtjaWNpMbt8PTECFZg8FNO7c4vbBKcaJB1yCknDEGzss
80A5bV4Exfd1H+E3NqdrVj3WEDWly2ub8ogH3qpfffk4aminiNyflEQUDaEfJkUutrUnmij1/Jw2
IUE8bDFc0niodAqAwJujQU81wGpTRgJR9iqL2dzilvKneWojofzdSr5VCq8tIUrv6faXga1Fb68n
aegr/Y7OQNxCK9TCu2XaMo/2edne8DcFhwd4fezfbK2BxFc8dNdRvS3K0e1Hn1Y7FqzBwKSc6cxD
obIPiLufw1WkEsroQcvS9FOtPP9e2hoKmIUUHTwNVbmMiKwFfVlSwE64WyIDZTOpMTLYy1YmjHfR
gDC5rOj2M0T/+L1rZ4SUfG7k3AFVsB82WG3aTjTBrCL081noeWWiVaFjmtaa6gjiuUuonAL/bPyt
JxKxLzhyWodz8yDiLRf+DgjgRuTCuEHtDWpNfioy3GsV4aILiO28QOcPRFp1K7vY23wpuo/XaPL9
qafn0Y0TeYvRM3s/inz0ldi/Md/qUOMb3iDp21IWsxfe4lrP61bGNToXHUGpgIBN95slYn8TqZV9
D1LsC14bbcYNk2JaWa9WKRgSHJooj3+UgvGYVu8Fo08TxO9sQa6TYbc3WhgKewBS7NQzq2X7gBEF
t4IjLf85HEGaLsoSusgvPjs//GQhxVjaLhaxGO61YWIKRBB/DDnjJUO628LbeoZebjTteuEGvAQm
TeZh30ugSIarDuLh4oOryQ1/lxBHCse0DLHhsmJEsxtknuuQ5k4/Aq8+xLV/5KjC2cldHFbkjQDA
lZD8EH3yZjemCHJOGx4eOkKD/HsAetOUsk4IsEop2WWQ0+P5AdrSAtBT9vujh7SoKt8FhcG2tgXX
7tdL9GO9yxRqx1KxFvuaKKvBPTd6KiZYBLSIgwl8Qw/bATQ+ASgfsJq3VarYL5Pcc1CF8yt7lcUK
euuYoVDQpuAAiunB7fslMJic5HJ3ZoMU4I40cMJqndc16rr37/hZJHq8Hu9a+YERDXEaa6pv/mrW
O84RlrRlkeI35kdaiTJb3+xzV96ippzwJbQgprIvc9TOJkd9DCBeE9jpCLb77p3yTFjKzxJFC9K0
DMkSPle7XM3oKGbhJ/0ftlZFtgomP+PO+n6WuOexaWKwgL80azNq/h6AGSq9Noz+HX6UIgK0PsxR
VOIto5SBGKAlZh8qSzZRTs0jdt6zfNhdwUkrMrgkW3kiiO0kGsIzRdBs/kl4yfE+zlzuqIwDxpfe
zVJO8mi+EbeSCwYyyYGlq1WEYRo1g78exO4IQ3xippc5tvFU20hYSWTyQ5LIx4og6RKaCZKf8/xR
hYI9tPMhkkRYNLsIFH4jUUvQG+xkLseY4M5yiwLipk2/IzN5y9fW0OsvDDgUPuBREE17tRSeJip6
KPjq3v5v/s3rC55ff/0+QUzmJsXNU4sEPTd4TX4Rih+iDn3G2fR/OacfyQ74tM89TvA0WT9PdDJ2
+heV7u88NE8gpuxl06fg2LgG3wQ6GdY8rQg7WP0lp6kzDqppK3dkEhJ0Biza3LLKZyn2iwyqjbWQ
0I+i5xg3VjqXO4gTeCSTITES05KsvqITjfFVocK88Bfd7+zTv6xQob2XMxqnjgOVdEHlB6oyUJkp
qLtOE/Ksc6B6r9Eo2UObOd2Heta0aNE3nI3pgdW6rYVfzgOsAoqV4AHYQYqQWHVpAsro9rQiGBlM
m7CsB4xHjT8jArg7RWA4YAJ65xySbR3++paXoAhdnv6NYSOiJUzXo+n7uf+YwpmMbkfwW9Ui8iQH
4Vl8Zy8a4pGxwz4W2GwyiVkZD2AH0bS5KkTvthOa+zE6PJsxoRbV4vty7eSve1EpTnzbkkVG2O+U
4Lh1I64m/hOwEhWkGWXDxcr4Nx4yt31aHvjHN0i60xAZjRoA/07WbM7kOSEwF0QaphHpibHqS7jE
JtjTHsOfs63B6l7MYCnYmVU10Wno6VRqm5gAX2CO/wsMkI2xVYWWqwruZ+b2cRBYE8Y7HwX8ifNU
3Hg0U3TX9zHd1xYTafCNxTh+UUGXCsp+ugeTfGLJjPLoasMclyjelYGZJo8BtGG0TXDT0z9EWvDs
+mwF8Q1MzYYQxBeZFEdHBpPB74EY0jPqCncUYrsaGIJayCONpa65fq7P2AwJjMpJ3xBt1s2CoMwc
y9NG6QY7z32qmqQkI/iTmYQscp4oRaAm9Tmp5FL2pK0H4ZSq+ld0xMNCOfMeZfowuN/cMv1vzEKM
gmmVf6POEkKQWNGoLeXrwVIl/m5XMJf/9R4P/XVLaBWkR9n9F6n7DcDWUrfKpIDI6GaiyK0yPGTa
prS7bvaBqbG8jmSxJqIZ0l3CeBJfTU01DduVsw1wCplXk8Mnry/v7LO38EiuBEpzbTNef39a4wTg
I+TMMJSoKmS/JYZwc8NiHqHtUrSx3pw1R6bw7D9o5ypCwAMihF6+jnFwxREua8kV0LHimt7boUhs
dKRxxcpsnhqg+Pe4noGFiD63Ok66nLc4jkYKtwlZ+1gzP8F/nShLe3Wi2c2wabi6bTM4cAmHetBt
G5YM/TjVWmcOpw+6qXeEJmtni86PdeRmjThTTnno9jqD7A2hCPTOeU40kZGdmKHOoDPNtmCz5AAP
mT/63Du6d9UIDAUKRw4r0YJo+wx+eHzs9hn+aRBA1kP1fvjtXKpEhDr8WMrNmdkPXEiUUjoTfWwu
LQ59Rj02FBm17OEsNARttRygV4dfqKsHN7hj8k/MsnDE/MLes9+U0c/6UJ+JrAuCtzZd7GS3x57F
DaUmgMc4DgFO6zim4eaSgoqFdVtIHwb4BprNAVef9c64KOMOdjD8fzmUo7+aR1WDSCVKeNMMVkaj
98emgL3ZSEULx6WD3L8y7RHNwrOR8DzMAjq5gZbtNal/l4FDfC+KzbBTlgwqwIjUVWWt4GyU5uzo
R1Z8582TEQBMvMLOcMoyJSpTNywFe4W9NUR40eiZ+u8DiIoCR/DpMG9zWp+F4rY/XEYrGO8ep/s7
+4nLqEuL1Cjpb8j/LfxW8GBW6n8p76qDzlevZbY9Ls0/cxk3PMb4AuiC4qQosA6WcWseBmT9l2xe
UG7rTUisc/f0VMURYcEBYw6HXQNl7prB/G86tyErWkSjBEG9rGk9tzzNmG1c2aYYIlDd2CXGwYP8
ExoKtUqNS20CcEiKduUSdfrssz82Efvtnmn0G7VjciONJy39ryj/tUwD0dPjCll8k+yZg3uFwwxd
mZGMEDURHRy/1DSXvrgMJms5XMZqzGKH2HztjyLALv1wG2NHkWGmlVMe35GoiLle8gfLKh7PQxYf
9GspPkx+eHS9vlbvbb7dc448smlWOG07MAOYydKkdYOQnOaA2b4ygiT3faMUH+FFhg5q3LEx+8eI
S7lmQMvipn0wlRaMRZtUgpQGFMiYuMxjFs/qIho5/jQruwJV1VlkePIC4Jr+GLZH8mixwwy+6JiT
w/Ip4t4OJmfR3YtfG4XaV+cKoRlZZvJPUNmGwTLR38UznqRuATq75auRhAO/TcWpBmOgBFG9qz7I
KehoEvJG+oI32Q4VApDSaKwCLktGY5j0TGS9szNvLkr98O2xaweArQbpPuicdxngl5qmR9viU37A
n5Q4Ssw5CXWLfdcsUx+bMpnLKj21EoJklrBZHxrYkIrgBUJO9U4jQZKvgkrVYin0r6kEgxvlwFB7
R26O3a/oY6XCPLrHwZIADsrRt5N9Uh1nqwZxmJj4ML+R2LTUfBNeO5HGO5qNKQC+zq9SQDtzrVSK
hh+sEqT9S+NwGizjyHO4ycaH0g9jeZjoTZBqhFtL1kdJDILJ25MJzrmGZXMJzp8akGSIUlPljYNm
QY9KAyV71xvMG6NchLvukTgj06omjSHIRramluApXYsORaBuE8Mb8xgtyeTFlNemavyKU9a02K40
ayMLB7S5Xt3q9CN3nZzwYL5TlFMS55uMItXG7DkNKW69TogHyeZHWfgcUdgqO7KiWYpvjd/Y8EkI
RkaK3RWl7PC0UwA7Ck18xUb2rqb7GkVQZOWm5uWTqMnGIoZaHYu/YypSEIZ+Bo/WbdmE1QLRYzTl
BllpafCuRhW//Dww6X9wFTSY1E9Zt5xpTclpVyFP9Xawmda7KryuryrhkQ5LhfYLZ919PrseMHn9
p3LrkOJctDyx4DN23qjUTVb4h402xNoZIduU+2WbS5bZ+aSQZCYmMEYTrrRdzGEIJKhRYk09WP9h
RCl1l9Hp0fVW20S26l9L+evZQ/g/FMrZAfikxdrxjdUu0atZwyk+hE+QVoCRKTJaevL8cfn7AR7W
kwT4VyfI4Lzerj/UMbVPpH7JePEpeywJtzShRqCtK+QnlNa+HaM5qAJd9uZNUHFnG9ml+3lS8yzD
A3C+iMWNBxGvzlHK46wn4I+PJbg8uFbZguL2dRzn3n+yPgVL0xiuEYS/Kb/YCGqQVcgHlUzV620R
O5VNDwwkBreTdGTVzuCSMJiBTPqdbPCn1/5+CZJJRWU2jKoaYMftYAHRSs6xL5Yt3tHWM9huzwOb
tK9aLKVhvqOIEHLQBaaIllphGCKtrhuey1bs2wDab8v2TpzoGi/0JwuIKXACA93WvH5qvBECAcr8
bLB2bGYswfCJJwrhIa66C1OjC7KMr3l2Ex6pD010S8lMi8m0QfTM+PnfXofEPLimHfnRLGvdGIlO
O4rR1veRBnNAjBB6npjqyqkxEFtkmb7rMUmpD5p8qnvcFxNXfhe4op4HXExGeQmdkDWE20Gkj6Vs
TBs3RMhjh0M+ONaJikAx0oFfjtTJZA93NaCaPpy7/dTFVUPBV3b2TPWXc+fgQOIF8xGPeMQP/zWx
ed9oePz5Mm2O3tPk7ep3J6EEb89FzGULPppaZmwZLoy+vLYIg/kLklcMHaIH1zvhftnISLPEcTTJ
hA9sLIpTpq3zL/Uj2sRT9YAu6trmY2AlChhRMYqbzyuB7YaVJiWs4Yka2lt9noSYfdqg+KtK6Puu
6TZHBvOd/VMlUz5kNoCpuTKVSqYpfFPE5LHE9Yy6PHbzdP9bkbDpmh5pUPT6wT8JI97hmy8PNL29
sE0qIF0o5JDVjySi3XfqaXgcfHftSBKikm/77W3g/A4bgx6FtVr1NkTcjG8GNUt8s5eFjMu2m5aN
qf23XUVQplOxhHYaYRpEvcFnSdtH4n9g0ID7PqTFOEyM6X7Rvs6+dwsU8etUQBDGShnAngIQkBPF
teQabfivQgv+810Ef0ZcWqqTr0F0eeBfyBa/gdaYgQTUMLtk5u5SPR9uY/y9EdgwgNPuY7YRf0/8
YyNsoAEFbsZ/VuxXM4g5XtkPVDZP8bXbna9MNkBcJzGksaffkRmB5/o3467RHhgd2NTYfrKGC7OU
5x99uuQTgxmiM/TlJtEQAM62xZj67s9rdrMXBsJ8ZGPrrMKMBuZ0knDuVLjaV+WnO1+PRpJ0Cpg3
gi1/ZYMEPJun3ufdIPh9v3daSmI9L6ibgkY4ccqHK8UXWUwmJcszjOf8spfSP8WfbhY8aOb8itmp
hifeStYdq4gs5kOx0EKWlm8WjR7y9Ta4M98GCanzAdAGvH9GZjWLTxL2v+6Oa7dr2IpHXRw84zgs
yrD57ESvdxzeVn0Ra7gf/hQO1PQ4DsbXqZvEmDCRQGXVBszQGncnuYOWRQV0CVXnVODZ4VJQvxZR
Oe8RScF+9oS3xPUCg/iHZ5wB33Z3x++FXkbe9eU9APtG2TBGiBeZ/E9JihCtB0N9OSAMM54EPTYi
hpid6/TEB4SHzxWzWvnr+uLM8pOlu6DQ/U6RZHdICeTjLacaEThL1s9dtS9Fj55rU52Y+WI+OGzd
gi2Oe0TrAwoH92ZLTloNlh9HPOu1Xd4sZcA8iL2j8pSIk98nAMxXwWPSpRhXHKOkvKW2Akdr7K/I
W2jBDmYhW79R9t8myfyLBBfPYcWCkvh8MoRuFo2ZF+DRSuTy6wlQ+J2j0PAHeY0BRRJHP9YBN8BW
+RAtDP6W3rdw3GvAnDYyg23bXZH44l+DH0EriHTlYgyzBwzL2JUQzFm6F0Cloo+j8miFnz4ncSZA
TBTtjevy8A3l9Ed1MSvv+QBggZdO0siFjrWWagcSCE11CDXLwZ8M6fsCWkoJh0p9et+nkW0if3xY
xyw4dhw4+I9Uioy6GHPFDRJT6GraeAW71SmcjdSurOSmzAo6CjVTb0EsHOwTH1BlQXYvDCK/wkyi
iinrU9u1ewUxykXbDfIPzpLkGFy1CjFA7tJhm5qq12//45ka+2AO+MdI/HUXKuSk2Hbpz5Cu9Ubf
Pvl45HYZ9UCsFIFaywG+eVs5MDHUfzqIqkAMRAOYgpMxcedy1jcD9Trcc4Q+pBrErbyMVgQLV56e
J9RhxQPVxTvbAGwvns25fvxXfpuOqZxFDTHpDoSbb/V1LIDlkMvFVZNPFamVt+ykPq5QI+ksB1BW
DAkOC0IIVCVMzJkDCX01trBF5kr5uZGqiaEWCDaWpZ8Oy+qeBNc5zyZlwVbwnM40wWAnkpf2dNYI
Tdtspx9qa4iIlUVpQ938+942x7Qnk5dp0/sU8/4SiINXXeiU1KcPwOZwgLWcltPWgi/G2xBZYdpZ
0D31t0couQHZRVNzNbrbaI43cnLG0OOi1meRABGFmdNtm5at607I/bwqQ4aD2OKSL0kvGYLum4/n
TS6bLzkIaEr4TU3E9pFkr7fzhU6vTpwI/p27/Yjyilu+cvbBo5UDBt0sqLzDgXOxHSGdxKunzN2K
JHicVtUHywmPrpLcOFbQ13fZK74MMw0qiVVt+FYin2RsyH0m87or5j8IkS9U6TG9wmir8OCpZ8uK
sszd4WhnUKqZqORzVpzWkp0ffNAdyJuxxL4ZlqeROKmzhMP9DAl117DKLnBR1vZiomrnm3DNje/b
Jq9UgtYTldvmp3QhqzB2rg6lZubopLVUDReizPzDaKUgbSeRzRRFXoV68ljYPGWo9N8HQVxWfyHJ
XbCqsp7Z1lFnu1raVBUZDDSl88I+luQPattRqlcK/G6gmIaEbprawDDV6AZBa8psoVS79kCzW5tB
NkNiX4I2Qq8b4e01jHoDcP4mNR4YVyKEqjlwyVbD3vE9VVZdOFFTOgHiHqU5LKu7XojVRUrlNslS
bw7aD5dRsiykEltGxrPkKp9IHGk6N1DJdY06FcxBuw7rDNo/Ik+U7GQ3VRuw5ONi2oikZDgC0dzK
nXQVqahXcp/Jl78aftj542FAlfYHJ4qc3AOpur46W/K+xMIbCYZ2SjxuMzlVZU53kIrWXm1bqVQa
NC8bJdaLQCw8oZRPi4NoUD8oBD7sq2e0yP3BjuU5V9XSSnLf4OWusk3aExcnpaEDK2bNHV2EFewB
qetv5hlyKCAdVcz36uIG+CLNjEkz+GnHa9o1bLAWf7yUE8DJDDz+aRtvEl9WIEWcpcufub99mTcY
0a2U9Aka9PmoZUCPwb2i75DCxSb7xrSro0GZgLAK5kyCncwYxxi3my5NCXvtujJ6VNiSDK+ub1Yf
l0p77EPnscuoJ1wnkJvMRWQDFdJ1lkoNSffdpHAhVL/C5zEt5j7AevRvec5s5g24nRcFPxXaY7cN
k7lHPelEmWrZqbXAoebeOge35dWvNp5bUgOpEXhjpAwbHTX0ucVfI28NWSaMGFOtNi1Uyduwo98M
k9XW5JPEv63zFFDfF9xt6dfErcFwfKN9DZSH5nk9nWKHMHBW2Wp4DMgkmiP7SCVanb1XSh3Sv7i9
xm9WxUsI8pGy8ugSkUA9Q7hXdfUrGwyUx1QE5ePl+1DukBnvit8svFLargwL8wCmU2FfD1GjK/vl
5rbofggw05F8xdE0W6PL4VwLdGRq04ZeM0UB+Nf4/IABHZ/UYAOujblIuudbJD1wjdnBmfTk6WFv
nOR970e8OWTmrnPQiZ0gr/pjFRJ+uJw8tSBejLScc5OLLMbmHMl+g82Da+5ISVWc3KpICb+7Rl49
vm7nOYJUgao51FNSeKQ+9TvyG86tolj35fncgN3/eMETKKBRpdIaqY+svDjLXofgyvV3eFa8KEPf
pfrpXaJ6THcaKHgPcBt5k5Lfx9Woq5IUF44l+sIZvsnut/hinryESwEjJixqRIrEoQJQWxDNQ/SZ
FaPVcsIpUG7/o414yIJALYu1vUU8MzttYVfxnzuO42RWDADVgp4DVX5L++sximgXTbU4cpG1dY6W
l+DdDE/N372/ASioKCrcPBnY2lSJbQcaF4Lv0M5CFWIllsPhckdIPpXG1WmNx8iLTmJrnIBU0fz9
l0pTInCxFlDKQ455v2vz7BVDkqVNu7NDnn4XUXOIBbfjpEKhjIDFMmwJrgqVCWF8s9CAg7PwRxPz
SWH8UoKm8GxrK3DkJfz4/Nc1n75xZGLCpfUXYiAoC3HkDFNoDcRH9j3r8Rk2JSi2a70lbQmpxE4J
q0cfEDcREyWkkWRT7WFQ7aqUhvIuSZOIYrofHICkw8zfhTzqiP1EVD3akhWT3hH069/CYZ2sKJQt
iYpddFGb5bMwvDi01A5Oq9iw+tc/U0uKX/ky7GRAXVmru6LeX1ABoc3WFGtxk0zKJoakTZUHLtZR
KRiviEQCP6mLiXzWV4JrQTqLbRicvKOnJyjn3gIIcTbS3N1FULsct2Oj++0DcWQI1Ofzm7W7cfA0
dfpjILZBYprGPDKoCcrzkEUmVame5MAGNeYj8V9Fh7g1fmmjQHW/75INq2bwtTkBpANuxgBSkuN2
SHHJ8C5mQnF2O4M25BLk8QTbArzlVE6+u5drt/djuKeo3n77gXDbXPVZCJdxauUCjE6Lk/YTMhF7
L4WGRi3D8+D1JaGa5UGppf0jHXLDaDs0X4YXjJ6IDVYh0fdw+4SUVJyxH3ATYs7RXcdqROrnMhjE
xBF89hilkl3y26WkN4p65SaUtdBIgvWSSteumFEzyS9ANcr6vlhqbNojBMaTIuwS9F3/yWtFJp91
MC/fl20ZFd40ZdGQf+mImW9oDUadtFT8ku4mr0+1a4Hh9cy7vTVGJzOiKACrArOyt1HJkatu/MAD
0cf/5/gSekkH9f+8/WLMA5qJwtSY5Npz6Ov8pkY2n6yDhQN6MNdbJhMSaYZLAqKrJd/X0rnPe7S4
x9ROuAUDxx+8PHyD2DTfPrMUEzaJ70Z+vqVR4gO67EGL16U5vc8MId8XEC+2fztMG09UaL20ohYH
e5n2pfgkSbRWv2r46jgVXpAIn3baGQP61dmxqtEacvoGD/MIZ20h27bimEpjS1tuRdUF2WdCJ5tW
uXqyUZLIih0rOS3+cmk+l8gjIy9aGvO/zQ81zSQN/EEYk6exgkrIPh/krfp/Ihx4OemRw8qzyuHi
b/hlii5GLe25o/IR2T7MR6J9lnS4i+qJyynNb9dXpCG3IdnfqOCzQuu2pk6Ljl1R7HfzyFUJKVuy
p41i3k7YZld4HT1YGXUrsl1RJPsJ58PSM6hJXBOACtBpFPlgKTFAs5N6YXGkY6RSM2uBm2perbBb
FnoYnkyLz4Je4W8x9cbctzR6TTZlRQQb86ldqlAYoy0ERs9YtvBk7u5BlW62+DPrJFY/RgzbtV22
vMN+PhHrege8Am+HlOPWBWTqb7lHjgX+D22cp4ChXCjBdl9LjWzeCylHMtu+X5n3k5Ut746YR7nB
QJxeR40Z9M7K4HNiHw4wqx18pYP/SsnDJmGadgBZuh5damyRO5iG7JPKf6D4RcwGGeURLueVW+bB
L+ZR/wWEaXQqa2cdkAl6BzCKly62bS1CeWli2qzPJz106tfWyNEq4B4dvku/lGp18KjswFN4iH6C
9ilMYBSuSQjxifm0KvN5FbUVAhtvf8D1iEbfMqrV7NzlqqjRthysEdIWuCPHtlluYMBUNHs008Pg
7zf2ghYbwXXX7hJmtlLR1TUthT98ZOVCi3VEiZaKTOrUtbUzHakvBUQ+ZKXtK3cIueLXxap8rI7s
1IPTYh7fLpgQPajKZmXzea9o1pBfuWP8CWqhQU/hPuHDHaXmJpJrB0NeFF2i294XQ7LZ7UyG3WMY
sQhFcVD7ZgVLclaNcHD7cdlPZNJImv7e5nULTOhFcyRySqiIDJ+U0CuAft1JFAQp3GrGP0Hlmmrq
lbok0ZJfmetTnSBQQqpAfyFAgVP3DHXM3ziwQ6lnZ3IyzzMrmWakA02TH6NrliI/VzAxcLqQVaXn
5ly7nYW9htpfgH4k942Et9amkSY8WjmBvpCVBCLnFiTJQcmIpENTDs0vl/+V3m5EhdmayaOYxuLs
FvYYRh8a7cA+tK1ccBuHfd72A9hRjXlb1VbHgYbDskBo1rTEpgfusNFCrakrC/HEmx3CQWdYhyhF
YGJvxAGIBx5EF3PJRiRJhGRqSy49maRsLsGCsQOpWh0JrIu4m1ujE4/D7qLiNoIundWyqYFuZKLY
7dy85YTO7eVLrsphwEQ434zMq2x8rIU6lwnnoq5geB75/l1PXVeNmC2CyI69qNS6MmFBzrtOHtoU
ZK5Axbxtm+WdOstnQtRBtk1Mq8HwCdogEjYMWyDcXjHErSiQHUCmzNGcSTKCY9D3f3paV2s2NGXW
BX4mvecEAaVwWADU2kilA1GGYXM5HyyQ1y832qmr5cHvpI8EXMYQgr6ZX4+gHjBZX+6QrAjoICPp
Y9m1sjFSbnswqb0FaasfL9SblWFZN0+/ZiubrcshygXNWdI2cYpG97urKVDMlt5iTJcODIjSyIjA
aYcvIMhII15TJDRXBW0i5gNQP/pqCAiakfzoBk4i+kFHnK1BcuOKfG8ksAdt/pVeg+Z3KabXhkkh
iJGKjj5vCUNQeMqJRx0Wt4AEZshCEhlWCTlV+HCuiQvKmPkILhqBn8ojfLc+QQcI9VpeiQlzmZHG
h0zRPzWWGHbwA9tvRbt8rNQORThl6T+rmcERjUsIKYJqOmwv4/0L9LKCDqNyN8g9EDdQKFjcUkSN
9eb3cE+XltwZDBno6tQhYbFjrJSFofhdQbD+CbDJ05EzFyhqMGM+FfzERCkbpQ1nAnA4h9iz6m0c
saJfwI30S3Gmxa4S7kyWC8ldPuR7673UPubyjI0Z/clQbSGx7rwiDYaXF9WXSby2s4cBdXNk6OV9
XMgzaoFUu+9Y3JnGlrxkIqGYIRqGkx56B8uX+FkAU1PHJU+xMRobXb8cQ2y8GDewTTvXOOeyNdCh
GyYumUlmLKrhlKGS47NrobhKBY0JgjFlXpuvTTw5q5C1c2R+eL7+VWwu1081E5ofY/0ogFPm56oH
cPL6G4TNG0dCBfgIv+mV2WUpblfpyIhu0WH6ASIgpjSjLR9ya/CnrSjrEwhwn/AofffUgejwYZ+B
2Hzeh+Hsv4+sVOWLZf35Tq6eMWhppaLkf2L4wnYS6OznJIVHY1vzbJDB3ORZJU4YYJDfZrw2Smd9
2SfUEnau7KzmBIIjYVJRL7pEMjrI0/ZQXgdd4tHHC09ROW1h30QXL5QYN0yfJnPoCwFQT4IZrzYI
U0fYKTMDfQPvqlK0Zh/FG6vr12+12uJXNs747EaH0B1IeWGABkckqccyg3oqOXk5GMCYvUErmNKE
dEWgiXDOz2RLIjkSw5opOEz00G53npnDaUUXBH8FeHKieNif7LKUvXtJiTymgcYzqtOWb+/WQ2sf
J3U/nOfin3ipoHSJYsomm/SmppW28FCoSJmoaCcF5JjlLwjj/cSkcAuLnnmPGxN9romgfpvs6fGy
0haXEIihDMre9EBA5O4IzIdUUVK/zaDgc5YxZP8dK7K9jO5arJEgclpgS4ylGkHfTYHbE+4lKUE6
L35fozZRCn/1TQX7UZVss+5wUW1KxShutoMJJjKJTDVAGGbqJ+kmMsbossau/gFXmeysqyPX1kXl
JNHmIFnNR1xk4l6d6uiYBzRt1rZeyRJNyCPrFmIUSiV6FxZdNEBwLNwI+/hLZbrlbxP8L2IDX8SJ
QKgkaMuuImwcvzqspIowJTJ184TBZ9O53Ktpz9bdMegkmyFQXUR0z8cop360MhVAUOgEJ+gp2XtM
v54pw3ln3GYNe6DCX94ddP7hUrO7DnlOvZ5pQzqB1UHv34f+bJzAoo6tuP9HA5gBfUZTgnwSEdD9
yi8ONpLYO0OBYP8iY1KWP4dIQWYHFz/qAiXz9SoE8v922gi880OKAw8fk7APZfpFH431slTsifrX
iRdfuiQoh3Mc3R/pfGIVJqJwq+3X2a3z8wGmMwk+gNSZr+0+U+qqW+zmNpjwQlmOVUAQ6lQT0JUS
JfPZKVrLTDMuT/NqUBLUNKHOr0NiDl5Re+/acrrxD9Sdfl6qamBflMgq2vExNZ6nJBZwuRTAtOqu
eByiO1jdNcRN0EtexEqUSEpTdBFW56TcV7ysLv3UuGveO+EQg7lFvLWKUYCNStomlGs8y5UPzp9v
5En3wrjsMk6MPdPuS+sgKzCo6tjOcaQAoPBWrqR+zEmiinju+9ZytM7+sWylI+EQAGw6JEke4QM8
a0w0gR+sUGUp8QueETqUByjh+mIZpwtyEHTklrhD9af67nQNprdsGLSJfneRJfTi95uHV/yujGW4
L2a66krO/Z3HTjwtZ26mrb4hhDGuegI2vxdd34UFijVlLHBodIJFIis6tFGyBqD6jAkNq00Zt/g2
r320Bssb73jtxnMRp4UmS0EmYx0EPRq/TTeLnjozPDAMqObNXP1Nyvj0QuXK+nFstIU31PazCmrt
EooB8n2+AMc1mx1rDApQ9Glu2PdPQ7IbX/CVg40LuXXHfKegR02CjmfL6ZBi3yxIfbJdZPpG+DZ9
Lw7hfv7NXWjDCvsLUTW7LtgaE2EAciQBvilQf9F/TmO20lBJPphZVR9FTRUZ/6Qn4dVuEIKpXqSQ
bWPhF5Ro7bi0QoiGl62pp+0+vIK5eyADUB5RqmxZwtEwrAh2FJSjYOEOln13iz+46JJoeeP5ff2V
+AAoUdXREm/VM9brGEXj5SAL1dL32WB3uxNaR+8xysCNq3uER7St4WdrJVHEb24uai7CI3bh8joe
xKLmQ0yNCPZOFdjU7gfcwVDkX7RMoFjkrWAZHzc5vfsCLxGAfpmk7Kz2TUtPHyUlcZrhbKEdQH/J
AjB1A9Opimp+9B7XEj5vh9h5C7WRAsmnK+k+lFWYJ9Duh1MisHnzzxxORfwyIBjFVHB/lcuysl6D
+IvZ0Xcf2Ey0sU7AcmguJcxdv2BwY2dJx0M/SAhvdAz1O7bufUuLZ9q9s2EvkG9VLOjOrvCLnBk4
PhIntDudaRzj6Nz+Zud/KD0jFyfuS1nNfRXIvMrErZ2JO6YkYM+d4ecZqXP3AJliCypVdXJZkMlP
7ceS081ghio5DyL14//1cxanSBRwFcMwDgYLNg11BmAXywpgsHDpXlzvGy1bGGxDthww9us2MmDu
bGEk0Ul8hu246v7Mrrju9QHpag93pEiL+RDRHyCaKzk0nl0Klphxh8BFHE4SOUMEEJHiSSgINJU8
QcLPMEw1L53pQKjqkQ9L/a8JzE7hT8/TsY9Lj41kenLRapME0EVxdTz+xTbCF9rf1m3SttIShTCS
NzpOqsC4xPHJXrUkGJVaM69u69Z7a5eVJ5dkRzfvX19jShy1gxQzjwgPNfgq2MmwpTRM8iFDSIHO
JvPYa0Bp9lwcvd9SuEF1z2fONLQEFix2z/mAZoFo8JB7qf1rhU/dtkrRxP9yrMiejFCcy81Be/fk
C+qKIbSIqX7wFeclUTd8ihqF7suggiKau1DLgGtka4y1iuLoliFONs7J4vJfQHDXLyLYa1RcxgF0
apYvmHx30qvHAL2T3fNeC47p3Ft66Re8iveNL4g8KrOJtkK66fjnVHVASnBS+hpy3kr08EwJyTYl
1fQCMvLHYn4XfeF/84aRzP65AIPOfejJgG/GuLr5WY7rq0m1rm3DhWyPH7rWNgqiz3Gk+lpopDQZ
RH80M9wn2oJpVdR1PWNXz6f96k5X7DgJj5xll8LkV/ZmeJfpgeqYot3kHa5jamgsue5r3TH42Ej6
8jGZ6V82Gqn80puFjQaUC6paJC1tjCUmvzRLmW6hoxOBZAPmty0F11WiJgl3Zej/b3q4EU7Z3egX
LuhtmRB22lKChAmgW2yjd6nYbU+0WgqD63rlq6lTQ/fqXoI2a19xaoQ0fvYJiw+qG51ivJR8ZqHr
tin27S/AOIS08O7W+nhJasGXusnZtpnu1ygGHMwMn7uwV+ZQX8miW7cYN4mA3pEVjmHJK4DAwW5K
VCOuU1Rv3fTrQSqj3kGJtV4dnq+puVp/+RLJbMl6oOsndDlHxF0qjgMrpzzvCekJ9gqQbWv5XV/H
wFbqX4sZGlobcjRavMGTb/eVshgn39myWhBu6t5GrW92GkvFoQQk3Jen2D9OCUJ1hxEXnyltFPyi
kvVUI3KbaeS/JC4IEssNndvqduZpDRsTJaOlpkNrOOzzBGH+AMn+hDma96Q4if2Rz+/vrSF26cIW
xNrhDtfL9HOPncaN5YluKlyu/qZ1SiDSmUIqkpX5qTmBOlyQFtEQID6ZGtxRGNMwbONnteqSOyq1
d/McVr6rdCsuSIh1Hir/+EgTJnoox6/wAPCJmRZ1HLNtUME5ozivti9S8pXbBwG3NwHK3LzXCZ9w
cJ3vwZuLhWJVjmNa5M094ouUyKxldCxbOQHYGX9r0ULZtW0dmjfifHsVb8U38E/2MdV/BUpJSCpI
e6OxYwmw+4bfzzQOkW+Xtjn6lxLTejKR5m2jsAdiMb/1Q9oLTO9zl/Zr3AxxM3P51eCJ79LqdkRQ
pymEr6COpY3UPm1GKWymopFFmBf1jTu0EvxBAPQhsxDPfudHLQ0C9CYA6eyzF5P3MU381U+8JVzf
g4Bba4hDRbKH/H9cFkY/quUkXw8i672KBBCBp9eSeWI8H07wtm/X30txJOY4HfzlEBRBim7YnqWo
Rt2TVx9+tpaGAj4jRa0Q+J8ex22TKuibn9Nt8gGzdDcwfH40GtGp8bh9S45Kq/e9yLLZfJywNgH5
ULHbLmQ2r20KgPNMEyh9IsGLsmCrUC7doNI0POHo7HSpb1sZfYmC9/1RvWmOEjG437/ZnSnlfHao
A887KPLvcD0Jod17FzbfPCgDdHOopi1Bwvtyvil2py05gXDq0IMU/aIBWr/Usm/Qpu9xEgQcWmyP
Lu2AaRB6vs/mpsRgSopWUIzNDhD0UHhXzJlK73h2HeLz6hyog8YmtXGpnNd0uY8PGIDCLGj7FEqz
3aOcTzatHkEkujtzrtdfzamkM6dsJpFylzFlDgmhSMIHVV4hmr3myIpnYVVGLrSwaSKSQsC+Rzci
A79HhsN1idXSpqnC1ioiXyV42eFXPw9qPIZhbAbfujpKPaCQveOC8o1DB0ynSloI0bQi7/TxcuJE
SQzkiUmgpfN5/y3OUdMPsl0JIN/0s/rA6nePhtBMI4JUIBXeas5uSB+F9ZFvZwC4ktT5M8OlvpCf
vEoMIUEXjXoaykMvNgxEM0Uq99UYSZBeMha3j2G2O+ht3T7fmD6AT8FcjCuLQtADSAZy+reo9ka7
tsxKShCPfhwaCtTvVz6RonTup5FLZnhhilKLTWWjmDm8fE+NCKW2CLFLBihGGeWx5uZYvhM47SHX
DzJ+hao3TRG2uEZDUSymRzxRuYAB3uC9irFo94NjLZnl1xsCUGS3RVmV8kPlkmOOKXcq4G/s5ZBx
aLI8ocBAWIH90cBylxqN6IDnt80JKD2T7mRECmIOFdzDdbAR95nsrHzUGkp3bn5e9ru3WcYi0kFl
tHbegPxkFYCjNlsVIqRU3qJYzrV/FwGzshaiVCJ0Ph4wnQMaGeQpmyNGSbbGPHLqgHMOuvb57iCT
e9O7oAMcDteEtS/JvnrLVbHEYfxDcbSvUVzKOS50fdNF0D8lMe5ONbLhFPkYInrwHs8y/zR+gm5q
cJNOdc1uHZIXdsPQGTqnATW7wr0GxU9qjcHPSQ/nEQgagspYUUs0jklz2LKLYBjGtUtvU9Uul33w
TpJERMTfXA2cmUhEdWqSGPVF64xTsOjntplOY6MaALgtYi3uCWDi9BiqnYTu5PQAAjw6lJq/OV54
vHwLOAtWzOfOK+Z59dqnzRolMZucnFGznsZWfrIrkY2v7+AIZElbrxxYkMc3oXruJ4pt069M1Riw
aEL1fmZJr8yNAPpLrKxLSurPmiBzgXiG0uQcVbEP90UgvJlXZUpMFCRlcYpL1W/a/A1KbfRaLx/T
TEY13tQuthLoUyKtpo5bvBda2zPQFHVnBC7W5h5Pcx/NIiU9D0yxDncMWgGbtDOq76sjS0KzGQzF
8zePwoLCfMsbVyRsVaaPvlA7a13uoMJnHlB3hntTkUAi4BddecwbxJ83kVQfJKt0lvUODzrgkaqf
+Q8SlIjt9NAGiXqAngPS0wdTeUOmjqzLL2My5QeAAUHdjxKbBEjojLsQfWaIBT2Rku2AN2+VCj8I
tqqAiBgsgxCtR7+nld6VvBnHH/+f15Xg/zLf+Et+1Bs7IYfEBEglBLs2Em9HD4yzpkjOBuIlr6I3
cocXKx6xhJfxZY9zX8RhIUOFiS+cLhWedOQpDKCKmbyAPrRC0WwHbhUPKnGxmnCb3OrhAr1C2X30
60e8gdQPLrd9kFcxXxfOSXFbvZwmcoq1lx2LzPJa5kTu3BsHIevH0mdg0vXmKroWQdsKsv3vDmqC
IzclOkiZer7lt7NsW7mHgNYH5owGuFGtpHyA9WyIHtfayavdGhF1vgXons/CpiOH8lJaGxSZ5nlM
V2zWmmUCu7UMN6mUphZqoCAhW2sziYlEYP/vnzUwfX+O9aMk1s0m5hSh3y6zv+yyX4faHVzW2vif
aR1KZmnIfDF7ugiifgOv8Mwmc3Ijh/At1NNysZZ437YT50UMLjHED5XyJN8Jy9rf9zPyIKVybJ9x
2VQo5hvkXnxzWR/JihFFSB4uJnw+uLaMOvL+5IeUzH14xTql3Yj9Nm2/PwimWz2wXqAbBHeNq574
/xU4dwDJdrYwecEU05garqxV1d9CyT+q6p2XDi2Edi8i1MtcIVYbIk7REgOqbeb4uCXYJYWidFYi
/Wmd8ivwwF0cvniZfcAv82FvUBqhSdOo7Xy5Cw5NLjLh/ESUIaUpE1vZOqpZ8HRqx7s/nQMMIdEC
5gWjvpaRaKi5VSUr8fASNsQf96PRWEA5E18pMhN1iB9UdQvqnvNCfFt8AKAv/jPvBlbt4aMX9iEc
pxhF7goQN5acGBCFFJiCR//0abQlYx3N3a2g/jBr/UUfA4t2qv924XsZzdsgyg70ROo66m3JNqj0
h8zCCrqrsgayfQWYOCcqBJQ+4pr+WG1Kd2wN5L2Xie7zjEZK2pDB550X0I1Pkg2bFnytg1RuFOM5
mtbPt3NYl9+9Fms1aQG2v+WZqyWjmhKEAHuzmA3zj2wQpY+6XFqv7XMuTSW3cwPB8/EAPGjLslVM
xS/YOQmYPPMD7JyD5TnmmXWqbblRsb5qPn2CsfdD0t2kFebyq7ovXDjZK1UmvPf97BahZWTMLhhF
gWpy5+QZ6HU6gCVCYlyNyhjjk4DH4jHLloO1ou6uKQk4k9EL3svK7VhH2mF34UvtAselR2IPULN3
9VlQUpdVVHYmbW2HMOW/P+27zaEdXpGYfbmRlsl8kG6ps+TXJvs9VDAWTu2e4li4GY4p+zKZ3zUq
AJCMYMl+4SBqWCuz+5pK4/NhnFY2NttGq+ikkQHadO3E+wWzqnU4lDW23EblIAVbaSaLEzKYIlPC
xa/MoU2pt/bcotV7e+O+I5YXvdYbeNqd60WDQi5A7JkcfxvKot3A3nBgdRqWoTgonzPtXYnM1KK4
z6tRMSBB5x11p/0WlIVH9cM8X44XVWWcmBDDiNwLwLuuV2yX+ildTMlSCq2HCgYNJwueHnPOvJGO
OmKB9NhkLegFu2MZ7eQzphkv5APrCLr40NFI8u4QfAvECj4ODW44H9P59H4UwsNqhORkrWeJrUq1
+j7wavPSX5odl9UhkE/giPgmxwcTsMEBnYuZwSzcz8cktMfjZJsizWHiWPJkIfvju/Lu40Cmf66h
3dBAYernv6ofzUdszmYvpjyP8sHuVg8kTVEDdARZB+1jOWyNjcI4wqYFbT9Omm53ueLD7i6but3a
eo9R4n3QlLumcukbvxDEw5OBkUXtjlfYFI75W9hIlrgmKS919IH+XMagB+x/8OfUhNQmlCHeO8ri
h3tXnwkOP88i+Bidi1zE0YGelxlQ7RkYuMC4MTWROxEM2bIVU9Kvao8PfUvN9SRyAlca7kmjs5E5
KnRPc9MVb0UUH0PN+C45A86AIEiSwAhHTNH1asqczugzP69aMUyM/aWEGXTjz5ZiVyzUPmmbDWz6
TCoA8wVBz8imiw5fCU8aVoNhr3oKmha6iAQSPHCZH0J0viTtjRw3DjueUe7cnApEuYzIpNGrmHHi
/p8iEVRG7Jv8Nsu1Ufoj7s/QCBJVO+mFZ5vYGhd1KZ1jZvSywsT5XcuzzTxJce6uRSnFJ0pZUMPB
aDEclPZUHOjXd7BIJuxOeAWJEzjadIUwjwFL9UfBerMXxrSFdS84WUE50El1OwR7XpsAY3JQSS18
1wnT4CrmAkY8qTT64K9Se2omp2+vWa5iS+dhFbMUSXU9X+EvpV2v0ZIgCuMuth+L5YhdVXUBfZLC
NOWYy2ACgEVqMNxjGj5jwQpMcC0nyd85T3rrRxZL9JoBO/vxybtHjU4+eg4h3f1xeq2e7tBjGEEh
t7gjG/+GFAHrf/77bb5lsYQxrxNAXX1pzUPSiYS5F0O5PzalAEzarG7pOxJbVndKmzTog289SJAe
E90ZGHni36ThTRaS50foVxPVaCLk3xdOJcrTe46qgr1Py2zYqV/GzzfN4UEj/e0F9MwcRHO98Len
bJ0F51KQsceb2UjPG9C5e/hf4OtOsFvWU/AseQr47DzsA80ZXFBag1P10X3vuopZmTIbdYAderMH
yb6DS/ggJbocJ/Blhn/qsqx+TMk2RTJbJBfJhBs5Fl/987wHe+vZvFBYYe0juPIFuQvPi175oO5j
1SOPdCNUaNKBbiCLDEztO70tivgWm2potBtki/0kWHBoVOMI8kxPI1D6+XjJ8CWhF/6QPfGbseZf
L7I7bqSbip2c2eW4VcXtSCEbk28PivH58xgQ+PgvsNIHCJk2ElfwqIc7hM//z3yJiqI99nOYcv7n
1FavioTWUmTBWorgkGy4tEjrKYQNkwWgTMj8eYY9OTxu6062hqadXDaF1hH2FPc51mLuaHh3ooxI
+Yxa7ur/5xqxrPMUuOpo60bovyyAMvdIPj2SMMHxwcZYcAopBjjIsFIb5foQ+Q+SUXsGJkFWv68x
ip7zQ67/dbQWXv/iEVCpQvcYUo/r+71uUFu/lizEM/tuVox5FUgxHp2e/WDraMWVJUvQnKksROcd
fArLbGprnLLN2s3pXUKhDwCg1iEwW/nfWS+Nhv7S/nh7W1YnswX52nZZVjJ4XmI5/MQJg6gv7pWO
BYgICTjBmeZAUvd0e1hYHBV3mgcqX45zDLo4pJ3ZTaN9HXT69wD/m1Z/CRJxwYn65077UjumPxWt
czd9aU9Qzr4iscopWAK9Ozf2QDL0m1xjl9STxDEiJx76Rfa8y/KM25TWCH1YkjPzemhbfV4xx6FK
seOHlg97nfNUy3q/b++wlIy2qJe9IOeHmpMxo252ri8/5tnmVOWpz/vJNbr/MFW2jgt7cnnAkqXS
kBu5opobbH8ZqfNBJ6BKKaL2QAmKix9SpMm6GBUEYmWFlpqTawpagpJntGL//fNJMZARsjeLhavZ
dJD5kLNLOj+t3OJKXtglKu6jaRsZhUVLssxbN0/uGg1qR5HGw7TTAWKbq/VixtGb8Eo2uLJ4Z4l1
AccYJAFnVDx6jCQXBdyuCnNyboFziqpVBymMTefmQX5jH5F2H/wSlNeKfhlmtCwvkcK9bbKz2S7k
kw1JLvpHIJHwjPkHtjYXUJnO35wGF8G8cBAD2+uJpB4DEc+Y5Kr8GHZcq0Ny1PbK+OM3EfEcSPac
Hyk5o/0dR1T/dNvFe9ZsY6DTiQ9XxuPb9w1a/ponAvhSoQKifq3t2hIytY2G5UOtZf/kz9FqoEcV
/+fxmZcyoBlOBlQoRtU9ytJlmbbePBxpSjWlMUsEcIsZ6iF+b5ffC1SMfHGPRgOrLXZGUFLXfgam
wP8Q6owbGXn+ujBWwlOP9vtzJQ7jmQpsGyVWlcRxIDIe2aGZCTovUmyS9a9flOn5dDpa3RNTUsIB
UQ46Ry6ZQwIR0dMvCccpcPM9n65YVuLJHfShGxpU7h00V2h4YqCysCkHmJjyvnFabAvNbhhFfSu5
nbvgzqbFJZk2p9+pIILVUqoX77v5NNxIE9iVB9sAJ+hByH6B3lQ/AxI1VlpWwFW/F/V2SfD48Hwk
OuXtsRl61PT6FkQM2Mr7ShsbTkQxlHfE9UkiLVDLOezH7azLau/hS7t5UkndoD9L8J9IFCzuH53O
0/JwQZUSr2KmOZdjIDrH7tAeezTKS4dSm+weaM/SZMKTy24s2y7Ew7U0TaIl6IXRrivR1OHOcxPY
ypo2F+Z/nbmQIyvgY9EpvYpVMe/qWINZUFD7B58mAgsVOzpLxSot7jc2QY0JonHAo1AAWLK7Gh30
/FZ1CsF7ur3xMA2TKDfSmTWEEWWTDYP986XyWRuLid5Bs2odXogchPY0QxMfRbVp4Gf9+DVG9BEQ
zS5nWy8xXZhNPg4f5NN1LP8vmuFeKpWqvaojYH+XjdxHCShJOuFSqDjHPMZfk2igB4trdM/1V5gl
pcjv8vdKCPynIgj6+WGydwIPxBg5GfyCYNoNjxaQMvwe7+A9lM/v/BqmTRhFpr2MxFUlKZho4mtj
FsdwxOcgQiwOh45AxVs8rJRc8Tr7bV4HRnSH9zNv8lh6a0Jf5+lJAjnxntrvYOVU5vY9sLJ1AVvp
a5Foqxg4quFaD0J72mEbTLY9wXQFnhZPe+6ipK5jICBsBfPgcJmlfQvkXI3nHytYEYWb55eMBoIK
/CuZ7bUpB7S92dyPtKrpA83l3bVq+9QOpCXEbaebhf49cqWcsYBG2Eqz5OKijQw8WsXthNV/pn3t
9f/+potOjIUALsmiMbBjpChjX5U8AcxhwTbD06llAuruUGUCNSLTOYQOm1aqTuuOkxkcH33BUI2W
VlS2XNj5w88z3MR6aD3Wze4NEh+wiTfrFo6KPuM1z4kBbsk73HZLS0ZLSoGH3aR0uU3jcv1u7s1H
uSjYYaXZtwGH0ZSHkCFAjb2aVNuQbH1z9dzv4mbah8v17CumMFc6rdu2Z11HF+henFiZBzmngWRR
7HBXfOH92k8qfRdiOHSLOeXufbbCGOFgW1dYyZgvGtteqpCE3M+a6ToJIXNSX9guuVu3sXgwbGnx
w4uigtO/U+9npB4Us4ibHYqnoIswwSC0TCZLvmiwK7yKG6Y6j00sN+iiQiWrfRaGGGBLrMhK5INh
JVKIOz4ozTvlSBbqOXfVYsgEDmhRWXbiA+46cDb0IT8V1ew8QOjQzV6srFecfxgFJq3+YcXFNvjf
Qp4ijkI0veZAd1hfG3I0ap3TkS9K7ieaPDc1hVJcKUnE850/PtOLzFU2VZhj573/ks10GaBIZe3/
i+EWBiY9KqJzyuj/jbzstSqE101SqdF5qK6ILULQ0v9c9p9qCmrzQ1AUTWNS6MBb6+5U9OfZthuC
+nloQe6eU4h4aZEucDJh6BltGcOBZu0MxCbxzpFM0WIBHQyMY5MDyxokJNjHQsjKQP/ci8zRcQYy
kG9YraSBiNNt78m36n28NN7wqJaE4weimgkljJ7TRJ3PfkPwgb9ggWfYyQcv5aE66ov/NL9xDXNo
fAF1munNzreAMfPOpKf8lG6/LK256EiPprokBWEGA2aZHTuM/3sb/0+MKofjEx/yt0+j72nlMoQg
zHEaEJT8gXiv4KxILtilkMurLj+MVhfd5CLLPAnTumhwpXCQqqJUK3x9wn1iQ9sZiwsUwydZsQvK
BuKBt5z44Evl+PjUJsYQmOO3DILA3aZoeiuE7Mm8r2nabVYhCn/rx/oPVDvdQ/lGQem1uTLEVQpD
HlqOpozQYMbn9dDA6+tLqew3APnYDFQ3ysUqerhVFhmc9ODZLd+/qoZPOt6yIp+FhgEMMNqkPBZ6
gBbfuHyiujqgOU3HEjx7cKc9HCB9X/4md3Yu+V1JKB8c4OG85pkwqIlYFSh0MInEQ8veHfMOTSWq
2DYzljN2evs/Twz+SgebNtzesIbTlp7mVqVqrlblPcRlVqxzsFrFaqr47jQ8a0aaNYIi5apOUfac
KjH4rojQFiAwvLmaPALTR+aX2lfWT80Y8Aij3qOogZwHRbVyRBvD9xEPWwHM6/2WTrFlO6CoZLsj
oVmf8AGDKhxBKDMPVMUHfJylEYlXLabnOZ0s09Y/Eni98yauQyHBZ4kb/GXoY1RdYIJj5tQUxIOK
M4tZvdc+V0Cc2NvagGxbOscG6qdTuIrgRmJp6axGh1XhsciS1oMM1LfiU7xpV+nq0XF1VfNSI9Ij
kjWmig5/erlfAO/zfJ+GIO5jih0KVH1/IDb3ExfbmsGAyqvqN0GwdKdwLOlUEcURnA5uXv3rkNMg
WpAkC1S2yxaFpG6tDEeYb6s6ZCsmthipghPlQ1iDVp5nGRqorii6E2QU1L/pcxMFhWC9L90FSCUu
LwP+ynNi3TmiJhWGBe5aRhESSpunetv/3XnsuEtLjYM+SGovT3eQCENLJAtF7QetG7l1N6aGWjTz
TJ0+qFr7R/MzaFcUrVRVXQQ9HXyuHx9W/0v2ZndxcRtfXMJT1Sw7kaffx/rN8C+gjv0x7CldooW5
hWwoYpXTd1a9MYXtNArbiF7nZmRMHE/SUJIrU/j/o608qQ99QeOF//ts7A0/0QhcviA1XksjKis1
9NlcT8VSfrVcXwxJd0646u76/f1cgOz57+U2NLboDA5Lsfsb3bRRT2w+cW7fHmypUdlZxQMuB1T/
K2WjxubnpAznIsQUdX6yJhmqu5OuHozCBkYCmMew/5YopvvbNjBB3kGKgHPDNP7PmTSIi9jbaMEP
f8ZMvB+/gAh0PGUbxcV2CXOEo/DfyUTwi3Htw9HnEp4dJxsU8TC2PmU0BFnKk71jGpU37K5frpxk
FNmhLdguDG1P3Uqj2zC631bDm9F8KUFNNnxZbG/LZDTR2rfu3Z64iLIT8EuQkv86hb7DUDP9DfwO
4r5gz8Eyex/QN1um27u/E+yXxVnlr8zHNpYONh2epDbP8ZyXgnlbgt3IIr4W57p60DYym6bml9QI
zi3e0kFjXmsm4Q7T7BAqIRvwuAzIMWiRIb9TYCKSsPF8jrUCAwvnMT7KzE8nAYgRqhMufDf1EYV2
XByaGwVWVq65HTfrZgZcgOoKPk9lbFf0WxKAEoUxUAk+UHZQz1kjYyP7gRHpAWyZZf9+FyrHgm6y
MCUHhbCplIaY+oKSskIBEj8ferq0hnPRtPmC0rJCwBpHazeyWHtoEV1SDcvP+tOpHiB4uoU0COWu
lNIPTB6WwSeBE722pqItZfeRB1m018WdlaJw4nAl46N9FRh8R30Y12ke08ix/ssIfoQ0+QmOxwpU
rLfmcKYD+D7B4/sOjQxkFs6K+QyV26iFMyPZftL7Y5c66keHDc9tmzynqhd5sFFS1geiyyS3Mq8a
G0EAwGKhAX9AQwo1HcK5ajKT2rzXKvHzY0nrzevsK+/aGj/1x1BozrPlKvszeyOfMMmgJvkJ0B+Y
IB4mLzMA3N9hj5dh0wIm/HacvubRPwt3GflYfSxzkWgJlLdwaDCV5ROVy77NdW4Ry41SdsP/CrcE
PiDq+SEPTUjsYXQtIFUKAMA+8E7kdovN8qpOjNzVzoELEU7v5A0vbCCDZZqcTMAS6DB4jHvFd1hG
LxLIGUxZj3COgJHlLVJ92JT2gu1bkmZJ4Aim8Ar+xM0rAb1damLeLYYZ0V/TnDBaDdZH7u7mlJpA
Wm6j2gAw2xVB6WwPLkxKKe/Pp2eNVwzzk9VrIw/4+LFHYGfY70k10at7XAdjHfnS+ga1IY+5QC46
ldue41iBI+GdiKMBwAJFzbEqFBLuFUvn6xWteF8o8Wu8Qppg+OvGk1AuQW0X4/ZWv8UaqaGOKJqm
2XQozi9zZUP2aoRlnVUwUJgJTE8CCidyYdhW4GFudvvk+A0sKt0mY1OObLhLMI/sgzA6nG3/AjqY
be4M4hCvrQ0bQmcDDjiKNAWQaAMcmjeBy3P7Acqf3/oQuw/De+C0Si4qMP8Q/U0ox0tdMCDaoKlp
dDPEMfSrPElQkMBh1bserMFZEXauaDkOF6ZjMxl8FAHwcVXjXR7eJulMnuYpzNH0GkDabImWBF0U
CtBVMB74s0mX7yvSaxuNQJYOwvLXrm7zhKE2i+1I1bZ78/Z4RAwHjaOnBeqRBg+ghcphB/KZGsyX
IhUTUuprIKCdNqaDiagWY/GvK38Y5tdFtVz21kC5sm25PH1vw8G1dvaxWWtWK73hHVW3Md+zUWpW
5iTF9knKaoZjPqVPNiZzpzquw89TY1Fjgbs7IBNyXd8D15wwKL/0VkkN9v4ac6b7td+eSqjyfog7
bft0J/bfBD213W/jPpzLNDuQrctRgV3XpMOgCuobd9ni4rQ/0DuGL26ibkSpfuOOvpJCuMAP5zKi
WDKn9vGqgXfzPcQbyv6Yl36/DfzR9vM+ZRxqyJ85Dw6riHilyw77TvWKX1lbzvkVFAKn5WKLjIY8
TDRKS4g/de4vtHyv2/uIcRMp0Efodm4R3TXad7k5RNzyJiL3/ylUpxfvignopSE3if80vnSNpPuM
iQsx1ZiwMaIOaz1kfDHOmM2Lwld8ue4PTEY291OE2dkF2eBME/OF6zh6On4A6Rz3hmbRuNCIWPkW
HGs0dqYHC4te7k0O6MlY6ccw/EtZkptnLzh3ov0rDHMqpbHPMxCWyOSZo3kKAO/cxCflqYzebLhT
myX59sreBATEutNw8Lbbi7YususJfGZFPph4q6jMNNr4PehmU1bnQyjRBLLsRbA/dxD3Bm+rGKPC
LMnqTwtYM4YSJASKshvWVnmyNaOHpRFmyTKQCM+s8+8QF/dHTMmazyCKC3wvaO1KWePJt1G2GZhh
br1AO9LYkaCCZBEFtXloya1TjZBFsN69hnKlN42ukt3ObH7IIZMUQC1/hS9+NYT/ZiJBCwE5/wln
D4pyGgKHLsbyd/Ykdefn2bu/vcqXbsgce2X7wAUSb6yDnoZ7h0zv6tuFlTou2hRhWVS+Tx9A4snu
iUL3mLvWffD+fOSAjDL7lL7pjUSFiz5VVH8T0V9/DdiK1pfun8Wj1cRR+geJ/6NaErKyd7pWmACm
YnLzQVqKYLbRFg8xvpnStoo0f2ltcoEyDPTHqra786EOn+UUXynNIKw6lBsBMJfMD7VksK1rXk3C
Fb8F0BUZnWhUZ0/nSdQXy/ctUkV/R6pIStQGZnf8+8Fd2zApCrYvjQTlKFPsKQuidG3B1rdDysAJ
oaTk8gOUTxUQb0iO+dftK+06GC+0+pifoJ5x/MLFJsDrEhDS9g1rvBJXiqxMKn/gFoubYu/wg031
kl1UOadlBGpWUEaz6k4rSsj8y1XHxw1AYB/zrNIMH7DHbGphR2RPZuP7tce4U2G6jZeb1uuiYGuO
RZ1rVdGzkI9v5auWdvpygIb8R5bscOoeixhKA7F3h7FHR9+Q1bQ5Lx8XEcToJvRPc1AQs8hwk2qf
GP4dpOIS+CzfW0tqclCCQt8QqLaZAGq2kvH6DdTDLkRzESTPVnHP2TFCiBlGGCl2x08d2Hc6LAGF
dSswe65BTU8LCbwFSnz0m3uYVhRD7hjRURCnAE8yFKBm2+1RIKolpidiGJNdLBsZZh0jyYXf+ojP
gMTeTldngH+nfKdJI9FG+FmHVUbpDTydpTJsh3NHi581Fk+rcyJEb/HzO6UsjU2EuMzHcfqQ6bbN
A9vp8nVHfXqSZirKZPuJ+HQGz53BuSEu8pSggXMXPpcr3TW8IkN/0bP9aB+BsSgBuLD9tUrpCiQL
qv5vHszMTVHIuwyfR6wqca32/M8UsN3I6xD8pwHEaGC+gj46wwnD2k4Il2wkaChPzYjJdadgiOxl
aL/z2kV/Rf4hSwFXVxU7H00I7U/VSI9yoO3A2Q8JkRpp55Mb35dL8fYjPLx0JuTsXjgWsCw3mgN1
2j82key4GUomRNB9D7RRcAurpooWPXdtjdxzsO3kV9Dlu/ziOTkhP8hXJSh0XKCzLuOcbld77J2R
2SQmSQ2ln+/1Npe7CTJAgPPVevk+n5iDbhsEoGUK/UwAVB0w7Oa/PFiG5FgKWGtG00O3bHQlmX70
oOl1x1dmEGQJA4bbikurCwj87y6vUaEKOurZkXOeDoHIrBUAfXyahajyjpaid42R1D//prTluK2n
LlkIiDebkLFw6Ku2cvTeUZG14ErS8ZLcX8oKi1a6gXZDvlGHBR9E/pV5NsIBH+h7qCft8mkwvqFR
k8zMYD6G4JHf33rvk9e5aarQvhSGJVTWlbZtDNCtC38LAOIKC7rfxRwbDyG0v1EunvxcRRQBNk97
3oBPfxzfYTL2bGXaa/Qdtm+7Ehg3jdzl571KhXywVnXn3P681ENCvbnAINNeVX8H4Y5q4KJi4LPf
uoz38iDh9O6ozKFjxIPz1e09ph9or93kx6oEss6lM1miaEWoiWN1w6SGJWBL6TsZ2NlfFKpMxao9
RciGZdsn79+7AxtiRrNxBh4tCmrENfCeeJ4lbciKaQIZL3y7aj/Fvz1mIjCZP4OleezuF8HGJvrQ
vggWhqabYlh0unt6AK9ESLXiKGzWXQgjbjz6pxA5yzShsxnQOfP3DFpfiS+o2vqPPC9SzGot56qY
d772muR2NTKG4Fg5prH+usphe0Gv5R+FVOicUaYuyO53jjJ7I3tNBmJs02fA17ftHjFJQFrgtCu6
w8JuA3JdfR5vmJKDY6q1d4RB/ZcgpKHDhBrmKC+cleP8JPpW/KDVCFRGqRJJZS4gE/5Ygt5AgdEW
2vTOUcrJQ0p/mdk707bV02FQmErCqySIpySSmQ2g1/89VpFVY4CkGv9QzOcSXHd+Lw/ikRBiAQly
9d+DevV8ScGlgUorz4omzuyGVebdfkshMggslL7J/WebE1J9IIreAV6QlqShiurFfw07AEZ3IQOi
yzHdV3Mhj9a7sO0y+a+huNElZA4Tep4UoT5lqiOUlVz4g4fwKndlTKqTa6sGnXVIh4gaugDZUDs6
ym9Dv7qHDlOJ5i6dZDekc1SFAmS9/bWj9tsmiCEkxY+MyJ7lwJDYlO+8yDYK0EuPyI+x4+xXDTCr
Y2iQmYI8sNBt9ckVT4qrNZRh3XaWy3yYFV56LqORfBiRg1B7NjADLO2AmMzbLmD53R+iN7yvv5X8
HOK8yHcRpGTjD/qXaCzz9wVAsWXgRAIvuEmjLDi0iml9ERhKFxt9EqLkH/elUItQQ2H2NvxF3c5k
4cNSAl4C1ntJhg1DzO76zlKrBb3N8F+a5SkfHfzSTPZdIREM0QAPkRS5ENW4/Jb+tOwfdTOFHQKv
hPBjuuHwW1YM25rOPvEXWfGC6T9dZ3gcpzbuzTnbSRMBcWM3gkkqJ9Y6/7MpZf2ju8xeJ5U0PhdU
yKC2sgv+bFy43agDehrDfjPinWzVpGjmPG+KwHkbykPyvewUZrJXKbJfPe/0ePs0t+ecVgu9I35s
3lrPN6FYUwDRYs45DU0mJ5diMmp3Sz2f2/jnfl3pIlHyGPksJ279juv7muiO05CizGQjeRQwxaU+
asPceL48XgHsOXGZSysYqE/sX9j0TZU4Q72KxLaRKyUgztvstvlpKAcWR3Hy7h9rkVOPhn54Cz92
hWKOetZ1j70nVIUBbMO8GAUovUP/qCg/WJ0dk/7b5g15b5g0zFx6VEuDGifohdDmwqZsLQnMwgif
DbCTQVAsYecOamDUSy+7yrQQz26YPDB14FgWXyMAAYkfsJzst1d/J3r5p2lmMTzxkhDUIyxf1c9Y
3/SAMQ5vwQl03O5qPVjWudguvL3aik8GbEUb9EJpGALfoYBgkxWNJMFySNNhrGEtb88NJx+I8JTb
OZbfw10WL/g+g1EDYvm6hyd/83W5Pr290xPBVMtYjh4tIio9Eo/9AqNaOTCkE7l0SOaxSG75+ROW
Q3qB7oguqfM0N1SNsqKFzDkhzlWnbB6B/XkPZ9EeeGbEHxbC3RY7QRHG0qOQDcnF3ZEM79YZH+kY
t8SrZsNddlwpYDaQdzSZI5pTVokVNqe6EeG8WhL2U+6si28UvWe47Vgn3AGwhfk3WE5StwZYo5Tj
LIQ4qPTEEVkGy7DQ5RzZsbiY6wfUN9X6KOOLIbgIA6XGkmUvYMmPvo1jb9GIOCI2B3Q9Bb1ZyqEa
RwCDl31guzkZPCy/Z//HL/pwW8AN/sDRS+a4P+X9WJnfHPgG0QXD7GM47HnJh/Ks9Q2g2rHl4XP6
4zb7xPmPhXb7PITyDGS1DcpXm5v5N79Ue7d/58po8dPE900Q2DMxqlFN5puOLq1MeOyLf51eXcTs
OqqHKbMAbTYut2ak/454Ay64T4WO6MR3RgT+bFBHCPIexwr9RXzARvTyawRQjiAdfgR2NuLcw/Fb
0q30dOk+XfAXzXfiYxxr9wserCk8o65S9/IDRsir67usVz3MDDJPKffih1uJZDTBG/y0Fdh8MFlO
UZrcsKaqIxtFHhjrYvq4OYYZfeG4ywaZZP9EnzAoVRIu4BZZqJ4OCRxSRoFQjU68B30qAnCQREQn
OSQoOgkCA/Fwb2gFBMOJbQAg1ZyGrBu10IJXwEg7ebVe1GqFrYnmEvrQgcbe89TcLsWr+oqhYyZV
9O+MiuaGqsHW60JAOsEhDv68+gNWCE11CKyWyK2PJgGipA4jXcYrqobMZYh2pa4Qo7dO8Ww/RTC5
TkFw1Nk3L9lvug0SJZsll0pzAy+cvOnC3w7PhICkQZ/u3cjXWzfDmgcx1BG760/4BERJXzxo0Let
vEAUqPhuDf4e0sN1SMuHAkdBSnq1gFuU58ezudkvqh/AJSfHYXyku43J5BxZPQVmH7pYUMv5Y1hy
lJuHpRZNc2k4zjhvpqe6zSoFegONKbf3YXGV6GiH6lFnJY9hLyChRt8pGKLesNJIYBv7O3+z+Z6B
1hJT65ISj0v5oNpHFeymtfdi61LGQVXvl6Ep0X8iLTDeX+aoYtU3G0QwzBYF4OVpRK2W8yolZ3U1
mdNF1Yy2+K0XhBpz0PCAux57jvc3ByC6ua1mmVZ2UuOTIKmwTSgMF8roq5hTpopsfRnxapRGI3ei
Wp2jDNfK7VlqG/tYBUGqfXDFubpjfhQ8gCD/RMNAhz65B5jziC/qzCKRWeZn0K8X37wRUzPNRuFi
mQ/eQb6Nzyo1Up5oYmxNKbsRabui5H3fbEBbwbt+9s95QNBW9OZ2VrlpAYKb6RbQ9IWw6hnAMXJD
Kx2PxcIE/BFoFySIZ0Ibo22B5nCEAj8TdfUm0EN0n8Ug0xCrKChQhTjf2IuYqxe++tCWnVjqi4xd
ZrqFIIOPDARCT3iSsyad43gufZG5UUbgHFWxKdQt3yyUa6qIA/40LWWcCOYkYLFGtUmN0zVgJoph
H6dhi2n4Qj5rJ3dL0UkJ+hDSmK3tXJb3pU83XPKEiLvo1P0LkeIdSx0iqLHSvOMGpkAN8TMc85Ew
g/ETv7jIsSoQtKWb6cHDHocoe9Z8aUqEwQiCt3VjE8yaHGMbmpecEyOa1na30sPO06W/QPb+HeRj
KYy1kfItahqv/XyjHCSrPddeV2B/TQO1ulhI3oGWmwyAP+CjTKMFwtTfeZmH2A7Dlw4b6ejgnqSf
aqv17t8jUpix8YlvfqUBzJr22eZt1txKHMO6NbzR+Xrjbu7xlCsc3OTLZMIxYSK16UjlWSS9xTUW
DpRNG8ZYaEdn3iP36zX+1M/eD1q8gWts2TQ9SKPjN5aiNk1oGv+TYdyRuYSjjBkgUms5qP29P93f
DIS96lRuVu9bYNH3eK6EdZwydgHVEmJh7l0IDK+Ea73TiMnqshRpGti3Ju7YG2Ou/EjV2O1jWVn7
mrpIAvljVJdq31E2ZdE+WMAtz6ygqBaDd0/KVCF69cO+aTKVi10pMlkNSSFG8saVOuEraPXX3E7r
cFSqaAxG6N96bkQfTA01dZ4tS4EmJ85otIpIiRuhE/QPpITOEQ5jm2oVjvZZuJ8YrLfW7o4niFvD
9IWg3PR+YHhLDEkldb1yQiKHKbjOFarEQL4QV1ninDusJxIciikt3P8PI2lE513xG+11k36byQ0Z
xPn0xpcg31jR0jW0JobZW5Qyu0Ns4z6kZA72Idqg4xOYsgRm+Xz+T9qTDdm0u4g9+hr+UY0ZmP1L
2o5ZjmrYfX/IumRFd2+KsfIk9Tb4DE1YzawQv5rW2KEYfZNijxgR3b3+YqCN9Bui78zm9A1FttR4
nI9GsAjpuyEsSFrTCQbpy56zXuw16wACpg/r6uGfvsAJSjFQhvXLMLFfk2hpLVteR2F8eKF442Hx
KdUbeJu2J306eqYLJ2k6CyEU3va5yeSJKB0NBQ+qAkF87E4hB01JYT5tqbBioCp0VXSc6W3Ni0Wv
FqRvmhUI+LjMe033vqLgxmqBq800MPD6QYCQuhCvGw6/a0tWhLuXTHO2TBcU7mC3DjKbUEPqKMXJ
vGLTuhDf1Fi3ox7uU9wsr3GEVdGu58/zcK1FV4JbeaUwwhtvJWcy6lYiCVU2MBq6gyih/n7M1GMz
+SwKlYlSrSSy/DGkV1Pd664ETw8KyNsb2ONrzfc7GUwusmoIyjKeaQi9SZ3Q+GNa1Lb5p+lYRDUO
g6rvQEmiOhFlMvCVSsGWaVmho8l7XyFNVNUmxk02hlOe9mGgVtql9ZvjbDkGgdJcCeN3iy1aa7dL
i+f+AyHUqjTjV+MwJTFLoOEyyncN2KPJMyaNV0GaiF9lF0mYznmfw7dIUhFptT56jn49yslkpPym
7Yj5/y3UXRZ2jROATb8i5pUeUd5E3G551GdlxPyFN54JhzH8w+e3vL/Q1g1Yfifj3vi3tLzUHGlJ
Ta8C1eAKzV0BzFdc5Qr4HxNtzd27CkAdGpD7cUOf0j1dejtkN4jiffhQb/ObJFjUjlJ3iG1t1Vh5
N/5R3npvnVKcyapDYPZGGvlHVUBfrhKvKJy1Vq8hJZU3+pM2/ZYCC9c7F6DAml/6yMlOTAfJd1HZ
L78cC/R26WGlTE0bihEwF8aMQ9kczZSIg8SxPBAmjXn/JjMnqlRmakwrgq/YZYDA96aoTxGO9djs
UGj11wvGHPLswtffrNaLaHIsg3scEsGvFQcc1We2pk6aeTQbgle7XCVGG2hiuEvtxZW1YAmmVwLv
iN/vsYrusBsZ9PmnMvtwmHssz0dSR4yfnZrrErE36x4qZJdcZUQugJhuQvECsZtTgMVvJZ8IbWLV
efbhk9oHsr5MEk+aIXmKEnlA5D1su8S2QHRIiJTHc533sEQR5wGj785nePsn5+zQ7L1DMpnYK5oi
1Z0vmfsfjzMI5yf8y5QwzfB84FK0/wS7+RQItnwrEbRuMQMs2RQfLgttZgapsMFzybz025Cq76YF
k/sasVEtJPGG1IRIU03+SS0fHjZm8tunBT04uht50nHgNlW61NVLt1GquqfViL+mVp2AGlBVXOe4
dOzvCflQahmrXKafFLWUdQgbMhUeOAJAjBOOX96mME6vea6J1cHZgI2rKp1isKJyRQAcenoAmFeg
ssgCdwzvfmHbjQPt23Zw0w1GgVoeCoMTwCXWq/Ok6Ht8r9Hd4MfxDlEeP5UglZkq4jN57HQYw4QT
8s9ZDNOv6bFw8AOY1J27NOTfdRaUFVWY+fFCuJl6FuC4Yh34NhiJgikScDPkQ83Zz9UdUulXH9MJ
m8x/3xX907RX+/uGDMXhoplL65ViXbL2ExnXxyxWXt5WCGCfynczLaGRGdHALgk9AC2pE8Brqpra
v/zgM7KcKgeqGdK7G0gIaumULm2TrjCPawIWQJCso4iUvixrdtRuKvNHsDf9SE2dKNTUcvnsdMI4
OLI2b/Hkzoq8dTySsM4RMc0UJRgfyw89Zv/x2p7wp3+tYQmUDN5nq8cc4yMEOTy4eB0IF3EOPTKf
jPRFksF2kL/muyG/ZLTItSIrAEEimd4YQz9aHFjsIkQ12hPc9qBqSKLzM2Y8BRv6Xyg1lKD5XskL
p1/2wVbC+4KXmPV0A4gqJps+OdSCp6zrxt4SGAx9CUukEeGsrc6rrN95Wanuv7YqXa+lWhe19uxz
vTwO50S7RoodmhqMm39kufWy0VmnBrgiNHOKqOnyJiCYIE6wpGGApqy6XClAw1A3KELWn9vLcZOy
/PrAt9sil9xVUGr7eNdW7fxjc+il1POgWkhX+n08AHQis4VsdJcY/Wx7OPLIIzv7PpEMoJUhj8J0
9N7VTQ5j9vTXS09ISAVlca69CWdcUQDijMvSi/hW48RKxIJNYvXtVqw9hqfBUv8gdPHJL7Fhsk//
S6CyauIr8NY0gy8SfWq3YLmq13jEjQpGeB1Io7FkSqxmkOGg96YWPYbEJCTV9pndDMb+HtIQI5nz
uDg5FxJ8QWbHVsofHJIWUcnRMYvcTk9NyhZ+CngX1CaKYjhyX4eHEHc71XCBEDtx385fgvY7jIhP
Odf9J9vXY2knEFb5lanTAbWHN9hBtwJo7+g1ER6XXUrw0imXRrYOdEe5VoHysYQZAE9s69LOEcd1
nIeUBKAs8+UIlucgRqXaupKZNShIWyUq1wk0dAUs4a0KR2qjIVPVw5WzEnJF0EKJwI0lEq2mqfVw
ITM/yOviywcVSFWpBIoPmYJLzyaz0nI+EmGXM2ihLahpU/AJ9uGXNuhmjmKKEDl0ouPSmkKTCZNF
j2L5bp7CQv4t7PAY7xcpfagiG2IePalQohyFpcUBJQdPbZDdE4iBfqEKKB4ElZhTAlZPLDE1UCyQ
j4UueSNDGohIrqQqGwdeSd1vGqKHKvwIb8cKuSKnN1NALG0omXL8tXC9gLsWzppbCIMmsf7ci9EO
Vn14+HxVAJ115lpH7S+FPFA6/6v9bywYevQtYXnaboNgfr917NQ6GLk1iCiKJbUZANG0cJKfL6tM
KFvKirNIgbjSBMDB1/VqiUlfS6oE3P90osymTtVRypT6pfVTKFeO0zs1r8XxgkRCwQD9nqACO+WK
FkzAIALV9cxghhCmGV3nKHwQ0kHqkGMjFvuecBgWO9zyTNgbgj/pDB+Yyi9EhKv4AhXmqp22EEO1
pScuUwAM01u/h5kdzdQofKw/Pj1xgPni/Zmt8ql3wfLlPHtd9UQeo/5E1ZWcNv9N4akBH5ISijRZ
8Ahl+nZNwLyGSLO5t6FPfnu7kOb5twnfuM/K4Pyn3FAHfWVavMUPaa0Rup6HXAWdssP1zXGDD649
vI1VMfMAqB/lAH54wY+CLfJAmrM8LXeFff4kOtb6kH9b7f7dIdIPK80pEY8gFApjjivPrqVwgsU9
eJUabJqtO7KEzdOy0W1hSeOPXRiATR1G6x4ZuSRxZk2YOY/HjXsiyzqqt2iwguQ5ADN3jpUUcFxN
1tKK5D1wSW6kYkm5npV9Z3h/6BjA4W10A1nTB2A/OMwtYzehfIwa/ttAR4Y9auoE/xvAYXCyYIJR
e/8jjQbZ4B/BJN3qkysl7fbo/MBiokvVDhTwzUk+VHh9zw0RwdF9nwkTPUxpsRLQq2/V1S6UnKXC
K5r1cdIJofG+H56dF2GsTucLFhqWv6RJSwq2TByJ7R4RBqgaSBFMBco6/Oh49482zXe1IxH4WRw2
lwxVW2nTpJ6g5WldYAkINMncJyzbPubOarYkxnyWkn1Or8nUr9mY9tgXRNaf3GB/mj2jSl6cU2Nw
ffKHuvrUJzijz932Rewx+3vD5EY7f7YYpajl2WoDq4BX2AH1gHzhnwVewvognbofgHshQ/bBQLTX
6ChchEU5TGSnDi+Cc7HP1bOnm7j1SfSNHsl3z3zh4c9K1qAh0np2UcaBS/pMWQwFwruC2+E/0fY2
UIQOwlOlQm2GD6YLnm0/a5uihJKEOfyvJ9meeuFXzoQSjPvI/id84gb4JI2IZ6APC1kF96jx3cVR
DmwimsmmRMlGDYtdjT1ppC3ZMG3UF494WOp0HuO1Qy3bej958zgfyfLgocZBu802wFop25vE4y2P
MRMWx1aUyRVL8tkSqm6XUGkpkfHgSzfQjWr6Jqdav+DHqxRVcGDK77OWVQuYuAcPSLl/xVn57wrN
Rrr71pDtoRlT2Fq6RJlbOZ71enLAnA5eLek+49R6jDk+Oik5WUOTLNwtkjuCwLwEEKtoIGloQAI7
kvhhscuQIfq8bTo0Vfx1iU6ZRiPTlDuyxjfa/ikySArcY3Fwgsk6ksodTP41Eub3x4ofaQuc36So
iYm+JRc9AiC6JatkUkpb8d71JsFJ30BB5iP38K2BWZn7HVdeO5y9QrSHr8eJqABA8qTnjXYiR3io
CPA+zwZvaifYfHVVZZWU1ICJnmObuaH3zQJyuIVGf2YLvdQ9Wqmv425+/d9HttdX2l+uJBERLfa+
4pC3NFROym4vNZMUlOFiehjG1fnFj/ZOc2m+8en/Gx4Glg7Y0kpLSRr48M6EDCPe+v/3m/i14UoG
TlA7y2YgFFQvXErUngeLKGSnCwrnxQf1hNX+sA/Qfhzhm2E95XTwrjEVrgxYrQL7MeByQFzXr94L
jZaPcGq2sONlBfEUF9amd5cmoZiGywb6KdUxSHZ1JoE+xGH2YJZKkAO7c8NFJpJwquQ8gTVb4zA2
2QzT0z6cDYzwr8ALtWIzmp3XqskGlL3br0YeAPRn3mD5VyeJ+OhsFixp9zzlfdT8I7KdpdTNle2P
JkYhIQWatHgu3Z8k6/XdKumX4kirapKwncA+/Iop0dWxV8wtzPgAkrV51Uk/1soaDZSOfCJWsF/G
WkMXHo8fjsi9LBIg8yXNhYHMgUMNhltOOm8fwHHDTfBYH4Xm/vQQKzSy0fRIWmYTsPVXCeUVzvbt
r7p49A5zpeex7x1sPjOlXm5eRoQYvdkfar2bZLdYB2YrSNyu/bLywDqQokfwK1z3y/zDTFRIhYDr
7tEJ2MOlEOSkOesMNXMKlv/O/AkT8Eb4+UZKT+LXm0v6LOKsPZiOi/KVBUtPAWyiCExk+8EIzZpS
M7iVRNieE4Rlq8DesT7NYkO+R5osM/ZZGSBb7B2pFQm5Cc8qN8t0vK8+0PSJxq9KLq5l5nf8s+Fj
PvvHpjGON2mp+VbDUn8/7/IGxN0I4qyPOCePAqjYC2ocd0M8cwdqGHuyrOxHSNpMAAhlbLP4Ojbs
YtMhPI2PQaLV82xRV5h/6SqsMBINo6515hrJID6Xbiz5KWwjPrXO4Ea8Y8sMk/Hz8Fm4EjfSHxxw
LsPJKGUudTQBnQtW9M2tf0TeZSNvpUYdvfgBrX25xN0dRrdV4MlZC47kWWsd+C6fCKkfVfBdIstA
59XC9G0J/W0OiuNG85yzcGwR6yLbEsAZeq9Q5yKzuAMvvFKdCfxc8rgL6B4jPwN3WubL7NkTNdbH
Wk1yE3u36qy+ujQAV7V1s7HrhkegI+L1bvnZw9hgAmlx+6cOLr2RWT3wZxhHbis3DvC/8Ygo+ISr
/RVzASoTir4iV676QH9jhERjcgCXv/haMea1xSin+Q3ie7WgeFOTWvV8cVF5OSHeCIGfVwHOsEj5
6LYFnKsR+0HJvi4MfscuwIRxTIiIXEUnyzix3OoR7YOj6OJMgZpi4yr+TkV2ZbLIMdOGKeeY0jiz
5q/fwXOpYvN3oJh78jPVju/f94Ry36l4QeSXZqpwOUMCMRYI6mMuHrwU6gfnLQgd/BCqFa8fOpv6
wYJqoc43CeQg/cJU9TjdYlHOCBdPWU/owtZIAB8tDhb3sufwoqbf2ciLejo3P+SvohfGHw3F+l/I
RA0/GYlhgwEn3Hfu1xt+TfHibx/xD7AolHAt41yKYTSBypQuCuG4Jtsf1pKsKMDWq+C8lbmKc2UC
/oYHNWZ2TpZt2fxu0zwmXkfBeidlP7abaZ7b2gu5fP1W+rqZ5B2HHJ6xz/uJkzL+iURv8idlsgTs
JV2dWnJObw812peaJ2bB8gyHqmp57Icdip+4FT4x97kIXoVGnHLV5583NFmmsJHk2k7Y89u8ulZw
rbxwUqY20D+BUDAkd/Muzp5m/s83MVp5nunZdbPA60qVDMARiUykBNvv5qgqXFveLwt0b46PkwZ4
O9w9NwSXZngLlCUfIdPUhUpBea6FncKlqjhYnn/H6QICrvIp1usuqdRukRKiqZgnKowWyZv+7vCh
fPOgExGzgX1H4jJnMO9t/bPpwM4DyW2uBBB9aDvWn86jwIVJY1ojwiiZfvFvtBsBmwTzFeZ8XcXF
YewfyzjSjaCVOMXsEnLgTk3KJv1xpeBdFyVD2kRAMCsKt/EqIiYhS2pnLMnTVIbO6wjQMMVmnuUe
7RW5Uzq1la2AFr7ASFFxb6iW+Jp/OX2vWxM/ScTO7eYXJELnSixGvsYgaXgyCRNBsaSfe4iikDi1
rXqUi3SNsv9OBULIj51R1s0wMn5j8Y+f/XLGaZ2SmXTQxRYp2XG52vbilRJBiDYQmdM9Z50RHR18
WM99agO9bzMMGornYityIxuOZZnSPnLTyCVFk86EAQB6/PaVNpdy1oOotyNHqJCr52iP/c69BMIJ
SKS1F+BG2vz0tvDN9XrllLxy8bYexP0UemP05kYkuE/BhdtEi/1cnthi/6PjTs/rswcmNAWxAxf0
cLSc+qCzzq2YAc1oeN0fjIsjHMMmiAmYijhWFUgoaY531zgluprtvLhdNGusFOksUZTUmmH2CuEs
6R7IHsoP6guJhagqtIk/Xr5xIzpR9Y1NBz2qJRa+c9HpYotAjrIa70mqVrbwf3HRoKgllwbvEKLp
pH8dpKgSYeD0JmnY8OVHpAX4dC69e7ur0sDQJ4rbejmjTkEC92jIsPwWISrmeBdWP3x0xJjzMsOz
5zLK7oOn4iXwqGuiectRcSd4f057BlpAO4N0jM0UHjUU4R3g3bTMmNXKPdXkqRROc6K4g9y7uNsE
7hrdmHQKNN4QlwvowPmVdvahWU/woDZdKVsYCCkf0193tWgQYTNCTe/+2v7ux2VZZ1uiwFGEacJ+
rydMZxRzWblEIOeZamLS2eMKlLlhFpSLilKzytfXCYkxs7wpFXDqVm3ExVmmxg+d/kvgPxqd9oyP
aQ3FyiJAGfl+VEwHZpKZaOJEngl76lWSw45wmZy6Zkl14T1PFU7sIidxjNJLrVYcWISRw95KIMXG
PwpgSFCytimzq8ziPCSAwtgz4eJxmxkRp0+NihiVVWRyXgS07xV6slDc8l0uumvtEGW0cfE9BZsX
J6HFi5PViglE0g7v5xA6zyUgwlIjELH89EptkyMZ9ulRnShmEEwJYtUCRf028pzXay0pFRiBhJON
C2MogxqFB+BMLBGgd92cgjppFVD7qsDAJZ1JY6ci9oP6csgOz+PgSHUOmrrMBWalY3W/OFPzFoMR
FSAYc5+iPT4YfTH03G7x88hAn6t8YyrwM3P34ELdUp0qQyMLUbDR+xontuv7WDcCHilPmS1LlCF+
EqtxFmMjc70qyGW83q4LSjkHBKKNUlgW0q4WhRGHz4UYAFfqZexwFJBnfmzFL9lVTU8/sksCEeVZ
nesU5n6qN0nbpzUFGpGi2pAoR0eGMV97TX0oFdMy84ZgP3Id03+97u28M45/raDPh9wFiBdg1MKj
UcaQW5U21urJXtrytpgjxqQq3BvyJGRofWHlf4nDtkRiHklNdGB5dX8hW92j4woLLXRuM5UM9pBd
tA+mnLqTn2mkYM5N8d8jLm8YbKrpeo6jmIPidmq/mHWoy4TnapNTdaIWb8RDD4oD4lOfBbVh8J6K
j4wlx7QNOc7aMjeNxG4naXMkW2FCzYLgptDBc6Rm9GKU9QEqAAAqRaMQX2HuqyLsYWqHMZbXEmSM
4gmrKQKbdHC272YIc09Mo7uSgGg3b/kqDfLWNsP84gouQLhk37bKkTcEaUUBeOgSvJkxTfbxB5YE
tB88a2ysJIv9rRNV1dcRzufKehe38J5QmKCr3zLEVLM0biyyg/5BDmlb0PPptXTEP2zCAIbRQ4hY
V1+VRpIMuIYncpeNeksbkwjHNssWh32yx1aIRb1Zfd8/PUPZOcva+QUtWPIaU6KT9VP5ejw6xotz
rrtpAMzzT98lgGZ7sgNDjNdO1alwUENRu6ayYwdYqWlht7ctP5FwZaIsML4a7lljXw6kShjpyy54
jLIHvual08LZeSI3nEBLBGUbZbHaeWxFrBx3kklMKK0AP8iQEo9lTCl2+Z1wHl45pY+eXWR9BKrs
ucVWlDxdeuTYsVKtgXt6lpS/lCX05gR9nKfWFWoNLzn0R4K2sPG8VwnsYZlFJx2sBxz4L8V7bUVK
EKb68ST8uioSXO5RztLG51LTNcxBhG0KTR6J/97DlmFdKV6pmLS2WuX1Es+mMs8C4BWGJyLWQ7TO
aaSmeuTMUm8aflkZzVfUl83ZUHSrie4wIODHS0RETLTSPeFpVKLeeeW+djWK2D88ygrwl5Ds39Th
9a/t/9apcydobvDsVQZoPYMDeGjQHxchBzqYxzLJsXzMtbxHZ790ykpnKSZS6k3eZc8IVLgfW8KT
e06fk2uVCiiyVs+TAt7+PhYlTuooD1zbbhIqfLE9LZGK5Xp18PB33pTSM92TXpwE13mfQZ9rD/rP
xeQ1I4bmjbQLobok6yBaSI1XgmAoH0bxXbpy5FXHa4uBLhvP3p1ETEYpgYt9cAw05xXFU65w58UE
CeXjPdzcQHs9qxVEzpa31PA66dCiNXUElRaevxY8JKsOidUHsW5Cz8j9wTCtzaTFh3wFDDRzmWYZ
w57d4FkFJcr6OK2BKnfRGC5LLB0Cci1XAm2zBzyjCHCmwXuaqEQaVNr/p/eJpokHqpqniAQ1U+n+
nNjEdhZBO8c0P27Gk2L+fOztYnTeLCNfc9DtDeDczn9i8rLOKa/i+meX+RGj8tAmI/PNvlqrHZXw
o59ADsDis73N94ucRu1YmEyeEEPTmAmyQK8BaIiFir9ZY9mFYMZ5zL5UvItpJUe2C3hJhq1Logfe
2LXGA663G7h/WMUtRiPDmaESqEWD2c6TvRC9TPC38sXxGV6YfdFBljDrPmHdP4qizMmSYuJ7nAns
b6qeY7E0+hFzgMrJ+fWD06RVZcrf78nYB4cfvIguuta9BXhiC516fFI8px5C/Ix6aL9c/VcknTyP
jEzPMU72nBsbMm4XwaB3MWAGUiAVqXFpurkLWG3Jqvks6O5toAdSKk+E2odFfisNgn06iBwu2y1a
BbonjNtQkQW2F5ExMK8Vr5yG43pn6WYiy78+oBRH05SSrP0+MDNPoi7D4vm1NUr+XiccBqiQ99s7
6eP+9oYp8RH+5AtrtkOSMNfg2JhXHv2GRNOyb9EHj/8rnPyaVctxuz1TEFfWmpkYPgW0KD9sBWoj
PJrtx5m/59W5fEvvCYPWMsECM5vYJA6f/3k8BNA387fb+tmfPxRLD1KBBCe8RHl7Wkg6+aZca/uu
onoelKjNzBGX3BIUHM4sMBik5LcjyGhNFfIEfwsN062esYHugBHJF2LPh7TlGV2iA3tOUcMb3Mmb
SatoqLQdWZln2lZ1WF6WPq/3xPbkg7KP6rM4Fkaj1VA64+MAjO6XJbdNzOFlybrQn2Pyt5pVgTkK
na+AA7bYyEkRUSPhpdQBDOstm0H71O0n2ezaC2oKylCpIjVcmz4tA+yRDOYlw66oujsbnCQh4i0H
1Cw5bzNNAU1OTqKo9mYuZhomx5NgdTiUXEOoX5HrFtSYv+91Tmr7feSYodEhfgaK0npt6BA7PUfx
g9CDAUY3sAryRyQ1fbvy+qURBFXbMcgEt9YJ7CNkl5H4xAUhax1wC/xxkeB9tqnemWdf1FbaF/hI
3teOJUx9rBwTyZz76QmFEAfhdqPqFGKnHDd5k64mI2EXLp8PgiA0MYunUIGF7RYNh7zP0WhIYXgw
kiBUKzcK25A7HMVCMgPAXrYmh7cnsYp9NMnbIkCxcWi0sdb2QLdCNEc2aLX6Y6VBWHae2oX/33UQ
mTOBuLi7QGIKm93XNxIoYeyFoyx8ixCz1MkQdmWd9wMtCNzeb2uhIAPe/uSW5uPnTPhj7LRbGA9y
KoYq/3xyj1GERhI1hnanF6KMCJTt0vzUR3xjd6LkZYOtpB7NvtevfOUPeAFGLrOEYMC+zaOWjR8R
hct6ZCA9tngPgmQDIzvfx+C4as/1EmE/H7tbm+EtUXettn9GQlHE5uicTBnE9U3bkvcZq0gi9kQo
M6rugCzfn9FCB31DRlDb6QVsQ+pKVdcyHO2fLsjbhi4+gZOdbkuisvuoiOQ00VUwGoHw4av6QWPB
ZFaz6c50U/jq+vuWMdevPqUUahrn1lR+QkkpT4UkfsZls6QJINcqefJueqy2BqbVviVAUq5qB84L
a2RdKrv9pBRuGBJor5t780dWzGuf/d5To66Gdv0BMZUtYKxA7V0M/RCvf7UNURETQfJEwqFBSAUo
yIibkUAvdZFQqb2ens+vSo3zMbEY+mkPAshecj6sQsi8KAe1zZSR0gQozV62Ho8hAkv7n37vJcOv
x7Onf8JKsf4wUdNj/25leHUhOtkk2maclfaSB9xjfDVe7FNLo7uiCrb2HC7S7vUNH7NcsHS47OGc
M8xw+ixHH5AykmikI/RBpkyTjEZXhgsTZshjJovtK7+82Tnfeemnz0DK+5JStYRckybG5/diVFum
pBqKXtU2vs38W/hfJKA6N+OKnyafXKepo4zAQScHMbHBQ0c+Y9FWYuBOg5Q1lEituP0knNVZn2R7
9ElcsRt3pNQ7YN2yjsHrzvk7ANwOzd/NoMEajGlLnylGKWCzmsOiLPGCfCiN8oHtRAJCZE5jHwOt
xXQzyMIqsCqX7qe5mOhJIflW47Cdi/NcwC7JCQG+FRHdKnX7vEjVSgDauAxJQLjclIb3Afyrko2d
WRG9KS8cfFdWqHizLZtuPdKz40mtR0+/PGLGAG+ZbDdC8YQb6AX0WIaJxSNkYerqVrP8B7QBuJv6
RPjchz7nTAavCaoTYXmcfRanxV9uqORVFmH7U+krf25E5MoRJvUx1PGk/jO9TOC2iNJCcH9hMp2A
tLn4/TlQaycR3/9V/jbIY7NvX3b5sroMRHw2euNpEbeUVmjcQM29vJzAWtHrvkzAvSmwQp1Rc70j
uB8M47AOCHeWvO5QQ0EowU6sPU9NCPoivhPiAEaWyzd3dHCFPs5tUFHzlAdrUXedVy0rmZpuTm72
q6DccfKNb0yEl7ktMrDih21jVEvpyBvfV8Ofw8Sd3snpH/8WTzlz0D//CP+p5EPRpKsMo040DODq
kFnTq49IGKZCLjRAvc6VppDj2Gcl4Jgmmr4FfZ/gnwPZmHYNxHBV76U7bmZrdeB8bdmjbpniRFZS
k1A7YVWZWuJpTqpE3oAmK9i6wUi4LJmjOzJ02+okxyj/o0K2Z9VmVdO/47j8OEby3ToxRO1jR2cX
PNkCWC0xM8yYerBIxKklKq8Msen1y/QD/v2MLbmlRQGYboc8dOl/cINWDJfIFqEiwjfP9Al/KQ3A
zuSxs8XYphPWPokebzAkda9bRKzTNSgDTSl1UMMZA0g6da/3bFw0zM8NjGu/bvJ6dKgQ+2NxwAQR
dkzTv1jlGb+x/eDHvaidjU08PiteFaphrk93S+IBr387wScGtzdjCb2PDHHbtThTTjAFC7/gpzEj
mh03MUClnWGH4RaPb9RK46nM5sR4up4UFoWH2+UWu6xDnLN4tmC+dItosJeoHP+zBDgVfI8pxSdD
W2wJjQrW6FP0XKcHGXad09LCJ3rBUvOxUbAOTiZpLXkIp+F2RghLQHsZQaZrEFb92y6USL2wK+hZ
/X5t+OpEmDpexb8AzNKW7cDlkKYM3ZyMxvXwfEQMf0n21WRySdGFrwWA8U02YWaQEkwpNxAqVM70
sb+MyPwohsnEGzr8DZpup2C8UDBXCO6kep0iZqLPrSIOmkCgDqjny69QtBJUo7UZSB83ppIkCkai
s7Q4QlW2wo52yyEtXpEpPSyWMs/tYQlItxubhhYgYKfWk3gc4nlcarYb5QYCLsYwyQBs2BOV/4I1
KpFx0arvP32Rhh2ozFIfvLx8r2DpZO2uzwTYT3y0JQ44NhYeDFP/doxzemtxLWR3EczsEtag9LYB
yZOV9/EYb8x9NXEL9UjILizbjPlEORYuKR70wB1UYqx7bD93Mz34yKaLMeoMXDlySpcVTyqZCR0T
/wav7uXXxfMlY8Ic8NIgfQ30JwB56/df0dewxTcA+IgoBshCYjeU2PfaGHIltkt5s6zGD6IBhvjo
22T5BZ7hF6oAg4UMrspGtF+qIVVjdd2258ktxVFPtLkkoatb9Fd/P6X/Hk+eKlCw/wDDH2C+pS2s
yf2BEzk53fN3aXraf8oq30ggTzWQM9L9ecp95zGM5eKnJk/tnOD4g0LlbfZgwX/rUto6KTVHSUb8
od1XxkHRtMVjBJR2c0GDXgV3QzNHeBnnH2OTOWRtTiW19INs430bvHBAyEns6Q0ZkSYk6tq7X+Py
vOB00RJLWDMXETJPBwfT48dFpBy2hHnwewz/6ZbDDY9m6XN3MiiFHEFBSo/uU3I39qNZr/pM6kLu
W/fhrGt6o+TZJynQYG1F+xK5xwOjbLsmjG65cMOsZVWDFfCLb35UGLWDpX98TXZ6Phsyi/u2sReX
bYdyFJJlvReAH+VZCSlo+xZUoqwfNDHXf64Z+EqlnfQOS2KIQDWiPUKZ9Ne5d8L2Ob6ULUVeBLqs
bp0QbFfd1FhQIHP3sbVsqoBzdXa8SORD6j+DBd5/mSIWEsLnELmg/5xqs/Tc0EOtuxWxB9qbuAeF
CKJN/w3SRe99+Ar829CwcfaOzLXpCWcwxuWE7shgaLaH5+XwYUcJRm3Lvmyot1W4eUi7K5ot2mSs
nGr37da210qI3F5nLeC9WPtvrUZ8BJL8gnLuY2VNwigvXj2iAm+c1f65CoGmg1upJ3fmSSZV2dK2
sOGXVtTiEwNRostBsWe+5hz2v/XJKrUQobKphaNZUpy6cVfg932G1N1toN2JmWRrwH+m60x/IHHa
mDGg6AIkQhPESWF6rXGJA2x+u6e+6gyYcWJXMwShVE91bS/VSvTnqT5B4krur+4oYyedkVCD14Mt
P4Rz2xFZUnqIN4LtZMlQfMmQEbvSzLMJ0RcKUxwd7GeYABACi0pmGcawQhOvnjWI39bJtc/mgzdc
PhXNgb+KYMNTmMd4D/CGzEKhiNh+Khtzi8jS50NPe+3AYh1zmECVveYJt7NkNIe/WkTKYIlPbtnR
oD7q/sbbhi6HkmiuRfQxZADvnZR6rYIiROijWqo9JWc3rTB343KfVcS3v9iaQ/SCfVYxDSRGJX/m
B2VPaKCuS7ks1m111uAuZlr0YW3x8DItg59/J6DqCj+CpOo7jziFYQoUfRjVU5Z8MpKvw9118MyM
csCVsowg3RFjWDDlXZL/net6gTBpfn/ZxPINV0wU3VN9CyeeA1VLcpVUtbXJcXqs9PkfeE6/bb1g
wjJh4isS1r/F1j3+LlaDu2yA4u6zxogGUPTh7t1fXly2M/9Jx1Hl2WOp6kdr8/s1kiiTXlv/HJnN
3ZXrKyxpKon7dF8/NnnJHZ/3yOh9ZKQHzppiNjsaPrmQACtJvDskyU1RriUPYH803ld4R6Zg/O0o
/pQS/YNaKsYp5RBWjjHe6IB7xf2k2gFQIJ89XWVC4ToQsZHw5xBWKLvFF+CWtfq/6RXx1UkXChHe
8W68jsY7Mz8SCPa7fVcCqVB/ihJ9WctUPjbt1D+cFDVGFvr6sM4doqtjEL8PbIQcr7JrO0+z6OvS
flRGZUhdL5n9cE8QcAra5sBCRz3BRZ/sbNi8RSB8578drymrtg3ToQDoCuTb9jnmVrq0WumONEd/
xqjTdyH4N4cFn2qt1RXlheYiDD5SwezyxHy60ayhLGp6/8XL/f7ygMkpXAr7839dsIQnRd2/jQAv
np4I6dPDCC3HCHn7AkDSPvshVVopuA8P1b0lQGn6xU478mI/S7K/bwYKWJd8HSYwI6eliBrX1qiP
Kl2GZ+nEI152JZBrjZelBOOacAcbpXNpNzQnNtZ3uzrw9yB1gdMNNPj5NAnN7E/0iDTqn/Qe5N4M
Um+5NouCdKyThUiJZEPvPeQVs+XJTiGnb7AUzWYje+0NMM4HwleAhz92x8/H2+hFrXLaVqEUlirM
6gf09VpPSGql8rsK9DDGlTeP4ptkJcBeRumHSUDJcXYOz8SKD4ZVrWkSJijvKe8vxUrNY1d8UP3F
IjYAW2WMG+SNIY/MOuPaWF1v/0cn9DxsPAwFdW16AauMzbznIYBMiWkqYfeb5AyBII/0FVaDdmw6
PN9pQG5bvLaTuD5xpYOZsZamPMOHBFJWtYbLOWU4SQ1/vIgFOPKSaBg38wO/MJP5fvo7Dfm1iMVx
sEfru7cJ+UZJe2Lskh12lrG4KZF5DUDy5mRsuPLbdbwdSt0fYoSnBZBvNoaMxZWu/q5nlWX1vyE8
rpJ9ucBjvZHqdLhitpZfxSOfG9xwS/lJ9wJmN7RG+1+4czkTlg4+tMoR1is+OY1bUSGOklK9f90g
pdevv+LN/KhEDAvCjNKThIjPHvHK2Q4HfQC4xEWGDgVF7Ow/t+blWSDw8vy7MIBuPnv31shkTjhC
f0F3Eaxs527FuVEjB2EgrCVmPUmm8mY0WmLpt0hOa/nAsVVn0Fv2VaDEdh6dKSInRMFLD9B2QcCa
isM6CUyHxoFPkBo+5cOh2ieme2P90Dfd++rTQmAdNqHRhf6BdEuXsj7+xRIjUWeGMaOMvRaH12iG
IaVjd8LYOwKkQx5dW4YrbO7KcBkdmBHIeD948jmx//F6+cuDb05GRBNY1WdPsbG9Ji2BTcw+WTFO
nwlxjTSmIgDU4F7/2e3WqDkEFtgu87Lv0SiJaJmjAeTg+l+HEh6fiu3aABymbVWw3/uY3KBE+Ovt
VrEdAI6XxD1M/OnGzB7f0L9VkrGOllUYSSb2phovSnWlT76p7p3iefEmC0GnljGtPfnFeoFSo1on
m1LA7ygxg26nw81TBKiWwizQbQ0weZnNtSzttmHsuB7VIcvN1+QIF6Q8s+jpcZmdt0Ok0Bxnalru
EcIsOcdqnmCKIXnpKnagn25zieIAgdcOP303CCzm3aAvbW7zrYMAejKFUnK+0G3VgNlee3EIaDmK
dOvj7R+gcRvvz0zx/y+E844FhNibL7mI7hiAaVdrerlXoTcBAimRRx/+VcMxk7KMMPrHviAOPdx4
JgLR8L8iMr2MvDAC7KZ7zdOD5y8CjhLXd36gNedF8yZT1iuA0z9MzNlWJt2K8HMDrOFxkwbOdc8X
HHQLug7ziKW41yw6WhXVN/KhJgZPRTuVg4Jl6BpA5BnVMJcE8pdyeaUMLgSZyj7tFqdDN5aS3Tit
dptwZmVzAuGRqWmjGgfFdliWoAzYUcx2RuVoYdtWpcRdQM+oDMEKqZuiYASU5jjUEWVGteAq87ch
+ntGKswgH3ch6CMRnmtWeRZ9GkC533+cC1wDudki//eOKqrEAzCLcN1DrXMDXCNsIfAFzW8NHw74
wsOX7vbX08Z47q6likbENJQeHRnJobskxNebSGF78ttzztHPuMQeSGDKkuhvf17E0Cf3JVylsWjc
y6qyUoIcb2NT4ZzPKuwnsyyzIMDr9Ml+MFU56C8g/uaNE88uFCxItwNSvXiswwtII7sJa++rK4Sg
CS/GoCvLeu3Wqfoi2w3mzAOq/kVx++oE7TDpn0ZmRpE5eSAgVwZXJgbfJ+ePFIa+uQTZFtIgGB3q
WO4CB2vBHo5RtnQv+jwzhAXQfRdKSskhOS6/rTaI6nxSpXAXlU+bo3Nw9GnRKaY9vrJ5ejepqo25
cpoL5ht7WctVIlllBIY7WNqpV5rRngg1twFvaoTtWvK4k9RvS2zjaYThQbLe+ljxK+jru4mogrpK
H8Rc+FnAN6B/d/2VWyRHDsnnfFs+Y+xOkzcEgrTt/q+HMQu5TYYp/mMi+uSxLcmxJWxL/C8SXd44
rZfaR2A1NzBFVKWKgXk9npTBi2tzMDgKyqQcTvhgjmE7z6CBMpb98B+oPl9+E56/ZEQt1Uo0TEwv
bN/D82qYJVrTdVyonZK9phnhlgcTkzNU5HS/BvYOp5jy6mBMdvgCoLpy4cFI69ymWDywJn5WgO4U
mh6oNePEot5yIQk9TC0JEHHpTjDlSsrH49YdjK3J+PBdl2sMAGh+wNq1tfXUEFWTbKI82NEs6TZo
c+YAlOJOOqGfbIv12If6Hn7BOy55NI7xb+YpR+qGQG3UrHImj5zW9pyyrfyVZzJStUNjoWit2U/4
FUEaGcwroKQUMn1Q0/vkAnLpZEZOSIV6llRHqhXtX1SsZp67o0snPuOUkPgavQpTDdIga/ZQ4JyX
dxFy5ktBJ83UZ9dRk7moJ34D1aegDwZ+Ch78xIZSDeyWh+4W9qjZos7LSZHGyOmRvpiVlH0Dv0Nk
HP9+jLmfpRwbzDUB7E+mZsFHlUqHLbEt1vfO/Axpw7GaEi9YDMFaZLITPM6sEVbPSi8no858FBpe
RrygorORavtXZV8YeBPKymdINm8RnyiakbyRJ4vFxriX6WN8duHf9fU26t0mHCEFTeMDwlT1b0a6
ddriHMlPTmtJkjaoWY1H0kaZl5uF1ky7/j5mmo7+sZ/yeaYF12b/uMRjXsy/sSe/MwB6Hq+hhqdd
8NsY+rqdqzmuVr6e0VsInLq3bp06l+j7Cd1CvQ1dvc5c5NCtcTPuqSd9SPqPE7apLUAGveRi5Jlv
sKnms8ui3daciOYMc7hajdq6kQ6OKlTB1cVN9fupQxAd10dkXjPFjvJXD6ciOuTc/JiYmoxup/sZ
IF9EVRiw2MZNGNsNUyeq1kM24j9UBZHUWdipEUb8+oTsvh5qCLDlBlc4wc1iTFrqOiuag3gxx9Ry
odEyOdMBOcQWj1iE4VQEcUjNTBcwPO0g+hImYgR8pTRhkEpTCLmmE0EZ+D9Y4SsJUfwNBssYYvTO
h+mmbWqBwvpXAXvK0oyXGRlWmAvcSn9H0KoiV7LiKd7263S4eEWllXp3UNa4p1dqgBH/5Vb4QQ/X
vgDY/zjVrF3pHMZIEpneFou5u+mATsRUL6Gf8GYXIYJOl40HCN5z5boldM7cLB3uM0KuVNg4rDAO
yWTmUNgIXpDovJs1nrCsvdLQammhSNCUkWMaFK/5wlWTkJSFLmP4+WoFZ5juBQblqYxnMg4XDtUr
IpVJPtluG1CZyK/KWXWlkn8i9pzLI/d2VeRQFJ/zTOYYpU5LkbqaDfet665Nub1L9zN36mNte7bg
eNko/Ei6GLEViZDmPmSCa5Jbi1+RdWwb3EQvISQ+RcOJTc7/XZtv5vg8+tEpOC0dvRG5+Eo/bToh
r4fIKWnkr4re05n0YfgSE0/+4lrabACaRXrpV+G1wo1Qq443s434iipyFOXQTDpccYU/NYZF+e/u
tqX7XsCgU7a3HrEt/SIcGH76+W8JkCzfOpNEx2/frd/gBfizF42f+GrVHnnTWuQvXIxDP0R1X4GZ
ZFIDA5LJ92ayH5yrlkXxX+p8zSmdxifYsQNs8PuZ3oZHVaAb9Nr9QvnMBkjos/N3yOTG1CBm82pq
1hlVgo85Gh4HuVxUDw6zMoJPASzvoOawcxBklPBJqBJ3v/zsH8o6D3262c34TfXMKtKVoMJ7hxnW
Qd21ds31ZYthnn4yOMmNPH05dP1pDhauckway3tJ5yLKK7GkIEipBDC0aHJl1EN9ifVcInVAvMsQ
BzcrToEA2u5ujIUmo0NnpOPqG7mjfbVtEcpyxZDUPJf3BWVS/9Rauk626DgVXJcRsxGdFWUL/yQn
T841t2e23IpT8po22cG1AVrGHOT46A9quVbuiRcjKPIccNd3IEQHUBiI+M+/+rUk3i6L/Z0/dkSD
EPlnKnybH0DP/ES23lDv9V3smWmmq0CRjszw5/S1Az1O2UpICH1nlvU8EKhM6FsdmdC+/yfIoXR7
5x4BObG5fnybx23Vu5VunWz+0i2Xs6mJE1m9Pjns9H4iMxN/4yW9LW/3cFAqnA6a9tdC8Z6Hb00h
j8lrYOwrWpACmjtore6b2DSvEHoE7QUNHPRJFgnE1/iaKbxr+Kbqv6Zm84aUSUfrM57eceaB/eFZ
bsuUTaa1OUaxkPJ/wf/8uYJFoAdSpxXrDGDAp2R5HMPtAlbZcV8VlYV5yjZCtcGahGouB1Zh/d/N
D2RpJtQUSfs/E8Wdtcm2tEKPQOTgI7neSh4Nscjt94ziIVwjQngCA7HVKXgo3BLlHxZJT09oETZU
QrEX1GTwYPYysWJBmk18IZZvPEvvLWJ4GknoLIFPQC8O+VRo9QFKkc0nx88KC2IrymO/izGgAW5d
bcR7IbN3jEJ0nSOw1+w+buBunnl6gfy+E7+OWLNaGUrZq35QagYDtPBqICVCBf7i57CAAnQ/8n5f
otaCZxNMiT3WcS1PWTr8LHL1Im5THeV8ptOIKEwsGQ4fKJlQfdeawk/YeeJbtuZfyb8O9uN3F64r
mIpO9LIAjmXWkb8QNQg1cZEygbfVRbPMRuEbIJsQxPy8P45AlLUTneLfizx6Uno5AXQ/AhdQMSvV
bsahCeFW9DzxOOl/9rz27sId0R4fOmZ8M33AL1L33dkCKXBSLme12YgA7fgJFDmY3PqvXHMDYRH7
iwGpLYrIXVa9BgZjwxcHcle8+zdNmGwPie80SJg8JrtSa1WKIKm5X2qQ1MjXTRu2T1zZprFRvBXg
vMmdruvd1MfySCsqVow8nSqEr5CM6xuLqgWVeQqblVYmu9g08a2YY3FtwoWT2Lm7cEopYeEOwe4x
H286lbJS86PICtLwPpvZp6QWKMYvy5VRUggmFWx6lF0bh3un+Gl2NT/fxKDLrpK257cllAukinMy
52eQ3Y2W0oilgu9taR81VtuwwkJZxM7f6MEysZytqlu9VPUJuHEBsXFjy5E0tX3BYTbIzpF9m1Xf
8wynmwXsJcduNPv0EiERNJEyYOwpW1DbqNHhlBdvwzvGJzKhdqo7EbRVScRGrTkhvRt7XLXu9nLR
kyZ0sUog8OibvUovkY2uXO6+F9vpIpo0YsT4Z6HSVX2YjXfGlsMtgq+X8FOzmb2DCvgOhWKxSK8g
98FDZx5Gz3hFs/3RybB+S8xcPur4uQQTfjDyzjxCEkZoSDpF2jEDw0H6zHC/zLulP4L45aU/kLKh
4zdi/t4ClhIlwaIB6mruI5Ir8PwrMcfVvaHbNvcMYgI8SXmjdhDvPmVsZLQd8gikNaruKKPBlTrE
QfdRP67VtbkN+20VkRSwXz3C9Z8G6W4Meytf8K1Ps8x+zKACfGtZc/P2HOlqeJDfU4k6oXhtBj6/
mPm6LvPPZZ3fy+dyqKk4E7u0uFBw2PYBzt1Q82V+TdzqAC8mpdkzR1j/8JY0PCBQrsZ8ZbS8tPNZ
57X4LAIF7tCYlHP4zfZyE9CLvXwxIBcgHNKI636e5eKrvwxfdWE8ctXjWk9fuOL+CphiObb1eJNS
Wpf29UJa8OBoxdwtazhEhoYy9WmdorjbLr4xOm8ybrqhT/GpK2YIxWVpM5qpz+xFxg92TrzjrQuX
jermSAlJ4mBp7/vLAg0qmCruHJQF2zoYNaJBsCoGRTKm1bC/W5OeoLyU0qCCq8kvR/QV3nWaxqzR
076fgV16CLnolIrSW4Tc/Ibfi+jlFPRBm1ce/IJPe9WLgskmu6NlCOplZ8uurOvOlx6Foi9fUjTF
G03l4CWdXvXl9VjlNCRBXpCgeMlxKhMwiob002GKnDor75eVO5KgG1MjHTdTxJqvOZA97PzBTpDf
bwg1SeaUx0VoqE9glQw6m6erL3TFxw8NZHCtOvzozUwmqZNF8+dUYPKL1Bi15BdKts0tw5gW3rC0
GrTBYunUOyv2+vmTK6oJp0TAUzHdtu4qBO65ORt48HETbR3Dk1l6OPErBLo8BBtgm5EkWiUdxdaG
tb1GgawiadHbjNq2kBjh8XJfo6nGJ+Z1IEV0xQpzF3fYFdjKzxafr2ZEbiT67FPEd/kU/ljwTAof
ITEDfbK8u/pRAXoU4bv0MO3HFWNIshb5+9hPGahSC2QiczmKcQ9EZnkLtktPAB/YcGuJOEBu/6YH
RxrxejSsPaA73EzNxWXQTm+LfqPeOHitP4P+UhVW01G5y+/14xYCuuqI2dJ8jyBvsVRYP49P2qRu
RSEA14AsgOjukwFSlnZ1qd1/UGnQNo5s+DF9a3XgqVXIZZRWHaK5dL9t3ebg0JjYPd5z/JS049iY
ztiiUXP09lcTSQLIaC8Cs4oqowmXf/9nY/nfsD/7gd/32AGQQaMTsQKtbVdN9uNRUW3Z2BntxzEe
rQYSsTA1MtzACgIglm5cxdg/mGiScar+erkcxjg08CnYdkcr0blghgL837d/f1BPLkj8W0i2wnsW
w2saJhPIMX6CLpuTfVptClQHoAy5PSJ7RrsA7qIQ/NlPHrRrFZlvNj73w5GNEnGw7T5znPRYlk5W
ULyJJPGGjfeB9FJFNPh39ZX/Z3/dWkYq5EwuSXmsJdYXemJstd/W+keDZKpleP1wRoW8RzZ6ws8a
y82/5W28OU1QDDCESgFvJ0d/ogc7VG027+MiPhUYiUhv0ye1zcJIBILheuOQCMm25eHnnMIzb5sE
p+NHiestfrx9dzN3OV01GPjIPoUpYn1YC/1Exh/9iO9P3bKpbUaAJSVuopeOIrozIS0b0cVvgqZ6
I7+ZWEyIoUS39vzQyym73Ruoi0Sz1BFq1qsT5Otu+hs/VVJvHDk+9ohcMBoYiQHXk44a+5WszMM6
5MS1d6CssD9+BaosgTiSj7ipOB597rXrrtmI4fKG8nCSp4hrlWZqUXyI6EuJvqNokos9x4pix+rD
7OtDvGXLRUPzOb0Fsm7QnKUQ7515NrTYtUOoqWdBYGH8GAF1bu9cC9mbEIm+3NnDQ5Fftpa4y2Nq
oObDMJnd+lk1GvP86Oj8a+CNHGcS7Q+5mVoX7ngXJTYF20NtYUtbWoQxIJxg1PPoF+C+SqqQmBZD
yMZxMXBNSeDZ6kZYUKmE8GxO5sRMrF8bGa7E4LkVnLs5NwfOl7a+jOb5VhfTcg26132RpG6VblMb
R3LHnwuWNdRqStWvbcb2UahXUF+2ElpMXCWgqXYDhcp2hUOSO7ffYdJz6shZtVNtwu4icqQC90Jl
oJ/aH6cTHIoe4JfMV/cStY0qzRnVz8kVDZzjitUbW4+KkLUwViv/2MYYAav0d2e56kpDllgfX45V
NTsdFDcWNZtKqtLjtcGvCx3EhVX5ZDnaSeD/1bopYedrWS7KOrlMCUIudiG6oSB8FHdn7Or5rJBV
nm2OGVqO7Uo8kUXOmftWsu3R9DQof/ADrdbhD/2SHPNZlwvn8fRbiZJHbYMUgbFxEM7BwzAP7aAA
RNf/W07je9+TWg8Z0eHbRwlBHzGFT7ihm/yDXRi84mKjdeZ4T9Un/Gql+7PmJok5+y3bNoSGCzUK
EFrCOugpl6O40VZN+XzhqXHVyyKt9+Yd5Yk5aq3CYnuPaXMBWOepjiZDIjIgHxRSizzLevz3vwG3
AzJJ8zfODE73JlV9LAdDinh5LOkM0Zi5THZlv6AmtZt4QYDafrUOmdNakXdSt0/gpPmCexq8LzeZ
9SoTjuTkqhRLpqgDCExEIIHyw0MSqA3yWzd26dCJWMNZow4mXeJuyuGHLfHGqyYVE7m815jDd1U7
l3xrX/RiwFSTcEk21aDdapnDO+JE/hWjic7aUBfdXJK5C92kkMDBcPJsE3tJ8J5Rpt2UjIcfFknO
BFuUFOf+Gi87b/Unp6IZbqLUDOA/5wm3SdEn6cogX4lZ4GcRBwXgxwgMG2KoBMd3nvKGU7aDDwvW
pXWeZzoa6q9xhKLSHDxmULux9/NWHoXjdy9ayq13Vd8cHgxnImZGRm8efYcErL2cwxrhq3e6GpYE
y9MMTrnnXOzGmqTmwlzIdFvGZYKIAc6MC7soL5W7FvHoHfPsIYOWjXSlwbqvHRK1rLAbto+xYX61
dHX8qJZ08i9TA0ildQSeNvaFO+RvwnGsdzeWkK27LX9fY0OfpdZFBfvHDk5KdIK+bKev8aJIwVvF
2EkoXqK4DHKv2VxVb2a/f0lydwYTLMhbSvu8b5OuYxAEZOcH8Ps4HQcOAIreu9hfLRyTEoi9V7g8
mijAZfreCy1WDsq+xqBxiZU5GoCPEsTHAFEG5Dg+iDgrUqmyLqVT1xx31L4If1YtEzFNuK0/5DzM
+EY5KDUYjMLjggwwuQvNb4aNl6/OxWD3RFNoYgNZGiMyKAXs3fw8eVlqtZBALLxWou7pWTdSFekd
TvxenK+AOLCTZIR16yGcLn4sgUwNMUe6UgwIAHbwkMV7KMxDrm5PE3+c1Or5XEnw9uXpwOMnvV0l
FhtXFllMtTvsGHYmmJxul81sIpc02z94E1Zyl8/D05rvPXzvsLS+d6MkicMsB8UXQMNNr+lcwxE7
Pxh426hkY6bKP1rSFJWSkD8MZ6CEC7WTVS3JlsLEKkdJ0fpLjwlq02JA6UtgoctjYdBIjUSOEbR9
ZVh5cQ9VoQvxOwtkrrX7WraifBjYJM2BJA/l8nes3Qpzp3tzN5GvpXBIRV/XxTSZsnZ+BQoocTBE
RXsSihI/CtuLj8PUd2pKWW96gOdLmPMKmf1jqPP0OUSHiOpVBCfcnwnLc4xOvkF/2j5WLa1B3XC3
UcRpzlC864lqqEqLILiJGQEzqPDobSLd68eDOgtjRLts/zPvC9EObCliZX471HisU3Dgy95f9jjY
ExQzbHOrUQCXPwGkkDcACWGIME7uLX8pmb26EaPeyYjC0OEbO7BFEJh//AEuOzMwxO9OQ6MoZRW/
TxRvJMdjVNTvK/PrsikxIg5moRWUsNzL+ywbXVOIHBvuDcl6rc7M/7NrrdgiW6ae9lgxCBDA4iza
SyblnETCeuDMXN7UZuVFTBjzb8gyMO8vm6Rs743jYwUiECjllI+jTcSmRsSKAd9hZENDHC5F6SIg
O6ePwqByYIQQWrP2BZGqxGeyjzHNQHlyLjSKZgZgqetqUjaiKafwX13fX7tzU/Ew+d9nEBVReriK
jSFnNrIip734D3ohH8x165xubcxyB8jHduhlwVUu2JkXU2OaR3ThDtynAttad3Wsah7rLKrAz2To
lcW4SC7X/QF4L6U6qE1CJ8yO3alge1TLptoi2rp8DPc4+H3fM9BzN6/r8LPsExzSXnx8fBLoVNqU
XSLPooO5NjIkGRbjVJhuV7jp6zHJsE7b5LXXgj6Lv2VGRsb2wdYg+CkcPRpaBs/9SCt0RC7f8HjG
8ii2G/hRrO59zeH3XemoXzkS8cXBtebaz0cYsC4J+xbQqySSElTCNgwly9jZMTZYu6k2SnZM4DbZ
Fw+4afj6nODAw3pj4rUHx+ACuycruU9/hvelZdIeHlh0jTtEapfn3SIyW8X5X16Gaq4lBJUKNUW5
ggkYJHIvvq+anl++br8ItyZJwzmjVZuFxoqFUoHznKTFX28xwLujfVM3zUW7j3vNRkmmFYjhutB/
piTjfR4oaDWqb2fiR3sIqzcwrPpBxweXP6HD6s0OlaPzn2qdTRtNoRyJLvyMHWvRGMIiFu6cBZWg
DbayDsgPXqw2vX5+TW76uQelMWnz1H8BmsL6Taltv3v3MWjpxEgLsY1HNxu9W+TeFyuChzyalKyX
Yl3kdkAVvp5yaIDD0bIO4G2uabh3q8LC/sxh4Bd3xjAfcmwPm51K9nMTgLsRvCOWsxt8TS3atcWQ
/iVlV5tFKkPjiVxu3qQinMtW3eYDN6T7u6I8NuRnWpAJxwLWda5jpbheuwBjtjxXw4AiqV2Y4EA7
wE1sL8qCsYMfClUbgFgNIfN9mSejRVWEBcgAlkB5cuozsOeHLmq8QE/HRo8sue5sZStr64BZdjOT
6OqRg3f+xoERURi5CVus/zTa71Y7F2EhAuSSxSnqzTVEdSxg2jgdUdR5pvdqHB5IUcQM7xsaSY29
Aqo0+dMWvr7HVv+CWXpQN6Vr0g6VRwJhxhqr+tJ76pQhdZQVQ1GCCbMfMGGSO8yb6eZWdIl0yE/M
rdlXA/FJkvw3+aU+McX7VQwIjDgnQMNup4+pcgDyg0AnNQ/lyFh0BZm2OEaEq1cD34cvKovWJOrs
OxzyxzraaWFyJKkKG62NTT9ygdeFjY8iEgTk70Ic8DbsmDbwLMLPdZMIt7TKc2IeatG8afln3Fyu
yHCkCizr7gyDuFCgIifu01bB6Qv9+lgtiLJe/TvD9/MNlH91nvzvUvPqg9SO1WWfiYo4iW7lvAWz
osPW8XCtYKRan+/nAq1y0At+MasOZce0UClNH1lryRPkT+HuNpbFkYr/VNAyJYi1uZd8kXNlb1/j
Hx+JfR+65OF7Zg9RgOxFdwJSb3MRuqRhYDLtMoTdW6LTTXpBu4No9stpMaX3oPhkhOfe8RmZ9Oos
HzCHcGuXuUJHzlvuYNnUZZkyIEHNEu6h2taNu2uiR9YOiuSvprZDcsDl1sKEbTKQ3XH24znfdP0j
zAeBUJbhHxf5CyMOU0We3yBhVrRUztvId7f5hEIBJLq6c6RCw+1Mus4aI9z+fxKxNe8vMMv2HWI1
KhgvUU/ShHAOvtrh2bfEj/um6jjiM8AvKTRVhZPmFLjf8EqUG+Iyg9iYykNi3vEaRx+4zWAsCaNA
KxcDEI93croMvH5a9odAU+YW8Y6VvM2Bv3zoGqa/qgxTbZWUdy7PS2RiQD7wWWD0+ErloAea2IIM
1m1mdH399y6R498Vmjs1trWM7v3rNAiFTzK7h7Qyt2K85ibdNOmLrFpeHcUvbag4cEyamMCIRZUX
XTVbb07xFyLAY5exAnaK9Tb/EyAgqxbc4gp3S+M5pxoVv9T4oNlHDTiRKjlO9PvpA/Xw+0uHNmaM
la20S36x5wsVsF8drLVrp5CpUweY1ZngfVinYVQupAvGOBT7XB0qVtMWyRqO7H+gZ1HCFShi530+
UrHSsSCYGxkMaP8TWE344b5NcTpklChLQYIiHK+hUK0sxlORTDsM9+cVVDR21t2KQ4tryNsaMgo1
uGUcxJHMY7PujQBpnAjbLr+y8W8matJnjFZqBELhvbso+2cO9ZuvmTYyG4wWikIEA2bEBF4UMcYm
Lx6TabJdccHlXur7lxImR4p2ABzzGTRq5xsUq8DGAv7u1hv+qmzdYRzTDDxw8b5PTEMwhmBEuPNZ
aiUe7jRcHIVx38GdrFTfmY1Jw2j7VuJp1nv954LwmXB9b7/iskRGmncmkKK1Llb0Ae9BMHaWjRPl
S9VOHOuXEJHUAfLA48R2JXU0W6uEPyjZfdOWpY5dNWDek0CymsUieKcZc6kO7Loa28v+lYOh262i
NRqqVUxdrb0rNpsdoN0aiV9zQsO93q0lH5kGwZ5zi4UiubYT4ivORbFXEQ0s7NicY6FG6GVQW5MB
vl+90naocyGPU7cJMNI0xW4HxsIXV4fr52jAi1H7h8TfpylDBBm9fj8XLyFAqML4NnFDBJEMRXxS
jaCZm2vlyibfyorM8ZAR4hUGeQauXf9ctDzGlVJPPitMrpjl8YbcNwCu0eXm233AHxLJrq0bu29P
0W4tY64eNFWMIf83glNNhAp/HO+hlqtE3N+tii2AZRg9qRyaOfvMYrbnrSDwRzDhrH1cf+yw9Nhc
vmQwCqgU9+OPrNQzKCJ/ROe3rPOFzboJuqVE1kY8yhevM4OGussstaDhxUr89/pDjD06pPNnj5IO
J7R8mDgv35ze1kmyfAJeMKNiXbwHmy6xW0Htagjb9GYReZmw6Q+1iPQWrXe2DUIorM5cSvf8cNWN
ds9V1GWKLNTNzHihGLQMB0Zx1jbwv6ykx2mT47MmoskTID9w1YN5kkdzwMm4CmPIbRao/B7rF/yu
3sLi8zs3CpTfucHgfBF5gyL+036vlrg0/Tk5sA/3dFgEFIje98meyqOQST93fh1lLOzo0x1WFeLj
jU2TSgDua8pHgWV68gymMuXJdqjTwUPblNV0LIAjV8f+MR5oaCpXoL/hCUfQy8PwidV/V6dBvE+c
1TBrwyGRAnkDIavgTPqDeAsEvXkg6CGs4i+fNKlevpbHIxAy9mVDdisafcDo+aJl22PeEDxxWiko
zPIytlYkDEkrtuArDlkIl1pjmHWsxaU9NgW0ePg0d/o2Lseo7v/tcRUARUE2x82AlOAZbXxg4RF3
xqLsOow2FrFwbbG1TIBKa8lecrRaeDQFEiwS0ZIYbEPfqgcfaU+Xuix8NhbwJuvVZZnJW30fIou2
rHeUsPU7f1tovsx2k6pu0QqMskomK1Q4tOvW+2vcQ8imfc7I8QLhD2L8lZwHBNcYu3USxgM9j8MY
kBbe397F4aQ/SEfw23yDv1MK4dBL6qBORZ0nB30oN4i3Zb4nIsRERLbDTRWk6Td6klB6lTRjGyO7
gOjMoLvHAjiBIyOi9rNLdsuz6WTh7eebP0hMN8CMHtVKKvAHOjFF66mYlmmifNz3Cs9Y7YN+nPyP
i2H8GL05b9kfmUZbfhmpAp2fi7P3Gk+D+z8vg0S4kLclGXQwai9eDEvWw+Nifia7ZEhuSfhbfYAM
6yDUHAFjhLRwl5e11+GPAx69qaDsD4XByqoFud2d7zyb7skdFE6ELqx+S3tIRCqZBsvulrqKqlg7
iy95Ls+IC6bhXB0KM6fIdBo62N2OVgzWq0dC5z8X8hfxLOiCuVcrRM5ai9NdB5EmY9Lq5povfCkz
dJqxQcGV99J2Tox+k6zvVaeT4neMVWVGvmtjU1vJ2h9H11KDI1uuoGqj3BAeckz9LdnUmL7zje7K
kfpE6Rt4iI48A8eMXZ40Kk09j6pFE929imLWWnVVXDNkbxe6WRhPgmtYvO++T/SRS7tpj06EgZ5B
LOfH72U6/aUt/Rc9L7BC1wcJcwAtJ/8nhKaZ5vhJ7aubd5W/+CJngwB8WViPdWM7Iyiv+PBzewIq
tojJTWrDCe2CIv/SGJmZoCVU2RPqxxWaOS29+E0nf29fgAqgS90kl91SqzAGdJiu0Zj7lpxx/CA+
b5nIkgkFY9TE9eo0YFDHlmOFXKrwcewBdbuAD8dJV9YhFH8OwrOj+5mr5AULmp+lBbGyxeBoz4Hf
uhxGAxHnj5hL6cJ8fUNr1UlTW2sfs88iXtTNM6gDXLpsF/ja2r8Q5xSErxETOxfnUSzrCgCKxshu
240c296Mh+Wj7iTLWko7VZlskVLImGQXnfo93rwoj4kCYShaukY5vdtyglFZkOg1xZ3pokzrbs6w
Zaqv7qzeZKbQ22JJ4RJQLesuJyoa9bb6+IvrQSi1lhmCQF9ZFbAWxNVcrt/N5Ba2cSXz+NLdrjH4
M8ZS53ulkIddfns9zsbyMS7ASSJHM5nPCdhJC9peyAvEg+3u7X6ntUaS9FZ4gvtZOx1qose6bSW1
4f2FJnJ+yxxqRGseV4vL8PzilIEHaXReVaZTKfsi1I+sciv+Rvp6WD8Jz5Ec7Vah2o848ayi0up8
4NV24PX6bJtZqOJCf/vFbw4nulLOO4YEbRh1IRrzTiN++XEtBEfZPZPnGdJC+sNJqkopZ2+oBGjM
mw0T3Cip5Rjc9IB8yxo5Ra7P7OGcYHqcM8C2cqawAFrNZzxNRnGHkn7t2f5Rlz6f17vPh6RGlPnv
HHgsAY3iQunjpESh7ae3ZLw8gq7JRnizwv1fb3YTqi+3BEYOm5uJrV6/dzz0BJujfkFLLS2lOQix
NwTARKtkCN4PTemC2HBWpEWJH2HGBsiAFmH6PCyhstkp5HZlVaXDs/GSQ0cYOvoBccE60KwjPVPX
hKbGa7gPoCKeb1B8Ce2kF3Z7BZ4CQBHIHImBE1qO0dxPyOItTFbRK98k9RPq5XK5z+VKRovoFeaq
6w/Q0YOwt5wrrA/w8H17xD3zO0Fqi+r8ccte/B5d8vhNkrVme8iOaAA/62o+qANDmVptdcxz649B
lOpE47yTSKN/h1UvA/sWcCKgXKguLgHG3o/415g94KYzaNmH4TtQmMHQaYl5ioA5unprDQSt7gUW
etQVV2MVGgD1G1Nu7trH/9HRodhtz0vs/5D/3DheN0eZNzqRTA5nwYB27+Q286McjpQwMDdp83vb
sESBEL7clrSyhmO+C17EhWyuHFGkar5ctZ/WC0VqmL6qJx0+165ChIufvC1PvnoQcNvasm0k6Pjf
TTAS8Gk5AoErRFTvKl5QqlX924KRClTDQbUdm0/5fiAmtfWBFoDg7dzX7tA7IAkOzyJ/GNMXOYve
KRphiW2Yna+0HFV+DLkYqTtxvobYJgQnBO7veE6DYN3LVsJ/nF3dwPJrFcNxCQV4SIKD5DHdnaJn
jH1K2whGNIJz1ss6GENV0cdUkpdrzvDCAkbl3GPtF9QjGlle3zfHDwJ7XX2CnfLMlMGJSPdvUDha
9sCymcAz2zM7ULBvvgeM21FdaJR51H81aOB2eOKiyGvRub+po4aAvrND8E/pTbYzSD3ITNVS+RUQ
zxoGrYA2Vl8A60/osLVm3kufyXlqyc9DRG845YCWytQddR/M6l174oeVbHTUepibyaYQZk1u9kMX
poxRaWUxjN5H2PttLgMTjhWJQqNc7GnolZ5+vla9DYRvGHXP3p5EscnhWUrTzVxFi1SlOVPFnjaA
9yLLp8Qx7ua1d7CNRSH2S1N7EtjoDAmHhceREk9soaQzrHCN2eG0IymECtxu5bJFTWfYV7zTSUpI
imdCzPNVUIBv+73xxAsCTjQMq8e0jFN2og662SzWMCq34B43x1qBC3GkvSvh0//glEJAjd8XZJWy
KIjq7QPyvkZsmu8U7Bc4pBrccUxes0QE0IEBz30Jgd/CXROxV5aM4c1K26Gze1BNIaX6wTqz0lW/
qk8Mu7jstsWYSShx4Eg3ywqG7nTif5zxoa26F3zoOT/SKIWELOEvCw2VcXjWpEvWJ7kEyvJpFUy9
8nfLA9IB3z4Z43aA5aPCLjWftumUqvPlJ3PWvIK0zwMbiGzNvu7JzHat1Wbo6PY1acQjFNj9QLgM
Z5jI5AHs0vClxYM1FEdyXjfiF0bSHrZar7D9jDGXeJrX4UMKQP/ajBvYaR3GehLtfaVpnVYXG8zX
Xnj/nbxJmekwLDZXlBx0utxR3JI/IR/4Efmox9SUqfAghTJS8EU64ibBcj1hSZ4foLN1qz0NX1AK
hPK6X+3onm6LmKjwraP8q3DCVTp52/joICx5AsDyVRXfiCUksSdtdniHZ0aEd2NFH0quGt1FRtBF
PmF6CsgZGGZNh9r1c9kaMZaCNShWe7PiRTIcrxVo7bV0meAdvPcHvRVEhM1foH0LWJJX2rUoHmr+
VGyRn2RMmb6D5lAKpTXMKokZOtzjTRM1XATph770p35je2OYtUJCS+VOqM+o5DfhWIQVTxPzM4PP
wPCPkbRZw2jrrmnoJUHA3X/nPZBUO/EbD+uc/Jtz0P2rDAd1SDtr9Lz2Mq7PE5Py8zGMaqd5dsbn
rQgtlkw0WNxKwm+AjkM5FpOr+JIsoM0iX6hQOBtfQ0JkZlTRTGJuVtWJSp5CHx7zvT7Y5sUarCwn
Rm769myJN+9cKPLlLSiOXMfn6zptzu/t44QIlWYZzkLief7nKFpNJjJEGudr6zdfaFk+TvdW6N/s
BilZs3WOcmJc852CgvCo386KY/TGz/Q0yFcsMpyNqLGoFSlkeWjVuYmL0jbZycx+RYTRgL6yifE3
ClDRB9YxPN+BxapOHU/PreLwU9WGYGpPiMX465N23FYRoYEE1kyLYrVgY5wlBr1fTpyyUHVYeAYf
VuOBL/2Nkk1Ms4NxpwN7RUZj9eypwiq9/9QIw+5atrNaTwkdp7G+3gGrS29j2KdlzIw4MkSStLP8
Bf47qV9Gxd9HefJhvp/F+k5ZZdaoKBlPtuHgaeJzRv2ZbP/Z75dxYgC9Gsh3nFrVXF2M2DEQO63R
YWTNjBG+NM2cSJNXnRMR2L33WeC3CtNpqJuDk2k6XfDtcnlpBKzJu9iR61hKijU1SiCvNHTh7H3X
t31UC27nz8zBAIQpBxX9PLV3HqxMetrd2T5mnpBjJg2MqYU3udFa38BXVxqMNKXDfAhxSN899ujY
PtuHdOf8px1nEHrsHgnxEDdq4FL7V+24PCmyAoXEP46GOVspOpK1Zh13/sqp/F5/FP5/7YQnAMJy
2P4VEYr331VGloUo/z9w8UOu7TElBGU5/cBvmDPYCGPcOA8Q0rA4uLny/+uO96uF0SDvSR7nRmwH
VhpOi4lTMbVkj9le7AG0EPs+6tiDXOjBMJUmKM96A/Cgu1pt4Usp5WanVzdZYIbiDTtqpfS1h+s0
UZVFFohElE2vET2O5tiM+tnLlNbSKp3s8Udwv6ygBNQCk5XLtFfbCOwz8z/y0DqfGHxOjtiOfV9i
ecoCdkpuGzMyXcww86uyv+PUvv7Uw3HqJZ5tX9h0h8yEkKRMpwdfviUB/AYywnlIbRJ2SlqFLXQe
WZ529aaVWCtchkrIyB2yoZ9IfGnZJGg5Se+99+To1rh/flcaQOr471Jgex9a7oz5sko70wJyc4BK
b+SgSOfN2AjXyVPvtLouKLeya+4wJLrdmXDZvh0nMLvYfyRLojVtPLT9p/JXjcwZ2vnIpO15SXZI
in8A7pszZmW63rIIodZ4NSAafTS1ng+WgDeVKV+INZfwt3dj9rR9+sI9bC5agMbWQmyOhUbNsQAU
0pyVyTf8vx/69UILoFw8kRoskbDOSWJoT5oP1adVVJy2e4bCDL8J1tetmzVxZJ0DrpHH9ZoD/2x3
FahofAtm1eo2sGICWkQB7nnpB5EsRiIMoxrD6aSjozhPz6rQCpbETJVjfNKRxt9iT35aMD8fW+7X
B/pzqp9vx+DbzHSHSNNEM6i9LvDzI7Ga1KGHvYX9muWMtL1flr2WKzDY1+QYRkR7FI2abPfPF1/l
3tHYh3lmM3NwPBRpDUX+OrLlvfWVDwnBQGm/EBTRWdjAIZ3XcpWAYLdolvbNhNJ6V982zdMdf4SE
C6rDF3m+qt0KKlZydb+7pdV0p9zDTY8up/oBKnOsYIto2l/vtAOduxMdEuDTh/6MOiwze6D5xjzb
Tx4Btm3L4/dHYmOw6rM2L90frXm4RRQ5safk9TmEfXz9j0TZOnLIgwhkVkumdIyv5F3IQ0SV5HsE
48Fg7+wKbtiPA2N/9IBxDUZGY4J7wgXZmAOWlbrK1YioUpK3sJpVQS6NTYSn4P4/2eOvGIWuXIxa
TfspqWK9//gYaVV9dgvPPzxt/E2t4j5jivHBt/nHAmNlGvg0z075x8hLvwN5x17Mimmm/L9BPSFh
Lih5QZJJ3ostS/Dv9fU2MIvIfWtAjmifShMZroNbpRupTf7L9v9Hcq91PjyZYiJn/IjznCHiKf02
UPf4PL/dLs4oRkXzHckG4oK120x3Jn41gdj/JfW/Yna1TsjMzzi2yJ6EFGFfPzPVnLCFJpaIxXwe
lG0qSRe/lUEFxs8koNw3ozI+B54lE8B+qdW6J0SflbspPNAKc+Iy3F5c8seZHDZm8qg7ks2o3uHU
0NVlAWV6yrG0j8Xq7hhdF1s9BHoa/FP/1zO8pXPbfDlOln4FQPrF7GPJ79zzqmCGYkd078DrrUYf
Eze60lizP9qKTqaGOGTYeFiRekemcSkF8HSk3tTlTe5JDxORB9mMV4+MyMba+kZbY/uUtsGoI+1I
Y4eBDKd5uySz+bxIwUWCoAbX6p3yQjYPMe8Ty1i3X+Lt7tbRjBLle8BocqRjG3Kyg4T1rV0s0uwJ
nuVLmcvzF66Xq+Eq5o5AB89sAj9Bf9NvgBYjIECh5xGSCFxbNLifojVVEScWULsaortxIwYm9PvC
IhukAxerXXfQfNPAa8p5srICeZ3HEAXUrcHTQ33UO+QokZjjsn5hfDXAUa4d7wIRPUSSjNjRfakw
RzJbN1hqukxJahPNx1J9DoVpVyuT4wC+UcBXZ7idjaO9xV6oMKX05BlLRWzUAqxi8Nw5qhpXxNJ7
e/hHLS8nzosTxjA0rpAJeKg5SHPSV9xmk0ti2cWLPXHIIztGztQ3AITnEx2suFuncjLpvB/SUKJ4
SRVmQpE4fp/bz53JUzjyXACOYWrp6REdk3SPw+LJoMj2RlFl7q0vklFeCA9ujVf34l7zZNuf+qaH
NVUL1z4jmeHbpAiUGwVSA95Jcx8t7ugKSKKmln0kkhzSLJm5oBZG4E6hNIwqD/vVwywWmUXoRWNc
cnDQYDX0LZZHnN7ngdApCuTpmu/hbmAIqC7EU5hy7KtHd+BR1NkO7xbUzEEuSX63R3B3BqYsBLmF
1SbxXkOuXBnB8e1BPCyZ7QwbAFer/I3yK6NU95LfEPzQXqMe23JHIEBZutpWFwzoz3QUhTd+rUU0
RJ+qo+R1xEUamvlORhgMHfrspVJY0ddwkRipO4iVq7xw9kV43E3UbrBM85OhO0xrnmgQa0wKoQy4
H82llHu+pkaIuTSPN2tjIaZwbYBDBjs/tMK78In1fG+51OviKowsjl9rNwh07tmjvf7+ZMSQaG4p
UbqHGwazm65n6qn1O0q7im91Zkq1TKp50cV/8UUo0hW5TMITw22SuNTtzqqiMOTkd5vPdHHjDaHP
nnvOmAdNFrFHBmrlJqzdrfUGrgNFIi5ARay4cfMtSH+axOKYuLInP+bCtAygMIMHJW88fXXACNgu
V/I2bIFKo8nUOfUFZF2TeugGSsNgyXC+uieBqKUj00zn9FNTKgagguTC7g7q4T66uN/a/nXj2WeX
RLU5EeIEdDaGL8Aj5PLr4RCLAg3zmIZecrxe9XebiEW8ME2bR8AtH4xhI4C6RRNuUgeN+4UXsbYx
pTpCcq2H/FR+4M/YVVw3nbut6xOCwfndjAi7PLIA5LRLcL23V9HAtxtuOwmqdbBbv9d0qP8tv2XK
defQzM1VtCMdTFawk3mPUSGXf2jt9sOn3iEwi0QvUHhPwsFRdsTBV3pKG4HQuk5RjndBkP0bMdSS
496cdtJ+WtOZKRnpUbmflvDBtHEBqqrPEGfvOCHbW/hF6SO7Nq2BlAuHpNvdVHc9sP1Rr2LSR/Ma
eAtZ00SaG2JmciUkgP+PRPUHqUvKRY77iX+C6pDezRVHzIrys/Jikg0R/CpDymx/ICXvaH9MHajH
RwMIhCFT1sowLnCYsvM+fA5qPL2lrYH/R8oKOYKnsrm50LoPSJJtYw9dvu02/pb/2GaelfbIK5kV
mYvkF6gdxn1YtlZUphaCPv4zLVrZb78XvvBPXHmuGp4MA0KFwHI1Le/q8VxuLDIGvxnc8KVFXC/O
sD97Mc2j4+TDQhOrkZXvsn0SBITbgvIvG3S3PZY97JbCu5FXnodjtSmw7xj8OWJHPmIAZA8B/nEm
VInOxgLtJO/2uoxLOOEaqIsfvM/O+FTnxFpIu+6RMLavweTAmK26vikVMir/lS6fRE5k5tFGyfrn
r6/eO0xcenRknRoq1DNzHKYfsC602/cM4Q+CpozfcObs5PvdCxm8TZ5we5sGOAVKYaM2+s9xmK66
fBoJaXQTu8UQqcFV7Gy6GpjXAr6ot3PDzPO/fdq10tazUaAlG5kindiaGyY9t3AlF0nM70be3lBK
HOXcYQ7ISx0/DdZIMp+olkuBlaiqGl/SYZqOSZaloyblKaOb3Zlnma0M8gwitJExqzRPgQXiuRNm
sN7IopjtrmFU8swBrZrJaUr7AhCk1DkMBZeuANh5KZ3MBRHonRGvpotcSTQbgXO5ZJUDbTlM2c30
xACtTe9hf+VOuyUoDJ2cVvwFR7c+mBGaOCSTSR1ORSTARDwWmm/wcZOGmzMyzjixMOdVx3hzcCmy
A+P6OW0u95L3GqSFG5KLmlfCTRP1eKMQA4XvN+96aK8mmiyAtHBCWqc6EsPzxSTXpMpHVx9iUy5E
gVi0OSdfA6HABZvPxOSNwocXQwO/GKFRq92AT0w6ocxnikWp7MfIjfcTxPHHPmkT3S9eQGCyRaZ9
GmSMOlmwDvgtsvA9DEeTdesTCloifxPrCfQVvzUxvRdX20L5lBzSIBkjSPh0VZBjDlosQ4gbw96t
gx3NBLUxuGYT2HLQCrtlaj0hyGc4ylZTc0vpa+7BWCuQU8eGIgJeTWgDmMxT7dj5vXQ/EwufaQ1L
p0G6VYGXKkppZn1MXbuJ4yonO1lhCM8MvEOqx0uvycPUfT5vE0QRtxrQKxY/iAm6mX/B5ts1aBdl
ykcVVE6sqGA2opwEecLOkywnNqC7PQDUo//xKwwhRnJruwZbOtXTZRSUJEgNUPlj/lI82qlQ9v3A
rr1gwbjuIY50vKExC29LdaUQaz8xfc/qq7dUuyeDwv4YHYfRTnVJYsPJDUFejobxTvDvAY6HfHB8
HqafK7UWuzsECmJVZtoRQcd83naT64Q9/aCdN8lJbtU+7u4VOVevgqDead9N3UIQtNxZOULY+5y9
pz20OBg5Q3Xm1beSJz1f3iagrePNX63oNhvKwDC48NZtrMZH8ThxZPkoVS5fpvvbXZVhihDYqo+N
+KiWJ3LpdlO1cN47ZNKC7okUm1O7XOtu1sKTDSDIGqLbzGliWL1bnnk2tbkB6KyuB+s6nNJvVE1N
JF0EjAfv09wBrBBSABjrAEj0kIKu3nkstZMAv30k734LPj95Pcp5RGpejuIzQIN5z9vfehdGJF0H
PUuW9OhoAQ8zM1Ln2iIrfwga3Gej8+H8a53KyoWsclOfaMnAZDVQDpdwhNp7rYIuXqq+Ybg99PQ7
mlV3DT4Z5y5r0BAryomkQXDYlAH6cX6HwY4F+Ww86RyH85ZSh9gBncinTUYBazoWP0TyOf9fqwSJ
iqBpnf7D/Ta6JkXdIPhtFIZOdJlw8fbt5Ab+MfMWRVo67xd77c+UTSaeZcJzKeqiDQQXUCrEZzts
/dW/77OrAeYReDI/3Y73D6Dn6UxnE7X8UpVY0m12hPS7pW0YRC746RG1RMLxSBhqipcgWBu8d2a/
OTZk01Q0soX2VnFq3SyeJex2gIhtTF2fpKrqbGgd3088c2HWhXA4e0tRSKLm0EQP8/4YzmR7BNoW
Sa5n2ZVBDx3R6KjIhkzy/a7oTfLugNd3SYBDoMf+ZeBNZOmxuASG7IGL8NwNKuUTr5EQpENbKZbv
30QbugfhOTs7+OohGhnDW7LMf6ufltITE0bSkhdxK5B7LrfzjIshA5wWnq8dAvyRxRfmLRUlcCua
B559KYxJkNPR2Wm4RzpDkf1w6r7G48KefZjbp4Zrke3n/gcPVm014h3U5HxnFuyXqUl5jN8sTlGU
fqQJVkJJPKYA+XFPNRcL6/jTxrIBIQStLhYnWvZexqa106EorUCUR5rQHqAt8FcIRKOegtYGgifi
psbQL9UVQ1IdatmrC3sUFJrQ7xFzM9bHZHbe4Cp7ftfElPD4Xs6uviJs4FX/I75glUMTzILbtKdf
4G7+cKVJQK07IB704QkSQWG1Pcy2SIjjYMHstJFI6ndpg1GdGT5kS0KANwWLzAwBuLjp1caiscmt
I8N4htb0AHm5jOppTvzzIyWlPYeygU64KcPbWJ4mIqLgH1AvtWJZdjewJl6EP8VYQUQHbr5W4uzz
UK4nMl/axtuaZc5gqYwhpEkTLDKgI8A0na5WtckpK75gCO/2V3mMp6wTqJElRlS1vQNJzZuLCQyy
7CRd1eGrqnVzgryfSTAPDYbQjzhczvJaeoSTLwhwmP/Ox0MGJ1TCACslXhTseqAKIhlE+APmmqzd
1eSCXbFgw5IMwoSRCUl87Jl58D6OOc4UEfxTpA9mY3Cm/GYyMUWTS5O36EjnyJ6b0Qqm7ppr5+Cc
FMtcaLbI9TIRZy0MlNz4Ec59NGvHjyhJWPLKW1RGgJysRofu/Xwb0lPh+R8zSjlrXVpi682Ar8A2
i21vM+R5ubkEmaz69ZhrTcXFB4BAVu/uikgGppMqJPk7HbcxJvOvphWbk6d9zFQFEiCjIfI3LbT0
useTRLHYM06juYNJRc74U9CImWy2TCDKBrTsKW5sOR6eGNiYxnNIsHe8CB1LLTF3dK7nvNhf8vHh
CSHSf5LEY9tfulZnDA4lca9NQWEIOeuQHs20tlYa4sU11f/6XLEUQAIQyJzzhj/HlSnoY/gKLyYm
nQx7F2tEQKK6inMXcEPJZLAcEXGZhFVfvmv2DL2qgwq2biaA7g35H4MRWuCtcgix84BOBG+bSrAo
lyOQwgTs8rdyn0aL2Wevl18WHz2aeUTOvzaIRecZFWbQGGyS+ixp5IX8BmlHysWLtux3FuTRaeix
AxPurHIP1KI0RQlLPjsucLdScNvlWaep8/r+aN5qkdWtMboazhXCymvHSbFs8AyTKXawRpNUSOkc
TnvRVzK4tOL1NW/Q76+RjPpkiS9mZQDEqW9pCthmEf+L23cdcUMKbOtWIgAiGgV9iBJaFe/Fq/ZY
zyx6eUOs2Djh1kXe3xPLVoq3AALnmHhYx4wdk7y9vbMUGpEytHSH3Il4K8aopHRsvhQeW5Dt6l3e
J5FZpHf6lGmTrN+eTnEsLZmRLb99ksZpgf86rBfzrZ0x+5p5zkOy5Ucyi5IiaFKces1RdIfuKb4S
Cv+BShH0kLaxghlITsRSezOZr48SfucvZxIOt6mTI7LXz1AV0NDI6BSs005rPoNMqvcOshQas3IO
O1Y+vMtnuoOTDShZF3ktMn+S2/CKRllY38JwJs6VliyPr6FxeQDyqXjCW6Hk/nmN2M90GRKSQUyu
eRE4BrGO25I9wqpGj4iaGTEMRXjl2YF3rn0FEjbt7+JSKoze7QpZ3E9EUYSxVIxVEPqxg2Kz7qUI
cGgv/xsIOsosCBeH4ZyeFPYjecXIQlemngmjroAuCp1Vfd/7YNpQ9KbUCXqC7yUKtQD/YLwpFd9/
nZeaHY6EH1s/fzP39fsq6hdXRwGksEOb599UIeQ8aPfur8vWnisWctiCxXE8gk1gPj575D66MV28
d3Q9qa9qcZwEIIfB+9Y+TKpYvF20kNL5DXJm003GurtvU78kBIX96LqnQPgKQla/APpzx39VhZsS
FdkXiFw7/JTCY006uHs0LQP/KJYRRGW1jobNJC7jZflQPHhXcN8O+tvbIQJNgOhXVTyGem4AT5Le
wCFVS7C/xHpPHjkCvm6s4eWJbbtaoeh6sU+5It5EI+YeiN8JifvGjSozO7VyXIHWIE09DG4iw8KZ
FzrQko2Da9+jxnGD+ze0/Yltx6jHyBnibs7ssjXo4hCOixH4IcCxl3s2IaFoYEKr4OvkdqnE7dad
hLNCv/df9iUvTtdnmIdLFxRupo7DgMgyV6QzmzAU5RlCKNI+WTiAgxeN04CoMjyHqNkIEcr0aqQb
o0mk8DMO2Hd5kZ9B3cEZ0fZtAT971rj8ePdD6cSBSSe9YrZIYDg9EhYSHLh/8oBrkCvCj6Ci72MA
nk4WYgMPAodG8hI0m1N+6/2Ae3Zln9qBSN/rGJLv4xlwjjx8oc1qFg6C5hKVU3bgt3WJgXtzb6xC
zNxWuSvJct0xt/YgA0gkq0dWCKUX5kc9DlTOODoxDUXNk4W2BMeM+hiplzZs8lk+gLFbWvFZe9b1
NvxCZn3ZBLC4tHOjvubcx+9xrAHr2wsqWnEyCCUO/8S6NMjUKOsJHqwexrIwk4i5NK8wtwnNPNG5
MVI1LJtsywbnV/Mnve1Bj5NggPE1n9Zyh0RyX9dbbBXD3Ebwc1CuXE3NkkJcmA/JGpkLEBAxE7bM
tGsxGBmdbgrfymPvgQGEw+UZDs/oUEbnWzCIhcanSYBFqSdPGCu/f3On0QaHaI3xMD0xUbnguLnK
hcF9ptRpHaOjR8fa4CKCgW0rt2XtqNZRd0nyDu3Q2d9KyiQvw4zKcr/k5tZuLPThZqokT9UCSBnt
tIUC44Kl8kteR49uoCczaGsfb2bkzBkM3YmEyht2u5r1dqa/jLLOv9rwm9AWs0ecJvKNZI04Swmg
kJ4C/u7sYgv1Z7Q804HBnHvTeCpZiyLen+EkqPRl84gkB5bxD/UrQxTVuzRncBWQJkGYeJBgRsM1
nnSfXQLdzwUMd+t7XuLKEeqUok7FFHMEX4W3tvqlp519FB23KRE9k1G4vBWAkAx091NgOgCA6LA7
kF7Md0CDzrUuXs/wb9h/qy8cZvDpvda2No75XIquOLAoB7Q5sD0MIBLGlPhYFz2CyYomMPjpST/y
qlieRziTlk3KIGx+8LldfUavPQc7YiFvE2uLF6vGsNwzii4Pb41Glk4bcWlySwf7I5GNqS5hrtFs
n7yx45RJpDFE1/YABMyDwpwV/ByiHZul1Bqr5kUfB0FyeeaVFjISKUZj5bSMmREqN2iC7+G4ufhk
1dx9FlHHm0e4jjwWh1wqDww1VMfgkDbviNx4nj4g3A8GLj21opYwXDkRSNBCc2UVwah/Zoafxs1p
C6g7j+QQPUVyg2lcZKWLZ5yXRMCiH929bon6m+40zvPtoo7Sd/amW78H7d8cXpSrrJ+Se1DU8Z/o
vjjc6DUrlxJLH6IUVVdgjqDJYLWyidI9eX5/8xH6P7Bvr3Blcy4/frtPhgmsTzUiHEAfTXrtCt6h
WnmHgkHPeescbuMME2d9o5OA38uVLAbCRRgBsOp+7VTz5dvn2zc0Is3CiL/JFhiaQVHs+wjAeo+Z
kHS5chg1yayXc+3JntvIq/yC7lZGgTEnHG878roHjNzJBLy7Wg0JJuLtP9JQu2BlgxkocV2BJQqa
gud2tCMC3vAiMjOMH8ALPCTjVPKqQNJMzrnNATPE/331dxjdbYWd2x2v6WQTMSRlVi4IJ7k6jlaK
MjzJMXT+0XEGEigLMNtev9FeKFsd122ah1p01eoR9V+8vjZh1lgDoaY5E8bADlueycCZ06a568MW
KmfNW0WL0srWIC8NnQy7SBO4okVtkr3ha0zRnCgjAwRVxuEElIoRS3bzt6xthaF/wEwzQZOv/y0I
Mz6fQ4iAUPXzeGzr4+YblCm08JrXHcbTr1i/PTOwJ3NRp5GOsS08RkZxz9U/z6JfeEMK1jW3qMho
bBfCWEiGaY87jgwkQ/pGzvxlrXXVVHdiUqcQ/VsHCkrpp1b4sspGQnARWWSTzWfCmsiSoG2pWiEm
q6oDLjylE4vz75AcqfrHOO2U8k2hA4Ob+qKbqnMqrxLeo4zZU1KXXGDgF8W5FLQB95tUjTg5XeWD
F1PK0K86JJDx+gvoDUOQ6XXeRxDA2RHuuT/qid+jpH/w8ZS+f5QpyLChvbaK/LYQJWML0qoWqZrc
3Ytm57di23GLD7n7EK75OQK+2FWgXT6KWmcoRacbYA7i/NRlZHaLrQwNeIaREatgHd2kH8DEaPfm
Y1QxOZ/KSEvQ7GB3ks/0QdwbFGkVuXy+XO89Zt3VyEeglP3GwdGeqSxitw/l5jBIXMFvEzL6GITN
wIVHCOX2hJC46+PHTlso7VsFZaw3qR1Szph/Qh8DgRO0H3cLxDKW/2fmqQds1hltIA1PvHf93ntY
lJKrSOoLfEoGfeYB7Lc35XbRh7dLtChrDOj7Djacdb4eTVYLXe/meWwZiSgTf3L9JWS9/RsSXNrP
Kgl6aUynPJvXHR2+dMVDsV3wp83/9LHnPmv8pFZ6WHeags+WRQGgbBKDWde7EqixfyWAVY3QPeWS
5RlOam8nAjE7apz3Z2ArR0CpVt7SNNz0RJBPNMRxuU0khCmPxK0xGWK0cYmAPg5HCqtsKoVCIV5G
nMxN79gSjQCQ6YCMD0pPjHdkes/2e83CM3zKuIJ9m50ATSVakb5prAemLe9X9Jf+BO7ND4y3+cm2
PV9Pdklje3svpvV2KKKsAqH7J+BNKQQN2VxeBPuGElGFA1Kqcyk83h3XEE6r+O+vgPZNj2mA55xU
h05PTK4nxiV2YDAltta7QhGmardyj26iXah6K8IzPHh5VRZNHjv37jSp1ehuv7sIeA8QgjTFlYTr
4JW4IdzeXAdFC7aUQB8m9qv+oUrqFUfWT3TaeCRK0bMlGXcqJkiECGa0mam3xalzzD956GmPfuw9
88KuzJ0C+4A2F0HBuNPHBtKreMyjKecrSsfB0+80T8rbrH3jl4sgmtBKhBlyWhThKHZC/Cc8SbQt
VZl8JxLKVcT0piivJ0A9oRirt5f5J89W+e+aAUwSy8k2qIg7DX0imM3zCYjTnGAaUh/be7qrahN9
pYTb+L/muY+L7eAzFf/vAqO32mMzQRFF1VRBnIRkmLugSBSxuv9LRyYqT25Jvd3f6/H8PDrqcztu
e/Qbl3PD6W4oQ65dj+OItZsMDuaXQLE44OlIwFJIQB8iNZ07o5oSdkOYH3gljXVO5TF3fk2RtTVq
e3upVlR6w9xGY3/Dah7KEOM9fJeRGnHiEFmq3P9U2ubtZRMq2ii0KugU5CBpoF/6lAALswppk2p0
UqHPbR6Z6WIGsUCx0kladpK9gwA9qx+zwexat67OtZwpAiwg+61eiuBal+XXYl/mDQait9J/y8iX
QIq9YbcqN6hKjK+4MEu9TSsZid4qdWcApkVabjEac5WmCVXSeu0oJXTvh/TNzI5qHvgBNANiNjTR
RfI4urOYLAj/FkgDgFSu+qB53z6GzD68nsSgS8GtVv4FXpcHtANLt8Nc4Wzi/51Bz7BIxsr1I58e
mCjxUPOUrcjD74iZ/tfCsVMiZYLQxTq/A7zqN2ZMVvW6mgSk2b3WRjRgxD1Knq49SJVqxzgsry+9
M4nX5l1N6eoKYVRcQVDlTFZV35Bqx2rcATCS2cReLYZZfv5pBXoq+sGnKGB6T1Vh/UdSfDkle8s6
TJatbflKdad6cNx8kN44BiGx4wCXn1J6C7te6YyA3CLQJWXBJQYfgSid7iDoJAlHPjPiHD37+GJd
31vfJ9r11T4M+9H0L5G2HkRJIWu+92gjjQg3HX4EzQtHAzxuv2JwlzfH7Q/ksSvPpDlkxnYrmpQk
OMYdeLJt44+Vi3Sy3RQRXzvSQIymOPPjoeGgIRVxIc5xulUubbVCirzUoeKUnEiNDsyRU7OTl3ov
S5+YbeRFf+wHs4haasPxziU/qdycvJB/vdzmlA4tVFTuPl1j6m9riuqJgVbkqLx8H2kN6hkbuKA4
Mb4G4afFMAKgfwtnXu3Y8wAnOS3pj/1ycyWUyMsUV/lJLim2M80KqttM9/r/50ZCtKAIoYuvBcvK
wDzXJCnZINZLgSnhtLhOKfOP9aReYqzEkDvU5iF7AoU4y3haDFpbTBouD4/wgomsbP9Lyu3Ldt1N
sRHTjSzvXR7muZr4ZjG2FeQ8rBKgrxRVhXj5X4563kEHeEdHQjK1R1CcQTzokW/4LkngL58c4I6D
UGbQrgmptLCFreUL+VLrE4qCVA1xm9tQhjs03v5RkkAAgRWDpPGd09d6szCeW1lJtg0/yZEiBL3E
t3xGT4VRQX0Mu4lsWA8zDujhGQAz36SfSxbdAKzqdYDk8JxbB+btAOf0gaIDZZWliX7wA9wyIEU7
oGDPnvsHQmqzUktaCr8BSWOV/GCnIEGWfZfTv/3K49inQBsg2+es5r5uYvXPTIw5XzYvf/YUgrvT
2lGj8pnoAonjs9irx3c5NCFdGFOHJ6UHKZhuIcxV3GfT3VR8sV+6vzGm6x1OYMs6tbep/RvLfWIP
3SY7OR/Py9DbzVYZY7cI5FK+9oMvvuluWz+1SG0dChOg58L2ruQ+J+BkWWyA9+sHZ7WDYhsHs5RG
mn5tDvmGM7gy6aSbeDn8lg+6LoFvCsxi8VpxavE1a8Lo8maf5kzn0XQ3OlEPbiSBVLETCzcspvrY
QvwouGoJ6eJPhGeKyJMYM/j+HMiDNwc5hIvthwZOXH0xK1gHXBIb5Hz9XtJPk5r0ruHET+vzB+EN
q1YaQyNHKWrY3O2Dt4oeziZG5HwW1uuD0H4MoGiDY7Hyri7zZC/s99kboM+RF0RRt2QhILxypcZI
Bd2U6ua+HY+yymxRKqULyGeWXH0HpH1zqCMJIDCOvMDmNnWrnkgMnBPOps42cnzPV0ed5ciC4S0a
8HvA0sxix5r0QO8k5bx6MgVOyrkc+oFsLAFFOnoyo6pTutqB8a1hQSuHJ99IoMmAesX6kE9SFzo7
/lsBHRZEO5tZMHu0QxNHuLnbbY1JEIDneJi0K7Y8xZlX2kwjadanaw8r35qHELOKl5VsByIjwRJ1
c99lKse/yE8wGkR470hE+GXXu9jCx2rpKZgj+hsqWp3gMu+opgLdExHpy1mt6+vhxHM3GZj0M8n7
WKDgk8bDN86uAlltBRxGY57ZUrgBTJzGt9nqu9/w1zBKIrCBo7fvavE3tToolBvzzV+FStsJN+Mi
FhsZ87u4RufejhBoHmZVXQwkcazhK1j5HSF5jm+wUhyjRQIJvnMHPJCI4RlV8WPdG9ZDLd3c7MJJ
jw6ROws79SY3mVW5xXlSrgvm6mKRDpBfW6QXRXqAK52CO6xt6WLBEUOPVu/APN4DnBceaEW6MG6T
WRHHe1Wcp3yYHeAUHxrdwc1hqj9dRAxv0PUVwm26CPSX4ZFzHX29SI8LLbly83jbSUr4ux730uhQ
T8cWWqQTlqBa3pHrzfyZIOYW420jmfDeNHMGQvHzI35Mt5SnMCVyfimFdmh54Duaxdco9Sfo/Kl0
kdnwK+AS3hEr5zdpMLmJJocKN9WenO7n+bgVO70riq8ym4kd1zn2YsmCxDnvmA2xp2gMhaBj9khg
OdpY9G5G4V3VNFDcO1SrrEPHk0Ys2pAexh+uBx7xnjQ1AgJ75I8S8gIextbPgJ6yIBcTiWSVg0GR
8D5Nd34TwrUg290aipmcauiqCcCD8YWYhrsnapNU0kMssXH06Kz6eIvSYOWzLpJf3sbO6Vb8e91b
S4/fRfSPjPvQ7Ql0R0mDo1bliX+RJxKBwQFjZQW/DaLE+iiFLh1vJO3mSEq266Ajzl/Nezd84sq1
ZlEgt6YMe9hAiZ+SkwaKSGouanNkZB6nzzdLpH1yiOpVmqJiadFafZ6G+8vK/J3rxEanbBunpBbf
bvNCtiQAOkpNlvzDFAfulHk64jNyPqKowyWGGWW01RD2qAefwUSEWDBDzeHMgnYt164gEU0rU2RE
AWZHyz8bFpDABhGofeeXB3Y9RdJNL5E/KXeQsAK7T7PNaSkGR+8gZSNvE51AWQ8LIBIcFW/3x1bW
D9+1MulzZs25VES4Uwk0ZdI8rx9IfGL7YAokvWaOFZX1/8vlWoL07wT2qNpEXDwwnNFiJ1hPmJ/e
Z0Qbkq0iH6u1VUJSm/Azbx4WmfbjY384K2FWzCX6sHa2ej+YZvI3pVQKIZlrAOiU2Moy6KPDWN1f
rE4JLraI999tTkMHYovZA+4HUNAz13fR9a+ryEttgR7hpHL9M7C2v4tFLdNKHb0sYWjvoZaLjYrP
R8AK7zmMiHcanwxZ/ZUeLV0D8z628ETxwZZpd4IIQ2Q8eGgOwLFxeC/ukW0Jclny3ZV/R+M0d83i
cVbRt4b00gG/vN+/6LEUE7EriaYbRSBhLiqsiXI0C1Ci1/cBA20fMOBgT09Zvr9Prosnl34tkd48
37Xv+Z71kBaXtq4Vi6/eXzWB/3nFbSCD3Slz3mPhj2Z0Ggt32aYg92bzkyZqtFhd2ex3ovlDdWf/
pP/tkTSoF8IAc/5gyz3gmy5QJLPPTDxCfeDyHfOuWVfSpDTcS+TikRulYRqRP09M9TQd/PlwVSJP
NCVXF9zMiT6bA3FKgTi5P3mMr2EcC2j6x2njKxqAgrYLn4vLCqaC3OyGMOZV+N2XK1FZTIOXgUH3
qMx++PgEmInPwyjf1LWxDDZ7zl4o35bkP+9Il2iA57kq9nfrd0xKVeSUowf0h1LXpj+l+JL8csma
rqoAr+yvUds+BJtIQmFyNJDZjMvyQJ3Ozr8dZ3F1bc9f+YPRE9+aoI7GQUf7uGDxuN0uEfFyrE0d
qJv+M9C8CgxrrH7J7J53Wi4eg0tOXkslebJsd8KkZbtwUoNbrnsLeYnpedG4cPP+GwNl0aucftbv
neOIs9Hs5qUCmmLXq1s5DQ1PU1+bc23kPAPrzPO1T4Rw4MTBn8BH+daK5eYrCgeW8vhDMeuGvO2Z
JYpCbWlFlfMHzIIwRDccsmOdHrnADZReqSa6vJ2cjRdo7HwmiRaU3SvMQxyatVMeAJ7EgXJA2Cly
ZrMxLpFy9Q/qQKVsBaVvJbPInT4xr3i8Lmcat7jSUzgHIYwCpEKSPKTFA2QrXJ7N6bAvSdRmcJWr
c11sf2lVR8C8jMfyEuEm77pmZ3A9WmvPJkAMxYRN2koW4cf+RfqiXzhwq8/ogdGQjBqg/na2IJvq
Ijr4r9scR36raonlzyLlAyWh/rNhiDKyp2iFd0dmI/RZNerYItOUdG2yJjQniZVBrsUzovt6C3QF
g2pCskoZj+eqQPQu9uwDwtZfa5lSV/FN4t2iBHoi8Ru3N2ai+IeJd8CNCT/BofZfdu1qTOaBmAyt
P3FtPcy7l/0njAkqtUZQJMHMTlpda72pwrp4Mn4P9LfAOR+rKN/rBKRR3Ic2IXZpFIDwrTu4c+0w
W1Bk7r6cext+gVouN3hGTVPePHos41bZnNw3ZgfW3ICymZYAQBbAdB7ux7VvgVx69nbR9jcabZZn
jvQRz2/wKB11/RKXIFjI7aCw/3QKRQZ68tmUmhtN+xOiLo3MZ1sw8RBpRY+dkR1XMEoTJ6IySCee
byPL7rKtuXj6X2Eu7A1MxjktYB/CZkn5M5+3IT+DmKBtUTEy9gPahkUU+WI+robCDpvZf+dGuV/o
+soc6KnTGsc2VEDtXXIMeQi+4LdVffG+p975PeCRoq9opT6fRhHklIWApSF0GPwdYesNncOaoK9C
Ihb1EYK103dfWADSrR/hA5C0SaZ8kuYdA23o7uH1tdQSSnAOjdwoQ96d8D8TK8Wac2yYUOkuxc5q
TrVl1fwrp5HB4bNxDh5ygDvwJ/kGy6MR7INBBKbpTHhXAsycibMJfUZ546yENcT2U0jtdNwZniBg
z46m0gFHbxBcyJqoUqSqBhR4pJxjjJs/nnHtAjzw8LQ3d25/junTQXR250cPY7ymDmvaIss9tWPP
8nT7e9tG+biUHYIvZq87tneAynRPfg7oHKsxvk5jHth59YzXLvvsHKvhVCQKHy2nbWbnfOBBRtob
CFoQeHpLiE1vDMdcGzc95VQX1k0CuaNQlfWWYn2gEA9l3J3sov1/J1gDp+WUtnJ5/lqMEHKDCfVu
JaZtEyIxAjZE8mHhH6jznbCIsxL+sL5RXTDFumlNhOfxW0SBNALzxy1t2poNkGigtfc+ibMbc0Um
A3Ut5Os84NfMyTN292M1/95/0Oo3ZF6HYwERf+mUSq5lSN7Xbeaxafpc87G+eNzoE+8fWyuB9eZm
UG9rxPiViPU8KOST/L5uB21vCKwHsS6wd3XMKKxgyTwGU3TZctIqpUEcJ0/XSc/VqVbm98VpN7Dr
E9dnTiowtt3vOP9ZPA7WTwGrTO5/Q17Qa3e4Y61u1m/goZ4gTVhTcWiR46fBOfkgFlAAyS8oMGPM
Z32/ppnxATiAvFw+l6jBlyrYktqGwv93vdbFDRbTIpNFkugcwfARMBl5rzUlE0Xu+e1LJnGF5Q9+
12+7IiuDp/viQhWJKIsPm5pTh/oJgvyvMI5/PuQ5jqvQnCtg49u2NM0ky6HcjtjYBlhG/XscU8Mg
gPBEyRaXBXkNElVZrCs6SA3xSeCcoKJwGBuJdEPSOB5K3ZHZMZxUFMZFFSJnxD5NpKzepj8I4A6z
nvuUF9vSnVJUUbVGOp8rv+4hvbOcy668UbD475QaIF4lKQIhVn1LTfUuTVNm7lav8HRRmJGtoxVk
kCuEdWRgwWCxXLed0T4Eqwic9DJxPxbZ5GaqZSaYhBtqM4INm1t5ys/RQnq7TP3scaN1rHeLYcRK
nu7YsQn+1Ob7YBkXN18mxWDDKNu7eROVn4GEPFVurKtprwWEivAjIhdT8j13vlILunn80EHvzr0A
Kxs18Hdpczx9gZoMjPiAuGNZS4/YkkPzsbsJpPem8TrQNkZuTnLPVDMR8bp6jB55rQ8tTE7dSPsk
fjF3Bx33/nPRzazgzoYrkDEhEUnE69IDBWnYjUHdHZR0TNWJReO7zj1ZPx4MN2RP40/7wsEs2/NG
5oK6GXUv8CuHbadGBOgPxhBoHF2ZyjndSl2Lt0BtlPsqG6BSsKm7JY8giDqET/98DVWb4zyQ7F/m
wAEZ8hs+hu8mFmPeUe6Dqmh7hs6iMdRdESiPK/8pgDs/qHDzzgfaV6txGHXlZaaMnN+923LhyWnX
L0UbcKIqsPYrn0sDvbvaqVLwgrYnbNxSkLsTzyHxlVHhizyob0YHBqgfk7XdND4Tu4sJI9uengvJ
7cZTPVTxUqVYAOZPjcXNBjj2i+cDmMbjwwRiTgj1aNuqEZqXEiqSk4P/E9H2T7alv5gWH9mGbnlJ
+TOt2SQ10J/RVEd2wE/Gu1rhFj/69LnO/EyaAhJRzu+JJGi2zJk7h0elpoAGNO54o9Zl6EO/qSgO
T6Tp/pku08K2W463sspVkZ9ltJL6gttX15pbvmzELo3GYXDw8+2rqC6QOolf1PUjkERL9XDcaUmM
nfEvQGA5n2zVEqpoZgJgwyF6Sm9aFQ5B1lHETHj6m5esVA7bJ++pqgpULh9HpxtNdAVaeL/KsJjE
Gj0y/JGxnQkAkwY3MZw2wrDPNOpIXt6H8pj9iAkrvy8EPHfSKefX8soHvlC0IakV+0FMd2Dn5rmy
sjP2Ylb401+WGpSjBCvapZ6oITQAWauPl2+gjj2NchUfgeha5tuRZVhgvGUCHlcjcohqG24XQfdK
ESWBf9aySEnH+X1XAAy+nxJMvIklwMC4YM7/bqMBcxRbQgk4SHVoTeSc9e8ZOsvhwbJacu5aN8RZ
zznMCl6YXeDtyM7Ko83JGwsi/bAZoAbuYiWDBMleIB5BDEcgd4UPRPoCLIGa25Ug3sj/r/3XcP7O
+nuu13Z7ywSvR7BpBjNKmvc40yYPpKcn3RclpzIean6qwQh7e5iZXQRS3Qh5Xz2eAVBmLJbYl+ld
tp4t/+wURH3OuSD5jy6y1G5qjJBZJwPNVOYsp96o4oDRKJ0l59yhNRB1+3tr6418N44W49noKOBM
fCw1pMShRA+USOkkW7WvR3uS2TTRqS+Z5tCBdUcEBlApF+LAASeXoyLs0nfcKLWO9ee1zA42Aaq9
XOcwWKnqC4zzQm6T+iejISq2hcE0hmuh6PF8QuRbD6ROH8+ZZrpVE5rRVoFwLmHs9+imMve7bsn/
cygQ1TTRtSsbMvyYXUOXJ9G+x7YBfqwpBvXudwM2uBCXCmhKlgQuwskCYmz4EsxJ129yff3GJnCc
DjxhEOBQY6WJ0Fa510LQLrrlQLUAWX3h63IpRsNWY1rgfuH6T5ZAVSY7bXntIHonA+/e3Yiz64zD
DUfsIPeW8PBcTLnuh/Wh1NB41PG8hCJ1Eaoi0KUhgPAd56dPzLDlkZB4bPU1BuZZQIiQCG51Ep6n
rnACfBK0QS8aKsyVvnuAiFq8TXd98e4Agxc9H9apjherdwIJReJEsD6t8VlEd6o3HbO0zTNiVHnu
yGROt9LZAW8y1yw8fbT4xR1/lgNct3Tbg5+qOwtXWd8GC78nptE3Ees/eL3cx5XwvqM4G+45TV6k
vIZPGt7auhuj5TwvZOTHLxwvsFK5LjzU9rZF5w4I0AaNsPgBOpxnioMVgm0mtNVZ/QEMK0zVwbMI
jHNMIXny12szSXEKUg3mIRLA0UchP7upXhqky/6Ox2Imk0VHVvkuXj3L4YH+qtKh7sOm/w9w/RXY
weeYFVfi4X59+DM+woquPYDM/Nk9t9ZhAlqUYrtSsAk1pYN/D84i6dcdwEQ+jtiO3UWbVjpdRML+
OdiGSxAXo0Wa5CMl416+CzdR7vStVmk/6qnx04VnJA31x/KGCt3k9HaSXLYNY3Y5Ju++Sd8rCuQ/
jhRcogJ43mj4t2ra8OnX4XYBPNJO35/MryeOmoavmEPVKj1whp7XeDZxVfcrxPOUnfoLM3O9kJMN
hFF4JcLc1kkTArXIZdeAie+5kmY9LmhyaepNuWYNhjXv6QUedpjMy3F4/+09Sag/KnRjB7cmxTXS
RYojmzg5BBAleU1D54H5Eu2AOof4jA1AWcXGnS0GcltwDg6YPQVmRAtWjMeLwsSZtF+ftgvByW7k
7lM6Kk7vWbH+VKvgBnvVOM9eZHC0uWDfit7FQEHMCEr9t9Ilmh7ofhE6jfahmQjkfnB67oUa2uek
H1CIxGUIQ0T2O6ygMOVi+GvtCeks3wFc/OsZKoLljmS3e8P36ux2vkbrIb1MfpYFostlvbjtclIj
gG2SR04Nrkx07T9Ak3uDgvTWplZCDr7LG47dm0tgG3VN8m+oI6ncYCHFd84j3Ia1eFBIvlcU7Vok
DbFHjvqeSlOnAQTzwuVxMonJc2VWVVW6LrYcZI85WIIJPbq1ixRiifJoICTu7UHPZvXhr8QAM4bp
bobzNgIkRNB+/OhXzRqZ+mGsVnwsJOfba40E7bpeGJQkLrh4dh69fEp45DObZP7WICW7tT016T8T
ytJrHz9mlsbk42TxEnZRruaUeT+6fz7hUsvsML/Tavwn/Folo2JwsTYod884vxoTdEaXT3XtIhQv
D7Vm+NcrD+lT0ItKKxobbHhSrKMEq12+V+LSyoppbnUPL6OtjJIAy3aoxA5rKs2zgEwzQC7TFGSW
6lJpwr2fp797xOaDIGign08lSK54vjnz0RTFNtmFAAMIhVnUxe1mNFtc8kwGlY0hOvvxFeaxvVIF
r5fwFHQ3RFR38WP+dtfVGlzpn6vtb6jwZ3rva4hXa7KLnSqZeheyDfm/eC3MmmJrunGtmwopnulb
D5YIskPrad13DIoo5LXG5/ouzko+KG/H96bo1o6xpcpEL2jUb+Vf+KDbtTDj6dvpnxIS/o/Y7A7T
Lza0DE5RvaJvyhKrI/v+/ohUus6py0aOpPuLdYnpmzYoAoq3Q+/BAS9nEiXpalh2xvDEa4sv0E1y
LebMP71MkdwQGQseY5je+Htqc3B0gNJoEKWmb62byfKUio7iYR/vNtuOr9MuQCJFZEDbiPhT3GxD
Q5F1DxmDxydPw9zmgoecose4gtIjFNobgadFLWNRMX5ZIwaba9FJvduhAA+5G3mc0gG4dWvKK+sD
lR/GiBar7brevE10hrmQrnAhIOtSaXGJgSmc+hZKs5rhNLqE22UCj8v0gkzEkrTsK241/JJzoSut
UIZFxzSZ/pFYH2cBif5x4AISE+hZs2mbkSVJtw1gVOYtWeDBVoburNf8xINIQmW7ovfOXkCxeyuk
HK+w2igpWhNa8dtZ5Nnqrsz0R/gtSFtb/42AXYNVkhjFlIw64FDdDMbcfFrP/r5r162Wrhsnv90C
yzVXeELoSSsYyMlPGe5ucYt033GCgEjF1kJUwzOuDmNdh27gGP8nsyBlvmQhNkeuxwpeeh0P+Ytf
fnOwSDby1thxvy9GgNHrrUhu5eKupfULUiaK4ZfrflqkwOHou1Vo10zTuceAeaItc6F96HS3y/UN
r+jfPx+PbY0sh1Di9I7wvIWBKfMdpjL5+LYC15jXQbkU/Kjcw548Q8EqpLXG/c66xpq8h8wld0Dj
bI+PNCsVBgw+9F/gz85W7xhbxRKmDcDc5dPRWVHcnu3C1UhuJTZ8S+/blTZVWLNOSM8pRGzAZWTW
TySOL7oAmLNoBqj0iXqqDSGpEpvmI0SbGiunPprJnpTNu35ZojyKAxmLokv8vg2RgmnGp4BVsEZ0
QzeO5J0xy7pSVNasR3/TGsB0sd+9ujsoBj/HR1k3I9NZQVyGXPfwDVVc3R9CcAEGK9P4WNezqaXb
ahu2TLbg7f5cIngTJvdo+SI++e9DJZudJ1B5Gjf9krLFvT/L4UBbxzzVV5wrFWbXfJzdTMy/z/Ha
l5W3Y3htBeEh4Ywyyub36QskwptMHmohSTxo0lYCC1xvd7NeMx8mSUS4Ry+7WdcCbXYJ4SHqXWZs
EZCplTiZEzYfLjhFoyD21uzrAf5Cv4ryLbx0qIBrU2pTzwFSV1xWTZgKUvn1Uet1HtCs5Dij+dH6
bSHC7eU0vS/Zv7U5/iO8wpX9Zk5pVUBcE2GPOf8WH3zbR5ojO/+awJI8/CV9A/60n/j4Wr0uYgcB
h34hig22T+j/CvqslSz0W6/9gIUdTKgezaieWG4S8Z8yP12LRtCWtKu7dyNaf1cYnB8Gtp2UFx/g
UngtHy5BpkxayXRdOXJtlMNX2EcU88+/aCKc0zm562fPkyVswJMKhqyis0NxAnZjdnzVryJ4vEgO
ESNhiFajgZjR1BE+QfNZA9/TO+k8VuMnPqQ01IxVENMnFE8TqgA3RpKlcFgXSgZJ404L54tzbkzT
DErS1t1Eouqt3xbMA2jg29czUtINaOyn2VpuMa+a6MmnN3PEZd/81xwuI91DqkG0/qlMR3QfE82W
3LnjsUV6Whr0MaI1PBRuxALbGjY6RtCKxuiZyxEUE5XN53yvu8BY0XkZz/GXmhMLC9oCQy/pO/LX
6tN3R5lyXh2kteVgW9rFrg6DjzLLs2O309JMEKKRj1g33EO6dYGK+Rt4dk0uE5Ef9mlAjfsVF//8
hOh8cUcDJTGvvyLVptnrY+8WTSprxLdCtfyN8IiR8jhaMW5B073AtqJkAgXiqNHXm0YMKx8kd9l4
BLdkYz8t+HbpGmUXvf1FABNdT9R9n4LeyLQRU4fo7gci3OiuxHA9EVSy+5Ox2W1xH5+CpB8yGi6K
5qmRn/Wunz3E7ir76P2bxVB4tHr9LBIEA9YhJdQP+wVsSqCcVaPXOfct/6PL6Ri1nwI0wzRapDO+
DIQDFTYpmsF+nlXocVybQi52ejfieTLfx8Y3F4yQeH/CHeDsO5Y0xFj10+VsgiSypu4AII5CbOwi
0JPDL/RuEOl2nAsi8wdOmez/1gGTXfz0a4vQl1HZwioaofUTDa+4XHHAUUOHaWT1mRINdIxiqGP/
rpOBuTGq51/bYyncLo6cQjNaPTIAiyieSHRhUdoVYYThGjjmA2yMn3Akmk9pNOXCwvaPPQQGMcn3
TBVSe0wQ4pwfE+hI+ejcSCVFgm4KjyhWGClxj/DTYBHi/35vxTJJoUh+/loNnWCfZh2hbVS9GnVS
gR9AJ4VcYG+gBWo/Rr6fTqcFtZ45WGxvTPWd+FrhrTzGaTegOmj21b+wcGnz5kaGgedzqWFWe3ky
6wFtJmVGL6zXWaYqMs8uOEgRBAleAp3kj3Jb0M5zSzzlzeOQS6ZcQ3D0nLI9RKM2DzHY9otwfdIP
tJpNXTfTF3PFMjRg8QyL9IzawgwEU6l7lgh7uLq8lzCY3nv1/vU9OuUgBOm4viwN0JLWKbwu73+h
4nvyqhDo6ShSk8Ap5IWGu1vSY6TD5agGEJ6JzsEGFmhhnzu7maM0Qe3Z6auzgXga6e16gOd5Pxfy
hmrYoZYh5XwN/vdEciPRb/9EJn/2HqOBECEGsPo45a4UmbcQUStP77L3Dv7et8MfAfvaX6i+YJ6b
GySgM3gCjWuEqzGTW2lANxYOu25MGtPKafDeC5tiNCpVcOunNsi5IbIvERjKwtMXpIVs37aDwHQN
nCvP1jDuJ+7Iop0NqPFqbWvUWr4FnPp4+rFxFj7sHQCpLHv5sfl0KxaNcUwuJz2yyrtVs+9nzz2p
tAAkLSI1Jkl/pWX1s5zWley5o6V7MjpX8ZhI9JJtc/C79HWSKVIOgjZGpHbEIrwLaMtpIbe/2b9q
utIQcjyog6jo+EjnHBZbMbwz0Hq40wgIDkeGpkw07s0VJRJx440qiLhTR2LjBuaePg+puRNVSMd+
pcQyGSZ6PejClqjB5cOZ9mvxW/7BX04jiok2oNLcxGc8UUi0/YfZsYLkWT+wCCKejInU228Et3g8
5UEcYt6hxbjGiDLxhsoNm9YWLvg4UwFz4r2cANnZDkeqaEsl5xE3+LW+S1tEDIMViabwzn+9xb9U
DrmE9CXUBTZb0LjqiNRwjoSwV7v4kYsXo/jXXDbnjfCMDRRMj4pMwklVRJqaL7gF5gMQyyX8La/v
pOo6OzNFnUNlbXbD9Aqnf/6foCBCwZ5B1U168qLnT8P1KbHOAFqKQpfLtSeDBAA0JGspxIVJuTVF
ZyuruGAPmhAn9V3umOW8inRuMwt44348EmZT1TKmc1nHFk3gjh3tH+ifXEEzIcn10g48WPoAOAzO
xSYXLPq/wMmVHlcLyEM3UMnNaZDX8H/G2vprYEtFRC2pm7tq6uiJcq6BeegZG6v97JAqPz5pWH5i
ina8iUmhRNzgb+GEzJm9EZh6jUSm10kUqZIGeSi3HaJHmLV9ohSzXfkhS17w3KJ0zbEEPjXZo6YZ
TZUr7MUfThfY8cOTgeG70b+lNChWta7EwPeo/7kNG80rJzEsKW6THkLVTMWnFyU8lujTPTm/WNlM
rE4p4dX24VM5iHmpm8KAStpitQQmp3BToBN2L9Jbwur2XYfcKjHzV61nqRaemaK7H6yvqeHn9J+Q
86Cp/znx4x7L5flMBeRMRdwzOUZGh8Wlse4NBVluqmJcm2CpWLjw4zXmpMDcPZJ8ZCyso7jLGV4x
eG5C8WIRlfmzZINS2UWDOXlQjjVnJauvXHMpAgZBz1Uhb0sDfE6awXtuT/ed46eahNzAuUQVlJd3
IxFtfq2RVGsqpuNvDRgMO81/ihWGD2cmoIAHoh40scF6HfXgl9JuXLVPTZ7kS1N3vYiQxE3CVXbW
TmNZyPiUATrWkwJcwFBaqhxM4Aa8Pebp2n9DKKdLfosNrDVQFysY6J4SUf/K8185dhb5K02GhSuh
dxmRWMiHI+8Z8Ew91jY2GKVVIdrxOMdYMsA0nKL394cRT+DKshx1ujVKmzlGVjFPEXJFHxxvt1xm
VMWttsDLy2pp5MuZU/Zv37Ej9gMkeEB6fea4lpPig9zjwEHKvbD14yrqi4wuY6B2h6zx96dVwXI0
TevmEWNATcRyITNuFAu6PzeitCdWDHjktcnNlY0/DAkw3bjr8iN+trhlcTNQKTAMAes0658TajWI
LAFtWiZIj1vb+IWabAx5Vt5g1il6W4s/3Wx60JFJ49FosL1NIIK4RK5R7BEeddyC+P5KJHpk7Dwc
EhiSjEX++8jnzopN49OzkWOlTCpr/oSRkCwdUKc0yilHAZWgegarqFb/ADvrMFTwjANHcc9Yupd0
yLaijWzw0LMIfGJNSU/jCCetM3Sgvyyj9Sp264Nt9rGNhHjNdfUHFAgGdd7qZjRqtrgBhXUwuWOd
kpS6WW+3ZLBBUEz0Qp/iiBHtRkPYvMcyOAxZCsZam6iwJTomQ8ozOg+mSqu/1LOWiYjZqSR1tmuf
w65iU8IiDVSkdvqRr/HqV65rDYNYgS9FvdHeDjuUICZHYW4P0rd3brYksSJAb9DXk7fRhZxcxfxj
Nhbatqh+OHXxJFLxCzT6Q5i3q19AqFiLxVL/h9JZ6XY5tp8N7Z2kimaeA89xHgfq4mTVSRVRvZaK
0kO2oRtA0A+stMHofw4Be0W5teMBQmbdcYsl7Hm5RpRPzOfgqjD1k58dQEkaiYuNCsvxY0xOGu5P
nQt9OcNABhjMLKrmanI4VWfEjP2r+ZZnZcT96XtJpyco4iNTWRgyobBiUmjtebyCi+1ntMnPmUMR
l0i2XYazpvYd9mkRjM5joRpGSA/c0XuzIW8bvxEWRVmc6HUa8mnBF+lk3VCZT/3poM80k35EGe8c
ciqxvooA98Y3Y9+4qwU4BZudNUwr4NpdfE/thtOKzrcJyEq1Mu1bkIpXtfTgcmCQES0zVUqKIpn4
YYhGwFW9IW3QWWCDafLMiv8LF8CKDQS8zGfc4hBkGSQTuPJlFDoKQjelG2m79qLex9e6p0U+TLtN
B5vrsNKTo69Dw3OoICVrf1HpEfUR9szHfUtf6kd0dridFNzqbaSA0liB0uxbqC9lnZDeh+uavAKe
LX2h7TpQK6fIzI9nbLePMykJoSd0zbw0ARXPTdrfETdt1LrEKo4UDYmKMMU3kuKOO8AVBkDpHMQc
vbaqVxOUCX7IQjnmpMKQgh2nMOqxEDbSLoR/pIhBY6J/fOFtQgjCW9S9utsLM2Jld6sDO9ODC9JX
5KtN9AGnKtOIGZDuLZ5A0DzXjRwSoFHWXnIBbrRI7/xbh9klbwGpHABJPlRLHU+o4ZjN8N/ZwXnb
riTQC1XoFj6D198/95/zdLUWH307wiDWOcVt21diyBw1yoifa+0TDBmGmBizQHRctwpaNmxkgoRQ
HsR3okYAdNJpx8kiyruCkhfxRf8xHJxI9rgAX19M2NB0yb42IKJqueQGiQCyET+mhmRFv/WxwB4T
5R9hFFUT22bDYVS2wVAJ5cLF5BcTA2N8y4TYUHkfSxC2WxTIo60xuIDbuLI8y59wMOQ9geohWNKw
PAbPEuWG2ajKfQlIYDo+yVsCltS1vxxUCnxaDGlxlJkGN3NMFAI47audXBN/cY0vTga2WanAY1Da
h7DJezrJXcQKPYRjLaUoOEZR+moV6eO4a57bBGaetVjqfNDXoZd1NijK+VKzBtaIKh2Wvk7IP83l
Z8WY4unABL+22CSDXDltd4JjT8nr41qb9FmGKe8kiaDov7X4QSllkMj+p5sZ6BREPE2i9XZKonX4
54fMJ4vyiTk8hlGoqyIgq4+TvlgIOPCgXzCbzzQYjV9CgP3a03i6XrmFxrUU2oB4GBIF/gCH2Kok
vsfJ/atUaH46U2Q9HU5wDL7fy1swJJIu9CLNvmcUgKU/PMBRIhTl9QYMjzmbob0OHxqbnEhizH4e
1JTrN7huoQUfYs47axTXMrlL6bwdMhzvbMljOKaCHw0iZByUPHZmzRSXwFTnljtr2jjitZA/Hvo1
VYbfqV3rJxC6KuUVkzK4t8LlZ2SZoDmBAsAKdFKItXtYX9qITI7fHmoXyBpWRt+dMj0sSPaS3/Jy
OmIBQnkoF2cpZr/aVbZBLaBQHVhL3cdD5yT8gnioaPjbPMoeatp+sCje7wYPwtQnHeYbsBQt6Alo
y/BP6X1kL4VnVPz8r9UtxgtUkit8IWF3/sj1LreUMO8meNYf9iKqmjNt4kVpi/LVgZc1mY8N0b3t
ylDUF6exrx1OyajF3H+9tUfOWnq6MpKZAc1Yud6iOLNw5m8aDkSOqL1F2wuQK/EIF9lion9ixoB4
qrDP7KEIvxRKorG3NaYu9j31jQYsY37Zc38rqpQBMxbEbK952v8rLQq6vYOMJ88FY3qRXSsdjBi5
1zwTbys+im2YKLqRC4eFxYniatbfmnd6j0w42RhiThtDadcYwaQrtu6pWDqS2XyosLoZ4gq2gPSL
1r06AYwK2BZTN84to5hz1gp3wtBqze0Pm4kZk9sojdHOX85vdlXjE/hhNCNNRO0pIuQ6N06QFQTk
bN7fmXWi8SrgtDw0HUOFsciVGxErH/qZVrNHVTS7HxHhUDqEEIm5XSmqSUY17dg7NzzRiEL9I2so
tr3TXcmkA1uVLhvqs7JbNDDsO0qSkR+SyUExbku1L82Mlk54MQZ5n8Bv9gAZ15cmPXWyjnJDQNMp
MJSy0JwADt9EGJG7ckjFnsCt185UVthJsOAr3+P4nnXaqr9ra1/V6jm2qpDtEtMS+ae+zIR9y/Yt
qIz41NUDQgrzYvj3SEcfdFSdydSiR3dtiwBjpA39kUu2KTrVM4YMBAPNAF3pNPfwdhP8hus8uyh9
UovagrR7jM1xAHShx55gqwgmPgbExCPWVVbB1Yvv+r5n9oebGDC/z/AcSzUJCrbwpuFn2sfPifMW
0RjGMJUvMANUerDYnZvdExbxCI2rpqOxazg4yzG0CZDfP1Umbl5kH3Pkn4XWAmOweW4sicyMKUAA
2JA+Sjyp9Amr0ISVnw7bCnKEXsm0DfAoamWNQHBCvEvmspCJapK7+WtqZInLxScHagHgWsaTyzps
MLJ+JbmLVhgbEsM0sZpjAlcXPSX3EqpsN3soWTh7nc2oyRNgaifmIZPlar7Xmd+3GingzNr2Lk9B
NzexitFLwN26yGEklFa6YYTPwprjgkagsYrdeCiuU2q1L2XBJERDC5o+018j4e6YLcQB54Usmkcm
eYaGfwabHFOdp7QMhleTuR8NW4EqFd/7+sHjhyvL17NMXCvkmusO4069PxVJ1t3Lc0IXlxTrZWf2
2kpMxQ+9s9LIrFSheOUOcNZOpSZBf54odzBjck8NR2iTREPuwMntAeMCKi0j2Wl7U+tuKvHUdMBu
pzQVoS8ElpfcCU47VX1Xsnv3BkuY0+u1IB8DXfXsRr38lnzJtNmVgD5ozdKPD2VzmeMFO8Q5HKOR
KRxDje9BinU8XN6EUXlKKj4sRmdvGyd/mcNqlG0klrezqbB0y+d2OvYgndDMZNBIBqGOb1DRyUsA
YHXhpqHZbCht2L6bM6lM87U677V11g9F89Lqeb/3qKZRUyDo1vABcCS1rw1Vm35woGW4s45SGymo
bzSPveRKcqsR+ycORFlzFBrap1VYttRoXxIIL7Kn5xum0Omk6b9VoKfvqfbac1CSQ0TpyQJtKO8F
cJa7SOJPIcaOwu8UEQv+uPoTAqO7KdwFyvlc4fmCmYbgneijyQGfQOegLey4eRPKOJ2g/kfxiAV1
DH05uXtxPfg7fP/Z9Jxq1zyY1RsaSpmuw891wwp5c0J7oXNbXZfOx9ECl1bA8U9Fb3WiwnjaGq80
yRzAMPbZrjpYAe+vJdBQW6TArq05gPQ1HkRz14wSTmG5x0LSIoz+ojUrBs3ST/SaKD9kWJEm1aSl
sDmUTnbp+X78/BsnJsyjSPXBSUlowsRd588h4EoQg4d6R9YD0m0yO6CENkhTa7K4A8tIvD+zwlMs
944e6Fqqkls+4hVckGBkVqKYZ7bckhtTa6XNdtZlv5B3X7bP4cVyC2O/kCWP8OcCRQHc0wWRHHsh
ixSlFxSO665vJIrVvEvFPH+evrVT9tFwv+EdC/IfCJ81W5htHSmisjMA0Z8n2KBd4eUVSAhg5ODw
OOpfh6PDv0Vg7m1ZwB2wIa0BTxungK28cs8ipf1PfKOVZn+rfopp0AUp+shmwdaOnvqje/uNV+rA
JuU1MvMVRit4V3YVqt2KtMTrijoDhhASF6ZZKt/FAejZCgkqtFnd11StQhMO0IWdaS9Ke6z+WybP
556NRZ/Nnzukq8V9bA02jzcz7RSqBcE/m329YbR6iAmSJR9YRQLMtPyIHDW+bU0sm8NPHlxCrTLO
gzzQp9L/kmmmyirZCdT/+3VECR3NOYaY+rpdKlPfLioVZ+i2WjQ68QmhskpPtyZGp5/yb8U8gIIw
NNhJwvPL5nbBR6/5oD1XVhmnh8Npjyz3LGWRX3R7ond3FLHYT5o+bkGS8T4ZkNbn1SY3yYAO+unr
zNhmGXOEuAd/sp1eEHdAmjT8hI4pYTWbVmnUBkK6QpL6qwOvJgCIimXpN5rAXvCQtphVpV2xGC8J
yFg0J4BWaARK4BhFYayoh9vEUF5GK/gSJfWcrlQSsPy0E2R6x5/WZjtgmxE17YPPu8IqvnYBWQVD
k2FU5Sw04N4LkQSHoZ6HK0yGLG8lUsPGMaZISwlzni4H3RuRZNIdCFI/QTHLM4//ddiMLeoFOx7w
T3g7Ka/LSChP3+5roXjdSRUACvKO+vdF7XB1pqARpWVtI6IBH1RAclPYuiqeZ4B9WEbb8/jz/aJF
5KrKT2IHaVaw/jrzUUy3ceWPGLjFIUim4JmV/e95mj6ytP/XOf+l9VgjvTzturWDog8FmrUKugjS
VbD3nU4T0f5mVsYkTQO/Zbd4J9+ULla9zLXPiq3MpeAnnhnmKyF4YFo3f6vOCcN2J90EX0NhOusD
uAm0p4sVoupz/4MI2/Nlh3be9QCX9sh1iCSmx3Mt5b0NzTB4iel5WWjA9U05sbOPvPRulCvfNSMX
P5ZCsySOIFWQhXVdcbzT1shF8FZh5TN6LYNlukf57ikmA/RsmtajNTVEEAn0RrqCzuINR3kRd6YU
nOkIlErrWevD0YpdKqP2Wl2jr1P6BgYjCLGgYc5LaOMgoXb9qKNOlcfbiBAjx6v62fOm53tBiptC
B104tV/wG9KHlK25fE811cVizp14DQic8vceIaCVLyLB3iSjPUtGzJVPZBg2VRF+OoliC8nzm8Ll
r48owMl/0legsBqWC4+9SkBUMC0c+2i4PgsUklU6KDtKbRETMYWj0EIY6j8/XUexpsZsRzes9SFp
stecmKItOZ/63zcVrBXiYIILmsyaPktCn7t9RPZd2E3k+ueqBhSfkIdKUq/4CRZd0wcRsClp3YTj
ere4Hilfc1Zgj25dsSb+oLzxohW9LREJ9sqZT+dK18WiRJqCG47IUpy0eZUjLDj/3+RfYqfcSG85
cuVrg29/MafawMcUHEXBy1HVaSQGl5ywEZLEnaKdljqP2d7wQOKeOJYFc4yF0US8MvBekyNO3gIM
sFbMtfEFFaFroy81aWQjhW51mfHkZUhxNxC1CtmneBU6MzPXbBz7Q65rCDLxK7343bXGA+MZuJkE
YXyz7aJ2l2Swp+jRlWMOu0hSuzbkoQeVmIuPQFTgOhLasRW1kswqLmGexvq7pRXWN0JWeI6VrAqj
bB7YFN4ReEluNCjF2aL8JJhB1S4oH/EzYwIpw68q+0yJFiHFTfQh2IhN/YsTzTE5XgycXTAwyauT
YqGUz3KTloToduWTkFTtf1ZfXfuWe+2AnGeQJi/gTin96hNFVn1Z4JKuAhMF1NHWtHedaXuZ5DAN
g9e76RM4QvGeOASz2Wdpu6b1x6BFvUPuCWDTGVaOruL9P0Sk2iwnN0iDtYpnBm1W47XYROnnMWdZ
eLVRAtdNpC6SzD2McPFVLdNRj89ET7toPRC6PtpXEq4R0clU8RT+zZN3+bYpGxRKoITxYaPeXcuG
mxpHUbcqpK9ph0knYxxG2O7ZFRyHu6i8ieAFOgGw+DP2p7SnheeDL3XvBNZyU1pOh0cfYGDePfke
hdiDR9JnDS9laYPiOXVR6t0uMz5ubJNu2v5a03cwXLPEDlJvuac31U6Sg0A2kP0mWIoUwoYSsBNX
XYlble0UchShaYaw9Iix36JQ+KoZrdI1VULUvV9fv7zsy0x7H1v5+Su3xBk95DG/sOYF+EEsKAXd
oDsQjvkfPIPhODnHi7A92k+j+LGmDm7NHiqGYQ+dOU4G13mwvkEpyIh8m/vHl6H9FimFXwANXu+H
cs49rdnmj9xGn4Ta+/+cBXgd2fV8C8j+IYB+u2tla5lLo7B6o2Mb0QiBZarSkzq86+/YFTBpY2A4
/Dsbw2Aaz/qkYBbLoJcvsh6U6oJevOytpvbUzR0aNznZeZZkeQp5GRJ9df3n7dCfG4tgJ1OvR2FD
AM9P/byfccqsa52J4Po3pivf7WPyyQhHfKb+o6LckqEvBNClmrvMk4BjZv4JZ8TU6u347E95TR5k
0YyqqkRRXnOqlgZJ29RdSX9Woq6IdkD4dvjwrrc8N3W0ZraBEgYemSXuME5xNrXwGTbwNHoLlYg3
MvOJ5KWHEE7LQ3EAlcyFvilnxXKxwuqrmX7Ed/akeSr4neacCz+xdXhEERM3ATkk863abfusOwnF
glu8B6J8DYlwsFXMFIZQCOhBUrS3bGQCKxEIaGph/jLAVcgj6AtUJE+fvS7whDyCjHvq75nad8RO
GzxdQROrq05QBGm5pcWMw3SftPCTKnLJP3wE6OAvdwg9lKn9FPnczagJL7LwBfBJcVqvg4J2HIYg
cXQIHmfkUkLZYRbIvkvHKaIxonZskkE+2c8H9UDAOnLOU5fMK5ZL0CyRzztQ07vXuGkhIE8HBlXj
kUG2SPW8A7wCwh2YK6arzZvatiMjPMHTQyI6/rgZZ5jvg4N89bAsp4l3boJUCNAHuif1KbKicE+M
tDWviZLpi/4orTbGzjqWy40EEODmMVrI49xpeyFpNpDW6uyjWAB2TTtHzQ4tSIRSu5/HGcDdOa97
VegdlLAjcApsE9DfiSWEtAgN8DD//wrah29a8cBoj1+SMap269K8puDSNBiYR+xeg1Puap78DTZn
pHdX1d4g8HVHwfqSNs1+WGjBeaMspDgBfJ6olRkfG6R6jttNnF9LjtPQPJrGcqsc+sRtI+rwX1SA
g2OPrt81R9j4XkqMDMaAMKZPeRSLAsPZlaQDeragvSAYKCatYqy+4s9Uh8GKizP3bch5rWqLMkmk
c1zux187VK46D0rLl44R7jNPEcre/WqFdxX6k3lBrSWPVK7v4vj87jQudvx5xevxvd7Dum4MRz1K
sl6H1sZn6+/nVTDKew9GVdxJYZ+hiVMc69Giz8Px6cspCVzV/zrwWs/5msGrFnY45UKDOQExorZP
sXrRCqrZejQbVmcv2mjlYKiFv4tUcUvbwEDLE+PsL8rlcobyBsaVYhGnGFIb/zchzcnMXMiy6lNe
6v8XvMV0QsnxXra1TIjvZRlXHLQmFg5QmX7NgveOqqw+DDFJQkT13Gj0PjsS7UCov6cjxU2XX+y4
MtGDLRhLGLZbvmLok4t3QzsMxPh+KSlyRfIy4HsivRnseCwtTaOlc5W3OBfT1xOO7i4zG4h7mSAY
QH3CZ7GIdprA7E6CMhUibgEJFsu901HHWPCchxuei9vcesVmM4TZPiwS9A+i4Kd4Bt0upFCvnoif
gAt2vyefXW+XnNUhPokUw+L3HxTg0Hq7sb5NVT123LzRdgwCniPt45zW8Yiiy5CwQQQdsCIZ0XeS
WR7A7lt4KehlvqhFi96KOf3hQ4QCDnF/TmP1hF0dbcXQr+Pe9l7ySveCsnl7Vb0WoiKCToU3/q4T
FQIZiJIUnHsVzHDc+2rTuxSyDo5aRAPkUAq/r0uJrOo0+RiJ8KynlTJfQbu7fHhQATnrrMERsvNl
LenIvimVNE3ncWoCi04ZFqpE5yjg4HWKzMLtxWhHnCiz+6qasi5eVJVoaprA/uluKy/i7lcvO3Mx
LOkn2runaLSwXDppi8xGmoyGZGaWwYOHc+FvTOAC4dmyMlTYHLu/JQb95L3r3ZWRKaNZONUH9BNO
2Y5nlT/Pb5UD+kIYoz0xhhs4r8h64K8UmpupLdAUwv4rfLhGVhr68389vMqdXzk3HnkvfckJZ4QI
cRLSvVgI+vOqi0YyiEG5qLrp54X7uX8SJO5lg/26X/cCesAc5PNbDL071n5K4hugJE6FYgW5223T
HgWQHIhhu5Zz2By4kQFXS4Ej9+GAV//LBzEHueSh/jBwK4s6y/cE6pjy7gM45kp+CDYtklrI8Dp1
XDWOg5r112rOTB3kDJUfeO0lReLsYfOatigTNANViM1bscb4zAwiGvVz3bftDHLVmccphxvipACI
7JZRlDJYMHspW4pqkDCCJho41WnjDbXnHHBLiBmqQwq9bnKb0oA+ser1M4hQ4k2b2xEb9fuiQc7z
M84ifUfTsDawXrIuXdeNcjCWU4Q89J+11Vu/qW8IKX22jYOEOJxzje9hCT1998mbHwEG3t6xjB+a
r0OcyXF2qE93Ev9xiAHb+AcrfvrHWCO6lXo/H55kxVv9aX05Iwujn+IQmX6mEKxpz0uWskbDsJBs
FM3UJpHTrZBGeVbJ5omF0Uz/k5qN55p3dYVhptBIk2IM2HylUbv8AFu0Hsip7Y0Ub3DJu/3A/gVr
xt3dOc0w+jKTTDPUi34iv6o5d0mE5r7WhEv4PBsfuR9JgJ/xb2b6wrgAp63M9oe9Kq714mMzWQMT
fMEjbxiWDYY90gpeul/s8RsmRgkSqymJ8PQQYt/9fa2fFEYypqnO/ThbIGt+iyCDK2g+3rM5lVns
t2ioPZPgkG8N4mWlNqd81YUJhdEbE2X1dCXfyCH/NaZ0iMsZNIxcRlYaquwU4+cLCxdEbYdhKzyt
VJGYIW7hJMVEuFQQ/nxjgvjAWzWLBspugRRaAgSJVTA9MQlCdHh9zceN5uw8pr+5nUhCwpPYYQf2
73qE//ftAT+Q2L1rTtMIVVJNeSoHfMUl6XtgHX5E9k7pHEaAzATixfY+xDdUBYRXstEShaMLQ8Av
SeLn2lJsor+njW6tYDcnmfl0HiihTD2I7+p1ZUXtQYvYtJaE6PpkXuvX1RsUYPxB5Y4c/C7a2b0s
5r5wdvnXWKd0FiV1QWjCI2bdfUUiStRr5LzcUewMiRCgXb4/3kPSQfhtGGlpwnRnDXDcVEm2WdhH
cxK1lw3AlajzlO7NJMf7EXh0FLF3nuGBp2TW64bfRlNUTlsKOcxVseoJ2vGUORocJGBXkD9e2cec
0eU2+A8jMS8xX8G9K6/s6zKOfujEwZwov1TSRWVLA/6nx9/vc8ipYUmf8X3SHt84v7lCbcY8cAGY
tFN2AybeyLMnrAiScBIM4MrIvZgDDDa7EBZZ5yjuZABxWanDBahQAl9ZTQ3boYN9dnhnHtoL3Ueq
2sxjdc4fuzWMPCES/rkN3q4F0fVMURWezJSCmidI9S37lQLbxn89QQ3gqfEk0E0s5YxJEm97w1jY
qXbNAPDAE9t5ow4fTbpx02a6O9idzFmzJXXj23kw4Rjnr766Ga0IO8SIBwF2Ui1s7CzMl/yboC3m
n36KdM/UsITyj3tboxM7WBxGjHH+ycfkuZAJkHjmEd9/siFp3BA2OpS3j/sLW/e4EBXjKhTtQUwm
MdNYYV/rIjLEBlnWB/+Kca0acGu4+yZNb/P6kjVw6G/Ge3CEXjunwFmt7622vQ1XeC0nORmQcjsX
Btj/3anl/IQMmNFvTwDBeCRfVwLcMc0V+J6UH8wshXGNX2+KGELw0Y4thuVJLejyIk+lLgSFcVBA
epSJPd3egU7POcpR+BmblpSQ0PnT3sJafGsJ7T/o5nVHuzYKBN3fFEVQVw/vg2nIXpvoBRF0Bnkn
Kyi4/HH5pZUtFtEJg0eQpqUJZ0BlqPI1RBWFj4Izp1xKEGN20P20z2A7I9bqGawrUTN7KgPW3UUq
TBEyrt+rpIYXQPW6lDpETcOln1paMrNcu0QU2A/jM6/SvwxkRXWU/L5KMh+X4d3eggVDGOguyvQJ
n/ubLHmJbd5pkee+B6BmyvGe4t2S7FDwkM0SDAxouHyN/TXRv5iZ1JU0Lw3sbsQwBDL9fQsWtOxP
HRxTEAfEVaqL5VRQySqbekOkyzNdzOZktlwdolkHmY+etQnNwU8QJMhUh7IMgS/68DLGiRvUXInz
2lnkEcDBj6unjlHS8OrMWcGKwANUTUWKzgbkK9GcRn8IHpbmY0uutShhCNOieYNwAvs+1a/Spi3U
Lr6fsjSM9SMZR8cWtg62mIlHZoCG7zl85T4ZpPkBveXrLrX0tbmQ20AF8CDGwybesbsay8IYBF17
PoQlaZ+OmeYm2Q1EZe6kPfbgslfpFIzgx0409oFjg2e7T8kTzc4trRoSYfZZYmwlI7qQtRgJbJfi
j4uRHE6GfEfW+GZkvxn9f8qjKBQ7+OwLYkdEgqa1xEsN5FvZute5zJb/bQbrvt/jdGePygx2ECKd
IJoH81KF/c3y6/MEixvlXeSiARttQ6iX3sgdWlhbARwUblzTfTE6Zze2z1PNvEoqLHzneWQz38+S
g8pmqJrcB8hsKbWKtcyuFWd/8fIg0YxdbXugHVfZm1tSMI0H9gAt/WuJxBBkU/BKXscdRjRTMneN
dKOHm3geCz+RDMVGbdba2N4eJGZD5pPYVKVAoDnEnLz+XI5y0mSnsnQPhTG2DbJ/VmlFTkjPd7sD
VWuvea2fDFYj34N5CtPCO8qHGDqXtPZS+bn6RWCTxFzAbcKLBDXXhTWHMqwHwTW2h9cID/WeYLKy
v8q4xt6cFfSzL+rPEZ3qyCQQ6KtsAbKDwmG7h4YAv6f0TTM8z9lOHHmK7FLJpb2eZYT+koEi2JWA
UFNnI7oormniY5i+dY/07reaQ6ZQGV82+OAvJBw9A1LfPYeUrZHWDFEu5PjshjaBycT0wjq/QaPy
l5+RlcbnknpJNB3TcWmcSXxpdypwhrXrthz0OJOBSSbWe8WUl5MCe57Df9zm4sLgBKdSHleOwb5q
R2nx3NPMsKOGaHBDPhnviQ/0PAXmHkJ0CIr40/xI7ClD/CEnb0mlu9R3Ir6w444xVnKNjzhB/1y8
ghqh967tiIs/kaKLbBcG2VqWp6vWZnZXUyR30+0BUwJKmBIH1eORD3/RQ4kvl2RZDlkzYLaB3Au2
ghEHI+WaZMgJrK811zrHA2bT3lUlx1C5Pyr/rfJJRCB8ScPXODtgop2nXvoGiRl97Z7Sw5F5Uu1i
RcXlBlGfp9OlR0xTdlTjjK8JumKAywEhKIdAMaCPAs2LvzwPZLxKbt5iy7jNeUdLMKtsA2mmD2UU
66GuPmujJsRw+4+MOQ6GNv6ZQaAQrTdCJ2RTGJaiU6SPfz989iEXX/NIytEigTrolxFTM+D/CXti
UustMU9eDgGgoP4NB+vkfNYAEjo7KSrWVDTU/7pjs9mgXkGfA/i5Vf+u+ksUpbJdu4bUCXfrdstk
K1W/JaeszizOipSGZlEmGCG/QT9DjoImLmVhCEOrMzUm2Q9OmE65kHLowDxoiwoDbc4fiTpyWArR
kydyVGv/TRJv5MD0ZSZkD/m+PqVPV4kdNacCQfVFmtKmgiYIqyKm3bKKdVgKOH/1+gO2Wmb8DqGw
WfVsl3jcuE/F66kfGpD9LKecdd56xuzWzZOPBdyLaBbqL6vGpHaFgAs/AaPcuMBoQ3OoWJ4xE9Tz
Dutn7a4wvGscQ6rygxQwMfhuO3BPmkAbm5Ec7knIT6WWkVcPn1rYGIlcfxwmH94QROMKrmvGcr4X
9eeRPpadnreNu4Xfr+2dBZL648mH2EubIhfJGm6rlYeIhiGaWxS+B10O51Hcz9p37ZBstJ0AA6Ts
rgwMiaQidtbfnJl0TI7lxH7RGH2EW3Y6cStwprkV32Ex/EKsTGyNzs7mJFgeOP/KIU5G1XQOO4aJ
Clwe+xEjsyalKt1hltMYE6CTtF6UDKE4wIRB3HPEvnk6ijIg3a/P3JLYMYQTAmygaGJOQs8ZvnjN
xM1kuXy91lD3ycP8BMb+E97YqFkohue2FlFquPoyUc/vqfZyLnjjDuEDxKHJQ/l4yliOlsdXmGay
kveUvs5c/VvOqjsabp8p4bK8Uu1+y9CLOBBkdSWG9Om40ggq54ukSO07lw8Ua4hKmcUf1/wrgNNl
SsDtdwP4e4dDhV6hC61+qTC1Ss3P/PCOQvsTsRY7n4IjMLbwbO2eI3fr9BQ0f7HmnJ98jkVdXMsz
gp9EiDOa11IukxZLykf3qExO8DlYVFe7jW098w7wB62yICgK+RpFdkJrAhIJM77l/Ic1uvraMBJf
1GAFYASHdlXLVqqQefKEdQJAdGAHNE1U8q+C7CuRgv7Ps4i8mF3LT5o4hKfA4OSjheyNyFkcCJdy
163hI9t4amko8idqAM3VowmMXjAvsNozGR2eRsLypSrM1ilaoH2CXOpVnPYelMY1I+9FTGSWi/nP
QmClDHGpbxmLACUSwd5t3gVDD7hRKEyjN72FVF1ViX9mTZHuHg6vXTA2Cs6jHHIIMG+kWv1JjbZo
YJlzt+UV2IMwN86UTKRIH13xJQEwKqVKT0drGlDxUdqsnjmZDv+qsEBh5qcrwLV5PvQaATV8f6GS
Mq3BDCDPWRQ1dASufliNX3Pm+QOfqshKpd9+bh2aoCJ4hYAwJ/EbDouPTDyDQsbkKUstjJUFWr9g
MGXMUBqAquNsZvC3abozSfjaG2nbq0KXivBzy9d+a092AlEEd4s63uJtpoWffTVoRVhsFmXLDx12
mPICzNw6nA0L3MpS4s9E/QiW7KYf7x6EJ0deYTQmkrA3GMtP4x2qDZTmfXhjz6+hyGKAKG/vIAas
ZOu4v23hOfF3otQWUqjxcCwM8HLwUb73aQGXf5rdPwydpqPVXRmA3Jp9wkmH0kXtV9A+LN0ufuJw
arPByF7XUnuPMQvxAOn7x18O63ZZ6YWuUhW3SolzeMww/vrdqFhmpgS7us7ViYP1NNrFUx4tRw6y
mUOcWgbR2RiQWf2gFE3qHn44EzD5tf6D7JiQdVni5GgheYpCFcetFyGZQqJhjigeIXbY1HS61w6/
q8z0H3pZGGFiNbU3NDo6XHnxYmiRyx+0+L0D2ttxMl3Wa8RMu52op1CtgI7FTo9G88ZAn7JFiDmJ
F0iSE5gf7pKfzWgsKhJt8X3r9+3wMZwSg2sPZ3mhPTE2sRRaTBFp5X0NPOarMMc9Mdu/+Z4v6lw/
iWO+S/YH5Vi8jILxBg/hl453TP++S+1GruVNHElNP2K/GS7ujlMq8t93LiB54xoSmVPuC6JfvBOM
vOwt3QOOmdPAmKhpLosdbJd1ZS7tGO24kQIytcv0nVX1YpeKHUw2f3cRpSL1jd7u5Td798Dggscn
vrLKfiW+bz6yu7MXRQVKarL+xooaYm9kVhQC5Nm6LiNJCKvlTyC62Yi1YAU9pgm9+N1Hi/YqxjnZ
EDoyubFoiVgEOywGYiYTMc+MdxzZU1E7FrBqp6s9HAndD9OPKtkmWWsgKsdy475sVQKmgRcaSMIF
/NDSADjs2N0A8rn71RWoK2ZOIrXNukup4rsy++zPXGCCKW9I9mCQq00F5KAAORdySqSf94rxBP+h
cNOWs5qVTPXKzjGqBGBULPIcrQxy7/fGr8SrGkremRU8HwKa59/5Q6be6+hIy2WDN6eDs/0Ag9y4
a3ydDdXy98oHblUksP5QDMw7NzfzC0gqSuI21xJXjetCBCEI8DH6q+zcl3y43y8b5FayfLeRSwy7
apVf+oXs6ZbwVj5g/qeAJ089Ku4dVJsN0QIhUnbyeI3BLcR2amAO8AIlPbeN37G0Na0gkEgSmCvk
YavWWI0QOglj3NymQgZIdiPUc0FinATAqPSYqUsH0KmsLUzdpqYgbRZn1z1yIJqVkaiwnKUZCyeF
5WMycgGGQ4XBUVp621QegxOkRACQTsB19fP7M3JLW0IWfVEoFgqroHx8WCEVQ5EsxmajF+Wmn9t5
/OCC2m5VoKPUiNumBtGOnA6j/pS50S+9mptiFG0VWp7eaf4wCQVY0K+3SWKFcAXfR7PmXxS6+bLh
pfpkzMWc4OQU1fG3A9rPdu8obAhZ4AnyZYoq+XD/SL7zz1Tf/1E/4hSr/3QEoIxx5//YGB6o86W5
zXYLHc/hnbNUZzItRa01P868DiGM2ywM/GgAYfgL/eIOzBR6YWz9JMRuJ8njx4wbkTjn87+1cPKw
/3MvrHKz4DGN/Et4bMZBVoaCT3BUXzW6vcDk4O7n132zwgN5xYoFnuoWUPcCFTRAoYFbZkqujDjQ
xFFjTRFNiFDj36+hckDiOAhOoRwmkyJMK3Gl+oYFCgujpMs9w3xRHnVgQKzxqrJGMwfpzMrOQjqD
l58q0xxoItxfuOSqbrn85eNmgyOGr1rJylO3heowPZo7p08HBzB1RrzBG3xzCESpONKtETKR+gjs
4TSyHo9i55QIQfieJqCKa8P6IjnKb4gfCCudqJR5jkRZRZadfynofeHSrXg+Wmcv5bkXjSwDuECz
YyDAGR81LN8LZ9kLYxt5t169tx5cpMCLvfGK/62dlhDDdmhG7Fr6V5wrfIV50kMy47RfxwbM83Ms
AujdAQzzEybVaJq/EVIX4HR4JcQQ5D7bLs50IYa4r3Aiaf3/jO5qiHMRwzE0xcWOwK946og8NGjs
KBk/t7r2nGAsrdKSIYHbnOtFYYPYGYoMGnkbUDu0dcm+IP1+VgQHPx+YS0fCF8bQxUmn9epgu+Tt
1dn+7eVx86gkdxpBv+esYm8WA/7VOw/IrHyavEzZgpYaAt/RtWO9ygm5AHCXIsBzfjXA9vFaTdUE
fmUaABwLGXEBMjNjx3QfcwKjt8LqFkxc8kcJk8kjJgDEYe6MeaI9QSOD671d8S4eQMezYvsw4X/b
iQPgjFQenjG4ln6/HWrpCq0HniBcheLqSX3Ny2t/AI0FIC94jJl/6KqY1gBZ6f30h0QlnPh89kxS
DLWaVDoXNvtNSEsafsp86VG7+o0fWUm2UXLUClFhGYJgRwq95nDnPk/f456ZOG/VsAGvcQ0Dz5e8
vgriVN1sgXUFYR/hP1WI5u+OuP+R/PIhEzQ6V7I+9ip6TgdIDoG/EapAkVXDXr/+sQGujOPia6rc
Q6BUBuXn/SgOIaFa++lfhVDE3Wlp+GGAK2Hz+92pxHIOUgIb95rMS7C5+vaYxmAOAKPLuJh0Hvsn
Sk8uYvGHXgMlYT3l1ZS0PcNoQsACgZj5unOHUUC7WyBp263AO+EoLorMXerNnVtsfxiy7hPRr0uV
2UfglzqgLH45fsWzgJTdXkeIg2DWnRe+mvwtO9PMO04r2WFgXfIR/seQtVzV4RsxwitTPRGG7qiz
od64FSS+B+XcJPkSKffPb8m9XskrZN4zppCkmT/08t/IL9cifQR/DJ6khq+d4fEvsTr7t8Rx8Au7
HfDYpiRJ49jWEEag75tjsu+/3w1ovsReGrkxmcWT0Oxy5seFA8Eu1Emy9IjwqPjIPnwsFofFzEY7
kW0nGCtij16mxISnXfI4AYDae7nYX5ZdLrQ0rvH8F0U6LMp4wbzweO6iSM8Wl8rMVRWL1GXV3HPs
npG1gmtsjUZL9OD964ugW8yFoNtR5TQmSFdLA9GvwqXMECk63PPYOWWnBbbCLM7TqWk8M2AXgCQx
YoQoFKmaIn572uj/vnu6AaFEtAXubOSjP2u9Vo298OR/5hWPsR0zBYC7UcKFu+Y+olJhMYNYt26k
H5LsucqzewlOPMSK4YIS/jV7dsTIqFXvwzZqTRJIhrttaunqwBF8i1mb5GyQLMFt6bQ2PTaXlIKj
lPClwnW1MikDuO9efxLSwtTUo7LLJ8bA8hi+oTn+X+30Hj4P2RCc5YPgLP2LG4SjQZ9DGZeavEWL
tw5VNzeO04I/1vxO5ieA4FPvySDqNOpI7+y3EsLMCtWGhNwtGu84GjY5GaWoPMcRCq0rBfa4uQZB
Ik0UcKesfw+pncpZWXTmKmDC6T2LMOab75PCteEmjgC10/dQ98U71uDflWwacm/A30jKsfMMH31M
jhw5us4AkNHmCxJfDcQbCYzIDyJE+blUu+Yq4+MTGLDn5jZXdlA6i0+jXQROMdu+pfjEf8Aljndo
wB+0MiiEdeiqK9W3ubrYMYGcMEHu9SC3WDed+zimJql8ephC7DNpaqWWkrzNpVujC9Jdnhu0fo2r
qFNx4KyG7CBcWAOHtsnCMlBlGsXXYfnKIwlTI8n7LMESZWsziFElURUcxfeQiEeZRqoGbrjXYoqN
/sBu2iHnxkFJyE5lDs48aqOrZHA8pgnO5GlC3jGvZ0Q67o2Pzq16yedEjOywipSW0oMLF1tmkxCD
qVXpL4EPyCMTM8+sh6uvTWCgb5gzSZQ7bDIm9RuOFJ0pcL7UAd+Vq+DOdhnJ3nQVO3dtfbxbpwna
O4uUN2Dcfh3F1kDSdlFEWJY5D578Dwv1yIxuM8KoiHIAMUr25ivD3i64IPX9tupm+yuqwuhJD7nB
HVko8fTp7NAChGsoi+AvHejQUWvpI6QlphigOuuXy0JOtSQ1b9WNsQ5SQVln1rbhJs5ytDfPryES
nICjl9HL0HOMZD/RRuQw4sTm+EYL//RUHlTOb6tnkHjmC1bCuOkCFUfYhzcSzxs/SSTTJuM8n0HT
ZLQg99tjYipw/rbtB4ybLgtON1r6jl1s56Tuwm29C3MQKAbtKoADjrlrYnPkpoS4q2HiOvPgA0wL
VKE7IQcs39duQwGzlBND+MDpElv3v1WTsfiLI9JwUtTUReMfUV8Nt/2dM8NbzoiTJjK0tQ2ogn6X
2nU1ySLtiaVHn3s+gGMZ5sXPTRHnS7PJh8utCEq/QYZpHvDSlvK8UpGvAVtbD4SqINAYoVHKi5Zj
GmgSZ2NJFo8XylryFsCdS2U0hxLO29MfMfJATlMxJFHSkxlEYfQgjJD/IOF4u+xz0f4Vgs2lF/H2
8cNeBTr9imuCMGM5xXFccH9uCnNM7VLs+3Cip97t5tlQ1piU1Mjm+BzRPm/i/0w7Y+fcyT10dvQN
XQe+Qf7rxOVE4TEnFi25vSVsmFe9izPVkzLVI8Ar4TGUqaT3A/uiml9bywH6EbuH4YG5RJ8rW7vH
lOBjs/mdIv8JgSQXTvN00wet2is+bbO6ZUP7WcJu2e3PNfNHu2pHT2vURnIWArMXRZyqmYDyBFZd
2X338r57sVFOab4pISeL7VVUeRkU5gE33wurAo2jxyd/t6JsIG4jHfDb/YzuBHIVwL2MHvfT7c+Z
UKvtXRKPldzDZremwtglDhWVMYBRCwYKvvfW8Q90bHztbwqcSDr9LAECi9W/kWQ6WQrSYpaR1AkW
F5+D7jiQKSeAHoXoWLgMVw/082MZViyLDtz2/FcQWhZ3ilgpYgrpWiSa+02KL/0doGtELFFlzRif
pOhM26r8Iy1wndohkUFdQFD3V2AYHza5YVCvDoXNOLTU17mIAAm94v68h9K04ikXxonUoQmzr8YY
/MmmlY/nlg5foh6KhDNRjzrW/c7g8s6G01R5DXtOHAPsWQWHUPHo0F4PBm5UjKvl2WcaR5fPHtFl
NMVEd6dbxgb3eKTG+e2zhjo/1z6bzYo2sKr4NyVfbnfpyscp71HHcNhuJIpdVwR1e+BoNuyyqvk8
6a6mFBoLH0e22leq/goIqHVbHJKPHI4J2g9h2m2XsAUJdhrLG51hukIJ/p5Ejyg+nKdinCpRIDR2
oLN0NzZAeJFeOYt44EVHEQVpR8IBGCYdYOXvUtqkIxZZzd5GC4EjpoQwjij3eNnIpegSimeFij4E
GQzJh0ShIZ4n0IXTAyzZ//BrCwaLdWRalOdHXer/ZUfb1wUsYOlI8dhip3Tr7szGQ5U2+mgwcCMF
8aDAQGHeA5KOg6ABI/6wpWEcK3fNoPOQHPb52/t8vHuJMSNlL3Wm30YB3WXiXRYfDXi71kdzJyNH
lOu0o3p4PgdDQfiwZYgYFDtU+fMKGDqGV/blsDXrjVd69v9LXeBiAYIdXaE0loye/8b1OzdmCYYN
9ZgtrqUVQ7ZdRJqEmxJUx9x2gxQZhNcwMwWKiobR+HhUogcIHnCevCQAuhW04eSuIG8DrmfYljlU
cEmk27qwrNT+TVb/14ED37ns9BxLqaMb4nPLo+mWgkIF9PFmeu2nNiCVRvMMQJgtIPX9YmiesUb+
45WAddsaGCF8/AHQkTQyV4oQnDnEk79GsKqIHhpy8qc4HatCrXjEI1OjIW5k3neykZxUOKDQft29
Slc8D5se8MwpFazajIwhn+eHe0cN/7Jw/KcF8JF4vMwwI87jkCCjNC7B8NCUTDCYlyqMxUlmJGvZ
iGSkYOKqib9okZuvfbal4Im6DRo95qlT3NrMPZhIHRXCr+Xr9la4zXIW+/IcpzSxxekitLlLepmR
8IOHNrNPSeW/KpcwbwBG/qxbtAizIgDfT/13ay5ik8r9okEyorPkhZla4JPY091fWZNawTaGhX4D
gTxblAjlpIZqmIIYS3WU0GGOanS/3hCdAYmahT6E3k7Ay2GY4nlHicp0q3LBQLqCHTEYf/6wJVvO
tQSLu9Y/Y+1EJmPOHNhM4rdEFCSN1+kksQgU8PsRDCLjGWFF93hj/j4k7Yp1UFH9luyLEIABm2J7
0rsHZ1AOnUkYs+eOEW/PqQzg3qN/Nc3leCgsCFauVimjJW8qUJ/SQO/AkEen+dEg0Yc0+TIPb0Ga
fg31h8R0EJDKooqXYQsS+dAcSLDcvfSQtAhRklB8eFj+9+9glWzDvBMMPF2xV7D3j4wI7Ia5WOkD
9FOE0moC+8G8kFODZOvXrVMzuZQ9Rfn7+QfCQVVaOe3uRNhZkmw7N0c1A/Ra+ayDH+f1j8AAUbal
iFAqEXnIdNQmspGjogLLApK+JfDV1nvjv0BNb8k8GX6ykBbPPYzMZo/aaWgugLnFIZMjcOmAWDn/
B4v+KZtSM4uEsE+nFxfnXzAtDUNUuBdRdP5xyg/xKZYwINH3DU1Q2ZYkGNC5W3pWPqdkei+GGhAE
wyogkE8GmJ977t8dm8hedUAHxpAVsWfH0FMYxAr9D10xJ6K5g7IoqXKQlJozOmmm/hHwmRw0g4ds
U+BZf2B6l0hjvMCjpGa1QB5IF1bbkGP4FhZcDOR7s9+QdpPxbMb9hZMi+hMrLIdM2VrWfcE5+oW1
fUxxwlLD93UmZpYoz2qB62KJOYpa/njgiMz6wuqB2YyR7ob/7QSrKIBPic2C0SvNp3/2t4y6Se8h
as28+gkXNEZacLj8xgIjUTqZ1K1sN1mAvMJJbIHZIzx9qkmUxkMkB8ZRlhcpviqwBWatWiD8tOSj
ANQ6NdKspLmxS5j0s0dmX6lxNuELkSR0VSCkWKMJ9EU2RObNYUsdCMlBybNSOWyz47UlQo35qS8S
VdHGsV6b941ZPfaiYZgZ+G6cR04uHqmn2uGqQAG8NF/n6EYfponlBotY9IppeVINxEevJ3ohfeLN
WyuHl7If/EVIKvpdZKOE8rueW+Sw+bnR94kMUZ5SMXndbbjXDWJNVOC2nSc4rUqIfD+Hp2W6fKKM
sx8n4toqlgITH26ZSRZpWHaKv88VX4evhXcKvx1e/BhQKcQKbW78bqh0GrXES15GVuKnKMGnZf7f
Um0ZxPPVcdNa2Efc4dFJT6soKlW5A+IwUk34mLp9Xxk57iltbPHoCHdFfDwUCJFJSmR19XsOkeGI
FF0aibPlCQx+jsdo0vO0OESz/6+9kB6W/05qQKuxJgmAmSD5FDTWodep2azc07JrcUalmLvLyu6l
XF7zyqBxJvxBLmHd8T2wQEYwz54UcEmNGsGf89ADYAZL43pXTHYrdRm3O1jZHL/GBa6Kouk6BuI3
+bU4tDE9EJV0Xcvgg+1p6brW2JQCQ9JimuAb45JwIjoGaPIq8omowqw6MqX7YLb3OhrIaqLfK90U
/BI5ggAZN+GfsT8FfouprR6d6/ZHjobITYlvebaNqp7FCNnKBJQlfVcto/PvkEYCymH1ZUPwDm3e
UVS/jxcc9MRzA8DBjdjc5zsLsY/UATcz/VuAM/Y9SPhacAwHSw29VlXS/mJKQlMFAwr1T3bO6UxH
USqj4UQYAQAegkBHu3IKMOe7F1nM+z51j4eTMs7HwOSJr9jj/FIHnEom10TG5hIET5EEwg+ObDGB
smxZQKGrfMcELeB6LwjGhjmxcgREa2+ovgHys6yrdxKpI0ylDYQJucKkVnpyiEOeBwxS2rQ+rl9q
s+qTKgMt3WmB+e/dLn+f1Xc3UffaWn/1zmM7prN8itHkLsq15TUJFWwY+55TpqPUfuU6bi4P/s/a
8alHhIE9aUd7VFLKVsjncey19aUdNFoubpeKeLbvg9zVXQ2XXBH4b1Q5YA+TKVpgz0AGiHDrRpLb
gXAgpVPS9/BLmusid/qE+z4CLt7/BiWrA8feqqA3BGlium6+ZIg/VDNj3HUuCmRttF0I6pR2pKT8
PF5m03qJQTVb4qrn5HMFzmdHuHS7P5AgN2kIa5yIC278gtyP9ubJgYjuLlEkbAKMJzekCdU7PQpD
7aST+nCQHR67sHu2u0RiUB8OdGOlMwDKcicC425zsZ8yjrfHVBh5rSLkgeVl4JfvulJyb8rLQoTH
/JfeY3+mEDkpynd/KnLt4dg6z1p3G3W5y36+VjOnjqLa41Si9OgBUeO2ZbRMfCb0PDcWVK2sRkRv
BFduAvTVBtXptM/3KTpDwd6AoTxCDNWbKuZ3N3ZWyfl5ARsD1fOEBhyZoG5bhvD4kH0tFYtWm75d
LshHsxN673IYTqoTZ6TwjoGgNoKIS8pBZjk6J1VvCzhv4TbZ7bXOI3YsCPDrMZ8feuiwn7CxxwcZ
+UisTKtEIlfi6ZK8RZJJW9T3Ept3Vcu1IC7XG6gyQLh1uM+7zwBztVw6kKs61BW5l2N5zKqtsaKq
byJiFVE7O/Yo3ENzcnq8Bc/ehyGZkcb5aJ7+whXI5xHF/22SxQhWSbEQw182kAn5EGH6btkOAqUg
Lh3En1MDdcDKfInbUx9srUsSSFQCrfds4VUs5psVqBITEgHdOwxVinmGTabmTGKeFLbRgVN+EAt9
c1j/wL4HOdoKPKHWYkqNSgeQWilaAZ+/L8SiAFJqFdZtPttIfnVYZXiQXqDMqiqPfMm8CWgtbOqS
ojF823T4MJTk8Lo9hrkM0uX19nkI2LDjSH6bo7idD3Ub2bo2JyeTXd9aG7rGc/CK5mO55fPmTfyf
rLM9E18vMi1A+jm6jo6W7qy5/PDooX4c1IzsL2/s70hqGXy44yRjhSgHgVqJtZDnAfQTLnCPw/dz
fciC4iVm5252O8Txb54NOXbhxDw7NB2PSpfHUvwW6GD1sDCSzjQYCTmzDtSgq/KTa728/ookKZIs
mFsFbLgGew/ontomgDtOj1aupqafY8Tg+dhEfkNjpScSnlxLiuL8fu6ar74JcL9XkJCq+A0nvSwG
nDxgVA5GCCrf3MaYOd08z5UInoNdsTHFlVBOPp0PgOQN1FPa8nRGeQ7er8tl8YJTSk2fPeSYiz+P
d/RxLB5/4bXbf81pmgyRQaSkpKX8sRfIfb3l0B/8Ys/SHTtdIdhcyrQF0o1oE39eUbCzqSV3zHfh
3Ffo04AJKYWNkPjsNjeMLDJLoxeMPIAxbIGcM1/IcPaqPiWag56dIKaeBxdu+MmNNfpBB2WMyQEh
oBnikMdI4B2/dEz3xOxDgpraIcMA8CQ8UH/4gWqxIlcDg3U89NLDPPhNiP8tlK2/a9+lmW+L257e
6BOK5EigWcDWyw4+uSere3hd6Ud2zupwtj0OUlJHeL5uZWmMy5dHsFnrww9qJvqJeOonCo1LaKFe
cqEKlSL5Sb3sccj3uNVamWlEEJ5U2ofH4EqnG3ROawcuazkbRw4nk3LNWeQWERkmamg0B0Mz98Tn
rZwezGgac7/HiR+fKhy/wAQsal2Ae91pq6c4i0fsfmohkYDPthf9isnQ0XNKu0XU4wC8ug9pzAHU
48BVzNYGnstI4c5ql4i92UyBub0SPMWdMu7byKTK++HgaTX4DSRSji0eNqNEDi+4ta/NlHYzSha+
mUQQL2mP9plGjfmhkOtaEKajSIgdSVdVAYBZa+OsULbOOkjJzh1a/h+s3RQs+Yv08qRtHYqOcYwd
3qQJKoI8E5z7dr3GisIa3J9oqLgSKPGVf8dbYrDPupa1zbFkc/nTiEO5J6au+1ma8NrZAkwh/rR8
J9kcHO8Y3tYmBQT6hJlxzqGrzhXcMi2JYK5zb338/91yYo7+/xQeOfeS0g4iI9jnXoIi3qzbiVqJ
LlfgDLJQJlGhSP79/v3H6+m2VL6mjn8hRo8t5LtcsdIufBfbjRsIvzxkpO1l56chjQmK11SY+K85
n8QqkupwrdDCUUgqY6Va4HA1wUAW7yHanYaW2hSYWWBZYFdl2A46CT6g7yk7IVan8u2STBF1i6EM
drHb7RFCByhXbhjVoJne75VkEwakL0KgeAsMZGuA5YnL9Jpfr/1X2BBlxFoc5JpEXiWd2yViQKWS
wnfPfA65UdwFFxLuhUF1CMFpwa7eo3MEpIS03tnxYs7trVPpPhIbaliYdvKpvIUKnucGU327RvF4
oTxhdfqZjEKX/xItu9eMy3N2laKT6vXxXn3zTHsf5sihRonAwAtzXofe+MG9wmjFPRT9dglLD8nE
TqI/u2QVH+lc2vbEVq7+oN0AYjOR7mpu1aBD6JjcZ6hHb+zLDdo6EDQQuXww3LU1DrSV9MIRY8k8
GZ1r2GE8o3QG5qUqeAzBbySVtFxmkfWn+jZeh461Ol0entud1akKIVJwCQaL5WweDwcl3tklH6m6
EPSv7N3AfrMvYSrOIhBETrycIkneVFcsDLXmP8BghW+23LG/oOZCLA61KH9APlcN7QP4zcVGViNJ
iXJSv4c/htzoaN/9jx2L6VSB1Wjn7813z5kC4DOawG81eXpoIgCPuZ7+aIqA3Yj8tZ92bCenZact
VZPxbc9gfcPY5lFFSLSfvmgFibvikS/ogKL0lFjGxc6A1u2s2Oo2P+kgGDW+ceSP+jkz6loa7WtM
ts3gnLtjyAIryF4gugjsaCMRlmNAbqoysioVSIxhBuv9szZu1onMy5O4RDYr0PbFNVv+MVO9org0
oxaT/iMFlk/aXrULXkR+yA6xjJRHL8gaH88G/qceynu1U5SYEYfsHBVqTQ41rWyqzWTsVcJt9gOh
xyMaDFCJiZ8jzfs8OyOBLjSiwOIki6fzPnzHDRsKxoaz7K1FFbKtbztUiZQDKnGIKbYX1FllWGoy
h1m7d0GYOMwakatT4l/NV2imKMm5i5tEJ7PJl2tFlhDPA9O31psrY24ijBYjNbVdVN95mjVFzn1l
vaZCNuk7pzkQ5V4fZxFt/vbFaV3zaGrCBhzSKBM16HZJkTdEukqHGTtvfofX4+/iZCv3Jbxm0+lL
2V8CNpaFbl8dsTdiS1fFqM8vVBjpiJTKhZUvydplbQzkszADKE1iy5a1RgpyeS2N/C93kKdXmiyN
/61RQjQZGu4ZEG0AAp+bmTcAV81wzJz+cRAJ4VsnKihb5OPAOkpXDmK5frYUxzHbP+VboUF77FPu
pMJsYFM8Jh06Iv9FdKOplVumbTAdy+7xAMCu0WiiVFFyFgbB3njOqjPAb/VDnO/AkvfVcMBdh89T
EK6cTlv5zQFcK88LyDEkM+yM4OhbnbcqCEtlUr4XFKLU2aRLfHKpAdjZJ3PNFDJTpUILkK6WJ6XK
72QfHDeXR4hIKaweZmakD21zPuD1CVqzWy8TYywTLILDxgwm6NhOucypjjCuWtWZKyXxE36iwBhT
JKc/OqomrQfvYKbq/COLKt4S5AgPpYxlD8X69bfKXEF+boB7lUdc2DSPtQylhTaMnbYnkInKoBMC
FKajztxxBOV+FexIQNrKoWlnisiQmvE0jCq9/edIjRQ7KdpvzBVOV1GnBxMq06D6g33R28fXFPkD
lbly81hFyfh6+9bN9SdN/qFVufDYLL0oRTLoFXUhC6F1n4Hyy6gxywKFmafweq7x2J6LPfguQkMO
eMZNJAxuABeTLOmp/8Y4CgZqllMKDxAVLCeAcFKY/RBU7h2SR95SrcQ8F6wtmM5i8AsXjMpLXGrA
Bwgm/8u1sJQD0ufQijL5batIxRjg4C+GK86L52vwJc8bqnBYuxdPzRkA5pm/h0wbxMaYmRXyAR9v
SnmJqmjon9Gs2LtaAvMMZ1/vrJXtPdBBks8E5QET2spNUVcZkOH6XIsGO+Hs+IM9FM+7ckYLO0RS
7povW4EAs6fB7Cb8simRsfYGWdhqtHjzDUW/U+QlCHloX5VFyeUeGcoCeTrfjlof6Uc+Pug8/k1i
N/GcOzxCA8LY9XW94GqfooD/kUoLIq78uUOTMv30r1ZpHcHT5DQU2A1xa0xahgFluDiqF+5sl3j1
iiMFBigu1olHdnZvYsVgQb7pZOKgX6BCNfXS4yHHLfM94Cs6MyrXI+uxmA+q62fL1iW1/Dmm7vdt
51I1A5xJCfw0zBgGMykUF+oetxunQClXT+JZl4c1giM5gjysw8/UM4VHxlh8KBdP3w6LvHEWLjLz
2BoUQr7eun2rT/8qC4qoP4+2B2aHXf2UiFxsBq7zqMxUcEwtMHGiLiI0iOZTtNwExwaDSBLmTX5e
cJ4qqyyl7ZfyVUap0xsBUstN2D5cA6pzPrQhtIvN1S++n7QY82IaexqrGEf+MxrlynyiLdImt5hv
I/6gPpEzaws4M/ec4HlfKoAflMjEalp/Gr9OTjXKN0z12+g688HT6+zgKcVWeHSevHttp2QDrLAX
BbKtec8T6l8sdNBpKofsp32FiYlR1NepEfKRgOxRvkZesYYxU3H7JRmSQV3GIo+guqiS27fx/R3y
Qhdmwux1URwy2x3bxAaPXRLtdUok76GUrnrlidxNeMAzY5pehzG/PzEOA9NEk0YjwcZWRvxq3IIi
DEo6ZLFXWI/Zg6NVfZRoBFMfHTWcOCi988iEu1ufU8flyu/iW6Br3JdD46GUSrbkLiWew0UKjmNa
wwBjUsLpmQyix8/hebzSDPTn3FUrdcRvp5Sm+HgITHgXvEv37OZjPgbx+YdFd3NtExDeL9XAJ8zs
eBS2hDnUh0Prj5ZbMIvFDBJm3TQUmtsKbUXa7eIFgDhf6MZb9yjWdueK1rWHfqCPPDdKUdj6D2P9
JzVUatrwfyAUosIcu8g6IYX5IELBYM67QlhYr8POPTzVrXJ99cqpdILIf1eXZcdx5HBDg7tl/GDS
CgJsGkewJKetvFaklQBKxK3T00aricN6XNYakJ2ElG//hF2XSRKts60Bck15h7TJm91MzJz2OuBv
A2LuZztkyHfJIX5/r+dk36fwzdihmNElDYkDQJv+d+LrUm4drqwgq1R1abTt7xlKb1Kdqt/quA6I
pWJKh1jgvlbG3ZPgwoApfLuEGsol8gxbmWEVyRekjSD6KWlhNA49V2WoHY7KH9yPjjzBIn2mYVLX
5qAebmdQxrzH1JA/ZBBQLEps5TjuQ5dPZcelP6ulOgnKwjOKq2aXjRLwx9hhIiZBKzvpVgUReT4q
daFvLSnMOuRwsXxoar8jbWN2oTRbab9ELNKBPP/bWhv8HBFkLpg5STT+cxIqVq5hxXV9Bu/vGpcD
ey1InSdu+taOwkkqFymIy030kTtuPZVeQWx12f/jlnAgMA0ujKNclNlhsBXLWxs2XOUVklfxhNgr
80eyu46ZEpYVBbh+v+GtDrj9HWKKqxwRnNTR+p5LzQWq7Jm8xwG1iN+3IDn9Y3zS1jfUyLZD0Lkc
VOBYli4Io7HODBBlX2ZZRRXRG5ACZ159BrNXPuP9VaT82nAgmIFKEOkYeaHaMAo0xtkESoZCGlNH
M5Ct98gLYNfa6rpXEZB3C4B88U3rrAf2aBjMaDzfb2pjMHEq1S/p8aNAt041nqxydMwidLPqr/GL
7oGdGYLC2IQ0KfgLYxpYCYFnV0y5iV/aiT6rPRNRp1MzD9hXvolMOECj/foklmp4eN5Q919aR+bQ
BXh/c6wWok2eWTpyzHe6XTF5BBR4uHFNJ6xS3hP2mC/L2WWG1NjTMJDaGW2MFcKBMKU4jn8hXm6X
bybKggS2gTI3kbQ3fAZXCuQ49qrU7E6/g0dJWa8T7P669X1CPLE1jsYV1iW6/KWbGkdziyanDNjg
gQrNqSq7aXj67214ZyMHEMC4VUfQJd3jCFQ3QMIEa6E2g+EDlk1nCEMkRJrBfMHHlfkN00XQayI8
icMdmJku1ZyYaOB/2GU2/8OP/8yQiTWxzCmpazw1cErdwQ8APSU/DwEZE2zjd/EvOJH8ubmff9Wy
UxR+8wMM4ye1enj0+ovNVTN2ld1civNnFCpZorDscfupxLdG5mSHVmY83XaoJ1Xu84h7+xTsCuaB
Qh7TXbapIKX1z9D4Zz9wWt522Y/prOGT9WLgjqihjIicpLmp+JWuzhH6/NyCVkW2px1P8SaGrzYV
1KeAwh+T/LzcEfGIZL3JSyaIv8XAONIZTbmKwifPp2eGemFeEwca5su8KBegIFT9wTt8kUZSFCY5
F3VHextMTtLxXhzRi0w7UYt55JgqKbkXU9hChniD6t/Znvmp9OZHEudZQyMw/+IYM5wr3UToTduS
OmYELwMZEfv4gqt1gwa57BHlFaFF3JnMfkfK/HwBbhG7mzsGEFJqv3HR0K3CfmCb1aokR76cC9iz
hcs3sYP6VhbaTkbsXwtTJna9MWNEOLdEuZJ9vdsVfY/M+UuIwUM4bTwZqpWs5cs51oHEFNVCR+eN
LkvNAcGlf9CE7Jis1mzBL/8aWSOHZXsm6dMQ64tJ39wGc99cpgiUemzTKDTVrsa3RzD9xaEXqzoR
Hp7yQm4aEVLlLaV9i+0RV7kQkSVJXoDsDvTm+ZLcSKDxJGKEv25Dz61ImT7JcWvZHb1E2jolR8St
iAN2DRfpa8Ded7tlOtqDysn2uPv1WnEK+gdvc5fJ3KmZoEEa47c5DB02hET0sIhPEWkTLJe9knR/
swW0csaQocgr4ljQIRADUn9x2V9X9X1R6LBBs6V83o0sXZgl5Cb92kiDsqrE0NKaQ10UziVDk/m4
vMf5yeSsEw4mn9m8nnAdbX80h+u1o5ODHyAzoyRFVGdNoNNKR4XBk2m3woYx9hDJxToWcHiV9smj
eFMH6qKjV2xGdH7U6slFTRI/9k081Jooas+KlD0miLQAg5qirBRyQkoFaMhtEB9TW2Hj3EslSJ5+
jg8exnByeOeHPFVCZPjDnk7teArNQ7YH/I5I14Xi/3SstcPHaXnYhdWtBsI5Y4995XJn+VpPGRSe
apOZMrv7lMSss5fmb0n7ZoBi+z181Ze2xL0u5IqT/9PScwJNVJrOyNVEAkfSooYG5LDS5DZ753CO
Ng2WD3Z13M/VvfLshPNgDae5gy3BRpxMdzj6W4zN2w52/V7wyNm6Hpwi8MDP4r8clIONpYJaSGLT
uFa9R2sTjId9sF3ulX8zGyKhg7LacDbZdGRPSw7trk4jKoLv0v3KRl3se7rrUG5NqGFPaWARHXbV
peNnxE+9pbO2teCCg+wHhWBmrACVEnp2FRXYqbQPHCARNpcUk69Zj9NtgmgiZIqSIMNkDecUGxpn
xcJEajXEPZqqndRi9xWGbb4DWx4MPFfZMCNymM+AXKRmnBrA9nMQULm2SkcMOiul3cvHkOnF9ykO
MzGxuzrEY6pB3otT3n7fq24hq/hW0uzR9ax/gdpg/nWFtSiO88kwzSZgMnhhH/EY+O39kRoZJj9l
9OkhS9hCEuDXg3pt/nWq2kFOravzqjhCHE37HiV7WVZcTZbDe710E2w4iXGy8KMpXpIUM3sRwWaH
jVwm5o5F2opY624j55Xdl1GP/BaE0F6d7Qr0wONIW7DhUAdekKtgMzrKGH1KAqf6rxWshQNRiLXo
6EDbLyYsYsmxHvmTI4I/FZArKOtk6ZyTVlddXc5GyaiB/tbOlCtkU0eOo3VNzxGFr80CKmSem3qG
QWgVQMyaYJTLQ6nuQNTpy1Td013Py6Gh8J0RfGIi5zpNQQZ8ULFflWaw2MpUmPHNHnv6yRQZuLww
hFt4WwoKZbCSZ8U6aBEYz6nwNWGPJA8AjNrYievQg/4/3jU4c7S1RFf9K01z1Wpdkh5j0GOhIW66
q54PC/wTnrxWFv2jCDGjaemAtiHSK3aZKlG3zlQuw7cFBTOGZyZulp2VUdWRK7bMnenGXE3Q8QTE
iGV8Sm9z8rs0DZrxbA+XDUFl2uEoSWWnAZ+0Xy/BF9dsjMQIcyWXGGK3m+aswHswtyJEB3dg3++r
ZwatpzzvGlqH1Z1OBXSU/oLSmPcGHdyIW4kQ8xt1XAHyx6I/HOGgHAueoxsfalhTOTBEGs6UXwcN
hCyKZd+BW6HNoeu27xvzNgkQLkXXAb2OCKiwJKGc8Ue/dXm8M++jHmJp+u5NKw6HPCu5VuOJbKOl
iDmoZoo2Rdy5DpJO2DbUUrwCNV3jfh/E7A5/PqCZ3oz3/IuQlBpHRS860BgJBl4EgQZQ6djDx3qY
boBN3HdaCavBD1qS0UtYI71OtWpB4PacW4dMloDmTXz/8r/5eeRl6ZdKfpqxVqX85/km6kEXrkU9
ckaoSBY5LGFI/MgFafMTeo4UU6NkdRM1tMAV69KvrJ9g3ye1EJasUwVf0g3NLl5UDSYQqDNvwY5k
85w/sP0zPYJHH/yeur+7wBMgnBW2Pbx9sADAD+ugkYnZSLlOcSKaMAFWtJcmjO1Jhy0aXVYObPzN
Ffrksk/Fp6wNUXTUa+Jg0TSe5j5Qwbp4BXZ5KS7rrxKR0VN+9adNeVMikbKj3SVf8+xNK/unU2Hm
dsZnxEr0aXnOE5KugmqFsc72E3ilHeRgj6UFHQxuq612O6cHzGZE2EKfqSL8IC2cWoaVdbtlP7Q2
yzraf/RUsvWKzL0tmxAy8jjuyT/MltjapNMp9cvsjUA4XXZCaBseY3PEB/TsTLCXL0jES/xV0nV2
nvzH46ywgBbLvNo1lOg7dHOZCVuWQ1g5TPtSFyFl3Ho8V5cfUFwQVZJrWI+5a0jMUZmrzL3dkMTp
bzA9RVcA45+wYIE1eqXMgvRBFzr/ZIlRLfPXAyLlP5nNO2iee7Yx48QM8Aqjx6dRuT4+OOkQMY3A
wloNhqtCN21ZauHmHaOOsReSNSA19t9kJXhgj32Cz5Boo3qooxCt56Oj2UM2FswADyXY024OxGQS
VB425tXtUamU8BlMRPkiDnf5kCLZdaJlJu5pSS6cBQJYETQolOiJDW1UWR6+JkBq3//3YPIvvPB+
ataNFUQjFx2K95jL1xuncy8aERcAU5OU619dkfdtwnU5rZE0ShC8zykXnHPSa6uoejPaQD4rNkeA
MgrrOve2ty8M4gwEzDF8tUcWgPM8S0r5p8A0D0ndke2HxxSXo33arxjHrVrksIGRtOLknONCD/H5
zPlapy4XrY/aO3mTwMNRCelsTEs4l2srX0HCG38Hm6IKP1iJB5DPfZyi52lHX+wRa4Sk8RAdsbG4
zGDzZHsQMHlHR5LnV05pGf2XT50HHQ2HIP5vdNgjG8TNx7Ke6cd37GKQvNzQznJFEGDFyibqrtfm
eZjfebZNvPf+MrnEoP/0QUt3aG6rCoZYi4D6mBr1ndaMyTscrmFbaGKx+0/qjD2eKR2LX9mNLB5R
5I2PBO9XRZ2z5P63ra5VgCRUdbeOMt42Z0kQCWALiT8S3VGGY1c7s2b7ls6Ya1qgxP/4FdrkpNyG
qMahExp0DPjgE8EavqhsPlZjzXbuEWDJRaRGQmaI2kC8KVP3j0RjqNwmkqt7rOAQL9baSyMuftdp
x+G71MGD5hkB85gQxJWAhNw/3W09KMEImuU8tBTJF8XejNr4H0CCsYVMlTEKwc3qPU2SHYFOd4ji
TBCKGvR39ZAoQKqHk0NMONn2fpkKlh83zicOEJ4Gb+GmO+dB0hCPcaT8CNo+vzuaEHZ9J4fvPyfT
U+iyjVmulPzvKjfdKXepo8VmktsekuFQfLDVJtEhtjdOi58K04W75KFLTTwBFc+Kk4oyC7QuQlki
MDeAwIm5P1zeGo+h6066xMkaliQoDB4zlXOZUcFQ0bruWHujl65+lsyxlsb7KojUB/LhF8U+uViO
qXulRyENB2jxS9tly4KnpOvjIlEPBuyF+xPhisKzxxLPHGsGZbXZG07ABaRuYeLH9S9XtQOZLfJ2
W5ttH6ghFUJ0AMiESEmOWEL9+iNXEpJ/ciFE4OTP3qroVacM/a0j0cpei8G6ORaBri018K+n+YDi
PP6k+QcPdVWe1dfruo0VsygY6GNuw+mbZzPlIkKHHNEvm0YF6t2F6vU94mAw4wnyBmcacXIAvLRF
NjEHa4ycV5Y5imD1mJ223XHeWqKsc/gEAB/u1qCtkDpzYujxkI2TJrKKcEEUPjc68pVqW6FZ7wdb
TVuudEeeXv14CnTd1jYo68qjWRr7uc0YPQLv8J/uG+B4HnRjhNlYhuETPBnDc+OKnVVVxCTzUtUk
cxDcNiuN1MLlYBkeXAusdyqqiwdCqtaVxDwuE3WzSL3rnA1SAoUr4ZWFHxJrcFtN5uQXwsjCy0jz
P9jWdGMRPPv6VC+2lSA8Rss9doKddG4K+Lrz76a4xi3xeMLzfYFKsTm2c9Q6r6p6hjNIcC4NM0L7
EPqvFlMiLMZidUPIJH7k7XcSc8cHjER7Im+lK9wiUilEUW985c4FMQa4BzbaFFIHai8ltHZcMg2c
ii6zQ3SDItoub9htE1GX4lnC7cnxQz3dmtLV6yhyEMNlDa9jUk4Gmanhz1M4T46rIQIULtOSGkHN
ioNO8fX9BZv3E2gEbYgWZvJcflKx0XiBZes7IRkwmtGnL4Ab8BA3YKgEA44NT+A9jYr5bHUpgkCG
yGTH0ujVAMLYqfw+5hljvHZMLHqnh92hz/O/FgDgvpz5fOn2IEH75t28kpilUSpI24LBTrbol8o5
TuJTwr1yUxh1CXEzNKtegrSqVPBb3+vn0aqHeOkSgBE9DUscizB/mD9L+Q7dip4pHmXHncqEs1Ve
MHFcNK11MGq1VRfwaNWr7CQ/OxMcH/Cv+N/7yQK+2Z6FKOh35gnT7Az8tIWl58djdy+MRDbK6jxx
SMVoaH1ITxEVC8jGLIsvNt7aX/kJv43U9tTrsDufANoZrK9oy+HqBy5pJYfL1pYEAdhQ97ZyldFs
v6Ckb8IRqs/eLIYa8rpYiXEezcgtduJMXOKnbGgz6oH9qpn1mtVmbTsBVJqP7QeK0U5DHLDzmtSd
dpahREqGJ0YIe6p6wIHIuYZEvZtYcr9rPt1ymw0//aD0d1vnYwQViuqXSyQAO9KUGfDU6EorDKEg
zqHsgQ5KqZnba5iuze8gZOz9iJf5f6CjFez1GtBIUjGVuz8RVsCmDa7EZf9Q+Z97ZC15e/VfqTVp
ZXuZ/Z3kJjTGPAayiHxSQ6oGHQ3Bre1Y+pN4XfgjzF/ciZYeiKOj5TsOP5qyqsT1fe3PrYzPbWwA
c6GizfeSyWQxa2IAtQgBfW6Rqv6YzrGnvCoAGtSVm7P2lhaZwxQaMEnNdb8UAgzwHYtJWfr3mumH
RpkF9acOfmOfYA7/mPiwvVjRs4EpeZbJPdk6Vz24RWUki2Q/J0X9ZGMBEAgHoBxhYfLGJr23P5CK
68US0g4hzJQ1DR46a2mgGHadY4fISS8jT/0giBSfxqBMKRdIGOiPGjnncThZYCoLE5w6r5ifhtbG
1KhomscS2AoGBw9C+gAQRxOS2DxHAdoVQzzYLFIPt9t9AGI0bIqGiYSfn16eSjmqxPJ3m3ReIKWL
X3MMUNwl/oH5PusOPWcycaZl5DWNOcJEdAVhbNM0IkKaJjOzdlnjlgRdGM/dgUdwwoUtPE6/XLHx
Hi+BdEU9SS8arfMk8DkIhkYWN28CHwa2dYg9gxssBz6KZC3FTc0uZ0HqOK94Tbv6CoCR5pEEyYLB
NaeXbOHJNav5NuJW0HqMxzt9tcJobHyKfjO44KKti+QP6iBYcZK2jTiEF4UD58ilXJswfdI4uFMT
V0uxM/ZDnfzi6q8KwHtXKrBpf+f4CsddBvPbuAdgW06YGM2K+CrOnZMMwfiPb+3OIG0l86ot6bjp
nl9maIVtjUw0Kng/4n2/i/QMXghLoJmCSS50bmGEl9nh2+RfD6l02KmATx/WURKXWgJILOiiz4Ep
Py+zBTMgBxuE92TsQpf43kb+uFAeG0aQ5QzALiP0qXAMMHp3j1fruyVxdBwgnvJ202SVXfds1WnH
d3+j4+X+kB7tCImQaJ1+g/+Bu9kjfiOonAQGS920N8MoZvkyUKbo3/olXGi3CVnFlFMvYhZ6u4Za
UP6rQVZo/t+hLwY9YntdYkCJhPED3iiK1tO39o13Ya5/wtsJMW9kmGyDUoSdSsAWMih6sa+S8zkH
n1FtYbwJN2T+hNeAIhQDw6BcJKT+trssJxW2BodEioRznNofXWPiZgcnFSCQscO+nGJlVKAX/cbY
AWP4mpczrvPKlFj79hb1yTk8JnGnuHmmxAk9LijRcjfYCav5b9mCP9g/TY1Ku02lIKzpUy9+mKeS
3E0TWCr6QLbYompvfOABALX8hQ7wji5fCZkGA4hScxbatucRCf7lLkA0bk6SWhyiKThR5xTgwuKp
TC1ocNHwGMKBZvbiIXkmRQxJ+92XF9P+MJq5r/84O8axXDvl8268mOhvzSBq2400DNeck+iyvtPT
k0FfcYZFG3xVM8kKOB0QWmwt5Pm5YxzyXTZL0XrUFuIcZECOfxLRFyDfuw/b4j61oEI9XsrwvOW2
7nmC7L71QUWOEXLvzQKVq/R2BUqLMKOWwPfo8r4y/dHlSq9U9Qex2g7+9gsZJ1m2ULrPGHuxJaB2
RfKT3dYc1Kxh0B2+BJm57yj8F32G3MgJBdJ7XLxDscEiVn8g34nHXIbwZn326KESfvhsamJpvMjd
7vfeXddGCabkrAYHN8CUXc1j7QfF1BX/nWCKJhiuKlhFy/s+BhVsaFdve1J2/NANak8u9brQOWDy
Pt46473gzZ0DYjdDPASB8js0h127HP1W7jrrmvKqP/NbZeUWD8Dc3xfMX/Dsdxcwt4QomgpcbSoV
NHX+RfeCk5XQhucBc1/x7JzsUgPLDarQYsDeR2e8G9e5+37uzy3vEjqSwtDIHW/qreUQIlv5Bwm0
LjQTv1Mk6Y4IXaXLztFZq916IHcMlLB0fPnl8oxm5xEicFRebrKrQcAvVa/hMEGtLan5DQRrWqU3
vzj12pkEY98H5tzp2TV/W0yAmKjy/OIEIwHtVlUNNAXd/BVCJgE94DiIsluHPoN3jIblJvqJfHEb
QrBordcJMkTwAYWvkkGNutXP0FUsBiw8sWCDlbxTJ4E+msaapHvgf5MrYYjY38A4nYrKqFx/Lx9d
/WNOPbrCFcK1ls5VHjNMxXVJO6XU6TbeiREVYSElGvXAWUHG/aZrdA+05J8fzgUi86kd2TgUDw4T
iKn9WuKF/93reQy9zI9NFNAaYskbqMns+gV8u5BJY0iO81FMFcTZKVdgrMxTH4IEdjkTaRyb9FCh
oS65ur2vhVX8kRIWApTOytA5EEo03yK3eTsM6I8DvxKmySvdVFc9i33W06GdLmWI3AwqxY7vTzWN
Jc72egwrdUtn+VckpIobTCedmZBmtltforRTBFuQ5DTuiVonHFpXgak1dlOdrYiYIbkb6mr/bwhd
7yL3v/Hnjya/Jlt0eqFMME8i0WKhzautkut9TJmaB8XltwAbIKPrViZCUH96umvtGgqvUGEMcfT0
TTteceepgTG1sZnDf593tvGt3AnaZxlst9ORDW7HTmfwwRXYO5/2poFQVXBhSZWm8jXdxeYpAVL1
L2M17CafIlS8ja9SInbfFlvYyTTmIP12b5qXlMKrOzkwDAIzHPe0NMx3xPA7pY+6PKUG3hgnmBKS
pLRSXLlVd76B1eOZM4KvyFBW4AJzYcuLOK0BFk4VvNrzk+36mGtVT0fRact58ZdEJLdXxc284CG7
SkU+YA/Qn5Uw0gcI+iy147vIYOxi57T2BcMMXazhGWetB2hfZDJOu8Za6QvpwGDMELxeUJMSLNp4
yNu4Eg+DCqsfJGgOIJ7YXMcqTNTg50uaIvOISp4OSmstKOnE4QICq4kbEhs/QL5T+8Q8s1h07EL4
SJ1+6Zep6MY5GArMyP/BV9N2zR3xxE2TlgYCRL3E9wO7WTeeLJrmpPwKV/gK1AHI5ghOvXJZslPG
jxibcmILUE+4VyyT9sOh/jxX4cCVlkOEkDiQc0OdEsAyp+3V5D5CcQ68E1Vn1vrZ5w+xCVu51k1n
TOxTMukVLV6+4efKr+7KmkyoNZdlNjVSYjEzZB7P0rzAlIVk9UgQlagj23KMLWbsXSgGGGHEpaEy
UbS5NDpuKwc2pjGwTpCprV6RFISDqRdZRBezaIAy5eVmJPsvfgv2dSaXjXjNKj1NinTIoJ50Vwi7
+fAKhx7bTMDnlyNYZdVtSVK5fJLQhVC85ijvfWjK/HSJTibIySfxaUjoKjOBsZ56dWUbVO4tWSYp
kYECU/d2Ryfaw78DuyBB9WTSM6zbZjXyRd0qrpI3Nchb4rV7UITCIWAy6KFM2mptk3kmvb8sMQkL
IEn2NMS9EgLXkKSWQOb1UlhU13ML1c+coPwXVlxiY1VQHRr9eH17JW9vOx/eL1qajy0Mgkyr1bEh
lbKPJTF8SbrCogsamyzgSVFOGjofCqTfwmP/Zcs9H+O8UsJ5rWR4mqNM7OdRijYM6Pw2U0SHX0zn
zoX+m47ic+wImO+ioAqqSqAQA7wvHcv4TMUO7EBnDNHtvu1BRgpvvKk9enBMX6FTW/Wrur4eF1Hw
2jPQ3uAAtNKXVLmUeeyG6Aip9klyqB+jBqqvL2Sm/Am4+HqwG96cHlqKglEj7nqH0QSqLufBNAd8
JeAi4V8vJ2Iiv7B+W4eTOOkuwYk5U/gwbyI3dnH6yOKFbTbrXHCntdj98TxDRLK3LpkLJUVqBXSD
DzhCiw40qhyWQy6INpHlF4FmsjbEcWNrf24O/hHIcfqUPpoXDaVEwvC7/A+HaMX7/tqHloSiKDjF
eK2UR71kQQwBEOkjVg0eW6FA+V7sbq3oza6UJBDaGhTSGg5ea1y91YSuvv65ozLeIG85h9/POpvX
DFecUkhlKglqdl3YKOaLRjlZiJivBCmnBr48KaEVZTIn/gl5qc4nNPauos5mA/vkkypo/VoOiIrR
BNxnQD5jo1GqQujRTL4I/AdBvQuPlQeDhUtTkUJ1/j2FXf1CptMR43Qg3IP2TL3CBUYBxwLjIVsd
BpZDnx9RvVvRxE5bYR+X97gq4HYypoYtNITGNTqelQtNNm/sMd1cBDElbu2C8XrBX4zy6duYoODz
Kv500jh34HnArZLaHaujv5WssQs2Aa42cHou8gRcR8PAYAxLAWDn2szxpQ0uv6snf7gTIwOytsob
aq260fFLEaCCziqSWCJreNQA6xAuO1WG9ImwEuzjs/A6+KIKNwL6WCud1XEhdCzO92HDc90bnoFq
uz9YzSfS4DUyZQioK7fwJIswi+uE5gglmkbNi8DtYmt/lg7viLIbJ98bOkPy5RkR/N2l5kD6Ieq8
cF/yFKXrKLPWLayFhVZY1BTT2Goj5MOPqOFHd0LaskpJiILtxN3ALB9R0DC4+RbzT7lHsLPGtCa3
c43inbIonMTM4y3WXGT012XbyT+nTf8f7ygtQciUX62VYhxO82mwxdb4f3rx0Uz+xYlNqqSjs5Un
BCD6VGR2zDylbdmVQF3L1IHTq+xnAOzganz+1gRbkpHi4lnL7iM1gciFx9erONyWEaVIN7850lCL
iueeIWZAxJsdg5rXE+LCrsApIUhcj4EKmnKtPdbGm0BJlVombDi6U7iB31Q80WQWIbkx/80SIaMz
visV+867JJ6GXUU/uE2iZAUPTzD0O3kxosSmT3J4CA8NWorOnDLz4bd4i8y5XU7x2tYmfApT9ZsN
AUPC5jbdRSR+Voqy58Pnx46xIPNzspMaOp5RkwHcRarQ2qk6vixwNLbTBjI91vhJSQBR4dD05uLz
C8BCoqjjXadVuCxt0kRnv3gNMHlaXHh0lfQnvAvkUKtbeDmtAp6yHLaeCAGeSoscaBvulZXvzwLR
5Cr7Z0atEWTH+wVD0+cR2VSOsZvGZqqMHHLJTHG2+yWOU3m2Gx6uZwAavfTtjzqcHB46+r+TxhHG
fM8EHRRSpzUll0/LBQYfYwfLRqHBue5yWMoicbhnLRGMMOZu7pRL1cEjGopG4VtGkWAsdeS9Dlft
CstE+asBWiWzr/vpwjuA9JtJeHg9seb5w2IAgPB/+vjTdhCaTyso1SoGC8ZBFnOQ8o107CVIOZW6
sMPGZMfsUjXIgo4VzvdRl3EqhQ+BmSpYipIiT/1RoBAhfKZnaDnk13bV3aAKl7q1JwL1wFf3fz1I
nyu73MDcRCZK3vHgKp7L6/ofZGpdNQX6VBlEOYvxuq3Ae9jlSuw2bBm52+HPYf35b2YT21qluQ7G
Laxo5LKOoqkGaStOgdw9jYNp4JAGDp4KhaFU9zGmrvxr8+g2A6MOdYM/FIT879Nhnv2oMkUAAOzg
DTnpH06pOQu5kD9KAHV79HntXySMSXS7pMjffkxEq7orQqcFh6IMfkB6GDc7vdIGCH4Tw/Ca6Hp6
Xxo+1P/72k148gGpDIKikiBnTWON3wfcgwJG8AicU+C5zAnRUw9+oGLEmI6aVURuU9pLtEEk0O+5
t4sFjvNdB0VdS0H/6A7dbJrhAcGHXkjMghJ/8QyU1ttahqcNlXg4nwyi1uhFiN+NBBY1Hlczxm1W
+W8Ih8abBhi9oVON/ignTOJgTSTh0NBHU30/cbGQGxdCJvpfL1chffS29uavL30VyLmgtbmnvrGM
ibLLqXADVpt5gEZ0GFz/E2elliNJUZulE2E6j8A4lDnX1/xnd9JF4Ot2tw+G2XLLOxlr/+LqXOZI
UzIqIFsBZLulXAOTTXeqTADrUnGX4NfdD/8QXAfQqNFTRPh/lrI2qyC991L0Xa6cUE/q972CBB39
rHJLTbYYYvbTnZNs3wxBdAryj6185ylZPH6G7YZxLd4YwFzArlJSI5LdDxUtIQono0J+4DqzJcLN
S/EEzt0Q7YsKaHpBD7PQ8FIsoJEMJf2dvoT815C2Vmi/kQW4NKzXmz/qhAf5Q0H/BMSJ8OqASm8h
LWfEoZ52kpLTNK0pFHVkFEtFwpzjLiSVG/Igzo8evO1K4ILOMukxfM8WiKIafrdY36/YudxgFr8R
XCg7pz9ljpc044SyyRKxUlyc7VpwIYXMyzAq3DBSpDtRJC4U23SLqlQ1/cpTwcV93c6cMlMKKWFt
I07LdjcN9Sm+NRLOxKeVRbNiHgN3WnB2iuaeY+7msRCUsN9rgh7M8n7RmiXE3g694cRWZgYU1vhU
gTIQXgM1Nxlm8Fj+kbfhzblZT92hnif5hB+cbeq59wuY1Hy+vpWWVjwUZRlI3MkFg1wm5QM/Xx/r
KHIYq1r8s5NAg9bxWLPms3dGf2T/ga8rVvRPzf3KT1P8Npjgqcht2CytyDIpvb5U0Ro8de8koYOB
IN/EZkKUDDqjNP2l1u4PHBRwtaO02grEKLCCLCxYJl/LbjcpVoF3w/EdsIBYpcQkhvluCFgOm76v
r3VwcCG6IrTz4SyvqeSKM1+pv5uHizuQmBmc3C+WrsKzO7MOjUEyGumaOD7Q2/9capT+2cEgY+Py
VYNu2Ymh/x616sGuLReSqIC+O2ma2uFQMCcevqGMSfEUtsdOy6tYINTP0nNDCVqdZ7zsLH0qqXzp
mLbbK1MXmmOsyxNLnHBKUu7JDK62ZxyEBX0xzOZKS6WZHCT+rc2Sr4hkP5DFkW8t6GD8gRoryucw
AXvPN3mf1+XCD1q36zlTtY8IenQd5jEoVuzc2sKj6OjwB+6iKhaIodhxtODQI7vnZY3QHxwDe6Pm
HylAkEGJuMV/ZjtGeOic8yLJu+6m48PzNwDMCub0K4wgMwl+Lxqx9wGn2Bp8Nwu/eJuMy3BO/mi1
cpVqzybTkKmaVr5XEsYQDoRRa7j/JEgyKxivBVQDa1q1/7NPJb6Y898xEbkLUV3PZjy5oDSUht8m
YazQ1OX0KtLhQRwGZ055n8KWBKrgHtgYxxXvPCDrwb89eLuEcoYc4r4oINaXdzqvwICIsuoulLwk
vnNH8jqvZ55VUnZK1bp3h+7dczQQplQknnNFcvzeVi9J/6KBGVjCQTC2StHsmsfJpYWCAw20RFoq
QnrCBOO4/L3wWehdNW3psb7j01EKkKN8NOjFh1ImN25aS538nmNObOZ4cDcBrAZOLRs8x1a55ZZt
q3zsWQCQKzCyyJPiW2h8aoOQdV6kErR1yEQJcYTGJzSJgjRf+0qB5BG+YqlZ6dTu/hiOriJ5kir9
k4ryrdZpJCGcsc+Tqd4ANZXxHA5iExuDHKhZBJkHoXKJ8rOnMlr+Wb5R6Zmfd6f/E9j9SK3ZDBga
PdJ0UvOq/c8Cld5Yrplp1ihkp2NmOxzMoy6Sgi/fxP7FGOhwKigF+llutpiya382amH8s/QkR28I
4ACh+uJLZZpVLRVil5xaEyJjmBXLDyZgmAFw6R2u9QlOvZDJ1s/Y7wr8EBDEhewAxRuBHWZ833iw
qWEpGI4dsxgLHmlXSg0zT6u9owrSblaoj6l4kQLq7oD3kYRH9tHFP476lo/xGiIhYMJD1hDlBTCm
dkpX29+w96EQVRh746ABSW3DMaWi0NbtV788U6sbOEEXoIRPEJAnRtyB/QNpfgXS8Ff7QgRXjPes
gSjBG6ePBpC15bZx+Ld/GVpwhqOYHt5uwQhv+99Qny5n6tTZ9ynp4H/f4kQsGQtskKM96OEiNqOH
fN1vFrWYAjh5IWBtoGc6x7SHZIgegb+ZarbARvvp8u15u9z6q0TkGnisGDjtlC/cH69gl/wnLwV0
b6SsgVMiGtygCIywSgIZzoOGLqA78KtR9nudX4WBHXdKgmbIzAliVmH1xUKY9UzLyzAXCmePYAE6
ai8YRmbDR3746JKCmmRiMO7KCNWQSxWBugvxzwY4gkHFmBli1aTCkG4o7OLDz9tBiN3lsqxlI8cQ
9tzp50ez5IxJ8trJIHGR2R6RGx1Y8xwbcHqduj9tgxjWPjrzzLUrQFYTv1Zmt5XAadXH5XpsJeyM
IHN+rFqPV/aKZ7IPgD0YKT6R1jcDa6rchN4rmbwhG5X4g4Wp0J8RPFpg1YI6mrNUfvE2Te2qVvX7
TW5YAvjhspgS56tGsuvKOhg7Do21nw9PijMqOJSfb9WqW6wOZ3Rbtf2/ftnFZf5h2wdgHCd9V3FQ
aBhU/5INYjY4cWmi88cDQIK3on9bRBH0ynAgIKxJL8/2WimWbWYc/0MCGvLCtmWK7VJ9u9gos2KM
Jf3ypeW+DkjRlRj/26o02Aap4f22V8Hrel8w4jkgL6b2jxeR1KSzejTf0/t2i2EWDVKvY1iUl3ot
h4RWDwCe4CSyoWw7aw+0NiRmhKwbr4xpzOtKcXSwg0R2IM/j4uvBZhTE1+67sIo6fZM5f9WPjWnR
Yh5Wj6EdyNQUOgf3TFHxNBCZltFjVpRAOoHswBGvhD0+SYpbaF22BkB/flVI9DZ1aAbo7NtIx7lg
Yy5CcE+PSzDN5C4JOnriVmuiei1ByMc4QC/j+JCd/ryk7zKITm0RtPF56VkM4AZol6MpgobXJTWW
2k2TwQSIjk49aJkadY9JdzfsbEHhalxxYmGEHhlLozfbzJxgEDQ9vyGh7ManA3Cc1j7STvjyHLTc
0aoBzf6YGDh5mQ7mVXHc86ZOdrq94Q5SYWUxAUBiAVB7A3VgbXJEbcWdFnUvJxDlJgikn+WEHouu
3TZt18GV5Vl4UXQSGThYhs+6Y+Z825hCaFPV3ct8GFCSk+fwl6a2k65cJfIbWWn/2FblzG5Esp3G
JhBplMjbBedMR5TPlOox6xiEXnwxg1VI1+EOHtrhbScg/so9nzYnnaAgrCR710q8FTZQ5JCOdZQ4
X7lwIkm3OJITFRCI6nJpxUpkkoQl8W2fhkGuLdR6ksTqd8H67R8DlGj2aNNQOJlHPfc1tofSB5QG
CkXF6kHT52DZwT3qoCvySdr18e7We6PESMhhB0Zv9Q7KGorcY7EiP7n7dsnT4jowv3b9XKV4/XJ2
ivbqv+j5F6OV9b5ZQ0Oljp7i7+ZqsnAeTLtzAQDD0IzVKrw1+W5trfG4lKgS5JU5/yoSrQnDKrQ+
Y4CE2oKSD4YzIsAD+lOeKQmmJIrh1ZiQ3JMd+BaAeSY/UmPg0tl6fFrUnkMlpHFTLuNcaPkFsf2y
7ZO7xRHkKn5Rvij9ZrL8NQtq1d9VtMUspRDPYtvkp8nLvWzsEuIMiW8EQ5iRk9c5flvVt4dIV99O
WGBT6LiYksJWBhcyLSC05flDqJWkOgyPwXwWTX0z6SxcYiy0FF36X5aR3Qho6wUfgXoWpPnTz+NN
RvHd61rEF3H1gmtKEzEeVm9WHl13g2IkrIXaK4fSU9Y3jxsRIZvipZcC5IYruRS9A0mEp+b3bWh/
GPj1Lrv5qcOkUwMw2g/mKowqppmXK57mroTkZJBFa5eplfk/fvcM2rDQ3trfc1dMlQ8UhvBftGIx
RdMTZ34rI6Ad0eecfG0xanXTPMLXX25Iwci91A+DaF16Hp83tg4SWrmUZ1UlREA0eFrsvQMzf88o
K5pEcfy1ceaZENUkT2NUaMZ5vCNFqtyXB57V+7Yjtz0yy3yKlXQ9561XRJEXNzoiZWrXIvcMCN43
pzq5Tlj3j1rCf+c8GwSzDHeQlT8Y/07ZiESoOFbsYMO2Zirum6+3G6/pOvq7hYrWSpKCm3w3KooN
xF62eTxHU23Hoxx+VnXtiuuoeDjGyqaA2KQiQibR2r8SVInP+o8pkevmybT53uEN+iXlVEgV4x6K
xr7KRVKByZOTtNoCVyhCWlb8oLF2nguuGxhqwYT91kASCCMuesBBRgDH3XJjLYeEHc98ZFw/D8rB
eQVNX3qVA+NsErN1IwbKq9SS945H/9Q3u7cL9O0qD/5YeBa/MX0JFrEgw6yQjh6fw1mVAUZ4PN0A
fIxUwyrFEFyX3wLfCrWhb2YTm+lJkVgHKo/ssSOOVF6pvK6jvw7Dvp19eJayyixWoRPk25vEBbte
ohhfw1QOMGhpBf0637m9MuDUn4236jwyPEAGl1t7KK8ELlLXMQWQYpZ5AIL6ruKMOPANxaY+RJ4U
ZZ66AQbxYER+zTQW6PWNhJK6+UMmqysP3aDhWL8sFrh4wnJZtdsVnbVRjCPzwimibVkRJbe2LftA
wZFFNrPM2TIfNU7S8lGSGNJL8SXgsMCXjtdcqML9wxf+SA4/DG5H1WhvZyEfQlXa3rI054gdPfOn
9ZEI7m5NrHl/xIudxuaew2ZiPD47AgD5LfRFuzfZKgnL/KGTLf4kZMF0dNR0YguTrH/pRvm8/iPq
S9mrRqVasvMmTbCS3WgOYpSvlp5iG2eU/VhpL0sSUNiPbaWkcK3+0f59VHux2e2d0Q+2F64r2aOv
sTX2zHqThPPr0KOi4ADMcfLWY9E2GDCZCGWzwQ+KqEa6Z5ZjmjtNLvzYTdLTsfmck31Fk6LOiM4Y
2CdA3bH6KtHbMeYZB3OV4jyE7AWEYL1veyQmiNZ2xz6GE1jtHAJJAjp1DRav/L2H438HbnwnwlNj
GCxa2Jel5YgQ1MQHYv3YOe9tFS71qFb/phWDe2Lr7uu343FaJX452POFZ8kA4Pj6yD0FNn1XGlIM
3y+BlslzFpft6Szwlfk/4pyRRXwcuoyu/mAGt63QcuIso1U/xPWdxq7DSnCrouEvVeFyjjZTKW4U
KSnOfcQpjvBsV9x/CB1KUQQd0ARoFC1O00knaH6k8Qd0TL2dwVeSxr/byF07/soLZ2+DctQHszlp
i4LYYfD809ug1sYsmbR5laogADwXpuxbcXxzVWeIbGWKrkTYQFpAnJc/kSK5vNyCqoIuJJ50CZKZ
Jl1UmYbGU7XkNLNIE0AbjArAv0GJdiX0BsQqO0fCm3QXxxDoZIiIWeZcnjjgxBK9N7Kg1BJxeh90
g78FDLaTc/vV3vBdt9bMiW/2q1YOlPDCUI6Pv1mkbBPKGIM9cHqJgosQSSbKs9KctdO5VhTKIXcf
X6lNjil3PGw2fN6h1dle+7kxQm9R54jamG4DCPomyUm2PMkA8id96cq5Msgrf/byMHa+s6o6xqN6
iYPMUcj+wjWRP//lHn78VsTZBiDs0JpYXUljWhjYf0KCr5O6POb6h+MGEf4k9Bl12VC8dThweLJo
VjgcDr/NYpEO7OsQV/oy6paVva1KNNPFQ4E2KoQ9DXcKjTvEcnTf21Xpey0MdjXq9CAL0HdbYiRe
gX8vq43FXV78547ydpCVsmoWn5k4xolkOBqRGINsPp8YiSXzEoBXffWLBsS+bWVon7Be4zlaKVFF
udzkmIAg35LAeKT3b4dBPFmWqDB6s3AeElU45cyYggiGKvzF6w9LupeK+9kxazY0OwBiU6uVPFby
4l31kTxSOilqnefbOfcSEM+S2CUw4QBKWULxFtqSVGPh4TaoA923RnoIwtJSQe4a6qPzZYqT1Knl
ztc/Eo3cpI1OIRqa7UfM0fCmzTRYGae5KhlMy7IVYOV+fw3R13ydWeehd9YGdzfNkzWEEzIajczH
+a/8jNsnSK1bt6RJiIro+85qTUfsNAvdPYXEBOEw6GLtoA1gn1lDkqN1VxSZk70AmEbQxQmUi2GH
/xmI8Pg3NtTafG3LlQIeCCQaJM3Jcy9loi6jMmWRDW22AiLPag89twT/OYdo45ZdagiW5zCLsKoM
GgCjIdrzfmC36X08YFbl5Gu3j6uwdnaA76aDjJjSZi/0tT6HSbi48Mj0W/PHEIDDQb0K6HcHAQvk
AQDCRe+GzMcm55ZKrZFbQx+HJRo9jssjrQnqTbwqpTAUxjb+Vf6KCywkp3YtYkhM+PXWex+CVfXK
/eOehLlVH3plVOe4LFsnFREeYnp1HbVNj3NR9X3f0poSlD7TKTMT7g9dfXcwalZ2WcT9X2X4aw7Z
wKP2orDJ4hJAUWQqFDmD9Pdidtm6TijHLcZNI6AARYf4b4i/hee57Be49qUifOUpmFP9X2l3VrlR
08xeKcJxmt2sZzGfctMQ2+R8O6z5pLQAyXAbVncuEa2bjlD2flmd5+fVxdBNZkS0aZFzDpDq3+m/
3LscssyYjISlU24Nf5EMLZhVGP74gupcDn2j/zqotgWpZfvtCq84FhrblbIV+PMBzuIsjj8FOnW0
9/on1AfrZnZ25OjTF46+7o89HVgAxP0huInZvm5Izg8Qz5vGzJ0OA7CLTUGeyHNxGbTXNlpFVpJk
RVexwbMy5yESyJ+rBw5IQSeRJXtnlQebLpntzE/MFVeaBEm46Zcl4lYYCjCK6uZzI+E9F8au0gqx
VyrHIT0caA7EMHLWqLX9zxE3O7BR7YpPbVoJUyR44QOio5II0c8+bg+OxXYRNB6dTFSG8fGBcgx7
/Ocyw71LbWjH1aJijoZUMMBcw2q4VHGAtk0N5tQhqJlyPgdul/JcJqTfmQ1mQ6vpkkGNycLY4FBT
lS7tbxe+XCyc4LQPSt8qWGPVhqajzFAZ2NsFzxUK8n3je5koH4OjONrrLQOhTHGJDzgR00t2d/wR
3Cc9LdKpn/JPouChrUA9QXUxFsz9aaf7+BWxxym7oPUQ9gnKgjaJswvyrQVt248vL3ByfCxU1XRI
DY0Mpx4KBALLSoKNYNMwu0ZBGiIkwE/lAuW+7QiRLYNW+F0p+mROyg63fFg65C6XLJ2pbtEpX334
qXsG7QoDsNKnpz4j1TboH5Hv/gqEM/8SOTbS7IosHeWxOfEwF48hpjjEYV0QExp6CzNI+uAt8+xZ
JQfoatD+RenSzznpLh+iu+8TQg5/8tsr+hVHxVgknR0WcVc7yo7FxqWh9nMV6Wk0K+qUE/sFd2Cw
lRQB4vfRlsTUw6yrQsRLpD6uR8yzLx7ZAPaVBfLj9gQ96+B+7YTgRZE0QlQXZa8WhlRqs8cDJ101
5Ofbu6uc/ef/kIgBXCJ3wwLbePdqpGrQZFhL1IiPVkLR7pfstIqZUjv3LNCdbjAwKzPDpkgKp/iB
KrEKRtWEKY4F0n/awb5cIkYFAIL+uZQCXexVTZE/N6Wvqzs56dFaTwVXhy5E56RK1wPFNLSSnZE+
y4iwi3apajaXMQMRbZrRYE8bFX5rqK1vTw1H4eSJKP4Fu+/0TGgPXfZAvbIcXU4eerufoZpRhc2h
n0CbIQVrqyCoXmR1WawwOi7TCzX9uPYbAZ/683tQekW1Oc6jjXMk7MqJ5Gm3+BlQZ0tV1GPHtApD
7G0FcJsrWKhcofdY9QzgxwPMnbTxRXYfBEiIC2TBowVok8HRk3M4mxDX9KRXa8vDKKe7ZxaMvJFE
VVeZGwBWuSnHe8xz2z0VZCJJ5iASJdhBENsYSeK2tgP6rfC53gZUn1G+gJnboS30rCC+f+b0a2fO
zD7fVMc3MEombEzp8UAeVlgg5NgOjF6U29J8OefPJV5ZYQXYu+HPj5eWZLfeZVmeJa3GTeMmuiVA
BC5G3Vnzlv3cxe7ofMuDKvaEpfpD9fvo+MOkzph7TDzfKw24MUDzYPYgOj59BrdHJb+0vOOgGOjE
uZF7CJk1DTmlz04sK3sVuiS7Wq9pLoSkRD0q60SYGvdnERd3MxRpAOA7iAjFV6k+uvx45RxXQeab
V830HNzbqbSaxRQ8r76AGm5DAeZJXK8QztOhBdaqYyq0n3NO3eEPGWT+Yt6jaYXkroCcsytraKW+
VUIHLImQNuY1vt/H4J1zauY+SCCM3N8jk7jumc9mXMNkxA63bhd4GdreqQGZ/8qCYWWXPAi46tDN
yRou6PSrnKAQYr40Q7N1f6KQzONtl1iQLk4No0JCSk8TCOY4SaZmm4Yu9WwZtcXf+2Ps6S2884N5
1dUw8Ons45QPZIWZGoN/3COpwA2H6fY8NEKUR1gIcI4Mgx0RgivvL7fBxy2wyTv2UBr2mrquXocJ
8NRcSlw4x8neQF921z23yiVi61SAIvqsgsJa4ldjpfxxnMG9hh4u+b1PI6u+oW6rL9nP2GQz32SH
+INd1FcYMIqXy+kFRfO/JLbXzuwtH7uVkHoflbbQI79H+769/MowwD/zBTsetoPdcb8O1DXp8YjJ
VlDnDt+a2hUbU52S3SsGIeXbqZaC+wiD7yAaJyAdZ4wJNpwCIcfPuw9nFUMkvF+hxtuTQdxA34ni
4eg3DApWParlQc8OdQX2DzNQEQT3MJwIi/4/k5rF/MwTWtos8jvvQEYwVVqA8TYPCF2XoTjF45rW
b+pplGtaUBFk/UXwTgsbWPKQxNv92DHtcvy2vMTA2I8a8660TIpKfnxroag5WHHJXUTVTT2OLR4L
eB59SgGPimePd0wqeqKdjCxihXjYG6J43SwI8sTBn4scgkOGdxa2WRw3z7L/kH6cSk1ogPperLcC
yU7Av80TFOnjUlKftOqO/jM0XDD8L5SYZrK4ZfMde6srs6n6gdQ6ATSFQK5URy01k3p008A8OxJc
5DD8qsrdGG3rityggFYG216lmbB+cFVIEK6vMxy7+LWWdhqt0JYN8w5Hgudluh2fSsVgt83ZAfzc
7QIGUdxrAuWZMetFhO+st+5e57/rfKSrdEFJz4Ke3Cuj0OrELBF3K3ULth0W1L04pDCeROgBhGrM
IKIu8uwwJABgQrKlKdNNxmglC65wOFyLzluMcTNODrgOt4hjZTAvyY729wAzzaYKk/5fb2BWTeqo
uIiU+ty1j1d6fxwdUnu3UMzhEIDaB6jRhZ2O7QW1JhCPkci6oP1OxKDKmlrKAMqmgfudLfzcLKVm
nUk0Y7ekbkxAlrRTYkykK7OwLKAwRJZEDIIao8QaXeGIlXiOkGTx4G5GiYHVbOhmYjh9m9sIc/zw
3RN8p2cxBKupHX9KOG1D6I9Q+BvGgvP4VhjMwSneC82C0xfQBFKXFFPMqPxKLS3T0A+QoDL4whUo
KItDIymifd80S/y8X1OhlfmoNKfZiWtrbM7uX9lZs0wS0Ok5LDPqCxTI3TXM5mylB2PkPBMddb5+
Nl5Lp1DX04fr6u5c4SCQmz0e9Dt0nvKm0iYbqQTP+diW3M+FyEFGdnyXP+oZQO/hCyKGuQteeGlm
iEGdZ8T7kBFGzg8YPKkA7K89qdoOFaYA4YR2l28bgESzfwm1GGd1lGuFapiy2fwjNJf7XXCKI3VK
Y9PTlKY23qruLr/i9DU5u9D5GwnnWQ/bLsG2FS0mgef0p6e8krAoaG3N82abz3KHu1/Ylt0yVriY
nZTM0j7qmD8qZySS22JFc8MF5Rzvtemx4rJbwQ2i9eBWgw8w8f9i4AsSckPY98YFDz/fqrXTBdQY
0TFnX7u5EySQRKDW7reAePcvvkZYjMgrJIZBWPUmhjD75HN43/T2mA0wUPpN6wMojNTGL1LSV79B
TKrmrNf50n5/zO1isG4aWFGck6SmTvvxbilY64WMygaIrQzFw2meEpSuHS75GFxz9SxSwWT0hn0j
rBeGOPAzmNHNv1gmHsHWrYUXnIjovQuH//PDA3Idgt6kOEfB69LNI30k8FnrwnJrMPN/sULvCHrq
ItWtq7dAOelWSn3xOeL/n3oRFJZwNMzhMinTFpwK9oGMzTBmXnKrh8Cuast3xaHgRe7Th/RfyL96
EYfD0uq0jVIVNqzqdV/GiqMwya8A2KkL66Xzn0N9AdVUL1OuGNNNkGxUjlXdGLKdmgpjA/nt0ZxW
ROw3yDXmnmKhmzixWiyS7u5JnaAQ1+5AH8HcqPHXCGyU90j/LJjnC2pock0AnlmqthZU4UmvIVgI
Ak4NyoJwj6LlnxzF6GySGsxugpLyo+TMNaQZLlXbWG3EZkEMuURCW6EYhov7Ea8jgM29vZ6dN37W
0eOatr0BhqpOo5+xROFSuCUsRQY95am0zVX07MMU2Z7SsaDNbCYxR0mcM338kk1UainDqUQ4wwO4
JCqOCfBFK0NffeyzUJSXj4efgdeLPAYoAe26aE+/yd9Il9WmGVVIsia8UlzCGVw1Vh2Kit7SXvDk
BbIuKpwQy8AG876pn2vz4AMjK0cz2lgSaXcxuoyiY2PoQktxo7P/89OAxYZmbOCHxuAS6jW1vYxq
SP1NgvvyK2sB1in7wV2fGCmaq1gIT6xygcrd53kP+QlqnAZH0qt+x3yy1lauP7eKo+nrQXVYRc9q
NGpOHEVeMborZHaAyxD7a4X5bFZzcFFBFsTsCwOS+iAz7TGi1KW/siLdBzwKQ5FzK1m2f2wJDc2H
B3pJsNtf7KPZUPyZvNPi68n8BP3C+ZPua63+6mWQ5sPDiJJIQexRVQs/qse7s0EfrdgbdgpSIsVX
XOGieYI0vd3lfjjHuPG8t5P95PlBGKZp6L3VxpR4sQzXM4Q/Q1BBS5cwQuHGjR+63ri52awAOAA5
iUhWgJw/RoQX2dC6NiFxe1hUQS37DEs//GkWO21Q8D+jW2JlpdbLETbxaGoYNLiORa6NXRy2P4ui
b0/UPWwny8HV21zro+VblaaUzZ3OPIFe6n7zPO+bEl5swmWYa6wLaQCqQ4cxidqfM2AUvaq/dEfI
lBeOM8OYQObiDUg+lnCB65JH+dcmWCevPO57N1jG7bBFEQ3hvf28gJLwNKwHdzmp5sT50vR+AA6E
d+ntpv5Zt5HRbh0bKF2EHRVKPOVp4HMbdC2fe/Ow4IoZ37ng7VGpGyfET+EWh3UYj2BgENwLq5X1
EaHYTwnadzc/30PYroZ439d3Xiob0zMAhEl13AEIZo5wXJs82isEHgAxkyC8RHznA6E0gFWtn8Yy
bAa8Swo2nq+bojE0U9RJdvPwVlXl3U2vMDKnqWFgYfGwScj9Rf0JAnT+KffjWBYcun52xjNC4THG
g12MIxJJXjLSbSWJxlTlFQKM/kVQXcVRB/jwF+wlZJhdrUkke4RYBWPxmrBKrEzKImFs9N0XGlT1
NeUuoE50ZtgZkCNs4Ym4VjM8XW33lwqok0Rzr8bUtfHLl0cURjsoMMwfw/gRCob3mk8Jxg14bV0e
Y9h2mXXQbRH0h+s6dSHtTuDXreWO0bTGWKqgCuBIWe+CXtkqYPhlH1m2SJjI/cMgj7Dn6ynpOk20
A2QUOLb6RdLL9NhBY+2W5xnyFvawGWQX8ZiGz5HBTWu+cecfduwJ+15efhDCse5AopAALPw/nqtZ
kqhe8dXtOlxSZgn7TwxxXjmGBlDkB9tevuM9wGnigjZkkjiS1BQ2+DF5QNAQiYbkFhMcxT4ZlLaG
FTqVBjZ6smbTM4d2eM0vBXuvlNp2oSynjzofhfH47MoTJLh3oqfuHQYfPtaJUygq2BhvAww9PSmj
A+7yWwa7+X11iHYHh5795m6V4fC+xgv4V5Dmda8GEOp7OJlUezJM6CO69DCB8urFhcRvpvph2vgX
Wed17HuvqvlLObxQUnXziQOtnX0gJRN75A2lzOTeEhUxFKyyubUBaufN5tQqlCiPYeSXztkbFlTj
Vyq4RhvIhY+PQmsAKu4e7Md1OcnIcH5IFfqZng0mobDAdZ//HZV640FxtzDOF3n/iEueLloZMuYU
2ubGbp7cSL6yX+/ginFFIcZP7JPXHaCo/36n1ME0kAW6KVCKheiG4syNzExPnk/54BKdV9aL1PTr
hRT8UzWU4fnOlPZLFF22Ov956POLzm5+6W/lqs5gTp4tNm7fdyZPrfhRtLlNB7+BB5H3n58WRqup
grz2QS+VoMZ/xRsBEsHjWyZFOEOyLnjvtuXjeAUkq21owSiBeqgFAZ9aTm9mzz+hAGBzlEkYCHWQ
ThIDZoOtO5rS5KUVzvUc8v3BgyOzAObr5e4SWbujNe/hj2siFE9vH9s8nJjik27NgG8Lqtqo9vgC
6v6Nk6qDoWn7hJWdYUAGqLkKtmNAV+PRF9p6rZoBsp5KkhDLM6UnQTofSPHbRWeJqKWwCZExCbS+
7/iO+kKCipTXUrBjV0wffRwMrcUys3K0euEDhtQZuDU1uKsu93A2jnLHWFxD/kqu+s9mbW6z4RPE
ZvpCQrHUj6dpVui/WIs7k84PMm94zfdInh5cxUyRYgSLRCJ8oGXsGPDKl9WC+EdQVvjVCagk4Ame
AgZR3SrQCkpl4vwle+Y3wMkgtv2fEpsDPnm1SzqCVKLM+KHKhFUi5t+EOjCOztf16LbbBAsuBR3Y
pQFA2Odvb/gR1rtbbtBWfQsq2iE7Ic2jz26RMIWFcH5get3jy1mM8zsLQZIwdU3VSNdcitM5PzNm
SZAHmDO8XiUQgg0ZZBmPZnExVadX3EOtYeYdqXuthDyXHpu4n5bwNAYYcMCeJKy0hH+kuMLZ45gM
nHmCIgd0cUJWcHL5Wmmuun60ndxURSwZFKv6UH9mLRWYv38lvZDaaEFCaoRPpAcHh0SxIMcqKjwF
WzQXHkPJ41siBIKk1pDFA9//9ub0p+ZMKUPBR/0J6Lgl7jquGOvpRdSNM058LVtug6OKf3NVyVow
uE8g+Am0r5hO0K5VHHAAlaLjcaP+eEq7aKpRFvCMurIWITjf0sRwPHMaFdJrLuhfOaYJxBynqPFU
rA/h2XAuF+to4ppTpzZM9/nA++w5YiP/+ZLvaV8KFWVRzxtCMI6+nv01N27doQD3wHw5roEZ/ul7
U/KqF72RCKEDlkzcA6XN+tgwujE6DqlSzUIRXzzwr53ze2UWIZtM6Buq2pKlWNMcOcoyR1baTDCw
7JbGr5BGmq3B9nq1buHbg1R4DW+QzRqsiJwP6UHs+OkgXUQvtLl+ne5z/IhIj4h1SjTXqcrnf5s7
3jk0ct89XdjkqX9ECYKl+NTtCemg3gE2DGgMoDDKqbrFzT7FbU5l8t3K3zwqq/Y7Ixs5YCEaQoed
gfd8k7MJlCawBN5fydjVJ2llqYYJnbBsEPPu5SpSpIOj7lvHGBgse0Tgqz0m97cTGfwkI+ZJdLr8
xACKzbxj6yzf+jlAGeDzojomCsklQaPdSNrOcwxBuI4KWWr/Fr7BHLLBdFIfGMnVIQ0ml/KZzTnk
Dj6MPI20gfUw6uUUlQFUI0rbTAn7o6GbidYQA4dio0lqg5YKVgS091t2mmAmm5z7gVsZGENmIuId
gCpOXRqNa4arif4okEAFQtf0HGAThzTd8rLLIixSALBu3+2Jaqx3lBX/bvEfvK1izoQtHfHxkkCH
UEpcpjuiPbVe1HnwdafZBrSP0tqbKziu7q4Dl7PCMUBGqDmD/Mx6izv3o9ngGjZYzO5m4/utsllf
AugDxPu6B4JUoEBzWbUa0Iv6r84nCbMO+nYqskGVwJLLpQOjMtBYO8MiJyLvDcZil1bp4clEVyht
PyS9iVFtCKyXrBQ3J2eRsKoYDjyhf8E6T476sFN5c8SO/iKKR9bGWlFbPt8aFok4SI0MRib8MLEp
TCR8EXQR6485PoQhT1ab7Wp5GK4O+OaVKb+WRtC2uVa2dgCbphvInKeiV/6/an8fLe7/hgUqsbek
S3fR/LcsGTi73yIOcFJigK8Q9OdZLuDeHLfzI6C6SRqfleTrT65v1sHAwbhSoZ/YO7UGMB9Tbasy
iUbOtmk67MrcLVmWFsp9sGGwt8dltfAFIGqyRfu9PMDZ10bObfrvWayYSxIc3vrJfj2LYv+IsaaE
NKYN3Y+JgdK16VbDKO2fQD9Q6dW6EGLDY7ThV8BdXWin1UzjYZhGQ5ACEw4SkEJ0vc10Upj36kpx
4RjqBTWkZSmNgSddaO2uzoW5wwmZG98dojgoBTIpP0DgxMdEkcqBZFw6HGdmOohrLBTGHsdh0Xn5
mwdbPgmFQdp9JJbjb1ugfMdM0+h0bu7JYVCJy+VLBc1ksXDhybocUkL/iy/OTuwN1HfKsbBMiRkv
QrAugvkih3rOFmzAaIJxbNPQMUqVFPWiyY/E0TZSnlQx+8mSliWHgsFTNpdoQc0iwlYJVayKWeDn
9FKbI4X6HUarj5ex95xaXD7qx/T8iadqU412KpO01D/gitarGL8L16owZnSzHock6RfxNyJsGeO7
G41SK5kS5qJv1kyVuoeqh7y1USwnC4OpMAY9vUTZGN+O4yWx2/9hScwjNBFkCkWa6uMDKOrTYd+u
jnnTZYwVKxUwBpM1qHanBWicMNxNoljZ9X+LDn+3XxxmUV1+my5lj0UG6A6J6XOuwfJevNRj/LWE
RYA3z95Usv91RZxAunEyEp0kxpjf5mX9EoO2vlS+lbwCRl8aIc4OZ/01khW84hSr5kMYkmG6WSAg
pIGqA4lPivwY0cIg4AGmsRWZOHUHTpsdsdOJ5kTreXkIS0aXBqwWrH0CXVnLteo7jqZ1Vl2iWiZ5
AJQqSraLVoNo3WYbRSg48BiHEIC7sViFQsU+SGHjTbQtPeoPYdI7aTV4tg3oD0CI5PvPI6gEX2hz
VlYXPV0cgxxYj/6DKanSlXihtP3QudTAZJ0YbPgGr6erkVx7lGcWuD7sJPt/r5FoXBcq221chjnf
Cw1EK7S8Sbn/zItea0SeiwOLWGew46E6tv9oIRXx1iyZS5fc6+e3WtJeiE1p6LZqb4gaqDN1UvE1
X2jrLmBfAgqJj9HPZCy0Avx0yNToYxa+d0OhYG+rZFXCop8L+/DCP96w3Xv/dDP83yZHND2acN2i
0AM7RHW0h0Rjqxtq91SvFGJ6ownFK64fqFxdrGMFehMmLN36Fz/VdBaWphSYzCt4X7AENZJAiYpW
2vvU94C1endxVAz1Xg6yXMVqyMJqUAO3SETN7Qjpwtldk8vrTOIGJxi6KSo8WTOelDxxHivMn0YA
MhXDeLgB5Bi8FRHJX2CfM26rd+tEgK2vtAW//b8NvyxCgp29RUrpcLOGMLlrzH7BLBFqGlzvdY3V
nEEfwFo4UVMLbDCN9OMPoRc8ak20XVpyiUOZ1U8tWWOxTiiORF92vSV713x/ftJGuJNDUPx50ASm
llKRHe0//Rd4RSLEl7n7BpthENA3Oz6SvpJdeXuuxm+XjTWASUEOk95oi72UAvfix6R/hEyZ8JK7
UBcCUoWQe9f3pLo1PF2sby8XM74Of/jJ6tLEaP2i7/XQ5b4OF8T/xuJv0XPah0/CSVL5u13BBdD9
AdER4l6HOBAEWBex946bgcNDsHm8/P9n8lVqqqeXE3bLv5wxr64hJNYfnU7a1bon3rFtaoEQWoJ8
b7cInEdrdJn9MGse2/1HByWB8EaYCfOcEwYNoxi72v0l8fhWlm0GJi3yjRQK68UHHmzH+i/DOPgM
qjg6r3rDBHoY+BwiWDLSLvkkIdy2jD7kRxJN23gpUsN80pmQnXpm6n05/1uhU3Vy4K6fFcUezYvw
UR/zwUj0AIhqp0BXAKMmbq2gBzu21ExZSHjQdZIfSMLIs/jDAfNPVY0C+A5EqNrpLWQ5umR1H5h6
eOeNe/+CvhQCn4zfqiIuStkE1QvR3/d4ZGyPh+YbCCZWbfmFxbo06z0d4UZqKOTJuqe/kQMKe+RT
PNgjPEP4kuFrm1mYvN9Mkvryn7yXt97bReIjD9KAFKjTgezeP8UZhQ4q4DqghE8ZFGzFZpUUFN31
IUAOKQ93mCMNaZBuxQM0Sktb42rNdWbiYDNjppcyxYAZsAdeEpyqSD9BczxCEFssQk+uXCdtuowI
DxcVGTv1RmJNqhcwo9M6pDDuTGGCnNoaq4BS7V8lMgycWh7MR9TIWNarAohsSSWQ6vD7S2IGbD/l
7XHKg+Uv6xy2Ulmx2uOUpsYvOINzu84+v4CYvPBsCmpJJ/8LPoa79MP1VqSG2tbNQicGVRCMqSDv
sQbupYSf1NYHKEDDwBAnVBcUsviQ2okLsEKumzwE9buvfGWJ8/KJIrrHMsECFle37Hh/te9sBDBf
GFTWNT/PfMienUXNy1ahREkQUx4rtZDkS6KjTuLIw7W7Zz737YXhHRNYIk5kL/AgfJ/JfWjWmssa
6cls3oVgP3RZxFHx6TpIQgIW9gPxWRc6a42BR37xm203tfORdN1PCNmj/HUDP7Ob9g/VZRrfE4o4
ODBNsaSgaUcegPRhpiN2hyJNOmfGktoKtDw7BoiCjxUflhPbApHD2vmC2hYRSQ1FzySuNV1ooViJ
7kXXzJxSjNzqYWjZB1S1+HWT2FlRfNyJN3niUezX6jcIK+d9on+FPo/njLyz1Q+VPWwdwGrzMmxj
rKsH+fH0dCsI8u8fG1BEuky///A+FChXtE9tThT5BKklaOqe6JnF4OPXipPS3c42Hbv48MCu52M0
Cq+tUChdc0UsqqQBMeS+GMkj1t1+tl/2SVzFvsG5Xiz0FdeTlvxSH4CTPUKf2CUvPjPjQgXsnNhF
1oiEvUhurhQtFhzOECjM60qZwHPmojfVgdBP8wm4xtRYIphb8e4VHNCL6FXTsZagrfQ7305u97JB
rAimEa/+2stW69ozRkB9ecvQs+Jo8fra0/AXt15QiTE09bG1BG0Fy/OmsAXJRGUc6LV9mWnBXUiS
tG2n6Go7S6KBaZA3ku9DEhlRwYWdMfG2zqPZDsM6AWdvjun/4myLcv/Xy/9iUtS9WrP7aKcMocR/
xA4WEuMIOPbensph+x6HHh6kbFWWEGOmITk9R3iMNPWv6e3+wcXiCrEGpUhUiJFsZXeIcPEWvXKm
fCY6WdmXkmZAShOUBqcxGGBoXGdlsCtIOfuFat9ZGYLO1djkTRyLHrgqzXndHZd7k3bFtu7nhVX4
++mdmddVoFvIH+qAUDIvy+oz39uDiKIlOyO3s6Lv4q2V163ijvTHDHAyzdZtW1yaCozwczZZIvTn
vc70H0Der9Ieq7J0SdUQZ0F7ZquFP1c+6YRU/jvpvHFg1LA8g9wGKg6TDfn7eVGEqyOgnVAbd6To
zK4+FzEN5ZoVUaK/LWule9NgwMHosWMcTkJ0Z42hdRJozZOHQhGCDqbiXS2vnBRjMJJnjL6hczW8
s0qR9plytmi29NCJ+GDqnboWLRqfuoUYxxU5RpzzycznmM63sbreJG6gzPVjqjWDDNJq5YKicpum
LPF0S2MD4vI19WcvH8VuASPcoCJdrhUjS4/POi01U7ZNnt4ZnkasEcwpYtMjUKnC1dZLCmRyTA8G
qF1kytrwsvrKaCshOsBnnmzMST5OVX8eE/7TV+iGvNIlAydCdR6+07ys7k2oO2dJBaKAnUtQIQRm
oeOfQYh8OA5lhu3P1orZi6gAwYfcrE0FFnScZ566RRMmm4HAeWKDSH+smCz8gmP0+fU/2WhdqzSP
hs7ewIdilNEKaozPgm/H+39gC2vQTeHbjemKXcue6VwoIDhr+X09DLqSZya1G2Yj/pOouxcr+nhy
2hMPvHv+9fAvgzIZr6Y1qOU+mj6dE8v563WJWmFsLwfH1UIb/MWxeN3koGrWqeORPtczNVyPQsth
8Oq5257f1mj4J5Mjr8zTL3EJ+BRxTSgq4/vArg0D4rh6forg/dAKggP5Gk5qWDGj1vIerJ12A3KD
KINOFvqEtXBoBxXJaIpkfO6px0Qa9YLelcO7ScpUBpTHO5ht77ek3BC3zrHrFwcuVOmde840tUby
K0ttwvg2pLOxk0tW8Jee8LZ+9pG4k0Yrg9TmvFZN1GLdsCAgLOe3qlH/7PUo1H452fuFBE20L+tq
cewQJ/Npt9QgS/GrR/+iGpmIz57amflyalPLjpBm2DyiU8YJB08yriPSsG+F5/3RYl+7JRZ/EJV8
Aum8azNweu9T9awIclCMSnvsTPjqkHxLisllC6MbsRbUBCj7lv5nWBtqmcRtZh6WUqRXO8T8TdRT
pD4ZMF+4xI+hTw755K28tGfmq+UsE/ILhLiL+PO0oBHE9myUH8NrU+wxIhT2s0bjZlpbZRaRv0dV
CfP69g9XZsYwne8OGUu/Yfyp++4/N2YQHCpdTPUFwO4aekI7Yp36EUkvaUJXqne3oJ+gcrdm9t0s
rqxGqGiVgGelNlvyvvEUO3PAW9DUYTTpoYtm23ncCkC03UoK5EnyCuuRIxa10txSwLVr5Jialbrc
ILZargVRlmcctQsM11W3pZh8ybVIEHYa26gMoZYni2P066hdBFQGkFYGYqVqVxT5xWeFcppWRq4D
TjsNsL80yw27uzToqGxxmjqxTg818CBN7pNp8KDha36hXh5pZIR31RCqFbM8dubWeryh8s3SwYTV
U7LLz/pa1TFlvHobHfECSqxWAKLkcBRVGCrya2P4pAhPBHnTV1qJJ3hs/bQffMfbsOsuEO8FeaxQ
IKa2lkGMFRDtXH1MPV3y3eokqUw7M/y+Imb7M4kMft2oxiyXlRhh0zqo4PaWAGKIqj1+BMrsXEWx
kZEHSQk7q0nSpvj++iczNW+SOuq9/nedG0KJetnH1//GX0Q0ynhuL2kJWp/1XCV8pVyM7I66djB7
IQYOMN1BR4bv1CNQWVro0giACCmxjQ5Ffm/+MAPub+aqp+9WraNXCO9l6J/rcJ/Tw0TbEqSdxuJv
/fE2lTraB7zni2MRONq6/1RFNI/iYF1dd8X++kOOO6CiBT7tAfWMdxLR1n6hoOrLoxMcBjwSQxxQ
25tL49k3Ik0oeKcJeVgnfyB8XMJwd5LpFk3iT7ILMiMNO7NdhMcz8VHrBrwbGL+StoFBOQRb1A1G
owNiYeaS00h4HB8LGIiypYRcZUmSlx36wR/Khn6JAbcoG7EFdumVVRJkviGnl7F6oRJxVmW82OLF
SkiiCCbISNwueNBYXsqcSYaKuewx6hCDFcqepxtNcogQoziRp4W6PLeIsw0T6/JS99O5sCXdvZzy
8jJJuQov/dq8+KEsjn5zLpOisA3awiB7mdaSMJJXFszGVPvt653vDB8+eiK6Laxm9npZ85R2LVcT
oyYK3X5H4KhkP34OQZPd16u5dgJkTErPF4H5eUNo/wYkzfC8pZ2QdHin8emvbdpZz1MeS+h6XmBb
kc7CzPztLOkska7yUZ1X6EM4T0JI9T11FXmQcg0ipW7r3ffh7cAuXSBYQk5fbfQwabzodO5kKXju
WT43f77dZibR+uqPswUTo01+TGCEjDyi/iU5O73fjiWqr5nyQYDLH91+jlBH1/IqXThP91LAlbUg
2sKQrQwJMYSMsybS/lppFWSw6l6quKK9NwhC0H9mvYU9sH5oOx7RcHXy/aVtREFS96UEoWyBxmiq
B3Rk1moiE5FGGmjHw+2QZprVewPrpzRkTcxKcsqeSknJ/b0JH3fWNJ2x2WP7bBxkCofS7ywd2r5a
eFzSiJuMJo4C8W/Cc7zW/8L/fQ51V/cLBcdkyKorvmhQEEuGKk2htsIIaSkc1hniE2y6mLyvqopZ
24kFHyWGVktguHdSA4xXW04244mW9q+EiOddjub7VMlh+muUGaEnfBRkc32sJILYUNMZ0oLlc5VX
YDHTcRjb8aigubeNnqAxeAnb83kwwH8WvR9d8D/Fw/7YuC8Iz4whguWaDA2WnFpjtKlv8zQ27yJs
BU1dHmC+l9g4FE8ui7vsFbWX1zbJHc2Y0v9zAv3peLEy84dIVzhXOrUDOnvJBh9qrwGnFER6LMaZ
H2yUPO5JjyUa5jiDAbIIdy7LlRBsdV//jeIh5EMTkzABflPMdom61C4uks44RDOTk9Qi7bd6oWpG
lxETVjD/sd2IIk7hvskSmvfgCYuwmRZ9xaHYVuXLB7k7o+S/cA/c6gv4697d6x1hTjArRYzmBNBP
phVjSAGP+nlX0eabu8w0dm3wRdOkUFciNQj9o2U1mS2+NdhOouByc58htpaWjq+z1/g2vcWMB/im
A5w9PqcYtX7lmffSvdtzDDRp9O79Po8nstdmWxK62Iu8rNS7OR7mpDH8kenNW1TqVF+MQud3fDZF
PSCCKoWHygSQ1H/BHAWt5amPnfvo845CQ90VCVu7+oS+Y3nlsx2fNusCMNqgSAB2xwhpe3BRN9Kr
FaE1T6NKTMn8oziQpQRFHf+v7Rl9OMng6D5q6lBbBEAYl47D7721T6Do+ObYCmZX4IIuJekCAT9m
r23AaHfkv6bID54TSwWTF/yrNiClM2ZaajP7mMdafFBmoI64Ht8BUvNtii1EoA3+YUTbpoo6/dMs
WHDHzI1hCUEEuF5/RXHl32exIFtu58f2Cxnm0WePC2b36RJ+g5+t6SFq/fJ5mLjsEt8vpAA4Hvpn
FbllWlLCl+fzJSEbK7I/skFQR0CL70w2G3g15L7QUfPwhSy0AtSWrc3tRMr18pt8eIna2cWqSPzu
DUumNpdj9EOfoxtmsGOQ6McO96vUv4FTnzTbnAAI0U6fWqg//QUUoCR+8T5RmYsccgj7cZgCVLOS
vrf6oezo0iu68iHDksr5H7Piri3mBBKRxKbLAIU7TIgqekn0OcE0ArhWtE8Yk0GAUDYckqH81wkO
5fjJkUD7EHNYwBYwiZsb5Zq4cqJdqYx3i799EF2zfWgBE1gBfBAV4CIkplk99Fs2P4QNq2GvdLXJ
WZoP/Tl88R1ibW50K4LAFLGsn47vwHuTg7AT8WxGh4YovsyQSZJs9UReD9wStxaNy0+prfhhR366
Pb9qa1abBaWrMvV24v/r+Z9AjLFx50jj4Obl0x8Goh4eQyCa1vojyqtuTMOPynCd5q4/xMBA38VQ
HSPrHHZd4328KtgU48ec+mw3uYYqCv0MU9nNoF/AMvKxCXqOcRquHtQmw6WX5r4sDyW/fZKGpqd+
XJqS3zPXh1i9iB7tWOmgWmc8e3+oLbBO/wbQ8HQ7yrjD4wIovSYbhG2rKOxTjMMpJT3H2vOvvHSh
9njeotohsTEaAdDwGY40fk8SBWWLHXbL5MUkyDtnOEFvSA5cOqy2TIgFaVF9zVA6L7OxvEZkwdZI
aMSy/Sqr/CC/4syQwDfM511p7h1aMEvXqM2X2Vdfpg5SVMKL5b2Pmgi29UioDI4Rh404rccxkh3x
OC6pnvTqB6ITyat8c80as+UdBRj3brzxoVBH6H0BH9NEeNGtmKfkA/yx5EIo8Th5k77dPQthuKz0
7YDZwFMO1Q3E1oI+gr7E1IMqjEz02KjPtm9xleG676vGDfd5o5UVca3n1SAMUHrFuQO3vwi6B+7q
S38gz4chKBvUE6PiCCnOLbBFvWqQY8E5mys7fk3VUkIadoFWhfwmDVl5HEe4v2JuBKBl9WkRUMm2
I7BZ6avCXHSHmpOZOCRQcB33MjmaCWpSyu9naZ8frAJw9HB6EZjrVPlWj+D6ZFyEOkGSEq72lJVi
qRuJHdrn5q1MIRRAfANR/Qv2OBYGbqeP/3ZLY4WESXuajecE8wy6YN5dA3ZusIywAoEfoYZ+P8bO
tMoHjm+15LV9F2kppx9/eghNzyrMMxwA+b4DHDHMAVq72HlVMu+jwDv1HDZdUyGBT9k2x9EYfoG8
O/XBEOP9zAruyHHFQKPRKpFrhF59ZHv1YoYAEkbK6tBeRH5jdQVq7L6L5zvjV+r6CBqD7MBRrjbD
4maTFB1YzmFuXN/miKUndVQ1lTDk8gW+n+Zyd99YMgfY6tpmRiiZyigYlPA3CTVFx3LitSqnoT13
XWN97LAv2l+gdEYgN6rTjst0tEK8pzB2E5a5cxl2L69D418z8hFWP7uEVbRC/pyesgSCIOsiAu/d
rjOUl69Z5zFRbMu28VqM+elUWtwBendf2klTA6uT3KG+43H62QThNFnLk/i4LE4ylI3Vzie3gXGa
tgv9F0BhNFhkFRKlcPV/1NQGKAInBHSkaSw0OpTt539i5GVV5Z4peBg3rg7A3Ilocbn1K7CirQoI
9uTGhVFBlGTnxuIYRY/dJiyQxtwy3wTVCEuMSuz0txKKw5Jk20yuPWVGBiSe8ARnFssv1AEOHRdA
qALaRHpKHWWZ4Tggzw6s7miELHhxJg/LlkB4lTR8HM0TuUXK6sNkzPlrifghT9HeMiSO7boI/nyE
rgGsbMlnD077aHfYVV5L1nUEpqtiGUA4qDdIlZMvFnF8rzsZlkeG3rD0zw+6+oUPgn95yjVjyE4W
ur1ipOTPg/ckIvo+ARc4RZdQAE21hueszTc4DZRsU0qZKQWyl+UW0L/nY8CqVVEIoIeiwfTBPEdj
XmrJWYPZRIfVnzB349GmObxnoIDmxEfdLZRY5VR+LdbcV7Q49bLXkD1KXZVUBcrvv60t4WAgPTAZ
uPqC30AkMAVALcN1B61JIlT4kCgcTkaYkN/8U6uOKAmRV6TqP8SQIDLrFd54xrmh2Ro6vl4VS0lj
6S8FYkmqn8w8mrP52kL0fRsbp8+owkvaNQl/bS8RtYDdFDd04N7YW0ISS5/aYJb5vvH93KTwdICY
hvQ20ojyXWPHCcyGZK2euRKt++MMDp4U1jf/kFbG1UsA9qUyK7b+dcDFD8WtE+jITDH2qROqxnyv
D7Z0y5q8IBv7GsLnrQOiPmtx7WWcl5kRhuJ8r1VSXwKbrtg4kmwJLAV05TQRwcm2AntX5fbDyd4V
/Fo9mZh3VA769XZtaucqwIoHjO3wog6XwTJSgd4xVEET2RC6kV9/BLWxbY8AWSJ2BUBfp3AVNefx
AT4ySL88Vkfs8G0p6dys2ZMymgAtkNrNihXRCYvlj5B8R67xJsphUSxH1zFmwyzuGkmVc/du81Wu
AlGybsHNwxBlIAeG44nb7x1cdo0cQzNfGXng9RFWdH6aNGlKER19hYbKV/kGzwvuWIcr590jcQ3Q
Qqq3P8miKX1cPWjfG4aHHONTbIo9uhfdeNshfpd5vydYuYO5ZP0kw2h8WzNMVWC+sY+CMZh2PQMm
j0iu5/U/rcIZodJPHrCDGlh9NhQTdKv/GyS+ykg11JiHtg1Fv/EtDWQKzfy22DFqiuA0uklV1RfR
fNzKkh6EClm+T1aAJjYlPCwkEE5dcUT4DCOrYEWUTuAKchyf89JOgDZZhGgIuQholsjrH8W6T7LC
XlRneER8HBq2NdvNo0Gcn0YlCdaQcGW7JBJcMj63EFsZ+N5+92Ege0O2yrnnIwDsZZ+2+mzhHZKM
lM2jx3ijbxTnGu9ufytW4uxeIB4c7afpGrJzpVqhiGwmy1nRIDzuD0Wqd+Lb45/Ph1+pdJMX66GR
lBlaCoQC8AMLjgX4E4++I9HD3VJ1xyQOkqJpHj4LOBJ6IWw1Hqk2tEOTKFj5zY8WDPHVK2fZ/mB/
ay+n4ZfM+/I1hFhKdHDSrRZVdFHbTitBW2gCjxBmGL74F4Q9CE7BXl80x5HSt7EZWkqI1g1PCict
G+1fuCKmayQJlBUPQmPnJjk83WMErMR+PzqJBEEetfxm8crvZOgpl5T8IUc/rkc7lK3WEnbDkZLY
O0jf51TsAhqu6fz1INz4oBilA5clhnGCoMAgQDWqct1eej+uqXHHirT/xA07KlxLnJH75gTkHR+Z
qWK0FdtPk4D8B4uXy/bQ9Wdc0FzSvo0MaAkj5u0W5L9kFfQof4LawmyIeennllvx/6VvcgT84mD1
KejU3tC57sWgYU9jbIK0RVzy9eim8WIMyiHIDwHCVLvGzNLWkUDrYgCDdGibKhESwjgDJc7aRd1H
vn/Cto9qKLkc6Wa1BHHZYHJ7KoIUBl1M2f/bwdOsTi7Gv19Sq+6uk/7qPbTAdEGI/02u7DJ423hp
H6mcgQtm4bgZltZVTGOCsI+XhNoIpA556BWq0BN2M8Vkm82m2oGUvQOVDJ8bVhfOAa0nE8mMvjL8
QHHWUsEfuYhvIigyCLEpsVMOBY4rzMoa8Qx0gpWumBZ35iHVxbQJACfRPMJlbGn+izzXp0iCJFIj
HOJ6Z3btceIkZjS6BiYjaj+hHDFlO9Asf1rqsUvtnt4Musoa5a3bemMCaAV4efArTv20Ek9M9zwT
jNagoZklJO+LKu8M6NVSLvi2r/CFv9mUHwvOWztyWnJMyq4EgVCpz4Jcupi7567qcN4Q2nhk8q/c
fflvXosvbunuHG/DeBgB4kcaL62KV8JpbD/WZ9JVHfSoZzHsCJXHjKvjpSYr9L5uDOM7biyCU8rF
rwKrDAlqy8CBPX2Q0WuB/uvUIhQnC81G9LLiFpmEkPkE+xkfyzzt1ILP0+gtPxJsGSSIMUlhlR6k
iwL60/KLbviM8oHYDPDbEqkKzFyAPxSqTDyghxKUh26RcvPOblBb0nz4w5TVTyh2mpOUkFWASRUF
roSJC0g4O8zWQOj4rvRnBaDdYEGJdyA5BR7HKeyxWUIgeelAhrc7mgKwLoLLoj3oByCBpo6kNN6Y
FzczpIfFQuBwKEafKCX3pRbWABzsWEy6xStRfkmlpZUNI11ucDFdLjuOH8V87G3LBjfcrT2QKPL8
q3QKS8J2AAiZwlcWsMnZGDuWH3nSPl0BfZEcQ1bmgahGe194BZ1MtPJrzgObr4fxWKUxan2iP3W0
Eqp6LKHrGZpkNwQy/mM/roBFB9PO1iOTqVVy+4/9Zz8s5Pw/VYwoh0zH3jHOXLbiw3xav28718rd
gXsYJlkBk8OWfinb+T6yU2n0gPju+29uXHnzOuURpw6ZD1TH/ndX3JCmYBK2DaHdwZzSPy4+586w
nED5hBEMB9oNa7aeWTUJi+NeYCCuajFSK8UcIxU5m8Zm4KjMC4HdUBoV/aTF4S4hLPS6F/xsLT+N
ZFZzZTz3zkR6UbFEFoJe84JZyFZPaFc7UztCKV9OF95TBkU9BEM7yHtBHDp6bKnUqyz4COMV8epA
uP90nN0KloWUlQ6v6GykQFNaDxFhds8wy5boZr/prB1s063xd0OCY3GGIwRzWH6lYPII+sNnL31g
QHcJazdCmbxvBc9GZANUiEFWfErIJFvnU2V28f4Sok8LVkA/+GQKF9tnpaZcs+0+ADnkTcEFWhmZ
Cj197Zal/kq4fcnnL9PMYc/nh5mMuOpF8WIf9+Nwhl9tM0fwwj1XbsvFt1GfFialLWAk7aMZsNJL
0T3syvuiN4PPgz22aOwJMo41DOd6o9qugfiaO0IE/thCdWGimQSsHeLkQqgi4m8dNJG7qTjtvEic
Gn6GbTg58C6yNicFFhuzE1nDjYQRupShAbZMcNf1EEce5Ol9PMq+Bccesz5ynl8PV/UXjINn1Uz6
zJGxdgrXiUm27rsmfH3ovPDsj7CrHwsGIP+/RN29gtiGdXMrebPov8qjW3okRhIe72bZ6GTzT/1a
2BM1YUPx3Iyqy3KU7ThuKe6fSeuoEtKzPioIhLe/O6UdbPVh4hBLjibqg+hEYVlOeOcCstnMFI4D
E/Y+tWa93QSSld58PnpNhIvnITyTg5GFi84A48LiY4+G0HgrIu/YZpiXCujBUVzAEWNPqGSl8cRQ
k626nCwRvAkN+2UjgvGhwJbDOkyo0N6E0e9ObD/iN6ThB8HB/+rIl9Ukg+ydFoe8fTb7r/gy+9Su
G2sdGwsYwHduTnwR3uTapf5SKffAF0wxLeAOIdOACpx6xvBW3kizGdjzSwpKneUcTtaReKML24bl
uMXEM0hofHpTF5lba5iR4WJvgTdMbaGyREkkgJZXmBxdOGPv4dTTCAlb/75ZuKHZYpo/CqEmvgb5
sSTO2M+30WvxuBEEZftimNwnM+aLrL5fJqDqB1OZZKHZ4lNRfkcNon2/j6BZN7WgmEhGlv1GywN+
1ry5qILA9vsgUctAS8tpsjDIKQjsb9WUGAnaI4wHbEvo+bBoM1oDOp/j/HTNtHYGz2X8r0ilJwLg
xxmBK1jjGqk2fppG5MZFKSZC6nN8qJfKjVVhvj2BtijkZ2XoUxVD11MiPzPsFxSf4fX33mF12u9v
wbmsuKnrfebwX/qkbzz4ulZa6TEMI6xC8LilNpkGpTHgPuKaIUUAft67WUNBiPYiIg5hHVBITCJX
wp8+zGPyUidno1Zc9RZ/+nFZV7YlqdgP3q3FF1nCTTEPcTXqUV67+qACpXGBa+p8jW5C8vcf23HT
U8yD2b8faomYVif5KFDS9PoZYR2Ht+gOmaDuuimy0Y8rL40OJF4nNqXnS7PKRCm6dfRUpCMC/kmv
h/bv12nccMlhBo1XHENqWVR4LTWy6Hkk9+f1MR8vjU/NOngLEq1+lsTNeakynIg9Hw97dRuu96SR
H5MkTHpQO6AEhBbdJZYflPsf8wvHH5yxy2VlXDVSvLL0zBBFcNkH5D4LD9m6t82z0MEsJN54zfrn
gduVtEpEhnTHUrQf8nSbDkr8TS1O8cs3RPGtuxFpn0X77rCdCnLlgOKlkNMpNsepQCzOY+B1wWwp
krn/tbf0iOeupCOAOURnYgd2/Yd9Nqg0vvbZUtIjxUasxe3dO1OBmb1EyjetvEVRLjYG2SRQ7iqH
95W1xTBlMv5CCSWjFbZHhwNEotHqG1U+9pWY2rnzzm+vBYOF/FOoTKnALmyJ5rcLmNf832Ig4d8H
o1QXbHSF8bKAyyWANuD3vnltU/Gbado8lNRn+odK6MRn92qIJm/Q4JowWvSVLbcVO8ArvCNxHhf8
YZRNpdPKu9NgHlt9aC19L6qhmiVfHPCwFuvk0Bjpp90JhD5BvPJt41w0Basi9SrwENfC+ATU9Dw7
ngXcNCgYX41Oif28QL6aMw+J3QxLYmxqI4tQEfZdPovZAQPxckWSOOZNXXyGSkEBhkiLRO6w8WoH
0LZ4iU8vtR5Yd5HnqOU2CpEHGV1AgBuUzXAnh+xvDssVKCJxpDDNt4bEMqvNwdvZUhmqvlTIq3Vl
ByKUWh/AUp1RPu0hQZoEc5pnNCvthdTSuio+dhOJppjka7JfBHTUlvIqZ86EHPSfKLFtIlJIuirp
+kATNqSiOv6R6X+tcGF06mR6MsMCwFSi4Ct6jk6vKXcjwJXm/h7iWibVlGKfIUxBXTgroS8G6diN
GXH35tciRMcKBYypXky6rmK/UL2jwkCAOvCk8YbPlu5YWc8SYEJiyE6AcGY/1kZVtXIlLC/o9z8J
e796uL8t84geySQeD/Vt79I6kNYG4HLtqt9FF/+lylZHX76POrPnffQXVlMrsAm1mLBmaR2k9rLU
Vl2kMO448ofaluhwepkcGomaKTNqwWZhJA5DhIdhkBBHQecEa06UIt4F1VMstJ/xxLJW7MNop+94
RrAQLmtqCOkPPvFmRVK2V00U9KTe7e9BMScQcQzxtwFwK7M/zGj1AqYlyKZIjLtU9KVPCKHuyAoJ
mD9xjiqrnRtlvsS3C2gxOcs8r2YICDJjHf1mFZXn+xXa9W7Ik+PecS8Jm9cioHjkzB4uCKLr88r3
kQ1XChdTtnwySTBYEmrLaURlI5qhtgwJLBAgy4atSQSsfzxB/f2NeMVaFZ4xZ6+Ve6mT4wZ7gD0D
C6Y4EnhHZ1BIivaHZnkZzqTwJWVDF1U78wmTiCQ5361R0SXuRRF3WKZBv8V6XxQQ4OgksTc5f/TF
qvSqxDnkyRGpACU0kPmpbw6F/w/4/kWBQ9tpPp0dXHAMAiPFvQxchaMuGyXdlw841hxQZK5r4G0d
ytosslHWmjlbSjSR6teXmaYhJALnKLLxBcfMeZiaTlW2HRuxrLmsb347jmarkY3BmKDOwXs9NkLO
hSO2IAF8VjpEEmWPK8ILQNnSEdLGz5b+yc4Be1bnZxT/bvIktVwjvCabguVa0Ol87LCV27LHbmug
YpMZUM53N0nrDPe3yvS0cSjX5amf7w83tUlR6RXvU8IbBhzz36HKkHvU8vCIq+ZWJXbe1katTehQ
CpziQrwP8u7tJ2prHmb+/B/1wnO/H4m8/xb4vg71G7FXONgchpd+W5dA+A7rtoAJoatJpbTJ9i16
Zy6xi5HO4F+Q5aEF4yJqRvza+GDHrTRrDl5ConWoJem43O/eOeHa7c0fRIiHWysftms6zJ5+nUX7
m/N+vLPaj/e1yzuoe7t+Eq4UIGUsrnRPuBWdMJ7+of0a9j8/JdmUw5tHGG+kyUOELbYpgxYIT+Oz
MS2C4H2PcJAvEDlAIBkhf3UGNUDAmEF6F21ixdujZbwAvls/lU1JnqTWMMBQRK8fhV22JHnpAaSq
+kN1OhUQEIR/N+80GTrLtKYaT59uP7dedwk1sAxJhYP1CEE9V4TD5AJcWq7agQcyKFZwUarEs3ks
J69m+wjcPsKG5vmCIHfXgG1ImsgJ28SgDUs787sJC2XDt2/ytqyNTfNeK5w9Xv/ullXIUARYesJQ
xmZZxL22y6kJEhBQpWCpyi971J1H4fEd3oXp47I4vPyGewpIeBULQDlz++zVnfcu2tP3FUaB4o9V
JByXwI85nGbcJLLq0VX+4ctHpxOiMTeZ+fXYPbS1ocqVWH5SxtP9w8nJHiVjiBwNUnOdXv+VZfyu
3uDXABT6yZRop/TbOWcg2iWYOE7/YtlBqqxopKjiTg8p7fqz7P5EELFnjuzbS1anjHu0bo/DG5Zw
L84lRX/KQKj1CkqaJSjRWH/l9nd2nhkwU7/BbDFiPW9bmbWGyXx7HLMFLQiEPL9eRyKPSkQqlUkd
VdAAoXvUgJd/jY9GmqePAqtkuwN7qH+M1TMw5+u4z7Jq8Uow5klmjYC+O30YL/ZKApRS8aD3Vc6u
u11pWBwb0n69i+aFOdAtlvXtYj9m1jYU6rfWPXWvahV3zuUIAPjFjuVWpH75TC8DXwjOKzv3jDNu
n5UN2GTv+UXjfpZPRMgqOQAH5XwMMMD5IenKzuAOdZcU2BkcjMrLRl2KxbBauSRd70BRpkwdbU7B
MxNIXgfXF2Alkf/9td0GMHTiYzQ77A6592KDn5xNnDC0bJW5T4ZnhgFLxwVb7XBVUSe2jGZgXePJ
5hcjN585iLjDwHI9iZYCPD9AM8xJyLtnCc2Ra/PCPQEohm1jJfn0V+CkjS4bhw+wDO183K08h1BR
RNhMfCvgu5VF+RI/LSaMHLcunOOm9s1zHT1uwEtROTCgWBuFITuCd610ArOEFRnFYOHIoHw7Kh59
7pPKwmVbhuu33ZlZa+kT22oyzF41JT27+dNITDRzfvZvK1LNfkHpL55lLE/GeQxAz0D9lQpy5Swf
a2h245TCd8e8ZCPutJ6Cles0gW3BGV1NqnHWks7lapZMT71fYbgjxdpeJuLxyUQxc5auaUWrYIQb
ANCppfH7MehC1NxximEgcWB+aSxhamkCYlqURMWort9Ap++mffs/s9zsn8jUBHh+ByXThwPgwZVj
BJMKQHXsEKSn39bV/H5mIoWoXGRjmZkseYVK0A0s7jn1eDXddbUksfdD2p+88jEWlQyXhVzhGYmu
jSAnJuB7wmISEAUJN8rvTJ9j7+4NvTSFXoQGrZw4SK2R7SNnUFnR7dxaI9Ct1vs23JbRHXpa8Omb
DJiaUnvZFZqIkCkaHdSiLEwSNiZX+YDKqZ19noPvpt9MVSJUcxu1gJ5vHJ6jRNU87eYxQ8ZgS0yt
EIi4MVCQ01hZ4ad/Y++PBGURYEuuFNexsh/+sY52fuiw1mwo33fmMTuoVjSnKQ2Apoq0emjf0znv
uOXXi/PZPWe0C4puKYdRLp0h9qE4WbEuJ+OCmqiFe0uV/qoRAHjNr3wnUjGCG0wb24YzM2wtLTOh
ERFlHb6Bejy+r2qLCwczGn3mBiupCMZJt/sHwzid/wGblubu4U0wCnI/CKTZ0+1yUnaNoV29aS10
Cq0ynJbQIWKxjXiFIppzQEiVMOa4IqsnqfyGovxca2OBQBmdVaOSQXH8fLthehLzXTnwKkh3P5wp
VEs5noKfm5I0IzcJagCW0AX6SEkbTRsRco2dtUfvxWORS4mvX8y3BYr75m6JYoOlbLYILWljUC2S
cevAS0FHtpqayT9qVK5ejbm3uhfN8+5svJaFq/a/Bs3iS209EVARz1zmDQS4WcDVl+tkJBAG+KbX
lfBhZJia2QcNIHYRQxpu5eQIAmQiC7vSUcF3TbcDKUIX4r8bZOtfYLjiBmmpYQvmZANelKF6Vv6p
be5aP5zKvVhrbORHgglgqZreZChnjsl4zK+Pr6VMxchyz7VUWXj/7PMq7CivbZg1GUAprIH/O1Te
m3ZnTNGS7g0z/8adcyK9crMuyqC0Tym+tMDA2TEnpuzsDZdy0/Ml1qigY1gIRmY63i1mUD3f1Q0P
R90sbvSKLxKZQkxBw7sCHrODEJneWYkm9+75q/z4GCYkt2UzuoWxIO2XwkkYCqZGltATIwCTaS5l
MpBe0zknoiFF/e9NhBMCxacTjKvYK2p+qr0hZ5v+0JxMS/ihf5obWkZ1ooy+FZSHKqMvKgC4Ul+M
YPSWP57VNFEgbcjYJhwhgAsNQTiDL5IFb0wwa+RPCuleJjgEaBv9tJabPGqF1HgVJXawaWuyUWPU
QalF0zyiC36yeJL7BWKJhSOes82+N2DSY5sEWkORGHpYOCjwJlKHgHckm8bONvwvWO+C9W1OkwBg
Ytq39scFF+rimbfx/IHbVpjwr2zKYMWVBlfvNCuZb0aFeYLgye9vuoIJcFrbAIAa8T0Bl1+cDOV1
CuOf6nOwGY+7qET84Ysd27+fpWh2Q1N57n2/TKjPsnoZ2GNGvpKUlgzxZLphLDjEB/ysM0qoVQ7F
eENn96WzSb9n5RTuipYrr782FUPSabhcTVNiO1+Q3kZ1qnPb4QLqyHtKoUd7VL3SRFFN5sqF1Izy
lzx4AgAeYdpbg4Ujf1l3nNJkIBjauVO7z8zGg5csWYecYim38dhCDN6Y6HlWlcr2bqSURjv1pZxw
/lQX8xa9crK+EAon8b5UP37j2vQcHuBeXa2Du2QnLurWj79Fb0kGIhhp+Vo59BFuNQBcYUGpnkQ2
rTHhfHKYT5olm0N1CSIMDLqJ69j/Wwk6Jx/JE3TQAPhCAealnH8Xy2AUic+B+tEOH/Bl0mIuJbp/
wmAzQTORsdwdxdvFAAyPS8n2umeGfxDoZvxhBL64u3lt8aiVtMKyMUr2GptgtD/Ou9RQPuZqKe6P
Fdq/624jaENB8t18OLXfm/QWn12VvsqIJXCCs6CU4bDgWZOUOOjgx7fmg61HVw6xRB8ep+1q7iX4
EPkBNM32Mo7QFsc+KxkGcwPdWHxuStMbjIC8WyQoBcil8OAU3BdrxxvE396rqE6b0BXQ4nfm+f4x
fOE+4ITHG/LyKhqJaEGRCN3GzX7yIVipL+NmXgQFbQ/ttcSjmzm0KPJtLTx5rYj9TfJJ5S/S5cwh
5YlIEyKZR7EXaB+FfaTR/g3cCnNGqdw6ie2xZYtefywJ6iIuM12Xx7isbNcwckgU+YY0rfVW0vFs
J5+j+rHvs/bAUoncTUGLlUv9ufvHgtNQLP1FbeyATCQjJiQC8/z+SLMxj+RnuCZhkYOqi953hmt9
l32izDWNDIyRGgYMxonTid9fpGZKCIgCnNni9Ejp9h69t9PTGlYckK7vmFrFv6+MoN0g4391/P+8
Qh/94gox/1dmOn1qxvE6veqz44MeyUF4tWQuBkqrlYIcxN9i005+sMMDT6J/2tK3IbuyUmYHg8Kn
kRsWyLk3mVQoHeLpWK/F/dl+mIYCC5oeS5fXVnktOh4CuEqbRtIscbJxDEFAeTr1XtiGBebkXh+z
f6qQxhEe4YxnWcjdfTA9sAaI3KWR7IrVRa0hZ13jkbKhek/65WeV9TeUldyIvLvNQMsBTUlAYDEC
SS4bZWbmGFr5jZ/F3MalQA2BwswTfB3CCQkH9U/ETVQSSbpmH6HYjNtAdlwzlaPFqCapUnc6TrRI
nMQo+WfNBMPqbYNuAwi7aQOXOiXPLHB5Q+srLdfRo6aRUWKLpyXuHIoQiJ3xznAk8hybkjSeNboN
G+j55TFWmyLeN5mupESs7AS0k90U9VsAHfWGpKRABeDLi4xL7wpq/nVcPAPuJ6aUKHGB1HSZX7cv
tzsheppAa9uOXzdFtYMhfLhgFUpAOeWkU/9F+PQJXxzYtrkBiJSYlKZ8s963GTYtv9zAcEyjeqhm
nR53004Sm85OOYDLiqZshF/loxBaX7dJ3BiNWhKp9BLXhoZbDkfMf9l17fAcWv+JGqN8QgH3+bmR
aMC/GeT1sgTQL7ILRd5ndKDApxRc5McxoM+cDKDVDArLhA2t0qySrS1GEYAyF31cMth2geInL68U
E7ViNUeLEo6Ai9MDTJgOmj61zNFX3N3LF54YtcCasQ2/APY/184rGaxt/WirQU4r6R5CXG9+5TwP
p8Vde+VP1+ELyT31NSTVBm7EFxM6DpPcI2uoue6rFJlrauv4UqySuNUeUmTTjAUFHbOCw7Q4RIwj
JRp7hcF8Ue4imbJUbbMwisDNzORBRB5OotuQK6QgsxaJbNcyW2VOjPtlEPdFX613h15BcOVqGIUs
sBW0UIu33j2vuMASb+teW0oOBaggNx++7Mx7sQjXftUk+jDgsCp9KkkfAO/y7YNLTBdUrgbXtlqp
t+PMmX0WqStRYBLF6sigCShxJvTikuzcYQKENZrRLG1q8n5kcVC+/34Wcak0nDp65E84E8ANp8/p
Lu0FumymqlbiNp9LmcVeVtIxn57wxiVD8P88GCtnFp9cr5/TjUAux/HTogYTtWYYtvgv4OVjze2q
mIe+eFB0s552D9WyXO9lJ+nXs9PV4Tuw8pb7Rd1L17ktlG2fbAcOJ89tZOYXaoLdZ3CofLp7qIli
MO/QF9Wj9KkG531GHOg+FYbnXpbpOEceGOt1Gt+utFLM3DZ7vbBfekux6QDffKHUCrqKhgnPKIDg
jmVGViEQfL/UoujcOigXCf6x2yYBPTptsRrtU/xVHH+NG8hBnG6DvU+KDcerc9AO4KKlOOMdndMr
DTOCwybWlasYx4F5BcwEA52cEsZ+xNM1YVMHDi70NbRXZrFc9WFekkhij/fuRxkoxhlKPXhuK83l
Xb1xBdBcaXmyqHWZRYzw/iln3i6ZilBPDDe6Pqs0muWgoCK7wZaAUJ6mA70oIjBCEtOn2K7qFC2Q
LXDYEO669TZfv6+UobFjvNhTSnZygyhNIoio3DsV+bb1QC4HUJgsGe483TxIBVTBltRowxe+hUpW
DDlufGfNxYAuSychWA67Dnz7H8ptBit+DaVVm933tKfeLyuqlcsTXxYSsU5JxHi0w3TuUNx1zieU
1A8/LN862llcZAbAi3iIQQxqz0kJU6BuJtyWOTllg1M0e72BUB3al6ZieE9X+oBbzaBzuFxbLUy6
ZBo3wWHGqHPaIXGwoVXfGR/OdO4WzXUV3SkRBB/in6Q5bebb1AeR8H7rr1wCOsEAzb7nvRDvxQjr
7cE/Z/KXYQE4p/esP0o00NfLtcMK+tka7fyYyrELTNVJwekmbFk2qqjRWOtxeHLJlgiF8U6W6Fdi
6n2ccfJaxR1wQVmOjmjehQPBQzfTCbCaq9fNFRHwLuVu/iP5qsFjWfxAu6dTQ4iOXjilNaOU10v2
VEOJV762LK/KO6zs73Muq5MglesLVwfIF8KZ9s0MlM8bFoLrZFVO4DP/NZ6aQXV3ezFm8PCLm06I
NEHvps4nZkps+M91sDmVx0PnDa0M+H3+aYqd22apTZQvka5dNj8mKR8Au41ihiAQFt8Wntsfm/Ha
U7baqdILiP+I5y09q7Yj3PArN8OquBCO8+naRcd/T5RNcv9JGH7aq+rQGsuxpHwcj8UbQzJBhpty
cHCYderM5puTatrVjQRj+V1MMNNnucK9dQnY4fo1QfKUGRgt/fOVTwgYYWKthqMpFDkUAfTM22vE
fSrZamt2TM7djOrmqqcHij6CC86t0gm9gT/iHEWNW0iEiw/3bROvWClsLaozhkBHoKBFKTngcA1S
xPt8PTXI0Zur7YUMOlVxtC1vb5v81/rJRI3ZDpwEEWRilr+eeQjzUjnJF85BmS5Nrn78uTrWOMWw
DToZc0+gPZmm7atGDUHBWDHpjAuSYgtP9L4AwbIVpC9Ovh9ObzUQmzqgmgWJauAkgLSMZfGsqmWt
lZe9q63lGaFsJphpifR5ySIPkUTGcdUekDitu4ZYVZQ7DILpyM6Nq7DqqB9FDH6soMyYArfIfrtu
1CHU9QQ5OStmjndH2hJwTYfpmJwRbyWSl21sp4vSUgLAgo4bQXxekObhKG3aS/N0B3My1LGoDAof
VHym9EThqKi6XJ8tG1R2CPhWekrpxCVsBS3AiQ0I57RJ75oeGkcdIxv9O7yU7w1gntzrn8+dzSYM
SJYchXdyZCD178bacVMWjlEYiuVptXHMek0ZuMs3LPtRNQ4uym/6DxUM2HO8QBJLS4nUVXemjCoJ
Aqgx9NcF+wn9madB1Hdsio/bEIyrjw882whnelTqNXh2xXLMSIBbjC2YgVcHEHjwG2WdwWuGLuqE
Qmu/56gc5+Dq5ioctkZbEu4xdLdbTAB9MgIe7RR4Sm8O3mV4S7AXXMuYfoUNWFt62UlbWC8SrXIb
LhcKeGbmEfkvmJH7TnCVTDWJlC8CVfUcjrBGnFps1tgIVCIvUx/xhEGACWOixSByGcnQCVR8qd2T
TPV4KZTwDvjZ3SWU6Tw2peABVMfZ8/goXOAECcp8xOV+J9IO5qqICDN/Ta/RbJbVv8snJ3lrPrtV
aWTVk04tVHgVGUtTeO9ElUU5WBFdBeB6t/w4NBXcNEQ/5BS8FOXIv8LUv0ES0o9eZXoEwVHtHbZg
N9Y+mqdIHisKWStDw551ZZKU193EiE5vW8WN1dZfWeerQIe+YVBhbRDoSsX8xy7mE5s3r7GXoCGI
QOD4cPz2ibAlKUHA7qR7oUwdaBEPDzUJO0AxT8mO3Y97hqOegfOGyZRtZhS5pjrCmmv6TqB2muGU
TpOvByGDfdnP4B+rMzSM1U8shuRIWSNpwNGXES97b6jgpFCWpaVZShYpsqCF/0HXwRi36ZEhXGwL
YvsdWofMCRh4BjJj56o/k0rKkiJXIwXnoRV/St0lVXbNh27l0e8AYGdE98WspuzvBxc3sKGJdU0E
XzZ6eJp3k6HKUh11wsooM01lHPQ1pFNYg672cCpTV3F8B6KjgeYs78dowB+k+7F/zs38uJUpTFLM
y1HbQiLbHO0yDlH4WPwC1QF9P639J/tFvcdr53Y8HheRZgYhQ6pejbjy560eT1n4mLJPcvHZwcyL
9Icjy0LV/Z4HeL/9fYp2Bdzf51daj1qNvPEBGlbfYf5z/E2BziPhslHaEqXerTtcjuXqKLiQojhO
u+t3UGMIBJCR4i3BBOokjIQsddsWTItkQY3vuLm8C//pVWvD80C269lXHy89UGsqtPTPT5oEXX9O
iOa66eK263DziJMtEWevtShgDOJpwCJec0VkMhyr8ZDg0DCfQAZAJ97VgMyXMXRZdctXkZvt1gqi
o4oITyPJaD0KMf/XUoNrwEoBU69dY5RPTifw6ZqFi8LY9SqhmVeNuhjZwuoo5MBJdhk8paq/T5p4
WINsT+aMO6LOr22UsTC2jGI/T5ZDRB90WTm9oWWM9F9yXbO2nsljywxAUctV5z6RGoDnpHKUeF1R
lD8b5QNOA9dOnOJGeL0DLbxQX7y3asmBqyFvVpJrduwfswX1iGF7XLlUZHYbv9aTiod2fjnXXHIn
3S/uBZXYJY9KHBjvQibU1HvSiGFXWFSlUB0g7IpQb4VeTc/G4qV7Sl65Qtt+Hb/yQatmFQ4JDX9J
30onufhHwpQ6nEITaasXCHFcP+UULDUx9JqNttvMHZi5Dxp+3CNI1007Q7qEYfRUAWyoX/D8spQZ
NR4IHvSclomprAUYnoaiL2ybBh35E8RsWXTLPmqMjNX9iDgaqsbd3EjM+dWTCAOMJkUZ6Gwn1t5F
5oh17zcsgn1efMh2HZaIgZK8wI12QUvcrQOzudhrziVFLeV/dSNKxDcAxF8gcE8ly1OJa2AohT8k
IYT+VmmQdhqG3MdhSucgU5fClQPLw8ENBisiSviiDVmfaat8MFgD+a2oK4imm7BQoMAhcXFINd3y
Y80tlrhdGSDUxkTt60UKjZuuGs09H1ydAXONkHznxkzEm8cuR6X52mZY5ktk4n0ov3yiAvf7Uc5x
u9TRE0SGd1l3Yv12+UhzbBS9zOg2JWNhgTWnWGA++sL4WfMc1KJSMO+2sF5652RDff5mJNmgdQft
FHB8RyW9MFcg4DGDgAg/kPb4gm0hJZzoBAW3nx4FYxiv3Zkq/eYTZ9ciwSmRSLecuZBN0OX7Mep6
0IEC1Kw7JBylo1q5bZCu89EMlWnmylg/Fj035n9SDh7p6kMqOyFOVKU48MJ6SL5ClbipDx3X6qH+
xyn1Y0AwByGwmBYd31hof8xZoSF8IDAgQVrmn3wh3nPpkyI6fwT96DaBdMhXOOYGfbHTpEKOnHHR
XUPC5LigA80VJLQeeYXGSg+yeJXEqZLs9vjPTgKcX5fHUR2SKiCM0AYIcc73U6wkKt2Bbnhoc1Pw
4dxCWR+9yD/akMaTxxEq2KNPJUb6Aci3ss13Tn+Bv0Co6fUuKI9cBdtCMedv/yZqTQ/upVpI74eX
XYQdbEXxzBO41dmoC7Jfw91jmJnvl9F5yX/Zo17T1kfDmBnWdvfYSvVjXuSw1ggQLuFMlYvjmXWR
pu1IwcLIcjUaAukwWgN+H+fxIXpCCb5G/hPkXK2QnKqy8+HKPkn1XA2XfXwRwp1ErrlO60kh1aOC
nPxz6SyYAVauBQVwDUQh8T8dXYYQgyswZD04IVewxW37sTOu5NREH1Mw18i2mErtHfbEYOC26cYz
W6ZLF1v64bmS95VzkWOJpqhOCRHPsJsql7Ir5lM0866clJ5Smxhvfe2HqiWMap6bYsy5gESH+TBD
7QlkFVSfjTVnoDeQVd8WawBVV9oyc/9XejkaBsowm+vufepuBZGP5TVjwoDXw28woBkMV4RsVzWl
dhIHIT/DyBhMCmr+CHqQt5Og/9zJqe20S/nzz03eEjPr48hFsg2sUiHuJEZxj8w+/knpBA6sZAxi
6K8FGOARMQGwP4Fob5qhl8WUfKi324nWojAuZ0HvgsGpeMpq+j4mO4KhRcL4TI9K1bIfNUyBnCSG
VrCYqGdsa2sAoIsbU0N1/QYn8P5iIf1O8ow2Qz+Q2dhAi+FIGfjhiYURg063FqPxIixAZVqMb4lF
8dudHQJ5SJShqaQU8lkt6gmNyAatqXUAPwNjHy0/fmdXNphBkB8jFOUfDZxA1v3ekP/72Lsm2pZC
iLo0QiGp2y6k2/quaxLGyTqPjvxjavZzL7Wt+xTnbL5MjxNIeBTFCsjd4KePtrNsYe5HoIBt/5e/
+BWpp/ybMQIqwxG8LY9d7dMkMfNGOJx0cw+rwsYMxIt/wyijCUnYDzOKd2FwFFX47Kk8/kQBaEKe
e9zOPrh+OC+eiVvpT9CBvqU/0gA5eL8Jm4sHOTqQtzz5+Z/PizoKp/6qILuJ9GPOwUD24TATS/z6
QnfZoddxFD54q/At2WOkEy3wAYelSRbBHYJohxHn9uirO/8t0kRhDpXqJhxNQXwku1dNuePVDPf+
LXHVjPm8ubG2OP2SaBKBTePfOhphBwvBGIP7eQhltHp/QeL2u8JLiGRnqdmOzUgl/YkQpI+e0Y2K
OXRNbMvlUtun/ltJ8mqUcqNFsBmdD0xY1/wE6+JsG8cXrgpuxbnrFjlPqH+9Wrn+RmwxAHd69QEC
UOVunS3qAEl8QfMm9u+41N+XZCUz0dBlYmBtPTM9u5bsqNy6JUoClXr8k446rAKVdkm9ly7VXZOg
CK5S9tT9ImsrClfrR2rJBJv/0OYjDk6UZpr8VMxffIjMJXupRbRLLc7Fk888E75uiJQ+U0P/ot1K
caciVy2ZZG/G/zluhmhES1woiNbRvLquSan21+GlzafR6goP37pUeXgKhSoMKntJtJU8zoC7yVu5
SP2U4CcB/Z6toiWMz1/nLzs/aJYAmnPEAmpokYHcRkKNcrzRn73+7OD/3WBVa4ZD2ncpY7k5xFF+
9Til5iWkdklMrbqBPW1Up6jRNEzqXAQQdMeUOVb/Is8o2laljOzVzTxK893SP9Z1s9878xALXTId
0hp+z+VvbUDpAKnBAB04MTaxJrKfYzEBKhXobYER6y32aPPCTdqtDQxMfC1/vI2g2U7opHSNtEK5
HvhfP8sk6IlG13jwIL9/219LsBE5THvtI3Fe7JVXHBWv1csB0QuURfTR8n4RcAp8NiDjG+A6JPrz
UL/C9vJgI4YqeUuDJ2mUQgrvzfY1o9GjP7UUdgvFjZHlA6j3HRSRsY6Kc9LBZbcnS6STncbcTdxO
asNF03hpEvX7MGGDo3nC71q54Opfj7S3FLvPa/bTOCeLL6c5aynXhQJPYOWg3KYj5astTm0KUi30
RAE2+c+m72iENVmrK1LTFY/CYZvFZI6FMVX0aVlK+4swzUjxuYOJkmevzC2jlCMvLSDDHwlNUZwZ
Ru2UecDhNFscrvjUWDdUFDRC4EwnQxVCQiQe5Nxt5oBM30WLBklYd1wiUUV7A7+STXToe2YlLvGB
5GXlOyaanfTgXlGa4+AvQshVyAGngfSPWG+aqtl/3P3oAX8P83p0IPlyIGf/dwC8oY9eapWXRbD2
r/Z1rTMLJ5JzI9rAqMZLK1oSn5Kk6HCCEGLbwRzBzjG3hO+vGa/QqgQH0Y9vGvq60lzaSJOH5oPN
BwF6o4fOCcVfHciLEZkQu63YAMSopprU255okajgVeJdKfPqm+58T4Qjx/JyBcTr4l7q0Z7I1PWW
OvcEQJmYf7qPfWsX2Oq3WySuJscAUIUCd3JjuYHOpIojHyqSQYPcADuagNnZX/H0fWbJxYCObY+x
bhRi8kwKS6Xe/ot5iak/hR11BLAStc8qD5lNvFwopd/FgmBLzr9Sy0dIVT7OUzoOL0b4O1TGgkEh
/tzn1CvIXB4Y6m/dsB4R63rgglW1qE8oN6JcJ8/n2LrpxhbN+cnUaz1ksME260kKrP7AFQx5Vzoe
J8Vf8P9oUZOJdPlb80/Yo/4stdqod7e25cUKzM7aTkB2LSA+94UY/h9iHtwCrjVmh9FMYL8KJdmE
QFhHhr1x9nAZMTuTwysBolKgRcrROvuzhO8dDxZ44aPVnt53CZ83m/j0dJeeirysey9zjtMZOiqM
fdFiGjegreEia6eJwWlAB05Gy9rYq6tQpsWw64RddRNMhFCH4wqQmTSlfF0zB1lcC/Hl2rjwkHXK
kpbLKcvyFigUfqwMHoDzB73q2vieCz7XQgohrkMFsqFnV0/pY7c3xucRoh4slRXiKey+G93mGRco
cjVIr2RS2R7pCTzdvK/i40oVjRXY4k8IRg2YCr35zHRzbXudxiqvcgHP6cURx2BF6egxGTQaRh3/
qIRtE9r2D1MT2qcz0qgd7eHStKDaj8R7eAhuS5gw+gpzztdZLHFKEAkTjUEqE2J0wH9V/WqXtJWB
1XhiAJ1sb3ba9d6pmqca+ZEBITwbbXp+qre/zG/ylQkzXPdOx1m/3H4Yt7H5uEAKX+IINzFMDATA
sudwpZkKYjNom0GiINDgX6mgi9LAqasx8ydmaknRTvwAaWtwS1vdm3PbK0ja47LJldIUy1LQgXuE
Q6dsbkXqLLVJabKCTpg4M0cgntQt0TGbJzlQ+Dqz5gNX7GXLaihEoNT0tFY7Xq8dpYN/nlq0JvpV
LnI5I5eHPHjZb85ED65/t7a7wNpqM+NxKsTBFKeVhLwMb56jvbfo08YqsshD7z1sTQe8VfMgmfg5
eY0mOB8Nx3h+tAukIhDq2Csha8OY+uhSPsCMU03z4AE+x/T/G9ROGsuGnpUjufzHFqs8jWtPN67d
gY2BgszsAZOW4uI/zIDVPpkm167imEFyJcOLe8oiF29CLxj78vko8WCN31TWu/bwgB7DIWf1b9nH
Xo8lG7EMCxcP8Pc9gDiIyzCAuaLJ2ub87thznq2wYedVHZ3UNLDXD2tDkGVb4aBfgtW12+D8sbuh
cAY1NCArHAirN+4G/6G2+a4E9Y2BeA4PaXoVUy+WKqKb1WypEthsHPhpPckGWVIl1n7MHgFUZGnv
sVy4D+uIDOSAyVmlgiDV0Dl5No8M0OD3tRp1lv1VFHzvVI6RCfV2mvkzsrncSiPpDEFVS1Sl6iAC
TaFZsaUz2JDCbwB4RcnkIET8vLedETaML+dXyL/eFLaNmllcTTnlxrwkLzSIOvba+gH15fgO84xp
te8W/EVTPnuBEYF4pEMh4jDr05RX/srQwzs7+7rZ0J+sA/3EhkVEeamElllCSxnfEnyjhs+eJ34C
6gRAEbA/+UZ23wpcpOSaZXPVlLgdpMBjlLufM7jjPQa/gv5TVE20Dq1AVkB3/giCs3tU6hbw+Ijq
A3T7tV727fFEtlNRGWPt0q2slABuCLP7zA5P1Pfg7Hsq7HIKIHY+U9PORLocrOms+YkmCkyojhWB
/+S7UaHoqUbim9qAlpmhT4fSdIe+8tjtKCQz0xTephBUh3vPrDt7ZQqWfqgMvJGni0SEmbV9obr9
TVVfm04mj27jDCG2faGsM4z0dc7o50uD6u365TmtGu6oA7iQovfvcgZ7S0tcMycOuhE/Bt4XbKSZ
sJeI9Nh0NlZUfwCr/aSjIqoIDfMNOYrwVss9Yf9RSDcSD6NjPxe2k/oQR7oeKX+IW2LgUsq8PNM0
PQMTiBh7jc+AVlA86NO3+IVdWHT7lUbbkcj9qau/NdVTwQ00vvFxzJnwf4J4ujwLqWdHsw7Yw7Lo
w0+pFPFuavyNsaqGiHuyvbT4wN3tRulySiifbM0zYdXp8W3RciwPnHwLLPTQhelKRYA25lQfGnzp
F941OC0fmH5LiXvH2dcyEILqw1r+MOYPhI5zmKfYhZ89LH7zF25cOxAVeVUluUP7lEQDqVYBgiuo
BAR35q+Du0CIFwoFziGANAkemn8gy5tzdJvaQLNCPBNTLVWV4dIrFF44Wmr7kkTYPbudhpluu37p
ByHL3FNveMogn1cztAZtY4mZFVHL0yzEZ1y1g65VAD5xwT/7oX6/Isr8l9ObFOeF5YWSxBaeEZW+
kEgUfsu72m8TXit783kyr+liqPam+h96z8LnsUxvpgAM4hFu7Pj3pr/PmgGfb50KMi7SCBCzeAOg
kU249blyj985xwOrYIXEc2dWwgR4E1Szg7NdtWNieME+XdeoqwNr7do5tBVuFq3+Pxkcn/8fjqFJ
MaJEGgpDL7NpS9YtoH2yTDoEqTs3EF2WYjCluXtrIewIsvR71/Xc0jMt9maRrfrZQ2kZ4/PrUXw/
iBgK74dGFsosKixlXOT8ZCeQ3sSGsG8Y3qZiBHEkEVfcFmYCM01FiBs4C0dsBZih6PWdQUXZLzQy
ixLLi0tQMw6RcIJeIM6YoHhINMi3rJBXv41Lf9wmtg3AZQF0EqrMkoxV+qQbmF2tFRmNqhJaVh/n
aZRGFC3RUOlFFNQIOk2mABm/EzH8KytHDUWMiQJR170TOER9GSdruwrTXP/ovPkK5vPZ58Z28T1Q
Vp9kSbXwzZbA6Fn6TYTesrfV1KvjlHqAGULhhhSeuQNuwYL08xxSknFpWFXcEenKVsAq6H2E/It3
pfXq06pac2Zelun89OD2TQRF2lNVQAfkdJKiWmWf0Myy+ZU8NPmyUk/s5cjZ0v8OgfYSbsvBXNrF
qms33NcKuIV5v7jvbFmcBk3ZqZoqvnUftJIfcQFiDNr9CGMeEbLdrFFq4rxkxSerrESyx+3QYqH2
ZjpkX8qM/D+Rzv/6BEPYnFcnN5NZOkLdoP7gnttUnK7ZKCzk3SmwNNYse9N9pUyEpWapmY+p1xAi
Gxwur0SpX5axMJMFy5IjJDfhD11FlqmddwOaoyk1224RfeYpgaBeS3nUJwFMHDWUE3/bCLl4oVLA
VZNNEGODYcg9kIkHuwLvQLriv1/qzyjblsjxNY1nhv411nRdSIrTZ+ao8UWynu57LDVbEOe6p0se
YcDemIzszQIV6dn3afd3T7wvrtxWIbSV18160+5WBDQvS4ihqGOG2JGvhpUWa8nPbbnmfHTFBw/A
eIBqlv867x7NTHmHP5S2x/Lf1FQcwc2zrOSodtY1W2cM2TbM/xtwfm8I7njD+MyKHUXTwCT2YOl0
6lJeEpNLgo+9fNPzsfpdD71v2mvZWfeEr+L97ZzUnQn0AFNlK5hmYQzn70p/tqZQaPmromiG1biT
Zljmmpp1d8xqrgLvY5R62CIJHl4+FnU90woH94Eego1oa+5bmiWYDrVAQ/SDraRfGiPv/B5HW/aF
hd8bWE92jVR5mfMzJq9yqOwGKpuPrw8jIO50Sea33gFgiAi7ibhb327rIUCSvVeMSpF/bUuw2WZT
BUCnPOBwzrzYAgP9u9M3ENalA/iuzrsdsaTUZMnDLiGTzUR8tKWG+9Qln1YOmATAuMUtOsx+AHVs
fcQscwFgmEM/d8H+2gcMRoRakLny2QNyjM7wC1s0Xm0jLVbONZAXhVuTO6Do+PvIsf3vNlMj0MSf
+eOvWITNMNObJPNxYz1j7C2kVxb7FKren1HAKIC4GLW1DF8yhPRUdjSFacqaQIZ0Iu8AdzY8XaON
DxO45IX6ib/vpa1XoeFoV9QimA+ANRZ++WI3RhNhTJ05ho+g5yaq7NClqtdCowiEN8ZWMwnCfaMP
5C32fveUgUl9A4icuY+8zoUnklV0zgtSBO36WHFEFlYrJlu6NsL+wuAnvOqunU+fyuojemKtze4f
h4i0uaw00gbUwItqPLbxrCTt+LrL8UKDkX7O8bvdgkEvaJYfcp0HfrEdFTc1Uvp4/Er9TCZsBqcS
WhdF4B0r+4tQXWZvs99faNT9MPD1UxDkYgT5DTnVHbEBLAMrkZKpe9hQJ+/ogXQ+oseq/PKG7XU3
II19MU1U+4QIt8q/4hqiGuxctK3ULKM8/HPzAUiOERxp7Ki4JWXxZEsZtTINKdqlJHnOXnfPTcCG
j0xdxVSAYrR2VKDBhljcwjBhEZlMOzwGluSRvWnLUbyfbQgfUs4HoU/nBKWc+jHvHWuWxcd0Q2Ao
4uQVAQLxwsJmEl5WvG7AwA+gopCjueFHoiRv1r/tZ5pzvi+GBxjPHWccPb+gurXhPRW95Cw2nX0J
+/sA7vVVCs0QeryeQTMoP0A/M5BkedxwcN+bjv1v/hCmBI+xnlOD4LWHCg83DQBr36B/W/c0ihKV
w9yXGcTfXpdDUWorv8XaXtrzDGfZP3rjQrX+Hit1Lq7eujR2ET4wTMqRhqtgdhTr+eE74sLfpok5
xn6nvCXUDCF4uzYngJo5wyilu96ayc9o7BKWRS5KwPjegVpTiKUwu5QYWs7NO1ZeB2w/lNTeDj9J
YOdgxtWed9PRrn5dIscaDNYsKVDqgtcR44sXwONk9EGQHkPtPjNGNN2g0M4tEKeR+OPVMdryZoW2
v29Dnt/vypJ7iT9Geg8l14e8DIse0XrpSD/FR3pN/7zm8Q4FFJnwKG+j9EWEbzlB90+DwaMVIXa1
lIjoxQePwHHGWRn/f6wP/3r45jVw12RgoymN1Qj1byI626Q9i+GIbL/Qe9VEZQg8Rck4u5qlvmok
Y4dSmR5f1/9oKIYGhoM9Fs0ueLNC0UI6cSlPr4znrgJKcfmPHvd6A8sCC0b7IyDEW6P0sbp64Rb5
yjfr0DJgenyUWc491aAjkQ0w92UD5azUBnildbKua4wX8rVhEwBX8nfO0WsSLsptzWbNvgtw3ExK
Fim1xvCqHvywLRcdPIqLq3GN+3xEJbo0CQQTNht/rWxlOLBdx9MX8a1ew6FpcMKkNM/Mv/2Ndyc1
KJ193359ySW3E7OSXrQJyg7xLI7gRkv8iUfP/+WVeboUcSXxnDzoTYxnlwl8wv3q9VpxL8qb1x1l
UAczbScOvGd0O+qpF/wjIpYeaQsYg1u7UNh8+wtcNTEs2ul0FIeGac/E0tWXOqUTJBZkgCgJHnTs
iAzGMmMQ+NQ2uuHKtSm0qUVMUgcsl1t9ShhRv7ekKP9ITW/1T9KSwoUVIGD/98TalrDIrB2P9bld
eFZBlp2CNPG/m3hnraWxgE9c9fJC/rJ32UHL0lQDgrXZi8sER91KkvjcqFdQ5jZXdPVAkOFI8gYa
49kyCgu0x/PNqRvUb4qn7CtQdkL7FC3NlZ9NwcgUkq1P5exxOaP+VLMhB7zF+cwpILi3gHO89CCT
UNoPfP6NyUq+GLviaTgboqbTO/64p/WkO1Vm2s3itWLLdP29O60JlFL/3UrirW6tD+Sq5QMZcKgA
5k8skibhICx1Z1gTt1uEbz/VOvKmQXQ+euPhSb38AAxaiw+qx4gvCp6Y6eXOVRYglq3RvkAEHhx9
ADNKcyeOL1PA97HQt0kBE/q++OGzTkPwwcRJsIX2BjnccFGtXWAv6Acevo80b4/g7DHlfOwZ4ajT
g8p/QJplGwL4ssgK0PO1rSArpldsP/H6SsJ9xPnzv29sFAfVJulg3w5te+KjHxDD5B9poByVJNb3
40IWVQnj83veHMAwnL0IpHo7AJTU58COQLSMOfS+VW8CmlELyjRPs8LKTjTrSA8NjKv0K90woRto
A2waoA6lHDA6kvS17cItn+wZTP86+JXrvLfd4SAh0Cr1Frr5FDJJOrbq2F/AQgv0MclsiiSatfK1
D6AZjDrrRN/APewZEeAco11JDL11CPzv1rOQY+8SqAHc1Z8DDkFOIQqCK9nPioO68elRMCrWJcpR
5hUahRe9DbGi+5ByI0CpoMHvJp2wBoGIDmgtqF0GVuyLJabtD56KdGSZZkApARB4+q0vvFiUbbep
clVn3yGVj6UNS17s4E7pZhFwQ1YrsalFxA5JPOBdb3STlx/im77BDEL4J8D9PURWWm0mv+geFjAO
jHNW7KD/w/20LvtlK1MNvTcocP4BV4FGtnji8Hrhy+XzrFlYw5+RcmOynpsZ56pahTI/XDLC4QtM
AFnvfUvERCtC13ta+LR6z+mh0fZZ6yvF+TusrgiN+4frTXbug64ipf7SSx0eCdOX4/bvcjstSRbf
6/aNM+pGvf2RgOzYyDGchXOMDV+CsgVWXFMV0YwjOq7JrkctcX4Qyng3hK+PO1sjE17HylLeyBiS
dIx0O9pHGg7rRqsoseyV24ktXIfct0m4X97Df96n63Xq8RSwx2lTalczkw7fc4sMrgvzfGbZq4Ra
7wVMXZWDM1w4EEQAahx3goTe3z0lLakMfHhEpOxuHDX1MVX5rRaW+Zs3bc8qqo9/fPdsrlQGYS2g
J7dDGVc38cyxy3NNzfXdcjMdo7IAuEHOawROrsUnfGzSbwfMuk/fImZAYOSIr/W0HQ0cL8pQ1wuN
toa4iQk7VPdt/0w4JmQVq17hgVySBjzhlwaQXnERWtLkuYq12G+LK4R+f4P/RNssE2j6Nrfty3kP
MTEDUgz1u6ZyPdtGhJWdquUzCV2FAnpaM2Hw9+JnYD7+3tpllQOurTXOAS23Fn6pcD5WuNE7iGf/
E/IfBZh1JxGByIIEo+nn7EQ3IbQTCLHzYczvAlQlWVJnrdHEkhgA93R/0MfI/br2+062r95gOcZ2
CduYYIf/fKbL/HfN0bLTpbw1S2/WI58Yt6l5Ap1bBNSA881uaKH4lACceuyrOYKK0SwrpeXQMrFP
P/uy5A/Nx/WI2uZRcdho0ITdetyy1ltZ4ZKJMfhzvBE21nLB7jXz2nA0SIpzJsVebWMJOhq/0X7U
VDoWt7bH4ZHA4YThc5RAqa6UNjtthOzfw1d1kCx0b9F/CnWkXGkVZCPVkh63gi7AutvWmMbUyCjP
A1wpUv1wfcMGlpWpaEIFcZMEIK99FSIkgDSTOCj8UZHRFTKy39BRSgah4duTbFCc9S2DLVFqwbNA
MhMlQY4bZJIhsuO116R8KC5OasYRGMdFvL++ZoZL8Fbxr3jP/Xm6yfH2VgOdWblggHSWNRt8yIO5
quMrcTaOJICbvXz3i4uH1P3lEGXA49B+qNVR3mv5/pM6rpDWEouF++taWUSVHDZhUGK37Zf7I81q
y/oKmn1eTtDMPd/2x3XJ7AlV1lVTp08jIq7LZ4jPZI90jPChrtJhE66jLppF5mz6baempc0imUU1
Km7WzGJC0f7VmXuoX5p7AVeIoEfQMhfeQEGeYSbnzJ6cbIySUPL3fHsQfUevOvKrxYBSq/82Ta5J
ihOjz8Qo+D0cWVqwPZrWmJDh4warY7ygeLVL4Xfzc3DtyuclL9RkFhuHS6orLsZyOZJo6Db0TgrM
T36eBaiU7ALXrf6c6Faxo/guwuwd8xXEM31CRMl2LeBUWnAvfbw2UnRC1nbN5NY2TliHf7zg0x0N
+sN1nCZUW0Xuc/NhSvntikqpDmwSZBF+xpj/Mdhfdtkz6DvIJP8Twxh5MYVeaP/egafdx+75/x2k
gCahyruEwaJqsUWzNK68RehcWAM8aPcwY1Tp/oK8fUL8i9pm8A86ZSlV8/szP3spJTVn8ceu+aw2
7ft3eY9WTp6WsHDFcZeIsSC2drzjDXxpPVRsA/h22Ns6dHYrRP1x6oksX+2xMY2LfzuNnSaKv6P+
tXe6mfIfUXkmnrRGOW8EUd/DMKjQsDz+XycuXLSS00YnTOcRFLwWVKFNVrTkXIaY0PyajqDYvvxW
/nJ/7PLroslpHDGOl5CVutqK4ubnaKjRury5tU17O/OuB2PvGHnB+2czuMhw9P0ptZkoKkHLKzRN
bW3+7cKkg7gMP/b5rI7pDC3tOSSkVx6OAlfRxH6ox6n+ragC1YJ9BOja/JL42OKsbYgyqK6Enajv
KDHLWSnQZ12aB527mQgtN0NQ9kWJ5j+/IMmh31Xj5UefNsDQV3L7hoSvH5CSAWWkMl/uFcNw6FoS
RvIGBT8BQBTOybsiKjBVm3uti4tr2Ur4M4z8CqTznByqBCyVQCEvHvuNyh4R+WQwZIwW8Qbn6Owa
+sCLaMxYdOlTgfrCxt2aFRYfTVHUvdgAj9m8tFwgYXkzNqRg30MKJo//q5KjUJb4u0jKOc+xhixa
lTk+pJtrJqQnRjYJHMrEC2pbWUnRbBGDbeXH1Y2QdkSP7QCi/u63OaR8778oWH1DMtA1hX/g8BZt
A0wLLHYEvTeTLnnRWpnvx1Z/qHP72BtCStPSKTJhBZtC1HuhLEf8iGBicRK34IYp3qYH2T/69w6Q
Fsq8a7q3hqmi4unWbLjL+f0EXZUJ81OY4w4yLwEgFnzcxTiN6+68c5NQRnyevQySf9u7VXBvT1np
lLri3kEPh/lHWXOeA9CV6glp4qIjpjdgcLSAXPyFQAco/s+F46JyBLDd3eXJ0Nzc9RjsRxX9HNva
GLlLYC5hzicvu6/HnQHnSQj3RFZdfpLkXSCvjSo/zGGRKL8oTv7rmx2aaxQSrpSNHn7HaydWgOE2
/W92G0hBxZxAkzstd2PQiOY75gSd2rmiH7Uqc2iRLcjAyLThsUXRWdnSjSJ9grZL/Vuesc8gqUW6
5gqq+WZZomiWLQLkAnKvxyfVmP5yJaRMZGT99SFEvKsodn5tquJet/ipRjCHrEuTxSBc41EG9P9M
vi/jUw/SrQ3Robp2L7SUsAtfaFpeexRB0lTkY4t/bQ8xFaPgTIIyfH64XBEpGzwi8BZgk4s7sWk5
RYSt7oXJzlQ7WjyIzovdO/s/XUKC/ns2fEU2QxV/obF0iVkxVJkP30o8CM410yWEb/pVRmrwQzTm
nBblWOxZKPYHx5Lk3PWd78sA/ChqIeDJfT6V3V2eM5AZgFAxyz9q2yzoGHS07I/4BV0QtvjSrNEC
pFwaB5CSYPEtSjl9kAYB+CAI0bJN2Tm0zJcVDxMs6ASi3+LhsdJv4L0kTZNgFgf5V2QJVvBrVTXQ
QjJcx1OxF29jh8dmzSOZsWrcdy4B5EjglI5fG4iw9bmjSJpeR5sB7EplSqRjlf6fIvb4x3S2GL73
RnZa3kffu94UmIru6J73NonASzLCU2u4oMo9cS5i2C3LYd0m+xgL+TuYaHbC4XBne6aIOjlBzUHk
XfAe6LgDeTPk/2MrSMjePYrSdGLMDK1jIoxTc+YV/rmMSrzLPn5Y5GT6GqLlPmxKdJtdLF8P1d+V
LhGMRTE0kWWS5Y1eNkWhf62oKV2kHHPf1K3QMma5+R7G+XBuT0DQLH9wmeyQuVrhD3U4TDnJxhFv
GEvromIi3sxyBqBKjWnUP6NuZqMIImMlqIr3YBi7QlXMZhxUYXZBadXayR5cGx/ZiSynL6rsAeQ/
b+B1D+UsDjgXiuR+U1G54MsKV7qOmWD+tTAfz0wejqBZWQTF8Ic4JUrFFJwZJ/FXGcuXYhODtvx3
GrMtVfn603vT9X+uR/A7D62cIeJyuLAedWJsG3sFF/+9JktQHAl5unVwQHEk8mkx8vzYWVMrbexi
/qbgZSOMALS9Rx6ZLld0SVDIai85vnD5c0kxLaQD/o8Cei1tq0GLi9GcsnIThcNa6kWpy45H+bkR
adRPMxrik82BvJs3TbPHySU38jru1tdzrJYFP+DEY005lwRhAThHZccERRbsZwfbszVQFmD72Gny
Uerk3H5FSa/3t5t42viTOIT/5js8gV8n9bGkk34998EgrWxX6Cp/gwpg/SjYuzBd+4ULs8yOaqO0
XR7T5wg+N1/Jb2jHFP+52iJXCmxjfPFe3wIr18q+b6yykvQn+ecJhtUWe4Zo4mJYu8evWDOqf1SD
lBeVmpQ+ig4lrn/xQL7KeMIqxbN9+pxsb3vQG437RQc40r/oB+NjANEXdyXhj2Jk6/+nrgRsAheL
SBLx5Cnxdc5rX9AHZn1a0iU9EzxJwcpdk3ZwHYtCEOPQ7ipeos1CCKltBnrad/oNX7sTFy0HWkbc
PsLPqL3YrUbZ5dzvXKFFi8u+f7MjvhOn0ViENiKyk9mgMO2IZT0OiR8MLtDi0Czv5xfj59JbNzmS
+eAQDRL/13fhXPSh24ww3nriFAYn10LFt5nOS+4T3p7YJ3n/QeiD7BOS4pgAzUl7QMZ0vJIm/uqW
KcRPo8jc5GYjFVeY5Te3TufTadKMqyRxwAFKPrRGeX/9901TUkM4xHyIQIs8j/sclEScnSsyyyY3
NL+iIRphI2CTJj4SaJlChm6zJyJnr8QwZBboyPcDvUA9Z8eGhcjutnJ35C1GfiG79Vvzdq40kzwa
W3KuulyvhJ+6kpPp5qtrj2IrZZeag1x8c+C/ihokk0LysiP4yuG4ccsw0uve5R7n7+YWvdYHhJnv
KLdVtIKaGAcJU/ytFQLnuvyCUwYf8AlwIQJKUkGUdiia+nXl2NqcHrI5/sbMXexlETERyTNpQx0t
RuMlv+n34Sm+e5/kj6JEfg0cPp81SlnnmT3+/m6Jja7N4Go2OYh6O0FlX+HmhbvBMqybtsF1WOMT
zf1uZ23+Dk0io35RHPFBP21TjgS1AHN4qqr4/yKsppW7j65cmR5vQZXL/jiCUVRBKOPPQfOWgICx
XqrAAGvqqx9nUScpiQg5ys3q7SV+TiI8nOdgKDpG+ywT+k021LuzjGo1wEc786YYCR2Ik1GwPLM0
7ebUTOhY+pmVeJn5Mk1wAjNCjya/qV6OR+QYFCgf/M1UZIwaGRMuLFb9VjhD6ieqk7ffVkPdyOCM
0jIDgI4HVdTRW38JvchDG8hUOmJrywKoT5lKOXdlZn+axgbRLizGix+H51euL62e3l6kj4pUcprC
GqHX5ULJEpE2vKFhJN5QpIQoCmIjOz/SX4WdO7jOpjqjD9AZAowYi/HhWp2p+M2+iggq/8g1zKWK
YT0S21XvTvrZ9vyih9BvUt9GqGZ4WcWkgMocAScAyxsn+xh++A9EFPpQv5lol3+BLG6Rz3EaJloi
LlIyqL7tFWZekjceq9w2zurawFxyWHtcAEtVwouzUg7qutRNvJStMjWGblHBaZh4zB8QOwGCSkFI
GCcwuG0fBUpMEPTQcKHJpfAmERLs9hwH9VrZYBEuXXJsJ0+cssoYRuoK8DqMTEGNV0wqz0ScqOY1
FIwUjRPi89ErUaVF/Br5T56QKq89M9J6hhJIRJbx7HJfLSr6RiOfc8MqU/Q62ycfbmT97be63DZk
5cRhjOh1gRzEEB40ni1bmTxGqT9vKgQdQWaCUcN3QQ/11KPQ4aJjEjITkW721MjnhURaNFnWpOKo
o9e6KMULKcA31hbB2dhdiCwYmjCRj+5rFyOnc7mBDzR3yna6TRhD1un0zQS1LMn93iX8+rJ5qdrn
4PrK8mz8Eh4ourbq7Nmplh4DYa/CNTwbQeoxS474tmKJ1qViTu4pGFaeipivsFs82OyymSI0gK2n
om4sipCpAob/r8UnqZ8duDj2pSo9CooZiiRRj89k4E8FweVWZ5X2K13bJe0QzAZlFtMBhdKPl3Tz
EdYZwOHJedSxb9jNhh9NL4BVq38YIU4AHqBFpmUDaBGCAMUapiaFY+MjiiA9YCQ7YSkHnPtAvFIL
BCm/i0hdp+NcuJpC5sbgYiOVNWMoOLb5xXwsMZGOY+bHOJmRpvhUWj1BNUsP34pITTwZcKt3S9JG
Wb81sQPnhOWQpZ5yOrAVRiQGpxCCxEqPH6B9Lokzjgd4nXEDS2os65rcv6UZBw4bjF/dxhOt46jN
q9EMJxhvoJqMNdefROJ2apnaaq1gsfWtDEStTWWiHy+AUETzTzLFRgAyxhMyTHdwO+qNMwOy8dPJ
9Z+otk8UVB6wY8iqd9Luv8F7/mEHtSvGCqjxjGGMIH4YoAwew2qklwq1oT91QhJOX2UHuQWl2NGu
OiFwJ6TBD+UKgCQxQvGM3VPz2RtVXpEEcZDt72YMa9W8XxIebkGCJpMlZAhqHYTODuQ8yFq5KClt
tkJjQSgMErZLGtXq275hlgB1E4Td1xqGSsqgUcKpb03xA/boF/7O4/nII+MdWMGzOxozAuvmk08J
6HgFs4WJBneMUv2L6DkPecZQe+UPRUYDwnGgmWfdvBUwdQJ4RyaLKTvoXFT+Ca/vz/quhTAS2diA
WIF7qWyCkfsOBRZ/Nw2/TljC/9Szb3OMc5QfWNcYZyivufM4zVTSH++/9IsO7IRpzUG2wnBzJRW0
h9UpjghKmuwolrMs334qpqfxc3gPUG/kmtHBoO73M7IS3Z4grKhYDVOixuzNYL0/v+HB5eXJRwS5
ANxV3djmFhtFEd0MQmdourLKT7cQ02UEvWl9OroRo9TEW7aYMLjKT5TGI9/6p+NEwpXLJFdYeBLN
dznpfemvszo6fQBqgTs22wZPZxa+CGZ1VHy/tnfgdFNhNrxh0+EqwNv5AUBNCA7JznLPozksx1LX
KeX7+gtKRXsoUkZVBD+j4X+ePKJfK5MvKJcShJ1LgCT3ydhxxRFEYeZcZltBzuN0PCyawrV+C/Ms
SFQjW8QvyvHZlHKFXAA+TIK4bHiBquExmHRiVrk/IUnUXa1lDt8Ke/wl8YuIc40FUvZGcAtYO64T
B7PxVh9CdniNl5/O8BKUBJmqo8xXV4l6AFcFa5kfooKYxsNWIwVfFcDd1dR4frCCSiUaepg1e1Uv
Un/ViyJ8nPckZy4WGgzQQN4WW/l/Uea8BRmvjDGefuf3Dr30ZF6Qe/eoRG0CcDHQdwrl5Eo15OZw
tRGCxY556RNOUFjjTijdS72yZa0v+U1Gynkw04/I1CwFEyYEwnPnc3lst+W6/pisCVYq/xi69l3p
0LUXyrgVmoSV9AGp3n6WkhPsGaoqOl6oA9nuLonV3PRvRhZxKNadqr+4DvjlcXzzZu+LgiisRko8
Z+CyBGra++fPzamt4ssn4n0qXI5oAUrkzjw2CwHYfmx7WBWWiWezN/ZIj4JQv6mv3jqFapx80i6g
BX8DNZKeZFcAQFkZWOZBPGDzHsYOh8UmED1+v31ggMdyJSs2DKGX98CiGeF2UfOJt1i5Gby2DiE9
g9r/viRuYE9zhDZWj5JuLeAxbD0rQqigKAH5Yy6jhv0PBcn5hZZL3dYsEyQDqlStmGEi0A8zRgx5
BNwAhrB0RZKnuhDZAhoiXGwkknYyFu/c9+YYw9fjlYb4hB3sCbK9PAJ5j2m0vIUr85bxaFiY1fSK
wzowYh1U+1pOVy30PR0d8a3gNSVYXOHJ6/Ez9I5BHDJO/xDs4pGdZn3ytQtjakaD+5OMvqRDimIF
sCt7csZjFkjpSD0z6WQP93qoU5JjBbyC41KcgTIwxCUF860LsyQba5Dut48KRPLWkKgHF0ocLYsP
w1LukWLmhwKSlwtHjtiCTMQIt/a9rFJsCbkBxduk95UXxKakrCfdFnVHOLX7lyzXd1+nINggS5r7
ZPgCFA5bmhbMsqS8i2JY8c8BPmqDNKkp41XvQ212N+G+qfTylvBMll3Qxf9YBTdXFb0H58WL2o+J
4yNfLBgeYpWtWA7sJF+23hg1MvXRM6J8TjdB5JJIg8qeOuzJPjkgVgOvh0tKn/riBqMbJ01v8mOP
+D3a2AZ1OXzpXi70pHVSrZeigkQ6aNHTyUgnOZgOMWsyWA2cLPb+efKW1jaHdIrQ/Sa/hMc4kFQh
sVcMrCwMVRxPAvDDM7aWIfn20ghajg03+3UvmErzRU/wKJoWeLukBnIZspYde+C9AzNXPJNkKPEE
C4f1mdFIq+Bvf8XH8GhKn41jNxxpp8Twt/vNXjH0y2zlwQuBci5M2YmLVA9C4QP4b066QcCTri0d
HALH0autzbdLMFQW89G6UxkjIUEI4UBu16Vk16af46hxkdPk7CRU9yw88/K48Tj3bAIcpgikgG88
zBcQwye7bMrY6bM6ibBAon2r/8TCXmxY+1haMaw0MhHKCUZFeS36VFyjrMDTaJ36TPtkYKsxPTdS
EprdDXwu0j/RhaMsJDbW7y7SZad7P4dVkH1b9WWTxhUnGlX21YFJ7o7So+0Xs/yxqUE035/D/AB5
XOYKfotFEdL1t2Hh58/b7PlBR4EUrTuevw+tp8dv31307ZAfTAzB8EdNpPHky92oXLcLz8CXFosu
6SmbsDZ04oRuXPZzPGLeTjqdSOV7ZqAW1wtvWq+QoJMKN/TI/vxThVH2lvEmg5fyvlZ1UUdQuXzi
FD8f0DnrHerHj8lRCM7s6SQfrkrkOkgm5YmcvJIeIKLyb/FatGUaANEWv7pCCxmyEiZMb4IBCQxM
ukb7N35Of0MaNj5gVHH54qLeHWTcgmYwvrEbFlHSAE+4+RSV7YJNc9v94qQc+QGkZ153cW1erxIw
VSxMimrGJTxOz+i7Ui1X/W9CZJPcku7WrfDI54Er6LWNji5vsgQz8V1KNDPp3H01MhIn9L/z7Ub7
qg1cMIgf27oyEZlGRlOKzZW5ceXdQYW7gdXXwZjsySH46h0WVqRR/xF1h78A5eymzzzAZQtJA3Nl
Y1VcXnw2xqbp1jwAl0Wotz29AKeQox7cynEEsVVIKVXg94XkLtL8tYetYkUrHgF1zRc+3imNhOe9
W741vQL8oqR+TxNMzBueLOGgHhtKu+bYa18V8+2LGs7GOnqMYxxZmlvHWh3PRi/H11IHsF/x+GYF
nqu/tdAAgvjNiKArfnHZurJlPFIUVTp7tx3elVMAgdjIZqwihpfWBoSX82ImBppC/Ly89aTcrt5m
Z177Emm/wnfxS3OfLuMMlq8kJCb1Lw654XlNbM3KtP+hO2p/xHvXF0ZpJMKGXD/0gWYanov0Ddp2
OyhRXoiH1E7YaFXsSfpwICkPkk4OJas3AypoZLhu1jdKhJNRXNxoC05DB7ylIh6IOFgZIgKkn2wY
C0JQV3ZizaSUyzp/PXaUHmYTeZFq4m+hEb7oYO0t0E5W5eDL37BYrTd24I38qT+u43ua0Hz/xVTX
BBKOHXLQnq/0vXmdo9Sn3L+FjtmTT7+X6vZ3ewK8NbKZEeQlBHTVL7MAXCuZFSHWIHGj/k9LIfyY
EfvG3R7cJbf498OngQ50tCGGo0ilo4qykFISD4JMDBAvgZG2MICn5bLvgv1LypkA0MlN7ACIK0Yu
rHa2EtL8G3esYvKkxhF0AdPX2Ip+Fa+j8VnlqEkSqhKshqFbplfSYFwUb4nPfNY/P/d70PO4SeqZ
aeeLvXmV2lOc61fB0zT4qmh0rOxah8NYeN+ISrsU263grN3clzcjKHK4yHcdnY0WeGV0HO3811rh
VefxL/fkfTK9dZyF1/PqGVlDZZ7tw6oiYRfxNAfUwlkAp7CwnBAACKN/+mmyEeDUJ1EPcv0NgRqI
zEoYlfszFOu0cgBC+sUDk8bdTVInMV2mzsVZAF4bw7bT1oFNk0x1CBcttGaQQbIJo3caqH3BPgdP
i+Owswi1Vv2MhxYuuIR17buOrj9LJNeEkpI1DV8YvR7bxPhJpTKQWQFL1NYaufMTDQdy45HGK/6c
oRCXAsIuEh7+rKUrKk1oaNjy39YzyVaAfEoMkUO0apwiHdeYsQeAAvRaVqpbmcU0Im2gI4xT9c8G
KiNCbAnzUdVqPF+2uWojGkBjUsc3C3Aos6ZT6E6yyVDNZVppJ6o4s7bFWo6NJM3atf3WRc7VEpk9
D4+GYCVEurGRQIjLuNFE8diJywWSyATBUkCCGZ0F2TEhvTWErqZ5xGxsbDGunL85npvB5/ugekP8
ZncSNkgyLdlVAehTKlZtdfFUwwI6FYvHlFY+aObFtyTql9Sm7YLXoUVG44TT9Kq2yrAjaHBv/2f3
4Cidt8P+wc5PnMVJocCF8PaH8A2EnMESMXva+M32R8RCIgW30QPxlqcnWZXq+/gZtDPIRXdVfg+u
IQ7ae0z1EsCMJBFcmMs6SIDik2uKadx7YvuJEXU71w6HCD5KtlIv9gcSL06gzlHB5xRvXGvR8nCr
jmMFa1gTaDnfxV0fqJbAFmY8cwnO+MdxUVb3G01HvK9/6vc9b/wIiSr/DNcuWaYfK8/at4850WbB
tSsecr3YsdOzmE7TA4D3zfg660QlEWrS8natkAG4UfdZTBMUdIzEWC3Rwr5ouspjFq56N7KCh+gv
JRGet+LU3vxBfL0wkQyShlS4SV3XG+TIcPrRBqiutG4D45be+jwRNY8oemkAYrbvKLtPm2xgahCM
lWhSzJAn+Gnsw+JwwksziM+zyaQCUncpWDIKek84ECEp4kK1ud36aZOeYQhOarT2+6B/hwp0En4S
VtVezbxh+3acWutRtXbZ9Ug3cnHVbJMxjqRwNLtcNIZ3v3bN2sawmrPUGH8aOd1W6L0gymJfi+LO
4fkWZH3p+WwcDpnIZjWYz0VGDUA9oUSTiFAKMPAd+qZFcMsOiZjOIk0CCYkBS5GLHJoTAUdO2OoR
cf+268rtwn+yF0YRqzXhYbGHjzMkMrBao5skRQxs7o4GgO8Y4tI64A+NjfbBKd1Z4fHS9NPJM23j
bWqvKfVy5/A9lfbUQ+yGSQsFQ8OfC5urpTupaSGZTK6YRQ4K9qsN8qEN1tGe8uUyLQJATyl9W0Qp
/dOn21BzAOk6CpL2b3kzhxwm5M8tlsu5177JIYvwIPUGt8iIDWnywfK49PNLWNr83scBZtLAeUUD
kuWorvtw+HjrnipHqOHvCnRyEzRUiVhqASf+Xjb+yhOrGy6ify6CuP3fSBB+dEpcVMo8X2V9HJEK
fH/hhaHHA2GLvkp5ckAHmPVCbEBdKBNLi57sn/N+wkoS3xz5fpGADEFXqDfAekY4dgP5aGcrrLBm
C8ZH/ydN6XNutQ+wCiDR9oYCjfZ/E0LZZjf9OgsMOg0SAME4I9EufmXJFzW+u998ToybErjht1Ke
22YvgD6zyZJrWwMKg5oKqP/Ii/d9/RtDftTtmUAZ4kqKvOlqOW94KQCfDsBUoPYeYobc/goH26vI
nO7llEW2lAouY7Nc/OpNuNqR5z8mQqhWnqfHRpG9Ph89eVs6/GzI645DH17hEArukDDpO+6kq1LZ
xpGCvzhMWmiKeF9pR6XCSG4nkK0SZ21PZQWiK5B2458SSX0W9CujshYFG7hB3wWbCxHUlS6E53e5
UMmwdJDJsPJIn4VJb5vWUVbLPEGq+brxe4pirYwt8EjGrz/+qtVBxrEk/zX4HN2S2d8jJcSoshA3
+xYuUJ5zgaO4G0wIwyzLR/MXBkKZvcfS6M4eg7Y1qdAy79Ksp+SCioLEztitL8w2ClMA7rl4i0lk
SD+w+EMbyqyPdX3tPy6I/3bdydbq0qgNrjFgKLXSXvr9uwyvRcTpgkTkdOaFOACUPBmeBKpItEuJ
9+M757DhY7Hp5yMKlXmKmpTCgVM96sUYECIEneDCIve86gYXNOcHxLtMDH+vc/k4OJJBaD6NEpe3
pYaswQbfeKJa8DNvccDAC95dlcjj8hyGouMn/CHEpiOjMqF8CaZGsZLt4H3WtISep/uKQ7dhvn4w
oFSf+BHKvLsQCgAmq8GaD1CApe2Um7/RdO3XAWzQN0YSLFv1/+a/vonRi3426edzP+XFfOW4WlmA
0lhwj2GWAhegacGMSxNMw/PXUAX3p3qcg46ieI7iJTqsPK20Ux1Ln4diaR3KJKPlKbRODVeoLfRz
nhGeZEifedR7m0u/WZ23Q1pe7RDqrO3WcrfTri0yeUiDnEXhKVm/ledDLjfUeHTF4Qs3iduWL0zm
eOvb/j2UM87KgJKGsXT3+FT96l06hfUuLovC7KGVMtp+JjcRx2Nr6pUVOV4KAeFcSF/IWXAjG9EG
ZNSp7xRLJMq0LGVVp/26uHY43N87UsWDJQF1S4uqEfECeb3jAe3HXbAj1b+diatDN814bGNXfbhM
I4+dXVqt7kIjXSVkpE3D3prKTZwUPlWLkOdGNefDhwaLTmEocUxM6zn98LGqeHCvb6TL1FTpKcPM
66wdhIKCbtjEQIT7NkqaC/NbGBRSZicfmgOvcAmqLR9sFlRRmJ3BehXyg72RgUXbsGsqRNBlZBmK
6DcPsGXmgNlceKmrtnifO8E6fjjoGPBavqxAI6bXyC5qxEVkAedKByNDdZrvNyQ1CVSSWAwg9vdW
el1xQ2P692jNqfVEaAUABPy2xH88W61vH2EOcKR61yKvyQb8NctH4l9OYWb6Ccv1wJSXmKRH6VUa
vB55q9CO8OHPtz/DYqKVve5FEmFYaEAler4v/9BCKgeAhH3H5OXSiQXPrBZ3gc36LpaUeW/ea1Eg
y4ZJQ7XBs8ICKu97njp9mjDbS9k9BSBupR560ACjV8oO3k8EJltkdYkhzZJVLVVr44CYXpf62P63
/Nw0d0/FK39t3nZYTElRcSVJqdjbxC3m5K5KStrZy/jWJOaq4NPi/7nucMFK6nFhRcbi23fuGaAM
z4FIP5+loa6I37q523jYEuBGZ7ANfBBsNwG11h/D7bOWNmmnGTHcHYzXNJ9T+PFsAj+zAl0foJgA
gGI4JyvsJdZyI70CSeOyN81ZO4PrQIHDrdmGDMeHOQyqv3Pla7VeVVzHY/SIknII58XQnh/MQJNV
KzsfbKXFuDl/Lv956AOiJYUmv/IegqWeI6O5SmWfNXfgrG0qx9eFdqYT6EcHD09XiDihspNX2xFQ
pfZS5w5EAczzEhEhB/pO0iWDf/F8cPsJD4jvYMgsughodn52emgXwFUsoCySrsxFpYiq/l0YqMCS
R0jmMMeBc47YdV2rxK9bppErOa3a8VHMA9WOR8nIMLnYj+e41uXsV/USJGugImWXodZWJdXRZNPs
z7Xay13i3fhguyFclG32V4oXThO+toXjQuNMSxBPbZvtpL/oEUcNUgO6/F8dBxlK7HQMBS7+FjZB
YhjWs9AeJfmL/8dhyVcz5sxbHlOgwC05NoxjAqIcuTEG7mcm2ZhBS570iriBla5kKSblzKn0Zvby
+Tlx4xal7JG+WngORxzJ2AHe30Jdn0d4defG2iTE9HByWKqzTRGL2vL0R6uAJCqk/HbN4eOG4vu6
cnpReEodAyKARYhyZyoPY29jGv7HovZqLrqlToXs1NOUtRmV9edZcd7bGwVsvokQ1pxCXRlcszqH
1Yiw4B5DeVdA+IrKg2QVFcg42igOe4L82LqNFE/DV5uftJb9gx5y94ew/T59my8RYFrB5rURhZMu
f6tKHfoGuDL+oPLrYTu2rAun6KwubZw4C/H12Gdj+nfW7vKW0tmMwSv7ouBDrbgOX9eYV4V/DE4z
8GyfA8eh1w1jk/ahp7bIxyufJuR0LHtrVAaboPuj+fxguZ0ZbaBVsredSxLlbj1i90KTRJYOJd/C
PbrCG/u6uegk18kGu5bn/w5HDtIHx5oQsvnUQ+Squ6u4IypOOXW7natcdryBcMauPTiCO6Dbxxw7
n+6kmHHE67+2GwykDrW2vbNoKzj7O8ElZvfNlQXThQxb8tZdlCAVdBF5fSKIJJfpvHduxvT2OT+Y
FwscJhZRqLPITEDMs0O3xBp+mff3gK4Yo3UmKqvn1hpsHMdGaWr/OOfFvl7AKBrQcqoMuqKJ9ntY
Sd8r93n1n97s6C9fJ+GlOsaoWpVC2SJkgOw00syMeZkhkFiJQPtgwZUaflB3K8gbe2VFB7lqI/eC
0DyukgAg4z6uvEyXtvMP/G0CUcvrI/wgtCfs2iWg7Xpdot9YTar3wqFdf9C5uHvh+J3gx2qAXs7T
1NKnFpzytZRd2FcF7VUUWuzDMe8vLSLex7j2IkPbo6NMiGAslGjvdIt7iYxgdbcAzRe9ivmE4rxt
JDdmBXAWcOs2zrDVrB82/2V79eWks+5MtR+hLOn7NVFnbwVh/bAYDShV01hhRK8HCuaNpTkhoTzk
XGXeOZ9Q2B5l2s491qmxQd4cupZuIzdpoTeHcHeVHkO4xPJeh2xTI674c8orvKRvi3N7bwB4gNX/
A3KHcjuclvFpwQt/KFEoDX2bmUQkHcXsKDAd9oQOvRIdW+geJIC6hHkPuXxP5XqM4oxGWK5RCU5y
72FtX05WRpTF605PzphykKSxP9giolNvM4Q3xvclJnumMvnOVGrVwVTChDSMFwjJPNOYwrcoX0cr
MEWOmbfj+4c1prtiv5OD4dJFkt/dvU6XxuqOE87gzd5e/kntJo1W4cxUeTv86Z+a2Wb7qswH+uHr
tn4aP/e0jfKzadLjb7IGOUX/ZNnCu1aR6YzBIlFJp7WOoOaTdY6XmothsS5Fo+06oP0rOJin8h83
c1z/X+ouVSEoY2xFs0e1krQGssCtKdf8kIB7hq5Y26m0s3qKB6G0dU3r32R5SRqKp/h/NJPKNOCr
bbYgQD16oBOOxWMJIpPP0pMZFaihf2U7iZdk0DiulZXNX/XLu00R4DCF1Q9le39obPoX+r/zqgi+
YrCM7H1mVryz7mUYrJI88y/5Lyu3dAkpMPKHxZhFAhjYNtycr2TpxT43zS9T4cklhffFGRfD7uUK
EOCAmP2njXpvvH/WtfsZZULn/v+vaG6RVA7xs2rZCuEXfPxDXVVCB5BK3wCdEjvp5Nc3xK8vp4as
mU26Xkz8cM/VnLIVSEXx1aN65VbKNwS71px2LOzgVpk1uSj17icXTaLT+SVHOlPfvjlH8uxEh7bF
YkQbrKNrBY0zO5YD3IEzYsd14m4/4giWn/V6CqIZ4jGNz5ixxZ/VkusQHLS5D+EKObHdomz4+3ai
9gkfeqcR8YTxRnJZ5dzwY13+Xe5qvuOpXTL3rgWZa6xPdNy/S510fOrnb84qJMbGIDt9ePy9zdnb
lF6ZKSSiljAK62NmnIgcSrgxbTmOOfUtdv4zftF7+6JYnB5ekWbmreH4HLKTJqm9OHrkefTbgja4
tVX1cuDQR2VwJQ2QwlPpqt65gxwqkC29boi/Vthc2R37UpwFw2XG34o26pFB1CJfhWvjSOxSsxHH
cxoKfIPuVL/LpXkXdqL4OrHGSQj2GAegz4ENCTn0HQYZF1TDomFnniTs0gf68ry3lb8KAkbVc52s
C/6J1RGVkb0/RnDK57fkGikR3hc7tGHnLUYeIhgmI1y98u6DMdjZ93ZYZ3fNzxwtLcGH/nGAvzgI
QhWzEo0ixVYwkwdD5Dw36abpTciPmrdZNTprVKL5UO1rIP+RbTO5fwXnKw/GUKSWzQSU1qa9/LxZ
o9mAQZwsz4HYvU0FtRMDE3PoTuWbH1enl5+j5MXPNUV0bd0FMTgNA3qBixGvI5+OtfR89OUdcwnc
E2ckKfsAdbJaxm9yxtXhuHvinS2QSPxGFYOY44J+2nxcu2xWHof8yvsno0Xi6mSk6xga1OjZ9601
f4WmWAb9z6ZaiV/BBX3/4DrsOK5EG3mj3P+3RCwy+yHDk4AIFZ0wHG5KQqQBKVaBDghsuw7It7vA
SNVFjWKBsxUX0L5cDwCgMB8g2O0wy0UaAHRMlatq3E4QqYSLkVkET9nzAaboMchDquWTuvnlreYr
pKNetPcDWp1dn3lTVu7KF655cVlT/DfVNOtCkLoOtHFgJfHwn+hq5vvZvaja/k0K1xPHfmjQgIh/
P1GLlWA6RmREV4MbrENuwm8wSpmnnsM3vnxGSANjgUfzgOfWQWT6II0vn3SqY4XXg7C9J1LWi2d5
DXxI32ZkDC4rLbxei3T1qf5YDnIFM5yYDvzIGkFg3mKwnzkLNzHnqHP7L8IUwwBUZAtZdiH4tAFP
Y7mjV50CHN8bprSGUOhED/T99OuEZc5Qll94q+e3dshB+LgFCCIbiA+ZAAZ/124vjep6UXyLIKdz
DeXSI0b+EQVAYCrXsD53DXpn8OZCil3foasddoP/eWZI/A1Xwnr/U0TjLB6p97RBEtbTV7l0dV1O
HJoZjQ5ZDqlI8sY8OqlohvOSd3oH4ILig1RmLDpn7oImHqIocBs47LmjoiUtHnDj0DvG86ilzLse
bSsiwwnoiBUVm68HTe7cuid3x9qzVB45S2CAoPzhJYX78C7xOYsryIecB4QNo4sg+rNpwcYpbptz
bTF6OcVdKQhL5MXC3mCicGZ2YVx4s1VaeCKloEZoiHXNiXtdvnzAB6WvU+1WtuPSeOempqDVUDm4
aU7toH9ci4gjbuahUwHsl6WV1EynuAqP/l1u80HT86fW9B++iMqDAFZ0sB3Tg079GWjSvX9MqAwE
uZkdd3OmN5xbzqYONrarXO5WdvXAy3mA9NowtkfRjJglMVwjtW9vSDaeFFUFTu0db3nUhd9ve+eE
YF89Bhz6ZvQWl2EvfIWf0htTv02QCx6mBxRkNA2LQaNP0N5l3aRiUIKoQoV5efYlQjL68InffCzh
V/psC3Mzj4/PCY71t4i08wDe7Cbt+qzeS/gD/XQl7xVH2t9pVkCuCGMM7DfrV7b13FLVE9G/OSPi
pPpGEz1VdHksZnrl9ccn+eFWzLYlbZjrk6gM8RtnOHnfz08NzzJqaS7+OGEBkKHEX5GD+x3HBuSC
3yIPZKXxDPYD8GuJxTtcPOUVmgG52Sd37yRIfNxzkKB4vGyswWbj54EIVOw2QclByL88En56tkgt
F/q/GdPuHVLifjs77j77WVgoTX+uRx5vzJCgU6uefMSTMdXgPd7QAjJDks9AIb7qFc4b7IRY/R7s
68OZl/lrlvcjPlBThzukrRchorZ6F5DIzTP71nyK3oTIcbJK+4vuZRMy9/XR8UPUhe/YO4HupOCP
wxDYo60qu9QWpaiSN6eQ67p/EbF8gbT78MFTrJgp6fB2v7wNsNXImiDWMh0KCfihrmzmzd8YOxFo
7Xt8teMjYykZkMhR/CdITquDzayVMqDgCo8TD8qJvXGW20b7JX6U3UnsEsx8i/qdrnfvpRbJ9QZC
62qvm9RdpzRFGAwU+Fe+U5uZYZDiPIu+GTa+pBpBhSrFHJdIiqpk2cDtdoP059bh8hyDwjzb6Csv
gsuIILHibjLk2HCBl9TMwIcO06HVOYTIJUnOiq+74+XFlUyt05ZWxGFZhO3be8HaKkykAi8D1RMf
lknKr0ZVNtFHa90Ar1OxHumFA1jDSU2TiKJtZPXqzuU17q+jr1076Tb/bP29Ro/ZyhNO9BmJJk7j
tE1Fv0m4TgXRiXtBtzK7FVb/3M5Md7b/KPsDfMIrs2asoq6tBHd8VSeB7bVLZy+RjKCzNM3vscTM
chguZzIgydKOtdWI5SNMyvnGE/J6UqUCHmkb+LNPvnrjyKxK/LbuReP0PhkUEcYpzSXrPWfu3S5X
xApxIXcEyVT7uFJv9sc8L5L2vwkrfJb1V0aK6H9Gn137SL+mdB/gZu7mGpedAAfNWtyYTrauynSi
U1GIu21EK5aXZQXYj2alNXgQ3cpApv9ZZUnNTB2RYi1c0kzwLEt42Q1VIyyqooPODjhu8Z2o4LZ7
sZ4O2AiFdHqGZPD5gHeOU1Di5b3iDZ5+ciuefdRG+RGEpnniqUTbfu3vORPSiFwrmVntqATkxv09
hB/P1YPtXpTKtVlpwPk4W3sw8EAW06AFT7qNbr9+yfNM2Gm1CXPmod9ihBN02hqZf7RNRP6bOJTR
Pn2BSMV+7/Vfw6FciJ3Gg371MJq7ra9hDPnWUp2AXvrfx3TUbUCFbpUKxTLlXNGS0x/lVHr0lMPG
Bn0IgjkfB4viOX5o/FYyat9q1mK0pRTH63ssJq6dBX+uhbU8bg4w442X5z4xA5MVuXeF4dBycnYU
y2+psg7vnJ9ibuI82G7gGmtnoy5E5GoeqxA8PpXZVoTwm++FmwbK3omgAVfZd5mrB8Inqf8Bxehb
Uj8NydqgYUifpYwRTdSxVEiwmWqbQVwOsl73pd2SawppEfggqwQ2FswpVjItT5B/8eZ+wgsTtlr9
a8i1mKYas+skP3rfF4oIH/ps3Uaun/iB+9CyI4QTedlNug4PPY1UALZTzAY+VtxUApnbtj0eAfA8
ZczzUuHZiQLSmC6svP1JelkFWjvGgxTNpligr00JVHWFvQvhTNCMogCOiwsB/6UE5m+92/u554Ix
ZfUElvNldbKh0CJX3K/r+E1DmCCQ9s5noo3817LZLsqzKMjY1TJUc7EcybQOmLpJhiDZYSbsfABA
oTaRtKndZmMlI1EaeUqTvRiyDzdzgO9e9lyrqGkyIKIz7o3jCYNgOT8I5X6QX7ljGiLaLXp9iqIx
5OI1sk66YsQgPfvAv+h24ED6yTOW7y30Mxb1nXe5fX9ULzEJv5OQVdjBQ3LM9cw80pk2MEAJE6gk
Oa4gaN9oJ4C/uPdWhjKcn4F/cVF4AMEPwUjGvE23Tl8vbpZMytNhDBPzmV4FEsf4tB9YbGY50HR3
EQ9iiYgPA+fCZes3coeknqxkt8jZj7pNHq07ijN+DE8ur8zMxu+mBIN1Z5dTnRKqvjFtsNZYtTTK
C271MO8Zkco9F2GE4t6g9gYzUBziMD9LDt9538wnT8mwotP7ynkMunFMtau3PEQ8rmXRLql0Jble
NDBL2Llc15FUQnkikzUUd4Mo48/1rkQetRSFOzkFgjCahEIb/rA77VKOpCDjJCCL+isHMxl8gYTX
+LDNSnI7BEoaHKD9ZrIQ9bLuKCDSZycF5rR3dUIE6xN0AlM/jH1X0uAgCKwP3yTWxH2znv6BzPB8
BMCw+Bz35QiF3RrO2HrHYxn6rHkk8SocAz4FOsGPeoquPhWMzXwH6BU292wNxUktKS8CRQN2V5y1
aOlJEIiEQCoHseyEjitarAbTto3nuWH64kapMNUQYcWTQHkzwa8yhcjVCnAVeCcoqZHGQ3J1rXVu
hjYdasaxxoX3IdBQj4DecbwoQQxkr1uTyxn+oBGRD26TyOf/Q58tFBoz7tKaHVhMrDTMxs+576km
ECd68T68l2EqLIgqZhtx96OVwhxdA2MklTAU+W/U5DdlzvHlRWEOZjfND+y0CkSUUjhH7P/Az1xc
5MVraZgw8x/7/lt9mb2IxMnQm55qWlOs5rS43TvjMZP1dapndnmoHZAhFmHtwsVRLl7HMBAlbWP1
BLqV97Fo9ArsQJ5X5QQXoCm9DhChe3G1X5R5s5xyqSnXcs0tb521T/50jXcZfYxKKTfheNcpjo8n
4zGXMdU6JoycesClKWDdKgxjcReuan6L2f4akj8k1fLGhsaBd/KijBS68gSPfxcrMTyqN0TajqDF
Df6Mibpnb7qj6LxhiM1TWYvwZUUwPBO1IRpefCRwTc5JDkyMtfcuJrnDlHEaeOkj+aWFUt6azRWN
lnCeOR5/YoXG617RGVb/vnOq3VKn61f7W79MdCWLGy0PSLKUIgllvED2A9iY0tAsl0jKqLpOroQc
ZSqJigLTLFrSZZKaPjsBL37HFtltpc9Ch4rNfif5GDZ0klbtYDySAbtNTp3SrFcWVBvDxwMfMN53
cqMwaMdJo5tMWI/2gfnXRDrSicClUHrcpL8aa6fHTEiVQXPjCzAqvNmEMhIUx+GYAJ0rgOM1KkD8
UUfZz8ceEcT9jlGcNf9opdL+wlXMeOWEUBFRXwkTV7NlyWbY5fGcBpsIvCJGXJd7QX0AlwXKUjUG
Sggu9GAnY3bhyYZAj5PR7WP4mNlX9NU2o9EXA0gkjXSPvBdh3XZrxTgYfwpmIlU9BAK3qT9/LNLO
A9MzPfPjagCAexjyAC/r1SxKGEvvyvOvJXFUjpbjqsh8AliF4pnohPqhLim8r7J+x7qhKzP4r2IP
bhzGIyxAmDkA5K+OD/nO4/Egf7Bmnr6N5vnPalG82Vv6SNk+2tfJmScngX144zpkNxB29VNVbFc7
vlIc2u+l7+ZXanhgy4EFHS3J6CAjWN+rtiHYKeDsUnQ8hcL+5M34q41lLfn6zFn9WMFsgFHlhMjX
HMmkI5gmRNvvgiHf4gaTH5nRE2DuZpt8sDk15DP5ZYVQ6WogVSDnUJzivSCRRx1J7nA+OEBVYwqM
Lrbont0y7hHlQliFiqkucKerasif5kIGllJ4JK8DEMo93UfInL4++oTvGNOJDpnmU2So5xANPaXm
xY9xwhtGKYYaq5HpdtCrNWqS1F5Nw2rmO2jpDA3TBc+k4ZOfahgg/4Y8pgBVOqVYScbGctL22X8J
j4kGz6CF+0BJIVfUWfv6HZYOuYmZFfS7TLsxpbKyUIiRB1TBIpFK/lyLBGInStOz13sVrXfAkO6A
rPAClArnstq7ewqd1gdKFAtsSVHAe9i3053gB4F1GWmDyWkxcg625cF88Gqy0JB49gCJZATTp54Q
7twN6FxHL0+K09ZvcOPCDeW1LpT3gJi0g5F4RG4GpjkXlfUxcCQmf4h0ZjS3tHfTF4AZXbBFsnUX
Ug9dH7rjY613Am6vHs/RwJypKWXPsssPnjrC9SxbP7CJeZKe8dQg2xJp9OLQDsMWRJrKjNw38Ucr
/1HWl9PqeYl7tHNQHq/jXYQmjQPsY2MWa4TS9AhmzOcPrDm5LuzUo/fQxdOsZzkb1ttvhx+CgJJc
ZYdwvxAEuQsRpc9PVen0GE1bz7nD1Ls20JFaqaOG+KTAmF5+TgeBLO4mZzqVJs1xf7LqrLAwZPiK
NTV0OeaIXod+q51zToCaWLp+iq2GazTd5YYE/2E7VmHmyg7NpWOqwrj59/bydcoV2uot+3Jm6/eY
CZmcvxmbLVjzscMoC+6b9/lCcm3AXqGf4Fa8VFmtUFlRqasup6P7cYzs1/G7nMmybihlGtdlzUMt
7rShX+MpDejIbrM55SCqrqa3tShSarJLLb3edBS6ir/WqTbe6FMgPYBxGqEAtiraOOyXc3M25pD5
IhyRSBCi41IJzh9K2YFjUu7YWR0vuGVdTwdZs75MA/tC61yhSgfH6Rmuq5xEnTEMf84KzjGLaFfV
hh1pK7lqSGHR+T7z5GyHa6tYtrFfHdYDx5c1yyGp+QVDLyQfPFQoktip6NGXHGqHqex8GbuNQLTS
OFpfUHCDa98P8xTWHkf9NbPNYrZt1lkKFfEsrABUoNsiZmm5ItRfn7lTE1mw0y3d3g3TK97PiWvk
q3WZnGT8R9xQOZGOhOKMLWnhKmGxM4F8l3PVavS2iaFOYhtzMbpX6dg3Ve++AlfnTQAp022FRtx0
Uwp3/WKHiFkk2VhQHLHRCDXRZ4RKslREk6teXYFMHH6lbkO7BdOWALO2TZvIOBrLYOM3FVijm+gB
Y9YvDIwrYOZvYt8JoyO208imSCznL0wvnuH9Vk6K8EkBL/VfzblmYLwTihEc9rMkZlXNHPGpf2bb
j0+ZT1qyA5s5wlpJ9b01MJpJM9aYMujPqkSOqVKGJCivWYED2ThnuhamL4XIZN216j/xjX+snShY
+vgjvFHQT1bfGKunKr0IHQsL2o7pAMPmTSrINHeI8VeTWGS0NCzAlBmVSsKwlkRtTpXChyyE6gZZ
8KOcmzWNdVnNgxTAvWm8PNLnHHtz1UmttrI16+5/idLWpeUCjaUC60DLX/CHnQXhSzZLNOj28Zqm
hv2MYqxzSfn/Y89LW5Cbqief5RUPz4Rex6iumpcq+9ZIv4gLmxTR4+fnm23KankrAQ5l51PTgkH+
25RyUVuM64yr5narcx4eerXDai607eRwKKs/tmB73Bzlg13zGMQmPopryXXg+FZwilzyLr2ByREI
KBV/dnkhOxeFzlDbTCOc7GQQ3bvcf3nLcM8qu1GV/NtohMuc3Cs0uDABChWGwaoa3zk1lwsS3JpH
SHveVnWAofeRiIiCZ4R5MXRWMzq5sZyxImQlQvF7IvWEtl8g295zooqt8P5NfOVJQ18nUJy6tBD1
dJbOT7LemqX0e35FSpPEQ+aNCaSPHLVjGsyjBA/P6zRX8uOK+t9lwYrL2Ldt36DgNZBBdCZoevIn
Fo9m8O/a5cDo+WWavqiIzky8MDH9XZzI1q5H++lBYqsvX7XQnaHDLNhUlxLHw2JPv22A2JRrW7eS
BmKikTQEbi3KCZj00zJr2EtpwH9soB97xCxCwcaa6NgW7lIwp1In/pVIBsPBH2vdE622SHUfKhLF
UC/UoFm7Z/cWZMWMhogYHU7UcEJIuWPG4h7Nlnpd7LRD20hKvHaV9LZI4n0o1VXtciDhw1v10UmT
vJk8UAqZWfO7tO8bj1fqyl4jIoL/mzKLbw67GA9orR7x+6mHYtC1OQfnECYambI8zdkv8r1YRu8U
lSj7uEmaeLXqHFynZA9HNF0IWXSMhIfHJtOv54Yx/VSCTJy4WjZrwAT0HLnrGZ7eOJcQb9nseMFM
5RdD+9oWfGn3q65IvsSp+QQ/sG9KmgsqR3um7KA6J+S9y+HJQzHZj0vYBjf1z4szYbsNABbIiicc
EXWNY9N6r9zi986Ij30tCOl3XXBuXyKcUNoiBXZNTSJrGlEFVj1o9cdz/IWjuYeUNatyaUElRNFi
MA07fYYxltr+r/UD7Pqr4/iHpZkbiCu5apzQZWWsxRefJhlwxeAp+AvJrhbuS08kS9AHJdEJQfJl
oVigkmWOm1MfZxq1szpjFVfCRS+78x+NYaM842hWdiqbdB2DOZp9h0w/fhu0wjgIh8hj+vXw/M86
LbzjDfvaiq1sbfg86JtK+D7g0NGHePX5IXIpTsNKsmPv9Wr9BZVE9UUUqM6WzW/HZA7XY1Nzd9BR
fuGWRZ19ARTcVdJccD0Vd3Ium54zMG5ZcLp3IqdfZX6sKemxNEAcHVhjABRDflUtr+gLgH7DTIRX
y1uvrm5iSnniEIiTI0ANhB5l/vicanDoIa5eRG4arvhUl/6hBgshUTv04F/9q8bwFYqdQVOdBR0n
/bBKserfoxd5AhZ8fX9s6a9ZLtMAjfuiweg8jmVI+lIlb/mWkKmbxZzr6KRPmCPzNGGuwEoQxA6A
sdiz8IiPR9op2baHI/9zK+Tsq59jtA9cayoKrjTAZZmBjyfZYrtDG9z2YNLUM3QZ2rV/JZotn+m5
IyaLH1Ax6MQkOiWNtaWkjYtLwb44v05Wg+5Wf4GaHeU/XF0hGtewHn8bIrCF8xLYq4ky7+5N8O+O
4eYV6psNniwqX8g0QH62rYuvVBH1f7LPjqkraFxuf7hCIMksmYgCs0rAmlyudn8uk6iXlpTIgPIY
ihvVAzmyIgGS592XZ5q59pl1KYervx8Wlc+IDYrlIfOI7xUTajyJGfrM6E7kfNuyKuMrIq0iUypF
nCfg/Uf4ipfi9aGPpmD7U5P2E+xlWwGDCU73wI2yj2AshQGPM3zJcKlLjM/b/DODsMRw3M1QbOpA
h1oHaSYv1uUVJ2VHXcEpRC4e5fy3E9FH6rfr6xmx2i5AtwM28oSCwlAvWB+HCvd87oWkcxC/8kPZ
5S+rz4NMnWoHKvKu8mMoNWrZx055nIIHCUwSDAwBfNwYUEdUi94xpBT5N324RgN0hpAX2qtRhoay
l8Bls+GhRd3c2+UVWzz9jdc1d75bDghlLpnxbd6wFhzo0wE6sfgGmQEhVUdRoqyCAvXi5qrsR9OU
91hjvPNcgvMDcom03IzTzh9AXdAERxzkMDVOKOCOi19zBAIcpUijb6u5fjiHXRxRSVdG1dtXFuZx
i0Uqd8bJIO3vZ5Wtb8OrLWvVdvgD0Ilp+2LUUHXMt/6xoLoHYFq+mzVqnK9vtvz2lRQ8Bs2+llv+
8XIp0utbfTaPbKWJX3qzORh1I0uBKz1Fhx4RexgnUExo9DJhu0gYUSK2UOWaB9paA6TRWLuv1MrH
jxS2/9gV5SLkfWPzkU3bqL1PYBJxlEperfdPVKKj3GnT5db6yQrMIbmoQbgFmQdebfQIy9q0geR1
FRtP3luPHAjyCygm1jZeGAtTJoIKAvDWXkIICz1ijiz6l8sWj6XFjvhczCufom6vh0mNjy8l+tRw
MAoItjpc3hqWdHeUv1LYC70kFDvUpGsbsxSe0TdxRt4LqL1uTXvyCVzVyc17zxGNA4Pht3Uirr5T
yUKkotyEJkbhSWxWgAOq11V2VhKE07BviicYIrZauq5umadhrh4/dwrO2dJ0V/rOilze3m/SV5Nk
6g74vhXGDBK1JlXFvCxy2rdQMRMvyWJytDcW8QerVPR32IaDzV5BxtpCj75meY4AXLr9FAfLznAz
MGMCl6x63gBdB6EttyIcGKnWppzxk35FYz47r5FM/eEFE97m7MEMiGKRcwjvOvQXX+g/e72lJYaX
iLPTC2E/ePub19GyjYp03D/wnMT8HwBk0t9Bf41mzr80pak2fIXJNOsd6Au5DIixHE/35WIry7ed
KINfOsL6HctLLH1DtWdgRG9DlVGAfsvYckhvzuUfEYIEg6a/0BkeBGRdJXWFgCtBoKyuI1Eur4db
IDCgSlKPqTnhT/eWdleVqmBtw+e2wxkO8Jv/2aCsOJW/L87GKfCToIOpfsKfGGFqDV3Kz7P0OxiJ
tQlgcCJ2/qhRINlEMDGEoYlIVfdL71qq1ljA6Y+6REYgRoZYk3sAVFC11gBz04+TiZ/ulXJjYksQ
tSBOATPAq3q61NrdyF9IaHlVWOKsKGsyHdvVYdLTjK7vkifep+uE0HNI6i5MOUhbV5U8f8aV8y+E
/dK7UkUYvygk2bfsyIKJcILcvCg7sPRQXodQGp4n82TelBoOwF73VO2JPusYFem0HOUxYlYUe1yn
0m5p15Mj4WuhvBa2sL4Nx5Eu+KdfkkCHDpiHtoPtoupcdxdyqxhGKDyV1uG5VC08vcwDBepBm1Op
jVMFsautYhqvmnZO3PQaZ1IWx7cyc/AD7j3OCfXn+T3chs9YttZPgnr24hcASBYRF+rmZGkdeMt4
uUBoeXsHr2uLNXRLO5AO4n9JliCoZIHcDNpXSmFTbr83iNpMG0w8YOgiL2Z4+S4CaZZkzT1TfJeh
ektQ3qPMZSGCXKVucEh/h0jj41RrU6WDgmmQGCbI4jYZb2JRZ9Z+t7bsQCURRvM1BMh+yjDgLpmi
DCPTSVhKeRcAUhWfv1tu57FQJIHxp04kXs7D9A9b+DVmaLgW5t9AAlc2Kst3v/WpqJVVTmb9mNUC
b8StaHOtr6ZAGFz5pvHtoAVK/JUxt6rhKuEvncE2KXHX6FNFG71rf3vIptm9KBr5LqRMWI9iCDh7
+2830tehQdopVoSy6W5p+v8+Eff6GVHaJbbpO/cjduiF4ba+5F50eRtnRxjYAO17WGHecZoknIPw
q0m9lWIqXGz94/n9PvKZETuLFs1F5BWv2f4vpzkykyE4tNPYNQ+ngTO8nrhLqyvbvXXaxQLypc1u
lGqJePQGWN2g1h4x1GcH/SQLyCbml+zhLIImo7bekEChSUlltlDKp8g5ylnLcqL/sQbF/SVsztQW
R3hwr/pDm34oFN4In8+nmLQVb2ytwJL5hzDNwQgGj4wQgzCF5CR+I8vbzWPTSpu1K1WSMIEdI+GB
YorPhQAzNeLoKaRjgHOxczz1fXDf9T089KOOHCQtYl4r0qf/anwVuqy0+xJqAu7ox1WQtsJjJtzU
UWkAb3mJCPICaOkY7uxZi23/zcKjZRi9Ns6PUEC4cIpGcOTcXuxswcYWSsu96Fki60rpViFVLhbw
eQl2rrAMnkkmMc5KhV4siShC91U441A4yXnKBtdP+6HchQzpvEgcc8dMT+f2To4R71E7nJfnZbT2
fK6d6WDWzzVgHPuNNxBHr+t7sGYdVp+cC0JMTwny0drHKJRMWt2wkqU0eGk6SSA6WkTUU+kVl+0n
6EXYUvAMwvltpI5bZreJMN+WFuyPd2iYU+wCzTsrvewe6hOQTdKYh8j7ZXROFhb1O9c3XSHcTdJw
JANIKG+AdCgSY8lKZfDFgiysF5nOmEMdGl6xsTB2MyW8qKrFUoQBBE5KwlUcIwfXl0HEbcikSFIV
9IBOs23a6cV2goT4hLQsk8JmjJUzgphkX2f6d5IMZAgq+8/E5oCPt0A0uOab6DdA2qu33wXmp30N
MRyr0tWf4PtRR8DRTXIdjTQ0BFRAo+6crOePrscK2AJlaytGXgoSil5+5rRBetQPtED8ZONbM/Wr
Sc7akzAAg6Om0+YdYjWlrzed5VNfq3Q5YZSjnf2nVnk3RIo1QEMbtTplUymT5wy6Goa9Sa2JWWXf
sSI0VsSSrBhRBnwEkyZLcuEFafNlXgOTFQsQApL4QOCR/KnF2acFdyU6o3Jqp41dTokx2zf+mWyN
CKaGdTp40tCcNH+nDlM9AIcifwxJcjJI4nKD1vzs4U//ktsHp3EVAC9qzw9uhFoZa4vaf+/JeHIs
cHME0Y9tr8NYxLH4scMFO6x2OxANsii5pRe5iefCOpXsSBX4U6lgGdjGQRUN8g89/OljrjoOH7rl
g93rHRDgYq9MhhnyUS5wTdCbnCw/sLJMtDeINA5aaakSi4z0hEjTRPbqDGvshDxrmurxMGdSf+Hq
E6Jo46DlrjhBTlaSiYV2WMLMgmhmF1hnS9Mioj1c0cXWYMN74MWKED8u91dbc2NmgNBSKkJwJnea
/V9CQMBrXVxtE8R+Tljo9TxsrZtr5AhUdtwJek/Nauahwyrwi2F8lN1oOYu5BXoc+0whgx0uNpQ8
RLre4xxYqbAPF4tfGi3JokvICKCX0QjnrG88Xs4elZs9zdT0C1vCzW58as/g/O/A4jsYEa4jeA9d
FGDG3C3zpGnRvbt3AXb3ZyWsrPcaTvhx6vMk7ycbQNw+W6moPmphCEQF5WeDOnZrTDR7x1f3ViRM
FQll/g16KGuP7h/RJ887yIvkXeIex220wPeN8Rvhp4phIUI+YdQJ8MXcQP5C5Le5vW2rWwrEqN13
g3nZ25WV0g3lMMfOB0qpMy+7RCE6kIFZKQ9ld8gCfnKPDjoG38sU4Y5N6l2J8D5ub70LY/jIg3VB
K8A5M6rYo6Lxbs5fFFhLnoAAoXLfBvWE0BBuuFPmvfJLVdVwhFTULdkHV2alGkKlS6rHRP/jyDii
TkVnhfTs2NjUd54CoPj/putVKhVtmtDBJHtNQ1FZklkF8lIE/c1fYMZ9k2PObR/t3kzlpTmWz5+Q
rKGUcSYg6A6WJ7NR4OyDl8mVJ2BBZIeTmoiRGJ+raVHSk8YyrHZNoseBcn5aD3fFtgmZUP6eZv0T
R2ujJgNmmV/KQ45FDZJBEkYzkgflNkUWNic3W++Eoqr2YQ2D8CINaDlBzoHXQY2pjRcbDFgbqlmD
9xI9n9k1SiuoqZxk+crv55CILoXvg3GvwkG59zyz5zpG34Q7aJh7AVQU0/MFGuvr7UwjNM/lbb3T
5Xd0EFG4Oo41SENi1B0pEHRPpfTcyug24hVoFPjKz3h9n5QvjTWaSvoXjinM74WpttkGuEEInn37
h2BApiZot3lp95m5mWT7xvQIFd6MVFg5qbrdHqMeuXJ9TSu9UQOOyEFDP8rYqa0V7BknyNJXcwem
dLAf80dvmFA2Dpyoo3T3Ed2LgIOVcIuUjysVwiW1BHClCHhwYkDa/uld/jBXtiCKgqGgXbrseKQM
9tRGjSzo3O5Z0hp0QbYhyYPBRncYN2xYQjliwEBLloQjAfwzQ+XPfjDH9pR/6hmXnAb73wbqFpUT
CrHdG/7TjXgV0ICR2pLeXOE5H6jYF/XtFMZWBPw9FLG2B2diYAkzi/ZWCRpn+nFc7rqg4AykBpW8
vSjSQ5Yexg2ZNXSlNV1yOq5c0zBA2GJZrh78864za05LYzlwW0sbRMDgtYKZJw7tTnQ9UWDQxPUY
NEgY+1i2IzFxlkJ69yUijMU2dz9sldesQpdT8UQM4FSYs5laPbS4ivZ0m1AW6o0rcUCrcGaqOtoX
j3bz62bwRncldtY+wnFk3pkbwZnLKSPlpiqg/Szxzaf648VFPEkmX6zJLzFdu8MpmpxFaTeFebRV
BH/mQQJKEcLdCENf9eSxlSN/WscmeZ09qCf95VnketP6pvu40sxMqvmWWdiGM3zJQD81anV+eI1q
BCYxkByBarfSV6m175g9CKinm8gMcZZRtbCQ+qYHVGW/hxTku/HtZ36I0Gc0gEXpdiS1YRSpRGiY
x4ZzHAyE3NBMDQO0QduWyB+zOXnc9uDd56UXELK9w+mNn8ly414y+6XRz4E/SVNdiyP79Kx728FB
yGiqip85x2X8hjBTfq4XVAdEuALACpEtr38KoCBHNZnCmrQOQ4NI466lu0VqxHrU2Ui2emNFZHq5
SenhStSuv74M/MZtCRmH+9a+aTcVNYIxomJ1UQpORbrQFuh3W9LGBGWJdggcoKz+b7Vm6Y2Ljt6q
Wx9ehD+e72Jx5hFq42F4ACDLVK0TqqAhe11Fhi9GzJ3rNexUSGO9/sd5p2VjIxOKQWPxwybohbYU
WxdapGtenkoRbf42GXq7HJw7IdezPzttys9M7cd3rqdFwgNoJVKngK27DJ/N5FSq/2+UOe4Ip3zf
esXRKQnlPa7CPon+dp/tOb2JEyCopkY62L6DttNN3wyGMpzRjhd35SyctracEB/Q1y0LMOrpj5FP
mj0K6yazMQg3I4uhWvfbalcux4/9Ow4A9jCz2T47AnMY9fPxd+Qx1jO2vebqzniqCOsCxD71CVkQ
DKxaGCkTYUceWFqT4Z1c2bgP0H5CfPPidddoGOUIwc178t4uRTN0WzDD7iJK2+ty3P8DU4P4YVsL
JeMk7lfaF1K1ZKASIIvG1ap7Uio44bkS+Qgu6MiSRRXr++1pXAjqarNAX2lSF9zImx4AhX0aPa86
01d08r46+G0/2pIwzOlwxIJYU54eJGwIIczg0Lzq29dNmK5aM5E0Dd8H6j258hBV85Lyna4CEjDp
Fs+W4281wBOdfz0YpwP76XEbaJEG0+nqtVMVkCs1HkxRvTiXrUix5h1AKwWsRStuWfTrer7Xf83P
Txw8d8Q0F9/xazOkDKWgn0IBpWTUv4oNvP8rZSb2o1XVrJOQOZiTzQl2lI12iUzI+MGwBslJ6c2Y
lSrwVatRQUBfzfhJa79nXWdhwZ+uXFjVgpdMo9leAGe5q9m0lRaBp0iaLy66vmfq6HbZmP61ULjH
7k11WTpHvoO8r8uYs38lVWgGaxb87TZQucZu1E96i5gDzU3AzF9ee5uz8TE1oow3F+feMpkbTlWi
BeeWa2qONun2bS1b4X4elxR54CLBie41LXvKF29MIC8TFnxMzBcOhztucSntorcQuhv5tuHBEJYd
hmMTrlWbYogLh6aNUMm1w+HyEXlQg31UDtA7mCjSUVhpy9dF4ZJ7Yl5jrSdA+AOXjsfR69EpPH2i
R+4xU2+TzXFWfTLxDG1FV9Ixr76iib32r0JH3g+hxtHgttz4pVfvXUXUvt26FujRKqwSBA5iQRxk
ApJp66E8QGN+nCjOuwaVfKf1Uxp59X3NjAVD4BjPzfPTyx+w0HNyxJY67kATY2bHUVJR5VcJeg16
YYL1BIypeeG95kHkFcDEpf1aTivj7nmE3NWqDDNPgh0QViGwWX3gC1jbewv8JPApyyNpVA2HDEiP
P35E0p3CIChC/Ef/2WY9uYnaVDLhD0PbxdC4DEOyfWIc73x9ZXXfUiwS2xBnyB7CP7y2W1VpE/zx
3OLCL+ynskRPS0Hz4qU30nb7MSYQ3/hhYH1drkI3Fj1CTVotDRNCPjf4iEfwL7pbozCf3+Yof7/C
hkCayHVdioVFdBQ9H0X4yYtmuxFeDjknPXXh7WflRkSip+swsxl0N7CGwUislfAMGMUc8NEOTMcF
5bOZM/26OMxAjRmjw3f0Sbic7ou41LTAC5CRmY6HoGJQDc6jTHhgwxl7YL4vxKeYO3PLzBHo+A9x
+JnfddIdKwxLF0hETJHJP/MjKqGAnTPHp6aSwCGRRVFAfVF32hENWIVs6rydX0dFvQWC2QsD/+Mg
lczjM/PdCZKT47jXLs1Dmsb4rpg5IonhTzoKBO0YuesGliX4EDplIHf+Em3b4B41nOT8LQ3JUyPs
7ogUxEoc7tyqPTWp78ntHs55HgsrXiHtGTWT5bwS9BSvzhn/qP7Sa9GLivLfDm4vRakKlANhTFzJ
XhsoDLLWd+Imq3lRT2lEszCr/cnUFC3bpAEk+ljkF3WIY/i+y5HWsfDPIdGwQ6Gc0zxc0QL29cxm
ADr8O7VKl7RbIxv4oq75JEdBuClWNWtmSFoiDvvppW7O24xShbO3NBAg/gWSjwTP8j5Oz1tu+Uur
wZZvK0jprhwMZU7m3gdLYNGzL6fd7j+ZKmBFx3G+ux2Sl+USBdKwXil1tmFodV5TAi5jp7ssjYP0
CfKd9wpKiEO2kyR+b/0RNSWNwvheBf33dZ86eD3M7Gu5W0LU65JcLnOwXtSj2qxaEFPK9XqnCqS0
AJRAinMhJU1URUcE/KmPuatRu4m8zHpnkE7817xKZGbePgZP985HuPpA8Wn1rWonurbEuUqLByR6
2ClUXETSXysshaPwJ3TMY/jCmu1aPlIqXcI6gH9dSNYGAUuMmDP71KUGYFhLEwOehBChkOfxoOjR
01wJG7+QfK3Rsydyn3hYkSvZ93B7whfYsewEV5Mpj80U7ismirgXMqULMhCEykmpkV0CZ47iVQ+z
5TcRH6ZKsHzf83o56WSUd3A0LMiioQSM8PmMi8rEi1Iq0e2sarYeSAke+tCZuqApqUUo5PyMQB5p
jbbV5cRMft4GTQu6gZgx0GDuZ9BHLKiHCzeaaxD85Ka9h1aEHaRxkSb67if3qisnrIavbtYO2Svw
+tNFIMkKFndYDv1CgQv4/z0+Hd/Eoa7OxBGC4cq1SU/1C2/zf/MJmiU+1RpZVQQQmvtbtuKJ3rWb
iSAGuZsaD5ulISKnzbuGYmd4ortNgIqvX6oQaqRN+ctUzjxX/e7S+JdrR3p7ZtwIQQ+M10z4skr1
fa3yUhQ0TguSfZVP2+wqWB0PqUSu3mizKDNfreF1ye3FLoaVIcnfhjDsnWfHecG9ebbfe5quJlvI
K/H7RG2YSnwH4GvcK3jI89Ezmg6EuJyiY8yfpxLmUWGjqDyRJDtQLi+GKcMoohUOZjWnkvx1D7ym
k5ZGLTDBImQiwumBhL7uas1s9PcOJQpHtPqvoevq8huvdc/49nSzXO+4ux5KP3zSSsBmEGtXNH/T
64fBh3xTKZEJbY7UnyS+irFxVC/b0hHOqZOmk4jR/p9drtjxG0z4H0Dds1jKfPcM2xriW8Ka/Xqm
l3p4u8fMzqRJuWgD0JqcoKsFczkjxsyPQrN3i8j0CeaT1BhrMwbcAtCrTg1UFrG66MrhgAJ2heW0
u6U31q33YoNSz/vAdVspj4fJt3YjUuQ7FlRLoQAKJ3X0fP0q65pGWU7CThwP/psAa3o2rvR4Hp3B
yMKxlklP0ePPFozzoASeMBxoZFXIW27TVaIHsOrbgg2aPB/Q/O3FUbKQqVA4lqdzXfZHUZuBtD2J
/6EiQVMQozH2T9PUTteXjUXsQGE5f+z/aTZjF5Ux2uvgvGGG+b4vSKEILYORbt/uGpkqgDVEvRUJ
O5v8h4sQlQytkxS5tKlnjmDjhME1NF6ydlM4WPFJ0jQlLoKMWW7is7kJ4c/ktq3UNwRnjLNi0Wq/
o0n86oRKjO2DOlHruKVYstD3YSC65yq6jdDN/lmhsEtJYxbQeQNbxPH9AzfS6y1/EcTTzGvQruc2
PXnGVkJ3cqrUeEFlMw1pHyfnDoq8LAGH8VaIvDWDkIbp/Q43gUT+W92nH9desVXhrP0PHSAVt4t1
pzIqOPufI/+lgGEZD0qj/9AU+Is5QWmbYQ+5GEChhRt1rga/6lBPneCpqZbxl4m1o/w3fZS2ZP8I
YSlYeptw2jxcsN2PgCmvIF8HqRi35XbYWITH22i+dGEgtdpUtoP5j6EVkGmtrO+HDX9AkAZ/ZDUF
Wbb5qA2+RyEIRJqxK/Vw0ycltgF3COWgsLRDyc1mUd/YBfylswQSIDSIiiXymPoczwC+rioaprza
PrpPj690qza/5eRxZxIMJA3GhxoOg8kprgui0GJvhodCUYax3SgLf0bQ4RISCL+63CY5kzw4F+sh
ukLwbcPCWuC8Hn2B7B2ovG7zB3VxY2hNKUvsKI2aqPUIgAoY7s12z4BWsa8h82eOEE1/xGlkbtGn
nYgBxAovGGneU8XmPuCBm3wpixga6oVnsP5aLG6C26kldxfbU1TYp5XGQ0SoEE7gjrefnoFv8L2f
mCGufWA0vHrms/2O/PM/wMsV2rEt0rZ+wAMwnm7OrmIL1/OwcJtJ+hD9Le1NHVwcaiS7zaHm3CDq
x4J2gGTl3Fv3uEMXDJyiERmNQwCFNAn7YSgLUDqEHhjjnHXpGcNbvFUbFUxZeXINewTxfBoXkPv5
crg5q9EzrvbJjHa43sKkwsJBIrcdon4xerw+OQLA2ku1h2QWOo7UASVNHr4cajOaQ49lg0YkMSPd
al0U+zCzXTIjrOx297MkGA4rEaKqOjRv0spwqlrmBF6+TTfBAD1YtDZdkhAISnzQwuXCJ7Ub6Z6N
LvFLUYyElhVL+x87bUDp5xo9a53L1DYWyjCbtJY1z9xAwX2yIwtyuevO9u4NdTMvNbX/9g9uZbWJ
qIr7+k2ed1lyWbeS7u+nk+jDULLDoGeTrvVMNOTgb5pEfrBjw8nP3EIA0osi4KjAKvgaddbExOJA
YA9MliTXazcd2BHHl95E8UDffX31VktVXtM1sod0NpQx1f7PwWsx50TGEJ7C7CjmpmPYa4vRkHvG
G+at8w1JipoqB6anoP83FrWwkGPISXTlElBROxtGtZGTtLUXWgk/zce/j2uDXThMJ3TDgGwcMDUe
VUiSCSW0vz+cCtXQCJuXau70hvj0RlPClXO52npxI72pT+T5CKOydLBkoou2bC6/FDl6NvcnPE1+
CzPtN+2wOy5SmeKUV0WsXayvJO+LIxk4NTBc0fWkApmJVs3TDOiOfhzKsAI7WyOo/MlI1Ek3TEUM
yCJ/xnmljjMSpjZDRdgsXyvI/xT6l3B0Kg/C4f/rm3Jvx41qU1agaxgLyjir2/jJ9CfKmw6YWhaS
Y+QT1VjlSLxb1soVGAlh/+/N+segf9e0PuqVWpuvV1j3Fhmzeyk0qDU/ArpjCrmcvPN5dk2c9J8A
mV+61jywVKTfhFLgCe3TP77VM6of5KMi1fUo80dJlfTRv0pG842CJzOQbjmCl/gDwGwB64XZVVVO
KqFv0jh5OWZgGrdr8Ewj4a730g5QFFeVPEaG4FcKv9Du5aTpu3tOUEo2XBOm5U2lJ9A7rWE3AAgP
shrjzwYuSppwieI7hvQBNiMZU7RBlHpQypNhWvWZIDGs7xldb1qRZuweVIebN/sWzf1XMzO6SJXH
5mMC1m2H64E6DrW6gJozVwzZYQIfyK1QGA9m5QrVHBRL4+t8+hgAFs3c6v3U013DIsHPXM//eTOt
UTfstCoK+pJh1ZfzgGGgVg8+h4c8RuSjb66VBgdcpDrAPRbKVEiD6O4eTuLl59c9GhS1k52jB5fg
oNCOr0OSKVwjsDeSy4dI+QbSj30bk5zEBrpuN5+MXACjEsPAriYibYl/RnRQxOiVK3DgOHhxS5jM
8cPov53GDe/4pmXB4fN2c3Fjp7agf1REr0qQrzKkHpbYEj7STjlIQwems9kGq6ZDM4M6JFaCywlL
6ypdyG5YUb4q+T2MZR+PrBGAI8yqAkVUM8ok+S4vmkFqzIs1QZZ1+yQcwJUnfYnIg+zAtz/f7TpJ
MKrT/nsL5KKFnI8nRTI3XAoFt1NA22KDqRiwgz7QUxEJgNMMUdwDSFBEgJkU9fTWWvnBxZifOAeJ
Tj/1bEDwEvD6Mr57wx+CtlgA9OBf5dwanNZLK6oz0aLU9U/KyFQHAeWFmb1xtPOYv7MvVfJ7pECh
95Ch+j/recMU6Kq5X4butpShNmyKqkW/LUCHVHYgsmXmD5oLZuRjjRBFpVyGOSfZD7frIjCKK0y2
iDrf5VV+ca09voYijgZVQBr4gQjQ8ZAjDUPPDs2tUDTaf/wokm0FHuUTEFI5mgK7tONrg89bIqzz
W13Jh1mmMV7q2STxIBMuTdYeNkHnwdgE5x/PkLUw+RR3Za8mg9i5VjJAdlMSrsVw+8BnjzFJnG4S
/g810bkSpRkk6FWssCJnpwB7k7Sws88ZS6vozWetlAimncmYvCqcTT8JrOC5CyvOH42QFVoOJ/Sw
4wrj/SibJ/jxkKJVGcSNuMhTwypmTE4C3NOs2DqiiDzDD3hGxlhDMNLiuqe3/lmHpAD5Cf97cTtE
c21eJK3QXbbIYQTX77Lt6E6SZUJhlqPMFpWI9CcFDQ96+UwH0FofClZ6berfeXSgQscWf8v3M+lR
//8qK8/AZqedYiTCYwzTOs3uXgd8B4G9ntOrhQgHBCOemVpq341hd1SevyeP1WxF7couxb2QoD2l
S3evVA4DqzrXec9l1i7ueZVz821AmVp6/kZB10ksauGYzyA917+UxlLcX/ZfBofYs2AaKARl94c+
dPdmFyLvJPiTDGM7NBhleqJTcIb1OoheWabDOo8GuKI6e7SrHoi7/g/ECVDXPXPOOznj8w4u/mlx
639+YNgpQg3aLX/Rsath4R5Z/H5hXX0sT4vRjrNXe4q2kkxpwxazMxsZZVcH4NSeg9fblx3mu9So
4FVuYDk82sz25Z0aLheu6Cim3Gx3rd/OH0fCEUof1uj1T4D/jYvCAXRz3PzSHXMWciX0QHoz8MFo
Nn2dli/yvqWfd6lRylL1+DCauOU+1hkz/snlEg5+bVQ7/xZU9D3xaVdFyxUaeTcdGCCMFSVT3zJj
wpScdbVvyGXXzk4CZGE5gAgf+CovItTFpnxoKXBoUMO6lKB0EN2mg2JADAqcakC0CSqfUesn409b
4Rc6D422Glj6sX2HOTbDNPP2x+NGyxKpXgCFyGGn9Zt5D0SfxI4xrXemzCpE4F440IrunutkDxRw
h273u06LZCNkmVzZANYNK4Fjdj6LoBq95zuDIIyvmjHstOL8DHCZTCtmZqGRn3ocAOhit9UrkFJg
4IPFJbONPnY/hHt153em/BXFIvapMZOXdBmkBP4dI2Cno42gEUbBFyUDxqfaeq7zZVOdCGKlgWYH
W7i05KHNUQVP4iE/bs8yzP7aHT6iAeUBxHdSfCaB0ANuXK96ZFLPCnsXtFEFSdZjBmdd2zcRrgl/
O5pzBlqWEul807sKc48SkiXnXQQzmZyt9abs0p64zWweYMAL0TRjyBKNzDGKsUDa+pRCSnfxnPCK
zuJHyzIVNvO9KCEk3hPBLgKx2YTyKu1pgjmK6su4biU2RrYtOPLxHytLevzY/o7o/8tksf6tEGAb
YSiX2dZpbR90fqoj6BMKxw9r+ACZHNttHuFbeJtQdJnXrg/8VntemwxYhiNEgHjtud5+LdPDotNK
V3L7nso5kFSJsvXvupW21ya8THeGv/mJk+KOcJiRI428KhUkWuQ23aC2nYHJWWWuQDMZyXr8yz0R
scH0bnUyvxzZdJ3b5ktFdv5RTcHsPuryhgHtQZstLNr00/JwnM0dvvR/mp6XiPIFLCvAH8zDalSZ
+vzNnELYTzQecjEd7Op8zVBJbpgtxvXkcl2qRqiSA/kP52+tjfYA903p/cmrGuCQ2KdafZVVPVLg
vF6+Ml6XJMmJ8ix2PwdDwgzHPB0MW51mrxSIK4QOz+kvgD901k6mvBSXc7a57n51cenTDIs4IoHc
W5r4/8KKjjdJOWlRIdO7ef6C0XHahLnbmkr4ZHZAhDtO+P5Au8wf0rFqgj8kUYvbRJaMkIjWCm+Y
hv68yv9Hy+8CgODiVzXaERFadb+T2kh8NcUJ1oCyWz/q79G91CUjYGTh6ijz4knuFhlkFqR0X0nK
FFZeIrWdhJCqw+XICXX2bgW8gcViI/fzUSIdiOmMPMndaHqFxcn6SMlzZg6AXMNTbDAxFKPFkOAG
xz2vIMQSS3xgE531LHHvouNCG1YPK2YoOuppPYNSRoA+wJncQrt3tqK7F+9FxF+ybZx5wBn8ISIz
5E0vG00mr7EIjenw2xnzAYyux73C67/BI0Q0psrALrf/6D5tdO9s673dhz29GMkRWt0Ny+/czLUR
AP6HosevfMTrPyROjyKRXK33sebCqeFM8bPPu7eJwrgx4AnwFk8TbtZv4Fk54O7AQByQK/M71PO0
QSnXEziIAyr9FCEKE9p2qOrXHGy1nj6xN/cHMEzV8ucHil1YxfPNTesJfLvFJ3pCqBxMFUvDJ+wl
EJ10bKnfv7NTTgqEvZXtW92i5I0hB2Gpo4ofHlmc8G+8L7Tg3rMphljNZwH2hEtyuF3v7P8xkpBK
jfIf9c1LArenOJAHrgZVJpZM74CecXWYEU9ZZ+JkRxSalOloRPCHi1CJs/FjEc+kVGvaym4/j33X
AfCQpuBMlwdFh9ffw2Oc8P+LnVADhev4Maa0IF+b8yQFOBR5k4mCwyY+LR9xpvbOeG6JBrXt3AUO
ZUKYjP1VAT7Q/fYOF6RwQ4162Bb60+X0/FoDQ78YxPtvD3MjT62sX6MNZAMNusyuaIoYa7HP9PMJ
hQKEi1BFAguBBA8nG6K8gZiYXthZPVX5PLGKaY998mrECMPxZS3wM6QetOvuPC0IQ7Vh9NIfhyGA
eLsYs3rqvXgyN9nl2PcWd6VF3LefGwOZUzR97yjSoLcBk2Lh5xfriQ/tQWvxm4IL2dE/EGG42f+4
GpfxBYYDGHCTmG+Cms5EEDH6njF3/G0XVZQcsd0+69/XHwnKCBkJje2hRPMYxJFlBRWU7szm5BNN
exf+KuuU9p+ZEGeuISoIb5MX2sLn3L38Yxz9jGI3Zf64z8fn5Cc6C9KEXJgRz+NfmqVsUpRXPUbK
LcQhNCocS5WzDks+4BdyUWYPK3R84FpLBBV3aK5Idx/h/TWq9CrD+2RiUakLOQmE+xBHUFLOmEXK
56kjqhyuCQGU2/F448H/jet0FJr56IscKsDRGxs6fcNkNA9dOTsGi9Ad8e1Av5C2xfCzyVq3747X
lAxal9QNXbUrdj9hc5JaUGdoN0lgLMqNtE0L2oouS/g/TEfuN8SwI7bphNqZNNbHj4eLvIy+MEJ0
I3tHLOzXaxQz6lUFSreOTXHCUsF0t83+VmKTk9VCLTDTr0MMOp+llO77ufsg3x9mwsHlrRGZIJv2
Q/VToD1jdLc6v6Hd4qCH+3QGh0Ee9Qz9zc+uxbNQNePSkYnVX16/37cq3TAkhixUfBQEEaB2tr8G
yavXn9OuD3c48OhNJo0eB/nlfizpgplQ/lBJrbCN7IH52LskRO5LK49z2R1i1cOkg7OIVU70GJba
eXexj+oE7Nnl7kBCOdnX2XWmE7pLeaK5TDC04MuGnpS+tCi/jBJrzvSHrOV12Ail/IYfLvJ1+l8n
otjo2rtu9sqoYlK9VSlItDI8+sw7GCAizWRLt4J/SvGfyZzkaQKRaM/0obqpcqH7mJ1qxI9WZNWh
hXhPme1rm6+P+1bDEYn+1YbY3a2MsG/wUWSp4n0Up9cVoAUGIp4YTjMvFyK8/piOkt6i7Zjo1kVV
+frqjGS66MSkU0rMvtq8EfV5N5iAo/zpb3cFhvI1iQvx2wCwHB5SKhv7WeSJRnDnZiGWw5pIq2Y0
Kqqq9iLEeYHPsk318DOtx2QMEqbAZjXTMhyy17dgUA9K9MntbUKSQBfGJ1fY+57WffSiwuPbsdV2
1BaCPPtzDZUYCHcSaRH1oLyIiHNaALSWdgueoy4S2gFsTUjySoYDPHxYEvKgkjJtFUN4gIQ1dAuV
ZypEsYnQURQpKHmFZSePHYPxPHRSfA76DpqzN0fjZUAyn9AWWCZ0t8ry9M5jGPQm7Jq8gebwKIXL
Ba+k1DlZR/1pa/vEsjV8NdPhYmgiNu0gujh1406ui0RcNb6tRX0AW/fz84r1caIrfzEICtGRZJgR
/z2bu+AFrkKM3mwOZ6uq1wfkC4FGhBxwT+8lD7aVoWwCiP/W6lImQGc/XXiT5LRtreEzuC2v8hvH
7yFptwiKvHKgfZnI7uLKaR/WHia4WUFFL1iNS0cLv46ukoBI2D16hterwOy/oP0BXfiips6EXNME
y1YYHMRLIb82PLE7hfDFhi3LVdfHDYBNVBs5cBTJjpBGyGTiiAObY3A573xk/G7BKo60naj4l7ox
KH30jFR/WH3nAWXLKIX/2cnY4NzSsnBo3Gm14eoZnltIDF+4UsUaezM0clK1jpuG2Tf9+QCqo8Du
AiaFWSEYxrv2lK7l0EIaRGCd9RcTcBA7H21XhnRvD1m2z+quuGyUykjSD6spT2OnP2xyCptxnVOM
0TU5j1HmVCVkVz2tGS0FGn3Yk1AoU5SCyAdddbAUZNk3/ebXiG0l7xcTpIoKVFhiHc3R2kqbNuGM
4APA/Bm4qsIgOt6ViQC+/nIcTB1V+JM6ZjfuPaLPiZ0mk31X9xLps9B3wQlk8lALpggB5w/Lf6zB
bkPv6VGpYDVG1LJWI8A20QuftofTkMYlWBzVQV5Vcf5nChnwuEr2fbnNTtuy/2G83xHSzAzxj67a
MDJPsQiVhH076Yg5Rlm4JxgetZKaVUSXYiI6pP64IW2mFB02GjnBZpCG9b0x2ksDZLKB3iCdBO6e
+MC7WdnJRiGfO1fhxB4LxtjaYqp6irFdEnQaxWT66Mx0hexL3pgVCHVd8FyAM56aF72eO8KGk4gO
I6U0g0JqAB6y2cJacWUr3HiHfxDok0QcwpDh9DVK+sHi4YoODe+TOwgGNfcZPbIKG+exR5moGzj2
2zsmqQxLEfOo1T5BfwUcqr6SgxadWYWB4CZv22Qt/V789FVrCDrKNqdFbgNQhS2+P7LcDafjKEts
8U0cKFYKvqaCA/Jb9fwJ3dblSdjgXBnJBDg8ihewW6f9dlQS5WJo+5bly820C4muDNaNGQJy/n9n
ZXvAiCdXCSyZ2TJMxtU2VQvxCwVXwk1ItPL7JlIo97uV00Y9qZ6Ihr7OV/CQ1oJI/ULxtwFwaNkm
IvaTM4/e+Q1qA3al5f2rmaQ+0TyRIFVpNx1Tw7hS0NopOlYK9IYTExtRgli4cyUz3QmP2qrjaqcP
Mj0bcX6diEYDBkbdMwtAglq/7XRR+oz1XWUgg47qiVTTHO6ZZTc2EQbddkDDn3wPE3WEWWSYzDNm
KTLKPsAL+LCoSAFCKD+MZgLdnNe9J3dyCYYHSjB7plllku9bXr3c1F5DDe5B2EmRcD6aXFhn7hj8
jCN1+rWw6Nc2LINj4SGGCi34FVzdfYMsfZILbzUuYs/Q+M8wRGnuhYisOXUne9l5LNLyXnM9C7tJ
vkaGqeM8cbT9VDybwM58C+rnjS+xLqlo2DEFlIN8k4nmOr3zUAbpcImI7EWFPeK4pc3/xA3cU0MN
8P9u9UHDxp6KC/TxPS93msmJ0dAinu4yg3ir3/sHfxAO7cmPOyExdVEjWYFT+fC/DWABETLtFvxP
A3cWJncieCfBekvXnPnsX9orJ/4DKTmdRO3imjQPENnFhl+NbrAK3Z7VdM1yOZo5ZQiDOV/B4NL9
A3fuxoviHxUlcdueU7RmrPi7jCgOC1etwwTfsBELIpRITDOBZsDT4voaXQeDu9KCslXF2DIaexcx
Ey1OkeWGovahkrCmsfRfNs+e/ALc0sIxAPk3IdbCA1scm/vsZr/B/Ah6MkemnKM4DWZ9NfM3dtVU
5rG+6pS9KJeaI9pezbOS6h1CWscrZKHssSC0CO+PsTMqzlD8IB3YPiaw6vIW2PDWBSBh+yemM+6h
t8rf5WtCKwOw/WtmX2hFfiOLxRv0bvi656pBXbM8T/1b0C98xKiJwCJ1yQoQw9z2o8Ajmx/lATr2
9WvjEqTfGX3bfPM1xdKlrcdsJek0TZ6Jb5syAUUhom/zRnmBln90pdDNuF7fmQjQJgDeXjSyxD1S
pGm1DA8LxT9gTkEmvnlh3dw919Ca1hnQ4vipw9d/T/7u5cv0LFBxiNS0n5Kjmf7sMF2kOD0u0teZ
tjE5WbEVha2uxHjbE/H6B0r756gciBscWr2AKYkQ55/TU743TMlje98TCFzSSvn8ZnIFZbMck70B
Tqeaf3nGbbXEmIC+4uSXl74eJx/3CmzNWs7qhj60Dn+T+W9B3EF5Xvs040AZg26WCH5G0fNIsxzE
KlKzMXGUhWemXaHseH3CaIV4NYRVFZh33YnvXhkkP8hwIR1eElyHFe59rD/nV33zQ31HnuUOWXjw
Q8mLUPUNI1taPuBU4Z3apDgtEtnlFCQan9Ls7lQ6UQLkeRSUI5GAbyX8i4JLhmi0Hh7eau9vf/20
sbGkPayCRw6DBpgkOtLvx7odBLNAh/4mo+jmLoXUA3FjXiWPvv4xd5A6KumlUaNHAL3teyseIGnb
VZJ1jH48E3cPUcpdISC/caeDakFVQQyYvBsiKjsVPy2kyQYXYju2SNtCeqt5gPlXmXopVEVNZFRi
jRsG2Insyux/L0EN1EpdUXNOM+NVdLGAaK/0JcNl/FZUulEg1CG6GkxvxbrIALqF3GTwrmM1i1m3
UYJ7SAnIQxejSMoIn4WJJU/OdYCaZ4Tf+madRkE8OchSqbwKqghYB0Qh1NpqCzsRthF85idLhwzI
Evvd3WLMwA7+1SO6ZAanxs9csLYERC3pAcZKSz/jYrzXdbOR+MZyM8FoIPnOjlUTt48o8VEXj6tL
/r/g21Tv8Sc3gOqyGORTs4yv0GrzTCuZx5wbs9QvB/YSog7y8YxE2a4QG3eCb8/0x+xXxRHQPqT5
fVOs+eNba/vouDGMe2fIhUNLc4IAPvKCdk8iBNzFbQ2j6xhLTMa54i+sVfYoG/LkhvcTMHuL3mQi
xZlo8H2B9819WkhbIXu3WYaNzJl9HFWu+2Wfb6yRH1Vmg18jHPDYavEwGAF9aGd/HJRaNMnoIJnW
8k/JO4M+M9k56LsJGla9WJgEaCOvUxkhKV2ua1Zm2BJhDaV2d3PM7+GSxFZJh2f9AtMPbgVIVyLc
o6o3BgVApQ2ySJbiGx9HE78Jl4jDE63jISqjXDGjQ5vBITjdV6PFtCsYXk962MTdpHJXQkj2FHC4
K/MkDQemVMV7F4AliJSrS3B/gHN2BZHU3crDMCPa4C7rIw4n2u83we1WRIsPKrL3WfX1EA36/WEi
XFP+gqCZHQIXWU0d0Na9Kyr731jLxFkJFgwwA3y7TA7CsoHmsr7F0Xfvn9lefjVvHtYUPQ2c4GZp
bmySR/pqorIWBuUKiF/K4oYsNXQlXDcXoENTSx0C36Eu9SpeePS3Ixmjv5j1wF55UJrI4fBXEEFW
/N925p8zWAdDcovQ4WYAujeLLDZoVg/6PJhqsAibMs1w0HJ1Ik/muszAYKq1t5JJAVSqGFZel5QZ
+LfSItji9HQeWRQ9toZWOnzAxbejNg0zMyZKpqxxaPqbj26ASw7OivrIZ8pWUjb4PxqzaLumYOrw
7IAN2czo88h/t/EMV/pr0FVYwWrcedV2sLc3MjdtsLY8Fkv0Zz8UGiVsTL2jtqyHUz8bVpyn3Hqx
i26PthfZ4zQKie+vkoTJRduCGyCw89HV1f79dk7tQFV94Rov1KZo9ZoFL0PFYh3TaE26PiTHWE6j
8xA3wEDHwADBT2rXUJcILL39WDczx7HOzlW8ASsJEV4Ycfe9tXlBR/368oiY/tthfjZm7zGz70BH
Xf+KikXPSFJAP43Kh1HZoidTnTfbEidQ0/p4cLi2xRk8ckF9rmFdEIxQfvJLLnhjdUIlJ3j9UH60
VnOKtqafmbifVa5PfPgMlw1rd/1X8udB5MB/T0Zq4afMA2yy1+INKuoOD3qJHYhhD+v6jFwqyGPp
3ONKlsIqqifJ9zuZYwiW97kKzzu5fYLTXhnVvMO0+Jfo3FB8QGcBMfsb+rwl0aHRTZFmvU9kJVEO
lHkUjQcd0DQZV2HwRvjYk53WnH+Vs7LHMekcmI9imTPe+hNI8Y0BklZAY4fa6Vur+IMYsrP+KtV6
/Wj+jBQLv9JASftbo6LsB18R9cGHv9DAmfcoZboGC9FjiKkxFX7Veo0kZH1b97Nqggl1cYbFgxCH
ii/qidztG9Sy/E7tieEwZsHgbqOQC/DU3p67zXhEPpoRAd4940TaeQ9DgT6oSEcEyTCZdptG74OE
eAvlTCW3KBvBMRucXNg5Z1+EcW9rVBGZYODxDyAZ9ESoOP5Hq44OPTsFiQFdUhzXMPTsoFB93dUC
W5noINs7uDP2bzT4tq8VcgEkLExPdXppTdhJ/jmpOUl/lBIMcraRIwMsVz86gqHgIhZeaui/HtDZ
MKLd5i4sDXXzsjcSNW1Kz46c5/G646Ul/TDni3rodTzlgT4eYgAl+UnBWJULIPKfhc4Pc/86dkyn
dyo3ICEsfBZfI58OyKHULtsVRtcPV0JwfeImj/Upl+QOisNSqGv8x+V2ppmg8PE1p7iJRtEQ6VAv
uoH+dDLmJnZEjHEy18OL84mO+VZFfWMY3XiH7wngCLp6co1FOAcGChQ+IiCv8P0EhKittniOj2IA
E1zGSFMs7mRR2PD5QuTzqKbAkPCI0UmmFLpaNWAOswV0sYUVDcOms7ofWwzsIQd3Dd3jGYQ7lbfH
rOzlDrC9LhwRvUFKjYxwibxu7gGNTiK4H+pJPvwWwyHezF2L4y8rnboDgcHX/J6krCVIVG51ZO+Z
uLNmx/3x6fDm8c2k5Y9Rdi8lyrixokUgpQ8QcWlb5h8kfD/JxJADNDgPGec/fNScyNYUBgoQbodo
giubrFaGhniHtnqRx04xLk68/k0d2JraN0J6D3560gEkVNfa+sDlKPUqp5ptq0V91fliDuFt/2Ro
X++0OqaJk0w1JhTM4cXE1Tv3uZDmRM7hT33/TjXz1krIE7B3AJM6HTe8h19hLL2/XJk5TbGPm2sW
Fa0+aCCYJrwAz52QtGfBZU+mrkEBtK4mYWhlvjSJDIhYKfaU3WH7pumHWacLA+S8Yarz85KB54Co
axsjnxgeGT0u3vzSerWKsQoc1AMD/xPUIEU+/xoWd7Y7ocjTEgT27lofuGqvcNNgrzw9UGd0tgNs
uxZrv6ZYzEgSEuX6TJSCa7xGNGcS+NYmxiO0A3zZx3PML7PTiwdsU5OJNkaGIFxhAdNB/Cwcx5H3
qxLNCHdmG/Gjt+c7nDBzjh2BcqO8YE/of4vlFBfAyItX+0ZA/VVdZT7B6d+AiRHcwWQ7g4WbNrTf
1vCehyMXzRmPiyKj4JyDSW8esZO3kSm+9newlS3u5to8IUpYbg9s4SAJsUs+jTDdUSC37BDnuICj
D+N628i8RV1Cl0iODDxHlrRvhTUVu6hEJcB3WgHRBZ8EnmOY0UQ4dpfHWY0idRL6bXXTDaXrjHbn
kj9dxYyitd/8ZZS/jUmIbc1hdtukYTPnCVJfGBgqlHJKL/eTehLKGO1Zr8rstL+J0u1SRoVQ2Uv+
3ZnkzyMOZR+XnNQwJaxQZKFMqG732TuT6qKt2NqHD7xPaSVXmTsBicMzh9s6Gpje3L4FfYxsz1ww
cIvnqkQXCt4ksSP32Y1chYSaiU92HCeXll8MEMOPh7harAI/78dJBih8MmOzwqatd+Smj/uNdMW0
gsXVIDvacBp6VyBDAVO+FuTjI23TQ8dOvsTnrlLN4X8JC7B/dCn2tNPFeqUedwtB0loGwvbiSyrI
ww8gJHUTSpiBusVWoCVkSuV9si7nXwCG3jy5tsa7+UzBijdEqBEQcs59BcMRoFr5ZQYagEjEuUVQ
UoYstFRuEzzw4O0ccZZ21YnK3ApzfiwErCwlS8zKYRxxJ3hI4gTT+T8SYgzHW4miSzoZFFpcgzm+
Vr1EzqbefmTB84Th+gOO3g1IP7UwwMgvK5hGpy0bmyMKYQ4r8imMu70hRo1ynEqXPAEVH1pSpHZj
nVWB0FUwxyDGqvyFNLglaN4zCU48fGdzSfwjBGvCKWzQmTX1pZWPQPVMjfOEaumBDfs+X5MEah0l
dGdD0LW6+a4lcuv776QN5F+0kvc0GDBF1Qsuo1tlUDaQJADbpZSkDRFyIvVdR90pHrQqfqI9X4Uc
VatYaI2nJ28NcIPPsFz6okACDnlVBBu6+ko9n8tkm7vjjL20KvLUY8F2+ULiEmd090X/0QNC16Ak
sOpLA8ICCgLWYbTpq2s69L/LUS1nWXPJFoxVM1QvfCNsvDM8r9R4ujSmAvnPiZcZA//el5/qtH8W
WaSBGkhNGwIVqS1gDmVTA/l811kBClDP4UBcmZp/c7TAhrrt731QMCIB2ECMrXwyNO2YsJCgYbZV
csYj/BejeW8+3OwsX2OzehAEJ9SnLxJv2Vgk6DyrwRo+t8YO3JVP5K0rpm/ES4gglEG34UhOhCZR
Qw9n6BmdRSC0qNQjxThMfW5Op02Kc+i09Sb91AiXlwqfxEOP2KB+0PfRS7bj2o9TUn3R/aHeRM16
rlXgPMeAELCKGeCnw0jzBOcJZi97cFXeyZrKnXFT+FEWbMnocNZf6XVpSDp6zKozjChbK0+xK15w
fb8MeV8LtfEQiKW107etNhMnYeo8oDMVx+GlgEUdBznUUaLey3iOnPDIUZCavKc0DRAlmGPiFZRw
QOvYDlpUCn3e71bQIJJ7NCKBE+c+gf7aYjifxfnSqsVxVXCv5n9Vocw84f0rQsLF8m+kSK87otxZ
18AdfWa4LGY6RqaVdw/MYi7JaAM3fu0sJKAu44Co7JP4uU1p0gMbadRKi3Sesv6OL5zXSMSS6MUl
8VeyFamZOy4mXlRZSH5W51UGbyI4hs+KKC8UzrSsGQRLIVcgEyb043wKNSiPGUyb2efRbEsCtQ9v
xRlcjFz5zTdkqt47QOVdfjP2KGVX3LguRpu9nPwCWg2j8YHii4DgLfPbjjTomwh5Op4can95ghOu
180rtqHuab2YaMJnNq1too5oJbUxfemBoV9AUSmFw1ywSvWMeifwWaaBQehDFVReNUztCqWoxKMA
trydCXDcX6Vm+ZsSobj/FLF704vyHTRvS2sWPi6/6t8LhR/F2DearbUKNWadoMz1lQ7+akgs0pzX
ooxVci4RF7PhqMyF5LPuzK8/iVIwG58XxYgJnSwpYrlIrwIO1iEFSi2wSBkjuvB5vacl4rL140DU
IwnMCgKhFN8cKakng+2eli6nwgNk77pUNZGBDR/MtY6mqonM1KI2HdJMsum2edUwKoTq6F4hJAch
htp1fVhT6tlVWXfjNgH6+V3FbEVYBBlJRn4Ht1i/OdM+kux5i9blNizz29xRe6NfWrPIa2KfOtAZ
1DpygYGYgAQsQ1xhYUw1cRP0qRAeDgJBRzwn7TTwdZMtthuSzIPGL0YztxqAa6VokcqitVILEjJJ
PTuRsNKiz+bL2zGiC0931LE+r/sowt9cn7j6no8J5Pil6L7o1LGwpVC/Q/hWz72YnmZMFr/0vAsq
OVUmyqkQDfTAObbvSDYoLeVlysqyHHkS22WFRe3EBOIPjTXOApSKkRnehLK0pFSPlEwagFzU99TH
xCSdgwtETT1KekeKc4b9EslIWliNLKVg5Wau+UWvr4gzDHA4DQYxTNPnpjnDnG4HxcoRfi+Xx8QB
nvualuOHnxv0qZY2t004VIOhqBnh+ymeTTkDqdMd7i2rfQtN2buxwNOM3TKmjbmo42IeWh3xUVuN
nBPNxUe3fcNWyOVFE4mqIiMmyGHm/33/LuYoEKSzdu9G7f+TVcDZuyV4OFy/pwiKkYvz9TJ91LKi
d+UjGGD1EYB5U+CufFHb0+v3y5e8GnN8s7GdHfoJFSeoM8NDL5ByeDDqv01fZRcVspPXqzPrZtNZ
hlSO9lPcXys2e2votuLojxIfLA3bZ2Zk33BWPn/2ZXkxPiavFvE6z4H9wxfRbT2VzQPlQN/tzbPZ
WNEBPX4jqKfE1jdPjPR3kwmQW2sfzS+5D8Z9IFiVVF2Bptpabm+oUwUe2B0canB69gR4t3yeGjyz
Zvr3MjxbpIzrt4S+2R0qPr7We7I1Bq+YmdXbCjPfj/cxzfDk9QjAzBg0iAfB14tay2Wj0fvNzFms
Ekm7n25PyipqY08m2U15yEAZLcg/vUo265OQ7907ldpjgGJaABnr2UOLnDGB8NYP5s9YilILHjb3
btdAXqB3KTyTCrUpDorNvr+6vXKpWdQcQpZmhyUWwbgI8X5CCE8quIRT4ynrI0wK5FQM3WrzllUO
LNHltU8b9qYkXlUclVkmuUAN3z2yvdVhy2A89x8zmYBrb1dbBsgyCtebRxfrwYxTxrHPmavfFTzM
GLyGXp1Wl9ug9l6AA6qx4bcfJwWw1eHJjbmB+LHkBkj02RIQhLh+pgOonnPNI+n36uTpiud8sXAo
352ejhQ8QUdJ6SQP1ehmFTCEek7Py/CLQan8JSIApnSdPq8BwFL7N8SOL/oH6ZWEkfz1dAVpFVmM
mKNX1WW5Btzvp4peBi1SjJ6CO269moIJld2KpJoTxbmNXTHeHv/hT7o1uqbQS7UD/1hGauq0xN2i
h3JGBBYJUZSSH2aIlanE+exB7WZLa4n/B7VY4k42j4o48qii6FVOYugMd+3fgFFdTE0vXU6z+f+v
6w0pkLuwlQH4JeACnUzj4WACSWW2kMib0j8BDrpQPWnAFxgTjWXgvMAJF8x2cW4lHooijEQtSFkq
jYzPZnf6OrOqU6ebsFYjcsJZHm71Tv9q4GygC/4BBpRW2hTQhCV0r4w8xKhimtuTiqv+EGb4m52r
1MbR8FgNSljTDFvxs4qibE+txhlfjEWmKi+JRRZjpJDQqwMaAgi5QceBcPIpkKyEpOz1M73NtBnk
GnQLlhdfKCi7dHEg+lXAL6+6fqaYgytO4NjX7jzYOVh3dIFrYBNVjOFQSx6TLyi5Ik/MDz9qoPdN
1Il08kBottUI0lMU2MmealL9+BUMPfzDxACKYCXa3vVLURGD9qox8gkWfdTW9kc7PMisCXI9kox7
u7T3jj/BzOkect/ID0LXv0GVEYt2cpltZZ7fdysy7U4ED/6h4iyooJ1JTlIHTSwbyP/bvvKfjIxa
8g5E+9EWAbECt9oE+lediYcqobvx7EyNogDRD9ROjb0NPTXr70SjryQxC0B3Bdr01ucTAF+4xDQ/
9W1roYPIJ9/gBtx5o+9+/ajBPj7RpFU9AYvrlIKM5cPv2+3mBv1BKoL+eysbJds3LefptBtNPQkI
YLqU3EEc8FL0ZyfGSu8iU3d7bOgh+yn7xOhrgxvclhP5BZDXnaGq8gJIvq1kFLy5hE/dUXOsy9+m
HgnxTcgExrB++N/fKQZVh4vH5oroqNbMESz+HmJcYGlQ+6nh2/1sK1O/iGZXyjNTMiWKJe7cW9XM
lhOWlLLmEa30ujSwOxY/yrFDVBhdLFnly0FcyZPrtrKK7oZHt1f6Hl3Dr5PndHDWl+EJJPV9NnW2
vYJ6NV3SzXrJGwjmClZBdiB5WmplxACRbbjHw7bALwGKA/w3WrwMl+2RnPLTcpCnyBsLZcp8PuOe
f6A31WIe/D7pnWS/on/IQO61KwENyT1tcJNWbVU6aaeAwTVL6ud2DimKJ0bFIFZz4QkTvK2/1zI2
UnX8Dx0L+LsWhFCtq61FtlmlHJ8Wads2RmZOcnToHWI86hnx94xnyigsq3rQ/zd0QkfH9qoeaz0y
TJJb2KzGRG9BFm6sjlTk4wcjrbqkCf1n55SagbgbaQGXNNfOYKD2BxS4exR9utl+TCKgs85l4DFE
83eMVgK8phe/8Id4tytx+3H+0eE/7+ZRnXAyWV23BYdovbvl0EujEqoXF7OvGRh0iNx/eT34Nx48
bYn8uxB2QReA8h4Thk6Oyo6xyKbfacPBqBl5i00Od8hMMvJEz80js9/Re+CijkRk+jH+A/xmrP+Y
zAbAwcbWzpz/JZmiW69zzwmcEvZSN8ocaMLVwnYmfvE7meeQcD9/jTYLLdRy5Z2U8YixNvZmXCJj
u1dyGP9UebOtinJyz1feDMZ4BtRMv49Uo6b9RQTVbFW24QLVzVezZEYswyaVcHVNa8gDRnJVt9Xq
bJp+SSBV6baGrK6IG5IsXgqlS80mIldvpjMccPb1Ef5JMv4Qyh/3fE34ii+VzNoO5tT2A0BVv2pw
aN05DLkzSgCK6RgCug/GRHpCpAFIK8KRDI9M0Z1h8/MaAo9w1OYP2WgdakgkLSJoehHQsB0GEuRP
jXqV1NDDVzc1X6S4mCJwy18FG1rt3BpxvI7eTaQMypUOVFpUbj9/VcnWW9H4VrJavFlMPxszc6LL
oUr9wbKNaWqBTFQpiQwYKDmgsVw8BXSzlcbj8i5hDy71I5hqhXFzDDV+5lOLhWXpfk1Xq5qg1j1D
ijlOJQLFbZhNivRzKwjkG2waXNNWH/eAG5KFgb6nIE7wa8SrgkFOZ6NrzpEeOTdrvbBbDRtVYaKK
5pS8fRNjU9fh5kvZbQg0QHsxFRW6nU1sPT6/p0r4gvA3xqE3BkEh/5mKVpn0Ab3uqSq3ydPbgcmj
Vm45oQoqA3/dsZWF7RjcrXOinwWpO1R2IVWZspuGrjt4vbV6hDccIw2N+XU2jb+ZO9g/eZCCT2ex
UHx7/CS+vLkxugBljC1CVrXMkmijK8gJ1RhqYQosDgn6mqwZ9xRkmbc94eMp05RitLf55Yn8gxfB
gfRazmMCWDUO2hgSnPymNAkN+X04cES7qsD5h69cquMDOQUcF+zLgnEKOtKjtBErwpZNJMlseVwO
kITUjyZJ9YpnqnDJsC0b3OT4nvIvKeBK2H/9GqpbazvfeVXAahB4rhapqnC2XBpG+hmuFXFbizvp
H/99yblaWDxjHgR89anFFI02I+p3UQ7MR9Nhf7XzDgEr0aANQIyTvR63ch7G+ueKRs3wXKYZ2roY
1A9iKyd+Q0PMiUzYtVYgtjUUGBVL2dOA+uDnESQr+cIJOhb5RemQfpNVbEp5lDmdkmCLoG93AKvi
J86JtN9cxiElhuiAXP4W6oya/5/G3jgT2tH5PzMl1KMYOIdB/E+dc3RXooYdyMDrTdWh2cVtEcmx
IbbgadItkQQ8cyNjSQhXqvWp7SBnUBqx5kLDV3DidLc8Zk+PZe/gqVrD1oRmIAo98drmg91aR4zz
5TRatbOTD2ZI183t7hmKuKQx5rdHNPLjGbaPdcPaOkQVn8w4Zfe5KJYBQH6aiRMK4T/YllbGk3tp
yT3ehC2Gpx+X75Jx9Hk1GzPKVtrkOBusuVVkoWZZqvGe1FMDPFejd0yHbvqy+qqwBDcztJDMFh6y
M3jzXPekTcVm0vPH/yRGBQbGZKTCzIxCHvEXUR+VTQ2F0Sw1al/gxtHz4/EHNW8YCbRuohZucolg
w2b7zyjX5Sfshdy993xk6CenJfaVTzOdQaLhnJUzv4nlkV/nBaDvApNilDYdwJnT2r0+BVci6xFk
BF9Pa08MtV6IU7HOtTXrm5VZk7zWkCTF4ENsDY4GoffLfgMBDOcB7kdk2WmzZN0iJoFN9Q971ehh
vXdNC0trpX5rNWCWmjbmhL3zqWif7res+E3OYoS3w8Vn+wmDTtgJ5ni6DXYlUhQwCs+ZiLI7EMXT
WCLW7aw+us3Qq5baqNdKp+wBLzixBdO72IO80uspSf3Q4nYRxGJ4yQtMdWkD2feKKgtTvqxQf3vc
v5rRF0Cnd1TwlFX1t3+E1Z4CR5iqOppqGvSBB7nW/BYrYkk6EyJuZHFHpJu4YwO5WKAF3UbhWSoa
OKT3U6ZDQxC9E0B13G8+2T+Q4ah/YlnQD3Zz9YUvyacC6Jj4QOK+FhJo3+bMOMZioas/pUloYsVR
NL2grPRRsIJ4zIzQOX5DfSkkCgkz7s2o8C/mx1QN7tCQmZP9phLFSzpem0gjKmIm3EAwEfou4gjl
EAD5JmY2WTll90QGHn/wZlq1sOTqRVaB2qskQrrwsdgqMvdumo2ykqBPjlGjjouDOeRA44MAGbr2
x/Y/k0PWbEFd1hK8bbIQT2GQcsHHH8vklRO69U57j7dfh7HtsasY62l+5q8oEno2GgeCytUc8zTo
NDji8H+Y59Jl1wbcsvP19FV9UDjofo9nOpgycXsMHXhMSmx0hhauFinRdyy9qKAi7E+6nzUR0/oA
MZxihfb8IUUGWgdIw6sXoY19iOaK0aKjd9gDr6KWMvJAejf5ttuRBuz33dwl98/Vvu6JfeDXobE4
sXSg0FkkdF9YUtv4SSJKoikPvbI/C+3wVXEqZMeU5tnCVuH9dCTregECfdsjCSnL9AaHGQMlJ/yE
c8Qd/Cywns46fk4Y1GWdBNYr/6m/slHPn86CXKMZKcihsyAlozG+/szmi3yEe8hOjpgDkAtH3Pr8
S1DlcX0IbS+QKsE1WOA7WaW+wk2osb3+fdOZJSVvaeJCiv7oJ9jPkh66Z3y614ngZoacN2eG5yqX
EEDaJluDRm2v3uYfWFN1reMsM12gVB3Pu0fZvhiUoy7GsUUCwS9Q+DrvecvVkLJ9sfv5FDIsTL5B
qjLo+xAg8r8Z4UJVqh/Rd/MGbFTFLJI8ccqi7x+CU9pLZoOEH/YrMhNBXcGJW6ahjw9BH/iEoIhV
jRB7Od9Xsrg+VrhR1CxnZSXQgXYFoUaRGQZ/sqTa6VlPX4LSE3cHg0jPPb4ZN9HZ8hxci0DfnibH
JcNSjp1RL3ImBYAtqR3SNNgAhcW6F8SwqV9/yv+dgRAIW7n3WHB6ZGHrQzHO3JpvKI5OlS7MHWK3
CcdAsGKNqL7dGV37ZFZeEtz+Otxd/Ls/QryNhYXdY29+s2D6b4fMprvDA5LWZlL8GJ5TWwTVFfxI
LPvZRkLLu0vFbpWGpsK0h6+LwuWrNP6eGlR80x7Y9sVRQv9yUVkGLe/1Csv12wO/SsSo7G7soDGP
24ZxblmBF5jX5HPH7gv85/Ug4jSrLKvQ6KrmKH98MUSXqxROJJQkbM4RyEjrhMVl9Sf0Ka7N5p33
uEGC9VyILqOfxfH4SfinR7+A7ddpM4tI8W1PMD6HSjPHAjqjoUcabIhaUaiSrnHh0YRYchr0ohWW
X1ee1jlQi7PTANhmS+GdGIlvioj9iyb3l4HB9paTI0IPBRwBrGfjVA0zdUISTem7NONwcutIpNRo
Iw7wq9vwpnt3OUq6cjY9VKBbz52zMaoYY75wQBu5Lude4k0t3yjiXGExWCk4nLjyBXWqOTNtJr0T
zm0TP1Eyaiupj6eNxCa8sx8IR4ikQTVnAJaXqZHdQSeXteZJwKUvZXdW0UjhouWtfSLWac672oOA
BJHe/RmXF4yOXEycsOwiw30+iZ3cVnXoxgaMP7+OnbPvAPYVWXIMvHtWFE7gQ4k2pvnTFbpJoYdK
mA+4Wtpg+4cQzPHRDp+PQ0KmBBepVLnjQljH4bdb0hzfIzwp95Q60QCGGBzM0eS8y76nT0DZOXSR
taNvG8bLshhYF3KJrVIAAlBxiDvgBh8JXbJiB1yKi+B8LBQ5G5oYxg0MDCXsVl/egOipdiE+fcOx
DflGvnfsrJBbI1EFwvYJahugTRcBjxAeJcGem4h8CDDG1NLn5MdLzdX3+W+fPpTXC0li6t429bfI
n1qf96nXhC5W/a6CvDRfqMzmrYREavIN6uKQKMTVXRPGQlV6UNE6K+33zCWSUYJr4pr/63RjxYyd
II3xawXhGqJfSCXyIfd3V816JhLeZ6WVTrSAXD/qmWWOK9aQG2ZfRRYGPEK2y2cR+AF2r1r5u/4q
q3ZVfGYysiO9DOhL3PMUKTJpMvB5096yIbilnvW9ziGTfBJz99igdttD73DWmOA1KsmqBw6mko1k
jFnKjMFnAR52d9q6vbceqBp7xo/s8W9l/vZ3Bx23LhDRwHorP6urtz0d6bqBhFb7KgnaYXKVGB4F
YprXA+MxoUFty3GdK/bcapws/fgHZjxrovJ6c1SG2ehINY4tOwqOmWJ7811vf6zcpzQGqgPIg37b
P65PdsoMCofLXba2OBK6tz0srxqQA4NIkoBlHM+vK3AHZS/nPZqMyYOTK0Od8rayhTx6z6baVsDP
FwyyncIKG+Fdf/dpicALdIVrydQ+pw+1NGrO2YMNgUj2OMGJz+scksRARr6xRRofK7QBIAURBqNM
jEFKD2Qs6PSA08WxYh+PvUeCUANuQkOQXXTTCes4p485OpwjPR1IFnPnuwcUY7GaVErQrWT7pIDH
E/kou42GWx67Nk3Kx31P23SviLgs0n/vJIuckfTD6hiJebHDlXz6Lg3oWCDJgDUNG4LODYCI8E2R
2Cx2F7nXdgwdhvCdHFBiqm2Eop/9ERC17vNUJb4kVpWfPHrG9mTN6tYgaVbRSYwyRcQjXBg3kP10
BJ4OVqL0m6y8nyg17K4Fk10zFSBeMTmWfYX81uUfZo6UxxkQhNij/SxOtYX+0s92XHglP/SGlJgq
WTrofaZKf8cz7PjDE+nF3vcn6rsIkwWU5t9p8Fp1uZ+hUbSnvGNff5d09FL70MExeGIFooIO5bg5
Ho7uXGNBV01xvZTK5jF2u70SRP0WMIdn82frUKt903ekg3+PoNJBWaByE1ziP1lNoQOz4+B0gJlL
PH9xaceAgO15kPb1lbJ6Vwye5QKKIoDEb1hEvFWJv8PyjsxlXR+3FslchCVDdo6cC6/BsbJg9720
RlKV9otZVgJcDCEhlga6VKFCi7oty/6isbqsSdBeVej5CQuRyd6QgNZ7i2meW+pf4BWwaW/0Y3RT
sF8m5HeGqAfMLI9Pxj7M/1AUbZ50odkOCPldIRgqqOPepQj+SAtn2BhpLFM0GUGlTdEwhIo6dysA
GIjhcXodsfe8d20wb/zAUCMp+1fYrwOeTXJ9zrCiWYc+6KW6mVAjyY0JbuO+cEN3CaQ9Jk0HZJtl
/LQ5iIWXROEabw8ymeUagXsyZn3r4Z0usol2dO4Vp8jllv/062cwe6DqswTdMEsOmLPgZnJOl1o5
j6WyfCEPpR24qr3sdlA5nSGx7NyL6sSjGdLQ9qbrzK4WYF/F7TRoL1Ao2os3FZX6VEKZD28pKX5X
YR92bo6irbhAy7U1u5HXeE0DeVYb+R0B3wsJv5jWjB8ROVY3aenX1z1s0F6mN/71MaL74BpgaUu1
SglPmFJZxoDBhJP0jBIqqN6AKHJ8bHXM8jF93zKHE2PVxxVNejp6XSvLqquQ03psb0G04kXgrsui
r13EE0bIrDo+ZlsWZRd/BjSmw3Md+LpMtrbsGjjtDk/2ruWGQQg3iq8WvH2ibjF4lXbp/a5000ON
kD8SMFZzsj1xWyf2B2HO+ojYMnjMXRem36J0n1wSfeZLYgfQANHbsYiDzXICtUdl2w+jH54SHWYf
b53y3Xwshzj6xLG4MfMjXfkPdcOWLlOepyxB1aYdKuSa0ANg3DTMqHgZ4pW8MEvKpdcbGoHRv3LB
xT5MVnczJNnz9vvnCdW+fXadfgqPeRlynAkS13nqNuClpq4nJt3uoKrMNrYGUUnIjOfEbMI1jVlI
SKW8ZX9jdtDGdVOo0eZW7cXWoSuHeom1vpkeOr8DsUZc/6d0aRQ6+48hNFQAXB8SfJZJc/ZPBLZH
QBS7LboJWk5KSwhFZ0nvPRfClBCwV+o3aOw3gq34bNNJJuQfScUpiFtYz6BnLbE9iuFQOVkm/cfj
t9UIpZwwdtjlAGqMnrvGYqEftOPHA8zb3c2OaXFX4U/zmNSpLc36orfwW40kGFttpiGYw/xxjHlR
Hf7TEjck3Ak/yIE6wY3YCZis/XIkTaNL07BvXFpyP8Uby9GCyl/44Hue4Ou2HyyGsM7+WZKkWL0H
WMZVxEKj8OYTOXGMHoxCFXta8/PeOhp+SVsxItZvj0yoekYl4s5chAI4CvpzNZhrwY0/iwORJyjW
QuK4Uu5gprpirsuGFsRxc3t6c0+4hB7O9d5qrBW6/8nUrV6ELfd3tSXEGmDN4fme2CVhGayksRxv
gZ/Ut6yp/culjJDat8ZttOO/I9hAi1968+6A0Ce6FLLBgIDpz+CXMcePasmg6bInP2YZ4Kn0nHNa
23x7YscqBV3VyCmZwfqPwzV57I5w+I0pu5qnCqT/R/FO6X4Tq/PS3Vz42D1tPua+nGSKoYYrm4sG
HemtkKjuCQ1SMu23hTTQnteYIGjULFk8BjfHZPq1+/BE26NnIKtJEZJPUeP45NFdDeO1xVEDOal0
EEM822yX90btPaQd0wCH3etL/ZBOP1gen7x9QG3cq1vYGAR1gFyStGvUXWUJS+/ZX39MRwgacMXl
6P4UOK9FlFGUZu/wsBlMlKn4EZwEqvnOZOUi9o2tXJVKRHeXZcGTJjaN2oCg7ARDj1zxZbOjQdu3
4n8zAgV7Hok4pcnqfQLuDufiDLExc+Bo/2dW1D8JzsodgdkCqEq9WLzgakoYHwTUNX2BEcOSLIf8
/HTBOrx1BWWj6ZybRVZSxuMC2g2wxd0F4iQTiYIMEZ4sJyjIr/WJuOalpbnk9C+BYfQT3IQWCfBH
ycXxRV7Ze2l4wFdi/fuQzLBRQ+8LHPZCjfzPpxmTtoZLznaf16uAwH1a05dRmkRcur6bOlmpQoN9
H1EcrgGg9hhbG8AVRwHzu0BYm12pVgBKrhX8aAAMyH6lHdJivAHbFoEYzXanpBTlVAOW+vyN15Nf
ADoSnAQCJU7BhwdEHZg27i20KsLLb27UXkm5H1oLOT6/blVju7PKup2lBz5sAJ6ZQguhgiOyrQhp
PHmkLXe815RglakunZeMzY1DplpNRFlJ6H5GGxyJ3reBjFnprS6hiBUwGwEKLfFL5WSesmhfW7wt
oigYEQ+qCkQnltwevmCI1nFNoQwDXn5DBSbotyx9bjEZNNTgFNyGpqhPKeUkPcEZXuSyeZWJdDkj
1bqLMT0Q/K1gyeH9q/mzD6M+XeysnX+t+0QYo523ZZfTKvfclNmhLFQ3CZnXRlMs5rRuZtzcM2mY
f61EAchMBXG7414Vtjr+OruK0uLCd+rqF4WsQiVzlP216eq6PxU+g7jQWx/v/UuGJEYQowmgRuKI
QAdCdJk/Dhz1Sv+O1UMIShzrh50M1wniQcJygfp0N107cXITQKaozBOHKsROFEBJYu5OuCbq+0+b
yziAGx+FVkyAbx2r+kTNgq+4HLLyfF3gIO1Vd3c05zoG2q6NXboPLUIfgW3JD/2Aby0zMNmFQnEN
YN3GV8m8Pexaxs+B+cbJb60vJY+0jnBE3OSq3WAYYAphZYYtue8unxW1ds+vMUBwurRkRf5NVv9U
QM6XOo2uoZwNbQOFlLHwIwSvSJ33a4tU5oJKLiq48Qcu4a831pIgsoNF+NTaUF5SUtZ8LLq3chSj
O9lxbEeKL0A2jWwmu1A9dYezK1zY1DUKooL2FpiKX6Y4Nb4/Lhb7QkvhTDM94mvJ/DjleGZmGtLh
WYL6EObN/IVXT0YMBX8jZ8ZCmGui6gbyWm6J8fvvC2UgZrg9Z+g+3GCDKVwuzYSORT2gFltmB6ou
adCO1wBrliq37bOuMGJTG1eutcaQe06G9HBM0IaQZqhKkY0fgbYOeBzCA0yPNNOKBShgESlqNKyn
E4xNJtz0LGrJzeTfrCR3reFVARrCiGVJaCbdm//fp70E8aiS1wY/ozWcZYwqRXh2AAdqODAX2f9s
G+I0zvSWFK71kzFSu3V2BtE+AvYhC1g0Zti0rOye2fXK7vUZoqJ76mTbz/Ma5WnC0BRAjReZizKA
IRyUq8u9AB1N5aiE/qacrCh8INpFaXrjpNPOKTWvGq7kpvqiYj9rVrDcyltYqqdTRDOfuoE/aLeu
8E8dvbOmatVFsxASKt9LqTLhOc7HIi5oj5/DOlke1XL2YAdWavoE5Hczc9ORScl4TzJzeIxEgrv6
/z/5MjXidziEowG/sJ6WQkf5p2r24vIeOLf0nxo67PUF9ZFZOj/QW9YeRsdTeUG9P9KASisZYq5B
Sbx+XQsvo086kCjVd4il8hxgxgHFdELUBU0SnDEh8HAc4V/58lxXzHXxKoLSIZ0YTiA6rkbMCnQZ
ZZFpPjLx8aDS8L6IapQwl65nK5rh7F/y6RmZmY1YNc99xXvSjmutPcz6z3vjivNiH2bi3CPUAECi
XyK3w+BtMQvPLNxzylN/TmaNlxc+Op/o+pB1AGIGu1qBPfuZv/ITiGvY+RwAsstFTKqIGaau8eBt
FBACN7ZECh/1bSfNyJi/ZFRza4ewbjczOkoGXPDTHGCv/niecFQcxk/cpWBd4kgBBqpwgA2AVgSL
9GMKkb3+o93hOZxsS3I5f7HvShznATGYq1W5YKZR5jIR2IdlffbB4jHZ89NMHiwNTFIUz3W+w03n
xWkbI1ifCySnJjCK88QHd0/3O2ZiADMHyo4ZWqQTmpi2y97i03R0k7fenF2HaawPmCtChnbijajr
hU2DePKvneoQ8WhCu6hxR5PqyLryQUkikZAXLoDt9vgZrZ2jDC1sRIHfogO/zD74JshYJwiuqj9P
UTGqxsiU3YNG7wyYhbbQ/eBcmxeLn3UVup9X6EOEq/H+XFECeZ8Aovikc0hkirTECCK2F4xmveSV
g5yUlVgA0F55tfOoEYnpvZ7DlklIkuyO3hPlAcwue6f6CR8klh2h7yaJu/hKDM+eX+IAtEktS27S
h9TocQjbyCET8FAmgn6fcToLfZlQ4mNEB4Pc3qQs4PQV0NAo6F4SoNynbWFmj70AMPgK0zvKEovq
4CTNCmGDiHBq5hbrXtSnVOOg4TTna1T9OQd14Y+z7LGEPXEzhaTtlgi1qCkapzuojHB6QIs/n7bP
J2NDdSDdRQWitYPi2iAPKGHZ8Z0QkdyxSgS+mrcQ18VzOJPAQ+TKfI8grQqN9S7fkx0LH2RGW8uf
IiKNgDO4azvmfTIb+7p46Pg5GBr1pGTl4jZp5eX3tcQMcaUPhGL3YkJFvPRlmRzSTSJUfCMun9m4
Sk53bLruuHrtYXcvKV8ietQPSdgTrjGSU50v/7buoPxpcaIKEoCV7tM3Fcjh64EPXCevnuIpLZky
HAP4bv14OwTP/UuXU5SdLy50XEYy4SpAcsARcgM36T6qJpLIj8ggtatWaz6O6Msv2z98xLPjct7j
g+O2wH3iWlXYwdUrGvJxQLt+LsvHkDjUanZzBAbLL4hCF5C3tgsjPVY809Y8Pew3+Re/TTPRrs1Y
W9xLFXsCn+K08v/1kBeuX+wgm9dZgoWywwG7bNJMmCgnRN5eRgsRhpeh+Ee//cNokQxJA0H0mwah
s3tfN7meOcD+RwC0o+eJ9eT4LVTXkDEnmHIuvCVQdPfIFd7HugumYS880ZOM3FrljQb4oeinmuY2
mI1kveLbHKl12kkQEndg6UaYMfpjj0X+5GIMts5v/XfK6kid2uKv7Xvla/4aKxWZNAypYJP89h/K
C5gOaS+ikKfM13DtsScfO0FV32RosF7/1lB1WM5zS5sLgPm8dh6+bpwYrjwQF2pVioHddEdyr9Y6
3uhBTRH97TzzxMS3xQcyyLiJPVgCI5KTC50rUY7wJSGShb1MzMbbgfwc9tNkb2L7kYQKqsGClsx9
hsbVQz2a8qVGTNi2mfUEC2kSAX7IphatRp6a3S5tbEfEZhhRB8vgHTUbyAh5jRHkuVwOkzYFRgKk
MNodi58YSxJGwazlE3AqIWXkYJfIrMr4IsbZr3USiUkDwLPyfY3mkJsr1xmfJVN6kWgZt7kQRDaj
l5N2f7nPMahurDlHBtVNf+XYP/6hK/Ti8t+fYZeIWJHPdQNpcuXPYk2WkMbwtnlIM91/omysOTBc
3cKswF54KdBymrEsTMpQmC2/S98EgjiLnQbtjG+xFBxjAyIT/MF0QcGAbrNCpBSQmNZ8tNYz+ukK
xxnpA0ARyiYTnjSHp+3cMsP+usa67/NEtIlwRx5EgT3A9sjiWCH0mVoQ2Pd7WE94QenBsy5mtuiQ
SABkQ/vrNVUyoG9a2Zdt3qIb8leKqukLGhB/HmmcU7v5L8PBodO6RtmJ8q1BsbrMNN6XFGfqNBMb
T2jfUIbck8on2c0hokGX8W57kg+HhU8m4T15UJ7U5BiiMix4yeMkkaZ+tdyr3mw/Fz+MAnT/GJQ2
9OVPU48qIOQI85Pytno6G2WsRSK8Rq/NIviMmrBBN2sDB0YXhXeIqa+/3FOpZnKz+cx93zXdaNTM
VwzbHTKZOlir0zzuxWEnIZJkoqi3OCKuzGpHBLvkIvKm4J8V/fVS7RuK0PSGDnd2Q/4uO+liXyU+
bm914vIw9QLNr7S53eA37czG67jgzcEVZO1BOvo627LrpJahP1oIL0z15PsYwHCAut0tWBGnC4pM
f9GwIk3RnOJJ8d1iEJyLAsso0925xeaKC0i7dCDbeK1AHyDPl2HGBEkt9N35nZPxhuV4Q1zHGkP1
BJi5I7LVr33Bq/ds+X10rRID8k2pDHMGcCNnpl1zsiIxBQcm7K/tnO9dfUzlob8DzIJ5ujhj2wds
Aj4d8cUnc0HVhGNTKCPVUmkrNQjAmN1neT3AVy0z13JibBobJpA3j2daVcm3eNP5rZ5ExhjxgrDg
QvKB5gw/+5PkiFa1g3jBNvvd0Wcsfvs4tEciGmK2C+LWsvEKUlCGQXSWozi0mCLgEaNAZoshh9UF
B4/DQniiRmwiCkB5dTHfjfsyV9MmQjS1Y6CUZ/0+DYlP55GEcPaPQGENOO4+BXeP2+GrO6ZyRBC/
fQaDy3KJgxt7H5qUKmccxbU9GuSPTPc6gb4yJzhsggzFoig7Vg50wxOdSUIaMlMSXo2gT2hdjFv7
Ra3CKt9jDqN0pBnsQFHtVo4Hd3d1XxoqBixxGyRJQZC7eBYJ9fJcnnuiALKon+kzUWEUGj2a7K+3
CGbuKZH2v7u/wsJnx3853hFeZbgQeGQe0PcGNHniqitZRvc+khk2eWrmaSUlhCVjfG6YuPitkZps
9D53lOdx6xIafrwOmfkISmzC05CiWfrYf6NH5GTWi81XglypTXrDrpBlrNauyX4Un0JSmb9ntjnK
C3vix0QunzhlXgrXZgd/l5YdVx92LPqr9SzfidzsLTN3/rOFTjMUdD3TU0YQ+s0EbR36Su7125rv
D1PaaGVRdm+BYV00DXk6BiRxMbK3cFUeOwV2f/yrIyo3dykSVI2xyGd18vqZUOS+Ca/fZqyfso59
Rik7OaxQJ2heF4ASdWuEG0Jlaw0XBb6oteHnx4csj3R8exaTpjKvti9OUDkBt4PtR77lWtBS1pra
0QaGXArQ7GiZEpzJk6uYrebedNAtfW7yrHovWd/dr57YsRXdY9B1jGFQ7FtJ5HwcBb7K3cfSTcF9
s9BML/GSh0WnIAml1FoIk9fKodM36oO2m2HSFKH4vU4V9YNkA6RGUPpG5Kw4HG5fPSIi3jsfEhFv
d55hGDVSlbErS+j6WLiGx2Wwg4OQnYWlnQ+khEZ+wlueLm3ItYpuFuGpW0LIHVEJRIkdPp7mFekY
1tvZnbmQvckFz2KOxvy8srl+YDEqN44pC6ixciuWzYF2wDtSM9zQ8QjBP62vdQ97VOr5oPdQ7beU
dgCIRIKzNtPL4dpjjOO97RP4tJRnTNuH+Ziud3eDfElQDfEmxfArZKpK3K+StCNQosykoqiBuzCQ
f5HSRPkXNlOcE7An26JqlG0AkRCBg+ThmnERYmXX4mdbIjshZy8W0PsjQWQTnOCYBrDHxXA4JinQ
ULmgi70vOTUzo/qRcmWl9YlQSdzGM2zP7Wcx/PHtq8x0HMd04A1G7P2AVEEumtC6qcsoK2z0sXue
b7mSFKi3IsKNH/OWlMFh5n6JQZIGnufu1CJkOucR4d2sIA3mdFBGMUbHU1VguCOGHUXBYnHfkWj1
f7MEQ8VPwEI5OL+4aaV5aApwa/GhlO9c3mTYYAnxKoTl2QKYYpZrn3NQggd3CLb0ed1PpK9JFN3L
HO701YZSHvuL+o4fDM3I7dGLuN15qsvnG3taJO6XgjS0hhBDPGWzjejREgaaxuqR6TRkkTYyVIuE
y06HUDcuBz48afPED5ITQP6/5BdP/nDRwDuVLAOpwKiv2A1Wd2wyT9Ymg2X0PIgCIZNri3Wt08OA
oSHbHJtDLK+wxHKP3kTt28Wzpk106N8A0w8PmgD/OL+miaF+/nzi3snhqd+foqRI3GKV+rBW9bTI
tn32jmX1/YNeyyqw/asiTMlbU1pR7AUaQZxO7GSVLR26k0T06o7n2Bvpv49CtECuzyBYnAPseWye
bmzZkqFd1OKg5kzUMw1O5tWQ20T/ahfBKOdS3TV/4L7RFjRJwcPAvAvtoEQFByaNciynJE/DKqMC
Kj++enyiF4fRKEUKyPVFrHy+HZb1PRysU84QHlbC39BKMeiG8y31C4t9Q+FoUXZnVcpSncmH87ye
5h5/KDgRQasVJCBWEpmSKqyz5i7X7RwisO+TquY1jg+EceChPmxlYhKOlLoX8/geOuNkPkAuY64/
2g8dL0DbprJDcKeGq30QUItR9BIY60VjMpjUyOaJ//yUFAc/ssf9yumG5F/eHP1S9jEtB58qhafE
Kl79aCX/rd79USQzIgJ2J81sdpYaZbIt0Fs9xJBgyRe7E8ADZXavtX4WLxQlEA+PfVW8WSa/hc/A
q+n3nLyh7wT8sNdPLLknrEG57lhYOVoxf/VK1ly16i75/eyP0SustH+PaV8n1OSs0UiD/x7NNIY7
nFW21Le7IXBOk9G4SygBT8b9N+15Xs/Guu11WpAnG4PWg2qV7dLlmQ75IPru0NSTf7Kf85XlBgjo
0r9oc/EU9lly1uuSiOhaN4fTPJU0ia1weMmIyjffcuCDyiajyLmOx3sl1KbUKbrSjnQIrFL5edYz
+r9jYxG1b97JGSKr/HTTqw9aVhvuVXJ0KZBAnPBc/rGO1ZoeFytvbTiOPuRhZeLqsKM9O0a9Y4zD
U+O5zj9Q4RKFat+O1lzMRSkoVjpQzfhF4GT9yHGNupHLUtoumrutdkqHarDUXdgcoNNhf9FUMgQd
teExDZnfjqxmMxWe1iLQfQs2raoS3GB69cR6zDe8xv+uWZT9Y2G+fLiA2drL8clIe9L4z73yn4Yr
E8evjVn5cz7mbzJa7J7z338SrKz8vvHfCvCoUXyDSs8Zfh58EzzDu1qHDIKihrO14w/S/McjP1YK
6NNaockfDylqmPGhitWEZyfARTo/zDpHPzz/b8D6DviyFX66JJH0TDZMMdzTXFhFWNozDWDTJQw0
pezpW9/xitZGBuvx97oYYPc0YIPWz1T8uz2bC7bVSKfWm+9mZAR4S9d8CZnFztHzN+K4IEeK9BhL
J2D1IrA/6Vm924E84igARHPZjFwwax+1ptUNuNqfnOhztOkWwHAB3b5ghOyzdJ2z2tQR98DeGdr/
Jr1iCDbZc8mNJqXk+gKilgHGSPMhJDPqYjqdMgmIlvIVsN55tMlOmoH4mnO5f4x7gqeRa+9enMQc
F7Tm4709WosJWMShP8FMbpvuphPlItcb2hDVW10azCiL4Wz9soH8q+kjRMhcwylXOpDYnbj0bHyP
CeP277yz0pBOrgQAD4Qog1zAooDNYt1BAhvZYHMru5iP5G9SjE/2+gaAdBIGfJYG0We/JnlS8xtD
4KKH1DFVzrOTdvhB3XoRty4x7Tim7qVv89uKVnuwYmXfhYXJbNCEF2o49nRy9CnVO4ee4M6OhOx+
v7XNvY8Nx5SpOObLYotfj7S4cSqPLx12/Az0UvZ3hb5oXvgbbn36aiyQ5HRWxY+4uy05wDjgGBJr
T29TLxUvmBl20/ORPQSaDtvpCVon6XHXnpSvCCs/6QZgGm4AEaRKveOS759FMiHTloYnhpjnC8GH
I7Xoc/G6EIK1zrd4PTmvYDQpCnANC+HLNSHWYIw49gXig+rV+hmv6rnI80S2nn0yoxQTt94l4jTM
X5P9NAY3CM+g6gBjgQVa6w5Mv8pwvO4JX3AS8m6ugPZ6fP3wPiGvc4HDUS79bqYb2r5ZidRyXjU0
VT8CtVoGJtALUnE2jKAQBxIO3yK4A4OMVQuoHXCjbV9nVjTlUG/y4hI8iVuz3/nqLhQNg15FmVKN
226DLfXMHxUICOJEIjoaRccRBfAIVhJWPPJosAgxVq7zy660tEI53GPwuMjC1HBj/lzNq+h7njwm
rQvLxTPpk9ydhbNQcG83VrgSzonrDbmTW+JdmvHdB/ExfMs6qpRbdO4QxeNiGx4gZLg3SzVRI7SL
rU1FIWJgTptEZtJoYt34N4XVY87+qGLiJy/tOvgHmnrXkAau/iCRQvuPvpO5DybksVKrSXY10qfJ
rwkz5FnIyl82H4WxL2IA/G8Wk1ALXAyhScyWgLAzmIgvojUN4OzCILugG0Rz+SPBh+bdSkDsSl+w
nkWA5CUZIae8F8Rr8JM4w9t7HvLyFbDmM5D+FrzmT3S4Wy7ql+oDshFI00o6LOSGIazv92cbwSy0
hZ2qx4fZzKQBp+AK4pK/pHR4juI6pvQHyUdNgWfd7tyqX7XLlml7qJWbL6ALB4ERdzVk2GZu5aRc
4w9EkYCK1PbIuNk6WcYunhXrP2dcSzmZjUQv0VGh7tkiMQCHQUqaBtXdI7qazP/liHs4DQ3QKNbA
W5ZFlQyHMiH3DUCw+04CeVprGQjbHCgrQjsg/1Ni9GOxyW8eAKX5XdAtcdPHZSgUrqAt+gTEwos8
FcPRmfPQ1TXbeXupKHK47B1PBm6dxVnyUApv8BwYlx2Z4jsTbr1DoTViZ0gp8jr2wh5nFZb12/83
LQaClZNeLVgn+halTDvTX0OmwfNRH8vjHlTIMfsqRDAns3jPdG50yV7Fx9y+ZgCM/D1B9IAhDuVo
OM3Kroz6SxL5ovCJ/RU04z3A60LX2duw65HbC4hiaheD/f81VKOmYrhaT+XEGdl8H/np/RMdeRhs
bEUtG1K2pPjv00+J0S8yEVmIv/m6EHTNQpB9EMTI330JbZb/P7hDpQbQCVBBeghMD6se3/mLLyXr
WEJrTEGDACwSMf3ShXpIL9/bQdHUqdj+iN/Xz0Aq4a3P1JvEe8Ud5c+4cK7pyl1B0r2XpxCTyGjh
8ljuqLEnBAJkkxUKQHcdopSRNtu3DCZOYYH/y2eVmc4Nitiuc+VGVXaC4fLbc5dvCONhwhDCUlpN
RLvvrz4+M/tIxBrbbIqbMFvlccluO/kkF2Z+3rlpyRmP76Cdi5sNjm5LZKWf94n4dkVr2ngILDmk
A9t0/tWO3cBn2k2ttOtSg3j1gU4DARVE3JUuztWo5xOH0uZD2IfYaXOnfoESuBOUKr3A4r9BXaIO
83uCav5k2RE1lHh5IrPShRxm6OuT1BvPpLzO2I9rLvmTtK5OCrXBJpLfiwk/zMoshmCevEE7T0Gl
HSxyKYKANcaxDOs/L5lV1mdFyfxfyjo7q1YFBd+Wj6NVoLDZNYRW7tpezoVPNFBuE+sDtN00T3Lq
rFgQOLJSYnvllo9pZNRBVQQjm0/uv/RW/ry7Jff6wYHmdImg+xRVv7rfuuhUIF5T7QT5Z4nuSwQ7
FR5QdL9VV9d0BKx7BxFFHrShqKqlQcK4Zx3hyQsqPySBV4C9fjyNFovWb4bsPxlkME50CmaCVWVq
76aoylOD6FWLs+mv3Yhj1exc9IPUGPfrn5rXHBvF9ohd/ntAbRWJycRqk0qhTfw0/8R+b40GuVxw
+fmRySjNemfHJ3oOVo68b4PhS+Qw9HkaZF3DjcIcdraP3yPpTbWGpMh4oPU7OdJhvP9DLQVo4Ur9
hqD+0UV1FuI+8VVCIF4glYj72l3fKPHXOfBnLGkew/dVxjj0TmSMH3VktvRSs+vzOrfDBvm6yOoU
Vlsk6Pog6FbYErBKlH5fRnhvZ6Cgk+qXQu8ojf6lShvM3PiHgHpr4mFv1duB3NJRNipetjaW0Xk2
8dYYvr3EKBTl2tzUmw1wHwN8CS1vJH9gKS4Vg/ipVVKMXlk3pPw5s80frCpDpkUS6MZo1ii9IxU3
5HSdmum1IErLOfZDRICZZTpprqIJ9hmknZvCHVw7flsJGGbpaGTPChgYYMg+EvBoywCERJvzgTKy
0xN4b+onlsfLSR+sP7dPgA2xDZ1VKq11c62qznH7HpoK9plZe0+ya72DY9eOkxd5mDBvua7xp8KP
0S5jw1hjHKq4mU6jbjmkA+TOBEa3fZ4+PwxS3c/GhfBIYD0gKd7npL3sjAID+DFghKOxkConn9g3
5MEUtjasoirEmdFVgTHwzChQ3OkE/skSvi4HaNNKg/13+7QBZZdtceg9Yzx0JPZkKF8D3IsIwOq/
7PekOcVTrtUPGqRHka33JO1TZKu6WEkCn0HEel88AYlXg3b48TnDpLCjVvca9gd8X9uTNaX1adRq
EETLnaBmMiW1hWuE2x0B7IX1dhz3k8lwPVsD8jHdELo1g0u0XlUy0bqrcx5zbiZO8gSIe1RWviu8
yS/vZ18x6FUOyuQwHO+LReO9LZqHIZB3ucbKmkxhBYj043W2Bcx8bFCZA5bvrQgk1YnTBqEl+jPE
1y6VPyk0b6/9+fXKQM7pdJtsHHqmKWCthwefxeFCDHh06m7DvlYVyRDcF3H24lp1hRyVMj8BerKM
QXavV3DqxVX4ikVylFXnab98En43h8IrzT2K1oVKCB6LohFWWJNRAPm5t1E9ONnWyEQhxJuJENA2
f9Aslbtukfm+jCBR6s6gypULzvEW4SVkfvs49EIhh4ALXRFtrlqeLEzQCfyFyURnQMVjHWUcjYSR
pzN8bhhT1kBScPbKdMEJjb+trZOh6NHMXOzeuNDV3z+jrgezzke8oOMipzfGTLOtn2KFxAwIbgGA
UqKrBLWrN5ExWNjWPOmtDv+zDNVwWFQY74h+kPBOasaA1avtMV8gL70o3/bCPPjvrEZpNP/zYUHE
UZFwPxxORKYkAMPneEuXZqihZCrMyXdJDwKsb2DcAtvyjMMY5HNy9L2EA0xH038PJigb7ap/vtvG
LyTxNkkN98MR46oyqV9xhN65LpPjwKEIbKsf0CrxXOKsxTKoY/PeX9lmm93Hg1O9SOuKi7r3LP4A
4e9pVM76Y2Sh1kM9f6K9S40Qe7kzniavn/B8+leuHTYMv1ZNH7KZkyuo2gKVZudHQnwOg4bHxG4K
vpqnHOyYudGled1RgkuyAFPsCSGN84IdQs1sJqLZuX1Wr6aWJIyWfsag5DX4lIB9ZNnU0hlh7IXU
Fhjjve8/3Bm2tSt4cRTKuIwa8xAw0sTiWHQL+Xm0W4Fx5jyVTBu7Lb9OsfU92FeGXfAieSukJO2B
pYwIZEYFhuh4/kXIvv2evZZi2U0WFFfHGpr/Ah5Tea8srZSt+OMdyPWtkRnHeqGBIQ1DMUzBDZg2
RU182kNkfF8ZTt+SN9ZbiavRBelXHBVH3rcHDjKYojkUGiHgLfB2g/Qaj7F/uWXQZCl96C/K4wSv
uLb4tUiLeK8ajyRnwoihsbos266eT23Oae0bVeZgtb0PFkm3ojU2XgZeen86uoL8jSay3YEn/JBl
wDVoLxkthpwUyxauqZ+4Tm4E46zKt2LoTmdzglWT1aT3hliHz5QHZK8teMpihNKhxoDeHbCGZEeE
h7z1eDBFhzZzMxohXny597QdmuVsiDZla90JrsLH9ogbGec+tqyjlmKOtF1PMkMwvHHNGZS5fW4M
jVcMwFByYo3YucpdDBKC23rs7/7kzWTzqvcFs/R7c2OPXPOrINl5NOgcdtlQk8RYyBNyn450ZnAa
ZePjlHtxrv/fF8AZX+EQNuNNLYDy8MZOBaDu8h30VHTj3sIyMNJ2yY7k6rlQ01E8lA8/TQWNAxEy
B+ZhHMQHCp+shEFe5ct8uHS1n2At4SN5XXT1nO+DD0X2gniPostE+9vJENdeKwuUM2ZpwOLcBAVn
roqMcBAiKaRqybarorfVA3MdOPylQlq8TKYPlsxaWQCVtaXZ7YqHzVWF+TOkycoU2V20xjTEG3Ms
FjBhOI/PYeoYXLjUK193F9n597VCSjaDm+EceM28Q2XprDrYizRruzjnbZzp3Pp4ODZlUA3UgDRf
okR4Qqkmo2jwNse3Pw4uyQudl/NnEpzGz4G+FB6Tt1EsKBSBYaxI2tzF8nPRbdDfvp/X0EWj7FU6
032UxcBjFYEcrBUa+6PR4xGLIvHLH70rSCPahKl5ilGN1b/veVXW/3OKx+vEzaofpa4Ntwa+wKpF
gbBjgfLUVattqfSbqkdq9k32QYNm2wsfdnkXQ5DSzHZ6G4eL88zdWtx0OR7PdQCaXVGPoLm8nESY
wBClwUyG8Xm6ThWsgQ4d5a4JvcpPzWutKORXPahWXjDftXbHa+bM90Fp25VNfE+I54SNVTQRXDJ7
GRWduyYAyzEYkPo3BYbI0lyFntLCI+3Xq60jPFYL5+pM3guAug7HTMQ9XqslhrY/3wqhg7Cq+meV
O/M2LidubqyoeOvNItqhITQpDK+/P/CWtZir8bJIIPwir8FyAgeiUdB81O8DcyHhz7k/sz8Vnttm
2C+PITrUU2fBbwnRGhl19wFyIg6je1G+XHx4BqZ1Duknx1AC0sa8b70VthK1IjvRKwrbeMiknQb+
GzwXRTDAZRL255JDmqoGlc8d6SpsAj5WPjwG/SfXgOkxh785uQe3G9csJrMYtwKc+EuVOmSHs9Cr
jm4guYNH3Ys9HrBEgSdgmNh2Cpai42DlrxCzoxWRYPW5NBm/K6R1/2RMIjQxPhP5aSz/nEbQmeZe
TRYN0/PaK6ZWzt/Lscpj3WTdpwpaBFAVS/GJR9GaXxTOLI2h+AJkj5Vssjb7KrgVBvDFUeaP3i66
nUH5q4EpPrWGPZKYSxz9OJzDRg/+T7OLGofb1f6eSaLrcG20HADVseqOIrTl9wYDfpAu3u8EbVUQ
OH1Q7rdLgr7XfOYqc6AjCXbcQZpnFTL3QCksbFlRat3b1s5xkobNYuV7IURGmwU1WQ0T/92ALsVW
iiJGDa8Pe50aPPe5+O37gpsbZqcsdV3XO1wnRXzAIFfpdl6ETW98Tgzn7YwqbdiAsDca/CN37VLp
3FbWStNJxuuMTNjdRpsLhwv0MxRFYNI5VQWtcjhuPnsBQ0/PfPjSSnMcitGvPghtPw+IaRUCAcin
HY+hytoCY8Ghp7iXt3yHscUtqsd2W7ZnTRSOwzP4dPhiEdsmsccbi51ECtcT/aYt22LNhCxUAl30
giblEbsU0avMIrwkppDlGShflAdpAWKcJhU7nXYBDYnsN3BI4e+kX1TSQpd/CSRjjLjS15YDfH0k
FkywsNU2mQbjeUmTMww6YDbBS3ud44mDfUlt6w2hmBFeKULA6q0FWZSiGAEmMG+MwjPhtRt0mB0I
Ls5RRWLy4zIaVY2y5Zs71Z0eMtlVbRM5X+soclAmcZOG+3DizZdRI3hT/9TJp0HP/0HH05fNmPJi
4GeLG1a24lPI0ka5/nQUFxZv59yIpmNKLhbZpIXvofLWd3F4DL9np9nrxcmenQSgTfxpDg5b2Ma/
YLnsel/ivan+QDI1AoUkD5OsVflMylR+gFP+XZrYGauKCxMB5rW2tUL4u23qgvrP6KK+MIBMyAXd
L3hZD58PYHRE4MaUzMV2zyXV7TQQwTiomb9L6H15EsX36OOthZ7yWHND6r8Fn/jOsij+uyYO57zK
8chdsQ4VsEzyxxqV4qkED4quJleIEHxTCdcxPwwILb74XhiaZzNRH8b7kAYQTCO1kCKSlafFEHMZ
zmlqJGMrfOuid0q3epaLjxBnoMRc8C4OSVxiR6uwAEIOUvbcd8fh0D0q4dU32gUFovq/MkS+bYuX
RdBuIrfXwS9O1m9XhlPxjUZgipZ6EMrVfjsF3bLMH7ZDhpon6oWmHTAWKK4Pscz9+NzQezvjYZnF
ZYNbcrSW64SRXUb2gxCsFzXfb2wybjt9DkMMAPQfbI4jj3LVrwsNGVpKxRtuVSlZb+wEgWojRViX
6bnDpP5dg6URPK3ehElbDruOdZJ6BuRuODJTov6VTUCY87GKEBXZ8hLawHJRkYy//7FfZxDBwvM/
qVYRJkUrkZgEgws1pdD+xo8bg6z5dwZeo/pgjIZPS213kJL8HSOv7dtLe/VMXQp3aPXfAv2cGzzK
wCHg6/EanQkAGptDquEJsCPvflKt52M9zpYUxKG8hzlQ3bQSeZwz1bo2y3OQO3nF83GHsq3XWD/J
ZPs0Tui0X7inrqmmLn4y9jXTnshcThcNoiRxoziDbYdMYWeb0Sz75nOKhfNlv9FqERYihhMnDhwb
QLLF6t+TAhnolBJfkwF60xsc7LOOafwVfWrkGxmhOPA9EPA/8nMf67j/4QoNTTRhHe6VlvOKEWZf
YoJZQjvJY/60xxdB6R2OVwhmAesEWzCXvFLRjDoSkwx4mcLeNgNMXKbOtm0LrcuGhrHdqUg0ryrO
P1QpFEnaldzxGRqjyZcfphPj0m+gX+UGa/QLZWfFeW8H0nsSIgMXjRIKsCx1Nw9FMN11UdjwJJni
lPdaOva+sAQl76p2httH0l18DC7nQyEQ6oYjoiHGqiHyrzBYHFtT+/a5NOcdyrkNQrsgdVT2FhPI
HY2Jk69i/BuES/ijoErdMeZNYJtonHTeQKPaCSZOXhUB3nzTk/H0VOTS/VuapHaotM/mm/NER9PI
/j1RXsek0vglwR1DIqkUy8jHdXr1YJ8TIdQye2ywYsZPh2NYhy2UdonWgXgJXEoL1Uev7g/ZwzI0
6NjUrxxDQdyYBjMdbrDr3mMI2QsSVT35SVXQdVnuQVSPBUgVPs2DHfHKplZMAHCYuvqVt3ukujTz
lopZujkzI/1jjUPey8VuDm3+7sSyhGPkna9ndBdP089rXOlHHnGf+rS24XA66YdBou0NL7baYhzp
+l6OfjqMTa8/NAx5KIClIDOOkURxc4iJIaLU3FIp6UaUR5JO3tFUzdXQqZh96HKKcLyfZiR8vl7E
AyLK9WlDajJHRIHaSxOZxdpr29M7YIQ2j3t+muT+s+iGcb1dz1ONfO0gRKsSQa6ttV+E7mYkb7zg
E1kLa0GJPfdBUSUuXKz/BX+ins2x6NTF5BCWr2lrMMLGclBOWNp61rM98iNQjHgxrAWW/ZTbQwpr
EO+ocqW2f6Qrson/BWeitOFzyXYTEq+jFFt05GamNQKW7IsGAhummzbmbx8dVHXnKcg0nKiJpVMv
jMspn3Vhr1CTGpKkFifIxMP3nrJw+UcZhsG0p2UP72+bpnbXZQMo7iG3uDtL0KdMJp9pF+EEYH4o
YazezXGInyUPILSUpNBZq8nqmG9Qbw8HCH+5tS6INRQZuTNzeH6eL33/QtemZPGPZ55xEp3iRBmh
Qp0G1CGaYfzwUSbd8aQqBd0ru9elGF+BXKvccTOwFtnO+Q12Mvxs5TkQbeS1KwuL2CaQTmdlUZgh
GCag0uxJJVgVyi5DA04h7mneENMMKUVW5XPAPpO39x68fYKECWBoBoiXIsHRVYqelvF+wCwJyw2T
FMVICCcRmZXsQsGuYLHTfHW6Lb2/T7s14zDe9ANpPS3CyopAcygPrvdI8MUKyt1J0LXWvuqEKvAN
vnRkNNvYVa96wgyw6j32OvJEhSJDYSB3ZLruTi5TnUU6qOjCS8VlJvJR/+OBR/Ok/Cq/0EVSeWmo
oH/2RvF8kgOgqs3MvYnvl02oZZNREuCkZpBV2wienz0psljZ48T++u1C5xmF25FmteK1v0uQvqJu
n8hEEqcUFLKObnXlsNG+Aho437KFdWJR7GmSqDs39bukTkD7zFO+xxIPZ6oWZg8z+WLrcwkauK+T
rueEXlgVcU03PpPSTdEnSyi84MrBgvSpxzKRvG74wEBy8peRITk1hd5mMRfQB74/gD1fk8y/oi19
KK5W1nZS91pN4dd3vZF/N3oV9nbUvukpdLiBnm4z058+vafvg40uBtxNec1gRHiNEiedMHNPf3R8
+bzXAd73sXv7T/PwZQWvL9Fj8ZGko0EJATvB+rbqLDM/0tJpdSBM7uXEI2RZiEi6aDUbK8KUF39Y
E5tUx15A0S+XwPiGTlQWE9SJSgj9CMmkGe7JYfyiOtMRAifBjLqvrg6Ht6dN51FdKqmGwJbibkK4
9E1tb7vh0V1TMVKHZuf6YiOiT14rKXUrlv7bKlcqWgQeSvGhqvtx6fyjdo/HTRMrVIJYUT2gzFJy
2LAYaW1E4/pg0U291+TkRYTxuMggJak0TJ6EweP1KC8fUZK21l/lxuzAh72kpWCQX4EvDjoYZ04r
V1/oE1EBWMIqZ+OprneeIU7x90Q+sNFcfeH+JYSFlaBaXQo8MBZ6Rp281r96JoyvW4ujl+flIr1T
3/WAktUgp1iBjZ6Oo+rc6H1GplQgRZtsxqTPsyDt6ozNuWjYdNQMhL9HMdTJ3CZCYzq59Sx40mQ9
qo9+8q/s1/xH5peFSidfGXYzfUEvkgwCNJSMtCM1KKQmN13tHQ9mOnDkItmHjOileQ+tnyKxLrUD
vmiSJyQuw49qd5k6XHs67ONxkOUNTvJ96FgAbVlp4o6F3c728Hi78lLwmYpcVm5vfxeYu5+cZ+39
Twh729yTEsI7uCviU1q1PXyiS+uiWEe6eoSbVuB2KvcZxp95z8kwcRFmVJWeC8pxe/5MltP3eqoH
pyZEe1iuTTWoJr+GiQKvRws0NRVU9GZBex0YCt8D6dXXVH0xQERXZkI8GoLPAYXJL8wka4lu4bbc
ANml3C8FsFoWZiaELwZmGVTgXSyiDGfKUq6HUTtVDVhIdcZvZYo2NLJfKHoy/0Tvp12y81Rmq1Sw
pqUhkVFN4ZLSWP7qGCjfuTJIDOh2mU3IItGgt5Ts5DW+sWMjFd27lQkug91YygiiQkfP2/ZRTR3V
tc7+YWC2ZQmHiR/1ORMvPj65B6+kMpyk/qnpQXTJ5/hi6U6aExVSXMXi5I7rKVsdQhWA9B6479dl
S79z+vivyatbyatgT8pRfDl/UK+8KDi+9aNkQPUhbpI/P+d2tpBsBpLCCs6Sx1tyh9di6yq84t49
oktF4bSvbcPdiBUDSvt5BcU9dm4x5laLU99e9kcTXdQikbIFTE3FD3fFFlZ0A6S+wHqPwLHSBDGJ
Wz98rsFpBKogfrDQAG10bowAoG+SN5O+sMuDdjxMiPvmI9e5bq3YNGmYhA6Z5DfFiJ/uB5LartY8
/GIhafd0G7CVtofFxhx6nGIFDzJkLVve0jhzWHkYyVgHxwNe/zzQj3ABpw6l35SR+6OTzpiG6sMy
PZrkTalECGjGXFN0/VpmkrUjEQX/UMvBGdjKh3OM4ZqEHJSZvt1sLbWIvi6ygU8MRwEq2Pe8cs1P
4BHgwVZy7yTbkDirTNpgDqAC3zNCdZsHzWwKBll8AzRBnK4rNHA3JdZX/FvOsXRf1A9k9T4aBQKN
v6GGquI/wqSOhUq0grUd6EryW320nF3OjnWbcWQCuyI1D+U4zsgszQEj3dyOvUeywts6IuFFijwJ
qpp2EErtD9kVfVa7OFJ/WQPuZgJnQmx1Pw1EtzZwD8sqzZsnGuHBeiaLsmB4q7JRD5rVWb6q3+al
nwbzyz7M6IAuSCN1shJTQd4Ve3IZYaF9NxGsE4HJidzMEynWIrYhvaki8SXd3FdrNHWw4l2dUFet
KhUwv31tWwEjQ8ZK5ONukSQXgat8UlPLUX2w10Mv3upZxw84yVTjp6NTiwXEcWfR2/yi8/1uOW5L
UB2O0euJMToMQzYEhmrFKkKhMwpU6xXdDKC2N/DmwgePACIogpy9pUQy9Tyvju2VDJWswkCUR8Bf
4S7caOWjm0YVZvMiD36XwUm+ZShOa3q8yoyQcZ9yXKoaoZUMXu+hPe4Qvp4u2SQjl4p472GwYPPh
qPFCYsOM/QbqBfhRdCZgnydvi7glyEEUrKGxvK8o8YgQxs5Ug3slt6NiVIUJr1jwdQtLma8a6PtG
3TIJ1UnkidcFvaGg9P98AjAe7XJwNNeZGXBXBnQ8aj2EYgEkFqx+XyzXeCiUOq+HtbyoxjjpIshH
98FUdoB+rklXUJWmmjdKjCEIT/Sm0t/YAS7lwuGyijMv5mQGqKm5idQCE5TEPXH3Lj5kG+2KhdJp
r5mKpXyXQJnTPll+8h3a0J3WhEIrzkO9fpJNAFF7syTxBTnW+vctfIxHDCmj0ZMmsxCEuXcuMLMS
tNrZlsFAnqNCX66CU3IuFdBqZoi6bgkcX5TntDz9eLN7Ro1lbWDZ/kpTOVi90TCsOznDxjXXMWZE
pOD2LybCXKbMRtK7/e34PK2/2ts7+wdUYSZRXAPfmf3jP9Cu42X3Hvq729422jTlCc18rxyr5JqA
iRJmmGo10AaU9cd3TJ3QwdjySjK6hKc2MreiNCIuK937edXOe2Z2ds0bHB7ORyfPKTpo3WH02Lj9
IvL1QsQaCsPJ2F49DbyN1+IioZtW2FDIZ2qzav4QiE4ECGNIL4GaimIHH3ikn8lDuHQG+MRSXkTh
BmzEjwJq2BRnCBEVcXv3FLChhZTSsR3ijAYw9t69MdjemqcUMB950V0OssKDmsuZfOM570/aBAR1
3U0ZgYRqi9TlwP40n1CXQ77ftMz/4FtLhuSMWtvjnrdI4536D0eX90VtOB4ZYjOdKJCMvLWnP6lu
0pg2aI9LnI05e8Sufi+SPZnZ6yCEVhUO8dbWpcqZWQ2lEGpzaZCz+BmAkGbKbO9VowNrPngIiIox
XyVROwb7eYUy6SGscz4/8315rGfr/47sCo739f4d95Ll1l1gpsnSAk2MH/QN30TWmIrwzYctXhyC
fD8s0PdXFsiH6rTYBBMYeQoghd4j25ENSoNrymtjQ7jOAguWaiTiSX7zM9RQCU9uBP6/daDYxH81
YnbMOaVy+bpfJFpgCXnzzkRs5XcSuc5/Eq+lQL1zeFxXQyt9UvYrmttmbIybyFSEX2uFrx4YQ4WF
+4cRxgWZG2T2UXmP/PLmAtmXuYlPuyL8mIyIuiBg+QzgaGVehTYlWHTegEes2Wh1k+oYIE+V0lys
zwR7VNHiEWW90CNdFHes8jsud7KZbL5C2KskQtepADYjcuvk7aEg7M8EwWiTnojxcVuO65FGtauS
Ac4ehvq1fnSUEyyqD3JKSraf20/NBLoSo/uc6jmGLTJnH5hHLNqQUcZ0LY/p3v39piRRLCgMzB+t
o1n61db+A5jbPBvKWnwMUdd9SLOsUW5SwpxJgdfH+SQ7oAC/2Bmzmi0BvrHHO17QQMujfNUx0QCE
BOCqRybtJMfxs66UXfLVP+TnBF0uWi53F3Q3IOUMNW4CUaPsihAZtTgMt3mXl9lvefpHOKQ18aoR
diHomnIPXF2GXaEqf7ILlK9KAGDzyLFWDqwp9Ijt6lTEVncZaJzsgQP2kUMj7Hzq5le1OZ7T1fGF
w7hQzQQC5ez7lx9utVaypQNVT7v4tTydgjYwtGeCbVWg8YK6JTjpYcdY8XAWn44gRjcPQtktMUAE
z+mgc61yDPdCgatK/jU7Dxbm93JttAoX1BoGe8WfuKXTCUgr5TgPSBK4KWjCNAxNdtmN91jTOJ2/
lKDhjhGZUaPeomww4CV8weYU3S93y3IDzY3bqjqf/2KUMANLjsCjCMiTYRIUomaez0kFRd7uR9vA
hFEiuBsgtHV4yyyI7YDrW10+4kiNLmFj89zZIKuFykbO2RQC5cKawS6NkOnsJqXyk7s/abpqt1p5
8faSoZZA0/RW+cLL9ceoywgwD0vcAEYWRyt1A6vu8SGpTo/nCA3rYTXXplUGbM3feZPrmu6tO1+K
sO3KLj7S6U9XWHlufnFUlUsgYJm0I5zyHwh8+8f4jyo/FMwiGOxXuDJxXhYixAMdTEAz5d9i4MoQ
XZ/pzNJCc0AHZXtDCuK0SNXjZTgwhOxzfPfzBDIKw9OwdQob5GWH/JebOM6EAbFFRucyX64btbNg
5J1oBtLDdk4/L7JTNL2/XLWoKqfIvI25I3f6q0sVVISe/B0KvtOoZxhEsLA6UAskWAzpvfgDtqsm
I2ei8rWJmtDa08xkx5vxjC3w3DBUi/oKmJZkj295uyAV982ca+aHMvL4M5OVhJrtNrRAVzHVDkXp
Zb7U5IuplfCMwf1mCcTtNghgvao4xAX+l6zFAKRm5RfAvRqkQG9DyE4wuccm4s+mBfKblaeQYpz0
QBpNTkvJte9JGQKee77JXQymJqHlyfvCNElYbHT8kcbC3/UKQCBatR38Jg5njOBUSKQfuwj18Seu
HGsPYhcrICWeKn7KwrwTTRTtDzMdFvRVuIRqGOMzxmBJQud+kfKYc9vjFl9CO2Dj4B7QB+WgWb8D
8yNHyKhFRZ5cm4IMuGPfYyQ/XgEe2hrN3nZLrwNQqiFtl4OGAqOLaHCnFRG+3erJrB+6eGANrHjl
03BBzD627VaxjtfxT2qfuez1ozjQjSkIKJIP3oM2EQwliht3IUvboHvUlwDISnVOpXcpV+TIv+gE
O9A2C21QBR6AeZ4RV3HeW6UwWngDhsB9JH+D1Ew/yXSyirvoAE3Ml7jZMK2Tm1FcRxZQ494brXzB
cbdo6XEarX0VuqQCJd1yfhrb6xPjKlkbSLNxJ9BbukV8vYnEYSZ3Xu1CozOt2jCQV2nzy3eWYhkl
82fk8n1WkalUSirv884NxaskiW58KBYFb+U78ytcuscuAFZm+Cqt6KMcaKTR9JNb7tx0nJuIluPq
6mOwcfFZfw45VGYqMUCQhzdSerFDdvj14lAJwZ2104KWTuoh754yIt6F/7oPM9KmETWYUtbJ2eah
+oOy3slyQ4Z0qfusdy/4ibYQEoSDT4oPG9meYQeY278aAkxhf1uenaFV+GNXsDGkFgCc3dJx7hMj
UmzMDX3tAyKQs/zMtT6yKDHvU692qmEaneK0X3Kc0qd0zFJ3JCZTcbE3+1lMU6mZII6YxjqvSIiA
gVQEYBZ74xtLzbL+x/iJQ42fSze8mSUl2Ue8XeHS+rRe27R9Nc3bGNAJpuuKoyyii7xPOHbjnrat
5fwxV2ET1oC3OU4OrGhcKFrj4JReNQJqX0wTaEh9V+5seEUOtDoS6EuGYQIxXsVup9SQzsNwCOBu
itD/ybfwKhcDRoQWk4sBvBkxwEXnDZOhqEEPc+tSIvmLOcklkf9DOKtaKK0GlVEFSyfnIW3iaZgu
UTG2QnatgbYEoOeQE/1nT9JXYAjC+hYNLSdbQC0pH3YoIC+nJMM8pf5+8qVOwGDckbvYZM6Unnk4
fDiul1ZRI0w/nNefbeSHvrZcOt905XtvPuoaq6tsQK5tVLAFZM1zku2sRYhB1LLFkyxk0j9sSLWR
nrGGmuFNOPGH1uoqRmNN2gMUfnTt8lMxKL3BSrK2AD44NtJ2aqvNRSZY+mAL2LznlTDg+th0/9hs
iTQpIN9X3tpv0/Dy7hW9BIDs1rG0FkscRFSLXNxLMKRtPrTF2Q0fRL3efxE7ZloRCheCl3SzGtXs
NuTeeaY/ESTVT5eLzr0VhPdhSzKHGzjfVdP98PAKE73Gywm98dxgFQ724l+DOMjY/a67oltemM4M
+59npn4z8SE9jbGUpF3QIZSe7T4Nbd8EumdKKVsULy7RU0zsOvX2o7SlXPoB6+cJvsSWRGzlc/nc
m8l81MJ/zqB/qX2TxA+QEQvi8fsGTZhMi/bsjjSq+f4BEtJtGh/9I11qAq302acLBdEaADNz814t
juwpgAhF+u1zeyKb8hCg70479cm8+Miz3VkRcVDCP3AGtpP8Vahz1P0mUaiA2YpALIIqLTNedriK
t6iMOCOLWdPmBciLqaX3+IPmh01Hpe1wNdKJTRimBEje0G8/k92v0IhNfMqfJtdJqzZzLxBYkw4q
pslkQUiYiCH3cbrLNAk2vHF7lZYnXQlYcNzmqKrohI+rLNnOGsJR9m5edssi9KNJbi3yAI727buN
94fN+4VSOyOrQDbndkORw+Wh3wDXVkaDh7yHINIdSmCgjWBnO3nd8Yu0F6a/Xnv57amjsXJ0hHZ6
Qb8LjDw6Jpe2HOimb2vGxYcx/xZ8gPuowUEFj0zy+iM4+QO3VS69AkdLprhA5ffsh4IEpQP/8FLN
/jv4ofoIapGTwStjitJOqCP8xx8jzrf1i8pHSgnvkLTYipTufIUwdEbtdYU7C0Z64UyviZEu49Hr
X4fsNOa0e7b6g5qh4dqC9zoIK4ca2AJ/M+0Qf/7O6n8C0x4MxKHt+HTgGJB//cTgQZ7LveYDy33M
H5sYU7bXsbbh0jUsjIySgylwHXJ+NWdF1Q2GdaxXr7edbq4I+UEwGss/6u4Q2ksAqJVpasblzS2o
0In/9Ng2AA1xCb5JjPMWw7nsE/mUAGikwM+qMVpiQeGB4g3UES1S2uQJB5KMLOOl4VSF3VHHgnN/
YG/rJ3d/tYWa/1L/1d9cxRsKDLqSdpdnmIcjQc5eOchxWVx0U0KVjXR7YlZNvw8Gin924Ap3FeNE
yVF3qDKPfSAOo2CHnj0Wngtpee64guuSUIZnjFtWBUkY9ocflysjKf2mQ7worrL2klRAKIYQj6b+
OyOAJij+rXm4ZxKXz155UubU7zqZYDJ00mOue7Y0IkxY8vbawBjJFZHkQ0pcDPyAcDfP1oYoH25v
bis/0yaywl78zuNeI2//ig6jGyuESkZXN0ISc9gShLlFO4bsoCqbdGVc37VRSETDfVOiwuetBnHD
dP5MEq9uuKlVutE31zNdUe3OvYv/9s9spp32K3wb9o4L0jwF6n52c2MdgmY3SDTrSBjZibHumRYc
qKELdM+qvtpeKkrrjWdGgjYYiif7Bi7q6/6a9F8nR8wRWSrgomjDgJ30I2gQg9pUN3DqCCTmvtup
KLTAmTKQOjUVgsXtuxCEuLZoG+EMjY8vcoyGIxFZtsznsSWVly3GF33RCco4p6pCNhqTVdhqOZX3
+BfdqJqBIMVMVC0KypU17IK65VksU6jQ8+5+23RTEAuLzP6/YOG0PTzK9SNL2ZrGpFx8ciJsg+9/
vNMYkzlgurYifduVpV/KoF+EH04HyJ0+J0nzV7VUoAl4832pKcnM4nOZZj4NP7JOA6IyYALVQXhC
hkPibgEwcfA/SIdS6ixBmFc8guNp7Yu0O9ZvAMYg70wV88Efl1n4OGCuTW+S8zbmUJAFeCU7JLr6
bTAwJlHsIeBno0M3QgZ+/ILU6hJ+pFRvglgltMDQCZ0/5IUXj5pFc7Dzn6ym1hmnoorijp/VKOFG
phQ/d55vEUsOA4JQoGzmqlrFGV0GYr9kPP2z+/cljnyfRZfYwNDo7gAn4Y418EnVR72GO9MHYWKW
FJjzXcbzHQdNBnmmlzYn+TiO76g0q5856GNa3QWB/OEtXtFbKnyOghLKAKBPK//cyFXBXadUULxn
Escw7k1big1oGcFeJpnx6ySWN/5Khz2wbQV+ms84f1mNiARsfkc55iEO8FNZmz7XfShMscDCR7p0
flvnMOI6KlpoB+BY2DHVDA1nQovJHY9ibZzurnPUXdn8DqXf/sQpQHkZ8ElP8wIleYM+GDUdrBft
tqwV39YDZIw1zZCGDnThfv8uJQ8eyS3+7c0D1+koZu86IraEo4kjgncdxfZzFstxOLZMRrfc158E
UzAT0HnfCn8d2zG8Z6Zs1ppc4RwABK9eWG8pRHeLquiKJV6NRMD7XwCJxGSnu1vrtdkdBg0CfXdK
Qb0KNBcrbdQ4MQx+fjcUJ+0V219vu5APeXJH6v6b+BqdqHxPdKaPxjKY++cShcPVUz28WnpN34sF
ijAZDK0qdz/qJe3wQOye/ZBiMrfUUMxb7TzlBLpL6HU6tV+2lf2XPMZygI1+CvluVje2xUk+ql2W
jBo+a3zNxGTNr6Ao3L3UVv4EtsYUtgW4hy0xsw2v6mK4gquzuGKYTzjQT4agUmIg2NAQrgGPDZH0
XM0upZFP8s1GOM9i32ttc2SQoAKofkKS8SOdWihHylbnP1FZXFnmIffA9XXPkIqdNa8Dohp2fcU3
dO6ppzJ5JwOq7ny37+BYCaJm853OF0B/Sk/4Q3ntjavQzMMFKNbvfV1YXlvN/T3gqX62Hoql+deA
dhva6FfCV1TNsbgZ3xUTq5WZElXRRFtiM5JctNCAriO71XMaWug4dI/GSKBHsuuNuCDrp62dD0wk
7DdUbNTimbxMkw+iEjT6F7lEZt3FekhwOdxRbQD/Om4HDS3dT9HLHXCTMwtazVkBU40INgnjsZ+r
e6UCUxcqrKgDCuzJhijOyGeuhAcTCIBHea1UPdjWptCcnsfgWVJq9+6SMp7bFDLYXSrbTd08tPH7
GI3gkzo5rPZ8gd229uufP23oyeGDvFRZr8p7mVywJnqWBzKB+DoiNaS+uMMftwqDhRDMFbnsy3gz
lZzq243aGvu4wmLK5LxMz4RlR7swvgclN1kskuouDRmOKh8qm0rUFXMXWPtqoVAkcGgj/LfvswUE
wVqawtCurJvQbNvJdQnZTLTinWEv0/fZ8R3xZ/EBajEuB22SvoRNp4Bf6HojRSWdlpDIN7xcP1XR
AOGAWc9+24HHaQbjaN83NsA3DPuOcCh2MuGKNQqu8qNOKcN5N7f4iBFJkmP6LHYmj9cDLr2pI5rB
cp4nxfqr9w0Gq1WKUP81+mGajWtTc9iGshAfStGzNJTblcdkOIh+YfAkLfX38Fo7K/KesDgmk464
4SOQA4G7PToAZAu9cTeOszywymqgEp3LXaRWZlCiOenJBxQrcItFY4mFEA/fj3FWdG43SW7A9D/M
cJP/peyEISHDWAIOFdxS4A+fo/R1rOTrcEqs3K0eZgPZfcT8HiUiREP384oERvdft9hpc6Jb5/cR
MsG47x92RS8L709sIBN19HOKtXPaKbTChhLKBCSntdDAzrG2NtNoaCfgLnW0PUY9LmlXVNsyhKAN
q0iIpAwp/57FGgc8uLOnS0QTUzNPrIAUnsKT+pFmBrut2JwLgDZmzqX01BGyb4kFtDh76wHrYPvC
hpvwS86vK950P30Xxrr1sZj9eoqEPA8RijzMZLzIKAJmzSp25LwkDTg3hBrUabf1wJfzy7QlANzP
KzjNy6FNiXEjzMK4HJAv57gfwsPIctGEn+9r1DEwKQhqdpXxY9Zl+t8AtSilGdLzMNGEw8//TpJ+
3WZuZov34Dvlqk5Or3+FQrCcmqLjWuXHArx5nW29623iSM4oP6fprSqL3z+xSj7HuQg5zuF00M7C
+Zr2edWi5fg1YChh1sqZmgjjQ4nLySx3v6TGUaw7mUIZpavxmic0RPmaT5Yr5c6HGGyy/HPNEjFt
J46Y/ngftH7MwzUEKydF9t+A7p+N1m+Hbnw8BUH8NoIvJSB8+w99uacYwrC6h10lHjq9E51pbEk2
zPQJLhFckdYfV3kTVmSRC1WmzB1bBKLf4fCVWR82auGgnFMp8ya29onFQVUVegK9XlhVWJKnQtKM
WzhqM3tufnZpDxzNGn0rWuG3YbeBHwjUgTDjjBBKr9//HFfjh7DDg6fTcwjCVyVl31AsGw+wouGs
d/dNZFdYq1VfpEfwUm1usHY5WaHLOdxUHKwvEJcwvCmkBm0kgTwPYMcEr1+V/vsCXpXuu8xCpHR7
DmDFgXtO/KjxfUNpE5ZgowI/B5ahFELZYin5b76QyOR6WJQJFDedaDGOAnVEAvJynpl30aGEl2KP
eAsEVPXgpGirj0OlXh0t+sdkIibwjRzocp7dBsaXr5LVrDNVnaH4tdDaYotQzxBKkMcdsNvtI6Q5
pfl01CHuKUKrRbHii+N2AB5FAdM15RaqHTtw4chIB1DAKvK4M+Dl02M23rGW+Km0AElPqyoz0PtW
x5PNxzXimlTa0s6KPy3D4t54qRUJIDRo6L7taDh4rFz2q0EUA3JLOwENLKkbTPPtwlUHUEwSHhFB
tuFHkH5zPt9zkloTKYXWaMOqccz7XA/pAjGlZmS3Uy/62F+fED3TvKPFBss2lovkvxPLt1p6U5iz
xd3O7bPvThX4Wq0+ZpydeHKbtjyBtMeie3CN18yqegfOJK2MbTjSJ+aHyXreLH5F+4ba4VeszXoy
QGc3cj6JR8OLkw1kRH34rMu8MM1MMKLqeWk9VWSzX2ERw4cS5usVK3ScFXg33TwPJ8joxkFBAM1F
/QQk2lW3P0GZ7qZVj4mpWK2dwC34n0OQsamHALEQu6s6ygE4VR8FoNQV8KGWmBwZNf98n/l5l8cU
voBtnFfE1ZG80h5u+CkxdrJB3b2K8BPN0jcpzuNDe4IP1l3Vw0t6CZtF2TYhJylO6D8jDzy/hfzp
1iAfEP4BgS9PbAM7HpMNh4COW+RNM5T0vesF/kmkPS1JCfQL4/fm8OcfHhb4BWtDLCtljrL4/0hC
sBNXQ5jkL/8DQbb9CFkaHnx1ToUJ0rALe9+jt3M0ra+/DPRFEIT1sn/4TMW7IQW8cTKeti5MIlyh
AaT+PxfmlytdV9M4kjsbF+ldJ2EYQ7VditWASEUjpXTNraIs1plpXt+Gzsz8F2wHloGb8EHDLMBV
+/bruEnhI0cV0fvqyQenyUuIgSK0Ye3HOgFXra0yiTtZ3ZeBoGlLOhOKZ65glEODFayKJdVu0MBe
NJHohfb4OF9qr2ISdut3qg9wwU5ms3DPF11dYq4jv46CjjOEuaQ0/NbfefFKOV+v73HeKqAb5iUJ
F7/q/cijFRpaK/15oW2HMrnKj2zpOO+vx7FaeVWN04OQKrL9T3KRThpzc+wi7rddlCeSS1S/Pzq2
+mjlFyq7TKNSZFGCbMAWGslxsETcTxPxblZC/FXX+Eabem3grbOE2ruAKyq+auuiQNMgzb9W90D1
GYCtr7o9QSJAnKY2gHSNWqZew8CR8Ir45CZQMJ6DQRYRgY4zozYkAF9gtQW4/kdrQew3iTre61G2
qjDqFNcm21wTYCAKqA7974Un8S564gIQ4rsyJC6DcRoi10x8rzWhuIP6IsnPxY6v7wskq6e7cYLx
wSEPvJqvXTfesQwP7hfOtiB+ADejxMK3LICpAV5bQUINy91PgyAmWAENcooPQGYX+YaWxTViK1sB
WanqgdJfq/HJ2xWWMEoadH7raHD9zkujfSygi9FNBdbd43Fzi3rTJueDinRuIKl3Tme7WBxxkf/i
VsORwkzQf0P5MfAMnO+FR+3BR+5HFxosQLC3uJtXWCe136ZUKpYOZe53qdIXvG6UncmSK7SC13rd
bKLH2NazGGGhxVHQUfe09kWynCFNv833izOwlpniSNWfFcALEAa/60rqmhq2nly2wZXR3DuMh72K
tzBLocSueby/H/lCriOb9MRp+huc6wNSc25s/39Ps4Nds1ewbfUDoEyB0IUE13+otab+RxyPBeGL
7MWTGhwovnAZNvqa5sFIoVFE7w84R1IssOQSoaz/UMec++ebN5BG8e9SzXn2olwWwv5z00eipwWU
NTUEgCEginm9wW69iG3yc872Hlx/0PGeIS5LtUP/cp+HkUhtyyGO3ckUMp6PpXWINcUAp045CNZp
Vrhtz9Q07tCA2QgKL1F2/zwIGxzN0B3KnnqRh9VZOyfKI8X61IaZrUdEGw3eGykYjF3xaJdhowLv
nsuWDw1lEjtXUaTCZpKAbRgJD0UvzNQ0eVR/9GY80MW9ugE1bdi6Z+GR5AvZEYSLxMleOLQ80Te1
n3QInOdmwHqZZcDSOYmaVQDX5aPYhPmVF0631XVdIVkCanDMwUa/uA0oY/O/HKiptYCmFSX4M6ev
kpeZu1TeI2eZOpvu8P/1ZqhQzSryND2IFoKPnWOm9078cnoVkWeXj8CbTZ9+5x5UFoJbICW98yts
zvUViWnXNbi3F4KwPlebCCDWOXusBveS1nPufqDDA038aPJo0k+LI2YQqCndgRW+Oi0h5ZXeteMc
RGBobI9V/taG1B3Fnp2AoTc13tENTza9aE+/16nr8an6Uwb3IVKPNwwHI7RS2OStPirf5f1XwniJ
974Vtip4/7Fa+UailFUCiW7PN9vwuHTRKE0Fl41d2tIlK7OwIOKGbP1ce9X7ReX/QjT4otPohbqM
IQjYwjealSH9EP57zdXKkjXGNK2qRPKUe+Ja81JYWJIVbsa3BuTeMze2KAj6bxV2wYkaYbJ6ZCdp
+r20p33lutKLDTThIPINq/zPuXCef/hLMx/pp3AJM5tSLOIrdKfFE9Gc7aZEaQpcOLzjbbrP5763
gIuvpvnr2pM3/8K8jvEiiFZgIrF5Wb8W3NpyQV7mU3aEn5VJkdgKuJS4TLxAs94H62jfyASRHsh8
ipu6RwD5JvuJs3SC2PVC44dTD7gPWU9Rv/yXHpc3GnChjnaMBemFpXziQJGeWCK8MrfAkYM2QwnO
66g8eoEGYZhoQJ75SvA9hwAa11DHf0zFoUshi3xepyDxWikUELOnuDzp9xlVlVPzn9jZV9CSzL1+
wl3k3NtGiPdYLA+ers1KpriTnTrMkrcc581DWRoZ5eqR0vKR6BB2fpocXqrBz41/gWYVOxd8Ux7I
QvEsDxPBK2DXxp9DhrNH4HkQ1HqVeCnYRPTcKAg4716T/5ou8D+oP7s5I9e9nxVxfzb3bm6KazcO
pw+MF/QA0XDskQmmK966sZMKFhTFTnGF06fSbwYMWgaW6f/aF4zoe5sEypoDwzk7jQESgJEBa3GX
rfk9jlBJuXB8w2xP8TgIV47uikNC2GsjXzQ9JCi7hQU//ZFEJzfnp30EuLbndQA2UO5+B1KzLFIR
qaxK+PKOcK7gF9cizBl9+ZPUK0NSD2M9/ICIClQ1uhXFHYN4YaIThn94ObhR3IRlHtVN9OgxwzBQ
zpvwJ1VX0GhUGLpEvO9ChkK6MB8DvCPdNDP2y8vwKnYYtHRFzHKZov+8H849618eqmajtw0Y6GJA
1QhU4fW48h0g1SCXBa0XxvQowCFK6eu61if/UFptCHy/vzLa2kKHwJ7bbck0GXNYBpCVAaLLE2d2
nM8oAjPccfi0pnT/ww5Q320R5V/HU8qrtgiXdu3G9qrQQryHv2XR3gFYhN9vvk8Ur8yGE0MrNbir
QdczEAtqb3vkxBym6Hm0HwACbhTY/dk7GKlLfgjwBQyy193fYPqfwpRtxbr16uR2Wyycsq3KNkQW
lDduHlY87B4DsBukAq1/KDjpnMk+fs6Trqi+e2237yQuQV/Cw+Xqo7WMJlg2coMl61wOXF5/58as
/Xu0/X+Ghe4+TrH3Xd/mn0xycXpZ+e1DCfFWnym/M6o8nQUPFJYXfy5d2un+fIYy+d5okFgtU9z0
ztFhGjgA2iT4FIxrCGholszVbwI260GcKgqkPHgO3EQEbiK55QokTGnDyUyLG+QjktSCaojbzVdS
/OMIysJ15fGBkIU7S4wpXYeyKGe8hmc5Zds6Zg07s0KKZ0a+TkAR6FaSvpU8dRL8mxkqfwuT27Zv
GpB82Y8UYVV6Vvb3Nyk3WsahZQ46x4vieYLiXaIwXgn1MLeKvSpR3SCWvdebqDbnhqQjoe9he6HC
hM1tTbKMAkFCVsz0ZPma9449GqUSdjdS1QY84A85rH2a6i7akH4g37ldFD5AtZGik8b2EdgN1hEM
koYmlYRSiQVa2w3cl2sdhdJHDc1soJ5s2jLBtZOQH1rjU49k8g6MQYCHgYinf5VsPJ3QfnvXxEps
K+cQLiIX2uu0+V01jLEaIW2PJyJHjelJi9zy7OTHwJdm0C8fhQxJfbYmWULnEeWRmIHB1WAKs4EF
bVCutSEzsY7smVrpKoj+jdoYs2WbjGbvQVwWqH5SUy5AnDpiXIsSH9imM7Sep6TTGuLulClfHTpL
lIMbxpELzAV58TmfZ5+Ul87ZMpXtMRhrKffZG/IAotz1d7439WGTLCtQ5pmxXOVWncB73EQo+bwc
H/8MK/vORh8T/0Ad4FpZnyx7lh5tGyFlyKauSGhkELqpXyUMC/pX1o9qyfBZGFiODcqBZdShckxi
t9/XbEhVHgpwie1A+ccKYxk9MSSExrQUxDqaltkmybNhxVZkwAh04DhFbgD5R4WDuzGG4UyhgPQL
bV2bFnvA9hVG3FKu+4rhqB46hA4DjpMYtz/OGaGmEvWNd/7AwQ5S8XrOuUC75cTGNrUaPzDJ8NGM
Xuv7Cy//zREWU68uyAdFnNCMrhBEH2Jdkwsv1gUQtXQjRhNUQiXworD0pxu7BfuFQi/ZJL5/5UrN
XD2MfSTdtlYSk71IfnIFjzD/xORJLqwxB1C5f/fmr//ewlnOqhr8F2evXFZ8kp82Y04BJpF6RTmu
4VwCg4oCtTI3sHQ8L4v2kgIlN8qy68LtuuRtk09wCVCNLqk1a5khOUOgVu59cxIA7SKUMEc6ZRVq
Z5qPVJDYfI7buOKHBaxxYN0hkfsc0GpOBxDmb6O1LY4OogKPILMlwyXII3KF6pyQr8CoE7uM9o7b
B62/EI9XvEYm00Z3EEXyeEP0t/fTetVSPd38OOzm2nr3k2Uroywi5r+asT52oGSL8MM3H0TS71Ky
KZvscDyPGXzvIGMs5OcWgHjFUzUEl07synD6upo7CMqIiZUpmfPVvO+wuEPNt0Azipi+bWDaRIZa
LQX36rjD9BC1PLxntsGHwsHdv/XLCD+MUJQYfftocE3cOvjn1bNSKkW4cssL5Go+vEYSy+Iyff0D
kST2dPrZ8iOQM5zukJDuET2hcMCSe34Vkg02kY7oexYsF8MXzTI9HwaCIR5ZCQ2Kt0RDG2SWpQ19
5Vg23qPhLFmvjt4Ng2pST/WMdxzzVi8323jcLOHbvgHT+T8alOz8GTV42CwnjiGh5eAr8StwfG9W
LeqR0yfCqwzFR9Fgi6hL3XVbJdqD3aPz68IkKW74+zCKApeBSzux5Ou8/xtsQMzxqjUfglulaktb
jufVp3SdjKRD6ZwUh8XtA+C4ZAhT/K6bNjIxgqG4xrpg042L+wjx5UspJHzJkWgkTa2NztKzJ7Zv
l4aQwdtBuOP/x05Ao0v/pXuOP+6z6VNgKpYmBSr7CzubxNz4yULtrC3mWjQWZNASEXSY/lkj7AXG
ap9NftF9JB4QrVBATmzVubEwfce8thsHuLIkclYQ/dpEzzgHD4qkBmU664+J4kOSInr06e9Gc12w
v+XHC/aMuiM4fdHOy9hd5rZ/AiD0wMWMpws7zsuiUV7gi66t7IudMg28eraul4bZi+E6PFhZgINF
eFOJvmJMzOXpK1GS8Ma81h9sTVtLKmAONPFROva8HeSBTNNikVybz1McGOrUbgWNe546D93jhXJN
T6UtsIhpAuN6NB2YZCJ4fIQFHiKmkHrustz9hdNNksutHYEaB+iFhIknL5Ku4aIdXREIq6VLV8of
2R+LiYvmSiuiJiZCXcXdsD5aiNAPLTTYwE7/92utO9gqL3PqmvWbwRZ8XmLK1Jms1e+CQeV6Sdxa
M+4+y2sbYkM93n7LU3g6UDOqutkDbnCu+wV2vhLZKHFSL2I8ScfQ6klNG17PfMmLmlc9tV7650b6
qHGC6UchI8UfBOx09tuU1jw9AMJ1Ed5xeymEQ2PfP4MJ0wCaHZdSszQzOxjjhiRzmMA0RNZ6YeZy
LQ0yml6X774umXSaAiP3Yd9+wrtDX8CiSYksoj0og9KIFo8n4eTtSZZrYctKA0CP+p6QUQnbZdHx
x5QBIv8ne8qjI/yUtRIUGKcXYdbVaYweHVkMlkKSAY9YdJSHwCk+qpfuOYZAunlgM53yQ1Cr02g+
qtR2Req0xLlSxhejnleAyUdjJ43AxrcCGtayp9mzIxhxJuT4frTC6mk79XafDpH1wipCxht4Pay8
xfhV9XA4hVSGuXxdVk/O5pglUyUImtQ6xAsHHE+7rKvmnTPnwxySDkGFq/pbNY8i6cfcckChf6Q0
EIonQeXNig3bHb3HLf/eJ/EGCtp/V7OezVKaMBbg66bYVipVN8kuZb03e/2C4KZ8mrvOOsoq6xqu
tjexCyUHdGVdFCl3OFFSnHGjY0E+pqW88UOJoFiD6o27JCquhPIvhIvcJy3ARvMKvNONEBhIwzWj
qDSBsetu6o7GycGT92MrVY4uo8hvN6YeJpSZvbwqMusRQHiSw8QyHefpZXsmZsFymEldd079PfoL
OTyGt+6RWr8LYWYQYBW9KsOir+seYBql+ikrsxrs4gY4DL7ZEq2TSdEcabQhGKFxv+ZeUeojH2Bw
zNBEb+e2AQ8uWtmGgIGbS+zGyBTIpMKlxa2TD6z1ZU8qe/b/lE8oPGCIX/DHZLHJ6g6dAnMCkCJ0
PVbJYl55UjTbmQDt4xjGgdhQdMIfxKyGFNZ0IoGTvjXxWvngmE8FqKbIvPSjGarl0sWthzoA0iiF
sp1leWlPB2tn+SkP3lPhvyvybWdd7kwtSRN4BJ//sbMWBiwoYZCscC5Er+uC4GDe9bHObq0jb60e
iWPYsAEdC/J1zpkZ6I7nojjQYU2oI0ueHrY93Xk7B4eb/RpFJXyWSh7o/1hFljrUxIlBIjhkR0ns
2Lm+1Cr+T9G/CipYwRHlERkEdDgTUygpIGd1HHF4xBX28Pk/QALObYs+1yAf7+IU9QsOi5j+UhRA
nHXpMlKSAto4OxUGxPKPh9GfrljWCh723LCsRfHY34rP2dKxmHcz/FGffWN1YTn3ysVX0gynzSxf
xJ4eCElIAR82rFAXFDDfmjXxObLVGl6Dl8377XGksmVQuhPmOAF3+E/3PcaTCtEKFL9sjEtIdFGg
oFmNXV+IPQi4WWyLUar+BnoXMwhIhuqTBfLOi+v7vmzUzSBcTCpGHOFUn8LFxh21r59J/s49W4LM
jhUgvdTYJjFQXZPDm7rmtCjdRHwjRBcPuvbtufvlOXiVuAT0gkUANV/ObEGMXRL0HeyETVYouTm8
gvPfmguH0Y8b2tK7RaGrhB7uKTPmbx4k8uJXYqk5UKMIWYql6cdM9rjy2YZGkNL+Y8DznZRjZv3v
to2x/EaSZUNAZ5b9lDvDeuTn0yPTo0BNNpdZXWbFeB3csOUZ4zw+O0iWZppx57dMCvG7d/WygId7
eVn6ZSUxlvCA3S69pX/K8j93sifRDYMVr0v09nnYgFfMwPNVRFBqU2eQw6hsXmC/CULiQmjURGhj
q6gPgKtIz3eqobstIg1VfdXLmcK/1e5j12oj5YdvCRRGXmMcKTyRnfiwygA53KVtZu2tfMggJnLb
6cHzQkidmmn3WiCsQBSoWm2MtycGwvcrF+GW81P/PlnBIllvBHD1hV2NHiChMDMgmjkBbxT4siZJ
4kFqn9PT2FFzuqKQU79nv1VvpDmBNCM93UiLXzByR6BzXFkERu3c1jgHFXdfMvCqDlS2wbqxNu9d
A/qVVl4jHKS7zBhuosPSBo6qapEZYembDqs3Fd5KUlz/RxcoMJO6PvUpBoAlemd2jfBuN7UN8lze
8pZOn+TIGciBa0BdWvP62i1VeaIUbcHnz3gxbC0PKND2dFMZD065Q8jfofGWY1Hd4wef0q+rN4Z+
DKXSIsJTVy1tsOmJzP3XC+FSAEC0y76Zku+RTI5rzPoiIq975J2WNasw14uIN2IUMwCs8BPrbqwt
zBy/s7X55FNua+9sG0SohctsqIAXq3w1HD/zd3L51l7GrrCHt1vRAyqLyUM5IEtysDJHzckAZmKe
85kB24WN7hJA1kWr+g6MOpPWow3oW6wzDuzT4xlmJuWg1XKoCG9uuDENFAx6xq9CeyuoysYp0kok
G0pUbGXmBkZXyW+oyiU+8TpZ6RyOn1f81fU+kWyMLSpJT343TnT9LnXujaSdjyo3V1OxS1nqWJJE
0rX0KCq97hD9GirCK1jvaGSU1JI20PoLreNVcFrc6nX5+8HWHvFG4FBf65HGABlmUHow0xwTTw5H
wBtiTDVvyddRT8+H6yZfHybEh0l4eoh40mWq7Dqd3biHb+Z+SYhXPwtQckd7hfpNAql86B8t4ebq
1lzyOTU7W43ZbgkJt5Q3uyQYguhooZjzmrQGfiWzGJ1Znro3AUl0N7qqvKeU2paQBYeNBey9SLd4
hKuE8qeXbyGj5N6l/ceMgakFMp+ss97tdPi6b3BTtvUoOnPQRNQXMORN37Fwkng8eQu96CBzRj/b
hd8cc+Ca7Rdqr4lwsrMwbBpo1tCH+RVKELLuhhG+HDoU7/DZ40s5yl5FHsWEiBzymjHf/+r1z8ll
9E0+U871Eny5bCB222CST3wT5w+2sbQtCkYae5R+hQZ/duRRPkpQC3wusNFm+hTurQt5IarQqsu8
Cy7Y7SjqbzpgQ4Mi6Dx8/iK/N57TwGbUo9oU4fMlTv6sZTneEnnH/H3FFOqfGnaxWYwFE6/eRCOw
ScTRlEO+J3On9Y/26hB7kBGPHbgsDUH7f4vIDvDmO/n9uYHQvJhAkbLdWojhUk8SBuaEUK6QLLHy
CeoLrIuI6AGDPNTWkUI9SBQIC0umHWwlXSdmlo+S5ctgXthjEu/Jdp5qpDHJGJm0bUQ1lg0OX6kM
cm+B62aOtY59kNIzQ8YzZ4mX3LZWd5IjejHKbeNpFCBcMEnsc+cOtYY7dEUaU4SjcMYPeuic55w+
GFKXrDIoY2yEtZ0K+Al7jvrD6UlEaJbjcwZleG0ii7dhQRGZxRLmaqHbAVr6j0LQg9Il4BpQ+YYX
9pdovu2WEwHCzOYmNwueh++iEHWcrCOo7Km58l2wi8JLUvdDQ6B9CDjS2iWguc6ScPKST/sqRCx/
cdm0Yp+/5gJ9lP7lvJQAatw5rt6ZCxYL3RvBwgKWDHL2prlrUoTRzWdBykstynzeyiFvb30bk07X
WLnRTjCiiQ4kaT6HGkDpPyiy/QlcKw1LTuKy9RUtHkQmIYPIY8CBBCO44bO0Z+kWKNJgXQCjaoWl
v9AR0Pz6l+P4cPbZmDIF0SY3hySLmVknRQ5PpMjJJ2VbQTvV0AnILE/OUgj+NQuj2cxU5OXjDTMS
6vbc//gdC1txIXhDTUwGEUE7E1FG9oBRnMAJBVcT3OQqCfoXZGQLYy/hUlQOO77mj/LJ+K3C5I/S
+zYr74YIfFQslenZ6eyTJ5q81cDEZgavp9jH+g62KKc5i0fOQ4PQ4nHyFHp4dcwJx09ZMWkRnPXO
tkOxeDbpWGp285s9TFsqkVMfVFMwpPiMrAYpo8OWPllbQjL+Rlhp7epNczdQYgThzQAzmDIxDeWW
6tmhBH8lWSwSBJS3rfjPsL3vlbbA8CqxmpqWmdgUjhnJXLiYM2Zy+QJkudsJV6OKcmfJ3Fy8qMfi
+ZUHfaD4e36j25lTKAsUtQHm4HpgcI9une1i6JgnX+9d5etQmb8wntOXsiSB3GlJ8Yhv6RpOAYgn
Fqpl2fEENiNTa3gsZPsU9tyGDYJHnMdghxTuJJAKjhwgtyPk+ipWRe1aCOIWt2QuLi6uUWLsueQS
D22NzD/T4UOfp0ghgNFtLjh9TMX5TXf5d9K0DtP1ZUagbIuzsTP8TwQQREI60kYGQzkiOaNKLwxJ
xypxMUzs3wwHqv/NeYPLjKiLClqGjZo4r73Zru0n6BTIZ5QcU9LLzUBrqQAOtthbuS9dC/6FbW6l
1gpURbwmfSpsyZqDXOedGcfYjPMXul/+uCAoIEqnhxwM74S7blEol7g2Rp3jRjkYKOH2EESrNe8/
TsuGHq3x149FwllrkkTaloKNB5KBg21J6moTliVklZw0CTbL9WWrJH6GLKiG/jPuJI7LflxgqTCL
GRPEnGVIqWaS15gn2fon5mpDQ6YzCENZJai2PbZxYj0TUETZhqX92I3PV8vgZgkOrxYO4rFvlBV6
yF5OmMVS7tgS7RzsBW7ThXmIpyLT+s4ezJd8OJh4c56fNhU/wBtqNlpTXe2BrKKqr/kaNQIac3MX
ISmBK7rV+pKc++A57H27k9fNrButhfwkuwO1qLBqyFaBbTQYQtGwmqXb4GIisHNeQrmVFMC8Z25/
FeCpqfVXxL2ZjBjmF3icFfCTq5eS7VDiWxQ/T1hrTSnt3TaK/nFVSX3N5TXgDvrZAe5IyGyWBDuq
ca+7FMI1alP1LwhSlL0Q4+zvvQi6f9U2kEVG99Hd0YYEHG418H0jqjGlLr36GkLljytpt0ObWC49
zXcY5rnzxDKSUGjwGYjarC/3nRO66D7qExX5xaI+ht3Lpj02CsXHK+UzhN2P50f8i50yQUAP1lE6
8e51/ozi8UsXBEj7ZEjblhRlhnI37UGSIjRg5YjSCLgTKczXiyiHxJ8OYkwRag+x60OrqBeOKerf
GqK5AbY56J3PtQ1jJyAa8QMuUvPDUnZnLK+rVm0EaqfjPWT/Lw/h9JLl3noxePY+MAJiieUw0tL+
TTuRN9kCe7M/a9sPswI6OPjRmK2m3HJv6E3L11VEhwTwPHp14iUtY2cjHOc2kgSRJl0j3NOgEWth
sjFM2iBab0V02NH8mbVY2xVWYDJ6nofiocN0zAojX+3XCJVny6ZCcFxsVPN/xSbiWzw4zJnM7ktR
3LdujKXHtfdbGiADj0RzDJK6iQ8SrtSivFzOmOetBAdazCAyCuSgyvseG6hXeh13J1O1eddxdw9x
7S+OvOR0b46UQ4g+ai2l8pK1USkv7RelYtJ5zxkOcMSP4wDxyS2QrXmJdaY+lph/Hr5qXcXdRo6B
BpJZKp4x+KJhazMzDY35oUMk50qiiEFIqQ3Jdrti8AVZNIcL98gtX7BVx8DdIsuIR927Q+Rlv0rH
BnVxNCSUd4JN4ZQNnKGFSA8hw9yMo3/or3SsdKYcV/WTXAFxdUFV6dtizFMVb01PQGP/bnkTBDF5
4M7ZAO6nhGRoMc1dNZyiutHzikZRGyvzXAJfm0CWgt1JKAZYX+u2dBchkZxDVAOZFUwwHHQhUD0S
uP1k/8d7Hm/qFI/yTPRSHHbbKZZ5EoqECjgt5MI4hAhvXA7zvzYbLXuWw2/kzJ7b/bMiJGGbic7t
BjV0B6h06ArrW3/n2sPpQGm1EUvZIikYaaIb5kia3rGimvgFMevMqWoO6ppwyDs0rksOatPXqjXZ
HPFndUepLW3Lo7xO/Dt8wFyfJwGFetubwLzor1RrrYxDsOijKFjacxPZN7LtLQjTSlY4daALhuQw
6IKyH9jWMri5MDZ496cRNuAKOHqzI1CY4O3ycaGpmDNGgeYvoltpkslNa/jTGMoCyC1AHF5be2Bn
kylVOy+5rsf917ijCs21eZT00FFBU+AcdFxzLPu6hpVzQj72tsc+8UxZETyX69nmOs4Q9f4wDZCI
dCIHzo5+qBi4j4ttE3OOwnugcu2laoiI3UYalvR7z0IZjCkG45ScQSVkU9iH1tQ+4CSyiu2ICgSW
vTFaLXfr5ilZ1PBEeC+T5H6+6kQED7kafxdRnMVWTXMDilXWHobQmH2e3SvpE2sZmkWv1wpbnp6x
Wc8KJaipHkowyql4VLMBxYoSaHJca168PW8tx64atWEwwbF7G1Nvujp1qbXcySbqF4FSPo+Dz8ou
GBK+RTf7Hnjgpudgs0s8y4/WlRXkaLAOpLeFYqhFa6bM6D449De44rAWKpDBzgld9ncCaCVc8d4r
GKjA+28DjhPQdDqj8UBPrGPf65ZUrloYTYNcdNLwoM0+L1Lq0ULwmedYg467PTd+6iEt1iasM2Lw
I6mIs2wzHvjHAG9fxvcbBSOXn+AE4Bj4rCwMEAPqwJfJNBZK65wwl6WBGCku7LV6dZqUsYii2fO8
vtgx5GOF231v98ghvw/Z53FIGg4MO2GJhdHgQfrRU/vHGU3v6uCg5WHhfB1eoFmm4BPVr8Az99WS
k+AXVqEPh4mrxSvha0D4Ac7RdtNERTtqar7py5stB/Mxgy8tXadmr8hItT+fPwCUu1ZdFxGFIkT2
nnkkI9n0ZPM+N3yOzC4sONPvfDKufdKv41nLtGyhkZ33X63BkPSYd0UCm0ng9sXdYlZQrm/i7VS8
NvuaciLvf9civ7Ttzh+yDSmWiDYrrGfsezgP2AXWCxudB7Jlw9PVin1H9naPINOasRNiWvKlqVN7
2TUhIfwyrPEORUrbV9GYmH82jgBkfDbgUs4i24l7IdKOfJ1QURTOxSNX2HKqUvG87A1mwqq6w/tl
2BRk4xBGuRbTbXcRzQv+EdqjlvPPvu4eq9sbpnKCypGFgMHnu5pqdmPqOmdOCbyPbjp1iibCdzDY
nM06Q62sp0En/EmosmhrC6+5VvpleZUgmH/TOQ6fRGGSGYODLDtk2QWkLXMicBWiIzNxBpfptgZn
IiV6VFqPlKC6UpBpLrg1XOkafJwSDdVKn8ix+0gZ1nowyoldryDYck1t4bRyK1/nmaXRUe7G4dRC
n1gUaqp0Iamornt+AAiKP6Fl4WwUJZnSytawlZqRYd8eXltD0F1aAJEuGkHXn1oNa61Ahddt13b9
kGBFDocR+esxsFnNaENpgXLd74NMY26nATAil4YImLNEwdZutpUP2IuF/ar2lQs+o7Fn/VRQ9kca
JnuLDBiaggku1Uk1MIyLOJqv4EGw4DLBahGbvMPXRD3wr7fxNJzcXDKm0wqCmOU2jGZoTfcNjZLa
tZWmLEogXAG/oddFuFXKvz4dGFc1Vk0PKy+26pBtDWPQQsMAHwJlAD88jCNIeOqnFEtwKMterkwz
bkQuodtelm8nb5VW7HJdd7YK1lrJ4zoV81PU/soO6wtJ8JbnHdcMnmBDegENlxV11ReoXorM7ho2
pmgEdbf42e5qlFE+8CrGrPJTliVeffxDLZgoT7xLcgaAVXAPfi5LVQ2VL0fm/AnxWo21P8AVXigD
MPWtOCxhHGMUgKREUoWe4lOscQUaj6hhteqfAY0nm92rbWVeIDbuw64lfMeZYrF4HjLheNxyyT1p
tQxj8HK4RGW7+CU+WetKp+j4UTEAZNasg9+ZsVwa2b14+r6hb6i4RZ2iCn/kIIMr2iNcwGNk4OSg
rBJfah1JXuogTUIPa9L1hMm8S9id2SzJef/gY4Kjg1CjqFL9iOmccrlFFduj5qhlN9+1owy8r5hY
qKuKPJlN6R56IF19unExSwuzIzloXXwPMwWUJUasQuNU7G3vgQAJ6JflTnSkiDeVqh+GpbkQ+nhc
MjbSneJ7zxy/5el+/M1WVhU/isQrLGD1uOaFWIB3iymF/xdaXJXUkMHHSpdyiI/JFd0pshCgsixG
Zm9KeeekTewOZ6eiFMI1fC/oo5TXw/b02To+eE990/oseujLtFZYtoRqgQFH0g6pjH2s39DZCAjJ
OFZ2zDYFVQkATqpgUp6b8dqfuP02nYd5M3UtOJphvgSZgUT/Lws8peJYydW/RJmaakSPZilYGVxD
pFINuqlxCbzXbogDZH4lfJP5CnM8xog+SAVtMqHirmemuwHN42E+kRpeTBaNm/DK3IpFUMxM9TJ6
eL3lttXjpuqt4i1m+0s2CJ/YPtOYkMm/Sz6ObrE8XEzz0foRkgVfYQS+VUaWjPDpRh+sUdvMbcKk
f6hXLKlmtlIuQIcssmp1zV+co3574R/si++cPdgkHUjlptK4reJD4jtEyhz1sIUW8xEHRnP0q7Lh
/+MRD65iF15/9Aps1crGHdoLPe7os4Vkk60LUJDAM6ATouEVo+F+qHSYTIVTrNu8G9ksll+Rn5eg
BS0MxvSCE++wyXnY3OyDbx/HGZKEntehjW6LRAoAIcY/3OCjzxwl3WC5vuOB2036XbCOPQXUkVOm
69DaoCORj/qBcrez4xcUhOeazo2VIhvLPGouTHGJXj+u3YxFUwVmn7v0Xde20Vd8mU1k3hBsZLTc
1go7wy3nHSz2ThstvtV6+UMm5JdIFW6e8wzpRri4ah+WbffkMrki37o0+Vdpopd/kmLk3CVjK5sc
U6hMgt4guw2rB3Y9JczMdyfN0oVAsU8ULxaLLcwtSD6/ZCZw+oe7WHTVq/+xW83IwCHgpKjKP/8E
yMuHxsxsVTxM2J43rlBgguZYaT1+MFQTfGrHtdZsHeb9R+JqxJa7aE6r2/Op+GipFba+0AbHPuW0
vgXxgjS8AAaoXewXRe6JOmKygda5IpBbGB07y2Wf2PB2sTqxqb/QsbW0xSOSHtqt/S4RyBDdLjXO
FjFZrLPNMg0GSXbO3qBLH7DPNVhfxWdzvws7EQb33VzUCybXxZlaAjnH7CfXGVVdJlUkvtMKbZaK
rO1fSfh1VdbFQvr+J2jaj1REJjbqazwvukituZDZgTyQMXJDGAYJhwFl6VTCumFni21f8Vh7RjqR
O597mI16LIJm7VXIs+IdHCYMiaR6PXLchMRYtqTQrwzaKmiU7S9IgT58v4EPkd4x3Cak/uLwroh7
VcG+9qYhehMsRue3wwIe3gF8H7uTp0XRKjHEpXr6rLYCgUyPrbJU1WrW3On4eq80o9V/be/p40/A
RYwX1iaMglteD6VOvUsv+/joYRxFoDWHw0el3sVDXH1DV8XJTfZ7ZpK2JQ4TEJ0PYCmWmu6geE3G
/P8Hrlr5xG0CIeZQyeOqEPnntfqhoKLvWeaJsrhoy3qMUrc1ra0vhUXrXhJw4ptyZUhjY3rSHa/L
BpVlHSOPUIYmnlKXYVy/L15gIjIyca+OO7EIIyErw+Sl54sE0mfoG+s/+LWKBNQg9ApCvt16VcLC
tRITyRU7nUvrFxieZqBeYXJpuZSBy3WDTYhKyj4QsUbd/muR1KBBDILyoyx9I03Twfx5k2rP75ds
ATODST/4b+IM7TO35nfRPRm9uxSF1Ebr8fsZil02sHdfSnwWZES2tWuOio7fZ5le2fFj1plLz7FP
Nk1Yfj+mLn/xVJtc1p5paqmxvgpkn2Zo28sceTNMkNGLX7RC6C/7wxjjOQ20gebzIoFt+uWlUx70
5NyVPswU3Nzjx4I0E96jVKALFlGlV0dv8HdOT5qfxt5pcfWflhjah9WZLA92V58/sF9Yi0vH+Ujn
4D02K6P/kFKGeiRPtenvCK2IYU42AffNrqCKv1oHnfnWXJY3OxN7/uoVXuq3QZbRtXIsTQ05JKj2
3zqltfhUvT7pi8BDNPstlXgX9Wp2mk0B/9IxZUCQAbstwcTWtwFSlv+r4NAG1FbZNXilvebn4lQU
emAbSbtsiboF7R7n5hW+4Iek6pRuGhSIle9nfvAMisFTChfWlETfKMwf6mUVb/ZV7KwdcGtRSprq
H9VHcAePtpi+VfDiHBHONr6r2Idp6bZLb87xI9f0uI7UlzB5jPGSBC+1RqJfA26XL1gYs7zMtOSg
CCGopqD1TC58pyQMLe/MeYGZeACeMfoxSx9D8XHGHfZv4WXydRGW6t8HJUYDhrSJGSzqiFNP2Ojc
L0vNX9xaKfWJIUvqbMQhk91jHXnBozgvTWK8XWivqATBEylqbJTK6VJLn3+5N3aY54rQpqlgUEW9
Yb+GmSVDDv2SLi+EQMHmEj/CYR8xZwFZV3C7M4tDvutvtDg4zgw5BCGrV3GvD1li+We99Sz8XRJU
kZQoUEIqtlhjPaI0D36l7sesV2FpwzgerKpIZ4ACaTVyVC/nFuX1LjoCkQgTxg8oaNzvkaR9H5VF
CW1F00fGeF56l7ExNY6fa9r3Sg5gERI7FpEIY0FmIqEhuJ3UzlKxP+pNC9+kh8xuo6NmfxYqoY9L
GyBCpZ4JWNn/D0Z4hNZvefgrwjWp/wu0ybS9KqhMYSv9C7kwm0LkkSCCE1izjzkUaNCDwEeXD+xT
e5NpdXVTbOLa59CYQMTyGG7QGatkpw4KkgAms2sEDBQ4RWH4AyDVQObEn9SUgCdlEXCHoOCARFa5
HYtbJ5LPEtvCouwQhWylfoPiKIWthpsMBkVD6RfnIvhHWROsNZ03YW5xAXIaZzooNO1oEifZEWvj
dfjR4kFZIXWEjUq66AZ2ctXVJn6L4ItWsDJZR9URbwsSaWSqpk10gwOrLW18TVwsrL8dN1HhOArk
HMq0/gPSxck5qO9lW47ZIYir5qZMfl7ahLrt9Cl13Rwt4KFxcYRpgHn3oXKlEREBEDB/98JewzN6
sQBns5dzxUJkp2dYO9Q4jFBHC/eap8FB1Isa5okgQVZel0lq6qqxc/iujzsVZ8+vxacsrFT726/U
xcajkneDN2nwG7MdbqI33CDhnxwTU2Tq3+VcOuqzA1YdkaUeq7ikrpJ+agogG19cs4xbBXBMaE7E
o0VRQUos9mHoo0MRABctcs2K5wM1SaGl5CzaqAmSPQ7sd03PiUqQy6MWx0dubQW3YbeWUaSaOlmb
hgPCJnE7teYTNC5HzG8xYwrjiNNOJ9N46m8mU/Dmt21o4RO9tJ8/297y26CNR8t+/Nevmftp8MYI
bk/7vOeUEFVTT1hqqKR4VU0iHcBfrlKhx6SR7b/t6aSIjjkDRZUp7ID5bugnidfQBdSCD2cxH/Fk
+MmXpb7Wy/zaUHByZmJVE/vWuglXL5sYLJ70JVr6D6DLSph/8EQ91tW2n5cNqy37cc0n9xb9+btH
NYRr558+b4d1QVju8bTmtlnm/qr9uHwNROhGklK9DDCzp90LGQbsykIR+QAfZiq/U1HdiNpIt4ga
iCzxS4OBFzscWMylK50C0WXzgVnNSI/uqEbCGV+CSnEdIX7isHL7JiHsKzg0oy+rJeApDaGI2+bq
WGtnFZ15iVSR/aiQuCibdQxij/0svDbC6luQceXbjBtrmIILaeukp9H0zGgCljNbCWEGDDUC03Ph
e5c4VUWsg3I4wSeiIBBJuw5+wXbOd59+J/XkZblruylyAS4THWh8OzB5L/2S5AdkEDZcRMnRI9rt
OnMtM5XznG5IE6ivUAo1aKjXwPb3oUYDM7fxj8DTL/GvxhhRam+65Eh/UjZ800pdzlUxL8r1/WuG
qw4nbheXCX0Hn+MB6QW8VEAuMS3ok4H1NQT/7z96IgzJLFDhzG/zVLuUKoGn0kf88MhBJmw7zZrR
LTUeL2naRWaVFOmYc9LmyIlF8YTZ4mEBS3/4kH1h3UshZGVJ74QtRWtXjp5FcqPpqVUxJUDaNE8/
gzFhFZouzuFDnudU1VyfoTXWRL5ZQ2MclGpaCGh8OJxqBqA3+hk4/s0o5v7/CoL5pwMCMFDK91bt
h9WVYmZfZjK6d4gFPWlMcDyMJI8JcezF69mtYeMIGwq8uhgGMEiSAG3B7CT5AQKP7zZbLde+eDHm
myWAN8UNeXeU/eEAAKhaWQkW5qcgbDc4lnRWy1uDgi3GmqEtClNQ31Ut5+swW6yjbAGd1YejteJK
uM9ta3sHTO5vuJNfKGwhrujpdqbmL/4ndYMGkDnL9zIMN3+Z61AeU/vVjP6ie8jId0HqSjV91kai
uDDDkcKLmekcv9AornNKZAVPsHQ80tGwvnVGlvXHeJ1iqXZf5BucTZgq12QBck1kYSvpUf5pqZko
i6TAepFWT/X7ped1mDzEL17EbygCB8ObpN3qVQf9UsJdqIXp1n2TxRGSZuI4sN92SOf/8oLGSnAh
bhVxj2TEsxoYCnUOPyKawjHf+gSpg5OAcC06Gsr1ziBVolM2xm3KkKfRYdv17DoYugTMA0s4ywcF
xyA4+n7vglCd9VrlK4W+EqldSwrC7+AY7YNZZtnnY00g4mgkBmEEh0g5rsCWOOHPzGjDjRgltCb9
CikJVAxOQD4pCZ+643iGhHpKCtt2RQWoARyJuRzJPIoctCOivR64wzSI7N3jn7/1pmy4jCmVVVSz
n+Hw+mTStTbVX9305veWgtz/rDRnvt1C/SwOtW/1GbyRl5p6nYQCXEkPoUbLAKcoSsUMsYLZYgCI
HJ/tgjPWT7TaNC0o3NJ6kMxU6AfqEm9TbR/2ErA+xL10JXNttob+dnvdEUC7TIXLxyERuktby+FD
8Ll0oqDkacZjikgT767eZelLMClHj4tb5V3MeGPjlKIWPxh/jrdkA8q+s9HzxSYsuVbYa7Ig2SCh
Wu9GKWfI2IQh2ADwkTiOmOM7lfFZdyNAAfx3AeD7W8JUHmZo0pYjfdqThos75yEIp9rzc2E0iZma
TAxaxnkfgtcIVWVtMCX3dgGFKB+Gw1MjK2QgdxAB0sB3hSlxwWnbOCN7jJ87b3Xr70FAVD6FLHNP
PUvyIh/E6QE5BmT4AAiXoP48sQ4/fbwiWjnYznRwBxB3DU8B2zEbvVFipDrVT66ys9yc3iMiIMex
pqf7h3gpWZihENVCALPLWYysJq8w26kNuCITSab3pcGApiUyKWq4K/pF5o7ptRvo/uT//MlPUztd
FJBe/R7aBi0aQLN4nSTVpXLRY8Xw7VXjILmLny/n7VA9ugNEm7SFsXXw8YOc+1y1M/3MU1QBnzGX
I+4NvJDt6X6eD9SV3pKAnPvRwaPssB8z5ShQpTcxW0DIWsmafHBHJV7r9OShMgthX3mxCnph5r/5
LZNOarKATJEDVapQuVAG7UIVuJTyga20nSxgKjOXd3Yr1zThZvlp+ldmKlNW/eLztMlUGa+QNmq9
3aoirMkLtyaFuZBPfRJ5EKiDmFPnB38XhtR9vVp7a1/wCjIQH69uzcbvh9O/ukIADuRbyBuwc9dY
ialOoHVwI8x6EOaedcRNjlC99v5UAPwX03CPrLN/1eFyNYGUwf8UeE9nH1sj1YM8sQiO9IMmGYcT
QMcwXj0+g8xCQ+6UdDLGbIm9najDic50ppEG9EksXpCM0avaf43oBjUozHoXcNYmbBA/rPF1D9e1
vRDC8SxDc91IXxSxpjCmXwAEbVtL1oySsQkWGFJREEdVnfUE6Pys5mrUrymRPVw+Uqm82rctefWH
dQRUtNJSyVTzok3d0hSBbrDnbFSAZIECG1Jk/7/URXrSXLFqNdIeuyFDMLZfejk9JOiCgt32poVj
9c2a96SXQa3GwsP4ABIEvtHV9G2/N1CwR3YNG/UPoIDJ9KuuUnSJSQfm+i42ouLOiWeZmIHaD6yY
1miOz158VJdcvn70xk6b/cJeWUGWw7LNlgmzoICZfODOVBzUYggTzrJMym8Aq9OeoI2pP1Pib1O7
smz0sQlHPrmj0lOmkcIOuMAA8fzfMrANluPkSbm8dSuCaJ1BR+x9utbiE7NBWMjFqDLxg18Fa3nT
LeZqM1z9NLMI8LyVzDWdzsVdJ7uzYML1puZ+IyXOjlS0qizWZ45s3JcmA2KraWdsONg8TTtTLr1h
ySdmmRRY2hDfn8yOy9RgJZPEyIMVd50KM3/+1bxm67R/Trb0Eck1+XBZ4E6ia15o4JWZjDc8OhLs
iFUEJ4dWsufBOYlMa/s6jlC6juea0BIkb4wOYdJWme4x+VL+MPezb9nXoUJbkmP+4XyIjYtZNYzI
La/VDuAx9q5oRrEG8DkiUQ9Xo361a6PU9cAYBx9vPt6N5FJs0PUB7Yulu5TtTteA/yqsWtsjJjiL
kvTYXsCHuXxnn9q1m295EccAccb4mjmYCKs9jcRYEuld9ufES5IGbqXywDjNqKtHcEQ8Jl24QiHJ
O2oR9CHp7rjun3t23y26DLIXfQugUQ8yv/nHr3ftVzb0yVl40TZXxUZQRsI3VAZA8nOabpWQgkTy
sSSx0ooulNz14MorjwVztmo5HDsjInRIoivfDpAjVlkSYGkDzavNiOlQVW6IGBY6QakuhJCdYG/2
0Wdn4gLZUPvUeyMZORDgmfuH4ZZJJvp9KhIddmQM55fRhj7AzJdDOm6IxGBMt5cmR+8LdfrFhnuP
H9aFum42+p/8zpny5+fv3yO0IbcTFCi3VjrMouWQczi4RsbbcbLgGX3mOIZKME+2Ac82bP+8wIPI
nFbBCZnQURHhcVADqOLLIihBgHdGHAw+/pETK/2Artys+Z4yThcQ5IuJu9464vS/vqH1pFQSuOC2
K9unMNQTId5MXnQYFORjs8EzSbF6OsDXwdUPhAhrrw0gGyTrfBgm0DfuOA4J0YP6dl8uYI0BSVZR
BBmo6BhUez4uPMpicL/u5QZgfqNbAstxCWu5kmiPpzf7v1lcg+XTiWJz2B0+XAFfmngMLT9kWeev
jGgjZ3hAxFDM4E7wa5dg+uQ6R/Cxr4X1pylrDOTKtmjzR0FmS3hWck04jlpQIT0i5rHNE85LNgcW
OYJ8010wee5HNJkmW5rm7GhucL3kcCNGGmeaZgHA3oZY+rZ8N2BCHaNQcTjK9kWsBDsEO5UlQCT8
3WmqKkkX/Duqooat+SD1qg7W8OK5ZZG6GZ6E89GMPMG4nkatT1WeK4gb6tNy2jdA6yXkNeUnPuQ5
9w8WJJNqM0cvDYvTltdAa8GcSKcn1n9aBymRle606RMEQAwEGrEwLYk8iG8cuk2ERc6Z4olyFT9Y
s5MEhK/GLL9CBKWJm2nPlZ/qe20X0cOtnkPg++LSUkIzH6U3ZNmsMsi8l7wuw+C0zZBmhe0GfPy/
66006Y9HEeLgve5cSZpD94lT/wV5uZvyqfjTDPlJDTYwHMmcc7UvmZxGBFfj9PZ01I8FqXOYOENs
GqFEJTD2whQfFJYw0kKwUvRE9GjERJyyIwsepB44Yw2vfb+ZTY/ZgjViTTqia7vrm1jOTqawYpdo
Wn5NtqTJTpRxqhsgwQd7DOGGUqD5jodidmg2gpk31mnVujrsqCCojF/MTDfw6nS8fFOlwZmqYDOS
cs5ltLiipz1jGQ5qy5AZMPI7SibJsZiHe8YFQ3IfbViVzmUzGOjBbzMBI2kAqu8NA5bQMvKSYYxw
x16czLBOjLy/6du7/o8FtnxjTUC/pMMOWExznrfiU7IYYCXevOMsMwBx10Wcg5lXrf/NDpyKJwl5
ozttHYdmH1MHgk7Q+Ft9xLRWzMKQleczRP9Z+icSsKOrWYi4Ifx1rE5szQGR6uW/Y5wNWj8814K8
6ttIVW2iuzBu0+IOHl0MutMo4SXxSOjGq+UOnzUGBiPMLJoOvfbQWffOUWYRulm+w9rRXgevlpOC
IYCsYnDmaBtjGGCXCTWivzCOFWEGC2IbOYMBNpaWQBqNLZQ/gm/yX2G8OWy1b+3LlJ/n6otN30DS
dEShWQrrj0MqaRAFgplppdBFqJHEHS+sXP7F7E/Xvojw3VP5mpW4rbG8iIlquUNvZiWXG74hGXph
h2sgp0Em/oxzAq7QXP0dnwMCo2BpBN60HWyPxh2inKMcO/1eakh1xt6icAaoWnrIvp53btwIKq0A
skwvcqqMIc6QJxReejEzz+QxRsNQJD3aiCO++sNoJNOCr+bq40dKccg5Scjfz8eBwPrjdcTynVht
PaCeTpemFWCJdqj4FSb0mARYXnwMjogg2bRDELcqeFrY3ZjRc8HSV2rFZpmdavIgPQB3bwf6xWmd
YL6veI1R83qDM57Lb/zZEPykJI+EWRS1nyWevtmQWOPd6jXaTMnwj9JQeDGCfo5Tcy6inNpB03H9
7iwgTquf9O/1TAOAY5wH75eiJqyGzYbJPjS3lsZdCi/ALa5grZhMmbpbBn7oco3Hqob+Z9oBdS+m
95Tj888CD5THRZ3DX13H9bbkIeLB22v8scQFqKQB6XtDSvx2zYH78OPStn+bGMl4+jpgirAHfHQv
FlgonaBmzJrvLl72QL1CdXEn0eHnlY/XKq+AhfzdvqBbmuPnv8xVO7X/Rt8jKQ9zbh16gifOxV58
vaoDJAfiwTBg4abNffz80F+biHW2BErKQ8yHcHXPYuGcU4/2vdj1WvPOx4vg2he9zGpPakCTyuJM
s0rbyTWsphcXqrhLax6rZnT6T+Ou5A15YvVGYEYdxWvgD+JJocsxre1YHhclnHHJd3g9/5yCnFM3
PJoFAYwJXlMIXLHdeWGE3awqZI2Jei+Ko8tu1mrby/QJkJqBpPx38QDxNKJpgBCQf/nL7N40QjqQ
XlEc7wyrpQ7Nx8tKy1IVrDl19E/ShEPaOl99aGTc0RO7e9xQ89L5tryAxa2fICnbRhaUdIZwYnFo
B6W4BzVYfvOXVNd6CdqtaYxCKPkkp0/cjOW0f4Zt2RRdFDYVg2DwPyjjBnhLLZF3g7QB4iM/vSqj
JFyc4j1LPjs3FjoxfuugRQVzKbyNp4NEf75hD+6zVt4Oy0sRxX3vssyaj2b6glwNtl0U66qTzd3g
YsQiSCn+a1eaLXQro9x7zaXcqjuRemI0G6YyqfiPm5nNPKN3ZnZYUFHDzPok8rNx7ZydLW24iT6s
GXJc2xLwXF+2o2i5rGv/EFapiyKuAegJK92RkujjboybUKPUPSuUpnVtju0iX1sUKb/XP1xJI+db
RrdP7HFFy5KL0L0C2GLiGNEXIwOQN9zUVx2d5x2yA630zbR+XOuISw+hYREU3yttE7lqzZ98MAxx
JyKjctPYeytRPFzsVC32scoLVFpGyavhAGBp2LIIofQJnVM5xW2DMHE3czdJVF+uZHg1BGZ/dH31
tattU2frtnwzG2QBRbllHE9lcJXivqlBBm4/REQtHCEBb5vB/kS/umyioaNX0iHv5bxzLftaTczZ
IwKH/S6RPa7GFCI7pm/avf0P6mwREIi+lPa8Sl7b5tBKEiu3MKME7bVhPYlrIFmuPueJ1QoIAIUF
rrxeUKGF3j+4x/OhJkgUI1Jil2qK5afPSVKhWRdPdsj56wPDctea4y8uqbX77LSB0oleulnSJEBz
D9NByY9AgDG5Q6HO5MgC2KEGdsy5QjjFPfGuiD2skuI2UgZzHqmhyXaq7Es7Mkqa7bVsb/W7DaPc
nKZm/53qqRMG7MPewC9O6GuP/gBs5A+BmwmquODlQ67so3p/Jd2RvwSiGPoruP2XlyOcmCg7Wn8g
hgqDOBoY5dXY0vOgQ3aPvjyeOL8sHls4gx4/wHdXylrFHIe3PUE/5GcJv8BIFJdWTV/vhYOwcTQc
4QedpUbUnRH6Vr9RnSI/ww4h3y/lKc2saC5iXMqX4Z2RjbS1xFEyywX0XFzETF0Nht5UHR0rJErd
kIu/EnwXu5YpGB83qK3K1OQj4BnbCB37ChWEc9pBSSG0xJzqG17vhflb216lukCAcg5MBK5VbNKG
QMqvycABagAQaCoLcJ7nSkT0/3BvqVYlG+SH3sHBo3vT18msIS67Im71Dhp95wSFsNC3L095zwTC
T4KhYVKXZvW1BBy2CM5kvLEIxzlncnJwITdYto3BgLyvk9M+N5EaHmaiI1iqJrfFvERXqlF54xfW
8GiU210TMBcYsAwYBys6yfoyAIZdNIDuf56w5NKeV0ASpUcKqmdX5dVps/ojTVB6IHNGcEo5kzhm
TGzlEnNFCcTXdd4NzctwTqBQne18r5WqN7Mdp7Ff9oc6qYFI3jYXhyU4QaW45PdWLFYsGEggCZHF
NlD5twPwpLRyau+sSDMeI2BSmx0GRwjp0yqkpzmnc5rRs4wMLHTHNEAkLZTc9h/5hLrkGv4VEMye
Ivb4NdPlreGAcN445WtYOsFpPT8DMyKgjSAuAjoguMhBExb728ZzSJ8fh2RwgRvL8YwYN+Q3G8Dq
SAffjFUFPS3gkyolIKx9x/5DJ5AvNdKYqekrD286F5TSonV+B8dLhR2Wsym+qW3IY6dJntLe0CcY
hpGWdEz4nL/zpYStN1naX1MTB4UsOB8L5vN9yzzXp7557U718ez6BKTC6AoAayBSFma5gCXWM/FM
L3eBCyxSX6pT/4upfcyVvLgjW+fD+gO5wxN3yvbd4JRyEHUXBmyT3wX0m2wavtQzrHVdjhjEESRU
YsDHEpyLgENr1bjlBld0KUJryhEdlGpANEp4S+KaIns2j+Y8VBksKOOVjmAJMo/rFS4DINxX5r/u
wJ5y7/832KBkVeBmB99Ie+KfKYRxKXqSwdz1ND6pzZ96uGDHTnc/exUvtn5OINMI0CqQiOEcyY62
z2HNUVWQ+94d2gHHOwB4Qq4Th7/fRW00WGsF3xC6VtsxB01aXYTrO2JfqH1dnAsyDBD1EpyKoIbb
Zt/NYCSIYoBprjARYyQYMTL5aBHgdDjDzVAiTsdapc0WjZItz5qOWzXq1RR9x6Smy3JDiU4qxPxc
ct/9ejv4QdwgW74OEFNWZDHnGq5NBgepiYUYUxd/g+cEP6sAuiqS75P6wXnOvIjHIDz2kcpdrx8q
jgmYySVIT/UTpdwa40Cmd8TJwtNw7lnXuIxll3m7m7YM0NY6FpjHPc/s8Qns4644Gyd+ZaglRECs
1rna4GaGqDqCgOqmJTpXcuLW6dgiYTlteXAofNpb9bt5kju/PHv4Amy63a8jdrofGBfK6TyTOVkf
ELE9H0yKmw1FWHVHtpNIcsTE0+gQ8RoSMaC4GN+l2ncIlhVAk2fAqqammxooPx3MwM+1P+76Kl0u
PoB/9sAv/1dUX0TKQW33eQr2eDLiYF4iQhruQM+aM44aOdODLyG2dFNO3oF5/SLf4670DIf74t3u
eG1SCjqnsYWkUeuhVlcsqT/ibACTSsq+a6VsmS/+O/9PlgIHO7vW+XlXF0kL+HVhxN4GGt2puRhy
QVkwBzC1pEuvIFxgV17iCt599V4C+6VwYZtDJM4AJijRg3qwsqMxzAqEt1QoiI4UB+H6JI0QyHqc
LERdeuEBzrd0LzO25HgiQWYgX1tYf4dATFXDGWMprWjsFeXUl0MSkxGxT9rL3svqgz2EFaWoj99X
UJ7Z3LbEOKOcZ9QTFBTU/svzVSXpBT12zpyMFQ/Nr2cyBverOLYzhF+sJbwKG508NhLcDl4bTE3v
TMnQT1tgnLznSr4WHrIHtqVHifZeKA3vzhaSC79p1iGz5RjisC5s3Of4joZWgdUwTHElr5q78p+B
DNiowcB6PfLUSZP5FvhWxNDJpD0vH/k7wNkJRbn6Wruym47W+40KCko4c3rpp5q8VQMPp7SLaR4h
/4qNIgPIOKPQudt+H9QUNzAeQwOKTMHTa42aHiHuGMPa9yDcL517dKE107oW0pCJ8okr1iJA/9kc
+bGjgtFQpp+5gpEEWfhynCrDVUThMj7mwVXkJ37AiIgsh47iPiaBmyBMWrBQwfuSplais0lfg3lM
ALotrI4czVE6MM7Nhx3OW0E3mB55Nsla4ApVK7NhB9a1A6U+J/Qu1L7ecxR2Mus7bQhYKtdHTv6M
KFj3IMhb8ecdbNrEAJS9vxd/ytM4TL0wd3IqXsQTb046pfHCesywVL8VgfBkxBPm0mlFBcS7eSeh
2ski/d24JOXUuKks965jolDS2WVYupEvguKnJ4nJSdLDfAW7Ql9h43vpYxNNBChFacrll4J3/yDd
m0SZEH4aGWDJ/zyWSMRVE4BuMeMXYzrEzxVMzdGLywKkemmCCPTrSZhRIeHq6kXoO94Oja+b/hx2
M9jusyXTX15puKlaQ5y9Am89GrPbqvvQlGps/6TWfsf+QQ7+qGssHdEhNn7/jjcL+tbBGE1DRHPp
dsuPLBmyqMSYmntQ5WwBbc9Vi+kcWRFXlW0DP/e++51R676KV7Y7NTTrwgqdrHsD5lpPSXScwLQF
BLharTcVP7MzVYfJfrs3gGIxmlrvA+B9DK704StQG7o2ikmYtie3GREWHGpR2pxnamFYqeAgz1/5
WHaZDpdd40rlpE0adWRkSq/EDEtHh8EV3laKMPMkU9/pQl5kvVYGjTAbVBrtIYGTvsY5xdpR8wtX
AWop/vFVcv1KUi/tTvlPg7zJeKB1nb6GPD/a3znzDUdLFz5yzZwv4J5ZNIX/V+vUDPSchT28BHhn
mNHR+1eQ2Gn6TBM7mCUkT1fI8ogIw8fzyzHsbCQLP/77jB4MRD77OdeTB30STS2t481CdB7CBLEt
HjCfo668xJLlev2JJ5KYm1vuPjgyCRmWHPsfv+HuWwnibowNMyONu3rkf7ykQ+plBPSYeH7FlUjp
R/vLXjmf6+R44hQdhQZYqz8SN4KZuHjFSIvsdok1c4Sqr5NYf+U/n2ktmnOMUXCJMbczMau2FVVM
cYlKsdpZ8NISXc21dOhlO8C0S3+oPhHEvWIb9MnDtyfBRigAFTyy8MwWHA8HDuQyOw72VnelOFFx
ESr99eXDVQPomxs28tyqc3AJCRSFKpOUn369epCnc5YY/VpC5kEAEMwLhLdf3fDTlVX+eVE79xI8
lN3UO/1tRIjkn6lITlP8jfuhWvKRuaZHajd//LJAcm9st8XQoP93g8iruZWkMzZNun7gbyWNF2dg
po/4LT/UoiJL2L9SeLEbePwsboKLtVpZCQhG/b4N7hPLSReL2xto+75OR+Nuj7kq+iQpwaegVT6/
XRDZtyHGdZCy14nw3JaECIiN1vpzJO2uENJh7WFlGxGNpFhuvBtkxDjv7czyqlLnlFPup0R73Hhg
5qFWySaL8AOvpzTT3oSt1bLmou+3+p36CYFEtZbltvlLHAA3ro8703cGrVie8wad5i0uRfs4+Pjd
0F2hc1m9R1/wvpA4cVSl+pmh1R5NjbYV99F6rJUut76ccQBqHoJjq1uFMUG3bpa4R3luRx4r7Bkv
2Ap6AtBl5Zq7m0Zk5F+FtNrsnB7vXTPRuauG0LQUHTP2eSK6ge2DqgyCKgTxxSD9IFLM+fZpRUTu
b1UnjrUP30Fp0ObDc5fueEbIYYnOk6xovRRzTO4EcVaFjv86n12dxaZyTj5pdnkSkz/YpvnmRZch
C4PbEaRF+e+DrY/qwb5GoaZQpVL6y6yO5I+TyfvDMQv33OdptLC2Mhebfb1ILSZ2VUlQmUyYXExq
71izgMXC2feKfhfHfA8Txno48OS84VRijzDH7moGfCJqM8zAH4KPn5Q+P0oxaeXUuPXH06DmlXl5
gSc0W7JEjQjEs0Ks9O/yGdgegvBqmaDjAxdePYloBMzPOtAxbFhLx5VR2kTlnaz90n/qR3uBqXW6
b+QA9VMG8AP1QsnHxSVUQNRIwvo7MTW5zNpVcRrMlDNvsyXhv2Y2HRcd4nR07sPtUx5dzPyH+QBP
nYnHDaeX8P2ZjyShcFcZnxcKycmCkUUzx8GzMS9SRtVn7yg0vNVkiZqbcDCMFkcxKPxJpxcmUfHV
/XOOsLGbT8V2eHM79YfZ84TVSHQLcAQMzFlTZUsuXSj7WbJYCHDR5td1jzBM0mGADRfce4Mz0Dt0
m1bxDERtrIz+PNWNFiSwe9pWNTKVtkvO3KW/6rNbhH+rFEcNoWX8MIrny4YhmqB1GshK04xhOGaB
pZdlKkUYZS1UtYjEk7SVoncrXqxsOlS2xKCG7QH/sfBSDnvaPNZjiJlB+c7oIPMhkETYFQqrsitY
/l3ikfqlm9zJdfzlTX8Fwb7hhNL1yodl82iZzQgfdzCghkK15hZP2ODEevJfFqXiIVBWzcg3lkWJ
2/bXoTS2J82fl0GD01gyfFt77URUumlbefBfk51VntFBU5F4kCYwXph8O1TmhVBBvQwtUabtyg4O
W/TBdlvtaWx/RPQ3aAUe/n+Ez6JXdiIHGWJREqhKslydl8j60jy7Au1tdNIOksscWL/ioBxws+e4
aBRWRV8tSu3NiQzyBXsDOvPKPFNTCSN6WL21E/I8xovjKtuNLyBenJb5QjJVf4oOokA6Q2j+wI7u
fTkH7lnMv5fr2zxxpL5xCZtdNAW+KHCb7Buzko3n+qJKKD0NsZJdp30/Em88vigG59+P+WaKiiEi
rRGY7YgGrIG73ZWU3Q96b3ci33bcU9SVPFQTbwkUvl6R0WdO+gj7iD8yR+b5LPN7yuh5Hhdign6s
3B9V/LB2mzwahnF4bmixbQStxHY5Nmy+K8bTVP4E0ZdOXr4RfRo4qocwkz/VzsLWoy4N62xN55rt
KGU3fPX7QUWCV2Wm13xZm6ZnWKmqMP0h++xQfU5N7IAxVZybpa+olQlrx4d0ksXd35nUdDW4SM9G
R4IqpRX3JJIT5erxfItoqP+Ar9SASXv3VGTmghC7aLaUsH1jgyHkPPBG5Ii7hEHspGqR6wzmvsTr
oJfNadHV95t+BGKTj8ATfE0UEo+0nJ8fPiPu6xAz2pZKBiKrydP64K846r13ZM18tWdCNQIcPAlJ
Qp7zYlNIxbc5moBjZEecC+sSvUQ1areZAVRtc5km/k64GzOD+lG88SdCI4uebnQrAmpbTSDVJv0Y
q49C9/lkJUP9Hp/BenQJ9XyVbfKfeO5j2uQ8OnhJV61LYFNIRPuTWIgOP9DdnWOOijm4RxBWwDUy
E7KDgSaZFM3BxxVw3M2wIH+bHfPmJRTceCEdllrD4ojiYmbKiCYwT+x9qVJRK83flrahl0TzmSDn
lHcX3Urn50HugMKTvUvbUzeSp7tGMoe3lc9x8/s4ZmkoNfsfmNJ9gp8gSkduzd0jLVHHqO/+dm4n
LZTqZdPvzytTGgoPHg90C13y9HkVZmYnWjJm+GyCzdNcAMwpA28f/6Gz5mlHfT8r+0FMzF0L/ErE
wKEoVSC+ZS0aCYekEFyl4GDcazq6xuEqqpoayEpXPYw5V5rs1AJCJUo5kaYXMVlBQDS42a45o92Y
dCYaPmbHI2XY7UFlOWsyOfFZtBfQs0edZU97/GPC9fCd1rHsf2l4MQIDXvev4AR+YXdkIumVovkz
gaieF+1Ws9wpM0Q5nwcfMLcYNox359RVZ8NDcFR6PSFwEjjXjQMBWsbP2qdcnc1y3ZaE4s5mXpo8
lDUWVA8N/DG/RScG6TlRehP8Noo/R0+CHSYKSm8Av1bqrLYQBRZAD0pS40A/t4cisB1kXG3JcbGA
HiKqQfXiHvK4ufN/j+q8++gbfMWgMi4a1W5xw43p22jM6F9ip9C7PuZMECGY5+0t+NHZcoMtcB1k
wG+Uh+FvksUChsHJCxahxOVShFNz9GT/r3mEfOSX5mfXy+1rxZ7boAegCQWYJOC0geaNMUVkqSva
i9MWp9o4AvAEOBiAYQC/7a4xK7BRKkvBAONo+sIinnjawne9PPXBUoTlzFS8Zz01J+XIjFL03gXY
39bfmafXsbqmOSt+LpJqpyGaD8bUb5SG//t20ZEsIK8h9jTxgi960SHqwxbtKyPypRzcfEmq+Y7Q
7SSBqEnGnXJzfnHX1jDv3G/KFx4H9T1Jatlw3zlBerkYDnEKIaBmXP2qUlNmZYNXFwvckIzFupeu
iom/teS6FSjae1a0CKiP8IK+LqDMXq3BMktgFf3YyhzMzjtsSF3SnRTWwg+iAqlP68eF5s2go5U5
sX4kZJUXV3kLA9ZXCRgIwYSIVmXWQZMl2rN6Aost/DE7WPCd5v75nGBXMPzGRn/s78qBtIMcuLIm
TInrNvyU0XO69hGd3ljQS+qRg2acE6dj7nvCP8j7x3fW3/ruk0P2/guCmYTmlpjiywzs1hAMZQU4
iJGK+MzhmeNbrsGqgezfz9fy/SefF0kr8h18PoC+ViugjogogvNXfMBDvREhOZMtrHL2W03v3JMW
Nd+x8mYnD9Mh05YIAx/B34tLNM/f+vyld9JlWssk/xaUkkJ8fN1OtifNytUyvw2umSxNu6V11TIL
xc8icYd0LRSxw0b+7AvlSDU3WM+bu+LVi22vXW2+TzFgF+QcBe5zUbjT9TakMaUkhqLCmX8/sBvI
nP+ula4QLu7mybssRaTorc0tOU3SKKwnMqypucTHAIiHY63/3fg0SqHNL7pVoERaAHogBVOObADY
XrwY6k2NtTx5iUz3OSTznjIXppX4JO+Vuo01uQfiADlSmkMIBQxFR1L4hszJ/k/fN0rrx576Wbg0
BGoMqhZ2aVQfffOdOk/FgzgpBmjgdtBN6c/aM7E/Cl9ory0mwsM/vktbjeOX7QjdruUoiMIYgyPf
ciASHj0UsYlat28/i/T+dyWpZYr+LJL5b6kgOykqteiHL7JTS5aNwrgbSpuJgyhB2fOzYBWElrQ8
WIi6EZ8TD3kN+cQiR536UtMSygO1FK7SFSBoXttF2CSCQHcamZOd+iRu1JxJ4Dn81Nkem56HJgB2
E89LCidM2VZyaTtTCvEjqrwLFcWpXS76730U8CUyf7n+EqXeT8AxNNOPHVjrKacxJgO/sNvoY/HA
fIOjinM0sMfwfectt68SFwtBldKCHi9V8WWCZrw4Go4+t6w7VDBevYnHBJxl5mblNIeOtsr6R54B
cOYLbTqqxEsKvKWhAhOh4p1H24ACDlzBTqyQsf+QWGpf0jgal9sGIhnDH2avezixk9X6DjLKBcqR
wGZ1EbgGWcqsnz20r93KEyxgFDNKVhB7KAls2v8Cb4yfLRFgh/gFsFWVy5pPzr20vuSZshKi+rkX
/nGRjBhsKyjE1DD4yZNNWvL4MpMaCmee20BQPZ9EeWJ3xqu1MAZC6iIxPCH/yQSbBYeYukmU667C
z7P0xQG4XR9OsUJQlCgaiCwoc5d7fCRYMIDlX3tQDdYhULrdIYb18ElJYZXloXBdJfqVdDS3wRXM
QZCbUgFvgI9+i48hVM0hXGURCWyd6yjXyyikkOCaJN6xtyozGNgUGzYy3eB49/eXk3uagwErmNkY
2qYVGxHky85mxTHRt6149re16X9zUzyCIqjCPcct76usm6qhGvRh2AJ2AfVGRLsV2Sg3cZbfMTIR
mDya7ibVLptNRPWi3EYB2lsUvqHaj6PhwxcAaoNVBzz2l1tL1qGdGID86q6BWoZs/Q93GqqVByRi
ZfvLy1wi2CXu8t0xnwc0/7/S0xMqeA8ZCYIeQE+bUj4k0ScJw1Nt0UC+exDEIReMn88pozLP0LYp
paKz9XJinvmT/H9V1tH4q3dnRUWikrITXIBMZTiGMClDs/gxfpoHSI1jJxXYcsx3it9B1NwOr8oN
auCkX3Z0r3YrgdZsJvQxvenlHxEBp+927lRvMj2PcX+hRCZuD5wG2MuySD8mzJDmd1+vKebDYuju
qjkZYewvBsfvT2LU45YPUe9+tsZfQTTKC9VrqoRGpmQIKAzdHGvcFsoVF+QXa3c98m9n9ugmVYaf
ZJ1tbSlzAyH1A46TSi38CmB3khNRBkeLcDV9IxwA1+KH33TQW39XiEB8B8Iut/j/yCt5bbjyDMyF
mg8ILspvJenHNYrr1N08/ca5ANJjSmXh5ueAYvmGzP2lKmyWELhDdeQxWrpAaPPHe2T9Rndiocu0
wAd4iXzqs03koSnbvXHtx7uqA6tJMZj7YMHnYS3Fhuc+2/rQphJJZt884Nl0oqoquG5k7TeZ/AfQ
y2Jh6E9puEeHtyKcIGr/zZ0IE/xKxFODgPJ0kDCl8rg2tThIqX4vR2SXDpWLUsS/hkqpqq0G0NY3
IUWPi6g1g2g9QtGQUdfwrBlPqtIcnzx5rOj6kWzMZ7cowyBktjPUVWpOkSYWUiB8LcxKm4sxcnoi
Ee31Zv0cxc+2EdH9zbh/RnZurDL1p2mpnjJY0q4ktMnNNhm15Qe9HO8lkMMFQiiEVO41+Kr2YgRF
G4k7NwXuH1QJw6TkdLbeVa5Hd6T8fydyrZUtokRjdPjgz+R/5WSF66Dy07Xvk5hFGmsEVPF5Au05
i4K9xdTVXsDCOVdEcsR5PqNPcfbSGEFpm9NPk+v5qpZgNTsJkS2W1zsr5ZXKw+ZefCWm4w7UFCJ1
a/c8MawnI+BV3u02vuvlGATd+FV/4iaSso8KL9+RqKbuzXBC349l3EONfSCKLgMxrOxH/ZRnUhZX
OyRbdpcwDnzTn01QGZLxNWasMynkx2ZjOm7KQVG4NXo4ZBREUcsZWAelHgMPnyVn0x/AcrvAWCkK
3Y2J+D3Uaqvf/XFnZ5D6D5ziBG/HPWdAeb2TbRkayIN7cpEXvABcjOCHNAfdp30sHtJSlbsXxJ2N
6elx0mkq/OqJPNMoZPxkMrcWszre+XEJNa+8ZvhsZRgFH2Zhmg7Q4ciN4eTBtv+7d0jM3zltCv3g
OTHuonkysjB9WsQ/H7u+Ni5onL8UrYmjz+VjIcNd4y3DdT7rr9PKPkTUTtRJqtpLPHFdENXfUgtX
0xYKYW2rm/LG4/T7DKF2Y2Ql8k2UwI0VwuwACxWsYnckuDIyZUYenlVbXjHSuYzP67MfMeZdnaIY
KZQuX7OmTJ/FWCxSuMltafxd1FMhg4MSoxljYHijsUjG7E4BhpW/t7ltnHX2nxAMhxnyoi0R0+C2
Up7Inv/HLgiXwo4jvuOfhc4elQRERpLUTy87N3uxSSee/rXbUxngISCRpRH1VbR+oOWPVRFVxLzX
8t5sPgBMZwXWJk7vMX1MwNxwWXmjuUzk7WpMMqc0jK7oke7bq6p3vG+3FN8da8J+nd8+I2jk8ODA
kh9K4YOwMRrfw1astzLAiOcZbIfkmJMsaqso90/V8ylkk6CfK7qMX3bNlTfDNjAtVyUB2d6CEmO5
ObC0d2U0/NZrWiYkvewyx4iJuk4guwsbTIYhbZd/IV0Qvq0IPhmAn+cXbjlwAQnQPtqRAfYlgfGu
p6p7EBzPjbifImHv6i4bBT3xuzr9nqk0XmbWEu9SIcgnC5mBSEkj4yXA1ioUhBT2uwsrmKXssH7R
WI+QsRllQ6aXn2zV3aJDiNTpgpN8SitCKeMNM6PUHaizlX074nHKnjggyE0di1cvmmqBXk8SHQw3
bNrYN5ekPJeisdcBAokok/i94eE/ZsE0enjEeDOGLmUXhd1TdOazpyBPRy9AVON2uX9cUv4zRHPV
uefmDaPjjKJIv2ueTtQorS3taNt7JHt/rHP7ov+trHe21BrGj/Tz/46Wmuy5LrAzehB0trzCYVnN
1Kdh00dsXdiIJr3erd/BHibLPwhK+8+KzSDaAsa6rS8tOB2N8Y8OicgIA/HyR1mwe19yBZrFrG8P
Zp/B/AYoo9honuRwE446utck64kyAGLviXPB/UvQAgIiYzh3XM3twyEXsJXaq6d8oLb3pu4Sz1Qn
Sa1ClZ6FP1OnPG64FZTyifbD2+5yIXoZcSmejkcI7p+71ZDoQctki1z8k9yAEy17Ufzh14P91R8W
Q1TYsLXROqVpZKO6J3cbilzQCZzOm1QjixS+W9Dmtys9e19GHIYv/Q6aWuBw2sz8iyrRYMUKczZo
bqUTTBjUijbN2PEfiAaP3jRoMA8AWSlpaM0Ie+KMWrOMfnHvIRs7umhJlIBXljwjbe0DcshBhjLg
m/IXTyj1urUR2W8ZS2UqUa2vEgVF6xSHcnd2Vo6Cg8wxsmq/pn0UyEGZb3/8RudaKdFpWFTE7zS6
ALePCYUEgbqp35q+LhDaUpH/elpzsvKEenzc7TjHqXRZSpQDKiqwVBpqy2WiMyXcqjJQ7S0G+hov
YyKOw2qvCZQIbaQw7Mr6cURBtWyGYjiuw3wm4i/aJLSAVwI3kdw1kgqar+SwZuSHbbY2fNatWCS0
LdSMnQnytujGaluCpW+vEVLR4NiyWYMjf7aXfD5qijwkxYvMyZVTTXmn4WZvMRqrV4XKh+jIlo9n
nrk3mfWhTMC7vmT813vwtq1DgO+FAkx0ePTNcy1iPoBCCi3rNbUF2rzxRLOb6sa8P0UDuKe3SkM5
vosr5KLP6VIFNCLdMvwPYGWAl4yuuGCXu7UU35gA+LKEmetfenU32OpRrfcc+Ysrv3lijLCFuqUY
HKhAAsPi/uNoaHF5zi0LQWsIQCibYZesSDFl6lAL0ZLmviffh7BGfT9KI5S+4iUDagF4ZKCLNW0T
PdafKcUaC38Cocs7jYtNJwMioiZqKsIIL/5XhPmmRAXmcwlKXsqJ+wfaMd5Mj3t1SKdtiOTI7j5I
yX6pOdD4M5nu0n2Lnn0VjcOovIi1MXBtl6Bwdcqb1hTy2TP8T48s908BcxA+XtPZW/ItdPlDxzVt
Pukj8Zm3jxnlSy2DxUyRcsq50jd/4mVk4L9LbFrhIoljJ1r6gl1EM4IpVOuC6gazMCCeostT7qOm
A00dbqCOPKkSG60eQ5mXjqp34YrCyc3lAQaxI0NzxFdk/ZaEBEkG/zr1wKQIKXoRNUhKLuED2cVH
ale2/32cJLo0sXQe9pJkoFEKoAg5xwptyt+jw21TCPzkQj5CDfaiOWheyG/9EeZchG9dOEXLlq3L
zmVCv6pUHCWMvrDuSPOdk5+9Rxt1Aa1099FOb2AF28r5H0GpAzBpRLRy8dHsDKzbuUxSyI/kB9He
mFTOQDsnpNIOtt4gje2d+tjmRZnoAtxjCySddUIa0TnBnJ9FLPpcuOdTLsWxxK7MjQabT4D+pAHx
P9Cg4dhbleUduulN6njckrFmtND+h8cUJJwkzrXfJneq2MCppXrpXB1lzcR4sFEGXq7x/xpKbSWl
SrHUQU1dc76udJHWW1VnMmeCLGfAQLJ5vBaWDC2szVo1hqRndY3o+5Oe+fsCkParIsSSLijFDxBo
OorfmoGXQ4/VyWJ18KpGEvL7/8wNrUZfGVRxvOG3V4f4v9RgS6MpfKOkN0gY3TM+uKQp7yNTApRg
qaXHbML0Ya4RHY9LKahFpJCA4Zqa97iFFDCv0iVXHUwauMzXnW/Mk3l8cCCElgvUb/BFHFOqPbfm
5ik2ES1H87odf0NSrQmGRbXrpdQe1dG4oki4tbZHyF1QJIy0T4U3eI3CMwtecEKFFIogLaH5lwYf
oNivR3Q5q0sqVi74Ul+8UC7Q7K0qzDy677uEVGPJf9w6ete9XWinsJJqqEk8iPbxTnk43S79nnM9
fE1YHlHSF2I6Y/rcxE0bZyYgQT0VQp1CWxjU8gdSw3Pyde56cOf6qVaKzQlyqpkRQ+SshSH9RAcK
BSG6y2w5WmUBhFXr331j1qNyddHoGwPTwviBYfmPuA1FblH7+JuLK3CpduLdd57CGank9CQTdf2B
91E2obZTalduHK/cUc0s9wYkQL4/CSoKNvv9itQZohHwfYK7wEg0t8Al9pF1VKF+oy3kKCjjHeKN
Z2cTFYW1rmgTX2e9Y3HEih6NHYoeDMG961CiaUpEiULyeAJj2fB/TKXNsCML+I9xw4u4t84TvVVZ
04rYzGFIexDGMV3zVkLLcsaWLLaf3ikFWT8lXEozNiraaYv9wpDqIuPVcH1F9t/p5j+arH190LHU
p5UXJWwkpOlpTLr7wffqKw1XCy8lQiKvJ0hhxnV0q5rt0NAB/DUvt963AosWAXo+ub0aGnHYc4J9
qR0VjgJuBx07gvAjTHfPXI7eOc4kMmu2UFm8j+fj9sb9QCmmg4kyeOhiUYo7J3Ii2YFFeXCV3pz6
LmwEBkUGeRA8bmZK43MZeKQSP8GXcmAWvxZdaaZhEzGIt1Iq1riwu+FXCDnT1WcGstGnGbijmOhC
DSaqXHgDCH7NxN5w3AeMW4Kfmky4itJmjXMOgc0ldkbQJhPmbu27EmK4a3JB0Hnobp8Tp4x707s0
Ut3STmLBDTHbQrM2GmO/h9SaUpUdOHP1r3wLO0d7RZ09m7K05ezG6qWL312JU5Fb085WYFjCdGiz
pbqddFQUiK0ditecMJU0aaeoYNBgKPpXHHyvKdrTdO8NAMD1vBmLldqKQDKKDPihJRnTDZKshqTc
d9Syan7i2VXiclgTXuBllih4046/5AcOhjpvnjlcbCPzRFdxRtaNnlag+WVWeNxaTYluqCA3sqOz
6KPnTAIPVeHRqpMMueIktGzAXGe5olu3a6jQe8mlTwwfTBv8eemoeFhB78Taf0f9S2gXMoadskGE
WxRXEzi6SFnE9/IJo5qygEF639ARqWOVhOQLPVEHgKTkmuzkz4HVJziQGqxNp9SPAYM1pTb3DYTo
Yx4P1v1iGbjvxTTldNvVQIUgRdibbhmbT3qeds5cWvlKFkGo41Le86/hqhuET6F/8ld1t47kUHnh
obQCr4I3xaWygntbCQ4gt9W5ndXCP7IYs565EtAsU0PUf2AveXk0/ZmEB1VjS7koAwFns4X5Bnjr
P9mSFNNWMsVSSMnOkWIkImc1YuSLZeL1itPCccF73ANrCgoLa9WR1XqSDvmKWZHbfO5meDGj5u2F
KNGfmRpmFx4rfb9dmqoRo/m0NAkSmEDBHrBQdxLMQhed63ORcJY7XCwSBoGRAbugiqS5IE1zJShV
N5FJQOtnof6ihtIEUydekHRo5+ZAi03V8Zl7+WwnY3JlWjh18xdvxGsKNkDVt6Xabic1GMCpuYoP
sVpGnBgOn+uMgsnupAgJkrJLutex5fMuwOv6/fFcFNHU9llGmDAvOLiNiqiFLP6ke8XgZHzcTY6C
8O7v+Amg0JzKGTL8O2anbPzd8xPxh66qsxZcPYV3t1pIinJe4F5AJOlnLlO14GM0bKLV9C/Tsb+n
mSzyFwybubZAmAsQPksO54VH5k0NxGLuMS6tpwtP55lDzWvO68hKzYBoLikeFbJ6YUwfu259aUrT
QSQO9YEHjMKZj1e5HTDYKf1nJ5nMM43nwwYEyOZrUymIvzmPukx6tBNF002JvU9If7+V05jgb39a
GI/YP1ma05mAVbaNJ4ApjUxslmczFhwDjkqVpdyvO6gIrD135fZzdt/mfCG/9+/Of2zPvh5IyBli
4hpUbJVfvVlsvrFLTOkTD/oEMBy96qv7BLCGOWYNfpF/6mIb9oJEdWDy942NrLmW/k1YSx8D4ne1
x+epLD0tjIXSULKVuWKx9CrgJrkYTZx9Kec0PLrl6AStYit+7CaDMcZhITa8oL93y7twWW9Y4qqR
BYv4epRI6Xw+tYAcjSa3ZseIxP7exAtCSXFub2kytKZdH8vg+pMqkFxe0/OZzZQoh1LmZ/lot5JD
SthezU3kPSTIQA0noQbFbFcsPQJyBFqHydH3dHdYPiq1O4KZP3TVG9m8h3a6vsrlkFgkGD9dYvcj
5VpNBpSU/cHh04pbbCWUhZTVrU9LN0xVjX3VvIaJq/saPAyaYyDgqzYLXN0nS1Vm1z2/FJw60jxL
J/sXCq+LsIWbk80zjy0WhMQLwNvGtQ81QcTUpy/oNZb2GXogqU8FAQltKURbQuBIUqoVxYvjGlOk
3RBCOhbAvKqVuzUs+YfIdc6gUeyhaGY01SelJ25cUs18vg/ZZwudLChvv0Y0+ywvHeZjD0iojufn
KXeTUbSRJ24wSobmLaOneraChI5LmxBZCNduNL3Pl/3XL0rZH7AJsXXZT9e1ILg5YRhRrBFPrhjo
ZQ3QW170FpYJpQrvrBx5w4Yk7ouXp81lgLdEFFmHwk67psWLH+Ivv6IkgqR/ly2Xsz4eMa2wr8NZ
U/J6mfG5zbRTlT1B+QuGfyX8Re9cLuS8TJjXxjKnQNaqC1R1lvNAzpkCFe+CV9RuA6rPixB38uFg
6glrapzNPdpp4q1lyCPxJRybYMwEy1euPU32KYnxT05UNQLNrzMGUMsqtc4KS6BLlvrDk4JJbn3b
i+dPcyKm8AgOuJpw4Aqgycm6uPM0d0KMVGmMBY8/sIILd2aPChoOfI8Xq7Aj5ikvjmKbOMEjp6gw
795XEKGPuheDwUKcwvtW1PK0UFo/Tm3q8326lgEckvVxA0pJ2RMC7EoNhb4YOS73d56OqLRe87+0
ZSg3mgyd3NtQ4a5GAdODWVhQyZTTN8WnaRj6hdF3oA66oUVPn02f/CnmFM+pR3cB3eLKk04xUE+y
YLfw8jWnb93ZHOASzkH4EH8Y82oxZJCRX4r0T0HL2u8nj81uQZD8d4LBX69nygOyr/eG69IuqfQK
5Uw8y6Wf6BmHWxx8fbTrCQ2e+wVRsDIljcs9RxdmSD/XM5WbkpuIlaaAYfGbaUnT+iwO8y+tli3V
06I5bAiYekz0QEstyMkCQuZzAcV+Yyq9T5PsJyl3P9DNFPGC1fm7Uz8Jnqlt3y5Y396bR5jIQkU4
jLOqwTbPWZLfImp9S0EcBNFG2HnC9y7FrFXEGawU1r/9dWZ528SEOL1gEo1A1xXEd9buDkWktuDX
PG123wTOyZ+kuFOA2UcuuB9fJLXWS79P9WWzNwQMdUr7fvoaaOMVfC8fP+IWjzuPpC/g2fyq4/kf
hFNaWWqtYPD/QG1Vi0L75nlVZ5fh+TZ2MoNJKxn41EtiTkHNeJ7DvxOJa5a/XLBLTpBlb2SC+MPg
Em05IiweHmO/IZ+sikdgUuFYaCNjZeit0k2jPTgzwBT+UsPt9xTGoxGONnclYpr5JQA/yg3w0EGn
xwbKhtNGLmDeV75xIS+0PBEN6L5TbzvExyuZ6M20duVil5F6fQ0hZq0v4i7mpLoW+vmYjSiy/O4X
XmCtt+8bkqm6m1cnn7aP1QCtluHjvAOvqoMGqTG/JYc2QTToiQnsWiZlC+efQjEf6ZxjycZUeJA6
5cnH8Apg8q9qNoq9L2WMOSRE7tcBAERT+RLQt0P12Oj72bOw3R+N0sJlSUf+Lxdne7uHv1LIiU4u
z1Wl14I7+r4O2dN41G6CR42XI4+7wUWmldovu7Y/UY5P99Qlah+qvXv1qiCO4Qh9EXLFt/nDOWZz
ML8RCBW7BBXQMIKVj0gv75B+FI/p64B+U5Ek3FHmP8mwnjL8/Sp8l4BDJunM2H1iSLQxP77Z1z5W
VJS+S4HYROg2HrgduEHh+5dnWXPvzmpLxZe4h6ypLh/XRAbQYFriRFmFqb7pRRbgufEnLAqJmw+y
aaLGw4Qk+T4DoHQKsd9mYgfW0mEbHI/21+1bZJeWSYIyY/LKDBOxW+XspmncAjPlzJeVZYBwBbej
9TQkbRqDXAxVnJdyROYGDPBb6ZpyVYMFXY+/LrGNgGlbaTdH4asWOylx9AYx8P6zB1g+Ursop+Wx
TIHfEogqFedUU2FM5Rl/6Y3Tzl/CJHUYSzV6pTpAG/+H5So0Cvr0e2kUTIYVrtRZBJPprlQbWpNz
BgdYVKu7SeurPMf8Iow+CoMJZmgrUxst+MGcfry2VZYYf+YowX6bybot4daL1SPn4U5Fdqv3jBPX
MfB8v2QsbkmiIdyE5GZeD6DUcXtf4lEPAoAAyg1FVvXlfw8zFnm49Of259dlE47aypd7Ge5RSsol
WwzyXylGOogpFvCq1up8AK3HyCvguWTV42XF3WEjQb8LFw4yrRmhg5oSJWJ2cKhQtDiqFjlKXZCs
zqHABrusmOyJrcbfd2vrue9FmtqTMIIWS2OvB7WfEUaC0SVBuMIsOgiowZAy9R8FftJMAUEcAQd4
Np7CCaJeXToS2p5SKd7J2qL2Px0JvtuKRQrINonRtp+PiXn1fpD0h8M1x7c0Ml3lAR43gnhHAB7S
rCMKWkG5mZg8cgWbZB6yDUy8iRgXlSrVchkzkIM2agwKUNW5N1huGaeWoN/WZtVHTRruS92sf8rq
CNMui+PSmL7jdnrYKmMo3+K+CQW0i5LkWQa5zH8hDQ7ZkjOcEIwkWZZZoXy50Nauf2d8bfh7huCu
9ZyI9HlVSdVm5KAd/S74Ec10aybG+JVLvJNgWTqTjvXDdcipFX7/gzMPd97RZ+Z+/nra8ySpt7J7
rSz2W/aTcphiwWouP1Y7oASobC5maqnhjXNG9ij4nHpAX3WAaSIxpe+hzhbC/GNdTiAluKD4wcEj
Z16WIBkFTUKpvtQFOSeQ20yJ8nGrHGbiBlTu52CYqmcJy++98zE5wBOAhpUWK9fSLWtklFtaVAOE
Cj2Q8JE/TZwuc+JPNGrkw9C2dIiRJagO0Soo6e+Fqw/qKbJzs4nMW1YriTmGDuBPBWTF4Ji8dKcA
hCRes/jW7Vf5kcUEruzZ9QIUaYUT7JdAz2s8OnAmBFJl5vpGF+UiZyw0/Fm++fPeOvkIdschx5at
Jq5gxfxhiwAGkwBie6Yh6OT9d6KLWWfF9uqAK786BQNE1M+z54z6qJMzVAM6rtwKqiXkiLveVW1B
njLbcQJUbQMYgfvCM22Lp6fKU2clKg3sGcx4p1abY/IPakPJsDNXLrGwfCCUczsUtOBfsdxTcO6K
u50mE9VTR8+/Jbq3xPP4Eg7kCdrqGfbmHt1ojp8rMdSefOeX5E2JtkIep1Y6newV2tCWl5kZL5CA
Ev5MSSqP7fmeRXLd2vN2/qPYeRtZ+SXZWdRJSt5rzZKLzxEuDiqLuoHcLLPSMhi93OwoykjZgGZl
BO18WqyKdbfDlEofwwyOGfm7/1CesFOGc5xPxvT5T3wIfLjMb8m5E451606dfalWln4B66iR3l2M
N+UoylLJyCEJ6ygB2eGfvK7SvFMiCRx9EJuDWb6ryWqpjtm5gXyKF6AvhMgrHXXFs/mP9+kDZ7hD
fZnJkEMy3cLjBfKhJuth/bwhgZj4vR7PSBgdOWRHvEhUf0if4QGVv8jKKpLiNmoWZKZigiFJlQLC
J7D93WYsAdIMhZddns99zsHuijiOQzbR2Zos6WbfQ32Ng84/LRf0qVJhnoQMKv2UYKU3Q9pNsZG6
dVTm6c9rBmDwkGWNjeeilFPJebFddTvaL+CZ/wt6WIuYPN855RoT8eqzFMcqedj2uTzxEfNrSoVw
XuRugaCsgZ0Gl4dZFiIEznfo5Bf7WbXmLe7gEHVzirqSMwEKiYzHXKSqaN7IdvPLigo1qJjiuDK6
2m6+UPdbTgCGoFC6aVp6IaUth1CXYzz0umvq6QjpRwYthIoRFYVJr83oQC0memu1f/16mI3aF5q5
CPNOeNfeCRGOOC4FyZ0EnCF94iffdeK2VnxUDro33VECyyH2YUKamNjTQIskVbu/27qNT25OGJD4
T/WPNB1NUFI42AIisWB8twT4CenkPuL32tCMoKjYSyeI5ofoDI9cvFfo2stU2F+eX+Q9c35ZbusP
TktXG7iQm6juyI2DyjTxS5H1FIFkK2J7GvnPn34VVwzKe1Av/aLkVfaDfH4FD0zBvyt4bR+s1L0m
+tZjr6TxXkjkRvlQthGtUxv22Axu4MvTAA0Dimqhk66aqtCV0Y8Jcq06nxzvweLN4e1zaS68fo/Z
f+RUP0tIK7W3rc6BPLoX2RA0/7DSUWMfAWus7xchoDfgTnY41LTvbdWROZFD4WatuxR2fFdanAOv
3N/kvCicrD19uoJBHXa6ZKrHarcMjsjbqbCdYWIFpIUhIQE6cgvy3vXbixfciF6kIRUQDa/MMNGQ
pHutW7tYsaFU6x+n3iAHO6bvddJ75nhj4JEwUgPJU0tfvdffnzkHcLJF8wum20gO2c/hHCXM/jlM
i/H+ZFaJUD42hakDC3mSaG2k7K4zMpOCy5p7PYQhYO8eVH4hzXssnL0uXExpquQFI5a7GaC+WZD0
QeP7vQSHOonhu5w6staGZe5+/EHpOZtdSt5nEfAztzRefFA3nzuLHiWcEIxI5OheCmAeCheGIn/b
WvnquTl6WkotlsxnNia6mls8vWDdFjoiBltSEXmX+RhSteePoc51hivvdB+/d9Ex907WcLOQtf5b
KKoWk4vgiqEQfGRKChSWIHEjC/PKqUp18O+YWdnh/p/kWOjwM5OI53iirJ36zQZQFKERKFj48QoC
8ckeQP1Qlir0k/Z+5snlg48DCEwvaSRdV2XRTjDc8BRZtSXrdMAcgvLGa1ckB6cbIFBc0Ooups19
GHfrNjYIHchw4YaFqNEAcXytd2Mzp239jrBNoHTb/+xtuJhqhUg6kb3qONcypeeMy0quZ7sro7u9
86UeEDhWo4HBqRG3262aY4+wAzr3Y6woRRG74w4U/cCWQYu32QG9vmaOs9puwBxA0n4lGGP0EAd1
H3g7fShsvjFRGHgzYvymGtyBxiOVV40BqI7YfL6FDtM1OcBFH0HPLkN+3g9PpI6mycP/WZ6H/gYZ
XwkHoRO5yExbp/nSFubwyhiDucrU4eoyb0Pnd6MnRhc6Ace34ZmSby0g0gxTgMbOnKhbmD4BDQoF
ygkHgkXtT36RBlDbpPm9FwT7W/HbD6XWfBfAdgEYYZEDTro2m2OOS87qZtcfH8lLpsW1H1MmryP/
ot2YjLpDh7xiZUyaJF5+SnrEImMByCtomPo+AGIMYB6A/ZpStepGtTRNV8IG6NLaOiQKjEJUy4uy
dYJN0Cg18e7ZrYPaH7y5XtwkAv/5fH/tNOxFK2fBiSxW5jrUPWuyesf7XAuxzthboBsm+xVL3wBM
XBWxRf3p4UMMOaObZTl+ZSiU+8IyVTOC4QpdzE3DjmbRYq2Hr00UNh7pbCxQBEkDS4TbXnIP89jq
5QIyF7yrn9Zyt2wR8ATw8OsrwA/YuBEO03Q9wuiYin3SldRaRFwo2Ti/dFuErjCbVue2cHAmegWn
cnxepxQdmoB0xSEZNfT9PfvL6hhXDt/V5gCt/OFN8QPXJl04WpMmlyHNVQQhy89wnNuJthv+XGvh
lhU761textgxaeja8zLErprMPyauCOQ0RWBPRdQ99rgHGPIDPdjpgZEiwncp1PCyjBTv3f6vMUNz
J8QNLW/g28yb5tiHLE3+/BXtbBQlgziQ0z/46mRG4s+sVCh6H6J9ZIN2njbvHMsdpCgA2GeKUp6S
4ydFTr8drhOj/kSYZCUZJlE7rkwxTXHTZTBwNWp7pIpV+us5DrbAQ0irOPVOdvqg7q26nZ3/T/bm
OPqdz9oCqQ8h/IKbKlxpc5+tAKbHQbVbv+YXCWPQSQ2EdXCxzHSp3bqT7HL2742kRXsYtAyKRruU
lRtJLDUoUL/UOxbxFcqkv+4YFF3ZrHZD+5N0AY+KLbwUoWNifJ2wpKGnMxKcYbuM2lwe21DvaAM9
m7UIkmkwv1i6qgHHhgPEpckfeGl2Y6OI7l29JIO62/vPXRFFtDhlAmu+jsy1+5U8n5s48pGvZkzT
nnBS1MI3irmmEwGWhYJxfOB+/FyTEbFYWBr77i4FPAaTKiLHjlEjPXhhSw9IjvDPzIwinm7JlCAM
cEp3BfcqGCs2dRKBWjU7yv1aldC0/7zLcGPu8Y46pHpMdI7BP0/1xdPbrPS9+GUxh2kLBdeeVlHn
N4IQ6AQxzAMQ/qsf1UbTeqqz4EJiJHxlyWjNMN+VfGRATWfr1bM+L++vyVotv7Z5xgJRMeaFmZSB
KVsN/SeaiSlbU+RUxTuJZvF6ETAe6m4vOJV82+vW1mpaXxa0TzqLj1NRa5gK5sFwut7F9pmJwFkn
UfBOsjAtmFB3stxPN8glB3PRf34m28e7YWWS8RDvwwuxXKOAJcPisLSAymY0sMIu2ltDKIWGv2AP
eQdrluDtd33VJIT51CM9wG6JrcDa9YMkIGyOFr12VhSP9FUZmgrp5iZn9E4xDrC/2exjHo5Px/WD
eHjU97QmgFsnH/9bR6z4MWYtxk3e48f1u1ZVIN1iP9p/RcELHUoLhqgM3y6hBBk7sHy2ff892iME
RdgHl2cn1U2JCx+5Ewi8FvQAlOGe4ngWfiWUvCnBRxLtyaqh4iMaVt8EFfFyB30QJYbk4xJN7Cdo
gDRERmEzbS4EdgUYaI7+t+cpEttt+tvbyx+vVUqJarZ1Kcbu0vnjZ1+ypsAxLZI3yHpXcj/QPyGO
QWc9Lrd4NTg8iBVl8m7WR6cRJDLExcVle5IGMDs5oL5XsZnZrF7OTZtwEEoPO9SYc2x/xSdBjk0a
Wy5yEe3vzxmm6oeh7JDv1eqEeIIQplRE6tpTdg5BHmEKKGKJ4yBmVjvzjuwgQ2VsiTdV5cSbRaJa
LWAlu4eqcDWW4iPfMS7hl7AGkD073KOr0BBUP2VC6C1hxjA/1h3xKM3jz7ADm+tpWI/xDkzBohY9
0e6zK2PX75Cti2ASHJbopH4l7eLvuuTtfYl5KuiBKRSK1RipGFxhKkPFhNaYlxhGdVHgZ06Yw8M5
7Hf4OqTi3yNZQZNZDPciwnHxGxFxeevT6logz6pANQiaI1uZUP/f3zXbDCc9fXML9uAMDsM/L2/v
rf/MEPqUCf4/+FxV07Pry3eDOeXGSCQGTxVxzX8CX9/3xWma21rTj7zGN5PBRRt4+zmWugTuZkKe
cx5bd0z6oYWz2N5WcMnXnz2tY2AdQZ0Pg9rWxcA4479ld8doe/93FPV1ykig6C0ilWMerYA5AXde
t5qxlJdWxLUDsMblgyR1/a6FsdLBMbelSh+nzht/3EzEFLkmhq691d9/tZdeID3K0QRHzfcQZLt6
uG1lckz6RpM8OwQf6GxZYHTTGB4SLuauAZZdAyAiyxAwpeoQmFHaSw93e2X4h4LYpVVUVWDMKd2F
CKMni03j2Aw9aM+lmuPRPH8WRyG73a0IneaJN2x+vkQgCJj5A4ct3OuH8xdDZD9EVHMQ0Ff6dlVi
SILwafv56PYQs9yTnLoEvGVgUP8460ILDJgptucu99SiXDSgctE8j/SfTxgJoS0Gyl//SBmBWOfP
h+5uRMscQgXKQBMyHYg0F9e+SOKaqWN9Do6m+edzuaUR0+PhuMKNT+mmIpzf0C7QuI1h37A9cr+E
2F1BpfgH7g+TahXzOiO2SqTibWRoFCyt/NmxrhZ3dFXBUqAwE5kxZYhKDRUcCUroPOYdp0iAlzJU
uq5s4+tdaxGhjJCb7N4Wp7Ol3Fqy2KFRIZ3zHLAf4ASJcfOexQYof508hmsY7Lo7zDb6z9M+5oln
rIieM7oPtjTbD192u0QxT9N7jSkviFbIJ6L+vl2CSOIEqzWnwMrqeK1T/0Yolb1qvOukAYwZ63/D
B3NfuwdmI2iPYq4SvPcVye4tHYBozHZdxN40Y9/17oWbsBje1rpqm+ABmng0xNaxI//Pe//yDxmp
ZWjyEAH+y1Yd1pICed2cwar4YLMqgBTicBb2HbqngOcUnFEVJ2nYYxu6f3QGNQtTiEjN+nH32HUt
2rfur5t9Vk/kK791dySOxijd0QprCtab+f6J80OCyrxGKWVRe6IVnZdXamVfw9Huj5btV0XCWGcb
WZH703TPn4eTD0S0gLd3moltezmLMsZJEgLkFKN8bZ18oRKwCoYwA19WrLZaPkYq/Yz3UdgaDBZj
2McXUmVHrjm8PgQFCv1J4Hkch5iKF/u+Qis6ebrH9tO0TwvUFf4X32zhvCltSqb2ruSZ1qeGd+1n
9Igf8WZ/T6zTi0xGHgAJkIQisfzMNZD9RLbYGp/gsX86/amEb8pEKzXnpjNl6xQUABz9ULsTnJBZ
OniHpf50pml/ieaH7F+WcRkPTKMsXDOhdrkhGPnPWfoVP/VmQpvC+U9yY6ZSdqPD+qa4SrM8NaKe
KFtLXF8Wypi/fGc5x1RTnn95jTluvDe9tp7DKL59MZ9cGU2iTUssadwH7sp8+EdjA7ZS7F0UZgQO
JvB3U36Hp/3SxuQbuCB+gTx7tABLCs+vLcncZWEA0bYKvXhitsTnFGLuCoXUdZ+uTMksnT2MI/I4
lbFWnWWDSBhQ/1OuI6HLkVBm8Vc7QWNK+FoFKOBXU4HPRXkdrRWrMaqZIPk4SB7nxzavYePpNfcb
f56UYG4AIunTRz7NnmSpX7XBJM8w6NYvJG50VnEejCWGvnJ1prGTFM0GFVmtodGgKZHZYftlgGne
AJklgo6wTzfiJWrRpg+3pqWGwyXYYbQ70N224DjjVSWOhjT/jWgjzfhdZZYFlaCa5us9o788aypF
AT+LqGlUAw+gSh4Y+nW81Iq9a689r3qhxCFduIr8pSIEInpZhghdh1obUYwkR823pdPdNpzajMCO
fMRGPeQWemrFKEnAY0xWR6tEMhjzrb70YYUTV5WOCLTozppn6zoZLZx7P638B8diplN+yWu94jAQ
gRx3wgg0MD6QPtsCqc8ZrnW8nmZSqEhXPzQfmEB1TnQDJ/CNFq+zn4ld6jocWdcR8E8nYI541FBn
T6Emi6bKeXFM733M3BH8VXbokm0wVM2HXynlZBQ5NoHFF8azKitvXAXhfTyCnRaWGX/nbLt+NxRc
p9mOhylM/beWA3S57ygmMCc+Ww+Fe5P+YLh+rVp7EwXrN5Ix9asOMB+un2eDCHlBwiHhCiRz5tGz
gVTh+zLrx+Hg2xNzzTu2HofbS7jPVLOKRJxBYJ2PsZKDh7vkKho83teXFN0yk1645QolMDYF5LPY
2RnHxHM2LNv/02XkuhieyNC77HvWka81JRcguNdHPyZyG/jDkBZygKnS0y/P3edGxMSWn195ARGq
lLM237dpv220zGvZZH1ekN0SZttIca0SxYPjaWSC1dHLteNgrR2M+tH+nKbsOBFMzJdkucGcESi4
DNycHATqffH9xe2z6Pr++Aiu4Nt56jubtE8ga9d+mYQWLnSCONvOi3a3zrnVyWu58jTPE7noSqIQ
pHhJgmF+s0ZpGTvlJbF1Al6YtvgXPuR1LTQpHuK69cJK0A3FRlGfeMXF0M3VteGA/FrCgShREIUm
LI3+xWk5v6bqzsfoXR8hCTR5JU44D1w2mVz7OdGawciBhusBrnF4SkM00X3LgfewSP7eraxHelKv
WgJ/kWMog9CLgPdF37Smb0Ba9ux4oQ0WlOiRipXzdXIiprUgnheM1CFhU/idLahvroV9gqS5fLZw
9d4tTjT2ygptDjJ/EUcctJu04JLW/74YSGsohd9eChd80WJeTr5Y//siLRxYoBG8S8e8NRuZ+6qQ
LYi2B25+omSACmRqPLs+TVtG8ts0Rxh/DHh+qdaBHW1AJPCyykJ2ba9Crd7cSMkG2HiI4NkrJwUl
hltIrwn4ngjfKOGc2Cw1Uumt4T2SZA47tb2YBRaeCRTWpFx1iWSNg9HfiuFn1jYPwG3ghxvFLwrC
lh8OOEHVM+Qd67HaXxC58wy9HQa6p69Xl/woY0A2chDdnraMjqn586KWJ01Hpx7DQ20eDaBRBIZU
hbF42vmlS3/wvZXEd5IKMo5RXDgdRk9H6SFxJG7BcvTFjmFI0Yilig2rXn6NjHeizWTFe824P3Md
7NchFnVA0ziJYFbRJJV18aCz1nPPUDqbb2OjAs7NeuBYNoRjJsCRO4MGTgsDFq3VBNPjAKaf4i0J
0S/TUD3qejbaOCpT8jNpDbxJX27TaxkQni3lAFe/Pib6tQ4NCMHF1oWOoQ4hZib5leilbeQb1rnB
MxgqebqzIsTH5L6UB6ksEq5UpBe50EXQVLIaYLeVjE4DlXcOKgItzYm6jG9oP+J7mVkxSuSOgzyt
OAez/JKsC9l1P/+MnUENVod7NraU8zcHM05nyqgfH+5+Vly6Ej+dEhD6QfDza4xx4L8dw4C1rD/S
Tw6g0i40QlVdAdigaolhKwJddvEmsZ5ttqBWOVi21DdMlMK7AuuDwf9v0Y1WZSvTEdDFZWzt9Xxt
tqtz7OsxTQ7wHhOSzAeljw/gQzUj1OLK1xVC/qdhZEweF9D8CkajBsfApL4sup/QIF/I2JFwk5EA
mNK3gLWvXlaRFgOxwHGq4suz5F20+zEMotJgiCd7ffbYIEndgrLD0g5Ijvn6V9MGHir9RQxUxNiq
yrypZCBsLhvMg5qlEdDTWqnYNCW9lXDHv+dji7DkleKyVZMXCkfeKoy8bIEBMpkZXpUaALJexjZA
P3M9NIDArTAlBj0OfanIMVKz6VQ4IPsO2uo9BIuYUAXh0OeOaGRa8oawScEb5NTiKCtwhb2+CjF/
bcaYiieBGMa/v7AJgEvVADj+uFu1dIz1vOBchG8IGm8F9/AAbboZFL62jgq7pPuNV+tbv4xBY8gq
kVoj+Yvj5O013qxqzhLJOxjhD1ck9xD7MUazVQI0dhl7GpX4pyMovvne+ZkFeVzUv2wnludGAOUn
wErRB86+VslIyyvBUIv9/Uf/P1eSJxhiCpiHjp0NpOdAirxuQMbKusBNnlC48ic1F1ZlpmoS+EWO
+xybjkqpzL2uEj9mr5QoxaFTleF98mGLJM4t9zmaMa0im4VYr942Kd6VYmhRVKoQjfWun9BoUsKl
3CIXMVgPyh+FPTeH257QAMOHAjaEmeb9GtwsQqvyccGtUn4bfZ+h4lVMTY8fzJrMmiAOfxCP8a6e
iI16lPq6ogMUZuc7cTkyumnzSddu2QW2zFDSveLZzraUmJkylw90+2PPPk//9H+q8INAyE/lHA7r
T4eGj8sgqK6MTEP5ShQxxxZNdt07t1c5En78V8Qp+T105Xn+K3S/JaWTO0FlCR/J6mAf0aMdWKxh
iEYXpRUYl1rAxtCMeo4QJ/lKjhXK6uMk7HajzCa/Q5RGeyjDLSKDXlKQs0WT3sV3UkVFiz27FX+1
Td3rlsV3oc7ix51KE6G+uqx612Gil4YT9cC2IlJfMQr7vLdE/OuZW1xMBzZWrZpi8XrSLE+fVfee
37XG2jWWkaRJjB1ClnB+mqCBzCdq5Yew4JEWBYPEYJOcM3m/gIdpxOWZdkOP3PXVBUqjaOulKlkz
9QiRIyqtEY0/0Cxt8CreQTwhS30j5i4ir/lO5StqmyzwveKbX+GPDz1RCPZfSDvFvEKPgv8IjDy4
qMvVCtGwyAIn2kV/4nKeIzar+1vzONG/iQ+JbSnaP12bnaQKpxedYSGddVCsy6/H+4vV+7ddDqaP
ZBLOnPSoZDm0KNGiy9YDCy903GeSwVuvhCY9KZUyJeiMZ/9XIv2j7SUUArBAJDfQEDlHkvxc8MMs
ugQFY/rCnCoHLEtjvMXKab3YTmZ8cClR13otmZd8/j+NfP9h1hJIssIsv7kU/Ia5DVX+3BPuSpv3
5J9f82+SZd8zDs7+Q00jTY0+2vrkHrfvPjUvbvAXX4pDTXwjGpVT3/1DGy/BywKz2fX9Lp7W7Lem
3DlOvIADC1zqlGDbGbjOmTeTC5O3P3MRHYlytZnKz1+hGYoyvdiVhv2j7mOdcJHRq+nT/yOzzp62
R07G2VpO6NUJbSc6hXGUaytqUCNvNCtcTZfM6SqubUjYbO2C4O1cwmAQsulzNIKxzhGzn57Rusx7
xjbokdtmIJBXOEyrfm+NSUYfyoqDQSZRGitWkOXxwsacmZWu7Be5zOHOReopUR3u2JTRT59zTIMM
1CvswVKMI/VIFlMOkciQd4QIOzDYwgi2X//FTUTGrY6sztPknEQCQw6QGK+R2iZ/wNe38T8i8CD/
ZWo4Hvybv8Kc40otJYLAkugEAejJY0LV/RoxSm/FCr8yQf6saqNPS69E1c6lTy6ItyZctjEKf4jZ
TAZmIeRQeM/DpOSzJpLeC5hYaBSCA3ZCE2zbV7OT1z9To3rdBq+GyM9o7Ga4XqrBV6/bDjKgsBaL
Lao6B854OqjFnLtm9H5fmvO5d457vzlrfPKZ7OnrM6UBzec4vpV28kq4cvBo4vy0QTGKy1n89fx7
TicuOQpp3TLrPo4XdsA2V7huYSBkKS8OduMZ0z+xzLY7QVI857+lZXRUy+ssuaCraMr48Jo43CdV
ZeskHNFuzQvJIJ1sW4LrzJqKH1VTpk+HlKsLDieE6GJyTGD0GwZ+wel05xwCOJ9Eyewfo8QHuROs
6xlwN7n4xXp+mmXIOf5Gmw6El4cxYj2eCCznfTwqC82IdnSB9aLWXgRMeCF3eq8L9qIPnyunjjuY
J5bKXu1t5EF/ktCciRSOCSpYnDhu/uIrUqjs6iFNh4jeevLtwubEWvCN2//23fH3fEY70xy91BTU
uRwA0wa2TGYmY+PHiqrwb96SrmZJsdcSv7hYgRdMInmTW9BSn43nzCJagoVw2ChTQHtroPbzCjXZ
GhdLtGFssF+CICkc8SKKY7kTAVhvFzeiGn/HmTfo2bT5CN4aV4Bfmzwveqk26Uuxn6gHPHkIin5H
uiFBpzFhClDkGDNP4m/2Phj0WGQAqUhUFYvw1k4oaKtWb+ox0pBarRvZ+WgGPkvoMqAcawrmwc+E
RbC8FNYRABXzCZZihPcemvIQtrm4O6kRlsr9Lc+9zjr4x6ZRe8VIeE6i6givTGTK9zQVsHd5+r9Q
NZr5WJiL0+eWlJcMafcZ/Au2zD1gRCIzjZbEftB9pvtq5CIUkvc/hEuuGakyhSELL1h5HglEdEdT
gMVZOYHxdmOgfSQfiMzeieJduKnFxFYMdAeDO2hp/fcbZG9J7E6v/Sj2en3ROJ6MZeKtyK9G3U+f
IXGEyXqtTqvXRKkBjnsSRRlqxeQQOctSuE7AnLfTLvIxLs1tnwSl4qERdTibJLutZk5rI7G8Xfb2
KngQQ+n+dIC6KtqMDIZWMgmYFjjlzeEtd9iAWO3YaHaWuHjPcVbIqRS9JBQ5uk8yczjNWnhVvn/4
aSitGw75JaAMFW+v/8vnKO63W3iwJUn+5rQDSE6JyLXfjZ6Cc2lxMQSZOcTCYZaqOJ8XAbqlSl75
FeWbl55eEJ1HYmudb9ZnVxcuN7EiURLHB23jUYtm7DEsojZTh3nh9ZUP7IriM6EuL5bLSCxytLcg
eH0hXtdpvecdtnMr58Gz7gQxePJBAvSsTIspfZUjhOy6UmwawAHEqzD6skCVnPVp0sqgBcfKb6Bo
Q9yhDKZWD9yv6qZsBEYc/S0vqtiQ+C1vILr+R0OLo1hrvP6Grc9yAjiA2t3Tjoun7vMk+9ZuzslO
ZeLgjFjxdcEi7LNBtlC9PnwxVcDoBxk7+DCsW9f0zIvPrWgzzOI2wxbNFGtQVmXyPXhxZDCqZN0y
A2fKeIvASvImTsA2Tnc1hurab5XtZ+yAcstRLE8slEr+xbGAS54jzH5Ts4CTPddV7fKKU/2sU4K5
UEQUQx6VIrfNwxNd0mqoQVOS/Nosq4+PgDdeRUPRjp9WbG00W94wA2k7Mtdztcp2A6B6isBBO1lA
ISCnT4xh2PkXD1f93n84gFnMb/0HKsE42YOksM9ptiT54Wm7m4mah4K+s5QzE34gups9A069kDQ7
gatviNYS/ZVno07wO4xXXLb2VHO2mYzs0l+8bnCC9rZ8Ap75kqjlMlo5hiDzv8PxHjn8Rl6l0eax
Df/GmGjfSTjMWCVmDU70xgFznDYjebRdKoKKoDzyIw/895OCnYIa7eaUhFH1Fw+ZeCslvxjAsfHM
CMa54bVxfQBDS48NNMCGifoYaIfl4dTjnQSij5J1psk9pD3hHDKEEibe/M5XxSJxNuXulARIAIwD
wF4EiKuhuD0pQEz1IZPsJ61kG54FFoZ9kBABxRrk8mu5t/9t7tNQ8M1Ggh9oKmUOcRAiKvUS9wsc
sOXM8Zhljx22TVFlpXlghIxTeuIcpEmGo2ywMN6g10M9pGfwFoJFKLbUUhW/J9eiDUF+hAsF6RaF
JOe4YU4dnNBkJ6t3GvqK+84r74RYpTRCBX24p1C2ZAqEzeqn0SJ1SxahzXQUlrVNciIQ263DINcQ
J1K0YrBdqPfZ8OYpj/R764BwworHuwDBZmIymm5N+XrmVSGoVwSo/1bEvlLa5HcNZ4BLaAw5ZK9I
ulZ0nFcHPL4J80b6imp7D/mNp3Zt7N2gjKDdFHi0/QCeH1ijPIjrVFrMp42b+klnxzKuQ6jU+DpA
wiVwx6GoVDdohxUjtz2fKknJqa3qS4TW3Z079ibJNyzXgLa9uF/9qkPwc2vTogXbnvomc3R2SqqQ
1Ol5QKpDXdrsqRXNs2czO3jHUMic+f7ff9YPk2CUx7mnYPgsXGpZYd/U4SE4f60SW9gXunGXPpRj
wZM6y3aUVXxz+XH1OD8lCYhzIHX+Ej5tj5VRO9xSZ9JrSw6c466NreyvSrRKtMp4R1pgupPSm5Xg
KopzOgw4CMeSFUgLuwI0nLsAzCAqIdMkk93ZXI4bhFxDGgNdVaYmoef3jEYKgIjpNURXKd8NllGI
jKPmUYIQuz6UjWL2BPy29Tq94aX8sDUXBXL1yMpIJnvNZk5v9l1fm7FKBNA4rSje1+W/ipR3PNG0
py+qdkCW+7yZrsTKz6BpDo94EZLeItDqZGV5UlwPBL/+RbtUb3/lfmKw40iaKkZa26Bhfk2U9ySc
nTq2lYiIKzcaiGZHu2pWUHcrdnE9RnY1FfNIVA7H2AJwicMj6N2sQNsFQbiwLKOILJUKz6Vv92Nl
1Qx+L8cF0VWfGjeL/YSK1IjI8OWNWR4Zsin6OtasvCmaT7KttfczzfBSMt5I3khZBRqT8KTKR9II
mFqptwBPhPE7lmaEjw0LTWKhQrFiK+6vp2pqvz8sSFohyOGjGStsHqTL9IyZmkhWWL5ULZN2/LD9
b/VPxoBBmwIartwRMV39Ox0lh0CqVZBJ/MS0GatwjKZzkS1et+YHY3BXgmwXOwSX/4eQVXyfGG3Q
EzLL3b7F8U+SyUKajubNoa532Usc4Cuf4r6UIvvc/5ZN26G5mUnF1XbnXeq+22/PPZcH5WX9OLp7
9rVRc64spKOznDk5UO6fenJNh+Y+M7nLF15wkltrVY/GgRJksA8Ufa03L9Lab9t3qJ9Y+qKIzxmp
pJy3Mr4P0HPxP+Pjqk+HA/xGT14ZY3VYeuEeO4/zkmYLu+PvFBxUdNsLvQxcHTmi+FV1ehaxjOLr
Q1MwOgEF8qq5TjySNhZgO9foCTcfUBkNLs57agc97k2+VVjWTc2UHfqAe7eZNiPbSyZcdehRtu5b
cVND20BAZapGhRzIIlSd4LCrWs6lhOc74zWqcnRhxCwKG+DsaXrziQbB/sBk0cFuhiimT2R7dL/Z
uo0uIjzYix85nTOPw5+YTnBWdB4Xdzr+bNnkQNYH3P2MDUiS8ZC5p0LRt9SZFUML0cVF5bWgGxr8
rcBGU25r2dnQNjIJ+rSGin0ydq/dohjA26ZN3v5NCTx3xlaKEVbBy+zGsl+7HrgPZy9tSQII/V5y
6T0LR64Q76y1XPISX8VqStRNOanVn0JJxsVAWBD5i6lzx2+JrNrdwx83tz83hWvgIdElzqSSinvg
2girF98J6djf79PRWaDbLKEnLVShsH4rbm+EfHwY+QnvMbKCGWYCNlyGOHoDY6X18NpogNI9yo6p
CBaStXQq0BK+bfRpAjUItzH1OECxCBOvBy6tb6v6pMrBBw9O9qx5Vd+jCroB/h+UUsqyp+sXxe+y
GPvmEB0sy3pE1bRWrOIJ4x4+Ic8Q400zy9YKq+aW4Ao2gsklfkCo8NehD6KK6hfdUJu0UxBpLDFL
0yCP/PJFcLlvcz7EFvor2kMWd7CB4LyamO/laUD7ZHxFqXN3Db+KPdcGPM/JGq7XlgCc+7nJwrX4
cilUiJ88GbLkwP7Q7AUgz2MJjVSjp7eBZFDmOQi0igd/Tw+/vVi3ZsFzJbAC+I68UlqpZ2piujgO
ANJ/skCSeJBJfz0fVyJ2/gWlirsORde7N5zXzd9yN2f5IrDum0F/8ncUoUwCi0ciqmneqIYNNlxt
Bb3rpO6k/NjGLfYpKl8wsvN9XjQn4w91esLCV0hzNLEsyir1/HRxzPkWMrD3XCamJ8rsfC2guaUf
4Lp08umCgBgtZrBLK2CmlwaBQEu50ZSPPTaO9VfuAoZjemerU5VgMPdcNrT6Nv0Dd+cVLzvwsnTI
GVL16JeGWurBdOACWFkRBWUiwDjYsMKrQcKKqVM0z/k5JIuM2HiuceekLhc/CEnzccbSqt6DOTT+
HCdKm6XxmnIguGDPozp5/V7cFHzeA39RI1IsAUs7q/cm8a6qp1F701zgydSrGkxLEFDl3cUni/Ay
RdmN0CRjoyWQ7Pqbbn8g6mHBMlnL6OhpJAjA2b2N6NFxORYj2NH8omjNUb1LEiR2DrZNUIMsi64/
WJq/LihlFYfUhU7kI/BtsKd/5BEQVE0ChzlfA97iij/nKMFAdwedzWu0VMxnOhHue5xC0uHHK1pm
PZIK6cUeuTYjQqtOw87gpDClgniUBGzpE0l+xqQTgn/5iyr5q2angWBnlTRK0YqA30xRxKkyF87J
sFQygRY3ZGBv+ey50wbIxk3WBJmHEwssk2z2dqX8USRSEA8QoZjpp/EHp3EDV797cHOHXqEKZm1p
eJJkgdNkwsDX+nBVppY1W/gaDpQDV4hx8WrGrkvlbLQlGAtCOYHdYkLZrv/pBrCFQyGKvySB8eck
W8schOcJaDfYqSmAvtEihxAGk03egd8VRAiT/16u5auMNKeTl45fJWXhZU+1B8jxDfk67INloDQs
yCTAR72I0htb04/epEb8CXmzl+Fj+o9LxwGvBZ7tpxU2fMThO2QTZxrZWRazVMFlvYIlc9CTenkH
MVjUxAx16jCs+3omDcpGhGAtZybxjJD23mNdMnB6/zygBJJP46j3sCy9QLDo5fF+fTqEKcoFyrHe
GTPBfsqYm62lY59jZ6EhYyFp4Vf8VTfYX5qv/DO50qoeHrFZscer78B5XgJWCj5X2/aB6uBWia+i
qdi8N6YfhcApcrWCJGfm8xROEMup1ueACSQLx+TPyhEdVvXyFARCb2/T0Slm+gTo5o5Ob7GnNgF7
Pwm7PoAMu2GH9DHL4LIP1SrYn6eSShNgpvOz+lrW0DhDkP4Eq1wloxYpZq96tQZBrDVaSqQgxRPA
PNUD/nzEa2s7Yk9u5dDhjdzZOdCVd7czJsI0OrwRN2eINzsudZDMFGSTrd1Hw2F2QJUzLA8wnq0X
t6uHLAMJL4Oy8SRPTz8jiJvPJbYIWFRYyN46QHD+IcBHyKR98fAtNoX7RvkqARei9YEQD98kQaEz
y6gRLt0Jds8+h3M3HOegWFKQd2AV89gxb8JjQY6RQAsvXox3lYGLUN2R9DaP3pmuQVA0jkaPn3Xe
o5ql30GnwvJHD5RUkJzONR8D4NDTSmqIGrpAA1Zdg5ym1e/HZ3hXmWM0bPdCRToQUUWFpYbVrJEz
N3COudJmayCxyRMkt+RLkCRJsHM5duaQ1/PusIajJQpqQDp3NSqWWbJk7FpBdkunbOREC0Re6yeg
u6wESgCkxXFTdrfpedJfkgMlDdcJoEcrrzprexgQrO2VHBs1uaDKHDmgOx9yR4zM2USctDlWrnBB
V9YcEUu5FqNJ/3HdoW/tqZGYYCs14ZNAcZVPnI2pD/vbUQRP4+BiFXIOPAE8EjXQ3Q9+1JxCHfRe
cj8CaRhBB7eGlZC1/dAsZX+21kkoZ1evAP4Y4U/4MTNhmKG6H3jQSjR2aTZtokbjV8YelwujIcdQ
c/OAsEGa4tXDjRDMaCiZ9CW6Gwm6o+8u7NvEvJHDB407VNzMqzVxL5Hox5LvTDF7OPIy9/rZ3+DJ
qE1uQxfufcyP2puCwti89mkye/MMtUIsXq1Wt03nxFJ+UiKdS7A1QphZmHMdWxuEdQAJrEdJSWCL
2x+JtouPLJXDPIxSxzRY+D+YYajsyYDlsFFbOoey62peXH5b4Anf0JovPlsL47xN5Ebf8PqoXz3+
YY+YGJH1IsyjK2r7YNJxg2IyjimIxXFfj/5JoF0TSynkW5o4RPE0e2eN07cBcRD9i7lxjfFB4Zg5
THtsP7727HnXleU85uz6DfqZkFN8L5FrIK5Z9yIpD+6DMmCwmbH+bN9v/4a7JAKqAUK5rQ2in2Og
O3mFuWO79lVV5s/1/d222nSQr0yuZr9PX/mchO0wlfJtdic+cYuT2y6jvDaKJMhzVCXYReE9KkIq
vqzJxNYCMSKk7EKuzfnOvLZUBtsephoVLQZf8CKfT58fi0j9QDLe9I0hH/gZINh+bMf5ryyhm7mb
0WGcxJPgfMFxqihuSoEMahO3VD1j5Zu0J+xXgutxDvA7nm5scpxZtjmaP6eYQ6sQHTdkU5GKWu7j
qLWoNs23j8vwEBlzyIUQMFFpTXvnUm0WCxmRPIUZcJBZQDUoD1PyE9HPSH2Rb197Z0drVUvU8LPZ
rHJDp1Uis5dT8JdazEIZwCcHU+oqgHWIg3JCp9edelEXvY+xpJYdnXSwjSYUwpCiv/yByPZObjw7
MwK879zQXtiykLFhl3md2KFKhMRVDBQGpK6X8OruhlWAUVzpKxqBG8tsGFjbuIN2Y3DFHvfqsEnW
nnPjCFzXejTKjC4CbPQwywIShoFeSR7dH8SPtF5A/hrHAmcYT8CDVOHYKpNAJlShP8KMgL8HnRVO
q+Ym4//YFMv1eUd/W3wiY3tzncCIKTH2brXKBAytJOksG5F8DxozRc9on/0MfRDrKROUzig5nDUa
oyjIymLJdjNt+88zlGPw0WvUTNxxJ1H0HSa4b2sbDoKh3Mof+xhVW8BDbBKCG98poli4HslfZfkZ
5qDFsDrJ+ByD4FVJeyRPYoVZ0EuDxoAPiOuWzA8NaxGCXfIZoyQYRnFylHo2W3D2IrDF2B/99MNI
me0OMxco2md5kw7jBbwM+CNEHh/kKGX8+pnmUzorOfrjfAZChlHAzlV3aMgoJN1AqHJpjyUzqafs
s/n1DWQ/hZgaDQ46K+4KM1/aYR4NefRnIJg4frzMoSwVTD2g0VNhGRCec8J3qqx+OU8oK7sZuKlG
JtwiLcvpSLKxazFkAei5w7o4laEMafkYrPcEFpPwPYg/tLG6KzIt1Pp4f82B7H/86nzZfZt/+QwZ
Zc0U8rqPzp03pJGUWZfLQ+cY2+L3SEqUk1cM3mxVtmcdrL7Db1avpSLA4gwxKElDloQCgVx/1thT
uYQYcyZwL8SNgEb3e4Hwmo+LwQxPwu7dKEx2S23lCJQZwDwWQrc6jHrVMXYUZEl+YOyU6qVanrpE
owMhkzhqrggK85MQB51FgSuMtL4L5dSUENh32cUf9NxoJZLYMr/zZwbjMYEq774+XaAuLq/SCGK8
PraLX9dKiZZ5Me2LuYZzkL/6+lMMGsU9QctVgrO3hgZJcdpmE+EsFcyUWnyJI/UBHPK20qj6z/xF
cZ4aYv23T0fwsQ+twrd8nPTcv3dth8YPjsrI0Aj13u8IuKZWGgQ6veqR9G5WheyTulvXgbCrfMgE
62+6Uu1HR2527U0M1vObRxsZa/5JPCuQw+WOApEAMiKxSe/mN30diIMEULY9l3v9pTbDBFkrjO82
MoAPfrrXWT6kXP8Km68lok/KfaV2YU26tFcV/VQqqus3zhMYFT9Dib8jcmS9+34tx75Tw5SeqKWB
R4k+eZ+mCH6lxDxYMMWX4EmwcSFhLv918YxK5ZHGE83rFdX2qRrMlznE6lXN+w1b889YhfEXQtiM
LOpULFw/rerCbFeHDI1LQKZKZ6cRLZF5Ngo/lZ32I6vCOlJGT0BgNrjnO3jFlLasXAeuYZqh1nAG
XBWdYgSIZUhrV1aeIBcxAddOdbxg0CVF/vuFy+t4oieGsOglU7rnUq1hREeY14ism5S2g2iAMAIZ
tZb+SZHFyi8KI2RkUrEAh2KZZj7UFZlP2QtX0ID5BdAl42tdEPnpd0HlgSIwhxgUQeq1gDTf83zs
hYvTYe7VFbGCQ7v8W+zmPlP/9ixv4GKhJ449Ms2MaKKTgJCG7L2Pic0S+VrAlYhEm7jeuXmKBhiF
k3FctqwLGlwoyE39Y5+JCMUSiVcAMatvVJw72ppauCWCXgmfFoj9a8IEj7+pYy+ttQ00rW37ELA0
oFk7/d8VV81l9srln/yQI4wI5rJ5bu+Z8oAhSOpDX2Bm1WUs9Jh/a83uOdLBskmqXBKzdVm7MkH+
IkdkNIiRpZMg0t2IQAyae9KWXS3bMR7HLoP4oqqsENUk1z4b+p3ll6jrZVTVugjPmOda1QQX4hVV
hoyRn9BHqUxougO5WxsAW96rMnq8E2OTAv7I5qfy+BQ6XIqTKq4fS/noDdG0JRZXNqC/Bwug9wq0
MbXDivv0BxZqw3INWStyymKODbU/VE6Une/2+OFUoc+oNB6rIkWpSGF8XCODPGeqsBc85cyAbEK/
l0ziAWNOcgcE7TDLeNJTKd+MlmW5ISVwCds1lbY0ex/jPy450yk5NvBGTNkicLxCJJNL5DiVItyi
912agC/H/DqmqCfNDaZWJyUR+B1nMX/uUtb1G1JFSSmO2qcNM/RG6nAnffDvMALfkJFgAUiPLjnq
TsKu+mfafR39GxpX/4BNKE3roWwRvQDqyqBjlfhRccfr+zmy5I/dkw2BU8GlZA5jKs+S7iCmLiNp
r6rEK0fpqu+0bCxXY39220CMgfzvrVFIA8SbChcEinNRYKbz5bMfP8IqSPdpUqOFRwNUfT5kPpHn
X2VYNkxq0LkXySJtgtC5QKAypu7dIcHmofVNMlAG5Z0nfJ9YlGCbxyyZOhgytOOCaNe5zOLcNOzp
IXtWZ0pa8bhzaFpeLNLTJ8uA/Sit+6L8hL0VJgnl2EaYfTKEw6PpKR4ffx5lXKjPB1YLv62AqDwa
MbzAkWE2IWIZDCIepwgJ0No/douPXYELJwERkYr9MHaCAzkpW7hlCEw1QExlYXF494ebKySgh1N6
f5u+gorLd7oR5x+ZwsaZhMTDLBUWV70TcEkr1rD0bx/Iq7+6axh4VxSlt3hDMvAV7l3dE2t0R5Jc
ztuCurvH05X1DBkLl5ibp26Tleq5v4uVPnT0O/yaj6EVRDBcundzXi5eqEDGIZA7hyz1vij10t9f
wPbyG/36Dd6GDO9PGMxCvjn2PnE0oXdzcj6pot/0Co391JQiNT4mdZHHhdk/JVQYkmZB0soR0kXC
fsYbHC0KOd6vRFKvWjOTCAUkhcG2nEJpCRqmysHd4u/8hgowcispG3hEnAEbaqa0sHRWY1YTSr27
V4C3r1KGxOUq5TAIsMUDdXdBZdqLdNeqzqgVEoerC7Z1CHyPeZRtrsXGiIfnK6UACH5kfn7iHXOq
Yats9Yty5X2gBk72XVsMSsDRe3SAm8qrsazl8WoVgSMvQ8vlWJ8SPjymhnyyLLO7D7QqDFlHCnJw
A4162g20Wz0pKxev7OTVf3q4UibKk4/Um1b842OTraAgAVhF/GsGYgJ3oTg1NMUacb/VQYvBV2KB
k4ijyMNSYeVk1IsY8gkctA+ntGsnSK7VlQOtH2b00wywqlup+djF+aiFtksGfhn6SXdjgOaSjg7j
43Jlj/K4MYUCCpj+RrOXxEfF4a/TbwuV1PW0Toi0Iz9aFItcJaHE0G1g8cbsvsX+yhcrm59DMe1c
I7m4D2CztJX2aMzEz3+WqtuiQa+v9LFha9GKb+1xn5wIT8k3PXQ25al8p8mdqtWErOrcbIuGBp5f
VUnYxLeP1f0O3nsnr2OFqf1ORpeQ9qsDANGXP5gZzOuL7zmEmrosXwg6TMU3ZCpbdnVNbxRJ9nTh
VozB1xmlU7+uZGhSOEkQ8kFWEu1jpgP7WdwZD2R5bziSncNOVCd58t+/YLEr3Aw0SoPtAUJUmgd4
NLR/yTkfAdHeooHkPdynecmUcR3Okh8j5jtOw/h0n0feza8Ttdlag9WNeuz3xDrxrWXVAucep5UD
scJDKSPNwv7A8iINIB7XbbjiNMj9ck7DB3aiR9JzNKGGW1IlVaLz9ZZnhy/MnwZ4eh/YvgCnTvY3
StYD7sF3ZR81LNBEF4GToIafxzjC86iDJVy8GZ3g9GivNT9eZpMcIW4gJGsuJDy6hBcgXXB8FDhk
7kQv3NOXmqpVB2IbGICEVktvvGlZQTAPWKahALz+6mjjSRZkG55TWs9medYD5INOX1F76VbJfG+3
IbFOJzhWrJbOpzjlcLHoQESLfg0OZ5G05jFl3hU8cyMwfJI9/jhxmgqiW2TtcBH/dPeotoqfG1da
Y8XAfYGKl0ppbAIldw7VbFHLSS73ZWQFG5aK2iegO15w4QlNnDF+b0A13FTXXTIzhVwEWL5t2Wbd
cYw0BsxE6MMYRThHgdsjIOmg+vzt5Y4c6gZUQThXPzPd48nwlYQT7f6YRX7oiwjEc92ZsQlzEad5
LmrCIQyRSzm8B/+MSzhZ8rlaNuJ4hh/zm4Dd/Dj154nIMcjmfeDDmZymh4W1Zan0FdHGyKj/0h0R
WNYfqSZIKJ2v/koW65teG7xgmzW6Lzt5fO4iHfiyq9QYYUwJtZO9O1f/sp35h4Cgm42ApKJEu9Ju
j5fXdG6hBgsjJsB5Fgf/cPJXm2TfA82mCHqvA5+nUja2u5Kejk0lVNHDsGA71WGHg4rHHYHRA3K9
JAqatL1rcU7iMIOIcPWB7l5dt4NsyDp8AypTRYIg7YOsu2e4F8YEORo6PROtwse6G7rl9IKBzf7U
X9B0jH7kkDUuzKpa5fRHZ9l5MP/b3oC/WL7Hdkv+ZSEjfvmyzhBXQpf2FHrbpQgII2Ifyg4BaTq+
K+sWPOqeq+gAcRFlhKw0jU/xpHIDWmLvk6W1kq+F0Y7KJsvpDobgbTGEFEx1dC9xSgshwESPZJ+H
U4BLp42rVWKT0/qp7Sm1eel688zVPOGDwXSIWsc1ICwIc7GXYaAzh4Iw+dSaPZVDeCSSkk/dg936
pqrAm3rcgxveEKaMgGfEABChbQLhPtmiYgitaaMyty+aEwTlC2chA5z0ihwrAp8TXI7BzyfqSd8i
EEuRu97QhDzy4jA7YnM+CQcVNg2PUCY6oZveZolScFcA8CwPsaOJ+UtGI7ecK8E2t+i9QNMxwQcL
2M8Tf8H0uWcr4gjrslKtotKS4We6Kt5kRJXHdkqw8NUBXGUjp/SiaUshBu/h9W9H7Anp1G33UwoX
MdRQ5yF/k1MSXBsiMpaUo3A5L+jNNdIEqDVhO7zGfbFsa2AeUeCyKMaeItL+o3WShZ3sishetKkI
gFD/k1QHzYIameUCs5HYHI1LohrO7kRwwSAd3/GIsbSEfR0eT12JIaKb4IeYKpIgmtkegeMFTiZX
GebOmv4doIRAWMLIR/ZY4noR4F1P2qJMNgUqW3gUpY1yphBmz7f9I/bXLvgnyI0atAxy5pmM7I2Z
l4fsLrMOZLmNez8OgGet+YHVi6UcvtIyWirkb66xTmprzggCIlnnFqoY6VYQeQfGscgC10TUdwhl
xM7Kpf2tQ8Y2c1Qi25kMIVuhfcXGtex3XpqZuVCLPO20Mf4WLEVyBMktvCG2447LcAylkDI/pc+E
SEvkJIQp5vJjjz6+3tziltzpTSZkpbP6Tu+zhOAFr1nsrxxW21IJmSfRQjH8iQx8q/sEWz5tNYd2
2orMItISqlZOtAt0KmzME+7Imqe+yLLGy7RNEmRhqtiNmgoO6MA0XtTcV7KnXLrJqm69q1TlY0G6
HfqGuwvnChrpTOfAbEfS10QwsCYJfsp8sUMmqkBri4LvFWdXopuRUxh0fqBjobF5tYzL+FpUN0eh
DceSdAlDRBB2x6ldS3+0gNR/mEGev9eBUKOu8C2WN9lAJabORb/64oT2bg431b3Egt9CSU76UYN4
L6jLYC3aDE6f2ufMGrYsHnWkTlmvH6S9RXlLSG5COYeQf+MdK6xLQfvshM1gtYgJrU+3c1jMzN6L
6uLRS+QK4vqzbOdFrWVi/4wvaQvET8UJDzS5TUmAcOxnPEzHMrB84zlIxzX7BuvBhNgzlGgs31fn
qCOq7KJXI63CaTci7XFWT3twh1FEoPFPzq77PfkWkGRVmUQ9Cmq2ShS57M7t/tugSmXGGCepIP3M
+JuGdeo44prXS3bsBiMTCXuyWVsV6Fg4ZlwHbruoLO3RMY6aUdICnDiH+CNEtL5NSlRymZJU4TBY
b39CRe2hXtFIWYd1Z77f5QPbCpmmpuSBK6DZW0ATc1/6ERfnSiqfkXNPbpNWfRaTBrmzEatC9D2Q
AuJKWp11dGKHGOP1YTzbOa0HWRGo42yeGj0SzuV33jfSiwx8E3gAAprpQyAfZEmVB8fEI3vYDB45
NPQFPUcc7Zf3I6Hm2ZsWqJnuR7RzQjiUI8fJdRWSMi39Av1WTe/JvYMYt+zoCGdtIbSg1nsTUTpc
zKu7Q17VB86kBt0wOPUphmsF8q7w8AtCT84ShR8yPf5VMIB3tmxKe6bS6OZqBf0dpWk2euQs7wc8
zdGL3qKPiCJBA+nqFttOsMrHtAfeTTG8okH6AVjVZpTblh34iwDppa5esi7doxDAijYDvcH3vzUA
cZsCGlR6gxsH3Swl0POw2lI0dcw6jRdmE4YgFWerg0rlp40xnUPpmYajGYJKRIHRUbveRNG2jKJG
i6VbcWslzHmBnb2hTH9JjBpkS0Ayw3IlJyl523IS7II4oj9eka2Wge0n1U1NsAeqVaI8+S17uwld
Sr1PFEODJgNGMfPWCkK0BGrHaSZpetHRW8kcNZypANAsTk/ArC722e4I3rTnfturjuS3QikLfAmh
iVfDCcD/vylev5x+2FO8los9dUeTFqmKwzt135qZeENqOABVxWtBKeIC2kw0vM9iYo446bcZHfud
4r3vAmreLK9tf5PURMzWnHqoPwygGeAzf2DxTqfNnI7r148TFicLb61M/Q9EH/3Jr9lW3AfW6sd/
LjAgJc0Lzfc1o3l1vL7Kew8jB4djNned/hisTKB2aUMpLcrsHHQPDU/gzAyR0kU8/V+1F+jkSov0
CM7R/1bnkUDRlBoSAA08e0HnsCAOTxXHewfmGgE4NCkzZ5BotERu8X0fhcUgnBUKV3z5SR06KFL0
iHeuz2eFV9mgeXa35uFuxKTadcUnqyYWdiaFgbAnfboX3Ofe/ztfdwkCqF5sqFvxeqfZ+zl+9jX+
37U5TMVvwMAY3R1k7mfMCoLx58gzThGL+0hbH1wXBD6BeCwBk+/AZlGoy/Lrxh/jQkwI8P1BcbDe
lU8DDV1Qj4Gb/Rnl0OxPrkm3H+9QU5Bl8JuKIHcq2pFnsPyaq3D1TUpmkOq4wL0Tv27el5k480Pm
2lHRcjqDtDUuxS9pZDs9GBIwX/JWI3iAwv60sukMyWJreOl9k/8qrF776OpmmwQsUPTvejBDTYGr
3EF5b0PtxziFYHK7iGR5+D98T1WJ9S3g6Jkgfemo3Bs5YtDWaujzohMQ46CMDRtRd2I7yNsGn7WE
tao8aOO+3AOV307NiE48hCR1wu7EYbrnMXq3UJp31jl5MUp+mkoJA4zpXwW6EUPgrEkusVF9BTzc
T8n3tVk3M9YNVQaJWTsYq5UX/iXtvUaU1w5gig8NF7cjIW7s1NJtS04HKSuX1+QY4ww9uxMPS5rH
fanXI/AotsGt69u4wL85M0/eKld2dbFyVYFT014Q6GTikyU81wuBhLXsYJNN5OtegDPjYx4lzOQj
bpbu/YTujO6j1J44vY7Kjn0RiP6maU429eA/5X3etXIwJJ+UFL6K3/O0JNaYcPqD0DyZxTV7tsg1
uZn7XkTeA4SUjzzXyEAHfZJsNQ5EFCXxa+m3RpIgu4ygd6PECXpfC3lCHA+7HsMuWZouF3ehBJzp
Eis6CnfZp/S6SniJ6Q0hEnhjLx9IcARPHNWaNYc16C/cdki+S5RvskazAY0PsSbF6EJCeHdIIynj
AkKhNXQz1omQf3aJ0w0swgCJhGjoO+fRgz9Qu3yDeJQFqbT1uBIMNOIItiL9bYLJrB/gGKWg37fh
eUohlc2Yn9fitCXZLu6WdUvCJgKi6uP3l+cMXl2PHMchHf5/e8lRFE2vDBUd+67XlteXgl9sQ4ov
lVhNUuYEMwtw6RJpYwjC9FYE067FVkd9nwCjE3qLB65RB2RKEITFzSNCRtxBNuAqsL1a1aM1DngI
mneMBc/vDTtNfEgVHRgYTu8G0PYprHp+fkjRkQ4vRwx+acpFDoNpn9reE6K/ZLId3/0YhvQpvim9
DfbSm/SNUOxDMdN0hiimYo1o/l7gRW1tUnrgrjNJl9jf1g1lOGE0d7RdxEjtkWet2WqWN52sGY0Y
077XMvviCfedNTG/h6G9IoWNl12zIOFrqxrT0k8Kndy4iB8D+GWOtTbbA0jTChMeO5m1UmzWo7Yl
JrCH9QwYKZJvL/FUnxF7Q37htHfM1/g+c/KPOGVhHhR82+BvjcLK4wfcenpoTLXtBG37YU8fh6Ul
kWwN4on9pyAQe8aq3xrQSwckD7kaD9CPdzMO4u5z1pBmThBrgy/TXrj9QmHLG0mqmTBargWbqMT2
fSrY3bQRHj/JvsrTwGaWYOWI0ag/f13eVy5BboAdkGAaPKBCd681IyS4uwi/AQUnB/rIajuLawuW
lq2tomiFtlXTliRdacBr3JXIkYrcHJPbMj+zP8smSNmZHZt8vrhZeyqoY/7j0KUfC8MgMIfV4Ymz
ztVkf8/VSel9Yg4hoDDXUm4kxc0o2rUqsZUEwI/6EQNC8yni/njLU23+58tUFrcUtT1Klqk+xrCz
zZjSsye5B6XZtw1+TNDU8GrXF3PiDi0lkuwvU3xhBiW4UvT/7kpx0spg4GH3Gmd5AkF9SptZJTMy
dZ1PvnkI3N+VLIzxF0taL+JrXK2yRM/EXB79tIdQpl+BEEjiGF5ltUeFF+7bkGshe2ba4j62yVit
E05U+SiBES1I9yjUykyufewhJs9FPDkE43G2acyQEjHZiVx4p0Ng+SUOx/TkOftwGFps16YD+a1X
n+4qN1MqfP5phnhbVI6HE+thS7BOd3BHhL9bLW1fu6t27nXyc7o3queL6YpPRmFYllkZz3fCXdEi
BdWun/PDFkVL/nqATC3dtX85aA4o6D6SYp3TFZiIHxw9YRkcnTKasv6Ff7poBlF2aV68B4GY+tJd
Bp51BEHzl42/OQWJZqvogBUShVfUF0FISvPPmqWo/j9/pk4J0IkAzOeCbrFoPLx9mxtXPGtHLHi2
F+cn7fb32fthPxNT+n/GpJNn8QllUJFUUpNVq0Qp80pkCTQ4KqnbtmkA+JOtsm5PRmHTCH8CR5AP
Gur+VVrpRyqVxJbgRPEAmPTKLRy1F0Bkkj85Pmp6nVyFpezErCuktLgHUpXjjm4av7zbut/GO4vJ
rp2nO+gt5EREFq0KLKKrbfxwV60paAAuXrSXw2oQ/j+JH5G4IuMK5A52ew4mTvHMUlMBgSguuzVQ
R5kS2YkTFrATnO90ttXQaMtsQDfvpDC//niAsHLgV02TfJw7XdyH1C+/KdN+tkLesjrMEtXBAxdK
/jnW9fvWrF/Vu7r4g99Q+zlWDgd8Yinj1UgXyNykL2qDxITPcmkyXtUFXzoGuXJq49qpQqGBH3j6
kKMsqGsFjTTRHlW2/sj8zsK7Wnuiy9CFl31VZw267rrb+APB4l5v3wfonE43eY3ps4H8d1lv4C1s
I2qR//CbNKiATfVXOVR2ubufG7qt+zBKDIWs+LE9641mC2Mgwh9/NfywjcnRDh17vTyJc8mdZnjD
0VbYdVL7jyKGQ/FfaN2leG9/1jd/zK95tupqc56ah8NyTOg7Wk6HMbUSLpJ98+w6/8LiVCJopkf/
nwMUS8zd5X3Npp5enTKsHrteuBz1R0/8P2ZO3FcDl3CZfs79XOb7OIjRFixtFNVV+6SSrNB0ViW3
4PcrBg3wYEUIXF/Q/9W2QOrChBMqlY7bDxkcFmN5vbpuQbzyIbU8uDCnP8VEnkRYZxOxG7GM9/oa
RsOHHiFdbbdos5tR3sDZINa/5d1qWnDkdrlgOA7hh7wKWOpzTVbPoauLn1ThxzaSWa2cKiq5M3AQ
xF8eo5cTRDoCuWBWkdHs7b3lz7MOLpv5XyCoeOljtpxCB+t8PjAZVA9XK+Pyrq+J5T6qqbxttVlM
2JrjsbSv/b3JkeQCz571tVrjo9bWUsb0mlCFyPH1K0Psi1FLJ4hG+e9qERbvBux8bAPySqmk3m5q
9/exmginp633J23/G096wvUyOe/cLmhH11X/47kr70cQlrRAxFiFg037RS34E11+hrB/dWVl32zf
LjBA1++N87of4CnURMwR5sL5zev24BFOr8imhXp2qZFqaCuJU/fnrcFyi35/b8sD8yO1qBYVpqF5
EZHA9U6yKvB9dzMFNc2s252RwUhGQq5Z+LQnhqN1JXKkMNs5tDKmGpG8P7jLUruRJYxuCkDhZm35
3Z8QEueU7On5LzDzVpWZV19NlA+MgEgvYNHwCoz3f/L5Yu1de6B5ppdjC6ehf07VsdCBX6K9yO3Z
5YeEf2MMnhsI/gBRVy+qXfkqS4BymjwkMu8eXyj3BK74VEixsT3Dgin/L7PXTt10sDeh0f2r8BNi
Pozm524xDyd2ANXw32gIxy/9T4CmGvI39vten0WrKD9fbxt4Lu5MK6IS9IA62SvtnVodfLF7ebEs
OnXZWIcHTSaG157YmaQzE12Ae33N1HJe6iIwmSHsggBxS/vzZmtz06OeyZDyPmpXSeK3XdlDQUp8
8qrNJUCYbItvOXg9qTFj8hRLM8dYdGfs0FuVivOFvz/Me4Fjr+3/3eiX/odOPxVYX7NfVmznRaRI
iUo+x/USf4lexD2e2oZnotIu+xgyiOkdymSOND2Gel49Xj12dSOaXTK17GQyPin9l4/S2wQ9um9k
uFw6u1781mrWBE9jjG7ggakDgAtqq5Gnm9CSq0a5SQsWCKB6F1LFa42qYWkBBsJe6T6tf/XQJwIQ
j/JB6fiklV7KMtkY+Sngl40ylYzYkfoBU9nTyxBOYRU2+AjLmBuAlq3Fg48jpK3FCnGGdS0svB+0
VfvN0XGDWRZLH9e8gm/OBl5b87AR8vmrMWmmgcNZPP1F/tj8y5V31XsbnDz3YRKWeMq0H6a4mtzk
sEo/i4S1i6Tszj0FdmuLSOmoj7wK6r2PYOTb66Jucw4ydMJlVY8gKzRnAGyGA5koLFz5ZBWIFJiI
tgXgta4Y+jDUjZ+Z5I4gEni0qsEUm2/YHst/xSp9Fra0Yzrz74IF5k5o3uFh50zOTYbjEht5ldN7
LlRfSV6Sd66yn6LUPy/cLDdkr1kxsE1BCEouprdsixEkIb3wle5DRRtdCcJ2fc4CqR+JJ77jcR19
ho0CrNaLhaN5/1tmoHpYSg4COGIHrSjZhGS7mD72bbSemO6InChNTTRWgP42Jcp7GVGbrJE7znME
/+Ys/6i0f9G7iGIU39K6sYLtcme5j31tu6XZ07MREPK4XC5PjuBsCZ3M4CrTRZCl6g6Oefi0UV+c
u5Fas2YxF4G2dYjuJMqNEjz4IVzltQSFIW8rCDW7PAXKomxNlklIvybuuCL7OuJkmIjcRrq5z2lV
Mq/1wb3ZzWLFZx7RLecQe3K+Aa9QioJwbAyp4SmPf8zdccQ46xU4qetCma22l5ZX/ksDPqEHawQN
dNkU+132P7TK76Lchx59xtLlTuWqQY7lCc2p5NZ50ih4/cUs4yweP09rZTh9AmgloQb2gtm04noH
ZgRaXXgyz65pARZW/E4J6UnizNHXnX0eMnCs7PU0OK0yQFqSWZfDczQ2Xr+7H4phXyyXXRYU4YDo
Ysy97+QgsH67TofCAAQdIKpcn8veSedOd6XRyxJH8wqbOiibUmeE0hS6TPVr4izuszbUMW2eJLv1
EfkulJaX2lwVdQfJWgPHS9VRoOSKka66x8aSO8zBD00BWO6TdMJ3KMW2sCgnKogzW2GZvP8CJchG
ejiP4rHbuo8aAd6YN3Ieh8LKOaMfNWUOA8KHGqGcvpxy8Y4csV5+fd9oOmbVxrm1uz7PxnwYK8lK
qbAn9BZcW4lZhyqYKgie2eT+oD5MEG7lZficT8g2WQUZN3XGqYCKGHudvKVEStRkdPRB0ag5nbUh
7NzMM/+ac9/JB2DtbrKV4868B48LdtOZpewOV+4CmVHu6YZuiSkm465N/7CrBYnTAK8Y2Lz7h5QB
8ZrVnjPLZ4fm8qA4yzbjtiEYDNNvPGgf4FfCjs9LRpZj2sT0qIawZMOjp7pWXV+y3Er1P6v5GGFC
lelz5kiVJnY3sHNjYsSMhyHWgPaqkWI0onq5SbLEY/LtCblIsg18eIDwHYF2PibmZq1hji0+bA47
tUW+/c12by94DV0lUhU87LoS2XeJ3G7IzfhN2+bWOVWdKGSAg30fD3qmD8+oqZbupNI27FlSdwFq
IlcABVfqWALtQ/QqOoA6IK8DJYztBL6dHyeMU2wxRCLhph/PGpc3GeDJguh/WH0F1K2O9qEUmfah
klVnila8678jd3+u9HTV/mZ/Tn2CpAoPi4pgW0IptH9vaoGSqYV7vl01YVNxEFEcX7rwyHuxYUFK
QQs5EybGxIOmoqxYdYwbcGV7BlkkLNi54vajUO4xbuBxrH2Q3b3Y56BhR5iM9rLDCC3q3fLENdE6
8NIEe5ojwr1cgfSIxUTRetslzi/1GwWJSkwT+1NOuE8DcsgVK14YHPp0LyypjQ42r6SBCWadh8xF
Cj1Wm3RjKOFyt+ZFjatXxYKgcY3u7Dn7QvCb/tV0/sU6kGRewGhrgR14CfTqo91HZGUi+7N1I7pd
jHfRJzkoKnMSrHXy0XagitFRfd+IPD3xeMf1qBszjbjeOIENxweIMDj8KAeT03Dit89PAGf7K4eT
kGjCE3NtQlGJxaAVQNz9+XExxo+HVD9XJkmjY3iXmekQm2pv2voYvo+/ca62HIDHVwj17LdX7vio
s9YyLHzIzGZ2zb7/E3WU6lVJ9t/vjKKlAIFPPiZig/fgzb4SUznIW8g7u6DemhBcbLw/Tfyzrtkn
A0GNTlJLpuKg91cSxDfCYdjwrUIW9ctB+tmd19amnJYrSe1QZNihdpylUU+KebJLR8ZvthNt/7ie
1Lw5tVsesBPJloNIb0ObX2lcGZ4YLLsbRDD5ceBfub1Glj/fj2w+dHCFiUy/AsygYwp94ai7aTuf
lMJwW2DeAtJC1TzXB2m3Y1fZY0JIWs9rRldTMy4b78DaKoQ93mjCJVgGh2JGLp/XNEbYq2XhXpff
62OedaHcC8kKLAFlSmOVvCZD7Mv12fggWIvU0f9piGf2xo1KL8LFUZ0LQBcJcL5Qysnq+rhulLq2
It6Ill8Wcs3Pniioaz+HIazNvuGt4hkZlyV3NauzaSX2Jmt0vVEkzFMCYLbI+h05FTU1c8Z0qNjG
P9C2mpZ5du22dSothI542MfRmRTbkThZc9FuI210ZSDQwedsJ1QFqa766hiX87DXiaupNGGpugV6
2RG0xEFbkN9sHK6t30ZYJ2NQR3xBUVnA3WzsOz7ZlsCdeHxQ3hMBH3NkNtTo22jdwghpSNW3k6Rw
Wn5xLW5m5BNtIJOWu/F928kMHUahQtBoNLWSBDu+lvgStM23V8DiUplNLsGjsPO7ZzhwyqMUQ53g
dlh3qYrEoEBknDdfKgDVnL2ajrzwyWHyffYM/QH4hr+khbzf3oYKGhSo/SmlUuTJHeAAAv8fhxPp
YfQ1pYqHDmQ+8nLWrLhYgGOD/J3s9/Fl4TVXOGSCmRAT1IzJlolcZrDDtgvbQ1X2Ix0PrADcPwsS
6iHd3R/XgFAwHcRzqxCW9hVQs9kfFAt8Eh/Zw9gObMGIZdkm8/CIAM+seUQHHkxk4mMO7WS1hm3Z
bRmiMKRUbPmsa2X8+q93EaocTZucjGFMlWK97k/IpF9/WHN33TRdCzy6bVo0CkkDV7ItklZTMPZM
U/Lt8o1AwaflOWQUbuMkOimwF2w36/l2yQ0Jvjz1wsbZ4mqsJDtXjIfZoS++hk4VXmkRrTYMgkEz
P1KxtvpwYvtuHIhlHWjG/Qahxy00sNEvs7eJzYFBTUoozdI4Tk93qj0Ume978UYTr3pUigaxnBJt
7zH/wHl+uxu2NFTM5rLa1JtLsAjQ5+rmE3G6q9Kd+S/2wx/SJ/6jBw3M2rM4TAL1DDhKIyoH2djr
iyK0DOQ1JxAf9qe+MbQHZml3vniJVUBIuKTW2r8CQPIIFDTjTEgx6hFUBP2CBR1xsnGoJsCHizmk
7a8JRGBLHk7CnhcqRMSPm9Q9RCrC1RJha3x72Yhu9Mb+jWe41XcTEeQXsiJW6sxYDX9QLhZ0DxEz
51z2K/jdzmLAfHavLxoo+F0/F377uJLs0kJ1Skj5AZrZW1QyKnS1wJCZ/Be+oFULu0/IUWnBpBCy
sfYuMpJlhQj40EAEOkycdbosVaC9AxHQHjguzftm1HnE9nGd5Lk2UR2SRHQSYcch4YteTJuLyrli
Mm4t8JzgFpn42nojNa4GY5/FYZcdUYxCb1Tj1h9vc3Pu4F/sGl55nNWyLg2mIpuVyYIXLZkT+DtP
OmWg9L2BW/ccRb8XEpiBLyKfjC7QsaONzZ2Q2OPpoaPZBrcqtF8SXffToyPL1JUP/OYYlzClG/x3
faz79GY911iqY/CLs3lVRm4ISb5v7ydlLzEG7pttkRlDg2CbErmTHuZlLmSdaEGXaixw4+9BIu7m
CeDlklJdFUd57SD0YbKS0TI6HbKIJL4eC6m0yFY3t3QSUPMb2zBF1pMiLFsry8nzVVnxsZSSdFwq
4TuYSqPVRAG+WoqTrDhI/x0nWMnHZQvZi+9HEEeQon5Il9WNEIj1DxByWpt9/KgvXnurcU53VLNt
r/yjMeOVCgLD/dZlUKCgTcUGV2J1FRr8TOedgQZxG2QKEuBrJmRd7aTRcLph2yPIucoFt3f/p5G/
Z/4bdjLlMHND+CVprkWLUTUAQ990jaoNMvVdZrwgXMg0u1O09Wjejm1/lQl7aIwsqlF5e+XYG4NB
dG+tQd1xnq/Wn1kdwgNOjWbYVniifxX7qVW64rTPnwHQS4MyNyZ3CfLoE2Pl5gnSOBmfJxkV8lcP
TyYsrhf+5lZaAVF5oNspbDL38LLz7Rcaf4x/sNXNi2hIF855ewCdqg/SCl28lBzcWo3qCCCJquPB
nA2mcUYEKkZJdUD6NNo1lOTqjEuJZqXvtIRU99/hThtWNwm9/9qhpvSIf5lF4uW2vSpX7EdtHyzF
YetqJUSJWHMwQWVx8L67EPE4vYXQUlRWpvcd1eTXekEEO5AWOs5orzm2TFrDwdXhgNtQef26ZXT5
KccEXdqgLEGEL7I93764gzfZGMm4M6Ndc3PqUQYhQj6/GF6VQhJjZWUkvArnt8fN5Qc9GtOoDyAQ
1CFECz1BP1ulaw5KzrvwrsW6bBSPzCyEz6elTMXVmlA0UyOeSWdkB+8kzpSu/gbg4d0Kga7DcvXa
XajWW5mazjgVZFuoYeOkdOJxsqin9oGnDDFxIQSroGoRQxMPAsGR8ohgaSz6myI78WDK+3QbONns
pby/dlPGEf5X3P2yyrxwP31nJGl1XK7Yl0ASMBrApaKefH+D3g586VS/efCRjx3QpPBbLHnNHf01
gVlJ4oaRUDNnwyDJ6U2vOtcMCy2HZFuMSBwCZ1F9QxFCocb2g4433kYorZ1IHa2ehgL6AFcMKxps
WyqZKZ/37Vn/HkS8UDSmoP0d66jq/ut9RzNss+rWCrqsIc7iD5RBiVltL0A8sHbAFBjdpqYs4oMp
8/UJ/6VtxYN09RavsK/7yPhy+XSrDoSKgpPcDGRMILAcdQhQvShAUeEhK8wHbdVea9VinTrA0kmF
BvVkvzqr54X8xPs9sBTU58/ig96J8GX9pjtwEaE61D8JsyNWlRpTzRgq9oAZf7r0lsjlB11IYyH8
H9kb7y7n2YRQC6FW/ppoMBO9t1wp8QwqDbtX0V/e0o3+a45o6E6vOZ1LxOX7uxWPwy7xT8/XzJc4
0caH6YJFPXqVe0uWAbPjWgeCr1SQPf0OWYAXCBX6Fo8iuWF2cw9MIvjk9KgpNlw1Q15evMhXrHdd
IGiwOO8f5JGjCz33LfYU1pY+PzlJWZ82bNwQkXEGjHr/UOkHKlH3zM5heN6eqJ+QdGm7Oe5tW2Sm
FQlGFw+dJVkh7G1MaDWio9mojbnSP5Nsq/n/y0TPxMn6ZnCd/PFO1gxt/3Pl9c98OPSQ5Jo3eVCn
flHoVNPG8V2iShG8zdmjaNvgstoDNd2hzw08KNlzrWXk/9r4GMX1oISmy/Mnsi+I5kZGk29JM4L0
EdxPuX5Il16S9+HSVn8xVT79meX6extYQ3+x3nHHnftX6OZXYa7Vdv9L0Oy8STAqv9fHdwSNNtKX
Wfy5gmvzJIvDl1UjhItq1FPiB1JbxanwqnfQzRDF2vjyqyd/SoGP9lnEESgt27ixb2WpUzoSDnOx
9izDN1Zgf9VJmOx+2gkKTedPsj6jjzbEddrgQ7Qc/iUKQlEGb2j9hYEEGRs5Uphw2BcENQRed9gS
vznbO4QPshnL5i+CVI0mvMG1PMYn3p06RB4fiYYv81hjxCPjVDaRq+5Xm8ecNBcWQw2CTTjzzis0
TiMltM1ofiKwegcZqSiSx7orM8qASSkJidQtDhUq/iYrBnf90dAPAYbRo0qzchoQa899+gC6dfz6
EYDGO15hxmFPfYqFZkKVEWTYKGWge+WL2Uw9SvNNR8CcGxSVk5tDlkWnksPlHG52OP3B+XBokcuS
CzRFinIk7olp2/enlxV3hDQlrr5QMX0Y+sGkhaS4GHYPSSmL/psO51w1Pt7o8U/QghrxhKhNPf5p
CpXUNMfhlP2FzucoJMpW8YSDiZtlecoo0m6SwMfPau5GHN2d+nIgu0d54yK9htLayaOLokbUqvRx
D7BrqDC/ax8guPIG81FuC72BJwMvssMKpmrZBSjnyK7YI0H71nvV/4Zi0fL9mKo+CqTQ73riHuKw
ID7xuA8FAcf1tZVyR8Qz7wJ/g196t57fgoXzlXVwsDSSFlUum7s3nslJr7G16bVmDqRY7WoDAHUW
gsA1TjhkpRmBIBJbD6wUK7FW3TaiGif+D/ht8Zc4KLLYYNUYwZlB1GGfLxXTl2Ua49+iEvr/oFgo
RxJ8m5Tg1Kef9qrWliUYixk5/YYoWL9154CwKHLPpvasbRuaRV0atIvN+5etmfIE1F19zYGL8wac
rLJqJ4kOBoc2IOQViVIOglDiJfxZjGXzNrLrFKWoAoMZ316DWM22QRMpmm8d0b+RdPkhIcPx1ZBY
LUBx4x3H8xp9ltwYB1X+5rTPDj/ha64C0gJcgeEpyVkJzTuIh1zxIwmFdVbV8hYwStKSAg6/8qh3
Ba2NN+2IBXKL5kONU8hljD9Tl3dWmM++Idx1XiHveix3tKeujzqVX8oxv996MZPyAzNraHF0EbAw
5oKxpGF7/vwT2xpGSU1tS/1CnfZLsMMZ7GZ5RttZ8Xyo42y2xwoxLErPpeq2PPdiHl83VrAACj9W
+Csnslw3hHik6VirrvzaGYCKoj4+EybqNb1xmtQX4rtti8rL/MsYNaNMa2IY+4PmZWxl3Keash5a
rNrLfJ18d3WIJ5lgfmNmz3K6wAQKYkKl/p1/sUAWzFDnnT6Ki7EO+Wj806peZp14v87aXnkuiP8w
r9HHhyDpiS06XZujBbpWYDTZMdlNDLtRjCCzvY76+rUVDOVaehDDSesLICg+N2Pj6U8vTXqDEakk
TzSF8d67pnSuHwmV79jQUG3VGpL8K9iZw+VMUhgy9BhM6qQooDM2EKE2eBUKm0jK/VdwCzrWPcUD
1UU4yn0vxQPew9uMGDi2J9jE9tPEhTIr2nJFsNzp59zNweF0rJP61Qm+45y9t8DXmh9qL4MrpbcJ
9k36uNC5sVf1nVlv/eHFq2wdIMa0Ux/WkvlumeNzt4RP9j2gqWqAVWf81eviBPswtbUvS3Fc5CIJ
h6v42/btYQ9e9EeAdzkpAIYrFF7s3DEnplEP/GSaxN7zd0kbk4edZFUvDCC5QiNCvBc6DAeue+xI
3UH7UgvtWb+PNEdg2VnLGsXqiGtrdMPDakadnho2RqyQmv1eM4qry1TRNtQna4Zn95BwEHkieWoQ
9RZVePYwXbpazAnMC0+ZE3KpKeRCVAHf/VNl9v40rCay2uJ48P3AcoKUi8Fn66dgRXpvYtFPH0YX
LybKK5OXYyRLoiXUprLSQvqn6qdA1hweByIJq+d+PNcSTxnjlagCa5nvx+/hAGtFDo5/QVfEn6Kz
YcnEY/XT6lVxOeVZiPUtLl+7peItHKHyAs2HltTN5utDoXDSzacdDOGE/SkKLt4usr0992JVsdvc
wRZMEoPpOoSW39qgeEPzlWXY0wW3gSb1NFf4Cuo8o69Fmy8jeTxwpig8+msLuj2TGlLMBtfNU3jD
3PTG/0HLdkkXQ/x+ktiRSlsaLHABgqQfnwcXIbAslrbJftb+xlL0GfxZZZsfEt+K0Y00BEwxVCOF
QnqIVIRTZTBmOicZSxxcthEL0XMBzWQmyM2WDn3l84Q7jG5i4PR3NxyuGP7LZe6rTxNazAl2Q2Rh
BP2zmFk++OB+0qOg5kBz9Tl6l5AE35Tjb9+K6D43kqmykASRnlgqTu4l3N6wdBXnSXvE9g6HPOgG
RgeolMmQyYLNpwc9NudwvmW3PvSDEnWRZ0EMf05J9/WF2NDQLinoev2z/Ea6TXG9U7GaKqf/fqW9
GWE/Ng+UVUarVWQCrFNRMenQArOqssoU3uxqPdRF3WXcl0eMHS9eyW+Tlo+45SnYQJUqeDR3c+8O
NR5Ax7wrepkMA/u3ccCft+qnGuTadp6H4Dg/qtp8oO7DruLwhblmqBjTJrMJQ3Frz86KHpmU4qnE
cJYrndPXq2o7qxuh9TUQxSsE6IkgB+IQXEfVFO81jr360eKmku+pLsXhYbNsuJigmtpaAP+Sxwj4
ZjubhBJWCdsJglB84ayX97Q+aBIIvVWyqEtQ/9P1srvd00f9MzIQE0bxcAy25sxWE4882bgz2Qfn
nZQ8UzS664L7xjyxmciEqItNnY7fG92JmRRWs5Oo32JDKJymAlr7VUrJ7Bt4M6a1EB4kayeYMWp6
BpWUzv0xS7JD6gzxDTQIoaDdqvE8yLSPLctIbzRRuwOFZYH6bXCVc4A4CH4tvJgIIVccJRvWVbYD
DGktwxsKJQw/GVr/sQiNQOQfbXNpb0LOK8ljzyjIOvObl6zfmeEvgnv2OEjRY6BOAJam0B0LNc3T
9FMwRRJ5LARnCy7TFfv5C/Le5iymk38G5dC9j3+FnqVj+UhBX60U7u246UWb47r1W2az/XqzntZ/
RQtIVjEneTjo12q/lNUKMk16AkDXBUUXJWhH2wvAuid8wCi0uusAbmZma5+xcgM8OEP99LqAeZ3W
GROiGPzZDTbDWRehRRmLOtjnGs1z3Tj1URXCfv8WLRPqHep6c5tefNkCajP10ADH5acwEVLIaez6
6LodY0ex4pO5N/uyrpZmvJ9vOy/xoA/LLCIOJCdsyztWE+jMlI92AC9G0P9UUcAsEjL2m03jlbjF
Ha8+B0ZcNfD8pxC89GhTTGXgrdYvd5uX/BfkcKaK4Wf4khSoVMnWL0bRusRfShJBt+FO09kj1xQC
jeHRjNvZ0iGJK2mo+yBBToe5n8Qc5Nr5KCFjw2uR33Dm+cP/3iGiliQMyyhgivwTFMTIS6zBkxI0
z0bReNwEShCb1K/Ox0x7fysGsL4vFGShdGWsNBJg13TgD7tHhbFVfjCBAifW2P93P7wRknYEFhRw
0zzExt6OVzaEoq4nGhL4ygA8NMO+9IueAYxB/8Mlb0YhEM6ox83YG2sxs2aP9o1SwFF57PfCWcML
8FvblLwXgs4F8yQ1L3HJKGqQSge3voVRiJHqPssc3PA2nflB6wpLfHTfBcVxr2l4IuEfxt2oT8sV
jJBYywFW+gzsAzkdx6A7GUa3/JHbkAZOY4CqM3E1EK0o++Ux8dvn+iIKOPObcyWrtzH5fKMwYyAg
1ovxUJgVgCeSX4FRA0JkQByRCwZOS03VNcCMwZI9YI+NAPVzm79Kbn9n9t3I1p7GQKim2Z8p8Eej
RJdO346nwDZ4zMwcwc2QMh+riM/HjUBcoBAyN8MIp51qIDo+ie7Sjg9/lXzPOysUJKhQ6eE1P9dI
BZdjx7JLh3OADtyWED+8gt1AyKtmbgra7yWEZHT4lSVRUHfq63T8bJIuT9lo3lEX9uP9erb897L0
MOoq2Om3n7RCrgSMQFVKvsAJDtvGV02hCbkxyWjDNRoQbFDQ3Tkbb5GPFCgJ35R426lPx9/IIJH6
uLTwH3VYSrHL5LhrYvxvWJIkeJScSBKMSEehkjU61N8zbr/EmIO76oRtEmsAQ/zuBwbahTf08Lus
Z/Q469AnKvD0rOPIwREhUwvs9XKxtdFofgxxtlYTFNrV6c4W1Ty8GDudEcVFU3qVY7i+LUYwzK/L
o5W5ibo8r/Da4bbxPRf6RipiPWrjTMP34TtnMMObgLtLqfi+giQn2BOCkeMX4CbpfJNKrV75aEFT
5MjJooO/GNpUYdY5Z3oybjpSRORcL7p+GXlD6DRVAzH4EXKybGcJr00QbGTUquWOsqqKsZqaBwzs
VJPA+xp35W4Hw2dLfj8r3KnouKN3w8dFWmnXPiGTGZm/k7oVwdqU52lCszgBxxPChgKXVGKChabo
hlUANQ6FRNSnUOlgrTk2sCB0QRAdY1ZdVtiCL90xNWBcPhDyeXlwNyUMYHKCkhDLyY9gOtK70gsf
9lxLQLrGjGPaxTUIXsRZ1MfIO9ezBFTbBPvvDP87x6zl4oFnSVYqxzwj6N0M+JxYzO2G60BS4JG8
dti2fbKmDIl9b2AMTLjtdmX1EGirwdhMsCzDrs3jq9QtnY3SqKWjVXIgBMJpe3bJksy8FaWQ0/V0
N/Dt4ravFaACTn07SD82xr+bUhfb0iwUqMVpm95/qo9OUzjwTB0aEua0+bdrzeXnGAiRj7dRbDO0
zqh3x8zY9VeDDcVjSPaMnWcKXSqdDeKQ+CQNU5S/1hBRIccineoP05uWD4rZUSoT7uwzQoKXrJ+w
Qkrbp7AgnehFzMnlIJk+o8KP2mCv3K60yd2NJy3ZIS4Y/agaJXgHRdri5ZAlikYIZ3EkTQw2Pdt/
zKtZtLDkf2ECED0NpPBMFF6jISywEozRuz3WiOSQPV0DATlnZRQ/9Nj7TlumvSHBadc4Y+PPuEpk
NuJgwKgbnCN40xWMrjIl+di7DuRhYZQE66d8k2NLhjYG75usNiOtftWdzyI3BsQwYV9sEMFfV1HH
u1BE87QyWuqRRuhGypxxv7zqSAjYyElNtUTRpVYWolmJDGRgsDNwTK64ml6yBFEku/QUCxYCvKPh
lJ3JuvzYkRDyEm4No6nOT3O8PVxoViyVJPo0bivT/wuAnpK6hSxZyvl4so4veiCyUjSP4dfmyAdX
ZmYRUhwWw1y8rfHbyIXeIb6fXbTvHWZZyeR6D2rTba6KCaI8Oix2xjIeeqDmfTb30lkKukbLjKcW
Qptft2cU4EP8kcDifGujTylVHXIDErhEISti/1F/0lNdms7Oc5EKCbZP3GRqmob2bCGlzO0UviKF
oGOGN6n8vvzANOxtGs2miYc0v1coERmXeEZFq6u2IXOAIOBNZDtzCQw7ZTrmRxHKfmcVO1S4Jikf
+I29Daf/uqf8WZZTdwZ1sCxDJ/gFPsJES7DxwJ5auqVi+167YJbLDL+dgmb/48Qk/2tipCRbbwH5
Ov1lVzN92KR3ZbAuWRF6CPdHC4wEeIYdZcTb9bOQubtsULuukpFEIkX+adixEWIIdshzDR6XBjZO
XpUxdAEK7al6Af+mGR3tFAQT8Zm1TJuXMTEZE+e5YKlavu2Kp6hO1+lWQMNv6QlEn039452jU3vi
Q9NX/m1Ni3m1WqaWktSPpkDwQ47Q7uEHuTVJoRGOwIPq3FzhKjvjM6/20/UVJYjIGIpbtOEjI9z9
X77cmnhSSO8sQTtqjJfmz2lpzeUjgdMu8N1kldc/iW3E71EchD+3MAXKDPLnsielLkVRmeMWNZcp
OSJ3/VhqoYn9PKUxtfxj0bJwd9DEIABa9l3JXsLFlQG1j6Nzj3GNbtCRpjD1U7BJBSZtc0cAo9+N
0Iag0mTQ79uuCaAPIaRVyougtxalermmXLhSmL8jqQtgVI9ulFahbBLVC8jxQMppw04imZWqQd40
c6Ovo8wGvPs5WHRsNQeXteT2fqtZnfci4uFoCwJ6Ww7554NXFEi7hX7HZVrP/t8qv3y7VFO2Q6qX
6FWfotHZ2A8r8ZA8i7TGTf6nVQvgi5ff6Ub2OHG3m5o/fG+GIn2PxXFUuLXLORnPFl17PZAYtlmF
QyUYNDH3ZfsI7OQQHGOLgCy0Wf8i6XIfZJl6cgQzj7s3iloUxLI6Tq6z8sKSJ/hjc29IU5LLwA9D
ZS+/rfOlLrvRkmqWvvgLhGQywyod8axDl9srt8CZs4V2ztNG016w4frbuqRFAx0dw72bWU1WQ4wm
bPGRnhI4J5mXGsbdxM8eme0QsGAMd9wDgJepZezXcw1y93iXRSSaYgvmOGxZjQ7uyaInQK5/LlqT
oflHqMlnivMeQP4sv7zy4a1B8MsVsUA4moAdFCuXOT2MCXyPd2omYKTA1OH2IhlD+BwOIzzSFPd8
ktDghktQwYkgMKE5wjcR8KyInwakCG5mdA1AKL0aVV51Johfcd9CNSh0GRc2BRt+CWLvWgCEFs72
nGa+dRCpvLo/r4D2mAGJUUx7T/n18Qr9L2qQ7cWbVSBD2zNxDP3h7CUBUlm7wANyegEdrDTHOXeF
y/2F7SrvVdQ9yiW7XsEAi/JhHNMssoAr+YbvUbdL5LEogA6Z/mkA3J7qq+y7ear92svm73eAOeHX
PSVDIWOoAVUaCONHzIFyFm4VkScetHe81R2qG5etDVo66KmkvHCqHSkQPnAAva1MHhK6bENmikcp
vLlnT23BFcBiz2LPv/8QA9VFRBrVqevy9q+1kn2NtulJX0RfGYkknySMzmkZIVzvbp5cxTFGVI4Z
8sb6+79/ZQiCUql1FL/GgAn3H3lrQUaCVoaLAupGUS7n8mCSOLvgUKfKdCUTbJIQDBDMPjQaNsrb
GA7zBQZVyTurMxD7JKrpr7KKJ0dDX+H5VAFCk0NEUoC3pDFAcmM6ZU3Qh8HZIN31nmrkWi6FLwiN
Ge6wpN7tXeGcPUJVHn9dizEAd4VAwe2vhikSu16eB5voKuDNEV0NRwF1Os7QLUkazhUwF5/6zJzp
aZKU+OsuVhc4/7bEWkTYuJLF1DdSIX+QgaVYWYt0R+z1JAd5OoLkNP6Zvk+SGV7b+8lyamxK8dj9
+/WuXXLtubOyBrJcnenQNyMhFGxPqJeYXQWNeza6tJOG5m3yH5vegB3pGMarhBJNPiQyaZURVDl2
ya2UZBPlhxPvQ7iRbCZSZNo62RTQbKJR1uyowBpLyXzYYsEjfqKPb+cH419/sPcS+hFwASy8rq1M
gFdtV8XczWmjexzFoUmeC6iTkLGEyZBQPNmLFt4KRBqKznNLAphPyqh/kwV8wdhrshNbO1XR6Qy9
eSfxs5I94W+Kinrd+su6MwpfdPLu2gZ3qC9G0pHlFw1d68LsExii0hM+Vh1cOKIQsxLbTBGj8BhY
ySQ03HyQxW7kdWOaQiW7CT2B/SxEqGC57PBRjQ4zH2fkNDtOYVIKx/mpX+8F317UEjeSqwQIaOFm
dmzy0f7hvalWcg17uFSyQf+gVT922tMNag1NRdV2M1iHB0ahVUGUU4muukojjMKxJ7wEdYOx8Cdj
9MFd66zB4GNFUDDbE6hZcNy0OQ0JQ1nxVcd5oe07j8VnHBQUa+bmZ8rEILb4/o/tP0fPhm2bEUWN
taSgpCkxmPddHjj7iI9tEcud/gOaSjZFR1Nld8m31xwHUUWRiVn2V0zefpFnfeOmqK8SYf/2YXLm
z6/mWRTAB3qjxgJWiGEnTMnfEZHB/6dCVFOT2iYNXq2ktdi9B2otXOsfc/ofPLsKEdbGu2gqTq0/
fPz0TfUaIzwTOBJqAc7c2t66fZWWGHu55xujlGUyoovYodyub+91XnmGq6sSWpzBvrRTgm4URRV3
PJZHyzrhBaxWWqSIA7mrEEVilbzZlVdF4F2wkCZyGSaZO1zJKAorL3c/lbQTbBe6n57usPcMiwEa
IGOn84oj+/E8rB1E/IFEXGVDdY6tQF2xhYRKBgohdin9IT1AU8eu7iIhZD4axj4kr4eGPxJpNmLI
Zk2tUXrY0truFWvNKarlUSX7EP6jQZTi5pq6UZKrbAJy3qsxSYe59nJTczNkPVmR9b/Iu9HLLWoJ
xr7Gr6nD+2zQb5ROTDht4LTv13/cIYHaKtPeko71twnuwj4Z0NHLmNHQ+Fn/qBe5HP62V05hZvfQ
RiVi8FFG2vMOR4utnB/2MQj3z5Na8pvTPk5oBu5KP1+wPxdXR1rX269iF3VKF6TQ56VcHoVBJHeT
QvE4oTK9r7LC4jBV8NHmGkIXJfRpf1qyABxaHfQDGZ+xP4XpohyJrv9Tkvp5IB8v/9B4NXvbiesc
MFIHYbWf0Xs74++VPNKo7ibX8Tm00iHpYMr1BVMw+DiF8zpxmWd1t0Vrs5NrsKOmiySFMJ1QGZEG
QifnddvYstMhVMzqJQZdqQwjgo9lxhJbv5WrV/oaUce2jSTY6Jho8fTfDBK+SD28fJIEkNFarUP9
kwdpjCasJLLZhpTX7q0gicl1Xrap6618U5KOZ0rS6MOshFfrdvRJAmPoOw2uQzscVPNAsgifstUL
SRn+4IeHP2dKlRQowLphWmCuZmQg6+oY3t5E2FvthebzZ+AW/0798SoaNhWthEv+JPIPOE+Ol5bu
1oQBHda85yj7paQpKUKTQSdQlsoKDsOGA4aQKlUHztP8HX66594UVsYSB+h3cCGMC/ahst2FEVxw
B6axXwz/ktFUMYB5hhps6uTXPb4DFmY2Z2ePNCYSYYQ8lwDSrmp6FMasZskB5CcbRuwApOacKJK1
TxB6mg+t3OZQwOgwBjXvCiYtZkE3pf3QRte19qE0t446cxYHlhcrOXxJlTZAF+tTHN+Q8NKjWgZl
9fvNNvQq1AVPO/TiYNHOL7rA7YymHtBVGgJHjqxX6i4dsB/FJUxzToWjcpgCqFhSJWmiir2qk0Jv
IAy8yT7kL68LAMo3QEFL1s+4bmY+uUyhygD1rCmu9MUOKKw3wgdrS8zuDTf9ID1wrLvd6/qQ3UIF
166KuQWTECOVezpfq67VwJcYvxFWV5ypVxiCkPpNnrjW1BKK7+ZOb/x0Mi5vlFHCHtzS3uZ75BG0
yq+7iabf0ruA1tiLAg2Pqs0bRDn9g2BarImOhBN66Y6ip283fA5Gp/97IqpqIkaVQJFiHxhylu3V
9bpB1dnVYFshA7AVo7EpaWXgF+mcEiN5sQIhGZUIQgoOGuUy5oRe+G6VhmT2Y1sfCQxrQ32LT4EH
aV6pSZfhXTlR5Cvvx9IMRzdVotRy4DTH77Rq30NwJzu/IQX9qm2TN+myjPVZOT2qRJmlbZV1Ryqz
rFL7Qp2G7RJsPL3RkgCSuLT52yxXvT1GVW518RTcOV7xuiPOuWpZ4PUUNl/eH8u6+uR4nwUE4JRG
cO0AlEWFlhCT3xYGAZ4nCOYbexbRf3CYMMuIpnEU3mOwOMjGuFaOUicdbqqn6t8QOrR+Uz5rOJ6c
SUbEtyA18hpRw1d4sAuBwdiDYsyySLqNFdnUQAfeGbsacLPA2FtE43XxfKGXI9WrhzdFw+rZNVO3
11y+NWbKEOkFuvNmo1ruksUnyAVYcUZuP/Y9sDvNFab8LGSCX6pgafYq/H/8Z/aywXI7uWrpHA+x
FuTfjmL4CS554JLyK73Qb4ZHm0NirRMal5jHifapBBnsfNnnpDpsk0ydNM3dCAsNw0RXyuMDl3JW
xFPokJ25Rt7FkkqkEDCWtlhmfIZGzn52nJylYu0ZXSR3jCcpbHhu2di8GU6YdCsA8BIpszu5MmP/
DKR6YCYT87REivl8muzFCFwl29GVETOcj2lUEb1m8TBMqfrs4ThUHzf0N8cycU0kO1CSkLDg1mAw
OJaL3TQ/0Y4KFpXijrpxYjC2L7Nqm7/jxcnSBq0aYVdHswgi/Eo/ntZZ/lLFRnygLOsaUVWowsuu
LKDnDWCI/okvwU6ukbuUPrS6I5+d10Q97PypZIjjlHHygvJ2jmCFHNZN+X1OtitUJDJNoRJ0UKRO
bqAaIqnP8366Ba7AIN70EqpMzKbY6Pp77VNgjEVHh6oBvrosSx9680uWQL0g58iU9ymJ/033JdZq
+//PupQOM32PLMqL9FqOXn57KDsvG83N8Lj9rSMWJnNPHrQgmneTCK7twjWkZdI9xqeILexMR1u/
FA3m1aJAIGDzzLU9Tfim+eGq55nAb+lPcT4jw65afCx/UIzRMGZVv54+2WabVsX5lzZnpUrVecss
HXJONdX//IdjwoVjxY9+70vWOL3nQ4b9VNyVA+afjW076AvHr11R3pe2/1I8aXFOcf//IC68aqF8
8gJ+C3eCPHauYvGcX2/W+KgUSCktHA5fZ0t6tgIZ3VvbZ2UB2Ukwupnu/y2bj8pUWTETQe+c6srM
CbrpIl3VfA8GvQIr0lwtNV5zuRj84mTF4xO08HUOZdYhIR/zz52NLwx8cnWjo0ie0aICnycoM17P
pYFpdisEgbYCbYDqfngiHqpk+cCnKopOBiCXVVLCU5bcOPyhWECqGRU9eZA4baKW4bYiOyscFy3O
vArF8TAamqM3j09PAPr2Dy+1G9mqXNNDiDARyKwjDXn+vZOoe+D7nNUBr+7wPGBIvugcDCLU2taV
KQ9vX6TGHdSlYlf8E73uRHhubNi04B7B9vhm1YYY38qwXBu5j3+XlTR79B0P+yq076YRQmI0yKpq
TY13nNydtLq/NCIXtn2Dm+dg4mx6XK3zcS539YPwX3nEPeFYgVpjJf5ehEOd/rMGlqYtCYOjxPqI
aOgzlJ35uylYmWH7QknZ5Cm+L50N1WZsyEc3qcKCHj965rTtnNJzjxPlAr7tbaJMaokxDvVes7uB
j0CJdwaVERfPM3yYxx/B6CHkJdnSQ0NRD4KU6UyPvAT/8Sk9wudAt1cu7RKVK6XTMwjqliKg6fBM
B7Zr7+uJFSiepWgoSr3W3Xs8TXPGIKjVycoLqMpUL7zvKhaZ0GnecqaHZmN31o9v+p/izgTDs9dT
6pkU5WxmKPdIPaWkAmtKn+kAmDTq82295VnbKie9KTgdIdMUcyweD8PYHxLTWb85sb6yRBiP8Ynu
ntC3S9UDUbp8KBAVIngp84DWiTTB9WOCsvP50GbwB9MiOI4G/XmZaJnfIJhio7/OuO6nMOAwhncu
RRctP5xMjQcDg/W8Vie98bxwcQYjNVQ8RddzdL9/eMSjlvfKt7GdnlZvVSJfz4EVihNygB6mG9UZ
Cpa3TG0WMYvk2zggLQs7jZmSOl0QN1Isr+Mkj9ASZ6fc4QBaARNXWacFh5/Wwx/SuMOKw9+q7NiA
9ttmc2WC0SIjaReCDpPWn8m6l1LGOZhWNT+KB3GbAn/rhLX1EA/UgfNe66L8GUxPuR+DkKN2TIi0
7qmnjWu8LNaMpCWksqO9rhv2eW1oT2B/4vOOR/c7fgdTYUmORrr1zNLE3QNbcUh/wBsUehdVhhrm
m3BmOd6H9xD0OMf9X5oLKyDdln+Ok/qzR25sMISCCaeCs8vmarMJisrVTbWOf1fNM0PRsnJgBjJV
RvmXNXoEHhAEfPKxB6VvWyDLlf+20mdY8J8NhFtFKzbESKdUBLsDy26ZXS9LdKisC8P/25yLnfoH
W7RJ7UD1NZzA0hCGXCrMZjgXJCNUAC8THofYg9iOLMRNqi3LruTUpHgE54TXiopXvB3+pvF1Qoga
ETrO2oTXPPMAeUOWj2TZUu8BuIIx0OX/h16/7BTU7LRiyqGr06xsO6ok0/gslEfSTxEO0zAVNgee
P7Ml1j+hfbE34t3luoQTSnOMkW9ANTC4gtRDUXRGW2oK7zUlTdzCpYByiJosZo5QM1kIlvZ0vjPG
O21IIqWJzXu+vCJE5RbHYMWPA2YBpVj5MAjO8Vsst7M2v6CHK1PHQkUuCSbEPV5xU+5mRAMQS46J
g4ye17ieZDxCr8J7MuagR6qhsNbsYdesokD+jDwMPUb1WfNlLU+bOoE3zFhp0Xfw0f2mXIzxrAyD
T2B0B3zn9Cd8pVSjHAm0Bydo07J3mp0Ibh0p81mmTWIKdDrzFffWLuOyq5qdROWR4R2CzjWo8lvB
Hg45cHh0KVnES6Fhyyyaes3GRuTYsn3S7bV0RNsYmmxQXpaHxJc7EZohxg5IZuzzDFg3rRLXOO6I
lB3tCpjmePdr64WrUH4e67YvKZBN4+tUFE6tJMU78z3vHVrCeG51vDQ92ID9wnWkNtA/29JYAb1q
wIu6ftSN265+6gYqGR5f3F/exUdV7CYxbY9eJTqF97+lAiThMSWSdkaXsl2MmYhY1dJ0X0Br4kBh
qL/3X573oO+BoPz1rkrajrI1UMGxtypwDf2ft7F2x/H3FOZI6hTzjdfFIEQc8LTlLJZ5I1gqt+qI
MXt6YJmQI17rfUTy6nR8PJ1Hhgvp5wnJcweuOunalZjVPLu1U65YULsHs++0DS0+jJ4JqSGc/VM4
yLWqzN8JTXVJRi+HKS/4h9FkiYGfNji/alQcOSpiFeoM/SuLrT1gpiJsoyRQyuRZEhwC+NPlR+a7
l6pqqYdma5u4c+CNJxfSuGMg60m3ucHYbo8smMr3BYBSAAbcaG2znvtxgVopJG+WMGXmNRwM8TzR
DUmE5hfuvEqeFsTmNZkr/S/Zm50226etprN+J7L+rIpzJS1jJDkm5wZw8aNaemZ8Z9pAngedvncL
pS/5KeBO4WxGPgW/h90cuvuLAzvdBtXl0CgPQ1fLq6Esob06l3jH67M/HN7KndUXxCjXsXPbk/Lk
E+/wSpN1Et7h+bG9KtGKnX2Uvn0QFP8YVB4+Vj1maHlcl+inzREYktZsMetF9fN8cIc5Mvcx089O
LCBdIktmZXWAdXkQMlBLXlG2kBUUz0bmFY0Mt1JkbR9fgYchROq+2Z5TULSkuVFFDzzgW+e5rb/1
7zl70oGPn02Nv3UHik9vnevQmAkNCIP7pKHtty7HrdqjHxYHqSP//2QRmWdX5sNsoOPBPv6rIjJj
LSdd8dpDNrNqRl2JAGtHAiNsB/whszAPQ283r749AoB/4SIU7OnuQ7Tt9CaRC5tg6MOcSVDSNnil
/M9XpglsQAZiNoq94lChZO63+KVrx+kRIkUe6OzwT4d+iCkL5TDBYccM4WY83T4nwm1GklEPep5j
q7flzT7HFTtWAHUbioXqVPprUJc131VjYNSanXc69sTxhSj2Q/4HvjdRToYUcYx4ZF2rQo+PvYU1
1yHzhY3FdQwHJBrznZ/IYBcye3AtHbaNoUANH+aBTTuUqBzwqq4WVNiGhD5rOAAz7YMcb7olLnU/
10nnztyOjxNDJnwCiMrlTmjWdBnLCv12jVWBJXDgZVcYVyeQt74lFnd7mk+dg2vUbxvStrN5QpQG
cuQx/i2BRxqK9q8nYYjP4Bd0zyLW+5cmNK/Oz3Oi1l2IVst8+dbAaF145RPlzPcgK/YJGlvElI+e
RJeGz4Q50ELaCP31A52syr8KQNHA9jDQ7TOwfZEWUW74EzwZtkUvNXcp9emrDdZLbvEhRnGCxsoX
jAqSVr6yw42YQUsKn0x8yPTctNB8CAbO8BO5+FkGjeR5MuUSeo5RiG+eUzpJI/8Z4NO+tIGaKBin
U6Zj84UiiNzbUnlZf7RWb2siVbWAAG79ZwQumLq+dqAm0PztvQWlrIMe3tBEddxwOq0fqi2XMO68
wqH892M/FbGMZVDDxcsW1ztfkeScUU1ndsomhUqHOiKNecilD9L8JhnEmQ4nDiFwuz/Ei66BSCdC
1mUfnBuRRxPgHX0SscULbhgi9z3HxmpfRJfADJ31DqcCMInWlEW49+ToK/14jUvwuQMdSlA2P5oT
2bfPX85dy1RpP9SjvvtTlM6xaH/Strqc8cVRZ/z/GK4WtOakTgcvw/Tc34nU1FrKj5IkVhCjpWO4
84TtMUWFl57+5jvtp19/5sI/3WoXeMx+DtXBsMu1Dspp/Ze6iUgbWMfpYNVRik31G4m7XW5ApssJ
EHCpWAyprQ1XliAQ7wjI6qNK+mxJCbnT/TTsA7rGJ9GcWI6TDQG9UlRvxHVWo6nGTuU88wdY/Mnz
SNSuCAtEVaYpEBIhZt6efdhFtzzZNcg9Xlc9cYMzpQu2Omq1Hq9h2rp8sVSjXrOTxQ3KEYvkcyNM
hmjkqxWfwgACaGvwpukvQRlj7Dxrww8eY5VrSFFU/eChDjItjuxDjWspmdna7C3JZBMMTmBeZegI
xyfItm7Hn4x04rxjMS5axVjyUASRPq6lxn5ud+7Pm3Tif+1jZT1ZpeMqlsDhnkg91cPXQBtTND/8
ZTah0kj8S7PSmYz+t7MY1V76rc2ente3COzdVGvhgkorgkYyBahrSaVM9WQbCFuX4cAC40DXp4pg
xpKGPjSImsr9tW1P3rsveccDPBEGudPnD7qa2rIgxH040SrOeTtp5zW8MdnfgJ92duRYBkBTBTNi
6kO9bxbCnwZakOKipX9TYhfut/5Rhade3b0hk92HhrFddQxcZSdoENwoWaBxGx02pOB2INjnS1rI
HPg4QGsJnsF/epnbCtSDQBpu8lgVhsHDFOpLPyOWvmaNWF2KTK+AwcDLg3FujckZwg2zkRBDU22I
DZvBueHsiIrqIEtXiEaSUAGtZ3m0oFesTJUvUHG+Km142hHX4YZrl3xml4ktTQyaaitji+IdjkIE
y4MTU+GRqfyom1np1pGMMi8HZkqc5Mr3GUJIx/NmHby/ts16nhAzODwu2CFvlElzfm9CJmM46mqI
m3YI841YfuoN+YzVqzugchFHwaYG5aBwLJvubREYSOm+MCC2rN+xci7o47O8FcMw9q6xB4mBt38f
x5VC1kuqe3SOyNodElVQQOnSsDDSX0SWcU3vKzMis4b5DugrH8Yix8BbK7g40OIJexKYF/AA6mdZ
fl7AZZolUCxGRTMqAAlwQkh8M94dj2zPgSoO5unzgUMf4mc+QlZGeR18SM02qrmWZ3funrYHMoyy
nU03blcd+LlR1eR4Vuwh0TY9LsoSG0OBochngRw8zAkvfnKcCM9n+BNAP6q38vl9OLgXbmdj6sK8
1pu+V58wV1ULJMc8xBkqhHHza4KPl4oQqcAmZGU4r/G9R8Dk48lWXDNBKHHuauh7EcREXfcL2YrL
QJuk5+2S9jBc+eTW1sI4t/UP6UXpV8C80zuwYUaeT6CkBpXXYtD8zqMUJVMpokuwlRuFSgj/HPUO
vVDSqAWlYUircyb7inGxgT9m3hW/X1bD6NJfmyEerJZ4d5Ep4okJwTvDdte4/KXvcAypDbA8ioo6
hzt12FaNK44wSue/KY0RBGlc4/KLGKR2QE53kE3+ap6gAomTzAa85GnzwfLLTmo4kkpnv8EDuVJA
mSyPhEOFt9OtHzM6DoDtUdp1UR0WZ5kX6Xuj2gMbKrAhDjmWF8c3ks/pSwbCKnWfY+ejbO/rG8zw
fnL4TBr1JSqx2gfQUZkteyaBZeWXxQIA3+HlMeVUZfwQ70QjwoUDS0Kvtaq9vuYuoOjJJOy/XjqI
+JjYS9hKFC9MN0iyHcUec+bNsUz/5sQiVtZShnyKEHyJSw2NLJ1KOywSp2ALfJDKCsQqnX/5Ttt/
SAziMeBUTra4c+2T9epxf0+i/5tjvmEQkLhC8vA/Oqd7zwT5M1PLgmJJ78OoLPXb+SYr1hMpAYAo
NjZAX+Cxj1/4veByTnNHVKztpKRxWTN7RR6VdMs7p2SMxdFNnWapskzLZjLxSunDE25LHxTfJYCF
E9K9+adS4rzZeIBEXw1pKMdImKzYukf86wpYg/RM75tHmh/2N5eC3c1oR8kb2LifN1E8PkC6aNu4
ChhHoSwIG0adZr8iOZ+7F1Kij34YtHVhOPHSiHemBQiya56vbGesLk9TB94FuCzSOfB92+5ybEN7
Y3Xsbvl6VhcqlgLxtLecWQ054VYG2vu+dl0XXcvqEljlH061L4SrmbvMJZgQY2FcRZSBNDKjcNJu
GzST/AXjfRzdmC2n6juBhVg8cdK8syR57uhT3+tVrtqGCkICyuBkv/jFcPpkhVW1LfonjRXioh+A
kaYOudBHWOW+qZFYaSp/OkstN4emtjsXQl8aEymka5iwuSmMYcKOG4jVDyMkwK4+4kaMxLwMSIg8
+SLoQUc4eaozp3nh0Tf0eZAzlIfJGtd1g0vxC7fBbHvtGI7kQpILwa4C0qyjrTW+GPXiFOUhHjMX
sTsTIG5EqXYw7l4UcBONS4qw+ouyeUEngoD80DMm4oDN058g2O2igyjAyJ8s5U0eQcpW9Jae4wm6
XpoGVVXzZJhLit7Ve2HH+L+GgZIX+t8P7IoyrfqKUYLXOEDBP9Mf1XnIDhLPXpGNGwcQ8/a0OgKf
4z+JpYtLjHKbUUZYbu3phOt6JbRW3vDxuXnxILZ3sAoGmKdwnueFTc+YjILPMKYFrYBZpiDVAiyv
Hleh0VzcX6BX8ftoTqnA4wOVqzjrSBb2vJwdvrjqyIwcjwM0tMdus4R6FZdUfVqEp7F6nTRMe/l9
R0NlRHHdhqenud4WhzCqtFmZxKtrHoRhjDNxmbvOf27GpHotXkhCFJyUpFXLRU3FBwyVAflTsQRt
Rv32R2aOA8Mn9QPYby0UmMGa3NSljW1UhYqyWOMxfWl5i5B7hZms7NGst5RQ7NhFzZV1V0KjiHKk
bnh7pKD+WZixXz0K5rpK04N6aVIjPXbLCq+L51rzyTpdYRpWtZ/ZwDm2qmC/e+1MA37cQTje4aYZ
orfpr4xnPc+rKK4iin+6itd+0PS4/rFZgW1YL8dq+i6OG8D7RF+4KwZrvsQFySkRRIvHEjT96m5t
+sT97mk+iRx5NQYA3yhf477CHMUM0ML5gof3K6/B4a7icv6K7TZAptT+eIboa/32WG7E87GnOFkd
c3TgY3uPG+Cxuha7pxzRb31p3KDfUxZTW3bjBxQGiRPwCs1Kr60YIcJm2qrIqWme0rxNMkofQSDv
n6bMibBwiZzPFPVMuJBxQr034qaUuD4Wb/RFzSC84f8WZa2UADTsiNAnduW+HKSPtkQkzXudWfgE
/5797VgjoUBEPzDnz+Cx6102BkGDQQCcx14s7jm6qnVwqWmaDVgr815jLfDSWe5cVM+xkg/5FF2U
cigEZps+CLmoQY3YVXQoE2KZmTKlFEQAUQfHqmjwlDN3MobH8mkL5ZoPaQDMhWS8fp21NU3jLT0u
ac8DJUsN5rEGmQpPFKOGGdlMlWEvvf1IPstKWsYY1xRw60cEuFRhN5GGQ97oyFdegImiLVzB9boA
N+Bjp72pj+l6/LnP0+VuhOvhjj3hk3PRvw9hDP6rOPEAripytIwDk8pmlj0m7/c5OgoFBOY9jh62
HOwbwaK4JISz/2hupflEr7YFcZ9QE7zXNWZ5VODBfflrTp9lnohRyixQRRdQdMPhk4v/qAARxDdV
TdD8DyTDTxFnLGBB1OZdjT8G/dnBLk7EXTs1qDR3ECJDxHWZdfZFW3hfUvCHHTTqX8AUwpmGSkl1
F8OmNXBqjQ9xiXS0YQazntlwdbDYmw/XTkO5//iiHpLUyks863Wp0pn9KRm+V/T6Ps0IYAE1V2zs
b485Ltf0lWlY1EDnaEyvHc9nr2jsbqzNiZXlOxer06yz6R1OcbjBJISfdZlXJMwv7gLfHxQiq1FA
UdIFsVIRNDMQXZm1xo//0eyBa90ymD8DkY6Vwjxi33MVHN2CGHqhbt/oHm9HrlrgdndPNsXPP+Cw
UaBtHsis7ZHhBweQeeR3fJfNuRS0j0eere1dfjefe4LbE8zAm8nABXxRE7qGnbrwPrggcphPGywL
1oHu/JxqOwyHQmXCWJIQMjdeK7vjGarVQYcjhu51NInQxTJ3BCMjIs390ZWTj4I4DtTU/1Fso4T7
s8tmEXtz6NjzhR347LIgoP1hHEwqNnPoiDarwz6IraO/z1+nHbgZquHJRtwrYPtTDLawTHHlM0u4
7L0mYz79aCSFFbXP9dWJ15F41qJBhouBRyOrAfh6ep6xpQxtPm9O6m/brpJlkj4U9OBhOcyETTbK
ucA16AZJw/RhgKAULG9TK+djEeU0cabrY1rQ2yn+YXc46Xx5G3kLn9QqPaoMvB3jBTbC6eBo4VJe
l+rLOJLw1Gc7h8aTMqAKh8n5UlwzWvj9qjazQ1DDFlZRC4+X1YqUEetQ7a8/zl1cP3KzhYNhggNM
M51WgYw00ly8WjHfZ3tNPMebLC01d9RIGhXN6gorwGfaXIyen7EZzh6mXc+d7ZuiZIZ/FeNm5xh4
xYbCytHCk1vM1R4qFdxPqkfaZ8VJzRMIBkZvECcHdrWPTZenh7C29EV7QKgaQWzo/UqxPjNxZiUG
l4gQCrM7Qmy32obdSPdDV5flBuxJJepX+X0AQslK9vvUydYUsv0D9aFKUWUcVnTcLEDIMWmI6YxG
9xNcxDXVZHkQRSaiOWGC3LJHGDprbccLgjBRtQT6XJGBm7ov1SFuH4rIx6Q9fP73jcO36K02IoNt
YvqUFPfWPY0Y7M5JD4tw0G+QGLf9lksciWH2I6adJcQ+W1zDvtLiTYeTPAyUwZL0XTNXMliurOAc
ePrSmd5N/+zkfvI9W6XBpwywsBIKiqNNJ4aYrap84XClhqNOLURGgGI2y9Nf57cnKfk+xSQtNwDg
vgm98i+ikw01RMByCsfTKfXigSmI6t+/p46DHkDnUSw8Gzwdn/yif1mQXiaOIdyzSWEy2EU5OdRV
nWjVT0ASO1Ii8mx0+Zk2gavS1N7JaM3odwpQdlS0wGTudrQ/kihjnWTIjWJedYL8mKF9a1Ij7F36
phukdQlVHVO53hlasoihaEs6p5T5lPcz7RC/6lfNX/k9AiGf/R7mk0wJktvoGIC0o3gKZ8c8z5hJ
EnM5u3QDu+eoa/vbKCsGUWGE+uKkOx7O95Wv/NCTdkaRyxpKUp3Lp6v3Pm5PYx/p+r3oNIHZ3Faq
IGT3832S/ZzR2aA+X2ia4Q+ZA8Xu5YmpmA2lH4JfXt1NfntwD0LEazUDNsCh6uq6hMAg0p1hMIsj
qCmruuomQ7vNkYc4gjzxbUBvxXGR/108qy8Vx4dmnV7Yaq6X97be9cQW6UIsSIhLFxBqwoALbbpm
u3QfFg8r1qApL7DFscDkQTp8ldIxxOSAQheaMQGIeJgrv3M2wlpsbbccs7gw98DmF65O61p1JUOb
SoACV37p7n1AvPKAaqH2Z5r1lOFmqFGH8FFqMpo8h7QAfGughML6E5wVRWlsmX2o4VtjkXRvKYgO
oFycfAeAbjiszxJoBq2ohB5C+eat8GfbsS3KXgxadbgaf3dyAUAZ+DsVxnB+xOAbbBVAUO/oJsPS
FnEDP0FwK81ntYyVnd4HPW6q4CpjvM2rR+UjH4zpyE1QhaD4+p/W/G1na9uqiul8lgLAUf5GDn1P
AX5Z277Gbnps12D2D9wNAQ05/TYrd6NXigNFKemX+0Uthxq+Pa52vObfRbZTIjq8Ptk58upZBgYi
isHIhwN7DQSErefV9FAUzfvinaYiS2SIHLIoZ7U9nmyLZzCuTG1hMSzzY86e754gD0JXhPbLB/OR
QWmEf3G9Z7WB/1hOirF5UMbMAC9ol6ZfWa6tOtc1vHTEwgstTTp41iyuzeLjk19qr2xN7lHCBgMS
KeTkRTFWu0Q9D/78JjiSqCrBM84w37kOZNQuAPAoW2iuk/aWNe3te+eXa4pNXoXE/duCjjrWfGuE
I/QdDKacPa0m9AYMm3zhGCemErPCP+8EtlgVf3tOmfvZBxu/gtfMuMsexwlTD1uztQRaqGQ7dvHb
Rqi7QhAxQQYXSviX/6iT362afFZEO88tZ9ODZgqopikFhIYMCjJoQ1bCpPK4RR6iPDI5SEsqjqio
L1LsaHu6G/e0s6T7gfSac87xYY2ak8FWQeXcElYn0dcYVdgXCgTfcZgP8mhAiEmBvy1FZz+Iiw3M
m+NYK8TKMqLF1hxS0vZkxHFNg3Al/SVSmjCy7dvW9bGDSTMn6YToSP2GK4A7DeFMlXQv/evboB9y
dcsy+fxRk7RCfd14og1xt/Psz2OpPbAvNxsD8SY1Fae2fbe0RjMQatC2PBe89+Vsd3T6ipRZ9K35
yF8mGccSYEaQuXTmIpolUS5BikGIVEuwMhcOj/hhvAAVomLU+GpOrx/za3OOz6e0S9Wgqh7CQI+o
XtaTtdgWt6NQDtWMso0/Kfr5UuBWNL05itpLWexaUSvRG4eD7K4wlzYMwQX9cAlisiC11KvZWQ88
XMeRGtwuzyM4fc4poVnxc9zqGnlzJ4sdh/w/ow+/0pcaykmxrRfVM5q6+55RgJAXZwNWvfmphlV6
lvGP7a291pyPlt68ScyO8vlxo4zfuCl08DPCIt3OdbFlsCbd/aeBBILcQzyDZR9028OfZIzsvGmF
oDKR5iT6Ve2dMgR9B4YmAkiHbQJ5IYrkuuNsE/RxeIg16RY0e/6g1ks7DKlL5rO49OA9xmQ6+173
Bb6OmlQ2s62001RlwHIx14tO8MUyXrgs4XcqF5bKFIZGDK08df60G5J2BNHqN1GDqDMxcjympvDX
RLgeo7VP4ZPZGfy8Mp7mBqIWlWMtpmvWsJpMCJWnbkUN2q2yvYwiW/yibo0LeTKueuyCpP1aBWZe
//sswj5be5VJy333gdLVZ1jl6Pvfejlu43Gv4D7XwvilXQP4cTj4EHIgmJOzi0O66Qwxx4Jk3A3x
lkvVuCXEZvGheXpChh3frhih//SEmB7sYNJZCJOmK4MoHf7KVxSX2HlHZC3/UZjCgX7IVJxxMeX1
sjSrLuEOIxFXa2OQdPHZBEvxHV07v6wmW0BkCkdAAgSoSg+nDFgHd5P9gSYSSE31OFrex+MaRxL1
JfTfPMyajKGRFSt/67JLiQYVtXGSEFzoc137Wk9HOmg0iJsJXZKKIRfJ3lrCiDIJbKzN0m04dZzJ
nVJ8NxK+3bAdr8TwS2YcG56HLSbUsEq9vdEyMEJCZoIPlZ6+iMrQT4zA7RYGhL4saDIVf9EQjsvr
NcAsLNzGe+NnikhbSrw0ypru/3drG4N9JYtnxOi9ZAEHhRYMVFtvu4B0PI2Vn44ONsmBviNwQWMA
8593ImjwxGRYOf+6Fr+CWrEQ5sRUOhDixtN4PnuXmPXWwSZfX3rGLsfaxU6M8hVMOwn5giG3mZU9
dHFtNwgFsznW6z5WaGLza25T9yUjRX/1toJnsrSQ2TW4np3Gm2pHlkTvP0U0Z/NMKDGsgrtcFxg/
0ic0XxTbAUI1kmRDPMwKpDhx42jna39/N/AjWbqzaetxazJqYdW2NaqTYuM3pI7zzS0cxBOldfdE
R/tq9vA2fF6q4z49DTrsfZxP8NJh1NgC52d+qG0LB8B1KLrK9hP06aaJ1tUt/4meciLlH5irJrl6
4JGGU+QAU0bI0vXYBIKd6/FAPGKorEuajGR0LZl+3RnXnIwaUKZxx8fXvnuprU1LYu3YMDd3iD5L
+pW1lZJWGlsrRC2f+wQpG93+lTMKtwxvedXGsz6GKZ7i6i1XTtSWEopV/iwTb+XMD4F5MCfBI1++
B5IL7wmX9OVusGq6ba1SnoOMvtvO68Ly3f3qVN479kI5Wz8XblmZ+8E81nlP0X5gHXGRv7F6Ad5V
EVJmmgovDgpD5/WvvXN4rRdFrBr/wFLKsPcbwI+EcfaXVNYIwIsY1BBJnD5KCYaAooYVKv1rMcYL
/aFAW5JvjzFv3uyfQWsnFWf6LfBTOZM9RMIQjdbDezJsDbl5Q/bxsHB6+nJ9H98Aa3nmWAPd8qQT
7XUh8k9Je3rPNkG9+6/Cb1fHpOCg4PczmE3i+4UlJeJni95gfxIyy4jSxuwJ/enpT3k2YQrJuWgK
rfUWmgdHXJ4MZIlNkMjLP46sI1RtI/FqmOXjINgxsbGt95KE2fDdKCNjtZI/eeqL0xqissLSfpaf
SNluJW7UTuPSO/5O2Q5GDl7lI/KAswd76ar60HvQCugcQN8xwi0ts06nM6wk2sllOSoONZhXNaAn
Pzk5dFeXlbSXAr2LjWe75TTKeCTfoufGp/FMb8qHF+D6xkrfcx2K0eci5sygIvRBK5ACrggleNKf
2MXsDNMwDE6iihZDEj7hSBxBAZowYZk43qiBXQtQniAyXfjjuw0+xWJbDnTSTsF1poEMIeEpPiE0
8DsV7yEO/wxyauadRN7a6CSHQ40w3jic+gFQe09lo4T47TYjWCBocWdyb3HRLx3QLSrD7qk8WltH
380CUKZD2E38CjN9D4Tn+DE88E4dZkV8J+7VpqY4jFuabZov53siVCz1TaIRbuX/zcaYeZAGbLj4
aVQ3Zp0553wx6JEwJ+lskoRqQkDQCOPKaJxKx1stxMQ2VjMPjBs03P90OmpMka5uPxlln+vmNB9K
Tvres8ufuP0TmfFymSCio6rKJ567h3oqxwF02JRLaZ8V6ID6MRhcki3JB3I0attGqfsPsI4wwRS/
AIS5NdKwKeJkHrYVhS0Ylxpn/r8e6mZSbd1C8AKUQDVtQc2KN+ROgfqHAUfDy1yhCsoL6gC37skp
NTxVYF4qZiM+KabMb8UKioOmqd+K/5jjcsC0XwRvOgVGfZ5/XXrtAiz/YjhDkSdC+RnApBB+BEhr
Qp/G3fSipYI1exGpqFi5p4i4F8dkQzpFA4X0Z20Gwequr3zBohry6W+NXr5Xa7mrRavIWl4rJSIN
xoUmAkGf5WEYYZ8vCUY0CAqU7UNXEM+KC1oDfpRiltvcRrHeTazV4C4M+MklfR/Us8+F4FVb89qe
VaZdJ9cs+KNXk4boh7yxOwxJZ4bBB1O55gRr+8hyLjbU9opKpjbdt9WVRT7aqQw2LRxg2BvpZdgG
odeCDIu0M03HL6tRG3EsqcZrQJLwIldamq3EJMUAKYBoYQewEBLZnkArahfCGds0HvnQbrntKMu/
AJKcsM4dAcn6bwbsZ1bz8/2t3BkG/Emy5q28p0icloYCaCvyU4cRhGX3UPRCVo7FB8UIaQOTH8FO
DM9Km2vLKKh4iowi6jCHYFHu84DfmD3VjO39C0+pQyiEje+SytZNksDgtZj+2wEwi4Kxn2AEMF2i
oStKoh4y33Hs0GGSEDA+6ugg7nNiUfDImZm+qYwFEuA62Iox90a+RxAeeHPNGnRr2bE8BZr9nHpK
zPmEtahOAya6+uqqQcyDWkxSoZ/IKtiNE+h6Ff5l2ryWi8ttsPTQkGmLrzbJG3pXPttAiysL5w8J
RHDsliGtz9KZzVfRgdAs16g0zLkJfQ3wyJkYpp2Pw1w9KHWRK12ilYA8jMeZYN079PSsbYHDUNjV
Cv5hWkOc76Y6aFQtge75JXooz9XAhxEpmeZmbzScZoAFixWbCOinWUnGA73WOrvS9/Rn8QlIzDIC
191E0jV5hFynl2wG1k5efgkDj3N1WmJeimF4uxaFitjvGN3z8HYwS3sduX47P2K/igpFtMcmPgeg
6n6w4ZRbq27n6tdv67HH68XMW/4/pB6Tz3B0NOxD7M5PrjK7ZIER19SGx7POoGFKxoUjmg1WaXJh
EzldKka411OG0UgW3iLvDARvlld8F5LuKh7/AZ661ZnwVCRQyku2GODwnmlkOcmW5bV8Nos8BeSe
FpSjoxr1I87dEH8d/9R7W3EwsJNJiwaFfB+y9Z+Gglj7F0Ps2SuGmcZXed3l3mOA1I94LDe6wdIK
tn42T6SkyqofP0CPiIBtTKeyFwT2ibq7cCe25pNd1w0gu00un0al3+dF8/oRHeBWeKsqt6q4paG7
qvGtCRh34MY6VLm194ERc1oyQJbb4KLrdKdjpLViTp1JJ9sfImEmyXZ4aIu9AgbxuHOSbSC3tvcj
YG53t3lEqfM7K+eW1wsKVCERusqNMXna2Q9u8GMyVkNDC0TZsY/AIgflNisdqh8VelQmlta5nBy6
F54q3Qfu42jJ7kOpLRjJ9JQtiuNbHr/HNTZ3FKk6kX1vpQraZ9aYhvaTreAWOgbGKRsE4xhPuaIH
pos7MYy3qMjK6v0oWzD4HgYSX/6QSTVRNRDUSi5N2fuJ2aocy/6CCBvmfM2HGgSwwrDUP03BrgsM
v3ATUAwrsRq1pwV3Ufj+XdokVaOjSJQ+GTpvsnkWuR51o4abVhLox/yGlx/SDGFeFgwTjE3lZQug
IxHRkKYO1g7YjecSvJal/dONCJ9uNqD8dwcDWC9EqhGXcn9iAFpmaEdv2JkebecwDN0hRmWOrUHA
QVKCuaB2LNrgXRPpkU7wCOa/QGAJy5h1W+4dwbl1jkBzBqP70R93F8y/+qngrh5fbAJbbz+o6gBV
B9+aTyyVuWS7fWT5D/aSh5k3hLtKYI5m67UXDpfiq9sI0YmDRBJ1QogJ7uvG4kNI8rbcvL12NHeA
cR/zEw4FMY/dF5EXRi4mYVeEcXzySdmXEujN77id+LP/ECLaRwJ7u8biNTwNyNtOevBxYHmDQK9E
dhm1V+ErksoyZLMI8B0x/ZIIQ38QiDKDMLRCnEvwTFzy+RCv7nVef/gESIcH9IvdsKnXWvcTfaWV
aO8k+ndL/SKW6mcs47wWQ4vnq2zOBxeK5LWyylPYTr5OX6G+mkrzcKImP4KZUvIZkfKk3Z5zxJU9
sDXwtMU0S+/Fro7jV5fscyf1Gh0JCNzNofDU7kRX4g6qpHxoC0vzs27bxf8YesZEBjF47IUa3AFc
FMHi6Od9yPWOcSmTjCXVkQIHcjrCLQTzlHcUdqv3aMrYcXNJvvWG21gPEr3z+slZA6by0KytaCL8
hwySBLnT2+Ea/rwtOvK/Gstixn27gbRO2NNDPh0cJVzeK5DoCFKaYjz8SfVMCVe2n1xtDSJJjnzg
VfKSb5maLS7t7clUIcwwVvg0l0O5Qo4lebt/zVe6/4eiZlNvHi7Ur8ayQ4J58z/vbeRtXvccSMmW
bodjhalm8EwJJbvC3tSduhNWd+2OixPoB7sVLtCDHWEom6bUR93lPDWHAY8eAVEZwH0nIp5VNVjb
2snmwngoJY/xVVD/dlsq/aKdMtizOJWqPLKA511aN0CN0/LhiK+2x/mDmSTAmjX/p8LXW9GRJI5h
5NR1tnfhLsDXgUE8bmUOeyrxa3bG258nNUfXg2z49DUfLyU6I0Rdl/ae5ks6hzVrBZFrGrfWe/QT
Puje28vkq9Bcn/2/ZobdRPZAwpuLAX6pzrxD8saEvCskVmFJshKS+GRMoLj14H6qE1x+JC5UskVh
OYkTQ04TEMoqBUAGZ/Q0LURRV6QvaK9XerRsvEz5JGx9ypiTe4DA6IERaDbb5HZM3CvV1cR/krgj
b1vBlDYRwV1UmW5bCFdMHrkOzpNCGDK5t+CfMOp7I+J/TNSX7IpvQjpHZtzjd3ygqL3uAbomk6q8
QIsI7IhW/L0fOwFUFLO8FnlUC/OrT1eVHiSTAyNlzEOLpSmj2+1g0/GX1faSxUWADyNqfyHBSDFz
5pVZPEwvOaJppqJaZ/wkHd3rmct4RCrWY7ksab2famckYhffzPc56pVlHIunxQgPqNEGPKBj+ZWT
ClwsNaN3TpX1KpHghn6qufyxXadzsUyO8AotuzPJZE/rIb7LRg+XthH2F9nYImboAPPM5uQyWVV2
GCE0CcjJatkMuKpEFr5Dz9gaPDWALqQMoOci9XjeZdZPLrZi/NXG7j1Q7Dv8++kckfsqwNLvkaJx
u2R5hLfILD8mL1qQnUr8uWRKjm6tkBq8Ck8tEOoBjlbfEcENlVHkphQB4F9uqKfEBghFeUySo4Z1
3I6lSCDB8jIrvLGy05BD1/TzDLUd3MXgrAJM+e0d04CVIQzs2PvfFS4W1u+KMboOV2dgimFSO763
9PSc4u6c28+9ih889qcb36lZswtk5zJ/y3J/kJ+0Ca96mB1BFdakg081Z3bvzhrOo6tCq71e2tPK
4IZAJqZ+LkWvyz05veOs2o2YLP4adzin8EOZW0jzJ+xgMe/RS7EvbsyiNL7Ud5aGuAUiDLZUanIk
I3Sh1CsPw76qJKxOeUee244QhUrXqjSnFJtifFFL6PjaQjhYgGSa06dbXmOhEIgkXYdztWzIkhcV
f/xL0iwDj0Dp61UuT11x5vl8eVuaVtiJ4P+Mp/NiaN+19oWXleM6DtRarbKswneLtQkFSy7gBGC6
KMbLEk3FwWKTy1o8QRf3LtcSsclOOAW8y/R/jDm4Rwk0XjyuSMv5/b8tdfOyxPWwto0AE3jxiYqF
ps0sfiANK4EY9quZ56Bcgdnh59RPsquRZTjGGCFF4OiYA5jb0H8kxMXBKjqyynVBz3rjgX7S3eue
2LLcXsq9YFQXVV/fzT+L0fE9c8yi1RzZR3ssvtkkmHuDLrnxqeePX1phg7kxmiMRMxvlOJDpd0u2
VV8AZ4/cTE5SXc9/9DJsK1bTc5Ov5h0IMNQw9qXePVmDvSca8DmW8uR5C+8i6CdgJcVvt27EUuh2
cMNmKkogHLUWZ8+OISw4GPuAchiuirI/JyptuxF+SoImrQHAi8fApHBn+EsKu39OyefOu/f7TAwu
hRVOsNJdh/LKfaDlGYKzzmrJGg0JUQZUSQfgjRm2qCN/T47/OiWiGaLGHVeYQsSL5B4c0UuqRVh3
6r61FAjLc0MzrhVM7+9SZ0+H6kg9yNXHhPrxZum0J9Neucv+NI8EPzdi3fdaznc9FlmC5cdo/qH9
zkDub3CqsMMOx8NC3IGWdPgy31Ny71lAUyOUHVA47duvjOuDkU1vCqCd9dSrAA/h8rL5ayEs9I78
CBPl3couLhJnA1H87UYnM0gjzvkpV9YYvKMdjXUsYo+o199uS28ug/cYPRD8ktjPnfIBzEjXOhcf
d623EpX+Lf+Fz4vHKdeEjd0X1aBuXvh3bzAbX0BmzH4sWSkVD5dwoM9XkCkU0ZgLtaBEqclGul2s
k523d8E5fDNufFnFFD84kA2RWCsbR0f+do1Ja0UDx9nNOAoRxKEfqXppXSwkoJ7BNo+Aj/jBTiNX
XP1rcd0bmpn6aeewTOae61Z+k9WceZX49ABoZiG11fO3gVFaokDP5GeIl0CTeAdJ4xsxsiJkS3ED
j4sUuOXPenH679qWiZW8kYTuV115JeOeJV3/kwHMXPultGlvLpifkDt2iwMQBWtxZI15ovHC92fb
rJfT2wAXYG4mxIV4CS36HB01v2psTave8vzAIONDwAzz1BGPxES8+n91cOC25n1BLN1Z/Y24nwu+
U6qGs++YayAKWMxNcWRTSa2YM8vkPXKZ3Q9L3KgTtxH1Gll84C2RzFtJnqSmA4fTrbppx/5FrgDs
557YIthwQNNLyTm9An6Wb+nij77kFFAZcsMba8MyewiVqd7gs7+FEJLFzU9ULv0ipbE+p97TruNM
ao1/TQZG1Xy7GdaViJwNHIp5HG44i8m1e1sdkdVURoZdqht/+XajU4w7+77vuFlhX1XZcRryPrWN
4fPjq8699HnHACtOcxWjlnKK7j7f4nBPoYGnbCNxd0XbpuUJFm5QD9SDzwUJW+FWVrS/ksEriRAs
wkJguctAXgREfK1lL4bZgFU4IaTqYlPx9V5ccAEf77MMZhRu2VvnBALuRKlG3ttpFi1PqHM7q51a
YIuUhI0h7S91QHOj/fF6zSZAywZL2w5OvoGAuwEMLfuKv8cMTFT0ZB+0YtV9qXvsBmQAQTroBW6N
TVesmwzR2FwfmQqrDkJMj+3juZr9Iw2hAppecGu0VvN8OHSm9U31ky+nJRH/jAuv37/C84zi7T6U
1hWxad3pz5cmC/yCZmoZr5xxHtfLyeOi6+U8b2CGQRrA7yrs0sG5ULFW64DxydzBZxDlExmBQP7k
Cyzo02aCJmPtaf9GerIdg9yqQDka/y6+K7bEutIFtTXgu8fII9G9k91RPH4cL08uUwx1XCG2XRyC
MW5b90EVtrvuxon8Rc48/BquwiMwbn1jciuLjTxMeSBxzfBMd1JPohslQMOKn3CAaBftJRST6dTy
KAt/BSsoexToAiLLFO/mHjQ5NU03+OLTmf3v1SJWRjJCK4MaSCHlF/nrkLXraTfSVe64MsJweFfE
A7zbNiWuhQkfCZOB3a3ngZlXqXnrJEIUvq2YZ9ypq6dY8lBbgiQu5LhGBFu33eC0u9gJideNFIg/
0coyvSQZOO5QXNRriksq3C09mgyrqOtwcY63bY/C3eGFj8lrnriiWyW1JcOQCHTVvp7KygCgwhyg
XkjcQ6zzTrIjQ5eHP2eozA1MRw9eP+Fsv96SQvFCHdxqewZRG7XKLhvSO7vxadjCXsXZ50JYE2Sr
b5CPYuWwS1KZi6OqxOeadIqOBBhpYj64kQaq91EErl2drIJZnHEBPDH5Tg5A3ck0m8eFpOWpl3JW
YFjR1TeomyPWaFezMOPqboDPM6b2p34rGdb9uDJqkrp4gbg+qnnlha0Pz/5lNIzanC2nKrvOEKV/
HkEpg9y0TklPLyBKvRCQjrnRbCmXMrpaQrOjs3J74L4+NGGbsl6EfAOE62hc6Ps2WR1ixL1ZDQIT
LvwwSoT4MWtPTmyKKyNYvOm9+qOx/JNBcFQLWNqJxXzbHEnxCOZ8ptH/M/wCyQJ5MPvC8QHX8BZV
kdzyYkPNoi0Nt5sQWeIt+1To9+NkYM3DxP3dcezkdhBfA9h0T8GEaYuNETWFrUbSQ2Dl2FoQ6V5s
7paR98hMm34neq84UgFSv+CrbSBkzu+ra3ifqMII/T0JB/yo+Kk5waZdViSwXa8RgbEYlEZAX2wB
0AC0uwsOBydGUCCy+XQyuGUNaQTaiSXRxl5Zkft9P4//Va6SiCzvc9p+tJai2fTash4Gt+SBl1St
tuKHBLlfkLvy/c85OJT/LaKFX4MPNb/ICqtUiKse8KYJ0NNS5LzRsnXIUviM3rlBHk0c8U+ss+Up
T7kb+XQaLe3KH0wvTc9YIvfjVb5y8cBIcCnoIhsOaLsH5rP09rTGTx4MLoGwyQEm83NEDhV6EHVp
kZKfr1rN/+lfA70QDtp1wqoff+uA4XsvOWZenbr1Faxtfcwg1zybkfd+JXZWSkG6Olw2JL7LPbDj
52whngoYleW6lOH1ahCXd/T/pfRtwbgVNX2ZtBcdaPxdFF4EG/LIqdSYTuNrE9sILEAcS3UUQdZx
KXSfiZ/jUL14bYZHcL8CskjX+ECfZVWVPNq8oUdj/2C0kOtYRSb7Q7odKbvQ7jCuggpTMlwq08Zd
L2vIVeYwCaMLS+a+utdFkMe6jmovVRs0axEOEErp5d67hdSJ0bTdRhb/0OaE01uH3WxR2tyLmCiX
uzzr1l55SCzJ3vwzKGBoNVjIa8ieddUi6M8bthGGhDzzqwXf78f5ECbpWYukMJw0Uu2oP6g/0l/5
fc/geFqJl3miSWxlX6WydPx9JGOuV3qaRpAqIy31bc2j8qbAgE+xrm7+XcToENy8VQfiKGppnP7Z
IWXFRyDegJDnL40RovPWoV8S/WlpbQewBRk7tlw/+FgxiCX8DbVfdhxlTncaaVuPJVpTz011UT4Q
bq3zwflKYuF/Y6uRbQbQ3xfGkjnt35skhqvedN8qDTaaeuZc3pdlO7/WxtIlPeTQXPnOOZV0y0ZB
oe86LPkrqwIpF55s6neMZdbOoocZlQisL5GAhhpd/hKyzI8XOrhZrErw3Y6fd7WtgQPgw0UwkRyY
Ioagn7eZh87z4C3y7EWM7fg9fhP8NTzNac1hDdmNEyG79l+ea7WzQtnxLR6DQM2+KlQZV/1xWaq+
a49JNVVYszBNrLSGFnxEB2zVQwHs57mECdMmzwiQr1mGFomJB7LY72TwGWqIasuJNlnryqtBra6C
xWVIiCmOf3h17tRmxnj6VS7ipM6+fTDmYHuFhHto4Zjsg6+5jhqZOqF27zIh7n1HbtQ9iQ7BmHIB
GUNST9PnzUUZHXCG8iVI+SIYIjP9Sgx4xifgEswQ8P54ac74gJrdsWeOxq7vEIiDgfiBISmDr+PV
1d9RandNjvpxKsUNh7OkYkcYPmwbyRn00TXOzsa3XUZwukV9UYWArBM5/y/wfQvSI2a0dSyMXWGI
37sJP5eTS4mP2OTyoGD+znZzy2N3KwWOgq14vtVU0L/EciudZ4+6skTC4jW0+CDv4142uhYhiFef
eNabalBtawWzxBHPvZES0PScB4d/MqtHG9bcIS22sRqH0oLeK5TKPflsRsPfKA3epCRfl+YnikDf
bPPayvD7kMCyy2/UG4x+2n2gNleldszqpaVhl42n+0Vz5vYCb5E8W90BkBqXpxNvco4tV6oB06aY
5XQx1Q5cL2KMDANTuYQY/QcOvbrH4anOegkEnI5qdUKlMxTIeqaoENe31ZRV907V44cQ0OoZs6oj
SY/k1tUB8bY/pdQ3iH24/zCkzGBKp6vXryMNqdcgYaEauYOQDhsZjimVPfLkN9Cm432u/utz+NdX
IaulSN5B/SYlicgEIJBHZnU2VPguICwQ3DRWHzKbOQqDGxSbWMkLc5dQIX1rR8SiH/EZuIKcWuR2
la1MeDrdeOESOb2es4C7gyZw9wkffXY5vISmh2wI/84R7vBtGS6O2PvT7CpimxqI8mzKkNsoVyYu
WJF50B9zmHsa5QOeuKay7xJ8prA88pgtBc/1i7WURUnv4avR5EFVOuTJDYzqq3ZerqdMIvt/tdm4
cVuCG1aB6qtQJoR9cCSmTf4d0l3LniUXHNUGptDGYdSj2H/IFOT/BnLNCYrOfzNsftNC3Hke7bzC
j87iiLKBct1zscp5ey/u6gh8BHSw7p3yELFLMOTlCROC20R521i6I9A6XGDfN0sitn4Fk4wAhJXm
NGvXtg3sAOxPQHPZSmX8TdMLTwEHO3tOVz0MxXp7bm2NGGtr56r7F8H0txBQRg2ZDxvETj3bSzzK
Pzy85zbZ3IVog6gfQXimAf/Y6J4lAV6ZYOgxMyBAmBJvm+DYW1Rn3HSe91USln9tYEJta1cF6WuG
zMtuGPh2baCdJLRvMGLzW6bwGXvmNdcE+4VOlhED4xT237m9o46amvFmZ6+pw+UCXb5Gq0Bvp1/q
z6tFIsHGDD2oaNq9w4hqG9Qg/9YgPspDeT7SeZFvlHw+lhizyVJppz14cGsezX3d/k6rxTifJdF9
y3uQ5fwbxmmp3J+hc7ZCkcV6engFGxKn4abPh2D3Tl/b7m7WFiXntDi94EbL/05WXR4YoutYz+S5
m+XOSyaW2DunPgisCczeRzISb05rb9Yc0XvnC1r/bmHm7Qv3SquA/eeXoojgCTT6uxdC5mBYon5z
lQJkrURBU3aAmAW/Ztm+L5Gw852jedHJk1sG59f4D/0NO7rI2BuWHLYcCGgeVy8zuki/bwFZ5QPQ
/DFszYlOInjRk8lpMBbi3iMyVaDuU8nI4WsHnZaX7ZDYE1WR6z+ZPJiMgb/8yUfRZwyPAVI8Ci6T
2Xz+yS+YKGX+/bKKCMkj8w1OweUxF6/oTdXjSX4r4raJ7hVaeUkOvAMd/69wc9u2lcPO040j5M3n
S5Dnm2C4ZZjoQNXXO8uFk/gkgiwpAgxbjJ2ZxPQOm+IRa612k6UHflqVKwE6YBpCnl+Zmnl5IgSK
Ga5CgU3TwyBouTm8YJN52V027cnNlNKuqYSr7xSg7zFYrswb/WyDC83rhEeSccBwq784TeKi8Yyn
Uzo3GKzeJl+u4opawyTMYSIIabXV5alrkTfikI3zKn6XyaBlZ5IxdPrnoyb6CFkGh+GjlJSOO6bC
a7NhDxZiGSzcAkh9Wo3130C1LoGc+pXvM9mR6OtPk767xRrvxQYh8JXKrLB6oXy1q1dAVbyzjV3J
GSSW5M9/XAZdSEwE+xnvef3TGcpikWUaQNyvmYHbaOrAFclUZx1TB+/qSEWex9mLjAcmBuOd58rJ
ch2jrWE9oR9xvHfgGZMmcpby91cP3vnwVNbjL6bw4H5GlXj3s3WSEOGOeH9QPc0XDM5gJkrpTa9x
m46e5dS7VodohC/yNLxUMIB6OHm8/FLDXMIudTdwIIqnouXpi2ojf+UMDKNP/KeeBe9PKiVp1vwh
UOhUIz6G83g4TeQFrtqZ0lYRPcVwN4QqWY/fyA+eU2hXdZ5toPc9ps2H04Ha12c4P2k+QaAFzqGQ
VLNFxRPdfoUyZIAPYALmTpryedwvZQB+vEzLp6zQr2YvwZPhkS3SCSS9nPXQ3Oe7zv032JeEB8tH
gyvp/NjadP6N+re/yyQLYjVWFYSsSUmLJBNdmDrbEAXnxW/FTBWmOxnf9RVe/gO+vB8WcG+YEsB5
IYE9X9ljhwLnex4D18I7Hzy2n1wxxwxQvBL3OtSP06GELsGYMozgzJI/c+2PIdQfp4Ky8sWPAok8
N3GEcQLSEGI3i58x2GK6sctP7Q8FJc8CUDlL4jTvy8OVOqqHsE4FpcW+QiiRP+rFl6w+CgvHm2/f
2sK+telBZ7WJLVvV9Hb3EmpYH2DEPKp0Ft5a9nSAf6PX1DbLkyo4oejo221/67akzj9MODv8Zs3x
wr1Z9x8Ga4meagzDTA7FC3pznwe0bj1JYgY1NnLVBsTeh0rq9fvtmeXCKTaSAQSfnNC+Ntp5ppQX
fWfQySXs6yneWgaHn1ka9RxWZhSOuavCHBnRzw6MfXnOE0EN3+n2d1W4w5yxuUgCD7Q/0APFk5HW
Zivvx9NZJIX3Zub/0rwhcRx0D+Fk4QhcaY1QYXQmAZC6nwMJQ1Vtmfumnsa/ZErynCVayJr6pNT2
0kFGPb/tXmT7k79KAnOTqRwfxaaG3SYHpHxRlaZV/G7w5HHAP3q8slQ+ZlOvLxe4UAFhoiMzyUZ8
8JiduVq5w5FZEJOxg9ACAh5dnPqC+wVuXGUjmt8PsKcnBz9ZgqC9lgB4ESbpA4W+XE4UE2o1f+ba
AJ5toqsCuSp/upJugJzDr+xeLdW0sgsxX86Rrri2OGOPNwfxcDB4g34PlNNW4JqiUbGjoY8lO9Sg
KBE/9AHmYATozATI2gg6QQklVFQqbUrphbmk53B00OfMIE3i/JCMbD87Nnnsxc5lrSCpfkHEtU8M
FUlkCsAJa0uMWZzmgmYBuYYdGGHv6rd9vwWkXt+vrO7IWdlVmZsRKp62bNCwKP3kA2MFQQUWGRsX
XiFN2GaoMcO2SsSVtcfaKroNSv1+HJjtZpJUHVXVePLQ/tmwLYVFglzkdbZ07t+IHiw7vSczuOxX
B4w79qPulbIO7pHGt9gjUVnxjS04Kngmg2tx81ven84278de5isymmf+LlYdWmRDToIIEcaL99rA
JwoYRoe6yeQvKr8VNKXbutZWZlKFpxc0mz4pwU9TgWMmnRSsGhLXuSGqJ63Es3a/he7S/nXafcjJ
6uOOqCENa8UuqKqWsaIcDFhoESRCJQgAEgc+160LYLDerqUC71QfXMdJDRNp4o4mHy42AtkCPM26
gPv/JG/+AofiOTe/q4CsueKIpRBYLu73AgUshcykJ+8KrjcBLdUmefK9e4a9+H8rSQYBrahQBA0b
j1Z1D/A13ZFrF27XmBg+zM1xBhUO7IjPDn9/C/qvjD+P23N8uz7cV1oNrTZHarO8V8k1VNJQ9ToV
PZGzJ9sOZUCaPphbK6JUL5v1mfhYsMdl7D6uqgKJXoM4beGSyhvYApS/gXwjczgh+eR/MXCj4ruW
Rrs5GSyA5Me/A3Y3mTemOSX4sCjLSIrRFHygURnQmU8obgl6B5mJ/ubk0TuTYs1uPjqwaf27CM+J
2qOXEHgtLxTcKKhlR0EUP76LcP6jKozpW12tymPqLB+poh0A6VSynDtmNrxo6ZzfbtdRQkfHhvoN
kvHJHCZ+cQ+WL9mxffInp+M+Q17H34vvy33PE7XGu6gp1Mg+2NYG7DaIHT9lmSmM+ncpHNUhj/mC
b6aEXTfBR5IydtCtGgh2rWmjAAkiCFnERezB9ZYjMGTjjFL3d1PK19rSUb+I+wdALPNvLNQUx+ih
zbgh9SdNdRAEtb7e+13CmtRxnYw4TOULSy+Hr0nplVEhQPpc//Ydegbob5X9tdlapXKksIECPVHR
eC0qo9qvFiubDu9pNo/znyymrRyGZEx9zkcs2a+cI+K9P9uJYDq4m/r/aKngHR7aybdjyCha7DMs
ndz0J8EZqDpS76TUBQoU01tzjRkIOEKI03Ub0Kh6pqRny51bJb8jHZh3Vpf1+12DmY8fAcfw/V6h
TIMBBujb9DfubjkGVpPCLZZU7qXNWY+M8knKSdZM53VkEHRhxfy8V/gAS+BOFjWSWDzSpItPmch1
ioW4oxdmtoY2I1BfwK7g78jpqRn1k8ODf5Yz9AusbBGKxZIp2JQyp725W7n/CrPQRoh9D/FM73Si
b9xTPXtdV/vSNzbIzr+ueaBmZY6BLzIKNAXN/JVl2eigIyFJoMjysThi8R6Ql0lKcq+EzApS6hkQ
7OOyXqIy1i6/EO2qyI4xtPQy/3cLqJmUXdkRT0T6/1Yux1+XfRchCIxsWhgX/cDmwiNfzFIlxB04
0UURpNOjun2yLyIag1uA9zksmS8KU3P2klfX6jY0OAR+JrIcSSuX823NQXHcg/kkeCg5BQaFoDSi
lif5klxD+GNYhxcPoz7tujSi7dHqzotSCFbBl1pHPDuwF0mEH74bJN4iYhypCow9dhNeNF8zcSWY
YyH+vfrdxvpYcV/T5Sjdfrj0OQP5RSCyxcWzQK21pyJy5iXvvbsEwEL2TH60JTfCPAMk9c+6FEm+
5nV7AJC0a+wpuw/OG8jl76EkjpHTXBnBUE/suyJ91aNx/9RH8VlL9X3+XWz8TFL9mvNPqKmj5akh
vwsmoiMOy16caSwwwDS61Jm1h5D0L776+zhhfYK616iRurxsDZcPUb0rP68waImRmCMJA7iW62l/
ufjPozwrWN+vjBsVfKC28gN6GwBEG4H+RGXgJh82J9u592AxunLTJiFxkdxNBNEa13BktkxVGEDk
6DDtCeEri9VdsMHJIacFPKvdCkQGqi/MWvmHHzbdFcGRyJiDuMxXjI2k3OQWnbVDnVDajSL8uKTW
zTw5dIBjvb0T1aszgs0uXYgA+MAritReN+gAaOki9SsaPVuvfYbWr2M/tlXm61eBR+sD9W14vO6e
fV0h59VUW6lBf39BQvp95iDV0NobfbEb/LrjKpNH9qGFphswiPmJ5hKFSXptmBDbS0j4bPpywLGF
CwaMZIl9qX681KgAXFMUFY8YNXROR80IaRjMrZg5g3C5O8u1dn83slfOdiJmzI9v9QOMHjoFKAYn
GEGSwqmhHzq3SUvy+iXroxUpCrLCV9hDo8va0p52Stae6R0XE3i0yFMlohA+yBGE4IPo26DajmBH
6C1RI7VqDG1ISiGW7S9Xx8URuGwvZgvk+Qc24X6zCLjpt710NFA1sUfpOGMhMowHWqCVQudimaWo
jTTkfHcGw49Vhrr7vt8VcLiNePf39jlHmAeULXoBE5Av7R1pNz2ZBL5LY457fIzSRGmiEC7SOfI2
KfJqReE4k5w3eivX2z0LBQ+QhVRSDtmqLkptv+vKW+s9ivy905wjyoKxCbbpqTd6Aj4iGtPMpLxu
zSE6XMd9nuvYRXZ2UuEzwYezEFb8SGQfMOrZc8Tfrum0EDRgwZWBV9wPo1m6qXbKRO1NJVgoE0dF
us5aFqnoVQaccnr65W3s08UA5zrS+wGtIs40Pskava9ogiPFIrrrnI44XslmP0gJlu5tm3FH6IPd
j2bXBmIYkYxPvSbAIr3pFGSHSxPVlIetd3PC9Oq4T2Arba3QyR7731Td2GISLma7EFFMMLDcqsOQ
h6u98FZHCdRTyaO9dLFkW5D6HCWwEzLrr3PwIeXbXvEcKtm+wS8O3w7tiAEdpd/+oCXaeBl0kRnJ
8b0C83m/+KX0OCDqZiARiDAOnix6sG8esXOWsmIDc1D/xnvoPczTitcAW2muebf4DEqXaIKJ+DZ/
zEa+7AXJLx7YA7/6R44XXqCmaWu+xLwQp3sERnkkg3ItqVseA8oFEyViciNtZUin1N/ilpENib14
RetPZ4ZAackFOi3S5FDHDXYepv76bkXicX5yGwjHvDdxWTrPvPPkrbt98jo6FPjr7lzdizuQPgq1
p0tyYiAOOpbO2Q6gt2zMivjTsQfVP0Xvz4V2QUQTmb92xfh9Mq20yAEu/N1WDX/YNh1+gukiKNwS
zo5XDSzhBKNzLXB7oiOLt9MI8ujEprPX06sS8MNk+7kgOJBeGI+tdkDOVPJDuUYZi8HBevsLkkhN
X7Xqo84UO4ECwPdv+lti+d5+Hy0xt6B1bxSLvsiTuvINx/gC9Z6LPcWi0gIlrkoOXGm3ui/ONdpK
cq4xXWvlcW9+cZynyLyN5WExmcu4drk3yC5UyHaYf1o/rauOd2qYF/P4uBkl/FoI/ssVkP4vVE0Z
vJ1cJxp5u+oAGfcGsqWIHM0S83Poh8cFwaqEIDHn30LFN8S0/3+SpsQ/7mepJgIfEIu9T8feqPN/
fehvsfibQxYR011xn4ZUyHI5sXsviNGprIxFUTH/066jx7p5gNDTSnNu1FkZftNOZ3tbrCXLezKr
JSioD4wadyt/7UgMrv0mE7uup6RHTC12fD92udPy60DAgMDP271RN1UxAB0t5grTGdW4vpib9atr
RLRRXR7uTIH8xgOw8eAEG6jTF16hajm5fsqv9ELyaOaXqDbsVKyo0cZc7+bP5c7aJo6111/EJOKn
tOJUwnOew4AsRxLp4Q7DXCJ4av0Y3KBL2mq12bObSHaBAXDPt7L8znrBJ5AYa6DYfr3R3JwfkDxL
fzuKemxFlCoRva1nBhOhmd8YHHEOBHBu1+FW6a4rnCu4N7baDq65Uv11llIZlIfJfT8clRRjnlZP
4PS3nqelYprTUQm38VT4HqOJxamoDTSmJKoWoMlMqIC10rUT4b+gU//kZ/fVxkvgsjs2rCK4G6z+
a645qaydisFiAgSVdLkftGqa7saqIBbsN/rDAlblu2aw+nWaHjgNcXm7f+SXlImQStdxXRCznMNf
hGQjrRmvoRUKlxaZf0RFaguQV5LA06+KiyT+en+bz17j7JLoa3nY7P/CzloCDscwPmE5dHSh9dy8
hfmjtuZ6Km8VH5ZOarbeerC7Ds/45DU5c2OEnXsPpd7oatKCQtAMBfsd3a4LtXU1AvBWU5o1TdOb
n9kbx1oF1RYVJ7Qa+l1WdnogrzHjaODRPP5Y1F4ScJzOByeLOhZn/gjV6sUwIdDk94c3Oxck+rc3
lgtVLhfy43iFbg3IouxL9xoyZbF3ZnCzSgb8EcSa69/G1FfTYofZLAXWNp68r2q5RGg4vHMItmqg
Ami3dqEOmYGT9rkKWNcLM/AggFxjrUABbEg6hJyKMFJW/HXETDIVhV9Z/fhmdMvT3hMkE/luPH7i
2kI0YRsCtc+TWT/zHKsLesvHaos1X6MPzb2rKM62fqQRCr0wEexvOVUhcFLO3ABLULz4p6F/QOa3
reIct3tTVoMNmcwJKG7N3q/Nnkb5IvbFfA8x1V9iuoIcTA5vWvrk/d+L13p305uCwPuqL2qrJsu6
rRrXvf56UEL6pYOSDLrO8ukbNdPH6VqlHd1MNUAxRM96A5NZri9sjrIBg+Ja/aCboMyxJMGPv6hO
39iOZ4BiWZJFR98Lb4/OCOuHT4RfFHu/eUiLQM9Ridoi8bAYXyPwjrLBU1Vd0oWPwoTIFAOHQkPA
9HlMlH0hjJ6qNwu9tzmTio9e+6kdf74jwRovHai3lIjNMHN3QVtpoeRKTkeCYbtLwwY8t1zQ2k/Q
EPdgP2c99O5WkmdWnEWqOtchLtMzdcKZPlj6FTbieYeNYCKgv8kZBR9SkLv4BXOzpdoLjwVUcTY6
J4gCMPXDmAyw6ft1A0Ln3u/iKA9QundAzW2j58mVEo1mlQj8EBDCpOs5BaH+SPltOafXasdycEUy
m9mWGMFL7cnEVHMmGdtNOUFpc5D9Q2eQAgNjx5tBnX8uKt6faQ+aGurCnUjhRAl9Mz1YjXDeS8+/
3H/j6VEfomoPs4gRsV4GNZHAZne5dbYFzIxz8N9Jaz/dEc+FxgggRhrSVjMPfM2c/jI6CldCbomE
C+wZ2n/QH1mPrdB5pU7IdCoGBLRU1+ZZilvmKuNxzrE1jvXn7/edj88rxMDPgjhZKM3nArXBa8AJ
6hsUN2pjTUA23DYcLMtgue7OD5TygQcpbISsrbkujK/iF55dh2H/mr8IqcKUHOAk2VZTQ5Z59okb
7TH3/zkub+adrd4pMbHNE8nvr5RIRijR1QlJsVMqAbuO95myJAqujJdICRJoNVDDye7aGftUQw0p
ue927ulz2ILWyIU8q/8wfEzyMttvnPs2jev0lnNeg2trOxR9EIzAV5vN0wxJQvoMBRIPtJRHCFRC
BWHzNiQYHivTnw+AxqMjzdFQXJm5EueKGKWqh+rdQuNaXzUFXOIAq53y1reTWKsPT7lH8BMoZPzj
n3iq4O9FHcoJeUF9Us8/AUCpjK8bxh/c5XccwA7rbv5lCzy45KC0ytn+DC4hHk+n658X3TZLq7We
vXUThSYKmHEYxc86tW6jhaD3Ml1DhHY1XuphFxYEC3mvjnl92Vp4+VfMiphB50mJlX7B4ELR4fbF
kGTE7uIklG4N+8+pMyBkAagusQCTI+8cvQsqm3c21tr7tPaT+iJSHhyTU7LnxakFj3HwMxGAu+Hc
tTms/ep7HbPl68BysGoto3moJUQGlHRLl1bwxKIsxZVeR5XIFoSKzEo4EpG8QIf9Jxj8tktVDwbQ
Ob20nZ43AglsgWorJOW9SubHwxP5luJ8+h2e38RaDk3MBMU6tjw1e/GD8lljNUt2azs0vbwI2Gsh
8grl4uu/N/JIt2Jgk0qBqIGcdUkfHNjavcP1JO6zcbiH9xgusUsqNBXX3F3sl+S5kFwmOSRihk0E
zRhnaglZRfdS2eKfIIFBsLlPBEFPDvZh8zMgKF9PjgKNPfS0OGt/k4Isew2QCN6mAAiMU42M1IJk
nG6Epyw962K55VvCN7NtKiVO4xpG1Uo+VEooD8Q9epQhRTYWioX3gnSyIkQWUd5EhIKw0v425k8c
XI7QGlmP7DTzCEbe0saz6eLV9eTHE7dty3IRmbMsn7nYpPjVlO6DJVapYaQyWm8Z2Ryv9DEezsWk
XirLoE7oT41Y+OCc6RVO6OP3eTbCCTVaTchV0Ig+R6T4E8fAjyfho9fb1UdqgX3At3ObPFXZlpJV
OgX/RtABmmK2BmQCGdnrBZYEf9vxMNLO17jpVF6Z43irbYHwK1hnd0hqsvLMhL6twVsEU00quJlG
TYkT+gf0G0zkNg2zPR/ggBUlc9TVU5Pv5gHng0l85v0teCvNLqx+q7xwo2nr0fkJOf1d7HRVL+/t
nvjBK1fGCrqPknScfxI+Fw0IOy5/R5/4uiceKT0NxemydW3m6LaJm09g5T5YZ2fQGxdfMOGD9ZfR
v1hDWJbOxdoFumi+Shj4AZKDCIeIx7DLTbkXK4fvxa0C4wTTqNrMgOqDYnxzlXoyUPbXeyMg+/co
GZwILmqTh5hKLL6t1qzAWLEuTlix4ngGYBONgqM+b2oaXI/kyZOKZ9ezpQ/MGcZVFi95FS9OyYNt
dat8+dFxtyS8KC8XJK+3N5g9rsicCkJJNvjiS9Ebn/wkJ2+yErcb7J4M1Ca6kGn3twt2pkf77ViV
j6jWtAdv18g+8mFVnYn6kHnlceK51lsvfPNTarKMxYsxxSsy7N2e+klAO/1P9iwjEvlV7NTIeP1b
qk6Bua0++6gPnBq1oYNQCVtrNmpDcyxMhHFeWxARDg20a+qOk4lwg6ld0Y6LVUX5k2e55OfDWtpk
ieTQopiskgVVD4Ik5haJ3R9uHmlmhu6zl1rmb2Z/QepCnmnQ+JSYz1js4Ql9jqB6KgirG3uU4Gyq
gF703ltFeuzUfFDWiXmOuLoyLFnwOo//p9RhP+8yeyOilSie7HPI7tYwgIhJJ2Q7hS3deOkZtqkx
umPu3rJiuBrJG2n8H2Q/EHRmuySRl+yQGeT7rj0IfHjBU7vJBLCPFbcsGKaMcyp4PsLjuDo8AlDF
LUor0QLDLa9Z66nussGD1Js9XDMLRETwNceRS8XGnEKQiY7BobkVpFEDx2pPHX2id8ZOZASxeRoW
8lam4Um20FCOeybcJ/A3S7Lzj1jv+2YjlVMJ8gPsQiuT9nOw7Curyvn+juBzPqhQbw/hpK/3GcLE
z++jgV/qm34voukl3jl1JwcmME+X5i2kSGMdGQjtZ+itEf3nwI7Jo+s7uuJgcZfek3u6ob63w/YD
kbGdl86TEPU3YtP11Yc+Ex9IWZnrN+nBphCj9AC0ySfNgf/tRnZtPtZT1cmaVZ1rO3LPo9v206eN
Q1hxWyMfmnh1RvtSTnMm86+5TUZzSu8FPdv/gtsWhMl0XhyO932cDhkFYJ9VSSxoPClc5WsSnVN5
I09ufC0JBkq7QoqPMoizPx6wmiYm6VuSSXROOxKyfe4y9emkIycNGenzWHro5jZ14crBJsMdnUkY
MjBbyDPhRx24sciv7ldObuDoDVPJ1gBvPOg2zCRFP1nMdsPCwcVyxg3bk6xzJyJlpTxPzLjFVljP
Y+QIfqOlSo9Av063MKN/l+Bkm09Nud0+DATuj32pR5auShJppGFeMJ8duQpaPMS79ugMcRZt2VNv
g6zBZfhz0hnGxZwg0XGpK6rDf5nGNmxetqkeiDBpFlg8BTRdHKMyWEbfuz0dM+jhpbSKp7nolvSL
ukVg1bfnLdqNcI/P6VZ+2EWc23tGPa4Ma5+fXxPeupduXIFPISqptmI+1u8vmu11qwDsXe0q5RCb
xf8EvfCrKlTdBHyrf6TDDxTbew0h8LWOIWvUBd/LkS4Myxw3NN6lzcQ/ZHB2rK29zsKIpvP2LT0E
EGwkEeix8wZBukArkvpB5sEqX8k8/H+DB2pfIp8JRauZFBGW5UXft79RDVGXjxSqJknevmb58O2Q
IgHuHhMFnq406M/8+LXSysQG/4npnPOO+wbJgFElUuXYF0hegZQ8c1nM32pUPfNFRJIG3sea8Xv2
6f1XxGHYOkFBXpXEDEqHZc+8swQk+bpfjoiGeQbkZ/FF7Ocg5QEZNVLf9/QqlNfkNkhBBKKfbHfa
u5Q9lHgTEmsyfLu/6570eMu6uVQ6BTnJGGoOSIAVMdRLtlWSmuJ43tu0EqUCG5YmbJq2MEMYgn2z
x3MJeGsybueh/mQCcmc5Gu4eEg+tHrDOuZVOcJDxs7zzeG7U/ZKJl6ICzxZ6tXOPqUo6jIYPLMK/
aINfT7Yc5yCtfGqPsiOrxgdy1zAimeVJAa2jZSm3f/FewNPNrOsYYUPi0zL6rIi372VLYd5J43A9
Uw2Jzs02Jro+5pwVePmMQfqRnU2ZZm2s1NCFS0hFmByn0CKwNAw6JjdnpvBF6UcBdz1T9eveZZdj
JahLcvhBAkAX+0j8HIEjqZoU53TRxPomUnG3GC1x6jeDzIxIZN1BdI1+T5eSH4lE6FFHzEuw/J+H
lG0ABG1iHPV/8IncGcmP+Cz2Za4/ER5/WTOSOYw+my2VhENqO27ZiCWh9cTp2d5jb1l97UZVgHFp
45jxlMFNjv6hc+hPGARY7phuF9jCeMJFtvYmfmsEOfTMG9e9yqvS5hGMICT/gSXs7gHRufVZgypI
a9fYuPFocETdiv9fGlcD5fTxsIW1N09/ajml42wfVCLX+1bYmGwJD25wiPo+B2G7GTmPWLgLiqrQ
MbgNkbHXNANZ9s45bFKnN41FoYc6znWazB7TZnSBDgrUgi8ULrVCmShWex5U79v6Gqp8JRoVkEKZ
Ucr10XgTgPiEoPunFNNIX2YVLILE8z1k8/mB0zShTzCL/beX4O/71ei6n3A5CX9ryfw9d1AtYph3
x4KCQ+YrCJ6zAtAVjti/pDi0jq4EfkyMAZbvxKTIgg8e3C24VgQk5NtV1g+qKznAk38HZvFRv6v7
6vR8Jk8v/R225A5eSWr3ze8wFY027Ry72GdBuIBGeYQ2iaF10PSzEHK3EWQp54h/Az6/XbTI50HH
ZsIfm/68ViXUBcvlC/Goqc5s/e68PRSCzJa+GB0IpXD7ueJu/g1As6e8vqXfpNkHTD0xRF3TvVhx
zXTyiUBwr8Izn1b1ZP8sCwTZTnjDHtKnaN9mlctnOVqYdsGQCLgd0C9j9fSQbeHb5aK5IXRtGMrd
nFQdPlkydUYf3rB0F3ARGCVL4czAG8JO7/IwM3lUMS6LByzAWoIqpMCpcbDEMqw7SoSk8696vBRF
Htg0S0o1khpgdNPRa9/TjZrOFzzc8nvvYY8ctlxa3tZc0s4i1a/nK1kL8mHQ744sNyeZ2wdy4ySK
+lOqvm0KubYU0bWJ5xDFdVt1Xxo7La0BBnc+CH/BCAKvyGi28lV5fG6q2acYV9W114OIkpVVcB3L
PHcmcQw8YDyTakbkDvMcdBeb7ihjmIjebotTsKbyOpmodXx63gcbTZh9gDisW3jJcxMMBjWXTcP/
/fgiUmyoT6ciTo5vbwZncu/8eSfWYPVOjSDZvDDQNx0pnoXZXGAKhfYGpuhM54gkyOLwB2+JM8JY
Dmn9m9556PPydNwOqagaGKiV7w1zf3uY+Bx0uF33TcoSQX0iWwHue0g9LI94HECh/lzEVQopGLHG
DpTTY/rvUKihawiuXlQbuLyDAI7HZvTq9JnrMEgAS8ywHux0ixULoptniHTOl2+Yp4rY6iKRv92X
+Vx3yq+qQbtdfmH3+H6XXFI1eMZzbzaz2FJWFDn0Tdn+pmw9En21GP0K50nEZjlaf2MmutBPgPYH
sS9v0CO8wBD5ioqkJ5+gw04dCY53GYmVgPkWAa6G0GlBLpB1K/XZWFZVGLIcY39x3s4118i5tBTk
5YYOf7Fn1c4SQP8E1viKxIXDj+NSXkD0Vv58Mh2qKVsHZXoR+uBPTBCtkgwWX+gux7Dr/0IaSm5+
Mns7UJTiE1+nzEj2YgSyORjxFdxS9gyERhz/Wbhr7UYgIjWq2RAtdv2CIaW7N6bv6I98or9Z1LtY
uL6TO4Jmj+M4NrS1aWEEH6ea1NPpQtDjFqHfnYiDpb4ts3vc0vY60AWzbt46E64fyAc7Qed8vWpG
VkO7pasoWeCCXclLXI7qXNDQdGvytp8J+sLDRadJH3xZ0cF4Q9lWvu30I/F+XF/kXLxEiBBsRNiy
lzPlmkR5qFdZ8kgSyHvg2M50FZrV9EvBCT+BmJzbOuC9Qa5TopImKJntPaH9etEYY33S7avgdpV/
pLTb3VeTdYpPkk8EudwozzaYCCKrwL1l36A1mkeRR+13/uoKbxYqNNReq4jKO/tOBiVTaaJxyCQl
4/RD+docRGCgUi5/+5GbLOwUt0+42GeTNTnGKv3GVhDKMZoo9G/oxZc91z1JCU/l/s7tpGsZL9bM
5JgXFyQGyYtjLlF8dyS9zr2rD8m3EI0gO6J93rp5BWmqDZbglHizYPq8llqeI7j/g3oTxdNKIJll
+EiQiy1jwZVaD7gI2ZV3oQUDrHx/k5MjAaRH0R64Dm/mrkkuw6InonsMZmY0iybEnIFDkv/QwL3k
0V0goWpsV1ndT9R9EqIdJl5SJCqfpxmyOzbmIqcVv627BePc4920MX+YdaBM34XQSapdeFyP7rJ1
avb2GHzxeo402aAUTRvU3exLP8BLUTWpSd2is0ZsyHr90jaZG3FdmAVn2DRZsau1FEwe4Suya849
L9EL6uyElg23qkcZVJubKydnt/82M7RHhdRt0lGcSw0J3UKLJKLc0KSJQ4mDPi3MJTL9+uN1FG1J
aOQOsPWRGVOiLxrFHt45usEiXV2FWk/ZZ7s4zbXLEqN8SkXaw2oS9FVK4nZSOI+huX3Rxq25HxZl
xD6pgQQDR36DPjywQclnyLry6e4MlOuZKaFKzVAb5KoyzCurb0Cahf+lRcK/peLr25Nrcle8fKKG
cdhrFurzCWeC+AXm8VmmJ+P2pjM5DVa/GqbZRstWxzBYO+s/NmAjPtJ01fP7oScd4Ca/ZcucW8bB
IcJX0a7HvVfpUglOpckjXrws4V7LRw0DK95UlLTFdQeEfma7NyfnpZZaXSPV3JQ57j8YXKuw0xL6
hgUBRCRwi0sYcveov76ZfG+YJzWqBc6gZobaS+/NjigJgoMfrDw/Kfmzf1SE4cHOzlwiKuPQShb9
OGdA0dKTpcIP6CJeIhhL1EztsGvbZjDNWlb3NTYexTWJgbVZma6zxhq8wHL9Ux0iPwtSnkWhywmn
Y85Wsp6DR7YblFIJbYBPGnhmNXg8RECTo8cN/O1/eE6I22NUtDOSOJI6DFAtvW5jWMoD37mnGJeC
wrqnBT/PXpsGSKYxj1aDaf9T1QHmj02XR60HC3pVLv/7KcpfOZZrsU+fB/wHE99LfbikfYtTJjHW
vFSxzZADGOIeNbiPhl5za7QDMqG4KVWeFwZCgTu79tGgXvAu3jv0H9Phf3xmjkf3x/Je/6S9bz6w
Nbx27CuTzxxgRk4/B2i4976uQBdp56gra2uju7Jje4igIPRisQ7LoOPQHhmiJFuSnDT4u/SMtebU
2wnyvhFqy9N1HbsWEoNUlKLQRfnb7Ng07KeHE72+8qVnbV0WHgE9rXZ4jaPlCqZ+KFNqealu5r0B
RuEyrfnzxJR7KuU/Jmx3CSKRYMzxWdpGhsDVEpfe7sFFHlKY2e1d7NS7Yt29tbf/+7Bi5l8l+Dbw
G6ViYzRJHsf7Prvn16joORHWg532kQZH9sljTNYxTHCn0B5CPSLSRPANmxyJWGDGg3+D0aDyNHQJ
aD54jok5GbGWPC7P2hzcdMczR+2CgqlyBLP0paVnTbz0Hg/T6FOw4M5zBNlsZY4SVwBiXaecs6P8
sWM7GzcwHVviXX5m504l03mIZnIjmMhyXHP+UWsqPLGQrLrLjaAOEFINJYlJZ2cHu+Q0NwxrNrzj
AIzE2BOvl0qN/mdLE/viPB9jbY42zZxAaJlMp0DU70fMuo0c/2qVCip35n3rAC3huP0MTD9UZyqh
REoem0RFHgAOcTtXm+m7+B1uklw5qLHaCywgwd2zsa2DBfF6+8oUrUDoyfIWZ4JBAzq/KhmXx1BX
7fIgGo63cBlLde2EgQoScUd8w/W9UzYTKZ0oEW5wu1enTDnUd4uzNEt41gWnMKDgM3KfYXJPhroD
RbGTiuO8lagdYUr0e6AyKQu3riwQPUfEL+hPN9XFuymaP0d+hWEZqNHdCbkkaMK2Vas5dnClT3Zi
l5UCwoZwB6OwdqoBqKgUHSew+0qjDweRzg3kovH2Ldn3EEFr6t+lGUcAYTa55V453IWbZGzvlmtp
+Y7qEiO9GWx150jV3h9Xojwmae6A3o8TaN6j185QjpJRUhv53x+5S7FN7wqtx5v3x0rjdXIUYqwQ
wpUcwOCHPlvAU5u+AJ1tjihliZegCwwzew1nlVKyI7/YvavLx6EYLmCyIjARUN/U8eMtDA9gI2nR
ioVJW7Om+3p8Sbgj5jWIJDtq4XsSswOPBZfiwg5ngUmdX8WgIsp0VL+y7UsLxV7u5jxoLByxPB5W
O+26D7CO7pLBo5CGdjyaH9771f8h5s8Fn8V3vLDpIUgPjAmTNZylZC0X87fd7qwIxdo6tpCoqQqW
xDuIIK7M4KZWwwG0JP3cGJQ9Rr+n5xn+Q9EbfvRLN00fsa0a1yheDA1BEE0wH15G7UkDvn5s1u6z
habNkWtOyaX4EGAidWbGngAvEkNjglo5YXSXAcNMqfmgRv8lqA8me6IgMCQ+GrJ4o5JOfeolbfKa
Llfi7XPdC7bTTkgyydBWEg9ifPmfUjndrpgczkiGRiydzmOMp7cyABCmsO1Q1kKzOLWr/IhV2LjC
b1R0bFQEMchHNinnP7EtvlURcniUq8S1CrE6TgDb8xKEb6hVL2Wz58NV19UfaI3ocDeoFNuWy79I
PZfH6KdIKx2xkywP6P0Q+Q5SBbPoPgL20o9sYA57CPCa6LWGmTcGc89/JM4VX8Qvk9sO37PFZf/P
aM72UG3MIuOwH/SsVdGk39YzetgZsFt2YrhwrT4QlwRiwkWTZ/3k+r9oLs7UoNObIgkGBQiuuEgb
UPtJWIYb904mSXL9T7hVpjHYoC3PwoZD2yXq/TzSPeRPrOhgAzJok8xlPnGU0jkZVANu+xgDsQk9
S6d1D1+nyv6j7xvYG28E7fjnjrWqwFAAicY4QQTMggk/f6xamLXUYwXJxEWFQZ2K+N1pnMYTCCND
R+9DGqX4LkdV8SrRl/TAgXLKVdZf4Q7eW9hU0vMknBUVqHRoVSWkLyg/yu40ik/sJInWWv/anNmK
HtkLmT/ut3/ejZxcwpL6slrEmF9DzuZLFJJ0WEq8Na3qUXOe9hk4V0lmMaEU9PIE2Dbvzn/ohKNz
DxmeJXee0TisTtLURb8pOySzQBIVBcB22SpRKq9kV0EL9JpRx6v9VhDtf8Z4cPFqcMqrCvckbfHX
xjobC13WKZ+pYyWvfkfuGzlMEzrg7weHsH6fugl7eEJEFwmW3sJVw+8Kf2KInxvbEeKmnkEYF/fT
HV3H7ZstufnTJYu6ZyEnB86jKCMIJXPUi7iouYMWg/WjSxr5vEvnoGze3Uadtcu5e1yN/s+KJB3A
kX/zg21CxlUmastgVDWFr2CFjWbcUIscbQ257zO0tmUwxU2zaqTvxuMiQbp5nfn/Ikcxn2I5DWX+
uE6Shw7YksuALyVuViCfFt4xvdpUnuqAhCryHu/MeD3uQj4XFscCa2NQJYzocj/taHYYC4nXBsyL
XdvOGIzI6vX+1jegvxf1pX0ViSzTXnbT6hc0MRt8Nqs/HWmAJ8Mjpwysu77MgEuSc20ilfG9Mu3f
yEKwRlkwWDuD2IwPqbZqAAfZKzLwUv5D0KW69v02EkI76VLCDbeHevgOb16aMeOWkgm+XdpATjGS
EOCqwnl93VtVbBNHi1140nzSDiUMJbKjL06+BXJNc/RmqJ+GO4ztgpX8OrdhJRXvBelTFHtxAmPP
dlTIQMEjOcKj57mN/Hi+R3zonLXQJ8JA3UcIQKuoz/WIWjbuY0jZE55pv69HCrjlUh9bd6FLbAS0
Dx56bZzYzXTVyDd9eAPywXC0ztA3ea6FeI5RkKRVcr+M1PhG2XdjTUtFwvpSQrmgb3cM2tO2ISGS
8Rcc/+b0S/XBSzHGjzvu4U/HitA/l3SFz12nDiisgeWMsW5QAsQn7OvVN78UMfd5O9Nxkbuywv07
pERi1nmQRIlOMakRiYTzomMDwKszR/6sH+L+C0VsLkU1RGNZoF0rnT5cIOaOpDa5WuWIzM11ze9p
D7YcxpLhV6u1bAOOfGeN3UYco50h3PdMs1+J3ccEfoi6P3SOT9JL9uepR2ML+kJ+5wExAFeT2IoZ
OUJGhQYb8MRYaUOcibM0wwefuyJ27sG5F+V6hdWAiSY/Ck/b0tugZFIp/Aq2OzwChUFYg7Y0c8O/
fPRGwcjkR0XF5K4KjTeXuYRAzG6W4qt8mg7/Q+269il0Wcpgtjvp4atgKjmTy72bZ5femgBbqYCx
7p/RD62bT9MIyWH6zBbb3RL70NQrtRET9nqmihNDfIIxiUh8zgJwIkDEYdnIJlQw1eS5qbeaWEfC
sR5h3nACcucEUHoaTN2ABDt2L2JaPGHUQqkjzc3+AvhY4y1JLKbfkcGAUKTfkYwxQoVOE/fGuq+M
+rjjfD6wMDeyAkrxGTb84Ivu9QBsa0QzQg8eGTY4BeA9NHZHkHcQ3JN+IvYOmUFM/eCUFLgyZy3b
8Ih4yVqRAaHMoL08LKMIdyogsevHtAhItFr4PifHiqCs2c/02MomWVI9r2fIm6IqDNG3a3e7W0Mw
eklgYu5I6NbiDnG0aZq8lhcAF6DopUDKfTbFr9ts768bcAAUk8wbEOHKhr6WxXIte6t0NJL9hg7z
7Wn4Xf1H/Yz2UVTfSe/DZcvrZPi8rVUwVU3Em79+2i5fqTJ0sjp94UbMUuagAZhqwjrnrbjgvZb5
C7IdHUO0dR/0SnuFsk4sUJoig5D91unX/l2bZNHB7SeveGgY5Wo0yTDoCFv09sfgg1k2W8titkJo
nvraksZ4k4tqO6+yGDAmURofo2sgMCIWiqrAr2QuulVtSC+owJxApKe/NFM+8Tttar01nUl+Dtqf
MHa2g7SjsluqlVXS0TMhB1XyV0iJEFAclUW2IYeT3UT+b2AUsmZnL3T/skX7EIKwbTbyn1CUXhuh
AmxbcaS8zKkiIa/F9mt4sgVmHysLUyMwTKfjP+Y00s0NHRg77AOIRpT5uNC6ph6Dgy3+EegztuLx
DxtOuoxASrmdaf1PJH5e6VXXMfV/zeYjbzy7Tm9h0dLOm7vKAPYPt83bC8BZ8FVGOLphvCA9kge8
oJY7xbVnf4dusf/hjl9Hkra3drypuXHX1QMSE9liEtENILAy+p5bfQoxt2HRCXajfDucU7Ut9akn
7COsyCtmPh9SX+xWnE9jwsqst9FrzQu829mkeAgwt1KR3Doy2gUMXonNG48xk0zQhQa8V5v032fR
TntRX5lRc7GZ99JuKJXkO8p+CZ+8O9Kve7eSBLHeD83ot8XpBqeECvo0Ox0IUI2XNZueO8HpXEmE
2+X1V/rsrPjdR1BOpbuFn+tu5dxgdQoOhsQ0vXThcLkE8HtjffSvqG2UQZeUV9r8gX78ZGxsbTr3
muqqLquG7VQpj2Kqo1Ko72+92o+VL2OPRRn511Cgj8uLx5DsdCmxPLoayu9x3UbS1AumoJ+rPckH
6kzK4MVfD5mYdZbemxd4TBajm1NMcWBa7QjYcqzxcv/MzhevP/Cpsq9Kfk12x0GQayrgHDhke0sv
aPWlXmprJ7lr6OElZl5OZlC0M6Hm4zsHKGPfl2WcBOg2PUFup8d1+7DWqOAzZwlZ3VX8162CuerM
ypcvXc6HEkACBZqpoZl0CnvhbOkH/Ty7oPXKgFtfdjhOdvxlTNE+oDIlJ9hZaSv/ozaS99Kh+LK+
DTygmkY7LanejGMWutn++DHiGAgP4aXgHIv+aZvYEmtB1beWxzQ3+tC6BWWcHF++b5ssPpJILa5B
vmIomMtqhCGwPBAjKYM4aHnECzDTp2iqy36y42tL4Tk7Fl7UdDKfh2Ryxx3Lh54Nifdu+/RCj4cV
JpawL+iZk2janzQ5zReJgtB37G28VeBHd+JVFJm4y10PNs2njAg9rLtDpfXEQfw7iuze3iNDScQE
aDWn4ys4DyO1U/+NVEmKfsV1KhjadMBBx4MgjCZhEYHYweSjlfjevJnipJajE0OblTR9vR/1E9BA
CPhOs8kEKx83wj2D03T2pRQx78p5cwaULsCM8F0n5uLUVdQpZ4svTUyfSn+3jC7r1Hai3EYWQHa0
xiCfjTxq88udfqXDw9LyGuG6VmOMVdKe76zJy2e8IlWjSAtNxaF2R6whLreLaczMEZOAt9knKNZP
j4Ru1Gw79LzPH/y4KK6JauPSl/O7lPLoDT6DBp79n4aP2t2Mo8Zw0dg+g/tvc8xerg3GYt5Znw8w
84hih/9sj54NfO6nURVov0yQbiFc4181R4RC//X41gevruURmVoHpbcn0LIAsVYkbGVb2XzVSqLT
Me9u5jZXByr3mQ5vaAqQKsCEk53mYz+2tHcQbTiSe1O9ncf39lzsUFqtAv7Lz6AcNoiOLKhLO5FF
Gm4L+PdxhrRPs1GQVmOSn6xh+TaXUpQY1d75OidYNDszwdNhHGsm/nb1FTvDpbrghaOa4V7sSemp
iwFLbOPP9CMG+LpSESzrSZmA+Fm+ygSpDkpcAJuGVYlEtLeMy1ErJ0oITRVlSVzZDAWnvMUlV7Cn
+OVo6PeHbE3fKMZFPiJ6nMp3DhfznEXY3XdvR44YJGl5sUbr0MP9VniPZu5G8ZdAwogmmP7WTppR
ioSr+MTMmZh2Ps9n6jkQdS+5wwy91GGx2CLqCnRTm0eDBBWTgal9Nc3WFwIZ8mhLy3zZVlLZrLQ/
pIHpzNeHysgNt2cRCLCI5wMkvQ16a+kqwFpf/cGDKzyPrBSznjwnvgzwQvR99SvuKijejPfqCZZj
CW2TWOxjK1hfECbG5T+RGg+ewP4gmS32slGLs4IRhkqFaqZSFUmUEwppYv9oIOsuLYn6oOeoexTM
dqMBKmg2W1k5pkiOOx2NtzvzGmUo94SjfPPr97iKG1naoGyqSSHAGp47K7RPpubYJ1kMtB7tVWZ5
F5r/yDeoJJCdqoXTz8kIh67kj7BuTI3GdyLiPT/xIoxUmFyzgH0OtX17dzxz+ImGNIqPs0JcpbU0
gm1rxhCgUPPDHmn5bgFdeQWmTUQWSFGkv7tSyDZ091BfW1Wfuw3SRgyCBSTfD5Y1k7w6lKZA2IQe
Dc/OKikAV3Se1dBQraLgSN2YmOz/RQ0WoyuBlHDWySCxDscy09tqAWel0ttsvRNf2ZcEiebhf1xi
tlMLum6OZyf1D6Q3+mChb1eJt5CIS5ubkrdjcM5fmz9oBRXFsRny+mNG7WxprYArsoTHn39M+sGH
fkELVXQASmfWnOjwUxdTm1oaJZ6KM1+T7lrpX3qN1K451rknwBZKjlLKwZvEGZRwwP9qFLOaPMnG
BCCwTY8YvRIKFLT9dZZUvCMd6r6BM5IR6Si4nqGC7uhvVgNPtHrTQ8UHvQ/Z0543wcR8xs2HPq7Z
gUN8zm6hAIc7O1aKMxeDQFJMApybuxVPeKb7PANHoTkB7xDNePnyA1C9yzadRE7OmhOEzWem8s4A
u5xM0pSxXI9T9PHNjSuvCQRgv4A/7RxJNzRlTsZmZSc3SVjVAG4y7cjhmC30KWtR2tWS/kK3+7kQ
rZpSmQjq4gOiGknCpj7x2oVAOI7vfkohpuxXpoNQgG3BV33EdyGAqAu+jXyqAhh0puo3gjhGhXep
zam9C2onCLpclv7snKwQw8FcTVmLJola12+cd9PO17pElz7MXwnnzj4qsfTZyamEsrZyrn6f0ArW
xLWETDsJK7hRHnbg/5MtXB78fGKuDh3LwZtXClcrdWDUBdI5oj+WM2xD/hzn48xigyEViVRiezUR
JGwRqE6Z6PDjSVJE3CIvlY1O3p1SXOo8Kp5kHh/sxRcCytC6I376yRELOKDjjuPyxnUfSXqbf/9r
clDY6yQNfjvICD5n6L7snfxvlZbxT1eeNW4Rkv+8cEwDRLaC/mJeydDjRx9AxpaqzQ9hhZyyT4Ko
cCDRhs1v94Lpi/s+LlEFm0wqxC4P3aStvwI5H7tz1A+DT25kA6S8l1MPVfnb+Bs2t6SsSEIajTKf
YbPhM8Wv2yDTJCZQCv7Ycxutl2wEU5i3v5pytptgCDPMzN8y35wp0MlMoR69/zrysukzqLuzj2yG
j8vT0nZobETAB/98PLhD1Y+kRlxfyjXYLzitOreb2Kl1eE6kDzZ23F5KhwEqH9hNEO8hxbTnkeEc
mYUkkz9JfFcacQF2CkRfSbeM6BvfjZgI57RpoF8i8Vo0uIe6bdEq3RUv0NdpXCyYRulgw8DVt3EX
ISbJOc20v7qNG3O9lFF00yEKAk3yiQZILSx/uf+JEAwx0ufTRDLn7qhU+ef1C3NW9NNx+R3E6XQJ
h3li/Wpw+0mLLoqQjL67XwcDZO26f8UdLyNzZi7pvrc6LJtzP4Q9DVvoFynEFBToQrWr0RzU3P4k
Qc+66d3NHr0j9FHUG0IaT24N3IjT3gpk+dDeTS8WkBfBTZ8MOdemkayifazglxMkExCcJ0aJAu+2
E6OUlAOO1tmhopGhVySM7BHvvRD+XJr0blNbi8PCjPkfUGLuVlxnTz7pJZVgcHsmrcouWPPet43Z
8oOcUO64A38aYwtQalW5MMQh7DlerEaF7WmwVN2WX2nZTXamILQ3WD+m7lUAmnxC1VCiGVSkxk6/
LqSl3M4tIHn1L2CeXbjV0Q6MnVhKhuPpWKAgNsjFL+f2ZcCS0SabRf/90bX/RURRQbXtTbHBtmqG
vKDExFMWdEDejMhj/AG2l6Ag1OK5BA9KknZlhsRjqyn0hbnVWucF/+npbdjMDYFcjugXOea+vcHm
lP695xHgzd05mZfr4/5hZScdqPlfQ2CYj0WNKNlsrFHWRi/97C4NqlDJE4HCFRTQI15Tf0+o33aM
UCrOG+FdP6xsfXtCQNkbJ0zqz70r/igxUpQPRW1deV+p4bSCD2CsbSmrPXVox7rMzDm2CoxuceUq
dsvvjELfgF+EnTsj4A34YzeV9dRIScgFWqJVVncp7WN7bgtxzafQJqWn1JBFtRgJQGGhli31b6l5
s6TS6J1atBM+wHjzP43Y8z2+eVvWUcUxvbi4Gnmb9ovVtl9Be7vVd+FjRKG3wUf+x081U+bLdzfw
NpRk/CaiKglevWxHH3LnI0GYdQCB3rs6MBghBV+aCTpCvsfsdAJOd0V9QNFLIw0bds+9QbEn6ewU
yYUhMvfivIOpisGoFDpb8/apSr0NQyFMKETI9nYvbH4wAkN+nvn4sQLN5469AtxcpYwdIrdFWXYP
UnG9RDV5z3APRlwGzV2ED6x/n62ojv5PGvh07ViD9wHLSQ5jDJBk0OlphbuyNZqP7NP4NzWC8teo
CT6LSrTLmfbvnFeWFvjQBEY+jWEtEpT1HgpdJjm2etwM1IFH8goSnMp+xwiF5HaXsV2NAH0m+Y88
t67WLNFXa1tU5S+jzH7z63a+OPttWvF1Mma0PLF1wwxxP7a8KfJbvsfGHZjJz7eZ5Jno7fhn2Dpo
6Xgt/6qETOZ11wgrQmuAKz+9AnVOZ8JdTV3FETpHum6+EXurBFcHFmDHMjNsCvjr13lhk2LfIuVs
Vai34Z5+14H2055Y6sjyZgo/GbqJfFwSe+eJYTR5djXifY2kXGqObsWd7iogpZ9a0dKpG3Ap5WYd
AHgC6TfuZ4FkGBYd/62O5SzeO6KDSGBcr/sOkGvBwpkLwHHZrArMVEhyfm5Gdmzru4rC94At6r+k
+Nqq8/EoreMpkxIyPkolxkKr9zGclngXC9b7ApUrJ7ZN6HprLHwf5rmqRBb2PAE9dluX493KAlZv
Fl6ozRDbH8vEtNrgIi/BqYDyOLnc6skFFoUxb2oZAuEguAVt09nXRPOJCzPTjCZJVi/ASJkvbR4i
+2dAsDCJwAhcUpXYcsAEr+dHqf8tucHNOdfoxIq5ll1TX1TlE/dRGuOd5EYj947p1QZqC3E1O7Jy
67DOMpeLyt7jzs7Hr7URU7DivV7Jt7MzqYrKGp70Ho5+PvuDFoi1wEjCKj9IuuJ5KfctyXjoA8HL
UnrSlFthb1rhxmWQ+p1JrqDJle0boTUu95diwXOS9Q/f66G0SLEojMr5Ge7tsSshNRoIXiRt+hBy
hrbQEI1gs9R/+VyGKKcJVBplkpieN66/wu30/8pN6h5TkE/89zy6Cad1of1js64f+EAuKnmkDirz
wi2Q/9SfcgEEwrTrcse4t4ZdYGV2bfK+tTp1jnpbqcsDB8GtUB82nk7lN2kEjABbJbIwB8/j2rUt
xlMOs0eKXfNa43gZEs4Y6DXu+A5gLhdD+VwhceL91Q4yyBRtJMNMHqhHAEhQQny7C7qL83LhGpqz
tRHF4G/EKvjIivNfRKSSS2Iq+GkcraLY13gh5eILPsN+P9UeIWFW6594PZXDUpwAc92gZz/FIUad
GqspoTxovHvD8YnjXyHPJQVgSpj0FXyBXA0HHMOGK8bLDJ9WWnwNT6Bph00fokY1IWpH+iZSatVq
SUMjOVuZ4ayTUVKa3RNXvHbkjIThKomES0lSsBhXc5TP1TUbC65eBqExHTLzCDLJQQ2qc9ECkXH+
3D8+Xhrhl77YxrJa7pfOj6FOE9FtqsjUahL8r4knYDch4izgNWTliX2eSusJ8YoC6quotPLv66QC
WmF5AFQonasArgeniiC3f9RWrQ4DfLvLtkv35cezNxJm90SH/z4XSCTU04rZLTdf2BQy2vB5Lflm
WLOf8nDohbyykQk0dWOjVQbuZEjXQ8OSFsjNmOCbOTmIB14OL3XZFiFbjsNdm8rO+6PT9L4W5gEz
4dSjuhbUzWbtsiO/cUEhp+Xh5A9mb94SgWABqjYkNvC1MXc+cmLQywbLl6/pcTTjuOMzSZYoy+B0
tfwZnLw9S1W2YyBRT56zHNBKlXLJ/rSLy8l3lix8yPJ7vWq3E3v7aYYSwPyLr8qeDHyBrR9yHSFm
4R8XsUNvJ9tI1Lnnv66q91kW1PBgsTlrctQKKXmv7nj1bAUvMQMFuvJhI2Y9NWNJ7oUKNwCsaJ3O
0P1VLImxJUoNRtC4qpvQUT71t4OEuZOqbRskfO2cQgU7xujf7FQUahtNCuQeJJXcjO9j57FmRtSA
QNWvAeWgQZ3ettQHPEHdKqu3ObSAWubbkhd7ZA+MfiEDQL0AVLK/WDtf2b+3nhffnyXaMZBrxBU7
lJXJAYqytBw4iGtoBXQKaFhmkatvTJ0v6kUa06gh1Do589wds7WM2HP8aMzlwrPtB/gZCYK42WiW
dSrl6BbmqsNSqgced4N9/iwE6VH0yFJ0QPZ1hm5Z003qhHPIRz03mHpbrteyjbCWqmBX3w8Dj/1E
mzpLDm9FWFhUkf1gkslDEqRBerYen0GRmdANXT/N/PiFkR3BUrPl49zZibzXlhPjGI70fYe+k0rn
wSwmy9TTJrJt2rTE9U50PPvjL2dlAYsCs970CWu9Z5xg+22hgu8TAt7qpxxHK50A4ARBMYEFQPX7
7qJPPHsI/yhEqRVxJ958M2Q6zMI1P2tG7dzTS6tgNF7IdLAEmLjQqOx6Wm4KGBw6YSxOCOWnqZ8W
uO1FHl84dfHSWlCHurQYrvQkfkT5Cozv1k7rqXncyFkiV35OkwOW6xdDVxa7kC5ZmTe252RU9aNc
RGPs8Nx0fxqHV3wqiXJvKvRC5hAYKKnfTIBhcDFLHRtqZajpZpiCaOJT7J8QzECH3TpW3DMCvQIC
jx6BBRdF/XLgjyHsoil8F0spz2uFzlCxd5WzULWICpeul28vT8PMPdamYTEVHKIcFGdXcB25CDk5
YW9mX317vGhEmMDtnlcFu73puQihALSxtBaT4IYHpLPvGBqsxaDppRP9yP6kM1OPuzPQ5bJGXgq0
ptxB0Z0LNlmxA+J8QHwUE4hZKczN+pAswIjsTzR4Rugffuc+z8E03gKMSXmNmoR6t6enejGbV7wc
U/Hr55cZA18SMZYA7Byzl1S5FmvOVVBTpnISzBy76YdnPvkCwe1VYnjQfTmxPehGsg6/BPZJx9R0
nGSJFA0yORR+nbspEgHqVA03ya8T/B9D3Ig1bXI28H3JyoKaKtIw0peGXJ4nvNnb3Gbh+dnqwRsW
0ILD2Bi6qhkLjKVCCKV4ZzsE1lw/CThqHDP4iUgLtef6QahYM7ZxIRinuO8aJQx22mJqTInckki7
/CkGuUZeov0vpy9aB4AcjWEECxn1fQ2QXuMxgYGPjkpU6oZ7UqtsnIyykESAkw8NPNoHK5/nG3Tf
UPehJoEmHBQXLmOb7d6bL0bry6+ST7akrzG5HNUvyo5rgZoefq0am4e9qeznw6ocZ95NaaDUvDI+
Jpi9HWpbUyXQGH2SHVfbOUyHiCEyQtoSPWCvjyDD8Ylhig+dnrKH2iPkSmbkBzd9Iek1rWHwu45t
L2/uBERExfuBrXf+xOyGfsNVc4FhbW72DzMy6l2+xvpRjSo1dDLlmQ2gVK658HYneR+FAEwgHr+2
nI2+L6KMO4dovDHCrq2YGDQGFuYkOqWBctPMxJlekqHDjaDVMffoloMM4PQ9LRANB//KkvSgIjiq
j+D6BFGzAjvJRZ+qRbamIKV3pwK1nISJIZ9lsiBglC0NiKlVmYaYF4EV156ayObaK2B9Dk8f6sK9
LU3Scr/FbCMX/PJ/dVvQ7lX0CuO5MuHQFLbmUfI7tA+j+owegHzB44Z2qZWv+ZfqxrBjRBFSaLCL
6BtAAajlagW5bn/tyGK6db2ZZ4T6UDK5jonA1sws2SpyhLCIbat9CdaPQqBXM3r6VZ4bke7xFJNc
nULAKmMNVL3cUeadfVGgnuU7S2T3mjjQswCoRjVxcI/xkCF5nH4DiSUmU86pwsHANTMPPblZtR4e
NC9IHgL/DHcBOWye7lIInin9SkTWID/RK1paWDqZEhyRalJvzeDxYfXGb36TAkw3JsWXrvVyras+
pcKcoE6FjoPSY2/V2dYWb9v5/t9C6nS2xVrmdPFIJT4WE4y2JAPiF2afkNV5Jhzf/lIVsY6eryMn
W6a2DiOzU34l14G1rcNnkxd25oOL33/FON8G5M9zvDJ7PsZxLLFjlksHmdOdBy2G3ye4b/CWg2J8
3swffMqyTYADnI15tY+Wth0BhNa6xI+xY0Ns95NRi3ju+UTy7DLsZWEAZLMrw358AM+IcdnestqZ
0O9j06sCIARPfNAlKiYUxF46+KciSqZQ3mwTPLJEKbAdFjaq5Dn/MH8l5uAtAK0saR2myfPfsI7y
ekQwiaI8IAcq4mk9Kwo4KIM7DFWJOImmG5eT5MuGy85ARHWavynv+tOYlW3TCeFXq19zj6x8eRkk
C9r7ZKwkv1ZqX2MAlyq22glzm68aB8bV6U9duhyNcsZIMmk6VryA1JikK9+7EI0I/GKIh1PaeCL9
IjGDxowopkfcdirmSVRQooLkXknbEsvByBgWTjZshgAH67AN5R7+KjHqmsIWrjTn0UNZf1/kAkyj
Z5OYazoM1BRsy0wIm4bY5qm0HYFaV64aINytQpiGgmZADZoZlQo1411hQsqURkHWXoOKHwhEmjFB
oq7KAmMWbbtYzToul5sw+yLal+6yaddfjiHkth/m1sw61Olw8un1W+5jbZ9uXaJNgbmy9L1vcUAK
8iklj7nt6KtpF2BCe8pv+jrVGEjGoJ+osqSG6masnPfEYRvNOgb1zG9VBYDL8680nwor/uwfAs4s
hP1Ub8Db3OBy3aba9c1tF4QAQ104i55H2GaQE7TcPUKp1p9zQWTkhDSTRTAOnusiZXHzHtTfAhK2
nPt7h53xhUSUYrVKEP+uQ/L56mUeyoeEnbLRcEGMDn5x+FBpI/z7tSbQXghX2T5Z9ufp3yOziRVo
GjAHaogM6d0DPkJUH52ZSaiEQzNP7KL7PWFrvxruHkGaNyg5tfKpry6XIQrCZTxDQpl5DflZju5k
sugtoHrxaCchVresrpxX2kb8+LeScF893SVwkV3YG3oYFIlrzq6ph6CxhmKr+UqbV+PeYIw2UFxN
izj6oPuM90ElhHonmM8s9h4P//z3703ofP+qtt1s9aex0tG5jLK4VLp6Vat18+Z64PgCXfOLNyw/
9OdyN6jRs6g5RQ7l3FWWE2Ki6B1r5TwFG7ht9KqIAstSN/ITFeUhecLkPlhvjHlv0uJz4CRAnen9
0klCAZXceEr3XZFXLQ/SXVmw/69TvXZNPGPDMQdRac0/J2lyPVeJmA4kRve9+cFEcZy0nW2AEsV3
lkGGKW0jodU6rdskfpZGlIV7oAa7b7/HWkvku9sJEkjNFxIR8WKthIMZa3OvPB3OgJHYOKsuNTMF
B7hvdh6trl9qTLjWvvvXx1bHPakBzII1CJacesWY6idCYSm526sIlCcKdiWU4wlcz+GOxQo34hJ0
z1liEbkddfYJ7UWRbNxc/ibiyJvlgivbRo0HR0lBkrz18n9W1WJu1PimM8ZR67RTsApC9U6MIkZA
u/dCVnZtkpJC1pcjaa7pujnVhlqqeO/FykKSXKkDuSpdOsB1oXKr8YYFHxUHAvbwOvcJdM8CcGSY
oOackLZuKOMyL8okGtcbcZje7m5jkiwph56pildEW2qLEdSaKg/CBosRXLyrdwp4/T8We6jwny8u
s8W6/cPjOtpxjVEov8yyxMYOBpzVznv7zr78X2vwNKGCJyse8+87Ur3ByLanvKgcuezZZ+WOhae0
nnR4NaKpeTrhGNEYl2zwLJQE9eTpuoVBBZ15QEwqCK5FykhJ87rKZfCbI/1AT5X0ekZSdkwyS3JU
xZzJhWmIl0Qwc75na1OYMA2uTBWxyr68kyAa09gEGHR8RIMhCfstitzwyx/1Bk51/LcLWvH2p0HM
vUJSGTt+UJ79Y+Kvvw0Ke6upLz0SWxxQs2IHe6CVFpzrIc9oTOh8GHMKzg5NZfPFxMkdQ042MltM
SVjZyLBSCDjjYwsB3SwX6+tHWCyNd/M+9uKknKT8o2zOTZkVSTX16lU+c/ndceaHp3EHypO/DULk
EkOLmK38TMGA6MPQcP4tm0zBTXLvu3hlUZE7qoLxVQh0GTzVyA7RuWnQufg8SLf0/eLvbLAnl4KS
sYglpwVrd/FRu5VLDoK4PrGR1eMTQSVn4xP6e6a5VOk0UY+5Wj/8BJSEuCKW7W95Fd7mw/MT98IP
Im3zVNLcWV+afRTSHeFfrgzMH2UsdRw49wD7DxadNtUzqonTI0+t7etGcGMmelCcvPCUfwJKCus8
xmrM+xo5ZPbHu5a3xXpl3LRl1mX7C8FV2rcDCNTs62xO+budr99xgNKaVunPrIGkdsCDXVx6tNAQ
1q2B+IOO1nL9hKghMF/fWWmqSVpogZBCSKEvXwfpiUuwDssQ7xGifdcOtAdP5QcmdwPJFw7d8i0I
F04v5Ust+scOInz6Sv/yFBcowzd8kn5+UXTy5jRt+liMwRNn3G8KS7bOl7pE4kE6nbRFE2cCLchR
67QlZSvyHsvm8qQeoNZkRiEkZLkQXVH8GSJjl//O6NoPEi+EBVcE+VLrBIx4cBZQKDaDAQoliiGW
HoiHORHCM3QTkjJRsBzgn8U9tJS2Lqc4UFy81Wl8F3y4XZWmc8OwnuUrGG5cSoUNO1P5OSIJRSV5
zjOp/vCxHSejCk3vcgQc+xgr75QPLkFgn7pZQfjrx4GLy7U2AoEUFLxeSVHaAB/4BrmA7Fy7rn/G
DafxkONk5l3qpcJWc+IQG05fhh6q1YxJPnBpdu/WUsoVFRk5iWQzzpnzVLAp6BhuRa6yaZBqVqCq
+CDe1MkClXyAVLhgWyYHFWqnOPEqRgdFevcZ+cgHv+6u+R8mgohOTOTivvCI5LjhL+vb7lOnSg5G
J9FLnJ/yugsnJFI7CwQsTwbzyMoxnCiTKZsExZ8G75utJqyo8CKD+D4LsD0EYHQ0U05nIdSzBhBp
E5S4qDEB2wVpY4iBVcnX5SuENT1XQRHT3X45twdSxsc3c0F1+YKidh6Q27q3wDUIeyAuJtg7OZ+f
Ew5DelMRgTrYGkSDDN0lmWKyXttp7IANUJe1Yz+zqeD5KBwFjWax1ZiYARobiL6UuUbnNvDWjhpq
W2D3U3+AzxN15baho1FqXt/if53MmEpIAjuEdy1kjEk1Kpr7XViYzqMILOU+sxPIlZnYP0WjBdCQ
9/MojPjpN6AwSh9HswTDnChpf7qSmAwNegOqn6I+kY8a+5OvAeoA+IPXmrCetu2VqYBjADXbeKvJ
fC52wMQsN4RqqQ0Z4REuCIS0YZzSpzxMhWqGcpaphSsrHQ4Bm3zv9uBXi3AEE0mJ+qXYGPAR8qjL
W6UE6G8SwAWHMBMwA7hZUiAAyXiNNqS44f3CTDZiUxK1JMh2rilEV6C1QLWzRlWZqPRoqDCxW77D
PG6XS5PxVXIWbZovGELyOmUKwMnNnP978fTMgyivoQiM3xRuuTzAl2HabIicX06JD4dwbEJwY4sV
bxiiGkq+vVhdBMFsWH1pUgSq7cY2CEDEB3ZweEYGtD+rKRMApdaGjPXgAaV380fltIdXzK49GMHY
Tk8di0WCjMcKp182kutjOs+FY+dMS62t3fc08oV9JLD6KUWl1VWXYmp7JL0Gl4zAmRpgHrsHVIUf
XJdeht6+tYByojBvqjvmyCHC2/PRROuMThAOYUOooygdRYTo/iDMsTHAiCwiZpcgsxdxxkMhrghz
bONi1bZ7lIh5YIpg8oOF9EXQfawK6WImhEAM9i5nEo3eXyCzyYXZt/LCyMB+Rfbg3iJkHQJEojS5
ekxFqT2H98ChJGWsnn3fwqp2LY9KVUfB/OQiKJ71FVwjS1AxP6iGNBy3MEqAuR/Du6xnIKcB9UB+
CnMWHXTfE9yej1QHtq3iUP60eaPGotUVQHAieDnTnu/UFB6MrNd07lObP4RHVqiCCj41tESi9TWL
XiqhwUg38tM1FFibOR3bSDslwL4HyLv8+H1L8/vJvDiu9wvnb7jnxZguXUh2N6K+cEpXg65uM+4H
gfe8PnMZ4liMQedfpQm+ZiijubnKDqaOybmYzw8L1kKchzjiZFuiYVUAQ/wpRpIy0W4SVqAmV1s8
k1oGINbNRg5I8uLHIxjY7gce4PCht+7N0Yp5XO98KgHCi67odtTowUFYpJUGj7M3OM4Ca9g4CX63
WOMIJi90V0iOcVv1Ajqkz8FhVWt3B7W4JBsoo3ezbNNnxlETM76L0D3eIkMVMv/0JDFvwMJNpyBF
Q+QjliMB7RsMVL4qkO60+BelzVtS9R1S3bpKhSa3Ys0H+xYF60mQzic3zT05lQKA6RFmQ9jvQaU8
Vf0p2xZiuxq97UBK+MxhdTNbDqv0/qeCSqyWcCxg38KdGlWf7/DDKXKhuYWophbCfozbET8ay65L
FkrRu5FEDz5DJL5t673Usxn0Z4qrSZa+rJv2xeXnCDayacy72s6Q/prBi9/l78S3hnqVIoZvRglZ
Igx0ZXxyJSB79m0o0Tbja2GmYMqnmFGtAhuAz28JEo9GqSOBpTRUgkkxrELD4XB4c4jGXMMbq9Hc
lYdzRcIJWsU3/NhouxtMw2Tmk/md4CSAILLWzOtJBRico1HTkCoUviI3X3O/xNkvWw7MQ8ASkXNN
7v1kyP2cHl/hzqe2Elmmj1XRce+/7zl2QS6Tuh4YlFiRfzxC39BItFPsVCrfz7+dcDf8ZdB3KAEE
ZDUNj1ivcl1AJqFVMv2VHQb9SRgE2Q4Yj1wvy8gtp23ZTRBwyWvYBRndAyUVJp08/6cK82nHNUVv
7cFNiOSiHo4IkGZau6HlensII9pyBwJbzgSrnIZTYMwH9u+j0p/Int/66yFttsISw7OXMVcLzG5J
6CCeaM+K9bnXHz27N27kQUDZJaCVyqaEO+GxnUEXaP0PGl6gDNSUVd2v/knSwcHIBEZLN9z1/cXU
bo08T0goG9csnQZqJMfHdPGNZBZlPvA/29OTPk1b1lObfMyGSvZIj2FbTN1DSRW1aVEZnmtf7fUh
htid6z9/JTdYoO4EHoPeiOp41Kp5JpCoWCMEgwXFWqcLBsZmtiUIVdG7DlHH6Zd9Np/+D+CnUesn
6QkGOPmpRbVpWlXG5ytVq2lbKBHhIdN6N3D41fBpBSUCPXuk2XXRjMo+xvsYvQukz7aDo11mHKpH
AYteNJv+CJHsUtAdzySbb7I0u3AUcsRpkEuJ7r798R0uCZCb60vKncF56VNl+f6aeEAnIae9RErw
fkB47OUkSIZ+M9D+U1VbBN+iVMluwoKY4yGdIb18QrLgH285UUmW0xkrLDS+YkBXB/Afa2/qMEu9
sZ7Llfz7JdKgMErs3ZHt6+0M6ax8h2f0umzyEb997RvfG9IMedGx+h298DYh8j8Og7FFBXLtUsEy
pMX649QDtsw/TYVIEWmn9l+Tw84iDZFRm7rVLqXFHDVN5QB/HVNNfeF7rpvl41ZLnOWNKv/BPn24
kFZFZi7r/9o0dSbPJlknnZ7GBhJqA6obVQa88IopRB1k+j8YwItA+XBrk5aNMtQPSbRVPINWbvEw
sfn8DDFrVmE0EoPh/9kwxBpAxMWm5avEhKn+bPYUDCeiILWCXpq1xWgYgJs2gHO1oTJW1eCtPkxa
jL9dXHJm/Bcg7P7R+KH8MVBFj6t1wVIwoSvWtOhZb+96Z9zdm6Q/YT78IaEt1Mj0YrulmhOaIJXb
rogvhjyyESR6BdSu0z/cn+UO5pNioR5FxPk8pnrcP1WgxqHAREquWqsKxaXueyeq6eTJq8Pm6ft/
tp9FiX58ZHjCzWluNXcH4pH4HZKQ03s66vskQjlInqRQT1PU47hDQGSkr2LPjFi44As++oj5iXom
JB6OeYThXMTQOaeByn/VmOgB8RHYzkp6Egca0E743gYHX16Exw5UBOoHns0UbBWu8feuHRdA78we
i50KXDZB30Tb3xtJXEMPDv00XtU1eGij+mlWZTeI/3rslTRJuINCwukVKOiNRAhs9Fpv4BzM9ljw
hz0eJsArfYPp3Xi60Qwe+5GuzRV7aqvbyZtgvZxWPnnnwFD8QhAbHt8YGJ6i6TOPsfzRs+oKApT5
Vk+lyqfwX1tK1Hca4F1NB1y2ENIAeFPZvsh6S8AhWxbxZSos9GxdTZSR94g4a9tacIIzFmXVaByv
jRGAVFrJ6wtWsJQAQom+ErnU0LdfU84Xzf4xTQX03UaoTHWqXD62U+i/J9AxLd7Syz/ufnssWakj
OcWEenfs23zax9Y2MNToeVV8g3/fvojGbhSbCIYYseiR3q2ncpay8TZdODMG2blKiKBPfeyK4wF7
2HMRkWAk5wq30cshVNnyZYTcZgvm1y0HA+nIbD1ADX+uUbkS0DcK1LZd0hAplZzBKMVec+sHTbaP
+2WnKs+3dvSmxpJPTa1Cqg3NX13qwkhOs8ZYk/wNFPpd4Y/FUPBAaur0C2Ob3AWnavZ2S3okc556
MQ14wi3TtF+x+XL8UXdpkyR1veD65nNwbp4eeKqk7SEsmygJUyIz/EygtdssWcYCp+W6N6n7L3Uk
Ha0JEDO9Sc5TIjgs8kgGa5jdB8Q34uzyhQfRVbI/X3I0SqQrGRXY2iRQpmtUC/UngR5i7xYcFHni
qooONZ5DofICJPZXseLRBhrRZXpY9mcJSn1NdM2xwRzNze9k9ar8ISXKC0QtisCnT4oXsXZVEfG1
l5nEudYzAAUWkjGt8NW/h1DX+J6jTxBa1gpdfC0DRCoM2hDp3MihJnEFw9yiCk9K9GV1bpXEVJ/n
0tKQIuAZh8xfP++DDjXLOal53o1Fl8iGSMLlyUrBl8tIXGaa67/IfI7gBhHGdEoMQW7KV/7zWFyg
feWsgP7GQYAW8QRvRygBukD0LumWPn8sRPxanrsutp9XxwpGozeLfpzt4KZZRFCf9r4RNCJLtrnR
6kFS7UIj6OlMYL+RKsMAZKE12Q5QJGOuhKdgJy/NFf9ADmYIoe+A46zv/dFCPCUCnhsx5Powa2Sk
N0s6Fwx0yGJLN0sn+a+Rw/jTKM9Vs7wTdjKSo67CVokXv90MV63hWprUAgL+Q61Fyy1wpDQIIRxS
GoAOo00xznOlAECXm1mAL2NyrqQq8HjN9qt/KvYa3+8GC72F2b6RRY8zJ7dfaAu7AKoQ9R+gnFky
oAYPsqKq/28IR5EmW02cpBdVhHykYvgOaO0dh1r+PGT3JUS/rULd9HNZsvond7SH+S2gV5cwkqPA
ibR683jmzGg39JgQd+IRS1Yo3UeKW7Ob7k+dhodG/nWosGX3DfVQlN9hnCBVB9sg7xiA9s5rkUi6
Bj8lRD+087vhTG3teMnO3uLWx+ZvNLRENG1dvGyn4/chQA18I/G6hhly4jXOooM736NYC9v5hFzY
xYS8CkakYvyAlCIeAEDHvX7EPlMjESmuVR9O/xdKy3LcFDNVg116c3vfPVf70fDsokwVsfmeFxqf
owsZZrNSeB4O2LpgDVG+i3IlST1rT7qxSRU7xupNb5so2UCjEtQ04YkpRfL0eBd+hmgkLo/4Pl74
RNXjIYZDZ04++wzwpzyaCyrsqk+tAbOkf/rORVWXCeURF73i/EpFerigOUJIEr0Tr8BPeEnDBU4k
gD7ehv4kAlEZfGxb/ZROZRhoEeZkMvuXuO4JizYpefmPHg5QGJSaG4xJ7aCKMMFT/3bpEDIDBl+P
mj6c9nE+06ghIHYLb8KdWElJfI82YqBiF/ctVby9XyCg4Y8XBaVT8Haa0zGntIIFn8mi2B5FkjI/
TaN7zPwxju5HjyXTn7rMo5zczsrebgCEZ1QC0ZM7SS83asGkTXR50Tp2Tk2jEVfa/T+iOcGd1sYi
bu5UFp7jt0NY1Mk6R/YVGsk+hKAtcbAFTdIkaXw+zxSKLNVzT1QTFwm/wZhllNT3SNENbjpRDsJK
6chyyVtyvwCi9H7yMGBh8L/oHcDitGt8TAImuscgNhmT1PQbEDIMv51w7mjJBiGyeuRzzK3gM7Go
u6SrDX7cT0sBiJNyONsSYHT8fYKb7W9avKhk8r2V5SPBJ37zmcszlA//0VLjpFsi7Vl5p/BqDvAa
phIu8mkdtCl2J+dJRnGAD5PCh5QeVgmT6TmWxpFjfUUOhF5lVUC6pQQZaJiRZPk7/S2C+ixibkF0
mH3ZMNCs5iLKZCFsU2z9Myk/p1u17buIm3w2A7fPPncMCp3dXQ+tnALLYTfM2NrMYudDhOh+vKDl
DnHGUa+7DGXAb+jztMEwMwUfVmQ/HK+o9/vfN03HjEoN2/A6zUH0mLbgEeirrpCt7AgV0UBtZo/B
RkwEqVLu4rVu8GQ8qLswtUj4ftspBtJhXRKKVlZvbl7MQipmqhM9l9UVPCkCI9EFGvc7lf/q50Zb
RTGVtQtLARjm5E/+neCkswR4wntEo2BwiawnwK0IhiwcBloX2apDVQ0hBkOVSYbX0hISVm7SlVF+
J+9kl2JjgT7kjecvzGPYbrySTtqFu5/2zLm1be+se86xYU7Aq6YDnrlXIyMNtQ+cEmAG4lo3DKSo
kDV0gDeCa2reYVB8eP/kl7+kVh1uKk8cb0/aHXNpq6gA2+VGeA8UtYJ8H5c575168q8Pe4xOLeGY
QpYcIIM/neOiunaUH8G9VcXkouiNJtks17xjniW5HoX1hyteiRSzM/nZ9FSktY/Yq7GITMiyMv5W
gAV3p44oUD3LvND6XzauwroWjCw9yYkhuH/isbJ7+RXXae6RlqzW3RNTOqG5UKhpJW32BFnG1Sdb
fPV9N4G4Tl2nI1hmhOzOPc1y0Z69qY7Xf9nOxzv3/N4rXaTAo4E2XhJiclXNs9K23upD8hpFAt29
2MS6WjRB+0KxF6143+OqYKVNf/wTWOBTMj+NnM78DgJ0oudbnXnLIUr804BBHevpKDQ3gsmTBxau
bF0hYUpYhSLMTsTYvFYa72JhysNe7r2UsAp8T/V5fU40P1JTPcwz+Tq+x7R2VS1kuWs70e0mAQ9i
R6rgXDyZsq5+veYtwGyHgsEGDx/N+AHfoK0fapI2IqdbOXuzwhHtssYi7WPWj/an7EwGdtewFU/M
J8NBZQDpNRvJQWVSY0+Ow/07qqezVH8UBCH6oDkwXYsUGkZpVJLqB54kIZ62WlNt25EQAdnO2Xhu
ab1/Gllq4LBBgUlycZli8v5IQg48/ZKcpyEMiX9ljEiEgb4Y+yCj5EmpgBY8xc4Gl2ihzayxfgCN
eeMrEPa48iYW4qWQaxupr3BDyXR7LnZ0bfVYtRDKEwYN63fzSc5QNRhZMuuuAPi37mkzq6YB/Dhk
ldPrFVqPU8Hkn9u7C8rnGtjjOq8D5z/y/ApkmzDQMU3EclusO/VFvOGtBTI7NZnEVgTiojjnZ9+C
ytpBiJSEWdfK+9hx6zD98S9Q9H38aPrg6gaeptffX98r9GF5VFF4jFu+u8tTauu4wNSuPxsWZaP2
MmVcnkdOv4ykQJBhbztfapdu2ateh97RWo5V1s7wUODBT1fiouDnTC/o3CvrjYtdi85S+IRwDTab
aMwV9eKk+iwtUfjTU/4nZWcy+NOiVCM5E9m4CGBpBOzqT/2lwZaMhzYngJ8q+DPuOTRoT+ID816p
xbqaI9peEXcpXTeLrJad20UNKAvE8ITskrNruN0Foku/lpPUckaYFCR0kOidjVlApKCc/lA2cltj
lgjnj5r12TeJ+szBsjDUSuscQz68/aXwMDe3zh/mKz0+H2VVxG2lPZOnUW1EbBgOydvG0r779soa
ClnrT7bepQaLqVWrzw/ON9drgY09R5Z7qSp2204lDqASx73d0yq0VC7vvZ/ovBNaYWgNX2IXWLix
5daKLGgIbnhJtap+YovGKg4GUG/8GN/tXUKeLCD3odKh9rabe+PczOME0ogaGHyBPBJs9pdXaqYN
epUTKQMaYcbMvHKR/OUQPtDoFc7AOHWvjh8VnI6nWftZXUzsyPIY6Tl6sB6ku59tE2Do4vwD50Y3
kNe6WivgEfVBtxK4DZ+ncvEgHJ56Loc0k2Eih+ofe8HFWynHrVascIWF3+W3B1LVhCIP0wjamoen
Zd+La4GUcr8jf4WLXKh0xCGnmb8HjVMEfqQE/FHhmGzJSh7SimVvn7uXfKLlOM708/ZmNsEGHrEH
NKu5oHCEnO14+uv2eBeQa0XKJNo5FeXI0kIfaIsnDtenAzbhppMf3Ehqz3zZ/Equ/iRoLrh6rQMY
kLxDSX1EkD4AJCgAPMBJ+FeMSrqlTqtUK2p+XhGaZ+V2zfnu1SYFZYCYJtOkMwhZ7uTS6OV4Uxuo
P6OZdzVBakS1yO4XZh/TCSDh0kYodjdHJMj/8P/8X5waJGmPMiy5vE+ZjjrR+RJZjZt+BY7Ng1h7
mEEjf0OeiRhfSs2rmqDzFebDBQ092j+IIA900YN16jyAAzLs/BHf0GqYsqA4cziUTm9FsL4HQGTM
od2Tfckxts0M10rL1d5tTmK6Qxuq02zJbsk4LivdyNmWhbOf4RDdrWJvOo6JVqkcrCnn+2kieCb0
tvsqGp6G0ZKgxAmB24EkC0GCQGqp/1tCOuPIesojkJ4gyj+Zv2G5PTJryadixXkfr+A/4sinv9bA
cDMCVidc/W03hzc1MwbfEesoobhNRyrFsy+8oe4Adbc9ZooM1Z6A0uW0PmXXcE93G0Uws4vdkr8I
phgAZ4/WB8I0Cbju+CqU6p7j0wQ04uVR1UcroJEQ7XlddNkXSq2i8gvPaPZbMunFYEJVvmMFxcGM
3OlvpLm1QKljh0gJG/p13qt4Plhp5wKHkWVg5BCZxnoUdbA/kBFxR8LWMzxJePGH7lCEAuJmppr3
0mdawLanTDNIuXX7WljsnHVjdpIrXpGtbeFY7lcGq6Clh83nD4K69MKFlm2C1XXM/uAs6Yy2eRJC
XekuFFBBGxqEA0HfS2CO1DP6Jc+KEtHHtwrqvk1wtuMLgWSu/C6rrvlz+8ypAkPMnQAbCe20v8of
M2b+DAHwSHbS/q/UP5jKmHEoQjsq/E/hkHY/bvl8j1KQ37k2F6xQEtP9ujgvug7K9SZzfHv7KOTV
a5egaRTqJB7YbNIO9VHqlerPJDmCYxQ4FK/k50yN3o1t98WFz6dSV3Gy2gsw4sJFrhaEGyWD+6Bx
4RHnO/ilOTTUlTlsQYgpQ2NT8e7SBL+YldjuNu+D3CiCPUhZCVktnRoL16ah9ljeCnFe0fDXpLzV
xc/tA6wNcUQo3P3sy+N94zoTVHL+XtDo7+R3fsYaFYQiAUR7EKubmTqB5bnFyrieLmhavRS/iUSg
Gr2CFuaOm7zQT/ETYdObCWIxCm9gf9fK1mr7EKg4GeTKmRCOaD4l0CxqhiwUNUi7DRubWXZXNPwb
VwtZs77+YBmHO2uqQ+nEEgaJhllgwmT8IggdM5TUNl55Nj6mx1jtgBlclhfYtZk4YgDjrmMpHYzt
kDzkGez59j0uW9HH68yybQ2bQ8bemTRiA6cwN8cgeswO/uMa9PF8DC3vWQMlBic+hVNPL5hXpNVr
PQUxjjIu/U6TVCB9vYdhaThBtG4tp/cdKzO3mjcBCSUKRn8fbSWlWvq6KQiiC1oGndmR+G79u4Ad
udJ/C747MydMxp0UKen6er/vgsJEK1+7Ws722zOxEoKwWNYinx/kXCM2GbJxd5jgWB/BIJisuiv9
HWEeH0mCrmmWG9CbtbjYdVAXDMU/EdzmzQBQ/c/vgtRaOAicJk+LHdXCipeI/FtuLtgp7SRIlvO8
GSHMYZ4diwXgFDOQXFN2eciKLkQuXpzmpAOH9TnhnauiUEq6G/ZtE2wQp6uA8pZyogHZqNksIxQ4
mt5tnv01n2KlqTDa1Umr92+spDVbya2G8MjCtrl8Lml0oOcoN7kyKLoel4eNhh82HYGTqeLiHz9B
qAlqsDM8Ow2CLswJ2ZsfrWXVs91Sk1lLo+KUQdMlTFYbn+D56ZXWsrC5nYBLrwx3lJT0ZsGsC1E9
wqIfzGeW/YUOwVvmAYFHKUJPEdwL5HncmN5dK75lZju4mUValU6cTpk43PF35b620JxWyFw2FkS7
7Kqx46vK4cbj7oaI5hnBqd0Nxa1k0JzXzwV2Fcx4PyKvgS5I4nVNLYdx/22PZYoJt8oA0K4Ic2Se
30mdh3E/n7q490i+TDpVer7pTR1ZPqtHHRyqoB6QAZ/7r+rQA72xFFo8xK/DSWyyxi2QzLGi9o8t
FntjqAfl/bdqS7Ul7SM2Z6zR5IBWQdo8KmjyhaQ75plBZgQgv+p7tNL6lYYLbRhoLPHCUKCH2Vqu
Nb77gAEPiPOiNbf7y5Cgph042etVJtkQirxEHaDfk5YNmvxmp52DbOZ1JamDgLn4l2fFnlfoXAuA
sy1ojozqroIvl0VsVYQdLxDFYvxN1zAjRXrcFPopEWl/Xzgn6kf+IVWJ2pX6hzsY4d4blNVy58Oe
nOaMga0Zj8KaieLeFsb72GmD8OqJXgD0r8nr0QhiXnVjWHOJC6FiHwf5WSqbNRddvF9k5Vex9vBn
GS0lK27iXL4DjBoGK8Ic8UBJVn6gL4n5aY3oIFi46s0feEh5ZS2iuSn0rn6GneDW8iwjWa9ml8Ds
jsJRu6hXPy4AdRnwgbC0HrssEMJ2Uik07KlBVej+JbZhuQALf/yzE5/tNxMlICymZ/xjiCpb4X52
iE59aUOPqJ6PbzWkmAGboOMyX8kmpD5TrJUEAldoCyqViqQLpT9v7N13/+t+nDvjTIQjiRKdQpb7
IP6RPueQJRbJEv5O+x0KgRGV5e3ngPC8pveC89m6tZjfQn+bLi46jG3MmQ8Ljog6J9YgpIaWRcNe
GYZAMJZr5pcaW6+Y9QUqKt4UOmlLgt9ccEIv8qJlTkYgMKvgpAFBqTHAOIr0PixqL8e1zeEWolJO
YckOnP4yrOyYdTLKMzWfr6KvffYzj7amZN1rlpaYKmjEUXUwM+EYwEBt8G/8GzHio9/Mt6gHQvlA
tYq/NYdW17sVMQK1TdRDBkblPebRZdEcD89YKueKaOZBEUQF2wPZtd/d4OTeJMdg+QejzChb9U4I
NTTe1GhEueUE6V/U+es+aQeYJ6StFqWv1Th0P/qlBGJz9VVWMmEjemMxbh+sxOITODVpga6V1P7I
f7EtWt+NLiaGxdIP2DzLG4YIowC2nZvsZqRQ2FrXb/5NWhmH9ARst3BnLQTRuzJk9Qh9gLZ9klx1
Is0xqXhauhssPG9L+l90zIXcgPasVhbHeAYhiWCO3e5uxS9f2iMasv8TjzjFbmOVar90HtvdcxdP
3lsc7RIK5GC3wtuP131LSGY214pUuAaykhIn0eTQkWGu+HUxnYXwQak5lmQ5/iv7p7QMHjyoH5Zv
xcG4AmoD9STXjDVOtQzG9+Nca+OfM/kwgQEF9GAyCqYxZjvXu6++xxaxVLb9UvlW+UXCmgWcaatF
Fk6Qud47WEBcdohYb9D32vCooACJdN+I/2AG8xdAlcC2uiXhaf5cXyWTHP1EsI+pKZ0XhJ879EvW
arYiFQ+oExs9tqN8j4IpOYyqX0bFA4xMwGgKg0kSBx97gr+fbiFG5Lnz8njz593eK0hSDsWm0yDw
nQ/crQ0N7J1LkO+Bm+kn4BZCJyQdRQbn9oIHwJ1QWlmkVCcmfLhKCx6w7t+gz+f3ZNSLX58slx/C
MaS8ThRj1Zgtwg1gBvnw/YEbXP5fdPsb2BL0vbXheMkoj1Z6fYBvEI8zkkkEMBfbsZKEme5ToqaR
PgPTIDQIVtAtBPE/qhNiW1uwW7LlZberNR9Wp/pvjuTV3WIQXDgt8yVKJFV7IMuzpGomvuDFenBE
DqFlL+ITiytdjaq1rY5RYh9wUAubtLH87IzQSZLckE0W+kyQ2ZZAmCnTDuRazAxWjQUrenrrtaZ6
pO2mXSfqgVf/dUluwVFwm84YV6/rz5vhOghYPWlbsmxxT3YzYNrXMFCZQvXSMUpwHt7sSr0RLPV3
EIn61xMhxVjmup7bg0TiaE7TwyzjFf1lmowXT878wcOU8RDi4Qca4b6U044JEBaR8Ri4d9NG7vKv
HzHUZiPa8NorLZQYt25buc4zeiTyo5/ELLYxUW9D0fv7dSC4s4rNaNDqG/eCKKSXotdNDwJgwDsa
ufU7Z/CxpuFjKVsQW+9OzMfz3asX+1Byn482SYiPWnzsXP+MjAJCJLTi4Tt8XbvBVkZ2GH40mujx
1doFOJczO3p3c3wHW3IXS4B/TxJ2CkUz2WU3AgcSwmQxoog54W5Xsk7wLLAMCvIC6tESNvlzn7NK
EcQmFH8hHWKYhA73UYj7+POiCoQb2FcyTiLd47IhuvVORn5BazqMrtv5lDVeOgtKl2v8Z3qGsGgI
1v4/lhCUY62TmII4yid8uVCgcXIwdDNEdruRgb6bpgU6jtSCHyLEyXfQbFTub558HinaEirU6BXD
W/zcUBmJ6JjZauLinoZ46nu3QG9bU5v0gbCT5m5Tk5Pa5IZxW2yz85WudkQm0PyLpDOSFcHkH1kV
vqNuUzAXjD3G/YgxM2YDbdIosH1srkNz6fRwf6h3FhDTKbsX7B+d9y572m44YzZVZgV6Fwf488VH
dBiWnhTz2jItN3MGM1quF8eyjBXFduqfCZno39aNz1u90TjSEfgxQ1lieVSkCP/ZZJLs/+e4Ti+M
3NoH0pc8ZWHH/f3Vl2WH4H32PMbA3QmexQsy0IP69TDwQyoUVe/W0PME/QbU1HVxgxjin1Fvqe2y
0d3FwdsqGn6CIqc+iIveAdX3Ol8CLzFr0qmAoosEHx9iaC5N5HxGsg97hYXRjeWmBQrXeneuDduq
ucFatII/45zyJ3SXoSetyG71TnVk8IfF2+ZW+TiKRImI1dEFkcttckE8BHjfrtzRMnUo5we2mYwG
nZvyAcRpvw7HiwEY0ES/6U3fp/o+0kXAgBwz1QI4xlWJALKMD4teb7xYjxW4r8ybCzOx+BNJNE78
oitOTf4ZqcQissGck3k+o2hmNtCXdKLtZ/ZAUIo+7buKmJCOH1UExo0gAIXCM+dFRO5GvA4ONuGM
3Opp6j3sbCYRRH+gEP1Kb+q5aHjo94YsV2NAipWfJNEPRbr3bAhWg6bmSlqlW00DNzAVzp2uglvG
Z8k47i6wudadIaVQGIjQO8qbvBa+yJ6YocPmour5WdUSuqL08S4VvVabKpGsU+YNCGoeg5I/Vqte
OeWj3oPRlMvF7iRdSS3GqWY3Bcrow60ixIogklAQSLjG1VdB2QSsvYEAgGTb564m/cHqkjYpi60U
5E3I8g3UkpIz4XRKoe3nXQ3dI3fQdL3GWFDV/+Le0NWsUy/KuO8HJ5qMxe9B55ikPd8UC1P6VyYw
2k9OOcWTzc7yvNbMpnAvADEzxIWh3nwrCFS/3cD28eNHk0NH2SxOkYIF2cWxO/VpwL+waUOfq6V+
RgYT0qj0py/gHNA6xIDwItbj8/FNmLLG7VbYjqB4oqB5oUN+qVeo5WHuM2+OUME84lynzMhKGkFp
bBFlMnICTEt5m+ztPC+i23n7XGsjmr1y4Ydwsn91cFyhWc2qYqLj6XyoQ0z7pj2wgsgLjd6zJFez
5Z9TwaMHbhCEC3CAk79u3PaRJRkRyUbKdg19RDLbySnnzGlRp57HCA6uSzZ1KvNxxSe3KzPczm2K
mt1XfYmFn7YbS1bYJpFPjZfNa2sPb/huqegiN6SMb5LCVqfRGV3NI9G+pEuwwYoYArd6YyIqhfFR
Vyn9+0C6XnUa41YOs0UISVrz2UqerRFXkigJNjhlQPN+yPdKZWSF5QmqBgBIF7NZiNCdfqx6ozWa
1TjUUi1ZvbPLOCcGMJkVPczzgQcSFnqgPoGaVAP1Ih2JuGollq8wPRxRzF5yD/X9kC34GTgMlg+x
VMP5ZJjZTuC9MShppcCTjTPssMuGjsPxME3ftljkVK3NmsdHHXlKlEc7+7v1oeBGqETC3vMqZoiL
M0HdBGnZuE1btxXbzDvQlWa3OBEc3Z4NPnZdgLUC6tcvxn13SwKGVhmlfOnQFs6YBYHGR2dPq1cY
ep7fsxgNFKBZL2w4T2vVbLVOdS47KQEn/KP6BQ3kgHqXO/lTb+ZUQG6Cz8UDzmcG64H2VW7r/67G
b8XRtCPskzmFWyP8wSJcE+xEHnyEKexKZdy+mwbxl4Xo+UWlDORLDzOwLen1gs0toS2cULlWcxUb
fzDrTPLFTqtl4VNYj342CkL81v/7mWcMjcvDw5kGNOVsbC7QQgFb04U4Thw+LEb2ESpopKHJpYTw
ATojXqFM0PUVUqky7+GcvLEn8v6JWdwwSM9JD/BRmZ2UBDVmt4VuaPIG7uSyHLfzGfE84MsO0toG
XPtZ6E8cvFBrdBdneLrKHXg5DGzs2k4IFFfjK+MHhelRUSD5crY5Q29opXs8aljcB4CFcR+P/pm0
/ZkSISm+jkcRRBoO3llgvzYz6v77eUmNf4t5K87TT2TKQJynAuYrZcm4c3R5kFismaamc5Hi2ago
UtmS3+d3vUVPalBWeqfC7UbQ3Vo96QuP+s9IXaUs1QkFGpAFBnQSNOMka9uv34IWLo4MScVnEixa
DSS4nKhLPrzOGColB0v39HyzaDvOXaMyNxVeOAwFU/2CirZXKaMagwF0jLy3GtBt4XCylVKSkSAX
rg16MXgeNmcVS854qO1Mvnm+tJYUK8NJgcUVnsCppOW8EcQIfeXRLmZcvfhbDH5BgE5t70Cmstdb
qkk1eKLg7TKzrwctfeV4iwqsmEAzzeQitzew3Y/nGGjE02g8FxBfFoct29i7PTOpAGaF4zLt9mJR
Htyhg6yTlOHEEuA30wEJti7m+626KZ6bIVsECIGjFW2o83D2ZGLj7GqR/yeDYgh5EHUrwXSVc+xp
n9NihcV9yeHrhhO46NH02UoSpPE4Mqa56qTDZMO/ncsFD3DWkPFQUF6nReTRBMgZkNUleF9sDSeK
9OjvQ0guCngLHGTdPH4WxWVmrQhFMl5oOcYqTfYvDGhEMdoaBL8oGazXlWWXlR2LUjvqPj4ajqaR
xPH8OtYPLtzsGT2gXyd0qfq/LiuHv108qsgA2+GQsRHNYosS9KTUByEpkalPyWvnVHntqAC0nK4W
eG4egZpc0a6XcswxaEMur0JKNXY/7YCyzyO6I+vMmQW1yPpuapD7WUXKJP4nslStqDPbx2niRY6K
/0Jd+qjwVomLWt9WgqEARtdVvYPPMfckVkTOwtKu/7a7bVQtYOOWwgQK2ZBDB6pfehvhLpCiLeuJ
HTOHoiBDEqbiH2mYy9GysPo5jQ/FsrSTiWAiY4Vxydr3m86phGX8GOd5roQ2mZkOUxT/lXGHU5X5
W4gR5fid06+dkJYfXxuiYcjVS2zcY7xJoN34jvvjGFJqw0v5QQu/chExo4kqB3hXbsNliBu4S7HU
K3sXPY4+MntB5CZRlm7b/BY3YRU9AatVo+Xr/PICbpRhiyEOjpZSpU5lQrR5sldmknFPygxBuc9t
mh6ZBi4cfvbTsHOa6UE0ss/RuTNB/eZwpuaOJUshcsGgPkaNQwCcOTurvTMxnK11ISrNM3xu1sau
W+2mNE2YKP/0K1VFdVzI3gHPhrrIMSAr71V6Zv+t6W9OFasraKX5UaxU5DveOi4frxP6ySIdWFVe
bHf5MG2ybLgbnSETARrhlU1ZwZe3PjsRbC3BuYa27HcHfBSnp63CQ6KP+HC+NMiFyDeYhzlhm/uP
W5Sd93krpnIsRAXs/jcqR8amKgzEoYE2dAD8Ar6ntU2Ztis0dxb1f3EX2Rn5S+JttZ5WWNVPW3Rf
Gji8Xm695s2LLLRQxLXAf0T3WOQeepKbeZnNVt0dLDLL5YoRxmv6LD69/IwYdHJ0+VLeKuAfg0At
VLPTtgOS8sIef0OYDNPXZm6IavvmS0xeByBxew7PlI2+L4GlrWf5A6wX6+Ekp6YtKybO+l2sGclZ
xoj8pNXCHesU2Z+qKehZ8bdON14XUTTTSPqjKmYj6amnD4OPorjA8L2Z+IBfTye7ZGVpNiUe3jRY
S7xJwhRlGGHAIlxFLEQgod4HH/KgKryHrQ+POSHrGSRnYCuX1TMXOSE4zckECzdd6O6rV7HZTrdP
dC0VciSXKXwBkyTbmB9EqscjaAr7XKwmpBO7JsLNmYBOrsgAHqMrpPMsy4ScuLCG8aE3f9kfKJqT
6YQ4YhlwHYZhb+hhPNCVrOoGp3Gs5gcZeTa1ZyjKlmLvtqqfUWXCwWxs2kOpEF59z13tCeQkmj5f
KjCbd2UShjOjWEfT8LFdA5xsTuy0QuxLc5ElZA6Xp7hQQwYsChXgEnNcO4zQWzIbhDPEL+Z2smbj
q63rGzmkZJX1wkol7L3CcVVoSzxeSZqMtsjFlpcQRW6kcvhAxtHWAI8J6ZXg09xYHYnIvx6WamY6
oE1SSEWBeLsFdC7l84H3ywW0ChEVp2o1QZddwFmxJl4IOuurfrsqLeL3lo0TUSdXEr1BiJMfEFOD
xet6NGLp/c4YhkiC4YzhulIk9k/cmH2GGAIcdhto/E/zWq32YTBt6H+9b6RTO8gr6T6hmCQYo1wh
fL3kjE+Lm3a0l9Fq/tpep+InDtloYYUHm0ijyw3OQKCwrbNkzXsR7roWNllpPUDUiVxQFYK9A82d
KYMXkchUqgjP2LqmbEpKY1pkLttVlsyujwCCLlTPqL2NpfNmHZ9kTTH0Dq0UxbrPx8StG3W10n/d
0djFV2BajEfKvZyUGmNQv0NEWfaH5Vbltq53++vRvikUGGSquVLZic4N7+50tCK177gTLTgOer05
f9ig1uy7/x51ci6V8PE/EnMF0u82YK9atz75Z26b+qsZoXcjqJXyomQt5DQgN7SFw/h3VdtVfcEb
juhNnNwgVgQjr6g7YDsPQxVL3REOoOJxViS7LB9kC6lArD9FmTacMt5JC7LqtM03P4o/VuO//wrc
cS0RXdwLo10IrBfOioqrcdRxg4p++O1i9rPsGsyTRNQCqe+rdDZ21KwOcrmRlK/TMLs7nUkFnyCf
NkDfwBGrP+dmRnF7y1znyyYDKvwmsfMQ2YrvHxOjvnk2YIJedAVGZFVnu1RfXVWyh68hXpnb+5GI
7+Av3uyTJDFwo4i9cI/yVJmi/yrCclAiKPuE6r+bwf9/e3FS4oqFbeNzrIBVBKYV67oqSuCmcbQp
pmw4OGCJmIpDAxV9leLiyCdHbvMc+8IVTeU6cxCeKJslQIK6+VxzAxGpvu/uBLFisJgn0vPebd7j
SQqb8c7u4WB5ljL5ZhAQ6sA50RA3yesT76iAS43QpvOH6sYpdiRmggyj9IZ5L28t1Yo3tOJiaiMc
JUvWmjz8Zu7BsZI+/Mgl0xQ5y+uTHJBc7bcbkodRmteGDDLgFM0I15jG2y2TEQCb8aRLUDsl0xdr
vtCl3qTA+Ney2Mf7wMQMUAtqvyWjyWXUFM9rnD0eUVBsNXI1mkxLlmYSmTzw9fh6NseXkR8Rfm1r
7xbmMRJyae8g3yibs4HQeutWc8PrDDrml/2C2LYFbzBD5Fk+0dnyfXVVlZlbA4G9FRNHCsB8wnkf
aftC/YmnbHAnQgwf1/84NoOUDYc8kLhpCp/eMdzi7aA4/T0AkcGekZGiwNqf9ndiWrg2+1e5gnx4
M6eW729V+duUMXd/07XC+fnEFVEmp4oLdVlyWgBQTkdTppd+WjSbvgzPkWFQTHweK3DzDpMbgOo2
HD3Zp/eLPM7qQtOvpcOFUswDX89pL8/ykkeJp3Io6nRV+2OsOc6SYPx5B17XBa0x6XX/PF0xGuhG
KOa0pRFt0dkrKbEa3UpbosLg4fWPRdo317iTuOmg0iQtXwY9qe+lO/pz4Ys7SjuuZnwGYkHmw6Bg
Yi7RXXGdVRDtCdIGrXKaPZOk6CwmLiFK7Q1hTh3YiluT34YDcJdCsadIZnubeG9zj1Tksx1Cr1JP
HFmM0HTpPic9g29+etcLSsPNoY4Q+netI6ddqqhuHFqz1BwR6pln2SDse65OgzRiOfHiR57/4+b5
e5MppNKWqSD42PnbFEmZNOEZ2xSh7jnNY/D5xRi58Jxu7ezRS5LY29IJzsRRT3/GZMp1liTSejiq
UX+t5h0nJnhz5H3RVHzKaKhrRHIXhW/W611SFYgvfWCiIAr2M+IH36UhuoPTWrrGg4JLh6+kK7tN
GRnVy1KIBZ8k5RhxUrzflLkTMdCZJRSNuBJ6QKftiEe64bDvawmjgaY5lxdPMR5PDxGXyGg0EWfO
jJS6r0SuuKZr/81qgVE6qS4iP1OAEKmyeFDae7rcgArw12uvJ4euNuk0l/s7x7z5AYj4C3f30/Hv
WocPG1P/8zEiGRO/gfjioH9E4CCMPNbnwHQvv1OqfSJAZztiG9iww8ZVQRLjGg6JkqkI7fDt5fqa
CvXmRfmpjPj/MrjEiU9fy36bKAhDcFEDtBzyTvY/inlnlc4Ebs3X6iLKALw2LpVoQd635wcmqJZt
HQfrjs6plzRAa6/UE5cRwKVfZY+nHPwYiFSX1FwMi8DXw9idYs+TTdevHE8cM4R1jCT2tOvjFoGm
FPb/nyP2BpPPxGhPM5SLtTt0M9KSAlkONuVKge3jE3nKLGd/ykNSkQVaBf3UyiZx2Un/qaIqFX7K
1e/tOcTAzTeQ2iVkstQUdq8tY9MNPuFuBbyYJ6U0kKUCQUHpOuZ5EpdGqI/tUhmf2ASEPfpVIEvE
VGTeNY6zsoriLOZr2KmOFp/+bveXIITFqDwT0Zzl/e9QTZEB9xUbML6K5ghQITvUxIjJnnFwPGkN
xYN0tJDSosVunevQ1zwaaaXG/pBUzNpr2ZrsbZcqL/7ZXe7gvrns4pWeL0qfQ9/MQV8ArOFwQktb
eVcO+OrkQ1YEwsiwcts3RCQlKTKyqwiZpzwAt2m6lxlLkey6UhDFDHwkYpVbLT8Cp406bSxhzZnr
fCDRKzbAKXobRu+69bpqIabxy0Bb07G8AsZsoVyevOk2wrlB4wnduAD7BPuodieKomeh2JXa7axn
630iGHMi+HWQI8TL+mQAUR7Eb2agq/Fk76bvhUuLo5U6QR2QwH7aPG1/rK+E+VZrt/K+Z8mxiAH3
+LYBo1scvhE6JJbTnj0LDRFg+KqN1OTWB0C8xahC2giZdiAoh92XLk6g6ltHUiQqSaD/4k5Tk3k2
TvgYFSocD+/DGr66EHJbxMcKTBquThKsFrN6qdk9WPrAezIon/BF6pSJb6hYVkkmX8YBWcUyPqlL
n1yN+LgMfEnlw50ZPJEL2SPqaQRvAGEDqdve5s5XoUgm2hBxV95Fr6zupt7lCtY2yK5G39a2jD2W
NsP+LH6rhQKFzMJmfE7EayK12PaVUkBym2R9abI6TbwxEOc0AkGSvPPE42O1Yq6GsMOuA9pE+dMh
7s60AUdMIgHKTtR9Bv2luO6JAQdiBB+MiFafUfdJrIIFMaBXehkbVl8mgTAXFzlTbpce1ont3hjc
c44GUwAZJJ0wS2foHGtcW3VuL5gAik0L6SFGr+wpgmogfNw3SuoZKqrMP7To1jMtbkQ2ZHBnwDx9
KsLzCSEIej/0/GPuWDYCQITw/X5UBuahDf5ZBPxCm1wISwECse1ykssY1dVDyT4ju3xJgPLQcwRG
iK6h3umc4dWtuw/MfoRsM0F1/XTAUPSa+wPOc7wJSJpaW2Ekn/BCsetDb/Bhi5iYRQmKk/Feid59
PMpbSdJeYwRubnfF2OPI7LLjkpUc3jL85dAoszRi9Z2VOypyVaemI8K/KyYJlXtCnJxJssMH9iri
9yA7rk7DogFoFrDVMhH8YFh0L6t03F3BwdwOpW2rHd3TSbyu5x7GywhBArnKa3yNxyCphaeh2Pqj
ot4iN2Bi1LzLgZM90TAdEnnbYuCozjO9cMjp4eYu2OUMam0D0vkTX16YKWEzpf6M5CgOxsPEuMmC
GpZtjmPi8ZekHluLgt0Zm3AStvqGdeU6ZXzYc8HuscPoHePFwmdPAM8+Q7b8mD7h6OlVdQKcOTkh
Q6OrTnoYbfXpIqIdKV9BXlTTUpy6QdgYZjFqFPS979OgVy6g9BViIRB299LZOiVho6gGVmNF3XAC
M467C7eHov93FdT8vVikTO564Gl/Y+KgkB6Y+DlGPI5dTwylXlzB9602v9E0RbQo5s0QRvSqLTRj
78Tf3MqXY549fr+Zaeo90pjUwcmVPpuP4L4tnr23GHsAED6lYN4E+E1+D1Lbuj8XI9tvBsfn+Qcp
LPxYZgxm2LPiqKcVyx5zxKTGQ0kAys+OHtTLUwP3rYNVPj4meCJ8Fzh5gbhaSjgf/7XLifP2JpPw
MgVbPxV7jeoDtnU6+mfq1WUZsQ4tsm2vpT1T0ydg6aRy3dJtiw21n2vx7AWSQcFoJkKz1wwfX3JB
/JmiM6JAfIRG7I+W4s90qWmHJ+9CJm4VvR7k9vinsmC5o8Loc0S0IPqaN8ilm0Id0seQnO/lnUbP
8WTJpLNASMOypEame8q9LspX1GH/wpbEvkIoBdyJ/IScr5VsgW1L4AbYBVhTyOXtq5GmR27lplZ7
CWX5+v7+LHoctLWlW0lktinNE3k3njddyXoKe2CzTrcHN+gDme+Zv+QtjijVjZOic0FYXFndJjwA
m1RVPIMzCACz7PtfKZj4ik2EPqWinU30Z8rzSqb2zuqijVbocEvD25R8glrUDZ4NIvtV6HXHRs3S
Xj/DCAsZXGbelYydlYoYZy1EbUEdecQkcAn0vE7A7z6wpI9VT6GImC7wInacycIDQGVOZQVuz+LZ
0K9NUWLQPZowiwgpfuEMx4v3o3nzCkxnVrYkTX9/KZNIocla4PA+1tN5237tTVD/HQZVKPHLHLVx
3HwVBjR81J8upUH/UhgAkeF7E4CWx51IAaliwyM2zO1DtHguNr+do/nXAZnaYY0feVBPDMQhr6Da
59VIt9lZ4mcA4cgauxEXm5ZLBBjDe+5AuXqE16jPVQB+V1pCb3w5vZydApCALX2zMQHG2Hb8IrB5
6s6thcMiit/xoFVIx2FchGMNsfDHF4Z9QMjlBqqtLGZIMaz9FjeC4RHwtWqllBw1kUKfATv7CbLb
R+HrHvhBD/BRtXIEuZDKYOp5Mi5QSL1VKu2WlRix+7GO+7tAfBX+9TMByxcgExW8xF61LHnpS6BA
N8nuUEqSyu2j4U5zuEl6wW1JhOfTThANyo+UbYMuh4m8pspvuw8eG7zbdvRdPXlsm76OeHOaB5/y
mA2ZFM93ZZR8zk9f6hWyCpp0tC+mMKxeItHhO4TEYNbGloEISIMZ8JxgJBgOv795iot/dleiuqSS
Y3VitD8z1KDj6OSHH/T2iDse4z/M030bUF8G5nK5GuYO+obsBhdWeDbPwiDJG0bO8O0o/IYAzPo4
N4f3ELxAJ9nT7S2nHyfiUb37j4IRysag3nib086cOsrGvqfk79w8NEtIAf+Cz1acnuwT7tblvhJ+
oTmx75XSgBMBfoqOtw9t56tBJt4CYpq4yumM4QGUewztpsW9pRqdIg84cPk6lrWcdMOhrCFkyVzZ
DmTQTGqSEIQUXGNGBU7xnDinrHCnVnaWeBvSKUKhgaPClXIlGxzlaJCJWkBOjg9pxMcd7CYU3EfT
RSD2rojB4YNSgLSamNDeZSjYRgvURNniXHLTR7lvcpSr00elbgaiSkNSdhqZrcv8U5MREj8RiVjH
KRbGQJHjgJvlEFiwQmee6IdXpwUIDNpHO6qW4jt4PA8BvHjKU58BnqMJ9W8ZNdTRsLThV3jJBCgN
0tb2fBYTLL80vrPelEpAO4Inh/mLuxZIHn+4Ue3sdWx4CBQ1yRZvGxrydXF/v0MLG4idXrdCKUra
58jobLA7d1kzWhe9NUAy4Rm6LMJYED/6xu29hS5QtrdthNZhOlmLDnA0JMLEz122PZoA/L7e9Fl+
2wdlvWM3eUlfpMDEVvFnpnGNlvv94d+GTy1YSxcxeNHHI+Mim+v8mSOpAYCHtg3l4TEbg+ITswdo
pN8fU3nSVx4ncNXlwRLxh8Y1YCTE50CvD13T6q/LAr72Bk3mIT5UAuF8+O1WBoCK+OqhwdLX2YSH
lVh5T9Ij2eFO2K/KGpM5GTVeKusnc8GGTt9J2NZfC9AICit5GiSF+zuY3nmMqV8mb9aqyVpqs0Mr
n8KW28aw0hax/Cx5p50ZXC09xqUTAVloSrepQa39W2KqZ04XSno5n+GiASx6OyVAoMK26mQ9yF7S
B2KDsarE0n0fyJgW8KVjtoqpz9WUltHPuruhcGag8Nu3qT6fZiMKIjuAB/JG/y8dEK2wqjtzm1VP
Pt9jZZqdFV3D5KcnImtBzEGZRYC5tUCCgopnIDYhT+mpJvqjEZ+mjDjrXBUuKB3DbtfA2bK28J92
pL503Y91Fbbj1ORXY5QnFYR4pmD6gteZH0MNiDaTdDZwxrAJP+xFZuzkvHQsgliDWiTpSAPQboux
U2hUanSUTBYANXt5A76jucoYwfhRhKEym1OmneJHC3EAe0kbSjzXZaD/KUgV5tVk6tcJOsSy1nE6
LVbqk2Gv8thotox+WuXFs5o+S6sF5vVqxREP0gn1PJC9iiKhHTgVwijyzGBW++kXsnimtc02rGHp
IDN6im2XN0qII6P/JjjIhuymJ75hgOjw6dJCg4BqWu82yoZU9yIiiyPUGvI3yHh3chKWpNBI3OJE
1sceNUtbyYtqdiFysNSyX8N+eCJM9qWyMvlIWIHWo4o42Hi0W89oo8Vlni7A1+RvRGC8yIL753Dt
ri4mpolFAEPkSAz//uYokLSOtZmp+6Nm3s9a4nTN6cZPhDxJkpOvBTPmffS44XXNFzN8xBaTn7jA
0wgR48++PYMOxMV7sMWsvTLBU3I7qo/R3921mhgloyBiUw+S+UG3JM8+47PtJ37xb2b/khiIt1W4
34mGUkwYO9optIyvEuhHWi8UTDvk3Fe1jjUka45ZBrivAf76nUDskwWiog4RuN0PqArsCw/ha4IM
yBcdPQDP8S2DZphABNNUC027l5UjLRZNl8x5jwirNpBzfjGzzZXbIZTw4sUHaihwvEWdEg6E1jTp
B9w4ClU5LdnXTZTwParFhyG20JfKAeb373Lv3uIKZxII6U5Rch71yOsBK2OwXw34Zw+ReLSiWeN4
FPyVTomA4qciUk3TpWQaJWTy5CuswFDbsSy4F0rjsEPFvkQcDYv3pilkGc0PiJm2/zfOuLTy6bjQ
ou7z+aJ4cgZ1EWEhXsPd0tonwEn0GkqBF9rVkw7Omliitrq4QVSS4s2ILc5ArQwki4qnD+R7gx6U
3qNx/v3SaRhlGA3hevwy9xMdWqznG5ZjCCa+h3WOc+TUmsZ+MDZzuDJPGs9Y759RDLtb9e8n8g3h
LUXTOCasrAhI/c5C6GtQ265EQ16DPlpkm8RWdvLQOt2RPH2A1MeB2exDNB2RafnPBI1RTk4M48J8
lhSHPLgBsAuFA2u2omATEzfV9vpYSe7gxaTnMujANiN1IPHaeslGsjhtPo98sXaYEkBIle7P3y9W
KiJE9/9Ldcr11Blxmv1ZV6p6qTkBViiaORzXL/aELCigvNXFrJZ8fwyyYP2viVUenFoTr5EMTLdr
sppJSGnMitVFVdFs2RiDELUYCTLS2XUplukObQiZNDw1jBgAz8DUU9zURCOQqALOjjRv2Vz+TD0p
jAylELGzMt+aNAadBtg2XrhyeZcalMu8HTBNj0VIPBkQ4CT4S/sJFz8PdFrw+3qJ5oJIDHdF61Gw
QKX6N1TssitST7u3uomyiPq4brZSw3jda660061u5m5RIuu/JLkt7bb4fQh/RU8p4TfqraXvPPZM
Vszt3JH3mOfMTeTGyZ19hvhKmA6+uRXlZPJFI6VYheuoEdX12gneV/A9SjyRyvGcaqItK262v64W
M8S/p6KQerpIE/GZEXoPisa/kCWgSnetlLsapN/2zBB3fhR6OYEqLVGRrIxPcDlzUl1wlBIIk/+z
q6K4EEfE3YD79VP/3OBpnmzWilSLp9kqu7q9qyc7WJLe2rQvj5qQnwEFOIQaIOeuzNcy3Su0uGXf
QeixZQavGma9wxRF8PrOcLbS2/cTXtteaa9ix5sDmAOb5oF2SwekwguZXnYss3NU/09AWW9GmdM0
PqZ+SHRfjZgSRnqE6StWDtqEr8s2/X3U3oB4faVK7SPAVCgJCK5V/GobHDETPhLjC9NOOM8FsEsl
zq6u6RCWwUa+jaVVOILjDmNJpJaQQ3Wwj4s9PE87CaFkxK1Z8AUXRnjvP0Glp9MB9PFvtz4lhCFY
eUxxx2cFiIy6I56CAzKe1/qE0vXLp6NimvgPyoiOBk/2GxFGW1dbLevWY1UbAqGHbxYiQ6r97mR/
ZFdN/0myoPCgp2h7zHqLm9dR3To37z2xg6obg/Rxi580fRoXIBN8aqubqcWyTswGvgc8J64Hi4gE
iXMbDqSXWin63cDeW2smMfP8kFmxiEC4Aq53z/f3iRm71THao50pm1jXBHKegjcO3Gdr6/ViZQQI
E0GJHqQu5P7E9Ejml18sNkFodoxSPtEaXRjop6MLEFCzjTWXEJ9hrD6K0uN92DRdD2aSU9gx//xk
XGXw3Fe591FmnY9MGPpNUg/LL15EHm65jGazzg1OsH1vk+xwx9j27/Bp37iiHvWo3laHnx82MJcq
jWkSOoa2133mMC5ODM29qKlia7dXM0oFf1PDWAWPQw/g2KbKO7IV+/IFAvqU/XqcXXlE9Rxc3f3V
UaseR6Yx9snJrjbVB2Af+m/jJrgvlCxPvQIfZQw+pzMDpNPC7wF9/3KuQUQSUWDKjcZVNVClmAoi
TZLKEi3eiT1Yt+pTz+21kQL/uJXZTVRTRCskQrNQWKsbrSA2CzfBSlGBjDpDAcs7EbCmicAshb+h
JpsKM/grUReCFdexy3y8VCnikXgoFJRgdAiWBycJ5SUbh+990C0XU35AKWMhPuN90+vJd3hbG8e9
rcEj3cDSB6yEy3o6XEskyiykoJAI2sxNBXrxktnFvZ2S/WbV+KF3+AnFJGLo6GkHS8hz0fnOZh09
1+Zyjh0ZCWp9uGN7V95PrK9ftm9SWv2BiSRURaxlx6HNRlXkQwvfZJ0Cpo6/wKkEGqw1Pxqa9Zmo
+Xalaltam5nqAtsffOKOvWUyCYXXlfpzXfF5FGfVHrB0oEdyjEHa1l3ZFgaeKyASkamN5FzDYGn1
tjxRuu4/K+EISRRfMv3P6Y2WUaAGVZCxO1stvF4nbMzz+2y84FynsLkIJtfOYAR+3Uq5N3bOfqYy
OFxBd7gQWjJDPUinTEQFmCaVv5g8HG5A2pRWMFHzpPuhlUPIE0f2Qcn2syM5q4/BlPknqB0Bm//Y
65mHjPZh4Jw9hkQvK5W8MENHuZYKsbeXrJXvFqsKEpFbGCkGswb6BRk6dfoWLXRlIAfKD6/YU8r6
ahotMHjMGwF8+JysbM868HCvzZPCpy6Sh5bA8hDG5UtlunzzWLEPO4skogLfltlhwsWqnMMssghX
cnF93LXPs77H+q8N3v0hi31hyVusnyIm6t1OsIpGeCvWebdFl6cE+Tk56TYsbuYdA/CLdTmNDzJG
DJfJMKldfGpGcBa6xanRGbh5+kuYbTYIfcvfhoYky66Y1r4zxXFEAG9UajtB+gRDrizghcVhS3oR
ysMtLuFWjZuS00T0NAoYPzcH+2DAAT4P0288woEHhB3RlqIfnSLCdIlEFRtvT0wPC3XcJWSJBHjm
I1zBcNzwAq/pR5PPGEL/IP/CJTyTPF9b9bo51XzwAIli7WyfZ29+E8J2OVDkuaW55cZ+9FbivN8g
XMCfz+FmXsJezHew+TD69bMqvcgUJzhQ4PBUWJFW5ZlSR5LsO+iEAdohFedQC2UJNH3daP9M/6HF
hV3kQrcfPB46YFcBYn879vFO9qKQEs6LH+FmYmz5qeXXEu5ZLKCAMIwtZuZYssqI0OrCHTLaKfw8
zW4UmUugfFajtGNnjt2w4H/CLPTOgRR9E25Wno9IBYLrw6L3SXMnddWHvJuzMWyzRLReczbH949Y
vvmIkCb++8ROzMFcXgzPRArHwFm9M6/wViywzu9VVglZoS/5ybbzaRrBJjbQxl+wMPmStkRsX/x6
ieltzoukSK2Xe6vpCWNAHQ+OeleP4YJl5KHCyvCdnHu+e5mdY/6GgOY4gesms/ipakKWy5+gPZsW
+8btw610TVKzXvpKrG4K+7mPxXzjRJcizJlrlkIUuPiV9R8+lReqjwhasvkuyaHe2jzOI1Z1MJBl
Z9VVWMo+o6IjMLYj2Bs4sCuBIevdiMB0YcryXPQQPNnJAo2vfIhgey2Tl14iEsHrJZWl84EPOzMt
O7vDmuUaagUY+YCffcKiQG/QWWsa0SKsGHopzETZVtVhupx387UGy0aWvT6jOBRC2f3jZnqIkbd/
reE+5PMkuWxZY/Eu2D+2Gm/vKsutgt15lJ+lBBo11hSsELn8pmJRxw13RzF7ZKCsu4lJM6DoDODj
Vq7FylW0WPbF/HiwxKEQktuOMVfgOxH5lgj1uOrncWTz6u6oZ3LjGEZU8OWdPMLqyjxToSaiRrm9
bKzRfH1FkfZZAH2hHb990PtbiFlO24npMDGyQ+1YIbSLP0SCwdQYQ8btDjW5mXUdfoJAzHk6qNEg
2YIzLKqNQWqP2i3oqKm3T0Qa8yCngh+VNBONk0sM/q0yeAbK9fLG0N1E7H1fNKuXXhrCmJQ2JxDS
Zy53Vf4K18Kc5f6sobI0uXcVFyTn3vNclj3AUjrF1IQLmOaNxS6uwYrn9iINEhmidIa25+kStCj5
ua8dxxuct5xBX1y88di3j46w9VcI3ADFEUwJ1nDyqly25bDow7vX6hA5D1xZx7aKev7HUvKhkGxh
HY+qZjMXb1WY95Ht6U5hGS0hM97WW/Pp9wZR5cld/yvkaCGVJGpge/JSCuNxTpafYOQJIvIkwfBb
yBglwgfhPUHYOYqiDlrRXEdBUWU0jc4MUkf5eYJgqFCvODnJrF5EaxO3FrmPJxh5ad1up+ktfKCt
O+Omk0Qes60t5K5JV5/RLL5U4rzokHl7GQx22TRspVBFJMG8Rxff+ZjymY+vVA/pNTbZoFvt2Hy+
oyYoyHo4YZ5ts0PpBaBPOIiX+UJ/qrOKfEiNiLmlD3l2I5rSQSCwWTelrXhxxwpN8UISnin2reRj
o73NIzrdn3J9FU5f42HgZvEgRQWazu1mU3M4KEU9xlnrPf8nNiWO+fz4B7Ka3r/EIQvdJ0Q5q0FX
5WzqXa/j7TWkvRlY6ZNd+zBw+e6e39S5gTJw2FNFBOWwt2FoVoG70BCoCTIFvAVwWtYtptG8nuZc
FErxSlB6YUF9epFxkf7lrUZpGAJOIUuART50C/Uwyw/mCfGLZXQHmWrFtqm0o8eA1hYyCo+i8d5B
RsO3fkyu3V3k5CJTGR81NRo6u/DR1ZFOf1BrGMA9jKTy7VODfCPmRy/KOL2mBj0yVpjBIhZmG8f+
jIxiqXBuDU3b8DVk+Vd+SZ07UyiqDkBE4bD7/9BL+krYz7lDc0TDvoWq71TdDCgwKU2sgeJ8fD31
7cEiJUGB/M5r0dzEfxWIDNt1QLAa/IXKsVtu8PhqB+g9Js6N5bGNRCJtiigwlXCDJ242SHk3MZ+f
3curYVK0peKom5ZdG12uncKdie7jne/yl+5v/eFX930oafdlgQkyubTA3IDoFO+NL6m0Q5Fap7Yv
+IrqvAXxJi37BlsRqKMy3ER6+42QIQUPWrB3UbdudykV2eLkdTjeg7UN1FofhVU3/quZa1xXssTK
APPFVRqb/Lwy9IRkSSAq2eUHqiZHpV8DjztGredAvrZgpWkEz0wHlSQjoPTnPHWaYxJl2JOpkHNO
ylwR0DtUfBciuCv7r8w5HubAu3Ki1iaO7TJC2rWdEV9t4Dby13Bn0gPgTSk4t95u1ytnd76Lmx9q
tLvyqMC/tQ6XOmVD2V+8clqrjdvWO/sn8PofpDB41P0wM9xsttQAZHnGILfwx6Sx7o7aaoxD6+fg
O/VPzmKMejgTisUaXeeHx6T4Q6XOgpCIHVXdkWBefWAfOO9iGAYwMh3lXUN4I2dQva+DJMQjootJ
ofGwblRfTk1pMqr76BVsvAx7SIu17Q+UBPOWLB93kzAWdssgTXd7vLqWUQ06S+QORqACGOa4nBh6
Op1czBG1OVIZPcBEQUyK6zM3WsdJ9ClB9xunsc44ixEYlKX1tx26UvRQX0hrt8cOMv5Lp88W7sor
9TSckMeOU2EQT8ToiatqdHHtpHMcAHwUsegEyC23uxdnx/zfgu4i+QgoqrJIGMOwDeZJgPV3arWD
WaHt/VsXmN0dSqGYcswKyhWY0m0he0hz6c1k0afO5snand7WVnMCBCL3vAtLZgmMj7OX9j153dJD
rNpPaBQM8/h3sv2NTaGgsRg7AK4Fz5lj+JAIf9V/vwCiMYLE52/raq66q7X0bc7Dbg8XP2NKho8W
FSJraOUOXqLmIq4Sj3d9Jh4Uf4L06HfZ7AvcZ5nPumNct+T5YWEec71GE5Ci3StEoPwohOkllKkA
wdnONy5XXthAd9/hrofTIDl4ehkrByJL8InDzM9QMrAG3YwKsClYfqo6T1mCm0HdgRgHvkU+oj/K
dTed/wGEnkcM4elXUkmVZ/20lI9/Kis/3hZZmEuIDgM9s9GPMzldZ5lvlX1WHas/BlJ6XEUOMy4V
fjrL11nAutomDIA5YSpQHx2W25Fs8Tv+K8sFk+4FFIJbqES23fTb5OsBQ3zxPt9b4kdIjbe6zwHC
icvZ3PQg1fw9JhB8f9uYjmKqw+FZQ82XkLozs6niXeGmD07Lppm9hLnSZAtJX8meRf8bUDKdtebH
tsAm8spm6sNPd05o3FU3XCZ6vh245kzGzfDYjUMoE5AA5mDAno33jL3mCbcgMNV5pk79q0qUw9fS
vH7hNOaQx5vj4kKQu4vuk4qyA9/kn6IbmoBaZTT/ouq2bkaIJV6YAsUbIeAnxt0xvAFRMOONz1+m
OP8sW1kxF65sKbG2B96IhPN1iQ7+vapJvTDQP9zHNa6nAqJ8vkCI2CThYpWqK0+oJNgxhOguhlL7
guEItKBoKW7QumVieeausXBWjv+KdkeTNmSUKi0Fk39o/d/9hpfrn9tisUhQ1Fg61c81rEhHGWIj
5JYE/Q0NzS/oMXOfGRJMeqbRes/f+o6Vh6xYTongcqi/8B7LUQs6YSCX7TnrWAvIrMaTQes2TNjo
pPUHc0hCRvq1Nchu/uBvAU9KSftisjXtS+LOeXk7lhrJtpbzTuzMJjf5SvLKD+2U9RwcKTwBGio5
xq/MdPT3TzxRsLxekYF7c5JUimsB8RYqTWeBf6BG0H78HUWzEXCemnaloKpUcK8Ljr5OCv+PMu7u
GHZNNnqH8JmXTg2oW0rjwmnUz/fqS71zCT69CwS/7i/QSPPWfibRzW+tFNx/pzBdNnOFy/ichkeh
5wxWoazp7aQctyPJQ+K3834esk+jHaaPlZ7K+757lrRdyhZbri+zDZm1DOZk+15KobdfeVbhvMqx
yHMUH69aEY8MQEeu+oAH7UxJc65MxQ46u3cYJ9YEKtPFAy6j+Nans/bwkbZgkN4+6SaH78PCDHgj
5+wtR+pUwW2M+o3eDt+wG2owOLd7VtDraG1nYf1tOsZejJzEG63170KnMJuJzAr12XbnGZDfXFiP
rt8iT2d9v9Ojz6gFB6ByRzUdEV5Y3n3EiqRZL/MVD2UF9mF2rkuBxigT4M8bntUBxrODcSwbMgKI
60qkwEYKTUeLmf48GSjAiio+cdvVjZsPqgC0KOX8PgAfdOYKa93LcX/viuCuojgyyeuRZmbq/fXQ
XsFsmIp793Z6ZRKoDK3oQAwVW4wnbCDt1Te7gvPH7ZdtBDyQuWnvLS7wYPKMg99nSpO9cX8pyvHt
6oBRDRg+4CmA97CAw9dSt7gXMNKwSbz7gYyPwVt+z1z32z1EGhPLrqupu2NDfCzh1ko1BiBiaVRO
90ESu604BA0xaNzW6uJ23noqqDrk6PoxUqdXK8P4jWRuGWTsuvHdsrT2+H6vIOen+2fxmytIF4Er
d4nN9UILMaUEDw6dBXG6zThCUehFC1NeRNrwxNP4I00J7mhZaMBBTg3gOga3Pq60EzDAnmbzb/Jk
GtLvHg3GBmR4NBGAqQvuVfkV7rHe51MAstaaU6cWs1ZSAavBg+4a/6DO0uOr6UMxU0c99TfrcXmu
eHD/QrUqGt9oz1QwYVkr96J6sDaGjhbNjjy/eQFGAkoe8EnsHHlR22GTUjjVl3md1lQw1WiDtODm
OEbiN0co4xdTnqPO8GejtBnFzPAa0QzVBP6toA9fzxZUUwP50W2LIwHTp11MnBhQa2p256VJVD81
+DZRyjkX9sR/GT9VwSkD2reb4b92aH5bS4jyoDtSKrojmzMOgm9ZATid5QAw2arffKOcGznKqII7
ekEmANPJrTYn6HWKn6yOiXt12w0oSffUXF0LrPVMs5iEIHhFsbrfRg/7JJLN4qwaP6RWql0y3Nk6
PtimNeV14hOVFtFgbYhIgkgwSPHiPUTnpHpimqAbCgcH0+ey3liEgweF76p7T0uiQ7e0mRoI28ec
+7eTsuTHarOAazO4pxoDVgJRALJBplV++CPnM7BHNFBbVynT61hVtilaqOo/HoXghRAHZEpo8qu9
0iJNlK+dPV+d5LWn7GhhvHh3Cugs9BsSMzRMJcG4UHYQokqqBL9cF7Xp3/pY1pVqrwzgrRqnyLok
dRQovFjEFCIHMX6wYEbh1gdfMxu2ts1/rM5bgu/bO8OZXnIl1LM6M9G8HPQTNI7TlY9rDL3NOCGl
wZSm3y74WPcSfdPet/SKQujVDb955MTawJ49edqmFyL2NcyeamxSmqiFW78dQyMeujrv4lhtcFem
vUrcdIReyA1YtaQDNAUKX8FXXG7dmIbmh+FhGANBppxTsutCM9h9ju4MYOPfHOfbVAz5zn0qm+vt
3KAgf4KAW/nbJuebZs+pGAIYYqjJi1aQVswzbxdx5QIMPrR+3TT9zsuGAzL5YMSbNWMc420uDi8z
p67bxmcUZ95aG+aDIwKh9Zcq2Zf3UuzTgxYmP20LbSqFnhtBibF6b/ehJ8G9QsmEscRrA5F7OD42
agC03/GImQwmUuqYwSueSHm/cEyBLnYzFtACkxjn/SyOdmoNkJDKgDv137n9p2CKvHF55ylXMMMn
kJvyYPuopy5mMugI7MxjfJS05mLlffufDonlN/8V/p6JIt1EkCw9/9fms59WN793Ii+W/LF0BLkx
+JllzuOzCdFH5K5SF5uewjqE6yXoWQ9mcZPjx88MIsNarKmrrvDSdJt3xXDFjqUvtbvjpZz6YNIk
PCSc0Up0Nyb+v5J0AB4Ews7PRlbgqf91y+iAYA/5MUTj1mv7SNeV0zJHyQkGFavjsW+7DxB5RmGb
QZml8d5q9bRbx2c9xCw4PQ6tMDKgqRJw359xXhVpIW59zOqwflsJQR2h1b4JGI4tEYR3cCg5pDyc
7eRmSDtRsOYb+ZDYfOTprsMoPa+r2teUqw+V/kKVx3t1X0LIJJDK6mAvOtGL0H8jTOXChPA16NFW
O8RyPrB4nok4vQtE5NF7DwqRZzxKdJKgypkg4ue6ZzuMvcMcWdS1LCCqPSejtJX/SyKQfkZXd58t
XvnjaecQqYdmVIERGdDKQOriXcNe7/Knh+Y3nZN6BWEd+kCFd9PgsC0rs665wkJdZ/jvljlhuLWp
r3kklIdp8gLH5eJSQ6LOB+sleuTuGca6tJK1ZfuKZVqPKJDfQKrSc0VTmA2HsFXxVE6qE0hY2mD2
yyADOev3tuApoVPayr78kqNu7hqhkB221TkEM2H0ix0kT62AS9ZAPoXUZSLvhoIegUZxOg+zr+5G
wlKHMQf7Qsnz8gQRufmAtdBeD6sQOqdsj7EaoJbv1Jr3ia19cVmJ7WlI8K9Gc2C6ro5xOEbPQp1z
oeBeoNkS+R9CRD9Z5K6Q9qkNsyjM0H/ibnYxUVEQnw3IG//+e/m9we8vDqGl6P0AKID5c9r4Ya6V
r2o26mJlXq24MWpyXYbEaPpfGhH4Ggax44WW+K4htB5kBJtU0HJf5mNgGpLTl6RvZNOEVAot7wgk
OwjHuIl5Iou1donfLqOzHfwAkyT6gsIxLsrgRzwX2jqfZJuW56evsu6JizsU9GT8nVcPM2Cx3LRq
hI2v42Q6uJCVdMIYbP3gi/SRx0akO9wsF4ZUEsHNjo91pzbZFLibMrvqWeZ4h/fJDI/WT6RKR5Qv
XqNmdsdZtAnONI43amLf3MSuuh30ohPlmA0KNY5wfDlSm79xpvsc9+78d9Jt42yz4dmhuisreyaU
CQ1Hiskhrpn24Av/SyAC6mRnsuHho6ail739d7s1wC+9EOF968TqytXw2IMYcJ6yDjg5pHDdDuYy
iXorJTYIr7GPqy1ASPEpBZ4OQOv36SHPqnRlPUYS5Q/PlgQ4EZ3sekJ73CNYid/ZndymfCDG7g6H
P2x/DjEzHhp2tf1MhmHdQfiGl/o0/7BHIjH8AbEMShnFw2S1/zRU1OMlpPhrY26pHk/JCFAXHmSv
O+8U0zALYIodjgG228WD2W2uJlScxSm25y1dK1MBIwlGP8bikWpH54KcO/xZgCyIwtUY9v4SMelm
wM+fTFwVswzFOazQNgowBS5LSxCOv5RMT99r+t1O9JcWAd/8deykvRaAFHaP+vtUFMjEKdeVLruy
psEeBjHc/+Zmauf0kodnKP+QCvAAy5zdfuYqE0u9i3vakaohWVbv0WU0zTljGcQpGY/EOb/NfoAR
GFmr0hb8iH9XYpmMAtppxAnv7c4ccleELfmB5w+6nGlnhNXv89msB1oYIimIn6CKPQ/etM6nCSI6
rGYHRy2/iM3nmkNy0xIp3G+PInR3+rj3/YizWdEtaw0UhQX0N/nskr/FgFyE131Wz7xM/KMNTqvo
v7lJtEkIihtbv7uJdyhlCUHnHTy7rzE9xjdTR0LcrWLC5+DVIsAJxyC9UVfxQmRCcrb7v7JIE+PG
aQqONLtdUowRaWK9YGbzyip8GV+ohYezOroOvYlqvslbXtey1EEkLr8uonMnCLNyoptthA3Y2qDv
n7NcN0/ppuK7YSoiF1Qig4oPri1kYhdhuPc0WmNubqxlNQNNuT3EbIJ07jbgsUzbsH6+4ylqbb8T
WS5JIVcYBuONp6YoNRdCvYRgS8nhxzLBLIv/5jLqihsJNrH1sv61B7NiC1T+PwnCt4I1j53dhZSU
3XfnuuQaZiicoj0JFOsMUoliY0oA9OS19Y02FSrflupvdxkcBJqXnF/qhRYEC6TMJ1HqZolgazXY
9QpxQWFO/KL5OndB8HKfUgD3KC9+3coV2wiNEdd4Rz3w3RdConKg9H3LyDiMGzC6Ej3ZQDr8weAn
c+z71BgItY13uOFLxJCRogITs01aaOSngH1B1kbJwDmoFPFylKzX9TaCaJTXG12VmXd9B04dFraG
tOOYl8h+O65JcMgwf4tTimPc9Z77NncHz+ynXsQrPozsBls1r+2WgDRdpPYYNjXyZZkKBFiTC0KP
EwjimGlKhNysg5FOtlKEwaa5pXudyTCNUJG6MVUd9SGZ6jMb0GYpyDyd5ZRLmoG8pD7fk5O71lAj
shSrtV+fDHAJtw9X6SvgSnEeZkCY1m2mon//Ag3LeHWXpRwnD103E6PdLitJ0GrTsUMvsmWrVkuC
3+ZiinvD8X8eYZQPGdCh9U2YdlKdv9H0Yjjdq0GP7S0NwLeaOzZePTT4F3I8qKmkUxa7S3BFAjoq
MRmAik/+ADKG5XF4zxZY1XEKRWsEttQ8LW3qFvCu2enuJqD5OgYFFOqAgEQrTTTJHY1vxPYyqjS0
pQ1bH80E8ehi03p+yxdWZc7ZV4jg0MQNTzDjae/cAieBHUFUYRiTLn2oh2N7E1Me65+C0MUK3rFv
LSfzcR6M9Wj93/YVZZAlcngPTrAyJvWj3E6ePkcGtqhBPgW5FDGK9FDF0S3iq+9kLaGrrmgyGtAQ
fqU//CG1LxF1/DdfFbIpm1CmmH8zLliiz3Y5BgnIH6sPtg+y0tTNUjU9VLkbTK6VCunmN9i2TBgz
McCenzYSjltmZYAuA+iTK7ByFc3/7sq2irBoA6E93Wd4LYUEttZ4nSmTZE1KmmND9raQTM1bKhXt
yr/AcKnXGxRhZv4TJHYv4QXyxfW+sJ4WQ0XGmfj7FNMK04WUTo1EelLLXJZOj03G6ieeqlqg5gm+
ePI+jmagK6qJO2P+NQemxk5tx/MTrC4ClcQ4bJt2Ae5PsPpncUG2nXWHeKBeQemhq5XI1L4js4mW
n9+HJU3YZrCHbAHKs7xYOJCBi2Fz3UQFkdU9kTZlfoEyQbAyZ4GRhYX+HU673oJSlDdnUyOiptFA
iIk3U/gf8DhnBweuAFIL6B0abXVJAvZU64FLIT1RsQRwKlCuR26YiTdbWMLuRfyVKjO7ViE2eyet
r2xrCr3UtZw5Gy6TdbMARpGScHo34PJAUB1kkyv3uMYezrmyhyER7vx+uClVQ7aQ9W7VhSMqutuz
J8JTLemokY3b+dZ9G5QA9GMiZHuydxH82Dz9sWMpv0Hsy/cF5qv8PJNcNDlDKduDzPOFdHDvtMK6
YOeY5TBFhGvEF0WujkJeLjJ06MpV/mHGeTz8gOFn+W7yZ+Vr6P4TivCBZW6stVYaweyzSvZLbN6p
WX9XG2ilXaXJRBuYqGGCFjx4sCUxdPi09hGtxPykX5WN7QL1GfxDknpCyn51DDqsNzVlUdIBOKtx
OG2D0ELQIsOPbCAoidTMx90Hmb24lJexldUDhHaA8tcVQzmrCBXam8FipBkL8ZseqYAmlQ4v3FnH
gWXRI3Rx7wUzWjUeuKeCs+Dw4MyPZfwUNhFvteYewTl7EA1nx69WWAucHf3dK7ofozqgrcgnDcsO
d5mVjjN6Fqp1cNUk6efjJiMBAJe5bE704SvXpVBWtycp21UPykx8xxmDpJN59UJSv8yJMF2DubPd
tyJ09lwcET/ffB+yd9s6wsixRdQLWqmz2/urrL5p1T/sDVGkjUUAXpD4SNEqm56w0XbP7KGwwaYi
qyBH4FOgJckI/TjT9vIaHU2AJrK2JJ8UpZFT+0BlGsAvKLiksYD5ZCIFvyo5BMQhk+/Qi4zqGj5l
cZMmbp1oDWIel+5Ie6XE55hnR21XUyPsPwI6GHFTZ5Y4ZqR5TykTUVNJdGYOwBFJxmxNnxUg1w2E
4SPsO+dhPdap69O2V6W9dwDMi1EAfNW+PQCOoqZ52EuHDUUNVP52yQxvCk1pNrSiZCVHq78LnVLH
ZxXFQhTTs5VR8xWlVeohxS4LYaUB2s4gUfgHS74NGrGIJvqk2uZog1eE7sNRwfisHYr3fMMoKaZR
f0eNX9bDDDWH495p3HF5trHMnorX1x4Fj/YSqNxfl5oeqSXG52ZNls/oEYqpq39WnkgfAHsTdYT7
RnB1hUgq+7MI06YF8nnN6A0YAloGSD1/UMEAJwjYGqfApfAtC4U2gdiHJpqTUFnCFHMbqCM1jOUH
FrIq4MnIlNPyxi6valWm2aI+LQwepcF6+pdwPIV0YIf90kbu/7tqMRgO6TWsoL/cZbNeMTZyNvO/
s/ihgQvIOXCSz4Q+ZAd/2fZxW2OxpWHDw6SpMpdwU2FqUGJwv7ufipgGTU4jnC3LMEHuFw+SqHf8
dutS5sDiQJoRRfBbancRXr+36LBwwQygjb8mq5jfu5OJs+vrSnU+xdnVV3x9pLy/nGcergobRrDb
rZgMvGUgAhQewnowF73oxmZ+2iTvvWwMJAhfimBCe5Y1aSTKJTtIadRhm8XpfAMm4atiq/LoYqer
oGXBbjRRVvvhVQqnnUvjVPvoC+LQ9FuLgfM1SG7Lzt+cMw3w8rpbOknDyOl2Yx7OicWW+MD5O7+/
qgh1Vt8lWSsDgtKMhrEZqV4ddNAQifnqgKsMIFYHR0ZG/xIE2BB6SP4FfknqecmFRkHQGGenm1vG
4ASr0eN7NhkmMVhXDZXAkpBXNUHxtbGCzgwZ+7hPOEf6VFC9hLIyoGuQXfnVlHtzWX0cVfZBvqd2
HAB5mTSytpBv8ASIXYMJqkac4FgW4gIzooOF4wlevTVhZi/LQ0AZ35drDhHb8w6k2RwiBgZpustC
FRuve5VcLcgbdYYntN5zYDlpQd82pWTLp+J1yaxDIOAb9KsYtBCbhB24kvbLNGRfOTjQjK2BPBsA
9cZwlmhgGFuV1YLza22PA+TE+soR7DIaUZJ0Iw6mc5+Z5oDhlUoug+RpVZ+tgtMRBudWkxrZz5bT
N//7diK9Lcq3J65EzbCedPZ1C7kxvI1S0Hy7tGL+FGwUqmIhxGuyVl6XkQFJQnq7FnDsqOjNc40i
2zaZjaxUudU/iiitb9HHIB9UDGfcU/JO8Hw4mMYRAWYJ9ZB0gwSidxusgVpFvNyuUIfaKfZemivd
NQ0xV/10neWCrM1lkzjmlVbjaTL/msHHODLvdqovT4CFvsVhLdcVmdx91rIoB9waQoBk70J3sZMG
drIvRQ5nvkywbod5/jz5lStdUiWKMnpgxDsHN+z4de8BVk4OzcSo9BooDsu2mGK0q8POOqBThloA
J4aA907OsYk1o3XcA7IcyEuSSYBeGi75SqNAAuFhoBbshurAMsTtGHWEKIBO1HXtq5dp8u5gXJ/8
dT8auWLpTxrDvnA6leJUOKJYYXGkz96boInlqNzpOrExc+q/Msf3AZo+2Dp12nbJPimiPNucfCKa
cvjWaKklBoNabxusRsOH6NT0mKsbzBTMGWShCPfZJZK2vu6nb1BII75omEcEU6y2HxA4odSJEycA
Sz7ZUCac353ti13vHU5QW87I+zX94qJk4ytE+BPOZ86jfy3bRpdqApGNfdNLQibm2WdG1bHzKxQ9
03NelGgMFTn/IESxT7u/F3prDXVDaqJGcXMIX0nRqn8xLwV8nmWEle2+/x1mo6I44AGh9oEBwXqc
DJ0UboheY4oOu7JCF1YWw3O60KZ+JmxDwgU8BZASNLO1HdqB1jhWyeCP3xVCp7Cgl3KCSGEKM2L8
8r/R8qrv02mZzSEmHdl32sGl+idv0av51pgZsdRRTit0+1xue7qvOlftiBWI/5EayNBOkt0cVV7L
z+epPJA7lGl5/pHZUDzt8qJH9AAlKZkdBpu9YXZi+BGMpMdl7ZyvhXgYV7xJx84zjEkVOZJ+UiJQ
9+PSN8UjDGrZ/XA+bBwb3GYjmJEBk9qgBHNhLG0+/PlyIw2AtJDxWfbX2ntgozR/LGGI6bBZNbgR
0olceszXgCkvlJiSlOEyQZPH4MLH/1N3r1g/o8DHnj/kjb9/uSns8ebrllbALbBXjzyAy84PJ7j9
srjeK5g7Qiq98W15m4LQ00nTKLb6EbC+OSI2UB9STaSJThU7fowPSD7saOA+/hM+Mm75qkHEgX3M
auL0G4AsXrRwEBOWgikqGEWx7cIsbbXzwKZEQqV7yiuANNeXFt9Ghj5R3OvoxOzikkUOBs24lsIB
gqad2GijU0iVZcjiEAyCjeeIyqyczQbVDTq8CNCrHYvg+/9trUclI6Wjdxpltt/20e63tDLzAHau
DWZq2J9ttrFHNccHw1aqTQwu41qutR7AL2aTWofVtBrbmZ9uUSWoPoiJhrmsm1R0lYwXp0VniZHk
ni81+YqrfNcgIWP9Xt6Mj7IRAFe0/+6apkAZQ0ehbvE9wqwHBTmOFo/kM1H/MEmQ5HqDAZni1siJ
aSnZdKsyS6jP7LmgKS9R5zAh3Ky1YYE9i5thFUm1Jizoj2+qfWYeHhehLJyhidFCVdjOqOagzlWd
oLn9DcTWS50rCy8JI7dQejrWWtAASsLQOKBa/l+ygAT0bt2rQzl1RRrg0q+EwqpIaeMcfaN7MPSq
QDg6vUxpzJRvatqr2a8TdvD6nOjjf5SLVU648mkKFLpNJm/2TFRT2tKuqix5P+fvEdv146w9RTrG
9MYBannQMc6uhyeQxluWPo3Hz+gxpVLKiiJJfo90A+/4VbhCpHoeUPG4fuwKPz678E8IxbMTHlcA
v1tnpMhEtbUQoJAppT4GiBCFcamPTbB94u+WnhXi86J1mJz/ggCfSOQB+FxdMpN8sYTrESBKR6lV
3E0Um4eQHotpdWqEy8NexN/3L4+bubBGOPI54EcU8FZ5Y5RrkGpR93FaRvnWdLANqfTu1pFm+j9A
6HV54VPq35LTDiRNDifqVpkhf01UhFOvX+ln1X7DnusDC+PaM1fDI1dm/0jA60kfknq/mr+1E1v8
z8txJ8mjFk5DdlXPpfNv15ySXDZcIWYL/6BuTG7LWT4RTAaSYuzi5SseU3hQ/bVIS9gj3F/Yg6xz
UjfjQGkAJ79wJMmFCb5Qt1k64djR2R7KNG2bm1F3r9jJFp8CwkrPcRwzo+R7j4TgixbHOrKAeiQF
u9zegsq/8gq+u/6YiM6FTBCHHnPahGL/whksVkz5FmVyfGPPfL4ail0OCQKrx65W7e+/wTNVB54J
TW15yrUtt0kr9UZ6Y50XOYGMbF2SYOrvJjdO8R31vXNLuQCeHsZNzrECTT5ldNwwJOrwh3Qdt+o0
6xLRBJPGR0AQutLpi6Nfn7DXmDOsCeWlncjJ582Pnf8/hR6ZCmmfdOWeQLOxjFQDj4t0CjIWLqxx
ASllaM+XN0Pa/kWzZrPFAEqJgarbh0dz9oydJxXPqHQWok6eoOf1y0zAfk3gLL/OYwO9+P9+bytq
IUbq7mSYXU3hmddBDeTeuD9PIS2eg8RuDU1+6V8wzGDuqAxmNcL5SSAHKELIWuNIz6c8O39+FuZQ
hfDWKLedk+07Zwj/IaktFOkbwsuGzS8y4YYzF9/bx2oNY+7mCUeMjW1lGdu77QuDLJ5/wzUuX/mC
bgNPuB9BCs8CRQzsdOD8WqFkK3Su4t0JsbzS1LdZ3+zjYo1RfMmYg7Pt53ECaUzF91P0LqB2K1Q6
HQVmYsXGBXj81aEhUlI0l7A0iOLWR6JK6bq7F5lwI/OwxaND7eqd96E2ghLySWnj7Orv75Zli8v7
Mc2C5SZtzJr7876ZbDoEUT3Mxi2gspz4op+bu2K/WAOSZUaNIi4uK3x4Zg1XSDsyKoH6g0bbPiDU
nuOUL21nXgIpqF/w4Udh6PiReFp5nWW1qnFL3DQFP1YIXEW9/uP/2U9KXhVhDnZXker89EojytgT
4yoZUdaOQpK/PPfMUbCEMyXJ2TY7h/TjJuhigadKpjS4hmzedytZr7dtJfEcFMa+U3UeFCo5VCcp
WCkmNJJlsPaXWK36LKP9HHn/beeybnFkJdPdMUz91SZwhXKyozUrcyMu0PxRoqwXw2pceXbQRTRa
Q3PfevC4R2HxTcFBX1BZqpkxDBz6hP51iJQvPU/qsN6fZ52tvgaefnHCXNOHcJnzmxO0DJ+uGgbc
l66cJYxMQFNQsN046cNQaQvVv3X4z4lZ5rGRpkJ3QZ+WnLnBMPr7VuXrT/i0hTR5iimpc1A7obdF
tKbxhceFJqvYrJUnVRIQuI4JyMkfc4ICKFA3KQvjL35zJo2DSQWRFVFJlSSxcsmXJ1JY4t0xScUX
+HFa+GZmdURhuKSqBn0/5tkTEvNUSvE1TIND5QEYVotmvcRJAzAspRORvQxp9LV1j+NVmb2W/NYB
caxLZdhJko/KQvhR76xDEBMjIuqeWZX75GJgIEBfJGDlH4j0Uxp206SMC3XSrRdM2i5czq4hEWSd
9+q6wScIv42IL6Gh15F1ltiPr19yEpSXk0QH6ywQKoBCayWHIidHg5kzY2OEUtQ23VMyvojqRn6K
CVGfmG4sBAxBXkIAmtQdUGu1Ai3M9wxB0MoERa62SBzdFcNRVOD9AG7sEKJEVXGxDZ/bD+RIZJ14
focbb0WrkhTv0NOv8Ac1CUNgrv89onJC2pbGm3BJOY2KsBPrMko4rhlg/jFi5kbhLqbM1tEA9UpS
XbbqNmxLyeURdhiS3w5qEg5P5+MbGCbPXUNaWRPs1RLC4Q46RvsQDZ45RO2UrphOCKuMfWvNSs5B
Jaqdkyqxx+fhUVY+6fax0cMt3SCzFVcWj8zdQ+RcaVThpnIEb+fKXTWqfy+PZAWsm7z8sP5NTnYD
M8OcYv1X5zQyXT/aeBDw1GcWCKIDZ25VjeOYp+nhj72O2nOWvM+mfKfnTfiHIxGZzga/qoNq0w7N
YhCxaLnSblY8dXGoPBUIV3m1jQwreXwtKuyfgAcu6DpwZjX6QcfpwXjx1DWIalDibBY97kSaEWjs
cgJRHNK7i81QCBo6RM9PKVnXmwCCoU8mRzkUes2pnW4V7v1Z9BXtFgwRnsHryeUpHbkvepvtFwgp
yzkHj8nFQ3qM9m1PWFIWyd7P/da3yD7A1fytyGyKHrecBoO4MdgnAhf9FVQeV36jOoDwWB5+C963
bZture2Jw18NpqlIsn8sPCo7Y/mI0cR7SkmmbLPc9fhVqLDG7vQLiw7SJkgSzPZW9yPeRi/eW5j9
Q6ANifArTabHPHUHU/w2QOTm9u0HFhmriH9srsiWcWa8Hps8unE18OxxIGRc49o0y5zlPQt7poZe
lpXn5PIRcoVUNZsAohQZU4p/urxF33lxs5zXMtEs8v/vOioDuhdYnl/Djxsh69nk0qj2cDtg0Njh
zmgtp05XK29KWyLL6Eo9JD35fZKITIYeC4vxMpH+HiA/yCZA/5VyFGRjY2xT9a5a/nzGh3EJUZr2
F3+J3SfZK3u5W+VDymbpQFhJcV1Psu99ViKz0YckwS2G/DrnHkATeuUBJVTHF8o0UDDi6i3IeRCi
07+oAUoPMZLWzS6v8hD2dqq6+d0rXHGqpxmI9f1isf1UNMoFEXkhwCDKg0XX59p8r9frbTUuHs9Z
aT2axgYwl6weUHcS7w2/thDahZW3F7hKoGkf4ZhbjV/QOvHeXF56jT/VNYBu7q94+PoTwFQJSLp8
sD3nC1vAAK9W4q9mUBcqAdBNwr/1wrwSVCeYGRabiFy0jpgitnVtoj8qTDpewKS722K/wEx2n6Sx
wj60w97eogtPvvHdGJ5tGnd12RwHbjgDN0tqSTMY36C3/kSQoun3dD8CRhPwBCi8buh5e5bQNcSy
14xPA2mbmf6P2F+nq7a0YANPJE2XwOTtTSU2Xt3fSWYdoNUM3MISQ6J6trHIAJAdKohPn93Kb1X0
NfWKxgbGTvaktZqqcEo9MKpbuwAaE1D9oE7BpE44tJDAKsJpDnwFOlYdNdpcaQYFyhk3dPvGIeRc
m5sTe7cUytAyrfuaClsuwmhfh9F9bOAxjZtIT4DZ0ZUAmKR33MdLs50s9GqWMQU7rne6NmNizghw
qWb3NGVsFGZx5dfsjaef+dQ69ksPxw2ElxePiIG+tQg66zyjXvt6r5lfTR3B5divsNsoceSjge6m
0XVNKgtOEH3zXtMUrMfVmQPlRd5e7XFU4DHapctzzFrpYdwrJvHz2FWHo9S12HFRp4qIW/u6VJRl
oh0OE8SxI7mOuP/jPchF9wzkIqYwtlPJGWAAhbwV1RQcHa8wEYhkUahPwr8izs7UJ+6FeI4suiHi
SBbSUwdebyeiCMks4IiuWKLmXxeiCwqVfpYYiHlcJtq8de8U0tRaq4pkdEdCtPaeLc3WRnPLGeV0
cVPkLCjYBXpKjbe3s7JZNitLk5IdUi/Ai/+JZJhtTpqWUuXYFKYSPbdAvR2BFc9mQtFMBTRdQgyr
SM2pmUnQA+tOFAXE8UeTIIcAiEiULlMti2q8axv0J+arb2GYaAz1BykaKlWArgj4PMvUXqzjIIJ9
PearDXfeto+aNFYz+iLUULYZQ0B2PJ6afhljwmfEDi5lQvWTH053okIPlB9P4HAu6U0RQxsSpjs0
kuxTHnWVxbKue+sVY/qjQNxxgUlJ8q51ovckUMXj6GWCoGvqhl+rMhp7ZGQMMCSqS0yoUCqGcBoM
Kl2nJUqWMd/9D5rrGE6xkZVGFIzXtpBxWLaB4dH4I3Tf9bkNI39A5GJqFH2tmQwhjR0y+Wl4fPMi
CNNsh4J6H7OLyekVyqzox8dNS/9Y3lmm+iPdOmrlmgDAxkcr5R2pWtwN+JcNmlMPl4HwAwArXwtY
beU57pt8ZRqGqtD7nJy6pC8ElAzjLyRe2YzXjf27qT3HG8PFs1gUiaI6rsQ13SoK0kWf+aQp9EXJ
vggh24Ub9A6Sy6Z16SgypV6UqiaAsLRAJdjs3N90qyWs08b0HA/RKlMtWitbW+guk5eT/hJF0+N2
tgrod5aorUJrlyeoMFEheTr+QRz60KgDJ7NS0mOiAgEUr5DqkD80znKjFgWY4Mhyyjs1J3YVKJ2X
Fet7noS9HT0le3VHjeGCrgwYFkQ2MLX3X7iA1swvKsjm98up66qaCnTvFF8cD1MhByy9OabQu8bA
rWwNzUxGeyvqfKrpfgB305AhxCliIyk76IfFg8e+tU03KKYTGf0klMBpjpwy7cIM7zEmHVYlc5yC
1rKwZ9yCrN2LmLi3hNaw3R/mw6KR3a8o0fnhBENXRJRxOV95VBVZh68T1Gn8aZaViq3YUwTJ1iAp
fRGSJ+TYId8/OSkaECiQxxxwVmrF/kIidoCFtN+NrbHfM11LRpXE7n7gp4ZVtJaRwm5Xyq4IDDRb
Ts6Ic4Fy0t1/5wkn/8kxaHSbdOlJkgBkKypiQN/H9QxpCtidQHvM8u4+5updym8HkUfP/TmcnPmQ
pJpZ+QgxtVDkdjmVy6thNshCDRLhPjEx8ts8R/bYpbkn2Gn/nS7y4FczmGJfaEHqFgHepljS5IcT
3WtH+19wtl2Ov7iuf25fhcAx1XxghA9cWvediVq9uQQSF6D2y/nC2nbx9XMhZSjTBJ1lo10HkQZv
AemXmUTwiE6JtdKv7tM0JIKhuTHNAG8noUqcR8eSjVcpGmgdKkUCEtNoEeKKkO+YA7pt/KsuoEw7
yki8NJp2TqW1fJ7yXEW1dYd2fHuwkgL5G9ERWhvJzj7IVNZdsAZeoMkLg4LuafEDZRZR+HklNIn7
x/i8SwMVoFu7C5wEijhTcfSHv0qqcS+3Op4svpFqdw6gAmAtiTbNSf8dzIf1gMACEv5NBKSH2Are
SHXA7oRKBOhCOgOfia5vCD+KySf9SVov2bmEV2Y+UkfpgVxCI/Mlnb4VofGwU72017HVGqeVYqvC
1Qo+h6GN16bhCwPZCwllszuUWftdGQnJcxeJ6dSqAuOlNpT8c0SQVmu8nEZhwrfuIfVlMEtQdXEv
9g1tCrStrg+cIRkdu5Rlh17Msp22zKRUA42MuOj2yVWpenwsjAAs45eQabUfdlPqHeBeH+OoXs6u
gMWX9dZ91HBpf+7PtPGCatEd44yqw9FQAPzGhWrFCtXz6Kpe1r9p8BUGRxBPAS4lJ/Bw9rhc7wxQ
I3FWIrpir2PM/hq3c21Tn2DkkxoSxxOsZhX7OtG3mjPWWG841KLHKNg35pBcv1OByVheZ2mJ/Zwv
RY6IrpxtC6V7bNHUU8p0CcOBdDaSPlzVyzJUyBx2fGa4C7awOMLcXxHfNhTohS2A8MX1CsAPaDt+
JjBVzOo1Wdu6f4xntgUUNw0oOTtt+HladZjpbv21FZ9A0kMGapwL/53xWRKi/2B/fz2UiR1vbYeP
Q2tb/0hIQMLSkCXdokmLc8SZjkOGLChkiPFUKKAIL1T4xQQhEVsZPVtrB9kFSRn9pTAuAsXiqLvn
Z26phkiE7h5bWQTA8ccJWrc5BRF40VgJIhXe6bQzhmqfKincHUbmkVZSTEEho1P9Tb79gbr3qkPV
O5Zl7VR3Y7uCbsIbGrLBNZhJBHt+uxWsx3ik47ixAnbigOUocnNLN7ZtKX5IrRBdFuEcz8vTnqxh
63ZglDaZBuL350FnDWIhcBoJFWqCNBkeRkb+L5noSVQjuOapTgh0W9K0yupW2vOSZTEW34EVjKsS
3shYophSKl9qLUMUbQ3VAPG7JhFOHDd3WCmnv72RKBRwdnJt6HSB5umm8v4ahqH/TdBABwEQ6/Lf
dBLIjHYIB4lH8Hi7z1ke+eRxr3InSI0zgoMCfE6pc+B2YwZZVbHhPVLE3YaU5xrQUMoUC2mkVwul
XyjEWAiwdaia7DZ27U5vQDHuDDgEbcbG6EH22n/iKLU1z1QFIMmf1q62WsGaH+e7QnYmbIWnSymS
2U6ndkiFLtiPJE5EfZDcpj1fjmgasMfWbjn367J2xIZPZjjFeV2UJE2JNmaHq5opzTUPQYFSsFta
TTGhd4a2eGy4+Srw+12Q6ni6E9Af7W00Sd4zEyX2qRI6WbyRbkjEUbDsYja7RBJy4M0O+jIvqlB6
nOCd+CJhg7Pj3tWvSTwdFScp8c6yG/5OPLcGXmwZneaINZRYv6fUIIzzWvDA9PaH+XRCMjk46/pc
NUTWMwvrFRiCkOeARkeLPSCy2qOQRPvzo1pKV+26X4wWct+NP3p7+4nNSrr8xJ6nvLo/WVUKXOAQ
YmKWx4aqlFn2/JD+33keYQPR3zqJ6WxAVLdL+dea2FJHNHvglWQDwWrnwHQCOUrChRHNvUAmVaMp
RoejiKzEm5MHVUftUf0PiEwM5rM4Mc/5EVdjpK7bQMRUi4BOVTO43hm9K6GYyuDge42KDG+GDu2w
eAvcgFXUYArhr5srwxps+LlfgV0kjRUSeiLy0+PFCg9nVngrq+3v9nJWh67BwHLjrdnJoB+SRWaT
+83E9X0TfFtBDDwCDpX1zjhjcW2AGmbUTzR2RjKXwbJbRbOPFX+Jcu3SJvtOqT3/3Rqj5Ch8x83X
Bx34TpdiFShbU1tUti45AcER3QKZWGlseHd4b7Jou/BQ84dPgg/mKZby4vMvxt3sBhy034bdPMuJ
ZWydLtPQub9E+yR9PiHO86pSWkyMty7+c1oRgK9pNm3QD04Pc71ZJ46lQTa259gTxMrJx912LvrB
nTLDTT0yrDhnEibpWECFu5joyOFHX3PbBGjewgP+zF7mdeAnHqsp/nPxajZhwrfUbLbCUFqSBkWe
3nPD84xnPYnOD9yI1SAe4GAea27v555dg8wMrjEXYHfz+UyTiNH5A/HFP96EBz36ymneBomZ32lx
TlwRidifqTYeAZdOt5f6NUPn5E/AYWYVgNgVKpkcf3utZKVNEtmkJxCQ1lQ8UfwEf4E/jzKcoB9Y
vhfLC19CYAIt7/LOeu5IwLiHa0ywwIUzfUr9RKmxemKqOdQIAiu80NjaY+2xFJmnYxUDb3aOlfIk
dAkBNeQmCK5+PGoF+uEcdn2rUMQrpgewXTAwEz7dnN5P5VGnprpg5b3vxKrg7WPwpdJgV8I/HljD
1UX+W07WZNdfNsbUmKyvxh3qgESAQbZkizTLiRI6fwCdjuqoj7j8IFWuxDZnUIh6FOhhYt4/TkXl
XFSRfZ5kt71ijcEx2bpndgMx0eJ035QPq2eXJvyYsoTVE1+xFpCMISN8g6wbLrjW8YolznGjnbdn
GNa4KEUnDQklgFQuvQcofhgj51Gm/f8+nhA+n8WF2HwbJ8twFopiONwpVZuorjzklF6yc+vY0uBc
2IjczMzo+P6W1CyqefXwgai6hpMSIkAH9cYxCKVD1xwtzmyemUShzxI0sDn221Ar9xB7m0yWSaa+
ChNSeJ0YAurRUMm0/ykRqWltfMSLNVcsc2nlI070OU0OrBtv64wpLkZUwsFo1RDtTK7IB2E9AwFS
XBkKAFQAvLCP7EepXUJ9DWVFqGgc19wTZ1oUObVClLEehWF8bCu/JQzrMtAJ2cbVkpyQd7roxIvN
BJheu7HMIJSZ7fX+zirA0wDvoB/p9/mGQlhKJBzZVLtJwo7FADlDv9vJVcQAzHjXOpdDO8Labu1P
/JdLAj5dqAOLx1AJmVjKwwkRUWR4JNs+s8cjxsQmuOCpjEukO3lQ0oIQC/DvRaH2v021RZZ2S4sw
ACGMvsFfWGK9JdU7D04+8ixYm+UKOJrMaWgQ6/0Aa00bvG3VWNt0JeKsqukKZ/RRadoEZH13ASkN
wEmzoGsuNPqpY8ScWEht9N+b6Q0F23vafHW6wjVWy4ri7VK5q6KRBiKNi0Gq6tdkLRekYC28zrZK
e1r4pnljQT3DhLPn54+Dt3/Z40kyFxCMrFdh+3ZEaLiwh8lnBVIKwTLem/1KpD2zRAKJ7OEDQEzs
0VPIzxh5qnrE7SwtwVbny0jXm716JS0s4glmlWxwf3UdAJc1VJxrMX/kH9mfL+ZJuTBrWd5ecAif
1gQikFaipPVbwPEMzQy47hRwOvUWtWCH3yIQ+L52ZSKLaGE5TOmI0buxh+PzHdtnglufLQ3lJWkT
VfZw0oLltkpeeeSb/eoJX/WIEUx19sQgTmCRpbsCAx+/fPclmqYfeEZvWuqTqye2YC5s8me7jdHn
M2EdDFUv+VL63/AmWg2pn1gKRboDBtmj1snjz0og5x/5u+f4mWFT6iKb8EMipS9fwn5vR/GUxJbz
TXEcEnr2Ivyf3aP0Nf4PQVgR4xc3EvKgl/8sZWSgni1x3UmrYcm+D6cDNNL8k9YzQAvJMskDu1/1
MabIoF27nvxFahQHVuNELuyDNmv9hS/dAZlncMw0FBJTVItL1mfYFuJrkQK2+uKkcEAdsUi8HROu
9Qnh39tsCOmWPNUrTkoV14vPURZR0MpZpf6gzBgTcQe6pcR+JBU/MoiG0O7yFJK5rbEw7tBSsoJH
AXe4oHWRR4f5+7u9YaB9nEYxn6hiqGVc6Ru/WbyuyZ0z7Wp5qCkwinqkjGktJsKw1GakATM4Cr5j
6r8kmraBDdrbAISzEe/dT1dkcM3aIhfqRuc/Y9L70er++zuq7rK2ZP076QjGOAA7zTJxBMWccDYK
VuQzUaui+fljRnegEgG9hPF4r+NPoc9VT5ZhOSgUP59SBXPHoiSp7VqgcM+VvofIlkRtV4bhP4YD
abV6ouHcFVBPOdDZWf70DN7SCYJt1ymBhdbUYKP7QhqnC+GBbMO1Ax0q5fFqtcHb7uq4hp2kE6+P
oWxG/gRP5wNnxVM2HlWCAU9r5EdyL+BfoDQVwZpoPEkvbBYxqeN6RP/O4I6n/m6t2PXQbVZnvhVr
XexayajyvRAeLr4hXPhnNf6FilwsAM1qWmSKlDqfPavSvfnHqjTXKoWWDcQdGTd7gvnQKEM2Krvh
nxWrDGdj1m+3WKlh9SKfeWp7eDF2eFAdMohjgulHYG3Ee1qs8VE8MSFhWdS0KSBSF9MP3KsGZUc1
aIbwvBx2PUvTzV03ujJD+65MFDEN5vYPVujTKKi7dIL+d6E22JuGAFuG+hWi6fQG5PlM9CEhk2lq
dUhD24ILhEfyXVe5lvU8+lnKpEQolPm3xTv2YH0uMJa4va/AaaAI5L4vDs34QptjVbpQz85hXhk5
ZZxn3GPaIC9H2wjCvfSsIwpSU74FkZzI9J0vTLE33YzNa4bR1JtqubnVy4vLrWlr8BE+wp5Dnx63
56YM1cDZ3Yrfi9KVLv7f3gzOEpXzKDjUYmHFtiqidCntzl8nzsWG61OpeukM3MLRx4kdchP8porB
nDYUjQsuGkspD1jNdwFfMmYqmkJa20hffHSD/ALbUVivRZwS55wyi3hmjWiMO2aWr6TDOwsfFLmK
1hR5qvs7g05GZzNuZoL+AAnfcC95SeI2l5NNU50nt0H1D6pnvKp93v4omHai5iYtQUVYkNPHGoeg
O9SWYLK8QTfSsH4P305Nc4V/zwz6NKidTI+Nkf+ImUxXZe6ofU9rVCwVmKzF1tFaswfev8qpKlbk
KqZ92UofEhkRiAQPQ5jVDT7Q11fe139TkguA7cG7y3I2MTPdgSKjnle1je0gTNOCGNL5ftfQxvLt
UgyLZV/xJ7WzZ4qnrbwowW97715EkjENVx588944cc8mUlDoOB6mIckYKGNLLdXqQlRduCAorQU1
zfTLkUhqYZ9L+Qglao/YN+//YifmMNsThHdmlk+HCss2PkMtYC12rrKi3cXi+2eSjuH3R+a4LUl4
nJmJ09AgouJMMCN2XZi4n4qM4AC78HqyFwZ4eKBT2TLFrmz1ACh2X6aMa+/z4A+DI49fB5jUN2E4
1MnXKu0NaFGP5hVEeRDtNo5xb6o/ND07rqIrMrUfjwGj5MpW5KY+P+UGJ9F/cyJySw0CXFBdW5cm
ZbNIYLHz/MkINd0UhNjKPYKPUuv7vOSqPB8yO7Cqf1RGbnqPCGyy9qccYUw/wAdGvAVCsI/TebT2
uIfi2/Zjsoi2goT5kCyQC7Jm9813U06euCoKF0F1CjmIn0+doxE3KgEI4CGGl5oV5T6xUtmg2Pq4
JJ7GepasSmS1Srdu5qj9XBjugR8yS5xNhYHjXbHQrqtLwYCS869jCVlGIdXts2zzu6efmQNjBQge
623oHqjOa6ZZpVsAlaUTp8ZIxNYnWhq3uypyiA1fwiogbxTnFf6sqd+WWOic+TSJhkl9J6iAo2LE
iGYRy8/SmnuWRY1UCcmbTuii6BYXDa+mXbxm7aEl2//o0tOYODlbu1i9h362bfG6IqLJE/jv3mUl
Lig35zfPEW1D2AhQRPq4aWPPbVg1Xs2u2jbITM3brxn39hBr9n81upnbTbCrr0DYGWvWaWUavMgM
yqn26IzLkCGzBUAPgQBSittgmgbLFfl/TJFZDv4eFERAqDvz8NkbuZ8hgvpKvagORTiITkOqARCn
leAqx5IEStR0+Zib/EdmGuZfSbAbHkBvmUb6tool4NWu0DA8vn32HaqJmhhK/8UFfItD0yMKHZ4i
aMQOJ317SK/dVzeRqVHBMMS7JaQEhMd2NMYL+h0sE8LC1ELBz2ubMKHDOz0wwbjqNh+LYfAuP19P
7tii1+HQZf5Z0vVG36NB7+XlEfJtoEv1WYb+NpgOUYpblXPuN1YWNO7F6Ea3cwEILYIOojG+NwLS
Ah1BJXB+uolCYPiTNI5GPAkX9Dx5mS3HTuC4BfG/392PTlMC1qrgKygIHdsDe4Q5v6RbW+9O5UMm
i4Rkx4TIb1K15FWyXUR0o1mIvnIYCh5gOvOznfaGeRMZ1ez2mRacg8tN4MpQiGkRBeVZgp8Z8X9u
EKEg7rCzYrQoaFLx9bsZgWgkNm0cz7dmxuIrGqxnE/pyIrvipggLieBaQR4dMePS/jtQikSc+ZLI
QW1dhkNgHbCt6PY4yeNM2jVxrLsiUdP6mdRM3oIHR7IPDzD1FvGkKcJm1VS/mbEamv7RdEMPc+F1
Lw/3GtLilTtVvccDrCh1BTcq0uLGhzpoFpPqVngAft0AIOfiwb99ChmmjNewl0wI/MYUCXfTNS1h
hSzj4JZ9lJ0D7jzjLmODoP6wvPc6+fp/fnvj9qpqSMxcHS1FG9btWU0VNqdf+pvuYGm92V13BSf8
OnV7ynmE8vS6u/f062kwUb0d4oUWnnFeVo5MDZEw3/LQnlKBYghEwITCeH1BoOIoYQKwJuuLZX6m
x/aw7LA0CxbzhhBAVmELgHfoXxWfH38wb18xXXsBQ/JBG83i5O5FX3wItcyNpnMGwFEem/dtLAh2
0xqvP8wdnM7RaNvHzNJR1m3o4DiL8LhHszHd9BdZolpQLElwU20ea+b1H3xjpriqaiOdVuATAWCI
UhKs6S+rXMD/7SDXZdtI/7Lkj7DHA8o2IRNek4yXBlv52jIuZdFQ8glOq7QB8rTDPuDWrTfsUdzq
6gXD/uHOzgK8Z7RH7bzPvbj40J3MSz6Tvx2SXrv1w8IZa3cS1TGRwvifI8bEATaTuhNuHGKBRqU6
WMXB0StMGpQqwpzDeSezxtnkHfAwJX6JvjbsSFsyqJiF9VBFyNx0Wujav34aFFB1uVNwsj3W+ELv
DoWXvLSj/NcByNIM6UpPMWvx/zh0Xb9pzEnhFDTvGQlKGlAo4/jbbTydRIf1uYQ4VSG9bJNMXN2K
KioHws/iZUu4Qm6noIKN0xyVZA/h0yJuYBKkfrzHvDJ7Brg0iFIMNfYqX3UGjf96FIh4onAkICwB
UXA4tdkASahplLyTQDHPkzn5w7eGp8/DQBOpF80OJUcNQwJJOB0erCk+5Rxo35fD8OIcLQ8EsVJS
8mwJtXvuuDpE66t/cgQxDr/KHBc8YRgOKTG7dvO26mnKXUW6rYMDpUiRfJepHtNSfLwEUv2hH3N1
3Yo/4xfVenjAFARG9lQdDZuTcXrxf+YwbRou0JqdjrP8PBJ7L6DG2w/2nN273RvmjhvozMNdmpjq
GgautnOgArYZDVMWBQ1VBYRwzyCDtJgGE4oiPgst8iOLoPJTOMXg2uzrXj9a7uYVbnIZ++0i0tx5
OJWFcCQK0l121cAbbdBvPYxn134U+YE0Js+1VUfKsz2gsMzRfOMlFA1G4vWOc82tdP7aaHFyLLum
u9n7NG9CSq11+n3vq5gKNOqRND4SOdsnS7igy3cQwrPZ0pnPkqa7/kb04PtlYuHgEV7YXNOkXcEN
40G5BTZKpob6GsyXxkaN1TkhcmMwqHa16SWKvavJ5s1l7bdeWsa7RF8ADtIR8LMhf59cm9WyDDz1
xd0WDkhmwuH/otGsFMmjFwBR52jtSykyXfdUyC7C4VnfhoYB3lc4OjNWtENqDfZr4anMn87CHmRY
tL1yiuVjXy8yfiu+e7oM19TCiQDldt0Kb38ZMLmkFOtJsGsx+/qALfGVMAhB/dBE+NSG1QfN+r7N
baE7T6q2q6ovo6YTa3XptbQWufvwrtj3y8vPzswCMq0RVRtuJtJ3wp5VSpy5kb+fHJQURc6FaEIJ
BuXIPaty5WHPqMSmQGourqdG4WugJ0MCy+2BL0IBH0yDk4so0nRCo+/16V7mSiVn0FoYMSxDTR/C
UBjb69CZ0FzAMQpkc4frq/o3rjgrqDPbf7s+2i28ULtz9cSOcRP80MIOftCWubflI+eDRNP8/aRm
zgicmuKfYKbtpn3lcP8Oaz4wGjnbLAbUueDZ/32NooqdcfprkR3NuAuEGM6Cn7QKqrF2ChZ/AVbu
MH1/uU+Qo7bcjMBjNFvQmAoamcEzoE/ixh2Qe939ro1IEmLC8kIJi9fmabodtYbjqkQnZW9hVqEw
K7Lj7Hupw6MNXGdAwb2XVGbve5RntiIho2gQwfB3CX7SSMU8GTOkXNn/1d5+5JGRxZugf9nyeYDT
vAO+b5nkzmWxYQ5/+DGVzEPNoxBY4tgl9ImGS/p19vXr0B5e9ScDtT2tK7KRVl43kL1KGY5e7XtN
q+uUmbVSz0GMHP98HmUaL0nnVfczRRc/Ga2kukVnIFRqvCxOAKf/wZwuBxCCqXB90uRmHwaxwxmz
+EBWDdbHGEDwaWemYUDPXFSx2RqAIrAKnk0CeF2pzYjrepW4F6YImHfG24YzM6qEgopQOvOrxFoM
jF/H4TWItD23MXFJumnrl7robLqxHjWc/Faa9LXwZSfbPzL+eQyus2KjGXqkV9AILne+eyMH46s3
squV7Z0H1+kGxvthWilXMo+cGePcS/tYrfaS+7Yd75Tw0bDWw8fbkTF/H5Zh0kgvGjms1u49fVhz
icJr2iLlKWSKoaNKQVMuAmJwTy0ixLDNdNogX3NeFcAbKME5qmeOxUlpqFhJyWkhPZqxGJIDoJhR
9q+kF2jgiw03zN/nKHUvLZ+9UcGsBv/RoQ4z6UN49OJAzk5O4XzGtcckqOkVoGCNZ4hWyKcMle7t
sYTqrKMY6LnZtOeLExoyoi5Ll3IUAy8zXjynb/c2Jjy+MFbK4aez0G+OtOAhIext9PQWcMrQhgUi
HtbA2A6b3TpvmlB82omAhPmQrdO+1ZUTLDwYJeWpOI87KV4ull4YGX5E5U4I+J+BrnPMlbi0CiJ0
r49uk5jnLev/weP7B3fkx9N4JzIr1iSiDW6UkJvshCzoLNGhN9w0QJ5vU+hshoCc+6japKIdDpzW
J3KIlbV38LZv0P/FXbZRDEjKYqC/L4wa34weCdCaQGhYnCRDhNtzyfhC8VtWmfgJre5OgLfW32t1
M6JSircp0AHwxvPpbRcyMl2vHBw3pns+X0Zcna0brY5A84mJNJsMdUGVBb5eXyn97BRrp+YRUTO+
yIoBhzkQ6Fw7irxuoinZq8RIoAe5AIGjewEK6GHiCYitIOJUJWte/miHnza9AOKklUccGuUGjW45
dnsJvZZjZKkEdWoN4dYPHx8TmLNRvUA5cJ5fkQiaVHwDSkN/SZzKXCBOutL0BQ+cwiG4TvZBw1I7
GRpvmd+nYCC3vbudB1eyXlLS05CBOtGaLn6jcJfu9D8J6MTgWJd+jl4DBs1dAkh4PtmCopyuazQQ
SFsk39sCkRF3MWy+Q5DGt4SOgpVxJL5WSMsGNj4wr2RHMhDGc/ZDgYnRm11stsId6wlbr8Tj6mDq
JYc2iL/1MwWgvNv2DvtWCoq6KPSQiMMFm/W3Nau0Lfmk+W2vIogSgIPm7hpzF8+at/CgGPHKEvrq
5Al9Btew/4Us6kAF+HO7eCm9jXwjJZn+D3w7G60gK3gyAXy75nzMTVi7oGErvvj1raEZALhwOgXt
vg2UEfj99qCPBXzJVJohqFvP5Cae06ck1yZEmILfoak4c8TdEH6p12GKeg7oNVDocyACedqPWHZb
8hIaW4s60Df4T92kbpCGBnrPJFqoURd5yx/NuEqPffTPzJTHcH8r7JuKW73yN1bDI2URpkRBWmf+
BNy8981kpBJsCiJphqgYjzJfJIROUcsAAy1/sbACexaD5ZfyEl95nJYdkToawxh4JEsT14vxi/uF
X25DWvEGG0ZDsJbrXcbXRjR2trIL3rm4C7KNmj3QQG0KFZOPuoepswDgsx6gn6g/Ff7xB3suy4Oh
6IJjHK+gDb3N3bpBd41eYbCs+G+nXu2bhTO4U4T9TpFFLqDqc/OcgrV4IcAYisEO/euOjVuWBuo/
64J5sI93SpBilPHXoh4spa5mwnqhRjhefC8wH6PA+TjhzpvZGPYwoCNbpLpR+3/sfm7HBjzYN3rt
LEaGoLhfEZnkKMuhk3nW5J782gtc+Pw4FQ3Jpjgzht7Jwza26O5cSNFoipwAffQpIl6cJiHqrH9H
oiUHtCZ88WOcjTQHIJdvdYbbha7XDiZCWtM+KUojvwS74BmQGhMfn9ifcHDHedurmlEJomDuvfLb
ETL0Pj1lRQzfhvQH96UdWg4czkOXDiPrqcrevQG00EeMA81/cQaKNv0GRnpydZeKubpnIM3nqsCW
KIpg0nq4P0Bpp2pZ+gdbs0kp+TqLeL0S2w+TdJUF/d2b3N1UPZ5HlBFnwDlZzSw2uNi44PIJ0jyD
V3BWa5RXXmBnxX7dUflZmuSlDg3b1aGO2BbvpgfmJ92N4AoxFhL0X0mYXxy4xH/zuwcjz8rEAm2a
lc20HtSy1H02K21B4/3hEmbMy2sWHMoa85liZQWQ1leR6i/bFpRj14thbT4Fc+z8JwGpDqNoI60H
hK9VD22eViHWv/9WcUG88cMtlnGM5NFsRa+VD+s3rAqoAsbrhGz5ERqjuK7hmqQcXMrvtawhQ50i
183XGLymnBP0dCv7Np4dvxr3sPuPVXn3PfI6yujqw3c4vPFQIMpVmaKo3OS7Qo5W/u7GymLHejW6
1o17fkTWdJOc5/AFQqpaH1aFTTDC5A24vE4TgQTP5T8r+R7rvWPFDexBkQ06MbBIB0HBfuYQ/DU9
WuaeYHm4hsFaBpa+M7pNGgFfQztWHMABs5riEupplzy1yCA/HHKhILshVeXy8maqmm1F4pJxEw36
tEU43RmVBt5cPJxDcJ/CljS78fQZmgV2MkL5MUJ5Nzuo/TfOyO3MWBcbYsTkLRzCuShvFGreUTsN
tJjN9EZP2C6PC04O/FcGSZs4Y0hWutao9iLHbXYAVrZ02YTx8jcx1c4vGCLzLyARHrIwLJBzjeX5
HpjpWjTqASZUhjOlOSCf7de2z0ieXl2F1lWjLR22tHw+g/p38OaBKIloJBKmnu/s5SS85vLomzNO
qy/XSfYb9p9oaf6bSF9v046P1eeIzsKfuxQ4z5Gf2x8bvk94k3lVuMWvz+D7kfNVos9yIAV6zdOt
hnDnQzSx6gH/M4krKCTmSv0z4y072RAgbpmXUWVF2fRkg/QNCX0lytA+Ca1atOhCS+vhQgMpp38k
K6ySfOoOt7+mdtDn+rgsrwbqGPLyFxm+I0Yxdk7VUynDDknz6bel+kldmekj6wFvz1QJDuq5zSKi
eKHkdkZPxmWR4c54JxQs7UbwP38q4RF4ZadjYGGIxxEWkyIwdCWzqdmPqh78/ayjTbKhChSJgVER
zG4K5jnIGz20sSMh2uuYg2BLCQRZK8qCs1XXkj3Z2Lfp1rPlXKAxtRaErtxYDb9eACyNPwP5sxmQ
RuMk7VkAjkIIbLSGkmqsKFE/2L3vufIwS+1n/93E72Y5IGdPUN8ce+uyTGvRiFKIoF2P7chjZAW0
3jUNe7OttmEGb9JpoW6PD7Y6BiL4oUUf7PSK9dJFQnYE/v0/xHeF+bNaVPZWOKCtwmGXzv36XF6u
EEYBEtqAk/HrlIrGBl2sKughXammRxZ6IVzk2Y4a+9g89cVDmbCD2PjMWSDMUtIsz9amr0qsM6kN
BKYDNGKuH5sZEmJFDo0JhY2pJXSOm5SNupc25HhN5UMAcGhKf0eO91QjVYchrVAFR+XARAEp+tk0
oE5Dd1ZVsaM4cipMQupjhImHcf+jSTnc8B/PpzQJTRh4Yz973zkBfbLuUbqmq9ni78Kv7iE3pYGB
KTqerDVgq9LqMgZ5j7jjkcwdnU7umP24S5kA3VMA8A5iZjzmnXr3EfwK9eTjBGmPCT8pS9SEM9cF
eIYKyh1/OZBQeBVK+vMziSuJgf7UD1IFirN6CjhnBN9VMY/p/k8SVbZKemBnpLYZoWsVT48LtTqr
kNeOUVtWM7ZdpDRo4Zc+CMufCRx9wMLJcUL1UEG1qNO0jbXw79ZpLTJasoaIw0sDnF0RTcTJsTqh
Yh7Qf69x7Fn2suiyMTMtQiVZhiNlMmgzQbhXSMPE6LJPYIfHaJLi+LdTU66q+PHj+FVmdoa64D7o
ru1ifzSCOAUflMYkmGpkB9E26cwzdWRXz4+7jd4g2nh6MwN9kn5d7eVt4v5n6iTE2/zPJPNUvRmy
PgzsUaD6V4t8mdChyDHOolosmXQ0huXE+L13MHVEhdUDQe2JNb3HfgvNtqWNWitycly9aWf0oMKp
YhShw6vO1tdRu5/6dWfFsLl8FyR2IPGrx2I60c3/qc3nu6BRA6YbgoA3/INU4DANQDfVLTc0SyZC
vBgRFxOvxWzNxQwKKKOP85M/7C/kB0+MyceBT4FV6q1iS0KqoToYKC9cEPvU4mff8DnKvWZy9yeG
zn/+CoBvXX7DSGAubiAYxZ58L8A3B5M/ZozsBoGFO1o+uQGih7b4IXQQONptmQO3vfvGyrioViIw
DcqW3uSydJ3LM6whrUlXpocpByi9hX1+thZKaGA+rp+jnnHLI6WbxsQWOHs0BwOuOamHTo0AFd5g
6RLUZDnFRQ9gOd4BgNnp7+Q+9ODpma5/NBwivR+1vWX9zCfXWhaYLqMfG29GROoLKLqTQVDXhvlo
j+A65vK/ZFd0i1GCLwfIiSWW6r0toiDgeEuGcLjaU2G2iTcHAltaCN3KdJlnljgvSs3Zc+hwSOhc
sd8hmQYRVwfb7ucFCWXCCWPUi34Eg0XSSm8MqH3gqgcnA1WIxzl790zGak5bErrXsOWXw3Cde4cI
S/QJdInfJvsRLwTf8K7ETvVKg7ik99lxJagqNZQpjoagjMeYCfcc+1LMwUaVNAf/es3LgAIRlAdM
soyuHCM9vvBugPILi1Xt4JZyEP3wd1SOLkIH5ltLVCgrCsPPKP94jZ5sa54XkZ+Z5G47f4r4SOv6
gAiCL4tYO9g6OXXSNVRwXSWxu1ljT1xc7V5dnpPELsyWakfThgJLz3ACzkk0x3LWH205TBnC0ecd
iOBjLdvo0RG5Miy20KadSB0nJACDChDi1CcqPkw9doGK+PFygI5SpXSn4PjIFnuy8RDMIQg+tne5
klTkH61tLrqFQrBHSjLsKmeMcsY36NTjYnjiAD9YYXOhbCaRdg+8eZypHRqZVCDpwOtoS8nTB3hu
ySMYu56yymZ5qqIdGRbGMDYgLayVd3wes6saRd3SbY95sKficy7lMYU7u1PpEnSDVMt7sC4GksTX
4QmQVYAr/oTR6dL3VyAtuX+BXUsr/cVjdJD9oeB8MAA86uKNMLLiFHknygzQxNG+Gv94MT4mZgLL
KM9/jGtonLafQPw5NUzXoq+ABeb3vZo1KHn1qd2d3xmzvY+5UPzkCSnxjxqN2aZ+6DCOjbnAjPoZ
d/0cbwGfDysnUoWiKDA2cmRFKtkEN1wXTxcaWMJzyS2q9rvbr6DcQOX1AAZ0XZmH8yqP+/jQ6wjp
87buZTOtLhUqkCPd2hpfRLbZHyYpOmcwdUgV7i8N0G86FTGHcg2+QHfwYJ9L0Ik8b+N0QjItTJHy
XAAU5vwjSK6oCygbL7IWWPWMnumnC36BXlUe3KOGS+2lA+QrIRzFKBuqvDsB3IuUB1wkqhXOQifo
2dVcr7p7ChWL1k7pzKueEFF/OJyuRLPDim3sysp+1Oc1a2paFL99JLQhjLwv8UPUJRHeT5aRj5g3
HpwS0Y3MHLTSdrYFoVxeV0ZGyUQMeOeNcoZANSc90miVW1XKXaIJjqO9XK6vcR3IhcImir5pwndk
y9DzXdNcseyOf+YJBIXN8iGJ+0lVJmmNm0cG8U96+SJHWpzSHSgcm7bZ9Rg8cJjBbWpfahysChnD
HRAiymwRjAksk1G/jR/9HkIsFzYbsx2aRp3GpN2IM+3gbmDjSZexnWwb/1scdhW1JJzY+t8ao51S
oqjAxCoQ4qi50YxF/QPKSvoiz+ieVO6UM1d+NAujqc5w0mqCR0/LpKjhMzC7XCWzspnjrzipwseu
AgxisbOdiwqlzX1cyFWND7eQj43MNh2KpnbKs57wsdP//yBuD7Q/PDAXNbJzChjvjhoe6DgbyKoC
QYHl10QMtANQkFxBHJaY5T1sqB+dspdtsrPuaXbUQnpyKQQGxmaFe+YxArmSdzZiLezPN15IGuof
SBJ6w1F6YW0IkGzNWJM1hPoaE+MyWUV965LVZt/66x/6ke8XcLjdtuIlV5o0HIav5ZvSs5+gvaua
zLLu/NjbjBpKdmkWjAhFitIiB38iVe2YL+9LxLmHul8w+TH0ECGksEBa+WDNPMxgmkPwfXeTux9u
JjuwcY/FB2MPX8Tc4y8dZBv90ypkhJnPeHhk1rlyxrKQ9xicQJH4v4nqUJ0ANQAlJ6gVUcYAQNHk
8+aRMkZh4tVOQEH15VVx/Vp1NNKuG6mRnKKxvJxiJ/XoiV+c4X0iTQyMV4M7QiafXl7+JjuvGQsp
uc6EVt77610eCf7xjQF/ozpLS+v8tlADJvTZS1X2QLiqZKzUcnl2m8I8xqqKxSHI0/dDXcNYYyx1
nEZW8xgzXRPXG9pygRJYSkvO2LFOq0TvypAU6nGlb+G20kQbMQ5/Ax5UbHmU0bRU7v2d7lEmoSpB
VFGiWBz6d5tOmFL1zSzi/HfkIrObOd6+ymLOiBqUo3twu9P+v+9DVRFCcOdt1vFai9jhAYR8gs18
2eXphTlM2M53O/bSvJM8y0iK7u/dPADUKCKtFnkB+xxQUpUyPkC0MlO4gFIDGXLjR0MHzbt66Ryx
DesZsgeCgZ5yl1tDDZ06cTnN51mVMpJhAgd+pKRq4S+9VCBZJXvoqNLlQnwERG2XfJj+7zSTcyIw
dc8Ww2YJNmR7ZQtTuBu8ycOdpjP+gbGyX1mr2gMgKvyqjbNq4+3Afh6mES9isqG4iH393Nj9tzNd
8d/AxbH3tavyrE9z70+uMBNIqAP3gd2XgicDIBXxKdcOszkjG2L48RXNNnE8EY4eiFRUn+0EuL4t
78pyRe41MIklUmIHwvjU0Joobk8/Cbnna3Oc7Z7Olq0sCmc6rTM/txTjGwUJD3omSRNTcJ9hkL77
cg6dKfj3FP3lfyA+TuOtcs5xKOOaP5x/ZPCrZXEBHZHiWXZ7f37byVlz7Q53Tweam6NSPglABIss
joNffCm5pBMGp5rlW0+STRzPiNy4ksJMbhRBfzmH+BUvjbZdxm1QpwvCr6ZMCfNTd7kEuJzQfQXH
QLBsl5CGykyfympwNB3vQKLemDZ0IiF0KZiNuhF5a2hBbhw16WeAJb9+sZVZ914CLuZe6gtmdpv+
SClx85Ig55YVRiyMfaGFLJq4IXNhLZNobbRTUTDZ4yPiIFszd0pdrZhuog16HRtyAWmVm6LqLoeM
K9Gbie3kCokDwLyVJL34AZWqZhm5gAy0WTokSLi+bd41cQSLNJaR2+BNnORHw6DKSk05oVhJRHMR
hRv17cLvMdoiK2PfjUoGtLjIZggXwwroSANffFFg9zuJAMlYND//FdNxDmSgLJJygPjq3j4ui6S8
aXjfVDNVloaRaREALE9JcisuSQoXEB9w75xJm1c9YQyM0R1luQWzSE6O15mp3GRxXp+TQR9lWK1e
Amhy/RH5u44NF2C1CmZKjdCQuJfKaD85HYsBF3wxaN3zsF05ygoHLYnZTUwTrW8V9IFFsOd+qCWy
b3o0KWZ5VIsGW3XbSEzmOmdcljDB4uSZeIF/MSL5FZPH0Kz9Z7Yocuu3LX8d0eMBpJtjSbn/uU85
ZCbkgEm8fBpGpHoUUTqmAOW6mrbP5QhVp0fVw0yooSlP6HR4q1zl/kYavqtsMGEUHk8FkvBV8by8
0teg3Dp/NsSz2h71/DyVObT7ExDCYSFb/Z8QxwfTyeu18248IP82j7408bVURjt1IWSpYpG0pdj+
6aqaXF6pvMKywqEbwq+PKFDF8NwpKFfDeI7klG56dtQbzBtYAEUaXV/6OdgAL8e16QJmiax7RpRj
H0rXI3QM6nqaCpxLLFf45dcpD1mcyQN3YxFr5/qq22gDPCTbNhCG+gpFVm09jwCf37dIH19Xaq5o
8Q5MNeWFudg64pDKtXlmQjwRWizcT4IJsXMZYLNQOHf9eMYiTCM2osJ5+RfkuJ6Lb4SsWJx7cFTZ
juECRzi/f1Ah/PFTWzOz1N4IgCyyfUp7xwAKLePdfrzOM96k98n3zBE/NnqFX9vEOJhthVNFhzI1
kNs1jGZt2v3Kgru1TQ5E72pFC1r66RFnlqxqHfCpwLrKX29xsfk7An8NtckUDknfHIGlgFNvBDo/
J1oYNkOPGu9WZv6xJfFdk6xc8ItWv42WNWuvPNH0L8xbvTrlXyl7S5ZLsVDWUoJXTpGi4CjR5hLF
id530gKOBN8TywTQFJTH46ZdF2w+k6RS66vTKQ1nFaFPcrg99pgYzqx2DR5SXQqZt43qn8tXOoq+
uisLihwqOexDxGLi26Q7Y5PF3tyynP42qz+UKEI+/UWwmZMq1/obTMAUwYkQN4vJh3Yh+3stbAha
lwialtEK1dwGWslhPJUR2lUmgf5XqHowWgsNi8Bc6Tc1/JYp+SGAcaWvWokhUnYB3X0qQxvkQPpk
3NDX92FrNJ8gDoY66kimqyRUkLZTdBaVW3OAF/C/Z9Pj+anBewqG5fpl82cwzKL4H9VsSKVN9CDb
7W/6sKHMZ+9dYfKKAULi8hWxzrkSwm3SdbOQacIrST76gySHfg3U/3dFKuPv1ceJbEsYxjoT+Q+x
/UvakHXJmVxsHE3Y6hmrNRdVvq5E7QZMsgbXCMxCgysWbgXPB7YdjxsSgOICoXigRDP46OetRUKt
Js0hh2EicjIDcpsJR94IqBF61hvB9eyzsqeBhY5PeZVpOL1sv/c+UJqJPIMOf89nspVcCqQvnKel
q8ywf5/xSdyS/SiLDXgtQKyPNkY3Leb1lWPHBa68x1lkZxmFUsD6o9JteUlsfQBjm4NYsLJUMWHm
rgzf0PsI1GbC+jsX7mNTtIBfM/d+o13R+7lqxWv4yDqvd/RQ6TFGB7oFHZEwSWkPqqKvrUG8jBWH
Pn3iai4G9w0tpTCKPhMNXmTj6joZ4jLseZAqH7Eb/qo3D9W4zPODzzONB6CHuTwdfNy+0l4onop+
kl4iJXPSVjnesPhMlgGOTWiF1ZJ1ZnBP8jL28JB9Tv2TJY2G/k/e1ABNMfL+cNK5aOvYVUW7ZJnO
MYJNBeR4hpriVqjr6PlMKj7AvtH7AU/hXc1bm1vDNsHvjYraFOv2Jx9Bh3zBVXmds5hE/yfWYaNH
O5XWSkA1IJ9OUl0RfSYHXCAz7Dazf40hWUgTbyVZiWx8iFKfs1ha+imVbMKJjMZ/prA9nC/UMqrx
vujAg3WYSd6Rk5YhpH0ZwzPlrMjrDWBskRbh6tyWk/PtbPBM/TlQSfMkPHpa8a9VMccSeVa35Ybb
SI7dDtNBl+g7uKlgP7fxHvODWwyUv8HwP6bLZNJogp6bQLKkfOhxWxmg3q9j9Lnt1aaTgjd26MS8
cWl8Uo1dF1M1FJ37jsP9xalI2eknEqng3TyNKKspjWlaFsfwub3t2RhuNkng5xS7lwpQvajtq9iR
fcB6IN6GGaiq4kn6CcL2fNqv1m8b12WmW/6g8XUhr1a8osyWnZiqth0o7PdsCtTKIypMmerE/SQp
q/p7pEUCyzkD61Xwhw7ZiD/FTKuZ7m9RUQX0S5xGwCNsybtZkWJ5D0sxDjzDqVjvyhoQsxk3efDK
nQCdrJOV7LkI//kH9gfIF7WyZ8j64lLHWReoPmnK6m15deCvgocwEvz2EvU7TmBU1TyF+LGiNv2l
hCqueiN40r6mCjIsza/d3agWmBTOSjwK/sozYQSTu3DnYsnToSwzrCehh2MSB7WLM5Tt+fkw9HMt
UXr9rCSxJBdRZ3MLaQnD46U7wk82DkGgR8qDU2jSmQtx42veJNRwWiFWD6w49jz/jiDglpFHoPx7
Jv/leO34gQ3KwYwb7qDJuJWpH7z/gEKSC7bsZkMWjv4rptv57vqcUkMC6oMT3LE35QzEUrWSugw6
BWyucbr2oUBbESengUGXfbo9/rao5tQ6Ref78Jl9j+c8opvRKymXpUJNnsUgmJMscennZta0C/33
40IGPOtc/VC4SuGzSPq5Hdg9bSDcYlPlHA3NYwrr0o9swJCkm6uFxOdnfOBARccFbAmebOyhapfw
QZTQT0xDMD+nnEFmJ1tHs5420OncB0YeAP0PevF0EHRtFsRIDfWYhzfSuUnZFxf8162c1gVMuaFX
/7B4j0Tb/E6GQV66hufRKHCRI0qElS15YBdZ5RZLUAXrzC9HRok/Hwhmzmgj5Mb/xHxeSayX9Ogm
cPaNzxjH+XzuptrWm7Q4pt/gm5jyNDgsneerTbebPPlefB9YryK7LfMLmOrrXMKnTt8ShHt/7tBi
k/CztX0ah4JNdG0cU8bd2A0QGv2sBr63KntmMi7lP4OfEl3YRAR/x9eSeLHnkYkhEQLHc0F4VFgg
+amF+5zohAiNfD+KKJH9T35GDki0Thsn1YaCEflyY0Q540nPnuM5TTb52jql9pZae3kx8c0iv49n
IPjmj1/aW53eJYBNkLdN5KkJviOmPmIW6molExXtitppshuUkcpiVgVCKqSwxvucUMhO35MUZaQS
j1jYIxeAAkb/RTp11AkS2iuWUy63yhLM4T3RJshONIZZ0GKFJaUs1SY6EBINxUjYTTvIZTz7EIVQ
UXmEMC4jFdQ/SSc9gsYFQ3r2tSzJCImdDIYT0q+HuaXd9I+/SchJEZdqbIF3Xrcy1MG0psHny25C
YUjtxqAruPfe5g1vE4j7r4h8abQtmwMP/07/M+S2PQZxb4TgwNEfsiHDWvJN3pWwP/rYzVQ8jpGg
4jjop0v0RF1dO0OKHbO7TtSB1IIJo78ZT1r/pclagk7yVXM9o60dIZLg9wcuC26eq+x1wRLGASud
NfZEqdWVh6HBX8zeSeHzNdFxG+0BtGnF8+6WxbvjyrxlxaeNNvySEdjo7Tojpx3K5UyfZ1UWIyQ5
zBsGN9AFUVG0eKAQGqmAC4qbP7EBCYBB99ZT7qYbBRVMsF/V+CI8Z/f5IuCpBVzkgBUM5saAUuQx
iiMJjujjroHJLV/xVD9cQVcV1WnWHz53QKKr2dlIJwUNx/+4xAbRt2mstlTZxOElFB7XF+OvverC
kgYJjxBisvQk5rCZDjYAsUiLEt0U0W0W92jNXB0ad0Hy0OY7Xk3XDOz8wW6ylSIrxhS7EtH6hnxD
T9plFsMfKyvG7mk265l7aVZV3aqICneBQCj8T4vZt6a6vmPVJLdfOiuxqm8Q36mhHHCx5kYIRnrb
qaVfrrmuEkw0vbRjSe1zAGLW2A9f/xCbCyROez28LLtkkP9RFn6TDtF4I73QLZAL7yMqb2q+oKBH
AL9QAMDzQn5+Qb2nE62UDRIjfgkeoReU+W6nbFfLvtSsRvJLbBldhXgcm5o/cWZtuKKDxM8gCbaO
k+mk0OHwX6U3ClzFOceu5u2wNg8BiH7rrDRZMzAxhJXX30RD+1AYzUKBbtMZt54jijtetjpLbN8i
PHhuxnycaq74liB9TFa2H8VpNqGkBgZthW32nRRlkXQt9lSSkOb3uhAM1msE59OV+oFCLtVw9/2h
kGjtrzzbvXM9TTcL2jf2bgVRqK61YxtTH70o0PY1Ar8GyRKH1V3urJffGA02w6GP8P0kpxwLor7E
h1J9/NSBGNkhCkc/5fZ6+kbrNMtdDXMRHbShbFuHeODIPhr6CPqTIcBQSPQbeQPompsC+Qe7ZqF4
Q8iYh/YjOfjf12yb7gv5eiELhZ/iAG24OFNpFLkaYykPYkDFqd+aYotvofIJnkwhuDygw2g5QfVc
JPJ3y/nppjNxB3RpPUuNnWSa1FU5l9U14JOE+sdXh/S5HwjsFaf/GlGfGnaQolDbVIyXhKC3yyD2
X7gj+IAL4rQbs7+VDSq8sUQWqZMv/fSVnDtpOiJmmihXv93KIBBNYx6KMc9Xs+fe8W469Xe82aPs
9gNDqePn8Z+3tfiOkP3vIJRaPNXvkQ1AJsbR+LAzUPOElJQ8PENZ+O59OpJkaaZwzYjoCb8Sw+ws
DUJTCiR2nFCGniWP107zZID1H3u1MhOEhAn44tNm0eO0vD2mAjv2Y476vb+NLKoRWfFOApT53Q1N
C5NBMwYi8eQJf/VmulTYnZ4slQ9pRR0AoLHWWjFe1XguU/V0NXlv+YJFBfEb8w5mDs5JCtjBp/im
sjLgVa3Wo03vJ3pUjm1Obtg1KgrgSGbSgEj2ixPLggm5cJMiXOIDkuLaNf5CNxZkzxbdneUiF9e9
wOcrPSyiKAqNsDPgI4cI43HRVbQSWq0ulivt6WOJ1KkL1MjzwCAHVPhN7FMo5vTF4f6+myEk0Xgo
vXnZW4R+l3Tk8tgAQ/7qWq9b41c/xOED+I1qA7jBNe/b0KAXhDaZLSRsukX29/A4gC+wbfx2mqEs
MkiZBG5rdXiw6Y19nD2wG9iwTcxwn/sL4CzX2TOOH5a0HvVx0ICRZ1gpDMyDOfIpUKzlbk2C0zW2
YJ5uihVPT9Cy79bcBwapSRn9+kRDVh6ujuVx7mEdsaWgrfmBQzJ/NjNJ8BGfK2Uj+/SkF4Y1jO+M
U3fQ9poY10oAyd5fMy+PiKTStnSxCIXUGI/5VaYPGCIF4+xngfJ/6RZUpeWp1aU73GncNPyX4b42
hv4HE2+rPgkduc/tVv9cvY7pnXzy+FWUtLg4oyJxBTDCmrWMO0WLU+BOY+AORPzTKMk0pZ2goOCT
LC44FO039OF+TJbER2BGtuyCoY0+H+ppdbOEaCM7Gr0lSP93ait/EMaRGij/0j5etM+8Xokbsde/
2aegWWkOi0phjk8lv0f8nfRBAKnWxpIWbed469P5JAyfA5tITXCIDWNOVKbCesL32RVyp9KNAT+R
OfGOJY9DZPmfJohtuGIoir3/CVG1MsAEtUIg6pxDMn4ildxMLiPO1HMijOnRzOVAQxbYuYWHLaSY
7HjCLPDnF8JPzlQql4PvmRAO9Gc0OwwfsGmkukfZLlASDcv+iRY+L/CDCJj1zg4Jsufb6bhPTnt+
sEmP4/748wKES54e9GMMSrvacowbdfolQTHnSfaBcS9tOMxYLhsyhemhEzYUnXpAULEOkLBz0xmT
VzNCHALdBggerghpaNsx8OCTEfsjSLfWU/TBw0u+reflL+0xgz29S1UC3TbdL/ITXo/anjW3YjtF
TucCAhvEoRpUteWGwAepeVPN6p8Qze6f3VsAAnPh+n/Xr8wvW09YbxXZmb9GCUOpqE0wHMHNMRzl
O5Khq/0XWJvXh/eMZFkFhziqjQA4HkIGgwS17BvbayprCog+ZYm9gVy4UBmUXcwyAYQDzMHWslYo
js9hxHpp5EyEU6I80Dn+MUWQSvIBg8hXPvCi8LW1MWMwOYoarNOop+wOh8aP48lZqRquSbAtkNMf
tLOfA31oiLC7/PDGj+feaq93VH5B4045AT9l0dyzBSRVq19XPBjuIP+dSKTWVjFHuBKN2BBcHi56
zF0fKRkVzDLHs6E//hHqIx1odbquiVpDHFLgmoHvp9unuBYCj89g0JyOUA6GlLv8kI0J7KsKfVDh
Wwm1jmT1z890e0m05doHWvSpX4yWezBtfZ6rCroCBy88GhD+vNf6JhLFYGvB4Bk/G1rjhySpCvhq
KEyI49OKoBuTh6mk287ekNmsK3xNr9keUDESxUCLHrggKkkWNGzTlOeEuac6QIGty8eotlOkiuch
P4PDjSgFzrdu+AWOU/NtHHmeh3MNbMUxR/kvt92vcJ4u9vhC81MLlh332VoNzHulVApqsUz9c5xs
BQdBVHd1KkaRnvxp1nun8y9za0CKQdvpYqv2rAcGRCrONjfRTJvtlI3wOt98vUudwqte0JKrBDlz
wKLtypYg4jLhRUISk0X0nPQddQ4aBRcdImEIp1Hl8amR4I7pMpiMYriRdAccKziIEiUuBTTQYjaV
O9bQdzgv7NzbFlOqn9MdYAzDyHjV92lDKd1lhQLyis8lr3GLc9lKgcmsbxIPic8LxeYePsMsi68L
NKGOaByJhXwjVardwBErX7kkSuLFO2gz+7l/Snr7W2l2eRtEg1P/WLi87BRNe3zqmebk578OgcpA
QCnHm0pwhaRjmYE1UAvyrXuOTGnervgVMRafOOZbfNFJ5O1qkM1LlvUAxOAcAdTXv9DTqMjgcmtt
H93nn/ehQSVXGRQ8VGA20OHUYF0FmoMZRsRdyUPrqxF7jUD6BX1oQPKPmiJHv18SLoLfaRydU0S0
Rwv52kX7DCI2o6JCHMTqJo3CUxjwKjeM4C24Y91FGp0o0PrJk2c21uRgUJEzWEJpcnQjoethSgVl
kfEZ/I6O9kcK19g6K7HmrNHlA5ynYq5FSyRvqXOARqwkJ5m1lWa3AFAKrtkhahFowIXlAKbfRj7b
1rBMd2r0WBnaQjP5OGoA8I3SKQFPtO5D85K25ezR5cmh1JywkaGiYREtwcBP8deicrWoe9WKNR0b
1FWbRW7+NM7qRCkt4wx6wL2apjJSkUOGcO0E784DmVNaixLjPxSkWMID/NioCoWDg7AIa1aCjIRk
x+GZkzO9kcQCgtCmnCA5Em271hgetEFwvr2r7wk1fvXhI0gqgCmcIkElB/5ejZf1Uo3tm86YAIK+
CT4BXLita/bKfXqzkOi689leGdIwfpkCOKtl38pbEVVRUV6jcuuAkxQLoda5WG5DNqCAIJPd8GNc
gG/9ZqEvCp3ger4fD3Apl7eEQv9a8f8GBUwgJirBDVrNo8XECWQHgUXUcoftEqPPsZJ0pDZfWxzK
4ksbgx52/uKLNfDWos0gYAieZYS8l6Z+UQGg86OkKwlDlgK2oRArO5qOGg+XoyHzH4MZBZPOc0CL
4TSuwx8OaIlDxYkRv6GCuxVLIZgNoxT0/7GmP/QDzExmlNvfNZ2R4NQWipbeHBnmW2bD+8Ba2h0S
w1Bpa7z0NV00Vr/96znyP+URaeXZzubgtjATdKtOkMuvIPSLImxBVTs2aNRBd6dvz54xb8y8WA17
sxZE0HT9WypjDyn8/1JjRNYjemQLQvdcLhZ64NJyaWfVjtTV+r2Z09dysBYnDJGVq3yqMViG/C5e
UNRHZ9Ux77T+8cayJpvInaRQqISl0/X/gitxqjJlUkbr0RaCMgnQT1atSWb5AYI8zpUx4Ow/7s/D
5UchDaJqxhewWsGYCZZtNGfnwG0WdBGo00wKR9aMUZ+8ScVWfDxa25r3XKc1smAtEYTiqACoOnZV
k4djYT6iet81QNohkiEMrxZsVdwNAMaUo/bl1111PDprY7y4W5/n7ujjiPOu6cIIssk4zQLrmyD5
oclXGZNPr/csdvELONXH2Msjt/zM6RcZ5LWaBvvNdNTswP7E5PAAJVCwmarwE8f+2JQo2gtRmGLg
jiFzEpzla4sv+bHPEHcD8mLSGruNSZCWUb/9QD2RG7y6GUb24XZKv2chavSZT61K9n50/Um3tWbh
XK6e0naBiWRVRxhYErxD3+zG1Bd3w0W8MtPVmIjchLb4cIn2gLX6NO7OTTmtG49kkcm6J/9Q7URW
E0W2oDyvaHBHWkAH2FtBnZq92sgpG4acPp5+bF45sbmhqo7VW8QqkGuzBWQgen1Nz7ZhbPTL7L/K
UahD+SP+0MBqJJjZDr/2Vq+nZ9dEvSFRyHkoaMcJNqUuIIeSAJZm2VDT1AoRp97JZw7LbHDKPGYC
zQGH3zKBZ2LBZPy0rrddCSfzd7hToc5UJw9p3Z7hfHWjkzk8OCSfIkhnyM10tN4mDAmqU5c5+jmY
SU+H3BiB7TeymG03ZueWmfJmT+cQ4DYWThdwcFcYuo/VrLk+3/9S0yJmvjc0Pb3iNDh4Jd5N5MK4
qKxwvrjs4VWA13eY/MkhQXqoq0VJL54dm5Cy08KErM4jLVhKcOFWKRBCXmB+rPEJwR+zMkKJy1YQ
0vXmC91AoN94GFwkTsmJHIZvWlPsTmn6m4LT4zEtz743/JD3qWy107Pl1UM88RmRcuaPa4iBzPDh
huF54SKJGRSA+HAt9iSHruKCfQPHYJYg2ZtZtIct57EOkJ7CD+Nb4OPqFVpDfcWF5qCwz1AN3O2I
/lkPokHNe8IN/GHSEidX8AwuS7TxuneRW+RgRG0QgVCZcF+sfKjFzAJHcgMg7BlUfFgnUnc6VuTJ
5YA2XXnDKGHpWmyPELEbVM04F+f+DlHDYTBTFp0cHWohnWjxJuATLakoJRPB5qiNIMjIv6KbUYQl
J6u9noZFMn/+cnRkrsiVv84IwIon4wzRbe3W3a1HMT4411N6Lrj6SVZs0IrTrn/QXo4ByDYoBtGu
wYUFu08yvomML5WUncY2V2jCBe2p7vsPgsuXl/9XflcpU+npFW7DkoFFaUmBXfV0Lz3jSoS6iSeS
4duPxvfBma5NbzF7G/XVJIWXvFQq6S6Rq+54e+EN6Ua+el4MWucuYcApLr11JIGAtKcS/FfUg6vP
oHnFk8d1sC221icnDYYHyWpIERvCgmEGGuiORD2pnlSpupRPcCopNdjyIB9Hdip0pa8mpaxXtxYb
ZftNCOS1QwmBaLZiDDOGuGRQXSawyWk5Ke+zOwpfvM4KuSb5ujb1VS+cezQizHdiZv1IoQfqUhoj
F05qD9OT51AJZAXc16j2m+2N5X3PraPfAaeOCVbyNZ2PqAaRKN5bhDMe0ZdEFSm0LBmAhs4r911p
h5nlc3c7Gfkgw7ykjlUY3lEOMxY88x+c/HhhRh/MC3Jb27B2j8hKIQD3+0rCuil9WcudvLBCDICw
S297HB1Qu+u7paQt4b+zBDfqt+Fxe0metniNbilDLyta3xMUD1z/LyjvIGe+WbeXd4NTQ8ifxkEa
Uso68OZaQowFgiAfH7UHWiGd+JAaBXokBANszjaDi9XTouWjIU2CcT0h9DFds8s27p5sVXiIJWHZ
7j16iAU89SZoSxzSUDGp4CAln7Wo+vretbGKbavmRnRZ0w3D0giBmC6VEUDQU6aVLooy2UDf8iVz
nyqbNk0lb7anJWm0BGMsdaQV8lfNLQwRSTt8mR9AdejpMmpzqoaF4gyVNpzHnClDOCuN228QcgUK
PXkvJZWzuzO5oiz1rgiY1rhGMFmqHQNOJB3aObI4BkAFyo6/jmcMDatUeCNosiX2aC0NIfo9rhoo
JUlVqhfs50H1uoJx9kw9s5qllME/LueBI68Gw6yGS+Oj4n7wyXUWD8J1XKnOSosRk3F5bgKSIJHk
WduAxhujiuvmB93rrNFlCHS7nW/RrBwBPJT3SB9wlRH+MLYQGonHoVoxmwHxkEz4Z4IfVY1DBjJL
JQ8e8mXha4HQdgIvCQzdVKphoOppEX5PMCc65Zyf54c3E6JJK+GIOOX6tSSgDuUvNTnTmjdgYJms
yMU2jw7kgQUq4RQAexdGbZAwFJfmdKDk5aohTYpjKFnyaLcVJkR5X9WlBiNIoYNfCQiWbmmroQJb
EVJWsovqL1khi1fz1dJpXmTRjwvk62IN+DIqFxdUPyMEtJBa8PyjWLLCEaecvob42p78yOjMsbu2
S5aUei91er+3AlzejZJDyfjO5m2dC/a90/n79DqRGYrUBiSLdZe6LsnRFy2pEirQTFLs/w3Y3LZv
ubDqFqCFF/fB7R75Uwiuh+fjx0347zYX/Ws/27kjejRshorIMEIlhCi0quW7jvnZqzn6uVL+fxQ/
w0TbGYYm+I1WDIwUKHpm3JGRmmdIT6I27W1l0LLMv4LKrFPds6m+ZEfGbSwdjBfbDE4wqbKRL78I
zXJH9CKbi4J3N7qt8GJt4gC/ap30/61fjEs5zYdkcnHWdkGohrt3OXkROvTpjvT4YTlZvRBscRsC
TsIGTUQVLgeFaT5j0TZJ46gyF3CTafFWoKWvUdf6bx8W2W/W5AaYmKh3Q9sUWYNPVwtk+Gq2LahH
r5aA93DAJwDTlxC+rBSIGhJ+LhSmVNG32q+EGHP6Q5oyoDoFxzLW+/O7MdQdm4/KMsOkfuSZ8GCv
3wCQ605rC0PtdCpK/QPy/HhklB7SSKwgKx1qEIjJp0RW+EMTf49kemobS/6M9SWYsJZMiQvfmFwU
iOQIPaDjsI6ideCaqH6SOonWpkyUqCCZo/GOZ66+E59LqydVNUE3/tLOlkzl+7KadmNeDTVTXtSw
ERvIQc2u8EAltou02aqATsM8ZXO/3APmrqZPyBMjQOqZ/cb3k3SA+klTTjWIa+UXQE5smxc0+ErQ
wlN3Z8C3A2jrDmzzneF2IGcLcFoJhE7N/X+Xz10tatAuH5tcA039AITpXqZDr2FF6cHgj0HF4QLD
LEBaNG1DU1IH/lAjm6UhzhnSiiS3qVRNivWhMaEOpMnsNIiqftFhfn8K7aoQTXk00DJ818AZuVNx
q8tAjnf/Dgx5qXWeygYDNP3jiX9I/fr2uBL9VCfXWv0csWI9gmxwXCccoqvLPLf1V3mED5xTRwz/
1KjVryz4R9scbXZWCymfiNnFC5OsYGAc4fnsUVgwWzIv+9BmR2ppdjDHD7G50Up15Ld5qtt7Hcvr
gbwLzpbtFouiqQT3uf46Kh5Eg4jxrAXHplGidKU3vBpaW0gm47laDuOlEp+yOALUFx6MyYdS6bBt
uOP6MGG7Idct6TqKwpd3WMFajKvNzhWfuY4nCBvwad+9j7mxxxFAp6YvYAlLQjaT/cd9kkBbweB4
vyPqLX58UgQggmkGDyjiv6lPnHbyykmDQIC3Y75lpl3cWE9ABktgFK7E0+COZEMvVPVAnSKMPKO0
uakHZtphByzeaJohFSIid0u9Id1y7rdWK4nZB/CQ//jJ0wpBz0FCPFhD7UQ9UPC67V6JRFzQSjvn
5RdSlFeFTrQ53mGfljklTaPY/L7eFJWu9JBY7xV0zdOz6erwgsU+o/4Oz9S3CsUdriu4CuboBwCu
PEL2xb5Mr3QXvS+xPe8zTY8L16MRCkPgEU6WaH4vjmsZktjEA8VwGnPPPqq810PM5+UX4WcSCC5o
A1mW6A5JRGAQ7KwqfGCQjQinhA3ajnNi7cpKvVrfRWA5Li+uwY3xCJDwFvMemf8hWZY8J82yGxZv
KGG9GwLVnjQ4dCHOVnJJasezqbOLJNZDL2o4bv5TXSzPtcf2SFN2oTyRznpF6EdQkDel0pGaPZxe
eYueBCPukzv/lnw67fdX2KG1yybbrX4xJFho+pt2ESH6Mv1ya70znQrpHVljEQaBuIC5Q40rQZMz
Kiq6HEXXCL9qsLh2bVj4H55qgaAiJ5pX9jQvcmYQrangCG496FbprOz7yLRF8nJIKDogC+PrZB3v
69+Se/E/s79amBZjPC3gx5s3QbZfngs+mwdlDHlCkNG1JT9f31PP/6kiU9kSbdM6vmPacu1Ibuo8
PsSXrJH6ikHfpUq7uy9iVEt6qVry5k8FyqWY21GXuf+4/FuGvUjQZVznzCWY6QOGPDEk51HLrw+b
44TrTZ8Ad1E9zZ9UW3y4yzv4tjYCJalAB7AotMh2Kn9y+9Mps+RPivTR0/ep0+/zGxr5t9EnMoUG
jqop6U3XNPH+ifZGGMEXXffEZwq4GgQ5/62s+I10QvLwSHiuf1MYYG/L52Ys8tbZkQqlfwc6uRJe
EsDJ3NCWNl/NxxklrOWYsv9cU4k/w2wM+LhS7ijLKc86NomTApGGzr55j2Xk/02H29qWxRz2FrEL
gow8pDQnidAp3JMy3iTe6fMFc+ip2MtQa+SakteCZoM44qcexOT72oU2Bkf4Wiu2TChVINbn1AHp
qVhUL/mfHm95kYAdXeSG4pNrXd4W7J038pmFo2EmDsEiIddIdBUvZCItBJifk6zBBnJvH+c8RR7h
ercgdlhbgnrkxtHhOWbRcwwp+a6s4xAliF11zPtnxJ964yuOXLIij/k1jQ6ThFvnPERC4vMbif1Z
7C5tcXaHIJ45BUIqnmmCrKjBti2hss/IcPMbP3T6GuPx+g+tJaYR7U+dD0URec946WBA9ygzkXpd
floRy620zXHvFKAeEJpcpeF24Ni9rdxwv0AGWpdM0CYwIA2iioTIpp9pJ98Dz1LSbfKucMplWBpk
SzekbDTqYClxOdmmjAjfpj3Am3Rhu36FJsKFkgIL2UgFHUJ+Ab1owbva7MPitogCay2IORd+Npdl
JNfkip7jaJM0sJrnmsxOjMtkhx7gwM5g4MeTl5tKCcCmNQwXgVoeWcF0fcjN8B14zBG21uBniYED
vHrWWmBEk+61DKP83wPy9BgMaYMHOdQdu8dLUVWZUqMp7v2BiqcyWJJT2O6oK5wQTLtpn19qNoIA
I160JoeBJEeoBI6F+0mE09ATLqjpSji9inu3HhXeop1N/iNXm7RbSpXngz/N5I7KFaw5HXJkb2YP
YfdCHQ8d1tS+qunderZNl9UHvtHJAYyG+cJMO8yeJTvgC9UO/Q9tj5IVqbJ/TtPrdtLDngCKR6aI
u2y/ErNMKlFbVrL6WRJKnfm8Q8fpSrcYJSClkuhuefqn/m5/0J6xzHnYqyUTPVVkHycP8AMBqi/j
1gl5Aeral1TIhzZts4BLQjj2pklEQ9ugXw+GmRy15rmz67pkKdpaGNDFameIKbo5lmPXxEn/l6uj
AR5zHwZXXvfLXVW9n1N2DqqBaxGU+vGjEFVP33KYJw5wTKMOM/n2fF/rA82aZ0+kb5fPAyW9r/w/
nzeJg6uMn1KL5h1bJuX8pBeW6TDxLqZ9rrg6ek1p79HaFjvynWfms+vU0yci1hMWT+YnCWY2AbVL
JVNU2zIvDzmUrhzCxYeNDKEeImDsfpAO0LtjT6XXU8tGvnNg9zx2/Pv+rMOGuO1eVYsuJiw4Eq+D
k1myG7BOckIr6seD4/39KNpHUvVcgu+czH0EPDQZCzlWENO8pw+VrLoAUIXRmxqsVp7C6Hp4I3ak
N9NMDJuvKJCoqlnGPzMbXFp6h6QXK/rhxjztJSamaQmCiq1bL0cjqBpH6GpU3VdtM0QqnGwGTc3s
60Y0IKKUKakBTnDy3p81KJrU1cxRJLpHxR73VkwjdlDzNPE7qCAhjbAMN8Mh3FPRiIA/Z1a50D59
xX0J2FDyzJBmxbiIucCPMJSMC2aT5BSJNZg++6/9Qogvaz2DHJKSUnOWpd1az/oLI+/Nvc3i6Z5w
OSpwuGmehxJMjbrlD5zyHfpsbVfBUxb8VhM5WAtVKZqXmucR6WaOEDfBpPi04OqVlac5SXZPd3LQ
U09EmveJQ50njskcGZHxRMOFw9Wf/b6cDhIzCOEl739vLi37koAT6WfRN1ns5XNTAK+G92k6XErA
Y3mipGXyN7qOsTBPhRtXp0BuU+pOXBD0JdwyIBGwckrL4+6YF+GKKfgrG1SI5fNdZg5x+0y7v71q
F0HRKOFiYF/dt3ecdZQkYKS6PFk5+vsyGDm6+Y82+oLV9P8ZfN/WVFBBrJGUQChOuaWw3VcFgEUV
EQYQMxH4ZfscJg9ACaElDHdJKwK30Oacq79JFMk99oReuuffR30vPsrJQtas/dULJ/e0beQhntAw
guzpJpbE0ep3YpC6rWfHM3CK857Tda8WfK0+rDsl/SL27dVCeca3gXONTCuGW+/boN2ZTcc6tush
FTJFSvDVzUEDx/YVN9qBKB4W7AmwULDBs6btnD1OSZsaEcX6QvUICt5xC0eTJfn72s+b3/WOjvTs
C6YZabpoC9tsp0iYn2IJUBXn97nRh5fahanJPo1Y8F78fpg9NbdNqC5eq8MvArt0HrrWE7BzwRW1
qIMLhlb+CDqvAu2EdlnYj9a9KxYd7InO23N1czcNflRuYoLtYVZRrDACKxaiImd9y2ZzseUDbbSb
2wOn5+DuN0zIL7bGmf9LPv1VvKpl6r635JXKCyliU/IatRnTY+oYP8tXAThxWycU5QWhV67fmdRH
TxEyeFSKJ/wJM4J0WctjjzPlLHmjOpgZp5Ah109RKr1YA1T0zW0uuUiAYNfK1RVDApg68HPeu/XO
eibYbXgLyFJAYWWJ6eNARLgDmS0HbMACpOx+opuAIS4gArY0lpZBlOY3Xf1D6VBfPxmYBJbvilmM
GEcvxHdhaEQ1may61qcP5FPt439QxKHvt76Zn2k092Mo1+JyMAJIwJwsVY9d6u2HTny4aQLFo437
kUJgxNMo52VGPZ/0oxUlY5X5usWOsFoquQ25hzwTI+vyGqmk/ERgruzz2RANkbnNMZmPvesenG25
8eb0Pmontq8ab1HLKKrwLS5zXs3mpuBuxCERcyYgoktEJRUS32AafqmsVxT7/cISrnsZS7UVEX8X
2Bb/KmcfinfEh4qGQV/MJbHhbtr63r4Z7pEZOb7473lpMB9pqd2VS3CxfSWe6HAMI6xTtkgu2+r1
yCIVEBOBR1tJr/Psc3R9FdiMC8Eu+WztzDFCEXFGRZ0bq5L9dAJR/ohRw91XrLFkBrh87EPkdvFt
g0ww9roaFcbUDHmu9mxr8pG/GZh2ZsptnkZ2kp8Nv9p7AtoswKHXMrNnnVwWL5aeU+oprjd9i96/
xiXkFr+tPgO4jdIf893uvULxr93iE/0xqH/bwIthsArYyI7Hf4rGO9NPKgUilXHk+x2yM54HfJw1
HU2lbMrsB35lrWInwQCbPPC7viiLfYzOkxkuvNTQm/zeblp9jB+HGNNETFGkpUlTXWOH4YznD/6f
EfgqrWrYhzGd2DVRXd6coQXRTeccz8qWz/aUL6a8Tb46zEcQTakJT1vwSoCpqlO2jxwOns+3lbn8
dl9FIAl4XHHyYvKf6L92TH5DUgaciW/CC/qH4J6gfyWBJ9wv6DC+ZJJqKGYf+s7OBDA0A5KhCn++
Z4m0H7x/c/mmgG2aZigozeEdRRrL428yzzW4vJCznTloCVVp0dQz8szmfOnVll0hMVtbFlHy2hxW
9HEL5a9K6vRgt7/Z9qEux2f+DD1vagkTO94+Q7REiqimE9NgxhZSmwNMS0tJnTKT6f3i0ebZ+gzM
914akaoyZ/+rQNusuoNXdBO4wJX/y4ptCKBHa+1jAYJTixwmnGzQ8WyhxSSf+5nGad35+whkHGbm
8nHrIvewTSLK1qHJTVm60fcqyo9o4uYpykWwF9fBm4IYtJ1r6A+xZXdb57F4tlqLtRMVUwag0HYU
k39hCUJ6kih+mt/AETopuWk0weYEGdluc4QHsNvVYTH1KvVMAMZ1BUtMbTLXNn0JHZMRf2M1RVw8
2S322WvoC0pG5PxDeLfaM129E03PPQrWLy5dHdw5V0uXZ6xrzjscSikaoe7mIHZWwuOnnmw0dncL
cpGxrL2frSJ0s2T0ZCWCnDer1ba2lWkxeXMWXByAjjEDOH7RJSv/T0PSAhml1HmpLachCoaWmaVB
YsD+TtTqvgfL9OUJve2SBihNJ28FWIip/AKvAlAVZrzFE/ZfF3VfN2yjOvQVQ6y9kj0choNCu5G2
d9HUxYlwbSDy5B4eC76QYkJCZ+OfPanv3jpI8TnMYQFjTHu/sWMMbYobsZ1HrgFgkblG+pvtJMeB
hzZ1zhlm31+qGqfEYls8CesdwJCM/kkb+G5IiU6dPiQ3SYzqGcrWHeCpOSzQg6kQRikpjVMpBaeJ
gtTDKL+OTJMiNUFYawvf7oGlJd/K2b0HtAk3NOhD9Kw7ZG7mxEjh5Qwj5Ik0EKbzy+tjkfGRSmJ2
rcaAPXX0zSxNrvfcsps7rNbkfDdqgyr4CFrFNmbS8xcsmeFjun6S2zIIxnuW+Mh+qsJVdFwGw4eX
6eomMKxQcQtFfdxhujDRNwVVp+yQGcQR7M9p2yjLFr4ZgqXA22dpyFnBJffhP7hx6yl0ArrlWeHV
4dXXUZ+Cc8Jg39cfbCIy+iuT9wuo+sF4UGSKU+gQPVaPWGxrKL45VsauA4GtqPKprHfseALVlrE4
M/8jOLNcLTidOgs6+f04Pp56RMOdixKdj3BX+E1Yc3z7Uy/kRf+v02jHBFhmBchvEtYpW7OwWHRd
/s/EVgKhLaampLdT+8aFYa3Nse8Osv7Ij8fjd3TobD7W1/oQLUkcBhKoVIO7E2xHHtgKwThmeXMv
buRyNMXqujso+8u5cselTbwOT9iGAOvWLGACF0b5SuQ/6f6Z2o1Kaxm0Gs1kUDHkrCEuie6uGl3Q
cMgyrDdH243biuWReCooOdJ6r4dzsdb+c2Rf9k/8wSY6bATI2AYMouXaqM7tIqJMskvl1apNxO9K
UvNY6+QOq0GmCQrlw2Avy4I6MSpSl1wLWbDWMyRdqsAy+ipP047dL4yxDs1/i4BSHhye2+ymmRT/
39I7veXJnhhQUGyHirmqyfKsKdOKwVKJ20Mz2zfOSPz7kLnd6lC0hgbBp5h957xiitIm24QUQmKs
kes1gHGjBL4sVEnnnYVx/I1wCjjQcEJVqbOXbUpYzC2pQrSvGcgeVH67aG7bC/8P4xKPApwhxt4L
prEDcmk5RDxalgaSK8/iqF2lV9kBTNCuIIe0jnXlf6y8vmoUXibRtG5R0YKHqQJC5euN123Eq6XG
wa2SCXoR9Qai+1hIraYARv/U6lg0rAOauX7lLme03NSXodSv8BBawK6VeOznzrqLkdro95Yk6jW0
g9uxR3FhZGsN9qwhLoMWhmVApJTwIH3znDF0YT5pvPDFBuAGCgKbu0ecdpHEtENtcBZmglvcKOE9
lwIUkcw9K0x9nzeRzo6UYjz1ouCM1ZmfEVG2WW2d/MXBOVnh2EZXoShskipdQ2625oRtAAm8Buig
dvxjGRU/KVO6wHq90gKjYhzN/It5VGM4wcdTOQLK0icMK/2L6gWRO4K5O50bfGajfLdp/DhHZHo3
/39MCYruCvotw1sAytnZBmWrpTPGEle33Erxo65FFl3cJk3OOOdioA7W3RMjys4pwp5teDP4GxBi
3wR8rRB23DqM0lZm3ZM4JC3gJL/Vlqs2tl+AYr32FDToSOuH9YbDGvS+bGXYclxDsAJgr52Ib/1z
Yg6YXayMA8MH0xXlF6uQl1+kJ2KiuBDGLpggZm0NxnmXgyAIdW9wfobX4dojSXHEtg/TsxZ20uki
EiQUGbjEoX+LGNgDmwP16dKX/TYLhYHzXciPimK9Gb+rRRqFpdyAWBG6LDfrAq/CdfLaBxYfr+CR
WXs9kO0+ljSy5/mgJvnrkxUSkCgtXWRwaQ6qIA+QDjMzTjPI0x4Gu2bpcbRSVu78SqKsSJjikj4d
6ozjaHfRBnUxS7ZeM6e4ERPyhSGDHLx2VTIkcxaMpKeY9RrmH33WExSa5uMjOlmKZj9YHwjpeODL
Up4bInLux8Upo5YObUZXxklGtmjpJSjs5V/sJEnBhQK7ChstPR5ICsJyKSsi5EJ1F4qWbpmDYc+u
1OqMizkd6df6BMwgS8JnXVudxhYIaOUMKTsKRNL3znaoP+qU1caNzM8zwIYDlwGBqt/3JLspwnqZ
6HKA65znxz9aSCwWl4KFiJDeX9njby8Bz/i1eTIKn2lnCoUe7WeksR7VurgfMfWY1fSM2mDqUsF9
PnV85fO1oe/aslUD72Pox8eycECYpmCCKxaxDggQK1qAAHB9cWObt7pmYfMu1hB6rbQ/57Q6+rJO
ifPtgBl0TGtgRebruz5X/VMtxIBmeOTtlFV255LGbp2L/xeHk/9UDo1vxDM+XwdwTXQG2J9XMOUV
w5Sp3tSIBZoNSQV3I1y3yeb7mMostPMa+2J9g7baqqlsIC3/7ceiIBSl4y00OWC5gJscWiS30RUf
SgBrhN9nYMS8wr65fiWnbpmXaN1IQ35nCRz+i22P8LOPnnmNvfK3FAYDXbzQNxOZTsJI7ySIOBRH
PoKMwUwI52M0oGRI4EDn/VfVbtTa5R71jLayEQKv2Uwuxc7cMhxlWwx2REr3HCfPW4dGaULbi8UY
RkvjZwaKVLV5HN1g3i9bH+Zwx8uQ1uGTaW7bRKmEPjoFCMboW1qGxJ5ZWjKdv4TtLm5RhEgKh+ob
d/p5DLa/UX7sM7gEMAp1mHTR91t5BfI5r8c3CXoqGJYwPJXtyyvimIkuO8TMigdkX/nP5GYwQJ82
UhscFDj0PKs+2o9YcaQqtcB9Y7rpYAT42jJYgldqlPbsw2BH0fQGvTlRJWTgrZhl5Wiou2GJdBu/
KcrmgVmaCWIQkKEzpLPy8xHhtxZF/JyT00zqRbgEY3sPLDF7mR7RABqhRWYmrVe36Wd3ulyUWawZ
WIbH+U2vdyxAOcm+/PNuXYKgu0RPUJwbuTSLSBy/hlFa1sKvBC51uvAbc3F+vhZTsNuHnWSVp+0V
HnwzUBeSG7YKiiC6Fgqb/kDjs+99KnuNHXaAuvTS2JGQiletsyNgK5yOEnSf+CIiHUb4KJE3Xach
IB0AvQcqagC/+rGDBUjPufh+PfoG+d9x4vDlZX3LgFKbU8nLn7oS3II5tFI6owxmXrjNyBZ8UwoY
hhmRKpHCqc+l82owFFW6vX5ER2s3Bc6CyFwXKLXxqnycR30MoAYKxUsmOABG1vwbzza360ayUgn+
FVtCuihmpVhbDGRGHWgL9awZNEsII/YhpcVDi1j3xmja80KX5zvlbEMXc5FAkVV4tAnMcFGw0aZs
GhC0cKVgYhEBtoJUn4Jp14S2lUaUYpmwWpHHkO6wVdnE41NRjbJRwl5pyTL0FhOvLsBQxuT2R2UG
fAFZl90umrhdjyxa2cJb163wc20VZ3ILMZ2ctr0oEEJfgFJq6Mh8PL1l24nR6oJ312VMn3OIXDVv
QKp/cX9YBB51V77DuIS4Up6vX4H6FP9XbDZc2Axzk80Php8hx947VLVyz9KvAeiOG/XtJiv1aZIP
si852Nhh9l5pVoFjHFTshDlnAqqnOPMNW6JgBR3lI6EcAKgd0g5Kr8Be07Fqfmv1p/QX98sIHV1s
AWosl6Rzqik04Cqtv/KYNXW3amY8xbAYVad+m3MBytXKt27Vg0lpvGABT7bCJ0w1WIwaAdAR2fJ0
uDcs8zZBoh2u7eyYrooeTm39zBrpsSZGnLXiv53RMYm2wR4gkVTsFYbrw5/yG4NMK71vZco4O8q1
O5ENXWgCNXDPpnvxLiwRQ/upe4lA3ldLO1h63BlBXY26FM5CmPTSne7zAHRZuAKo4fsjnEJPAbdp
Jki3uwZ4U3Az9ZzRFrUpHbGBouS4BRDP2EBbMgIwVUWbt2P7I5RfT7q3xY5mpIZUMeoU4B9smg2D
x4Wuy6/h5RnY6mibbnxH7mtv2fVue8a4+GAOBMEDPArHaMV0L4MMf10qaomDS/SYTx78XZE6IS8/
lZ+W4v2DsbT2gHLIRC+KTtNfMhKymiksAD8uqcmRLx6sNVsa57YY1DyoDa7134yKyzVZaq1WR5Vp
jbLrKhbjPNBI2EPz2izUUOmkZmPLo5xCEOvqkgFNiI/1YXzBndvEJZk0bkF+wcmLET+WRTKs8KNW
Sfpjk8Sv+yU9UyvckQ/k/rVvqhgM7nx8RYX/XcTG2FP2errz7DjCbbbKTa8F8umyolV43MSCAt8M
64svnGdORcuijkGm/k179vmXQQhS4+Fp1fWcmkLulyCI4OIX0gXmHpCeyfP+EPzJjKyAFqngpmXD
9Cv5GDogTqEJqsr/h3LpfYjR+SwKZgPLet+Ck0fWheeCMl7U0DFdx7QXFb4Da9ecbrWYXFtNHth8
MDpbU7UUsuqKue6BiDzmrj/R0f5n0e4Twn9P+ypZo7xN4Vs5DJ9DyNhRIa0D0DhDrVk71phbVFXH
yc3vDBtgDKl+YXpxOaiRSNfDdpVF8tOgqAzrori9Uu8KTNI96IDUcDV6b917dCwvQu2zPf5UCIIA
F0+jA9jXhM+ock6bUG5St6RgsZnCP57QxVHUFUgIObniEBXaXqnKSC1bQ5aqI1S2yEmcfRmTFovP
e3aLdNCZHaMt9Pbiy3Rl5Ovm9i60cfM3//pVbh8dVXMxoOr9xSoauyKDtsxwDMf1j3dLrf2nUeE+
vZJZtPI6DzXzIHC6XJUQzkGjFdVRCeiPyN0piObnLG6bY3nwkwxSEs8Hlq/BiErxE5NTCVk7noZ2
yie5cTb/R6uCdhwv9Zud+f1FSuJAQ/nD3xRUWI8SpF1YUzBEm83SZ5cnfWjIoaLrIA+jxW26XaA/
udt9LBQjmFACTufw7g2gyRMdOEgiX2M0fgOcrHhuGdXtp2eSJKqpbolLzmlfDD17n8XgX1000i1Q
wkgDxzuYV6ynOUdudkY0STJ4jecqJliySLDqGZJaKbaSbNs0l6EwtMlDY6DDWcT7X3k4mD6Szx/a
7V7sIQStIfIXwfAsMucXJsuOdbRFzUZGQUolhNCQEZEyz+nm44EINrzRT814g+yUgV0oS3p6VxfG
XrnzHUFy6VQbkwJXzQbCIYHnxqArq/D/SCZg554o8FsgXtYKpY2a/yPbEr756i8eloR74QF96JAs
lpkv7ZEwM+KrNbMzH/hQ+TAoxYdl0Vhbzxy4CmhxMSf44Um1pOU4lsS9fWj7zP6wFRCG9XR4+M4v
fufk5GueAFaUUtmIJETQ8r6lpxlr79ysnuXfK7S9q/Kenhk9aL42Aa2T0+otMdMdF5tpaI7dESYV
pKL+7wO559r6u9EDDRd1WNP5vvc61gFZ1eUpV3b+wYUE/RjmRshjkqolGpfhKC+AelBRy2XPY9IM
A4z4xDCTPQQfP66y0FZ4/tPFyy4q1geyoTytqwCXZA/ZkoDLjCycFwTok9t8HB1n1AZAa+KBib5k
XYAM1/EwzBJF61NfCHF1MT/8+lSJRMlhuJE1vV/dlacZYSyMhABlKQBJyHO36SR8IqtYQD1HPxn6
o+shDac+921BiPFXg4tWxUj4g7GolgmY+Kd9ScUqKrWIbhufNRIrkzG34J7B5YNnHFi3gu/t9K46
OJER2zD5ddZN/CpSP9U/hKJzXZ+p9IoAJouJtv3xpHrJ8DT2NRRA3KcNZwwvqFu+FqNecUQasihe
00P/ka009JPS5OjgdDGgtpjTfqYjsHaTr3k3SvqbtnDhvqzm0jj6lEIJDEvXZ7pXARhLk8kCfayX
HsVoOOI9Wxv5v05uFaftjXMc8UXDWOCRSKa82fvRIQfR3bbei1NS3Fks84IJQTtOckxOKBlVm7VT
BR9Ui0/UEbIykrZ1rc9X5wP8ZT8KxFoU3YyQBqA3S25qLm1pQ4N+oxiYIm2FSlvEuoYAv+tl6whN
BEYDlXECAoWp6Sj+SqrRNPB/JOjCQMH3rqS9q9rASnQV7UM0S0eZEcMdQMsnP84G2Gsq0a9xevri
Eyef3KPH2iptZoHeKwxFS8qoG2NawQhipA0G/WRzPX6V2dgqcKuAnVcSFxyBWdgC7pDCeOx0Yba1
9/clS+V9285vk5dVWeUb3OAs81ZFe0PPXei9+ZIwWDAibuMNn4ItlEdVIepHgIvuKNzQQ6mi9HTB
q0hCir1Ha8mYxCQcyOwCB/N72jh52ulRHbkzcRv76x1/DGvj3fKLRlhO+ma9y+jQf3BymJKeFb2c
ekapfr01mzA/uhdjQg6/YGDAlVM0Sy/aEyLXWEpWDjLX1yHYRBWAM66YCVUu68y+BBqtHyrV+Dyg
oytGjV46hOmqFQoqa+7Uiu1eflRyLYlalRJGLj9dM94XZIzmdf/+Wk4GZkWKACQBp/z1P9MoTYN9
rg5XMaO+f8+5duFuKQ/M6Ys+YkFWn5sClClNN8jfLQ0xmKyrBcLESsQj9tmvEZQKnvS7Mr5QUpDl
u8tfG7pdWjnWcwJtzN0aIEsTKsv4Ou0vdWbAK/pJgxNNtiK1ELqrNH6MmerfoxCukWJINd3S190l
vL+h8XUpWMutBIGpui79VF1gbUlrVIrwb4KQdGa7+GTcAGyL/Xzm8o/+mEtHafHZPjeXdmsyPBJU
6ZP4/yQZRblJ8gVYyfXeU029AiS4g/FC2jWkYFs388/6shf3iqEi+DYa9Or7VC5rHlJo6YNfj4iW
qM9u+SbN+tjaypwVnDKzZtstEPg25ujuDO/TrvIQVGyD60wPiCMuY46WaZkcmhc1AZzCA2hwrIyy
IwMlUXEtOEcPofdUrrYCAnSPm5Ow+VssAkmgsCFdL5no3wP/jLy9ZP8bY+4flL5gz7JIslSoNb+q
KqxneHBv2saRhmu+7HM5NAikBNpYyFk2uCX4PPOoMHUuxrrfoOxvPLwwkG/fVBlZhVXy7YihAyHa
ycRGKSlQ0We8IYDpi5/H+z7bYgQ/72jzMgWHNc/RmlEoJFvCm/7ovZamFrGVf4NCBWrbmjMaSJfG
H2mY6Q9PBrrxHwuI3W5cyHlaGo9FwLa6RdknG0CySzr8/WR8TyNASWTnond/sROeS465gzymFxTB
8FHE2J606dSa3nECxI9fWikH5lnmB+e5mGtNT+2rcHryWnGvD1SNoFKsRrqVftqi2q+fVNGFV4HI
I3qJ9vA4ANN9GLDda1W+NX+9FUb6xnGGL9dxX++kexsoDGKxJeqRWgtQQjEvYMVfGR7Cvex5kjpc
vV2CKGl2LHbhJXjzIBrvWzA9oYv6iluQNtrwzyZGlR5zELGmk3xirDGvunbN5BHbJmboW/cRStg3
XTxJ7+tKYU6YoE36G427/bYR5qkjYFFx9pY3TjYqTLAG9nRwCIVoB3lMu4m7XVKMmMLe3zwGNqau
r0rPxf+0jqi5E0MA8MIcHOzmiJy6TbkGGkOWjV0W3PdklMb7j+/PqS586jzDJMwRQWq15QjGp6O8
RTNue/q9cW7ZBNNzcwsw9nTNRQE+5yBL4/xYGlQcju5f2lELAuaL5jAABSlUFX9ixo9+0lUGPUPK
W8iIh8cGh9jJB3JunG0uzw7LP0ThTi6yAqIw06putNJEnPUeZQHp2o9Q7tlN+pQL+ORXIfwA/T1s
l4SDWpOiFt03uoHokvJk4eW0aiP3Nu3klp99a44ZaY9RcrZCH+w5vBWlYDJR2RePT6Eg1UkuB83o
+IJKWEjk7li9gLvBktxhaHDaKl7wStFcol44/wn/8H8wgIyBGotZrEzxN8tXgVtaN2Am3BWyGuBf
OUwpWPBL7/7NPL40rrZ6VhiaLy4P1ot0gYki9OKpD7xZiY4B7eBFEJNm/6DO1wolF3oEfNTgzNdM
554bqPsXTPLObnoLEQxJSNbgdlH2gliC2gEXCHdCrkvkFMF48hRjB4+nxh093TrpiDIamabDaEsl
6zAaS+7270uGGkrK9XgTBwNWvy/5ot9gsoopgvDCl6jQcArNsDkA5g6p7GkwIROK/l2/lnM8pC7C
VxNLThHuRqu7zSaMA7qCjJmFMo1hiYXlqVu6tJzM1XjccQYMjGmAI5D2ZlhZHWK3rcSjBQd/dOD0
2lmzJrsATNxswKjzx25BdVHsAuwzlSwxGuQqbWLrpivV6+UEe7sr3BHH8tU6Q6GlTEOwGZIGfLl1
vVRpvukcC1FMCbXuz9bV4GrG2vWvnPyE4Cjygn8LIEZy+UQ5VYVUSNH9kzD80GMa1UN8MKJy/F1d
RQdlv2N1Gsa6c31R9TH71pVemXMawHlDr0i5rnXAzDnODIMUoJttw2TKsJ2dDB/v0vI4j4NN+Vy7
zjl2oTnQwCJfhMpOEKfojWUY8KSqrOvnH5qCv4YOCSrPTLSFrcIprCtmS7KOoTbio5Jtw37BTvA9
H+3UyZEEoGaCB+eO98GPiOoaD+2V+fGaOIogcfMUXOo6Rwo8cuAPUCAAdri2HuvLaD9tC0zLfHEz
wymYU2dGyDtFb5Q5qf1jYepcm/Cob7fyYb8vPd4/IEUKUf395+zgRq2sSqbTtzspx+LvAaFTLEso
4oHvjMWCPwzot7UEI28Z3tCAt2utpvvjny4oApCvCzS336pv0CJRDOfKB9NEHfsCjF4bl/uPDppo
FJA6wr1Lq9VdsF6uvuQ7HE0Ogwy5jr3MfoD6J9anzC7ygegs7cWPiIgXbXxTSe3AZ02xEHqPWyuk
JvOwIpqO5OwwjsB4Ek2T1zVG0LY5vpMgL6wK+5SMtWb08FSqDcRfwi7NdKjqzwzRzH+uMCg67L8x
95GEZiL0oD0WcuS1FKYBC0sRcGbloX4gSD6MiGk5mdU5ZznMkyd8tsMFWJ4ms3YSZQPqlFk2FtyA
570N+ezLdPv1c3n7xA3NxaSQLKxaH7aerpNYAngMXBfZ5DkbZRjbaBTRSQLW79UBz2QnZiS5JZrL
MyD05dL/NMWJjJlJf7T3xSQg4rqAXr0NDDrZSyW0v6IRUcLTqQRxkU5vs25Ckp14e3lKcbNxejJL
dBNeQwt7S2XK70pnYwiKgUEr/O80dovmz4CchjYmYH2WqkyoQ4ZHal8ATPjeLHoazNDdK70Yl3Hh
VJOGlUe6tinZ3wvKSXtE44gikcuI8X/Dnu0ODo+IelwBocYExv855eFk4ncSDO02OoifsAn6+s0B
6UW5nrpjE7HdqiSBZ0V6lPByZ0rn+ZU/i4nzTKLzGUeu0qo2Kdl76lKtELefgYRXMtXrhBAKSG1z
akNi8vw421iVtTdE9awnR0GfO9U+vtSy2kvUVywVqFTOWXhUrIfiIk/NycDx+PYEftj4KrCzL1Ex
uUky8en1JD55lFWh9x9LRcVGdLfhPyS0V3mItZ1HO3GlH/FCARcWO1zRW4XuOHCXEaPjnWrA5glG
MzjQT+0U7eHtywdvaA1cpcFolFmV5Vvcux7Z4MXfwadqUFI1FNm51V2Hw9gV/ImheUJVRQynTxpU
/FtQqVXlfFfXxmefgR7od83yOTbn0Df1CTvR+Lkyq/GUpU47wRQrm+kFT8crLIBsCUgT1o/dOKBd
PbapdkmtVmCQVU5cc0fMSXPd2E7mHp8OnU3OrN7p+KjRBPJLHVtu8QrwiV85LUb752gFJ9PncdOF
ChsUwUK0VJQKevgHUjkRJcfV/kMgUnokO2Tj4AbqbvbxTzVUs9WzkIETtq8B/JvAkkBKMQq8lyE5
N+Umc/68Hdq8NNpOHuIDac3Ea69q9Vb+uhwIvELuwIGEtQTaxoB+EJC1UQpFgFr/r8z8/UDIggpH
t88uSeKI5PoOJEQfhX6a9CKHEhqen8/NQMEPGrNX2IrYyM1ujsVLlELIqdLgwgmsbGPbLRerapy7
XCzmWL7utMw8HIusmFyBDzPZk+JKo76rrnSpHcJQX2xmKBBjIeJ5wCLYRDGCcl1QKsq8FUmau6H3
aH2YblIOpNXDLl97PRFFh9TopH4fUnj26x6C+hjlK8aQnpAnm1Zw9ACvaNh/A0tIv8hsyDsKLXfb
Xfru7Lq+PP2xHwhgFjowK4bhnP93EvUdzqSoEQubFHgE33JaqqFjtYG4LqNBbu66aUxlb99p07bc
xFeK8vjTXXTPnL2nW1NQ31VLDE+96e4g9WYiom+y4jT45Ot3Q49saVJCzzRxnFgRFOwUlrP2JN0d
AmL01rSBdtPLPXtzX6oM/Ao+vDgSsSMaT9fWNhVWI2pHIsxce6NdiqxKv+UFRtm/plvK6jDPnb/u
EmeNm9+6xtqCGchClGwJLbT2v2EmZrjgsbBO6Pm5JTRMWSMEDwylthWynDmK+12qN1Sy4P6xvGX+
T0WMzvzB8+elcXl6cYeOGZbYBAc6Y33mN4mWG/cnN5KTT+m6yyBRY/Y4d69OJ4x2huh5VaodUYZk
YHxn2Zn5MnF/YlHucGzRDWqBWNApnlbzPIB7buy5CO3mur078j3sxrfl3rn7XoXUayllBbbdmIYk
ovKHVFpWgVTmYbguRG5W9/3htJVCR1W5aL11LVvVx8ZcOKqJW+kdrhblV8k+sk38fcbnMxnn5MXn
PvDIxxcD38dT2fIlGk1h9gqTG9sdFYdkUMgIDA3KtZ8Xtb7FOYJWkmc9T41/rg3sqJWyPRG4NSQo
q7qcjI/PpfoFldV/urO5sF8tGsLLp7cWUkD7XLAtMztXNcLgZriWkdvq9WKZfnJF0OBfo4wMZcbg
RKFpslUoReCKulhq0tMcYbMom9VY/hrERRpe+aKtIjMeK91GATLuMI58AIvcPZLYlufnElusvqav
ONVJqzo46uWhz6tWHkYRYWh4Eh0a3JuS8byEB6nqPlYEaSkQJ/EGhCfw22KmYWN11m8E5WrBlCf9
HIgrU8fZ3eiUxB/X+dYjUyfkKMp2Yxpgvr5khhIk1iZTMCC12tSU+ty+PNIaAU9hJad7+izwuh7k
YpB+0oRWnwjVo/ztXJ9OYniDRJ/Bgo2yQSkM+M+5GiRYtWGdS2EbzTitqjaegu98EHRnY7kAcb29
bIX81zXxLjYONvgO8FEYPFDD+KKTQ0lxhw6+m2lALWt+otREtUV3wjeLpdi9u0FtHzeRTmXIqjQe
VNlXAhCpnDD/S+SYjFBK0nZ9kjKaDq1Y5+/UGC2X1laHA9GLDedgO2gUz8k3Kv0C94wrj3zbPyZC
ZgGdQ79BAhKoBaWOaruodl9Q7QZY0uhTFeRM/uc3U/k5F2HnCZT7fwul/fWpWt6n4UxcwnAYUb9P
1tUUFAtDYgXBORTSCvuHnb0C4dKLd04L+FxzqeKjt53oKeHP5sNYd0r7ikGBcsdaQr3PsNLcMdYo
eWzqnZNeup3QWY7gVGuzrkPbRKrWVcT9puI8po080EOSHpntKA6z/YWzBpXRKLn4ril7a324LewE
+nx7MokMzEZzrLRPQx4vUclvZ7gtYQF6zgguDJlySXsHcphEt6pc6mU1ZyLhfdn28GsrxPJYHwbN
ie0yr0i3ToDp/Nzg07wbJszgnIVeMD0HfGsV0KVeTWNI/ZgO7OmAAThDrSzq8JpRQO/ByPvt9bwc
W8RJdkzCz3vkkT0YJbbi62D81NAokYoR87ButHBzaFc29Ct/NO+7AtmtdXpkJmx4ZNj00gaYhZEe
9EDuc5NE7dq0jHpJv4K/SxVPfWAb1gWvetzaIos6xrUARYtowTgHrrYw0/Y0AAPXUMoeFpCaC7Kl
GCFeKQDsNWR/MQCYRPmOtDij8SZDLYE4iUfFC/uyFvyw+yoYlfGrIpPshbSvgb+3QSlUGfbECA4K
BYLsY9bnRLoKAypy1/QBRyP3CCGZeEGR/dvcH11q+2sX73AVPNnvHKyczQ/78SXjBYbpqsBi4JSg
Xk4ydwgmmYhZ9T1A0MQ2TmvjFcXDgE3Kk0YLKrV7wcaAuXKhlPCsp2dLcAtSEGHA2CVn4DpMXBXe
AqbH7rrcu0Bpu0yaWmZ0XoiAvk9HUu8yotLw7SPZua9A6/UTgfsHbgj5L1OU8I1hPWa3wEgwC0yb
NSmOYMVzUNLseSEuChFjFrow7q/NT3FOJAHUK0egq135ITRCkgn+z3Ed8CFD+QzUl5jtIDe0+RBs
mZAnUk17NP0/kVkIUPXkhTkFxq3hws8ZagfLFVw7/aOv2lUvkLzOJUodIWWpRKodfWx4pTYC9DAD
9mUfBXXji/2bY7HI9vG2cBTP+jsrhsgpslEEsYC/1sDBwLOIv2sa6S7R7T1ayTVCJRe9XV7PRoA7
TPIVs38b5pXKMRchb88w1inJuj6EmRWA0Gpf7M8R6Ofvr04delroBRBK2BN+AdnUbqUb+dvbOrXJ
3txkUnGjmm5LmsPnFe5853EYp8DBWLFMAVb+ZWvZJqZoGpWRPyOnlWLM3d3XCs0f3uhtiNROg0ho
GzThRvTr7yo4t4fCR3NVU7jge2J0tpK+FAIjvtVM5xjdO0RCh7iDo/DP1JsdzgJbXGbDV6TXiNJJ
LtXhIUm9wyAHor3T5BRAgjM5k+882tMxyLIEKa/dyTDzpe8neJ/I1qEszBHkEcp1mg9TT6dHTdUG
Irj0lEaSSttkhyK1C3x2c/yiDaGzzBkHVTV4AbGPdoXORbO4sL0Tts/hbnxTnkrgC6phSnBzAbih
u1EI9J6v8ZdpEyL+jzSHdOE4LqbD1istRtWo77HQwaj1L+LDm5ZLwRtaO08vauggc6ZFnv3ytgWn
VnvbRHT8CRA+DkSFKMwjj1lf7DktwqLTgMOu5f+fRjKecW6LtIYBRwehwZhgfjjfhLbHfvrT7k/K
FiEUiqrYNa7JFui6PpwAuUOojdXyfEpLLAePYlIJIacR1DayHk85EvXUuANWKex3CXp5CFaiR3q3
ZTrc3j/STkmzXMCntDF/1LAe6cZnf0vCBR0S8RO+K6225edAyQG9Wvhikpgv2zhXpVCR2I0DQOfJ
pFnkv4U5W6XwqPmFud2bgSHPFuf+IYcPJR5r9XAzO9ykHjx0LJd3D/LCkBnRCxdU4IEj//2k+w8z
8ShBVBHtW8ivAQMKSKCMpvHLwl2MuxBILmhj8akUA/0nVqBaAcjlWyPxXMRa7mMK5SKeYfOLMxA2
KqgY9OEDglhbfxTYZifKnRz5lRgvW3tO9Chy2H+4/nfYfQ+AbHeWy5q04EQhboJfiXsVyMHpCehr
B1qWCIo9pq7AVmQU4xc2kELJtVK6bKyjJXvknm/NsGvvAok8b8prSKsp8tn0M9gLIr8dHwNlVa4Q
hbGDNRn/IG3+mZEQMANStIi3f/6ngZvBMPa7X9GOsW4nJiUgp0xJR5Y0ZFQGmI30qgGTfW6ocfNN
Aw454zFe3MJ9QYj6BRs9w0NI847NFJp3c6iiG5VjAzc0g9NAfl9L+fmFrwBAvEES5ZkEW8AVOMPb
A8BjmkEr1VzUDaLVsrZ5G0F1Ho9oh4MmLfDmsyVqQe2XoLcwbdrScMEnsh25jVz+hxe+5MKV4FjC
BPuTJcwAZXoYz1Ygag8WDsorLi9nXhinCx49IDU1V92o9yqKf/un9Jc1nIRDtJ61rp5nSO2fSmr1
BT9WktQo5gtkW2mJr/aZCpsIKyvVWu5C0WOeH92Cum1Z0Vz97YY2msyYM7cW5M4+Dh0bTySmosGi
PnUquEIwFnyuNEmwyI9kJV1Sc6ApiMOlh5fFqu7yiA7MyXc5sZC1OB/5DulDuOGHzL8tJts/WxfX
wE5s/n4wtBSXNYFZsOqX4A9socGQmqMeA+FxCeI5Pf+tINhizwHGoWGvYCFPrtLouvJlN3wYoTBK
4ZmPMObgOWqf9ROiANyrke2qdEol1a32YhrwmwScadKj3IePne9ehPu4twy3ZTi17RZHkt8WIAUs
HHtM/Foet2rzdSJHXWd3qV6hmjp9N2xjwp22Fbid4ObFaKAUWh9PMn/gxRL3xVW9olZO3YFleOUo
nTc4fS5exbj9FCj7StbEut++d3MV0AuMZ6kyfOAm34b1w+/TZlLa8R2DwBs3XPrhka3hVnzt+/Zh
7a6W/9FgzPWK0zDV9w7McraPrhXGBPRZLE8YuxzCaVGpuHS4pQQnaDFFLjJzrl+3s45Sbw2iZdG8
JfStgzuDiCflfnpUQOHBqaf4mJ2rQudfoqmb20aMQmb+If32G+S0t23s6CvE3CJYEkuNm5En39/6
fRkb8nIMjkvsdDvb0J1z0uq1R8dhiLpr76ibbrzDPlZT//9OraDOLB/NyIK/3k+sBc3ME2posfGA
NcmE393ULfxAzyX3JYmt6gNkXoAqi70sREd4rkxsGG0vMyE0YH6/6nTxz3yWEBRS03pF4XCzTq3F
xYRQ31OoR8g0l26qZCN/kMlCw8LbK+/ixTtcgBM+VxTTOcN0Z7dqDF98Y5OVxa5YldfFm3/hAB41
C++AG3a967CmYShIkpUIKbGbHeCzg9hvxhCiRVZyl+0t6X4jXbTspUI7WyxD8etHy4rC7th5lE53
s8TI+72GEZN4wAp/Lbil7p1dS9hZr1cU1Z6U3/gNC2WDA38/Xb7G7x6vNDxydwlxITi61gGw4I+L
xv3oV+3XOt66u7+Zm/F2idYfZG0R4YzWN79QSXKR0OiyEL3hbJnCtI5Lg6PHp+x8RS1GN7tAklOZ
RR+Md4tS8JsycOAOX7GNt5hD+KgTfcjD+yFvPGhHeCYK6ISs6jWrDutlQg4iviP/Y7JKpsjiRjIk
ncvxQ8WSJo6nC3SMypZ4UWeAyrDAgZ7GMuhL0NgBp46pXy9+Bm5Zq6/CSUBXrwXG/Q85JbM4YXDJ
oDLbUyoemVArBpNwpDXGMzAYH/1inIxgxsWV7aoHwVWhqasRM8KSR8brVV1av0PhAjRM2ghSoQnN
VSmiPZlpskA9ShJtZzVNaLY/e4BY4HaHYs+S90jYAlT7htf2WmMYlfRLlmZVI1q5IXPHdGITa697
zU0pUSQF//su5PIXom5XMUI7ebxW5OL9h4y4XRllEnn251EnUu7Mlwr0Z+arMkg9Q/TubqoOHAiR
GXWl17UXh7ZDIHAwvB4BGBFVH43R0o1ITFS2J+tK77fpIhUh/KY1WVCA92vRisrn9wtF1gXubmkI
iXFfslOplBfDLMY85mo3ZVHtaOIVzFeIWqMF1lExNP7By/6adJMvkfhTZNuXUpz9uLZunIsllTkd
kelPXoBednk4cfFNeP/GzV/4y8BJh2r+W+hWtqCPNXqxRlJQpm68ucGv7rAkbgJl0sSSUGhPWkD6
E3PzgWkljuelVv2cEEFrEHtAZ/Vv5U4oFfBQ93nwXh0i4zeWuzk5XjoOpvAI4HnnkFOv6DrFpPA8
HRJJ5xb6JxYEpVKf36Tax/tdiuWkzt2NSga5QmhBox2AygNkWbcNcZQGdjmY+g9Ejh1SSsz+QhHM
/ZAybhK2OLVWBPDp5Cc9ONLs+HmiJLfAq4DRZ/AG/RHvcfsKBZaMcels/IR4XPF5atn6vUCnBE7r
nDKKCxYJls6wt408jcKoZMJtOi2B1/tel5AQlBXLNx0q+gZTYf7Xoo7AE9EN9AmR6hS9ifSOB3z8
6yJHAmiC0e+9tOwZqw3hanpVWyzaH1OIJKsx88k2utzZGVUckm3GCPLUXlzlAAxRpl+cogOR4A75
m4+Svs1sZlUSxYJGPjXxVeG8dMLTLJt2QfmKwDC2fe17lfOd7Qf3EP+nVIBjkXxVJcNqn/YqV4dQ
d1wt/5xERoNi/iLrUIxN8ZLtdoJ9HbapJw2bOeiFhBCQpcl2afwSGr50EmwqEj1v/Lzoqqj8+BsT
Slmb2q5OTWBlQ1cxukyzD2M8AwNwNQtzORQglouUoUuCBOMVZgz6Ley7O/z6wT2GXd0o/Q3g3M9L
eocJ9jgwt66vn6u45/Cxpah14UGELA2m3IxRSPIwdgFfhqR7skx9NBc4kP4kxYSQvJHuxmw11inC
RIvkYibJoE3gwJkITp/++7FJp84Xuoh5B1L+zkt6s7sgKXoe5U3Au/2ba2JiWA6V/squSFRuHCoQ
vuRL3ewz8rD3ZapLC5nhP+63RE4lAYyR4Mi057yJ7LMVwt1zDU+LSwQvznKkUOUjBm/bEHVFcG0F
eN/mBjifIdKZqeJd7V3UOFozVJZJRtYZPkXiXbUjQ65YIbJebP5ljtze1UVScvk+f4fJWnOa5phR
7JCUVR/rkWNrg1dLCJ+/NlQXNJkbazb2AJZJtrjbG+FKzj4GtcXzEmCtsfz0zeuGmxE05QIH1nFA
G9YmE/Xru7WjGUFwIx190lVAQmuex1XOBP5aIhmCQS6b/0kit09Pyv9TsprJshWSi76DO8NIMRrP
6xu+GyzaLZtf34DniaNXEbfTCbG8ZmCpuXPOrxUndmrgVRYxBWYEG/lBzfUFaLADumo7VLDGXV2w
gG71iqXj0HS26jfudvYDo2MW9X9vwMmxOhbNq3gFFfVslZCpts1xZD7WL8xGRZnv9TpJGtCFXGfe
xo5eIEZnHcianQdatJF7xh8cr/CO5rScklfTD0/ogDAppRJKtjs2obYqnN33MNUZr1kVE2Yd2scY
r3hmmbmLtjDEMXHs2ysCPZ1qo0lUZDXuYj5PrU+0uhNB7c7urceU2bO4Ry2F91vdlMcHV9CKEeKE
C5fjevxBk852pavtmz+b5wX+4WE8qEvexdjXYNAyPY/6r7NIZtcX+UAC3N+uZWj0ft+GoPHy7SR2
zvBhbDbVX9evquNPHGfYmtJ5kN2x2PPzM4IMQQwudNE5Mj1Dg7EmGZgc64YDPXq2q7ym6xAo7vZN
KLg79Ldq3lamRlYCAq5+cxRvE4ik31BfhMoZbC795Cnf+ID4EDFdhtoVN7dC3lPEVWZGtZrjdN5I
AdEe3a+KXYulIkhi45Xj+7KgvFb35sfOmXimSuVfnZ4uAJsl/huZSZydpaIbsriZulOB9YUrAJtk
xdaUgn7rt4lQ8u8wntIWbk9QKZ4xshDDNOJuarOEIirvP+mFW/6i9LO2cghc+0rXz0hSgATYQ2Xe
fDbXCNEfdd5VGUyITl0PA/b2FHlvIHikDwjmK6Sn9y14KOtGmEiX8448+IHwfUSXwFH7qcpiAvNY
05OM10sS+bC2wAMvWCwWTJdVZ0t+LqLOzl7q/N8LrGNummnCtgUk9yJJHmR0OTJhy9wMcNgVMIoT
5UMesMq8mRWkCOdL/eE+MOvtba6OxmuPLFI4RCU1EwPj0pza2IQtg08hjBnBAubeliiltTFMhBbk
WVjTVj5+zI6xa4pj7WcISZ8dCGC20iJlJbkmMSNp5eXOOPJUOqwvsOFRPNmgGN3K1E4FZpjw8Ocv
zdSpUT4IFeb1NBGLG/0RtrM1MWhOilUC6jYbZyhcr1Jxsa1rGvbFX8Dmywv7weRLU9jBewSd2aWn
TOmNC0066xE5Vlr7vapo51DIEk33OfmBc4Bn0/3Y4TcqwBxq+16nnLcMW+4Tq3QnpwdBbSIgMAgc
Apn4SLkQ2z73GvNKei5RFNMnzWZa85sz9VTBtzSNAO/WO03nsj2rn+nhrDEkTCmhAzJZYisCjFYM
aQtmMgcIz6heE87xs9x5mAphW7Qjgvp5OlUvsuGyWh7aiByyzk/f36ko65W7+1W9REffXyshxuC0
CLhGJ17fkKx8kTouPWGex/pQkJvFhFUmTWhgVyyM8pFtOuOlMUm4ghGpySzv4l8uCPJpGXgmDDtv
JJjUvibDSSO7jyCXyGNy+KIrHFpXzVmZIS0K5xc9XGOSGpLzURmvwonmZciiJgJ/9c7h2pfknHPx
kxGI2dFhQhe3IiID42ctaGeNwby9oOd0cQmkEfVcMMpZqMFPHDm5RJ1ZbDz+ErD5vDP1X6jzj1dq
jhAbQlUb5qeC7BjXMM92Nj+vf2d5be+Bn057yEQIvvbhB8dv53e+ssBikzaaraGOkUeS9zO83r/T
MpuonFTkgegoXWjpauoW/FMDVh9GV77iPou+v0vq5FEpGI73TgBrH9O5ZLBCPZ3GTM4z1H/8XbkQ
M+BTatm4VJtFKNgj2glHFfwUiCNe+rH+9lIrhAg6b/1MC6gR054BuLIf6JqCAccttZCJA32hjQkn
zdVhFF6fN3MCX4Cx5aY7SZeWjG424b9EBrN77i9U1j1Ws6x237kcif9tlgGyhay/OjUonfa8JSsz
RbDwh0+SOOQuA7v0AOruW89VTgmHR3l2qukSs7OlTEbi1AyHhAHh6/PeFCkFnHz+Lgji2ZYA62Pp
kjsxD5pgFcOD10EgaZ2gvmwOlkTe6rlRlSL6TH6uuHRmkQ8iYlyWoC4xz9ZvCYO3iNsbYP4L3W/H
fqp6V3jLbcNEPilhouROiBLb+yWhsSDvckTdMlxB8uRgzZLz9ALF4hWC5DN1XEdquPmuQo1Vj70r
b2o+eOsg0apWe7CQXBfEovVLekfYM4j+3O+OA3FCx5eBcM+VXMgmvCbxWbMF17r6HVA3pTBzYmRQ
CQHx9o2cKUQxlnvncXuATFw9w8TUYjW/ENhlWupGaqWlDJ1hBOBWE9Px4aQ4R2Jug4NHQW9ExrHA
Ujng/7Xr17ICpuhoMFeyNSjWsOBwGnAHpUk8ATk44TP0gbWGXliCXRb03l2kby3bcSZnhzyByXXE
nVSWfc+eFYgZaOOA1j5h5lyCCdd6IFBUZCbRtICaDtd2leykXPIqZ0BNHeVZuFZb4mdsAc+9YUSp
GkFAF7wzSaVN3IIdko4noDF1djXhYV/86Esmqntf9XoFIEE/1Fr76ygYoyQbkM8ub3OlzAbuGgXt
xMDXodzlgqxkuPeV53/1bOVkFw4DvmBRK7/62o+F3zXf4sRXRz+wcHvkVgR0wtYDMrgKz5qeow5Z
pIYnuIdSXMbYl83uI+Q39Iul0Njx1+oPAftxI9FMJNR1eUnCwWG/WcJnCGQFSEh0rq+CYgzdcsID
C2oCUf/j2IRuOnEUkRSxEY0FLWJOZXoNgGc+sEY1Odai/tzXoV1z+khf7Aqz2hCJGYvZN7D2axY5
8vffcjrUL9v9cHwuA9TTflU9RyF8mpY4XnA6DoRxz0AA6V4yoh7gMAa9p2ybu+9rjbLjZmILbHQV
hTJCR/cI5DJu6idwdJWEJ9F+sUo4GJ0G3zWZ1V6j52j00j7CCMDzGnRzyeXRHimdYJpLbWmPFwdd
LgyLP4/AFZj68uhOW0vaoePI7xXbpk0O2CPID9elhkTNzWAZSKY+lntM5d+cl7en3xxv37UxmXqZ
4iy4pKKbTx6jdD1pyQpmuWzTmTixjnWwuKJhs1wz8ucQNHx1zdhB6XRbRr6O8tLQxuS3vNkDicZU
MuuZHEMbrQrMO4LFAwCOzSD1OzWrBbBgJ7kZ5F9D8M3DjQJL96F/Il71vBSsig+799h1jfCp6JuN
9fKnGrAnLlVhwToSQpusAQOW4hWAWqiMFnCEqKjvDLXP3dVd68HtzyCx4xEcJNs7f6D1X4RtLDBW
EB09WXQt6L2+RgwXOam4FmJoYgm2Qh3mE+uzFLEwKxHj7AcdKiwOspWo70oeGRHRCKq15Q/9KLkO
6MWTpeCFV4AmFHuswf1lbaOatt3nWJ/f/0sI6kV1P7QsiyaHNaCBzHHD79+MkG5YUQ9XWimnKpZM
tEOzQqNzYZTkBdSsCM9p6GUmDpnKSq86oymSx2gxNpUEnHHtEkKt8M4lg1KtNJ1NQ4dU0ZY+BwVf
nkBaqNhneSnlu+ObWhcQLfLZW4zRlyfG9u8hHU4hzVrRys3GzY455VhdSp9/NkIHVO797ZgDWC2K
0D+0jNsLGG3FDPftoQ2I39Jy7MePora76PleWBM0IvAGQTZX7B7bLUQqq/tuEGCGG6zXAP+z3DJb
xzIDcOeQNavVlRIX4vdO7M4tRkXxeIzCE/4ruMChzejYFa1Y2s/LDN6CN2r3YVp11t6XUtMfsv3i
mLnFsHJCWD32A+q0Sg1QhwtBdfA4E2w+9ENhku28lHDBEhGKxP93QSP/LFpYTIKPT0UuIpSipJKJ
MNfgnwaD4TTTrWjfWKUFCkG1GECngh++Mb2Q82qwnl714uaN9IFRfA1KlK3qAB5Nq1ZqoqIE7uWX
U2p4SfdA2C2maN/AA5rQOjU5/JKn0TtPuxr5SPCATXPMAhKV3XiPWH0vKQn/Q7ZySwEz3hv5Pwyo
ArDMPtsoj0FLFYlg7yvJQHsah7udRmTQaMoYExVy46/Yrp5D7l558k6BVwNl9qqliJrSuTAE+M7j
hm8S6ZuU41RgeeEeY4KfDhxMGfrkSoNpMj3lfr3DRUxDzx+JyraDt/v/qiOv2nyiG6XoUI+JQQCG
6OQLnX+8h4A9THROe9QsNKyEkO34JWGkcJ4gCzbsHF66LKqHtULK1Lpka6CP5rH9/tCkluiNZMm0
3bU4qKdOl5x6CeQc0lfKOeqJGhne2Pp6sg2Hu40rY5L9VmVE1k7pUcNdUFfBaAc5wuS2U4ESvAj3
oc/7fxHDetfze7qbd5zqvI376d72Emb92pWfZMBV9UfFuO+5mnb1f6YacsmgamLY3tzP/TCOD1ld
a3pcFFuVHbi0JFv6RielvitAx4u3KGqtRSq2/i0KaOX9T1dYch7Ze6wfcKfVG0LmInwgLvLduuxW
hBdYJYbaWkMwIurlKFkOkYNUCszSujDvIyBVfoS9KuVKOZr94y2vunmYWMzWTnFj6cKy/UxOoW0f
umj0tMuoJ6ie/ccQaJX5npQ3ESIdrKmmmZOfES/pFFhfd/X9X+g6AXrQj3N8pIHMlGfNo+6y/7xA
68e1bHgrqKgTID5r+xDjlVYynV6/avoOX1b9MRDr2g3Gy/jwC/qvzqrr+px7M3HkuX3XtT9f9699
0S+uCXNA10JPgpnIt7Ukzc/PjSxOPOQz2EMV96JzCUf2p60QxpyzfbNB851V2JLZZr3nfWorMtXr
uItIVSmN3qdaRvTW5gJB1gYfm98JnrjisLxWSjTDJNhUJADj7TNgfaohT2TrS77Y/D2EaBoLwQ00
uiU/ytdSWAKgNj+Hcq/3qgtNpdYiP2Zn8mdHm4qKqnrKzBdj6n5m2P8494FFtAkISCekKrbUhL6H
SkwCMBbQPpHRGCuz880S4QhoiHAAdQ5BNQf8mgRl9tzIg2v1E/vsTNcI+yy7wZgnAg2linmEYxMH
i9L4YdhECp6AHGLgyQVuc/LlkKAHCgYef5M1A1bTHTyhks3/z/8x4OTDye14MNG4PuyNLyaCUiVv
4VRauM90CCzuiO2AT2hjCdMExWAvz5pGaCKPT3V4ueTEkqGjqCtuadlTbn7mos9blef0FQL51SGK
md7MuV1w5e1bcKHGh2IWCO/phsTLhcR11v0ZjKlfbgvjIv6ukzOzizqMELmQ5RehOrlduy5OLO+3
/j2piLdYPSVDuYYZxpZyXTtJfqQsJEuSRvbRpAuMPbQtuMCD6WyUhP2/LX4oKw97VJA7F9fJqnnu
ZQCEh/xwp3Iv1+ugiUbWeuuFcHlG13s19L+Zj+LHzx1TfX3uVpTsx4eCZGDqLpCGFkToN+jljohr
h1bCy4/JU75uV628u1ELTfVOSRJIyCpWGlRuSmxnP6K+c36Eq1SH/WGQpnPq8c9FlgJN2jIR3OD1
rrUldVVA+VwIn/IdO71K3eK9K+FXK13cU2H6X5ZIQtAnffm6DpGohMfpIJ6UtFHzhGkO/e1CHWoK
+FBC8FYOOUOTiwDjkRDuWLT/P03P3S83DK8AWUGQ/R/A5iwq5mCUDn7RpalCZpvvq9PBP62NxJT0
zHOagVgnNeNvX2eT7S1ebFR8JW1WGtI7+v337z1qfKu/5QJ/Tmda63R9c071UqyP9WfJGiSMWns2
cjJQepL8fivYbR4Sp593l23JmzNOWuu9VmJ1DZ+/3zMBYS3RZCktSdQTh2OMmJsg6Xmiu6B985t5
ZVh8bZDIhlSwgjlHQZLvRHM/gxHt6dYbf4Lwm5h8CwaRMa4ZiouU30aPyH6sGyuKrVhFIHYrz8g5
o/d7Nt6k9IVpN5fyvlDWn4nVNVNcK+PAFqyOmoxA332DJumDyhrwO8V14hJDvNUONV9CPkWYZPW1
RNW6TMOYxJQ+A9gEtWa0uvtFCeCgD3dFb+PDb9Rqmcrgw1nL6/7CttesQ2864/36QGk1JxXK/Aon
ezh36At+24E/MJ/Pdn7oXTvryCyur2PydeIxJZFXJscPnu35fv4/syBc2NKYSCnsK/uzqkH8/Coy
0zsQCgSPiniC3qKkugtT1AP5nUDZtA+oxerow0srvQqMWZdBeF1+k2sTRqIjr3bezCpqcSaXZhAn
to9pzaT3XJAGLUTMurUGaCOFhCAcjdIK1Ysi57dtnLBwrmG/enXbF1/h8DkdxqDSTHuZ13uS4nY4
4gZbxPVyLF26RNKbffDBAjyEfgXNp634SAAutxuTHprUB3dI8S+UvU8hrtWYOV8y6LEZTpzQwx5G
dr/O6bAXiCwh9HeA+SSAsrdRjJ5b5bykJbTUvcaDbP+1JcPVSFgDKkKsshkVoUdSOXW0yeWcMbjv
EZ1fadZpW/eQkJHBmTlm8inVhW6fM9jStFaweuSUQZXiwzGdYCfxnt5Y2QPn2Xcj3r27+umxUdd7
8S65QUZOzEazraeisDbL3mVkM+uugpK8EF6CuBnHQLNMBzQJPrz+YI+XStyq3QhmuJZSbwjT9g1W
s4oDiqBOjG/XpwivbY0Ppz6bYrKAmooB+SWbZDcL0er6aTy25iuqpYASUrBlrnjJX6cAfg5MsIcb
bUNkEflEX5l7i48ckQ461GkOxk3S2lD3Rdh6RFxeM8T+95cyTOfIDapsoAx3lkpjN0LrZoEgA40a
OKEK74eMqMLRjgWY4v/QU3V9ZlQGkozxV51k6bn9ISEKzw+o9m9cOqIFU0Ox8IW/yUDa/mHTPu0y
saaFM0fKwXt5svEYftvtVTCHcsHWRRhLrgHx6sydwDKyqTlEsBlP7SdBinWT9mPW1apK4oynSy/y
MwWevBYkvaCnysr109o7RJGqKLsVYEACKNoQeQWhiaWrYFkNcGR1MRkNXIGGbwu41oonsKkbzwhV
1rBYYnthliWdjvCs98nHCEstl3gn76woQrZoyf0lgGTPHHCc3Sgx1HxCXoo9f8oYUXvgAlDco1lj
+9isvCz+sMcChO0Q+fiUOiilDSEFyAtHIjOfV2UfwPi0zSmdtRgDom4ZmCImldU/An1igYqOr2PK
md5Jv5UVBrRC9dJEiCZ/NY5bEzJk3wlnekEpTLwlh+rgjP7qbxNp3GqFDe1vuLWJO967Co/SvkMK
w7qKX3ObHGb4X2oiYz1s9Gsn8pusOS522GFkHKiWkfPlbLn57BePcwpQlnrsbh0w6Fl1q2ePrOA9
5nN4M1ESGdvjd3yLAuAEhabedfxeRU6Tc96qfjhfxyEVuFb70c1mJgLbBccjaKCgnqdmkpSb+n+t
+grR3wIihYMu1Vv/+3EPNKFTUSAD1ok2iMa6UzB0CV7WR17y/zI/JGpVLB6WYuNbARqLdCZSRUma
X4GhxSSI0NHTyJZ9diyfL9LiNI8ScrRd1LqGx0mPiNmLoGbqC7u1rFL3o0Szkiax5k6KIX6lrft/
EtHzJApieSx7FX36tAgfYQSyKld6ys3ArrK9c3OiKQPfpjCMazel7LcgHTT/+LW/MZFYDBb6c2zc
z2ERWgSdWjGhWCbFpYLeoyAxCwXbR4ArvS4mQRNq+yrTqviYJz4Q/Tg4EkIbY33Iw6WD3gpTnRwt
ad+E2l6G+kYAzAuwjii2GIDLXkzRePqlrYPMHr3Vb9cKGDVI6YlLbuiSkJNXzjexQS6S/j3Abtux
NXVMakG9MYdVPGE9g6AkksQR3A5BGlnV2/Tq9GIVUKUEnrRbHdu0qwRmT+8e6Ere8yJGgc3dQMup
wBKc5CPRbUwv50vsYB1YZwlE8YXChXoE3dzulcbvW7YC7S/JnX4trHRfNaHLrO0Mk/r14r9yiE3r
1Gw+wZW3LTzyyYge3DZ8/YGgOE9V2i/3waDVXfGwQTVXq3dAagJyGUhLn6g15syBaWKfDAuAPvNS
u5Arp2jXE9VtvE6/dVnQq5vO2MU5L8F/7vCefdueoEbA/f/OUl/g//Ho2njjaSTP/zrvwkRXoEFA
cXRAQ6pJIWfzHOKsxhXstrGNxOTOgdbf8Z+MP2EwFY3+bRpa1jQW+ksoXC7bpaVNPKbf55krTvc7
hN+dPBszpiMRsxtwOJeb0R/zA+SZRqLld7UFL9q5mRh1R5Bd0WP735ecSsOVnZgSZ3ip261Q3WuC
Xh3CTR1w4xM5L3LuibluitCKYzDW6aLZE1LQVpFtL76vt3Nk1AGWQl76j05cbJnYVo9k/YbQTLti
qjEpzFWYDS3gQFtHvovIsTPGEPOnuBs+do0Fm7nhjZAFb2pVweppYId/lCKjfYTAVhwZ0CaZGNpz
/eeSDFLyBio4IiRaPxNWpEAJ+itKccyKS4/TPlCEENKzA92tCIre0w///CR7i78LgxDdtmGaJ0FU
JrMcGDxgfShbzxf0WPmpvdVSO8r9PNUTB/XhFavcbX47IEAqzW9pc4hRf7Bj2Sq7NRn0m16mWQxy
Kdt7372v+p40KQIchRBFqDSi18ehT5DWoxS0UQ7zMOO9MeKBmc8veG7u5yzTJuv8sZ052N4lFZAR
eCkVaArlS0rnpst++lqaJaPIvpk3gszrHKZg5pwZ7y/LqtOJV8+3eRv+dLjsZJQheUo3rJhxLSEF
TFH6zqXZXB/6t9py7eQ5OkEcNVv0b58Kp2jOtiL+kyjQgCyqJ5qDBv0XFkvYx8hBIw7JToJNXTeR
2SSsB0LMq7dY1mfoG0VXDOYSDUqPABTS6wAFAT9m/mM5tU0pQ49o6dj/sGZdzEdiFrGX2U20OuuI
M7+99MTDgldpxaC3xoSu2G064IKWh+2M2MZR6k6XBfohk2bCwz2tBU8dA5BTwUTb8OZ0RG9YmXgi
8S7wvZCH2SXV1hUDFMnLP1RJvOpGpvhT0MJriRE3jqwo2Ll01mb8DqqrmwWsodIgtt5sBzImx4CT
vG1o5MCHJgdMK/KU+oSb/i8K8ltOtZhJHLpVzl9QOim0QMDNlmaovDZYsUNfwD9J+f6H9QsHk05J
onJ2SuMrG9fBZXUk5IiXmCOr7/XjTZHZR1W+IA9/+SbxmZIRmQlMWnizxTDNOP1+uPQy/bXUPeQE
nzhc3N5zualJKsEsdmsxJrhwIBp0EgK+D+IVuRbiMTtZIjc5m2p2poPFoydCP8uFivae6pBFyKSK
vIHHUxtVuRa9ZD0dI07UBWtDPzpfqAXR89kiWBl2j+RA5gDF6vO4Oxf8K6LHKX8EEaVYtwHkhkuo
a8ah7GgD5gsI1jEP+hDl4AwdOeLeORDStk7fts40ASKoN7bUGWjiP5NPYvFX7c89Hf3WL5EALjxj
Od4S+geHUJtK6QT2J9ip/FsNqhCUrXhbf1I8NxmlufMByCcMWrWazKq3NyGEBAV9ND+EeteeGopZ
Rbu3YsYEM+dKe+GNSx3mZr64N46SWut7kAEMFDIoUEwc62pZb6n4ptVwp/r8H4DVvXGK/ObfP/RF
MEXOvroPMseoTotPFVGGFP0jGQJSw0BHNlrmsdCwBTZW9+qB1YG+Fz7dEcVxwBROEaHsWm2NKr/5
HaosDCL4fs8/+80xE2GMGREpEh5eSOyDf5tb4krgI+nMI/Pj5fj0XaBnoq2N64U+oJ1vy1dRctas
AitD/EdDl9ekuu8LRxtAbLN4HxLsQCXW2yQlNYN7M0jI1yArUGWIMOAv3MeBWnYZAmLXHoQ5p1bC
gDaEfJhAim0JkfUnp4EcmSXzy8JzwtEpx8oJe5OonYEDtz+JYyNUbEw68VQ9WK/2/SXWRlJRAvnY
RiXuX3CD629nVSbb7HTrU5AUVVR7v8hhCDvALKt1UrQJ94MBrC3AZKfoMu/pDHR1TIA5HG/TThbD
5w2K/AdPafFI5d882GkdN0yLg0D6IeNoEJmjbM3ZByemCfG/3Ybls53fkNwwdwuJd/kxFLjk+d9B
JB9CjsJQ3lH8x/Z0gOp7ASz/dXbl7/EzBpE/YbZKrB87oYrtlvGSwgvAPV8NqkHa4NvR6sdnDgkZ
T+JetgGRCQVebBqpX8KH3wnQLjgdtoR0WIsFyddps9iFjSvOLBrlobs8vXAFXIMFfjhITKeIAftq
N/d4OEzm5S3YcLMaj0DyvlfgDJvxvZ5w2d3q+uwYpVbqhZz126MRyZppRvNl1KGCM8TRKe2hs5Nn
Dq2U5G/xTxs+K3w3CnLnO67bidc+n6I5QTRQa16ULYmsTkvWk3+HjLDTj2HMzoYG9RYmp4CnTydH
dCOg7/qTdiusNXXKiykf0NynMVdhbD5XQiO+3wXXn0Y3uP9JyyZs4S2f3LyUBNVFFkn3el8jg+k9
snTsopH90xa/4eZW0uqGIinqR3SRSohJablOjhn77E95GnNNVNUcAXOtZ0lhXvwFsICdd6XcM1Ta
R8jjfmpU/B/qvdJAbNw1nZg8RCESLtbQdHvBSghD5x8EPMXATV1+8CBjfAFvUSLMCj0v4FIPer5J
sKMuHtLTM8cjZ+kVrKqcEnnZmf+T7e8uwrgkuq0WOmrO1w3UTt2fhSlekRbVB4VcaS4F+Gv8BSHe
NqJNbh3ia3rvS95FFpA/KGwgj7VgOsST00ZCm3+slVNE6kuMpsNtUEtInNgFBVQs4I8Xj1hMwgZq
njj/NqCR8RSg9oIVi8ax3WlrYmqYPNeone2SjR24f51EqZ/51nAvFuuWCBMhBJzOng1VSi6C0j3k
trHTLbMZuKkm+uQhKcyzhDJ1w2AyATOrC3+7vRhb+G9PcLZO6pDZMTLsBNr6m2b5HpCwiocOEtfY
kowIdPOA4APZ1yBn/6RwchV9YMM5rHtQarMBn37a0ePTkV5Uy8JMuGBv+akh1FbGiY8jMKw4fIt+
kdUn/GIwNag2BcKWpvzdn6NG9fAonXbTrhz68UnsQHa28pd1MCulw/HTzr46D0K4b2dfqzsvJ6d3
DbvHjOfg7MQwFpccjChflxJpvxIYYIBbaMDS1XNWbz4ceNlxhYUrLTb0ieUFjTTFbfLTAMKtvHIO
JQR+PXTrVs+9uZv5qUzIg5aLrXDrOhj99a1FVURwwL0bzdPgdp9i/pJ0IPY4Cx1zk5Cpabgy4ODO
yg6rpl3WuCXLzitz0WR6Nem3BdQoLxf/6iY/eCY6+1CXhuFR4Yz71gigJRgOfoezj6HmL2CrX6Sh
LujvpihYdMOXa6SmjUOZxS+sxa6Hn58b54ESeNQI+ILgGutyajWkZcuKDtUQ/NrDfnEPcPRadvY0
HcaYW4ojZR+KNFTX7iEReinDlFPrCRNljPWfqlX1YmrDezmQNMinIxwpV+41ShE4dyKRO0fQXWgK
nKMPr7jOiAfamqlzzZr5pflA/WE97u8+8nYWtjqtS9Ad4oVbdXUUvCwWeq0JuIOaMZNdcTC8LqNx
S3VcKlmdDoLKA3WNpfe+lFEjWai+mbVIfPLcLOulXDn5BtJYU7y3aVw4LSLj4PLD5pTaUe/Ltokf
Z65YE9visabVVExn9Ag9TLqNgIW0vck+9MZW2r5xK8b/CPIssrUlI9xjCR3tAChnWuHirTV1fzh1
iWsgF4340MbrnWaDUkiNuX00VmNbvHdPSLsMjkUTYdoxUqgYy+yuJ6msvWboqXQwlvNkYIYs55US
CiOlyQx+yINJ33r1Lr//2UXOT7ZMk8ANNBK+3cB3DfaHnef2Oc29K3wrDnDrSxsYFcpKK5nl0T+l
kHUYymJD3wQSFUtzz+T3cs9tsb1OtmgycGpm2fj043u4tMTkPOc5Oq1cd73PSZxW9zMsKlyYhyDe
OuXKqWVLxS+i9ZKXDcX87URUh1k+xbiJCjtmTU75qflF3W66gVeCxAxva6Aw2ImnrfWRJDm213QV
64BAbYMA+yUYsBLVI2VPlGfVox1nC4IIS08zIE/+Og2BKY92T+m0raMpPi022AGwhihwZU49ZfYg
R0NMXCIjKfKnKOKX2P6iTUqQSOOdU2/OhL3Xs5TGQdT5b1Ib3JQsDdKHY3NnWlLRU6u9CcRpDl7r
PrPMq4nNnLt0Phh7/whlwma+nmUr6CLe8RWYU7BTWOH49G+7XpwpGiFv3jnoX642bv2AKIebTsGW
jx9QSZfPJ9Woq7mNetzRpgdFu+C7GWVoxjee+HGPjTY3AWqXmXyxY86Vx62QN4cnGpLuOLJwkYvb
UOMOrtCWT9pzEys8nJ0r+cT20GmWLTdFV0EVd0owdihjkBl7s125AWsjEiCQP5AN7BKexpvphIK4
hKTN9fmZckeoN6EslkOH+ZbnhaLZLP933kYzNtbgfK4mOclL3xMPJbLHO/toUsX/fe1Az4xRm+hx
CU2tkMYNzqTbqqf4xu736EgtO68euKzbRsQH/5kYrPj2xmQDLM8lLNSIKlSV7Rs2IcBC1KwrWE9n
csory0XL5ff59/tK/QIYl4D72W8uPBSJNPVD7aaX1e1iSy14+Fhsj3rEUF6affcAoXqqty6KGprs
obpZi1e8s6TJ88nZUug6JyeHsvIynxGWivzspFt2s938xH7O88ZBiJu3P5fRxdwLUOeDt44z2pWC
2gvFrC6Hi/G0JvjX6T9NWZjoTcp0QnDjScosvw/9ERGzfMHWBevb21sbXhMG6u40E6g7nQoEzBBA
5uFNMm3qqX4ZK2vjwVhMhtRLp2y/5dA+/DULMRpFdusC5Za06R2OuHPWKwhGXwHGjYDVeWtKFcYu
FApKVhxFcDRd9iu3yCVgECk81CpZ6Gs18XSIQ+hbd20GsqoS284HXvOwsAur7lLQi/wxuYe1VGpN
O84/stZyoXfSXalO7cf0FB7NxYPu+klDFOY7p5naHdZ4XBej5tDrODOMUWKJDVP9FVWaAhslUgaE
158XZPpXpKaM2j0gKSzjV9WfnjC3Gb/dBKPv+zButRoiDX/LaKd6iWSl47JMYPNSuh1fsQPstgN6
k+gYBQNC7YyQM8YJ1mf3KQw3h9xDBKXvaa7SU78pClNAsVzOd7v+mTDPnjHYv4cTrWmILOmQsm/B
O1lKY8oLcJg4bMtmfEkwMr+6MzYB+P+D6jwv11/+SYyJykEJPKDFc9PDhVXr2RiuAawp0PFSRRRc
OZpDRtgpqkiBirkHmJDxpqvlqIFHohIUGkvbJ+IwMUZmMwCaNdghy55+aV27T59QUYBVQeyTyGp7
2tLkfiej6dmfVM/GAkF5bGHXyNZ9/li7JZnvtNvhNSUG0O4klKfyFGSDkCGEoI/EHE/cT0P3vTO/
RMGws5CXY69C7+1bmFruMBhBHhvPb+dDTSl2fo3rRiOoMWIuFBwiaMS63xeYBrL8J4FwuO1b+B6y
wHNCnnKWn8UWPbHwXF761Uo3XYT6HzRtIa+Wm/tFoIX21FbFIJw416LGs+5+m//AN9GeijNnN0hz
4HM4QVLTJu/Rk4tP/gOhxIyym+UVG/intS4bz/VA4ey0IO+97iiAq7NnFx8dfAQ80pVAm8d3Z7YL
7RZxk1k1E5MmCF2M+kRj1Yk2/j4rnjyDNt8aVd9ppvjEowW/MBWM+uQajnsDrkUui461iQZHT/R/
v+sShQKzZ6k0YcHzYMZTUo9Wm5FKY/nvELyVGE+g2jJTmiRhrX3Z9PJTl6ErZNuBEUBaeNbmnO3n
RuJyB8eqBgUl7LUT84geisvyhWzTgJQkDroMEvUFdZfhaok8p1Bt99S1J2nn4MYFrkU+bwZXeG44
bzkskuNl0KS/vN9moTCV891+1rfZs+69EqpGDtl7t5SHvMenPEwXurSaqmyMavSoDPhtAR4wJ17L
DB9WTafgwmk37RHcCp0AO/k9AYHDPoNcoz/cpAbnLw1QyWHPU5IhJW0+zLqp307EissKFIyJvk6o
nvsfyZY34x9HS53xYgTsUKWuwy4VEdTAVsmnpahNw9gKaK6MZoM+455NeN84C97ZPrxhh3GyVVTG
b9R/Urj680p9wK+eZzJAgclostJBuRo43suTAoIfF2uyqcw6djb65zwplgVfBJzjj9XVQK+SQzRV
WP8ZI9nrfwB8xC0jYffTO+4aF/0vfpVSThG/huJL6Q2g4FklsgEv4kg6nz1MYG1updiI6yadDHHf
xp14x2UHkglQoR9MojwWL7ahrl6CFnkyAjhSWJGQ4IOb9IYgeEs5wQb0Gg7TJzcqVoX1JngLkoBQ
Z1EfXUtwszpbAcDkDUWA9vY8tKC6VCv4V9Bzj2eaiV8Iri3t5xmnHLebXyFWd5eq6xAzHhviM4mn
u0ioCHTFhTnjt61i3tx5fpFCxIGaGwB93WMLQ3syiIETZaQXIFQ9M2Y2r2ybTHkj+OuoPH+RFm6r
kDO9IPe3kH1oI1sZUxuJcMjD8thCdZR/R3l1AHzUjIpRBCmVBCGrhTYjH426Ryr2kSPioebfRDIc
Sen98DKy+U+upLnDhbVZrWGpFSqLXKqqEKON+F1hl+BIDIEmWI6sieDhEz1zfP0nKi2mOuvXlF7E
ufNR/QKU2fB0TYdrOCjRTnJ6yWwXbv4YMkv/MtwsJAf9TljZ+3fxz9YMsaTJ7/Fe2r0FPhvbN61h
RBzYIbbfYL7g6sZEloSIA7qaIN6b/SvZbQ3ZHVZ83HGMJHqSlr4miLjNV6U4BF9fGvnYdMShw/1Q
I8uWi5Bf6Y9DakDZxeaQrlCDPdW/IMVgi5F3UreRfaHMAIXoKAiYSwNk3AmEak6jneWihrOA1nAs
xP2m0cja7mBQCHJghHZzOe/CSY+rokjwZ+nx3ZhCjpp7PUVEPDxKVOGXT7/q/LOzbQkg+r19swjQ
848QFhMe6qOLdkjY3yiira2jrKA/Zwe81Y4SLaC3pbxfugM8Cpy4C/iuHlAwADRSnn7hZ2Gh6X9I
94OSdW8eFjTga7rlO7RIO1ED1lYVFcdYFn9ei7HFUdattyCJca7/sa5ZZpFmSjW02OFdc7fp8rfD
XPjWLgM7E3OsOfGMSL1rv7y3msmb52L2b4zcDgR0Twe3Inf+iCLpkqTSXYIpYgwEiV7ypA+Qbdnc
fhPrYXPLf3+WJdYrJGVjPiPN/wtcrN2M2IVyqB82xGshRj/UGgKt2XENFK+XolSMVwxLuzBpE3z6
lFunUz1Hy0SvIlXj6O3iUWp1BY3IZ8F4i+LtZPbXXTnvHX13+QQG+AUJKvQ4qyyWy89VuHMPqmV7
TWhkI/Bx1WVW77eoO2faTgDJw/VB21YS5Wn+abOvfO1c2iou09Uj7Mtyy9kulFN81AAekRwjUzhc
gP79gwkYWdVDzV071a1Pd4j3qUiQdB5m3KZkl4tUqxF299Lkh2BGiEOVm/86zsnIBtHfEnyHopG5
tnPhf3iObu7mFHtGJMW8Y9JHHEDJQlZl7oMjRDszSFY/+GHEK33SQwJjNOoW6i8x3Sm6BuST1JIV
NMnmBmo1D0BFr41YQTOAqjt1wWRs5nWepwzv12JS8QuamZ7KPtgXNCKdeNwj8U3AgrU0ButsScx4
SAr0S5Kc7XyUnCvtFDRSUdrQiK0YhCmMSOGrSgvxjoQ/ur3v6iFYZLZM8ZUtNQfAm/oFH7+T2Y9i
kBDQc+PZT5Fw3ZDj8RswChTYqIb83b/2PaGJsKlYb9PM4FHcCO2DJ/jOdzanbEEhJKHxwHwK4jCE
b7uzHIrAXAQJNUV6L6lRWGg0gzzMPjHJ5HKawka3DZRpmTJ903RNH4uBY5ct2OtH5Eep6e57vxQK
Y4A3D9y8g6/odI5+86zR6GqUkpqVY31NMy7bbJ2PQyRt76MRr08k7dmbVBppYLTxMjOhTjPZ+5F5
RRHkbZhxGariq+5Y6dHvSQt7x8+ROQNKLmQ8DnE5sd9r4tjOR4C0pTUvPKn9OSNlJEec0wFGdapl
DYGmIhhENYs7GCXYyhn6LErYFLMpYdbYGGOt4jh8CWrGxeoUXNdS6R6/LReV2rfFlpVfpnrym6p6
sEXzr3kvNYwA7B7XhHMt7q5o3PnSX/H1+o+IMgS4TMuFaewFDwhKHFRkCW/76tkgRrNv3TK4n150
kedhw6BCCQZLJuGVOzQHdOa6jUTzAiroOOTLd8BKcNXfIsM3sd/yndCfn9jtazHf9+f0k8dnQNdK
6VJ9HJFdMDeJP/aUAS0SH4FyAlh3QTUb6U4Ub+Cx/T4sYsYBhFaLGbRxjVhgcm3lGpbzaLXgJOxQ
vbB3juNB3DO8e6c2MwRtRoqlYCRe59vlIux0NJsDXurtEeOTh0mbQn6PeK97Mq7xffj6WIkPUCB3
obuzsrP1XRx8T/Kn8JWSBDivzfN+DZrACMa19k9gmtHlRpSDHZSpj7GItJqZUF8PLssY2cvcG/To
fYONpP4GHqZodo8wrxjrxzx63NGt6/v6pdEoFn0VqlW8shVbTe6gYH3nI1wulqAtoAlAyIhEQuAw
jDj/VqAmyHjqpCgsNdsL/1lZmOSbLwiXW5AmsIbYZmfuyyPwEXsVog6IUqxvpI6+4g3zEwpYIIPU
2Ljzqs6xdw6pYO/GOPA2hEM/QHfB6uqGL8gZnfIwQb7uktwTaE1XBBj7G1B9z4MbYAtmLjSXjAnr
o4vX7y5TROE+4LuwV0u1nn3B2ujRAUQJU7KR6C4Hyo17+ANpY0UAOUt97j6rAeS3SP4Ieqj0K2IE
IXxeQGRMFlIyesgdxTiYv5wt+F5MdiwLxc6IqU8HQpYo+vGkVai6syIIMUVdMk3xghUW6xHB81+R
wPkoTMfbOmBNuHiS+cXSGHbFKJpb5RX1pEKwFtL8DxYEGWLX9gbzfpFP9W0dxLvoqYKnXWfsmE9E
fKJvkfyp+bsdbX4nBzvDZLXSVE56wLB/lufiDlZFT2Z4espLnrT1LI63hYepM2dDWvQDeL9WIesk
Fu7mRcuS/OYla/3ZaGTubDjt0MAMxVQEFZIQx1ivVbyOQlEHm/nyzOVe/UDO6u/k8AjOAcZnE7Ah
r7WPNXafcTk3MQQqDIr4ZQ3ZkuhukbGUvCw5BQ47mDti5+9e7YXI9nkiEAW/9Z4jPgPAf1WCWpMR
QC+6teh6EqW6fV8/0UD2auUnJyx0mzZDkMCCr1hgDQfq+yIdRWs/iXgDCl8bozVZgAXSYTG5yum2
RYlnJiw9X0WpGtjIk044UpXkP5pLIK5dI1kJADtDE57XfCYvTXzxIYh5ZCv0V1gmZPm3gansCjC6
8G+Xdyr4Mg14mDu2OflIMloCZhwFKx7ZuGvILWQjAw73BDONXwiZeN1/jzRmqnZ2VJFSln377QKy
5/f4M6QQGIDhE2wpgP/+SR91VIJ5X82I919UUrHX4toyem7hKkQsXkxhrHvvsMiz05zOIcJMTW9D
OOnp7NjxNgBCrWUqYpl8K5g7Ost9g9ce88mttQN+/4Hqo0UeNsjH9eevdVHikjUX6l+1tRISsc9X
FXGIetUk3zDHmQJfORxg34RnWsb4KEgjs2pOLtJHlvb9ttDh99vIVwYDlMQ0SvYqB9f/OCsBgXgk
rjhj4fO/xUID9E7DjlXYCXwucL3XyGyiwwN8xlU0TTfcXi6zxlslma540q1DP8qB+bs3IBY7LskK
pbMtpOXxF7MMD8Uw2H/e8y2DOpX6MJ3wcvJHXGtkSOEl7FjlOONDAxl4N4ycAMZ2CvoJoeumGWRR
dMT281r7BZgmkxYEjq05Ugr20sd9QnV/8Sluhf9wGDTQhqnp8m1uY6VPOe9BL/1CHmXXXTTx86J3
QOqz7G4d+STxe+eWEjJeInP3KTvXo2UiHOfR2SkFb3H9NxU334RTF8lx1R2rBMe1VWULqWm8xf0P
yRH64aAY1ij18ZBYPVLKk/8yMS9lmQg4U4j2OLY6YQDrVOanoQ4MIsd7oxZIZueOTS/JNL+SiIsm
Swa9dHe4TPtOZ56pMpZefIbPiOPRLB4O9a67wi+O8XQIdh1HYXi82htJWmnYJ4azEokdTX1TRW6z
YkDapgww6GCmy7hEd+raqTsgskRqW4ojWyniJVpvfxOmkwS79z58RvdPVdA/d4qBR/Pi8FcRaiV2
tb7pXMuFQkiGtBsvfBPXH/1WC3KMirgQX2aGKWJBmh2Ga//oThXGG/iy7EnZC/cF9K9AuNxsm81f
vV9OX9HxaBe/PQKpt2f6EngwaoOcNfaEdj7VucJUgC8tEo9RVKoQkFOkZofKs/MyL2S1N1BOi8Bq
hM4uELKmoAYvbgGkYX52T1AxVQWTmyFZJ7JmLdae3e1ofS/6+UG9rzIpYzSI3w0jMPdN8i9ZS43Z
8OP9U2rEFx8EcBnutrrKUYDoXwrqaN0sI/OKPAphOvM1ONny2TFBKSzykoOUpa8/ZTLhTvZFBJp/
+K+Ojn3A8Pk+nt14xorPwDgta+o8RAPU9WBsMa4TG5wgpK1XH/pT5Gr7GVvKm6obtk3nzuq5pfah
Uk4s8X5F8kNQt8panXi58ZbU6Em4V3La4sneArQeaQs13gXjMjw3kbS120BKLRCScMhzbqDKqBIP
esfeBLp+j6Ie4Nv5qvICqEMhFfc7+oUYg5tTO/9cN2Ial47Kom+PiaIZ4zqaiLU+/pBI73/vgRLF
37t51woHzhKpIsqxwNXZXy4GKM2bGM1mf2bvkzHzvmPmT6LRX9v2DzNjcVx4ITQPF/DPOwVaM6kX
+7pNLL6E0f2uzCWx0OEkLjIgPKGJPTlhfBz2RjkDHkeJ4qguUwuW7ADvtMaN5+XyQ/Gj92Bg4c3t
ZRWa80JlbD7IPeUbBuCPD5NZp38m8YL//8ocxFjF7mO2MbxGM/kfgg5zgy5dVuw1AYNQpJ4ksDeL
faumCuN3pO6lpC0QqiZ16fk5dyeu3tO994uprFv9/PwuW/d44QIKdPTNOFboq8kJeWV4oTtGKUWa
F2Tp+3b6T51U9mEYPnVaLTm6gbzE2DVKSOrS2nxphYYiTGI4dfQduV4ZqGnoQzpQr2fWOmvR5av0
cN47wXpX4ZQoz4bznunqYUMWpCJvLejfnnSnOu0BAkeIVsIFiSr8OKSymxqj7pX4A4Y+FqPJCRn7
m8V3kXzOthrWmsTMboqMCdz4W8n8PbYwhOhavtFno5QGR2thoWR4D50aTP1hxQOHRcmM/QoI1pt9
aHK4PZEnK1nlb0snjWRT5dmMEtSYf5YKMJ4jEnsLmXJAow2B6waLwh3ot+ebVAVYDszflf2Myk1f
OX1RRLv+077g3uDZ9716KizqQlgSSr4MCtLhrYTOGuPvTvRUghh3aLV7Cos35TzvIEhrcrEuOGOQ
A2YmIMmvXch1rPZSBDEiQeYEz3bb6mlntaCaG9UVIrtLmbY+fK3uJQLt5tqMzG0N6BnC0Th035EO
9NNZmIjFbjhLIJ4d8ulRl8E+do4xN6RIFgDgjWH6pz7d0X1pQYpcViBhz0nc7Hzx5pb7xpX5beml
dUgf7qUN7zZxmXU7xOWMGkLGjB9CawwwN/W4Kt30VAjLQ6Ya2x+4nxJSxYzGXpwgrf1CUce514B8
Q/DPjPhfYM08W6tMlhcKbIOUhZ7PzthRmUYgoXOprzK5+kiUZ2r8A/TkwqXFE01JROWPJmVOTSNs
7NNDx20MLXOnwDERqUwCUl3HN0ATv23w/7C0KHA8d0t28frOdVTMUyvUmr+qBIOqcyYmRI2qKh6F
2gROyNwu79+LjvwD24zMorNJQa9ONPVnSVd2cMametT5b9/YX4D/1mBrWcTn9vtoWqfHEYPI9VjA
XijSQDEFgAdGjF47gfYLLlsaS5Oyq9v94Z2+L/+Vv5y3U3xuyMZpKcdH05KeOkMmJZoieoZA5kWE
VtyRsj3B39ykm9CwGs5D2VqKaNGbYl2Z5bzGPOglkwW4OUPytGd/DEXAP06G/ssjEV6ldXIbYMwf
CMpk7AXYCUn6hHxSbWfDUIyHP0vfiRVWdKG+jJBiTyl08DLKkP+per2u2eby+3OYxdVPXiRwf+fx
uVVMGukM+pbli5qbJ9hMwY/werc9FwEzgC0sSDJDksYPx3LSq8zMTgt1t04yGnLG3px5nMmEzNMQ
7ec1z/osyEJIStUn5eq9SQmZgaftyJEknuUBjYKA5qPXJVXg9IbN4VZjM4cA+lNEZ14fSvBywd8g
nH+LFCFWtTPKEu2hhbI0PSzwQYW38HEIvJviKMUukNg9lIIcx+8dlcqgWYS6LIK16PgA4AcMvJfE
EQ0i/GNlFaoKlCDSvdVa9GQEgEhQTLTZnD0vgBQ7Hc3W73hoI2MKQb0dxg/200ecPU3ong4zpaRO
EQGWnoNy1I9FUGe/Lo1b4poevWdje/hOzlTWwi2NZ2C10oZ1H6a748Amv7LK3n37mdFfPLmzjdgE
NpBnp3otOcA8qt3LPeW+DpZ2zQIhc8qMmXLgn/iF2/D/QCk2L62ruiyRua2Z9iadSenmyLZaRQC7
bXJbJclZ08qFDPlnvcRzgBfdQmBo1jQ/fVM80uygBorVudFn0qnA0apeWmJeBjVSWH7zJLkBY3JF
hehk1fy4Myjgozdefu986aZxPgUuC6YTYyBv2pS7FwReWCNgxaxNz28Q3CIwZgZt9sV4wJpJIUwf
CYBqQzZ/RELfsfFsk3ORsJv9ztV9CHHkE6tWAM971+k0/5zMydVioQVnuan2yf7bGEK+eltSrPdr
mIoX1Rv7RKzQ0rETSILtpKM0XWaKSGNkaYD9T04wCtOtf/ubmaLV0pdDEQ/KYYHaCwy7OZnMS3gZ
JJCj29Xv6yxk4+oXhTg958YO8XVSSrzXNKC9UzI5eX7P/W4JcxqQBPFQ62wRUvYVHBWYTpgXm/A0
sXJLezOnQt9qd2AvTtNbLZrpOWZl/gLlqm4vdILsbm+z5YXvxxvogmYtEr/gJgrY0HbR2yoPrRRa
oABaMY6oAIC4PlxEH4BRytl4cm1vBeXwZ4ieDEeNQM3D5beIGlx25h3zTnlltk7yQwEYPBP83HFD
nHkiR43e6yzq4v6C9Nh0WqYJf3MWr9KXPQAmcqroRqQJGmrwFrnnogSq9yfOM9mJHV9h9PNDrIAy
aJcFpEX9NPaEbm0nneXsf0OI9EruX+jB9mHkKLtMz5wUHQC5/qSi5Dx55eRrY9RLnhCA1Kt2KyjG
XD1B0Lynq/PWlZ/JVm1LaV+rFsiGzqvdojwFpRVG077OD22ti/LoURvG8p4rfFW/KwgghYnIPMxI
nTpauldBUREbg3V3UP1cLbS6Rhttr7toXzXspD9kaY1Lccow8IV6LBU0xseOXIKdDlkhDPhro7PA
g4al9mROpTzLIhjKFYVHndlUQ4wEAiqW6cbqlFjC1tdzDzS7LMKrkJZ2XI9FhI2WqUlASPA+R0ER
pJYSrV9d7a1ZwSRp+0YkkmQtH80bdR8jOwcX4XmFbbhjsbo5AAz1eyb9ithSrrtSD2edjEc5oqWW
k/vhcwIcOKcRUPcWkFp6B8A2zpZz0LePkCJn0fMg10xipOf055J61vu6u9ICzb9TSn1SkMORVzEY
YfLKk43muB8MwD7PcUJ91Uj7KN29HxFPIrL0w9ppA2PNV2B0MQqRK580g9AJlyffRpHnSjZ2QrD9
c1sq7fH3YtKA7MOUXjbwhBuY9rtPGj2NKL5sGQ6o93crpLRmzLRCV7Y1HL0Rshza1G5MrlJ8gMmO
lBi01a6j4iGKf/1STudnGsQ8/JaY73NHdR0OwBy8MhlFNNxBurYoNqjrQZj1H7mMriOjPnVS2r8i
JXEkjSfpj4pGP4GnJxcTNwc8u/uXVVyPXLXwrXII4TM5xvPFr99gv0GVyMYLSzVQVCOmDcJ58B3o
NHXV6+s7dfI+XDUamzALvehGoBNiTHc6KwcuTAHKrnZNNjUedIZtmK0Qwpulr6ZMynZqkAgLEXmZ
ey7pfTXBGiDHV8GNQDDt00MmhpvtfLfaFgq52R0VwIYqO2CUGeGCfI5AlzcWA9at3nSDT0uMW6W/
WxwTY5HenRnzFcnVau5UFIEZZ93TbKqkYqZgQbCW7onrciXw/6SDlbvaIU4F4SOOMC/KsPRoUjDt
A+tVae6iDYEKVOmBCYrcJvHctsF/ibL4JU+3vnhtxp4KuAVHhH1b2J5DouJ/mtLoBTBD8pQUEZUm
f5KE700zPZ1q8xrs/aStWEsOL/7WFGhR0MV8E/s7to9NA31t9K+82H/tiYls7EqvIJDEUvnc4ZnW
b0jdpHcvsdtHmGcN/mbBvKLjwVNFd5NxsiCsEyDP30+LB6aJ3HVYv4jmBQWBDx62+MKt/2q9imIK
nbhGDjzw7W9OBNR4iIQ0TfziiJdLSUUw6wyVUd+zAtMRHaR6xRTsyjuqjJe7ZBmHc5JazmmT+amj
adWaeEkASB7pM2duP8oYl4HzeznfAmlqNJ7CbiqsTWl2bA7HJ2ecmW7JZlfDM5iYp3J/6vv/ZZAF
5FmCaD976fFyLhHFjQJd6iVzDeZzNWqoxTfG5vg3ZJ0BnUFLmqm6AjSFMokCXWjl0FWfxjSmwvDs
mBovz0l8TbyOQK9+1/u8zmWHgOpFR6YtfF4sNwXo/WKn6CVWSxFXHwgeyvTXew8Z9NNWTqa4Uzkh
722Ux8Rsti81/OOQRvdW8fDlu7IuI5GRp0+XL/tbR39bUBgxudt7Mxnwpx8EdISSQAMYBWzPWoTp
f52n0sPpC0GahGf2ebvxxVtHtOFO0aEDyEg6dbDGIARcHgLP1qRx6bquB+/1GeTOvQosL0l2FbCR
CVqmBOvwFp0c1cIHZ/+fwsJibIwbZiLrxrjtBoxnt0CuxFh92wc87ejTnwHbML+mB8woyRQRZtsH
cH68ymV8SKRmeWQz1zQGdSD6aj0ELc+J++nYhm+DYhk5BX6ywQX3PFtQ6oa/5rpyDCsy4uo443Gl
wA7aYPLpq8RsWj7kHPZJTtqw9uoM225BmO+MlR1/9L8MFt0cQ3w0agfDzChd51qJ4IIF+QcEDOHZ
UjFTIC7ookZnVq6cRVE4rDYDFjPpw5GbkDAtWLJs/UnMOTboWTTwKOLiFlbbfrmD+Kxqrcz/xj3H
TAKNz5eH7rc3Jv/01MawBXKGTx+jG7guKySd8K7P+gdLUKsoPT2ToRoS8uSMrTElyAxE4vi0WPh2
azoZ6kN83FWN4thL5jtxRs8b1GgROvWFckRAncIm/7Tyt7guvwrjJtGyZCEiUdi2XWj9ZSpuk10D
Ugs8EroPTgeojuWdKsFBARUxrSbJBfYNYbX0fvs7cp54WsTWGEmt4LqSM05/hX6iM5pvOUTT0xxr
GFo0R0MUNq3gjA4F4cxppF+ZTkje1qU/T3YlxAQGPNmx4EqwnnsM9J4zs6mHSbdPyKVkTdoRymfP
/buONATyRAfzr685yjFF6pg84jJU1rhrius7LQRJWW/9rD8jc9v4EvlOXZP+4E4pUBmCYHsqp20I
z3MIl4a1wFbeBQ65gWBHbrQHYvpsZ4bc3euP3F013VGY+zf5tvT7IY8vQT+f3pD//M3pYAPlGVqg
UgBXLh9AspSiEan+/W8qakWiZwrgVcGQOt16Zhy44MFvnE/xhmMftD/8H4BiyWUFhDWyAKYLEy92
0JtzeA1vs6P1/3wr6xJ6jL9m/GXzMYSKk/qldAQIv0hsma5Y6IQFq8kaRK8/A+tm5K/2/9LjBcdK
kRbpFyTN3WSoBQVVYO//hs70q3GCGBGUVrMxFqDB7WxbCw16bQGM+ysKQ8UzQe5o04XgpLBiI1Pr
DiWHsH3VcdZwgKyX5JSmcFANcGtVJEPwxX9x3QpnmFLHGW0NzbISk7V1qzjnvp3LZUNzwQbGh4d+
ZmnS4ZMpPxfHWw5sQmdfVuyQvM05byePS50EEcgwedYr0drgboV3Bmik78IW2CCDvNwN1WRDuUUJ
j07TQUkzCtZgkpF2Yapp2x+j6hZaAGHrlHKV0dqUfDOi8uMpIRpXh8zbSZBAlht2YNWGgCkKjO04
3eSQJM4Pat8muNd5kVk7L8Ma/SOWChEku2joFNx50xwgy63WVPVFLdWET00iOzioBDupjx9sKs4N
HKGrgfst6mcEZwLjwgyksa/8RMzcvUyeb2Zp0QAR7B+eX9xrBaQadBB5bB1MzwG4rbHopKHQoQkw
xGF5nlAp/39lMCOeAEhOHq5zx11FhyjCZ5gISM0cHGNwSdExCEOfP6PqJQK6s45V4lEDtMmVzxlt
7MIRP1IblhDoeq1XoxlwY7fVXxD37MrFdkYPKJQl7W2ra/W/mrF6v+G/i9pVopJG2jdAjXCu42Qw
WWUfwe3uZBemjQKJnNSS5lZqkq4p7MeIYwnZX4txClFTkr61Bf0NEP8t9wxQ6P8X+MpSqf/mq5oK
305NCq9ziiwuhHZT4jrx4TP1SBbdP2MsGQJYcM/Ei4F08LizjaBtDErfAQXnHsRIQZ3Zph381TOk
JOEbBHQ8zXORcnbVPCTP0oxrnULJWgf6mJQnrkyoUmQGOwbWrNj3BHySD+A+grWYXdjpDd8b1u1G
OWxZDFfpwVG7kZEUSCA+aR3VFkcc6lZEEp3bJhCcYdX7vp2F2tPVkUY6+wO8rOM6VQj0RugRfC6n
Azg5Nn+IvfAU2yYujNV8nINO3Cgc4y6auLNkMl2iL5BwS5GE1Di++AAK4CdytF+pl7CyIMas3Lt0
U1HjdJ0WG1pOBxWwGRXusoP94TQ2QTXJkt6YeXpQaY9GgessdwqA9pPA9qHtYbFMnzd+5YuO4cSC
9Jwjs9dAP3Jv1nYcZeMRpNU74cGLDz3lsyZ0HnyvREo8lUb73/i6lthM8LuXvGB/i6f9iRr/924B
biz/00YNCECt3ZWKKJfc0zfmpOTCxknnc3d7nto/5/VBGrnkJRjNmWAWjJTm+IeYsoLta1z36vB1
09VmQEBHtZAUQybPhqdhsvf7J9ZFuBblw3V5+bnrohYyt0Ylo6S21rkoSRBXYgV/9aN4SsZ4ag0D
K69X8aGViRNi44HKjXYpElG5Ry/F+k7rYKpSsNG8xjUILndQkZ5GyjQREIBDtr3dOiqh5/SwlxPI
tJoFJrpN45TSAxfHqn2hP4Mpgpo14diWvuurFNTGgT9zhhIBFT9dCYwolcHcTKakf6+K1l47FAZF
ghEV+jsCqUfTEB1TyNt2ZmZH9WBiPE6SNI4Ruw8ei3PMTkYVlTQr0bDMXuR7c2V8RzksX4thTwiG
OQ96APONNuin8x8jlDyHlyvCJWGAPYpsD0VHoIBtAm85FhLxZItuijODuj9oUm/aVExUoYCLkP4a
zZF3NRaXnIx4Qt5E16GM3NZXOLWqILDl/+8cvxbJpOVEt1uRXcwX6lk/4Xbo1ytni0K3jlgPF4Em
mvlydJbVzG0iOPT1LTtO/ArnKltz3WpG8O0go1aTusANI218xkkCkWvEssfWEQm4cY23zc+KcuMU
e4gYa2M1gZhP6mcrTvWtUzJAnAX3BxB++pKk84bJhM0LtCKPJGuhFLoo5BrvvzlUSgU59NZ9CLzd
lts9hUNzyzUVV8QLp+WXTS9Hw61ki1/xo5FNgOfSD4NVUDlLr3Dy1XsdeOy/0FONPfhXFBKZTuo9
taXUxwWmO07qjEHKsXl6suc2BYoRVcfsg+VVTMAyXlOVG3Y7jWwvuqdpOVZAjfiRt7Ms/yAHfRMe
HkWFRaYgC3sfROUsiRJ382IlR/emv1xPFwEYYOx8k45lU7BkC7yzGWPm9uKJ1DzIbL4/5/R/FAfk
J+OSD/fTWOKw5pwsam5rHnXvjd2xBtXypF1pJDH/6nJkylTb0cY1oOMLJKdGrgckQAy5gW3U/zOy
fHb62j47x4MrU6akcnaF7pak2lgQDQuLbD4JDmHo7EOZSIbngl4OgcZjZzGR+aBJFvSLr4oHMMgH
GU/SUg7xzbnSAVEQen2wgiqwZVXg/DPGglXlaXKnXV/sBUlHFi0R2ybCHMnxJFvL8B5Au4YGrf3E
k7gSVu3yzFuXmHbbxBS67GaTy9o1hWuOaLFFUN9VkZqJtOyroAAAiItW464fVUzDHu8FryXM8cfW
z4y1+o5ubwEBljt979Y6rLLRTqfhtIwZtP998mFvv4FTpeZ45mec0RzINwy/GP58OuaRqVi65+2C
Y2a5G8ePhvOmq4NbNnD8p2v3l6u5ImbtHp4da5uX0iommfHXh7FHUt7+DqGa1m7ORhccntcXbB/c
upkQ8e24vVg5A6p3tdsBah/rnmVQ1P2SLYGfcnBtJ3YuBLH7QOkEFE7PLEX2pjpESk9ZkuKFZEJt
golxIqiJYTPbgc01ESqg186xImDU1+x9Vz4UC0Bx3Es47wb9GdcLNT8at9MeU22wZWGXVMwa1EUs
FedVzBn9EeG/vxwiFoBfA+pknmfUIbfA3E8PxmmNxMmxmYy3hAxCRZDFql9Y/GjTzvd9W8bDavWg
nj1hKEt+BFRUtTNWKw8zScMGbCU6TfUnlxPTUqrfscQI/1e9A9nJcUrttJb869aJ1JfOL1m/Fysx
ME6IgmtOgb0rhL5ZCXb77+HqCPNSvLKwIb0OFJB2kBV9lXNsqXT8g6JrpL9kiN/xpApWXr7IIrfr
flE4KUE4+nRORSBdPok3ZlPhqSeumomsmO5wKhuc9boD9pBTTXVfXk9CpmLLOkrpe2P/JTMlYfkz
NF2bHR5QjeAPVdRPX6yMkg4fBVeFdME0nX+zyCby4nvl0sBourRZE/sBCzVlBBZDOqlcwZlY6NEM
PVQ/DluzdPiRQYJPxcHiXIEypEIBz8xtF52yhxzwvO9hEOTiGBhcwi15IAAU99+eIvMOG0s0lMQU
vgFK4U0vZ7m7IqaJQroAF3LCXvo3iP28T02uUjLsLd7Dj+fa/H6TIsk+yEqPDZIAgHOD752VhtX1
HI5SKyXY/TrYtHehV9Azbk/JN+2xpMV/g0knhO1oqehfBQQ99a8IEOkI4waM18TJ/XPDL3jDZ23H
5feoCTmO+WZdpfvKTbO+11bFBA9EYa7KHrbWuogTO7EXCXlhlrCajFDqbSofyl8GYzviyuK7Oq6G
vtU/8NF3V+hJ6F4rWRV2RpG6b0Tf9j4UzELdIXQKxyL5ENUUb6XQGeGH5NCp+4b5lKnCxDUSPp0W
UHgKoWNHnznMH0F09w+jp7GduZy35aoMxbCXRX+AfeynGwCoeEPjRpGNZc2o1KTsnR/oRTWq3h7z
U7y4GXerG6q3QA5tejncIELyQZGphfpwKkXlchlV/LnA7TfMD57hCXPZTcOypGMVXHaeJFnLnEvy
4u1O3pu4d6ndnWlsZXGmeSNrBvgwBS1kQ/NrEUwcEO4i8bcr3K5WKeP4z0L5ogdbumwIQK8VJwq2
lUlpyxzjDnsyUakR8wBRBdnY7Z5pTzq4in7SrM2HcQQOLzW4RHuZLA0rmA6FQOI7+siiIC+M7ql/
iCRnr+LfEh1Rr3YBbiCsaQ91z5FedwzSFtnzD+Oq13AzsBsJ/uK52j2fijlJdiBv73JXVW22IeJ6
6ggLwjZLdH3A0R4n+T8l0EmUsGBMFOJO6neUB++e7V/pVByjeVHWWdAkrJZXjvSm+GirVBeCFVXS
9yd0U7wCFyxUHObkOSYoj6eOssg5fHzLDEGugqny8xnEddhIFD9cOkZk6HZjMiPgxycA3bmTf9vk
9yiSSXK0sjqb3ZuLV3nnh8W7oDS1mam+KvyCYUNfHtX84WKb4GezqV6EW3erTynBkmvMCVBJUGGy
6Tm0agNU+CxEvlPudHA3cWTE/UhAFOsu5AMetfMgXAkmLE9hKyRmdZ5gDzl0CIWudI1Bq7xixCmu
HWJNxjTJPdLg/1G0AoKYoONaRuwReiBslwOvo0gQn1Yp2j/uhGDwqVshPTVMgp8jIbu/IVuSPcTh
FLxQ966OPl1xd1o6MyDNW8WnXJcJZQHE1rM/gwE1/BXEoXM8rpXGdNUixL+p1Icp3vWgczSKjKNt
NrQzfNczwMs+PVkJou/WbXlxzmmENhhuvl+XvAimRpcnWvX57C3m0FnjlWX7FL90SeGf0kpwjJ7D
lvhDVibubrPzMda3Fli309niZU42AYlsU+IFXg27ZPcq9RLzOOIxK7BFY/Jt/aGQ8gwjxVNgOFFd
vm4WMfU7Lcu1glpaR76I8jpsfhFoPIeVeq1a4wMDME4fE46e6EJZkvqGB78RLLduitNq1Ko+Et81
g7laF8a5vjkWpv9TWtPSzYZNqwPOD4j2fjbBfhUc6EBXw16Fvphvv+qPjMLlQlVp0m2oebgXq/As
orURbkbwbZlmxyuRJGVEkjOQLO/TfUJX3L9IE8qatev9D086/WicKOE0hXPkvoUhntC/UGIjyE+C
EuQnQldaZMw5jIPnEw74m9kS87p8sIBaLoMt5GHqe7ADAEgIq6muDt30wmaUz0kEY8453x8qu20q
lQ+1qhyM6ote/T467o1w2CyZhCYBnDaTKGigd2if6ppya1T0DrGm80xkTXSBtcVj/gurnQysB1wc
ED1QXDMJJClduj9iK9YFQy2YvLXSTt9VvE2SerU9KS9LruPynhhgXLWfkasbgM/bMsGWJ17iRj/7
wpB1Cz94pEPMnaRXr0uBSH2VJEPPgQzty0FH1YVcCY51ZJR8Oz3uK1Y5LUAHGVvP2IHuZ/PqWgP7
6zHqOKv0yC6442FSK4qPiebKhXv+xfsaalRrn/2OUcq24bPtxBGP0lI7b54T4hCmVCXldltLhNmG
qU7Mue5cvpqYluQ/QNlD0D/YZw7Jde4QM3E0V4FSo9UusTJOte4AVFcbuWrOAcq7DIG3a0513tNY
WNEnp17oTrzAOlAdDWnm1JsHDiMYgXlNd8R/MEsrwUBZtUqNH6JLCjHh0VzjX+fsQVMOMNVnFPhR
a8qAHK408ltdUFToRSnIaM4jAmtom1Sr75FY5wClrX6gnlU7M6U/kBq32L0O/MJM+g0QtVcl+Ax0
1BSxLgZE4wDEN3bnwHolw+PuwWkzDTE7bc42PxOkXnfA5/GGuZ5zh9C51UZMQ5jewf7HnTTsA0EQ
dlsq85MEFUGolcu5VUECv8FnwjDdz1IZNHXFiuZh1nJC+7c2f53LJPPwt2qR2sXaDEYk5CvVQ6fk
M0u8rCuJLRRmDR1pk8yHaP/WhDKTjNbwCtC0SQBAAPYKEQvHnGnH7T6PTPEgHb8IYsXCMp+U0jUj
ShOGGf582NN2KiEyJRS5bfslW90qYkpSillTjbdpqXbRg5v1vfsape10eyRv3hIAzGCOuRPA5wkC
ie0xG/otHoKxuYK4SH0B5P3fqgRr9NMG2Gl48GXHiDSTvStRktTkfwCT56+KqOk+OxHDPYv0Ee2m
8pK53PGbRmZmoXtRhQCFteZVDg2EFnT8/Hr9tfOiNpg7FV7iLLCPoXTDR1z15Z8riZDhgECZ10Hb
lj7Xr8MD+HODYykb7AbBMX1yijHnfAIjPPOh3+03ljfW+J18nfGHxsvO809PHu9QE8VGp0O4pEZx
NIWPerYb3T9jZfIHKQDmmKAiNlbqVjUBGZd2itPuycH5iJI/NWRBrvNQmhppROAO7IIPsMv9QVzn
1T4Z9sYCJ3fvrftieZOypnYwJYCng+kCQvSJzn/xpGCC08c5TLBAejtP0n7T8ne8Y8bJL+u6krNM
6zgU0SXnGy8FipdYeWoQeuO8Uw10w1sYV3+Uvfo0nCkODDug6y/riXyMwYGrngm9Oij5E3nlE+w0
br1evQhR9kpHrTUoJBeaFodg/w2d5luTvwQ6jlZE8RnONpC0P7sA6QYKeQJjs+sKztLaX2/oepzs
k9CPdkA7mG/Hc1uk34kFjRXiun8wfTmQXp8aah3968BNtBeq4kCIk0WRasZODCD7rHjbtZ97hrT+
lLKknmJ5VQ962KuYEhi1He3rHDJs2DEjNd63wtO6NSyPAeuG8lFLnVcaGg30EI2mkRa1zG4dF1Bv
aASwNtQ5W2qKvL+h1SsY8fZSzg22CxrevyVJxxGcfPGahygGXasyhg10EBZIEeqeLPVRSyxnvsci
SUIItRMqNDAxwhRboId3YOn+NP2zj6Q+4JmdTpapvXHTVlXstRwXOe/88hmsDZ6x5Uom69yfutJC
w0xsq01lU5CVvzAxJM+/gCDeejBEskNyEKPdl1TCwMDCywrumyrUbH7kLPRj6iYdKPtqplh7hm/U
jfx3s4dcDX+IQcD+ENoJGossFZVUDMqEYd9Kwu4trczLHUoaUHTTL0elxGE5eWmm//bH+WPIEFRL
YRtynr3Y+tMG61YBBTFt9FVIK52ppz8U3ziDv44AX5PPveBA0dZHlcDl530/PwWy+mzJmeRgfu0W
Tp3KOVWamw6ga2u4KdXaxs+m6p87DR1cSsU5LSXgKCS6enYMBx+yFFpqVb91Lx3oBDKW7ec10Xf3
+jdGOpMd68onynbuXHGXmzd4dj7yqXRpqhszT3lLjaxeXUtmllnmzHrwIG0GkOGgD/IQeXd9ikX+
Fg2exdscVcIEjPL49kylFfzlk1kVaK7seTVTevuEl0EANK24ygnbUVtxdiPz3H9O1y6Ey4qoDjmO
PAgb+GFhhWvpAOj8yFobgWB4NbgzS3+16UigC8fZNeH4nUw2bQGzQ3EBpVDy7bA0gFHeVhPRWYDE
9PlXgTFCj45QQGlkK58M9PG4UDJ6r1qS/zW7biOBKYUIty9dLOv7sXAIwUmFVzMI+E7Btjx4jAaj
2X+fa3hh2UijyhDnlDakI6udPAqqZgnAr4EwA+4lpgWXX04utuTgTzHR4WEPSL2dU3/877dw6Y/i
XELpVRkgPAwyWm83wOshGahg48t5ZcZNXr3nnOWCNIvnnj5y+GPMrzMAaFHkvZLQ5B4eDxO2Y3Gy
BTGbiaNIDLTUuz+gXV7fxSkTR4H41g6sFOBCIUlbh7uhv+8JzTrjpN3PyR9ZPzYxzlYK2TaqxcV3
PGSr21HDeN0CkTxqPHTDXPFNaNWs5M6XNNwxOqCvebGunHbzI/g+gKmMOmusTEMlDAHfwYA3WVFd
H9iubvMoRh+saaVrAMJik9I2BuWEHYudA5EXwz9hiwLLrd0ninx8VpTX7WtsRKuToFpeWar6CrA8
NnILhc0xGeHJoeeM7ZN7rdHMbLMB8xuSwBPNPUlZ4aSAKPNfr4uVAmPHQ3jxFqQaXWODfjHH1DVi
SeXn55JIofuPobagJJBdPWawzItHfdYtyvYpVlsqk0lGAEsqA/CRjmll1qDK+o7KUj2XSsvPppzI
SvXfFCHCq8ib5tZdHu5SleAbjq0rmFNyZOcIzac1MtCRRnb8j+3QjzlCgs10LWvr4lbPHk3lgPt0
1gUQI5mXGR0M2d/4I1Uoqtnp5iNQ4hExZbzchQpE3G+oQ7+gOk+6EXbkQ/yboccVHKoZDMV02A+m
UE2aeVPpK8Vkfro22WneWN+CSzJHNM9DiLTgXS/VSMWZcALeBa12W6u6VuU69yaI1wpevtZ3TxGg
veKqJkTxzqwzXH6Du5kSClEoHTNcIymIxX2WYSGJzcDSfelWMVFDxUNx+zfvtwPrinpgtdKcMhwQ
JpcpPeY5MI3vnnXTnQZOUXWCvEF32fvsL1MwYYsb3gnvHwFZdAp0IDzHvMzWSL//pMDPH2Bcr05E
i9yOdVpbD5r/phrJl0wRRyRRV62Aw4DfQIkTChcwLB4+2IVS1E/LFOl9oOC3OyGl12xzxLPT7STw
d9255xv7RiV6Y/th4siKU1cOxYHXwn9OrNFThjew3Bjid1ksD89FC2MJK8E1msKYTIWfzRyc5qZK
pUe+BpSbsogs+5mJbs4D5N/nNogRS+cQGQ3Lfj0M/odbDooS+oQOuJV5qyS/kMfMuJFtMmiU4bpW
Tv4rGgvFfqL32r+9m3NxWLH4uj5F0xscyFM4acXu2ehXO17VtHDesWX1JokG7yFgXbAgHL/BGHDN
lO6o+7+oE3BrTshULpvZ3ZJ8oqca3tgh2V1sc4jjxC4Ndvf9BYXxaiYjfCslJV8YTFblzUQe21Is
uO8R5cky/Va0kkr61kqcmQnyFOUMdMx8ABNUPH3gi3/VS5b5wacpVUFy4gins+ukLjCYeboNr6tT
Nkf+A6M3aNvNLDM7WlCKQFeS1lttHxUNNAbajv0mPDLC15mw25nqkL5rBrp24IjyOQ4e+pE6x14y
u/YUNGRl9GlGcGpLv7RMEz0mGZ19mRIh7s5iYrAV/nDf4ma1/lSkCiLyUXYpq96yMivdgPVcjEpK
attbYeUSXMTvU55Evxq+TEIq+wSjqLcmfKSqYcxx7ViRnyzPMF99UeLTGydhzbknP4g/g3aKn3TC
dDgW+m6H8aSNPeqJVGu690QGnoH3+d+cD52u+EXMBN6DogtcL0y6aj23a1G76sQTlzh0PvVhFO+q
cNMa0jrH1kgILHiLlFP7VgYgZDRqCT/xywPUsbrcjmUIWqDfgcTpiOJ9AsCmhh4rown2sESHrR+D
5mGLPuxMWY1bIHVApkU70DlPLvwuWwh5Id2NLBkpl8xmlTCG8oyRGxA2d9qoiqSxLh9Ylmxmzy79
XQsahd3iY54TWxiiyfVOFE+L+2sHwFepKYZUoiI8M2+9H3ddMnEAyTKkEy8NwymHjFVD3m/eg8mv
aC2w32iE9ai0MfbCB8GIa217AUfpqohlnhD7nDzDMIf3nhkGWAnfI7w7TXsfFbRJ+6Lzle8YxCs3
FvXgh7zQdvUeoQ9D2gUxgY7/O3KSIX4LDvXYwV4Y2elVMgRrTk2jC78YI4P7IiEqNjHpY8sOeedC
E8Un4iii+qWQb1YmfXnsnBkmBlI53DktBhNbr4Bvpnd6pEBhcOLfGwbe8PHRYaK4v6+Fw09hG77A
lC64uf50snBptl78OFRJEO2zHbhUdjSALAsPTWamwdvJLk2G03KfBDZ0bwTd5Gqx+rYwqZvGv5Bg
0KQ1rJ3G1/3YWnmhI8SAi3fc+lIq6S0CMt73rZ1f8FNaA8owTrw3bGlHDXmc+85A0OmmXj4CPVw5
GKhoXPxtIFEkcH1F3fcGGs8RAMw+U4vECouFn+J2qIzuk8Iafi1iivhmFEXm/iU0GjUWoKo8V1No
N3JlL+O9ZU+ACr8fruAh5PxyAN0SiVLF7XueikW90ujJh/NnsfKUIG3QvTtng1vTSUY7CL9zyVOK
DN9j5KDwPtYj/aRMrR1rIJbrcWNHOVfiIjpoQ51QTHm500dribxC4ApihOZPxija929kDLnaiAFp
VrgOO1HanYTbUOWZMwqkG9SomLJhKErXjevULjSw5/VUI82OQhyRigPzfRnlq9QNHqHX97EeyFkL
QqfQllZMT70i00r5lGJmMuqLr0Thd6Bq5d16ftdQMljg2LG7UD+c9T2SerCR4EA2YvdBsQpm+L67
2+hudghA9S4E7zlW9hXH6Lt5qEQQwXPVJQoXrlLiib2+8gRbuoOMTGuIU4xTqM1aD2sbVWwSJOBV
U3HW6NaelaI9w3wTfu6QdpKvoIaOjEivB1t/62BKFRx5zB1Oe2lMN67Hic05VonJOhNRDRUZPdhQ
nOhiYGSdPpAQp7fEmN+Pz4XKQFC5z4KvtFH1x/5CrRZHKwlk4172PJFIbvjx2qsbLOt043E+UIOO
mycelYN9BuEsMEjj+rKFRUstzZFjl5J7HrtQQz/7Csbub6yGrKUmPh3M1yTgtiQjSIboZqZfGrwr
2wPbh3xziNddgfpjxiaw8ZbV3qyHTTxgsvcrSpkk39DSQe4dAkTZMgy0cpHn+mmHQKhR8hrZH8c0
6yLYh8EJBImhMJVQNPVfpDH/t8OuHfLuP09vi+FvVtZaI3k3vyFT+xNheGigAxiOjdrTL1+tGgAr
n3KcExPGIdXvL/q6rhyxUGQV9SVjSGsjTX+s3v1oAXmIFnA3eUbtZ65d3t1az2vRra8jVhGGj08u
PbH46Ab2FfFrn9ge8xks4Bxqt+KW4p1qdT0u3vhzOZNzEqkecITzUXjXcOuU/tOf0BX8y0pOve7O
dIvKrbTDCWkSTAGnxhJzf4Yd64dGCiExoOvwzsZ54GlGjgjdz7+gzu6KmsSwLkOzISUjQopMKNoX
9fsKMsBICU/mv533rSlKT0Sa3gPfpne/D/UosGn1BqJU9KFo5YuDHirzcdd+AWnzEiR59Dyzdj75
xKxEBdIlo0wL0UFiFO/5yXscTtFtHiyArNt+RHpjxriYhlrP9QVStzfxEY7ovJl1pwsuwfhQK3x3
EqZr3Ca5N7WwXifJ8URWgrCzLun341iXyLniMkmcMF6gCYPIqY7RgfCV4+7w763ZTu8jFdauomBt
D3pmt54vsib7K62Y4Wd6smkZrkdXp/E4IoqTSqXbuxZNHUf0eKmbpb8bFSfkjXwQce7SECoC7MT0
Z/2tgQ4UoGtQuy9jfB3N4c+mrAf0M7eQyS5T91jBKuW7fiIpP5v68jFnLf/Zv19qkueb8RN4K0Dx
0btTpt8CTASUSvXAEOUx4imOPHo1nQ7p0+5w3QXwIFo2V26nyGKv3t0csPNzKMywa137c/XXdL6U
R9LgX0yUJr2GhJYfZchCRCvkUoFEPG/2wEiG3nWtOxWnoKeHV2tqBGxWgQZpWsEsXsWdIcmS+R3X
T/FOKrF0I3DEYfhOOJM5d18vMpqAX4LSW/KXQLn4AXWzTxfT61/haDYwCNe/znTj5BIOityiXR81
SfIfKdgVU278/GYobp7TfaCC1daRmJzYIScbQclYSYHyczEVLP8K462tIS8adgySPLB019pApgfo
KvVaifT1aFOluPRwv+RtCV8hAmikFL1+d0av57XqCwHU/1/CAj472NhP8vuES/NHheCTRtjOte9d
I2mS1yZ4c8Fx4FgXhEj8rHK2VgTNGyp8ce1RvNZ+arYkDaBV7pFL6Mgjxz8Gh0B6yKm1JWxW68tL
blH29BPCC/bF6cxFq4Mblo6rnegN8R9BLlB943fL2/cztpExbwWMboPil15UU0LM+Ihw0/KXRLvA
d16sjtoT7c7kQ7Ueg65z2vEjzWk06mY6vAEigsfAP44G8SGYnkIskc1MfpCeVQkHWujIZy1dcZI3
U9+HrV4Kqr8yqRSG8RPqdbZOL7AtSf5LqtkTkERDq0fxBGGUrsjSFOL3J+yzBuOlalPvPqNxRY+S
l0fpaKInfiG6ZEzB/gavIJuNOMjpCM2vkS3xRFouU/wyU+LPQml6YggSxPkXE/1MyQRtXRD8liob
QUcaZx0FEqOxRzrV2dmGmxp9roOBTMGrE4AAunIfvwXfA8X8uvzAfOLhoLanDir4AvE9dEYN0jln
4kwIYgu1OrxL+IEKdB0Z1e+1DgpHh6MEG6DIMsSjdzP/mRciTvQfMvusfkFsSWK4WG/drtsBN4vB
FnpuDXEyaZDtHi9DRXv0qQiulxZu0Je4G5S13i12KhssuOFwtodrwMG/sXlUME+8GnrreGH29oMb
3YaTx3fCxzOqtUQL7rkMUg3OOhUmb73Di7l13IFupbjWPIQO28iCjkDNMa3e7ILuuNiWN8dLKIvA
l+mzLAaQvEPa2Z8ZmwARpy2+WrzJoCO2gTTuExzYUqSKKtaZDsV9WD6HR937eDEazqiPHUPaiVSu
7QEYcrxKUpDF31/tDoQSFRHj1WbRmpvoTdNh/3gBdIFKDL/SD9oZYlPZ5Nvriqtmmk3PXpkxrTX1
9sWvYLcu/qoQsPTKkf0Z0Yj/JFSg31I1OfWn3iXW829jYp5zVnAxja0W3NwA4S5frM8kj6tICzx2
W0MNjyZvtuFxuHM2Y+w6z/ZxXbQJ+BARw37tVicfWUYrLFq9oO9kgu85xgSb6RpUrzxm5hAlg8NK
tuDDWI2QGDAjvWjd22Q3MVtAbh3QntGRcwDiekv19HcV7XcET/qeyAgTGwgyrRHUrmLdi7catGyG
1Ydr8VLFI0Xbt8h1W2fm4e5TpbVWl4NCINuZDRYZ+u1NLWr2enlv7jv2papMILl03G9umBotD3r4
u6s0MNPkmwz9eH6y6axvrqOUTzo1tp9vWoVUBuQWiqmI8+o9wFQmlmSawMlj3ftidT1rYkUdH8/w
TWIBZIdikosZNPNQCEnvsDtsSz4ML9SZrNKSvkvTD38zXRgZWEg7ynIpT5XD0WIIvq/4hZTTYylI
Uz+AM60eZ53U+j+kBhV+SLLKQIDgg9XRhcz8NLv7lngYykunorTejkD73pd9pM8w7WNmscUufAxb
RkhlSt5cIdzcw1pMoFSowy8mEZP4ReET7XnVWabtDtRvaCdSfAdDnPgr+NLCMPp0CR7jB1c7skI3
VPKJ8Ia0HQXjxlVE5J093LA0GTU1R2D7fXQN5y7ZFj1REIRvI3/v/RJ9vsCwTS7Yk/B//w4nO8IN
aL0aPtllp1OviA7kPW7LCFGcqF9Tr6ToL/3AVEpIIr4pbhhTpomx+GQbCfKet/iWSEZEcwZH3Epv
f4ReunmDI8sfheh8j1SJq3yTvPKXBHZahVuizu3gzeQnGWz5+EdU7ZZXXjOtdtrcCGMP56r/wL6Z
5+0KRdHatbD45c/2hTVFI3DzJVU//FQkvMgOJCEHjt8oipkjI/FeDsWZc5nl/a68KGiiSsVhrJf7
YCKZZaU7kjq1i+XRgZDNaZKKYz1tv/IrvMMNiartTg721L6MKjvqLXih6FiAt355+fk4rX7E4G4A
dk9LMRGKaLq0TjdqCYPgUePo81I/wcR/vonL2793L3eBW2A5jkIZiUk2ePadmbEyAymS5vIWCC9L
WqNtdKrQ7Bi9waLXXZKFV9XMPH0U55+BfJE5ajDaYmTFghZs4xUWOPggVTDwN9tvd4cliwlzKvYL
ORqUJVEybVyd2nemOzACKVXvyqpZMXtDym9jRXqVKsQYl4UtWBaMHPS57r0SCFPA9Q6cDE1ar1Jf
l0pPrBFc8Zp3yr2zruyTWnr3xJpMHv9CwBohBYoLZFtGNf9ay0Re6u63Iep/7OCx4FW0kqrxs9Ro
mFBYQthfzaMTGfyVJci98bXORvUqCRoPDqB9BvjfBGBleFXp1/pIcIl7hClwMzat8kOez+kMOUMk
eD7P4HfhlIxa35ib151+2jrSYHQDjZOlxQXg9A8KcAcCNVMpAf/nAK17EUUEwD6C3IYPOUaJRXf6
H4MvSGqevt00EHvxdiNNqMUuSDCpjrECS1D23VVhUKYSQ9Wsh4Um6HQWjaV6cVMPbQLsBRSGbXXI
LyDgxQllHW01mJv+zWhtBuLCrmBws1Nc2xqm7HUIDn0BLk6nSTSb3CsWvHru5ehhTriNOQGkQ4oN
AddU07fEvH1foji3fjMuVQoDwlhoirFIV1ftCUAAXS1NBh5fJAEMjmGpKdjB/A/yPp108m+0acO2
DLK7JuR8yVBJiHeZdsi2zMs+MUzmK3lEwhgC7Rqxxj6Me2tlc2AXfQ+jZ72m6zT12iMznUegm1nb
zJZtG/0PPqsmYzKn2x2O09UqekQqjB+2CKcO388la9rgSVjhgUxQPJGMLIl9quQz+/Izu+TROhOR
G8dPTcycpSGa8mvlH1x2mXdcN74QV+6muX9Q0usrENf5hep3DWjbNsdqbSUDrg/MJOBifehODYFS
EiVRKjQEQa+gACw68jmgo8jYMwHqwwDymKI9p4F+BhuC+dPzAfdC12VidIPkLsi2IbzHvVIFWgPM
Cqblv0Ro6HJ9UFerp6ZL1jcJ9axup+nAqRrYHe0R7bXdMxLcZRhsfM9ADt55g1q7zrxo9/2vZAXb
8PlXLSLOaY+ilqGZhNWvxAee7yDt0oRWAcRkjMRVm/EkZw0t6bF9LWxj1eH+qJh0ZYkcNz82ZMQB
PMEO6s717zqJklxyQs+3lqX78vRj8UWTwVbOP3eGWA4Uk2FFDXsnxGNcEIWk1cjykB0Xq41+1LTS
5E593VLLLNF4nhPnBC3uvhPnbI9MDdM53pZRe92pIdtcTV1apKIlX9HT4v8tgRVZ0kuaQdp6/SzY
iEntrJwm38LZmB6PEsgwD0XeVJGcxZK6EbByzLqpF77dr2rbvqZHEc92SXrQsJVqa5NYkfT/f8tc
dd1iWayhZsjc2X5CFLpMeceQ/PEs76VoCI16pzucY5bxTt2FxmQGKaxZc32mHFFoQRoFoqrAzInv
frA+AO7FCHKKkr455KUs01T1ClhtRPp8UriT5JZCJrm42Airptz7hi4k2lE5LAifW3hT9+7f4+yo
vfCC7ChnLJo/ElzyGe2vGimUYBs6HrXNjdiAqyHTaeG1eIuNGhx9vUsgZ++P2dHzisdmDr/T3jw0
wklInqVlBOk9Z6ZMD3rUuqzM+HJaSlAx4CAed9FFaQConFFC80vYYvYc6D3zQngUc3QBijo/07f0
2vg2ftX5K6K5iT74ayb0Jf2CE85tBpTmE+qtaqz/ZVp4CpPvM5dfA9J/NOAF/ByxQZ79+o2ZUD1f
weGM6Ayf7s90XssYs8mUUkBCRLlCFsr4ZMM7t7eaeg2rn+l3aK1CrjqX9FzslT2Y/DAPdv/IEH7o
W7VPyVDRd5TcNTdxZCKmx2Ee/fopA2EVZIcvUi3n/NISeb1oC2RDuZy+8YpAqRxvL+MTDxuHDeaW
GF1zaCzgfDVg4AaRTqH28ZWpVIoaRLaPMv/5FDIh5dQN8lBJ6RACf/fJJYUACLN9OiHOn6R7VfjY
e7AiiD//NnSCdN6QFih8maXzwcENkvzrojSps8vPwkFrChkaRDMjS6Uom53Jq8GYvvu360HndFpp
4Z6EOvcud8h42rpFAF9FdCeoFbIzO15S5U8Ki4fGA7AzHi+qJYgfTpidGp2S9uo3th02LTqvd5RL
KT65y+CktWFFqFSbZBFGaNue0S6pzKV7Winx/raqQ7Xzz6bm0Tpc8qgJ47DWmfeuAWnh3BkoQrFj
4+NPdjZoAJg1oSWcnkTHW+WfZpSkgmbluXgOKBjXvhTWqZrfLFh8Ck88yEZrc7XaJGN4Vc40CcC/
ygCfSstbvxC4lHzohQLoZibrnP+RL7XBCPK30VphVaQ6JfBOjDuq34sYTMrH713aAUFHKBULx0rI
OAzIV3WVmoQrNbMSszL/rrXpsmsuytmo0iIBdbqHOBIvP0fj9b6Q0haux4rIRRBStX73fBPFMf2W
wDuoLS2xoUm0lr97fzGvc92zxKtWS3TpEg7fCitDB1R66RPnKTTxFPDWdLtrA5H2Wdat9W+XIHaW
ThUyCwMf3e437OBlRWjKGtn+btPnaZkvBx0JMjfvJnBp8b33ZY3DT/V0yoAfm/ui9eTCH5J9b+Be
NjJxKeYnC4+R284Jhs08n1CVQ7YF/IozwExhHyL5SSZpO/QA0ENWld0+ZPteFVjdlChgjcmIsWzn
aCyPMIO7GsB1tnNzb1FMkcy6yYQqLbgd9WpM2lSkEl/fiMwqet14hxN3CKI74ExGptXwqQOASw19
dkok3d01qkS9neooZbhfgFUZCAYyaKuNHbiy3gx+YwGp+/PHePKOEjP5BxxBAyonCiMel+Uh3M7L
ZBfXaoiv0beciegDd25/rfOXZFLF94um2mDY1CQuXPlEPGdyGOFzvC+X5hzNayZ9aoDWV6MTRCZv
UZyX9PwIKUs7m3lP7JrrnNDmhbp/N+hfTqe0saET8rITddIsFNImuq6kiKvqJ/jI/D60PoOkIN1m
KnnQKp7qzK2x0LdEUgbZs4cnGPcjmU+qGfUY6+h1ptWrQISFKvp+iHmb5YmFEAge4XrIuVtHTewU
PQMSWQjsVul2z4pXEKcrWjdgEtyiflEarDSCl0AqrSrSa1+kN4Qw56j1ZsX3+N0yECP4eETVbgBe
HlANd8WixPeLK+OSyFrqS2R9Ufyoyre+nUIAYSio3cC614v6pgCflLIosx9yTda/TzK7S7NIxkUH
IHa4kntrZGQmMZ4TUwsifLQOWjSnivb5FP7TgN38cYJe7IVfDyTefvkKjJ0UH1Etqf0lv9zhPixy
6njwtjEJ9Ryey+sZYmJ55vMA+VnheM6g1n1GU6Wv5oKPvvNbFGlTjLO5yDcOYrjiiF4Dekr3nzXD
VkgBBpPCFCn+Rh+uSvYPGLVj5JexrH7eyQFTqHhdS9n87K6VIb4dMxCpr6irywpzjbtpA1t8MWea
Ym9Xc7Xo5bnqfROHYiqbNgOpJY2Qf0GmFeNbzGtw8X8eIXGlS+8uFOZlge0xXSZe7VlzNRljHVo4
wb+J+Wt6UNziba4mH2jVdrX49snUEb11xzB27ygaI+tFfjYYTFs+5Iyul29hck0nRz1tUa9exxKJ
/7w35UGfD3WXtZw/m88ONUXi+MJp3EuUBC6V/QcBXAOaYWcFZbPJ7ToFbkUCORsLPmm3t3JW0a9v
/GwC6B1mqAdNwO6XvoVr1gGzmG6nF8upIVsVF1TIihtOgLamKoWiogp4FxIWOlnMfHvIGjgz1d4x
PAe/BibGSEky4On6mjuUCYBio1M/xQ/gLUFgNnlKM75NKxr5SA56CsWO/O4tpernVIRwsCxm8yoX
yLfhXmCNkMlJimhWci3xYknRFpWXmW0adJoSIQCqPZRQ0kIRpI08+oTj+Xp4bh6O/0txTQDGFSOH
EMURgXpvFJD79Wq/iwIVkuQ28Kge7gNUZKUOnMQwECsn9WFC6B1aYv0NtC36f2qRhRHsK8R0pjnV
uVdpJqMQMWqDqQ+MVCICsvD8ImrPyhmchwk40l6qm9bJp+V9Ohf+IiM+FKAjGS+Iwt5PRFUMH29j
MnV3tgfS6i9eH4uTyGt0vitHBGJ0GLUVttB6QiDG8U1Aj9Fzf7VA/C31hpBcwPwMh3fbh22nfomY
YMvIJVERmn4dBtjCxAiXKqzNMgEIxZ1EseayIcQ4nodPsLiJhGyu7ruFemqkDWgIvLqMDx8Pdb8M
T0o3Z9if9c20truk6pjd/K5Li/Py6n18/5DmfoieWE9q8qEGQaZnJaSDpJ249vCc/j2FrCu6QdEl
RqnJ0kpeGSdPjxBooY7oUwtwlN4/hK1wLMqNJW4DXW7lzk75iUTdLP+lNgsqLfovEKlLnba9LEv0
dmHvWmRYx9vjoIHn2zeuj/EBviTgllrvRW8hEY7vFbbpEcb/8A05cpDJ8yn+og1UyUfM04dQernX
tIhAQSSJUJkDhOApVw+etNCmjEXABTC9wiB10VhUDYdmaqoYAyv0ZVjfKKH0T6dxRX2Jn5SDDX9o
FoHLARZcrn/MzfyUuY4pHf1DGSp5rEAWHfBmcpKibdfuwF/haIhOuz4i9yWI3OrTrfDQucNbIoW3
HObZ/ZXmGvv1s8gkAusy9EeBtxibq0izb1d5Kx5XuLDCBj2jtjy+TwFYjmtHUloun+Kb21DxduGc
wU6LaBCrtppi8P62YVT8mKguD1IdiBuUTIzkpf8fy8+jyUACZxKoRORNSAMDB3ddg/iD2b5eAK29
UxHjGqF7aim+k5V7NKRMzNJYL2e7YLPeiOiT6v3ZTOh4TG/av3O7IawCdv99mylOwajMCHNqbEGV
ORgIhq8hVuiTsmjpAFJjfFfV7cBMxiNiU78224HXA/KAaiHYs7dAaXqO/hgLTiTPHoLzfYpw4+NB
hIRJV1Ed8c0BEy0S4xqJb1XAnlAVU6QXSmgLCSxCBpxw9vySRK5h3/6gVmMADBvobKzZQjAPpVJp
Ur+VG0FbFai12NU0OTu6Pob6KsZjrtcBi4ZRw8fcUlyHWTK9r16S1bk3u70Z164xk9n2YkGk0UlS
NuBagSmg7yYQNzNWJiOMuQ6BJf7e6ZNz6NcGnNrNLphF4Xjul9R1X349if20qodHKI5MhlxTxjG4
19nSr0Yv2el/LvZOTj3EDAP4NUxnMLAocGhCTdAWpiAQ7/+l/Wsu21AY/xpOYRKHW60dZXB+rI+S
sTlwavaF/2VC5GSxmo3wqqePytEdqNV6zgULhTX5QO/ZwtgDtBTdXo1NCcwoyL7aa0HmewDDvQ7r
C+l8qxrk2t+NDBcaRjQ2oscNCHblK3RpJ7xKoQvfZ9JRkWLsQQkt5flDVS9MOiTWZJiAKGSAABLT
zE3Sy/whHIArGX0zJ/hCYwvHtnDt6sskUvEru42lDt8x2pqtzfbeAA6Nj6Od/J+s6hJZA4C3cDfu
Ch0emNVYtYn2E1S8Dzjf3mL/bpEGreHVIhR49/rJ2JVuAk+WMgKLlh58Z5tvVhhRgbfETjtZezU+
zyg963VI15q3kZfh/ldaxb0AcieZPHWrh6RFeFeGFB00Eg8+hsJCjQMG1m17EjnZFldo1/BxdF65
oZnyT187dtBIf94OpuBNHlt+jXvxZJilo0rGtIfB9QlGS3WRIhUTquHYCbO/BIwrhGJ1jS65kQsU
AhyA0M/CytrPB/YeI9iahkCRW8lzDll0G6r3x/vI7ZKGW3/TpCHRTeH1KEurdPqk2dixkrPPKyQh
znp9AnG+H460sVGGTiGA4wDbFF/EcpjJs7asn+fYvD7hjbP+TZaUfyk5TFMreVzNpSW5F9gInvdK
29+OegE2y8YGI+om2OOMuKMMcNrbT67MyB+mBjOj9DTyGasF32X/NRJ2SY88soh9PV5DyC1G2G3f
wPCwG3AuWOyfCpIKg0WdCD8KfU1X0gmvbdJZn1cxCNhTTThnEOZboTSMxPVXwscdS4ieenhM86ir
hrPFiKssru/J9TjVChTlLqNLD+S2/sL8V74aElr/aj3xmY+pLm73QY1VRUee/ZSsuL9WvKfn6V2f
hQS2Z9kuFceDlbHduIhneIFstU5d62Zd0VsCr9NigTXY1OXXIPucG1zsb9RCaZEWegUEOtQ8p7A5
7H5eroFL2JfnBEWELIFH/eK63yTuCZIcWwtfSIi3UI1ECvkAXPUFXR1+AGOVTb5nTYWWMtQHIhlg
yxh+2ZZz927t/UWy9QXYn8ZGgDc8TskLpYGXQsCISy/RrhNvduBG/Li5WCLQiLH62ZnyMwyI8cnc
jLOoWc77jmdjszaiaCFxbvhZWJBxeuoQn5mb5xNsR/7v7m/Rnh6Y1eFkqXSmtWvwF1ucRosFJdaT
CmIMUbx9sf/MFfEwNdgL0IX2UZ2G+fQIN8FE5HCOMPe1+3DJp4QopamYuVERd+KXxuDvcpiTYbS6
KuhS7NXjKTzkWGxJ6moFC/X3gKw2brEz2tsXWP79I+Foe23OXFg98n6BdgFCO52dLhOMyMvo+QPa
8BMuzK5HhGjv3SbjpzQ00obCiklbksCTmNpSl8l77LeCULlZX162CuBV+MtngBYHiOmjscUT0DsP
UW9Iu1vB6/R8aWG3+Jzdx8BLO4TVXiGPrQDBa3YRkIEWC/IWTy8teaRe6eUD3bq47RuDURyyof0G
KiAAgjES5Tlic9bT94YpKdS1MGiZKylxMCmGxhMtWdp8zveC2PK5vahrtZqsTR1XHme7YgnblhNN
ObIqz1pS4DmlMUGQ8XbPBwIa06ngSQ6HPlvkkOKTJl2VdXCQZvnJTiP732ykmd2e1F8cGgfXr+fT
5xNBSejnQvefYx2PuKsaoyueJDgUA1fmnsIUKpLj1V1l3mFtny1pKPkRJ9JlZbAWnB/rnS25TI6N
CtNtqmP9Z1V9WC0IY97z+6ylKdrZFOhlYz0fHV2yGXGTQTB1D+j5xViHDtJOyiw04CgGP6UTeNUB
9lC5AlaorGHAPo+6PJh4+92uSQU8NGPrklT+kV2Hmv9ob853DG8bEiL/ZE3W8uixTTlc1O15p/Au
HL/Ci6T4ir8TScXxsGzxJX2/l3jXwGspkhoevr3RzrF0uk11bIZgJ2y7mP1XFgn9vYFs5coay/1D
WFcodzNi3Z2HQ2YcL4PnfmKWJD4IRgjZjmjA1cIEtF6xbMskWkuH52wWvucHN/JwkLYi7NqEklEv
vN5QjAVyJ4R35vc5b0MMUkegN415zuccwY6s6d20GsvV9LM7jMtAmHe4tQ0d4C2+RxPM1SsiWATa
ODeQt+L8tuaIzfVYISkRCEA0G3Abe0L5gJlgsPpDQQh/ysW35+BUwqMSdK+Z2/D2MVJlYbCL5cjY
ODIdfN46N+ydLRPu6sIW6GW9pVDBPC+C3Zl7dcTRiz9IEm/QjPdDafvNiF2Wwf1L+L7qD5ZXGvv2
LRviu4k3JVz0aPl9wjAXrlk1Jt9+Vyt2jgLQ60zv9gyvlLRnkTX4R7jV/ZPmB5LdryYD17fOL55r
XiKM8aLyo8IywBxp4gNJ7T7DtevZHX4wgzSM8U5F7Ys1hCZAKQhbpnY5Bp2KAv2msxUDYJ8RwiHD
U5NuYiSgTaNimrSTWBMOCfQjGrPMB6piRdSoT7Dk+kFopK8CsYxu17i9NwR9WsnXnSOyoLVOyN8+
jKpWUEZhyU1b7eIoa4ZToGOX0ISFwmxKCJ9DcrSLyudvHq6SbUm0abH9kWgIBGXeTEv5qwhD6Kyg
Dy0625fwiYePQehJXx+w2xYJeQ2GgHO2R0gY1ffRD3+Nk0dm/q5/sAHNsgGWhWaR/cYLl+WjmkGO
UzkRh6KqR/HXiLkT186zF5yj+X0ZBpjRFn7T3JXfOQCmWX/3t9koOcUoT4Wc8xA8vLIQ2q1h6LXW
fwIDKLP+O4E5J/Od3KyC+WBFOXwYU56cFUXa7QI7JuUZbNBZysg8t+or9lBvP6vc3nAxoJDeJyKL
iP90trO2yjBBpX2GkLnv/NHo9qCEdfpvDYtaWK7ALFgZjWfkTzmZ7bOlrcKhwmJTDlZztIPWXnNo
ZvGEAMl9M5BqxP4Vj7FD05gMHPpNyKbGm6JUXosN3VyQ3ZBKyjEDvwOkAHYDvpNBATDE/WaEGD0k
eyFBF1LZGARMFY6GixSD7a6gG2Ra2WMFBpIecyDLsT/QPyRgpujNgQOICGYJa92NH2FT+o0r2yKB
iK8fYSZDo7EnM7O9NIB8FkPbhMtoqkVPI6RfDcfOkc42A/Intn08u34PzofXgRHeyg6yBpFo+Dny
g4q68oOaup0MS8NL++N05JzGCOt36b1upMaQ9t8ViK2/zSiCLrKuKp/5jLtsHuodrg//sXFlxpiA
1v8UJ8ER5PGv3fCRuna3RizkK4NJVylpoe3EFlYVP+kOg3CUdAwT1Hqgdt5UkyfpN/p4yBKDjqzH
oP/pOGOJpvCEwxysJMowGz9minqf5GPxy40Fmf69vT+v/6dIRunLKEQ231RVpRqu+K/cCenK5wYK
MMMPRVpVlgOwVcaYlG51NI2alQOqhVrvKc6bRShynFfVd/JTOiX5x35iEmPeHC3u7Lxg0naa0gOb
RZQFjUqUXpc02ZXCK+jfbEb5bH8MEzYkNmlJm9EH8qlR8lkUqKgr2oYvaMW58QiSufOL5f9odXxD
OLYwqTZN3xGm8OGAz6X4dNMt0DrBPRsy56ipfbqu6/68eAY48EKRiFjODWiBWF//Qalvg46jOhy8
IT9bI1HyLSGaXg5rW5z4VBhxFEsSmjDbyFqJZpiFUNnOAD85dX0zes+OlkZKaRblke4kObqFuouM
qPqAi69MVL9czrwFEHxM5oJXYv/SMCsQ6p2vF5s+ScapmmKiOs82EjNAtmdTZmg3YzSL+o8+F0AV
1D/UUzuFrIK9QL7+BUFZEwL9YRjFTFuutz2A1MEG5G6DxubzAppoGzr780SpU09klDgMOxbulmLn
SsgGLxHuI4LNn/+5oHctNHHJ0xOx7pLxfED86ROJBGnEO70DPb4UXg+fvUhPAfw3k2y2g9dMb4Tg
kE9/PjSSZI0jo9SxCSwovYFSvjAa0Cu7HaEoWnotyVDvwJ2t/ygHMv6aWuuqqBQQTFCr99x1os5x
F09EaV88BPhLd5nDUSkoD2tbnYhCm5Fk4Q9f9RGIpP2obdAnaksdTni/GVJxKRxhUe4z5YVfXUTQ
IBIiBXbIOpPraKQfJyd8jA20akbFr40YCB18mA90CdRkW5QQaqGb7RazsMPWwA1uoNs8ACpIRAJ1
ZFCFUZp/kH6wvaiAzeGWhBiSocwj0FUQlLGdcCxAzknPVg/5RTpF2ov+im58bOIHxtYLz1dR16o2
qwN2n21SUpdopjSQ2bxcPO6OPj3D+LVG8jUUQmwwUIqoTCZtVH+43KAnDM5SNY9ClRQgj0DXTGlH
wMcscju09v0HC5PbUgfDPEz23TiiTUOJZ7hkE5x41DoOjaJQI4CBM5k8b4y9NDUuKoz5kPGECdY/
bcU/cOZc1woqjS8Q7QCoY8xGChXNZTDemIYWtPoWsWK5i0298LVkpLeX649lnmi/I75dVmdGBb/X
XiYfhe22xc3RJIYoC1+C4gX/r0rVsLF3VwymYy/CAJkKPXJSw1pYuhOoLjmkCqCTb9zcxdqqmxAW
Cxou6E5PT5ip4XBPgJuvY5iILAQU89wwQFoR0AVHE6yfah80bUN0PWV15ylgjHOqHizNIqsXnG9M
798hmAs3JzIkWVyOfmmYyQ2IuYu40l6iAzUqT4ylRysyV/yyMzYIsqNZts6ZqjoecuMqhrlJ9DU8
ttMXNe247abVJz8hfsEoeq8Uaq+dkHXVeR8YkHntOpgYf/ftykGfAFxjZV7YbiYY+a4WusT2MVum
LY1ArgvbR5+tWtT5YqUpYVlD9PuVxbnQ8Mmlw97uHcUTElBn/bKGO3gUldAqAKXNBJmgOu0UBgbB
cfUn9omanTJyd9GIGpYfEsU8nEkaRCjU+hX0ufVRxfLG4t0Vn9/hkNXziF/xo7X3oKXBhUufAPz1
HRo8zkYivPlQF0K9fhMhOLbA/pnYnaH1j9Y1mk/WGNRXD5iiX273WwKC+2EJmgfFLRzYQUkJGh6o
Cvt6FpL+7FW1mPC3FmEqdbEE2MFUY4Q6nOJWHs0BkNXjluGMbhu4xTZsZVE/d5HxtvyY1ZQphP5y
98y3VTLcX/cUxUWjpKsWhkShvHuMUQGdrzwubDp2yfG8xSodn0JMNcT4OH3A9sV8teBI80OgZsTC
x8bqrmCxB+mrPAqTIHydfyixMeahYB/pswEw8aoAmFFY0K/HTr0vAKM0Bq6CnSE24oTDYzlOkUAj
3MgKKHYkIoXAaj2v0g7GNfWz5YnosTkabW4tP3PCJtYYKgJoxK7bqDC9FELoGY5uAOf+pqMAy+sV
u9WNvroH8i1H4rvyz2si91S5iwuLKWXIzZ4qYB2UiH1M6kxlNSvxgO740Fzs4/gIeCMw3Im+53Ma
EDteXD8sDThkEF2StRHAq2b/e2Gc8WRqVucm0NFBPJkQEqcHZCvk0Su1Q+6rViwM/Hr1Stzi75+z
ISxpQrSGai3ZX5E3UOxp4/6GjboOL5NWs3JDSPgVmlJVXqs/CiHFxECee4lVf2CyDthrw0Qzm4Kr
NC4fabYA3ZSdjZHjHXjrTQKR1JxlwV2vssWndm4foXvMsylAL8w564TG8gqIJx0WSTTyN/T/9UWN
89Fo9phM1l6CEIZk5Ajsv4x4n5dPsxpCSa2IwX3UB+bIpEHwuxBKN7bIr2wgy+ru55MKn9vezAYF
3wMgaAE3kk86fvKTyi8olsrxqR5hOTgj//HWGcJt+mnojixpnnVfFFQ0QLm1TxBNeEx3hrcXs+S6
cbrIGDEIbS2kSlq6Y/gnD9su7OOtCRjn3zuOSkTprAb9oM3wajH2CQ5yVdqRB6LhjKrUMN+tVbPP
XjKIV1Vu7ItCVcBfIpdazdegus8LWAz9WZkazqO8oKaoIoUigcG5LHN943qKU0nPSphmJ+UpiE0Z
FBZ8AnWKRG/ByChv0j6gFVohvfEAXCET4xiS4ZgvnRzPIkC/oSGUf3jcgUTaOZxb8xKCLZhEWbNS
6qI4ZVtB/YEa98+FpGuPYWbRGpJgps+v6gbMyGMCeNExkG01XXhNN6Cjih3HDeQx9d6NOW1dyEb2
z5PUxtCyaYRLsIZiRsVEcyZ3H6Dub8NFZ3xQQtpGBNVxE0uEU2CsawVmKzEwE3QUyb4TEKJ+0y8P
9yrNS5h5I/iVyqw0yoapc0LIUgf9KADszVdAncdd5VhayYO3ulmMVAYLUnt8ouKSrffdU/B/C8JD
J+kqRLnbf3mCN+1PnPxYZIAichwtXLm0iiDsay3pJMz1qLHNvqagie7plNQ1uI5Wg43NUhzbcWYl
WLh3bz7KXWqmhD2kMmOTmRVqCMrBG7pVzvAQnnXY+BUXeSDxJbMfYdfuMM8RH516NpwwWKB6TSNz
JfB7QWXFZQXfw/D+t0f7Di1BanSGwAmoIDg37FWkV7l3vs2ZFURPvJIqjHBLDef0vIMmJnsQ23rj
IrQywMs1TLhW4d9rbvYcECAkhgG0JnoI1tgLe8VSXrPFYwwk3eTU5e90ReANIgALmvtU+5htZIae
kixqUs/D9+eBKZrTpnEdxNtWEYOYmpqTygBSbP8fE3YChs1K5eLDaibWTJI6w/y4p6qOqKRWPcB9
rrVlG5iv0cD5oEIU5iJckY1h/G04C2efuJlmCShOLkWRS+IbdlPRs85AEcxfWX+f9w+sR96ddWA2
79Vyu1/BS5bxAwZwHi9FB+ai/Uvdg99kvehFZs4GYvFCu3Yv7f5TsHgec9dFOuHw3FZ8rd5X3rNR
FJCS6qIBUYjI1V63jH/bNnZn+1ne5JHOQE529e2ZkAkXUEFMLeaSvMVVXaMcr6jRETYjvc4+dK82
r0ILf1FSIrGPNA8mj5Rtz1X6SHa2pYCT3PLiZXDtJyb3wa4Qn+QPTD9nvQvJeE1Ae5/1EwZ5Hmg7
MjZItGuc/kgJ90BIZGoQJ96UqyqxmHQzMfFjs0vobdqT5U52foPWFDGtk4Fim9N/FoXQLFlr82u5
Pwc+fSD2qIYIo+6LmxITayFGFPtTshGptgog+YHs00nLvmCvwIeUI/86U5pJTcAmsvgVCj4Uz+Ta
zkESR5dsrIVCYe81t9Ij02DjwDTkQz0MLmxfG42PztmZYqMj2lnWfb9Ir8Mgi8nHuPARGUZSJ4RR
mPpgn+BRepAXeW4kI7I7RQa/44by4/j/JWQgCixu5PZzxPPLhYHk7ZM2kz8U+ys2lWMRUmVwcZqE
0m/XXDbnxEiiqxaG/Yf82Qwjv4PZGyUk6aH6jR0P4VihR6snDaCD//hkA3zBv9Ei4WaOJbRo50Nd
slM7W9+E17DAM1vy/N+lCM0AyNVDwOFvQwP5JpBTEMi0WfoaJ0njLWKeWTipq5WB49nVbQfg86N2
cWfdlv7KxhucG0jqHOZKpAUFBYeSTX5sE/NM9w87R8Aet4pv8cckTnRHZlTTK6gWskSl/c4tWN1q
KEFdUuEuK3v+gL01eX2Z8x66w/7LhGlzK/YlMYVf1FCTGxzzypy3l6ESEqkml6FyxXMaOcSogkIK
nObWD9/Ad8e6EI/nfFH1fz1fVkQkxnxXIUTEApfITEfK1mDhVLYrDMqKxhSrg3+KvsYAqLGBckFW
caBSzTGnd9VnkqVdMyqwzwtVB+s1URvHUBKDUInMmgpz3RNCtXKxQSVFtJ1GBp4USiXN7t6FxmeT
9kwcsx9h8bHWwylyp9bqwlROb3GsvqyFfM/HMhwGY53kklWbxKbztRnUQINUiwUPU9ILPn/6tljL
MtIIp6Cto0XLAS1p6tVn9czGv3Up9Yz0cuj5xm9xKGA5I6ESwdtnPKsGHuh/uyh4fwKAnPMT+8SJ
iq3ZXspIlqL/tz5FKfXzhOMBL+plcFhJgZg/pzNPv0YGC68dG7vljeE1qaIaOSgjNAu57THOmSXi
u6EpbV1am7uBmVTTlA8Mge20T1nyg8cGBZcXxyCS4pWdiQXKAZisHammC6QDw8cwfgTDumtzVskI
OZ3cvowPEai6QncSplVp7kOKRh8/yu2ektN02p7/Y21AsRF2A5B/bieZX/tb+JvslZY3xIuRU3tD
C4+IBnwCysON5UbLGTih1BYBbF9AZRr2x5wcZymwRJw/venuodzrZmKaZj0WUNOj3hVkxUAPDPXJ
7CjeyF8sXQwFGYycnlxWHCTrcAaBBnmuj8rLNXVy1f4ZK0tPCoDI5PdVJsvulO2vOgmcDuyt6WLK
gldg2u661apQaFh5EDQYalnv9rNE6V8kE0ZQjnFaFc56eKyh/QJpp3af46EcHxZMDiK0k/ezI3oe
OBH4EuggI/Mn1SQvORwpT1xKXt0RKg8CDnz1MIkinF5kGVORKcgA8tgJIOd6dk4bFeP9EwpqAvuI
eXYxM1x+5uEeAb1jaeY1NOTXxWNuIBOtDkcJVximGOUtQt1CnQTJfg2FtI/JjYGIP4dl/PRmRUW1
ULZ9zncco+IaV3k+VME2sM/nhm4qZYc5dnYMVYe2pWs7ZVoV40SscGPXRqcuUMIb/DAKbaVuqWAz
jUD/21aLhClsM7qn0QSCk4gYqNzrlG/xVe2ya12BCvqfqjUkjBWNVj0UDcOlJVkUasJrf+5cMOgy
dWihSgV04mt89hJyZD3Y2zqwb/2EpWc7CTmb9j3U/u0VTAqAUtscbnNC3TO4rmcXWPz51i/DLdHn
UBIGOioZr1BcyUZLhZkO3khKURyqpDXcbexMbEeO9XyL5YIbmRbyHHKfHBQjhDc7Wez1CTxN/QYF
lQq0o5bupvZFcPdcQ4Kk7e7o0Cybv20tR8O7yiWf0yj9PnbOaXufNFXm9WDPWKtRLE6xQ08A13lT
YeQFdv+PVFGBro/ohbOvngvikTufGWTPXoWxQ1kCISfSOJNim/HHUDIzZwhsWwJ0JTi5ENxNWW7M
4A2e3LqzFqjvD1r7ueVZ7G3bOXT8HFOxrCck/WSk9+WUh/dIAzRjvHnL5G7zMGpCGeczw7xshePp
Ujm0MpmRHN/MQM7ggEcOqz9t6Q7aOJlRzQ2iF5SdoJvxZlOO74LcFbSrPpR/vSjXwUs7cExoAibl
1s0mKVPJE0HZ1KuDv23lSFTrF+DvT5eERhzg1cw7gNR6KN4Rowm+8rio15dlhtu2C8/bQ4lEDBLS
aJP9AB8pI+NzD7hNJlFma5gfXTSOWgbCVxQ3CG56hNqNic6bfOGYu4bKahsMg0MIteILGCKZRJ5A
X9M8gg4DPnHExD9TVsQVd90rGBuu6YyigMz6bZ2y0IwKY7k2moxX5i9HQ3kBzLyomxu4Vof/ZO7U
aEr5RNQdIT1sgoEEvhPahk2dJjnMeFsp3U3xj0ApLD26LGBUZmaQHGlON6qfRoMW5n/BGCR62TKP
hPT2M9QboeIOvnnSRgjOm9Hv3mJN2BrgtpbgPBXOV2TbI9Fdk2+KPiCjg8EhjK4r37l60j+OSj3W
6gCY/F5Pbfzz89fgJssUCb6cBLxeWpZ+hJr7Bd9SBTU6T55+74cpw/9FZx4tbUMQOssWOa5xXRvt
SmhprJWGM/jLcQTjh1yScxtkJOseyyxJqUJMiE6fjl5oDH4p44t78rA2K5ACm6l4HBnD1dRux581
9L/zYqLrMOcmOI6/sFtp5LueXcOsudTDyKfFDe1P7weFTT+GXijn8wEagKtcfPuuQyv2CvGaXUof
L8NtpYhexyAV22+qd7EPNd2wAAVKkN0bk9gWgncjCuTA0Qp5lyMISxhvrkbK2FHEWYZf7QxKl4FI
wAmMnzwRKfQcJluwwYzol9AujmfyZy0F0Vbykr9E0GHux4DXY33NrgZPGIX2ipHJkyPfu9i5wIeq
JBR3CkqXbYHwLr8mya4WFIvcbBMEMMC6Zx2c+u4HHl4zRh5g6U5SNSLyPuz3BC2B6l6mHVwzURCW
Aq4Ljrp/4i98F9Pnkikc72o0yYiiif82SFY9YF3sIE2OUt9s45UN3syarf5oA1KcSaU1CkwNZhmp
XFmjlRlGe6SSQ6OMxtaN8CcF1vV64e/SprW/Ia1NN+pFPO2m9cuftoLKMuW1LWl5YhbZcb8VXEOk
kkftBd5M4P66H6s0wj92bTNqUNoxB3pP2WBN+1bM7yq1F1ATiwlEg4BV9k9nWMZMtwPEdhNMUdsX
awStsLlZJYDlQkTmh3NPIicJiU+56iGtWUHVL3D21CWFUbzRRI6ZzIq8oQ0GTBWJLGLmOqizdkdg
sxh1G5ooQmwm7UIbEiCEqeNjwzUjxsM1r86g4/ineqXhYgls7+LWAkyujj24/qAv0Si5COhn633u
o1nMVQvtB3bCel5KKtWPzKsF4cr2bTh3ORyGh7of1gpvWSpTbnwVIse2anMJNjaIZ7XGKawoKuYO
BW+L7t0vrkRKrl81wy3kFzrbdWFZ1n1WKZgya+fRdFqUY0jPCAiz45VWlGRgMlkGyKusU/Mc+gvK
1Mm8KDbihu6Y5SAd4xwU2s0FguuQPUBzV6Mo37jY+9tie8SKkCA92l1hocIy78SPDpg1EIvhFzDJ
lWX87HgG2YhhksROlwp/HJr8u2+Gah/Umac6po/JReN4c2G3B9fFk6oDWz6GntUqeSNls1lmpub0
biEGfSdoLzr7YMLYCuYiiumDRx792AUuKfii7KwR3JGuxsnBWQcNE7d3YC15xPeRDukW7GL0Ihqh
bN/q6sltINMmd+Ari17SW5CLzfuu0nREnwyz8S57gxKs1VYaro+bxwCtGjMByQtxL2VNBZWPjm9d
zvcilnnWLBk4n1d4dkAKhYF6O0OyEKvC2dQGy61ksTcokudv1xkHzqVCDX6hfjM9IU3Ozmri9bHV
AYZ3R7LV3BmWN3PtTsHuCGSZEYU5GK6EJzBkolFXF+J2tB6lqFdGC1+otMH/qnA6iV0UpajE/TDp
UZGMNlYVhI+21riKhSEehIYnaaVDvbxsLUESvZQ4zNRVg3EZ1Jv6Qfyrz2J6Mv9EfABefoEFKh2E
m3LMh0XD7pvxExWGG4HB1WiP+l5uZWDPJ24MVjS3WNfgL6b1GzhnmNHW8UlOWFzYQZH9L7PG6GNA
AIkZg/UAJEJqrEwb2kKtSG0QRXa+9lpdvEUMYYdr5y1aKbvVAlDhnPr/gDp9cGzRZ5CmRSrN1tYG
TKzF4iLtRVZDpqG+7ebxuwki0zC4x6R4E049iXEomSRMROslr5gc/zQnXaqjZTnXrSkwt44LZvO1
EoEWJile3iFqmU1rwq46SXv7InycE8xJvTmGzQmM6TRDrbv/H9CvEiDQ8634Rwi4b0xG8QLVsI/o
xf3mkY9mCqdL6F72iRF0dcPv6H03lGekcwAoVHLOi9boRHqLW1NJZmm07Ij+9K4soXALQsfHSVON
zSUVFedtdub2k6V8nf82WMVQRQSCjyISZ//Ewasfx0qxvFdeEog4ayRLJ92MgkySrWPLEvEAgJIB
5TCHlV6lAlj+7dfRX2StoF1ezwfwpH40w6o9oLayZnisQR7UevGICUDrykAkkBEKlSg8Da8Av0SJ
67KpimefcNM7aYCwlQUlRHoqWC0Q2a+gFQU9A/+zfu+oSZ9LeD5VoPQXgQ11mMAWWr4CvON6O4Z+
QqTt/uLvPzfbIhdK71/CNrsC5BoDnvW+VcM+Ylyy0KuhDaXTiUwMt7MQWL3k+SCeNTfVgKfPpiV4
KCqcKqnLksXKgOunS3owRNYPVuJ2EG1k+AT8h9FDxuRf7/XZfotncM8PVVnNjAC6nNxRvSLgdsFi
iek3tP0eGeSArlqmLbDeohWgycsgAuQjot3JX2XakEBoJb+AqO9B8ywpZRvdBFHg7iPmvgaCPUyt
3sIut5UVbYdAFU5GPyuBRtQuYOlJOj40Y/YFAdtlm6b8AaeiXPcxcAqoJ32Gj5eKa293TK/JFKag
+CteUsU+SWwIasxZMX4bKcPGVmu8v1FCBfPeaQhJ9IbUt6ioFnB0tcrZKWjSmgjXC6WmFOp6LoQV
Zn4G6aB50B7LsT1QnlrdidI41AnzT8EDLU8KrZxLa3rqvZsfuSXBUJXCrb5wiO4MkNXVTyAbfjyd
YqTX1c1PVc5/ilOuVqvCsZ0MOGbG2OIUPsP3D6STCmRcKMGMV1+cLoCt0DlFNbM45ojSmnzEvBSd
heUIQa5zXlXbTm+NQyU8nKAOOCnLLMUjzAjcCyLh16Qpi1YwhdEibztG/gQZqknBk7lhgeHN7QV8
I7xH2gPOaFcRbm8QNXq5NcTlD+rD4qO4LB+i5muloNfqblqjKnuNXHV1wtt1k327C1U0MF5ejcyJ
AngChZY7fivipdnEudzZj8nlcNxVQffPOSCpMuKmRoy2KOaJ99Y8yilhDBwM75FVhLVlCgFZcKnP
eC9GHhTSKEia6J1sQhIFyv/NyMPx3efBEUMQahjiO91rLgw+SMZ0RTZQTbZXEShlADMtDb0tSZ6g
/+/7rS3do/vA+VmT48IYEPD/YdgYAJ6UVf0g46FvOZf25ESgODaTsThfBckaDSmRULz5Ox9I66Re
kNIqi/06sbkwPihYgoSGKmGvNxcrECPTVFlkJDP6gd4UPzjGLe+AtOPeBrjxpANFu78HNsfNhVyK
24yjzrFgQG4I/QRjoeIZ6Dbe2qoyq8JUtzdGazHcPOWjiQUpH2lyP69uj8bAbTOMFaXg7FYBbu5j
i5BgN/o9pJWcg8SJmEHctY20bsp4gTGb5GbD7z5p9IXT1/UU7n0su7t62k9m/t6P4AfBbaniS+8k
xHSoHHL7kQKtaJv68iR9MhlFI3U1YQSMOnObY4ueuZahlapZrF/UNsEX04JiGXd7/tKVgrUBVULV
Bo241r2d2wZXeAEyXWWDp7u4y9WFJ3ieLvL9BdNR4W+/Yp7ibx6EXyOjLE+CHcENu2KifmwA8+Cm
5e03EmBYhrcjeUsDyVH6suGqL8Y5wcH4wTCva4Ev2bUYdG47ikFnyQoznOLIywhGr2PVmVEYCwBO
Nj51OlrAEbVWryMYI3gEzmgTnq7eZjeoLbkmx1TG0QsAt/bctC8wSSImSR11/+CSYQwx10Q1f3qm
muiqGfJ43wf/kEP1mUV/T567m6OEx4r6g4JhZ0XnVbOgo+gijMa+uy01ObCekjL/ozR5iZ/de1NC
bNleZ8LtMW5schsoJchYgj+alj/0zExJWuzGj6mKvVNLhdrahyTdsDgX4Y94lr0dScx5cNThiF9k
CBVbrT5RY2upLOG1YqJ5Y2y3D7uqJ+t/OYcAZNadrqNELnR7yQSHr4ZQ5nQOqPUd0M6L7XjBndR9
HW58v4YaDJNje7Dk1qdjHnC9tMt+qJdOP2qlWHKXgfE17QeuY/tETcUd8hEgfn0mVG/JaawQ6Jym
rk3bbfQODRikRb8vr0MHtIXTO6qivdRVu4DUkqSIsQgM1qtM87Lsz4fcIY3bk1JUA9TjWB0SJuqJ
k0ypWHMdk+mm7VSYvtpRgSOMJUEJvQyNV2q75BTP7h1gNlnocqntYGzgZ+UYycGbdZ3Pu8yyIe7Z
V6yg1rkrCM31a03ixGHLYLrkwqiTP+CtNCz1ttDo7Lcgut0YXXDZ9GLJkAOU8n+qpQX1dTzrark8
xTmyOwuOWJ5/AaN03Gl1utKOwBC4azD6id7bEGR8kF0hJXE7MVpnrARuBiE37NZlEEHAXLcNW9ur
V2AkMylT50HRH/jJ8PhW7wbq70TU8XfzeIF3kyNV80w2ECTtICQG8ERYKcdQTRVtLU5RfamAPJuM
gUJk2cCNQJCcXIk58nmGRaLWaYR/qHuTp1sv/Cn4QooS4elGQeL6e/aJsTcnDPysdTdBcNHjelOF
xsudmtu792iav4qcKYKr9pOJugH9biAY3lSIAJx7X0U4nmqnHPlhO3QUTP8WCAHVBi6H75sOPwrm
n6qAkvDEgi7ih70PCYqWk8LEGcLwvwJRcboSe2uCuQooWXe6cY/xH/v14T3XHlswXBepzbvshMfi
WBxPNyuucDSHG/h6Lerxx3JVCRLc6Z9//UJTuHw6xAondGFFOSDVRBOPjr3yL+R3oSSAeo5bC/VG
LwHktVlYUZkchsScZX4Sc0ju9Obeipd73ppl5YdqXVCOrnkjoPLy0EtFvKqXzHIi5WJHumqFzm/A
F5OiFkVoVgVrTE6oZMJdmGMXEFB5KAAwtsJFMB4G8jlYJWei9TXBvAJEDEGW2m/NQOpkEntZiOU8
BHuKgXHy9P9zH53KP4aIeEG6WQ6u9L5gbeQCR5766D+6SVMDUCNT/FOlW3kEBUSkxn2RhwXq4uYb
dTt0VYVBA0xXGLz93eHDnReoRofsR1q4s71dF997iqf+KsdvcEdbj/VZnRAzAEf5c8iwpy+T8xk8
YzE4uwejg8UE7sfX/sH4uhhh9VlDj9v20YhHTex7QsLsDnCVPccwmJ703YCGHwabV0q/Gwd2Q5Wj
Z6qCAn8yLDfFwMuzIZdC6eEL0GZlnwFu+83AJwKtTuhIRbtTM/ZqSkLXqIm718V3Z+Slvu9v9o89
jE5NNBK9mkCCAKRXzZ0RUgidi4g4mUvqiSl51tXl6DCl/dadHVtd5lX2b1JIEwafaJfXR4Duy/Nw
c/TWPQMu7ccULmplj6EnIAHy49O1dM1jzSt4nIoWub+x46rr1YZERtaJK8wq6UUcJDyvby+JN+uM
jzuIV+7an8kP65MQoUe5SU2B4MGqSioCvTJIgi1DHO8Zn1qSK5BUiQi6gqYy75wQBj7qn0vXyQ9B
jCX5zyvaIyRdLLeBkkElbnDrqI4SOR2+k9evorQZt+0HgDFJ9uRAmpUlwAFeYuBzEEwyduLQ8x7s
sAlhIDKG0Pbd7JJqOVkKW4i0+trOYRrJnfgzEuSSQWJ9/Jj624VwNupVRPMnd9Too4jVMAJP5a3/
3LzLNZmvphUa2VyNpOsAN+7fcg23EYhvhYGWq2kB8Wk23uoi24XHyTea2MS47BT9AL8TzHVqhIWc
/SOySb2DVczVp+ROeCi+ls8G2KWP7M2VnCo4P2twcfjSh4c+XcNSt7exIkD/g6TTfbEm9hbEkJfR
dVVxl3mGZTWYPqLkpBOo7puC4nNHaoobMsZdhontvN+WGwgm1W2Hc8bsZlRTYR8dKuaUV1boD/qc
IWahStGdtJA9vM/2D/C+faIDCac/tXi+UAMkpsbVE5jyzefqcsesje6xMPfofarb4NtrNYG41/c4
RWJK5Q/NCu0DSQtwY3jzy08B63L+H+/pleXQPNIPw2f/QFbisZKkCWHdDI29DGVkjeFdvf12SR0P
zZ7UrprXSkTfzjyTZVNQzd67UYO1P2+nU/+rpcQmHWI6AUjLCYddHQd8Zck4ciE9it5zV27dJUDa
Sb3qYYePi3SBzEK+M3Xo8SM9QXl0MpxPoUZcD6IBJ+Leyfw6nIBS9e5uQroS4DXsG1Dq7yYrEFWt
4Ggk/7fqIk1cvaxwW0SZ866ZvaH9Ke0m6cCIGtKzXDhaFCNQs4Zfz4V2hRAe5lNGYAzpf5RSx9s2
guGoBKUAJiHyQap6SS0W60m57k3cCBhRKnLgzSejV84GmRKUApCHh9Lj/xrpaoUyybhn4x6/umvq
spODHAvLidHAZBEaDDZOX9yewk8tDzr7aVWuIhcE/tCwDkhMawGnI85wRWx2FvdW2C+bWWwfuRw0
3RgcYpzv5gjGeTbt1XRj1W97cZKY4vxjgoL2+NqlnT1ZBRPbSZK6kwW2n5JXuH44OESRhXqNgodp
fjHPprQ8/P2OaE+zuNNDIAAg0h0xGQe2KJdqdaLf2Dacw8jZW99zP5UhtN3mwzkaWf+6GiDFBAgc
X6zwdrtlAB2Os+G618fT/anyPSe6nInRyN+dl1mj5rXXYMzvMkb0M6lhuNzdO6C4kok/DgU/jDyP
ekf83vJIxlzr+7oGbnlF02qQNnLRJ01gfyZCOLtp69SpZyy7CNgK2O1DSxrwNfxdlSLLK/Dv2TSv
jEEQVOaLmBQf4J1LGbsdjPOvHN672aVpNsbrYZdbFlfZj4rT9DjAJnc/+9RLAcIwjQfOWkHR7s/u
Y2/OsZnbK7RWyGRLmidwoHXhatZv1846qnVY8TMCBXy7baYujXC/9Nmfas/YNVHvjGHGdcl9ItJs
/OD7UQerL+hXjB5a5AfnOXjqhbvi3wjF6edIvBk5mImz+77tTmqMyWOfu4SRSyqO1jsM/0c+h+BQ
+bbpqiZqVB9qmHM+xhd8GVchnwjTqg1bRAQZULf/sQV6AyontTnQY6Ze7lL18IyLHv07CiUuo9V1
+0NI+4X/+b9G85mS7e+4C5ZxACUM95zzIEfG/muedUVJfQQJKz2EAEMX2JGtxXR+6Wg5U6fxYMdt
grLmmsJxTrJTnoZ5pxKSVEClqpmSRlPKpDkwzQk9Oe4BmmVvHOKg2oOVyBHnWkwbTk+mS5eZC92H
YauhV5iVVRPV5cgm+74i6wm7d+7n05G22roHS0Trw8Lge6AmmIsVyUSV4ElHgkNc6r+DqkTYkLEz
5WHshMg2WQ3zVZIhN+vHhcXpoWZ50DLArznszIwR+57DeygsazQqKvBzAxoNGBBtUfJlZ6QDUInd
1+6xsquUashVvf8bYmDj++rQX0UCdSsiIgLF2ROVMXyTEm34/8mBtLwTv8P7CK/mWJW4ZsfMu+3j
O7xjyVCBCl2+iXvPVr8lyimvOs0Mnum3wdMi4B+FA1DxKLz7av3kDMVidAxDtZsJdoa7tG9l4fsu
Pmue02NVeOkvgSG5AnumbYhzwyw5ijPz98qvgQ2X4tECFQdVJwrlJY2o9h6RsH+HMl/eeWSy/SFE
reAgNSYEBmrEejQJaX7f4KFW65Tns2cW/PprlzbB3EntAmFqGxh8FtNfl1iujtcewV1H1YjQjNop
lMmhXP6NpFbu4A/J9UoVZERBC5I0Kr7HTN5cU9VFzAo5n3hPs1L70GJ8ekuWly5fSYOzqJrUDcjO
iCMkCVvF6vvQHMOmXqRTjOtKvHGl23wTMPBz6SI6bsnYucDjPZhab2/4buNWzDuNq2Bh1gK5FIED
YUoBjnCL1sa36yal0kw3OGN/Fm9b4Npr3cy03mfY3Vu8DlheBI1WcuNumr5LD0RhV0eTNW8AWnlj
ZBWkd+Gh3rlkfSM3xF885XU02CR8WVOskWtoxtPTlhP+QqKMhFgVDC4A4fRroxIFqNBf5/DWNTsM
UB4lfDqPSd7EaCXxu5LmxMtW4ktEgTR9F2Vt3CB+iCH69oNFRfxy0gEpQtjndgYSG4Sc8v0i8sXd
6h2SPhCdgwvCaMhxEa6DQ3nUQ4tnmKX1J1ZGe5+Nyl+QB/50g5MUWsdW8KDjSGjuhGlkY3PyifhY
phD8H26FTIGAjfU3BxiUUKspuI+ZbLH+MSs9RSJBNnux9rwR0jz+eIG2O+7vmN7kGSW092TafsnC
muC0yzhz7wighefUADXBu67zmu/XVMm/g9+XAvyr/ujK7kNjaMayYz3kJ8aEolAAvEt21kvzrXWk
P1eykjLltXOpohMFKD72YW33WG+dg/v+TQtoVobq0qa4s0HEn7P25FAqywxJTaUo5GHRkZegXwY/
tbnfUe0E58sx/5AG9ipoFLg3U2r8J2pDSPVXkJjjWpJeAG2LzWBfgv5ecWB/Qq5jH44vwT3ZqgXW
Mz9roCKtb2WihhZmIREnPHGLYvJvcW8rV7Baj/EiBbJ+dHI+4Ia+q99im1RESwzePons3cdhewaI
vd7KHtsUsPNzdOof1mWm5Dtk2/itOmzgw7DP1V3l/IZeBVX3J6BHGU90MuSaNprpca/Qqs0QDGIP
C0VM5wu93/E0BZI0pa4esKkAUY0ronGVe0N4lPdi5ovFMPGxgjrG3yknS8VPcCazXbwqkj09Ak0l
DAwR0Chj6PWtB/ee0O/ejxeZ15rt+QM7Hv2G8J5CFMSPmyHPQjVYUqwLowFlBexnGaDamPpfgUDQ
70VztC4GyGQt9NtKqF73IGMgu0og1cYnNdKtATrSMZwE3ZHp8j491JTKTottIb0CSlGMj4Y8JvgK
4HHHhrUvyQvbYpQJX66DaCsC/6aNnHkGMuCACjpa+gAMVWN96s8H+Ouorvo8mkABBvCR0VLse4Mn
Q5jiERDmnmof9vrt1RzNJQWGTO0Hsq9CLMmqwbmtQp6/wgX40Oa2AHy1MiIVVHZCaqIml4Cp9fID
/+skLqtPZrRD2WwKazuWzGdrb2g8cRqwH77XFCDRMolGT715N5v+0w9AKcxT7aVDLsfsGlgGxGZk
YEcZdqrLMap+lTsDYUdG0vrhD/F6gGb+YZ0Ju3Phz50PvNl7ffZ/1CEpbCSUnOu0IHvY3hYPdei2
7Ki3zcJWrL4NfLQQpLn031hVUjtAxJKTlKu3fTQT8kfC2wIeDrcy+3KSQYw8IRWfF4IWMuYygMVu
qnsDUUTU7/49voovPc2Xopf7ARZfyUJPx+82MC7jOX+fg9yRVhq3MZ1iTNKLflj1ovLm//Zu2AJL
uq92bsaalUBlVmJy0iNcgJkP60xy65TbpPmo/+5GFSthOK+gPVI5RUkicafoQA70FAhnEJZuTRj3
3Fno8cVqYsyiBtBIhjOMNH9hh6D7/6NF9SzT7yqlRMRA3Yk07yy1dQMDaLLI/yV8SChCSeUpI/4V
XubnkWhiyEd0AbWQXdQiOnmHu/fRFSnKZW9R3d24rfstbysH/XPqlD4mmnHOUVvQgPyohK2u51sy
YQwUeQMOctJsLZQ9XGr9BfDFTb0aqpnQpoWiBDCd0KbjwFCR7t9mkeTuG5KsLNffKLd5/Ut9QReC
ZGinWgsgzqMJTGj1U5hZ3VzQbI6eygdR/T48SdxxH8UX6uGYU8PUoTjesFyOcyugHLgVFugRxIfn
8jl7eQ4Zd6US6w/5UHVNseGCJinNtk1mIFGO1rtE85pWoD730F5oxEyu0XN65rgtvt12DZ4MWDvs
ikkQNeut1B4prPP5tLESqQUUx0a62aU8H7BJ+gGB4KhfYoN9dkfpd1jHofppssSDyECqpBwVny8u
UJy+ld1//1yP235ymi+xzr8E4Z5YUFrcA/A65ulno3eH1fAtbjY+eZjlrhrgBmXPfoyPXZdyNwbD
OsgzLehRgEyRg+R7yzOWa6pkI3PhBlMYQgpPnVEhKYXd/ttm7iztQlOPB4T3kKZB3kWiIduvXS+t
l+RdMTWP3LYLzppXoOnMyT+eX2I1jsTAEe5tDzxJbwb1vxRVpdoIe9SupVaz2lR0X7wvYWbftCR1
pX877Il+ydNKb3/+EPBLOinPlf8L4CGw8IgeWRr8lCw5HHQoCH4QInT60PjAr95uVWHDlhm2UaFd
6UE+FIAcpzunBdoEdO4Kgc9ptDNjeNVN1HDvZ1N+dXCtlF3sA33mU6AfDV0qj0PFMOhBsagVespG
s7WUU+h+mtki4tN8oO9fBa3P7R/OyU8j2vlOfFbaVuxiEjP+sKlMx6jf/rcB2SAi8Ryg57SPgGka
/cbUIzOEMVruhKJNDjqa4E+fs7g+qbTKnVIRwvxTODRrAlV+oMA4KfPsvO8iotY7c25WhdpPPxXH
dCN9KozNLibD7pHZwt4afu2Csk1sACAdCOU2QbwZbpedRi3wkzTgRF37bk82j7RhYGc4U1xoHq+O
hXkhQl4eAfk2U4NtjKhkziWu2CqzBXS18dzYRLjzZGQWTgBbachMdicTUzahF8mXS4ChMW6+h5Nn
koQdJ3pyLyDwwW20JqjEMvgf0IWbkWDlhXWoZVLK5aHzU1G5xzVgHihdPTlxiayNff9R6dEm+/qp
joms+XAydo7MCFX1nAYmYp6UEVt7D5akIBPFIOXHK/nFLQiAVt6Yz5FdwKhi+ndYGT1utN1PQr0t
FJ2kEdzSuEMkDxaMacNshpAgwBmVDXiazHC6/O2zz1P2KWHPuc9si1ZPyImk0kwEeTshm70MC3P2
jstjn6RiZwElzdGjXO4efE3v97vPMW/5FK7ekkivDHnVaqpgVW+HtgAMiDCF9BTjXx+YEZIeGkpA
MG/Ja/z3OWxF8KokTBMj7281w8Ksu7jBHQT2u+RRv4pG5vUWlJW54bePDNH8EfV8+FdW1TXvoBAE
ecXLMCDPqq7Kfxkk9xIOleglDksqnP+EECxc0w87MENCdBfAThKaMWYpTRqKP2vaZD+eo4aWkISl
3cCfRa10HqEMGT4LykW/EWZjMDmOaJhu9mziexX3Qx+RNVxTAarYgncPIJ+hmkBeTkjgdcuIfjg3
6TvlQXxOMbj5JwnH88dXwmOa51Z7Ez+pYLAondBYJbcPYKVI+NYPuH+OO0BAHvb6KFd3e6bK6DPp
KQYoQ2bk6gRFUOUy0k0rFF1Q6aFCv47Tu0pxmE6dQf+ebvKmH0WaRXru1XvmYFuaYIWnR3L7W9uw
NWlzDLM1nrMwsc6Dm7CCZ1rCQKvXA5Er/TAjm7lF9QNJTB1nW7F0DE7W9uUbOpnUCL9iGdmVngzO
ESNUGQDEnXEqwlJSDFCObaukAMUmo6/Qk6Ei+mWPaZqSRVy77vHkMuKHtjF0YU2bIYRSz6/8Jnk1
HH/cse5MMGNM85ZthKqcblWLpg4/h4oBpgdhlfkAnPyI94e2O7nMHSZEjifjt86fCPS70qjNtHMI
1aQ3ANVbhFgW8lPje4lFi8Ad9B1z/3t37tgShjHkDcCOd2QmJn39Do6Ph+10lAamZz0bMX1tGDdW
7LALg8U4Qfgmlw6SYfiemEq/Mtyq8J2RpvtmCZeIDejmz/032/D4AS2DrhYmtNfpslcGkbBU6zQf
i/7Srf9aon7Xja5Qix6mSfZD/zzf50Sl8CuXic6LlWuIAJvrvpH/4PIK0FrNAUzGuFToP12BdGYE
35mblueLGMGEItk38DrspXJWHES1/181Vzw++eHFFRIK7ljvoInFO4iSKSIcTdPwr01FFVhWihFI
X4OdETgb/Vws9+x47JwVK0N65YYQaNER9KFUradpFnNkpE4qHcG07BFCRLAA7oOPs+7X7197MTPJ
aS1mPacUWo5fImrj1xC1LCbb+2Q5GnlFEWUMQgmcIOXfYBQ0/zV1A1thHxuqTegdrXE7/M3eScNo
rddIvLGh44epHtv9aqLlCi86v/ogtqCgRvQ1xgMhr7mIF37AmaxURhT3dQM4J0PihZcFTpzCSTDW
QbJO1QfquMP4WzR6J7h/2iVb8M+Oz/ilA5gD0FfP0QV6prunl3nBUwbZ/HkAtL+ioBXM+m3l+WJ/
5/ZJRkNdhPy8lceJvshuiWDkCAjTTlarLmI42KkdPhMRDqe6dmm8xNa2wNH8AQuupWHuvDUB9YZV
NDExOcC6/caMPll7Hp8aCrMF4N9rjg7TjQtgscHCsCZhHhfbQxgyn6LJ5VxwCFd3zkBR9p56UfPn
D2XtX4fjairey891sM0kz1eApeQebHLZAKAu22KBPI4/YFRagZmrb9rzxrN7yTmFt9XKlM0yPVy0
ancVhOIuG/cSipqRaJ9r/Qwhqn9uHZdcCcQwUhCsBpWvMNaorQ1ZtHHzXNoB1cT/mJZEmJmGsquU
aMGctBsvK+4VNK84fIrIgI77fBBsMscyxPoLiYabiavy7XYi2BR52wmVnGaNCV+xVtWhRfM2bGqk
YEDoLhpdIv45h+fkg3p3NeRhELZpq6f3yqokeNa6lxl0PTzAAtXBxKd8hNhvHtgqzQTJAwi4GvmZ
NFtr1g8Pa2gxFv5yEGkXmRlhZv61iU2XXQie4mGeFTGHRuauqMzw4ouOv4eQ//QHkoLmZk2rsM5D
GrNeFxPfAoHvkg9nrgCF6KBGDq8KETuoC915TWvmK5umHHdN9E/rGC+hiYcCXQGUTAy/bKBXDKTJ
EihQpfphLBD8RVqY/kvSmO/aOtAsUVL6kR3QphlARLLPLG/PdmT23gTdvBUBZAABiHMxMNTLU8mR
x5eJuVlwgrSARmxrkPHNfbfTyibF4+mvkGPsqN0hbB4V+d9Iexwtdtqclt6hfB+GoLW/nJ5eMeN5
G4k8LoGYzutT+QHxnF6RH1Xu3MxAv3j/q15NEvAuMeCpu1EoD/qgsegbgYM4epHmojaov0sGQqGd
9VHoHvpeEzeMhjZxeJIx54dZyzb8bOc9E2BNIok3dlVt1odKhChb8p8QI8Gjq/7Hmy7BuDTGlAWM
TE2JE4/3nevxHgYeD2xTssMt109uQluFQonCcIfGEfj4wQ3YgqEaL1BBtmeRYTEt8MtCsR9ysPd0
QxXapbUiROlHOWSha3I5CpkQ1mNjhhY7WQVjFKNtp7//sYCb6GfPowQhiq5t6pqB4RLsb7G96qo0
Fk8yOcRspL2ROGHHTGS8v76HPxbFMMQgEspmEVwe4F3As8PCEGSAIhf2bdgd4H1ZpzjINtDJG5VL
XZUE8Y9+Yt08urBOP3FvMihk6b3iii/h1ZoL9tg6QcQrkf4X7yhiv4ac3gv+DRui/bPj+8GFqdOO
k6T3uMmn+cTG0ny6bk3u2CllOYFdyk5H8DkMMouxkYVVXrHaoXAc1TXZ8RCcC3rRi8nDnk7Z4Z0y
s+Fb89qd7BSLANQidJ6YBqr71mB1fYaQzCuKASuwy03er8u2aMbY9an6JQvuyAZD6j9Xf7jlIc8h
5CVXssSN/MtVwwZxbWeZEc3rcvhkZn3pR9oEGkhfNm6dppSraEgJ3ET3e1caO8qSjICjhlF9e2PI
AFI1Ygn4auc9380OoqzxUfRTPzfxbvPEm84C2BVY7VNTMm0/+w9pTd/JiotSrsimagRHZ1oAbGZK
eiZXaRPRfUWX4G0LzQFxeGDoS55CYRtMB1AO1kUSISMpcEINWNqFfUUjc/SA16YxmQALrcjczrLS
JEkXuQ2a8JXv6DG8R2eU4ITYFPnnypTDiygRxEGJjrMJwwFF4WQuSPUnMNpBWd0iqnnvHiEShpxi
RWPDwyIcEn+24mc2AXgTefkkWPkRnEa4EtUdRBh5LsGfepn5WLx9oUah3ST4AxVYx4ZDtTHhXkdj
yuCNjeqHQuAKkHIufsi/PqrhSh9QBN4PD/iENNqaARkXyY9w4fAzJXFot34UUcdsW3GdMT5hSQg1
BYUx25aHPSYMc1bCDjkFNy3YCz9d6eIb+oo2h4cHZNZs+N4NtT33yZzwdVx6PHm1jmjTUK1AXdzL
STajle+LSVhfxgx/FSdsrHVujmmb5t6v4GNY+ZVlQ/dZyWnn4iMPVSGvene0mX4knsBNh2zSoTi3
AkUL3a1l+ezPKd9wQju160DCI03yzQyQj9FAmzJGSQM3gvbPTG4ZdDeb8bLdXiDmmkRWsffnFFy7
/poXOJ5SmwtV25vg21n2IytfIgFQUpe6woCF4h9FYK+kyy3sIQXK5gQBP248YW/d4xVyarJ/lYZ+
2TqONB8lGVvyIbkKH/0Qs1LrGoFdMRcPthA2EkBifwaZUohlE7uKsMmMM0PB2OdPLMQo84MqqZus
L7eVRyGl2XpfGxrbZFN2BOuUcyoegRJ4gnvGiNqB+nX5q4jBorIkAqTRWAG0vQAjT/p7VQLvOw07
FuFW1XVfzb3JOIgjD177CZD+xueuU7si06UcYCuP9zXy4F6WRwMPof67/Eq8r8Gm4EfOldfGCCSP
HBAUO4oIlUBXnLftYKmyY8qFp1S8rtZRzjWDNMBcDtcQB5I28EKjTl2GJumVYc4Hzp+zmcU6+xEH
Gko7UTeBh/3N66rSRXAk47+PY6AbEpS2dKFDCaWRcWE4zKSvnmTQRG00+Kqa/x9iTwyrkrjX68wG
iTeDTZ4Id+KVtrmQEDSVgfKbUwJUIJvP/JgL0MuJLnuvF2waW0PnF7WEffpVppxtpTRtqsQLL0p5
pHkUSjQOwDkbwffPaW1vLx/ptva9peCHRf2OmRy8nGpV1yA3MNEACF+C35rxoTYTbrP576/2l811
yl4xwQoSWTf6CrX8lvz2kXyYa9XxAhcVqn3uKkuylRCtlSYgsbxBc1MozMOkLZ2T6GC5/QrTI7kK
Eo1xch+cxRvpESdksqirQ221yvHg9tLxkNMM++TDG6CoS47DvCGfQow6ty+ZkAdzbFYf3l2HCkmn
2xch6OL1YoYhiFsXBsH+EiIhv7Y74j/6PcIB05to5u7lPT/d2eBN4py1sDpJDRhJK+ucNC3weA/C
W8IrBoVd/mKKgtTp4wUWS40S+Q4aaB5AuAr+opPdVRhTAL0yXwGPWsFJlJT3DqmOCa1jDTMzJ9qK
JSh5AnCd7XoHu5h8pwbsul0mOGbuuMlgEuOzfy5ORazm7UNMxHN22k3cqzG4aPrHYH9JvBdBSGqO
j+VHn9H/cYMKQEkb4NeXBBhd8YzGN9VHXq1gZjbo/TMoA5D4XTH2U1RVb9sqo5XzbRc5pxROboJG
lLSCWKwE7QdS0OHF8gckmaUSNt29JGIU+b0zz7qTksqiPxkQtwPiYhSN4ld/X6Um4OUcH+Oh+yog
+ct+HAU3/JvYdMQ77wU0mpJCH/N3DXtWfD7PogxVcdGCccXyFxZnaFREBDBCoaa64+A9aYYMao7O
5N34E+1QYbTLKo8esAIzQiCVHM0ZMXJ2TV1hYJdIiRWBXBM/x6GyUKmeZdIxM5/yMpCS6FajbCoI
38AIOn0rDFKlXx9+r7N6HqEpvDu0aVANjLA/E6d7gpLDPQwQPAL+jh1HhoBQwfNo7qEHtWe2oiHt
FBXuZAQuJVS6RI6ZlYRp3Mmvf5nlsRzIRLadOoTWepcEIZ0fl6vXlYVVfi6pY5jMqMCfXJA3S49e
QXI3T8rCTKi2LLFP54sGwtEVQQkpCXAqmXTY+mZv+cmFMHpKnXnKNumEGq4IDKlz6os/WHUj24fY
8Bq29CqhPr+LARPUe8gfbky0+ZMCul2tHuF6urIyxY/CHcPFgxCMSi44y/mGyYMuQBbIPsOVqLDU
umKdhlSkLPwwp8HwlA4g19wOksqHx11hTge0ivvw7+RKWm4V6f4qqMOZp7lXj01YEkCOFbLMcrUd
usAqA2FkpNoei7zq3NEtmBwy7PHaoP4/ezNyuYifP36VxU/FdXoyKGLwC0ELaem7gIi7yMAF5J+7
VC/9n/Fd+OzI515MzfnwetXw1bDiQ0vA7nL5uoA9DPQ25TXs56oa4Bsw2S46sSLB1ysvMfvkzash
04OZ1zKFYwmyCAYfEEuUxojIrHcPDin6256tVZhAVinOm5nRx+u5s5GOv29DrI9J+T2GGOYolBLT
/3ESlZmrsQep9PpWYzt8/kDkdsJDt19AbzSTNSkSqb57DD/a9QOobUXVA7FOGpBMgct0IGUyU1iw
I6/3roketK6yAxs8iaQwsdhJiZCiWFIj0wPDbWX7L7CWJLmngpr/jVUmxJd9IiCZdw2cMMmo4luf
Qu7FTLdbvp5vhK9h1vkuKrCq8I+J4b3EV3FGR0Doz+sMy68TkmYPj90F5QwxmrIXvXamIXpcGzFL
LWZ1j04/Oiz9oF5K1Ug+FdGOrREG9lJ7HMP2HRRYeoutVttD3isq/F+HZqtPJZff8TFP2NTkPBWk
AMmTrAXuQeExc1bpyyyIhk8MWRfMIRl3fqadSI00I5CjXoLIJve7f2IAK9bpHZd/w5lwAKjzF4Z0
4Vy+UnqHnk72eOVWukLJWx8Twbj3Oy6tG2TIohWP4NU/rE9We16UoiIN5YTISSEM2e6uqpya8JDg
7Kl6hoUcxhPXKafIxzrRSouyFLEDwHBTJ8cQ8Muhxgc7Xa7c7xFMrnyDbWkPyc4w2+w1qQu6cJ8p
nMm2F+KxSwfagkfvCUgSuRzYiI4cJUACPE/b1uffrNHlX7gih0os3TyT2Gi2AudgjusElJXfBotv
Pjtk2TEgIBJeqn9LPQ57vPs04V7kOLq/wHahRdOliyvLct+evlD+k3KBleH1QW9JJy6i67tEFV6K
IXAq7axxRd2gduU3eWK8l6kvw0gGBKuYkIxclPxsnRVoaW40bYp1bDkTFhr3efWHF97ox6Q3Qe9G
/hBOQut8IDrwCDXhex9GbYTj5pLW33T+Nq/T32MqbCCmKo2c07bKr59aP8vYsSZuKfT6h1pVpbVh
UXMZZmyJIL4xReXT7otBqvDCLu90Iexqky/7CwWjbxU2uY6wlr0NJzpDDEmQUBMeIKLnr92RwPhf
tXq95GrqY5pgKPuffVfl9Zu7G553m5Pb1wYp5QKh8xxzI4Q4be9ccdP3hhWkt7eHyalIv0rufR1C
TaG4ZVz04a4Y3gK1FXzQLTbbGNXhi+sI2+EF4yx7PtcyMl9OD88O3cEG15hA2Pz19AMYVGDVFY9j
zk/DIKjROziAsikeuAll5XJS8ejlxLyqISHsDe9n9NeJ4TlWqhGW/Ymbc+T93DwvWyMKHB1SJBsh
E+15a/kVaCNir+vDwm57kciS8aQf4A+HGyGvYcA58iAt/TPcnn2CZxjMwv+S8aClaZwctYjwAYJF
Q6/o7kQXb/SxZt51l9HkrLsLiZKi7oAch3jQxOQILTUtJtlEvyRqBAaG5CtE6wSnw/zUUtBUxZOe
Kll7+CPEKLNTi+6ahexOqfh0ytdGl203niSldUZkfGazn3fGZUdCq12ArGeajK4Et4GAr0Cp74+4
hOAPGATWqktGYzOgQ24gWXjIM3/Jkl/74P2vs2DSTRIHXUgA7Ux2D6AHhBvJ5EtbiBmPDxcu1Uvn
wZxXLj3smpxWDKTQGCZxlVpwIbnWKRKKbAoPD2ipJ/e1pwPe/zQWaL4AGfO6wZlj2sq4U5JY/uvV
7TlOEaaJ7tbRqEDijgF7QrGdDGLP6FqJiY5pqRMqFIaufbGS7Y/lJoM6BH/3jt3389ct4M1Zhp0m
wOu0R/NiuYG3vZgj7mQgDhdWzYNW93VJkYlP+XEOxUMiBei/nWgXRsz0y4q07SIMqYrbGpHVJ3Hy
W8R1m6Z/qEdlAa6ErhiR41oOwL/Bhcndpv0IYg2GBWdR2QW3LbosF0a7eq0UM4KehIWame1sp2E8
KqSc3ikt/IiaUqsbmsrRM3lYe3vFyeXHPrwHAzlQP3gxFQwEPb45A+XEQvVrqzjF+9qwJR+RzZQc
1pPGsTipYpUlw4S5RkpuV4RhWMoV41DwXdX9InaqC8EdtfITlOMJjnwrt656kMB0rZDElWMIaioI
FYfhvF3ARQDox1o92f32MtSevTcQ0ptbI/4pi4+myzwCY1wIDHPIR+39svt4h1X37OAXxu8D7ULK
P4yiHxKGVL3aV2h2z6VKcbqOK+qhfe5u/oBclCZS3BumwQ9kRhKpirUBOWBqS4zLVfYmg0L2VBZZ
vcvyrh1hZtWE5Xl6QOUWnIxzQ/nywhNWYevDL44xrN1D3QhY+vIgPZF/NmgEpL0WqbsL8iJ4mrfo
O38v3M1GcnEk6FYdvX8Un7xBlr0Wh1vLkBwWg2F84Dwwow1P6VU8Ttr+GMTQolBDpSSzlSFXjOWX
Jn4FoTR4YIh2yJpUv8PBf/Ni8961eX1VJkjHsPolmHPzqSe/U9iCCInHEq9MpSvko4Cy/9mL+1L5
rxPZ877jbFzsc/mbl6o4NRSWlSi+4yEYh0jBNdXfOMfg5B2px7Y9NEdmrIKwxyoR+72WWLTof4qF
W37wRn5VPbAg/0Rdg2wLz3c+/7fczlfh3oDZabkg4LJaMxnpAVIC0NbJh+ui3/chLmEGmInUl1UJ
fZBOZSfR0b1ucM1qslCqTuMxsbFZ2O/+BBFi9M+Aqc4WI1NNne28jdHdTVV2Q9i1ivfx2fpsIsRC
KE0O8md2lzXjWvYa0VIqo5jZ7cuCWdfB+RSET0Yw889CP+C6n0f5k7k/Wkq9xyL+ucqeBBi+eO9s
Y5Vk857KCbSFfjNI5APjaok5JO/PY6oR+HVf5EmXWFgIqpK0OIeyJbV3fwEp/XUfzpgU0hz20jtw
C+oPlK1lemp5HvAYAiAsEX4ZYZJTo/RhRbUa+iIc1jlEH+CPF6vv4YPKx0Ex5ZBMlsHlCwhP9MTq
3VwSt7tEummRKu+19ZLxyBvCs51mBoXI3s2xR2cBIa3iPIx48ZfHjEVXDlL1QCi1sS/sedvu/bIf
3WxRb2/PrhfHh9TEqVHNYajTny5Mo3IHDFoAsWv5+f1IBpDaHIA3fN6mORmeRix5TjJ0MovT2XBd
Gp0elbnXzR7R1gy4FGi1pbblIL40+Qqsrk+zCEdoTgz+aLjBFdS+gcJlr9MUk6Uk2VczimGnKqfh
8VGm/ItA0n4AY9qLsaTNfqj+SmennOcOmKGaLuIMayNQlq+FfxvQyD9Udifiy4/Pv6hXyCMXXB0i
rD7uiWmaJv+JYy55eHHiCYmUYFFoVa457K1sQsgDdp+EYf1TWMHUdZuxjHV6HQkyViz4F5vMRYtY
NgbpNXJHIOfN9FujZyqiyXiK63367sMYJGOHqut0WH/eUpB57ebGFlqjR1qEIUJSY/HTTCXgp1qG
g0e9qNvLozXEoE//iBPg0dKfWEZO0aZMPgVt8KGu6n7HNIc9u8ea6P8qW/kZopVSvM0tfzn+D+bR
Xzhs4sHo8IjITHmrApVcrWZXWn67yRS1sZj4zXXnZVHNEnsA8j+te9CUq6eh6eRJyL+psuVBugz7
9Dhle7/myUhf9i5iUVATrot+QXuFLeZxFAZQXoGjpN5sENFrWXukWJEqvPdffr4xDPEnIWndgt+r
lLo0LUtHZUaePl90ubpQ5jSXzfloYIToXMN5ocDv0eZ6meJxB21JodnYtyFLlaHjReJ5maEntzL5
rL9pmd3KPUKQDHLCfHtbRAh1RycdgCof4p7lFO5H1Mo1iVA8U2kTk9j8ucgExSrvo+3mdv65WHFT
gL6XKh3FD7hJ5zZMhgKxNA+xQyE7VvE/pZ8CGgHax0VYL4Etv2pXkiBSt3UvFptIOC72aKVBxtbd
jMyIyjC54VNHSJ4rfrcXz+QHBVHK2qfFCvjDPY8muWgPiey8x7ZC4ISL03s8h3R5h+dk4MEyGAfK
3M947TBXZ8o9+2AXF6js6K59slEnPHqOOQJzqU7f/eSewwe5yGEiVOcevEt+LogJPvh9cEZoau66
OardqfwCu+mXSGUF+ccsz81kxetPWPpeCYItVULGoqYdg4jOiOA2yXis335u529H0YNfQFg2Z0+w
t8UsgD89nB8fA3xCxrF4OnzcJc4MXE9bcogVfnRZu7RjzI3uDeDUDebYdCmWPaXN4Lt0h721wy/F
BLTgsTl0gQcK66T9EMWqZD9P4YblOD4puGAskQCwR99Qp7Kwb0ipRn0e7oWjoNDb5WoyHu4oS6E5
YmSkhUuHz5nxAbyuKgkyTcJiL9S4vjhy7wMa7+M31oS1fS7lNo0Qzzadl+UKo0xjNOk3BkYIX8ee
9KTai2zY6HIQVBmDixvoj9ZfEkfzrRa4KnnSgCE8fh9u+XQGhs1w4ynGAapDwAl7/h5/tx/8/TeF
y4sQPGt+fJa/IVzBQfpAiySJDAuYBQDICJ083xcRoB55XsbH8TNbhn2C0ma9yNaPIgpgWlGKczVn
BnDj+H0hZG+2/gUPykWR6am417qqCHAaNdFBcAs8ZmANxtMTbcUgRwAjyAXnEUeRnfuymysXi28a
VfxxHQu+FyQ7ZIEVyGRxlEDpLCNtYvJruyX24yZmvCTKkQ8q8J47K0FYSfxCPZ2mNmGIU+XLoQLX
OMyDlx/XyNQxXkUaA3GawwAwZhI5NkjVQFIWkJQHDRvGzabaWVy0OKRoyvmt6tSwl6iomuSzjOuj
stwQasGT2YWVKNsHeehDodNLJvABpnB1XBCBSZ1fyDB+EVfnKhj3sa+ClarVkLorLZkJPWhaRAae
3R438jo0Ks7uziU51wvbwsu4f9bdZraUE9FTg+7pT+LH4PfYbl9NcW01OlMIYFBrNGIdL+b2tqrq
sawCh7ODDpIH0K8zhmcOh0+nFqOdIzJW/1KBXB/UGRUL9p5zGKQZHTFpGSiKRDCgaIzPOKPXEgkW
4j3Xwa9CMrMb1C+zcz6/P+2yTkUDF4iwZScM8cSeIKchtLwcPzrMJcimFKfpx+dFVSkJIGaI+pgC
i0ymcj0PGj/p+fltL4IHP9MTePvZ3BKz+HjsEiLYXmsQe07qeG7r8ELtanRo8Emge2PhzrJ1Y4+G
5LKg69MRsGqLRykpwi/B0ElnK79enR2et+1sBrqZ/SmTe5S6ogPwAGgWQ1DZcTS99WMGdbEpUsXt
hoZYO2h7kr7o29pXQ1rG2Egtvsgn3sgfEJaQlSnn3kCrw94XPlh526CugraEFaHedqvhA4ZBz6vn
gumFvfETngpN7105YsvTsLAPyCtAmJZ+WWdPfmZOX2bjg4hWzpDdc49jRhUWZ2KC/kdN+vn7rVrV
ilVd7y6oi+d4jfQoADBSHbCAUjhPEOmCcXrNziopDraX+U7nAqUsTbYlw826DbPiABk0bdq3ZXi4
Jal02qKzlZQ5crspouqH4GpKUnwXtGW5yChTf48sS6RAM5NMR1JmTJsvt3xXIzsbEouFhZ8OMbse
oanFKL2DqUGJj02iqMtW/WJWNh5uInnT8SQHP8YKk9i4IrZELzdRhefrksckZWyaNJNb/PwcfiaA
ZKDFqnzwawH/ysiYGlMme4rPjexF8HkwhaE4scvvrtoCdJ61ssbJLuxiigguetBFhAnMeI0qc728
C1zOX/N5zfN/rf5LXTdduLREHIwY9mLUBTKbia+1pql/Ox+h6rOyZGOp6g1X4k8vUfWeyrmQ7yUE
IK2fcLXAsJSTatFm+jCXuAt7UWbeLJgr4bw7eOqQ+JZIZmNVC2GGn8x26rKabi3v3FRfpMVIp88G
hv5nI8G1VjDvfe0sjUuvYl1tHJ5Wl9SHQI4YI7EHzZhMNmdhgp6pOFNntoVu2HR61z7pTWje4OoT
/Xf9wpeJRIMTNP6MGULvz0h33OBH77Nj4l7Lkf35Ima3d3UccszrOkUJILGl3GWbT28BcbkSSOnN
FYYLzftn38llTbYD++UzNHsoLoSmyag3CerErmAdFqvjGNfVzGm0oLTdHEUJgGLOIayhu7QTF3T4
R0pU9KxtmuP2xY3Fx/b9yWcN3S8aihtmavD6x2jEkiZzYIjrSZ9peWtSh2KQE+cMBy4rhI6R5LmO
ZT1MkRO//f+035KjArOSUgque2saRAds/+W/9rhbxcdOFD0lVq1rt0NaLzF2rJQ5wWJjjAvLPrj4
3jxxFWRVBXt+Xmwbo5u4CP5UpEElslLVNMi4Np1x9OWBvtYvfTQ1z5Fbjql1snIF2q67xMY2UP/b
lnKgawaw6O4R2fI+uTJ9g6v8+90Cbr2E2J2rYS26qwtZKOIRUHU5ENtm7xbLVE5B4EeThU4S3V9z
wQ+3UmQjoJcmEHGD2WwqZY96LtO+C/fSl7wBw1rHjzp2fBX1imch2vkwJpdfKyOVqwe/uJcN3cds
9Pcm/5NlU7jy42LCM2eE0q5R5RabExC6+v3otHvHLGj2fqwhsWdGNvy43aYYkWQXICwikTnjEKkE
sxK2jRxsFeEDtfl6T3poTabaKqQiWxSiOpxRYOV9lRv5X1NTrNS0ZrgVy8htiZkURQnkhlIDhPM5
EwpQ4eg5OQe16OhEBktjFC/WXw/lkyQRO2W/3XV6/BbB3ULwrnKEBmmIvC1R9a095puRrc+lt/Qz
Y7miWu3Lfpx4N0Tm6QsX6Mg9SMAelwzPAMsjfydp0+FlWfxaFThIjaAZWM6RkddgFj/VcrodhEKZ
sq5x9R+NqjLKSFyrjlP+wJF3RDcMgupH8lz1QepWFJKG3f+kzLtFmBuOgkdoWZIA0oHir+Km8Uyw
/rO76k/q9Sk6jkXyoik3dwZSnBcKAa/xoOSr6eKn2LMakqyEcOtvodeUk55hUv7Six4GZBduzcNQ
nNdqWBh7TEjIHnTZu3pgbxXE6mwqKOZYfiCqK9sN5/5kzZuaACmsC1KeuMJiWUbgqhW/Zz9L6SYy
lNyq4ZDsiZpbWk+VWBdvlecEYFGy14hVLE4FCpgHfGWY3FWZvEET0Vb5beRCruLJhn3j7e4RYlaZ
x/vrwjNBsswbm2+GdRZaSZfQf9EON66f7iz72VlXvY64t69lsDYm24E7KuMBckvv7S/4m+aglt3Z
I/cK5JGVg8pZCBeRw5xfacwqwfl3/4zCkbu8EUVsOruwTrbFJRIAs82ZChxbO6DVKWsCzDDy0m7J
B5MOU/MGhdayJlrsw+DIVO67m0aFHw9jfSUO2QJiKWlBRO/sa/AA1N8mGAZu33VdCrpg8ZkyJDVX
ebqpf0m1xpUYg/Z4lq4+gOMbgTq6cdoWD68jPeZVM1SPQD4xGr1C90m85oGV56JuOxsj9NnNeLAJ
5s2KPbhlzC3tQuCwhbtzQs9HRJrc3CfnvRAl2ib+qeOwqJSbbuBxS10dF/GebWIzUxW3l/wDmn3z
8UQiG+oAcjQ8cm9wr9ebi1V5PXFIiBUUrulPFX4h9Lxn0VyiU3lWvz/yWonKBPKXznVB5F6ZObzD
QigELiwyrFj+BJ/VGqG79sd9pgmD+iQWosz7zC1TEF/9ngXYcizBsR56lZPJWWU5tCg+H8dwwFia
avuoNnK51b+THKOusFpnqDkcItCyJNOSIkK01MZMqp5LwBqknEbWbADmS5wuZE8CkNwui35zu2Yu
Iw3fQazMhOwFdDH8lZ756h1z+wDyQajsh9O5boJzMdhp/aCBA5QbOyAmWPSzsMIdbAxROZr4Kb75
fXObZTjX0GR80op2wtYIkbhrkErY3soOh6bGRufwlS9NBYNH7TmweV3u5M97RkRph5oqjAQmS3+0
EjMLFpfCQ1Q5vyy1iWPyN5upDq8ETNsWllV9rBJya68V/Xl+oNW2EKM9VB8KOXGrIYUq99iFvzef
EzfXcY6Pdnukl+Dap9cxjSsHiIeJeRTyClaAm4JDxiL73Pf53D7H9+4+TR6epKd7RPPzlV6EFuGb
K3B/ZZpjANjUz3l68fCc5MieP3n/VCCoEtGJ+NpPOtVEusCw0MaCM0RzGvw4qeGetD4kyM64Xd7j
DTQw5WcXZGqNWEZqC4DE4lXXU1TrOBzesktfRqwu++btuiApdY0MGIv8RBO71Sn0PBrEQ6nC3vHL
LlOrTE5nCWvE5Xgn8b7dm7n4KC1FI4MrrXD3XiETXYXoIQJCLdSPpcXRv5iiIlvDu3j2z1aZiREy
CVE7XiuikWK4ka9n3LLFhzGilMrHBcrrRXMd6P3pogqEzJ+PrYZxG7I67BMjii2xPgXJKMDQemHt
bbc2F3dJcwB/L9RpnxyiPDOIN6o857J/uUxelTECo2i8zDbyKRha9HJQ0C7YDbL6ZQEHWqUEiQNT
CxMfl8gpujebQ3Nlxd7DjnWmdAu5wJMWKEFxyFNAw/Rby5Hzh0hqTEIwx7b6tBXDc+m1Ykoae/LQ
JVqElwa3XpQeTUOkwS9NkWxShYAyMLsLQlfBBgLRGDttqE3aR+T2FkNSO1xq8Y+71PQdaOIuhioh
7yjepob22IDRT2brrcuSxBvcoMLm+HqRgzg8m2Kx2sKfMSNjhGrAtVcrnlypUxVTIXjcNK8RJOJ9
riBsdwJSDw9W3YXldh8EhgsVgqTeMU1URSyFjColwkgvx/yyLy25IMtqXDVbrHHFB8gsSdZlpna7
69fNThSMlEOYPaGA5JvVfqRVqakjJeY+ZAcN1A97jGepjIOUJX1tZQrpsmHbCjg+XJqu13TwzSt1
yp5MAyPmEYlytmlx6Im/XoRdhxoEdoBD8VJ05HXlDW1M4/gCvfxkoZPQHzX8w6WyROJ7xJeRXUQ1
usCgM0Ov12/kRtV3mojehhxip4h2Ibc/7fJGzaNv2E2Uf87QiMJfVaAIocsxKn9DUIRvkP/Kcv9o
cukSu6Ix6a8oiUiPkAlC/0PoeiT+yCvwvFpIfB/itRiMs0AE6EMs+hLXepxLCN5wmwF0YqVNbasD
XQwjFbr+N5HKw8BDLyrWKjk4qUGhmNOTSOaGMWYc9PkJ7Q8FRTXE0tckZxY2p+yKMuLlWm5lgn6L
vwArZmhbJnBjKm5Rh97/rq+H0l+girosLTNE/YHatFYtlmDrMtGLv2LooY+6TmtemLndZVTJpXy5
SMQ+JNsJWmY63an7uo9eigIRc65Q2Q/f7saDF+uKlUyNUy/6PDjOfmS4/xw8Kv2DAlWVBwWY6rCC
TQSmxycc0lIgbA2Xs4Q3CsX+vUctkXDJBvFGq4yn3cEEyViiAFIWc9KDqgOQgVbkke5zssioxDEm
oHevrg3WjjmFPuTYQExkqQ+pRdUjD3hwZO8KyHwjiknRB6SezaGo3jWIPZzZbi1G7ppBNi0m0GS1
Mby7/OjpPaF5AsAkSOB/i+AFEqGDKnhIf5VxAYzJx85/U+78tOGRpvyOHFqezTPCVtAwnBgO0iFI
TRGQctA0belaQbKQy5sBp8PqWyYVv8kjdLOwO8jOrjjXyTUZcmGTSCW7dm0CKXDV2yrz/1Fpqse+
Af2nXcx5PfSoOlGVZEhA2REpfIFbcK8s6dMAjVhkNuMtPepbdXHkuj8hPBnpLvZUYN+mg0UoesKX
KrwCBne/DkrdBoIed+5fUNMMMJIlWooLTANp1/IA+lbs/IgEwbz5hb1Jv++ShAfbEYoY5z/ayugD
mEdzQOl/89Nl1H79kwFZssOOPIdUPh5WnkFdKYE6fsD2f1LzCI5jZLITy3+diThaP2wrL0iYEGRM
YZO3ZEoBoxSt46qdECRQU3I9ry7Idny9agmjwti4scheTusGojmcmQljoE3bH984pSp8ljGm7T/s
T1Re3dCpDPZIXWynLxkiTfpkxjSfqZTKzkaypB+TPtQcYsUO3VnZyhmLtZ78JMom9FyxwV0WWxFo
PiS0hYsawpsBzZhPF44TiMJ+qAwqbi6FA70CVE6gt/ZCcCq/S+K7jHCzDM0omp5cq/2sOmTLlB5G
p53PWrALvlY3bliyPXz/SzOdyTvJVtCYIy9SC3zEb8lyaZBfNLQNPwehy2Yup58DDww22wK2AAYU
787aB3lGpsSJch6PdYbUpxx3jdQyotXXn7Ur31qKKmXuIVrYqOdwLHD5mhuxWlaZgaD0ucnhQeXE
GDYPMZGw3cfe1eT4NOOZCCpfDzickoIJa1Rhu7eBMQy0UJNsdaSE5Dx7vRW7b3PFh+TzbMXXswi8
06quPUNGYnoJVymGLLOTEf5/JoR/NPdkF4Emn668r2CwH5WQ+VhSfwbp/eT9KnIfzwj7YhGokSBl
H2imjnLT0QSBP+8W41+bvfCiIb+8J6dyFvt6sYfAeV4RgHuTyIkuCCVzOZbgU/kDzsGblBRnHjbr
Yh2Ak3iKNtPFAOxHHB2G8UJR7iiwxlbEiGpenS1D1he7MQ4QjEE+TG1NN07iC3mMjJygaQyjVk78
MiB9SnumebnpufeSF3SoqUpTMXMemXIs0QY9PRgimAgjUyoESNAdVDN2hr6GkKoP39RLmPn4CJ2y
wWkgXADgcQc1r1j6Fqza35xjyTCZZpmXbv/qDYw0evy6esI7UbKgHZqoeNMAxWt+vgy6q1lFLioB
cL9pocytDFrCvJuTKrYLjNZhZDYd7HQjl9z85nUGMyYdcTcKjoQwUMz/FeWIs8yCCdcje/dDfeUk
SjHWgAarqHqjBxIUNrDOClVRrXgiGt2ZS2m1IXqT2bULgNZq3tyRUkWCOvxclWMVLqU2PEzZUcGl
sHNIzuPzgLvbh5LrsWpnORsTtaLzM4N2C23zYH2d840idrFO6ROMVY2caH8HJNYKA7OeXGIFyK0Y
m0C/5Tj/xDOnpoGoDJfuvanTJkPS0EEUu5sSW8/qIVt1AQboJ8OmAn3hRVZRGi6P3XdPZTN6FWQ0
sb4XKQcKWB0nlLsMzh9Q+1du5klvvdh2HGUaOP1ePUL2QcIZrqagQcO8OOK3RJNaMBmuYG893lHO
FRmBcbAZaGJDXThjeHVJDyvmyWGTcqnW4ff9LsArJW6AF3SeDhS45q5K1Tp0teebAt+Q9W7SJ7L4
Rg71QcGlZ18qRr6ZZEdyoxb2ErLowyB5fcWJIH9QUvRcLkr/M2KhByGzv3pVLFg/CfmFiVErnzWm
a0zTCF82eAKQCy/aPZvF3pcSHuzyjEs8HiCd5QViNUWVgY4WsHYbYuYAl574qTwkedjj+EKEJJmA
4qFXtwjO3YzFv/jpn/c+EmJJKLDgoIGpjDclwvaFX6eplUtk1RZwMAHGvBD90Nhc5vNBQG1NNkKQ
8bMPnxWqno5mU5R+LDw0hp0GFbfm4GF4SGRmees2aO+HLzPDFqoQm/5/mplLH2bPqMJrpsKGw4a4
jVftm69kL9G+hKCgSliBTEA3oVR54mxombbutlARfEuLKVfzMi78XtkW+1AFsDQhaQ2AJgty7PL5
Lk4aacYsx4Nuvapi6IA0r0V/wDm9UPwtslFiPwilgM6Mad7cK9K7ViltzzQZbSDTvb1Th2/LB9zC
qjvf3b+xll/I+oVM/eCWtHWdtMHPOcxuVLhbEcuTDxayYYTGSZ6aEjKPVSN/6orHLozaOomrxaIj
2SpsXJjbQtyARxXEGDl7/3101DK5pFc2wPPGyyeLBW8MYiWeLEV1w+Xf/ybDlCYt6KpQejv/WZMc
va4btY2A9RnuBXYmMPPSZuIuQXnFt1q2yMg1qEiggpOLY2MA1gCXlNbLKbCn/zRM2bWPhkYiaQSM
B0CUaHI2h7Pfn1BB3igRKN60AP/w/8L8QugwWIb4L8kJAVdiJsNki6hZOPpBSpawMguY9Y6VQtH7
2eu1I1GGkM6hPVakRZ7pulih13Sn8bAdLljXO3HfO5q+RmmJZD2CKBaAfpxrWBZrbzB+tuApHl6l
S7/qMElQPNQTZhhouXyFjyrAumwAXkInXRSQTTNToGMDkZw6AE4nEnHXCJmtRS5mGkpjJcDCzi65
4EhcpGvJVqELCiEhr1qHV99x/P9rEcPS45vufQWaBfFO2ozRg6Qk7u8UPlEEV1OfmdQKV8MH0WZM
7AVnh23CqBluBuWlURzyRAsUvwO/x0mik3F9z2nRo3uthK0t9HS31+5ESm45/cDo22j3FrgpdFDI
MwGhVBvM9lcOv7+zg1oLuQBOwBQMncALBzXifn4xPQ4fF8tIJhFb4ld//+RWZIpbiieQsZd8mcAk
TkEEXg30a5biUVz/DMwgf4TmyyRu3sJ1/XS0KBJy+wdC8w9i8KGVsdnwLLytU9QK25nf29QO2fzZ
uDjgY0ht3BNMqC/vCK/goa2+xlwzhKPMIWLlI01bYawo4qgX9+hfXL9ZOhbHPD1T0sj8sCZaGEkz
qgMrFmN7yn4SiVnHER7CtpIDIuOrBaSnNM2lWWm+xtCiJizlER/Iz2PJ3B+ob7LZdjLPugm+DzcQ
jXe89adRlkB1nKwGW4qcL4dwwwahxKhtaP3QGLRaZ/acMZt51XCxLmmVrPsvutBkpXU2R+iFm+sr
tr6t2x7mOBXdotbuJQu96LahMq/x0++MBD30EmcLmYxZw/cZsD28GUpvv1buteWDHMS7wd+LjOfg
EAYuWu1GLU+Th/keJw8qbKGRK8E4HliEm7cE3J/0CwvuhLJCC7HHupn7h03ESQ8AoQyHHYyW/G/g
Y9sN0T8LJVZCY0Ned0f3BzdyAxd5CpkjrH4ogzAl+G2Uqt4dgKJ6UgQoZzIOjtz4HerAuy6YkID+
Ocun0UMmL2NLCnQfCK5slxRTZCfStWYwINsq8AE95kqu7/GzECSU8GMfa17bK6R3eepL4e7DkjK1
9sdrm4DNT1mOqaz81a+SQTOxg2GzaTtKS3fDnU66XIzTR1Me5XA3TyanF2XpU6FAIgSgg9o7UfHi
2UPjMIw4JG99V2joiW7RB7yEI1X+hDATcxv1MZIyLKUmteCdxpq0eiQyFY2VFzV7hh5dYRaNlkRK
EiIWfRESsaUOrSPqfl81jUSDAnJPahlDbpiZzQ1dIyT0GA1nno4bIdpsJz6zP4v/FJyXZ3Yw5B9+
8noYNPFhnXpKy0mFUd+QIoLIb+vs1cfOPQ8mtrUwS5edb//XIMWOChap42iBLM6jC9/c3+odf/K7
8UkACc4vrcOaTRB/FhYKhc2aSYLOAysOm7eQubBsudhhh2DpAUFqJgDoDyRwQ+VTTR44dbjhZsJ5
STfA5SdqrE9QulY4YKu/3SpZlhdy9IrCi+gWHoVzlGdwpj/NIvXLE89iNg/mHHkOJVCBUOG5W5Og
Msmymav33xEBjut0qrWGWJyeU+08NCrZZU9LJdaw78NMH6PLkcnlGJFO8Uf3B1zk0WlYw7N9mtnq
6wrs8KLkJsZD6LOPYywnkMoi1D99F0AhTqPSIJwVwEimHu5mzQ2BhRf1lNkZvn93mRcFCv1OpEVO
r7lrGHz6yj+GsQWmbSvRfyiBkD9cekK1rpzPva4DX0SwIZw2qCEGSWOLwH50BoWjThB+fs6SkVXH
PdYuR29VjC/QuqwkOJjEjOCnldkncyARwZiC0JBjc03Dq9NSje50fhBdLKWGBfJjkwtgULZoEGzR
KmNmvA4sEyb0Am7Y+z//tUMgHnj625iJIeMo9TatMkYMdOYeMCgviOsR+TrWrcpBRv3NGveNpSqh
SLTQLLu5aauoKcGvvqJJDJpZXVfk4n2i1DI6+/bor4vvRUNsXGEH1M+wCFZieJhTtzmeHvC677k/
SYX/c1nN7upYW4Fi8YMKvYORYi6jqX/E/mHWVyAlDNB6cz06woUzZRoctF/VcaAn25qsPGATU10Q
sIvdazweHVsSjFhz2+3cIxA19WoJpIzelIVMipiULwaxkmdsrErAh3v5ogZP+FZawW9mcWAgp8ZB
4kqKBIh4cSP3FhJ5MzgmC+KGHJVTdy7QzeWMC3Ro/ZxNhuuIFAiawLTkJgDq/nkBD9hilaVabnl4
ZlyVS9VI8jVTSOYvgyA4kbUyrxeyRKBAeqzo1rEIZZpcP9gNCMLrpORrvc9cEl407Fmt5eSKvE5q
HqmC5kBMNKvn+gPs7EEcCXB5rgXVsrVWWsFA5QW3Bu+6IbPoqwxOyfOVWiGfblgx8NuSU1njF4Tl
0WC6lyosywqJYkbnm1h1mrlkKtedGklZ5Em72bSlRotY+5/r77vKjRru4gFk/Oa1njXtfqhQP1zs
doI5dX3ipwBcnM8I/Pqd42sy/XTkjFK058HEg8ZHaYuTzKtUUbOyfUTapd5das/vGzvN7BoKOM/1
ejXFdG9lv8ilAAyZMPYPGcUO3psll29zmnMPT05hdrJAxnVynGi8GiHD4MAeFBloHn0jFB3xodoZ
vREHWT+Gogjm7Y7+KD25X9n1PgK1avlAQKznvBG1lLTiMV147/3+jnsw1a3/8eRU2GwkHmZjMPhN
4TdRnRkZ1dF0UECsQxDHWvk0BEwZGd7M3q0VROWuk4F19lw70NPYkXSNFUnxF4ES3UHSFuRXbdt3
uuQTAMl6aji3zJD3hm34aytzvPtfrqYIB/oIBw1Vi518Fs3vGbJf4PLOOz4jKWCt6VZKgB85XppJ
ORec7Jik8pPlKWp6aRbeSKNET8qwIOiRfiyORdCy58SBjd21yIJitZ8ZvOfk4YkkpCwGjEGT+4WW
Ga/TDS/vuZGV50YbG1gu9JB96Kj6jXEEXdFI87eBPSRnSa6/xRUjZxUtvhtwI+PflQ6EBy4ozNNh
sKt/LrrmIZn2Wvh6cL3FvrmjyUSoZcqLoqr7sZWqAgxP3LocP+7OrO5dAjD5Yy+9GwC4Lt05p+VK
8In6676ZOApV/PE2t/b2eRUoprsGje/r0YgZ/Ny9kRr65UKPREWPIZMUja6P43naiE/NobI7yIxw
dT1MdJbl6QR2uXs21Nd85BMo0V0X8Ko3GsGK7yXhXhHO9a+rZjcv//WaZLX1Pcz1xA52meVtjaN5
rj+NoC+pN1jj/yhrz7AbZylc/eAqfhdqkxe/nzdD6GczVTrIN33sUw7FJHILjFWWByBTnq30c5Ph
V/UzOsAvV9ja8OyBLiTQDxZuWlN3bdwH+hxPQSmfiAkkMFvB/4XULuVHAP2b6ZbY5/ykrZxhLFOF
xx0hXFKu0NlTyYAL8V5B3igH+tDVRAqMmNSLWK70X8tfWZHNMnSmbVHJgzeopan+GfDaKttHjWoF
7DV1kCJWDj+5AwmdINt+ww5dlTt1XywopM607h2qCe6KGkX8q/WSSFhAOQdWDF0kRoGc3r03atWk
278r3JWqmOQLDgtEc4vrQpFZBSWNVS4lxcCMZdUzHWV7IdjzDNhLkI6dhQabSf0+LUfyWn5LS0dP
hJRehzENo+xZyy52TJpGc374JfnxjenlvtzzfLTBtQsY5aM/vOd2ughgBelTZJGu70N8C966OyBD
IXmrNkCtJKoyoamysSdTvuHZ1V8w6w+3FSu96mYSA5ridqd/34Obt2wdgveXm2SY5LibW/pbEwK5
K0y/XgkT5n+vtyvT7nOqN2PR29UasMcbp28jPd7LcVr8A0JZRuBVHt9qJ5fA4WmlRUaMvbdVa39s
XND5KFyWLdnc/3v1OewDvld3JXf8ZwoawdOsfVUNB/DqyCjg0VF/Z2H8QqR3PjdM770WQhjezAt0
+UYn6MpVULsTMobLS28v1SKH+0UwXe4k31K+k2ojgmqrbCTuY/16s6VGziQAjNBt9lYa4KM5dCpb
Xqye3UzXSSQoxWRAZF66tVZrMKX1IvEgZC3ANBYJY9aBF++LoBoxbWHN/gCclipf1UlmkIKg01aF
BtrM3L22NbGgcfmh2P6GBDltglXWuKnFtUaGRZjQKnil51tGHj02gVzFhZkjLClTnmnHDF897zX2
TqtRYYPh59kVowkb7zWKKZ0KW1sgUTwM5GLvTqHqDdNpRIgQViH84Ox4OIdUudK2zktw2okbmdGL
hu2iz865NvQR5/MPO0PYpNyHngBF0eNVkOGqlZyx6jWPM4wc0AKuqx7XBJGT5zQfuthBGgXBrqa9
75NjXuILUNXaQ3utWqQ5yNOAQkHD0ncvZJJg38Dn7iiiUtek+HsU9RNa1eRHbjpzaNV9bxKst9XA
qnfhnowx94rQNZZjrkl4Nia2Qdk1JNavYTv2HtdUE1Qi9hoRedE7uTx17kJfUlcv5/hNSMlkL0Pj
fxqPw4AjYBtp6nZ7eGqaA2o0gvvMTF7E3tEEtwAJotkWUo/C18EP9t08HCnr2A95Ra0UKvFAreMq
dbDzhVZYpJhuw013DemoHTzVSNU7VLskLfaIizD09xfJ9t2hgE5hnujfLQpQVL0T0bhcoeD0MW5L
4/AQOFzQ0lR1X9mvSp+hZjmnIBD+DiUWBHlLdtplurQbpojnLaMUNQ3AE9sZFL3g5TqQgz0k+Efi
UhyvgfRGYzK75hXoq+Y+DGJsjMMOKA97QjxeaCcw18+0wynLmxViHQo7/WfebTa5/28VOeD/EZJV
kgjkQ6JdJlZq4jVGW8TYjakCS82Lx8zIavaqsTk+pmydSFftVQNn5GUPoq3JWgE0ZfaP10orrsmn
LpIYgyVUVEnKQLmJ1Vtz0By8j1m5z4Wup3gSarl4yMUgS5UDl6WVijBgP06ptrTGE52lb3QtI9WI
nXzqMlTTVD0JOZW+xD/OaoZ48Mj5j7idJmEHuybjWxnYh1LGRjCcM3pS4CWIFDlFmj33D2aT+SdP
eQmS8vKeI4yY54E/gstWp2dWbydidl/yx/1n95TYkGi3CYyF4tuwKr/0YVTSmFbOjCLHIsP1zocp
Vkknb/M1t289Z43FYI37sVaqr3AAziXJEm39jCY0sLtcKb+Smrs05VyDsPm0u0lNpsOwzAZjA24l
WljhC5/pEN4cG+ADua9zg9mePQwzzy4eUixVAK5B0zXW1hQRRauy2jUPow3Rlf/2EEUar3n4XWUO
PcApKf9KV4Ca8a21hZF9lx+qb3DzFZc14g/UfzdpTSDPz0GcKzPmvSK0Qfmw5SU7VX4Ao6/9mn63
oxzXOq48rfqb0RXQpT5SAM56aHFoOfKiByocZnfrzlcQcCxPY+k8rWvv3bxvfhuKUQv0XltF7uJ/
DUA/3pu6dJcccssZIYMtsmlJeZCqyrD3YtOXf2EVCUr4P7zETCd6Uv0e1uhmHaSvnDvNppQIhLDq
7tacwnpRiqfZJU+u03zclXl5kgPaDO/Q+AsROVl9yIcdbZGhQ1+ex/hvnsZtqXGVtT3hhF+PMVpH
UiP0lK4TCOL/OZttjk5k/b/zOeC9f1n93S97qWDtm2/fUWTA1TeNEaTWlMAfqX5I6kLDvKecstn8
7kiVeX4D5Iv3mtkCyKdUtn9B1Y/eWZiIV6cnx7tuYWb+TdBbkA9MzFus4Fp5BwFBoBZUMUBY/rKK
nQWZS8UxbvPE+bq9gJUsB5loxQ8cYeCA0JGY8Gkyp2uLEEY4R6BnroST2hwEdf+pde85HmBxDvU6
+Hvl6I4TlgNMQ7PaER2S2Lh3Bp6vogWai4GU/o9ZzMsUhZ47anFwg83khBWUJeiDcw8WkwJTix9F
zx90w5z8Nm9mQzIU/td9CYdR6UKpafZrw+GICrJjPQwJrTB2z1taHRRGyyxe2epnEzUwc63P5+q9
KqTtV/THBlJFEvLhHVuGzY1gpqqzlGdX2KTFUDVZ1OlbQlb+zHg/cs9zfjGz+QbqcAVEjCFyvbAq
+kqffc/sPKOaCLzJH+UZ8DCJT/SV7MJVYoDOs8o+bdXKgPr7ADMp1mm4JHLojhl6RIDj9jRWy7QR
OMlWa4OmjVXH6Ao7V4IlNvCHcGAsCR7cpiKqai24/RxqTfm3Y47W4aRJ7VFRRdc2wIJMlzlZehGG
UEBtb0ooeBv2pB5NjhnDoiT0GPBzPb8tKWgqh+WLUitnCFIqmmI61EtZwDTGKXeoWJsA9o5VLrW/
WzIBxegbXlSlb55dqH/ewydxCWxZjQyTk96z6JscAzIefOCrtsvCxt3wRMyAwWokbGYpab5jT8Nq
novNNlEbEHmL01B03pf1ofdd2e1Y/S3Sv1mjalGkjz3pPf6LXV1tSgX4GA5RT2JwPaM1G+BBw2ka
xSl+2tpBSgG8Ged40RJohOmHfLfPU5L5LG2QC/9A8FimFRdXnZmfd9vxSfVA6c1reIOATq+aLGNL
mbWRwAWG2pHBC/Dy+lS2tHEqr4ewVVkbzOraazABvc/Glo8o0C9EyYFAWbrdnOMQURjdueNBV0O+
zs5oP0XxpFBrxudnRUSzbxbR1euQBXQZrSHPYYPaL8V9ZNiMnMsft5m1Vm2JEYoVzk5WwWw+ceok
cf25wz46v5p6JNSq4L0074WlnTohQ4Wa9sPB9GB0xV2J1D1d/YREuJl6ay6i3EGsLFXsiiQbWdSc
zo1i/op3pl9xflAqMvQxKvcfgNXPuFPLmMfXmpGZ9uA7HmvoUQ7XXR0ieYnlllJfbG78hSMFh5jv
DXYbJMmq+YCFLXrvNxADFwSOIC3YMVr5GqXmXLvYMlRtrV4Ju/IY7WjQ9AVT5+XohM32lNFclvT+
QGsPJKFS/yIUg6OQRJ8OPl7DL3VGpFcp9Z/EKE7n0ReMKwU89aPuxW2FY8RmyMyL0KATMf9D/MJV
0Yhd6+TZeSdyUNk5ew/nhUBfD1CCYWcb0caREeH2r9GQ87mvZA8Z6WUop4LCi4s1qjVQoo5eLkwX
1zwYHOMGM5TDPitMzH8uWyqGbAzguG/ox+OeKrxsFSq8oPMD5TPHxF67MD/QbcFeng3V35PNFmoC
L06uY0OqyZb334Qe39Ip82O+9SjR9G9ieipsE4gBBTFk+e9wV1oXNfEqoi97BIohRRixENmf2MBY
QlV21XBoCH4IxhUiwtGOcT1WiZhufgSXkaD1HoVvPb4qhnZkqYYAmIhutTxOa4nsvqPiQb7Nm3wB
av0PeS3Bv7ijsQztr3Ie5IYm0xTjNCfGrByU6e7PR+4j/J7H3AftVUONWrVmCwAR3ipguWDSApBK
HbCq5NtukK/fU1NCvhi1gEFInXQHPp1sXXjvKB+w2GhqSioSGLmKm97pU8c6SaY4cVP/41lV/cbF
+p1Di/uNbrqMM8ZCWfuQAj75Xw1559bqQkrH6mirHAhpFHOPkIVa7O+/fBsejk/QiD51ow5/zCNi
QSy5+qWZ8Ti4E8MsB2DfxRFypGskrbWLVP/PX8xX0XKzFiLj/ZJRAd1uBR8N/iYU0KvXwyZXcCBk
2WvD8toKNfBupKlhQRj6HDK7VcIPAfl250pn5AyX4pQBbntXToRY88pO2sm8o2Awe7slMf0AaObk
+rTWgmqDmuSJl8z9ywJoKCLRe3fphzJy7rtKHV9Tbqy49iPQJZnmld5PKmEYZ+OxEoTpFcld7LaI
+vb7tz+3q2x67C4kYBA+EkcIrfQNoBcDqndtRmhnfkxkbzOXkRX51n2FPwSAAOBZO6xHZwwvO+Zy
+QpDPjO09vc2K8FpleFuH4gt99f9wsEPZpaieHVGnGAnEGJ0jQ2RdY8oW3KKft9xBEZmWEDW6gHe
xCrXf8II4ERIktUpzJAO9xx9uqfnbFyAF7t9Vl0+6OpPeEtXOqPkDIcCMib/mkEcgv8RC/pOWWbr
jvB8/VEFMFnHYGw/6W9xs4gBWzZDqX7m7oxYuvrsXGDhol2Ix76qqalM9p4E1MM9Sg8Ri+gG+zsD
+eUi/peDjKvKZTmpnBUmBf0Ld38MfCnQZh9TtFwYrXPBCWtaG/Ftq9fZCBPwoljUgCqUImQCXAOY
lR3QqTnjJZdo2aV7Y5EuQKtEBXr0mBF0E+bCjBR4ypPQLsdRfSszs89dPJKtixtAst/lIjd6/JNp
sQZ6TT+UdOEOvfK4PgJ9UhpaXWNNga6CVOWHZ6MfxflPcPT0TuWQWAEfe1cc+1qEExldhhUxSX+Q
VWcQif3Q2krGLwd3zYFZH2u6s/gm59fQbEt5KeKAI14kYusk3nC2vVFroEtQ/O8CAi/MgcM83URi
+xORwRnes/lmuflZTDDp+XwtHZd+DWemVrKW9jIiAoQHAVJuqRaXqyPxQrD0eR0lwsT0MKkfxzaq
iweNsoFHMFMSQn3lARFS8TTJSBBOwiMNwlroKZ8j7SUq1NyBq9bGzx/817j7U/rj9t4DesGSxg7S
FxxPHXXrOHUexIvgiRgq+DCuHEMJTwkwZsU01Sr78luSJigWoGeA9fdGhGptX/3HfMqgnivYMfV0
Msxg5f+mjSlNAH2kg7na75SDmnLQS6A8cZAXbDHXnnGMoPyApTSW4vAEc5/Ask/9eeAhr9CUeDMP
lCywPUFqer9lGeIQ2ZGas6T6F4hIjmWVi/fei9kUXv2jEawpU5VtfdO1KzXmTwVLpMpQ56U/eY7e
VlSM0lw6r1c9XTw+AQbzDDDAGwgYbv3pGX83kKoccWQUYxSG2hbovZvDZEBWippveUAHz8CiyA35
fcn8HkDmkxcy6m441gEdnXGBT2gIbHYymdDXO60dyRF5KueupCN6AQHyNVs2dS8fJMzWTPDSDvCd
++1BQe2huAWHOlhhazKI2aPsJXEbKo0hhwtd0gl4ZE3tp9Ljb2E7aHUxX758acG23T1X2KADFyyu
aNvn8GqYG3solxC7V8Fs5su5/UUwrDfBKOV9frKCGVw8TMWvoinO4k7kI48BXxx0hKh4Ccv82yKC
o6EFSPjXUVOaWwtLPv0TR/z4QNn4QAlGDkS22aZxyh5Bgch3TF9hcLQlWXraJ2o0JpLfIc++onEL
FblGy+mqc6gFsLydJw2Ku3cTnuqJvHZCGBPuSrU+VfEpuoMbBTEiGdus5jfGaHbySS0Qqe8nh9q0
EnBlHhry1P4k8CqB07z+qqXQLcS6lFzjcXWkFvU7FdhWCRgrC/WnmpQcJxxWrUHBFBSvdv4vAaqY
xDNPe5yXRuEbcQeopxD7uS0RSTK0tNSplWf/AnX1/ln9loGrfqgywaWprp/uqxaoKjcR5R60DzFR
Ssd1tIkRqwNgWbmise7tNmhKib3svdy3CdOFdNxs2JYnqFVUnawcJrLj3HkekcEAeSFCJqAG4ni4
//EhMu0Y7ugbu15U3ScTnzLQwu3qKCeLiaouKfg5F8kkx0VszLd5g0b6uDAHJYpgBx8dWFqWvGjv
ld4jQd2yTbBbUsu6/5QKtZdoCs81j3ZBI9EemyF2/z+fayX44A9mSq2dfmBYsf3ydKzcObucUsvg
sSGW2aW43ohvmZCjXrn/llQNfVXJJS4QJlD6r1z474IdB5KAmar2fKOEEOKT1ny0eFK/GsvFAKr8
YK8+m/anY3n8VcoS6q0ZEiyGR5sZfKFALyBU/fqovKeGKIjLlFycoezdkJUyT+c24j5WzdqAstyM
3Bk1GZHGBQxzlzp7Y6XXUq0rpkgrFPwq7utOLzOpGaL62+2b3usiuvDuX5I1gueN74HBZJC+7wiT
k3fsExNoDEknnKR/seE05HrAaXaeXfIZOtLmMubtgPnldiK4X6Zs7M/2Rr13+E+UDUOPefASqAht
t1xR8EUCFzG7H0rDE0RcRGTL+vJM95cIasqNFHV9lEz1VA8fHtZ5j4OB5vhLhY/uu3pLFgrpPlzS
EcM9sFfG5uX+lKUFHo7PbUtnQkBPkpHnfJ+j00K3Ra/9e6BH8khCXQ8vfqwYZQxWOaI8CS66Cp2l
LYD90sEbZI4kr7bp/r8/hWRszX6qk5UzFNISLagHiXW0nSdjH/zwLbXFeh7ClENQ4jZQJdC1SAX0
+bffw/kD5/n2PixdyLwvKYcP6n8Z32kO6WOJVLOoAm44ZolZGXc7l6ArlDlewEdpSE4as1v4oirs
Pr/MUNXYvkiLoleB093jVWGmMDETXd+X8mVaBKNFXJLWxWbUDXpobHw5Tg3Q2bvD37EtI1W24U61
U9zQHt3YaceoBAn4NQX1h1J+SPSgyEZ4zowLgI7O57ARRCINB7f1ginATr1UA0o2SbVz+W43z+CZ
G/M+4wxG0yUNVJdAxvsZx0MWf54P7zAEMz6X/yR3CePcSGHA8uS7cbQqocxphckEERJs2MKyKpuw
471k/f315K7/Ka8Ja1wwLogyeIJ9fjPgVCzz9GxlAZosNzeW8zGNGc1n3fJcuKruR2ShiT+dauXV
mjtc317VlZ++cxqQWB99wxVmT1bR9gd6Kwhe5fzFxTA3X3NBNaNO5Fa/Z0cIpHWnKkRJFQIQIWmz
IfTE8babS2Fi6YXdCBHK4ZWp0kQZ43KTnuFQAI5rmrNlu/M6U9r+QC1Fegd8jLdlhMicXh2vSJBE
3qxM6uFgAp7Re9cUAy6MwX45LxXZE/oReS3GtvNFQXYVKqqac1HG8n72wQK7RSTEoDNREx21i0Es
r+n0oAXWgI3WqD7Q0M5h9MH8UVwP1/CeFJj3YLGLnGMGMjR3oSxQvy4avvuj3LdlPjk2qAQc6lwf
ftntWfqyQDd0xhuwGYIehIndVY6uwzhC/chovgWwrBZ0qL+iYjV0P59yZz2JjOfAC5xo1ZTwwxY6
FEAz1BiZe+A7H4YTYdDLgEPaDJi10G1v3Ob68Sdg06QICbWqcREIsLrdvy+bZaytia9Y/9DASvIy
SRLShGUgBOLR4CkMZun7IZNcovc5+Pv3gxCj3WpxMSUt9Twmo+j8k3ensbvObZAEmxlPKPuNNUQY
lKCM+idGwXBLa1iAIHTMzrNWKG11dtTkYF8p/s/2PomIv9GgdWW/U13kEsRE24B6yZ4aeSysYjGv
7WKgpjMNsTnPCNOVsTDA1oSJggAOux8Fgy233/xfzXEMbD8bva/+QScxhTV1sQYsRlPM+6M6DpRi
Rzs9K6v4rk79buzl9h7hKGSMr86AeM5gqDZyvMRzhlR7VkYo3qfOpQNS+2hCCL/hAfReSFLneut2
QB5RRUJGzvWfnY6GXfys/vnIW3bVjQkaQxfTOYpcniymOq6GKSAUSX81NphBQUqo5nKOkkmuVDmi
2LWM+FKawTAOaw+spxw6QrXuai8DRw6o0PJYtj+9H1e1f5L1A1i6UH8hr74D5uO8GhpjLwi/osd/
t2rkQBbaMjvuP6Fv/UlpuJdaxZIkmB/SMOeLXU2JqtjiInnVanj1DFMb+Dz1HZ17fPNuNKHY/Hp9
fLLZRiMLHnyc7NbSqnYY5PcweK0+avjDh79llv8DMCg7jO3IXBR/DSuqSzbpHehQDqFNAyB18LgW
VvhQoJpiz9A2As9i5wlHjeQ0AoV9+gcTatleppjkBc4NeyzELQalvfFYdTroo6Aa2ppZs+MiG7bz
FkYygT0rpB2AIPoM7bg6OBwckBuxGseBDiIT/W2PON6pAt/MOcRE1AxBxnwTUxMerLsLwG792vYo
0uT6evhHT0gBE7pjccH6bUZvHZvHez9MM27UTMClEPYY0a2cEoS9u0lxUj88AJv5FHLiGkV2tbLm
bau7VXNdiCFCCyrf+0Uif09i0Q2s2Liow4T9VXEN/CeaAoWP4yTnl+LE3Ewe22RNi8cuy7tyzoBz
coz7sMhlq/tNu+0Hd6fsVXcaAbnCU2U4EGcHQHQERfiMB0uPkJTVmTK0M8YrhtUFMD9TOBIfHpr9
7nhWsjmiSUpfA7g8QD26tfw5DftvL5nDFe4tby1bHt6oY93HJK5hSPmdDYLBbTJljAggVN8sfSmC
ByUyQ5Wab3NyvHM7BKZpkdSEp44peKVv/YVTdp6EU7x0zhUbNkXm44+MPyxV4vMwr0qt82WdsXfw
BBAfvwQWJ/TnLOtzTqBu39CyuF8oz5nF/jr9frufvyRO7B3BnDgTwnZiD5ss+qtCYe51L13qTRmm
S+VCoUtWVH8GQNsaGdJKZKGjiW8YNJOQlgjMCHQEZC0190IqrZS+1vfDDSm2jWGv2A/vfUD3mvS5
uT3dnCgoFghuuseQpbCD9W9kkxYDNmHZYjM7olzup60pDU7I2gK2jlC3D3u4ujE0gRdqIh+HP/cr
GFtMhHi4hoc3JymjKNdl7FFq4KrqYIoK7tHzNgOanWl70hEuf0ROSA8r4w2ivcmZ5g1zBh/NZDS9
/11XmvM8Rds30b52NS1GJsZ9NnPSPMSEmvgOoB7mw6AWB6FUpx4shZ/hWPAMlIeiWcRtRgPswvth
5ieUB0+au4Vhy5BhHOIMfcWdNNfNx+VWz300K9sX66NNyO7apEa4pxQgq9pO8gQ0CN8ahaEfO3BP
WzGC+yaHDYTAf+nOwU7srFo14yLY7bBRY65F5m0HUJj0NHhHYcddxscA8Fd6XqD5MTMi8VIz0JNC
hBDemPxlr4yLDJw8hrwljEvDeCwH4X70kz417k/b15xYQufvY9atytEf1ClsvFYdwfMDXFLq90bi
1QPOe/Pg9Tq6gpNg/8ZN8s1rK4yRhG8BOmeCRBGzcZXyJfH5Zq+ePs+H5lbxi8AHvSzDdDxE04gA
phDRMePBdAOhj+CPMlg6zsTVcr4ztZiF7HMnO483W58e60fnm1umiy3QEy5CfPbFyXsSFx/uA3o2
MwEENgIuzWnvRYbhH+Uef8o1K/umRYZMsER9uWQrGCvJwRTWxLTL9DZF3W9TXHuoGeMoJ1Kt8bcv
BNmSCXEmMMgHyXuBs0CE8ZMu8CIu57kG6a0hxr1C/071UCXs7J/bkN9NHyjEMj2bszgBuPkFLc/g
ivoUW60DpFAHNJ2K1Ie/CepXAKmKzz3x6vlLN0xyyA2Vamz+Sk7KeFsTSK9aT+EsnyBtWAxyjYnN
M780wHHT4gGxZOV3fVz+z7Y/JYEtlIAna01RmgtJCTDPpFSlqE5FAW7m6eSU+zLbx3YU1gFrQe0X
nQJnQleU8fzdkgR92Nlvmuz2BXx7y/FZbYM5S32pEzp0nKiKEGTZIAai2FpV6VyrFoFGJ7ZqPrCY
+hjvnaw87eCKEIZgdqssf2GahrftpVD4LR4NasgKO3Wykex/BPhtyKmTv3MnKugCQoax2xIywORm
zFSAuWyFkxk9jjLJ08RYB2sE5fpht49hfkLa6oFc9v7RopkwAhRRD4lt1qNmZXoFLxkrYWu6+MFA
dFWiPDgiR2l24HlilXdzOmcUN56Dy0pAwMCmF3vHZOJZJv43SsuJpPfq9ChQYzws/CyeqVV+z7BV
4lWJ3TRUEPYhVKsPPaN7EUN69KufdV8ZZC190jGa1XviCKzo5qkIdYEp4yJOWAQ1dwAFuLBal4P0
sNcxCUki5fJ215evZYEiH1DdIYk0cOJMy7T+LyAgXeST3bQM7OEzAG2g4/ffatjxuZ4ceul0Y3D7
G/u7rZw2KAeYCC7QVShcJ1988BqR7B1XpLJh4OHI4O5t9UYYX5mhlJQvnB5tF4MEAIUuFZo6WQMc
JAfvEJgYeiyWfIS6UQZflLY+jL++tf5JOK8ciogzEYpBvnsYos6tsxy66ZWh4s7nWweDMhXkBErz
4nplO3AI57sc67VHPrme4tkwz1XqUkpp5ST+hnVbVhQI7szVaCCPl3A2IyuSmJeozpotbeyeyx2y
YsmnvXJLV7v7lBOF8OExKVkySdO/ymL7kOmM/8J2iiTp0FZtemmBOs/nicpywAVWJOo0JzjpTd1r
YVnb4RGaAxHbhuvan1rJa186StF8Im0BzrcceEhfPl7heO8qrxev/6VRk/+ZLCVm2Pkou8El3MIJ
vwfE8Qxv6SJxNj/te6iJF/w6lrY6Ywc1SHf89v5FsyThCkDkBvNhPy/ljJ7BCkzCEoSWgcnXh1tf
wpCVBBGX/h0orzw6zEp5xy2DRN96Q/HifJ1wgCN1FttfJv63tEXwMsbqXylehHpbTW3fNKF6fmKM
h9JrwmkKZ5Jj/Qk0AwdXQpi47FLnRM3rl6tvPZ90rRO7Z6WheDjMnzUHFKqyaBAlXHes2TVnAcNm
a1yPHyKW1I1YS6uO3S7VskeJlnIu+GTq276SrW1JiLbMFT2IYVZIjvDFEp1RzmKcU2phyjv7fcKR
wqk63OqFAwXmxiuT0aNhImFgGHEujDgGM3SnaACmmp/i1WGG5x70CrR2Y9tJUst+zq2LT1AM92HU
Mwn8/3w1e2uoYWGxLWftulxb4yd+tcwRTkY4RkdF4DzeVZaKx0Knto81m45RudXuUOTlm6c3OKQw
Eg9MVgXo1DvCpoYA4SE740wj7kw+J4Zp9vjJg9HCHj7LI8Ng/6ZeyxnDHsOiGcV+7nynbTeVRs39
L0R0Mg09IzJigiAr0khqK1PQ+65/J55iCXqqDhnZgdet8Fxg6z9nzut4cS/QqjgKIDvRmt4bei2Q
Dg9N9MbtB4VYbNWV38jCY3kO4GIIZanXuu/eBM2E5hLwEB4hhPKjq7ZLzE4lmn2D2RjuMKMIssrh
sOqUz5Pj9Th62ZJmvIgktTBe7Tor20DN4vvAidAgVQMh+2w7l8f58l6ChOnPndtmgLO58fpTlNRj
ZID2lIfYz9peaf/dr9Dffl5NvZUiGlg/PzqXVpKLwm62DBr5/TT6/dywEEXFs1we87DaZmvERZSZ
1USaT/RWIKvWQFzx6wDdsYDX5OIbLdbbGyni4t3Gs91NltN20HnjlYGjXPv04/BBehLy5ZTB5jHh
56O6C5c6IuyXdqBhS5mEhbPs5NcilKdBb6GAIaOv59PMujKu03UvtC8Y9zu+2t4zld/T8R8rLw/z
wOFp2t2Jd0Wmk4y2so4GERTZQSqdMFOySdvq/KTMl6fo7i69mmbn2qt3Zyg3LTACxA2BMO5aD4l5
HCIAaKpcgSjlgpQZYsjpHHPNnFFNegavCqaE4/t4T/i8UnSN3sVQylevy8QSTjWug44kEKPDJd2j
v6+oM3veURzMXSlLwGvtfh9qUtvou1yl0xXfZO3O8rgWXUR4CslDOjIBF5HOYqyT1MsxpAiVRKtd
zwx+yQc5wfGH7d440HrUAURTegdrytUOQVRFuVUbiChaDfG8k++jQOkygANkwro8P+L47Wbilg3u
3+G2RkOH9/QBzC66bjKKJ/vA1vZxRKlck3nM4OqyeTfzkPGcc0gmpVS13wCVxIerbCDsCv46o2JJ
Sp/P6xBpaWJXYtYbWbLm+YKVzz0SVzb/Kc6m79BR/6jflPL84cYtAxlflPp6uUmbeJdosQyjG0Sx
MGH04tl5/1+eAzN3m670gSn2vgw64KGQjEP9rLRlq/V2VAcCxUXgexvHBzMPQuVUeo1HIYBjVzxm
OTJ+EpzuQd8RG3v8WgVHPaHqXC9wT7BFdOSJH3N7i4VnEZN+5OMNyE38CSsggh75i3ixESpx0/b4
mt4jo4cpoPoUAWsehVx7cy5311SHhHbiarVM0cLrzXSkmNZRzHvbLSsHnHgGos0Og68LMVwrKQQ+
8B6Y9gSo8AiDYZpEH5AwcsoPm7EvYOzv10YnvwGB0b/geFM9dRuImfnXfLeTT2/pWkPgsUUdfdSO
ENJ8xysF1ALCWHtXKHpIFCfOeQ24gxlywnkhxASAMOG8rBu+WN2qqggAzBIqVA9qRjfGc0q08vtV
mgpX0GXUgke9BnSiwbXzQu82hnK3sd/FoL3vtweTexTT0MB+pI2HBVKrGbrNHLHlq/tIxYFV6QZt
oyoHpKdH9DqraxLu/XmhrL7/flYPRcA5P2PFhlfV64oIcIZ8b/b9Xw9oKt30OR0ZHudq6hzZmmFC
vvcJ2sVy/l+ybKN/wyZiyCXfOQXjFmNklxZDdgfqmyo8SPuhHj7wozRGpvBYz8tDBBPcyM8jYYcl
zR2b3X2z0b8RyMPO4dRUqR3Y9zq4zuOd+4ua7XKrFtLJLuFk3javkxhnDV06VrUayc7U1bWnx+yY
Zh7E9/XZVaWbTFmwEtExm1IR1TOIZGczFWkhEoBHxQ3xYIXruWan3KpL5H6JhnqY+JOETV9k52qB
FL6vKGr8kvSr5XCeEAk+C4U8dkF+N//SgwdG1u+nCe2Vwtgy8y7JkHvD6+l+Hnk1TzTTKme0pmUb
qhY4cmJ1mBOeIdrju+J7CaxFVJX1meeJTMQp7p1w58UYMgNUaYagkhZ+mu5gFazY7MuwCkV2yHCZ
Neyl8sf+ZPkevtI/vZTz/qc2Zp+fdrqz434WQ+vCcaLh2z7ARAqY48HHX3iiClZIi/fbyZmqPjbi
D5wDHCC8ovXv45r3tHCmvRKHHsDtm4LwW3/IRv0u8odfe4ObYQj3nsPlRT7DkqO35ZP1WJ4CYHgS
qocazrV/loaeZY6DAhJesgk8+WiAIaERJJm+HiatjxN8YI+ReD/GbNkJ//4bGjOF62FRnZFj5t17
Pz5uuE2GdzTAkUQh6cL9VcRn/gX71mwaG+Hnh5EIvNcSPy37zTdJ86P0dx7OTOE/XfeL744KQxCK
yy1Up2yGiHUh48q3ghFwI9Kb211dOj1ZH3hCxs9xjGmVtNuErQ6pT5t38phOOt5gBS6sxunvJM50
6IXvkXsek58FSpxGGMAegoAFS6Hv3UZIR4kyXtdbcoiMVlJXTiP3QB4c/rXTv8H+GghL7/ypfexE
UUGLLfr6jU9f/6qV9haZbjCUPMA5/cwIrusLGHdlH5yG7crupErPPmfRqxh3tg+i/jkN0Sy7FdV3
Bp28ev7snG4tQWiTw5dspze/A06hbZB56TnVhstkhKDfOgR4GfEArW2O6LwNjkZ0cGQNkZ5Ya1C+
fw7HpSFlCqJH7KPs5AJjkXweVbGh5zbKfca//fJNUd2scfnPGDX+GmdpQKmzbemoVK1zmSUa5ggo
qlNzepwCsJviVkUOIDmHYkozptyHZ6bp5v/kCFNT07Saupd8fv0uBj8IgLe3qjtVACavXNjea9bz
q/casM4FxWMLOTmiLQIVhZT7h9hsIMyuGNnjurXAhwwnawE+H3DMVzahJ6xHPWQw+grTAJwgWVC3
DdcAzXIoUEl9PLUxG4+TVu3IoBgRzCxuhWpfc/U8fm6W/+18d8k1SQeVPZ7/IM2Tci4Gw6x/z0tR
HJQUOpiSQWTqsF2Qk7nXTNrVZZL7GJtZ3qNK8Dfhnvu3IS69yB0YEHGKw/mmqEbHHOnlBzVD4eGK
SYvAiBxoiJKmW+1AQzp1qtWiw2zzYI2jbJPiBmdl5ZATAzY7hqiAeqeckcFwmJUelLtrYWQI7cl7
Ng+bKyd6qukvHZSEtYBvpbkk8nLlA4MWn/4LA0iaOyv0biyvL9MWzKCPqbPqoik+ajAVH1Q7Vs9U
Fh+96PB+/oMigGiwz4XSRub3lzeWfQxneTt/uJfIln5EE7197ooHbk8FKJ22aNrfNSkND4gufbKT
Cpg0yAgh73bZ2AxDLqbrkoNfsh3nXoYAOvJopF7hMyVgoaG+g7r/rYzprSUPQEaVU2vEueNZ9foy
PyKi4rNbzPKBu2kjlg94EKclB6ufJSzOWPdJser9TcPOf/WgyY1Di/MNL91+/2IjYVKxows2ZyiM
KAtRD0dyK7LtOx2bZMlSB/lO6jhjh1ppRB+kuROJhbVOvGA1/fV8n0KVrMw+eTG7kctDKIIkvmTs
KVXPBeQJBJNg+rTrLu61WIuaNrB9q9vGFbt2usV9+4iuFFtwx/qwgLwCeIoHRoEK72lWyatInKjZ
C0fwC9F3vUEB0WL5MnCDMwt6U5xCXdHgZdtHcEcqGhp0SnhB5nzWvWOS+M1lHw0ZbRn0x03+d9UE
t/EFpXKWO1q0B87RccwcLBkOfNkYJgI0GMZHwZn5R9NT4BJtvPjOyg9IQhbILlNj53cPo0SBlToZ
59Hp7LRv/zXNlxqOxkFSEtHWTafQmOWIj3GxxomZicmhFVC4xYg2T/Cfn510ISFaA2OTnK3Do5KU
idahW7rpH29qP8aK8onbpQFYHlQumVL5kbyl2oPoj8cHzhUltf1sVEOxqeMmrS3OeGWMKnhkI9k2
xXXI7IEZPbSEiuZUfJ2n9JHA41Sho7KNssfW/jMdT2WAPimS6ZBiEyin5IPpdG4eNA6NNhkGNHr4
SpHxEZUJoVr2IRGa0u42GfUYkTJA3fA+/g8onFCL8OExWAyoKtIXPovb8gDiRmoYnP1ME/Gmyvoz
fvqIzSrPtSDII0AbLPkc8c8RlRO3i/PsgoM/2yUUo8mx2idxMcGmWltGS+WjzQcuVpSo+y7jMQHM
ueZvD5TH++x6qlyxRvEqjEcV0k/ZiNW82+62g5KAReXL8Zz9WH0yVsdNq5Pv9DhoA+hBRMEo/v07
yWaucaenRT47u3e2mRDucCyYSTLsx06lhc/LGkfT2kbO96zAPTZsantNScXk5Psj1dqYjDgRn1NK
JZZuTv3oHz3DPXwlrKWsWCLGGw/BU3VfMkdocxU85jtw0494Ixz9avWOe6ApyxChMRahRgQqKLAh
06bdcdfacyZ5T65j/ONKt1I1G3BfYNT4goQNODZT4RsSB9wFUPkzU8fFC1SR8qO7mAUqGoSvlCkN
Kh4LeZaa6siCcut9ERwMVHeXxz5nFF8YwPWYbzT+hldWkod7WoU+eR4520x+iDA4jFUnSOfiYbuO
fvWJ/dm8/8Jto0g4YL4AKxxnR9sCZaEHR/D3+QkVEqX0IZwxgRQBW98pEhnOovvfU+Rxdfb3lRqq
aqB30DNgwJe//dUH/K23c3z/rLmye2jACNAr/2pvJV5iVCC43HhGb+Y07nArj0c0JitchgONQ3uW
+ibn0HVhfZbTvCn5cMbY5lD30HIR/L1Owuo3JdwHzeNUtW5aw56818TQng8T9wXdWQNXcq30NN5X
8PJJK+QNN/W63y53GeWzsSadoZYVqFj5QJHQ7qpmpj6VGetG0Zrhv2oDGWqMK9DjkEJCO33UUwPr
FsqRj7oVbluAx4wQosPFGPgH3WrQ1oIhNeHw5rZIYvpVN+FBIbUEUPwl5tlfxka1IT9AJ+Ca6bzm
FhMv+Us92PpXd4vJ5ETIIOTxVmkT+2oc6wRY6wXKpeyhHdEInNlXsiqh5B+ua2/kFWQkF2CSFc9H
A7OvE0bbAs+89X+0NJLy+p4ZS+tpHbv+Bjf94tYJUGwTKr1zq5GlMqIcIlgzIsFkdbrk+7WLcYd7
lC1rLj7rKvHJuo5difjqa5eKXgA1AC8Vhn+RRFTqU6zSWvRCFu8Gxcu/gHCD+EyJpYBpbO/BE7z4
wsMc3PsXMnnhwo713meofB0IT3s9iefU5CHG7o/WeVRdvFiFZ4JNS1nlWMg6WVjFuj8sAGOZlSt2
kHjJGjiqcC+8rbePmZcvWYktLTIvQEXuSOYqZfVYx6IPhqJMzOKvcBjwvrr6hKT89quznSRnSAuh
Q2kpg/kZT5yFl1s/56n2KWvD7+5pLx2+L0WHw7GlMu/7NNLEn/goq3tGRBPgt3O6WOZERsopBAHL
yzbUWrGDI4FgKZQKukZx6UGITa0LAKb5N9NTfB+6OA+syctc1c1ZGGUlH4vGGDZgzc19k2IrRfTA
Xxmr9jD49sdJ7AKzLA9CWF6ZumsJiHzkw3SD3tvqvtwMvljcqwV1NQSozmcUIFGbEQphKak/tAyN
65S6WKoMwyl3TPd4vOPf3pOgVrlX1lCRGuQ9HCvy73eD5W2NmTauX47x3cf72MODH1V1arXCl1we
G/WlUXrB7pKKKKr89whYOJG6Twx0429uYV1vnuqR/PERxeQP7m/ANxvI+T4K+KaKs860gjOy2hDp
OzCmwMheWWIewKlJp/ETavBplEUvRPt4LTvoT0zzSvgyG9vlZ6lKnfCrHlUfl5VgzqC/b9MLthGe
FllAtseOOoe4EW0q3ylAKL+yApkKNtHBpyIRMZiwnkRAHxiKZD8C9IaM0vlj7nZzmlM6eJhhaPo1
9IKymvAgrZxheq++ggb5eug24J9NoauiBKJ74q4XdadQzJUliczsDJqiGldaTUIkWMM5SwrLxCUi
MRd3lDQTRKh0736Go4aaAXP0nnAa72as2+YZHbS7+AKAW35q17La3K+vW10mVJmcWoRRex31Afuv
ULzciZ2KYxdezvi2wsVeB7llf8gY8+tEK5o8F5hD2aMUi2DITYkgDTaNK4k7987Gn9cwyicA/8Xz
udef6kvRClvzqkJovN14Bkel/g/mXKyuexzXr1ltNjHFjTxoHdB0hEC0QyIN1gzW7q91GFFwZgnQ
EwEIDMaNo9Ax3KOK3k1hN1R1rFeNTzV+Z9h5tLHv7lDL1oLDVzVYkiyKAypUaY4Uts9jOPGx7YrG
dGUBOM64fU2dp6yVGAAHuoRNe7Nvt/zb8USnGrSBRUxRYIeRsdXwZBhBVOjdX7Eg1X4MQ4/ORcSw
w5xrkz1MPCNYeeUAVyXJ27EYE5dDdcGKHBY6kcL2IX4zzR+bW4dw03j7OMFtwBn0gs4uMB4nD5c7
+E5qP5AHlVHOhKVfObShi7zcrwY+zTaf3V3qSCOSWJ3WV48xF0PifqpBqIhrNO+6+x9E+XZTgUF2
CWrAWj8aowr4bhFO/vtd+1vuEmPEhu1dgmz96bfkBmZsHUx4527j9tV2DiLj6xJks1kqbSP+SHvd
NeZTMpbFCUCpTOSS+K/4uMinG+/Noql6fb2NKT9bKJfT4tOtJy+KlE0W10rXHE/2AWnBTpiHipCy
Z2QIZ1IPFjfqYM+nmcVwDuaQ5XzNSjA/OB4R22tU7Mqk1DQbumPX+bW7Ybje+UqCHjLlcYVqTp4y
KkuP7m7uIt8Y0ZtrL1WXQeKs9q3ZMrMyqXt+8+0ofaF36csbGQKYCCKkji0iJs5QvgK99pSkN7iv
lvMu4jkRq/zGCE3/f5Ut6ytLD6JT2mbV3huELEWR2dhX4XyQ8pAUUpyERIcJunXSUGyhDhZ6Eu3g
RPjC7zMtHlUZc/e9poTzXnBwiPZJaPQQsb8X9o+ur0xSO9yxA9jR4iAuRce/ew92WfpVpDWsABB2
gTOEIqWQClGhW/MLKnHK7oMepJgXZ6+0j5o6FU4QwsskDJp4m9+StgfctIyvCp10sTxQAGlJKqzv
lpmY7nHa2iIoitRqT743xf6gyQpeUMY1OFxEO1PST8o+ywp+hnLvRm3RjQXItgJRoyChPf7KJQoU
ftblErUdbIil7jxGwh4BS5nq9IcHAXZKHU2KGbmTbR1+sLqEoaFYfFt1a8IpRmcyTNlh25l+oxfn
xzDLIywjtqDwIK7TX76J4nEch58NVo6zuXB3qxFunX9syc1+az6S2FbfxXWu4nqESBtvd39V9xCQ
RltaoV+zAJ1TlPL81jzBNI5MsNcDKx//9OsIWnXXEqmNl/F3cdBJU1czqkSoId63KVRaBh6dFdtT
VFLZsWAsGtu2Wjoe3o6zesdn4e2qF6EVKcg0N+0cR6KdlI7ao3Wl2ZJm1cg/veOzImDQTbOWnQqZ
VO4vI0VKnYACGe+nZlN3kh37Jj7AqLDvqIAEusoywRPhajCUNdQVxK0PLsmj1BBClhrtoRtToUuX
qKME1w7kyoLIKZ6BRnRDBIyRhDPrTwdOBGJWAQdybHVbC6BRubbU43FNjI29XHmw6jTlikAIxDZN
oWPF+V1yX7Hyn9t9VMkfxbmqDluGEWPRj/mZyDPncBXS+bR8siaO0LIfq8rgR7fIWBIwqa4bjFXk
HxXULeXf0wQpXNImReCskjpqfmhH+nl6gNn+h0TGDxLC8qLCVfTHzxKv3+/By2TOX/rKM0YIrJ/G
MLTATPf3O3AMIuYrd4KpCD7zKD74En+cFbGIqT3waYp++tSDI1Zy5Dc08U8iGPy6MuT8MLOc5Bn/
YxfT4FqEIFrT2GFdSjxeWzr4NiJGjdySe+7SI+hD6jbZtnxuyOnvNUg9BiM2aMgQ8Gxga65Rma0E
CmX5KuqQ+kglAlqmdoa6y840AMl6AKCFNQ0KrvtI7i7UISFLT2NgwpXDgVUGCns07BTcto5hZJPR
VSFTzQPxFnEjDsIIu4k8/kzly6fnYo8qIKUvCXe8nbkUxQWnRTGAvZ99dEsmCDjW5dRxFrSxKRux
ajH6mc6fvJmzq0EwOFItTLPNxRbZRjwsPQborFKurNvIzOPB1Yx0rzzm0v4O3oBDNT2ZGrrbPT89
kjRDlOb8aC834+iv6lGIbQGFRhb6QYI9AJH2lF5SGeXCKwVL9a2hEl9NljTE3A6n/DYlFDbjzasl
prlesIdtqq1VEu1yY3gS8eQlvOYDMWdAUSpDTfag5m4getHZBMzKi5Ph9GufNEePA2qBYnLXlhtv
sOPooN6if+Y1rl6XX045lnl8mSmCenvMA3Vy+LihJAkdHSilOvDfziIF4gOgzhq5o7XP5S1d3Bhd
Q20o7+ckXFNK9QAPQgToEij2CZj1OgCztlwW3/DXNILg+uTPuvUJ3RL5ss6YYnC70OegWFCkGyoj
TxNJvXs+NN+MHBd7oBWBgwaMLyo72U8MtfitBpexXUrEI3Rsnb2CBazMCJwk5PoTt7Qfhn45hnio
Me+nzi2+x/ZS0XZo1SKMv8J0zxfhHbToWSHDuKxb7pMqP+FaQNJGEE8xFDwxntVy0NsTiGH2Ary9
gaP16b1Xxn55LLEw7TUVwCuuAeqmjwBmvmkrgCYx3tNoAAOrCIVMSoQ1py7YjYRLkuoqzLPsSW/N
iCapk+71FVIoEp8CpJQRKXWU1sCey8PbxkGKBmsO4xTj85QdCUWaOeO+NcIqys7tWCHODSiowiLT
T/CF/b5vZSH3wkfckEuL4o1D4nEFRLFE34hzEuHp+R6Gf1jjBSAh9oYGRJUXBXTagSVea4BmbGu1
fJ9Pg4sxdhUPj2xF5dFFrz7u3zgdKePAD9xk2B5OmBmeQIxlASy/SIa7acNXAHCT9F8TXiMJCdyi
tR6WMYopj714+nY6Vln0ApsIDBGyGB3t97KN8rUezidUXKCm2EDTCAZL9gEmP3/RHUC4nVLVrh39
R6fibVcdfKQksRKXpZRb9xUiuyvXAx9GhMIwlSwYbmVF4lirW8b/KBQ9s5wQf4J6dlGkfcPbIrcZ
4X0U4cUWBOBGBYPo9ri+j6EEt8h81FhKdM+iHnBHYX1zzqdMdmVhkrhmk1gbmnOiQoI6DVFJW+Zn
ot7rNkXV0/TyFLj5CLy0V6VH5I2K74W8vJa33VVHmJtLV72XDAlxg5TZ6TAd0CNMjhRgNxXMGiVN
M+Rjc1Sii7MAXaTE6d7jsJtWdVusn/8STPKwZeWq1tahGrTcH8F2bsAyb4KUY09h59E21MvtkmTt
8fWfIQ1XFMJpQtJCJsuBX+dKtrZBSoHgAg2Nu6I/5/kBAeGvtfI6IoaIwg0ndjuwmWK6FDd0UEzm
3RzZpgc7O+KM/xzZMgOBP4fES5ZimJV6Ci/CpqHRWV4jMP+uSglJ3emr32BwpfIXQZ8wOjYREu3o
f0jFofN8KD7iQjbZeJmyf7YIGRT1sQ/VkDh5zL3qOOUVyc8CV8vahYWKDvPM868Fg8m8CbUEIHVw
0BtN/x/NEkn7tWYYNGvWYbb1PKo6HKI5g9KC492ukhIEf3VRyRwmEaJBl8UV44ullZK00w0KyitA
/QadEIM437rxIEEN8A/ThyBt9I1LhISzGINcZoFImzRh5cqaqGBrWzQmo3TD2YU16C2ZeOFwLwD+
8/pMiaBT5dhDvu/wprSEFJQsYfsVnegUq32s+2rvK9r8LcswWOoU1Vmhep15G6Ta8sKwCeNvz6JA
apaymD9HGKgI0rLLGPCF28Mdev4tm6j8qyxvrrgVdnQ2ierrASdC8E6H9bGhYElyXlWvYeF+6kme
SkODcZtQFYkx/d2b5iyMMaIE4XY/oBSn6T4QEyiRZNzC+LyucUA449oik4gcNJeC3zBHBBqVEpXr
QVHZqNqjXN5jIzy9PxPnGdDP2lmRjz4j8D2s/HAlGYL6bPCCiGTBe+X/kq7+dLiae2NxPXwHvc+G
g5YktcaF6r1GVZNJwCVfV3nLX28gChZ5f8QSFej+rE3Ll3fSIvSyDJXz+87HbVOq3owwIk2pc7Xz
oTJdcCdSYrsL6dxyjrvuP5nSdi0WZV4b0nLvB7hreONrMPooXymUUPjqfiFpJEENPLYl+y4iDJyy
Z9p0TTXnR+8i4y799bu479ssdWR8f6GQNkqNdut9GOzS2NAsEkh1+MmdjpM8400n6fC+ViDuzGG+
fbBMmsDYXP65Gqeudgr3HyanMbsuoA9vGpo61tNUndRtz1Xwrrw8zdTvMIM3GxSSQm7wHXWJUvCD
EeF8N0xRfuW5Cyq8w6uh+arrqxLzgJhC0SZzRkZyAPTBG9Ov1jVpKkpoCg8ujoTHXAyOmIwTuwRw
eAdIViNaP/UEumHOK7PAhorIhcb6mlV692W1kDE9mNU0TLgGI02h8OL/+AL4yobdePPvT2GLb1a6
oOHPnrn0rNvPkp3Sk994TagyS8yC58lP5lI88ldH6r07TODTiqzw5hLpRHfw6VENgdV+VdD3PXzy
0r+N9hlNWeWitR51uJvFlDaQ8e14uO1IA2ReSVHZbqqQV4Xxa0T+kbMO5+QfXbk8sLwC7GvBsH/2
xe4A1JqxMueE1JxU6HUSFxyC2eVlsDPq5IcORcKEliiYOx21kKPr/Q7tM81xAPDgWQoFQIXgzmnZ
VXweFTSewI06Ly3Mb2kRwxGdVIj7JyPQy2xCCG7zEbrfalpbiYXAXKuELAxYtNymuAN7QfWmRoCo
eW66nVRPt3cDsBKz/uoPXFoAAjjADXJ+bvXN6FVgCPPEIgnR3SFWIWY3UXjjGADN49vU1tFCIKP5
glMk05vna2SFrSGbJBg3lTey/iaY6HhjorQ5a/JiiTZXsPuiCAQQadnwixOb75EyQ3mIm+0KVYAc
ZX0WnxxX5mwDEoMSof0dKZn7qMGPK16Wnursi689skebjB045zvS+12tuCuLOC7TUALq3A76amMf
Y/gfDrrNYLFlAqSvehGjPCq89e4BKu2femXSUWyKnEcGOijjKlquUy3UGGBgylRf0fo1H7zGC0H5
7Gjoc/7R4ZLTTGmZes89Vx7JxtGrIAufximCjTcHokVWaQXeYsWsQT0vz3sUdUv6o0q+q7RFG/RE
/0qEBlGj/fJ2Tj7hTdriW9HGznHWX4gApZt0dy5pWFKEjiqJ+v6Lj2O0J3LpIkRYioMhpudKpquQ
s3F7bdnJqJnEqBNNFjnaFHiWxLgHPhSCo/PF4baTN/NkPAT6Nu4qUGpc9LtBu46+CtLZLgKlSxQa
pw8+M152bkvt8J3grCUgNf9VQtVniTZNNqi34ewLgYO/AfpvpCKBqmMpQp6hBQFBjs87ud50VXq2
F8Fpy8furItjS0JS42wKPz2+yuk1y+Xo0r2NSrEsNtkIFqQwsqtTZaM180zoRGNdNEsagcCxxC/a
uN2CzOw5r59iLtO6oflZMiOgak62vGjA1xw5ToSqJlS8biaTMGPMlx9pvGyM/bDwKzJsUNmUCJsd
KZdFJT9d59YGmsB96uOmylUf1CGivJlSuWmLO8KM35R8ByFAxxKW6eR2UH+adxiKHjOO7j/lOl/J
M+BdegBNDJQPhhCEBxt37ellkva9coLBcQVkmfX+J7SF6xkA8jv5qRvtuV0vooAWqyk7/8d2mGs6
gjSIqQv6MzqDl5YZoZ2ZZln6tyAx5o200zzTHf6DpYwYhX0aoLEJlM1zS8niV5zSGzp/vbO3auXP
wIYwa1EF9kSFH/oV9PxtB9NOSs0U98h6qrAksoQgpslK2YAa19l7WqBoFHNnd60UJEiMZKNmRiM2
kVTRFE6yNZm/lbAljUt5FZ6sN8v+Rf8pLthNGbF78KiUUhZWhtEtwCVe8vCbIbMC6fuExixTPdyK
hrR/jjAnaLDvBTLojLaA/cY9P5m0MuQHTT0JZLwBMBOHOvw1GsOjDOH5Y5eZ5LcFnd8QNu50axAF
UdJd7yUWR0fnMFamxHiXWfgWvxIQlw/zG++2hv6OrxFVnVzTrCGSUsY4zp5ABV9DkZLQy/Zaq2XD
hgSUAXGEHlc5iVux/CkBMylKud+euYUb+GLIGag466XlsgtSkGLMNsz/cNpzD2TYr2FKHno8H3oy
a+viTHdoVcXt+WxNE1RleJsTCb1HuK9rJgUApO1vrN4OVhXkz13HwKD5iW3gISr8ILxqzFhGhBtf
5YKypFlrSTSd025Hj2W+sFq7eHLDMB55BDqQmwTb2Yq3v/gLy94bBTpS6uwocnlrN+drmIu0vx87
5TNJi8x9CGBNLHGC0ko/3eEHq4eJSKwEsIqejBuXwbDxPxmrImefD+rXu8rOi2X1lXT6VTLeG3u1
zCksmvSsd+t+8w8tCp+Avusq2CTSp43M7e59xI+0fvbFt7j/hdgWB1NHcHiIJLeDqub7FSg5hCHX
r1JENSFz6/1L1i1SZ7DQMT2YQVDxo+uEdtPz8EOKU2L6mnrdjbjGffBoSVYQ9b/GeeHQRE8NKYfK
OS86ynxURlsIL86iLxLDmV49jZdIgnyX5Yur8Pe+5Q8Xx6vaYVqXTzzlG1miZ7paeJX8hF/zjjli
FmROj3yFvEMMatWLSEjyw1E/GnpHZMTuQ6yBzpSSD/LyVoHByKdQzPnMxK6tKRHuVZ5jh5SweJsJ
mz7C+l6oUfGpZE5lvr97WpLAW/HV/t36GkgWWXMb0gSupISAYnAcGPuhfbaj1SIDA8T64XCWy6sM
bRxpWTpdhC7XBEvk73wCg7Y4JAkqYrT3PaeFKsuwYsJZaFt+c4YDfDsoNjvpOaqp28LdrfOXBzXj
F182L/oncBhlhJY3n3f+zQxkZfKbHuLP3Es9b2OB9ecWmknj/LalO5iDwps1xvPXNClDFWd8/Ffi
HsGuvgF9VAfu13oMQRvDAqwVFpeD4SZKiMYk5g32dfCark6/V/iXj6Bs5GogsKjykVFuRdhpiIbN
HUzxDQZSRL9BoZO4FJ/WMSlp1be/vgDrCfugp4avAxW9RDf9LtCDAxb6qgX2q/sfMvCSYGjGQat+
75oIlSRdRKq8Lr0gTc8z9MB9d2OGCRcXa6qtag2qqU6h67GPW9swxGu5nxVLExIWEV/uYCxobk3i
70TKIyXID5nsOmsRPKT+IdXyUixadD5pydhXOUWgzbzzAGeaw7T4J2JFK7nCd+esbzz1WM4cETrE
JqavcW8Mk/6iLGHtENoyDUiGHxGJzuT77IZBNGghJnoIBY6TiBUZYmfyZJY19gvalPmwlSUHbDOe
XishG4YrRCf78Vh3P2rNKne3cBYjivW1SW+8/lbUrN8Mpk6t8xOoZkAaOIVQcn0q2JRRGiKhIxtb
zU1CatsT+sz8SZ33V+Yl6EwLHip05LvikW0L818HZL3C2QUFvVb2lTNHZieNrjv328AqQfcnKCLN
b/4sbmUeHvBH2tlfvCJlbdi2l/JMtNH3K7+fb3VSQoeCsPy98TRK/BaDTdlkWLM+YXBkwZK0j/vq
yGfBTCdr542UYakI9Rmvg6njVMwnIBx9myjX2e/pTdcmvTDbWqchXZWbIYG9K0jTdOvC4BsuHBDx
a6tCNY94HZWkFvW2eF3LAAG/5kvjGXLQ9dytGJ4EXlgeQaQyMzIpL6/+L1ZXqXvJuhoudYUeHgYY
WdmKCShQvQEZrICKpWp8pKuBqwS4ZI54wDL0qQ2quzYAEPM5FBieQCtgwCwWJPz7Tmq+7004wN8a
800s7mAdc+SB1Q2JHz1OGVwH7+DEl6fcDQBoLrgptP0CtOAlfrVgCur9RGbOVIvrFyHqZhLfTrVi
4S2ZmqVYSPDmI7RqQMkvdl08CmzeDB1GIkJaAh8CThM1KmyfJY7BizwZZ3fj5HhskH4v4R74lqX+
we2GP3M5pjv76AM5fMdo1QhD7Wzw6kwrnnEOxc2QKLteK042DIJGCPzH4g9fmEYjcn3Cn+OL6HxV
wKkEfwy7kczFRCuPWsqu5WOeiAOY/l77AgUd8GJo/PvIID0J8GP5P50U5hS5b1ag2HJFQlTLmkAc
AKkEk34q7yeSDqcE6dzqJXymvF2JNk51CERCoebcb8u7bVuFDxdVvlqxu8HQmCn1bEL7ToM1xtsL
zMlcCM+BRdtcSiHMmaeeW+G3dQf2FWB4ivAh7Pm5Li17HoFFL3QS0W5GNorIQ/kdkh6Zb/YWFyJn
JHPR337qKayxakVheLc9+awAR16o3kMqWoyjZJTnNlFExXEnigoXYIJc+rz+jtTq9rZMZcpryrpR
vH8b4Pm8h6H+QIgbdnb1aI9EVV2CdppmCD7IY+mtM78EhXibv+zfjXqhOmWfkA4GUlr6ZvPzx0bb
Cv6w0lvlcsnf02a+3jR25jI3Zz9JzxxeoVqCt4x4Datkx0/bdxtRaGQ+hJH9WvboyH2Y9b1NXiKN
CIn0SdiGiIsZ9DnPsgzIeN5zo4aMzZA0/oreNhJngLf/io8p1AjCRmb9UBLWRpEbLyTJRKN7A63s
sbXvCZ6hXBPEV8KY49YTu+4dz8c7DROEfsjA0xRNP+hgfgUTLII/HNq3fYcxe9taSU3siKWSS8HY
PbIwAVdkGMR5s1G/5nDQfyGkMXKaRqMvKFkW8VbFhSbCzhFrTVpcEr90bLHRhTs+h5SRnrK1PxtS
2w4hR3/zJvBX7bEbB4ccKMwTibzcwB3WW1PxQz8ELVQ+zxflm9sCJdIQ3jCLFvM5Y7EqnwxvISge
ECDWcfboR5m0PqOK78w6YJe3H7lj7lAFuwqXROlygtxHT8NMR/EloZyjx0syGObLC7K3s+6oWlf9
9IEc1Zsb5WYL5KZuO8dP1AOSOT4XE1Css4X7VfzLKmK/5bK3VLzDbDoTxCXTEz5vAg9PbWC49DNB
M82PPQ0u2H2vc1kJABW1TGvbBTS6XjXXkNgqePtrM2lk00toCWclIsgYgFKVLQ6qIRUPoAy9p03J
SB1E29/KJo8HLYTlLrS6gUd2Qm/dV/wCEa3oMniDg5JPBtG/LqiDvOsr9EGD+zWB70jJfaP7MWt2
xOUiPuiJjnOgNttQvrJoh7fz5M4JcSS/o/dBafSDXKahzzzE24F92jwotIWLi46HUe9MCkLwkbuf
nqb+eC83mH8+IfkxLLjSSfT+0XpyLkGXs58zp+ioXAYDg2sms9R6LeMId1leOiQBiKk4YFqIbswB
RvDFobnrorfvpEQ/MPCOAll+T08Le3850OZ+wzj5q5fGHRAuLaUIxOs/ajft2TNw7liKtB2xFX0/
S8n/IeskTgrTmsdFEgIGyBymLTCqv52zoJecT+jx80hN+Ag7vU/viP0RKARhXZUGDug+2ajmnzG0
sbSNpPm4ksHiydF2GVYlN0CxKylzBKjTJRr4IXVLIfEtRSXJK2FOFvNWRuwBN8e27bFbb7WKydkp
IYC3FnlFBc87xcw68k2hzI0K9zd6lMiVYQxFtonGlQ2m5CNQevt4EGBvdGj+jLpzUay+9eP0Es+F
oOEYILbYP2XzGsMrMBXj6UT5orwHoHUB8/1uvBASPl3udM0q4yJtPvVVUSTq0OUe1KiS/cor4q/Y
UQraoBOpjKymewwK+wgCmcGkr9VzofgHn8nDrdcPqnbLmhN3jtRJyyyqoTole8ntgiGkJCKNcd49
uRzkPFsaWiwJB/MlNZv2ihX95L3G5DK+809orVEb4ZWyoH5QrQqPd5W2vFLDaOaDppQhrCOBYPkQ
5A8eig/JcnuabjKfQPbc/p0g5IQb46O1TlbiC4Ml05NJergvQePUkIKeinZiP+mfybzUyO23xYbP
9fluxXxYuUNytHiiXZVNVjg3T/lNZQN0StPcn3BXrrXI3Oq4EE61aekdPkmc3vkjfsnmjpUR/mwU
LxjLGxTAht/HDLpvZy3RXZbXfae3BdktRRPLuLPp6ZoqEhmvBsJVVckpww0y7E/HWatKpWgYXCzt
Mpjc1FBEG099FNw7XCHD9ieY6cDWPWl/+Mi/B6koOT2TK4B8TQeU4LjvL91VnA+lwtRiYemIA2g8
bEqEZ5whgPossJ3qEtmzcT3aWfQGJbP+46rZY8yUc9tNTygoMMog3HURXiDxnK5+xpt1ZmJ6sQka
wNjowvj3DdAFKGVjIIjkerYFSMSJ+It1oSbAH8cpWyMel58yx8i9UZpYlRIENRE+b/V1JxF7hNbp
+HVhSutiurdGt0m5qcUuYsTNCAjYhC7c2s3iM4ipAqsI9fEjfrDVyYddD4iuwniq88GJtpZcFUoL
N6xa6XYg9XktYqZI1e1oqdA5+5qe6DRvSnOQkXohHvTI3dEPWpRLZA+S8nW0WsBGblyex+HzoJFw
dr6XZtl74NzCXNnrup+EFF/qAuFuu+dotS7PvlXZygaQKP4h7FRMjhs47HcrPpo/89YougWGR7Lr
GpwxQD74eKoa4wssvV7MdV92s7t4yHYPymmjLjbeFsD/X6grNu4g2rwsddghPhFn3kKdwpIkk6fo
fwn7uFJ0RUXsk6NKbuc1sYAq1fzWE1EMGDA3HsiQflx928NLcll2kYFuNLQXmgv1uP5KNEfHyF/T
YdUaNJsxJ/zUoJKIIrypV2mBD5cdG6awf2Sgud6o6j5QfdHt4DwQ8VflMRc7gm6FA+hfKhwsEYZh
ypEEq/2Qo2hFXWwiITt/ApjR03SSmPh9ZxzVP9O74qbkNm1PhvkTDLgDl8FGyTgeRju9O4OroRe2
I3hgxWJo+3FS8+jTycyG4f5pmDlNSP6eqQ4F8zFWZOnhuHMekCgOOAerGs942A54AWRITOAVQJ4G
Ym0ctbi43HUmM1arEgyvsMWLIZsJM3ftMxiAJbhwNRQ52sSIqcwbMddl5HR6JAZq5SX7/uysR2UF
7bcbgbehHgkM1wOno6tJaWFWYhoQd9OJonDl9+lqZK2PT5/IZZad1vnNZxLuLUHuf1jFfg3SEJfQ
5LRV70W9HDXvThvwGgFYCMHzn35Dbz8L0IiEZ6lRNERWFfLH4AW3Tu/t9UE9LmiU0XGcIC6So1Vn
LaOX863db/ECE0GGgUT+2bUUN6ir2KmGBGos6yDEYk8Uhzru+BjMDHIyb8IfIPwwYn2aNNVmVzTF
7pGm8xEU0MUtQIwA+bVfo77nSX3fs+GZu9JcIJd8UafGr7yx+X+EFI2sFvSYkO6yhsvlNHpTCxhA
k6zCYaqbHduxX4mRCaw9TqxS9pyfEMYtVwMhBposZPL3aMXUtITq6bOKJzkb24PwK7W2/WoXoKeh
0Q+4p7AurQRSZhpVkmISsjBeLblRzGHF7QorXBmq4RBNts2Dbo0Cd8NZDaD/CzCvGmHc50YRPg4S
Dm2ZQyzEROCQSYvzUiFdgR0XZScUcFlYjj0TOd8hJnqCiyxd5i8LrS0kCKmiVTuG8fthY3H0pxal
U4QTtLcKwsUC7kfK/4ExC7wZu0M1EjQOCdB+6z4TO49bGEpl+BELBcyuJhIv59JjD+LfpaQFj19k
6+51Sea1BWCdfUfjNK/QpzkWPHFq4Q1U5RNGEROcZbG9saWP7BSpAfTwtuY04n0FhEpAcut/2OcG
b0jO2NmZ4xPJnndESo7K1BINQRi1G3j52UgVzmx9XyGKWrQaxAT9B0yyT/ccTxH1uZNlksryt6bF
VxbXfbTzwTX3vAFfkKHR3I2Tygv48/c9EJ6EcXm4iXWRQbzA/UzTifNFT9hIsMIfYdiCZQYDuLFf
/+PFzIwj1/DME8zTC+IUpVsFCdQihloxMqt2eK/bXy13WxdnxGfLqBsOO4DYBJNQjf+BujYMcbXq
dJ+RU2r8Jdto9WXhhxoz65DQa+ZyPtGwgiXIM3uaatj1soSMauweYpEvf9+ysXW+cHrW3xcmTPeO
NL3kA8fygbX1dsCriIWlk2S+KZ4xdinf8gBhkUUl6xjDdqOnqK1dFT0QJBc2YjgqqYM+f8A4zBIi
pO2MlSuK/+tvyZt3krryz8WZtwb2U1AtdQPYpdQpk9TPxP4w5cCG5hGasOGa9Q1ubaprBuNIORF4
oGt2ZkVJD43jrlTWRoVjVzNdqaD/CBDJ2pgEyZuaXB56iYMd0WCBsjj34FNd5KV9byleuLnPTvdP
oCA6rz2Wd/2GubD1SGRVb2UZttj80IhoVrkREFkcOub3P1dyxTqHzvN7sOR3IjytyLP7S6OrTRzA
7VCrhykyr0kDToYULg9H2VfLnRcq5oxaT71DkpV8TuHFjGI5zWrGHPrsGSnV/wC650bM4Es875j3
PU50WhDx+BiVZq5xi8OHC7lA1a085350EwbNnVkv08e3mh+Trn09m7kbQtrg3B+1Jtc4DbMSwSu6
fD6MFvqh6fxGe5NJE8r2RahcR3NQS268pnm5wNBmqFtDQhQeKRSszvmG+vYrVxa5MaJRX+5Ro4zt
UX2rrDDGmWaAGF1qbND56KJ40CUSyDvXf+F2e6y53UiscdDS1zRh/EfWd5epKoLrc3LlpEupHHzm
8ZQN0ipS3QRuqPvQjOVIPW+M6akWJrCLstEkOSqL/NYRGctV7GiFQ9oCWsduno1e2AlTWqgo2pLX
v88+P/GWKqQgkZUbR+74M39mxlzBhVBOICKK8QE8H87+Q6GLc1iKLRxHUok/o08F2wo3j3Ek0zIi
rQk9Z9XDYLzXYNfXg5PNlkJRm+vXdZ8LysbsprNSpRlfP/dGX2XU9Z8RVZcV7rwzQqsN51zzH34w
K8OUJvGuIBs9soI5o782YKzqDlx62++iTMQoErau0YaOH1NSyqiTstkrgpi9I/TwSLJPPwvGSlLE
0+HRcYpKgwqakwXT+wYOFw/10w++kU4aAUIXK3h2e1UukndETLD1SVZdZqXZsg6LyvTtQnJThXfZ
7fkuJs4RH9IJhVPCXwU2ldldvsjJs3Zu4B6jJQrX3IcN7lF0qC1MCkwkcfUcd29S3ks5F+SLE3QY
bhIHCSDaxTnnNlvlZ/XMVxZFWq3usRNYNZ2IxoSVq8UjxKZ2jqneExFST6mg54eqBNrbDGt/EUkn
bnztdOvWJuB8a/lbWDVl5meWqLc98KGT2gTb+qjPkTS2KIEw+Z4VjYCBzag0rFhNTMoVwMwTXHFM
pNYHLOmyjLcNJYFt+UWtAW7VD8WyzGQ5eID26uhDjLQp3cS5k4DoeiabYS5n+z3n1IJECCI0dM97
7NJyyw4reDE+pp1XDY3C/Iu89/c9J5SlzEoXzsc19OKZf6F7gd5pu/2psGAwxRXEmq0j0liRW/cd
VaFpSOhVnq+xmqf5dFDV07snPKVVNLQkq4ZIuB8hw4TSOmzaLkXG4Jv3wLZkUfEguMXBF2ofNzhV
iWaLBagO2Z+c+5wc2TA12pwKSvEmG/R/vOg2vXimbA6Pr/L4rNmVc5wyjCjf8xMBl7oYxGPKv1bv
TfPeAXeSt26a5lyaq/HWQqmx3FqUpo2k81PultcIQ99YX2kFxcuUhFQ3CixCPEsvo5FL1t1Bmp6E
iZQKSZXs7YQdyfZPTk2FBYDHG7KzKK4svsUH9lLECggirlQzcoJuBSy760CpuWECFdERqMHDpA3W
p14+MfRniyhDic6EdWKP4gSM6HFMV2KVj2wD1UAUO2JcSXVArlU3O2RjkE8v4V/EuZ5jW9vLwsTv
L8TQGPQdRJeEw8qqE9gpaye5G1yqeWiJuywO3p4EO2/Z+b7HS8W6FxkQFRTLIY8fjMBnPN3k0xQ1
oy4MKSi5tECwMqzNd035HAFaaeo33j3f3AhFI0hahQGUMWPqOtmNfPk03JRBwOgET3YvE8p+HIRB
Mo5LrmHqY4BRQkIFtox0Ip4vvdCJSgFGmEOLQZq4f0F0cH18fBOjruInoZmNMPP+Px5pNSuOb2Ov
RBUtaXHTSfQggB1yQgDT0yolqngavONeicktomQuisYDBurImw79fFDbJbgKBfwWS9V6SdVUvLYP
4W/Yqi/ESXfQcN9Usr2YyGpPjKP6dl58+kBxEZnWUzuP+YV4QMW9ULxIC97klOi0DjfR6y0LliyV
n/YfnAEUvZlR62g6Yo9hliqj6w3MS3inZ14G9mXwcMgZbjsMOR67sVbaPQEqRlSALXW0M4e6zg9B
yXhi2S1F1iT57+KIHYmjA5eWvO3dXzvAyMUqwTwU2niOgvyeV979rB0rmwyG6AsGQCgHRwbOIfoC
3d3P25BmVjkD2ReUZzCIcfkb9X/EVMZ1P0VxyCHkEU5slWufG4kHiez/SxxY9jG0aCFKRlCuMgV2
ZXfiTALmO6cEsZ36RPMtmk1Zf7Gc1Erj5VzZeBiGWDyQg7XeceyRGIJgkGjfGK7yoLV3JQ8hlnPZ
B1uuQoxbEw61yfTvug+jUyQgkJdn4u7HT6vX+jAjhNAHDh5GrBdEO90WPfMiZttdcR+llSyOo5LR
d3Ja6o/aKRQTJOMpg0fgAyWk0WHvGx26lV20eBfLmK3yp6tlK0CpxAOB16OpAJpm7xVFl+tgPDg5
ATGnuYUowaKWsWeY19VIMkoTjPw+7/5+ct0Mf1LiGg5uNop3Ej/1Uf9XY/eL/Vp9TReX9bDT/Dt2
7yskCElCFsuJGppCh5I6BYSfHEcC/Oj/k5C1za7beATtH22drX5kxiyhIKivDFF49JCbNWp7YDGn
uVJ6Ct8RnadqEoHHl/6N5zoOV4BcIpSPwEY1mLEbzufPeFO6O9hkRNmgA82j7aeLPTQsqHf/iX0W
1rNfVgp+XwTQo6qVoUhjM9X4eMlwT/Doir4FKWxmJrxHJ5sDFXM8ka1aMfD0CeXXR1hOsgIuQBqS
9slE9ikYH+79B1n/UXbMemCyuz//XD2JBit7mObEuYMjjV4pduAxWmy5IgUYL8cRfRsUXXzSdKBv
fgA0Tfn22ctkjRa0Bcd8tWn0F1PsbocCNpe0H99PQ06OYAzwt+VBZwxmtZry3mT9NeWaQ+8Cbi60
Bty+cPqQumql7PYlzZK2bdNNE4SNbwMG8jE7YiAYoYiCyzEfL9TYwkdml81RzbIzZ41wC1dh67jW
ICtZYaylvOL/xTK4uaOm0xBx0lkH0t4Zp/18bKNuisedGOhrcfvvpA9RSL62CCe3bvcwpzrvjRy+
3/VeAL6l1KAAJWtNi/PS3FiCHDOqvWgRs2WrA9u91t7EFyMjZJ2HXVX/7vAfyLb4QAjawm4n/EFS
GEvd7XS/WqwyDn3Lu+8sRWZaUxUJTln6jyZ9faI1xqJIgMn6Ab+dYxdvGBpmmwoe1JCz2HhugDtW
VVBNyNk4wJAn1auZ9ggMPwhiBhiJoJ1rTdVHtEpH7JQFuSsDlUdn1IPYPml+pq9of8HgtfMif3Gu
Y5fEHBV3w8HHfn27mTLDmuZSwqhMtISO5515XPqPspZKZqI1mR6SiMBaC2RCunfwgl7Nh5OcfoeN
VwYFMAFY4J7YcYHroNOeZ/Y6EOEYNHLE6lWzSQ7Orod+4SVg2BxgOieVtN6SiBwtJ09O9+ZNbr+/
cvtdQidP4XIb4+AA8W/VoBsdzX+rC2mgK5SgJH++OoI46solFgP9LDVm725GDdItz5255QBDtOwi
mmEW6ZZBw9Yjp6iolcqBiuYRAf7a1PPmnjpXluUAsO6xI46fPcGtSHkVZRXYLVwNRGzzedsTscr2
lRKR2toWXbdrWZH26djlKZy9fUVJjehVdFQTPaBs8Jb2KcN5Cah+1Pcar0i7MKu6m7a08BZjAkAQ
2yEoQr3NWyo6c1hH4empT1mj58SCuko+5icUtTg4LpKwW0RQj9/cp9G4o//Plcm4W8hzwKyn0Kwg
k/tZja5DjzHP/O5vWGjsTOJEr91BqMYfFGJ5xxMgMpsZCJlP5a/eeAJLZ9oQUz/OZb0tZO2OrxYD
v/Drg+OSKPNmm6U1ylwVJxfeAEqEs4pxXa1GebxW/zk42ydmgm3X21XP90NgRxvkGsur4LBDYIKh
wRHa8Qo16AEk87ZYT+iuct3Jmvorkbk/JPtZGdTc+Ryg3b4bp23IDU7yXE0WZYQhBCsYZYG/Wjp2
53sBTeq9f1b47MqztCT6bPXUA+WY6qOJlXIQgoLNe5d3YxYLNjPL0xSiSaJOBpyc/VzweoLkFyZ4
fh8CC16F/RAJJ7/yzTqKmFwsA3rL/rlXgN13F/e7JmQZBOHdsTBS04Cm6iL3uc9SrtTKpHBqQGUh
FqVx6uNbMglP/qA5xH0m6pK5XTRydh3dBtKhZI7u86rFL+ueXBe0tDatF9Cjksde6mYwxuZusBnV
t6Y0v8O4Ljgo5zMydS40Egfsf9ZT81KFl/F6gHhxGbfThZZntzkZM2Nb/0o5BJC4Aig/aynvMuOL
mZZBgbCgiyVcs5OlUvBtJpo/vYEci8Daf6Adk/jqPfpJ9BbADAe1hViOMMjxeIfrFM59H6LWA4kW
lgT3NmBScOt79bxZtjF/WxH02r+hOk5QkM+HOrv0cr+SP0M5c1qM0Sq28HL1ReABLdLLjxycyNgG
qYx1LAPL5inWqk5OvWt/aR/rkeA6YZ2HTuhYshb8C0LfQw10DBogWBg5A6Yz0OA4UiXRP7vxzXBS
MvLUuWy3SoVBzxg982tM26cOt735yLMNuvT4UU/PLbK9hnaoCDoI/Q3kMyTR9GPwxe69kS+9zPHv
OJ0Ghoi6vRF9+1Pl/SogR6TkvtzTuEVhQFeGrexu2FH44AOsmdJt+DOD0FlUOYOt048fz9/VSQKj
cj7KrB3oNQGS2Cz3+Vj888dUKTzm8dpgSJ6TikomNor5TAHt13QXpk4UwHXhk1p7ZketUzO2rFw7
XV9uGt/xdJJgOKhwO0hlSsyWgZT8U4rINaozHlxfD0TYlZLYj77DaWhYvAWq+bFXok44gqY9JWcd
b0KEueBMASvqiITrvBvfbhc3WY6ZW/SbVQT7QUgiDr/qib/i/qfja4SZkPjH6IdWMRy0y9mq14Ld
NPiBL78sZcX2Xyv6bB9Pt+x9KBDxOmUJ84wuxD7VP7IfC7bPR/J8k8MT9gh6CP0eUn+6xXP4Fa08
wg0eRGt9wdStGsfe/dfJdPUO3ofw0WkxeCbRXq0jPGRsWql91OTspNsmiy95ILh6a8N7aEh73xdT
X/VDtg6TcxLBNAU0NVhS5Zoz+Be4+LKPENaeOfbDT5FWK+bg5L0mfRkM9FRvfb/lyfx0+IqZjZTv
sLSywuG1HYzTuggZuuW0VXZCJBs2F19DLo3noVoAMN9vpns0hiijOiRFfFfo2gJmlXZEa0iaiDjU
nh07eRK5wEQP/MEilzQhuAqp/kc9AjpE70mQpUxSOZG54XLcMuMir1prNYamvvmhrBZQJIrUwvfk
2vtMcmsfuOujv8T8+ZJdgVkPPdIaHqe1xWmfknzwMnfv+XM+4n3hLO7cqv2/Ah62e4g8L9mLNSgQ
LvDXCmiSu5MXLPXGrL26+m56mGKURc8OwZpdeDRarYir0UcDwIHs2dRwASdlc85+MT7uKUgH3Zlq
8sPpSHGDEl0stD/JKiRcVxOMuxrcged8ITMaveiYVLdJ73ZQmo2AqwetdWrhpxIMbObgegLRvFiK
Quc4poIYv3FhId0rFqSpZITL0sf56YQznL54gwhmMRsQ1c8da+9tcXL8Qqzrjnz8aGX5S9q3uCdp
4QtEMeogAP39XKz7W8XEgEfTIRBTIEUy8qEVAy5Lb6trCAENJd4cX0fklEsipmkJc9gmBYwSCwuv
Ok758r8jN7SNJGwITrjcAU9SDfUy59xRwpZC5dJsdpPFBAtWa0V5ChnQgfF9Drx28C3lcbK/bAR4
oK5zS4c/FOYyE7VXaPZxQTkKpAohDoIcTy5SNaJR/ZrONRJIAg4NpZjiRun3h/BsUigF2xIb7y1L
MQdvpWqIXUP5XFolWbiFrlyNMoE3HDeW1MmQ72CYoB+StMyauoWEjufsSbh3Y1JzgBVP2X+dfXoE
u+Yt5dklWjzY8D9RmiN9bFgNIFI6o+XtDWkY6LfxpVtbGUjsPyeRmFfOIhW1MT4xAX6Y+N6Z/r6+
aj0YBfWuQK32l6XEiV1DfcFAKEx1rt1XcV+pNQNmmiipckM6umt9RSEsuhAi75tM9dWj5+chFl/K
3jBJPsAhZQozlu77rsFGiJ5wAIxQ/5+b6ZIAEs9Y3kq9qVqSJAqG67MJlPCjNcI+nQ33AV99f/xU
rwj/95o+jezweyLSbLZ5bzF/L9jiezYz3/kBhPsJn2XGNYHEw3f0TzgID0+/D8LbF9PTILsnVXzL
FARWAr0J+/mWOWNRMIkFmy1YWI+MZht4zOjAGN9/CUPCI9SHJ3BzLP14W3myB4S0UY3ihHy0OcTN
KmVwy6QIU9XhvyuMrNZXbmkuQAnPuvAfSWEm0JzRS7zDJbK5ltxLGbJNAZf/ECqK4Nj2D1y2H9ah
/m0qUuLznCcTUce+Lye/LmjxytMkEfV/u9T7iK8FvyWNmEp7ykfv9v0qIkfRMoHtkMWecBt2AfYn
luhb4UK73yucnxg/C9xjQmTCBkZV2k8FlJC6yDVryMFB/yrzvxYeD5HDuWOgaUg/Sca0oGb56MEE
SP65RqFY/oUlBGiMj0OZlHCdapFomzI6lMmLymGO7j8rn/KhiYTU/B1aK7vd/pbcBN0GaVYLfU3K
Plw+0wtNqLadk+jCc6sDRt7fNT1888sxJ9kEol0Yg/cxBlrsbZ1dU0GMGMRidWcc+njeOXzCTJmy
OP1id/3WEFjj689fvq+i0L/nlfQD9R0G+UzW0MeOCIhG8On0pmIMdWRTZ3PcF0xUIojmZnXvC9hm
C6e0jApWtb3HWZ4Cj1sEWDPoonWdTkQJVYXaxnB8CmJJSR1/WeS2MdbP1yF5cAQbc5EGHNQF46Ic
YAxc1vnFCH6Fnq5kbiilqveU1XZgKOp1SJhY376n2B9Xnv89ipRTL89EoDa1SJIuu/4WIBFyRzYr
dgJjQKLF/Bfu/XrXXEm3faosXc+pyZ4lRmEbdavaJrhXR9ieU2hbMiwC+hwju6LoZTnA3AtWphLW
M8gBwojsJGlXJ53SY2hDXMNK1ccL6UnuRc0eRubjlhI5AmGN5FiplziuiNKP2zsZwC7UUhhlniJ6
k1/dEbuFqQJ70VnZm3qNGsV2xUTLP0bK9wTDkOgdxHiQMr9zXeVdQp/XsvMeN3lnPZhbWyW4qulJ
9vt/ngclTXnlR6Ym4P5P5y9ovUkMPj+N2epqSEOnpi8zZANSmfa+i3lxtLJsM1iyZ5GymxrFDKDo
5Itzv4ZdYoF+PQrDl3+5EV5KdZoznx7PKH8EG4IMrJGx/RBKYrScdY8923+bv5RTlJ+K73Vw39Cz
oElvdBviq2sJUXcXN9r/sbyA8VhFglvmUFQXUPI8eHqasEL7nLFJ+EFsmVbrhrQvZrl5Wjk85Vtl
y6Urd/VwTeJoqBGom33DXLAgnxCujlCUitKr9bGQ2+Hln1b6Ik+PNMaDIf2QX0ywItH2ewgUmnez
vMXo4r9zpX9HAggTPskaBx3aNPsFv6Crazf7cxDFL0hTHdTp69IAi+YmWbg0dyVNmN1CXF9llyzs
UoKfPIKSkObB4LhQJVnO3pAkmPVweq6MNeeMNKumge6RdXblwR1PaN4whrBWoaSzn5NHeYcodhwU
2ZTHWGnLGFh41Y+clj7NUwmpZtG1yZOaOXPUp2vASa8RItWM6WbsxtvOoGnqhhHnJgThC8sRMuOP
gl0va5X7qrzbLHq1FuibCap9/jJzz4j3oopqEbynGppueeUX14P8IICss/noqoK8MDkUFDoHOPdY
HbI2vCqy/ZtKdY21g//mJAb6RNs1OVrLLvHQNOcag3rPZmJ3mrW3T0o1n+l5ZheRbexIDwl6iZxZ
MVHTay4lkZczQdDSLkdYdF4JCrGDcnEyoskH67ZTKvOGXU8YwZJPWxV4jiB/7nItdU/ZCHPKbFdC
LhxhwfT04jX0S4QPk9oBdTJQO15jz1zzIEXrM5qIwiIqhL7f/UIUW6EqV9KH/EsoUc7xE56vzhnP
PHTPnh8aaIggsh5IGbNidvANFQRchbWXN9LD1bzxP5P8zcCRGUrsTkhQU2fTOPTxILazFgK6XJ0Y
S2JOocwKIC+2wl94g/e5lIqdUxTOg31URQZWaYKiu3Ex+PMs3T4bpmTb1FE9KJoI3ygwVU07Meph
wKZUbOFJm27dptOTezRd3J6HOymX9VfUYL2UoDY34nSNInfiQ3ihvBrgWP7l3xowCNQKj4gtVZgq
Fd1jXnkH/lH/kkK87qMkHuB6fE1XWYuqPzGiZB6qYKZpU999jt7WJmv8CurbCkF7PFqm1beLqsRF
Kg4owIbpciolkTourXhY2fqXRwJSxXvArilf/djjUkOHlTOmngB8AtvlHYI8exAogz+1q9NopVe0
nmp9PgwzUNmk/WOmCKDU6o5Wkv5Y1smzOTGGo80MmsNYJz+/9xGY0x98ZWqjDbGpAEvWG4FFx5JK
TFjyEIPiwsspTyPezYIWmQndvKpyzWqRNgZ9L5L6BOO5tlCnxhQfraKDEe2Yz6S7D3N8hmXlwrSu
haYd/pNHqK5sFVzndMLi/H6d1UFpbjV8Zis7msM6zyopRaw7e9k+3z1hVCw6vn05HG5tDOobZcA2
FssT9V3q9RCHqE5QfsE0z7WQsj451P4VCn6yUxmAkeshr1fwGE+ObuZmJOETdCoiaTUuALp3pz8U
B2CPpzRvLsk2U/OWttCyxslfOkzRnuLSm/q24CkidTJ7yArOODEtH2x2b18nZp0TJqYFIXPBHVll
5uG4nACBEIfeAY1JUmEL1XuduwilwRfN5bfZlnRIfJHW1Xa6ha7BTVfT91cH9pItOT3VRR/jxG3Q
+4i1eBIGbFUNReGOlTdI1soVkmbwVIcJ8MaJj4ZhEkKqEUFNZJ/yw4xZ2p1X9/uMyiU2+s7eXc8Q
kb7W0oJ4tzo6q1kZHgRDbCmKxXC9OiG/BAAverr7SnJmrFi95BqiwBB2HqxjBbH/Kmy3pttNyEEh
4ELINAFiIioIRl+dpP04yZRLLFjrkzi0YCRE10UXBxuD3HX2lEgU+7G7zYl8yIvKxuiuTrniZ0Xt
srf1d3xgx4RjdFBO7211FoQkbSaCs+BHErkg+qnskqYwNWyDLCOZ0zpDkEE80+atO7WM8XVI7ZnX
PKpV2rvjFyRF1mFNVf0opbzby9q9KB4pNncMlbz1aVWS0aPFdtX55vzsqMzdicP37qZeqKAKc89t
fo1NOH0In3wggHhjOS0Z/t0djKwYfqKtTujML1MJ2YyFzS99X4LAt9vCLtA52wCrq9GjpzF7LBfG
/B4ZRsY+r8zTZ4QE5w96k8XXdyZCUMkDGO+V2ciXp9x+xK0U5bgsOEE6pIieSjqsuuOdikrB85wC
LKHPsQpIorZU+R22jwAPWqCNOrQGOKhiwhQ2TU6JYznPieV1EUDyRohC2j6Te0OdtLYi/GAy4ckH
jPn2TzZWQwwvCAewFMHzGL5yuq05VrO4gFLq2PFjddUTvMvmHbNWoJSwDPC3n1ciVngo6dE7WJrv
HQCL4OLkopUZq+sXmppVw3GaSem78cuOTfr0/zQYh5tLl1PG6C93DFj2j8CaoiwwYn4GwX1etgUl
X316RvWB82MU57xAtfrJ7wc845Fqsj/zntDDh2Zx6CFrPpv3SclzQfrAzND6nxBP9PPRZS7gYImm
3uhuANRu73E1nngCTWq8nqqdUWRM8WMCsgQUNjx2dnr1/JCn8ZjZOElg1UQoqnJBNqvcYtzxdSS0
q9Vn5olV/l5iooIFArhPKms95sudxqL8PSpslgmvaQIKjrKYMdBukH3Ux4CtLgvWUTY18G5Ndy1s
XCTF1Ga1phBHn+c+/E82Y1JyZnt75I16VMgCW20i3DdDxb7+GBFwyR0wLowJYMobX0/LqrfdKCCN
eqWiLp2GTxzPf3GmnwPJQwMRCOo7a25XN57lb+qmItLi30afw8gGuXI5vnWrlVSAy9/hub39AaMK
biBkmQGf0Y//6zcgiaaFVLcgnPMggsXQJwWstdX/tGvI/bLyYPhj0mRVTicmHQo8dptaOoAJK5y+
wKUhR39d7ckh+z5YRHAzHf7SD3QMYGaa8MpgbUx33B2qiU0mFklI1r/phklgVT+hAt7aKDj2lpm/
hzfVDZMhDTxiXqjvUfUykGGkBgxGHepVOPhnI89teMpIcv0emspfqR3C2K9DUHg0RJV7wF2IJF5G
txACBdLEFbDzayB54ENV5WxSBeF2ICUtxeMAeDdYuqnDQTVzFoAGyd10okEEf5L4/v12xM1yR74m
bZSavJDLwOprzjgdnXIPFa5/sR/St+n7xWildw5bC0Mn6DFigr9gJn4DSj+Io1KnSeOMHsmuKhoJ
tK63g/zSG6xBO3XSUJjyYxxzNMUUD4BU3XsldSdwpiJTFgZRsICBOtycYVHCR+TNOmbxNd/EcCg/
ypMyug9oazj+0nC+qqkPW9bU8REIKtnpnijmli40uelPvbvvn4NYIeczGRPurcIsYIqw0XN9PHu5
PCC9beLIblOArKDO4BVmxJBn0BDN4YznBdI0qZ8OZsmUhZsI64UxqpKNZfAYG9xwMxj85qj68Vqr
aQIzcfhUZLIbK+WXL4ELRXZL+3bIcENAUw39F9D5IdR3fiz3qe383JFKUu8lxdmI68S1YIZC0+RN
LkJq+AnAoOgA8eKJKQmZ+AY6uhpB4YOK/5jhzE7ftIBNViDyzzybyBgXuhwLHp+/ZhX+RR41D7sz
DitsbwaYjdvlq4rW/OMuEwG/x5SDTiJ5IaCJN8rzrSS4Z7fL0Cj5DJ4TIB9frzd3S/CwgVce3Zxq
i54LAcLrZBzS1WjaBupVmaISzOgHbQNWRC/JkXyNiM2GN7G5lsfL1xzX4js5mcO4Vlz4uzXsVJ3A
q3qi7/brLvGkxPUkOUqN1CeYemy7HCE8esV3/olrzcvA6w/RkH7LY5GsIqys59Zz/2TrHaoCzXzg
4UQGZQHVsW7rMoKdqNjNdhtNjMF5JHLuGIrOzAvU7tjJG25UwQeEQdqZ3ayRfEVyvmBx+NHvTrvf
NhlfDH0GyltPe9trUSqzJVfs8PXwSASJ71bnFvcjfjNL+HYRZvjuK3z5t/TpVqAZwmszNH1Uk4ux
WXCkANRsEmh4R/b2iH6nNWtoAJrU1xiUgLuMm6Iub2W4KMPbOMh77zmhDDIdervlki8xfYMT58PR
slgBGoA1R4aYeRc6CsVTG7tZRyTR9ts+pSBRkEJR+l0NZcHdVIWXa5GLzx7ZBg6BhrzHz9hPUKsH
NbuJdP1+khJ4FZkeFhKDlt9NL0PW5+kETJWXjJ8zydFJtO4zTCe+gdc3Edv0zmFeRyrDbLPZiRp6
ORxQT6b2PfRe6f54G/wOeTcvXBa7HI5/X04xTWc4FaqQqg4L8SFU06mwXtZ6/p7F/WzlrArWY4rN
hYhX6gAcRqPJjVJ+Fdfdb9GIT0J98phAaJjuyHQmLSKjvtwoIiEkSB5sTy6pRD3F+9+lX2PBKeEY
7JMZvKVniopamhZBftK8JxEEsBbfZhJyjpfh9nr7ASOskB0l4M5Js98YDyrZvu5Q+RkLlDkhurYp
ZVT0h8icsAS9ynvLOI4twIOnnEBZvf0P6F7qhYnlUJ3l85TwxHxc1T+pXKjPD9DG0Xmw/vzlpo6I
W6e5JydkdJzAWlXh0m1QKZtHUrSbyhjcL+EFodB3U0hAlCku/bq0urGPpz6I0Ek6gGt9dEJXSEIG
8Aqpt8qOI/e0fN6UpytN7C05ZUq62yRcbPdGznMfES/+FRFHSwiVEXbVp7HYB4b9b41wvVi5negg
sDjIZ99jiGl6o2NTyHTeTbWkfootaHAawCc6AgP8E6SpYKnAKQgCrEdVm5cyI9PwgmvlcgaVuaGD
xQ7SWSS9CqbS/URIpfLmeWWyAyFhHbjffRlCZ9E0odNqDouHKWykY8JWKkcwL+U55uWkIBvVTHO2
Q8wLkZq9RMZID2OEle0eD6iCo9xj8WljKmobBLbJtOL5wgcqs/utaHbOaR1PD94bxzinL/RyMkur
yLoQhYL7nusncKx2dFRJslutQ4WfKb/lNfs2Ag+QTU4YcE8338lC0mqx0+UGb2HO5hPLYQUgS/cR
TnL0szRiAzJQeTr2ftDxih/UY/cCBwMrNJ8adgE8h/mq3YtZXqZEOJnFHWVMlrrg3w7F66creKxn
xlr92Twcf8ihvpuY2CdD9Pmcf6Zapw4cRhBgqCTbK0aSOB35u09Nt8vvGK4sxTOlU7Ubh0Gg0XJg
VSyLcZGvKygtDTXbm7+40hp7wp+d7O7cm0PQjeTgf8b8W1jT3j3WbF8yTvpxN1tpOl1vmiXrAw+x
/E2/nGOKjv1C8KnxH1GQZ+cnKLywIKpIs9kB+yOHynXVlEup68JNl74qcylg/l8cJSDhxRf7x9Y7
hxgA8pA5mM8P9xtAznngReWE4V+hngb7C5EAzrcq9zA5Szw4hy9Z1026mQE0N1RG2spt0mz6Xtlm
JYX2ko/JXiLivzp/d4OqWvG/KH5ZnjSNtUYvRNqbNXJ5LCb+wU/PY2NEDO2/1D8FFKz0LwTXkjX7
kiICiXdNJWmyUmQCpzLrgLQvoNo/cYPuwYmK+2Uae2q7mEg1RThOCvASMQnlcDTcFblSh+/bK1pb
A8uKSkihKKbHaBWtdfIyI2RcFj+7qCkWRTOcZOCa/RQWjky7cMxxNIkJM2rTbvfg6V4lsXm60f7v
lxWLCIrFi++stKH87ajZuvgCnbYeyrdZ5PHX1/D4Z0IDvefDn5XflG2xmGazZY+gV1Bro3zj6Psw
7Y18wkjXbNsVaSoEUG1W0R22np2rb+JZVYarRry4vSw4wL8XhiEONzwMzpNVlC0SrnSeMpAYYbnc
/ebr57SMltviqiw8rUd+fzgWw9Pc0b1QkoAy1NtiOru+E7DSaSnafmWqLsVDrGjvnqvyI4s0GWiT
6Zn/IXzKgnr/0N1A7g61RxRQsYPG0FL1SByyY0+Crq8AKYpiHOWwpIB7/QaevlhnheEbjfvTdopv
E6gdnaK5aiQqoGjnTA4wnmNs8hyVvf7+/k+U6rSlEKkfjVxV0p4Xi3RpGeZFcNw2Z289dstxdnAC
OmnXeJnbwum87QnyIFA8KLub91ps957j2NG1rbPe9Q/mGe6Mvmc2phKbOWWU0wkRXXnHMF9GHAqO
8YnfYHfbQX5g/Ad4ucObaIKDFKuWxzQ7HHxhlvIYME2TDX0G8JQfCzZF3skvsVN9A9fZ77ezDSW/
jolu+PqqfXQ3txdaUv8mw71szGPtHQNxvm2ZZySbKB5NoVdNooeSrTfTWSpjL86R6ukuHdMqsPwS
5mjEUBa+hoABXZuEImAsjPargFuHm+x4/rb67kX7HeYerX3h4hJF2FLNJ3IaTPLn2kIhc+NH63EN
tD6N+2M+P+jRk0hLtnAm0wyPsX+gQ37khMlGNVRCo94D5k5VxmkIiwRySZTkIvYiZLBj9MS+OhUK
XXjoHsfjqWInSf5CjX/NGuzNCcn01LZf+92yB65yetMwLrdFodYLcwJLmf8ztANRAGWC4GbEbl5l
8fu1BAWR0ilUU2eL7vg5Lv1vvWgdJVxemdr30e/O7ygXEqAdsRB2+Ym1s5pb1u/TtSJFCVjagFVQ
7iFoq5q2ZvTZuAK2Ausn3AnlY6oaWFx6Mqjs9tgu6W2qj83q+PGlmdo/0MM/2iahB6qd8xL8MQom
6HWXBwwURdUVkKabfUHUQyP7WY51SCmX5bDBZmY5bLW8Q58JhoV6D+fazrLvgAym9JQtlpeCt/tp
8VWTmwLDsxiTmk/SIZZotUg5IdarUDNM09AqvRKIQJJQxrZOj7Xm7NkibjblbC0PUxEhtdYOzrt4
sbqRgWkcCWu2TcPD0JSUqMkge4pRvU3foC4CmJvEfuehRsH5ujxX3QglSZgoHOo8Ahm0HARMlxgJ
XWkvGfrR7x9NyuX5Su83LikSAoL8YWRDVZIUyaO8V6Kwq3JiD7MgiUA/K1FLUx3IVH/P9aOpnAdh
cDuBtSNQeYZ2dYIgig6NoLGnxpvYw25x9UwqL/ejirW5NPS07tWv58RaHa77Bi+d9pPchejnB6A3
uAnR1lx4hr1Gef8ZKSXj6qtWCvI7Uj4ORFBbf7qBYxlYGtm7TH14s4HmYZnohjo7k5FJfdGXVcUO
BirhO5jZ5FzZQ2ozVQ7FktWZtsK7b+p/BYvtuO48HcM1qahRHpWOG8pCMri/5s6ds1xQTxHQh872
lsyFt5Gp5qfp2rpS46P+OnBOLWd0Dwke8qmZ9Vr8LgCqza/ejiJ7xfmAAo6Krk1lVfoj/Viv00Jb
vq4ZGk8byXarRZ9QWoc8jkY4+uuono7+U97b1TpVBmXWyHvG3h+gjCDsX2rBIUdhmxBC1wcIsKyW
35MlCY36rR38qFdyZV/qy+4sx9M4hFj8aigfN1lHuLfA9tH5ugaVYcKRkZnaCQkFExmbjC8CL6oj
U6vrfsVr7BZrcCJzi+XN2qisU3cQld8boK25Fs2chnGrrnPM2BrNQL88qGOuiUobd2GVE/ssLvvy
OwzsLjgji35E7KoSc9ZS/pIDg5V93itVokWrXLTiJUmaVoWjkQXAwMy7b0lV1JVaVdgXEpHtUZM3
Kc7xMDvH3xhvFQrb+UQkLTb+pnvsjo2xW04TIBwNzkbyjwIXyxABZnsVhbw7QvA4E+TEKP4tgxhC
CGdZuCmoLBsSUe0TeqVmEKoYbIfCNDdOHSVIpv54/N18vvatuhtulw+ZKGU7++bmgb2oES8LfAYS
cQ5h5tf1OVrRYthkOWExl6n1eu9LLkjW8XVNCS9QGaI+dv91u/Tu8jginaUBEbKUmyOQmFTkEQDh
c4nn2wTAcDEO9UiggN6GRw6IReiLq3nt544rL3Ge8afrMwEoTNrMKsJpvUXLbpRy8ifcMGxpRejK
s5son7AQj4pB/CDHXV2xG2N6do52ZFhp4SJzRXc2dCucN8qXNma3vDLWkWWCf9daT+vhrQiAlzGC
u4eQbJRl3Ed9AfNBeDd5qFQWk6fVho7k7y9Zimg8IfIq6266fTYHf5JDNVrfqkFrjQgiNXqTD+Yd
WCh7NdPFpueXJOoHUexTkWzKcGH4Ia9TXoEDwBRH7aTyvi5V5mTRP/pQQii44xHeJ39qK2PS3mIE
Ni+p8oCsFE7u/kPIEPs/ol5O3LJWoerIfB7RUGDyml7MDy/pc3r3eO1x1aj2Rt5+j9JUBrOAVnh0
QznuDGxxK8mT9/6g/hfW+SZ74ooWdqsZ/cqqo889KGmK9vsXz9gLOnlmsoVqaJmbbhgHejT2/2Zt
yYcPjlJPKsziVopVq7Grkb8wPJ1CFpau5uMjQNyGLPl8qk2kJDdNewmy3WYU9dS0sOsaqILZd33B
sN2KifQRaT1lrO4zjPg4dAVeNGhaP7rXGob/dTNhY447ORSm5frhQ7yszh48s/+T558Z2XSD3pR7
Yarqoor91XJ5Z2ng9D/kK1PjD3YKDMPjps+Tz61IHc0j34pbtJtAxBa04kVUuq6Xof/XfL9t7xID
d5rdTKrgVdXSEO2z3oMNQ+YqQS2apVx56FycTX6lIZGZ2GRyXM6qpufYyTb4SfzQyvTDB864bPWG
QJz1FIOODo+AL2DTRv1IckbfFaJ34CKu036tdbIuij50lvIvqgfoXf3IAlD6XFxZJV9kDBlDdWdZ
1hB4QDuv7TqDLvGWhhYFBlnepDSquxtlgw6S0rGmXWo0qCCdSZBqXOQOHwZEgJBdtvoTUcGrE51t
pOAbNbVlAGbxaQwSnS/G9q+5nIwJlcVN1326vau3OAYOH1vztiS3iMmUAN9ZnA47fB7c4G7wBjP+
6oOeRZhr1pQD3GYBTbv+4MfU6UTdVWmRpgwgkt9WCfKpEu0uZIdcfh6uvwK6DpMby0998V8oqPS3
Df0aSlmgIi7VbNv+2duv3mokXJ3z20f06ZAqeXuFNj+IT3Delht3jvEULCooVrLtaI2dmPYbAxXE
RjuyxYryOSkzOZ2NLFYCgRiuzGs+q7sYw3JkYPRcZY0LIGej7rvEZHKGMCo/PmkGbIAEFfXNRwPo
0qSZollRxzdYHvCjyT0+1r9hw25IOQ6Et1uNIl+5lVvV0msJ1++4L5qXwgCdBG1aKg3Y7Od9tpVp
kiyIHZlZnsuGCUKXb6yGOPpxlWlCTj+CtmFCw5As/qs13MHq5O1f67Uf0+yqPAJGxgkhSJvbx0Xj
AnDSMwZQhKpgCLjeEX6+ZEiDygLnOe/API9pxdS8DMFfunFDlQR/TfzkS2AjaupqgF5cPwuz/4gc
GoCHT89yKzauanNrhzm99CuY/NJFEmw6WRPhJN02v3I5P3JHWN8XY3lZp/jqnls15FIm9JHLcXnt
QckitLvfCGYMV0IpjoYlRgsoSpcMNASK9hnGizxljmAIZQ1E2sO5+weBMLUU0Q2R5t/gITDOOo9Q
U8NR4WNiJRYAsoz7fon7AP+SOU9nHeZz9H7cA96i230UmtuNQ5FWrhytod33MZoT1NPxeZpoNqDr
xoa0T43ufz+iVfx5XtS0SpoRzDspUpjsCbeE6nfHo9FR0HKHsVczYWVxN4TqzxvVw5S5fSrECrn8
olWpvRIkRbS/E8tkmaCCIiLFEgmqzI2SrW9dbpw5SLN2TgSWF/0rjNco6BDRGj8YHh8OEWutRZ+b
qUWflyB6deqElc49uYc4fPPW+yRgBeIiK7QqkoUOaUJv+HsQvK1tbXqrpzBiTkjrG82GF668LLOE
sETO4Vqa1vZCLn0qZ8tlQWFd3tirvY12Yv5ExmGMFInVqC2tlUHR2d7Ztu6DKFEMkmTUH/joMYpk
ZYSfm5gXz6N9p3z2ACigMI7wwKMmAq0zs+vLgHjdA41ByG8yK7syyTsFrJXQKCYJANhBeNZ4ifFc
I3ND8wWdcUS3NiBNDX+nNaqVHr5f+qcqCngcThd7u3zERE7TifAZqNCVDcJuZgSbzo+oaph89+EG
BW5DG6VmjUyM3HeVs4CZ/3NCeyyQzJvrSxThGWkCqoOo3IKYK+OJeBjBgqz+bWepsrQABN27sCfD
qsDtdStcghgEm61tXAV4bI1aqnBYHlRspgCmiDvTFUp4yMBagYgQ3TgSbo+TyYFDoGwy+dsKclKS
WwXrZnDeeh0KZSiQ5JHc6e6DMXH+U+gYfKheJ7fBHiDKez5hw7mfOeTm+GMlPUem3Vr0hEH/dDcO
fGPk1+2yCagXf30gkKgm1i/wJ5DovH2HQO66nDgjGlLglH0ADahpsAX0IPD0+SzmSr+Q16NrQTLs
acaRLUEjnyEtaog8RtC8agOKQiJMp91NdlR0CV5/PiZqBRIqIMh44yzqFhdxVtJxDZImbc0yaaT/
KOSmGPN9OFI0YpgXVEarvi9mBwWVQlj5nPAJ6aWqnr1/JKajY5+dWz4wq8ZGIepAU63+37pEMQr1
36a+0lSBOHYCezn1nlU1EygcX9VI1lfnZQFLYoIkp95vuVLbqtMyuvNWgLAFFvblRvtMJQfJ3Yxr
Q5qVQHEaEU4Qc8q4Yt8j3kFD4VYLtCnNDPom/cBCq1L0/xtL1anynheeQTNtHQj3O99fVKMlFdGY
0t738m6GnTMasFMVOAc5VDwhr3xCvTp559Xci4M4HBuw/B8NBX7dBaWGKifAYL/PMZ3Pwg+3gK1a
YSqtW2o7LkdLcJoieQlkjmx5comCj8gHOz3s88Uf1iAExo+ZWG7klkAYbEJ5oSVNO9fy0aG4kU0o
1CNbs1vsizkIbazFAxjPe6OQ5vgpTEpoEb+TiFGI+FVoXxIx84Gmr/yZ4aTMY3Yczy219TfzEGWQ
ILGjg9z2Vpm4ovunUZzMvqd4C67d8K31X0XpKgpJ4vBeon05O/xYedDatYqFJfWBXtHa9er73wcl
hAVONFfe88etyK6ehVlbOy9kPD1bBuYcun7Z9qL18nkPum1gHc740ZOvRDAYnRDZiUy5SGdEMfLY
Ctjf6YzSLqRxZFtaV6exBavD1emo8kaOgX/JrxclUojxMrxoJDAdBlFuHSpmTII/Yy3G+xWCRUca
oPNChzLX/d4/5zvNMvdefPF/O1GtRoNAXkYxnLwQScsJOmNdq22zBn+AKUNDBltRxHjt4ALW3mrw
H8f3Dek88wfUbyMTPFWJfrF1z5O+TrxlfjhWCkYvChogZE+p01xLBMZ6GRW5LnuKLEq21/mFaw1A
gFKjKH1auiaV+X49nR4NYZ+iDTL/TX48muIhXv0CsoeE0QlZkYzNXfVVgyqxrigqDvX+9Qu2U0fb
MyCPMUtYDZjqAdBJfxK22SzOY3tRvjd9w4EeO7RB0aGT0hLENpMt1ArAL0L/SoXZwfPhkZ6zePAm
+dAEYw06d/uMfbDCb9FLG6uJdfzFLUUMbR4R3Yl9EBXrd+ap0tiGkg8+7aGBLhzqDGIR8PT92otj
Xd/YLL1+Pd383TpoBAalYcnhWRzQ5/Q3kvBgp0DEShfqa6ccObuek+21K1UCRLqRs1wKd6y0MqUO
4j5QOVfwkfEioKGt6zNvRDHePzYBWgWwiSHp2T54WAFVK2Sv7S6FXDlzXUdvSP65t47CkebB9sP+
cKYHzfVAPRBsKUaiyP3a4iO+PLFfRy969r6lo7Q8ail0fR4B7bcEIwbTqMfpnYam+k6JFAiiYhwX
lDMgBtdVCNiPEri2mEKfgnNOZg/r311HashMB0HqGCXQ41QEedZWAE/vXtLGAZldyFYBRBreNjxE
3VEDohYA+kLeDUy8nFx8gRTuf9xOwuSlMN3Np1/K/8yUAu6rYULrXouy7W24AmffxHzEMQgRhjIG
PiedtOucnIcsFfLNMZplCcTtN0QqQr7sNd3qE26rtMH/7KBQhwIjjVT7iPCA5m/72QwmP0ae61hO
JZ/8OyFo+6NvaRWoasrnavPwVt9pQ4DXRODmQxjGN5Kwy3fHmFj3LKmj6DUxa4X7ZZJVQcyIhRTa
jRWSFZHKH64Ky2rKqoi+DLPtImU3CYffgnCZfHM/er0Z1WOKusHb5iZLFph6MLW8Wol0zkPtxek9
rBdaae+O6XlsOkNhVmSfOh4KCnV62UxGHmrbs8CCtd0YIYXcANU0U1zd63C9xgAL5j5GlT0lBjjI
TezD9nn/j49a5zsh61HUP4XdAwiDub+FjCN8iDrjLOP0vi2cBgU6fZ9FJVh1Ep0f0NlZ2pmqqenX
5SNA2Dn8+TeTMkhM9AMKanEyXUCOiItAuaq0dwKVJCy2bHzdRslGl+a36eVvsA+o0uKludODHm8H
s6Km1+r02ix0zbso03AIbBVPlOrroz4exe3Xx0q+mme5wSpWl8J+xMSU02L9XBFR6saqQIdTmxzd
8pXbc9Y7R9XC9+96sE2zZ6Baz6wlzQRCqPetyavn3QDaR/BkESi7WeSO6Mjhw/pezVY4jDBxrhm/
JI6lSvNwNk5EE0mXvGRBUKnnOZ3kzdr/ppmgMjWbCkepXt3Ob2R1g6t4F1XkxTHgomsRZ4sImsWo
SqPf9K2csNdPN38A/4GfXvaTGQRB4wHGTjDLNbbqeHqGSOxGIQp9H0PFMKSwsgd+eNaF5RKGzHoE
sC/E+uSHg6veAy1si7Co41MMV6IsHC6/5wbJHk2cQzYvV8hYx1D6TER3iJor6Y3gQKJ0rDeT4ixA
dnQXBwRJnzOYKmig0QYywYkzFiVUFMBXKjezVDArj6CqR0j/2In368rTiBo4XPaeH0GnEg3D6sfy
SIy/3sFQio4JmCAWfZhWiK9TOCR3iMqxguxFmhUpIH5nP7j/BcaFLYMYMS5NjEXRQPfUcmzyGV1o
x4M9bBeIiNjOSuNurSV9wv2fsy3685TFjavs9pZ2oOZndDIMxIvno7cRy60d1SIHc1cbmUNuGdL4
d5yDckyA8MwgMlYt3GepT0+jiuDzN/qfmCLlhknOWlNgrgLMuRng6BNvI1I7s0JHS+F6GUsqvP8M
e+vJ+mp2XzH9QoxPoBGdOIPlisC2AUStlYWSH7buiCKHBB/CNIpa7oCb2zsUnLdwN6arSpXalEnP
q089gr2iNJR1BoH2/EKdYMy5t/scaQCXUZ2ZsGIuzFswp1DvNy6SDsejPzciUNK30SyI05JVoumy
8Vs70cqIOM7k/AQ7IY5VnhbnzIA+O8LeVZtagxSXBFpChGeu6TzcZqiqcX8yWiFd028mYz5pnEJw
QbQj9aaQ/fs41nRoKz46N9mzVgkPXXb1p+SjZW+kDW+zGoAFzIGIS6UpSe9a59aspSMikck330Jf
GqEordGj8fIbuAn6K4A2jtRF+KHQ1t0cqum7Kz1JlrUoN5Rai8H/Q0Q5o8dpzQV3d7P6wkn2Zm29
I3N7EOnLLmhf7QJKcGhYE0K3KG+U2LLAGpfF7F4OVrKvfBo1/TMWS1KL7hnQyF55j2XeZlFy8+8h
yM45nbF/3c1zxMFLruyI/8FBGJFQQ2uOt5L9v/Zn06MtrP6CrSpFZExc2kgm9LNR77cfjR/xbmkv
BIPygso9dqXRb46PWqPTzI9qiUwlfEOQ7zMfEPqlX+FaSyW9wo2Np318LBJ+bs4btbRz7hmBAvlD
LVvG4uIvmVP86DNkLkheiI2+833DEPXTertz0z++FSAbchIyDVKyluoVQxEQnfRe+SjZ2nET6e/W
0LOT774mbgvcgebg8BpmbWtr4b0zUkrEB3rAwkgUARugyCHxjEK0HtMeGx/E7MxQOUPo5EDPzXHD
kGlYMPI1Z8N44y2pSt5TraU+0ED3EQWTm1dkLmy3e3bwSXRzWnxVW3sgn8vQocadYu0H/FUU9j2w
OzdbGa0rCeSw6QOzjtvch4NmHBcPYpycgJgv1V/C2jqZUBsjS+ZpQQmPUEZMGnM+7NU8dGcxcdmU
sYYt7aH/REVjGPebHuPW7Cz4F02IalwSvSdbI34VBZztvZz4BOHuBYW0uQonn/j6hU2NYxu9lfhK
jn16bcZ86Zr4k3Mwu195XV3LRUkCOnXPvR8Z59WBHHobNUGnMUPDxJJm7mIiB69NOtQ+O89+aWC4
A0qUoIAss+mIadyMZvk6YXs3mjACj3IVz3MQMclKh3COuSF/zBY96DhsAbxzy5wono/mLVIGqfPe
K0icte4HHgvVJxbmcABACVhw4mI8KSyjOEzG4MMV5CundVrhlI8EBqXs43bbLZZki3P5bczgenEg
vFhc69BAgyife63fSc3ZfUScrkWBHn9r7PoszJ1grhMR+rUfnYhZlowoTubyCh0TEgcShLbYqplB
devTdpwqoBSm0UrMEQacuAxiWNnByIFuCPndKYS1kCNdL+/YAD7i1r1YhoPrTPlM3BFDGvFdN5ru
bEViJsoCAaKHcq7eJ76fKJkAgeY5gnqyTZxwkKbm6kn1hYHiUEyJS1GiTT1xvsm2cSz9ezqTijNG
8LvzwOK4Bfm7ZdSbtpisCG6zzHhonjMjuDxA6xjSTAdBzKdrAmvUn5V7E49V1n1YhTFBirEtWmqy
HRkdaVIwWgONtAbk9S2WJ7K0Y2onNO5kHxo8caKVaDP/SXAt0mIaoYn11LkHPoWqZnVkz2X9cMDc
pOKz0ba72BzrRQeVRtzaJRC/8x1I/7zTt8bTltGQk/Bj9LxyKxzHJbQWxHNcaRB2a2vO5z+PcDrt
pouzLq0XnVOSyujK+QzBOXop/ld+k6plKNXAFFQGAP8G/1RkNf8gl7P5ZYwea5xKwQ0DD3tdnxZA
xWPWGMJBLD3kPP/ynu/gQcPgeSJZxvEsoVM36ir8mkANwgBb0cZ0JEM4G/WYEvAsNrtilU+V6AfV
vEvL8D7O6cyGiYs1rfebQig5jooIRgETOxsX+udIJWiM8Nx/AuWsmjaPpzX9eN7O1kraQSdqxHlv
zYFbLEueK6I2HDnEqZAUaOg1jY/JqnuUArdJGlucjRfg2dfzFJUXaMOKZC2UW4Ed9F6seLXX8FIS
YYSYkkF9PNhZKKMwh7BClOT2MHH90I8/MDIUaqbsY6Na11EBODp4oXxTFDoYezP+VDax1Wvyg3N/
6+dKLMEFQC76SKWxRBrKaxjPwg2oKg7ItdftKmMBe4PYACXUlCVgQq9ImYyQgX7gjW9Z0bkPMXs9
PdOQEYU3X4m6ZiV75C+0B+x+tV7zRp+GLEE+VoM1G4bqr1KHWCCP3GO9Nm3yKj3HYbz4WHb8GXuE
f0UwM9bGbVZkFgysefn0tceDh3OvhpShJIe24/M8IaN7jaNeJLl1H7PV3zM059R/MwgZ2wkpdygP
2bZ8TrundjxVJXKiUJQ2oAJbB+KCzW8UH6sZx0OVlsa7GMuEgjzrvPMUz2y0jQKXkWDYF5SFPN4V
1d3jGbyXwmUCCEyRSoREMLH3d3lZhMuzwTIznZ56gCW/oUd90+iWogcHsOyoM0B8bKiCFDcH3O6a
BTS6z4n50+ufQZdW+a1q+/Sj4JhkJDkBZlyQFvheom/PP4Aprwzbm2wXcJMPlZAaBUAVUw1pzrhC
Xm194tzlc7QFsZ2Kytfz94VzghiE2rcjxbi6W1xFHmT7bZJKOGhl3xK3UTbwyh8ZCPgfCLtBQFB6
ibrILNmPxvHc0LlPcIjKlyacF0GkZagx5eyePv2Or5hIxbEwpkRWdanIbRbbXBfQ72DuTxRmgFo0
/b3FhbmlgA7MJF59yI5fJZk/wdx5nAt1NWYyxNJqGnCDo9K+yc4k1V3NZ+xnHh++z/FeAmZ0hCRV
6LuDNz4VYj6nvkc4h4Tu0JDP8Q4Mna2maqa1mgHepFdlgdpB2keBXGaVRWnNv4Ko/VcAYlgMeIh8
k1hwGfmStdXpukSG31Y/SLh7YeFrXVJrzk6pxEnvD4UvQJlptnWFt0IKpyEtD71NRvHZQt64biRx
taEJwj7rPd8UYirmX+HMgsDaTf5ebyEf+BJAZ3/+Ozei72j5C+opd4r72ZVlaUsHMoCP5JFPtX8j
zW3upQIVjlrhlGMZGMyw6tLQ0T+yjrXomx5j8EqeouaOpLGqXyjpQg4d7Xq4QqZaRKPGJSiMNs4o
SDBK2Z2jbZw8Y+5SVWnyHrUkIG7g2K6rm7WhwzKHz8cFu5OIcyZ3fDTzkmtbPUAEvthdi+jQ5JBi
UI5AbC0ylA1RCTumWa62WwRa2Mee6JyZxMRAQ40oS2d1NIQcTWEOs/1+5B/WyWqC5UeYPeB60YSc
+CwQ84pBH2UGGP/Ux1JvToOvG90eWZRDGT3yIpAKyYH2TsBAeX+1F9+V8MULehBeakBOoZkN6fJU
5Gqar3iOeIcfmSMtoBYIpiV885lifxRi3D6Vn6SZ8/f1UbQVhIufqVcm0qm4h+31a+oUOwhC8/R+
f2RF/RX8bCnzvIXhO+Kfmekx8UJo+hQk3oXF5TOmxkBFm1iuXeA7RgsCWQM83gIA8ALDKu8pZpWM
qJ+t7ZH1tlP0I9ycezBrAhW26ORlcQABF24ezsTvcOFsZS40HxjOmiMsz5B5EA/p4ox4kw/GTX2l
+75Qj2nnOeRv3nCfkwnpvt6tPZG3qgIVQeCobNOv+KCgxcrAsgOdjNwoiNKKEDmpVQ52jBpB/95w
ng1QznksxtLyePjpH+jSOyCtoE9FDhmjjm07iF9BepvTT8rpaW36RDPilqoztetndu29bEj1oZZC
xPjUM4AkwnyCjGfifMHVliQA99BtNOjYDz50WVjrCkqI1Q0JyMYEzigiwJRUDk9J74MM04S12FGi
xDOfpk1C4qaBgdrb91MesoTNb9O9HsjYVZ4Z9RCcvbYRsfd74hco4WYMsZlcf/1krIQIw3F+D7E3
Yo6k6Whj/+oxMCqsJ4OU+JNan9cCVTaB8A3GHQSx9RY4qqPn5ZD5z6Qqd80HhmKxtJAHn9ESnUII
KfQ9fvjBvOxy9q7Hvky7KcN7QqjbJWd8lmrRHv4Ngn6jXYqXRcvS6VaCa+dRmhnVSQCgcs+OWv9F
wz6dMV/zvj76wEjLHsfv/VC3qF5RV2BK4N97zkKkAgnQN8A4jDCs3sLLu1qR9ZpgE8IBDy6p1xUf
NLd3ZXUBCIecDQwoobju75LPrRAusGLJPvBWxnBP9A3UE82L8+gI4HlvR+UncwVjA24eag8y+7UL
fSTREzWTELblry6/o5LG2qmqfdur1bQYkpUJDPBg45T7tqp89AhSc2sd868Z7rNDpxmZHRGS11t6
vvYy/DKp0ZJuas95Hye9LxXDOH3lwUvbmwzd0KgXIfEwLarpeUp+okhSyBhlZJOjoghBlnjU/00t
UhJi7txtdc8hEGlBffAlBlCJJOXI1xQTvvIiHXCaOtKrvpPmN5kbLgMgs5SETTPoedDt+wW1bTru
gIzFSHx8ozmwHG8JmryTqfn4HJj2N7b+IQCoLs0ZRsnwJfRFAj8SyKK+XnLDUwWsLIl/wm17cJVm
rhOnWhEs/nkQ6XTfRwjRMz4s1lhW6qlW/U/TtuBw0szRAkMgB9drg+YN6GY4mbhnTTiAX73tawxv
YW+rz6pjMC8wAOFuYdIejT7gKcJueuvy6j0APYArEwp4XlVdGA6+ag0CxyCtt65q+UUggpUJqyT1
+d0lr1IianI3Xj/ZHPcp0ci6TAkruLJXPM9TSa85psowRSgD4Lhg4Pwd3dvp71tWX0rAejEi3qss
mHMgOuXqwzrk/IzoWiCQUcEWZf0PwZlwXz6Ge/VaWkrl8PrKQ7GaWblGU0tOjKFbg61UBi25ffeS
4jOMa9czB0FG2+x+tiCTvW3wJvgiwOzN21qrPmoWwVbrOn2GlAzEPEsxvqJAjPeponowGSqpx0VF
ANFqpHyPFOWaBqKv/Dp1kOptTDWQmNvpGuTAaulYwkdfIoDJQjfaAQ6UCdCrr1jfKa24idXtr/OF
pNeCQw/kEw/jFFS2ieyJBD/2d4Gyw2Xx7mHb3WTjlXJJo6z44ah4eHLNTTMDjk43+4ahQ5IbCnIV
LeLcCbJgl1brX4uNTfGCQ/oqdlkymLdnkcPrEO0Nphb0PfnqmzTSp2MBr6KBHPZ3ffmpcOswTuvH
1fWF6nZhbT0umY0ziDzTaRORoOkX+DlWQ0mpshLM19B8nOqJQumXjpw/VAZv3XLcXEYdVqzqMQst
qULACXnVoRwKeu4c1CqNuXiTpmF3U3jrBIqLLXZKy+hG2PtzFn9g8xDNO/O90wg6nYpblWl4C05D
js1GaOiZjFslzPhDtcmNvBcFEzL0USK1x+NCp3Q0DLYJvDe6VXcGXyoAq2YCDOrveZJ8eTkT7FmB
5cEZQrWyUrqcrQ63JN+hlRrmvdC2B8mRzPnI3RlBHTSA3juyjFVBpmBd78xyyyyvo+nE2OIQxiqv
/y6/VfWgoMsg2N6XS9E4NK4cWXH9qj7zbgoTQ8gXjys2kdkscKvu0OjtuE7I2K3AzmxVz4mQ/lPZ
4AitORJFeBiyy0S0zDvL1omzRPWWZjcXuyKMu0do3+TZCANJjZQWgp00LS4LgfWbCIlc3SPBmG3m
NWUGD4sgrZyj2w/WcfBcMYo2ePaYn2cDbkKOKKYoGly6eLmg0s/JQilye23FcnwBJkT+d1XXFFHi
Typ8p3TT2DLxjk1y/MFZFZPxQNW3TOPzO6K4u9WBSK+oDk622KQXVcxLbDyYr7zAbtHLIir/il9A
TmPbft9dHP2efUq9NcwC9gLqRAlx3Olu+1frZNM2E+Hpoi1XjK/KnkOXoqDPkWEH9kGgjdVz4gzZ
/NOOFqdbLwLAc4RiRFrC3tET+e3U5/iNYH+o2fDdUHkLFHK34/vALABX8RUqHZP4b3TvU5UM7SVe
HIBN+5MqOK5iaW+bx+zWTGE1FnMgrjI405X+3m8cY8tD/9zSlazFTWdN5dqFVqUl//AuoKF7Qw9/
DFqbQPbLlcyrKXtsgUYXeyoW5HQd7Aqa9mpC7o+4XyUa8ZN+SJPbaw3FAwoLqwwSJ3WYnmR6xiWG
yq2gb9/Scmu/2kZ9WpmjyH7i95gZyylsch7/W26e8BGGyLLlP+EH/lH5fHQI8xpzo/QW53if7rZC
lMxsGhHJIjdVa9F5yn5s6/zgT62a2/NYbvTlWr41Bznws3h34w9SIDQoVul7sJgCkkuUXtSKZNUz
9dUum7Igz5EcEAYd2DFDitlGQ27LUmgbb7Qi8pZQqA1E1eW4IM7vQ5V2FdhHade2yFU4HuN1azhU
OKTh8/N2xiaumQVLbvYPUgqRhvZTE57MwC+4fQdoHaEA4lYPN+BYlUZn5Wow0p4g3/c+q8SBDzoK
sGEnyU7F8KXkJNJeUCAuxXYjqB20n4odT40SLZxhyntRM0tCCKnuLK8pyXSjdiHVuSGfifwIbwZp
lz4DAYB/bdeDAoDv2PnxRp3p3+caT/7Q+oKJUfcolnKmdoG2lLGMMBSCkINl0v7vNpk2HtWExErL
z255asCxFUlf3RRjVxedZY7joNiUgWVAUTFp+/+6ncw0VfdeS4KorzGCxqkbrq0IMsTzdHSDwfSq
QxiDp7LQyyLISfbMmrW1lXZ5EfnyQRSxaLwCTwK8Zm6ncpOjY7+C6NHcJqjEOXNftbfdm1Lyzwj5
Q5gSrk03OW5HMM95MKi2Cc+HaQjKA5xVkAWKqfGZX1poDQ8i4Npq7GQTU3zVucMb/EpQ6Kn+XpNS
N01S7Z8rADKIzr+ShaOTBBGq8uWgw2GQ1FIvcQ++B/Oo389VbLyD1T9TSsyz5F7LTxxrteuOf7tx
TXt0/pk7RveIOir1hX9mRSlFDkscHy935TgfxbP+937H52vWXhdUbE5nYHJ+51Fh7HoLHM0eO09j
+si637D51op9wBVIEYngtPwMJ292wdd1WFI7R/K88STT/KscWlT93BwRkCJiLpc52Mm8MY3DbWNx
s5ESjlxg/xq9aKWv7S4VDb6UWLTAlycFRkaIPz9pbqhvQAipc1/J9lx4Y2HnkiD4XZHhgP2Hs2sL
DJuOVcHhSA5leeVddnvr0Ohj0trieKrfJ2hz6+WCLKWCshIKjKlqaKVz8WblXcZyS4/z2Z7VeLfJ
QbC0GUxr5w/B5aMkdT1SvQKn7IPMiwcyMG+IDvAuyh9DXsr9LDgHL+gkRaVupxuAvVUwpkzu0qIk
U60hzcdI7doVYhOKk10hXmJassw637B3LOYQjbnMcBRzV/PXrJDJqJVwNaouGFdXg/r/QvnVviNZ
7oidRyFCwQAgMIncyYZ7yL0SQaZGyCEAJUSz+KkE1OxOA6uKYtDn2agz49FAcuwm2bYc3gqq0+TR
zG3yqpRDRKWFaw9ag/HD90Unhlnm4c2EMDGrijCOcfDTEwJzOEgIAFgyEsJH+ckZihRQuftQIMzn
Wlqw6jwDsS2xjRhUt8S7ZN2723kuyY0KZYpfz2jsiUqO4gO8P1gG4TLZGplCzloqwrBECE9vPlLN
j/0Di10a34jkJc2uIxm6uc9D2OK83ZUuvPjX2WrmaPyMAGkdAHhTXQ0YdikGZkQ8sOnx9iIYZla6
ArT8idqAFgKaLzXQIcZihMoYYJPtlVDNVZBJj3Ok8cUN9xByMWK3p9lpgVRX4f36cQPcTwC+P103
4saEG4OIqfoBZQcjOS8YpftQ5DpEKoUHvcOBZ7GDZ/j26Gv7/NQlQUHKkqm84+Wq3GBpwvRf4IQK
V6UlPPL8Bcxq5B1RwE1TdUoTqSGlO6126Kh9DPNcmskIv1zjxmwK0s9goXjXMkBqmnXRCYgzACGW
Qhraqoza+32VRe3Kv6S6o3k64GcI/8oO22P4UgzTYfSZmHNRST3l7tCVapd4ZGoRPWiDaHminBKa
CCzeWvV/j9zJRuOo2VU+3+elEr6AQAocA/USgMuaqf27/J8YpwHCm0zcx7SwiPgu8cKwgS3QCSiB
qTZm++FHPeJegdyJpmPfMHACucv8NKTs/o2K2MZJ9nauuA8c2fupqu6qHzHJPXzjiZMNiAwfXPuU
iDioFQUJa8+Yvvqn+ZzAimQvB6LazjSqXJRMzy6V4k5GfrRAw+l+rvrOMoud08qv9aHw1NFR+YWR
JtoPJqtIM8Px6PEi/VRYp57Tq7TzlJ2q2LGYf6ldNf4+ewS9Vz8FAib3ZetNKCEsTjIHAi2ulhKx
ZJbE6vb6zY8yj7TPKRnd7J+EEfd9jU1geNKjyxy+xnceqLRLjQnGSrlMEl/ciwBLVShZNrC/cARY
5rjAl8TpMK85H/fkWM4byq0O3dhoatRlj5BMTtsmYvA+Z9U9I7AKEovFOF18o9utzc2x7LtXCsoV
0M+FtQycI8dhBLtXsXyCfvK9Kh9HEhoaNizAAIDUcHQDGJuerHcU0Q2X0+h9ZomDYFvP6j23FBrm
KLJMV2bavbe9iSyCFZ2R02yH8P/4y7dIccQUUYmDgfdfGh8HPQj3tRyAE3dccnG3HCbCDdU4IJ3x
WHjLLrU+EUy2BfkoRll59hzoMAetHc8LvQUWlOo9DaPmYvLJBxtWbU9XMEnp5NnzHThEc8qtHBg8
VOnOup99l0wlXEWTMBRx+5NozptahdJL9Mb05moiZnXEKcy7jpkkUgmujMlhBwzWXFjD2cystfjl
9OaLbATbK1VuHqTn3Buf8dcHnxdt04KsDrF6TL9kkifkQ5SZhmGIeC5KepB2ZUG7WRNmFTA3+QYb
NRtrH8YtYYWQAOKi3X/sF21akmH4gsvQDPpxnOuBwwBLZPu7j28IQGlS45T0hK0lmgk10Tf+6gOG
8oCLC83cTbjAFB1HIAx6bw8MUEUMzkAsGcOemGqJp2AZl8/WZZ7VIpeG5/5BsmYhhpmdzD4gQyoO
asCTcQyse96Q+gKrtQ4+9BgfRKHPO8ztVIvtGNl0KoaFhPi4tIhbLyXmh8nJjxy83X6RsrIJBDpQ
OIrAv0gCnXxaUdmEaP/eg0jAcGI31u2PfWA3AgjwlT7Qzbts6diUj0hmvSSA+ykHsc4CnsdbwWbp
sbRebgO9M6JOUi/Ua1TvaswrHPatf1TgLTlkeKomjCeFY94zMMiMxwaPZXjWdOAHMfXw4uDWJ2xE
+bBMaKjD29GEplbsRQ3K16X+u7KH/d76UcDB+ktupDstq0xve8JPNmoDQzrK5epNmpJ9X7YP1deX
cze8fCHUkVlIsco0BIrm+buRqwgASMlK5pF57a4UrQU/ubrl7ZzMEUHM6sUSSOVRPxKngfyWvBau
Ov7+z6i94ShTv9Z9xVbc3AWrQv2boctPhmuuLXM05MBsi2Co+KREuyJkbE9nzN27EbvBYpmMmmDe
oRxM8dcY7bqpTkNPa01rV3hR7kBjBY25ejzjP+mOUoNulV/kZkge89YqbZYZhAIAmXyJkBF2qyJe
yHL3XsrjeG45b8y1RFR+FTDIVi1ouWZSQ4ULODDYA4G7bTeuBZO6KLrctI+QYgPXus1n2bdAy5/X
eAE7vTKlA7/5WAKlJXjXyZCIzV30hYp/iQiiTlbTHmZJ4Y/ymOgti8e+s2AnC59+9GmY05NqHwCE
hOH1RGmWUDJHdSQNZqnSo0W2dIj09a32BxGw3j6YuGQlmCy+c2mh1M2S9GR9vFWDeDH51/yXDPWT
/6ZhvN7nqbAuYIEb21uqrNAFhHJNQjLXFztWxBVX+WBgp6dW11gg2058UylAu53XDBR1nKKoV64H
SKF2EPh7crD/BaylnFtp/ZKteVNaQ0dheswoE1XHmCvo9WUGairXl1KI8APtP6SqF3caDhs1o/Hy
3ad0dihuVFxOKUISRJuy/iv3W9FtBP840B0PXRCiySCe4lhy/Dco/0ML8kArT/yoHo25pWY1L8kC
nAI6gTrf/I3TeWenoPnTmQh8Tx5DKx43hr58iRX2qyMHqkRX/9oAdmj+JkkWuoYOV8Ttr6TroA++
LQDKSFLcVFcfB56Yn6YJeaPucALSNtXbTSjCxuJPqgGygN0qm61q6AUIGCOZOmOri7AyRUyn6QLP
JvmOK0mATAdYyjZSp8dyUE2rNQ61D3eiO1IZs/Xw0XiTpTY+JebvhP9NPa+h89cMgMQf/NGw5y8H
O3SxUZvMvlZ0EYMQTDuDtrYpAxBg/3P2dPaVCiZNr48xgINfJMQejGh0PyZrcrFV+f+1O1GF2jMx
VljPihB1ylHoUYV6bkzj0xUVVssTiLEymEMRg0W11nZkYaCSmiz2qvhsaK7xQ9+AR9WFKLDTKKbd
hfGD8muBIs716NvN/LxUwCvHFR2RXpV1nOH7Ef4xG//O9/YqNJrati7c7cM1pRWeq+RJ2iqWgVVx
KoHp1NVWxNLEzUWduhCqHtFsK8IywbC1BxHX9T10NqIGZdKo3ViY3/Fa8CSmkNzwFKI5aT8eyzxT
9rTZ13BdFgvI7dRbagAfmL9dLpVgMyQ8iyNJM2WWWQu12LeeRu9xuoz5ihodYxIEwg+taB4F9yDg
joBX5ItwTqJYJOBm8e3gvucjXeL3thWA+ZL/itMwpA0TPej60ZxFrx24HIzVMyZuxl9eFtDN0Pw3
O/drcS4IL0DNup1tQrKcWqu02ukdGipAbo35+8B22u+y4TzhLgfosrnnuD2OqURBEPk1B7IxwDL+
LtIRsCX6ucUxoF0595OszRAA3RW70qU6oQ03+Dii09wosbCoUSlFf76d2nWFTFSd2Bdu0gNYNi7e
D30/ugP+yaOPclt6baVOAiEah8k/CUzgRJNqOURKQYGsQX7NDhC/1qRzgk6Jx0XcEeMqfEsDN31d
QMjk6nM0M3G44Nx/eUBn6vO+L4jgRFBnaQTTp2JR3A0MrMlFZzDHhViDRMgTVl7usFZEmg99XgHw
hBnRZqfG94lFL3Wg9WOpobtiS9JBGWHWyurSMpPoTgXfDpvIy6/2kDPWpWiI0M08Y1RoCSVVUBCO
TTT7NpvMrZyoMRr3AhFWBNq9MrE2l8qZ2nzFoT0GJyCHnDkK/0cL9tFf0HVRPSAEvJLnJIX0WkXI
MDG4PVvrySR8+R7yiaBrHgq6JbUL8iJyKXmY8SPBvhymhWbseJeqQOlbXIcqV23XZVatqcAJ8Er+
gGSTxhjBwml6nx/9RpLrawHWI7BuDCKDPsmRXMziQ1f9hxkhbf6R+ZJ+QOa2OmY3ID4kdSAn96aB
k8juS9rrvsOccThne24p5h8kOI7dbE6DnQsmGjQHO1NA7f3jRTOLCMPeYCisc8L6GjvVkva/yQCc
1/AwimRP7ZtLNT1M8AwGgbRt20f0RlaD0ih4MQVP421unO30xgqTCxVkXyvKpRdYUrNaicwKjTWD
cL9gK7LXpWPGtyWUWSVDHk/nyl+oigx44n0Rhbi92CxlETW9pL03C5bjiFNgoxNdYvu3Ff6gLLqr
IyYBruYhhaAq24UBksN4uxlFAh0Hqjwlt4zskr4unwbnKIdcAMz56cXzDsUfx5we1wtHNkCOPr8v
+7bOoaIMTT55imzXbIplhCZQl3RKDq4hCVudX1oiL7Aa/IWMqIU8rhui+rlL3L59eQW/7xjDGgGH
UknXElKrR5p+DK7b0d91fJXg+3Ji7oq0SNXdWWQT4qf8bQkqwaArt1M4REy6/tV1n9rXdJfPhSmR
sDx8Hh3SYIXh7sziuLAv4Wisik2oBKnA46uXNiPpoIPzwoUn017abEW/RSJaHa24a/I28tFsVlkh
LxL8ODj+u3TJC/DS7vR8bJqRnbR2ff7dEXmY6y2IlXmIeCF6fjOYMw1kPsWXXJqCY3F+wjlCuHSt
jCymtVE7u4dw0IhP8sS6IVZyMPqhmGh1y7/f9dZHlIvHi+h48TjRULElYPSnBzLizrq9/mU6z8V7
b1lvDdFgX6jO7VWd2TVkvSrHruTYljbPvqO98ESikuDNezFHivg9vqTGlejDpBE/2zRH5h8Iw3sA
l6oBesbFcfjmknI4mHnpCDAvKHwMDSDPKEip+GfNEuj2NCmVlrHeZWChfhbJJ08cYycFfkr2RXaF
eVYW2b0zB4liOFbDghYVHvb5y1lXWoY97CH6/UayAZ7rTQCY4RNZFo8utWaeeUg0GX1a+x4H4Wyn
u5H2Ksu9v8Jbt/G4thAM7PLHJjOXpynJ44jy8CNWqNEBkoTW/AZGGEtD7xjtULDG34+l54QWoqXR
VXoKaBBQlM6qgzRu0M/mQpsUYWbMB/4wUZzdWhGMiuRRt16GzVd8G913j4J9zXaIqtoal9ireBE5
NEwHPV5KhPRmjylc8w6ac7ukbLd6rofwuinN6fMuUuB7peTkrh7XZwj7kd+bkbk7gSv4RNIs20JA
clON7/KJWpuq1V60Dn6rb1czowVzROOu1MkcNcvUm0cI4MXfms8XN11wSZqZR3rW05JcXOlUFxRb
tiQqbb4cNh8TG/PajJgiJGfJdHE8mkFA1IeweGoy9u4f9KjFpcrnUUB5bmZXSEl67uAFASWbCZhO
WCJJnLBDI74uvahEQsViA2NNPEjNo4/Bv+sgHRrPQCKl/VinSCFSHUHQZ/Yswd+dFz2iNeQtIFNw
aMurMx94p7l/RrNVpymls9imndiXSaP8wwwCdJyI0aZXO7h/5ymX5oqlqOWhEo8oHLaaiSASRzJF
MTiftyuh7A4oYw56XVaVv8lUHGSlv6OZ+KRhvioRPrkV0OwTjhT5DCusFhr8RiDp8X1lxVaChWEP
EwXiGZhj2lRzwwsD3uNe9pQGkCUK2jAHdYjwOhRlxgoEWvRZ0Mw/KBdEcRR55qBWXDzaHUHOwiKE
kCt1YK8g3oWP1mXUL2dAaOn76V2IF3PZ7+1/QjG/akGSRPFDQx9KjVcSSk+e+kuW81BsBuQFl79W
C+A4GKAOQDC7SGoIoI1hSrzYjngOhGiMwSEiHvUU/5CI0AQ7i223nXzSGIMTjl0LDYgbtaRBy6hT
NZPB0bTCkZlOZw2jb70G5v1Z3iMruXCXiQ9CNipN7nIR4itOAUTx6NOh4+VpoaaPFBZcJLYU9WEB
Rmjvj2MO1vk0S2XwB7jDDYzcLTWV7B/4sVR2f/hESwtaVr3hd1j4G3WF2HjeYyRSyM4t/69KTijV
F9CwkHQhXx24i9EZUrGwqm8DgKISS6cg+5z0cBw6Sugc2d+Xu7dtNMtl/zQsRa+9qiWme/jE/NQs
zOjJFC9TYiy6Kp6NxcQ+MlmoARinKUP/zp0VLtfXBRKWxYAqJwWvWDGtv/Wt1NMTT5x6jOQNWHG2
uyQKBGlCBQULUl0VYUWqnh1OlmJWPAAuJ454ButvSO2kDVET0fdYmFiHH+32qOTFtCCxRQGFTlpI
qDVClKknPe5qtv+BhOIOGEvFN7XUT0pRA8HZcc7D5j7zN6vz05xC3RsZeD0PgFOrZPHl4iHp5PyU
DoGNRPmBjlOabaelEwXPHNnB3rMvCwQPZLs+5X/kYneK7Due73fg+T5Uxk8vJeBc33c54SN5Lnvw
Rr916zxQVVr1WYhSRv2bzhL1JZU6xVZy36B64k2vn8hb0Nf2uAZh8HwNCAbp49pknhesZBiEgD/m
qpn1VJ5UwzhQktzwmog/T1Y/ep64l6Tj+sU9QWemFqbIs34FBIAiuze7f8vfPWWzgCKo82NOeabr
+NvlZTxN+pG1noGvi8fkQ5sUG+z30jhhl3sCgU/iFvRTy0fDEvL9iGgqWP3zd1cZVtEAXEvRAivp
nYc5hDCKd16vYbGvKUB2k1QoXkaO4do25LWfPvGXO0yBg8aZH8AHDZAEwJRM6K9yT+mtIhqfNR0u
DN2uccOWEhDUDwWUERTsWpDYVnqipjLHvyKbjl7rqtsb5oT79jOPeTvMzXTjaUeGbFOTWUQdYDnl
Uu26wkLsWYF09AcXK1eEGhLyx3XiFpB6dLOdpTzO4EXFojko6qaRxjSLSt8SUDwLwc+JMyE2wyRx
agfXAmDBBqLcd8gKLmgdlaKrUTOa00WuVmALoa82y87J8fPMho3ofC549rwSIAsPgo+tLbdYkRrC
RQ5UlwVPM4WwMN2ouGXwqp1H+6FZK6iCDjqjw1g+x1KpIZkIBta8omDF2quAsSVWjLigOdXyoK6J
ByhzcDDWVXgQc2UZV+10RPSXv0YRu3ea+e7rPgrGWW2pIFDQBSndXNJ5dDFJDxYmPtcGW0c7U13f
4qYtD/k8gQK/wHgG3lV26GthH7ZXE510WphPA6bCGgMBuypaX71lq0kXGrJBdHdfIB661wUQmzIX
e6IymyqvlcSPPYV5x8OiWPJOhGZ05asDVPbEtAfWLrkvvEp0fTI/Cl0VAHzNIjcipfyoYGNVzwyP
eDS4CAWDuwLja03aI+0ijBJz3yV4JbyEyS4uXgyEJmQyTQlhJM3gBGPcNuP9wtSGuoWx2FFNWcof
nlq+kJydC3ZXSxawkM7qVasX1k6s4PQMhDCdXxho+BAuMFpwiwknuPFcndGIaoVa4rCtL4dpjk1C
o+EObvahJtwAi5lv4ApQ8TgHwL1rLOXTBqNpzixSjv0ObiCb57sA/0xSX5rEMl/sZr9wukQAYlfD
UaOs9tZ+UpJpEDG6rRd5cU/aH+wsgIpoDa3pT30HAzPqyD1cfmJxUfIWNtbML4zkP06mgMKBX1+T
dwdcva1BWaugRUyduXGZZ1mm97nmkMJdpuj38WsuNClL4FyAhL4Tfq3ppFnc65ja3tS5ObpO2i8R
kQ5zKmjtLJVpiSsr6Q9GRnmnIqCFElFSKkKGErNe4sVHggVvbhKg4RYg2pRZFWSOoCUIll23G/ar
tzJPHrB57vv2tkyuU72PZNP9lByDcBYIob0DDUJiAU4CzUBJulTGQL2ljZLo0SRlYktPiAQzj31S
hPBouigZeikCISKCm+OTFOF5D3rxhiX90vY/pNqTagMx96KaDNRPYVY5e2mpk5gT+vsaF3nktQyQ
phfCFyJX0QHx+QRTC1FjiWGyDONgPvCk1JljArgiUUcIMX+R+wxaYsDC5uJQ8kQBz749YEfDoUzT
QHYbHr7VseVuIRs7LLWNwW9xeTBuT/NU33N2nB6I4WgVKKgA6gaEgQ7MYEz8WG56dhYTD5+zJLRo
iczMDxor8zuQkb/btvGvpjk//xkBgRovVsvZBuDhZj8T4dsRTxW3NzD62XFwn2lZ2vR52C/EMgIE
kxgZHb5DTqq3jI2CiS48hztUADpk3ac6MSd9u3bKI2eHxFr2Rjl46XjyeYLFa2S9KoWoSN6h/1g0
wdzkvc981Zgg0M/gWQze02OcN+kjRg/+OLecszPc2mwJnsBO9UI6uyzmGUBX5h+gl7rGF68QC68N
mrR+/keIQLyZyOmEA5T7OwAaMrzLrQDCw2polJKkRLWB5FaCV3kIpP1yQ+88jhiM4irNWlQyULkD
wAUHeOihNeNPIJkIyTLygodD5QNXTAqX4kYQZNq4ElwuOX8V6Juu9u7rAWGS2Otkp4ulMaLDADdC
iugAa3SUxerDSY4McCHpqAhtiRCofBtiY05lvu3Brhw8A3RU22FNFJz0mm+Y6FnD/2ij67sAfgDZ
D64reNfzRjU4bozU5FCmUaxBP7klr3mMj0VnRZE+4DS1yH5QTCqGgaOu2bbrL98t3hZVgXed2zm4
d9x9rolheQxVFhtS1vPsv7K2lNPe9RoHGP2K/VHTsdeTrsanTcH1JTLWqAdZxo7DSo+UqA3liC+r
8rqehBg9XMfGCpNvq4fOp2aA6zbYTZI7eLxKER0fpxKZ/uFOxt013l+dBKV1GMTaMO/9ri+4ZaVW
HytZ+R48OKvSCoi7+hINI2b49P+IMPG8PZ/CUgz4X0l14cI/gSTPU1pYP5vCwTu/4+FEM5i2F6NG
GFBKayTb2mNP2oQJx2xJ+Bj+iAVJPBQdG1dIyO69zwG6nBqODfvmzhetYPzrwFmXE6/tngz1tyOO
2QOPG5bjD4TPCvhcPA/CpsC2waP2C3p/WY/Cb1mi2DQTVv/bksaBTCUQXPoG/Wtn16LsqGA7m3pB
6VwKmkhou2712tZPXE8dkzQGVaau7gDhIhs9kE5ebB3hxmqfEX5Wjbcfo0qV/FwaDeM/ycl/729b
KhGb6KOefZh9LVkyx3n4rYpQp3LwtydfXjMsD/KYqaviEJJ3MJbaLZnE/JX4jbmMrByKbxXpCBeA
u/WOVoab3s04FQheAM4F81+gWTEDJhEqXkcrCT7Snm8J9hXm5c1cJ7ciXtyZpHPe9PN7zVkUNrZv
Mn5UledeBBLRIFUmIgglq3UCa3ToB3dUg3CHjdSibrBugYyAhG+sawtTMPKb1LWz7ugidfFcNTSu
WcdnVlFcEXPjGcroCh4bXvOPNZnJzq9RBu/fk6hRiXg/4VdjkpP+ALHDvpZ5T1keow/SdylR7Uro
GEGNzdghyEpZYKrl5M2uSwpqk9Ffu4KzkndxmBRaNS9FY/0UAIY5a4JwlPEY//oLq/oSvbFXDEGd
gRw8Ajyg5tUTnogKmj/zc9WFWf2GsLHzeqncTgHfxRyYKLql1xvJ2aM2jP5vMJ8RpTS8mptcpcOh
7nqlHSfqN9OwQ4esHK/h0zGxr0RUGAEuz2C4qd3E5f4joPuAs43f3DWS2DhteWgzDPr6FZ/oVqdk
r9NavvN2gK3wMRtCn6vBzcya5faD2jwjcoiSGqVL6sZtoPdDL68GgH3aZnL2+a/YFOgPWub8tL+a
X7X2VSaNxhuEhe5pNS/uD8Ua97OmH8mMjgniZN+CAYrnfqMjon+fpMch7Qu0jJpm8lkvOyC4j6Cv
Jw7eYmglaAOtfTX4QfaIv01GcX18Lm65EosPyNcrh1/J2ooh1w/behLOdOS95jNd7qmbvFNhMz4F
R42mQeCM5dLzvrt4JVWzxVDedbND7Ax2NHImdXZTfA8VpUw20xZhiFPzWQY1Rkwa0dBGsuQQPgOf
Ri9JV7ZwfeKAGX1efq40GsZGBIdOoNW6bUjz8g8sNmOQkof5Ul//aGqQmrt8pCyUVi82TYHSeRQD
nWJktKKAYABtmj532Nw5Cgli04zuYwwPIEvgol6px8gx6l6kWqoeuDxA7cRL0ZD91/q5ACSK/9k0
0d1ioj6ZK+sZbj7am13IGB7KpJVI98aJIXSV8V5JFbcNmTveOhDCeJKmu7EtndwcHscCpR5pmM2s
Slh2fAwlh5cuUXIWACDJdikg2H+TzKT2tSfZ2VbJbPnhV03E6+BCsgpam0Oj3C+Wgn5J4JlBDhSx
sLSGLPvfGQLcdL9rHEvTELt4rDI4U8eaWMTDiQ8f/4RdqBLI4Z8HLwJd6nrclWiuMGZHgQQAnSlJ
IpHOW2zrffI7iGjJ8m8vC9d/cafP4Vjro0E1qLWKEQCoXCulzACEoC2K1CF7ipWK3DxbF+1fTccl
+bdioVuoZL5raoogDhflwrWMpkhD4V23IPGir5eDkPVT7qEMg3Q9Eco47SjdJsPgOD/NwR/o9AeB
PitWq17g+sjnyDH4N+88+TIZny56kQ5gfhOTxppW5CvwM30O2XrPxd9d+pBIBRwFsW9QGwMdFCgi
XO4I2symKsnUSabILBX7eEyL4l5aLw63Vc7TEEDFBkWHrqYrO39jQwG33klRCsdTxIwl8r//vdVC
HIsJLzA4XAUTWYY5u/CvNn3kbKXEg1kgs+00HExcP1Q32ljBo25HSkTOD3wR/XfRaNcH2jAmUv1G
WBiLBfgU7jC9JQmurOcAYPdEvy6xPswJqxitrK0htM610VgsBrPcINqo5SI8OVy8AYgr9IsOvRUi
wI8A8J0swn+h0m4DqUaOB4t3Pf6rD+xJTCyDFWP1Y39q9r0uACj9/ODfs5ALQldHuiXX6PBigsTz
dAGXjS32LS/HnDbSjhf63fzu72H1+WNJW03+Yw7ZLqZGz6hrWi3XkzwxyRZYiUAGlIv/3oVWtwGp
pGJUHVJecBqjxmplFSDeRXj22p4QNHx8eNatPB+u9IsGmBhabeGNYQs6HBl7N9HO85zp8zHJyvWP
2r/Y00wt04qeTvTqn16TmGaWAUadGRsYnabQPPk9VT0pkPMd6TK4HsLpmgyiz3hkXKuxy331iPEw
KPBGc9v3TGnf+J3G31oilYx1uFDofkttmCfGOpXPyJ8aoHGWbiAfHfRlKNRcnq+RIzGCEVa+Gz9k
tIcfwAlCgnEaPYka/fqtezYnqQl7MiW35TQE6iEoysi+1C+ByNjl22UMWa3X9K4wUvn+sIj8Nfex
G3NnezazsXu0s4qxsaL0q39BwG9Aimgy84xPvcjoWthlBY6qMDl6ol+OEiKmS9nlV267aiVdQUYw
iZYxKlNwuvDuWldg51fuDuUcHWIN0ELNftI1BceedmX8tSWEZM3sjQL6lnb+PYSho2R+rwvTvtEv
AoFqnsDlpIXaAxOaj94wfxQFW3AYOvUxL6D2ezqbXSJ9lyjO9t1ZQdrLAOo2sUTviii4PMl1L4Ls
4IGBxlgmPMX7Sw9pbI/GcAT8UojGXica46JJAAJF+HPNuq987gEyrHjXrtnqzERxBpW8kjFYH6vl
BjCjSKIktD57erQ7unXz/wwuaZ0lcxUdJt6o+Doo08mN1MRFcAmw2G8WlGItaQq1gmq2zGZb4+2z
dNzUNRK+bP5PpYY5Zu4utaJbS6uGV1zAupNHkTwC9av4iDn0YMQpwhJWwPuletauu6xztbY6b+AC
Lkr0bq9ZuF9BlBZDKFQqyw/vLc0agQlFb2OK4adIR9HzYjHWt2LD0u6NPMKvq8UgAIWmA38hSgHy
5JFpPmNYesWgchaxT7GX1KZp4xhZ8x0S2VmMFk2z+wXpGWoUhcPnfO5ZmmSHE1LL7YjN15LBy8TJ
CFOBJ7lflvYjXE75NOA2HPGB3F/4p6OL6T/UYoHrLtFqQy6ElBZcP9I7HqpaubtRvk4CLczkEPLU
+z1oGkbs+n+fN85WmA3/qIuxfjwle+nbT22cxnL1Uyk7vE3a6M1JXTxjJHH2ZSdZR9/41IF6j63O
F1W9TTpkmJFvx13phQgwIOOqPLRCinfOoxzZLFJjpVrlrQ7mf5nn5FjMGfX+bbeIQ4DaeNX28Mtn
dWdlWCFw5WnnVk0HGV2leBfhTFWTptCWWe2GhFMRpGZnYLdh0FLDwMy6qvvm8YyBMJlOWVYzYAhF
I/LAeJfPWSHBSVfFgYsPvGT7ChWpwpB7iAnsAlT5uYRF08nrS+oyNF7AMYJdG6AR7GG1kBQLq2dS
U/wPOFcRz0Y8swCK3Z18yLXVl0QSibGcwc4PqgCh1VWiKUGytyw4RC7VCmWMklnikXQUuue5j8F/
NqzUxxzm4mgKB58fI4vLOHiSyQs9SgX80ZGpw5IuxyAN4JmmLCr5yr/pEyRNf0hyhbaI9RgiUDSX
qLauNG4Wny5EW3fGdTHWay80m1my7DVDI/IH4Dx7NXeGRDbSl1H0QFnIJBh/vZZiUx1OJyi7QauH
/quca6ttBOb+vOXgfVBmNND6j8TQo0mDSH5Y2HXk2bVNThqKRGPcUCKfuJYhJcc5+8RKoFNvxBDM
LQYhAT/40ZTo6eY6tUL+61RLuv78RL9PdN5y/SRDq6yGX4dRPb+x5Rh8HW/6S7z1+02Jp13xyqvq
6qKRhMUGmFSZyig3e/7k1dkUJNhgW+YspZz8cSf0qBmoBfAJ0YkrOv8arUt1EWGXw3eZgkxTrnIj
5o8vGCtlPaMMIoBeXcGfQx07vl3NaIMjFNx3P8MR8fmBwoP0Lk6CPthSjFxGxKfn6UrDt6UopT4x
PH/aBn0erl/S5AuF9EuBb2qJd4o+dxmZVzDKgIIIXzO8+Hq48p/Bdj5JJEgXL3JHaHblCcRF4pJ2
GZ318KYZyKB/JmIZO8yegDU92T8/9x5mlvbSghIpgEsmc8/7E/V5ogzg/BP9H2wt2j5+vucqFqIK
mHzpyPyIhHnejAtQ9EB6SB4edxKbh9kq5rqvOJgnJKWeCmhg29kv7HF/LQ/3yM0uHEYw9mruTJco
VrJKbnND0AWaCvZoaZPn/bPRoYKj7WI2xrlZQOObj3fiCUxNLKKAugpFDKkJLff8781EJ36B5cpM
0qlJX7ZcwOZrIxt4GUycAY5jLdDX7sBaWYT+U/pVYTIQIXwXNWJUHqfq8oQlQcm3a0X5XjzbLoTi
2KDdwZn6JyyxYLLjWmx1wbiSpFNRUVft65GqqLBxM9AqsD43c2e5fvwfBCZ7DpybnyiFuhsuAY2K
17gmMl5HsQb84GZtD4pKfQMRWiHqN/SRQ5pZm9iUic+FHM1oN8Oo6xAdxbimKHQYNry+RdPIXOBP
jlfLxZ8F+N0C7+l9rpXz3hH+HN3VRP2zDAmReCbuYlbk/f/gu33RSK/MTJOLVdrnuGBGAcA2ApBa
UINt78An71s/bs73cmR0Pgcth1nLzS5OR3tikwiJ9LC+xj6lsIzYnNGx70gZLzUDwuTyl7zll5kh
uRofcEWLK4aq0AH5MdveX6LY4ZZeBWi+2FMc3UkG9jeIh2HEri98P2mft7zI8gGCeMQqLVmpRSrq
6rmQxw6ipaKdq6ZSDd7QlDl0IHc08HNof4r2frRmMMG8R8XJr+MFE+FLNWnEFHnWg9o1u1WS+10r
VtmiCInXaM0lpFhpiI13N+RTkclhEfwzYQmKmnAsat2BREiegm5WGgyy+TZe25NNLASsj+FmiQTv
6yWju948FEQAks5EjD2kGtFLV+gehIjIanP3bVFBenI+rGcj9oPLNhSLe/K8teUdCuUu2oA2MyUc
9aUoP+HAeDMGQBlSpXqGUgzDvYnYNftxpGIBfWSBMPpUBwtpHPTfjyJh6IpSvFVCa0oFcqHZz7sr
1TA07jphuOrwbvu4e12N/2jcYuv0N2232pbLjsO28okTUMS0H1ha+3XwlABEhxWtLi9+Nz1tyRc+
MVA8m/bJXQxqmBKb4rCSt0Q0JM7+lgaUoTvpb/ODWHKlhu4KIJqwdGme0TcBY4maExYdH2h3c4k8
tr3nh/F8a2C9wCXNLdclhHeZpcnJFLc8WOyTjSUtMRasHFqUxG8XkePxUaKMRz/dj+QI25CoP8Vu
OIyB8ZsMrpnAFtLSQfs29Ot5+AxIklAyDF6MMImTGPXpckyCRFnJAHuVEfMYicAnLhDcXIBuDc9K
nHezEI46/kjKp13uPGKGXPgxBTzQAnRZvpvkSCi3t1DG1mvOCBBdVbUaq3/2Su4byP5Zx7ugHROd
cHBvFzJGBbC7Ps3outFc7jnCEQ7TUB1r3GocOT81ONas/mP6YfS9xlKqfR2sXcFpTgOIFxZkkza1
io+Qc6p2BP2VHvNIrTGDXaaqAyUOwOuibiq+o39igudviIpFCqqrAEquxAyeFXoZT/4RtzYrRug+
6nTdD6zI2BSHqKJ47Zed0BZh/ZYtbtbetnjLy83koyrVT8y4dO50Yl2wY7xuoik9+ezAl7eaWq6a
S/B5y0dUBk9N8zDcvc5JnkO9Y+hLHgvNBqoaUaZyE5Kbl8uHGXYxgunjHi8RQk/Y4SbhsLnjVCEJ
ImrQyqYrODvx9e7j376TvgzcBNvY1KBJ7rNUj/I/8TS1xfjzXggTd3VKt9zc4DUQNF5PLZtkBifU
DY3qU8HZ7fA9lZd0aexvMfPcrLLaQXnZftKEdGhrdULpQkzNi1Tq4WOoax6Obc0x0+ovf8b4DK0+
S4cX5bNP2bUmriKkIJKNJmZw85h30dHUQNauPf4QZiYh/TeqVPRAcXc7d2rP4hmTlyKWXpPA+ZNi
wrUHj87FQI5teDixql3yXuWDQ9kN1AEuKDbBqP5WJMUSV3mGpC8o3YxAJ8vnxe7H/0Cm9L3x+aGY
Z4uEaKBYMT0C02tBS18Or+Exy/Q3wvWGNAUfwJhcCnC4Gy8FLyiZkdCVwiOTsMKWZx9ibGKRC4SH
ZqCaOLoaxEjPJZIHtArUM6uPlxD5fsYx0mhG9bcwWlr/lGnZbxKXG0PmNpccZiD7yl82Jv90IOHw
S6XiivQmd9Bm/+qtdk4RMk8WvsZAjzk8PmEuUtfx9HIdvm5Cu3CvEknIHyagbWWDADYqtXJ52dre
qSbwvYIKfLliHihqUS07lsYPW0AneOI520cUJpUzsylUeeK0xdHTF1n1jVuthhcFFzO3eG1BcoSM
tCnh6RiJDgzWKK4LugwUEM6EyUymY0dMCf7TUBMtPWvYaIJidUZNq63iyS0HSIPueOWWZ9ct8obO
mTqol88OBjwx0JA/XYjwweKalnEm2AUokzHVRL7zFlGyKkaksw2+0JDd9VALLE4D3vtLMq59uPoW
ltVgdATHVK9jt/ZC+n06rmLweB6CU2WPqT+GAd/n22RqVluifAofFQxvBQ8vC6OnWoqil5vpYZjC
KZCYX5/Hl/fp2UtIL9abtd/KMaigk28p5RXpZokJovFoRIty7jJC/eLrZ3Ux/VprstcsU5x3NMuw
RyvDzFoVZZN4PoTrPubxPxOly5NefRM2sPdk2WM5NPmj31kBh7C6N16iNLqbmotnxEIw4VR5o0oY
QPAEA2zJ5ws29R+oTJkakpWA/5VJKn6YxKpwAdO76nS+9inZwUiaFMMoXKjIKHPhqHsdEs07XROO
T23Y7p17Zczfw+Uw726OI8Lrp6xttTXWsotTgJGhoeK3yslN71e0Awjsfj1/lTk8wx7AcXUrGTqy
zSCmA37i1DJxz4DVCw20DmPK5v5pFsJcD8b9y+Si9NP2Dl2/Bk4jw3ZUAVv2UPeWSnByBhErrVU9
OhRiwY2NxSSJm1P7kELO0gQWwxfi0RkG4Qu5DJ/L/OfRiO4AlXrT4IiCLkYIww0wHmFwEz+YzUH2
c9DekynLykCzQnZxIJ2Id2ll3lFnZkpbp+/4jUg9nvkKCtigpZpwtcusauQSvXZb0Dq8SEeZAoWX
wopZ/j4b9yGvY3o/fn1Dve0qF9EkTGiNKIaQvQMYb9MwZKB2BRfzQhJlk+c8SZxudZ8F750SQoAA
tDPshnKokw/j5FMVDLdrw1330smfHdmVflhWNuAq40ddRQzgScjkU92iueOIoVdaC511plHHF9J3
NyUhXwsj4Sb71+Xk/3P4KL389nqp9ND+2Vj2WbpA09anZjpTjJFUXLSdX9mxx8yQtwfpUYyQ4qLL
xFE/i5reh/KxS+z1Tklx0amGJ2/UpoLi/4WTRo7NeTNCGOSEHse6sxbHsxwszWXdtSuuZgamfohc
pT15zJagoiro1Rq92ho5HXVlOpGuUM1ilazWP+90kQR3c6rly8kAWdnQJ4SyOdt5e3Z4V36R8FnB
XrUdtspxFtf4vUDlpZroxFhVSWJvVZ7KjlYpPV1lkWji3oEylj/2XhEvfOd0w7FAh21gUV2afHG4
i3AHWBuC5gEFY3mZn4apI6H9z1ylPZ4CzTbkFlgJyocvBlHpQEEwoaoYqBUmtU4PM8yt8RVM7Gt6
V4nzELnUX6IBLlongkIlHfNJl8De3DEWZwBwS3105oMVdku9AEpZ13MgcqVnIINwVSbGjpLfa78U
9yOU77d8BiH5pbAA5x391qCVrCb00jEGI4R35Y+fo26dIjHbP8ZNisgw+XCVS0KIcuX0UI/mglBK
QsxO89rfAw8AymcrhDL8qsHicuyn3WhJVANntp1kkO29offBuxVUTEaFAj+7e6C+pk4V0xIM27xu
rmuiKHyEwPkSYumdA/H9nusp7ozPAlRc1LmB3FHvniOpgKNak/58EMqVTTgM5bWRKyvYaHgBzxPX
TYFWHM1f9Bwqv6tcJ6GiUmC9nU0m/IqCQRiTVk236s9zwbMczN7O1EBQ2MY09iZK0i5iuFjYr6FD
W6BVRgptVO+GYdrMAJfNGLSuFGakWrfcyucLw9AQINhyfsDGJUDfmwAPmLu32OhoLusM2G5vPAO4
+/2jOG2yQpKp0a2IWOiXKjhIlAoq0O0FrkN2cAEd0Lrkb0qWNhTXMJ5axoisZ9gI9ZRKpLS3lUkS
8P1lhf0N+WgE81x1u1BbFy9PjX3PAWsxnZNCUOrqs329q2r4Og/PIwIqkJRLJuHFuCu+F6v0frLU
5EP0kSJYWXo8VFIhXBPGzgAS2KEGj+sTUVIPjGBn90V0jNEmjeYpQ6iokBDbFDhUii5eO/0m6N5g
dMJflj3GPzMEciH9ZKSDsA6m7/mq9GFUBWPpdiFQ1iTeoqYcrtaf81i0WWKAZUl3q5K527MyBhhx
SV0Sq3gu5eYs2Vp+XHCbGRYo12mgP5DkpeLPg3R0YFyiPW49FXPGEmgjUuGyiBntjjGL8HVYYnT/
ubYaxXt8N7MNr13pSbyNd7i/DKROheuTFbNcci8ziHBc0xGqRUufEQ3g22CknUtg7X3fCKHRE3mm
glnWuinMsQ6AxH+QfTAisUCRDLRr+DTADV9Gjg/jf8JlZvWU9f/5cwDQjeMbGxIX/m2f2wZKaU3o
j+iR9l8mPJlSIIfyE08OETefzppPXUIOUtLWmK98lIWljnaiSiIEp5GG3a8RGhIBg6o4K2a4BVA0
DD3Fhrqwrb6b0UpjIOLXL9M2LYQ5md0gyGz/mQlzVrMNWCcLrAEJENk4+gb1p7DcibdD39KuCozD
ybYS0bHpMVF4Cht1PWHwQxQylEqslyNk0cHodVU6AfH/kPm/bkBHi99QYLGOiJM6/x1BTeyd2lUg
Ec7ObVW1FdFot1aXmRSOA62jsJeMHjn71hHoXOT1qxiPq9akEBhA7cYdztTECTha0q9fDFji88Yi
tBb/eExSD86cGg9Swz9DSptu/m/xxn925/Skar7mNBZgbMue4Jebm781ibbX4KsZ4vJwyYJWZuWR
++cB3+XVkKM9sw8IEy4rIIISniUE3I/k9KYXewebqJ121TxwpoWgvY6MXCJELS/lFv0tXmGq9qpw
w5e1J5G4Gb+C9EN2b4AGDwMtekOGeUE0U/5Prr5tVFBogwGtWXZHxjuzmFq4NLEphUIfToMGYwtI
/4xo+WsbskbFFo9Oqe4LC/3yNXFdYbS1iVb7stOgjKXde4AEGbcCKbd0YJxrw1OOdX1QYFvMFGBf
aliCWLZSJoVGHStopU9EwqdcA0cH5zSPD0VAID1rq21d1FtEpLSGgr/lj+2FThdpbGt1WpyVMirZ
OJwCJezWnUYumxnVld2NGkNGwFmnHvvT7sMoUplc6Kb41dDlnVJcDrh16PkuWjK57w/qppYu7MDW
uj4hGmfxFU3TXpD72eUJtxmKkudPuDun5NdSdcfAYQd31Ik7JWvE8ZpY89czg3ZcXdhBrOqhHC6i
hcUpmXUcRKBBqWU0kO+FcC7W3SPkozpIP4eo2Clel4nR8+P/AhNgNNhlVDLNeKVPVcw1MRNrB59M
qXTowQKwx+50+h1Bu9xsE4207r8YgGGHWJtOm1VzMdekyDJ2AVjsakC5Qj6XugMLrXwh44EcrZgi
9cEcFn0VPziJWpq+sIfLsP9Ekjkc9XOkOqs1IxyBpIGd/aaXQmnscR3P2DpoAhKzAxVMmTqqw8zd
47+X4PfmDqfhkfmCr2x31InYT+dks8DsDJZ64c2jxmAeOyxJvSgk30UT7D1LsCmmuRAwQVri8Uov
rKOeK+ycqHoW0QVnV2clbeI735RHZqRcODftWM6TTGYDlxgfF99xcYCM663SqzuF++eZPOddwNjZ
5Wt5NH5VuvVKIkkSXM13obyZJFwnD050rtoh2FB/fzJTV2Tpr6+DtITa+OXWDYcf03xisaEluZyW
L+6X08RBS3ksKZgwGKSj0SdqGqavmnjOryza2yutiDjpNxZwjUHfHnAYEaS5V7fwF7s8a8HRFLK2
7zxrQsUfXv3zvXsWrkoYtuRhnC7j6GvWuc+xagt3wF0leoC91ThyHMy0159JRCS6hKf+UfxAIu67
oh1sDbZ7jVdIUCbzanPS7S+3Bd7bwLZSbW4QLk5LJt0VvU1pi6gqY5fezWURpfCg2Lh4Ji68W0iW
oKMCSI2xVOgL029r9QHJR4lUnvij1gzxXUAdPaEnYJ0lDDglb4yi/ywm+ueHcvcNGSJRBP+AOvwD
ebXdhvu5q7JektUXM2BmUEDa5m4bQWx2hNXpEIkKB75moa/4i95Gc9NzExzJJPhZRuW1iXM+bqdJ
ZDhmbZ0qzpsv6p5T3RFVOJgzJGLmoY+W4Y6zUWYP8RwB3UA78y9yn0WzpFuBdrdIq/sP2/I2Y+Th
2zH7Ix9a9bjOFrFn4EP7AunwFz7HPkO6h/YUhIy7lGkzHTNS4HnY5yOd3yz10h+0m7cvd8kYjWAJ
5xHQIUuD/f3hEQZhTh5Ly8Bah5XPfQGxlHvhFLW7H/dunLN86+OWZHKxCRDlbuF7gHBI4g11Qyrl
K7Ha6/tvTcPM2goUvLbvF9w3r4okW+i+9k/Xq2Gczz1ShgLJ5k3268HNs0WOZxWpsdqgqUGyS4kY
L2CXC1WDRXs6lQBteYcdTD7w8vq0ZHTeaSKP9E+FuRWZs2VtUTiQTbdqz83r6+ZntolfkyrbZ9nM
UkkjjspFpAtQlGCntjmqXwuZPnlW6Po475vIsWcsQeU7HKaHhuHwkIUWY0HR1fl+LqopeFqTg0BC
MrT3CuHs0TyrJ4YnOL9tmULg5J0bVbqU1zadRmNOxrp6kW9iLIRQbRRcbjC5O2A9AIjR14YVGm8+
OzMnvM8y+RMGHG7iyNiwphM0VfesoX5dHCHaTi2JnKcjwVRgEE6SPtnY7f4YwVBfCmsdTCjXclmn
abIjH96I2XlHG1BqbAFpYitU2lxcZLBZyAwgOUXfIAUPoBXC9twK6EGawUCgRAMKb+MdAiMWDFlV
yoKCXtd9hv4liTGedje6HGQ4kTZ9WGc6ueo6jbW6pN7qc0pynnKTjvC50+HW7g0wXWAxWQTKPQAA
dDO7cLeFjQPuuBs3FGFfExb1uBUZIIycdV61axYXseHoM/UbRjpxUppIU9S1U8GW0KrzJavgkiVV
2SMvGm+rL5VSBvUEypISbOCrTSo0FcRyqd+Olhs/NoKvrcKwcucuhjStlt9iVAHhrZ0FxXYK+DpC
m/+1wvJv/WdMnNSX8yRy3TyGX/AjOmDJIgmyNMboYdfYVU6jcmcsLcBQH03Q6CVvjN0KPGv+z0fP
WlhBNoY0SD+qeJdiV5cHlVSp7P+7n2+6EFqOx/2k7pBVlvvfACG4ozg3fMdL21Fs+XiePNuTGA90
gMpPhofgkLpIYHJY4qo5zum4rKaidbZZqJ8mhre1iRsKpSCtlWou+NjsO2bpZL3v7uP7Kh/1yLfI
A/Gb+jRTPwRO1oUk8rPHHn8awmh+TrazeA6gABw1kHNE1uvOgOtnwL2gmYWL6xTi9SHbiFohKEgS
uk+wp6sVF8qP2j6SVQbiOoVPgaVWXSfP50nJr8V1y/CTYrYoGBAlzyYZKTBxWxbpdu5z8F1miRyM
xB1Ml9BNzcDFOadBGabjbieoOMcL5q86JOcOZsh8FDp+IZnbPe9Hbg1MfC2lPlggSKcIlaftEBft
hxXDo6AsZZ1bFthnGVoo0JphYo7j2Lapsm0aXze2i8LZB16YSjdOP2IpxVC0v5jGaDA6K7G4gcTL
yFoC4erpm5gE1x0sv1VQgIuUZ8v0vpFvYSY9W0MPUz0SyTaGGlOI4JL3PNMrBKDvFrWJPqzM6t/R
FrDo6o9EzU57du73dx0RvcJegtZX3OPO3vq/Uk8iIJlSfLME3565cB80eV1J0FfPIxjpSr0dB6J0
3tTuZoITICSXjMUDthSyculJWQcps0gsYNNxm7qKykCYvvtoGGcPpO0mujooMtm8u5zubEcQjLws
B55XUBvmGroa6l0tciq/+ALWvbV1uHOC5E+nusSi+t5uN/WcmHc97V44pAqKhnPcGmE5Adh1DhMu
rJVWhPTQsPglmjYxSjwOj+nnyJtrjNLWI3JvPYsLES+EBDlMBbT0F9YPIUcx3FRoFfILMF59OzKf
wdPz1UcZx3o4WOf7Mz2rpydAZqY362tQ4v8UJdZvM+kW49KPZ//rNSY++1R8N/Zsk21eUePGMpOL
VZFl5Fpd11i8ZUOg1LWUl50klMZYs47vwb3D8Hr3I/A8T7fCZ/4dSexADLzZIn+NO7tFDJC4Z2zp
/4iYfOy78yZZMo4TCT+k9ax020SQRrC1B3VL+kYEf+AJyVbcxdIsHP/sjsIZyqCvsl7//Fy0SMGZ
AeMgbPN+s7S+qsvXMT96JFqh373aiTUlM6CjX6wtuJ5m3bkxKtsla/EsNKHH6Av+fMUR2bM+Yco6
Bk98Ud3+HGGCOxTQzwK41+lMdVJ5/PZ2ksDH0Xq08sk6fJUcsR63P+whUzDeQP4KX5w7zpUbulen
9zuGoye5jG8TSZLVrBD+4/n4dJNidbDA6UtxkN5T+3x54TiJ+lt8Usjh33KEdMQZr2WIxYo+5Msr
ADuHWJKlThUxCfl9IGLzNNR8bWvW5aTcfPHl20G77K/iqLF4Xz5IyeRyYfSzx4NeN3XS7mvBG6zV
Jka+u9B29/1OC1L+709y2gBF7HAkokCZQ343juwdLO9KztJ389lVadcVUNM0/SgcwbPkOzB8nl/c
pcn2JE+MXaszUa8DzuoIwokf1PvuCyqqPEUW3D0CP38B3oLd12BO8BJVXh75dHrv5gF6V37D7ApY
K6w8oRT43Jxdtavyv5PtpoDeHjJoJNoB9eAVdCWnLrrtRgT8BOVtO3JKKwgqbQQeBPJ6vbO9NlKo
bJVuvmiQoF/SnwIA29xFnl9AqDrBaYLa1DjoIMElEAiNUuCLAj1vqR0yZgqQd1ELVtRLbJCAirIf
IGVYNmysPfhTk6jDfIc1VBWLVtOapah17REVXa4tRa5FCi+gtaLe2KPwX220vIqdgbOV6kHvkXrP
mYbFZ+HpHv3Uswv/Q2U8VpH65jnKBTP6F/1rADeYiSWVBfYhlwWlQlzyiWawXXeRLD2+sGkqlFQg
P8jJT3rBAWGhvhRsb+ly1SiBUTKBWtnZEPtR420NB9542Ior1JZBEXxP74pUJ6NBgfByhZGFlj5z
n/VS5J5g2jFxTpXnqdqM+KxLnlXAVGVSvcfjJ6rR+y25OFD5XH6NNvVXKggowglH18wJhN3297Ca
c2BaBIQYNlqsbR8dvtz1klaPv1svOtmueMdPobQ6Q2HiymCBN9ECwCCsTwZFGdf5cVYQz0ZdH4rc
2aBtMd1n9lQFEBf8sypxIkQd01O0YOn0Td7NUn155jaR6tQBgNOXswf1iWy6nwn3wu6IOa/15GvG
IPUP9YD99pquWd6xFDKWRn7puNIwqz+sSiJBv/4JDT8eET2wBqgQMjKcMEdnBPpzU+fYjfuvYFnx
xP7scK19AQkJIQcsNm6CbLEbDSwweieMSFEsEzAWCuWcD6iq7TMn8dnL8zQ0YLDx0LwfDASFaC5O
yXTYp/powRsPOqC0FBXBTDkSSlOudKqyAPxo4RjQ3sRUKs30HnGCzfM6gCjZP0NFUEPOMHrvjTI1
mcCunwAPW18peXIaVwan6MfSyQbHPxBC8qaYBpykIUpN9VyGrYwbeU9oU7ojVX4lCLWpOyFm9ddg
oBTgc18RcxVoizPyItJW1CyjGfKEvIaHZEowMa0SWG+S2dpH5lqCTPQCcF6OW2g8UXdFZLkrXUrN
PSZ9p0NaXvrGdkdzjP1SLnC6CIFjLHmw5MoNY1wPDHz+wr2QMyTwEnnpfuxOYIGxJI58GrKk9rSR
8gzKwRTQqOeZmw2UvIs5L4MRC9or1UKYTGevPj/xyyJm2N08+Agk+M2xTXRTBvA30NXzowdR0KDq
hKduzswcc2G2hKLLhiC71eZ4aDTmn9arV6wfcvwCEfdf5WrAxXTq3Xyt0Ps7anpgVQq1ZkmlgOAG
ZRoaxfOepbR8aXvK8yGNF9j4yoRFQIhhr/6Lqg9Cw1mR8gd1p1umHPbbUSUvV3lDqM3xImAezoda
TVKRs7uPIGz/l93dvyueUQqRZwqyJCZjb9I3f3aIKvsiixcgcwFxJ3szeD3xwpzHqC/K+u2Po9zM
140QxdfmsddKyXpR7t6YOiPVAzEG9CfUCxBHBFTUWi9U+8ZQOppgBbi8kdYMuWLjz/qhdQIw01Ho
8gqTlitt71czFpA/0WykCesjAJEi/tpWsJv4ja5PmAmpr4Sm2SM3r4gBIg6aiEuAxx/xjzSRtPdO
iX4eWarDs7gQW/bGdloRXrSCyyGHRSqj9xO+Hlinh4M/nKXaBQnANYvkjx4A12CrCL5DG9szV3Ed
93ujMlnmPrLqVluqhgNkpFjbbcSLVRZyQbFjH9gPZCEYR1SPxsCCZ16TafMyelX0Q5lxXajUQIoc
Co5PskOzsuPISnIx6gRlBQU4Ut+U6Rskkl7Who9wvgwyjfputCYlxF70TC/hD6rH4X9YyYIptdOR
3UepO77cqOzZ9tIHmZ3FQ4JPYhu6pzgeAIsRaxlqOUrvnNjdOpguCaCj5s/Q6IQyaU78ZDn7n7q7
oME4Vch6iLMaLQlpoKTuHEQ0eXFf3LL2cU5Vl+SX3VhtJeLk4AlqMTVqYBbl88cCzbGQYbUTr6i9
Q0Ka1b/7nyO9/By/gSlnQxTqJ6Id36Ou6YFp1PWQhp98JPetvE6Mcbepr5Rr6WKuaMa8CMKAlxWG
U0HbZSiUuUYCatVZ9bJjacv6IREunWZi38q4wiOLnVJT8agpfysrb1aiANjdeWkhhY2d2jUoo5jc
NOvXp1I3POiIY3HgNtcTLVvtQwJlsVSED6gFrn/mysKdE42CpI7XMMMNaRcLEpBcIcdih0sCk8Jp
ZcesJf3xlio8vMhtiiss3XJAmkqs3TmY4V/pdYQuXl/7pRSPQH4wgqCovqSABC8jZHMoSl6xwA1v
xcxiMXAeSgo/z8JRznpvE1pBTJL5NgCuUFU/yoVhGNhEKpaXUJMoKgGCGivS9aBxXQf7CnBb7Zcn
Nkk1Y6OU207KbRaBhb2m5Ij5f6MNqTttirHdwY6JOpgM/6Q3HjFENX7OUv2i5FvHLfGxzviweVRK
sQTtQ5TJ4K1CnNWircXdWMs/jqtdFmPlpcBaF2Vmc7jkF3apqSC3ET+o6prpl4bXBQVVlVzwTsTa
UCuyAy90EZA5vvSZgb4r39yyPQlwst0AEbYGyiw5GGYbZb+DZ8/rStguE3EK2PTHtIgZp5Z8BnKo
trBC2YhJotq2c0JBKfMzCNCYLhjnFbU1KBuCAxdw8ynsJa1WQGMjPc+OY4bwEGWZw1Xf4GGibftp
J6tXG/UMr4QLzqXhr+tHSinjsXV1bLcmhZWbDPvLtKsh5qFAYd9FFEBs3nszNPhEws9VQz7kaV/B
SzvtrK4vzDrbM3IVEX36Sm4S0t+ECZ6/A/O0gZXVoGLlHUwp3AENJfo/T5UlLTaaArlG7nm0vDyL
VnTtutBCAceclo8+3hn5hPjGcDvvVOy9rGpDgKL2j4VgNZHbZfprKJdWHRbXXzkyjzj4u5bHXPNi
INZpxa4l0U0bxydiSfgAJReZqm/2bJUQE5fBUxglR2r2G2rEXosSxympBEx/iyYZxbGBrCcZBT9Y
OXIp6NpokKu4WTAzmtXyVifuCMWyX6RgOryW1EmkTj1Rj17j8heH6oQrIAZD8X7EMhwrzp5LBQr8
rCsaxdZZ02gTXhS2mAD1jj2LVF2Z/cXk+iTO3tRf+/uG8PIWJZIKGwHrmh83mYjdUWpicWxbYLBw
P3UP5AN8UyKb6qaZlM4X5uaT7iHrMWvaBsqX6fEzUZaCL5Ygb0WkpAw4So1kvBCpv4k4a5UzTRqU
SSZqkFNS2VcpbmauZb7JvZRw9mWH5DqdWtf3+T2a1mIovn501urWdjrxQ+8noSMwpoY4vPpZz8Qf
BDOuJsyjBPZCZ3Yjlch9gMidno0whtVooQ4I7lBOEO7J8iAAsmYgJ7//EutgLGoGxJF8AnCduO5p
SVMk6JKsy6Yniml5xgfUJ01NtwH60psEwdUoexWFSQcS7NgkMdXm9qWuU3wjUkz1XISojgojXv7Y
8adsgXmxAiPZqQOT/vJOgIP5J3WRSb31/TsVnpf+KoHWkoLIUUOOPJ0K9eNdIDd3Yf/bQ6zBP39P
cHaKXsNH9QV4sCl3R4zlAfgu38VsZJhOA8G3o2AX+gwQxAFkwmEpuxrUqxiugWmtBEaEKPaPlD2e
D61Uvl4v2wD3hzcq9GdlGXytF2oAHhVX2pozdq5ZRykpIUtNhYOUfhDcEE5FP8wwyLfD5PAInk+U
9QpgE6r90IT4PhifnOppEGnLsYqicnpaHU8Abh4Z1uFqm3y/ect1E37+/xtGkOaEnijFz/L71xzp
UihRmbgd25Kq5UuyWDJwJNY/yN/rUSVcFuvCo73AMjrx3rTHWoJs5UC7b9MRml8JoTgOvi6/Fio8
GkdQB25hjZqMn7A7G01isY4lpd+DykeWsl7ePq1OtuYyR7zjiTWi5Gn7XvV0fwbcSVVUtj8VUObp
w73ie2DxFVifDo0EHQCGlIPIHm85G/szWzA6LNcMESXmiqoQKUXwZokKXYWu0lMPzAopGBdarK9G
SIVMB6wJ4lgSzduAeNwozwdG5loUi2jEho09ddE+KnIllivsfdgNWSsSqo1FXyk9SRQXC2l8BzS8
Ml+Ax/8Rh8e8vJ3vYrdveC18/tHvGj/mdqnuCXZKciofNgd5hUUj+E5TInIRM7xnv4SVf/b6I/KV
z/4Dk8et+l6oj1uD+5a8hmKmwG7lAOweL8n1wz9S6xyp7mSv+uHQ7KPGth4ACxcbmTzJzgjYaEJM
6GIFWanxWO8IF49ZmSX2Ng9qHGGH++2zOhAUhAYi7stn8FuIbEaaRYzA9nvF/sewui0/opYoFL+2
zNg+gV+Ws0S1LubjeiSvfgj6TRW8qumXRUEWjBqwfPxLYvAzHYGyjPtgH0Ikv3KOPd3ioP1zFzk1
veRBOfdtm/iNrL2iEiXxkKCAoocp6HreX2s4Rmsv3xOgxaAxEI5ANqIsWzzjI6rgyeI+5fxcMGfS
z8Dvv32FpvqU9mix1zshDb/9RFUHvr1Z4q7vXkXNsYDfvl07UH8ExP9lMqkFGyf9kmqtbgfsuMf7
dP2pCn3Wtj/jMLey7PH+X7hMAsXAy6Fy+5dJEH7nowZmLowsDbKbUVnvHnlGGTRI7mmqGM4l7Llm
MZMmrOdZOxxCrE3iGQw9pFArz0cnGcf7bWal7JflZmbyVsyyNaYhNPyQdZ0oDpk31+l4pX7+nswG
8t741li9j5xFWg5HZXZ0YkrXA5H5AiL525YbdPJFoCSptpywN7TQyydt2sBbSccRsNklw920esRR
X9NIryaKFQ8b8ASfvNiNNwkd7kotLXxZm4tCeLg0+1t8g/pO1fKOo0ttHw37lMp8PxnJvL/641pP
KQ4tm0G6KhAE4V7WlpsWTdAl3IOnAqoiUrfGGfpidfspG/GogY/wD2Dgp9L4xPNgCvIlYSMqapYQ
byUJpoXpu/0XJ8yAjBkBAq5vzT9c0NVVrV8efYGfD0JS7R/T+LOAnTt9PIkfCO/X/wcFFXgrLYlo
vXqz4pMtRvlQ6WcjYRN2cnh563Es7q7ba21p/XkojDzqeu7C5e69pII8MruOwDFoOW2mhhqu9+tc
UziZ0Y8lsQFYX/+frAdjBvinX6ChVAbJLpa5SxxF1aVekq+ltBjRms3coi81w5T6QTMi+PlyuCWE
aQ3p8NvIDCAY4bvno6Z7w4w7naAYRhzuC+af0Agz6NOzIcNsxy+7pyadmjfbyGRHJb1knrVZmDe0
jwUhoTpYzL+jgAGblL8Tu/e0Me0O6Kb+KBVqPsfUAe1MgWGqaLdtq6Md97nvQA73/gMtXBZzwz5F
3kGAwW3W8FAou4rDToRbN2eASJQY+yglggkMSEHjwRp+HF0A3kc3BcJNEWx+MaTfn6eGfrBcVBbU
Dl+W0tCHXJICDAY3PwP7cQ6hh+9/XuFPQmwkpiU9fiVskIFS6lZlAcsau5qlWV3C99ISG9uHMH9S
iTGThcFPi1Qww0dYvKp7qYAtivhXsVzCh6e4su736UmXG1WMd9Z7ZqXkW/owmUUyvpLxseluDgDh
jbvIVgpwjMCjEUcCiH6brJRHUE5cJ8SQM+QYL+h/ZyXuLnhcW1OHhmDrQWFwU1GLnK2qkNo05slK
I6JiU58dScOWZ7/TJBcsTh8MCpY+Wmcyrwad0Pk4Vr+LTV2+5lNBIzmaYIbkP+QTaGKIgB//6kqS
Hx/l8bsPXiuLNiQ3FoXfqqGhd+Bt4BFwbtOdFJld3NiJt3My/nFhjQPHi8fw53TbSDaYXhaO2yc7
Gn8tskuQ/98WQWdKEL1QK3kV+FxlnVau8TYB7SHcQvi1GWaVJSP6LKMJB9/7baY86z57wmtamrwr
ufhDI21t8TWfzRTLncVgYoTrrn8lL55PC+9X0YS5VftFbhrW4UCXwrqh01SYLEn/fJtMfOzMKdVv
7GlcO0FmQvbDs1MG5pc5UT0UXOH+VAyZJDdY/LUnDQsZxFqd2I+Q8JRtQ3oeX3L8R0Ayw8plYd8K
+E/MtwAjB20YizL6p2Z7pf3ueY/o+ZIWPX8DdZOWgYWAkMN1JzzH17ftStNnEtZEEvP7CTDSwXr/
jiIVniVhbdTDpSIBau55JDxZVWUGyJoJsVAgKqTPhfrmXiWHMiYI9kuhwI9s66+uOJka+e9ZlF0J
xUYGnr62O7bwPV6thslLQEeYluSaCmsdYqeoHRskQgm45wRfsmBWy72SVv20v1a5X5SQb8lGHIJ5
cYf/iw2GI0JbXGxPPC68jjdsi0jSth9Zq7XxRE2AUS3GHIpUGGLJb9WOjLJ+j965Vtsu+SgrHgdP
dPjgm3xK9HULlchsq9xcqSf4Q5RXiuaS9AoilEhfqm9QIxaktdyaiMUl8Q4jEXX1VwGiIPYH0Syb
VVWI7+6PwZkcS9Rt4K0ApH7ebaQUIMwQ+SlXbSwyzeLhkSGy1qSSslqakRSa8igcfD7NHw/oXRuJ
56jP4k+eSrVU6iWWq+ySNCobEcNxCvnMJHzSvNq2I/5Pp3iHiWvKWsKKKdf46z0XXvvAN85gpnUn
z05rkWEA/Yy95OmlmTNzBgSS0J/fK8q28ltv5AzJnkA7S5RCenV9tszssHhykfa1lD/wM4KdqxIN
cyh4kbiS4nI3s93lWXnt8m/PQNm4Xmrf/vjJeZhsP8BuqcajzHXBV1npkHg/TGz93CyZORGbht1R
oan9mFywokrqNKytFbAO8UNGV90FXDv3iqJ4bXE3vDl787TXkrzhtt+icCMhFzkQYGeKk++mw3G2
8fh8rP/gBYiy6t60fMk8IqOOudme7b8dIsr7zhG0LyPjjzP2MdTJWrpW/iIlocXhi7n9ZzsSDi9o
mJSatjhAF8NXSqTB8v+h2A484uoqJvz5fgzeE2mhbziR59hAyRMprN3cB4qhT7uZo7SLbbWXuJra
WDJd4ivsIM2CUDaLCtrWMf5UczT0bozpweTSoFNGRKOmjr5muV2vIfM3deujFZNwy+3wtIpbv4a8
5glU2O22vV0ycF5Ast8rXebnmaPBLaI/c4NgiiULgE2KTUedH8ilqbvwnTezMimpUCOsv9lkISf4
X+ewfd3tBsXPuZ3kqskE/86NuW3Dxjsi08gcXAu+I1PrtIGKZxdb18utnIXfNSHeAvyN3nVwKdnt
ADUUrHoL+UiMKIUBwe7Ro52Uxq1he95WFdEbbDP0fg5nCuqHojmRg2bQmPHLxDdh+TcRktthqvc4
K+9Z+Airv93+V9z+DBpKvPWmAhDqFcGnlw5L/+uk1q81H1vS+ZK45Szr3PLwA3oNbLKCIjt2MmJt
eVwkI8H8rrKPpJJsaJuEUgG+tTCuf0FSkqyocQ4oQo9++qRmGVT0zty19yn16mCd96Q5FAiOeXoN
f8Pg2aKC/POwcwh4E2wfe8Rn8WGQy1NTht0LKvSEWMAqNwuGRsU38TzFvBzebkcsFfa67x9/IERR
fu8GSzVyaUOPf+YXH34ToujLjslEKWC/Z5xFFtuRzKU8FOvhggi5o3NY22Nkew5QEMCAhwLyaEGn
hF3PtmxUGKmXuAW41oRGZVGSn28lAMGwJ3aY+vkpoLI3rkcGQOZ19zjiFcNhkeET6IHUjHzslJ7L
X9blztKshtbStz2E3sNObSa/1ISRQ6xgKVBfVhH8baNIe92mIYyagtcX+GJhuqcjZwpAz0Q+XYPN
ZAGOHYWj6NiHnyT2pEBq2wz/IOO6mkWeC3aFdSQezhlZwh3BEb1/aaKwyGUXP5Hdqd7gRZUws4wo
i/p2DAi+J9WBKi718XnEqvdIExPmQNk47CNEjybhb/zmVWkD3gg0Ufhph6UD4fQzxwSV2QxR4ZgK
cnwgrnBluy4mbuJ58pnEMJT0zr7/LBo/SFPNMJWn956D6nhzeuvb4XZNk4eFB6FpktRdS5Ej/ETM
qJ8KsS/ZYFC84uRFa0l87/UULout1GR9Co2xSfSwQDGenIGKsuhmIUyVQfSUSOa6Z8hWvs5IqM3w
I+teVB74JoYAp9aBzJj7wqzdJgeGxPQlticlENTOgA7eYJ8zEfFjzzTBqSNAFmzfLdMbdtT1uMlH
g0S+5uRRbOMI5bEUp0xE4TCdvLsmL9ruuF75pBs7gfdO7PWF+42mrX1wRy7f4meAX2//fB0kc5ef
MJFvqbLHCbaZRZhB0VEMKDnjJLhnn9JNCY/00EIGbhFX4cNisVGs2NcXKsSxv0AQ/iXjfrCvLVjX
VfpEO4Hir7SlnX+OmkfzHrzobYGKN9FE6pYFQjSoyzGnDdpEx+k4pQpb75rnoLDGWfG+A18KScLr
amXDKvGSmIUucEJkZhxy2Y9HTVkSGQF7zNBamRAh/7Cj+a3PfgWvJ+vHqyHVWke3FFEyL2ZctK+k
vErCuILmkSf/Xirjp0Iw1WxguT7w6XioMFjIZ8cLpplxATp/mwBqnSHibGhBCpGHe9lBss7cDxun
wHqesL0Lvp1HxX7LXiOgZORlM6BPKSRB1zcI3jpKb6HtUgDaKVC1LV4g0Be2owZ0Q3rbsEa1BRGH
jFqkQVZKWMMJnnjsbf9SW8AeDwEJqd1eJHuohxvXp2E3CWasWvvmTM3Tu1w8UDeccgkk4QF+g2Uz
u5/dqt4vJLyhCoFQSPC9C6lAS1aeJLANkaqvqyRiSyJ3JCbrqCBrt3mij8YPc679OfV89005H2LG
FxjL9cS2a8NfRVBVkJZURo7sanput6t5p7GRx29MPT2zbW8JKDzHnX6Kp0fTrUe7gvKkmtFMjutL
4Uz4T/+o/erkX6bd1OnsxbAJTMYLSTHFrhjlmEa1dWsCbM0jjl6ZoQQFVEdJAGyERACw+kokxVu9
kBDzOFuPzSSQR4bT1FUfWp7xkdNCkExGP4gcN/kXLEGusYEo9QAUSP/tznBwl4gt4AKKZYHbKH0L
cR6L2GR1NEjWCEVZ6BFntwkwboVV+eqI5e28b8JIJr1lA7ZY6zv9HC+QXu31QdK8MumEA/+Fzjnp
BQ7j9ag+Vq2hOuZKhOXgQjlNJs9KHQzPJDtW4nhZIBw2+Y/H4yPmJ8zxkXGWJ1kcLL2WPlXLkrga
GLOVhhQamaxy1T3OxAo/X8hJUcifhm1t0yyCYaPw3/5EY0/qI24OzA2Ox6uWG1t0s0CR+wjDMwHU
TcTNRORKleXYxtFZALSFowlXdCUrjnuENLw9VIC4kCAR4Lv8NPdj58hk5wyti0LisU6qXyIrp3F7
LqMJ5jEbL9L8SqMs+SwmrX90El6ui/d+3fjLMCq6gUae5hA+N8LumpqQE8xIw3Jsq0RWiLSch7tC
4hqLL4G6+WSzKQueabK+Ff13V/s5dDF4YQDD49K9InxPW+dk74sstNEwB5pnyWJk6cWcmqOz+Jdy
MXQC1JwpAe6GbB4yF2C907tqbQRLz9q2bOLmmor7y5ue0l2ugeHjU3ZIZDzmCHZoDbsPCe+IvoWP
7vZrM6f42Eiy715shzbnkX6cT8+CUvdmTOuH1hAauFwz6vemLBB4/pQISJZqFjPyrFE7qTvIyFVo
K5VwV0wVf842aMQcrWEyVWJ9Sdjr3kXY5wGK5lJe6Y2yBgGfqTlWkRkOi/n7TfWxP61gvn3sj3dX
D2kPmKXLtY3RzGZrt7XgmHMzsUqq+FLIFUIfgd+PIuNdjlCRX5OMyslLwN2+Sy4ZSj4E74IrVbyj
88MVKDkyFpw7FGrzaJVYM6Kr8Qa7rZwoHqt9P2FVHuk+ayRnBwaYKdVBKhyAAiodqxgAqQMXg2aX
yRcbKBGZxtZ01rvO0JZ7f4IVKSrmT5+a+6XyIko8uYS11QhOf+MZI76IZO2b4owRrOTouf9tQ8ed
N5FCkyKcZfcfgm1OdD8VGhroKUOlYV8O2A3aUH0OodGPY1D6Mev1JZRGk8eQOyAspZDA0l6xbMkq
0dW4bgA8CxX0S0CpoDex1aCzjSRsNt2UktEQ0khew8im47K3KNJH2E5SFQwnyOBORVPUJzMyVvRP
01qAJRPMt5zq7tp3/ldCe5kOkO6+8yE6HkXfvaUuwo7qiAtYFgxf8CVbN9uOTY7BXJatve7rXJYf
2Ujx1P29pz864AFwhtLIcny2Y0cazLccs8S3vbL6EGNxRvmXoheyJuiHt5JPt0/N4APMKHtPOIsX
ERbBHmhLQhx052SEqbu4dLhqaYKm7V5skon2PSH7KdDAq+P+YZcw7fbrTkiyEAEC2LrI9N41Yo4A
gKdOQ+CzmQVm5bZiV6vRmNdbylE+HUQYO6FtvlsGVqfZV8nh+0FG8aV+q8aOJdQLe99QzswVdMpW
6Sf7vMjmp5y+Ao/r12Rs78qwB3gvU416wgJ8OgrcEOtxIwbxG3xcXAoA6Iv7EIFAnF86u22URfKl
Vxs7U7O8cDJY+U4FO6vu/tbJv1Gu+lPRuwuaNV0rwp6tXI9kkthIyf/rqKO0hNVV+0X1dnIvC+I7
iADjW/qXdnNydgsSM4YRHI1X/S7b7pYi9groh0vU++XSe0CcTxXHNGh+tmlnRGB3veipRE/TEGnj
1zDV/xt/UnFG5eO4pY1JF41XvJcJfvR9skDp2cSuldvviDKNHXDkuHXxgdGzJ5i8vALuQ72/8GSs
llFH4HGEh3d5tnam68EOpMRI1YFixjhfl7g/GHgJqvLr34YR/bVN8BNOvjEq4YVDYv6sonlWBhgQ
fu2c/k/FSGOnM4va1YmVxM+T28HYfpx8x0os6ViXF2vv/2k/oRdGmvhIl4hKoJj2QcROrBWipgXw
ZtLtfHdgUNdVK232l/1FZUYZgDVT7lGntoWWjlybn5bU8aWVHF9Gt2GB/8nwNpfTWdI543V3EeDM
UqbIHgOxa5cmJHHfwDzxC9b1RaabSYHPtJc7l35pC1FlwG3shcmDPD578V5afiI9YBOIF1WYuTN0
cTqpGrXckppcZ+I2fd8wyar5hTe3+LqH/n3dzVKLAgzK5F2naV082cCgCFcIKiB/jcAOoxGZparZ
JFJk4/tIvpIcqQ3INd7rCN/7VYliE7ZM37BlN5ZbMF4FNnjbw0bLlWoOfJ14VsOvQzsSLgfwIqZn
0XMNe+tFCijAwnKfvqlLflCIAUWAkgBNB65kp86apQa4VZtqC2RTGpFU/eZolGbiIdO36w/hffc5
j36Ye2i3XZeF05G7Ocy+qtwVUltgGbIyCXLrMUw3bWpBBwO/W43PNqqgRyM5EOxJnhHECK6IfVkE
OX9vbM6wwNHSdgLVLwb88+xFJOoVxNvpNcq+B/j45psjqM6Cs1qUOUJCPvBYuZrl9sqQC9uLv18A
E8o6YdFo2ZNbYNSwzXBXS5cElWZ/edGQURm/aXRqlmlCNXwGUrJoivRBg9cYMnomsBIxAtFl1cCf
jArOcDa11jmniDP99ZLjUXEb5T6ab7R2KK0HgfX5VtT/kRjfFXvcJR26fBNUfOoMh1I2GV1CCI5M
87vrTfLXS5uvesdmWlv7976dGemA81jqtlyy1vB8ld4X5sxjdJTOU/yxyIvtig9b+gRZTpxE2wT2
usakYfkWDs4XLWal37cZBsqXmIHkddN7K+Ihiy6SeQzEORohlUEFxLJrpGCB66Ep1OdRbyb4l5ob
EFBLz7dLxDWH9beS4hAX+pIwSFHaU3Nqok7Q9/ZpJsQzD88usW4x6Cf/7vLSxP+eEeY4lk3x+G9T
Dup+V5y4k4BNBDqA0wcegJlNzMfNBoPvO2vEisd1u/MwPTlAKyDFZwQrcXKMoclYzKIk48ILSQcX
pos1EVe23dmajJDT86tQWEaFvAecmwbdMk8SvL/1tD2FdDowSLuDnZ70KJshOMNGkEDO9R9DBmOF
Mh1bDkuXV9xPWiSi47lff1p4d45tbw38dGtDVD09Yvf01CINctl1Wbo8A0YtfWKtItNMidqDxXID
8S/h5jkzdlimzdPl+2U9rE7YcdQt7bLKD3XYW90P6RbLzTIdSIrvjwGYDlWHsX/WUhIXhGrwpoXI
Xa5p6Z1WYo7ln9EYLIYRyJo0gNntsxsgrlTurtM1z3sbnNHbwGZeqW1LTAtKCPhdNQhcYb9JJcVf
Iic+GVxKLXsl5Zgr7B+JEF0SFLIbHgeizHJbSqBei+4zkojBWsiFgEGn8Y9cLw7UYr/UKrUIEF7H
qopDCarsAZd/zS4cp6NY0mj4Vu1xCiVv8Ox8ZDc559DwoHvC2DfUcAQJx1Z5Wlg3jZDANZurFEH5
fk/jPHbSC09r/KxWhAz3JFlUR0cXEm6P0g0KtkRjS8OCyuDKWayIrSAWsi+OxegROn/Whmtp/Njd
//lQ5mkr0uBXZjsvRiN40NAKo3DomS/zbPqI5q1Q9rNFV9NqR3mhdaEJZMR18uxpK5SiTsm8Gavj
3ZnKFkBBHIXVoYeAQj64lgI6fk6RaY3AvnJDPz5RCEjpABTC25hBarh42DnrcATcJnPSSJhJG30+
8MXqwW8/78TNlaN4d+97jsA3+ClbRWKeNpaC4juvWJV1tkn+QoIiXxJDv4CjPoOe7UxRb1P9ifaX
d5E6ODaEc5Tysvh1PR7ixosZRhbKmip5dnHbqV620zn9CEoGgQFrT5bXJA8se7mtNFVr5ElezehX
DRozycZaiFBmEv0i2+zwXxAalnNrlK//Lrtk889g2s8wcGNOgZlGSxflY8zLNA6pi6s24ustWLGb
o2cC7pydNxBqNmnKsWqAmWRMVovI7og0DV3DyGJshkE1+7jkT4dIjFSTSgTqkDHhFT1xcmlKaMcs
bFKXQoYKZvd8KWqBMsaZ6WG+zRS8H/wFoVMYgXU5H+FscI1FNkyqDHN0Ii/e0+5mwWYDoHH9xCTj
3KyFhlS31NvH9pIKPd74A1ga+6LEaDeVDAzxeE0/iowSgd7moNlZqIYMxudRdN6dt0kXL9DNC49V
reJKePGu4R0VlHQu5Gqyc9v3x6MS9aMs3bs2IrDIMa13zoY4Nzq+bR0dN+X9g2VVSdFFBnw+CMSz
1Z6gRZmEuCYAVrqfpYrIoM9mSvD2cB/hYrtSG5kJA3dwlghfZ3EogejlkwZPreBcIzvIE3XZmPBn
WInuzaHnjlGfCgBifJ39LDqhsAE4LtmPOZ0qrx1KBevCULrXO5DVQyGSxqfBdW+vVFG9nY9uwTXU
zSi94rMVaVT9MpCQexQpdiqy5/SerSm9rTtsoDfe7NNFNFcNF7Zfo8JjI0aI9VjQYWWRJ7yw1RcJ
nw4/q56io0uJzN6M2Us6jYKPWifaiG3Toh+ZnsY9ZJKdQnvrp2WvZcJEkj8VzaHHRPRK7szY0P+x
2gB/xj17lomAehtH3Axm2rW+xdZaKukuaEq+IyDoKaB2y3sVOIFXnff4M9W6ZIu6uF8vaYfFp8vr
Jp9qAu3GhpC6yY09lNtlAYw0Yjx+zvS43h8R8CT8D4AnmM3qoV96kOLcbT5IFyGYkj4OFp3VcieO
RV1Ir5LC6giAHjmMgjtfMNQgWu3MOVlouDvcntvk5VZ3gJTd1S7IcVm6XGJrjpanqVg4v4GYgHFn
gb2iLvyzn1Fb42R3kv8jwmiqnOX8oZZRp9CeV/ECe5sqMq2/qvrCuFciU6lxkOAjQ/yxxBUsuE4a
feHI5MDcuyzhwyoSfmIq6WU0r38NrB8Z1Dbt2K1A9VFx4PR+MWOw0gY/AwOw5I1kSeQ4PMDMjTDY
2wmFnfLL9//WKhn7J4Sje71EjpT7+nGPOKDkVqJRDz0buceVJrK732u0R3PHDryCpNJRGzPAMEhc
xFCilT2Zhl56HKmgQ7VZvOqxo7Uaoo8dqEmfMkSF/AHDrdEZSEDRE6+X35JBQlVyQHEyl8TNJ5R4
RtnyTpnukBwjZhGBs8iKsGsSrN/jmcKXwF7XECh8zgfJxseHYUSJPdZ0wm9AVVnrnWAQXT3x2zy7
vfyV1WqBGQX72OkPOGC/X0rQHt3qm4pCYbIod9UhqYtZiBFPMxOjEnK1MZ+roLirXO9bWkecZ4e7
mN1iQf879TJb0RROUJpE49tChZEJO2PXXiswy5i2DbJmt5THG6PROW01DITk52jmWYJPAcu8Ev8Z
u/5OuQjNUmA3Y1C/N9LVRHZDdn8kXd+3Ssb+/QhpNS50/wq936kHbRRpJIZcnaCQ1Rs8YjHKLckc
KDGqQCwiEJWDhXTw0FzqqACPPuEnmoUIyVa7VQ5tcZLyNUvm/Lc2wIBd4gTbzrJA/n1zs2+8fbsP
AkmIvThH5zw9trbzvSlNAImvJOS7fQnTm1hequ/IOqQMvCJmMN6aupaNj6ULRV6vno7UQRd3Ndhe
aFGRoIk2qAZngND98ctoqVVySYH/aq+XkjorUddpcLQLeKrVx8PUyQxwWrEK1akZsbBXBudfNlfM
faymUu8+IR9+GB6OnOGvOOLTVPBBtAQiDCuT0gHCCoY7Y8C7kFIeGwIhCPsOmXaqQxlJKFEhZiih
CH/S37XN3lZ8qEKCT96RBZh24I5oAbAZOJmcmNDTY9UUCaVN8pumbssfRvRo5chyPeKfxMoHY6KS
l30MBc702ZhcFaSsFhKIt2XbpzBSmztQOuO6CetLXx3eJYCVoORmgJpj2XJ3K1W/7uU5KHUQI3Gc
3AXPFvVp52QL4vKyVJx36fef1u9X8RFYIOnA/YNvHuOWNX0U4uKDHS5gENC2Sl7ziEG8MEttaz7i
v0E7sGhfax3p9b+roypss3KQ1VgZJ4h1zsQPSi0gck+tN1tKVSWBONQqzit43VfSPCsJm4pn9av3
aAviobrPqK2WaGqMtfxsjImp5dsFfl+BHLsl01gptEcGc0s3nSWk6NTGA9vOAJrvFJrh3j0/u0/r
qSJ24e3aitH4970uNDDUCfVZyG7AO3/1pVNUKW13yZqREBPZDJ4S4iWmdG0jko/5eEGkHTDahIlL
HhnCMyaard8sWxX2t6k0AsP6axqVhDvw9ENTEf0DhAnFD4S+UM+ZSaVkxZYl2VBYErN4Lnez01F7
Sr/PafegsziBWS7cBF9m8RRUqJRrv3yGBskZ5zEnuePTlhcusgtJnj64LM2mb94+TNeqJbRWMOFi
k+7GGz4hoVYsYhaNKdkR6WFVz0InpoXoUO935BmIwZCv6oQ70ZpmDgcy2hqTkn2v4/CL0H4krBQ1
PFmgosSB40/hWiuoQakMGr3FNv5OIG6VdKNPqoSq8tOYN323/GKsrNEWtTPxUAPG4dFWm/AQ83QD
moVByCvoy2Ce1+q33R+IeoC1/cvKx4sjGGQLTiitIiG5Wz7ZNZXg2c05VeOhhQbnSLuEnlYibwHK
NN64xI2v+59PhlgvxhX1V6YnkFaDMm1bBjNWl8m241KvBr8J9/VcDVPiKeeTUZslUED0aZjqD4a1
niZt1sv59FJ1Vsie8Wixb6KMjYvNt4siN6O++jAs+JbGhaaZnbn7A53nHvCAogysXlDOORXCODJE
EYh8fEyODCwyKG9qOlAZPh4K9N01OStN+JwGltUXo3SvA7S7dAdAOjrBb4rxz6q1bO0V17KQ5X09
9xy0h0PVKDVCSheszdQDbQkL/Xaja5beaPuTG8m/dpUkQXCnhNAz6qqUFLwj0/cUYzh1Iq8dNw30
p9C31Xu0QI3sG2n2EIIuEXuc4vsmKiNKQz05ZvNNcXsf5r2gn2bsi+iEy7xFjwnY6o7v/1dxEJac
SmfRniDPysnGC1MD6T8y9lbAXGE90WPsed0oloFUySUklq1FlCVSkSrdqFbgU/BpsM9a66wLpNcs
56SThApJt7K+BcEON6Sty6rRugQhdw3cuTUH5gfiHX5eutk5eGLKjgs6cDzwQx3o+0ZYHhHqFtmu
PEHEVda1x+fa9JgxlxMf/5pf5K4UZsN+BhJ5o9ikzFJVZgB9LESwQL14ADD1tWfvwWaekzlbCq6p
O7fB4jCnqYhnQrmS1OI1EdUCl86YAhJ+NkhdAEk25QErxpqwYH2hkm6w0TwLP6X7edssAFg7Qxmj
2Uh6b4n50aWD7ZlzJAm5vKZ63zei7riI9Bw9sDDS9HmYDnGsgy8Ehow3Eivz7ad0EBX7dqGfKD87
m3vjI2cmSZUnVNmNdqCgB+t8bpHd7Hkk5kQFb3o5xZVyP7rNbkGHO9N67gnS9OS1H4p1T5kHNP4z
4a6wcKkCLXfj93TIpAnL3OSTNIEgZr1l6ukI4r4Sm5x38NlQ2jFBOxRdCF9DRHaD0FKs9ThngBfE
kq4yUVL1xsa6sgHHAqTK9329RZKGS27pGfItZQ/zabVNiueU2pG6BQ/smv+dRuMVwarn4pszK0yb
VIKAxosdkhFzeMpr8QReskgp3rhOFyFvsCxIIXNcIkbQnuekphGLLkqvd9dlUvWN5/gCk/6VHbII
KM0/dl0Bdej6Ogz1KZDhOA1PEuzey3eg5Eogw5IfuBNZUpxJqLw6g13luTLOCpu6H3ROn5h/CcwS
3+y6UQksJ4DLBEuXP2s9+9JRTL1i69iagym6ej8I4lZtDaV7ld160f3yShyx4z8z5EWwqyaCtLPS
Tw0qaF6609IYZJTaZGZh3+QGWRRVQuMI//gtWBzjA1Sa9/QwjZc4y0ywvQWopwEoHW/V0hm66cew
P9tor35MOTraofojy96jbigwVDd797OQvDoXIp49LKLchwQu+BzeZ+RV5rTVd8xJtiqMNWcpsI0K
2Edc0bVUgRKxEDgm2WNa2FOl/jC7QuL3pFDDFvkd4uSifSbfNE0HASWMv86k9hyxCSsAC/rcUh6q
wguOtaB7PfsrHe9SptTK4lXUR7f+rm4JiCJ8bv8zDqWx6ZlXFwJGtVahsImvIb3PDTT//r0fHGfg
kYkutVSF66mkihni2OOMbjcSgeCBmOanl/onA3Ufzlz4xfF3JZB/0PsQFh1OuTJd7R7pJBq7mWk/
q5TDc0dTBoRebGuK/D6bakiTkDPZx0loD5K0MTcCwFQlR40fE/CkxI+fUZlkhakwIafBBT0374aY
ofU/FJGC0b5C/TEJ95RLkLHv+Hcd7zGZ1SU3x17T/YaATKE3aKyKU+996WnBrmndatQs3fRXGb6e
nOi27nAkzUUIYDn/PB5MrBeb4RzgAgjbLyJ7qr1JrCuO5KnFm0u3C4hf9KbIYJ7tKXD2/WZsR3+f
6BLROPW1ofotTlMBjXd/9mkR7nCgNFpXy52rWX7irIp/CVyBckYERRL4+O/5QPIU9rD3tGevRErq
yxtkkAE04I2/YctXTsTFueLL8EE+ZLlwAmzXXOzrQLmTZ+CTXyMT3f3i/SASySvwq+YXvMMYz2qa
SgQvN8Uu1jrx/dwpHMgNNnGTQz98zU4zz1GoZ1jShCmqpv6Jj7H2rMHef1Y0a5M/sZVszVyemyWj
nw6A9UWFXIVdPEnFqBgFS7NPJNHtsyVcP07Newpnwg0gVdiRu2JjGSPUyuJWUzl2aV+QdL5EPrNm
EbFxAHNLCh/hyVrNoxVMhpe1kj476GeISLgIwc/kemcnxwltr5xZ7EFIxy2YGTf0m7XW2VwmDnqD
VjQNFWPPq8XqX7oJMSvrSYVVZCqz0dvN+RyYr9EYowAOw1hWEOC4G/BXIq2jgyAhr9fnm84x8BBz
YVtcrydlGAqvpAL2xneyQZE/tE98dnfRpSEZC0UCrgiPEqYgwWpDptko+azXVKII4wCNKScMxv4Y
hOuylf7FOV5P0Xanmk0YxZG/H72pok9ojLZFYFcMtfnNilFVXhIBOzSQXhNSB6TlNMkIggQlZxDI
VjEPUnoG34XKV8B/qq4cXGmEOi+QdyyuM6RNjKadTKZIFz5NculRnvNTdH6IIDvdyEuypiZYn7IY
SftnwyZG+mOuQ5Q3PbLmTKZ0SoMV9kRPGUI9rYRQKmAG1Tn4MXxpqPLmIEzFVOXSOfKJla8MGUhW
NR3Cm1yyTLucHQh6DZc7acrv4GAYNtMaKeK/vc3T/O6s8mi6OlP6aAFBxaCaNsiEHOA59HDrA5ps
D4GvZ6Xy5VyvzR75L0z8G714gTUZXCrpeQSzKsSUpyUye/KsxBDQG4sA48pvv4wLV7oOqfnRhmhh
dUk7IbVRj4bmoipRojxjCFl0Bx6mVXbkqhdsWjlPGwZSJX4njDNQ2Fc7cpguF96xBkBvsKewULQf
fsB8mnuX79iwXfBats1wO4WaRrgF3ehaAA1NfFnfCAehhhuwDd0mVdXG6Wykrq0/ZbQrGKIiKO1+
4YnzB1W/EKSUkd/S/TS8MNsXp19D9DS/BhpYYyiNk76x6wl8+jIV4vxnbKgN0hhrh4TpOwdCyANp
/1nkKC2TVe/2RZnOLrPukTGoD8/UkfbfE2OJQDz7pzPjfIDVKehsYgj2ao8ZBs4n+0gx5dUYs7mT
H+1aSJKb7M9WD+25YvHhjVMHcZztyiVT+URtM+WJI1a2k066JKiR/ZRwNhNUXtWUlq7b7hLfdVzi
sVX1NwnhDmuagotfUpiKS8EjsL2nBPQTHq3BSefAAUsYgGO+/TVC9V8A/uJs/jo3X5Iu7JG+mYZK
bezBMsYS5fLDl2Hkb+BelbP5NYOx7P8aYHY3itaA6Fh1iK/PpymnvuMVf1EseUqHs1Oqik5+4qqv
A98l0I4tEjxH1hTwvUnIU3a+RNgBXOCs8ytrrbWK6ijppU2BYbcC4V08xpf8dN+7Sgf82nLwfr9J
NtDchHo4FJB+QaBxLuGez8m9oaIlH3zH1VCudWIeI/9Iw2NheEFH+tNMrmCAg96/IoaDkndeae6s
a0/RPsFRLGd9krr5AwQk6aocwIMEfmp0vLeftjbkYAMp/xfw5Kpy208ot/zUhP6N/mFfa3eovA1i
bxkCCbuQ5HENmCBVTNViXxyZmES2lTpYu3jvH1mxz7t8SAcVvx5RrE2NcWVEeE9offo0Ay/4i+LD
RQwAd67NO9NYkaEvsw/EUJjVe40OP8tTMZhU16qhjv51pPpE7EGKwHt3kJFTrQX8dYDLP9BDpwXg
U+Svr1rVd3CpEkuTsxEqSRraSb3b9WAUE0S465EJ5F5uGAuadz+JV/tLZqKWT+Kzxy5AZagqfX9o
AuiL6pYc85TTZH0PWnJFYi4I0Pt1PHvRTeaKfCP4Yy8j3A2H0+S9/KR0/zc8vJL6gZYYqjYQL+TH
qqLZcM35zSzo08k70N0Q9x/++GWn50Lnc+PN6Mq1MGNEVHo4VBxrAvvJcgThAsWfvvGef+PxkwNA
VQATScHgCEwXFn5VQrJlqTw8dGgFkXnN7dp8HoI+KjJw4UZ9HXUUZeMAfxuZwMADf68ESDqPLLMS
HfDBdZCjB5revww3RhYn7xoi3wqshDjYCygLILpcUEeggDOO32ddCus/a0kw3PdvAwBtyEtn2xvq
iAXJtCnQPeiwNVe60p9mm+SMboAD4gI0YZbtK1fXX552+gTlpF+m1TWlCHQS2KbnNWq7RtKnmDnK
sTtJ0bR04mUenXM00A4HkziAk4fy0n5/G2leVvggWRzxtlwKTWP2vE0jI1O84jkDrdgQUj8ommJt
ViWqZQWEXvKTOb+wSmEiaiJdm9lZm9QqoXJcLJeBuiUQGuMD93CgAwJ49ISwwgUdy2lLYMPCgXSC
exq8x+XYsxeMeNKWs80Aj8jYB0XePSAgBEpsAii7NsneELOFf7hP9JP8I3BMMa9lMyx/6rtTJ/O+
KOVmqdx46f/4LGESMKc9GxV+8chWiAl100b8LzGp8qOR9ipZD0Lkk/Hb4tRLtiwpSan6gUm+ZTO8
3QrZq1rkRbfYlFw48+VNvJsv38grICXvMJ7MkwYjoYTA/yS9eJFllK+MvTwY17P1jqHQ9HKcDbLg
T0cSs62ktPtvp6UkWNyx+Fh4o5QSC4f6MebgndUq0MR+Muc/IBlB8OX1fPySOrHruoib2Fvkg2L1
BQIvYWOU4cgWjGXckP2/Ue18XCG5VHQPmSX+RMIsPbp7Owxa47yb5F8dkm0uVGNtD8tfvw8ljt3w
yYglLNilf5HGg965cNW4FijZYJS4KomVcmsbnKU76AXdqC/kukE7FzzKaqtZcSZE4XhogPONEolH
Q0Fo4fwhQ+9aVhUuN7s9MV+ZDEdqt7xWFz0i26RQR/EN/SuZuLN+LyIo/7zArGv+Ngz2WWD2XxLB
beI4iL/Ouo5s6YU9f16aoIyr4mmEVYXeyj/v3DF800hKfU+9/tkFWnyfMMDYvO5dboyrIUG3+b8H
NSsCMKcAbXR/MB9FQX1vtBolyXgedXdGXJFk2DYjOBcmrZiLIhUIkzXfyxqQFBMXTclgwSEIc0tq
dmYSaXYamUyEoz/yHYGIE5LbRDhZUcyMKZlkNi1hpwAxZk920ZyVC1OjcUBQgSPGxAaTCIl/O9k0
OqcpAFRrZRve8LQKquIv+9s+GvnIgHl63VwWnZDUcDZRZd9ULidu/Ti1TupoLFj9ktvjrqYo3MSg
JsBu9zHim9Ll+uEw9yEiAf8K0G5J2XqlwF/sCzZEEsyWwDdcBZNbClaR1DeQkGEw3L42B0UVPXlJ
dnNcfkAcQP2KBeto7MDd0t+pegFrJUgLWdQWUCqtxbrkEK+XC4IBwyMybWn5mrwT5yQ3HpPtGjmP
Rae5hZeEXLp7F7biK9D6c0KeAE9diI6crFZs2enYM7njAwjSi+4bpRfKcFJP0/cCVbfeCQK6VTXC
2Dz1i4+UyHjLil34NFkclki0Wn7Yx82wkMAbCKjvfzzvjJE3h7yQlMhZynWDYUJExatqZx3D9eZw
aEvuyrvMnWbSEtPUx9XNRCBgq52/qAqVS3Z8adQBxbbc/D8YRuuBTO27NQRFhRMrXIk4K9CJdU/C
skiEhsbsZyLt7Ljt4U27J+nMlEog/I6VbtG1BKNAuoxaJ6nnkpi0louLULXi27j6hO1u2rR0l+5g
VS/Cr/lyChVNO5pMj7COmVsC7c1Myq4tfhaguxsu3QMGvA5p1pR1z5S8jIzKC1IeNP1siA9Ok9T9
gjZdjV/YFfRvlsNMRMkfherI6OW+iw43v0UbWfmC2pkAGs7b9hmfyUpUCec/7peP//eNTUuhSfGj
zutBpFo8Zn4Jhfn9Ed44XgfFtQ3ft0enw+bikQd0mlbFzg/Aq3DCN3Wijtec2TaAupCRlwSBNIGg
vT6Nk2g+ixyiIjzqSjASMoT7hUcmTjIelRFLhkvkBpfeLIrFnPjGFoEYrzxLFKKnZclVdso0SMBo
ExfDStJfGpAJLEZL+jxDKA0up35sY/uTZurT1T5mIjPjee7d67Dnf//q4YGeHgI01tgf+LCN+GT+
OnuHLijIH6YHdgD4bgPuYKcxmCN3zQnUrWIf8XedQ3UismMEIR/zkvEeaxEUTh27FFpRnRXshLfw
h11a5mx/JjU+b+plXh+7JgAB+gZvrTHFLZ2PEiCkUUz6R9NCUCRCtmrYK0fp9DLGyT14qlXv3fCZ
OiDGmyrgjcyU0GAVn/jtTkMfnucrA2LqYJmo9hS/czXxiG9ZPH4bTafX/xhd4MYvD2x9Wk+f7MEZ
WFt2l0s2dRmQkNaFDjRWwvKwLNAxRoFD+Iyp2SfALV14TN0zWi71jkxaQ2drjlDrOmuW31oNopIP
SHc4ITJsZYKO4Q1hw3OoKATQsknJ1frlSHq3b5N34+SD10WY8kbM9gIiq0ynINrdY3Hk1mwRtR1W
bTjh0jTLrL/Dj7Yqa3pG0NhtClFpM2YcYf1P8h6y/Pq5m33rRxMiqZaNlKut19OCnjWS1ZbZV6bI
BYnrfmtdS4cES2oDYG02tf40RPEEXlL0enq0IIRvrg5CymM7teaxyznFwq9zuoTpqKq8LQsEdhhs
cUyPFlpWhTdWQCh4M8z/c3MZYd91aYYC6bX2WNYG4b8YhYIseEzb1+mHGQUSL/eCzuQde8Uw74mv
C+RtoAKyt2eP0lWQXsIyiT91C+1c0Ix5nJr9MXowfocE4o/dzg75kjO7XvBD1OS+O+E7Cit/eiho
iSrpcW/Z8Hnw7C0QywFTO3nkIJ29DJTogqamOMoJI+qVy0A4/Y57pjM89NudVvNEa0CnNBocLd89
xYa5GwTCSJRdGBxvRG/JhKqmcx39nj1K3/2Tg5200O7chRgKhrODHVy8gHE3vBM4Em4HL5xGya0I
GBdbG37Apwn/8cr0CbkfSkjJYC64X+jay8sN5U7vw/enz2MnRgNGyaZp8bAyyNCZ2t2EWxJRjChy
F+8dvOkoHJAS7xmZHP7te/l8GIh7c74TkxY1tmFRM2BrWVHZAUya1VToMlxPFbVKOSuaI3n7hKRN
/1ijtCAXcxFYCwvEHE2Kdus4C3HHgEUTc6MwYfs5ihRNbK54WBOTO0QeNclnSvdGn2dBz1Wk9sMR
heGT8KoseVXW3NbcvZXZcTiG0xoTqxenLmzfv+gPqChhsqR9D5NE+h8GrPfzD/GDrCtgtzdgCDJT
y+ZJBj4jm3TNdcVg+mj04vypxSwf3i1zouUzQoEfk1SW0rDOIk1QDdkCFnzIVPQvvvtpmEOP+v1J
FagL1k6JKpR0zvsBd10Yi4R6rmR1dcLYdVVpmUtpY+zWBtgW5ujOJvGBesqtY3r+UwoqO/NwUScc
i14exwawT0nFBpLnDfLsEV8VN+iI4j0AIjkK5R0YTnYYJOYhWJeTfITIy4bDXrKu7gze13089hMH
Swj5czzTJWP5Ql6kRRz2wNLA0B4BoGVpgf1tOeU7jY6Nld3CEHD3rhR6DM5hLNYOB9zQEJBseeYb
5sNiCRI4evPzIGWeSYrHl2r4kCeKWcaonvgYQ2Zcg5a8RCehnV4tOd8u7oF4fI9kTKT+Xd/XpltJ
IIUcT9t9BPvm5MOwwZoljeq/0VnLAosQK904/ql8Gixz8R2HGU97CLJto1we5hj2r3nZJbBF02Ke
f03X6PDesWMd/ypTeBsH5jqMIDFiywHilbaL4C+dvt2n8aAphwKq5tvOu0GF3/h4bpGYuFSqzxWb
95GQ3doLpMKcDKsKsDpE3iJbwvGpJX3GlsDRl13Uw72llN+UEchiv9mFkqmE7trct+RcO5GAMYQt
r84G7IpxyOsuE52/H/zrdJ/sy/ktk/GtRhYjkRo8IHzKQ61DLU6acEEj8D6poLVakIR+Z9w8v1mj
/k5A8P0v2wf/RXCe3Y8BahkeBJMqlVhHm8dmN/+Y9yKXZnXcpMWkudGP4oYD6YSq+l8LKrSw1Ecg
p7mQHU0yfZ1M2TMt15FRKepTrB3euPmnNGaDW4qp8tHt09lK0W+rBbEIA9TWtk3EkZ4M4020ALFz
k4cu88kUciUw9MKRONaJA4NigydmvPdptDfDcmsXdD/PaCj/m4FhZPGqyjKN/fZYjixyhPDccSi8
QRiiNTDX4/r615aHLm1BwdCLZAbobf4LCzh9xGLZo18lunbPogaJUi8Ni4cBMextHsivDvb7tnxx
W5cVI4ffkX6EVCYTOastwBXt4kxoWMW7jWs8/yQIXgNMXpFQmoED1ZiAXTMhEf9tutpv4Et3kHeb
0UPSjP29ECuo7e5WABR//2+XSo9iyqEYGGYiyQJtNZL7IXbyRkkajwMiZlAJPsc4rtGhig7gzUbR
yBGqqxU+B/02Snb6QWsT1aAZb5ztrZpkPZBzjchY8doW3rs0zDwd88JD6dm1vOqTuFMHENE0KsNt
NvUV/BYnGlZYSBPvY/PZM6av/qfBbx80IKJruHa736iZVfo56pjiSPJDvFxUvYQmbA89sj0BSRJc
HgJThlnGcDVdHgbJ7DbVnC8556I2DCxO0iLTdrk4pNl1vpd+r6zZUoBfQbxwhy3nfAs9g55RFkLF
L5bG6zapFmps8UhwVScB7k/UPFOS8sdEzMGu6HVKrTp10cgWJh1TBvN+kl522tgeFsLfhPlwbAoB
zgIZPM0ZCEPUWZBlCA5lm2LdtfgivjHyuQirImAgrN2ZKsV9mB5yanq3lhCVHRihTpBoPuzjDlqa
gOfa54xAGD9f1Le4YLCjlN8yIukdHrZw/5eTkkcee+8P/ioSVvv8oFmoDENOwsKuTpn+d0WHa7C0
DxwLNI+VcUmK6GSlqkImhnfLTh+RQookwpyZ+8hDPn5Tp11kC+NpRr11+pe7Eijjwq2KFf/snC+9
nZgZwchLle4SvK3BSSGCHfI+SWKaExWfsf9uDf9mw/FVTRy+ejrDZlpDsr2P1N3kSVAqlxNQQ++s
zN867IGQQDePIUEhyN5+cQcncojLe4c4zd5imWRBv9HDKZ9K9zcvLYmcqaTwKCohv3dhXWm8GSBx
pYAgGZ6o3JZHUUr02QkqbfP5joGhemHEOUQvxHeHIPCvKN54cVFgYzr8d2UR6uY3YHLmCdE7l+21
rgXbUbgGG/C7N3K6l8E1Cf3rgctUzspTlrDIulgD4Syx++2eOIzkMZLIYChAPUljgaWW36OKwevE
z9qp6RwUn4BEVYQUXjt+Hfl9yhUqB5kw0eB+pf0zTUWN3Cmgzbb6iMWRyUgDueIb68GfD4yA+RSW
Ld3Kma2rzb7N+W28PVMIPicCEiPXP5dovy2VeXZyA886rjOnBAXIGoKpKTMPVQ0E/EIhNI5GgLRp
GAsV3xTSry6yiQS8qzzpdKnJh6nLHU3T6KDw/gDueMARvAhcnnumzPi4FR+zTheuBdysRMlov+yA
+aXoCK6CLbm7LRs0sS7Un4vFproe9G5f9olnYrUVeiwetrzkyW8gSkv53hZKDYSyx1XcLCC7t2jf
ACAdJzZU6S8OTQbEdyLX6pBrsxd4iVzCXbfsviwUEO4dY9JtSY6JtPoXj/1yIBM2Pw/z8AMYb1QL
m7NxWnSZVlIGt0Uo5w04IkKAeZynPMUjxZ69igYIpw2ylRvORLw+wcLsbeNPuxcXj4JXRnZh3GqJ
saU+KYeZxmDoPsQ4m0QvQ29tXtmU4DNrC0G/3Mwt4wRrkvX8o54sc8MAVHVDVz48FF9efR5DNDs1
Wk6HMoaXvAZHnG8Mo1Xzrv5bVB29rnA6lYKbOBOq3WjjZQsK2DWT6O+F4sUBm3rKVis1Rltj7qlY
nAPTQuGhDKXLZ6Eo6cS6KqI9DJLXjCWRPXO4YbVVFF32rronI05GqPFfw3gxoJLsU6nl7oTV5n3l
0Sf3m/8uL75Zid1Ss1fhp/jILYIaNnbCXAkQAadvzq7eNbH0MUgkca7THiB6rXdDZn/Hr44WVcpZ
FwF4RiDBEA6eKClPYhJziKmrvID+oPtizCf1vkx/2fxqp5mJvS6T0cNoPyFgP7VM+POsjei6Jg90
KdQMTIGW5We+uTayu8Z/Suac7EiYO2iXGL8WjWPbsInbhg3K7ku9ZVUaVcexmZbydopCVRn8NJZF
qEet324a1WJqB3LBOcZBSQnpnbkKlZHqbFAR7M8oVqXIcX7IdqwK8FWr9prj2ydklFC8C+MicdWX
b3P6Gk5vHaSQFeukb4hrWhEqGoKKSO4EUYmNkkTaz6jpjuJBeWItOdl3Tso0mnKNZRsfA1XcZvRU
5gHLLxOXUMwwca4sP7K7BCutky+nxakbLRLKU7JyNmmIqXd6uoxt+iHAy2a8fucunrY1OMapvHhA
N2SCDS8g8PWCTx0LJ+TPA0ZywVFzMagNnlzMAIieep4wqZDED8+sUmJTwRP+oZ+8NLnL/qN9TMxi
me+ZQtdhOT4KLg27gSAhnosFjT8fp/NGBqFQWZfLlqpvajtC3X37c96afU7K2PNCFTZ5NimCMEpO
HXUvkAi6WtBSz0lFLf2cS7eTKi/inC49iXgwBvh+JanAmtmKty1BSlb2bGkvwoUa41N0j2D41Lly
JsOULit3/kvgr7Penv0QKde4dTTskMXdFCvSEiu4ba2FgMSZMKVTJaUHUiGBJopGF1otWRCuO2kA
8nkEYZ25Q9jPwO89gTriyIHngHWl9793zvbPi7plfL8qiT12FZrX1d+XhCaaOR+FPkzP7cqSkJpr
RIqcix2YKAdn2dIxnZVRAB1WI68mE4FiczJyhPa9uynrTTfL1TcfGWQojob2NygoLXGqMRMOo7ju
iQI0D755B65QzE8SEfynTKDlpZ4NC0FDqMvdkxXtIyu+A6ryEuOrTOEuguLcYmirXladnmiF1RO0
Eut0Tzo506Z44FLT9LsMr06r9xWOJvNXvGcKNd3bMWxrNKKetybsp6UmjPIUuXASDR5HM5xNCq8p
WvSSpwl0NePeuB3Ijo0vdl29k7Udb2HzMbXK8WdQwl7XfUSUR/G11LoYU2S+koUgN0qMj8woROXV
kS7GiLAdB/YulaR1vRcNYoRvmCzroE13K2e3Fxb7oVsJZa0UJm18bZ/BKjV5qtD8rrvHXVU32ULF
M3OsZI33/gXcatONCEBJw6V//HeD4Hsfw/Grau9tA65t9LNrwB2wRCq69KYwFD/A2+XUHSIUKyik
sBjgo5nEmPTFP/XJvCdzJql9qJlCUwiJRe4nbetA7hYKYeDoMblQOmZNZqUfwG/DJN0p+f02/i9g
Y0TDAsgY6AL6Nc4NVYUwA+RXhtqNy4mY2hebJDxOf00mWqnlMTppY2BvmYLcUEgAyWcSKDbfaKqs
oARHWgBIdxABA6QhBhqQh527ROYKCHVdfo0uowNUoMmgoJ9TuW64Kwr/oFfxDbh/T38GIXeQWNxl
nYtNNpMNHu2dhxZfvITUW+EVLKS+sMUobv7kDoiy2tEIkWnMocZ7a755NCcHIaCKaOvmycpvqPS2
hmCridWr2MLRNtxb+lQTJSvkoyomdXLgYaeSfYUsKEdjXa74vZtKFmqHSto7enEwvPpMxtghe4nI
Ndder3xbNwBJCeH6wcfP9Ja2jUbB19ojZIzoBi4ZvpwMUS/0fY52hTGku3uDeFZNKsQnaYltPCQJ
LIhRBRIKTuXWwuTL4m+oSFw2Ec5Orz5NAg/iJqu+z0Jf4kO14JqcHkhKTWy5AqPzn6PaAoOPLb4Y
U6ja7ARgK1IEw1Dl+U+XrCSkKjAQAk1NgKhVJ1MKqEImfuW6FBwKHZZPTDe0EdkrB6rf9Bmsbgf6
B4v2VGRETPmkY15yn4OhnbrOhcncxaIKPRMVeW4BEyOQKWMHu8LjqiL3pJBaxf2PrVNTc1LUFaAZ
pP4/zlf+QZzjPQWzBv5nzxFtdxYIpPrw7ML96F1WTQTvdaMW2APRkg8xHUb6Y7dFOx+EwVL8fmqS
5mxKQ4SlWd5hphLYqvaI5mzuqEBXmb6whAoFdB2ZJB3xzEjMWxk2afCP0if6/mn9FknYWAXvAi72
NMe5BxsAmaW3t/Ss8GzilkXWry38zLO/+pjfXeiKfWBXvcNT59lcJE38qFierqDwbw+srFMDu6xe
tYF4HJ+Ts1IQlgC1RGKp8RXZqVQB6Yjvq56wcC+8mdYCxO2KfAWscju1lmGZadxvQPUk0P8q1WFu
L3SML3fmzx2GoYp+JxxqE6AnHTagd/ZpzCYlzG0xh6QXHwIyifEl3TsEHAA+hvtazXFEO+YfjqQI
R0tIZy+y4eBmgIj+cMaJs2/dLd3w4ftRQy73BdYXzP1HrDjmTNpF7VWHq9m2PQpcL2YLeB4fNEbQ
8Z4Qyw45gX1/1o/BJaDkpCJdkkNn3roFUHIOS50l+YPMrMogbTgwI3yyVuU7BlExya7ShFXXvysV
G49FSnKvM5G/sdem6W+0ar6jvF5kTHGvxXHcSn12D0TfgYglM+qCfPz+dqjfKugrHN51sCjwErae
ALVkFSvHmmXew7+PLH5Esk+6VwNorXcZcawBVhZIcTMLfmhisE1xmM37nK9YIVWI1Cw2BmnggMkz
TF3uNboDFM4m8flrYF8k+GJ/cPbkiMrZ74taGiIS3dtuaXyYqxzV8W+isZYvbliGG5v9znEzRFO+
28n/wSKueBhKSkcTAyfJHftgfmBtds2jtxG62Kx03Mo5PT8cOYA7LJJNH2I4qMWRmMRAanuc3sTr
/pOMO1PuFte50ok9D87n7bU6YXalRJEt8l6Y3rdB5PnW02LipqrIq9YkK8M5Pd5d/R84JLk8Ea4g
32S1YASMJDz2wobePROBmtBHgcQ0fQDXYXtTG12b0+6+GK1ZQJ6C/YL2QzeQvQ6677lERuMVwrH3
SkBlhiLDznjetaBCeZxo3lAAZ08dogIA89cxpM7IFQoBfPsKDuHtpD/ADQIO4dJs2VJs5FF2PI1/
9iaVGeHgLIqO2HWQjc9Lolw/8w+1BtWrJn1soEM8EPn+aiogoELQH0K7p9F8HufkcGMYNW6dd4PW
MpzKVpqWMk8eTR/HKqNZViugBEo2sTesLfO8HVex8HJ7cb4lNozIENmuBHMDln2CfG/meDn0Y/Rx
h4alAhqO+dv/WDR2UreBD8wiQvjYVwegQ1x0Au2r78lQRVa3tCiuWpiL5eSCX1AkAFcdWDIMjLSr
w1wyLp36SBrHeUKzj8kgDpvsKo3WGo3pp66mv0XUFLeXZiTZFDqvBt2J0uT6E1+j8Pkt1Az14Hw/
hLqDldYO1peBbz1W3OLw19lwyFs2OaLnj4bG2ALtfcmdEemCpDBNDRmhK35uEToG5u5XQ/NWVEOQ
8S6NLTDUXhQ2ayQcaOlAXdt0qFrNKRXDbYyv+btzmiVuZn25bZ9t9+sAMeCK/a5uDlVBIQqMjW6g
uU9a+NjMCuNm1NybLr+hGs80zk9E5X5UT6CUFBXQF7jeDJbx1k08XXgGMdlmWEhy5p/4K5D1wbDm
+CR9GPSmZrghV58mzpB/psgcuMDPbkti/Tgs2gzOz3ESrNY5kPrrtSOwoQ+UTSee6tDebxoJnKtL
52TF/b2nzO9Ix2JEY0z9jG+oB11reb4FkOgQ5mjo6JFMJwnMrCuTV/PyqtjAnDnFQkeke1xnsagi
19NqDKUc77Uu0/2Nb/rXSYCxyCNQgHDWRFqYPR18YWjh+zcRlyw47U7CGs1N+FIiFHBiNgfVZLFS
B2LE6wwvqEnPSQQB126L/qgolgbmLFsAq5dKJdPX+HQ7l44A0G/vpCFCLJrBX1k38+OBZxcBTIGG
WJvVbiNTI1JMU8QhS9AlmlIBO85nfm3V8mDSRyM+mYDUKSlGf7NEtbMU33McmPLOchNJaRE/Z0qN
VuINe7jM5ROSMcwin7B7WvE4uekJGC5X+xYOCYdre7VGaTnVyglZdCJ4ZlyDydyzn19cC7hblcNg
JD5xNyMLOIDKcy5E70CJgaaYcB3qjLIk7naChkKkbUteJvcwcRCJ7+blmCWMv4+/13veQ539yX27
VEB3UL6T0SPvyLxfzq6k/4iZD4jEDmPkLwyOHisDihs+otoyJNx7/ST4COa+YzCFWC7mj/xa4uMK
B6gvqLgunppr+nVC1mJvN0k3rfdJYJQFV3tG8NA6FGxvQy6c0gII16Oa468hK73TLJfCbesB2c8j
UOpX4lLddqHvgPCOyGeNdV6GUmaQZQ82P1idUu0pc4D3VsD02IoTlUxfTWtVm/xrtxkkVVQprQFN
q4A0sEJIUZSkvAL+djPXu0FFfJJzrGW4c+Jt+ac1mSF6uBBCJ6I/ZLpUgJYcKI3atJG2HdqFWfkO
a3fC7cI8V7l/j/6ilAl7QIVGz1R/XnT9bZsGE1hsFimfH61Ptk55RfBGAuY/0iZxCqDEKiaG++ST
LRDfxfIpA0F3Oq4F9ESaLLwdy39xqdzl9LMQjiGaP2skAeCz0MW2pI3ubx2CqADKoW1NEavy5ADV
7WlauwMKtMVNBlqY63JPskx4UiBTxpyz4I8IIXf3HjWjtvAk4Zdm6ItZUFgOxqO6bOLnLYlaiar5
rOoAHOA7lmg+omE8+zv7h31F4r857pH7EA5R+AU0uzZC9JC9tHXcgv5CxX9Zr+U5g7x8l69w/wwN
QTdejeP3eqqmElKS3DBZ65hNZMo0ACB9c/YKZRhK7wkH5AH6qfpI7jz6TBTxU0slIH5+/phSUCiS
UvH+lLmYi/tFvipSKhByN2Sb9zQCLZKr67Dnp+qqCTseaFlNSNlZ81MMTtj4FMJoUs2bVNu/qZAU
g+MOSK2+5HFPWCvp4ghTardP4adoMBa0k/LMxceXglBXRmQtIWi36fDcHL2QqO+ro32zzewGoyqs
TxW7ay82BKBwH9i3WppQBN1FXv/ZEVFh6T7+Rv1K8CNUmw8sgeqMCbukTmSkC51ZohBaQE6CXxep
5z7XL0iYfEvAXSSh8schQfGlyKBGcUT3i4EwRo+aLdaYqlv3VMi+Yjo8qDj/g4PJg0HW5ZAz3cw1
bz2Ln0nqt5Obiqfd/FLzKTf3At+RCTC/T9Z6JSQEPpw7wlOvLArTdZPxgyKf0AtjYH0dihSWm2Fo
HTohrNgbE5oZ6M7EAcCyyaX1adiJJzMYNgiLa3uCB8a3cL2GwjSvvDMo2i81Q4H1xDMtXRCP6/sB
0TJr9RiGrKK7K25Cz5E/hE96Uc/rv5Hic0t/AiAsbbYpfcSUjvdaqzwwAQsS/PNEdM2rPI38dP1i
IW6zKxV1QPODmSYkQtiVS5EWfUOGiNZZk0EUr9x45LCoEpnySXsyesGwpK8fwJrwIR2ifjWrmr5t
h9/cgnXG9kI+jeR9B7Vlx0FovhCCSk42eP6moN9ikQe6UACKoJQYPPQgUTlJYDG8Ed/tp6LfWXSF
k+M+Uedw/FPVZBkayr5xFkItpiWFemKiWmEkQck1fDlI36ZPZgc3MvTnJwvzene/piI0biFkBd4m
1laD6STsqN3m1vCzNAASwDPOO6Omp4gYtO3VpEd0swgl2rzYjASiWXiVUWXwxDrNMSG4yzC8i4iI
wynGZgHHYL86R2ifFgmdPljqJ461cB9nMCuW3CMwc3TIp4TSvSca3K05nfoKrtJGHqECP0a5KEhB
1pfBlT2/Qr3c6j1Tz9NaTPgM34UqyELr5suTwPERJ6L459WNOSRKsyIhn9YtMzroGVS5FKiRSkwD
PU92/+/KKStGBjFEoPmGRWz0dhtQDlM0LCc1ixeqYXH7lYAx/jeDgx8BNylEDTJiQ8YLXRemBz4L
amMISPOb6bGCGMtBLVekHNsajE39InvCkbVLu9SGYA75Zgr34ODkT2K6i2AWFrc7ilFzyzfqZsbS
VtveVs3t6CdQxq4i7JRlq2RCsDrN73Igi16D2qjw74m2XB4nLSZ94lL1Z3r0/xLRqbrvNw7BS5WS
iZDm3iOGJZEocOnnZTsoB4y2FgdDbFBeUpWFIoc1nwMzw14uWrfdpYz9/imFeiHDKkQXArhqiSBO
T3dNu4FUnOOEZL0ULmPOfs4KCv42uaMoZPB7CluZeugyfusKRYJTkaGTU/E0zOyOqirE4aVtqdqp
iBiGanZNbOy5sQROgT8gPS2cToVONIxJfOFEJ4pxwGD0csvWNZjoeVjsNXd1ss7KwG7R/vc71K73
aJP523WM5Yx8EIWdiEgW2iLojiOhPKQAT/5u6cqd1wJd29OyDOC5Px2j1nTlrKFKt3gvdfRwOIDV
FbbDebKYndH0+WQ1FLsmg3bJyw8WENvOcuU6Uj3wT+7cEd8DktU4YjbVo6n4F4CC5oFoy/ZUX0Ni
Fk3iewtuvWQZtlxdkHb8u+uo1UoM595Ot43I8sg9pvdbwY8U+75ZhfMAxAISSkvrIVnakSRd9ruq
G/lu5FFdG+vR8AP8JV+AsDzsdkDmEhKGxAxJe5O7Bi3zfKGJjEoDHG4O7kB8SpojC9GxUgUgi7+2
ZEJw/7O62E/hW81WYhzSLQCvJ+6cn3VgEiWp3EoQCf8ox0P1sKeSDSdMF57mnI/dKqgQU8TVvB1l
8mQkj4NUTDoa0k+u+zaHvQVeRWHRP1As38mwRGHEVEAtWTWxD2eDm4/p8sBJC9NcQ3mBzOIdSE3L
2l2aw6WRvk/jXv8G2GrJCGVF1CvtnmlQJSoZ/Mkk82WeL6Tlf33XjZWT1hCDL9rSkNybHU3yf53V
XuW7Ljd51R6qqTp5JHQNdlAmbXPOQb+syDavnJLyJ6u/zCGuqCMGmoLSQ2BLhersNJA4gS/EvXXy
CFW8RzlZn/28phr5w4yZYxIopcpQ0RGwBdgaJbG3Cj0DO8zzk6T694D9XaW21UtqYMCKEmVwHVpW
Pdm4+9jMDr2Y4XEW89/uHuPaUpVRlxd1foqg0VJ8ITLdz019gJGVtBAYOmFyUPFSz2gi9w1p6qts
fT3GQHoUrlJGWkjgFESk1SkAKkBYYFWZ8rNx0qLQzzlJBm+OPjssqyzBHyBKKtQWv8634dqRGFXY
AJZeuOYjAcNeaUYNhQYPNPRBagEdk8rwjqAtGdtmNp62VNS5eKZ/nC74fLYJRFgVNNyLoGIJ55wr
tEO/HfgXrTAUjPQKVnf3gzld5szjTbFpPaODSeagE4FHKR9XYNId61BPEXC16XxFlM+2G6Y9pJRQ
8xUUvzJpWzlWxYeiWHET7d1g9ks4QgBtwC80YzkyHdgBd0kZk35W92FUWfWlhvYHY0qErfb8Limz
DJXbIe13ld7v1cNeSsg+hYIMVGL5G9Q/OcLcJSyqFuiuB6KREPIyfC2fAokosGHL5bMkrtAJEccV
wpVSCYlunINvvWbwN2I/qtGftqfRkufTXe+CtpDM2l1Ho0S4iq/SdCYDUkdtjZyvjQEeGeH7KhVY
SKdqSycHrdrkIGKZQvPLJsKS/GucStGWUMg314eaqMIbR2knRhsyo8DI7lDvuAu3+AM6Q/O2c0Qd
tH198oXHZAeqA2Q0Z457j1PXhokLCzhbD9wKtSVDQvCEysRqKKTeMHUKzXL7kgDa5UODDHpDSwN9
KnjrYyMlE9wMrW9V8Kb8EOZPivxF2yS9t91oKiRgkEAtFgKcRevMuBLbtxkYKVHd28W2hctzntXE
jgM419W8wdb1KBEGlc+hSmM/3oGDUy/EEb5UOmVNRZZxBK1rRYNmxPVQQ5RIWCuF/5jKmr6v4jCu
dPbgc1oNz2WBTRAfs947ZqcDEF6weMKynxpFH4UJyzQYLQ+uBcK741wPf19yoTLby/1Jc7rg89nk
Ae2ittcyOjwbX8CSU/1LivED8pk0wf+xZLWRIGJU6bhYH9Np0siJoOEsSMonyi0UTHv6KyPUN9q/
UtgQsyQ4M8oBq0oxLmc3nC5jayeAhk/OqiRYOBXCXng0L4Zfbrcoj15tHK4ndT+setPIrMPw99JK
vrVSelVyrvDb56NWjOU4s7Du7y12S+jUPxjx3ZP6282GNo3pATo4DhoO0rzaeFixgR6VTAc+SfzQ
ToU0LtyDVRotNCfUN3AGmGUQZXbGRwx34aTYCFSn00tbrjp8wkDGFNUdJrYrry1jZeshbopjix7B
51s7srTr2FJKvJeRFOwnLw0EaYRvTT6/DmLDAlN2mlN6Olr+lU0zmGfmcgUDfFUQn6Ap7a6EvKI+
anS/ZTauxmlH3Bip+coujEBdo2uXoALfVw1T9QPGRwp0hwvVUHrh0fSc6e+fzk1Unga9avJY29SW
0yAZPO7TsxRqw7nI4wNOSubIbnGrfQypVbDtorV92yCVK0og7Yl45oG0ZkryRZ0SXDIDeA3z1Hey
9lIk9FmNaJ3tsePY+lt4u7BG8dyGutu7jpVmB7qNtajhGZUU+MHxrnZ2+zAThEIdDfXiVjZW5pEY
NZWrIs7VYgf9EhmV1XJo8UBjjkTzdX6o/vJNBmAw9GXlnVmFXwd5NKdW8zep1VWKdvQe4G3I/jYp
/Dc8NJYw0XW1dcgazWj2UJ/gNV4U8BvRIP1S0gSpoDTkSGtCjiIubUofwY0Uur57b3vtQCj+5xIw
N1vlXSMJgLfv2QlUA06X8bljwQKjO2iT4uyjd8QRExGIJbaSl2Jkc07nPGJBGif0F9mEw2l9YCaz
EwsvTAcrbPXq/ZpZ11F64j4bN0/yAOc2m4klwTY78yYlevF7DHGevPIvsDkdvhhddeFj2w0jhSLl
1g8p3dcUbJz7xNEji7slSkrWvxXmbuDnVPA6D1vYqmWS7N/SkuK+JoFvoDXbAnmQaa+a4ApvNk1M
V3vp6F/sR6RI0OqIfluZmj44zwrl4+awo5tHHfcwNxwGhCSvuw0tGHmzyngq0hEw3gVEx54SjD+i
8FTjzBws5pa3rT4GIZwrADCpMHCOGxissmnGdYLVZZnTznSAAoeFxZ49TpicbrOU0AjZJuR5ghrC
yIeBHhmvJzu+zT2ajTIJe6vB5PAFqv0WAzlO+GO7jw5G0Pw03nNQxr6dxeTnoywILQ/keRsad8YB
NFjlYxNKasxi76kg2aS+SCELRYQz0doPz5kMn+iWfKmsaXJYfY8K3a7pE9fc+rMa2YXokC4MDmEs
117Z6AbVmk3gZrAsnyYHC4YU515M0mdmc4wKekHhuKvighEbPG+rE3OmWG/Z7X0sBl1mYAIbc6p2
RCsCJbUbNhDz9nxTFIjH2Ple57pAH5mJI8EW2tKWqyvSVfsORbRze4C0Z7o18ygCgkfhQWkt+bKh
EFXLLgQnWOm6Ap/yODu4dGftEdICzJhTOUF7mkMmOluaXWCJ0hg3YEtZqWwJLjezPtodojNv+OqA
qi+jPjdpRyLuWeMT+tqvGauHtFZ4RNG65/0R0KrM8ax8dedr2uziveor/Bdy0EnlrwOw1EFiKoAa
DwajB41Umd7IH9l60DeX471Djv8A72VYdaE4hzoeb/E8JuKUpq6PWA73nhmXOdt3XQuqjKl5/gGD
zxfDpBQ1XcoY0ImY275l1Mm/sr12CfiD9731jEui8AMml3Y2EoVdH3bI9Q5E8uqjyoy+l0WRlVN+
lv2CdSv4MHfx29yseVK0sgdwSWQ1Jm6aXgu7JuJhrCyxiO9ZKVOdSEpoZ/JIdcSWTF6/15MbZT4E
yFOMIdul3M0/EBAlPFtgmyvX4Hiwbi97lakghUHKn1uDTraMjnYUjPDTEXn4Ko1l/0UOS9htJ1Xb
67TI7VlR62xSwH/O+xL5qyKB68HVNHLrd4EqkspKJ5Inb3+K4Je35l5vb2tNiqxm3M0wt6P090fd
1yrT1YSiWdVlGfe37PCkr00UhVd5LQCyAFAd34VHZ2INCE8CJH69y/AIe71NBKvoft+TvpI+OieW
vM+3Xu0VE+GIfP0N2wmEVK2Tooy7kXuZ9gOuCgfP/nUG5leTkuveX5kY13nDPjmwK13F2dXoewXN
02qwBi2HIPmBF2uJo5oLQxfXFsdC1eW6LCblkKYS+V/bmBctLvzORXFG6CB4jC8XheWVsOjNUAM/
JWTnJyTvBWoSCk9oY7Q8McqrOJbUbmiT1Raji5dQ6hH6xumaiM+DYc020FAkUXPCFIx+TgXNPV0A
o4FzwECxXbB+vB9BgLJoRHWU+lrriFhvmi5acPrMgIv1/GHjkbFKCnb+KZSwNfZCYHQOwzipUblQ
aaiycC7MHnfr0L6hjPodD0gDLbtPdusEUZV8H6Ksi8V1kBSI/ANC7rd5c8x7ST00C7ZnAJp5oFL7
wZnRaDuAffpQH0Vm/WrFqQFH0ChdcwH7xupRNUkJAZYu9EmqA9qvUWnfsXrJGKpRt9Lk6mR6rM5/
JOS3mKDNqu7jWp6ZNq1V4VkI8D3DRD8ObPgighwIJ3yi0NFAVL4mOUjxrSC+347rHZMDQS6EMwKu
vTMSPrCBmY9NsJgzRB8LhaMF59WViT4kCRbIT+L1IZWWKKEGEJQQbUUy8YLVrAKb8nj2opiAFdzQ
hysD7o+L2x7YOsDC2WUqCmh03mtBzPyTnjhZYiyC72MtG5aneor/KVGy0VVeL66QC2tvc/U1lHAi
5D3dScSwJugCMcZ5lOO2Ff2ukqjKbVovYTYZ7xf+DbnMci7IrEXu51A8VYesHmPXWEVzHFN/ZkyS
6YbWPTMwqu4PJIjVuXWOmDbqRhfppwlXmFlv8aUz+yDu910V2dsK/6aAZODE99IT8Wbx5osNSFQe
XXJBEpLQJqeQSpMxOoBcYQhYRuc+X0NOOAiLiR1aNRwImjlI2gX+20GWGxcQVUgZX1L5YSU/bsnR
tvmv4Ok/Ig6FzrkDCU82St3IjudSb321LjFqBuTqAshnHVrH3FkO+scWAoDUsDseuwn/GkeJuAhL
SGKXIs41z4pCenJDxjoTa1HV+81VRM11QNcMMwdUQJKSXipbCeLdvInmuWZxKVOmouFZSJTu4AeI
dcgShqL1WUMvJ5w3uOC4p85ITOX9zfMlbD2il8q1A9KzsBYqbX9ADcMxj9FNDqGvU1sv7vIiLpZ5
w4udbKIENsrufm+39aZgrd3eTPsEOdWFaKqtb6VmNSuEd7gtx23KN0lUtWDXmP5ItxuexshiGCpp
k+nD5T/LFIWSffF/S9RBm9ojl8nFzSE/JY/sogl863OSafwmcBHpcqCbDq8Qq2+QfUTLGWdn6QnB
Zg/k8qP9oR12KxLQS15tJHhDhkehuZTwVGmCk80xizWqKaHLb3dCpP8leHbIxUjoQ0tX9swjV2Xt
Js7HuCoGOQbvZiVcUbfbeqbWgCkNT4/zAQImKurm9jJZ6zdqi1MdZ4hT/Eo3ANjtX2CKst/yZWMX
dUIXsQmI6o6QbBy1V6m75Dv1T9lUAF46AC/AepirP5zZleGD2RgSN8jDV07zMQh6EFFnns5FkUlp
QYS4kdbsHf61+OX6trsjCdOJZNQUMa2EF8zta/ytPIYb22NqeXBrPSxrlqpUQGcQtMPu8tihlN/U
DGpBnZEHvdAYOFTCywyGlDKH8FsxeRt7hJm+Db9iYJ0o5N43wAkfnkJ9H3iMNQGvEoiivurrK+/g
M2ut8DW3qP4FKdCaTXrWJdkcMlekfGzXVG3PikQusCUbO3uIeA9iYauOa5yN8ngekU66o5BbA8DC
ufKzqJR4HtbOKWQG7ibY0hbrGCz59FIXj8QtKkHBDvVC/fa6xlnQGn2Ekv7rIcm5VnCsy1oOodC5
TSM3l8MbHGlmxfZ25BhavQxBsQ8gq6T2HFapsNfjJzdqFMryzM2aposLMW0WtXxQTZCeUMEYIDvc
P3vVa/rp3qzcMjEntDlwbGHaTDPuOwxntP2gREXrzh9kv++D/20BKuE4nGq14hnX8XJ9MipfjBSH
GOadLqy5NoJFk7RlQnirFSeA5CDbXt67B0H2RuzQYg5AsP9Imyh9kXNyxMiL54+/RRsnNjl91MKl
XYwGYm+42TimVfOWPsPNvw46jwzB/LWRFxh78+18jotB9oA9wsBIspWgln5WL0aiyYm/S5WJE5pZ
FITba9IL+Qf8Zxns5oPeKIVomd10pZ4jWdDN7fTcs8+jAVipRNnmLS+Qnk3uWScyIwGD0yO15f1a
mpnHaya5GAgEKS49lkxD6F8PA4W5Sd8lNbuhh/iFity4qy+8hzgltYZf6+ezpxKv4Hy6XA2TxtHT
OzZy6CTo9zY7MeGtw/u3+jW4w5U3eNd2IX1H89fTCWvfn0aM6WLUXIj8grGoZX0tKyHi5kstutF0
PGX3gApSTNJLMn65auGUE/4f3TZmxZ4piJ1+oOWoBm+G2sJcBQw9QZthwivd3aBTjuZwHnmwESBu
R+Lzb3swS6hFquYhJfl5Qyf5BSdUw3Ww5ZlH+pd84HxK4iZmZTy1QoyKC/ft3B5JfqbDtHRgjKz6
tUDKmttwEk8rIZ1IsyVjtJEB1mWMwaeJ2iJvnazOrU6k/Y1YcLnq9guuJupWs8zs/g65n2SUr+8K
BpQ0E0fVyswW+L8ko+CRojR3yGr6plEzPPsT3/CMNttnz8SCJRdpDkYt3hvkznuBMeDa52pBP1I1
88ZI0NRs8Diao5XJ/5i9h4RrOrBdC7w02O9MKvIwbR9BE5B6dfr3lbAIudVLqvzlkvzOiQWiyffb
bhvhtohqpOlxiZm7DvxMXwl3Q8hvvH4YokOer22ua39mbY9X7MIGjSYUkn9MuT6DEwjpSnJT1Qi5
pNXqaWwz/aYaKtEpM0Y3NdDGQRJFiSgXAabSBwVsJR/qfbrfA04BxRGjFf/R9ItRAruAq2brE7us
J6wlRgj8yzK89f8xHYVuWzPqIK2atEsCveGDLa55qgEvVXwchprcc4yPuOXEUoC4ZmGE2LGhYsLr
ccZ3OZiqf/YSkfdGdPrlI17xKui2QegogUAui9cWKKbFAtZQM6RyZfeF4sbc8PS+VZZJYy89NcoE
6xcpJNecAN4gEQ+B9+j7mNw99RlhQn/MhiTI+InpEGgq6pK1PuUtBnKnGhETTg/TTQT7UtBrOS9f
sr2SQE1ndTFTcBfXamL/Ta4Ao9PN/e2fIVGm/gDXpanpM4qpDavVRUMMkYAfNBtViu53fJmMdcs1
F3YbcAsdUuXFkW8HL4PRjFTJO4GCPAOI44Nf/6dJi+JHitMfdphk2UXSRGj92p++/0XHTe1pFGnO
XsXhgTjlxHkESoJOcr0qHKdrZbcwaqWziPYSlFVx2f23RBhI1q/8hsZs3DqITJK+ILdhwagtsXly
SIrsciX5vrSuKitQqP3+k3hFqv/XAHxrSLy86t4jXpKA0lk54FMXPIky5oftDAbz9e+tY1Co2++s
6aC7oq5PB0YeX52FAFhB/+eIAEyqnAwIVXPU8LEVJPFFuI87bPxxx9EPeExFckYvlG/kiKPriaSm
EaacnDT8iUFEJFg68vLb7yZdzU4beGrcvDxYhYUZyvnyy+xCJ0xryDgRgzp4/ntqwowin0/aqBYK
GNtbuROqDe0lB4y0m6q8gAe5lJ9f0CCnNebYchpF8bNdef7ZoqDMaSuP8VdBXoEHc4L2dKkDaTHn
x7uaHTqnx16WAzrUtYApLfMBZfIPQX4RpItzEUTAeZKw9kbstEehLVsTbYJ09ThLY88cCiCthQAM
xodqCc8Fk5h9NtW3yQOenaTlWVcCrXpuulw5fzSFexaxCs48bh/L1h2dH2zvOa9D9W7k7vpghFk3
YHZztboM/RSB3np9OAl9MYeahGGhsIcQ9250j/rertcjRQO8iOASF2x1U0qN+4NqF/nLrB4mImJQ
6l0p49FILBw1aOM3cOuNB0U1J/TPXMrRvhc0EzINc8ThGCSgNuISL2qbRK5v8+d/lsxsiRaqE7AU
QuDpFymrmn8WQh+jDSZC1L2i/Ae9D3xjbi4CwqtADWLHGpL0FYUeOFqzHOouWk7jfqwqUaYalvzI
mWlBRtOAH2aqFjjmc2OQBUfH6sUIVCJA/Uc7w3UatucT+/PomKiol49yXtfDttUBKaxh9MZZAcXY
/+QIkmlkou02wROJ45IyZnm1lITTo3P7E2cLfbrZ3lMmsRorxj457IaGvTfeIOuOy3iRdMMxeEKZ
E+QVqfi+LaNuPjEh4VmZUW/9m6JXFI77g1G01kIqQVkekqa/d/EK7fcHXcuejDjXrX6/Gt6ttjgV
ti/X8EWyYgxaWoI0MN2fcko2ye65wABK4WsCJO+IkcPGbBcu32uzGqog4smf2Z4lCVhYt5bdkpVG
tkGGxjt6m2sEaFVM8YWfdqqS/jaTG/7oKZuQ4qVaW7gDkscTG0hFi0f0P6eq10dT6GKAxCdvHxTO
R+92gDyvi+QzPl9KIgVyEhGFATGV8cNPV8kebDvfh26L1zyh6Pe7//6/yxYkKhKlwuzoPvl2RwrX
kp0ZbfZ98NziYRn40Jgvpp0LJ3k2R2gk31E9S/WAq4myHJxIJQJf84FhILkw1hgJJa7xAvL1Tt+x
opITUOEoBgb+PJbWlFcLMstd5PBHaScmIhRebyQTIgr0uKOPCiR6YpLq3XgHcQ+WpyLE7XoxmQc9
RlMq3Hp0YYik935X7Bx/sEm1GY9gi6xI0oNCslqiHaMdMhB6RJZYl0B8t1mjbcxLWd4/KlMMPUek
QTrA+QbEpxYRnXtQu9P73VSKoZSVNM3BYcr1hgcj4olshkfIcjDbopGz2aLAw9Y/AmhUdHz0ixrJ
uMtH6X2yPf9mv4AFmROxJXWwbOvoeH8Y/MIYaK66EQNBGiFMlxALxJugN5wbDVIlk4VRojS7kUqw
q0kzPMxgcmxe+rMNl4yCqMhl5xgv/GQKpGPylARstGUUpU9yAWO+p76H0Pvk/jAD9oSC99XI5g5i
5ceyF636ofuiCGU8nvbuiXEbqDBJ4m3OVWqNaFfltZ6Zdfb2m/B82OPk8699F0juGdYo+KhpmHGB
ARvHRvlnff4OSi53SxHztBE7nWqMOJO4R9MKWmCSmHNpDI46Uzn5XXLuVncHJ3mKIPTittdE8HlT
W9i4GNUUhBWyheQ1oyLhfy115PJ6mLiWmcSqTLGH7ip5NNAt5LpC2onkcjuFqdWqYiQb0rJFh1iz
Omdj7GFVtlMx7pLpjLqskEVf8iExQ5HFMykd+b5rh3uUr2gEd+daBNIlrxlcpGxyWM3tscbSB++p
+n+kd4+UNAjh7ZMmPnyyOmd8bohzJjo437q41WY2Xi0pqcMbVnTE4SnUEI8lwwV4PEj/hviMJMaA
2NwdgNJyD5rbE03haCtg8gBEx2s6jeSC+f1a8IEGreRq2I/6mBLYEcQOwhUy028EbqkvZq2RPDpn
ILPAuAWRTPz744tUhSabuI2MKC9+7sEOzHHa8AgyTP0/kDtLJsebUub/UXZZco/wvhlP4DAnFzpW
Py98s5I0q6PR7EzqFDGxlz0U4TiKD+mKFTrwOw66WXCmSFOW4IZceKSsATGXkQKg620XG2wUIMpH
VNMhQKppjxiWH6W2KA8im8MnUMCwFE/BQVzCaN6bpTfoN1hKOXWpcXhvrLL0ZhC9EGNqfAKZDcsI
bka5SmHwe3PkUFlfHtkvnPRJ7TiS/GZFy7NnYewk7c8DvbAOBqwUQmucx78DmZ9uKuDZxw4h8wdx
aE+b9lQNujE1BWA7IG5Aq5Rc9bm7eHQUJxeDR9A3MrtANPbREcdSZPR6o2xuyxvoY+L+83BlelmO
9tcytA2QDouXuQrncq3fq52FBEo3QVYVVHEXUOngYBRBSkWKJVfRIrwgYDZE9kCawttBVXchP5bF
pyvpXDZ82XQS50kljT/6ZD4+F6CbtVg0KnQ7Wi3hTnHULH9sXnA8t0LKK74v0V0UGnpGgCU+vA2m
Jl9TZOy8gCh2XvC4rrEXJ92zaWwZJ+gVkrjFpfzhjuQwSLZHiMY6QilvlVHE7DaPm+oppYp8RLkF
/hCeF+3kpsYVmM9ZChAkm2nCsp01TA3SzEGoX0G7qvnOntptDp1joZWimfB5/7YdKjM4f5MJKJ27
KKqm2CQwnShJIaImkNqBldV+MNcIoIaiCRxLh3d8h9y46MgB734vLhhizpx1ITY/X8Eb38jWxvdz
I53gG5EoHIJMofX8gtn85GTOLYibGgCPAECV6bMIaSCaz24LSQPFncxC5RFYurlqgWK+bhFDj9lP
5nCuEPoyANbYdDAxQpOKFu4A0fiVREqqdsbe8bqMvN7THmrmQkB9j2UWjvuJ7rotLEcV8VLemjJG
bQ2EQk9w22Zl7dO7E4qle9beeiI9N4uFjpwmIEPO8ihRxet9Ts1ioP3WV2Lk+UVSqsZmKZZpk3hr
h3UP/BaQ4ihrLYAHs72ixMnVZP1Wrvxod3kTTSs9H/mR2rav8Ykz+0jtE1co+MUJsV4H7P0NKBaW
OoXWYQ0A+cqP1Eby2sUk5Ezez7XNfUaga4bTKKT/AM2ZPXf82UbjxQovXjSbv8GkMeWHjAfaakAN
8aY3JuFqfeGIAC4BTFvqaaQfvNLeVsnr9loHcAhL6JnmlspPVQZ8ApeZ37vMLiHOKOVIXGJKdkL1
tZauPmPWQal6j7Epq6oRBz23NO9CBhgd6pePObnJcTeUZnV547KwjkiDZDzwJDDz+0xQIs/7Hqcr
LwvCNv/BgTXzZckwX33dN+UsUDGlWz/XcEulQniwbbRjdOOfTPIBHI/1y0NAn+tNEU7fsDdQAacG
ZNZyjadQN/nN+4pG+hAUVFarTDJd3xUAKsSOyPu7+cXofa0Hrn2/4ygsvvnAqwQVHjol+EGZ9A7T
u9+XBGh47WFU75vTNVeKXHs8+O2IOOYSoonr29EInIOZF2/PwqsOubctUqcXmjsYoqy6IrVgJJRv
UbkE6BRz5BUg/KKcKacxaajl633IU0MDWAzs55HV6pykcLlLok16ZzsmrOyFpTscZx+D9lOyvc7m
SsTAgDgKTM0DAyqXBQu5h0K4d3npFHMJNYMK3Vy7xLyyWpEI1ax+p2I0poye8HuvIWf85MJiso9O
uap4vwCxOSW5JraZn+E8jhUj591a3olJvjn8GIYi/1grdgNfHa2B6t0IfUhuB2+rAJEjGiXVDXSH
Jrt7VdXWpAbH201K3PnWfY51hT1JDFu9SzUU4xK4qbYCplKKFeTOfCDiyD1fyXhKH4sYIA6DbRXx
DG7ck8vf+AhdsaePyAdwN86S63YJTEF3YixH556P7ad2WtCpEOYDqho8D88lpRpovyVvx58EcClM
ksWUueuxYMWv3YlSRfy3UrvGIaIKGAhwC+D/5h+phZPcjqCQWTu5VlVmK2ql2Cs63s4Zi2xbq2AN
q6EHy97GA2OhmX4ZczxOD86FT+Ip01krQLbJ8R/FubGJfGJvUL+dGirBX/olZpsHutqX4ReuSrbw
TPlC3YzLtQr7ECmLRbUI41UUZA91JsLR2lqmHgdSIZ6uyfYaqZuF84FntN5I53FaCS5bI1HNxAg9
88BWY9+/NhFKCDRrxNstBNv9U6RzIrn3jfZryn6+0DXDGO/TSpiWsxyQoAl7FDfnlsDwS1ASBHpE
Kkuz6oATmgjcTuZeWABss9KJVSfx2mhQAsMCXFJNPE3oQEHkSOEA3o7Q5SGcgI08HAPevDAhD4bg
SbSSMbLSwhodsx1QN79dO1kaFg3j5u0luI3V4ukrKI62ot8QezH1oIWg8+wRKThDyDCTloFhDsL4
N7oDfXr2e+n1F+RWDpv+FYJoppn6DFAZ9n5ZwmMLfl3mrC9a3XgiX8me11IAUSEAmYQr169tik9f
tiBZaGyynm3aa0QoIjJZlioSpA0WiEd3Qnnb9zNsSRhndc1OPgCVFTCxuDaqekcM+6/cvvHGHmbx
/U3EciMPgZFgBiOy2qRLu2hFzBe79CL5iIYe1X7PasLOFAi1LPn+GkGOI0/ZI8G+cGAz5JG4Jy1v
UOr0vjNAJTUbncDwjPXmcuVeDUjpQ53zDI6q5rhtr0OmqzVX/KXSrFI/PXvWgZ4EqvK9JHEMsrQT
emyoEcYd0dYsSd86bujXLB2OcKQxx1DUggOG+9mq807X8v1VBpUXmoSciAARUPwKI/l75FIkSdaQ
9gRHMGtQbnC+kL95w0ozqLmwtBU1JmiRLNOgrp+LR9GlHYJ6muITbKLOlRpOHfxGF3WojPAj6xhg
eMWTvpVEUuJ5Qo8iOIyg5WsNZkNITRAsWl65V6tk6JBOkB28riesJlu9JR+JqwOcoACuMifZXtEZ
WZ5ngLeYz/W62PMDVnro/YY1kjPkFCspHm4JYc/rGI8dgYCm7V3xR/yLTcRK86VuUVnQSONqzKO4
9mT0hHMKPHbBffjFuatYxhjLB7ubn8A9IqQ7vxrJ18I97Y9UpSitrh8EFdZBjnbIqMpWlYHQLlyI
bEkB199+qZkXPViuCsCwIGdh4iomoNAiig1jX1bpFDiaD4D76JvIYNg5gtPOshW7C/KzwPqUMaB8
gIbg97ltjO+tWmuRDBSd/Z0ZFJ9ST1iUgNkg0UOosza6PGh7P1lYcdjUb/Hy8Ld3TG1dy9UVvBEW
TAMuuwILXlxNfxW6J6By0kv8DzxcqehxKQK2rNRM8zDBXUSPx7r6nlghUA0CekTEQXb1hUp8Ulzi
kq6eKS56Ubeua1pBD8aWwGNsQZoRkLPYLBmkfg8jcAQM7OTSsHN/aYPNAKAihwjE2P1v/ubhls4i
r2j3v5f8eKciQ8rjE41n3wFJfOhTG8lIAg4zZOICrGuhg6tzUgd4Hm7zVqwIQvf7e0MAhl2i4cA5
5SK84UH6HzJ7EagtuOG1GMjn3eZ/XyrjlaGwqnetQHKBHH8UFWytUFiKoAUx+68Hh6YZaSQbiQ91
F6v2/59UaLkMj+hGj4hL6i7Fl3BSAbKM0RsE/zuHL0iJ2cG03sRtEDfhUF96rOdlGDocBPO8KAzd
HuS300Y6ISmSxBpjxVBi3m33pcEWl0h3CQh6VWsOntZIAdu7IHMybJJfjtnDaUhTLUWYEWLFEXeE
1jTTmHBo2nVRAI9HSJB1HFCGxMdgzMjcR5VlI4QIIiI5u8M+x9QhcszOMXfvtaIez9X5qm305vJQ
ynREOQPLKgN3MY4B+girgAiyO3DVRn4Xc0eBChCOHrQNVs58qrXYMYedoWCauYeaZnBNG4pymtnO
NIcysUeyYi5slqJ9XtcRt7ovOxv8z0iO/qfplzhDjnY3LE7es2oaHFYhDYo7CBEEKa/2IEwe2obV
nXI+ug4Tzi/Pp/0DyDFxPxHuySdRAn7JT1oqHj3xPVraRW6GAfVJxN57t7TDg5TNd4Z3l0xeJcLr
mZj34JXh/GaVaquYhNYm/0X9vTVMzohN6JtcLUJM04v4KYDXBpYPSmLBkHINngbz6yHUAQ3rY82u
yMRRp/FQqr8+0GRfnnozyEIvIyvQQK+GzW0Gg6rMQRNSZnbws1PwPlIJcBN/B+m0SbjtvyBDEyfR
St2rbxqxNVuoFo52dYAKSWARwT8NLDFzRgxNUSS+gJU0+wPWU5xJG/3NRvyjUnx6q4TmYWaOy6pA
x1LmQa7jvCSu6rGqfOhMAk0ce34OMrWYBgg5HEfA6wMn0fRmGQX1VMHLwGdlN4c8webGg79Ta3Ed
sYpRn/FD9FEA7k9jVOugJYHboo+LSNm02GcuxJZ3Vu+Cv+hyddR0J190ry/lHb/w8UsgnxrcKPji
nJEYbJDRfXu7hniUfip2OpSUcHSmcBnp+MEqkGzfZFJIKloh3JXtcHZNX2LOvTZka1PmD+1v74Xe
XmglBya04P4ZcPRtzluppqcuk4N6IywpOTdep1nB0Le3S43ucwH34q4NQKozicJ7dSgJJTDCS9Jn
yYQ++sOT3O05NUtn7gpwEufqGbYSokEXQgJ550KevZW1iI3FIchRFH8MG5psQ7HDcknwm0KoWTPl
ORauSa2qG8T4Lzt/z7eackkpTqhsNIOd476d18ug6tF7QCWIxyK6ySo3fBjN5f7m62agkB5kdH6R
GF+PtjMSUEGTOmo+wo/3Pe+deW8zPAzMJEUm3DrAUoy6bWTK+fIojP3Xe57OFASDrGrf7zPFGe2v
jcCHp/Pf8XAvOC7ZiyWw4c0TJMF/MBKrRiyUzsKpXYGFQpJpPIr7HxcRKyPHw4nTiGh4nTuLobQE
2POGPhlmyzqbhrJTcESWosod/OC9TabbECXur5GKaxAUjOCJtV4bVXqbNB4zLywPTJZLA5xsDXex
TMo8mX1ntii5+xWif0XCYCTHwflr5Zi3ag4HH8wBgiHMgJwP0yhaofze2znop9DlV4oT0q/4iMnQ
EmvviYfrhPJAKOeUwqcd3G/LkDLZ2G5HiuNaOJqOScARIDYJ3lkbsmyWrPw80cJDvufAdZJ00CFn
EwCntfduufqaX3EWNkuy7jHwR5BIZDQscy4tX75HlCKkB8QM6ChNjGIgndVjv9KuIHX5ZAK/IMAe
JVrRrJBZhvjtbxTy9lZwBp9NV8v16xBL7oJu6M5gTCXo5je6EjovaK2gkI4VN+DFpSui9FWzsGZl
Nvxm+lHSUto9t8QxGZJ7qiRgOhVQC7txrhy+CM/7K091+mwt9BApVm0EjmHSO8ezYMF/0B1YWv8u
ebc20h07CGkQyjJb9IOfZstllPoZTY2o7H6NfzJEHQP96aLL5+HlkgBbqEvizlzHvhG495lOJvt/
NAucFcj8CijACLI8Ey/YN3BILmyORUBeKFZFpucpd+owd7ZiQVZg3z1l3q5DXOzLdOiF9OyU4tMH
3MHa2Crar05mVVw+cu7XVI55PBApPxT6mpySBNOvGYfY+UVYPtFevDrDIyeU59fE7EBA4SESxyqi
gbMihEpfBgBhNeW2cpzmIBp3WbmPy/J+jW+YCyJZBxLAWlIdaGlCcq3Xkqbzo/Em7+q0kJcl+XDv
bdQbt8S0RWH02+t1LVOjw9fqEloLAhg5nueOzoj6LkTnOUaOihpj/ND2R/4ylaytwn6JLiCCXUhq
j8FFOF07Tg0PGM6ynRNCM8stwS7BBq1vieKwR325nKJkq7OS5uOnn8a9ke6Tg+LOZVBXTi9t92s3
KvKStkpupjl3AUIbrD8fcovUDCkjA5OTY+YaHg0omDH63/Qk0Vpv+DbUuzkjvkVtsuer2NSC4T22
BzCQVpxDPWWxdNJh7Kp61r5+35BwBm1Pj3DJVUV6OF0dYA+c6npBf1Artk6jS0XbUJ+mJSwX0VGm
t6gL35bnRn4iLV+lM4JgFNrNjh6Dh5BDW9COniZUof2B6+hHHVBnT7Tkcwx5BPpKTEqZ4VIix1JV
wpNjFqzfdiDh9diE7ZauU2PZo9GLQr/ZieKURbD73gSVXBEtTsHVX7nVjZj3J5+FHgVO65ObdUYY
DE4/+6r6WGfb1K9b+61LJVosvoxpNoGohPRM0uYbjYAEjUii2uAlk1OE+fDSc237MxBMBbPX6iqb
o1PJ2ZaxDSoaekYxgwm2h/BtQE78A5byUHil6Pg0fE/DKmzDN/CyU/YdgCgjRLbYLkX0jjIhGWLf
NMsI6qd5/4JsCAmz/CeUvYKrVYMC9pso/A6QTcSErKsOy7naC50eHQ3sWaV7eNFLiRHel61huICg
WU0VDjCPUweS5ohmvca4h2wl+KnTyns0LxzC1j4cjjsKTi1WKURQ09BUyVY3wTa8pbwhB8/BrLwh
a1Eg9RIolPmZ9nOZphmFEemf/fMSDm06ZRyKEWKlTklxdb/6YTDIGDe2VaiYqqlIvBj4ZQTBo1zn
3GAuwDSdTjUUeLSx1eMpCltlMjUfEZr8h8Ebc6p8DzUzGlgneowPpoa3g5262MnVJm+e72B23ZZ/
uNo0WKhN+w/gK2djJ/oSVVk6G/LXjLJJgf2xdcO9hhXkBkQ20VEnhr4H+bAWeNHWTc2TYiKMNYy+
5M6A0ieSh+8gHUfn+XxPbIZgZ1Abyrl1tTjNvx4pWTKTBvSvakI51dTP7GFxirJG7y405z+qUqqw
20iunIWiHONYJYP7aAdbwKYZ7YlZJqp/Mk2GnW+nyVHbxYk4X7xcw+HriJgvEg6U0vB2DggU/bqp
RsRKv2CPz0m5UbbaxP+PcBaeDK85t1gjaEIOt/hgLvjoEYUY33jsuOX0CloxhFs1LjTkojXxIPpt
Qfr5xcYbS9y/zidISJD4VQTAol+gQk1RmAMGIhKXmdmBh/O7JHsGotPQEes6iM0PmQ6+nLq8z89F
9J76z+waFKA8ZYUYQD7fVTdyc5DDl5GVWEJ9A0inTgSQJNgsd4wOmB1tHR/ddKF2R3qcvJdYFYJ9
KcX82uJJFAHBQu+DM9iTO8ha9HcUh3WpofmWQSQHdf0llltODB2cATPv7QuH2fDsh8n+3WtZ0QFj
/Xn2ga9wg+ebFL1hoN8N3IPREfluTqLDuSKmPyE702GYk3n19iA3POeQRLSo2U56+C6FAHhKAGTB
oNQFyktpXaBqWMvC3OUaQ/8BtxBBQXbt6VA6kbcxlS7ieDjw17v70Vr4WmzZ0XM/17XfUHWsI9a4
CMyw9ijIVb/YreuP4VFgb2Wa5RplNzw/BHhT++Yl+R9jLSuojwZXANvpGMVsNdHwNIR/B3YNq+J3
nFqyQKP5ulhyJ7wAL3sxm1nI4oKTXIGNvdY5aYgAPGy1IXiYFO2GNTsTUTkDtbobe859NyJH7C3T
/qs7YL71D2qJs8pT6tt1bGEfz4OU4WsCw3/Xlw62VyQg7lEsb9nI2lo8et5Zd4spMtU3W7fPJK5r
6ZXU4/Wac5Skz5jEaLw0CcY3lA+D74XSOSA95TBNnzOagUak+SKjXHd2/G+fu0CpiQvWhd2P9LUM
zU5Uyr3dLkSdhTgVCICFYzk6+mYKrv7pVkAikQpBnkADS6UYa7PPdieG4cCLKrAnEoQd3RBoSjBE
eMK7xlICXNxHspZ/bkcaHvQVB1wasWLJ/C+Ivqt8+jNxZqBoaHjm7evrKS2Sp3xoSGo6j9vqClKn
XXQZeEkDbU/F66AV557iX1oRgZIAac59D4Vj/l042TWJyR1RPiHyEcHIgrR/WCSANMMlqDX0OXWl
ET3zFL5XrjYL12iil0FdMlG9pY5JGPZGwv/vvzD26L1YTPWwUNGRMH2ncP99w4zKNXUD4YT9CxmQ
EosuBnLWf4HKZRN4c/sY091rB2W4q4CHLg8QAlqFz2y4TdM6oLohr1mPXe1np+DS67MLQMA6+mOI
yqGxlBwNJlGvOHbJJcFkTi2xa5WXNQ8GgdwVzenrdg42wXhKzA9LqckXvUDFdfv8gjip6GB+y/tM
wAtZDi6kJSAXXuIMooaLHhmN+fL6CgJGMq9t0nkc8GyDwCYq0TNfxtTmCqhrh5M9lDVjo/8LLMpp
YZUy6RQrjzePha5RWjrDtPC8uUu/LIM83XxOPWa++RMY6908maH0DyM4nNYbezXjXbCtJCqHpIeq
7evaZKYTc/hVG+kMzAkbDnjg3M218rb4nnzLHB0gCyZNI/ulRXqoz1HJiOKLyolI6C512E76iOgs
fwr1UN6Tg/xthQfAGQIlejrMeehAui1o6/ymYEsL3cENFJqon+Gut45Dgvs/V8lxGpDMlHorOL+u
EoCGwlXBKuZY1N31GiFTm95wsN23w3LXup7hKSRxs6WEpc5hIuhGy7s4e64n9qhyvYElu5V1WxWE
l0adMKLX/4JCNiz/nflj+7c9QwApBkquIZsJBeh6b43vazSzRNxIDwH9dhIPB1SqIAZe7o9FsoDu
Q95+zvaRIRi/APeVZwW7O5A6I8vAGidId53Pe+icKsp7ey1aFXUOl40vZkl4BjEX4LtLQcSTzbWW
xyOQ0ELFMJ+VtzQrlaZ4gTY8eF2ULv+ihX+RIgxe5tQ3o7qQHQt1oMLFyfibxbd1lXSjOrcGeWkd
FIA+ZH8nE6GV9Qw+nCWwKfbuYeiufMIMHNPGPB8LfoUtsCLT8DcCJ5Socuj6S9IVswlFW2HP5Ma1
0O0psZ9DCQUOIJTWJ1n4butBe2n70KfLKoQBb1DIri404z6EgkWNh+WVYI/TNgk52ZPZxHRuCVRU
BR16x9HQ5rPdHrn1zKRwKNWv5mbI2Za9ZTknqNAA8SqCZPyW7vOZCnn7bi4D5RD6mim+jodjr6/0
efEyWfMVDDgXPtZh7wdHb1Ex/VHhF+b3dt9qhecJkcL8srIwoD6y2IjJB9Iw5j9n5atPGdSiZb8X
m9Uc6lPs46lZEAfVCibgrOmRLu63vaEn2TegufXR8RTwMjAxoaOOfgDJydbSKr5SfhA1pYVJv3bU
6RX430Nl1Cwc1vnI4VfjZAzeEpHqWRvcj0P6VgTgDVGy0l7FswcpDyK5QF24RBg1JOGCPl1OZWNg
EKKMxyiv8cF1UlApkBPF+lEc5rWRAsnA963biNUURKBkBBEwOK35sSlLrccQexocyiCnDokS4Q/t
LDko3rF+qI52ME0MRK1abFyoH3NxoTMg9i1d/Uw5+WB1WI4lCSTlYupBCZJaNcT/9Hy/70caFEm8
yHQUqbdhTsBujP9yIUWQKuBMf34PUXJxMhAXlZtVWPg96nuMVqbYDgwYqjGcoWpNlMwHn/TDrInC
BTocvBQJuHx6gnMVq8mAFk6UhscyMsfj4ytmidTgT+TuQvPSBjqY5gBBjssuRyRwnGTdShFlSRzs
yXbb7ipiNQrV+wRx4K87PwvGu9j6GrivQdl6+bwwnmSwQoMufqxmFazHFHPW9pt/YgN/gHYOu/HV
bzhjgprlFn/Eq8euKdyBVgLHVRsSczoDMS7jnKMohm88ks2nbZj0chcpoyCbXobXSG6CF4O27F3c
1fCxikSdgOoCj28fSPxLJrPlu/smvMuVcGUaMmyZW56f9u1cOP8HWugYSU1NgbXUHpu9FXwATl2T
B6Xd/PnpxSAG6z1ZvzYWfBmuCeOGjdGmqaOKqDHD82bu45Ixq0+Dvdw9i/PDU9WMomsQoCMUrhtw
f3m9v1jIat8BAePZ3D9RsuG1U2v2Buv2Cqv7mYgE95yPRtKkuP37UTHvrqN6UL8Y1HNJ0FjdRFIb
Dl5rR7efoKuj2MDAoAEhyMMbmMc6Z8dlV0Acbxm4tainMlkJSRvEu7Gn9xsoZ4FkbKu3hdy/XBpk
qDIjSCXS878sA5VPVeRFXlYdZPD2dfxUb9R0Ikjn7BpJeBAsyUDAX0C41g1uT24TXoGtanW+KzPN
YHFbVip2WhuH/jDac1FH/gO2KSarsgje6+vjegPhqruzZ/AyAeEBLbY3KiY3mtFBOwcOvWt+GjZB
P18Y0Kk/8zVQNclUpDGyrBzQPJwn0NWHRUoI36A6BiEl0/jF7rAcTqmqAFKWErr+hogYZVSU19Xr
gC1qCQ0v61GDBf25TEw4eTEndOORzyvn80O5vcWSXV+6BtZ4zNrDynMIxJTsIXF6JA1sBsE7n8Xc
GEgnwI2fKv4ZCcpezCuhsoDIk2hRs2f1b91EDcjMZT1A3m98XfApA6QkwdIUit9cl0m54hUexiL1
Rg6kCpjUjaV8JWm5m1amPw8MvBTzuWaabnz/rbnmexyJuI/9s2mrE2w2Bmk7x/BA5X70+2+k4M9m
9VLSk8jSGCSHhFFJV+1j9sCRIKMDMBLngftV35UNyUvW19C6mHTgLmSmmfgycibuk61KtFxVg6fH
cctNFCukhH0pZQ2OkaZ6GuymN69JRbF5+Hzvo+7DzQ6CgeAXal0TpuoErrRSN4PdCzq7AA++ldzv
CWsNdYLtrPltILAtVAAvblcj0ZfBl3U++VAuF56LDZnOD6dgmez8Q0W9kjDyBGus0WPZRKwRefR0
NudxGjXB3RzTPll1q5ljFcgc0lyzpip/wjGAEVv7ZrWz0J0VhP/1U8gM/o0EKUtaO4UOdQgiwzYZ
74uFZeQak4c6OReoCjaE8v4mTXkDRzBv4vuJawrEkNW8z9pJXsF/GAKmEXf/mz0MKROc8Oi5r1C1
6iyuDnXwNgNrgQFpwBk1T1hYecSNv08GmGAcKs3Cn4qqrMD8Sin9oNCvgnPb0aaJzcxAqas6X7aq
ln3z2Iw5y+DH87p55lsMm3VtQqW4nARKJSZDvyG47l+LEGye2ZZW/0vNPHGV0+eyzwfDKP6S0I+Y
XaZwFet4lAlCS9X52XO1vAVkgzDl4Nq8Wi2EsyBkdbxMk5izazefuJijmFPaQ/9pHHMreomAW5n0
U9h3kaQpIrusDB6iZ5li751sXvd0NJ033PBzmIK2CWeB2Ofr7+t5jWXu+RDCzZvqgYTl3k/6WxbX
mVNaTjSFrU+oElGjYJa8CxhtSkLvv1DUVKnH5Ja1VaLT1GckyBZAE3H8Py5rajpZ4hsy9YzZHGXu
FNb93liMyaKkd7wjZegTXLD//Gp6w6DyJIwMulIDLer41NDRh5npjvBYTfRFGyjiVBo2c32d18H3
xaAGd3CC34OGq7N1TN3ZQaJEyzrDw4/DXAcpVxKpGXjzBqAeIA3qIxyA9ywaoPqQv8CogMh5uBGK
irUgiNx0ghEpt9vEVVBA030Yc6r7/vtFQ2M/DKmvrpJAW9IAEOA9bjjMha6zqiMdFid2F8P0jzqs
cPtd8qOj7vlvNKnAf9FOW4GDjSUa35KjeYPQ1yinQHnRqS/JC/wlpKusrDYMuhil/WskFaweQ/Wk
Rz6hCv3OntG/yIW9cL6DyvwA/eRR6rgOsl5foK924Qoa61cykyaE0x0qgeV/b3tcv+tAV3VLg7d6
4ZBVcG7WI9hSxnmnbDZITvOC5EwIbjPDS2b6sWpVOV4LAMBzLnoOhhKNCyLmE1W9XSjjbhOJHzzV
u84KpSQHcJmSWEYqCH1hJUs11BNU/88emNDjI4Aoc1XI7QBuFMEIyRgTc8TAykhytIZKH76H2jjS
PZrMqpOEFJYOewEpdl9DwytHZyDmnQVwXo8gLHsRluhV9ZocYNDX+b6fnryqwFbzgWPHRMRHm5KN
StLVbS45O0vx3dFdSDKekaxarCwZvdoQV/eNlEt7fdpYO7YZ9p0eneMz8SVUqwfEy45J3HrsMUGR
XY8lj/+dMP55nRrtEuGJXJQKH6iM1+U7ADuFtd7oEGeZ4wLBZIJIZJzs8tvbVixKgEv2CwxLqWw0
qZ0dkhTKhHXwKrIt19vgaP+Hf5tVUL95SXPHs3K1WrnPpX175PS78oJtB/SlDf3Wu47LhlDvCXee
RChXfTKEXAbFBboJiIW6/diV9mtf0V8OkdKnjhep6C488KEg7SsAaqzJbtDV2iMQ7ITxvUMghJUZ
rCDoeu1SYyDOPiD/bKbh5UOUV0A3rybN2WCaU6umV/dkNvbDKpKE09ogAtXgW/FdDoitPjDsoemz
TDf1i7aoqTanm1c88du2IWfgW9i55lOB1zpPsG4q8vnhP9zBYKZ/T5d35mVehrYW4C+HAXmWTBVs
nypaJuHHbdvCbbpY8eJs5NiGmGB0OcT4BCvtrpDWWu6IsytposudCEPISikOKwNJwSF5X7E9M40V
0uvFt5u2LRSF2xYuVPz3u4My0/j1mPXeu9OS3mzyTPYGZNUVB13JZcPYIgRnFeD2MrhG0BedGaHl
Dh/iLW9B9ljibVOlO/+ac3jveGj3HCjr8Zlx7dWc5/mJns3Ib+28M6i7kxvNN3U2ok5D5zfVpnOn
PzWRZfu8KvZ9cHYE85H2gvriYPggHmU1y7PtFj7uKC8gtbx45JKGMzSCOgLgcy+qzieSnNQsoZxN
Q5eWj5PcuDzJnUzPzBR9W9L3p7uLTDdGEKAaBvg7wpUe1rV+Pvyhkwu1w2ieUUrQBDNsXadShni7
TV2o7ovefkaEjcltMk+3SBVyiOp8icXrFjETshaWJrGxAYS8Bs09l4RjmPWth2iv3mhoh8D3MQ0U
GNutOQNoCbIFUFiCh1i6lbcrN45RN0VZ4d05VFdAzTvw0dh3W1ouysQye19cjqGEQUDVLTaF40Bs
HfbjeNXB+SMjrQUKnaofB65LcALUOL01L0C76gOI0Bt4KY7ywET5Mmzb/N1bpCXhnlE47Zqev/Dp
IH34lyWxTHVWhHh3lWW/eN3I1P5oidcDexAai3UPcOuvVx0lcFTImPbG2KLaeUkluKEFCAJJtOtf
2NZr0JbNyVtAfRfNYKdB/gOzP0h8B4Q0H1fEF1SAyr9nY/QucrE9argKuZKwQKB8Gk8u8ysuxRUJ
kV8wQs82aJljBoGRCRFFd458lqpmXvaZuvSFK9lHYDG4g2iiZIPGSQBKR2RZSE6UEmmUD8DWJ+r3
aibxZSHJ5sIpGD4CfX3AdfJ2SDkrU3FoOwRFwOVvn+PYJOvACLeqQYEENVyOAKyeiaYCGGtiiVf7
C2dTVdwVcL/Bvb4/+AdC4w/Krtu8w/+plhVdJlymWunuUC/N96QACklFDcrigaEgA4VXr4FnNtVZ
Hhj6x+wA9S9pu4c61lE/Mnm3d4ScyoHxjsJeLDA6TiVicKE4Vadq4HtA8TTVQdJORex6dlR4PsMk
mxEd5VPmVvhBMitHGdVjUMTkkfVj5HVgd2rsouXTTahHZzmQucuJ/8yoNwMZDE5cH4mTRRiANMFv
9AjjDK3bzic7IvCjxx81UumITA+ScMNHT9zC7M3JLGiAim9fOBCCPzt2gWb90IsLVs4IywP1PZAa
+e1qR3FloSIuxwl2LRZkVFPVKmMMbWMVt23IYTH5ECSnnzmYHjEw5GGtGv1kCm029FnStncGc5k6
oJ9WkVziafs8jtDulV8ejErd0S6/YVe7D2zCCjP+TlvPj6ziGQ/sOKz1hBrQrlsF+hy00rwOc+Oi
vtIm7C5CM06cQOkt+Z1kzovcF4Sm0GFYNoAzBSgQyMYQWccYuJK5lYgGVW0dZjlwzBZuvonkoCMt
ysc6xLfT/XbYmkQaIyJhHqelBjQt6cgX2Vn7/MefZ3alsIY2G39FBFMrxZNlmrdL1En2ZKi1LPau
jiaqYtlulKpYqQkxTohdheZPFj9wpbyDxOaDNYStyXDEJccZra0ztjw/XTqgZq6yMeMrnuIYTU7T
JcFQqg2s559NK5osh+vMMAdo285DuSb+EMhHFnOsRx0d01h3eD305iOQq0nc6SBM1mKWxI7OPu3e
AlvKEk2DhmZwhYt11t5TDHJavZ/u9wfHv/S3JcB8NRY/roFug26lIWEGRmZtd8VMU79l8A+ERo7/
6Jj1d8Vs1NRIWU9bSMitVedGAu8wQbgOp+kGdTgIvSu7dGxH3ss8O8aKRcUcsN8WnySfLqchJ3+s
m7xC8E9JtXTyU58QZXZdYL5K1dUEF/8PNifT+ySySb+HG6I56yvdVl5M0txXRhoyNLuVjMKbU6BO
10HIrs1CgzAeHrbpt28SJNMs/X/O8TgytrL8xAptj9SS7WtVckfC3ROkoW3Uhmidgp21hOnleiox
V6AHdZ0BU1H4/fOR5c+pLiXgJ53xEbrvj9T/rj1RkbEndGMKziAmhpbmuodDOURrtMvx4TD+lrwA
seFxQGAYTTfpBU0nVV2qbJTSO3V3ba7p21DDi15PR3n7qyxPXbiKmcgfyO3U7Kin9UuFo+oIWn0w
1LZfv6SheoIbmSWxXfR5KsBhCjyplA/T6m5ARaLWIa+TaEmoh5lBeNEYsUD6Hm3z4j6aa7fVUUPQ
dxb8BekKo3YLQueZKyTp6wKOUBW73H8ONhpqy4ussuNQg5bt3Ojq8qlOVnlI1eotyyphCfyNRHN+
s/LjfkMyse4ZCmfl5Uj8v0qeSgc/aR6rLK85a28TuTvJmrSuU6zp3SXiHDuyoIuGyL/leBpvpMf5
AJhOnRnrMUXenYbTLfR1UidcuLpAuD8JSmIb4ofO0t9thymDDTfyZApJRP+vK7oVlase8xp6lMSc
q+FoXbQtvRYaVtfNNsjJdL9FfzQfSCmZEOOpDzpFWSL8d2mmMYQDqptZLMnC5WxNLe68C5CQgMY2
e9BinsOWCu/jPBJEknTnpfVkC5YMalIoMYUdHn7Hcly0CX5RBBHZruCEE1AgissHNxdrt+uRDukC
s2Xo5d7CQ8r+szmhiq3aY9QUb0vVFd6yQld4KBfbBEki6NBvMOtaEIX/95/wu7O7eh7mMWa2bu+d
BSh3DabUf7ePZOiSTMcgl4Lnv2o1U8WRqQz4mFrHCeZcknksGUcKFVqHM/JW0N6MvaevoaiO1oLx
F+kLI6hsOMqQ29G7INJPsDXKduek/zNXW0gmSnk1oK6gq+l/lAGD5h1EhGgcKprD2AKHF7QUgKwU
bxRrpAs/7L/rqVfwIwZfpLmkLn5xPOvLVeNrVmeWH+25kppTwFsC9fa04lQLA+2mwLCjiOcYt3Y5
j5TZpXGJyONskaa9hXVdLqMXqHigWqe+Md6sjOjyy2P495AT2mTpLmMp1/d5x8A/2twfbuRd5/gd
hzPY0IvlpXDKNDXxZG47CA9VAVal0FUaC+LOhW1R4aIsXHA5xb+c0j+EIqipRFzLWfyABkDV+oo8
bB+JPQSVJoh3BxzImiPL3lk2bUBm2ZqqPxnhbGqsqkdM4gLYfn2SJfmE7hyR3hJkB0OJyzBFjBtM
486gGKAIiooqIFKamlW45e9DRzuckmaX1QOyQZg09awTDf+Awi3GPiuC8DgVoiCy5hElquChS+Zw
CuiT6V8ieMS3dPTvVBihwKnabeIUVggAKYPvkI5vlpHQ5FvKMiIFhWldPE5rVqJnd6He4f65F2cE
RjJkcj1QsDUOevDZHqQ/J0cmQwXfmlh3mylRtaSYXMERF04BlC5GQPV6SxQZu2N21kgl4+X2WZYo
Hes4/f2dcAX90I8/dJHYrUPIZqVALiellNRa2P0EVannllyHwI2NGKq96F9ri/O8uFo4hEoLH6Ft
YqfHhoV+Jsi7TPfNYm7KWEtczGcZXub4tAsk/rSirCLq79QFu6BXLsbfbbpF15MZ7EHfvtJ/NVnH
Twd6lbZu0Rk+1Pf/rCbuBeIG0frnp3B0CWc1hbbsaamGgYMsZzA6NeaHWf2w76Rscw43NziEBarP
gnXaes5ppmiHwHGDGZS7HLc4hGHQW42vXKDfAhCJ0MM3ZGGLxe94l7MY/PbKGmUW694ZySOFwzyO
fH1RrzddPLdUK3I3nUzE9CS54QIZDdE08Hcbao9UHhTFKtq4ByVNcONQfUiOX4ujws+TjYaQO8YM
+k6GdPH05TjzMtJRb09JcuaIDkkDeXE/xs6+6IXsraI+IbsKlKcf3zUqPR64AMYuZ26XvZ7WBHuH
mNzBi8oesz9e2DLGrQjFNHFwV7NJYdrvbGXg81AGU3nZsewFvsoVjC5dzEiWMCTMW1bSVfHuAj5o
Jg9wO8yMcGGlZjc0QFK1RWMyF2ychcOEdxlxVh+NYilg/CUyF/haWlK9AmBLED272VJHqqJHQ4q5
8ElGvQ+Os65QzyyzDlnbNG1jNr7GIS/RPxs48zpEh22sxktXUJVtvWMNmAMODOEJjl0pogXoCBzc
ZJkSNB1FGHi6pHytvZqBBSpTogIu5d5LLEowdI3rQfxh/H94n7Rr4yLJq7jPjFgSRPdtIbRO3grQ
xWcs+YmET80JRoeWBHzg5AWnxckQYqhBFr4FdFNuEa/DIJtZzt8ZyEBCfDqe1+ag3QJqDV/CiFUq
UqjgP2DxquIuKmW0YKxokLPBTR8ugP5nzLKyNLtciiEuOtBIIasXMp0DIEaFsCHFFAXx+uMuEJgz
7+Th8Qlt/HNGJdcYOInVnkKxyt8DQ77274zgWNOoTKaDD3fUSJLt3Y0NSaR4sTxIahlCSC7L2jtZ
QLX3nArLfYvF2KmYcGaL9tV/JDSmPIzE9RDxShBtLZF4oSEU9Y3kBn3LIGhL9XtXMj/SH6UU/rUH
adQaG8Bc33hOe9OxOkrso64GF9Ul0k8nrlsB7MSq6KKsx62oFrdWugjcXgeCH1q+57nSMNic1u1v
7Qvf36jeWkk4bf20uAMU1itXGUL6KVv9FRJHQAMaIx+svba9gPtQHnkfmw/joA9vbarTzQCRt0xm
KaPMIEoh+2hjDwT1tmmmRIxNKS8fm7UXmxJc01CUH01y4wjHEeSHfQtRcvtC3TwqJF6Zak+nAKmD
Gw+SOUbE4ZhwHpbb1GuZ6ve6lMFDrQpShBWrKgxgScJvTGmJqGC6Si1vNWNpNzEKNOVxzoXVloCw
tTPTPQGp1fYIHs3s5RzKkj/z2pl25Xrnh7uS1OeCHzOwJfVTg5ZEcDvNoIjzJmGTHCiU8dd4qYjR
AH+9VKOKlys3Owq1xLvx+H8mBPbHGZ1hbK/EUz2KJX1Ljt8PtMqveHj0QiVmd+33i5N5BsVen7hM
2fpqvaSJI30lyX2UVWHYlH5eAWjRatb5u2fXT4DExiteuKuw8Dmoii7wzlcjM1nT1WMLGOYeDUWb
zTEUiVKDJMu80/rElZAiUtWceiw921oHaa7kFkWxZ9xSdGYfbWCQ0er/aUn+KMBrCaOrt7Oh/3tQ
HUEk5q8/aH45BH6CIcj3zw1bYqwOBy6HLqb11j5I9RfkNFMAYnWq/CYFDUNnv1E/Xe+xpoup/aYl
Ci5QXcg65levH6Xh4K8i4Z8vOAuGoVq0l4OU3zz24NVTbi7eJqlcLm3AXHdjEVLJnpcgzz3CUQ11
uHpcTUw6dr4HUpQew02IHIc2Ggf9fmwcEAUQgaoBjhjWzjb/VPDdd5LnYXsJfCFQku8xOS9w+KKl
bb9+hBgmZw71ZKrQZAlfLR7NXzKE3jGuJndIR6Na+03JGLOhd4KCrwA9VnKC/EQ1dwR0GmgoBVv/
SfwnkhaNMlCBmTvfizFfTDX/oYpWDxWqjpLN5OhrF4iW3V0AgygCDDc06TPHN8QnD/Lzz8iVcGV0
aRMmVpDhDmmAY6hNwXVVHtt0sSN1/dGrf5BaS5oD9M+YHDx8f7fU0pAmH4mw7olM0ixzVxXFFA0C
ygOTrhfVG313y9RMlkT/sj3Cl1gSU97G9y6y6jFzcQ9WXZ/Xbj+JB28HPw/xxLR6TvhofcCfM1/N
XORQZ5cOSKppH3iQwBGIUSEA/uhLEqNj/uKO1jXVIXrjv33cwb1UqkmjrF224GRxHXeoU85EZd/e
w0Aae49yALBvJQVoZejQx/87jBThKPVWbMrjoJhq7btXo2KRngQaJ0tsUKiwa9OQOJiJfi9dFCAr
rnobeG16vo3zbKl+y6z29bjZhC9wnEsn614FOlmVWCt7TMA0JcSuVAYtsyehbXdzM6prjNr/CTgt
b15lnCUjBs+dIcYEeWPF6uW9tTlStwpaohzK12XseLvVmEc7Ou4NfMhG0sUO1ogiL63jdKQWXr7M
yiFwTuWZLQN2+sXpgVIglI7UQxsO9Vyo7sjGOI4oHkrNLELio05G1rXxpR6HwwXAlXPW4R++trTJ
OQlCjM9u9s8ZaiHZzPL+N5XXU+CDtUdjVbTbs0V/xUlb4WhNIbaL5tsnRUZZLsjtr1FYIowYwEI8
v3oCv47Y9qoMqg+kYDYcS3MOgMBk3nkjTaad62jNW8f/5OpiLRqD6XHLXb5VShT6sL0b7SGlKVX+
r9VhiAHH2zPDiQZAWKDeCcD4Lm4PNVzDg7Nzzn2ujvvgf2sVp0X+QxjOAZ1ifUNOODz3ljytPsaC
3bzMQ+uL+HK/fURCKRsMu1Z18GfR5eXvDYrrYkvQMbt9K/i4+NRbzeYO+2gfCB2jibVthHX9Ot43
at3S2+Vse7lB480+xvusjEF8YHw98M2D1FCMYDKOhBjfpfynypg5VqYLy0mI/Vs0R8jH0y2NznIY
x73OIvMIsDySmyT4uHEfwFdIWH6xKYUOKkqVurNc1RjybubeGqmNGEvApkc3mivqU2dZ4bKa43hl
EGylh9jskdErsgh/Rk3lF2qjZYOPP/rPU1u6CJUK1MaEYL9lJSTP2YvlqZp6T68bP9n9XOqwJQOZ
b1eYpNImguKWGnJmIm2U9JtvMM/K85KyEnK+cChHbiUiEmKlUQJXgCWbsRF6DvDLDoKmCz1PP3HO
tncfxsXazKRQMonlYZis+qzvuoy6qjsgNKWNfoRXWt2ueMnJgD3kRYByYdDhfPJJB5JgBKYBQxfh
gT2getGVZRka2SPWdQYT2b1z1ZpyUHV+7dUxg/hNHKDWvCrfVF2BNiiX7ZBrt7Tez09wsgNRJqH4
+2QFpIJPdkd+YfRajBfM/ORPE1i/OVtwb3t4A4ttbZISZbUzI8Lvpr3W66Sum3qeQaUx7Ax4L6e5
grLfEeIqQovB9TEV94M59Loh+pLhUGEoVS2isbqaYcbvS+GbxXNuOJ17JqHxl3uGMHRttBY2zx6M
ANXxdMAGeeSNGVZxolt6Wyx3FAvIfrHAwa6AP8JCFXVW5ouuQSHMAufhhStYOol8GoyTbJfqrIlb
i7R8/BkkXal3kfu0dEVnE7VYbNzyvuurOaaWpBj5X1tSYnaNiMskVG/P/6qomnwLMclU9ZVTacXs
ul3JBq/712tW+E04wqZfhyvgyfmcm/o8GnHNkuO/3AzSSzDdWadN0Cuv91iYtjyxa1RNbnTFDrC0
d6deZtbDqDggKDBTlcbtbwStMuE+2pZuUr6RT5vmyhpNAsegZsZ5nNiFZDA6gNbe3ht6SlKkZRHR
qhBVe0kJNoW6as0Sl6S+xidhw1Gsc9ro8KdnPpUwc+9+0OJvAI9QScZUedrgi+l0FYxxqqPWRQ69
eTY90m9Y5oGIv/5IMyD4gNsmaXn0DYgY4cSiAS8456x9fCwMzHUUBq6I7BQPGOtOkre/mvGCqwU6
4LuPNmUDEM3ROaud/J+LlJhM64Yla9Nv0pcRveJkS8dFyuNfviNBXHFz7S/OhmZFK4ipSFTTlLUo
TQ9UCLsLjX9jLUQKiuJtqAyIKa5agf9MSFf6fDoF23sd4e3zByc5D/ieZx5HJPvXPUC2i1zon2/u
ux6QLhnfRBIOVwMVZ5tBg9noyxcYhtf4mbz8MSc+QUpP3Scu5Ge/62XnD9A5zB9UDlJWYWteVyFr
+gFZ+5JkSpVsgWYXUYKzlmPzyLGNDdsNqeGdndwDoLSJPhdQ5B0W2xXi9GQxGPj8WqCKjNyhlKqn
4m0QdNO+1ykO4w028DP63kiIXEQPK0e/MRGED1I/Is0iAMsDLpF7lCs9iHB6cBUg8IEmO61JfqZm
13XMskxOgHQ5q+HU3xewOvfAtrVK6iCsjuQmH8EdjlE2AJjjW1O7Du2LNOdvsy92fdQG37sKBmFL
s2nNZNVGeAmzuGaMbULJSX4JmDJVlzOFHpq4jd8GUPMACOLS9QJ26xIRTLK+tDixbAoWu21XZY9l
yj3aTGci6eBnT58TPBWBLLP+nBIkkmeAH8OzPcl/dPFBwBAapbJoc3Z8SNqXSTWBZlUkLnnjumJT
ySQoWlWWFDN5dKRA9+cLu1vqhb+/stIrn6RqLX/8EGb7CfrPNLsZuIZVgBZvWk6wpjX9VDIls6ao
ZpeiU0UOPUWn6oueTo6vWG1U9fdh1xToMsIQZwLGl08It6Pr/GwF6mmcFau81XoMTRZCB47Bqycz
kQPu1EaeNQw+lLTvnre0bJ2vGTlgskw39GkcXwQxERomSuRu9kQVbwKiLXdCcMCrYwOPBd8s5U5f
NU5OZ0po/rZ2tu/TC4HYMn6qn0RzBCzLEXH/YB4H2nbEZ/WcitCOFYLLkcwvojmWZ3VzsziZMNfB
LwY5H+ujvtTBzT2Arx3f90k4x8cYkkLxKgPrrc4opKxaPU/a2fLmNsx+sNTLq92bLWohR+nu37ZS
siO6Hw2HS1OVSyZKBuM7tYOkj/y9KO/L+fbObpQsGTczJ/1sScY+o65NSOgXLuzmP7BiQZAsmAH1
OdYD45RqoFgVgmyKuF0KvnyqaYCdkL1l3fBPG4+lWNBvl27w/p5slMwTyfeNvXnKB7XQ/UPh1IHZ
7fseGmRSIMDETNHBHk+0JGypjYqXdWxF5D/rAXlp4e5EXWAuR+Q36FcL4seQIzdRq0FzG5pSz9tb
xKqhCeX9jS0OxNIhxi2o44vpwo7zYeP5W7UWSKSRy/M8bhLPWBsvwE3t9jXLxL7kj6zwaJUMdTej
Y2xXRakdZLgrU0VdoXi+AbHYUf7NAbx7HNAD3o5HZc08wdXcFot48I78/cfJ08pEftDaZQky+t7h
GKTYYCdw0rQirorsAep3pAqqiuoaqQF1KhoEhEMN3R+KB52Gf+yG5I2fqvgiJYOhkzDyDQI4BD1W
SLEfbol65U1/sondmcKSAFBOPWllxtlIRAI0+AjYijbWqjdiUPlXJEfEnxVoRq07QRqJGyKTzMPK
3cSbZJSiVgLdwMeV4mrmSy90OaKq4t+I7pyiDVB3aB2OcxfDJy4Vqv/lu7kSQVboh+WSZhxkHa9n
hKNZeP0kmdaP0h1Q6SZwpJaCc37feRsyKx5cwAadZCO/3IxXt91LdW70nQywEJ1WzHxg9eeCL97t
NjKGFjNmxCVea2prm88Pn5Lndtaoq9kYv3QGhUfgEmQ8B9ONIWupl925SgZtgns4PUvjbYoBnZdh
kcr+RnmICVz1VzNNi7LSWvFqmSZ0K6Hu38KFX2hC3V1VBSt/kSLztWo4JGmUHrrPUUt0eA5PWasr
GM2UIhCpzQpe8VmFAMDYzj9z70djuMqSLBkbzxuj41eMHHXs1zVbwOVJ+sDN8FFgIUo2wA2zXcsv
cD+EIIhkSowZN5KpOu5NszAG3q/5GSM8DC7IH6+d81+ZmyfNx+HZIWfy3n3QtQzRABx0Dnx1ZdxZ
Tcy408VHsN19emquwQCiDaZuydhS+ofaTfIxWH1Md9OaiJjslnqDcKAjX0hUlHbhgGm0ovLM4yZC
o25sLD1YsqfTpbkPrrjxiDf0W72AaKkJwKdRk9TRMxnPCgMKznfG5/Mix9wrtIeuWZ3zq3wnLN/1
sjAMhfLwEiq1T0Uz8jftbaVOG3SbuPuMdT7dysgzb+P6xcoN3M3HGdpYoA4clhqnOeX9LX/8luEq
8+8/GYEmofyJwBuMAclvJArZom7gmlALTWpSLNigNsRQX2i6KqRUo2LdgWvZtaCsYTxmJclFViXf
00UFnqnAjzMcDFZl6YzxCckiTMmGzcGt43SM+7jiIQdnc8ty3+N5B2tDfS+5zWK0x8ppXQzEiIE6
Bzj97FRCC6OZEDxO827AmZt7M0Ofvbb8uGftSBV9IhZ2U6m5hORvvhVTqWXXkf50pKxJsCfw1BGv
buEHVKYT0T6eQJZ+jwi51nNdjFUWO79aYGlufF44z9mn8F5y31DzDe2HqyHeHBvIsjsxewQs5sUf
KRQx3pabohgpIh3z625OpY27uUAfFVJVRSNI4RLaad/YG7U7v8xb+QOUfpwbzTfiwbhcAv2FrNzI
+27akv6xkMveBv9UhGMs2ppB7u4omqBkUnEJaHk7pZE8o1OogFBdMNDcYs6I4IqhVlKjRav+5ni7
/swm6V367loA6I8q561IVyclxRppfI2mrxlW+OGqodjf+0QxHpwhIQcAIk+isSsvx9UiYyrDMiog
bA7hsq6UV3NI5I5mIwfVzudKw9M9XIjRpLWCgvmfY7F/rKQhUZn43LS46GHJAMb833GMSUDvHVkk
SzoM6/VN8Pj+PbPwjvWExuEtMoIAJ+GZo+Zg3D3SgST48lL7Pg+82aS/mXZh6VaLwKcjt37MRSqd
bv8Fq12hGaaryk7cpYWhjwPx53/3flcEJGrylFEPxVuetz0MPrm8nCTxl5v9HnryyDjKgsU7aZo8
f92nFIuWFVjj36XAexni1r2npeEwVWNgjTcDuiT6ygI7fo8hQ16GvLnMlB6aVhJiSsEPOmd3C6U0
yXvEA+AUt9eagGk8LlLlr0pZ+hG3mSUcf3CURWqUoBn12bRJ3n9eWTgSIZ3r7oV5JgDES260vXVz
alWqWtMAhNEHcrXrjFVRiVnBIn3TrsP3XYSX2b2RF5pbw3HAwbCjpQmml0tfRPP3bJFYJhyzVaCl
WLfsRq//QzymMj0yy0ws5Aw9OyHwMgJPgwbPr0bwInuXSyIN1IAoPF/TQ8Ns0tUgnII9vTBe9YM3
Zka1st80nHkzGvUqHxC8kpVN/Swb4MBYZVh5PBaIZVmk2hOnoFFaINNmInSCnG3JHBspImvkbD0w
Yr0dqpVFQo3vEIC6X4baux2gOxiYDRnsYV0eXJbZnR9DGRSVzTx4YXbxsLP6GWpen38C1xWqs8tT
/97sYEIso2T8doTtkrXHoJnSCdmPZH0mZrpga51FDKDPoOC+ottkFTnng0l2ab4UnHuSBuO1QP2C
BJv6y0nfGnrkONYzZpdNUeWZQ4nFmfjskBZEzhIP/B2bLPXa2owgFXwW2GS4BTRyAV9BZ9qs9BKn
WeKEKnUY6zAKFlU0mRSg0u/0ZTwy1hN412vXWLmtjky55HM27bFNXHEqyJ9yAP3EpQew+Aas/ugV
/qaRvJa4J3Dy/HX+Capz95JiyGRnEImj828WJSjEybIedutXOSUC6ma0z4vjq0FQLVLUUiAKdFDn
95MSjQejmRTTJP/ITUYtLfh/BR60ZoHeYQY6m2CCI3dU4OfjGkRsSnQw+it3q3QQd4LH+Ic4brty
uQmVKa6UJXnVu4XK++tKmYAyTtCGDacPwiEbVh2H+PpuMSS6N7p88DknW760JvDeYkuYdPt3wuCa
ZtQL9BtcwOBaQRm5w85DShMlon28LNbq2gIRmDQlf8eJ/HWy/rllfV8EnUnw1NU+IdR09rvc+lIO
S03OF/MyNOUv3HvGFEdzirkQhvhmgGSdbzamkxzxp0VVT33K0hVf1j1H1l+KYbjFrSpW4Oevp6RV
5snorkLkXyjjmpE6M+c1f6eI8gwjYBmofTzVYPtnRQaioHhXG2SzqtX6mSX0bZove44SUujaDs5j
itSTN8hthL9venVUI3Ig6g8PwhXTxquHkg8hryAHUK6VlKjwJoKxB9YkNkaxLLvkFpfan8Mfz3LM
nq2zhNEnqoglb4+Jpcd3xZl8/GBmeZoZIgcRCwRaRLz+j7/NP0ulYAU0BM3uRwAlnpKz+nztQ6pR
uPDI/L3ZrkfaRiokf7JnUqf8pe80g3HCwoWqiq8kBXFYUcmnB92rFqrJNIBrtaX1JTJGNr6wOAgl
99BrAuyQ8hISlpTWlhXfdSEbA99tYOAZCE0RZKrtv4X7AK1E91c7PH0iB7e1gQwhTt+BoLd60TE4
Om32vPMxnEZmodwuhRLQOOx7zfPl9jPsTX0i/tjjqIG8Tqttd4t0VildzmkZZbWtkp9RS3bWoqZ2
VL2rK1WJkH8VecoTWr6TLUtNntvvqV3qNlwwW7nZRSb2oY4eV12hgPK+Pc+QJbZM/L9Hqqnv3tJg
JVL5QdmZXVf9Erf0CveoWTcZfmo2Z23uOFJkWkeOnkdrDclRrNevj8DDZMkpLnTsrN/GCg4WgOHS
uDzFz9to8ggfHMa2cmVEKqmNEtbo8hlNDcaJknlUxXiVkISGnflkcsDvc+YxABhFLDFwCg/hIRRA
TM/pAkA5DCJrkkxQstzed1VTnTNi+aH6N34suoc9cFf8BIRQcn23DGHH2nt+NUzCG+vNjH1sQ3eY
47CS7PPQjJWr3Hi7DWsHPemEpJ8OjtJa0gcqXfirbXxhG7KWir6VaUQrBt751rOLhBY08eHGYWZP
VyoYJS083zGNn67cYTlL2s4HHhFyxSiW8C8fq12ls9+JyjJa3NR0VpQQT62WRC/3G5drRF83cS8a
naO2nIQWoWRMQU8dGwykEdxV+Bb2X/k+HnFCa3mkTggi5kdMPPKom8a8zsN6fFzQ4Hne1eDjwnr8
Pwp0kD8X2FXPBITJWp7PcPOEtPDlEcFyaCTA+gqjg2SpckeRqgvVzww9+Yk/AJMpozs80N0nE8E1
JxmHyRY6p1sa2VYeMHS8mXtUkuu7lMz/e+TR3e4ZQAF1uKb7+DTVmYaCIksDnH9ERZiHG+aFXmHw
G360iamIjXrfYN2uK+VPhmQSrZ4p748PgTtQ5aoaBmelBsQikD+X+/fAa5Dt1dNIHg23+c7rweNx
EuxmAl9QOuKex1Bn2uvTzcnfvYi00ivPMBr6NcS8ZRXOloqZZq7InZZwMxyjkiJa+4d8m+tSmBDO
hqtMGle94wI4nIyaOOgLPM39H/wSSjquux5LZD704jUbO0B7/r4r20IVnEGrbHfBahn/GX+/RceG
TpGlYLIjWU/5+5lfuhsIepCQjpAUVTM/RY7uXRg91EuhRyi3QNLPkraIsfSVNr4aMrdXTACaoYzi
XsGwGqO/m5k8L0WM3sVEXbTy8DUwfffuN9eOUMUY6ch+onIKeMVd+bnNrEZEecmglqktIvaPRO46
xJnGR8YXKov6QBbreBz082bW9t7/gGKyo6SUYD0yK1uU0D+hhrI9XFcR9G1YhWuu1YE1aIk1Vlgi
4zMErKX3c2FtOK62/ugLakQt9++F67SsyXrIiwXiu0Tz6qP1Yo1L7g3ki8Q6KYsA3n3qMhzOqw1F
4JqPCQVcWDKytlBxfi4fHeXPRsYM3sjvqSDPcHu8UoN18RCi6zWA+k/FvZ3Agu9M03wbv+iXYzgq
ZB8E6Ph+fF/nIf42yLUZrreKJHOeYwEbElmP3Hn1zwGW4pafy1BLP+lxbEmzkkgSJJpsd/cbpsPK
eGk+quzJAgTOgfK19D5dRG0VrEzgGlVRmv0bd/HSMsS+moIYfoRRV7jSaN02I7q3zsyosR2GhtzN
9D8nJWF6384uhPHBcALDdLxlG4Y1H0FeQVCcOPW/bW+BfWQO0Sq9X3s16OcDpVvOIf9MaLd81scS
WexebqjJgZrJao4IU8mzdHYoM17gqQQEBYUhMfHtPqOmhtSB51qjAWIIJzb/yykzrA81/ypnP6OI
UBaq+6Ku1+LiDwCaWkmbRNNVdWoCbKobmIUq72R8+3BWl6LMFVCI9dp1Utzz3MG5dfSJQmFveFd3
XIvkLiRyT/RfY3Em227tTpeqLcRi3imlo+S57qfBPvzRqYN0EK7skrwqFgWQ4/wDIjyHum/BrVWi
9nb1zZhu+V0EO39fDK0HehidlL2WaS8FxNkvQ5EMYB+y2cWWmsF1Kj/gaY5E9vycDfJg/r5+s//W
xarpNVqBPBsC5Z2CaZMj9EOM08UM4/VKGsBWqgN2HIAwo9F1/EBbNYpKhR6sELVaiVlsybA8cZS0
8XwyMrLLOVV/ZtT7rzU9JZGvkS08vVuCjSpHTMHCTUG7oZlJxt45BtB9I+J439gqKRA8lcx3qe/j
KB457ju29D8zTKDH7YKvzI2powy0PETzp9lQW/bblye0WkvekUx6I9Gd5DXVBQ5A2LL6h/RUxKiM
qVQnjJmRaVE6rSoUQlvpqsnqD3rhLICRKnecLzy9vsigk2+szV4Hsgr3DGab4w6gSZRSB1YcQ+fF
NkkiN5+9eRRorzv1ltZpk+AskI1eoPc60Zr1URsDmoQzfDsYFLJVfjgl2u3sAul5CGJXXliMek6d
fgW7rEXUAKP24M5Y5UAKedwlBG4nzu7o+osaocJYa6irZlJu/qKVqvHzX9H3DSWMoKk9WlQM+fKS
VcoXfThDsJ6oA0oCcXq0ln7wGlAQ7cOcDvJ2pqkz4ALzwOWgIo7mGmV7q/qVjGpEUr0ebXokpgUJ
yLjTiqCXyqXxiasXW9UslhzjqrtLW8rUvJxHyF2VfCiA1rESWAjt0rpHOiIpZ7Df73fcIaaBgc5R
JvP9AGnJoGOTiw5jyRhSyDz62lgh7Qh9NyGMmJfcZ0jvGOnAN7Q6138pY3u23mH8IUwX5xmZJ0oB
qo8K9XNWelk1APswac/uXkA1+FpaiD9VExpdvGYw5blce2otNZgLTa4E25FjBxyXfeSozL/Ybecj
mx9KJjcVdeZOtiwkZdRpzhVAnrcU8yqBQ8zZHz/qxBrbwahI7ZxZ9g4aZ/alP78o0hjMFDr9DrTP
GIfZ3l3w7hYUPCsI2yjRdwDNEaNryaGkmcp1rC0yDPdG2zjFq9jDlLGlr4rrxF5fxVAMKeOYb6kX
c3ngedjhlzZRdQ1/or8zgCt5MKmQzHHERGtVzssYyWCrOU+RC1OKhY3ip9UlFeq/7FAn6XQR68xk
CcvttejsWadBqc+0xTFB/CJz7s/eV8D1JPNqOt7Yl8iSsm58YDUZv0zmloW4XYelu0ahcl8gr6Yn
1Ih6qu5fmQ6K/emZMAwX/o6RzWLVlC21g95zkrvtQxJ1s2xhRcUsO4me/1QDUwHSWAjbP1vWSP1E
9i+/hQBmYq88DLHQPJTHP+S6cd3YToyZLfyKp74es3fMZfrGG1Z2UqVHXEG0HJI19CH4HBhb/zgE
byPfoo4dMNjfKRhKbmeUG71/CQYAsBp2TabM9YxffNmGwoAelnD4fHnU0pY8HYib9IRLhWAYRi7p
DA7kAMVrnA/Sa/CjmQsEE1XgG+m5XdiYYUtP6E6DMDNwtgKuHFlj9Ll44KDPJYRc48HpFflE8FzT
/y2O8loPnKXI6GbfnDJ3u6CscTruSYgigPZAyX1ikMOeNtMJj4ByQzXEzsP58FYmSC1yKtqld9vP
/RUh1b5g+F8hXetgjkNrVvSFOrjfeuI/H9WpsVc3Q+2PogedECSnAP/AgEbOnNEl3GkoM8UVvns/
crZBnngwOG7KjtEbjyYtGlk1eltd1Q0cU5GFwXhfjyA/gQW9OTjBTQ7eQNhH7+T2hslhI62cq2Z8
DGT6NlH4EemSL14s1SSIa9WGZgHM6N5xCINiTsdCpvJF8kYq2q3lPAI11b722qHfCJli8DYfrDaK
q+Ml+cEI0rOTSDNqbKNvORAhw35Ga0SB2Qkx0xg6exmJBJH+FT4i2I0QraP2OwiLO6h9unBlJz41
zAV1n+IPaTjrwJaLyHvig7w7g7nuv8jqXoVF0Xr/KKUvnm4DKFsgsY3rO1bzKe4urvLWj6pso4bO
VXapDTUpp7Wex9K8VzCSst+LfeCxbBYXoZCyPUCTibh72ZyRxgkGAk65ZcQxGce4IBALFUUxH4A/
zeM3dEDm8ANEDIdyoh3rYkudicJocVBZZEL2yqNt1nuXzfrGRaUNdrDX86zfIPWVc+OflZ4Yv4A4
JkNtywFr55S+/N2t/rSUKQj/geKisH7VtR3uOCvHvHGVk1RAwblfaP23R/GiNPKfl82FvYf3EAXF
VaoPC2o4c54mGaMg5oB1MYdsR2n5Q9WYG1JUoWiLXx2L4WD0WUGydIy2J3vHlLl79yYLblBJ2rmr
30dnuDL2alVn7h1TrRYuvFOSdwzjvZvpaizN0Fzv7qvf7ZAvG2QK+T4TZJ9be6jDk3gKIaMx5XGS
zdcPwojONvYnkcC3ByLF+DpFlRK8BdndXIPbK7MG8mcHFx8iOUhLXHJWRGH4iqC0XZs02Y692J6y
/d9/0adpz8epGytecWWHDt8H9HL2z5TkZxCze8q8aP540h5x+nG94/21yu66+gR5Cl8Lvwmlk3cy
PK3jf4tz8ffD+0w95kdivDb7FeTLxbU4FysrSUaaiUt/Apic9/mFUPVOg4qfSGPHgUepK7MP52YT
l35RfB5jFlYPM+hrsykHBuXKnBIO3w9Maj6yCf2RPhsdUX1DCJBE+b0dkfVus2QLM3IzL3Ys1mbP
eM88bEYoxyGllhqMmT3kxa25V7/PgYlDjUhUH4L2Ogn/BbmMv9KgEwT8O1/MbYgEQcaGjwWnmEAR
f7GI46uTDF4IZi8NRZpuNU8ELIrvDUlTnAdq5j6o5wMncy+VpmERysQCCrLXuzKpBKLRwfGfxq0y
w5byVTUU1nXwEIvVoMsbC0go9rC33tM4gBDNkbGaoz/pS/qwpU8iZ/olGJGflN77BML54A0VylNZ
b5Rx1gJ/Wlwf0poLM4IDZdnF5xVPauyR7yxztxwCzH4go/hNwdU8HvX03q834tAHWiLNokHrlUkQ
7RFgYv6/I2rA0VWRfJYCTlB3CWNVjkfEHt22lkNBRDy54ObVggQFy+hTX56zBpGJ7GBd7pOiMKev
gV9QBBDMMLtZHPpkLo/hMAuV2jjHotGD8ymtGULs52QTfaEVyb4OmlDPQVRJzaywLikqXaOcI3+j
2xpnUBSxcx42T0QiP2y8tBfI5mvz8iEWnxJV85CflIYA504z0WfDXDJL4/96D4pMMYdxfkBU83BR
w35fTZNuyo2Pc3xAlsV76D6+sN7nOEfQJEqNrWytL+0Ebl+rvNnrTPu6SbPj5SdPyUy00qyZ705j
irPQCBxVkRu0bFnnpb7DSogwahRnEeMigepUjlM+vvIo09w5/y2jjei3zAgkvo7e3xSoTkDUR9L3
Fv7MikgOflrFLmxtjVaBCFaNYZTak4ojpJTCWI0lA8Fetg/GitRxcDzjuckcxRqInxxu+VqM6IkT
HXn2k6ZNX+fdkCOtfvj/4wkRNadmB4cMlYAM9DowaB9h3TRo4s+pxKskxmST5UQtgmmcKMOgcJMC
V3nwTREdXcEMIHn2q3v32XuHGBuxNhmWijfvjdco2nZZ7IFfm7wBcf93oa165x0R0tB4pN09FSUf
XuMYrIhZf64SBJ4pxPD5QyN0yurJI0T5NoFY/G2nEhalgsr9p0B/lu1yUMf137QXqGAUtIjbziQI
p61WPN9enUr6mwyyN0GikbhRSOOc2n38dGCrwpgl7srJ09eQyMPTSYsOzKJWc3gD6Fd77LvETE1j
jhKNhU20QHv8s5aVEVmkIcvBj2jrTorEf0N6fa2xOVBSeivweoSrdezbtjRhKCUPLmIETlsiNnNY
uAOKx6Pl/Pgr/8WXEIQswq3KwpLrYvmap3VfJL+MX++Wy+O9pAWcdq3BC3b/oIlvyYN2DHE8JHQT
JSeN2V7Lg0Bv+iKhMR/d6AdOvlBJiPdY27igoazQdz27mLdd0UEvPwSZ35EB2hIvaZyVrh/tvg/i
AIhA4IK6RV+RN3UmJTV+z3z4UbNFFa67KAgS0ONV5ZKwzJ39l4y6s615cjGyjiN3L8zjnWIMZCrs
ZhCVaXOvtz1T6HPkspyrb8hMxffbsYvaTxaF6njg4w7y6Ao5QtAQ9tfY+OrlLtU9sbI+YbY0UjE2
eLs3OxiIHsqsV3i6pcFHtkiaWy7DfWkHAjgZmRFvDf19b/96d9TTbexvz3oHTzKnSla2AXRr/MsU
cat9oEyfL/q9wuaLYTUuklc8XrHEk2f8u/D2gGQ6UiD0DixwNamVgzFKm3+9PwZ4A0BWVyVknZy5
3ylkQapEPOihYHR4+Hh7E7JsBmbMK/mtb08rqekicJO+dAvbbjDDsW6tD5mwCR+5s+XdlT6hI+pU
M3vhoLmgUF/Trei0dogJaszqzBn9QFxjRP8MVOhTTfIPNo1xC8lkDA/JFDkjqU6uhgg/BdK1J8/b
nCBjInC5slPcF88tjKzxsprNbfubN/IW4IfS4DZ/1Qa6i+lyGxJt3KMrbkU8XEVuLyic/4LPB+Gn
k9RI40fdb+NLI0TB+3ieO2nzWMAcDABzK1fUAqFtrEf4ot00D9cYidpncd8G4zcheovEZv/bHXro
rnHOsBiDdtaXINnuigZYnGgNOFpmkIc4iabvzWZ8vw/0can6ZKUQEJ4CBFAwuBMAPPJBu6I9N3td
ivsYLHZa06OOZnyrphZEtZekxstPpH8V8k6b/NTsgOHmC8mLnLKhYD2odYc5DWl+mDWhjk6Hf/De
YHiqH7y9HcJc80LI6i1SolnqlxOZD4Ly8xW7vfq2Q7vU3HK+1fxj5Q0UFN6IKr6ACEZow3B39Zu2
5VUkn8VEmMW+ZgJ5XTMDNflLbR+qxWYrBUDW31hDAKuQjMaZqRDtHShKoTyFFF7/Wh5er0i8R7CG
eb7jzRhzTDyfzqc1sipRUCO5Wx05YjCzN8cSrLH6C378P502SssvxlS8VAmuD5etjwwZbLW6Wdts
oclM/501mIpKdygBo2LKXU3Vof7JxRwkta5DvFF8IwpWYtU5fRNVd8UC+gpx0D5+/jz+KnqJX3ix
XDUdeLfqBPkB8IfWQT3UsoMH3VX19X9LEtnQdx9FFNfAWFosHWk0iQCQ0jUYh4fvZQW6pSuBA99Z
z79TceBtksEOm0jMx8sZx4i49H5WyoPG/RvtrBUDMOZgpXYYZPf/7mhkBmSETKD9p57Agb9SJE8H
cL7KiqU10/GinEYR6/r6g7gnaTp6DaRsHhXCOYPLK9QKFV7xBRqQwlAbcc8nlhZmDV4mzt+mYWzP
aAmrN+O0JUW/7oklUsmXX1dAQacLuEydGpAIziTpKWjHJOj/k9MrwUp/8kE6BC3Nwdqafb5URyjP
/AMJHumRPivP/rCzmRofTseCw6EC1nsPrNW+CvIDPYPwhPNnwV8SUAtZ5iTl9jZorqFf9ygAUW3j
w3Ey/1ozRW7FQ+i5GNaMJgdTsLifkVYi1NwJmg88oTN1w4yaU44HyQMiYfQPT2DXAXZRlWwCg/bk
A1/bsFBfwZpov2/X8qIIrE2G05GAA8jR8dmF5ztXX8qOlZP1eEvmblxTUpjhI2taaGmVTnZCnO5w
IROCLqC5HvNvpxSTbM/iu69zHHSIKw2ZcTPTkpB9Z8SrvsRsFwUn5CQfFBGriD2EMPDF3L0mHfuY
ff2IMcca9j3wlIGq6DCT3QC/dTs5VmBbjetG+r55Qo62B+wQTlH7Hnu0WcS/y5cXfUQ+c7Z7sc2s
SqFuRdrsUhvzBXoLD3BXK4QZJH0y9wjUUcpt3sMPhUr+jzbQSOUvQKIi+dRSLxGi2aHfGVc8G0By
jjE6RVTkVt2OuiZrEUrUvULT3ryC+PNCcfAfp4raj+5FvbyaB0qrVhLcfislqmH0V5NW1xivoYtn
JSmLLMOI2qPUcLtNFXR7piJbplc+hxBCDNKGe6hCPiiTxhl95xF3GjdU+HwtHRDJQYu+H//vr5BZ
vH17NNcAnxRACkC+utx/72YcIVRhl4XmVVINTKb0d7m8sNcDSflUyjKqFJytqqRLDmv9ySxaR+lE
iABj1piARmVvb4gR8xlsn0ybqHnm0nUib/XQqcv3amTmOctr1PyL0zrM7EewqYN+0o+0h9iR0UmW
UvCWO0MCK3fp38xw+XJKEsCSW1PvgsfVDcDEhb9SZ4h2qJswr99KWuXPqprflDmj/Ngq4ptHNzy1
h0R5NDZmNAwvF5RiQ9hQDXzTT3GyYfkqfOu/76VJbkErGf0uRvbeVQcEbRUAvAlD5Uh5PgHQezCb
cNULryG0Jv/Je506lio2B/oS00IMZ42Bv/D3/ILXihWnkR8FEjcQRe3J44ZXhuOX6K/pa81o2OdV
OH3HwvAB/lw8usQItmsKlZTyCPjACcOUB2lLCFWa4iuv2KmmDvtYD9V31f7QAITC9xVc7at0yOYh
u1UvoiMqJhnp+FnWY3aiJggaoVjbUjw53p4yHnPWIs2/H+n/+ozuZ0sel0U+IZd92AiyV5OyRd0v
FQg4BdEu0ehvZoYae+9vOV9jwCYscY3+l+PLeUV9lVLp0LSJMGQN1i5JVdL+rQ6guPRnX9b7Q5se
E65W7AajgMKk2vEZUQo6Ph1dP9zG05FMsKWGwYEk634u5aw8CfofkjWA7sxvlz53E0eL5ad+ehHn
sxMte9f+8g9HWo127td/NgbKXdg/UtAbFrnmVcXBXAVcpHgnwtQgjLhdoo1a5R+a0mcw893R9sXp
LhEpbN6h3H2yhcb80BsOVp3Fxq/HZm2d+TO6+RpfTGu1ZJbXiULHrXHxX40yliwwCGppyv+91jwh
fdRE9qYgKruRSuF723B3t3j2H5fiLFZLi9kWdwKqLfBvgC5jJKzudrf/fy/zhGxIROT9mPOGeJe5
liwIINEXIFgpOwl85pQ2wjLkZGzYL0XxvngwEL1XYmr1WG1bxB11/Tb/CIWkjqQgrWLq7Dsyuej6
oedvbx8SoBPP8sGC5R8EUaYctdRGiG0Mk+kgvcuGtSO9dkilgMNCZYrUZy5/s7nUxEKd8K1vhnoi
ULADAmX10sY8LVJ0jWRzDMB2rHPtDjx7vlCUo1Qb/RapSg4qKCBtJJ76WxgBJsUGzyoXcvn+/I0M
rZtRHvNgFAR/G8gyjRGnRNBb1fIa/5pos6ELEt+oboncBh5PNHUNX72ScZGDwXbjPATmsZiF8+IT
Lt7ED8HIuw+bqWMpKn4hpWx48SSKmSuPOdhY0YwNYMh1bh1B0jR6i9JsZWZbhoj8oVen0/9Scy1D
jXSWMLFggeL+7OhKls1WE+7QQHiFYXVsIyyU4NVm9WuQA8dYwyJ0Z/EVglFLQBtzIqWE+MF49kn8
5QL5bgu//RdQ0TzCOTnW9dsu71yKpVy9uKPyEwFAL9cv+Y5Zlm+YdSaIYclb7daKCfpz/1sacRP7
AN3acx9hwf57w9e639H+bPvagVzHEAno2ozafA+ytBZtdqywD7bganqptSfcpMTUEOscAEmyJmus
x8R5HjZy9OkMX58cx7oBJMcbSAaz7mXq+zbX5LRxFk0sV6IwGfgGrpAUdXBh9QYMwU1lWj1ETlYN
KAW+FxChr+odLRllpXSYQTfWawHKb7pTUV2zvYGgHzfKhsy4hUXu/49ln4NTnVJm4aqGbwtSLUW+
OPSEn2tM46h91myIEM4SvauDXpPdG1n57nF0a4FI14qmyNYyGpZg0HfbzJYXzCbEuwRWxPoZkuxD
WgWV//Q6EiwPgYuKFc5JMqQ4TqPVA3oLoOuCbIeIlXdr6kqqDZJAkCWYXNUqsSG37U9zZfM3kWo1
EgPC4ILbVmehY7F2vsZSBND69nl3/Yz+RkvrtjRJWU1q1EvST39iDNNvi9HciBanmDTR3y9Vogb7
evm3LeadAsesQs5N3vyxy5hj4VUBAfa4G76Umx71RFgrb1ujEU4W0iePlfsKTmxsEMpTjZLJhx+U
8/xcneeU1lqqCmnZ/76GKDrrcdQqAP9CySgKEi9c+FhbB0u4m6AGn52KOoxDcjhk0Cr7k2wNCQ4T
RWPSCKWF0uNwYpChVuc+86lSCGMukL7nqZbGsH42ptNlhRhk7MDKLQtdEM8t4DkoTbKOyJFQZAIO
MHj0+rdcuH+fuuQlcdIXKWbBmX6YKnizflgZasIGM0TlNTHVmTLs7Qbx3KKByEZm17MFxAQD3qtg
2X1zl7LIhHxY4tcBAD+Oy3mLGJErJPTbx4rAvI73XkXHcyy1+VY7SLxyMChW40ZAyBc+zi3+6uuj
cfxtN7fDh8NnO0z6G1Kg/81mK1/cJTEYwzwoPCT7fBvDbPZue8M4zoFlt92Q+iPe8lc7bv60/ADT
SjmOH/QvcXGZ9435zbQqeS4xoUr7yX7uOCCFL3lmXHPwByrzTxsNuSko3xYKt76al5HFJoco6cpT
yMEuO0dK2EjFR1ztNBX/xz+LJt4OOzb5wHBkOqhjAPiVFCVw/3YEbzMRKZQhVR7lEAwmYE/Vrib5
CVNtIXytgk8Fwb9FP3256poR+b4M89D8V+sFdyv2JfGArderT5iJB6mXQLiUNTvTbBw6J+bkisd8
IRJEkWpsA8CMJTuxA06xGEAn1PtRjnsJwCqMiZtRtNyC0D+zjDaI5c/hbg7VlH/ulT6NjgmvvgWC
YvdK6egE/orbZMBg43JK75utQzRfxQOLeoXb1pwnbPM1lu6WWKIz2bOPYQEtBU0oe3sMrDskFgLF
VITH5CNuH8q/l2MGLVzR2bPehjKy+nrWTdd2OLJzTBd4qFoa+chT7sEoPBW8loOBrQSj2InmtsaQ
LSye8ffWToEGY0sUBKXUSdjTIV7qa4KzQxVpmKUP1HeNEKWMH1sbb5d9TBfjSqSdt0FoSoSVyYzO
nfiacznnTk1KKUfl4lcok1RdylWouTDxSK1RhhQw/UmukSF2FN3hp41OX+TcwC+oIVgbiJLUCK5t
601Yo38ZaHTFixZqc55pWiyXD1QaVo64i9UcIWQlTw7pV+HFPE64M9k04M9rn7X4DJhwvoOWzY6j
aLv9Qsd0eGlnieFFOiYpYAW6r3+Sn9eZuKZMPC3E0825LPBS7p/S03NDWKl9jPEd/Nch7bB1OlaK
xQ3lBXLLjX7AhZcatAAlozbJncjprViuaNVC/rRUS4UxdD0xKU7D+MCbmnAe4tPu3XTB2YKpe43g
k/RP8eceRmxhSKsClTGYXZT3cC2AENArFcUvByigJGWgcHwZ+nK1JbHLA2ssECgkymEMEB4AOPru
xwx2ePj+oV5LcIu9TWLBh7osLIhDzCdpoPc/p1GUT4KjyUPVMSw207ATL1nEuZO4kJCYr2ul6qG4
fURnTZiuiHO2ku3XufyxZLAGIY/14A7N1qofxCWNBkFIzooA91d+Vg5Cx40b6ByowXUrMhwUlr0T
EzfuEqRlMsKIxcdjfRlCj2zJzRpZD9iLD/2ldS8id8pigSrpw2SdNlOEwPlRb8+y8gWFNaDyhy8T
Fn8ZKViH0MbDVl3/C6IOcQDrDNUMIXHUvExlyPgPzhVspoqXChl7mUio2BoWvL1yFJjX3yAmmO9R
z6ohz+MiUsKI+P9AIJPB7966FC9VttZji3n/wztvBPxt2IafcPZxO9eWgy5hkLs+SHwiyebXg6Pl
VJeS4V7pY9FzTNrAf0vMuEpTP/BuszX0RVlzSll/FBbOzsXp03XJIoZ8PMEJfRlU4yJs25lwxrsm
2p3hZE5UNxpeme16vBcb8RBJy83yB67wgGULofpcI5Uyfbup62V5Gq9dE7EcErcM261h7ghjYmbr
05QJdb9f7M0oZ8PRq9Q3OVg6bYVYaf/ICl7uFVEXN0JGehKFNszu8gMBe/bXjwqFA1JsVlixYC4X
zNr0PXUyVzVCe1foOZ+B1Zu4P1K7MzAxisMExEs+MvEcNWV3dR4i5hI0Zm5Vhetdd34LuUKtcbkU
OGa3AHI8RWPI6xS25DwnRdmeET1v6C8ofw9zXGeQyzbbloUS7X7j9w57aNmjFWW2p7LvZZLs7vF2
9vQM57O4k4Y/+tWK3h5A9f4wTeTcp1fu3boSLPW9quyu1p9C8AO12mDeaqCwjsmYDtFiPra29Yk4
KVZJbsTCp8I6sA1CkHBiGsMq1MzF9pzF0qagiOcgQ8+EFjdJwVKfARkxV34duerLI93x+L/nvtth
6B9IijkCsFU65o9uzVrq991ZHHRd4mQ/dAGAc/H/ZQ6d/28iis1SoLM36hUUWeE9Prgckjz/sZKl
Jzr7FXKymDVtScKHF1cFz4vLSwcbsWmS2B19gcbFPyuWlVu2d5Jv3fxXrB/RzaU/HJSG3Sp3h/a4
8xGDM07eiN/vrdxNwzMOYWYYmTHBsmjCYcIaym0itsuOgNu2H1cdfvH8QAhh4tdsWZELYMqBxQFa
zufrIOz5XwgvhS2jziej49lI6pvo42lO0JAidWxxJ+EObS5A2bS5xq0CUH9Bn6O/xndZIxh9VI+G
BP5qx4Wc3mSExNzQ5C4c/un7J+lTEsDTa+1Qy3gLLtyYzmjXrGecuu9gi6MV+m5R79l/j0l0Vsh3
71UsaYbJt2+SXqUoV/YjoF/WS9gtv6VqaZ4dcFlR33Ohu3MS8EXBxukMpAR2g9aBI2+USD/csaPH
9HtsOrs1vmh5c2+k2mLMAJJh1ndhL9f+wdvt2R3TWqOhsfzPnA3v5SH8mcsKkna8XMkyBNuZGn1l
/J4M6kvf78sCwCl+aaC4fYqpWs6ULLoWQSRuACpCnNBm+sPS8m6GeNDqvf5g8DS/3LckI6NEI30b
ZkVqYNwJZ9s3AWcFIS0MMoW+RSIl95qHhm0h8cZ//R17fnJxVYm1WuwixhGXCPXZpXqL15uZVpgE
D2KFJOVrgPj2LzibUnYJJFMbVphbW4cLDtnyAMPtufamtqNPRQ9zFA6WnZDowWI71CvlqFGqKlCO
fwgR0+7GB2/zwAybU2lbOtWIpMYhK/LFHnUbyl1Im094n0j+hGidcfQK+FGqMxLXY0v2Q+zYZsF6
AgT/gRocVcpN785xsgqAwhqyJrQ26q3H8KhQ6Z5v8DoBhikv42VE2BYLjrZGfd7dUQm+/LEre7wR
bhJpxkJkcUXAZIlW+aV5usZXuiko/VvqTpNZmrL3meE6SWrHRZv7cSKHyQ+Vgxjj6nwm9v8Jxn21
rqvfRe77EWHLs414/CA/cIl7yYWS8qNa5hjdVqan6vFAhh4FhibY5lepGMXjjq0TlSuka5o/dgoH
FH4YpKyhBkIm1Q1xHs7M7sLykYPEDMeM4fGiGXUWj9VC24AujdWbPuKljMzglTJTpnMjDtOPzUNE
/b0gPaGPFcr6DzzxQYLs03mhxU6RVOAnE/6/bkF8qGRoH8GRejcFEYRO0ldnWVSF30zOSfNrshBK
1yUMpr3LQ3GHtBHsVvPiETf1IRJhxE6Xy6fYFFz0YuD4vfySJ4se74N776IC5jRxb1HFUnzzVZBg
DwCXmnCYOLpQC0Od1ESS1FjrIIKAgEY/umV2ZbC657pd8u+L1W5r3fYw60aydI95owmnZif6W6pj
dWRsICIjfzAgQbeBQCtaCPpE2DARAlJIuekx0yFWnBDIOhYhcd+evzBPutz9fPHb+G/mN68pRaKP
tQvAS+DfzYlTPMAzoE/cvST5OAqDSNJx+r0UWibdG1NvDDttfIspuAIx6fuIob0hzAUADG1E+7kO
EJjA7BG5p/tRztcjLZ7qM2pELvPRq8PMshe11UWYnYkZuh1qg7dqb7d+yLXNAe+2S+vP9G/Zf1Nz
5aPmEJ8Ot/5LwzCDMvyd7V0u6/DQ0YDxYtDsEkCUuX13pAHV31P9Udt3yJeIg9Yd/5H0XhinGFu/
9apqmhW2nNrcKGQAb/E4fKRPglm0cyfKCHlEgKGp9MorWCpk3PxBWKFKqwkkunXk3WZg55GAD9RT
HZEILeraCYpeN0nQOVEsmIJcN0w9d4BCZmdU58E0CPIkg4+nqf05GaLXJzT1UR6rtXQa7ConOW61
EcrHqV15ZcTWS5nFmQe7i+X+4c1ZyGHFHTmVs32/4K2+vw/m9vZQSMrVBkFUpxWAl/IbI3gzkIfr
+jb+JWxfGeJbx7hCkTKja1wThCGdyp7mosITiJUL1kGdPPiN5s1x+3N69r/T9C/jGcvEZmmsY6qW
VRz+alhjE7zOHgR6BoGur3ZGFJaAsuerFOiOwzY4Lg/5j8AJdtPHlW7Qj71j/w0d4NeMb1cxr0Ou
NMZ9tnqaN4YGTGBdaZT4qEg2nSBaWnhQ74KPpzf82SFDlaUUaB/AoLVhawZGtfPqxyT2PqToxiJ6
6tsnXkMZJIL9KdYjiRn844DemwZWEPbME7ayDmVEEm/6Z8AMNma45pGazLAmfPiul1wG1cJeJ4X3
3x7plvWuDk6VYXQLWnj3WG+OP5UvQYHQIPGgqKfM8P/NQJ+lI9bNV5tsZooV0D80jGV/rEVIM/1w
6uogxggedX8z2TJrlb+b2I+lQ6WFCnybjC8brPKHCD5M48Qv8syXjWj36tl61GjozJE8exUY23kr
jrKlXNA7/87mFjnPN8j1byl8ka4Zr4EpnT71j/qyYF20K4vNKq+oYjwJAubK94mqK5RIJcr1L8I2
wwLmAC5J9vLOIwDKlZtY4VZU4ave6D5eu1iQCAfcMK4XJ9/kVbmFtwbTlyPzbnY0cP7qSBbblRXP
IDuzCbtCO7JL8xIm56oitUwR52WKNeRcoo6yMzCbkbbIK9ntt9VCwMH02CplpRxMTEKsKIJKku+V
v7wnBGzJsU7cUf/ddswEHNC3bAIOPn0Q5tPhv0Ug0YoR7xfjIkRgcJ+SJkjALsmDWmVReG+EcF4e
bruby5FofGEsPT8+Xq7pBpnknu8lOfIptALwTQnb5VmwKFlUjig6Wy//h5s7MY1tAvZrW4DUo8Ck
y1XYeoTCK+Br/8yD/IQokp59RtCkbHT9Pf1pM26GC74dSfrrZHPEq9XyMqDZ43LZRuBbmYvdyVvd
L8acVFAUsvUOAgZsw1INDeh0C5r7XAvjuN46jiFaVWwFnxVsa66NARV9tF1QSJmeqwAGgTygGAKb
l6Hvoj3xrx30SGXoGW/Kr7KPBmZxnZyTTjMt2tUd5LlLmTtNmBJr2eod8A2dC01Kt6ysJ7XvMQ4y
t9Z5dhAbCnVuDI19r9H0+YAk4RBPGPiKCzkWyVwXtB5ffBtkzmGC10+rhAo0rMtFjuL6xVloljch
bhxjffo8KkLhAURMTadK7e3AKXdRHApyG+Seop/DtLGgsFapoLe/djWCE5sP/VNRh8M+1+qs2I6n
9d9Y6q0HGyehCGRH4ztMoJsSJMS1xqGuPwHBFepJ7Z3sDBma/qnR2yOlvA7YKzuHE5huhivQcXEs
PdEJwXDIIGXedYlqAty+mu88xIRRjc06wEjtCz5LueCsQDsyoe2hl6ptLjhK3SXhkqEyEkF3Hh0k
v2D61CJBRJmMckDW1d8Sfc3Cxj83w+gL5RZL3dHx4SZZ1e6xbpbLkhnehSdNleECW0wzxU42vaP7
Vms3rthdywvDHPfURCqD9zojOJBEIrjVPJrdukMd7+C+GBmKSrX59RfDAymquxD2y2lZzZZFcO8X
YUF4HsVRGMZ4EqMm9unrGYznKioWh5ypUd8Rxynyl29Ywz3yR39M0Qo1HnvQph1fip5Hc1YRRr6l
0BHXUdw+vQdRFi0WaIR4Ib0nwKMbO2G0Hxzrpi0jdXWK9SvNbWypxvfi+lZS+go5OXu6prsO6Eyt
hR+rgS9xMQJg0YqTucJznEVkHPn57EYYGwb9kwWdVATHVx2bq+GnV5kNpPP/iNLLiHdNorsypY8G
YoL8xTauy8HBvWughEycQ01wzBpvVM//5CW5A2iqzf27dlyXRADj3ArT9oIXXpd1HDJbLe0l79Me
JFqiU/MXP6ZQYpysj4B6fme2iL0sd2iFF1P6iVxwldRkfKqabotIKniTvW9WYv4VUS6u06FUwQCK
IRL04r4Pudz3YaKK0k+7LPVIVtkNMeV50xmpSf+3sWdk1DM3Ip5GWRSuGsr1xisrUTmkJDAZYUzz
X18ilHk5GAyf/95MYFN7AE+rehqoOEuxMwg/zkJ/ykxrcRO41N70vP0k2h/u0lYptniXqwGDNrzK
aaKx2Qyc9DU0iyGxRSG1hv9CV+Bii7UGtUpje7HMGe7VWFfhNTBvhr6Q68ii4D90JH2k3sC8NBzc
ZAxNZQzwpMc+/3ZsDPErglyw4PkjleGnbpX/40bm7fzK7s9dtF9CuAucgiAPmjLnX8D4SY/bx1rC
ND3iNpz1Y/wP76PLRGGT/tsRFQdCyK82arayXdTDMFGQKf7lLQVq5wtOK3F8UkVKKRvXuguc6KoI
+fHu/Yxb7gkyfLC4p2ai9NxgL26umUjmH41QSTbkwElLFLeNU+yEeYsF6fNDOBIIWmfKNNtca9Wi
3kYyCw8ev+RSwXkLdaqW/hfCqg2OGPITbuZNk18FdaYSNs9jcStTY8y0UIwl61dInPyTOEqYdTRF
MNPwh5K0y1iRyqLqeEWPp5z8F3+tu7RHc2MGFSSpdK4TP5LX9op8SxEMOl0H8HTFmdxgAycaFE2w
Xt2UVRL5l40DXzLghtmghnbgVVYMzepJe1nzdqysc12N8bjvxcAtE73ECp123L1cmXDkcFTn3dMF
9PZ15RXr/IoezCnEQ6G8+itjCHZx331pWKTDkPHWtYJkker4/wGz0eKavEM4qNXEbu1USKhOIKk/
L3yDpzb6w9soco3omwFuaPvzjQkAqw9B6K+L9+5LH0/UEGJbZEIUvkdjkt0ZRSoWFsRKCAozRXbn
aa62zhd027WklB4oxekMyyO34c7tgx/qYorObGt0CdrjH1rNC/mYKJMbKf9AiGLghpefmUzP31jc
D55ALsvJf6X48rVk19lQ0OaIbRBmowHf7N5kmZnDggMAgnjknFWRzHwQ5bKkLl0eVLqWj/x+6we+
Zm6XdC4/UX0MPSnQD94xIcqRrVmg9GWVK34ATLggFIuR7BuKaqFFnAYImZnovnELEji+PVL6Hv2P
qNg+yTqtCaAaJ8CCR+yoPEHGR2lGfN+2dAXFCLuFow3Ed+3wCbaUjwG7TL6SCtfu+kY+VheKEoC/
T/hEWqkey46JudDJ6dfRKOA6gnHHZzpPN6FkPhwkkoCDY2OiMLhKh2wMrolpz+w1NOO85lFOaiVH
103nHw7hbN237rqVICe3zsuyctObHLqMgn2m8KBywxHEpppXC1qGGvzSKD0yQT3K4gCa7GySbiT8
GAQlWH9b7OFkzdGJZmG6suMgpSJE2XuyY2jcHyezeurw+Wu+5m9XKtoq23z2fnFrD1wcdAUe37BD
39dCEivhz+3YMJ+BLYFXHn/U6lv/PzH5UH7OYYNOGEw6ZQH9Ds7X37JFTK9F2whzjKqcDXlqaVip
Go9oI6r1IKZdDPZPp0+3nBBkx15F4scg9bSJgEzQOBz7SE/jLIr52Y5iAwhRU5RioWWl2/eNii2Q
P9Vbv6avbc+mhawLIPAidlMi3j/nedFV9VVcMhBcK/uFMtpFfheUuwmvccxSqjwvuNtj/EMjkiOY
sy2gQnvPdqPGlES5FvjcFdWHmxizagW68zdOU5M9BJMv7yfbkG9rnZnlzVgnDHOsCndCT3LTMp4o
WDlYaNz0NWghJt56YZl4LDCjabHFejC9R0UT4jQmwV3wbMyRV7L0CA2nuxVsBAQW7/n6MQrmq/qZ
9QlGBaan+N9IRxoYEZxicPnuxuvlOSSjhJuI0gvcHuBVUwpCJg3bhyMzAHrWLrT+AZKI7P6naWKA
oCKvCmOFy5jz44rR2bGzimwhwfHwxPcp5lFSMGLHXchAiCrYHIeCRRFABlcDRd2Y2O1dSIFY93jy
NvNXEPfp61hzHb9MV8Igw7RYCKnqiaRSzBtOhpRz22HL1gLv5ubf9TCz6V88Sm37OyQ2gk1iH2Bv
pHfuV/XurTP+rUucPPxpM+z2QQYa9x/ytFQKZR8sG5mopQnugfbC/FkqWcgUhCe22Nao7xVj+MMg
sZOIabX+58iWpUflpCk/nF7ryAhsdCTVvLy83cKLWONAdb8aJwh0r7j1FI8kBdGExQNCMZbM4Fuk
/0GBLr4ks74TebXwDTLLLnKdPhn3c9laO7KlaRTyXp4WALlX+Qh4YAQZUSbduKhP/RRBEZs6fVe9
NtPWpiqoLbdpdW6ZMaH+8e716VenWOqxUTDz3n+dc8ufVh65RVlESKpE4UK5jVy9/UGNA39HAJWB
+tYpFBMGZqx7Bh30aKZBoczmt3rsDQcW2XM2sr9sNt/tDySX66RmC3fyDKWAm4OxCS8CopOSQCUd
jmyWFMosq7L0016OGpGx6CbNjr3RRF2WE0+PrvoVjZGf5AjZ62ixCiFax+ZWu3zqNvZl9x1B963S
kHD3iSW06zX0gj8dZschrjLoVxPMcZxY3gAhnk3jXuVJBSFBJf63z/E8wwNiDICOB8E2F7N+vv35
oqUn6bs18epD4VBpa7XpTbkpTUyDOX4y4O9V4LWn8xiRz5st/xdN1UI5vYKxlAhEZJH4OxGGGv8x
LehTWXKMM0yYYeP/3e5u1LiG0P1aGMD9laW5s2+W5VjsfHAjhrF4m0Nnk3HxEVC4Me8F7zKu+5K6
ELk+fLBVE8+tc7Ul+83eWk7CRN5BYd1/9ZFjznNVdtN8zNbfAR5SHxWx18IOO0oiNumof4yiYPz7
+VRIb7Fucl3r6anqIUXkBzZzqFAU5eRfDavYgbL5JMcWbmErSVYy+D4OjU5QyNPndTrR1FESBj6h
z6ecww9lAjRSVAJRJaUVcB5pR3/TBF0HKihwpuAKHBFPSz7EvfJzUGd/yeiTjr1W5LZeIdCPXtpi
FE+dJ3L4GSHVGZ3JVsE785mSHQdLJJLnmiQ7qMxOpvEMaJlcfzubvs/h+ujyTLyO3SqyC5eLUxtv
BsgKm+ZmBxcT2CPX7WrHq3kRoehWaO72GgXjKBgthJG+YGMtHKhzXM2F4Xf5WfETIr74Y6w3Usqx
axQ57LnkXxTIJ9HAcQ+7aOs1aGon7chn7c5VvmBTSFoHTjR9rpevKD7U2lFzzTHxIX9ylyC6w96X
tlGz0ia3XecxKwmx7WwZXpSNnSBe4wdEvkW3EL7tysAa66TqS6UprPivPHimoKWzMB2rs/EIbpO3
w3HeUZMOnY2d8QeavIJV9L2DJJnQ0UJIgyCkiJNAnr/EUtLdZQ0AVFFVuHHPak6bNwvgr6LW5DEY
GephfpnRknB47+fENqnK7CT/fLf1WwxSo9DuiYIceyDuc7UfS4RVtu6ve+StBEKe/w0bLrXuJNaV
UKtGh7KovgmZ2encBnUJo4b4BEL2djQpn/k+VqhasaqNepCxlvN87gXGh06P/DGebD8TYQbC3LJx
SbTrLCVf4Jl9veAsRCEvteEDNE0jqUHNg7TQ3Xcyzz4bbPc5cALlYyjLXKt7PpnyHWfMVw0zQe1a
kn+M9YGZ91YbILaVflwEdf/wePFUXD+ULX+KYxsHjSrj6Hs1YQmwXOUiJropisYgI8/sQDPlx+Fz
EmliMQ2idGDV1RAX4TP0lL+9VrWJPIO6r15OnLcJLWboINeL2hkXlzq09N4bqmnS0IcjLxT04uMF
cpHh32RtvxGQsHYGZ0pEz5vs+RT4JGKtcDcKdcdp08UZnCsb9cgfIwaTUErCX+gZ3el5NtbhcSr4
ZjGJDFUQd1St5v4FVWbZ1bZis0vI4bLdlwpBa80GCvIdzEvFY1vlPqwmAxS4W8/ifeH7caauJJTv
0VRPWv2Zwis96VWCUrIP+SDAHZJT254nJCDLKtKLtE2+e1OazVQGxEiDyrKsPDfap5KHVWlMHKgH
oguDSBiwqTfk837+qls61xbmYSjigSHHJQPl2E0lgkUMOA259Rmqz+Jbi9ShI9LKGkBqmDM5LekE
AyqnhgW+dG/C9T+f1qsoN1nEyziWBMFOSDQYZqfe0x85l8v9JNiAM8bLRaycsepVoA4elPCgmAAc
sCKiUzIejaGDfPrxS/62wYhcI7sXXo7y3BNk2mHtYX0LWD9vp+lmL/VwfPXboSqmhwtmC9unYN2X
mDEpO9QaT5fYTV3y70hIubJjB5E+7OQIkIjYtx+j9h8W6D83l6SQKfsGeF1zfHOYZckw/+1MEdwy
YlgN5gX97WAJWl1xINuHqrXioMylvB1tBvLg+PkTcnSx0s+OryMKLf2JxEArVsKKtu4ZdxdTF240
+geqc1xK9E49qWWmoLs1Jrf1Guf9U232z3CrvLsEuS+DzxDIl10xspBszVT24/92bbnTc/ar80+s
uPy+A5PDerEcEN5prFWvQMmjobwOZLx4oFUg4UufhVJuKhH18q9sITETCjy+gPsdbhgxJI+pLV4c
dslBk3zH/pBnqpxiVUkuSJ7gCYrLypaGspZ8hk4cm8MUCteB48gcaPCYR5iSdSCAhWwaHft/4Dc1
BJrsUn7oxLe6Hk0BcHCHWPZ7AD5uUuZHNNxM/mDsofxZAO0YLk7XUjZqJkLONQG5fno54Tv8Ky1p
E0YjtqcGQd4HBAuILMTXYnpP9QuEqREolXHBNhycwzgq5bPh/bsEMdQxf2qclrvFSGx7JjjQPGcj
ptkyJSmEo9mD9NEC0ECT1LzG6hzHUeN4Y+/Ae6oxnYl7oRLEjwXsWkJBt/0XX3ddFqItzPLvxfGf
T2I0F7H+u7C0EqeTPYbU91cyOQ/ARwgZokIO7hRGrJ/yXoIX5lh4tWoWuGpvolhbeWbLMqMSaEPi
3TWPAqiScqVCnQZ+O8dOb8B56Q8p88efqmN7dSChxLI91kWq6frlq/60Tvwx9FqvVTYEDjxt8nnh
IGi9shb980QCc1+CXBOXiT/+xF0UsJazVQrZ949pNVRRUgouZFllIXlmx22yBlaLipHMy3ZKWJ42
3vFsYX4/wAxPi34/PCkyhdFC0xK4haowvcdN6DgmU/7ES96YSzoTNi9r5LmuPbWhAKGwtPqH/PxZ
sdrv7WSdemNt0qFuCnjuHAXmgioN4vpdwUf4TlZ2PQxJPf6GpF6u3uQEwIKvOR1hDEpO73tXTtgw
nwWrZX7HB8nY+/yCCimvRfzXM+7Qm3GXl7RfFfN4cd3vRsyK9anxLoKTCfOsc01hRu5gnkEIOlT8
lRzf7C1GysM0Z7rOY/3XOi09/o7ly7xFliEtzoziQ4VvSJLt8/ee6z3pb3HU/g1xa92NcgVcEwJI
Z4Vi9Y0zMGKH95alRqGwI77mX05vskg4q/YJO3LXx9zL266o6ok+EMP7JaaPOmAr3IsrMPSvc5xx
acGYqt72YD7fYTN2IjfnDxZCzZd6EiMPMx9Uq4SiWhKpoLUKPf/Yf0KSW5xXaE0DvzF3QPXA7Zef
OQ8ByOBQrr38pqwyLB6e9U97JG2uqx/49fxlA23BAs00WbaAJ63mf4roG2XLTDZJUXDl+cW2nn3C
fZfcUWPbe5cHqxR1ZA+cb0JxZn/L6KVo/HAHQTQVwS7Hh8vYyyS8qBgQQZ7idBbNd8zkPgA+KJo/
D1hFO8MOOg09IP7RkHCPnr8X21iz1/7TXEwZN1942sk4/4CIDMJvsQCfOgFBxVnZyi3eMPvP16Ow
B6o2HanNxpPVtziTSqBVMJ/FCzbDTioPS5n8KqknCiggcTvsv/oiqWu8dMLsnep3wg6wrmjWAtmR
7KI18vbjUS205PS/tpQ2A0FkVxXC8ir4guL+CqZv6sp65dRbQqOAp/j3VI8UEx1Io+10TzwtQjx1
IEIKoFesUyBoAmjI46rPf9+U+cdF7dc93WEhHIMuO2To4ERchV/S3hJkvVBX0TvkiOprwGtNaUKi
C1uwzgo9NDZi0YVfpQYLQxNd66ne23uuOZMWAXwm6YXy937gm9sGhIMAWazYLD8DEVVnSWc4REh+
2TujIikKd5mjxrWbnvqcpaOlu8Y2yvLHtSUvKcMiNOmj2NwPLjx4J3VLF5anvuxHcR/FvBIuB8M1
/L1wQ6Mz9tB8rz8EkJ3Iz0Wq6bGgKQYOFAh57uf46miIazzshzuj093mn1UOBm0nUzCvqAjGJrY/
CnsUoLNXeCUWj0Gk2odo4WHTWdOypKzTVtP7mJuFJEdlBAeUQnxbv5MmL9Iyph3yeEVBXbweJi5+
OemcVNYWWbZEwp7lfbZvic+pIV+lsUES/QoZCUA8ewiMub6+6xGtVcJvTzeMmk/oSDKxvuF2Axur
KrUfQh5rhCnTzdtu8ziK1ZW9wEX4x3Z90rpJ1vmyYsLMBwwuUuzc1UY32L5/BIGsddKM2/QCLn88
pKAiJCEN042L6CknA+KKX/ZhTDyCBINZv6FxWXiSujLSxEf6CTf6+oAzOnWfWlX+4r3dVe0aJze1
HkaUm7aUvYOIC3bozLbnbY9Kyq3md/2psKb26Tot/RFXwyTp+SaxXNatHOZ3/tojHdUb2+pfnAkt
hvh7fLaHiVh2fJLjnH1yvOBIK8IVKUN0j1v0bg+agTGkAReRKUObN8SePOFaaBAbqcy2AsGuYb7C
dVc4vmmujvTTcRePBGICi7QcYWTmFG6BCq2lkn+0aPrktN6KZetG8HYLxgUgtNFCGPgmViud3oiG
LkaYfGwtxQrG3Pp5HwEEwGH2JaBCGmdIKGO3VF6GvOuJ0bs8FOc6+SgVH2EEWa0GkSfN6kyKsJ6K
TH2JTTDIoPENfgs2TY26MhmFPcEGLxMKkklhVEoHU/KFYW+n1ByKMZulhYjH9sJkshrUiMRkYhRH
BmOJ1zoWOz236NFQ1CgNWKAwTg4L2LgI6OcjSezNlDWyIeb92QET9h+PA++GCImZKS31FF5GrVF3
ofyGHRYEbLfmS+IHFq/7bOXmq7hRcH7/QONrFtN84VZGua7mzg2j2dITVWrXYna6TRMNINMJBIdo
u2ZscLrkd1LbAH8ixqdR/iWIqYV6OSI/Dy9HigBBxl7uAfEijPQeRAACLDY9pWr1+w30Me3yiQiw
Hw87f7v3jDTq8HAjvf2QeU7LmxFaSrSRPYW9sUcSzAPHCvk8Clyz7No7nlhGN8V8x+SrsbgR4noj
hWn50meQHSFj7qunr5pXtT0xmpNJfM+5y8lsuJby3aZzm9TN+jNeJBO2JN7bwdWRSuEyhEvU+Cwm
VicbVdebY0hDRbtq7wWE65vqA0YFmZy25ejL5qheTU+BgkCSm5XgE4nqnYsKHHT+zPGspgskNJEJ
MTSpMDBSFbheC3RWhUnn3aSLBjvN4WsP/G4HElmJYQLgSyrBpD+am0yNpY7H5f3eTXnvW6TnvuRq
PoUgNd52qk9Cr/8D9lVeVCfu07NNRUR6bMnTAXiyxOJ8CvMMAJ4NvaNCNtuc74ZnRBkCaDqFm4aP
+S5ATFvgUvL8cvHs+pP7ANB7WBsO/GxPWW25dywaHbyC50LvtKK9n688ae2Y8RQ/o64CEr7rHBuz
IzF+UI43LxBtUQs/xRzucaYvnGeuO9RcbTqxGxj7thiHQvJZBqJ1fEofk5+7E+ZUPsQeB26AUDGK
cDC64FSGPFqppEQt8H4DoKItqBffdqOQsxZoksm55poRLF34OyA4Z4ysfYkP2rZkRvcvLNf1LjST
MLUtIknTAAbhaqSLMfVncRAzkEc34qIjVnwk8oNjIP2qIAiJ0UC9e7VmYGtDbzntC6XJFNaE3A7+
TXNu2sOqYF3tVJl7KULySJOsEE7s7US/LpNFNZDHV5cdu/xlmbfv8VpABEpwBaNNfEvvhdh9lzHN
Q2ns1hZseYoa8G/SBiNt8429a6VaHLVcaG6yXIZxoDgJGSBU9z+fZTRXrKzfyog66OI4FgvJjFSq
djT1q9Fkuc/dBXHr6Ps/Erc73PrD9TfjBjWA4jhbU52x96niJ1Cn931MR8Z++hKu5rs0bEECs12a
H+o+O8fk1QWRuAhETEfNDgbU1BKGwz/8VtR2OJfHeYkMIkmeSDR986ISzRPZGp6DNrPZpIjPH9RL
ciDVKEVMDIJAG75Ah5p0RJnQIue5FDVfibc0OjYqeYAbExqGdGF7f23W+quBObJoEBFfTPwleTsz
s/mNvqLoPkF2lmalUgsyV0WgM0lmwXkskYfg7o3kFcPZTPferIcFGqjy7UD6LPKqqQl7X9YBbpD1
veSt98YHF2lq/GOHK50bcQSDpdtG0p1KRjs3t04MPY2Qxtx7WPlePKx02E0IR8L8g92ByjZtASzC
DlXsZxvhuVGKHYBmSEQomdZgnL5NuC75r8L/IHvnPfOf0SahvwC2JuXx8/ZEbKvx8DKdwKDawbQv
QK/L8f3NnSQ3YjRK4CRC+nT7Fadqjyxwlz/CB0+rrmt+SKAWHDV3IlBeJecBXXAUMD36ZNzZRM8Z
SL1ceOJIBB69n6nQf7QSSyygdJoU3n26N0Z+OdO2Va41NHfj7U/Q0iXl/5leBrAUVqhRmiReNj47
6f6ppuwjDegY5nnt0v1qql38vomH7tPanFSF2xwGi/kB2YsvRk6WtUCsyQAtwGeAKw/6mzvCOmnM
x0UAAd+52Lq6ojt5HHOov+G9GBCkg6AzZZaqKkCEupvUpgqJohuFVPMGWEwIaSnbjjfGv9m5nH73
rswAkXCfBd8IP0PZJXbwzUHhw5dqT62dOSs2qXi//ztHfhs4CGtY1Wx/DWeVWD839y0Jr9NgFRPs
u4Q/Sfrs6LfdF0rcYTFRAAuuCPsxkTq9o5wgiC8ec5GeOy0Wx8p67hM00Zn9Gkw5VT3hFlEJ6aEC
Yt7UaA1kTiGrLA+I0Ip9lJKMQa8fued3WERU9UN/6iXEaQb4PAeJGFmCkBDDem2Gyjcmi2+2oCYB
uRsRNmgQmVJfbirkpLvfNhzfY+KxUyIFn8+jrniUTxoWlpK6avRjEBTYYRHjw6ADr+4wjfSQbOOR
Vx5ZV4f3U8oSmeRnrXOtPlBiRpuMVeoaGNyVFs54nh8Ctxw4GDV56L2o9/VyEi0ShBe6yW6QtYns
REELQhiOGS7SAIxKoJFlOQTd0PGHlHVhF/wy1+TpSpmhWjhvZqHz6MJzAvNbRVB2b5aViCpswRWQ
BD/x2sGa+MHsL9EJhRMHqvlFRWVIVBqtJIibTN18n+J+rfrqsLg0xYocKhnJbMpYdwtkjRmRGQIG
9uXEzHjcwU9Az9LLi/GDC6kb2Z+ueDUAgNIXWXhouq6S18ZFNuYXerIYtXg+5zDqi/UMmhZbTquk
nibNcBK0PrN+nN9QzjxpmWn/5hKNFyMJ2r/VJUkrblrooVDUDcEznPe2L+OP0+PrzyVNCNfr9sGA
u1uIukWmbbWzoDfiLxAPgADcnM4uq+7zuIuJtpFkyOs3L6meDfx3zJS8cW4WnGWEFA6QkBI4g/1n
JdiTaV4HnwoUlWUsnGlI7OnRViQJ7uJSHsHNGlH1Bj5FMRJqhKcpFSXOBPK4CzVWOywhfbn35aGu
NwFRZn5uusanyObRnqm4axhwy83jW9OO0FysiCCh4uBONUs0OA4x2vTpYRZAtzDz+iX07b9+Wsw0
gFO9D9+eve5hdlHhG05HsxCltl0SeErLTceclnG2BhlbV8EBQ8ATtMqTOVQdin87OzFS1jRB19uL
wjb11AgSnB8ml2M3yF8JtGa8QMd5UkQOGFL8vrQFYzGWkAJ/eYPNerNQDWqeS2AFN/FP+ba6Yx8z
PiDwOhVy2ezOUUZO1nNNg9NiS7iyG4/gZCngw6m4Ysyt5OvI6ObVva69Wo2miM7KdlYt2nwKscmn
fDRkExHKTag7/rplxgFfykKsNIQinFcf1GzJmyhwm9vT0iBJqWU4pyan+YSk8O2m2nM7brKBjpjB
CRtVV00VcjcTgfEd/3QBU79OtllWHSiiDOerDlda5rAzvz2ry0ZAqpZIU/FNGDzcqiHhoAkQaSd3
soG86rwo5Z10TGfwI8CorRdlDA1+g8F3sOr8CJw2mvRxOmKbUnYKGfJAhtxtEb2lfv2ARi06Vt8x
GawhUTo+G+gVqhddfVVtWVOl4D2khIPVUWOpnivVidWctemdwJnbiGg3U1ftnh60IlmaFqugvWma
pIjU7lMeyDzWPMRVeyNyJclCmADwdiMQwPf+tnyQdNiGRX8lBIQbmrFiSDmIcw6lsiQ9XOBUtvrW
hRqkjkTgyMfAoGEPJmBFXLAH5pkfl+RffgdFn+YFxfzyrDoT2RrUP8kcWYw6eNOfzpCPykvQu6dB
eh0kQExWozxjE1aYdruEW+H7XrVMbhqsklzA9/k3J/TkFYYJpR6sPVMXgFfEvLfz1csuDMG9M9j+
XCzpNVnqbXpHdbw+RXZ7wK9aUGfmqhx9SPZZLoOdDkoYO1d4D/JcTQyfidxByisuw7LLkpRc8CA1
j+rW4pjmzIaSNpPfq650UlCgmg9FbkvOS0C9U8EBL0bH6/6Je/iOhMG3AsYa4uIxVfixGjSCExOi
y0PFcngenxPp5nBb0IO/NyBNlG7LmZojjYkZBbQifR9pU/qL5dG5pApwf3cQhtBwxDJlFej4FuXc
spxKKfom7mxH3O+gyS7/m+kUxomlfFPOoBuN9Oo/uECBHSnzX2FEErOwdcag7HgR1mMTwqweov/q
xDbqt+PuPs+3QhtYdjgFpGmKL0oQe/4BHqy7J29wE/0jPl1R5PuIN97nt+I9dI6T9o3yQs4DBWMG
+3FmveZsIsnQ/qRjufmvN7w+fsS68iSDRExuo9W7W2uWWgmTL/xzuvGKEXrHXg+X4dbIA2dghkuQ
k/10406BmBW2H8b8Y9qcB+1dwKlz/A03PNLmVkAvY+BWvvDWSll9zhHSotLi4NXNIgDzWq5Fd8TJ
LCaXwfckt8JIp/ivcfxyrYlKTE+h9IWMS2KTGuTgqn/insVZPnuD0Z3Dg+z5P1pIi5ceg2s3e5jv
WLCQ0djhItoyxhxpmXLrTIIpWsRPNkqwCMznXn2Mc2x5rWdAkM9xwvlHf953tHKmUCnfaKfZfc5D
0wmMav0FPnRWrFynPL8+G+HWRlPGV9oBFJa5++Ualj2R/BHXYFW6y4Vzqctcg4GUjMhfWmxNHEej
pTDInZlDf2uXt4sbvroQgjyUrmD0aHmOk8wcdLFuYTg+tYi5w4m6QsQ+/v0OHsg0vZucDNWkbDr+
6I6siBEW8qDfSqrOOYVoiKnTV63F3vGYsTT5Dc8Iibr71mQiBEYwZ50zC/G/bhDe+893Xdz7b+l0
qq9QUWE75cdEjKURQd07wsptldbXbip67VjyI3oeSw0G/kLpcQK1IiFNZzGkp4Ph9gs/aNS8vK0r
DrLvL5slgo6xBvaPe7E4eeWSXE4WWIbmE5HrMlk6lPynj18/nm5bBJjSFs63eDmAli1kP4ALuUDj
XuI/M3i7kdVaAXi82HzPezw67pzUmiR7hJ2WWrn3UeDTQnSv302Php+C4Ndw1mz9Ac2CbKcjOS6F
lO9B+ogYffmq9naEWmIT+B+48szEW/BqgTYIcmyLqel2Yj8R2tHz8VSR56Ez11XQUqbSH8uYKEg8
gnJc4z+v0I/rAbL2YFy99hRj7bsPExEc2jce6nfGWIyuIvPk6cg14hYEM8guy03oGNZHVUdPZhTk
wMvZykaLSpNA0DGQaeElbUxfmdGQj+fq7LkjQ+3DEEhRVVaxoNSYxjn3MqP/LUcy4Ww7sK+uQzpT
00cUOjyZshSVRNDACSmMqaDIpTfx4tO5ZH4TN2F0vyTvqgZR1rnogFv0vq6/cm8gc4KFtNUUevbd
f86sy27LHs9sZDCVfAwfQqkvP3RaB4aExCo8wNmeApCPZm6C1lyx/LsGy0LddWIkn6IzM9Ejij2d
2T2nauEhqBpHOtiBTOTKuj4sQoIs+ALSd6QX3YnK5AE5+kcL83HlMVfi93IJi16gYaTbpQ6AAeOQ
bljde3F+o/55FcqH8WY/9y9xp/WmVXfcjoRyZ1ur3I8xPVl7oalrC0E86OVS6EaM5psgqPpwEXue
fFqH9XiWddnDDxPBESZSg1IhvXvgGnIIhl/K6XWnLAPBwkMDZV0s8K+Q0bcRqWk58zyCBaZytERq
8BFj/O+p/HDZXtIzr6b986fi7pI3IrhI++kzPkD372FhawrvaypSTAfOK65lxqtRTncb0+XkYQ0l
kPkGDH+wCoFYXJmezux9IZYU2SI0gxhZFMff8TcgcwKcv3z8V5yqVH0Zj1AtR++JkDHbs1YcU3FU
zvvp1mFIEF9FnZk+igj8+m85lalrk97DM74su7voeNJ1zR6Q9yoqB+AEGJOJnYUKBSp+mg+4sIoT
dZV+vgnQFwBfg1wjHjpOV07/MBVcPUbHq5j7xFzmuzjkzAbatyUQ/tTodLwC+KFvzkdYjVVOAOVH
4ydvAEy2wZw+W9Sob5QcuLDL2rIfVhPGU+OjNeoSwTH7a34FnKvPU7DI0UNp7xhf9Vw6sBxS09s3
24FT0rtiJgcE9h6nFzo8DD/FMJKGeqXfP/sY+RLMb4/RMY3odE3ljfs9R6YBZD3HRkO8wSoGJ+C9
ERVfyO3GAkE507Aq/b/KysUccRP2tA2YG4+s17UKo+wlrbOfqGvivXvt6CTV1JXT/ONnxAuloEW+
XsSDkGYVLLgUlA9bTZsQ6N4iHFS5/e4jxBh6cbD6boLe3x5TUySeFXRaaUehD/2gD//EAIX7jPV8
mWzJNF/w09Zu11tujQUBIbMquKPLsVZMkgEUQ0nwjgbt5XY55BN7Hpu0zyMSF0C1rhmHoEIKhy8G
aboO7jTLIntgt484e0MwjJjw9yJC9N8FS5P/FMTHQ2OmLAqB5D9EE0vMDZrmKk0RcbINPXQOvY6Q
IwEWOvIBCTJDMuSJnh1TQIv2BILtpAenEtJLGB/EvvimhAjIIKNZu8Yxf9kQ4SBjsBgDDhPVyn7q
Lf1wkOX4D8zwWMMFQ2kDKr+h2g8IlIqhqi2wbDbzihPapdBduR4qcxDRDhYYLOdpSv2TFyCbW3EN
sxRzb/xL7fgWCBLsSAYGwSKlsfmdvgouttwMNLmsIt30OhWuR0TNBeNvVziHF7lv7sW8Py2Jbuxq
+4G1a82pau1ABel7JXyxTDckpgw2SpLrZ0VZWuXPb1nMi/wlrtaHc19WDR6nWF8V8kI+wJL2qSXs
7mYoXkqnG0njiXR5wNEZ1CNlCY+CTfp34asDSmlpNpJLyfcCDbrFAAHNR99xUyugafZUEnHmsCPr
Vw6aL62OjKG6p9kIhE9aQBMLpHm9U3r2AgplOFSe+uqSFwN/8V6Tdn9gdThyLr423Kygzn+9oKzD
Ss3ddtVGzxPb1ua6oE0iQ54Rv/tgXiY/0rJuWg1Vli2t83WbkZ8BXisxVfOYN1VL1aE6bWrEsp7/
pObiAchS7RbHqRbolQPeu4pt1JHLTa4Ol8MzO10XCPudWTR9bI1s8qkJeWFGmbCGw2K5ge5pvVQH
RG0+iShZ5F7JEXse2wF+A0rAargmUpvhZflVe9JlnlpiVRB7l8Y7D0iFAl1SDZsZyqoWalgrHEPc
TdFNksQyoNJnjHq9d7V1Cs1Vy3SBjhLYvtVGsagwLOC3F5ZLMudVkTL9tBsj6yX8SpAGOscCZASr
dyzvnyUNbDY8JbZsQ10Lg7phlh587PHUBm0fxHp/pa8KDUwfQOxPrio+E95qCmlLva8f7tM6qA9P
fIARgIe3Dqru+R8UgIPF5zKCgxb1cHz/nu302/YxFDqNJyrqwZFO1DFOxYU9OJedqzRxh2zYPBo/
TOn+sDfrkrY01xCP1xP7kwavClreLbT43bZybMON9o+OICQKsL9YDFNi5sTgz5meJU6xRrUF6cBv
ErxX1gc3W4aonj/GlkX2aOLzqWAwRAT5VRtkd1yhnU2xuh7zVPtuRwusQvwQwFNHtHeakobcKXI/
vU/EsE+B3CbMqGZQyjcVy58pwpicvBLz/Bh0TjWIcvANY3jTzHMjfW9HsZAKdwqorI3atMTMX3FV
wk7t7OeKOobqSZ9yUswE/+4nhf1L/Ktie27Q+R8XyB3njEDbkYI2snY0yPMHtzenBa6Nb3YuHDb6
whs/WlOA2gcy5F7MP7VJNOz1HcTTi1A//3poGjIEPTNlrGBAE8xa7rCNitnU9HKEXpHg9l56ZNWp
GJ2FPir4AxpEr8Pwiz4FRdM8JDTRzrPbBrf5lROotk6Os43n4Z9GxiQFMCKoesJkifLsxUxhQRjW
5wOZg9Gp5ka5ELT/1HLVNTy8BC2R1X1I+jHKWYSYPKGyFTxV79Slh6+T5IwmXe16pXvJDSgKkRTJ
xwLhem7q+GHmDv+RduGLzWe5Zb3U6BqKswbR4wbNJjNbaAi4YS5hGDytm57dS9AA+D+GGEOp99px
+aG3RxvW7BAjEZrpx+57o678whNbpl/MafbljjM3aBiBRkOGHwmWkJ/bdqlKixr/sWubXB8OKDI/
pYzytZrrzT7lqdtTXoNqtpjCSR0xcIf4SgeWID2nTYZpPx2sTDZooB3y2OZwL+wO2EFDco0ZWIjt
DnMqeSdKhDe3ETJefeEdbRMsUVqO9gBXQnb2zObKYExEm+fLWWjjbneSvXNW0jeRV3tXQLT+fkjg
7CW3gBEhVZz6ajbTXHQin7S247FrHgtPSiMibpgo0HhnpuVDffkb1M/PAugv1Q4JmpgySGmWBehH
u7M6VDWCAujio5e/HCeeR64u7H8rKrhei6bycdffz2x/btwT7VL8rptXIGlg9NDGqQPKlC41ysLT
wCCNhpwBLELU8+t1L9iwAOORGBWeqiRIihS8X1Rmjg1+VVuyoOmJTiAcVIXs/AoyZ4QwCIWdl+z8
361+mmqtmWI/RDzgzyEoqLItHMLKku6+0Gpq1tEzTffTseWnKLIsVw4p4c0t/JTOG4UfbQo3aisM
toS9986g+oAF9FAMOkga2ceWCQvYI9jC05E3RUB4kDRA2me+NnQWBnebPNZy3lOuPNbUj5MCbd+z
d1qgxfPYndkzXarM11LqB5U9QeqTFWmvYkn90Mjogz/172TCyDKcK8IU2ZsPC2kT1KLltoVPsHKn
MmFxwWZEaMTW6R7auD4w8KsYpNIfSI/WTSWftOjRbtdWgHzfo0+fj+qjRFXcC079OCqe5uyGyBeq
LtdOR3ibEb5KVCswfc9/emHF0Omm5rkQbqQhUYYuia1hx2MZDHb1fTFca27rufmSJhT8hUalrT51
ZC9a5q8csGnTIYIb1D8QGsRf4JQNIZP4zp9dxI5Oe7a1pqLelziKw49mrZMW0skUN7BL6Rn3UmOi
9GYJNVWahP41P3FTWbLlgTGNF5paR/Pa3BayDGJz5bHkLTfDj2umnLzT8V0VkdjQPdvV/J6cW2YA
xjSnd8Hmbz2yELDr97rPV5paK5GEUjPRq/vqpeiOlKWMlzzo/wYZJS9bLfdiHkIekUGHT4ZhAD/M
vzN6NJGikNgx6qsdC3+l/+oSl8WqUGEgoEjfWtN6Bqi7pAz/4xK8TlvOPFKlmb5jsP7f06Na/no2
tAGVr8q0uilPaumWjTnKDPDNhCvYOYnCuecwDznSdsRsXR221/jmYnQngH2WyMMOkVyASvUafMV8
q8MmPL9ZkhzT2KVnyeQfZQJPrQfB96HAMt+0h931RDUbY10PcSS0lZ/NOL4/fZyrjTzU1p85fqFH
SJFFtSSxDRMvikdetqNRLIi87rD5hvwpMsz3lw1D8r1IxPasN3OV+TvSwnyYepUH1zfR4EkvZttF
uRcZ/VKFV1rjRwMBnlJxxRJtXbqfZRteRuHFeA50pnneutSd4Ye4zGeOnsmdp2kavPdvoay6PDGQ
x6fcenIxkkI8lfEAXGJjgtdfIRk/MC1UXhJnN7Mdga3s0RS4Jtl014uYw30IoFNLUDkHyChcR/kW
4HwfdusFfYrTtLiORfc/JanZR2+hrxWitZXLSV3abioYEeLEGBuQ3hvMRYnW6/bobeu2Jk8Q3KIK
CK7YT1gg3ZDPuKj7oVv8sASo3N7bjJR3Ue22qtpe34UrBWIAJt+YcqXfVQk1Wcm5pouEE/8FFEne
Y2ac1Luh1QQ8udeS2ppVXd6hKjscdNvpmXKaTAclXHbAbLLC4dMPYXRiK235XGaqPiS9yfqwOUuD
UO9b34O+ELerCrG2gpUP2XGz+bufceUzpJshbu4r8BajAoZ1TO/TjUkx+zGN+2GbiQJQsErNYwMa
5crKstDfFQbW/2Jil2+6dmNeFd5AhCthpbzJVq0W77y38/io+V1QSeAr6dPLQr+aoeQCw1CJgLV1
rjn8JTYpALl9kqxtAvMGQv5iH5HrC4NRyH7wPS2E7txKgVZbuD1mMFlDpbghnAhQ34X5c6FNFOtF
+fhBfVw9U3+BYPIlqeAuNdXW8IQAdbcxKGPWWj92TWHiVI1JDY3QYOrhTQRG3w70rhhgalJ6lgue
lGSbQaJPSCGD7Af2MKaiHVmVCzZuEHtl4szq0YSNnLxxmFK7JsZV7LLvWsz2uMx1np1re/8solrf
i7db3nnlE5BYp5FtzecQTfnBhJYdqRi6hNaWkec/5jEK2ygPwdUB851Lej7lIAVg5jgnOdvZQP1A
8p9zEu+rXUJeQws99OYXIeHL11CXptDVHkZ4Q3QSXsTyPdnS4PRZpwFVmEleTWC5lSx9ZPDwyr/p
RPdv8yzyO0diLm1ukwlDfjdTbwBWXL3Bk4C4WARL1OrqQQPoFQRZQeFzMdGdAZIPEFGHw0N1YHD5
ZfnKd3RHn8D40yLzrJwXPUgcRQjK7zTJZ8y6lR36PLyBpYTyUS49httEs9+D8ew/LOEM/oQIOloi
S3oPr74GRsD2y91tx/0d7pjenUsPsXkq5GcCAKwgQoIVZ+JNGk4W+YqZYycqXhL5bt45dzq+UfaP
iFD4fT2t9O7/cDqmYfGvDzgZWqSxJt6rBXtKlCZp0K6gIPSr5FgZtj8PIooqNAByKAqzGSkomB9i
rhdj/e0TwVHhrs8AtiHyXfbLA5HbwY/h7QCZj/MhHGB6NDtnE1xNBeA1I48Wrt7k4dincO83zqbb
nRItRLN1agFcV/urHJ1YwlZlePd/URU1E2mCZ7+mLrVRoUvl7CMhrE0T3dbeFDmFBuiIZbKLzHtf
XpfuE0twkJGjtIxbBhVEG34y7Xpw8evedDKAIBcQsibsGblc8yv33gNI5uMqLujQuyuQ64tZ+Tq+
2rTu6HbEHckXUhgO+/Jq3pjuHVxQ15VdTvKLtijfA0FqkZPrfMx29ItyNzJxFrUGSMm4LJ+lOpoL
gApwkMQ+TuZm5vWJECHfsDJXZRG0MpvEY9mo1rZUCPadFn2WQcu+Xn5EoalVOAvgEpfd6ZLFrbkG
aWqFwYlhTCFLr4Zdx1fVdMqErO/pFSUi8DyBUZ2zRq03/cO7US/GPZSXBWz5MnqQYBfwmfsKclGC
jHXFovf28+jeXcin/QvYO3ZSy6iJxQRd0p3qe7Gn4HnCdckxNLOqhMAexvhTos5OYQM5zP0QWlAB
Pja5yfjsTprIufmKrljMR6zAtxyFHKajw/ZCzeyM1/4nTyZIbUD7KrZLbo+Qu56oBrbM9TGqlGbO
PV7M+pJpvbtM6Sj7wnAUd1+AubP2HOilmEQGMTF28ae6OcJY4ATJXb6Ypn2PvfBB3oiMmWiweUqu
R7qffl+3bIFkALAcTj+RCr5FoTtay84Nj0rnSlCNcWR821wvsOWyp5tCCRNeCpjTHPx/P2gJ6xCM
HvcM9uLOgmtsbC3pUOqVPAfJmc4xjtznc7YvCVtFkwH1+t2WAVbDvlb0kQeaRGYrQkkKAiohxepB
IX34settpjVwj647tBKHxutcR1yJqwZSRWWS/5MTNn1D7YihAcu97Go8UwY5dHmxRh0zB8OHj8TF
RhMx112WXdWhzAa2ytJIJNAioPirGZbk5SFP6W20dIwtgLLF715ZnN+BuEzs9MbXfWttA85uLE6L
4HEUIpJq9gGwKAfv7xT2AKoj5Qmyw4kD1HIyF6C21ZtBuRLEhwmM0BMXf5IsO8rn9dw2NOZLKxN5
y52TdfeLc2fh7NUemvmlz62aAaqPVpeCzpxjsC+TC/8WIQoOvG9aEuweJAtBFWWzV4G1j0yXvwYZ
0SrUcLWHul+Opn8zSC9rI8Vjm6x5kss/waojbqBOFbfRUrKrSa9INVeVTzFTqgoHhR+K3wv7N8hw
Px8QOSULoyzdF46ezQgDkWLSYhXHL/AJ7CJZnist0TS++GpHNwlNa4HWRcGGYeNtSVAsnyHTWSqj
FyDBrtoxIZy0oSLGik2borbmBzmYj0g16U2h4LDg2RZ/HgugzfdnmhUemjvYX8eU72TOpHQgXbfA
2Wjl9OzWNHC+431k6Hf3J/NY1ccExm8vcywS36U4IWM41BoxAvjhgM8sJyeMynxWZ7r6gALVp23H
AvdlREHDAyQGL5S11e10dTvMiwbCfmDhNmKazxsUXFonrgvRJ7b3VYIQP65/pf+TiUET+LBWF9Jy
jQLWE6d6bWAkdGOjBufrImdSxTbfbltTGkTo+S8znU+tccgz98MhnggJEcHy8wTNi0PkttpLBBg5
Xjti2psHGeHvCofw7CuWYv1KcckFZFMxjK3sGcrm2mwfiIaZgBi5Fb3F5oceDxZleWdrIsD1a7+H
3d8IHIUfDOo9gPbYWMX8TI40xFvxjg20loE4K+1K3e9j4qP0N4Ck9+smf3Ct9dJYINjx8I4sGURH
zGqbW6JRJGHgcp0hQCxUW0ITgBZEtrBmg7CZCY8BG59qiabXz5hm5DERBsLKcJX3qLwegN8Y6Gzd
QB/po6PQgm79TJsMa20qzw2BEYjC2vFWnSiLMtuxuygj0uUMZicAZnQo58FDYKDiDyrZQNmGXCqx
Knsv4cVgMBBSNleouEkR8NPmSW6uoH3NvJJTPrHBR+TFPIka6AcLDdV0HteAirJfd/lBjZvAFy1O
k3BywysbvSskunXsEITUau2xUOSVBmJ4sKPHfOIpC/Vts+ALiCQLisVTSGWokrmbgDONz8zSETM+
ozc8Zq11wdTnUjXu0D4druKmtasmJjU167tR8fJSXmQNvf6FuIdLjz8jDj8b/ilmMijWYTvYGKzJ
mJn7iwiljIJ/MpcIJIn0XBDkCrBqNuD3wPpVVU09tJYuaeM8/GG70PAx7PglXtjwYCi20CneK5SX
88DVYoqPL1zyngksLMyu7s2HxQV0uqmpbXqvGWKkG9pLNOs60qv/0YGEizHYc3bbxi8046/iniIE
x2h9s7EVO4D8aIb7F5doVhkWJbz/GAX4zuUxSsf27pjydYGiD/8jBeV0taGzyL+giCr+vzce5EdY
oyLAK7QIdwQYzvd+jHbfMz1GK5CI8dyPbKGbcVIL+bwkHR/9infANQLKy9cPOMDLQ7lGw20UtMgK
/gof1A7mB39T9Txe5cwKo5kFI4sqE2+vrFqA31sT+KJfrn11LwxiUqSfmrlIZ26GIFWf0cmLH790
jnJliBIVYykhog8RDNe+dO9+1vssOnKnnixEd3gDZ7Tutz8sr5X6mTDgyMqPC3kty216DBttNDwl
CfsrjXfN02djOREQS2isip0UZ2e035ZuZGOYS650PXd8wdnnR1htaR1uX2wm7DoPvbnz4LcaD6Lr
1b3KZWNjDq6PWYzdJlaPlzY3SRms3drQhr2p6tWeDBXHVf/GA7oZonghvqJY10eXXXTI48mcYpPe
dKiPNsGJETTp3Kdtfxp1q8/0mLw2D4z6jbEN3L6T2wb9P4fYHqo4X8nHO98WASsp3Y0b/8aEdB8G
SecjbZdoT5Y1vFU+fyb5YeTMO3M4Avf0xTcM462X+7UT13nB7fTG06EoOH1SCeVX5GSSK+INQUoT
2NxfjaiLWFuGo5E4jebE6T4S7fBbe7EuAZoq8pdYSQs4iFp8b+lu9t/LJIXs9g+n4Jrt+t5HbnkM
0clZGVcJoQ0X7zZuH4Rb8RuI+EdqNZU8NfRkp2uPYMU9gc7hMHXRFh2AwKYoUxx0hwQJGhk2wVkD
7Lz2tn+ZPHxoIdjhRLaUsSrEfODhC7LTMkv9Y2+xzIbFNNlWgAdTO98YO3WS2Sqz/AwJs5/Nt/Xs
LqAbvOczWpbVOEsGbKYKVJfVbUamPIXccDLFW+ANznfhNdXuQ34tQXLwyPFXGC8Yce9vlTHHrGmH
nTuytnScf8tWsjZIne54ckm6Udxokzq2ds8cbCTBw9k1A2u2/WMQTGJz+89048qayZhGJxfrshbH
lLCjlXpD02qnv/GZmaH377hpmCHuYqKEt+xtwdKyf1yUQB3+jZ59eugZ08QCcQ9AWfvmUi9g8NlS
7SQmR/V0ocvXNQylJDHbfjbRsl1fmDwbqYBzXi/GRg+MwtKnMXUi6otRqOGEmiBwA2SAeE4MkZoO
w2PY6sTwUsPFynJ/S1Z76dnAzIuIu9n4FlApPmZTbwu5kKj6hFWG+envq75evI9t9/C81dOdAKVT
LnHlIhVjaE/ZLUNFBaQBx/zU7igdkxRZrXz2XTGyM+PNoeStG2FtcIIqlULhmp2Rt1g/jkWOiOmv
lxE4AibozNQRgMKOfbWLHNFQo3hBkEwJNJC1Tju17iKr5L5j8wD7kjxTvUGcT65CDltkMNwJzJ/J
s1xjTR8nBoNfpAxsxszvFeUJpdoMokRCoHZaQ9FwE2BcfPIi6FF9xTUt+pmfN/Az0aajxx8BQiep
JYQvkDDv/hbaY2uIOeNKXIk0LQI1qEJd2scSjwN508D8uD7MulG2rS0swbIl1nVA8Ae2toYYQKtH
SpGhSug3dJlJLdEJ6MbBGZqVFUgtyQGFFpm9STLcEsFKUwAVRPrWJZ8wgZZ34vzYJCjObJr8L45A
qF/zoXJmGywjzlD3WHU07T7Vbnx+6gXY+gcqBPZg2aghnKATnRjpQvOPSaLmfMQnZkJojHAE1/ob
1x11xN7MyRz7M7AFFhP2DT+7zYWar9NaCvWfImV08R8DfGTvTs+c0VVVEiBquIOCdvSCFNqTMAV2
8de6eIrVJQEWLxXZIUzZG+nMVzGOro9w93ejlr5I6UgxJUbDuJcoPj+tSaBTfqf3sPkZ9yXM6gcm
XxBfgLW6s6TjIq9949NXl9mO8zPrfuBwjIv8/RHBOCnyDcZKOQE0eUeeEocpSAF+ixSDksiPePNf
JS2EUv429B0R3IHn0W6XDSCnN/2eAG40XDr+Of1XiEr7n0+JMEb0d7Jn0v8seX5rvxk9kKU+6IoH
CexgABHyMhCxySWwu68U1206yh6/5Hr6YFtnWvxZyw1qF1rToFKKhlYjkZNStHW0sPxmd/1caDSi
meH3lXCynZVGea0PUvESnAssbGd7tZAuzFEln//uv+lHSwrLF9aB9w0TOmzQ7wxq/CZYwIm4vuWl
Y5518NStw510TpPCwEBKCHUTPl+hqFrtNkJ67/3s9L9tZrY0MpgML9mC1uA2RSAYAX1oHeezUTCk
jBxLeBjU1UuL0l7R/7u0ONg7T3GPPdj+sPMLCxdq9BUTGUIy5iGb4GnnS+oiXwtb764Y7MvUqw8n
cU6nezN5pedX2JP1o3ZOa+lYov777HPdvtvmBKycAnqQupFO7t4LF3uYD6e22JGc33HmuwBjDtyF
l18b1jBNiXFCz8GNmU+T9jrD6jspb4mIGMf5ClWwv34d9hDc3Ko00B8R0VYMj4SHL81RJplaiy0/
nBNzAp7t9dLEk+TXYWnLKnGHO2KUbB0r0+yrRrslLN4Q3Mr933wzSpUpaMXuVbNCJLdK99OWaPjj
414ehg456OARWfwyD16Xj3w2wf8smCDstmabW1prVtOB8Qb2tUkVjPTBN6yrSKG9do0Ghnl6oEyG
JGwk1zf9dRBTChgb3XC4w0mT+EjvFkpQdTW9qu/eqckY6ZAa2V34dxhc3ak0P1ZJbk0J24XEVA+R
gzyp/QnB9L1a2Gclym7ujOkPG8ksG539c8Nb8DyEAiwNwWMMnvFskUyQHbPBw0du/B9XBH2+ECwp
CyO8w7kT5pEgwdFu17xC0pmcbfGt5Kw8y0pwHq9aqV1Wnp3WlGrBOdzq8jGo3on8LwRoqSFSWuSw
LSPAA75PXo0kmyeJHLarKgttsbfLr1/w5NipwOVO57l7IO2ju/qh39SDaD42tF0FwMm2Q3KN/w4n
jWPPBnrm/GlPRv0jmEJIqTociVj8IrYeUjfG6lZt9hQHmBrhzlg8vXdR18BLC0sU91tE850vPaH/
3e66RLT+6HDYvh/PUN+Arq+97cP4Z1o1WJg+s8dckgoOTEapKXpeYeUiML6d9YYxYPuYxN4s0Q/p
myc+cViLfcaBALt2vl1+ApVhNknCS/YyAGHRYBM/yPys6YrWclLlGeMk9HTNyvFexBgRwL9rZxrR
wtFrIKuQdlAtjDAtRB8ZvEV9GbsHXOD/Yikm5aEUrIR24bRtXFlroqYvdw5cONE6Jt4g94ZiUs5K
d/Hn+LqWWcxsxPDjECqo4HsaoVXgq9TbTDI//LeYVw2TZ9NybEcLHOyHVRg6duc2hbNlJWplDXjQ
1XIaSiLXyTmQCwYQMDQL1zzssfwD823I7GR6FGTWOf7cg9loeAaRXaMhVVziQj4gyYzzk1W2rVxV
mQ4PSgcEVh3NwlQK7CxaGFPmszaKQvHud6eGE2z+oihLARF5SDDR784XgHabkNza3bAknT6W97Lj
s6Nd4/9Cex4hYmUm0MKWwCTdYFbgXRLSdb51sZODdrZNn/SZh6xZt5cl+VK20y/SxbTOWyET7Ezk
IaV1SXYDD1y0td384Y5+SKaHLZwzLy3kjeFqWNHcD567Umvb5GB3qlluIlYd0kpQN7Ye+rV8O9QB
cvooodiEKLh4roJygo3tn+cqQFGe0dgvAou10X6/0zD2x9k8UcMl2cMLvw5jeeHIjo79Ie6icOz3
3642GnlwgnEZhKbktBYSHbcD64wDpo78lLNXoDjsXttlAYfktn6FXyrR+kBKKiUtu2AGWeqJTWQ9
ZwD1C0OorOaSNEjVmF/ZQlnKGiSNktdMWKQzA0qzSYxn5jrIh6au8z2XHUp29CneILemWHfo1ttu
JcstY1j5dNII+C04DD8RvYCLafUH3l0KKpRX1MAS68xksB3q5vKebAaPTcgbWQPAZlfrZQe8ht/N
m5W5nMHKZGGlX3xDNx9K3wPcRtEH0iP1sZoP0krlbpXjgFQG2B/JctARcwzL4M95mNMFUhuBuPvC
SnNdxigMO/1H7QHuo2wqDjtMIRDShz5Z/VmmtXvGF6eY1CIQV3xK3X2n7nJpXkMsQl5sSPK54xRK
i9nmHF4/+yo6m3emdumqa8F79/BQjYv6fuL1UTIv/9BbMkFVZ9cDOfSAq+czpcbKeDHRDyOE62GO
q2lQpK4Xm9msmLXmGAh+Ac12XPwt9COTdpQU/hvvrBCBL5Fd/i/l9loYA+510VOgsmm8udc4F+nU
t3+Pe2nJbjkvx0vuHV8q+vrdfhxIuaPJq+BjCDsBUOXWZi+sK8RqfILBr1Ur+tUYql0wdvIYyiWU
IWb1Y4GVutHctEO3D8CYzBY83G4mbGLCCCT8mWBmFk1KCcUDMLcdtMVGiPrGaGGxyGMrIKI2l9Ua
Q7B0VAwh65TJC7ltuFdInueaUraDLG4rLP+2pVrS3KkLrDdU0ZtRZ/IFkxtymwNffEzK7uuSVm5A
gkWDiMOHNs8z6TADRsnbs5ajo8K5J6TdpR1bhrH5k983y7zhFn7MpxG9/2lcdPGigHnZi7+A6sev
9ST39MXTgfW3AE0vX3CHqr8HFbRrO/J1k8xUDNB3JpNlgjZXgyuJ0nofJZ6F0g34csCodbAZQdyX
ublWloAVSwjqBpm/SSf7c2muOcyYWmyYQ5yqAbo4MYzefvPgU1ixgXhyC8HEwz28oRNPlWBqSte9
1wUHC94XuJkiqjHJlvw7oFZjG8xxNUyfCQxPoPxsEDF2o+VGwWBOlX1i8WmrqOMxAh7/y8UHJd6s
mL/435Zts3PdrU2brDemJiQ91vFHZzolDc4cT/I9NG1eHR1wh+1fpjo6jX7dluIAz5YeysOQzSwf
2VTmE6zhLTKScNkqrkkcmltu5GyzYTokPe5eSynvJ1xEZdsVoHuHNS2b+m6tyb/H3IFYsp4FE0fE
/figmPV1uy/818OIx3pELVJiXSPPmpAWcnXoCYXmx4uE0IuP/ZZ/htbzC0s7Fy02uBzqdfV9+h8H
UvtunV7FBPNxOnhluvKH9V6prFmnNFGXE1cAc+wGJqP440j4tSs5BkqFSduu1qzJyxz8Hnckh/TS
oRzZ7cZAM305skD5wZYgGMsIVLBAhtl7F5ujBEXTwqsHOI7GEtD5TzzARpYNV22PT94LjNKlP0pn
HVuKAX8d0TUDyR82KSGPKY+4Fynt8uuSXpgn7mH+itrnn/iKqT6qJPGqfMPf5s3qY/Ok9WkMeBPB
0TsSQCVAGjImHyeoPqmb6tLFnhviFubUI8X4IyGelBQcWF1m2BqUsVmZ+rk3BZ+29VsaxbdwLSW6
hz0er41G2Up9xlHeVBc2R3bWgxymH8Mz+/poNh2YR72DgzQ45+xTlhzUM38OMt1DYNz4vDiAE6ek
y20smC/58V7AjbwFP949WTzQUJOZX+zkeRjMHe2fCFCRiaPPIReZC/8MjmH9A4snQ+4PSKySUg0U
saTOjQAXkLiRtwBifaUqVqwKNQ7WQ37LPht0g6rdsJCm92bwtWqL7KxzWaa55PI0E2p8kCjGp/rT
AfjFdngXiplzUWBUmhcgWBDP08VF2Nu9T3hi8+Fw+SO6c2/UUTt3BqLnYOfa1i96TfgVj9p1IRGE
LkCD3Wvkn0q22Yn+IFQlWvoX1cZTiKX/DBka9OW11pz4kOnM8+6+Wljd/sudOhgIxrJoU7b/J1ic
vXR4udXyLywrKh60nKQJo5vlUW0zvh7t31DoYemtaFdwefQmrVYRzFJBKJxFOHo64LM06SfNpF4y
T2Gkz8Dtu47dnlGgW1lBHWOVnFlLmC6x8/cGgd+dD0QZXyZTud96hOyKrtkiuD2jikymM9vc18z0
XX3qJ/A3munQSZVsdFtjBR5i3i1AdVlZhJMQheO8iBV6uNgTnDQ5XZ9MxeQtPlFkLMn1IDZnklY1
PFgnInhyucwPAqz4EyaJsNi7JC7/QwG2/Qtd74vu79h09L0TgYP0ii4H4/PXg0InqBEed0SFMIAn
X8ERo+A1rP5F+wsOC8YFuxEVXMvyD94BYQ3yzF5UkupXmfXlVvci/UFfdIje5uiHbCYvJ9BIAleD
VyNSr0iofnE6ekuGPMymObdbRxuO6Ja/zAPO8ipqxZexOTTbbc9q9JKyNXb7yop4bY+zH/kqLGBp
KKRR5C0dpSFh4cYxjRY/7G36TnUtLgm+gv9Q8WEYm+TtBdB991hE59V/UQvss9uXMMjdTrZrXbFp
NivTQ9id/0cM41JO+Jf45k7POPb++TsktQItKq3/1V183PtLI8lSybknZNKEfAZGHg6tPFBcaGDn
PRhhX1kjjnNtPwQiIjB0ekjmij2vVbqf4P5fjJpMuv+bEPZg60IASVBoBjTWFznVtJIy7uw62abY
zvoUOByfWLJ+H1dda68UQ7NLHzopniF7t/EyBafjST2Ofh9oZJEUMYE4JnyPoQNA0yR40O6ED6vW
ANZveVEXmNr+bcx6WQ4BpqUWC1B3jMdUwsvn8M/2cwHq+rgm1jb0JANV2+vuigdHEIJeX3bkjeYq
CYUEQv9LmU1Ld2bc9SbOb+Op0pA4Y8x4yntg8tmP63qX38jIEFiuaVPeeQB98cgcKiLQSKCCFk7N
I79Em3vhq6WdT4UvawFAYddLZd92aDGD86Dfn4dZtPDx8BTkMpg1uHdT9h9aO8nmzCdhjuODBiRy
TQmGwknheOd9jAX8XnDlTz2GC+rXDC/I+xfkW/0T27Ng4eVmrArqgqme80WNHRNEVVBLr3y6T6O6
8zKYX9tEL1vt/FayLxHmnOm7uwcxqBzS/j3XOKvBc0I2ocRvA9CYJ+d+jtueBzIIGwXwafCrJ6Ux
2ilJt82aiUNQ1CETCfLzfACWDWYngsHhMyB53oihRI+6Lv1cMzld/7N59B4OSGoi1VNCLSE23b8E
t/aGpXbWHxL5i8QVBt1BFaPB1117H+i1L+4r4gewdLjrjAH2YdQCsO3RVCAMZ9yMrsGBpIOam/ZP
Ydp9nMz6zWEitAL7qzp/zLmylG3tE1uhz2CQ4SyBHs0cx3aAtzZhZ0oswVG/D7vWwPhnFUnH6GX/
nbEStMWfRf0g+fVuDiImuHUy3ETwnvzQCEArmHQG2ugn4WFkv8xf7pNX3qmw+cI7NkQptViahRnA
fd2ZFazCLc9p4nrfMS6SWvoXFMvp5fCg5WpCcQcFSbZJamDuCFD8HJ5wJYdqEnuL3U+iJMp4DK8T
ihCRmuK5ZERbAcL3WhreOlD3S9IcBY2VSx7BR3FziEChv+9huzsjd3RjgCgw4MGwDV4myKRWOGZA
Lm3mZQZ/h5XuTKVzh42Qsg+V46qwe66ZGn3velwNEciMlemHd33sgcoJZV2PGFCQ+UrF4bzdiU5P
+mUM1vWPFkGPtGnk+y4pHpNb1HbN0iKwbDgI+SxdCpUVijhcQqU9xezpZhBN/ESAC01LiNNNi/Do
y5ftwnZfyjUVXKf1x+TJjyCrvLKKlUvnytFic8utFioQg3vlRUJuido0q2JhTRzl+EYA8pzS+3Z7
L2BURbRoL7eOtTnEN/ipltoyI7Ar+1i704U08WlewlwBT4XI1h7CmfGw26l7+QeOV8TBdjQBjv77
1YFABqs58tcgNHQGKKVeSWp70GmT1BM+nfuHJPqMgQA+0KraUSSzkTSdfp+0YWKut7tGaefVkcnD
LyoDSqV4Ky252HIKAHkj5pVjrWKCBJ2T5A4l2Q8aBJ293WvNZeX/nI1PdvyR9dlVleZDHqyFY4ZM
yK5N3YNKlL1rZiKMpff9kjNKYA/JM5KRgLzLO17YBCIUtFPGxnGZAFxMIrbTpwKx6UXQx9uF3HZ2
9vdwF6hNGEt6tIfSLx+JhKPDvReNVePAhKBvA6C10WfLnTbAzOrueFrVgrBx6x+JQ1ShzPdSLE+p
XkRSiSAVxZl2ZA4rup6PSB1vO+EYxKIu0dym43PfS8WYshI2ptxB48QEiXfMMbthZTcHFJ5vAP4a
4z/udU3seNnmPuiT5KFFYsG78NPE89ujVCwUGecUaDY7jSA0kkdS2LMqnEzo0NjljuBA+pzZHIsS
JGx0qHb+roB94TuytYskR4NK/xm7wBR1lKUbaxWvKx26PAO2L9qqVWv29GAY7ieFHT311vDzSMwd
vYC6vSOknCNyX7M1KBTxa4qmt/UqrjRhJdfE07TkzFJ4sp7vRoQTkGPwL0kxHGk3K9RezYoDFiNm
Cw8HB9sDL3GS+/Fy0GjZannmPObBnOyZdIQTOxk+GV045xVziN5jtfc+ttwxGmqHsTeL+tdHdihG
JO3JJqTdB5+S5KSpzcoaUGIA45jxAt3WTODFeAMc3yMgTqn5TtupRXBvaTi776kiMBsv1N6ePzdu
xBrYS2NJFDhpEMjBowqyTt0VVcZhAiw7mO7q5sJXg1+grfBk0Dbc/5RiAnmYAvjvApLtAOzYhmBz
UfubuHw0TZHhkfndjYS+CwyOuOB0wwEuiUjESbpENeGgife+PTdTFSpzJ7suI+ynxXbJeTMVs8eC
rwsbRO/TXayYZgY6KaBkW51mZzjNJfTWhTOtbKcSe/dxWLARp29F9aAZPS6wDTSQLnE/gt5u/pXd
btFWxPAryzFrq8JIHAtEaXEx+Px81lnmvZkaJaC+DifXzSfPSTOUWjgCSn4OKMPHE8yw4ibSBtcr
GeeiDBkBnyOi01+Nic42pnH1v7Sryg2ssR8n5LhrNcK80w7TODS2CI7VPzyJ+W9hILFB65bjRnze
lvGsgxvhneh/e46UxJhuDkMJEMD5ECwGbwhDzU+4r/Fc+3RA/jnuFY/ATczUFUjIhy+Dng8U0yBf
OYj3GBwDzqqRcJT9E6DWXcpWn5lNQurbSJXiWhZbhOUUyHZ125N7Djt1Q3Ye+kSLA2lGcKKikrQr
1i8ZFZLQuVTAtja4y2Ksh/jvplyMNg6nC6qaL2R9dQ9lyxKWGTefQrHkzqi/pe+SCOpCapt1jSNE
kaU7M/5y4o9yHpBd6333U/LoI+BTRTfiwqeHr0p5o8nyBJn+FS7cnI6VoSyYulmRC24oM1MlBlir
EDfCtxTF9hwFdMs7EBPVVu1pGXdM7GHe8+w6haYi6MrITBV2JsvEdK3pvf0RuViPXzFBCEE0on1g
FJEtnSb3iNsOsIqVTmcFLH0tyPPg86friWc8Nc4veNY64bT4TEo/2bPD0/C3lA/X41unj8aBhqEx
aAIbx5xPURm4uJDbZJDH9MjBU7FE1N/RZHmuqCu4Fe8nmfhG3z0LWcNWYd+p/xqEtb0tXKyN9XE4
XWknCI7Z5prb7irZK5uZSPDnpigb+zEtvlvJuBJneGgHUSGXQfE4EPLC7oizympIQy/Ogf0iT9JY
ovZFD1Vl8Jtzo5siU9RIr3x3gLJnbRw97fcx5KOQrIWCoX4EeNLtBtCgZMcadiPht8Oq91gHYm87
VDXROvUG3/RVgcQl0BbeYNdVY3gS3AZWokNlBwE896uY+kNCRVO16mTaBH64FJw/T1XTDaVASwe0
YMhDEu5Aoky/73/oRqnkgtA21P4ao7hucX26Vpu97P+2+dW3U4tB4jW0j6+A0CnfyZoc0oFE7BsA
lVaJc67bXLADfmOcSqPhblefZq3gFF/7Mi2bmRDRis9xVmTXlF+y4Y2gQgXyQU6zk+JEyE51iGGe
qzBmrBTjTzVWbj1t/ke8JGevO6t7hL+sNtcG9DsQkU60+/VvPSpWXR34pbmGgstiMSTNkJCOJtId
2e5rYwN+4Nn7g0OxcddpgBOuma9SjLFfnDzga7h9h63ygrGpGZ8/crFxsxcCW+KsteqXNe1i9z5A
HNl6a1PfqYqz55V/fIzsnnDEPOKjG90KuwpJX80NVzG+F1oG8j5n4ahiO+ZjPWtwopDBrsN4aaDb
cwzO0UFoOn26Ybbl+5Mn0ZsuIly8r527mvh9v26obLa+eSIzWanMEbbuhr/B+hztqd0/CnnY73H4
7wL2FpR2GXu50K5s/2QTkEIme7VUdFhe4GQZNszHc1qXO07HR4ZcGcu01ngXvv13D3QsZN5mhf1L
WXQidXIt83z6h7wiSBqVbT3nozZNl4rFYMMbEr+06L9w63Q1gyjB5laT2MlDzXzppg/NesLT2kOi
2NYI5MmgGR/DiNHTJF+duCh389bB/TObwQZJW+23qLBaU3gR7MV58x3gmWrM2x4ZjCvgxj8Z6iTo
3Vtc+DFtB4FLTm/9mkSA9onFaqQMS/OG45qweZaWWF+BeJUz/Qu5gdBbhMtxiB5N9uSa3Cga04tG
98TL77XJDEwwhpyOpvG92caND5g41BcqgFnrNzhTOJvse7AHqwAzz4WJiO+j64bF6Rpfk3UBRDkx
3yrvZDgMxbs0R8YZenG0m9ngSko7AfPoIJDR290rUpAt7lUjpYszKawylQdFAx6NNVrNALtV6+Jy
iU/tbFFALj2nq3SvFY3jfkmlzDJ1czTmKNmv7ib30Yrj78Y2icESbTall7P0hSGIHOwmIhxsNp3l
Jkjt9uYQCOUaU74MTEqjPp70WwfKLBxH96myFc4Vwo83kyzjiX0KSumcaGpZ+edk9ca5howrp2/+
raCXWcUJAMDgKkQReQqb4y+eryQFlidd1CC/DHuS0l2rTVT9P4GOZLnhd45AK9jPiddJpXEuyvZX
MKqhbMtuDSpe4eRlVh+p00aoPJ+zx2FN4/oXrp86XA7EOzR7t+dTMcLs4WLFJN+0VKZGbKnifkDB
ds95pwWzFg1jjr2AHRYVL28SL9l1aY2nUtwIETVMfwPr4CvToK8CTB2Fd2VmINg2GSTix/blQGqP
Vcbla9AUBQBwgUUUT4t2qnL4nS3kKhUk1AgYgr9S97eDxQ7UEZgooUJWrIJZtZkF+/kXoBEFv59L
XgQ0ZrE9/IrzOlmRP2pkN61lYJ6sZ8HItmBjcFhf0jmQQay1V26aRJS4d6GcxBTs8qZy6ORFpy/q
oKnrjsBn04ej74LfrcGcGxwbT3vSV8v0oG1TTb09t1Qc2kxqeYPUd3A1/GMc+n+xn5Mx9iKFlA+2
6PSgaXbM7UhIfsurGcQBFbochx5ia56CiWIt8XbpoYymEMin7u+voVD0BIcUtDnM4SofhrjqjRqS
6eVDlGHvDyjrTasVWYqmzuvpO+z6wQQ2Q/4+WLozHotFtY5t0jbBrmdS/WLW03ZoaOt5IL5FSaFy
TKtp49mcJADjd8SQVh60wbMYA1gEshggbCzucXqaZynX93yrDUwPAK1oT9vIsQ+VZGQXi3OVquK0
Nrp1TYHezNenhKt5jTv6Uea5QdYCGgwoUcjtAriMKN0GFi3XBR/uotoCpqheccIKP2G6O7jKv0Z4
KkiV9Q6jqf0u/5UqLojvBRoK9rAAFLAhm0BEpLyo5/qWDNtnrB4ktnDlnKuwsP6ZoGS1R6N0u9jE
CR5RJhPCpPKDWKTTSgTRB9dizAHuFW36tGI+N25D8DDJHmAwDhH0nPwyW0WIAGqlxIs7BikLTr/E
WIVDDAsiFj0OAzwzumcMfY7zXJhDmehLSsZe4W5GhfIXRnLwrZCdwv7JECRPcLHBSkznUISEfqS9
HJ1OL30n2T8mc/u86pdSluBcO3MPZmfw8dmT719DL6HgqsH+NRXSRVCXmw258RCc0ujkA4CexLKb
ZaEcc3lnwKSvhpE3OZnllnnSmWg3AHIn54VyKFoKMdwu/sA+S0lnUJDSGIRmK7a5Dsi7xhU5LP3V
n8wv8D2/DQVQrx0XY4oC0OMJ0y1mzoymM1PwLe7c2phrZ9sLvi6a2J9xRuLNPy5jwqwEO99mDIM7
b34B302UhU02exWejP5DB8H9nX2/2UkL2Hl/Aqv+/h2q5on6Up88HequD+GCQZqWwBU8bMyiWnhB
/RQIgS9EUwmpsm84AiEtZDgxSqSoLL9njUcn392YZclH0q1BrRurbX8DMlBLG/DLbzUts3P3UuAK
+beDX8KG7E6icOoW2avZcfAs3sq9BFFPhdyu9RzLfLIrctyZxn1Z1ERdSQhPilotr8rexj6O5KP5
32/B8J8JlMCuTixtqdwvVhQq+aRPZxeYfl2iJU9VvCWttuq6wirdF0Wf1bEtHKth3uwJlafiBHIp
QUXmBwpUfHFSBrpAg5i/G+VvvjR63v8VqSChE84lyVaYvM5buni3owEboBtsFlf4LOCCoaCAXOHv
W0lZ7iHy+2106lsDA8OCNCUKUQGHravtl4WnEw/dCgI9gd/okQBaZ+WvOplEng6X/f8YvqmqM67h
hMgOcMeN8CZ4rXhRz6DwXx/wob3zBjXyMDEGtohC7pYhUNlCU0D/m7skwTyRZgrKN4w+qCLVXbmJ
lois8yW0oWhbS/js8FL9hT/puSTgH4W+uWRK2o+G1nfrJwIrEy/Hk8LW2z2yJFFckTwUyEfOIN9V
zLR6ikc4wBw48G4QC/rewK0GAPnDwGlDTKyQsD4sPtQGAyZwwLsBh0jv8rFiUiawKoTK1IQEbL3I
fl1wkGiakS3oX+ihBo5caQaOPB3anGMtqeonOlaCUrtozF0IBwMTzBE8feXXwEi+9fCQL5RZJ2os
mxjn809bbr34EvPnc2AN/1Jyn9fiqqR9a9OJvbb7QX4ZOaiMNhqlzVgPZmPlhME/EHMUbZx4wxLc
NMvw8tmN4O1TmJ1zXUJgbH7hS+KkDU/YvKDZMhk+Ho+lqUPVdSY66oy3Zsg565M6oPsZMHkvKlet
byernM+FW78VOaT0hEj9o/vr3uyx5twZZ2tYdVQvHavEZgMehsHjNGM1/2c9doxxGWBBhhNNeOwJ
iQUj4zqbAG9X7E6/c0ZPKEuYdGmTyA2Zu0Uls7s8ub7O9tQtNtSny2xECEULJBzAS+tboyWp0EvS
kjYz7Qtv0u2WGkqfc05zNUD4TpYXbdy6JzRxehGU8o/srP7Qi95JSvJUO98BuZxMmpCK9hwiWAwy
Kfj/EJ65dm28fpAKHqAxTgMova67XHgPtR1HxU+z4ilkhvv8oNW2ix7KuT1IpWY/A0kaiAdBrYyL
ySM9V8lZSNwKkAJJANFe9Z4gHIl+l0XNXpBXPCOqdl3oHyd96IxDq+4qkEzKh6K7xZakNxVsRrML
HgUHUX5jAnyWg87WNnTXWfTUZ7ThkPoLhCMBlkbmbVMRF5wgso/cf0kDDXbZ7yjZY0QzxxqWi65I
yKmZvAluEW3u9MFGTT2zhlmw7cfQBAVZTK3cKWVzgExwkOeMWdedbELaEJisnLVL1CwTuUo/c7Vz
2lHmh1g0a/zeyg/4rZ+WRxae5YavIZBkQIkM0bPEnkLU/PRbXN/2TtidnJpESfbS4+elEDCaxIpn
jjIXr720o7S1GApcblFDl7KNZOJmPF2g+bgOaSLlA95Z+5oAsCSYVd374WK4Y5tsSSfFkXZWQVLy
fX4m6yGcacJWfMrIJjAcRz1yl7Wc4Pd0noPTxJlgpZnXOG8ZuVX3NOzvfjT4pqItcDYNqNFZzsuW
kDiHcaCIbs7oUDY7hqU5Kc1f8Qjj/icbxHo2fdbeYy9/EXBr9M9ELXgRQtx6cBNbT8xH71JZ6zFY
rf67rlnpdOTniq8hMHpotHM1r63LPp2yvrq6loFmzL9qmaRqbUZQLpVAEvXGCLeiGPBlKO/Le//x
c/CxWy1vINmpJGZdRpEghPtlOwd9xfSLqtWLLxnXBJ1dPbLgOLCtBvID1jj7SoR0sLZYaoE1H3z6
kTlmbSb8K+OvQ6b5lkL5tTudNVqW2Eiu+0v/+JyvRJpGWxcyhaG+ufTR+9A1MACmOB5om+wE9/Zq
CvwpFhzGDGp7ffn7/p+x22WXTsktVbgzMaoeYd+yB7YuRbd66tJtscZ9zQZDguN7kV/nWO0e68Tt
tF0ITMibzujD+yezmRQ/alv2Xm1zvvaEtIAepWByYAcpTIMnR9ZHxkc9OO4agLnUIfn3wWdlp9Ws
2+HEuLTBRP4iCrz+URUi0LV3gBy1vPVZnjnG9PyqwsRXxHZFxwyIASMwG6EN2jPk3jE1PXZPlRU6
WWqNyd8JQxei/eq4NLjIGpT65zondob6EPuMDFzhI5qNzC8fu/hKK2LRJBlg4LW1Fs4TJSxme0QN
mLUMCOdXcw/t7eX57OwClzRTnA9eMUW+ZzN1AtZd+OSYDphm6y9Bgg6scJj+b1wr1yhgTx0ai6dA
ESgnXDzeWeUXpCdDRQtINgOhKTCRPk7EZlCWzhmJsLAFVm+cEK1MlslseAcSxx5YdgCxgFbSBy9g
QGwU63s3s68bG5lepEeYWZJNi0OhS/lYY1++lf69x71aSWup+yFuOvxEmMQ+FhpgthIX6G+Z5Oj5
SzJ6QcO+IlFItrLqiM9umuIW76Wa2JM0RGgLWhudxz9XcBaRQ3KfWhbIkT9fvzEJsPC4O0QJRxGu
K24hV7gH7v2LjcNpNH2zbINb3jOj50VDZHyDIWqYNtGbo9F7brRSOhQ5zO/yd45snF/HD8qCqeRV
7IQLmSBgOB5AULSJ0ZKCFqNN6wBHAou4+gsYh2fKAPJGEcJBIBZReqk13jmAsznwInwtypfi2pql
fx/aYDHN3b0Z0eOY7pRDQQA1VzFwUI0IpcLdY//2KFuYVcWepDC+taisggKFrMLOn6erAXyJZ89z
ltEApEIW4/LaVMps6Jc8pTR2BGEV9/PF8wSBc6iAFS+iJ5WFB8ZJTUs2F+PjmeDXICi1a739z8h3
d6Br43VomYHdo/jhZyhnDmf55JlbgY0Ji7ZPQtttEkO0AMX66Dm5edaHjtFkTPeCBCgDHe0ZXNA4
dmBaRUzpRbsXJYtEVSbUDkgt9xQ9xp5234EoS+tP82R5Hb+9FKDldv6mo2kY1NhhwbfO9JED1GtI
bOPvWKHrJ95NiZHil04EgVpbb9xwVvj+sPWarBusYdrPZpBAp5kl6HUSfiGCujDSpScwIGEBMY4d
1nmUHFjEQ8g8bnWrStmHQNO6SK+M6j7LOADpzMJU5rk7YIGjI3Wbz1U62tKbGaYE5TKipTY+NQdq
2MNz9VnpB7ry7qFepqitJ3O4KxUU5vr+VKqXpP2fd77pq+JrTe/lJ6XQxAEF7RDtNjxm+7GHWe/U
SSAW6EpHduF9lRbAIUq3JAvXm429HV4Ae8Cx4ALzeZC5yUrQIe4Aq2nKnTTncUa6apkNhcES80Tz
ctR7Gd5xiWQ5EWt1f4NKMEZSW2q+ns03sq5Zf/BoEIF3h4dEa6Nv2aqZu78uBU50fSZDAxPo3Yuk
aaMaKYhEn6OAP2r6bob+jG3gSxMdwWIJdE23ZdKm/nwXbKGXZKBPxwRztk4Sw6qZUuDgAkJEGl14
C7Cl2UWEKfwEu+EQ5lHbZwSNuzeAgyhPs9eFWH7QXMvwqcHaqjTDfzlb0cctyKgsGYUufqiiO1ZR
jD7GU36YUHxzPegIMIs1TS18tC+z6/OL6/sBFHPwmEzXG/rNYjEboWevfjybG9gIfUPoBJZdXxYm
Dio0oDl2Xy5S814L0AjTXoETLCA2Mipb5xqHazEj6mK+F/88WfDclDDT19i6MCYXATD1wM8JeSBq
Zwb43G4U8bGEgbQBM5yP6pd8XKROc3IeH1nl10Gkqdpl7ut4SLxvGgHEGYRYUEF3cm04NnfN2wOI
TPh3E+DtXECJQL012eA+jnbXZxHDWFnnAlILnWh4mjj6TCwh0SVk178glB3FFJg1h39VZ0239JqU
t/Kr20WPevXZc+otDDjQawNL7U3fg54QPE3J8Eaj9REnig63q2jHdsMdPAkoSHuLsZxd+X2ugqnc
4K4jyoP07qvBB0o3SUsyGLRRn88seIsMyATbxFgQcaWpKu3La3WQZSPbS0uCu8rDYB/C853kGJAP
qwaBS2kw0amJ6+co8ZkqyCBAYcr8NVwvkDETnUesMr1QldWmtsXe/JdFNc/3bpERIBNRGZmTAOq0
T2b1npUSwogXgBAnr4q3qeh7T/YHQa94D1IndgTXaS1fxK2BNTvPw5JplbE68kShmxoVN0J2bd72
64TGy9ezCQTYZaAh3ANkYSzxewZbHkpMpK0CUBLyzPJwS37Yjcuo33FNwHQHi8b8NHXihXSyHZrk
IfS0n0ZoJPGo8Ist3+8LL7/xXooLTMnCd9HoEc/uX9Gd6H5A3A9UpBIAlqlSV97g8/LCJhZiptaG
+wQ6jxhtkP460nRvKLeyyGVVVknDowHS2+KnXuAaaklq6t4ImcGSesBXnKkZl5bvBfrLZSPlAGh1
ijxoIZVQmdk7W+T3uZ6741wPFhkAXg0mieWVjAH/E96tANrk3uhSwNViij8hDv2PCqIj9KnyyMbG
3vfHTZFlAvdZ8vu6prL9xTS1NTe6y11VHfBceANsdSxwoRT1Z2XfhiRk3Rk/dJbt3JawIZ97Fvs6
Lt7B9CPceEwgeWCM1AJrjQVbH8iLjTFD0T02rCh2h8rXKF/9QLWtKmFm9biGpo2TxTA2/VttQdvK
riMM5DoVsLJ5kYw5fTxV5KhTtxezH4zKFYfLLJDPfamtbOMjoxhPOSenWzOBSdjJJS2DAOeAbv98
u2SchjFu4Ffd67N+qs60/bIO4qCbrh0JOTPgZ1Hl7DkcYNih6Z+lpDk/K+x/8WdzJ4C8udvIkNfb
tAANNH5LJnBNQwKg48CQS2iE8Z53LLY/MVOsucG2MmhOt+Co3NVKSzirfbLvXiK/w2gtZLUdRFd+
xuydFHQsZEl+dzdbld69cZNVNcgXM+/+13K3hLeOGPIGzFXfAd8iTCug1MjrR5DxrAt+xr0rQWKR
eC+GBROWx31VVjMErH7sTJO9HmZ1/fZTLkixPbWgprwOhOCogL3JLvmxvVbYyizmlhDUjmqsPX4H
9yP61CNkJaiHr/RMp6SHlTkzwd9buYurWBOFN1qIEYoGmHdOAkKVQKEuJn9LUVUnU8LYPZXeWCi7
IGMDY7Efmg9qrtK0DZ8Sk3IjyU0SI6eYPGGkEKjpI0tf2cuFPDSsghcH0ZK6kBmx71jCLWX/ok8d
g/73DBeHJSGCaQ+N/3LCZSPUK9HPKsV9NliItfqrSPjlTOhncD/cvvCXH726O7BwRp5W22zFid7p
2TUK261RBnjQcsMyw0IaqbFCnplKxRe0bfMA3788BNpZcOfp+t+s1Po218eus5XeM1a69NneKPjH
uCWAHZHi3gDPq3jiN3nxJq03QaHPFCLdbAdyNE8+ad7TZhjqHcl0CxCOJuJOrZ5inRWIvOFl54sb
x1TX8tCDcIJW+0383LhWWqW2jTBiJMGGq8Grmq51Gg7ibQNV6+/9CSffnldL3eDXuV9BWGhdc17N
CL85QsTgIBsOtiwNAMOb3vqdyL5RY/zRYKubcdKoJygf8YHTk7YMNmlBUmwgD8Q4RIaB8ZjB63u7
3O8YyaqXcKMnvAFQq9v8EhAJOmjwdqvWwiibRIbAwJdITcV0fFCgx+foEekir/naxkuAsAzd9lMI
GgtZEDIqcDSN7tyNvc5RNRZS++/M32DkdKnX14ZbJpU+Gir0X0rwmYtxOhCVAk/OMM/tedaB2DYd
RcnaBAkXUpJnzXMcH3RyWfbfymXArcnJXD6O4atczKKkZhbd4c9DFUy7gCGgTcM94ogsrwnkarm6
2vYG9AG+rrhi1VnDt+C9AY9PqwtZAUuPDEymfjHtDX47mH3dF5KTc2RyaQC5y6JhuamSK7BpvT/G
fxsodXuJpRQr4Z2rADzDzDYlwnf/gEs8A80AZh7I1Vw5GbgMRpaqDYBN5QYLkYQ3ZzR76N1YqHgU
o0KMWpncn93YvCYSPi9JUW/scoQUVi/2d7fZC4UuGh7I2gTkFozkLUUgzqoUpy6B6EDaJDqJMQPb
ILWkh+hp6NG4h48SbeCItOlmHPlRZTjA3PqlttNMrqydsd5CpKK2fZQwj2O+YUg6fwLlVDRJJSZe
in1DvF7oIVxW+u0jR1hC+n1ifu0K7oW8WWX1DxWbmhVccKORfT9ferao5pEet1b2jAbi6B9aitX9
zhqHkYeIVN/X5QreIcMxwuErazFfC42HmaWkmZoOCBt47M4U4QGomyo5bmwCQEmHr/xDBomeBu44
YpWaGCn/KH1ir77c/WoW/B1Q57ISHeTv2Dcf+CXhygcJdn2K2ziQCFDFo97DmtkrCk5zR/0Lwoq6
+WCBNjhZTK4luoPfHYNRO/Qo/0hyRipaZm1cKfxe258mu9qGHwGBZGFKlvHjVkuNGgBzolsivWII
nhqfLw2N54wzq6ia1QCg7wxrdV/1BuBEXHxC37UkJ0ISNvSeQ9LWqUfF4BwL+xztJQH45+RidAMM
V8VVox/j2V8Csc0x9x5m0uIttg21CE7jd3o3NtlwcCNAtBHxv99x6+Hc9hLWQEBl0N9PNovXhCqA
RP0EJSBHHRe8Ek8qoTuZpB6fV5wHGC4yN2cOxkIK/DEV3f8XxbIwJYrOtF+2eDbQBSv9DZ36Ysm4
zvHxE0cbGrHTHbJ2PIyDz2uHZDFtcjDaiP8PQbPKrg6/v5UPE5W1/sFPVASvxcSyb5fH2P16jUug
ggcZ8KwVBh7qNKHlXACF2NrmPgZC4Fro1Ta3nSFWL/QuEm6GyeGuyuU89/0x+UYA1kdygeTekySw
Gu1+rJNm3P4oeLOsYmnpSSMznESiF42coxJMFuoqgVmAuQscpwT8+ZnUwPkwmhZ6xm3dekLL1hYQ
r9DCpyee1dhgrPFWWLjxqNb7qcyoT0z/91qfKY5UcxC0I2iEl9E7rHcIrMjYDh0A6Usw/K5wZAZW
N7kjRMhyjr+0nbkY8hoUMri977TXf6YCTNMBCXMLp/b/RnYyojrtih8GpKagjnF60NEyJvW63PG3
hvEAj8xgRwyn7QFePm2Z8a3+/K768BdXny2+ktDTV47zVRIVHvyNuV2UChEQJj66RaREZ1gb8qye
ALGIRGvoj6KzqLXp7yzZJYlIzAOWNzYNmdw+AEpNA+ZvjOjo96frG23TdpjFngfpdZcuS+VfvsK+
0Z63dm6ypl56+EP1qvgzRFvjDy//W50PdN5jDsiQtZqBm9YiUs3K+q/5hs1Wrj9+pbgk5qlj0Fej
W64xko5aP1G4ysTpNmJvcwF3dvb/Syz3lZDq5K6n0ep9foAmi4dxQwI4FhJUhFF0JDNW+crUJmuQ
teJ9LTBSprjUCNtuxNtuzR4QAOh5eS0By1wI6BSxAsprQwlKs6bvIGgSWFcHKcRmZIWYsDYEl+6a
Ewo6cfdUX5ZkItokWS6G5Dz13IEKsVgWi1/rjcZlUUPILdB6r0cDS3MfodEJXNmYl57Ec7ce06Zo
Gc4JQJ9T2WnK9z6Rd9hQkgFpuA/MyyfC7Nw5Cpyi6fnQu0dQuDcj+Qn50LbpcOyfuEpgc+/5gyVi
UDXSfLBdDu1MV3CkCSAwgEyxPAE3qTR6G6s6mkWmlM7f/7+ChRq94GgeVkRPMbC8TYNqCpgTMjKB
iSUtMB72NhZdfkp52C6iLVbkrv9/Bh78ncZkXNvmqk5yo3uH3IOdmbO+TydggbaxAv4wbNGRVYLS
yZ76/QlOT5kTVJRp4cFD+IL4OGT24RBeEU3D/TJ8vhVF/jxdPgjZuM4ZNMGEEe2reGgyMzwEWPQq
hA6FGTZIasqD5oHMbPXHZGsqaOW+xmTpXA6ay3vpAm5deUccHmYQkC9CW12ibX8MQKbZjKIe9M+N
47ZnrLSb8JkN14o1dhArhS7vI6K+17czAy0naH26WvvC2i+iPh1gfgpU3sRK17B4htA2iawEjCCe
9Xkk9ruTfN69sU8ncj7yjwa/n61iwbn+1SeQuaNCDtNQ8+eQQG95j+T1zD11A0Ul4of/GC0ioqzU
tWPyrn4htzReeF2ek4TH+CQbeCUKi7BIiVxtcibH0jx+Td29r9r0PlN5+sjeSSgEphnwj7MvfIJZ
EpJyipDnftIIMMRGGKxauecgOkuZ9+ut6teIUb/aTfYzdRdGq6qG8xRR1wo8V6B0IOS6HnzYHYv8
qNyYk4yQmy+FTHEsua9k1u/636jEJcdIYE7y8bwZ7pOi+KTN7k894zIMeLtSiqcJMXkRJDJQP2E1
Ti9CFq4lTj2XsKI+9bCF7KblG1B3MY3Omn0Ci43Gx1VXHqfAJ8BCG5RQp4n6z8XnyYXc0OfUvLOR
qLkiSqePwchEldG4HtiVpTOMkXfl7C/NUHnOiuU1V1VbqA/hk74gsOxdtW9lOxXUkWQneI6+omgq
PJiQy+D59WrqFY3ddhgKE3cIbPPKeI7DenBbU1gXHNpgUXPxyxT+DzQ2Y7gik2rdLdgWY7WOAgjz
6oEYrNm2382FJdMtC9fSDZZF+T8E1zAkj8mry108tTPAuKi9oRvhhFwwlPXzVd4iv7flds3wozlz
tTClAwJepUL0sjBErJPt3tZyvoDeLCrHWnTtLhwDBhEq/bscdNTMzIMiFlmBO17DV7sF14UCMCat
rT+O+fvE5Jm2wVJNnxI9uxQyD9B0T9dIaGApEYV4tbic83/U5yzerIe/SaFmLJIENFUScmWDc1Cm
GHRiMHLsEMAV0MzSdFCCEJ5E9/j9X5Ip8dwuntmyibzgqX27cxKn7O8kgMq1p5wRM783JtxAy3WH
uAT8TDpXFaTsDMkAv+C9sNMwmzbamSExAq5QsOMeWk1srkQxhPxohMfdNRRyGZNAaycGC4yw+vz0
T+ApL6j/HvBE0SVP8FBwB1Ycub4Yx1wlwlHU7lady3P1GDJkU9+L+4z4akd0B48LoErD6rjXuQmh
8Oe2/sdgGorH5EjSbKAde+2ff6aZHeoARngzuow8jGIIEpmQuYz8Q7yzzWcuGAqdVVfchh0mHfCD
PSL6k6T3f2W0M86o5XUm+XmctPmdLvJiESGQnkOOOVTX4b7YVdGWobugf2/sQFiwwCe+ZqJZRAxm
4lJO2pnfhyIFlYXQ+bOBqQVkn5jsRFoWWIi3/dKXxY1ELJoeOID5z0tIioVdnyqzVJvr4MlltwCl
Z+cq/nCpEq4HL0B9wZ4u+9QbL+jD+CGMG5lUZAlz0yJshbgDEeCn47eKeDCaJXbU2qAjn+TMPyBc
J66vwsGLg4Kax82UKGUKQcTFCjsYrMI6XpWbYiU1/OeaqUmyVMMV7CUheSI28ctqBZs51tzLJsXf
2+CD+YOY6nQPhc4D2hP8AXxdIY4G+H0Rxuk6m7nmz5edmTIp9T7qIbSym9GwXXZPNuDJ6DU9NlJ4
qdCx7T93LyyHjL4hLsVsvDxpMGbLhLcBpqkDMLnXkSOpIIlBRiEaUJu9P+6wd+7gn+GEJPIr6MqK
vzrisPw3h6Js9Mpipqz+MafyzMJRRgNWPllDC3/3rIgsTViZV/sVTmm/PFwmGG2xYwQi9R+jUPyA
9GCrbGnJZQQGMw/83Pw8O4VxU0/T4sIv/6ez6Zw4VvMFxqe2sjeLT4aoq8QKxRqRXK7xNC0FnJgh
DqDRS1Sng+tRLP/qRdfRFE6zLQ19WuufY9wJocaW30lZ166WSDAsmyAgPpliGZl7KIMV461vFO+z
GZVRDEbS38wYoKxUsHqcgn8ucC6FYN/vb8FXzphLd5rKf/7CjoicU12MoP5r1ZtMKHRugMWQRXYD
QOrHexXM8OK28MnQCTTg19z2TSy1Y4G0Gb/4ir7FClXob3jpruFEtecBVi5xMsD3oVyjjtGXaP6Z
h+IY2tNhpxKhfG0y4cb/EerjL56OjLIO4sgVmNjRk54BgdWrU8GV3vlpuo2A2xvgf6mV2k1aas09
j8m2+BwUeHKwpm+RCyxuF3R6cEIDgCtcGZ/hl1a4wdcoPTlx6GWT1vM297v2+8sgeUifse+KDnor
Y7JG1nA9oUIEkERhq6pxRxq+6qqfhLWaDN3I+w4WZTVExtqyJVtgQmLKoCujRzVrBQ+1DYiL2QOE
KOGv+SYNbt0O1ekR10Zv2lmq8yaS8ldzBHidLGKEJjbxd6VNhhuAaJ1v2JLmKGYtw4eqq4225Pfx
1kTacAc836G0btJC4atb4zE4RE4rUYthnIxzDBvStCtYP90Sg3WDZ22CEJ0blVdzr+u4ba0jlW2/
PiKAnlkJsOvvlisrqBGjUHPWtOJpMHHsQr3p8ORIqFvjO7IWGbXH/852hX1D0j6wFFJGvL3Fkevt
EzIHzzAxPb6CTGVzSFFTK2zDBF+CRtz1iwOTeyg5UF4QVea7j9tiw/Fp4qEEV19OBgDEE1tWw38/
jpylGQdB/QjM9h5TijfNiY35BLg+yoSWYD1IIXzQtMpvl7QJHi7f53wl8czi24iZEehln5Kz45/h
ORH0CIWCNiLIBpk7gROCjlELj/+Zove3foQUIgaWT1FDAe3VhowNi4N1feGnkDkvnDaQsucMNHtH
AMPA+J/dvlTBph2c16pnDvN3PGf5wVOdrMNHhkMRMTtDkDKJGv01ZEAuQGzlBiEbQSpTE7t4cz+X
kGjdHnzks8UEGKh+5eJGDMLvyGjZ7XIqUs8EZCILmFFyPT6jJSc+EiKrzmH9OOnE4Y6+giTlUqdd
GYVcqLi91nVQpnr5+5TM+s+9ebGbWWJMOAcM+xlAcoPRfIWSVQUR3KbVzZhJJpINGA0rxDXBEDqz
rrqApQigP8a3aauAXxhhinvSfhV6BBYRLwaZZjLEYdy++v5m7IuDAXYtO1KoHUjcC8XI8p3ajOjs
LVGk7gze7UnGqBzClO+2HFBQgu09edCT2amtRrLHSYG+QxcJxyogybLbSkN+120jW+9kS8rFFS0C
nJIiFD0OHSWWp9MsRg/2AR1ahKlnLazMM9tnEUdicouogM2kPFJbOmzltVXQBGXDiKKGPEBIxJ8S
hgox+c71pz6y4Z2May1lVy0cCKp1dY8VX2ir/ZSUskc8Dcx1Lqaw3y+ouK5eqG27WbR2BJtKU9BG
i3DYVYq3du9DNAULoCxhQng17tLHPT+PUldiz9LSbDeN7JCKaWwN5XXFWA1/cSOqf53V1sF/eHoy
K0jvDFonGIRYXTwCysG7YQ8oQnaP1QP3Qqcv8WvKDKqnMtPwd2cz56EuQM8X7UH0e0Vgx02zwfQ3
lP5fcNTCrSSiYY7kJaMueQZoCvplvQdS4Qwa24tsdu3kl4ch2WlwMxmikzES/MuFOHG6DS/K/G0D
/KYiGGywg5G1JE1Mcp0nqu0oXYvYM+nQG8EZrohhSAOwWuXrBzx7N+A2lLilBdZrGeOywlc5e4Qe
QlQ+4a2Lct/BWn1ECBUFE+mp5AsHfaz1uQu5giO5RoHnmjg1jvBqCB3ptJCuajii6y9hAhSNw8Bf
ZO3MeJAqUeWSkQ/Y/46ZKrqTPV8u0X+tk/4+4kEtnlV/ivw5pniZ0p05j+kQDjFe1zaM/+kt8HLk
nLqNI8R0XNOoI4qco86O7s5fPXAoSkmY1SFLO0QOTtudCagjQtjV7zWZeMhX2r856TR6sCP3iNPT
CQis28dNVgzeJmqp4IwkEKq/2YJsDdqvvqB6DI+pB2ELvkYoFHuz3DHkVeXUUT8ztpWUrQE9j9Tj
1rlgLZ78x8MR0d0+U2rmci0R2zStven46zGYK5xNsqDKPtiReMbyYYNMiRygj68IAEVu0rVwQnF0
b+vcwMN3cexZbDK2AmdQXH1Qr1dTHQ7Si0d/WVn5t9mIY4qSR8boCmUfa1XBpj7E2Lz0yskzBNq7
MIr8VrpNM3Dq41rMDIWJXmo6FCDNpq6aec7auie9wLwcB440uT9DGTMjrYuOtNElL4Y9R99Oncfj
PjICMvBv0BV2oxPZ1WW14TD7F2crxbbzKYD19KNSG4EEhd1OS6U5ZW/1TpTJJ7k1ges/tXyYvio/
pgG7UMErYLftmFj+erUkd6yqwnqKYstPq+Kg+R5YgB/clhdE2Wizycqzqp3uPnutKAeNOx6rrCxS
39axN7lvF/Vk2T4iLL7O41hQngPc1RUuh0Q8n03T9cn88RR9V/BtomQXlK2tXCyVkEcecMx36QNF
NC4MosQ9KZzCEhm0n5ISfwNNldTr6lGoW4BHCuM1VOIenM/0rJj/BYUtgisrvRR7FkyT7Z68pI5o
za9kam1NPaTGOcIxlEEPi4K3U/yGaBa4w4e0l33EqOPYRM3SpH58Vyv78aAH2W9fqtL67UojNDha
1NP1DikwvBxi5x8b6AlUgKKOl/WcIz5UClHsmK1FhAqXywEsdSb3UrWw2+GVz/xvU0u1fIBVbkJL
uRxRNWJowRHfQdx5oL5N/KHxUJacYz1YfyvqC5F8aQZyqQaHZ1VYeTaCJImcKb7LWljFLn6HvDDV
Q41JdDJfHc/fXXYxNK0VE4wuB2X1x3iR3no7yqc2YrS9pnh+ZhiTGiuQJiMWWLngje5d4WW8eqkn
3WfW+oQZ32iFwReCEpjZxDj1bLUXsbWtzjPKw4UOS6pYXfs8IAbDasGqBLj9mzihCId8ABZt9Jfs
RUDSrhLUyTw2JYrGFhGaHoWFX2s7mf2M9EZetkUPs6AwWJI2UIchtxeBfYJbPPtTfEA4MbmmBds/
NtcU9LNgAgyOWi9z4z5rgPfnULSud2hOypfP1NuWL7e7xaLslKDp6pd8pWfSeLgCCLPO79qWfPLl
+Dg3NAh5aoGEDeriKy5/LQ7CskJ9xBFAenhxhnS6cYA3L/Ul4Wfs0OHWvkxws+S7aNtJzgts2Xvf
7ZVomen5FTuxhOpHCjDvGIKODbrcEHp7VqEEzdooDVvv+DTDY5QnNFlzpxA9NngaImED731VNm+C
gvrHVLqfgtI3SBp5UyKo0FoR6YORxPLb85GEV4aOKofud9yAOp7uhRQODwdvxk0P9V/KiGgDzpWf
bS+/CrVnjbiZn9XcqksxeNDnqNlwUBpgJo/dah6yZvvf4ebI52EaVNHP3y/IH6p1AApuiSUirAUB
dmL9heX2PaQPEycjqXAoRY9t1XKDKYbOZo7XrppN5vGUz+lqFTcat9MAAKP3+f8O45+0mvK7NtI2
g4fT0/eOawhrm4kEGjpdmnRhzzAMw9Tu9/QXNldVITj58q8rX5bWXrm2OuMLvpnUfJaR0qjxskTe
WnnE/nJWM2clyHI73G8MrE0cPxy+KTH7AcUtF0MJRXTYaO22EhsvegkdgE339kUkkg6ygsU5ObA3
uEBWu6tRFPTsiEjIoI1ezjKAkl9jFsXxIs2FVszuZdMAFvRKSsPPrbtohbdBKhenIC2Xk7vFlarg
P8CPBJNj/9u9xA1BJ0NOgY5VP+OmMpHMnjBiXP5eJmyd1Fix/zF9wtT+hlcshgRCDxH7ush1t91u
spqRs8bj/pyzaHtu2tQKchGZwM5iGrKl1wMvWpewba9MLz5s/Z+RTY3v5vB4TwSHRve6n1itX6yA
16q0w4uX3c8HGDFKCK4h0dRqdsG8deT7x63YU4o4r/O+s5jA5XnHqm+g3LuozT5MJRVOwJ1Po/5U
V5JfGama5pm96virKbX98OqiqH3O+R9anh93Jhd+S8Orh0/YV4ZQgXdo8vIpTqmYRQntxA4A88Ni
79akOi6nh4N4gyZ9qS5uPzXKgPyiKer6Dw0dygKGWzvnb4FSgARpvqmDnNL0AOtvZ/vlTtz9iYlt
lEf/AQvP4gS7q+D2e77hIiIHgWPmvM6U3SLDknCOvKc3OEasmoC1As/CeC++O1rhA63HzQag2aWF
lIntGSj7IpbjVhKJm3hTkrS1ZgzJnMg3f3tYVlTw0OWKHDUv8Hk7Jc7d5p1FvkpiFqf4OKwCbbNi
7UPJ4MfJJmOQWPIBMzbc22Rr6qVLS0EvbWHKBGrN3xmTPjouE89WurvEFLco52+NAvxC/0W7JFIQ
mt3adj3wOpXdDSGlDAo2WK6IhY3TLDRjs8TgfDH/qf3+azd1o/SQ7VsuHLv1HVumHKi0aBZxGYPE
mLAQnM5UldTcciOCNXWw7tEqnRXTyBdnqSsmd+tB19h7uyw/IVAePCgCG9JMkM4Nu7dfBqpFlIHx
MxtZlRCbmTcSjGtHKnXtLXCujyxb0QQ4g1UYocHBEb15lJbXF8goqvkkta9z4YMot4UwGVZmTZO5
geET6oD0Akub4tVis37lbIC3yMQh+JuD8oU29yVnEclFDvkc1JL4bw8S/wR7dbDFaRu5Hrqpa161
XW86PMmprRQC0mqSOb/GGS8rx8ssk9tMX6hW7c0Ad72mBeWNT5lXMp8/5T5ZlVw1ctBasbPQYi2Q
BX0/AbSkonM0Rvps8SaourxYHdksjmWmeuXgIINkRtnM7KMYPyKfR4UaWkl1s18RGIPY0tSLSabD
82c6SBeMT5InT9r4gLZO7hQABlsfcrDlwlJwb35OLQy8PRQ1ywmuSPvd8xEDj02ZjcXPBtSpg0h0
Wmb5k7AH8/BnCQ5yT9OBLFfEAl6CMaS9FqOaYnHkiGxSlc8r+v+6mN3lGmNh3+HNY5kd44rhHN6h
aDA6aZEmmRfdqNIjU0+j5GhYpLym9k0m8IHIabJZ9QTRQ37fe+7N7w2Ni6p2PHOsPKcLKkcWrWM9
WsNRaH1klWdntYVZkG+raME1HaTpeV6eNSBsGKeuaAd5VFb5aBsld3fgIW6Li14CF6UTqcv+NA2e
SvgDsEE6fql7prr1tpalu4EIojes5w+7SI9Mx/U5q0UAsEMQj2cZzEWvINKSR5AFv0X/Qoaob1EU
3leBYPG/l7JyoeRAvJ1JzSC5D9i8NNmUgLsT8wTFLereDjXWkkG1ja6BURCNh+nQyENFb6ojck6Q
coy6rlwqZBDtPvdvcTueNjhw/4UjDPKM5zwYrWyUDzWBKf71mNHnvthoGYIdymPxijbMpgryk797
b2Nn9QFiq6guWnT7Lq/vfLrTcJN/TVvOzBNt2h12pQJIL6T+F098XmzhBxKvCO38iyb+FVisEFAr
Bl1F+R8J0XDqcQR+CkRFzqcqMrvl/5B1gU8JruTvYa0vqM6A3zI8egjNU7otpDbGmtc896/ieM7O
lvjRVDKWOphz4LjxcRnl+YNHfw2PGHRB7kA75LL7vplL7uFVQ2FA1zpfe3uw9jd+SPkvO8DcUetn
qTmY6NxSHpWROqrus4I/+y9E2E7wSHiAFSmFdUEd0gUUp+SFYWgTYCBU8WqRcit0zN4XkNJoTj9d
8oXUw5yTeqrS1LHz5V/wtTRkfFJkf0h5puQe/QG2unUh7qNsnjMOag3tyTmIul1O7rrjiPTLqhP5
isFa9AkrB6kA+NkMRgePADgMANOFGxpLtjr5Dko07X66wYy+lYPh/sLQOvy8EHl5rPP71iQcgu+T
6WLNPE8snMkWopJ/0MehTE0JY+29117Md/uWkSRRpGueFGAlLA+qhBFIwRHtWtUws0WA6TBchz5s
0ovhFRpL9rHmjcXkGhrcyUS1KTb2AQB+Nt3dZNeyM+JMuaazoVcldaeO+zDTTnUu3AOvWCr1fywV
HZGtTQnyArHR3TVCTk7Q3TLpgpR8V4i5zgPvVLRktRAsIvN792T9uY8V/wTEDlb7cQmdsQW5OeP/
fWyLX4KJR8mMn/AEnCgykjlaIJAF97POP1IcpsmNfsiQ7/7HJ/avbDjX6cXcRcKLxYqRPkZyL96u
X2M/wmWvtLhpqYtA1vM4I8lDv/WP6FfGEqplZ4vwmlJBSwgPLMTizus842iFYLG35ntN2HOC0gcE
jU+PqvnHqtCSe6BDUIbN8CinNxrGlx+o17389rdxRl/446gMjw0App5iqaLcrH4ZFpR2Jl6So5sF
5XSaDeyIIlIyCpEoSvmMZy3PTTdMR5CK+jL/e2S5CDdd7izBW9g0CMbIP+/mc+e6hs5vvzuiofiW
X+9C7qhQARGJedyoUP8TFPzSMo0IX395DoehcuG/ryxMJTZY717lu7eoP78gybg9FQlFo56jqAS4
i7/bOnTqDciDJwoif6OkzcyQ0DfldNAiKrRPkf9wZDXjmBv5cEa9LhA031iSNfW8tdzXgtdoQPxs
nHyhTCcosfthUZMbr+OYSZFH30+81AwNc6GLSnmIiAyqebIggAjyqDsuUzDkJCifeeiz5ZOJV1Qe
zTv4HBqVbvRKfl4T2xkT+DdI/lFBwD5mHacEB8DBEu/Obe2bEnn7Fbi1lEGv/8OmfJiI/cVlAtQz
dhQVeaXUot4QC9IqPlK70cODkmegm2OLWMbbBGlsf5gKGfdIKV7YSBzKG2zTo8Kdx6s0jFxGn0oy
XNM/pNhgekRHXfZDJkLCEqUltcOT0FewX7VVpz3zhz+4X3MQHumekjuxheXrTovGEQWMUZNDwrlT
72pSNpUtLbH+hYWIrLkZh7JhSDSATO2b8OLSG79hzQft1wsj7PtPBcZcRQMKh1NTwLWeV4hRcdvb
ZMv0kMt8hQicJkdHE62gL0jmKdq1wbA7jIT7JWiugrcCvhpl9ge96XSGzJwiKsR+MUfDGZfPGpok
CQBSWaIIPHsqUrH4ril0L2kp9ZHEaq4o/ApCnEzr5oNzKyf7+rrCu6Ve5cPxqBEE39Ff7iU/bf8a
7IpYpdZssiIGhR+6boFxwr98xBSRtNBYT51MGU0S1dpWY6nZ2uHJ8tsdmFsiQd8/2h4ofO/G2bwN
lQhIlEBPpaj1+uQwjgm16VpG8X2qCb+CzBXX362PjU4qFJobZSxYQIg+D6HX7RMjT8asEFyhMtNh
5rCyVSjbDeKOlke6En9xwK1O56LLcGJWA84nndlrFalEv6JDmihTFGGtg02kDTy6RTUNsOK9Hhrn
ShIzxaBrVPHhG3u0MUUbrOVX0sFmp41vJrcOcx7p51vc2wsrjYZnjdTuZtuihA5jzCjOvNZVybHe
PEEfXuTnRrFB+CQEPJKtrHCB+Znq+RA1uEEVJfUeSUrEYgsygefTBLUdVD5xlYkgZMVSxwvWNrSL
i/MWQtPHxIN92Hj1CPck/nW4lop2RbTIa1oPtDcgN9Hg0zBABjRSgr9/4QI06Ln1CumhFvyV/ybM
rPG+uVRDoE/DvSiUinjQyANTB/cNneTWkeOSwLz1lAzlCyerTUM061p3B6u/bDvnC0I4Rp3OSqkQ
Z9JRD4DAXS/ZbVamOu+vW9bmJ/rEhHuY164X1TtTs2QOWt5ZVfIoi8JA79D0Y7Y2An4wB624TBvw
+YODRYNax8IFBRADrAFR/TuaGKjvTQmD5E9NPSutv+VyBjyloQwc0BNKeRcZ6kqbEAAvFWDFu1/4
hRddHFPQ/6eUGxV7JDy1SAJHG1bySEt/2F8j3OMZoRhkhhWQC8+rCRWxR5ySPDZkF7VGwMavq/E3
geODl3AWT+SoVWNItud8CK+IDNMxbqnGjzJE7OmUZh4ebFHWl70uH4EnH4Oi0Fy3rXQxsuig2qlA
9mBs7iowbovriMYQtNa7c6d7nm9VWKzk/JA+DDWBh+4hjXOXb1G1s5k9Z4XXlTI1tD8zSzFINLsQ
/dFki3pOBmmgioeA1AJi7FbkIjc3jcJdZV9ji2D6DKOitWyCcuQC4CeD4+30E15BA720YXla4Nu1
D2duqWv0sV5gk7HM3E7DPz8QlHvBC8w+4UcWt5wqb8LI/zXO+dJs52qfUz4JUi56Omf3io2viE4n
cayy2N5ggXAssFlXD59+UNCbIzlA5Tse0t7a0IgvzFXjrUVZDSAr4mQ/mGUxj6Zft3aqJjIyCjJm
prcXlW6AFhaFOAW1KLlnRLC4JORExnYtsnegbG7TMluU4UFSBB+CpC7E8/QiB5jdcHaq6TLjFt2a
z3KjabOf424afPXD5/vuwqGr0wIPqSqK1TRKx48SD1B+elXKwourv6pKkHK/cUm5hSR4cy0q2PoS
3kvGna2Xd5EAYbhl4Dfem74p1LiC7U/JCZ3aGfVVWKrvXgd2TdZlIMUOPcGi0F8ms5LEReMfrMOr
I6wxAM3DFPbh/ELG6/MEJgX69tE73OMAgwZuk4XQQx9nvraT5hQxx6Ub+X+dRpD1VIiijnjp9ozb
smFXE6JxX7C4K0bc16G5IWAPV6vNyKNFDOoA3SwEb2pm2wRSjL7Rp3he9Hn9o3O0/ocBjqxG3jKp
Y8grblPMNEHOzYbAbUbuwKHYMp3vRC2ri0hTwHtjRqB2csIUm2oesviY8x6Y6cRuuP4oAICZQxve
amw8iVQF/rKNl1yWc8ThVAVh4Sl5l7K9J8A37EuVzewqZQ27odmJkX9TfWgn22uaBOFijzjtbUrJ
p0invUJ09kaPfI6lzFluYpux//oXr6A0lPZf1/7owm8WT6V+UL2fd1FBsq/dSx9vrPH1NN/BpvkJ
8ELiVPxEb8trsL7yY2ql1/jioUJRDxSYiGqlcCWfwPqR/YndMq3HwQ9qZWM4y8WXWOM+DPFAn/XH
DQkbbp8VwSXwrBI4S6GS8RQyU/z4Ie4RX+S2RDpKKdjlTS7Z0KO1yDDnqdpyzP6qmUFtEwbC3Iwp
FxCIWfn+GYvUFZQvxR6dQNvOuBfL4+l9Z5mWxLe9Wt6PWUMEnDGY6CubMeuNphtSdKu1SdJXOlV/
8ilqVmxYldapS8GJbwPimv1Owgk81mJNg3pEP1/3MYKERhKampmK4gW0Lkyo/dKw+GfJozR5bdSs
W9G5LtPoLjxTN3RokIK9G7SbkGUhZoBlBfYcAkk2AHBKuqEFmJcr7N/+prpiiUdYy7yfOEETtp06
WG56yG5O8isHJ+g67kLAPsseBLaYL0LNqbTBgwt/j2a8JwTQOMAbx+m/FXoSLo7qunVVUEgL8e7n
1yil1/hnBRBmTJxvPPk9XMyQZ/xFfJE1WV2NmATBfNXJ8q85zxxKg1nRfmX2LLaDxO3HBWpvYehN
nQuLRi+PBTKbKbqC2GfiOS2LORxk9d0Ih5ezy8shscq3xT3JDrjEVgK79PxJcLf1ldGlY0S4I1MX
aDu2SPHxdNVHRPoF4zphK2jSct0CM9pSaAzZYRh2PuYlAITxFUdTwUJhHWPiBXrwSMdUKubWwhJ4
yBQ26hGFpMwEIkFx61Skjw5EH0HWtteW/F+2Nsm103L9XeB1KwohiDcfvKAX8JO73hbl8Wa/mxQf
Pn7wYjxSy63U7wehZ4c8t6VPw4uD4qdQ0FUw08DVlpiq9EFIXorzM2HLp951/UabxPtStO6KKHdF
PxngGthN/O8Oggn4oSYeN1MJzk3mmxkEszt5fOUGdXFBqhqg8QPWHJy91k9VICfcMN8CkXNemENc
eJ9OBSLJSSZXP/Awi+aFc9GqN7qCE4GTC/Q25Fhe6p9pHSbHH6U9X+Ua5FG2oHEaQLPgytQBpGXY
mDjaqe0HUi6RFih+I0ntCP7ueEmrmjUuhSqNB7hZwH3FNkckVhUrQgAidm6PdELPM8evEdlMANu+
5t3ZQ0+8hnJk5DrBF8Ip4QwG/dwuZb2ZFYez5AUFvgt4LBCR4UcpfOvpcjGFxGVcYP35omrwoY2f
nFfnY6d4YHGAWcwFaYNhFh5s8yBQ4XKJOKl2hnZzuYegrjECcXU45ENvG4u4kAIYQUIpb02O6zVU
Z7mGAlYBumlgiDY7MuPC5rIqq51oAQW7i6BiZ+uawUsrYwCoJ9yYd08OeMfT0woeSO4M9j1iihJt
IW9YrWhpPpbA+xi9fKHiTJeAuuTGEDdWFt07Tn/JHIuCRglKoQF73kTii6ZKmxm1wPM5/BHeB/5w
ua4k35+l++LbaKREfYWpsEp1cnVnTMBOJ1MT0OCazO0Tu8n4jCNaTrqtlCtSH85lbze4t5nsLN8F
sjLLUpBliFubLsomk/DcaByQUwtybJzsWTDv2/+F70h4MqFOZ4Pfb0lBEjtlroM7age6ZJa+ZYHA
HE3L/S8CZBn4aU6EoMfEP/WHP4IA9P+RNZpcOAOmNTC6Bp/Gqh0MIPcadcU1TMEawl5CJ3JtiaEF
3Eom5Ivy7qnITHIk6lq15b7LGnfzOAnC1NYGEVWfU7G6zFyKeqHJ4xwNx6E95M1DidK3FkSgql0u
ajKZ/olTrmuhnTg9eue8Xy/3UaZ8xeRZkiR8fHTNt7KqOPZTEEd3DDeByLbVPCyiU4k8wkBst5dq
Pk0XODVls1+uesd6uSQ58AECVCVYy/S5AkX14vAWOZK7kYNPzICHKAHdV7TSFUwDDz6KgFjy1J5q
P/GfRlPtr/4X54HNHKEtwy9F2FlvtIo21fsiLQ8v4mCTgzqVKO7IsLTCH7K0XMjHmI53lsO0Ja2v
N3gmjt9qyzqU56lChZWb/G5sP1kUshxhNHM4m2JOVpDwtXynHZJ7nveHIeXP9/YimOvunvRlEKK/
0avWfOoonFlLDAQfpqut8qTo1D/EHZ48QqGRq4kUhFSea0AEc7NhrIoGWEM/UVjzH2/AxXcF5xsb
oEiB1IMxq5CXHgDo+KU0kZKnfZRJ4qjT7iEeSX5avnwpKN+pOgNTOI8QY9Kg4Wu06bgI9Z4Zfatm
dT8Hq7v1v/4dK2SKMaQuROMACX1OMV+trz1DKHkkOJPm33R2A6dj6GNQOSOZoMwN1KHaczwuYCtB
v8zUbz3ufN7nnAB7Hdei6Xwm2Epec0i+fLze87Z8pZhBK7ZYf5hz32K5+t1Brp5nh7s9hoVfCJw5
hJDUNaS6HGqyrihdW6N1ap+25mgmjyPZPWriNlHzwaIv7jXtQKTCI9ELyIamzDM6c2N+K6trWf5Z
mLiDc7uPB4EB2+SIqOH4LlScvL+Y3JRdkRi4xlS8Epp04QWheZYvH5RP/ofhiji5s/vRNZYdE3Di
efWWd8oi20xyR3hMvBMg/mRwmxHLH6tBQh0vfG9+WQhVJJGJEFLnNL7msnZdOh2HJfLsUNDWVMea
5LsQQ5Ib2oQ71C0USIzTw34/P9amp+cm34/LFK+hG4/Aqun8itJM7p0NS0gIA0TZ43oeuc4tHe3Z
JYwToBZV1m8m6Za1OeXwO2hHIunyH0B0PlCI5gl5z2a+EL1h5VBCJBbaLe6G9EjoEpf2O/Fvn9At
bfznK2WqnFB2lDdOBxI9pmeK8uxKaB88MTKIKXmI7v26uEYV06uhBPnvBVxXWfPZSjwLDJewSfqt
JzTWMtT25kE5FoWUGkWEsVDztMXBqLt1jayg/D1EYG46pOJ9lMhKiIrOaOMGQkdEFO/uq800LgqL
bXtb5iwq2iA2ZVD2VywljlhWQ1bYyibFcAVRSSey3se5VRheG2PDg/K8rE0uaAGcjoaScIoHbiVR
N7gy3ekZk3HVYkClo18MjWB+euQGobaAZu9ev0fK5zjknw+1g7O2NyFsunumSGWSz75gQ82w3est
yq8PKD3NkmfA6GydnBqt/0X20j7cUHbJfDzeOjSssz7jdJgoKgbt9h7BzUSmxF1uIUvl6/NhaV2E
mi2DcD74/a1TfmnxRRj+25om7I+PBxg+srH4qV/fpdz7prmLF56+xeX9ujpd9AfMy2UFpx1OFOpn
P9Ky8Gfpr5daJdS9vgLjL98T9fba5RGnVl85eQuZuGlrP400st16ZVOyD6LgzVXyMJsTAGSejhqN
q80PQN3X8US1rSZh4SNoAFHz8FumaAk6uGg0AOFXbeku8flNN857fkaOjISq2z88NUVxb710BRE7
xuLXX5ZX0/LpJmW/iRGOtNuqCw9HWxblhpA/Os4QZ3GFzFWj5RlSbepW1zsKO3NuBqQEFIUVmEKG
CcXhZf+usoVRJ5TwHLqXCpWBbIG6yHeFbDTRg+tw7YRiMJyZicidti+NgoeJg8IbGAG7uz3qcZM3
5fvg8VHQgFPQwWYEU1xU2QM+WYXBhKKRzJWNvtMb3A1jrpnB5h9HHI6Fv/M06qwq8WB9BmS8+nIa
D+AdlqgtyCvZCD5WF0fP35m7lPjCgBo+yEzohlz0mA5K+nvfkYMaaKRohk0ow3A1MxHTLg3YOxDB
jnPaIJZitkSz6IbBp6IqD1dg5z2yR/liTpa+Z36bd61WEVnb8hgE7AD95Iwvv+IbYTIKrNJUGxJ1
RDoPEMHBLM1VuOtEM91VLxPMlF6zeTTWSBeHq1H8mypipQcLHfTFfQE8denQDg3LF7QYWdbNsjBy
trP99uuE+8fV0xcako485kj97KhwKXFfZTBZkpJewMFj/ZgTQtkpV5cjm86+zRowZbWSehIC0C8p
DieTiSurrJr936VIlN/71pSukoacLWUhZgc0aAWgYUC2rrqsfVsTtrQWwS0KX4qEG4XZivQOjen9
vUTaqh0qbDA2NTnty+XYBZ0ucuYP0eJLov8u2ABa/3fWQeHppS0Zbi/CYSULcs1PF/x2Ldk4E+yC
V1KUO1+Ghb4hESVfJZGHk3ea51LRgcfoJ2tuY1zPPPU4IpSB6TyrPBrytKdjoOPHzc6y+aU2hZLp
udzzBsT9pqLrMgrfukC2MqX7/qYz+Ga2RkcC9b6Owpm+GPTdFYxWzTcq8QHlvzl2XVxRvEjfzkFP
X5I/InH3UZ8JHVuVwcJ+K177OKWbvyDyVRqbtsgwScTFpnKkvWSaWRd26Nw9q0R3qXFRm+5mmUIG
/DULBXP6MdFiXUYM51moFWzgH4rDhh0JOd6u4RdaufyywI1zZLtf4m+H8sNqC4cnKgv3L7bg2TZg
YXvR/br/CG7RBVq1PhJYDjhfxqcSuy/wo+mqGjULtH0wHHuduggvrQxgdLsuP2bnN0gxgNi/zmcX
7F3N1MPmPp9/1O9AjlK0gHZJofYjh5ufCQz8VwkGOTyvsaRpl7Pcp9o8joAoKfGa+3G3iLwNueLD
tJtPywd51hnzKAsNXUIB+iS1IQZnn59GmCwBmaRV3PdtcTg2Gzi58SS/rEACEDN5pr4UxMC/7yQm
gUQxNNpCyw+cGgQi+EpVtij43wbOQBgu9NrWxFCRW3AizQjdWfgip2U+jBjLVFZziLJmS6cVLB2n
oP2aAOBdMwRPxjYTR4TdTzpiXPSeM+qOzSXH+pXAA5GCSAuruzicjnay4rr+kw93Bteyxu7qzmSP
BxOle90zeutALxEBBgvauvkugqQsReEtEOsPvfspAftf1YpQgeoT2uxRP4KmuiJBXMbvKxae0Esp
GI76wfD3XAUe5FJNFbOV22gIddJO4LTR4X9eXv7MIZmnvU84PaZ4V5+gfyEjk4oEMlcZXuJ9ldQR
mLiBra5fkP2eWbvpUfLHEs4m7ny6k0mKAeP1NHiBd2RrVtT8J9G/50/ov4BtX2RyXxbwpJ5kCVFl
MpJQSBo9ESsCXBiIeSvklvomS38OnpWEN3HRKqKKSxyi6T4VcTi9alBBA7qWp8dezmPZKXk7yRYa
N4mcJ/cRkz4ZHWtts4m4vIzs6k9lS1wsmgKISBiQObdfLINuFIQk0n1IqQ+meDic9/Qxt+MslHl6
enb0Nk3Fl2jKmUTuTGtWOnhlQoWmp5YOYtY2ew7bzpa4m6ymgWs5glk4QdbjcHRVwu1DZsdH1+s8
vmKjhKItwv7Fqfe0G47ceykLGDz8EG5Jz7dZQJGoCCA872O+cWQCAGI8Qm0JW8Z6NGy1bfAwL1bf
JdwL9/6ReXHgw44m77tkmVeNuF7Vlvyooi4LCqq8ty7fbnm+kXeWeDCXbKsNCMODvm6Z7L5loCda
3bFkDtab0RdyA4w5Ct86EXAlZ9IhptDYNr7iaJZQp2a7GX3THCy84c8SblMgj/s4N2uvIINbFsBm
4IixQCA7v/LmmnS6D/dqS1xCUaFU/ehzPmPljU3tSZam2GriuZhol5Uv+eI5dxVnCZH7gYEe7bf9
g/axO03XesEjkMUt6suM9Rh6+hdJG0WGMKy42irWtyv3XSJtIlFTi12J09d2aKXyzgJasVAxb4Mi
/HccjN+mA2Huwzj4rdsHDR3Y13JLWzITjgVin/IIwKrjojwrWLZQr3wU1EkTEixllfSlkFs9VpEy
X4nvrfgsJoi3MqoSU5VAO9dgd0h2qYWTvGyQIbXeC/ZStMoClBS2HnNp8bye+wDBLlOvkCpodzCk
kPPx70swne1DODmr/yj/JkEc/bgCGFmTtBOeDUovJEQVM7te8vFMMtuN33HKRWS42c9w7PLJaCuo
DgEh363+9nPGwGmmaV0RewmZezj9ve8eX4ezAMH/H7RDtFZDa0PMzEGGScC6ahNRcs28W0ZQAy7b
lrU76RdMFhAQFvaPwPdFYEeUBZwqttPudr/uwfjROLC6DT2RuAvISy6ZgfGbVlGeBXVYJIBiH9cA
fx7gWqbK19lILyQi2Ak8C2FL0G7B8tGaR9Hk1oCIGkQ3WsPeVTUqR9k0DPBQRvUqb0b2viRIj7cY
kpxihQtwEd5phu/21wPtI7MoPVkpIdQ1iN3lVb55lEmuDB/zmM7aVmKsddpsFzO3gfQGphuA6ADc
8RuHJnt/LdO7PyvqIUL+4t+4fLAgGrydicNZ2pNTLsJSCqiPq7fzYtQt/zNDcN6cGc8SVXcA5UeO
ls0CNDd8lT1PbJKw65uyf5XcQnbsusEgBhH2K3td77e6Csj7CO61qMXFAkqjubJKekqI+rl+oVzM
SP6JDdpFv8Cd0X+Vjcp70xeQ9HPTqBHMr7DzifvmjsPK+MZ4LCGTad7oxPCRscnBVWFOMYXrSScK
q6OnS38GbrXYhfmf3TWPEt3AnbJ1RYBeupmMtE5VzBoyO+xIsantJ8hdYBYjuMTPFZLXqXoGiUl7
790La6nKy8pnD5cPhMGe1vg16z1EqZDTZx1WwAJhSXEIHWYakvwMEwqey6dsLBMPUJ+cqWCnZuS0
FU+REU3MA8SottTRQ2yH4982wM9KFgCDxiLYys0sSmzkP9QWCOqrsPVuGgzCld/3xDzM/5iAF263
O9FUYbjMbkOx3tCYKku6bmeylZqJTodw9ccBMYKVDj0PZbnXDHSPkPjt1fSVOSavT586utG2RF4/
bQlymoZl5Bybl2apx3Py6/Co20ua0/rdc7Yv6fOtr8Ox3pB5yvZSowFQ0oEG4v0jBJMWChbXbEko
nxx95JL4fBk+dBafttnIeCzhO0xdrvrOF+SPZ3+g6U7J2Iq2uaO6SsuhR8CCsDCynLLPUb3Y+MZV
57qCK53/UqTuZUeoskzl48VkdUYeZH95LAiLxL/YsSKNSatnG0BDMUtSW7TaYrRQ03ZPy2JKNqO+
ni6LxFD6S4gDsVe+vJHBQbsTdPDzwVmOWydHfZWcOlTc6f8GvVaCjXU39p7WfeMsbuqS6yPMsDYU
CDJdcPqjw8znIPhbTVgiwMFLye2dwyRoQZi9/Hm+9fKvB+iFb/Il40JeJa3XyGPTmRpZI13VkPb2
zBd6Q4It7bi+yF3LVdlK81e3K4uRFizLvgxjh+KUuljlkKPqZuwRZy1OFTawsPg75OHdJeFjqwLT
jlRNpHeR/DBY4XFEyHLDBaDMNRv4dij3zNbvu3uqhD0FGyEh+xlOp527TIV6gSyXPfSDEOmDZkUu
Tqln83oL5A4RmsJuGL85dZoGnnbySAWVz/bRb+Lb10U8UXjVWiI1XmuEPdz+Dtk1qvjaBEta2TFP
In2Hw6EiQkF83QLDFHq/CkA6zzbRjux1WISHeEJ2hhfE2/xEZtj+CQ3Epr1lM3xnBOFYEejgmyls
Xd/hdWiVbWY4tWEAyHUClTtop6sBJ1w3JZ+hH5GvR2WxkeB2UZTiRkoP88MmW0l6U/Af3AemR5gc
XpGHsMYL8/jwe8Lb8EpVKJHTZwVLYP/nmgC7EwsrB4YH0Th9dlr60ZHFJudpGdUUlLCuKsuk7rJa
b68TUAeVb2+7N7GUy5NSaoJqku+ghJNRFWkJVzJgIn4OETBrQFEGRcndsFyxGF/2Nhn93iWC+hU0
QHcTgr7wG8h3k+lbAKVuho87lIqHbzsXiK8wU9FXk3O+NHoC0oIuIvl9fO6G/4wVdWcbaH5RQLLX
r5rdaHrhpm8B1WbNZmLrTuTQAXTnBZwOhYJmTTzVcT9gmXQtXqt+DlDIG1tmGlp4QRUKTjQHm7Lk
jFfpfF8IpEsZ82A7GIR9ULdtJKzDe2yz42s0+nZFKVKn1Ue2ulNVtHIWojolRq0EQe7Oh7Zk9vzD
ApTzgmLTBd14ckw89MJg4heUWdaGqNRUcPR1/Rey0dT8Lavp65NlfSBq3DqG1IDGxSNzi8n8VGpV
l0pj29TiiLvvUyoorhO/WRN76Qnz3hoWCbSbonrkPM8LFMKf2DupSOQJ/np/vSe0r7JVKH9JoKnG
0FMHbVd8HWep3ukYMgnD4+cNgmlUjG0YBbaI6CYb7MLN2QdwtLuXVbriSAjI2Cvpr7oKveEc9+j2
4Agbejc8fO++oqFZj4uWAhSa1emBdebLniaq20YdFtK8bs4Y6p9NTxu5C2+mDmZ47HCmdHoHkC/S
gcQxHvTQroZS2a0DsMm7mYc5BxnI+oNPftK5aGngp6tlCuUcT2cVjOLz3YbY0FM7fEsDFbkaV6Hr
1eY/Vy9vuVvhr58uREpMOa9J4SUdf8FATdGLOy47c56t4Rvt50jpD8wPRAxDULcOY4OHcFYmdi/T
iBv6mqgt4mYjxWTSwijMV0b04j1BuQk/kDmdmmS1VzEa6G2uARqn35nKwDfeCyQm+BeTReA5efxV
tcU2aNP7Ep9FYINRBOVCEmfh5iswdpnLLjci5BqF6xcjyFcuG03x0Agl+tZrXr/szsfidEE06aJJ
TA8DZUvJlwyS/nP6USjFX81NbQkha1mUlNtX4kxF2tRKzahhZI2xFtk9gqr/kHvckAJUugXIHojR
A3MVGT9uoBoSRzFA6VCMzCVYcKoiLsPhEEGCKhDP4gpdJTBpZoeNW5f3dz0wV40HiVsSsChy9wVw
tGCpVbTssZCGRz1BNR95pauDUHGDGSp2Z3IGsTwCiyBW65jQ/3J4y5TMvpQ5SaaxkeSDpqNXDOlI
tjLPFi5MsXXBqeEBPLCVj1s2VgDvnwN3opAIXhMXBnHe3aJRmr9ueytVLsNdhPoRK0wa2PnjwR3t
YgT2UZALYATK6184raPv7jvszp7/BWhOZoEHEtHfuVuLxEWgrz1ghTXtOAayLg8iA0PXI8pgMu49
lSj/iE8wOBIvnjLHI6Db9Fqtf7e6uXMh7i5CI7rCaIhuue/c8fPeUbS25PE/fQzGNBxijMA1wOOv
TbiydnGq9NVt329yTQjb+WtEbvc8IPDuyIsSa+3nfVeVCURRp8+DY4HXOT4wDhuumiP3f0QE1OhH
c4yEiphgbWcHXzNd0BIbmySAcayXyje4rXVT6hg/GwHPLSZozSYMC9Xe5b3sYivrfJ1DhRVgqFPZ
pW+EDjC0RIzCY6slt0aJym/Wcf5+As5+lhdXArJ9Cyue1SF3iy3ewMphVI7y9jfRDcxpohLIk2x5
M9RO5jzM5W6Yhr954hpJncUzPCss/6y7Si4l0rUw8yfmBOqGu2PqvOF/TZYuxXDoNmvregHE0cLh
ml7D7LfMU+KIe6A3dEPiItMcAxTjtbbOlPAoHKxQo+6WIiH2LAJ1KQoPOING//Ir+53FSKJxjfIx
F4em/OwNQMevIVdkqybFpMgi0Q5ZjK2yFULwC2DcU/mg7iQCt1PvI7wQAhmeRRnBqIetz6WBc61p
9wxrTNyeXijfG8BoxZUTg6rWNhK7moPkQA010j8P0zW/v+z6OO5Zzwmqb61V++xZO1B2UGIJUjIC
ab9WHKD4jhBl+ViRmg6xIUWBN9EQVMGUU45rx+afJaL/bd2D4K4IVMYkodVc9u1VMnrXPQbQc5zV
D+rhZ5uRK4dfUzd4JgoBrrU73vWHUB+V05I5bLTS8fRSf//rDdrmS2QLk9wvoRTzu9/L0Oqnyimo
1cdvi6gg3wueQgMJTiyKSoEEr4x/Fvsv4LfzhsxxkVC0YOuwBZt7An0DAEVqDB1P0LwRoVdAp9ib
EY8w3RLrG0H7PFcm5AJgeMQMvjYXNDt7v5uGOH2m5M/Zw/9ipg8Ygv2k1oeR8Tc7UabMn3QG6r52
+6BP9P+ApGefgLrNl/EZOdK2qGbvVkAv3BbLZ7FsbHx0rhMV+N0XY8LQYVl8Z4VxOnci4rCl2oTK
ig4PV7EAQCBNmSSRMCEfKkx469euNisxT0cuaKf1WBAaBoGTrGO0j9+QQ4AgBucl0inGgDMDRyZf
bhCau+5uX448yj+jcfkD5jeUJgo/yx6fY6QAIjrivcnD8YE3DR5LtnzEcZ1q0bgGKGuFuWIOGTbq
URPTy+GBK+fK0voertDvlxFoMVWEPOfS1zNVnEQfknc6LZtLEpJ3a0T0fslGfdysUJKqe8uDxh1H
PGZWNQ5lBQwhQ5d4izN9mQ1ZXIoUbb/CrUH7poY2ZrVsci5/M5sxudmzOjjLlZbOvTIwxPIywA3f
MQllZ73yxu02ZCnTC7qx5600O6/dWKrDBG3kMachShX+5XCUxTgOshr15ws7pO0y8BuVGMYJY6J0
DW6HHXuzIeLsymmbP9jHIvSg/UAshqSWC6LAnbLkY5zHRvJ5Ol76Ke0D/z+nofCwuO5OlLLG27m5
897+ef3ZX2SuT8LXGAiNn+bPM3iHjfN3W+tneYwg68tC5+CucECh972wetJgdh+Pa2k5zrNnj9XU
1x0y91UrIr+3zbqbnJ/qEQyuR5ZNlkr73aFt/om6lgBo8hkZ74WfzONIkp30cI2A9aZ4VmmBQpHE
2Tq6CKwLUFUrbNqS6wYHcL1b0I6klQZBMX91mp3hhhnNLaw2mxVnlwVgmwWLzUjm9zcLTq+oS/tk
XOJwNk+5LPWUZUBIEWbXkxTJbBQPukFhrqACfW9qtZmmnJLIgRWMmTwYlO+QQkkprL4ItmxOZ8+2
cwDnRKKvxUn2BnPy94UZsGqNAfA40KCZGUF74bP6NF4YAp6dj1u20UHlJxsNI2uIQikWLsPViTMe
vKBvHBzvnMN43FtSi8oTYv+Sxqjy4y9kbt/PL64viOu0TE0/GnTYHYUzydSL1Do7AV7pK4GCMDPz
GsfD3h8HwBDHsblDp2x1trzOvxTAMGsjIqFz0oYd5Qm5v2Fjwz4F5LZN0DMFUyVcQ/HbWhd2+OgI
2XcM1xQ+ItmFjLHFFCt8xmR3pTRXnE3mDqZuVK5dpd3qlILw86IpAkl8mJvBHs9Z4ccVubCXzYIV
nFk9VKJ7elonUmOgqowT4rYRRuvKZGY8T9l3QKJpwGqvZY1GaCpqxSG5RgVD2NpZ2L0AqNdz5+rR
PWIRw/xWVEeHdsFGiHQAO0srTg6/ZpOJNeCgxuSVFbSLs5wabUwZmCKrg4w44RK20+HN4Ye53RAy
2SGhip4JIpkvfAT1muAtOUa6bksiV1xOL99jL39UHzRCS3payLcwKa3jxhkimvHU/TXmAC6lGI0H
gYyoos4MMzgFOfQe3Tyr9fOxbkU4p4GDiahp/wgxZ6ouyX+VTu57Qc2u/k+se5Nd5goNax0JIAtf
wXn+KgAakAc2ia+TNmJvbZSFl+PVdS9M4nUEvg28H3o5fkHDf5JXD6zfu64yp2ONuntz663phevg
7vhlNVJFNcXknhVk0/o3lojKY03DvntNN0FCca/Qzac9iBSzvMxpFfHBLFsHXtXA64f7nEJ24yn3
7EqavtWSzVTdYSURt1vjsZsn2LAkjkTtwHQjFXUAhagUiYw1fsUbKsNwp+ObujRSOD0Q7x9MTCZq
ENMzyzTZzkZchwTgZb+0xPazZTZtniF/FMvnkStx5ebihy0R3bwoJEs6/3WHo12fZSPR4Vsoc7Lw
sMdPnazlN2OAPLulJiECVj1tcO/b7n2wAFe2rnXa3zbMlI+YHx5sTQRFcgN5JyEtmilLFtBMpd8m
TESNbNGmJI5gys/b2DNVECzihSzIXjqndXn0nKRBb27ZhD2rk5pns/yYa+65iqQzXvNTMs+Fa3QT
hY8LpDIEYSdvPeFeTGl1Pn8ZX714cSpnnXAKN4bmZmVpcv92GrbbAJJedcwJqWS7lMGAfMjhU7/F
WdCoVbYaqyA2io9SAp9qmbcclTFo+FyjNB2kwHbh/XcupXSSMA2H+/k74RpFRU4spc+bE2syiWiE
Ae9CkpeEUF+OnVV7wycwNBIDmxAbC68PU9/9mYcePTGm5AJpWZWSUecwy2nQ5ALKHEdZOSxHw7wy
pdVFVVLfuzIocV58FooIhKhR0VNvSbnOKxA6/25KA6QNR5nyZhMODUShtIurZWLGdGGonn1dTZL/
Zlt66XFvFt1bB4adEtMa1JqNNvkFJNCXwb2eqnX44+LF4bAoeki/PCqd5hVlJnjaq4KrClvFy+8N
VJ6WBTym/VLB2bqMGEIsi2/MBIXv1hWq6v6q/Ibw8/JIfmyl9eywfImxw8Jf4cjELJnrRG9+3YBJ
IksYuAfEoh4uqqN7qosmteRcEyahPvsiRQLg+3UT4oyb65as+6H8bB8ZHIdxQ3Nz5qgpe/M0+ENV
dhd1qysQ6R+dfZH5jxqbHpCcaxNdosZCC7qZVBpl5txj0CN5NCvtZ78ZaewGYp73xgHZzEQC4VWd
0/Xg8mzJsIFKkDLvbXAC+djuYPd8+JIjgSXm5P0vUB/jq9K7iqCL+cBi7dwVUgfSUrDaERLjw6vj
lsMOqWF57U5QYc64fWJqsJK9bnR81cormZPrOGfPh5fbeE9XTrkZl6P+ePkE7hbpRT/QH8/v++hH
H3YCw7tlGSzqGPo+ME5o8w1jkFUoS3TnE0Xgqi1Xsa4TDzPxKMNr+B7GZK1vx2D810yidkUmcNs8
pnLd0Fwh2utBVumc8leZj6qBAct8dplZLaUMNGsVP+83fSJI4i49d5I1PC2eiDBMsu/B6YSF4tsN
FAprcXXVpmVDbszwEk+yEnt4L0bE44PmcNbWQa6W/RGF3HsDoSmqFyseHzwqmpVPhlRtPXOuRWq5
1FGYK6EeupzcO0DWcRhMVDyNpvGt/CkbO+jl5lar9MqD4vIQHiebZsD/r1ZAeWD07ovWqTFmx1UU
A1bUVkicnesEVQsjGf+nOXTpLp3brWlBU2x9e9MfEeWUI9miUy5OLWObgjncGlf9eQIDV1T5k1SZ
Q/iSqsKFuFxfr6qpeuafW8TUQH5T09u9Oy2IflB131cY3yxZ4aXu9H3y3pVgxFbaTTgfs4GbtS7S
oSLFHroqEzBLLmVIox29cPZQCuIEgdGNr5UaZ5JwMuQNHndVmb9zFRpszQ1WrJlTkZkjiyvgVOs5
lBK9ol4pEsf6iGncdOcXyDCtke4R0K6RPFUdVVaNIhFgUwXsNzkvMV/jeSuTpSK0O6JnNqNIEx9H
9W8a5WcrRGlM399t2GIDFczAyajEUGuTfnGE/sshlGUttOjRSxwroh28yuH3A5WPLdzrUzL/0244
716mAc1QE2aMj8ALmhwJ76DzEm6zzJGUksoqdylHquxiYjLFjbFAlUgLAIZFzssPjrppJ13bx4lr
Qooyo0E9q1KU8r9Z+FcXvIa37N+ZIQKiGaYJfyaFi9T3vfMQuV0CqBEH6v/yxXqvgAFJVkLmTsyR
3DqnGs7CRkkGkCnX/5q+BLQp3Aqs0KjHKU3ybe41OGtzDaZRHQ2glCg07DAMEMNVVXLLIGzrxP3k
K1RyLLOnQgpucJfoWml0g15fzLyyHoMnsLrZej05ywIhQolkcYKvu5R7WZBjFODgdGMaQdYt+EL5
z0AFz8XoOq1UH7amDjAQ12+HmjPnQ4hRsN8rWqrHTAU5mTpA0oHMb1AHhxVUvf2PGhsfoMo4jg8Q
hK0BvMWy258NmIG+hkGNc5tGzu19PTsqJbdOS2eQfk8LHlk1mvd8U2VOdE2bcnQTPLDVdovu5ISl
EOD11J8LihOAzWsydXCRRQE5whrODgaLuVOIH8iCaWiYK86Qz/i4Obax64Ruy42js+e1Y8UhG3Xs
/0COCTlSTDY/Bz5LQAVpowlGoIrrD2z1PnK9p7vDJFjPX9KhrEgA6BuhNHEynB33f8mI0CeFymB5
vutmtA4LuXIW+wur7/rh5mkR9dcsVSKd2P4WMgVWY1anoCpxGuLhlvwXnWpHMVRsSJEVCBrhcs9a
fFcSs+6NfDs/wavSV8/kTmmj95mZEMolSLjZ1ju2NswTn/ZumVka3WEj7s+07iAJ5uU+KqMA+cnK
NZMnqXjLJK9pZlYf4z3M9DILHdHV4onW99n0DkeC6lJcEZ+mvq75MmhetUba0Mm/SQmANiiDa5EX
6V23LFwWvUPV4pwMWYW2g1ODUUoiOyJVPoM+CuTyvo5p34G84zUgz481dBQjqr8QIB+l/LMta30m
jYbXow7s/wgWpd3ZxAloHrpEKQtp9AbrBwWziUQ04VzW8NKWkv85i935zeOPx6n7MXd9ECh87hAq
6+007OANF34culPciDf1fy6wfh99AgU2YOgcisxgu3XJK27XavrCgP/XEQH3wl/Jv8gN9hI9g53d
cNx2RzhV18YkMOFh41NiI6rreq/Sw9Aw1XPXiJ2HLiT7817CJ584YtNbwxbWUEioCfowtxKgoxc6
XSoikCavyCR3adVZSEXN1whwV0DLJ57g4PRjKEpPGVHT5AaA3a7FtyBgZSdQ3NiMo4+NS2iyIc5s
JePOqMMvqN/Oyy1GssHBueM87RXh1Mjjr3XY8k1RZaYaX3Kq+DLdDVBlV4+iow0v9TM/Upq5sISi
Mt2l+YY1GSfD8/cyl5OFVrTCb5bKp7EaABK4lHisc8c8C7cMl/22yZFZbPTsX4ZorcD8HD+6Lnvh
oz188Wkd1rnMWB+jkGADjFjefPugDZ9gqt2hjjSYd18i3xieWGWoMlZOvi5s0qiXT+vnRoHb5iUv
MzRCYjyGFzqu+92j/vhm+Z+lUb/0O83uRaKjbv8Rotm+jWtNAD7QUZy/9VbK4TcfW+00akspoOT3
Is7NLAVT9GNDK3tYHaKn1d+7Vd8o5LzTQsoVsFyaVHaGz3YB38pnYCJXuSB2JqTYZ37mueKzy6kZ
vFw4p1eiOc+l3zGy3ebZdicYL3lE6TVslRmbdRLs69K/r1RAqP4cSi7crm1+pGNOxSJBUScZBZn8
MTFdSMHdUTR+bvMw1XgaMJCP2l4f6SpgMiBShFdg3XnYuZ80DanjvD6/cAm9VpNHHNJrYi9qgZDd
AzLa3NNCNV5P49ggRb+X5Chv9/EXuCk37lWMXB9OaDHSZFqk40SMyQ+KSx9/mVWSweyHqsrpSSgi
75FtYibmnd3FwdawzOxKSIT+GmicVfOCTz/6vtCuaRTT6mSs0UxN6c7Q6xb27y6YHvvNpfP8IkAv
XySkrUbZEPrQJqLyvZOR54cYmy96mFCFx5Nw8PVWJIltZ9K25D2tNemr1S0pYcl/3e+Afgzm82nV
0umcv+JooBes4MgDw2suldw9uo5i0dTbgv8szWyBrCPBClSmTZJDqcXxr+iIk6r46j2ZbNX29yhU
MOIgNnK4j3PoZLf3YSLeAllWfX6uLJlmWo4S1gNzLFXOhSfz1O8JsSNuZBMZ1iOsgQgMOYtIoDXT
ZrKjmt9wkwhRb1E+mFncW7WcUN2FCbZzFItSfOr4RaBwe+Irr4TD9I5hdUa0gHRW3W09BADtD6M+
0Xi85jcwG1HwTf5WkSfHlrchwWNszY4BDNG0T7Gj3daK2+BIT/UELJXhwrrb/OXVX0AmZTocg8/Y
nj4f4HZQrvZwAceJAohbk3D5OM6Sy+8NmJ8okv441ByZJAU5l8A7h37YrrqCahBlRtbhY/heIrgv
TyhGhfE9JjJ+jSCaWZsKoyzVAS0xcoFezJW0TOb6DFEurozZJr8OuBq8wB3V3kKuEGCsMLymbQE6
TW9hYQW6SpHltyoGAQPH9aIMqRPm1chzMJ/HoJ6XWoBOqGtoqaLQWFLi1F5s7rjOSvk6ldfM96f9
RfubLPkFe6dNdZA/UKmijZdl2wKegpbrS2cJs4CEiWCNKP0GSUzOskKJ641Gq17mC3mJLkC2m2op
4hWERU0laQLLgXVtr0FyQtksA003dVlYPoyrIeo/VOO8XMBdEPvhG2B4gEJm2s25D46/Brk9+f6G
fnt2zw7MKdllx+Si5VSSOK6fsaZjFgF2qCXdZSjKRzeFKN8Lenynk0AtEUDj0LyzK6Ey3NRS/ixG
1gTGBRV4ThLAFfkC7Tv3FEExnc9w8Uf97kJK8gd1JpSybBx4d6Zro2PQ3czaKI9Cw73+y2mhp5XF
hPwYR1/W9BGD3qnpkhwPTcJ+Ob43jGlbf0MoG90DLYG8Y8nPMCKu3xxucn8+jo4s5gFnvKjyS62S
Al60gNeCPkG87cPsTUwT7PKjyMonGRhLV45MTkSnSwuLAlJU5epusmUzl68G9qfZLxoIEUBQIj1M
nXintfS5MTis7+HYxbijAMTVViT90lcW0VUVTdcE8n1RCN99CB/EU4y0u2ezjBjC18mDBd21jiJq
9fF1p+/IPMKo/pzY+GW2or6LAON/o72cD0SJRa2IvKMSc2iinI4irAPx12CoBZzYYLfkdLgd9Z9F
2XGCizagXLbLIHSf8Lm7yw8aPvalkqtPBwEpNCGmk25AM/m+t1biYdDr9ha8ZM2iryls4oQfCCY+
R17818KmYpMkHiZfUJuDXg1kEnu8jIQQ7ipFkQF7fhggY1DBdWWfC82hZUBRP3fkTJkdpFwf0rnA
KluztkioUqluGmNYNOKrrvWkCWnPLNGo+NauoQLRlwyKGqGloEuBiO+UJc+xIR1ejbRaJXU5WDyI
/mRjYCfxXXO4F+ELVosabGJqHG+TSpB7/F1HolmAKPd/tfhLHFpuLLTfKbLlrndHHSgkWSAw+obZ
mEt2lFqwW7Fi8Kmph/BW65xfSjFFTrlQcE4H0A+U45nurcSKr0yvGHOGj5L5eucHmZHHBVm26UHj
XFfVZrkKYlbN/vts1ms3neFDPlXc3Ozy2rjz3cRoXz86K/m3f4QyR5brFSe5TvOe92/cjqYef34b
0KmGs/skGLIlF1hCg+J9dNPXKC3lah4YAAEEbBE54gjmtoqRDbFCcoL2cFg+kOn/MFJDNEc394ZX
StK4fKncIEgy2+zXFVnLLGK9/EKTUo4O3pq+gxWxtu67vHVbdGqgyrnl9KiTi7udVmzaVw9lI+cu
QxKc4uCKt1v/1TfgvMUjPL+yYF9dtj+52PqKmxuHjbEZBTHMMO+1K2NFH7WbFsxYbTViJPIbglpn
B/yFzCYMBMttbo1RQTyQ9igdgkbKhy5lPMD6eLnoFw68AlBWCMFl+2DhocG5tZ7PJXRiORawGKx2
9kOqJlN7EuvNl+l12plMVHUxBu0kbnSM8r8lXi1f2RgG1eqNZgiEayDWt8OJ9Hq6mX7W0CQSlV4z
q07ckqARmSUCOa3M2x3ngHVvYSoZWyjybsTMeifGLNLn+cmUaCVlb7Q5cxl9kx21YwlycTxEJh7z
iDvgMON9cIYXcog2rVPL8gWpabJXxYOOqoPu23bo184KOu7+8+Q+xVUTZbqYmiq1WMhbQ5v12gbD
b+kLVL+DHqr+USQMSbuw2q5FwB3SAZ9HcqTlQeopb0RNwyXi7gMoB3u4KzPmf5DWt9blF2qtabrZ
iQjLpKcKl5AK+LSGf8pxOFSKAci6aIEAAhKU3bkNDzfGIsDHWzQW+1KZIBNWQBPmY5ts+5WPcjMH
N+n2x6C5dZ/OrbKbYp9UmOX7rsNV0+8gkLhqcsCi37xM09ti0LovBFX3ySkpIi7eq+cHsx/iP6wx
p3Ci71UjJUCgESHijt36Vre7ojoDtBIu69lWWv8RYXrEcxkYAm5p8NIgxBiJWzsrUz0F8+JcjwBO
ijxvKIWsi4f8fIqzGpyhDdsjIUHsuIYJwu2ffaaATyo8n5X3xIvgv3Zwwl/ZkF1NzPQhEd4hVm37
qzQcirSnETMnTpet2flfr2whN9eeKirO70uINHe71aUH3YsOzpsn82fsfV8X+StdTrEYkEKjx15D
mksmMeC2kZuSL7UOevWq8SmiuGfhb/tOeNzswl2JUvkJZzdFB12Uty9nxfLcSwmm/NiuedyZ2pQp
AkZ7MCfvFrGHfUi6WLJ4FigVzeSVxXOys9+9GOn2JZe+TRjGk6f5rxmJdRcvppcewGaV4JG5+5lR
832IQ+5BO8saQv/IzFuS39uoqWCRc+AneECdsMLLf7ZbbllRhDoWlx7b/Gkkxjx+b8kPekDZXy9A
SU7wCVocUq0la77qVvXKRGQSfXUCUypywz8PxwZ7Lu2AauV7q/AwsSBvvqgbBdwvwHfaKwn4J/r+
lzVbu2IniU4tgnQej7C7AUKWUj80DxFPpqcwyHaCBF07+0Rmy6Q7mg4Ewd3DKLhoQ3Cf4u7Abqad
l2oh6sYOeAJ02GkGx/99akJ/y4J2LHkVOzM8BWiE7Pv4pGPuOp8mGLmH0bhAEPBGO/F1cQoYF4kD
ygjh012qM2ROWi9EA0uymDfOVeNum5Y9D4WJ8EZUh/st6ByNentVgIALlQ6EHNFBuAyoLPGiUW23
dVhmKTnEWKqle71V8oMVHeE4Wdyekq3S4XTvGMuLdL8AWs5ZVevO0EYkR9XG+Fx5axZYauaNHcbY
LZo7FMbe3SsAkryaLpFKiwCwlwiNvrj4SGKxLOy6QNO11YNpX5gU6UQGW6n0OUxTT5tJbo5UeYz+
nFRHZ8B2ZV7zDYhVDl20e+xH4ncxTJAUa1L/LTvVsCt3Myi0uwdowcQB14aE8fDM6QAD58+YZW7A
AoV4IlH5Z0wc0RtNxBMb/pkPzyuCIRUvAzQgT1LV1xDblUrDgpxlXyPdruL5Tp47aX2xHRoDM8YX
1C7pruFh3E8gtOh8jKKdCZoiH8wOWPHYP3iFVPMBxh5AcCeQNrgIApR7WPssKaWlIsqTAea1KPtx
KgLi3OSz9QRq6HwDJw8sCURncUakz3M6pEviMVzF07WQYUkBH5iG/VBASSf0aE2hsYZMSdu8d/d0
GNguLNyb2asWu3VW4y8V/CuMdUIDUKehCT/WVvCSgue3ydQ2bOcgg7Irz7UgBvJE7h7WdAeSJRIE
qBdOD6ewcWRHnsCTNr5V2B6ZroAH8sjlAydpNP2aFrRCo4uEeDFXITd4I/Unt83OhVU+U/ZioOIL
zUwLeaU8qUKfVoQ7ZA1N4mGRcEfoBLG7XIjCtne5PTBfj5nX9qCcACn/hGHH2Jsciy0GjTqJwHY6
skJUYdJOUaRyFBKylU0swywP/bfiPPX+g9rjGtCBlsXL2L7P/DVu/WOryp9SSoUFIuCCzgLuKfPa
6+zVTKj1tDl9E3eYw3mu4pDbRB+1gvs5s8BN5SC1y6gplY1IssT+fi2PyEPlJM7/NsuuDxT/PyL8
rSP2jYR8gnVqHw2RKwIX6iM/aZdw/cyGzqr6hXuRPfYWcdC2IVqzeFKXjjhHkQVqCd1KlUu4ZPJF
hBf5gc+hHl0Aic86pM8+ncM5Ru8OwCE57QRJ6q65ynXS0kuGmGeo6NNsVOwn/B8vL5B3ExXieZcU
FvJBTeSqnwPwQLAGHH51TIhek5A1UIf6jhJVhvMCXL6Yzz9MXLixZ4gbgA76Iqv49F34jnZKJ5Xx
GmmeqDlJ6Z1AUXHcdTP9CyUewTnu+WwMFUpgVKn37V8WliOV78DP/NhvffWtI5xnc3QXb2l7czuI
x/2vKwbu69dF1WPCun5g1nhAAgdjJp6UD+u9FWlgRBi3hsn+SajpYcUG4NqYvLA7kCUJbAjyWU5T
Ci67Kmm4ZHw1lT16JEzgvGJvWDoT3ltZ6327iVq1KWfD4BFulwZh64M6nTJTf8WkIYc0aC1zwUUb
Kqpp0LlV1vkbsPOJKIkWDi+rQ58XEhqeKtKdvVzITU8rxPqLF183xl5veryhy1pfxrPzPxxuVDMw
HBYvl88FzCTMhN3nj+XxorH8Eec11ShhmZnrchaffF/g9KSowsXRDsgjmfcSO2YJrfDP/597GBDD
quMPbIHoo7CfxVbFN/HTXMlE7K8LcFhozKXtOVZfdZwQkHwebwP9q1pEmeKUy1X4j61K3EZvqBFp
JJOmdkwl8RWy4ZsASMVdB3G+WjkXWcorgzQwRIoMuHO5864M14rzJTXZ2n+YNac8xWKgtj3xlncW
+xVl17gs8AGBn/eCeqlhmYylWQoKgMSLwN0wVcAW6xe9AOQM0ZiEilyMch55ai4a1hJr2H95pEtk
aavtmvAcEdphqjbSJFpvB1MxVd2ogqa+BJseO4l7DKSjeT54Wed737EMLxfYt9Eqn0WxPEcZsaKm
Gckq55DTEQiFPyRvXuilF9zNdq/UCmN0G31iDtgVW/LJY2hGh1yhzy7VfIn9Bw+2f1sxvSfqM42g
QoDFwp3VBxxlvxmrpM7AuUCYfOo7rcvsIc8pKEcU+4q8RAqsS4WcWnK788XMouu76ZKLE06U0/Mk
nE6CS86Qmny+HoEVhX46zZCsHRCd6SLN57GF9teyDka4sNkncx1k3hJKW87IjDgGeWmS6/DcPVzl
WF5Veixg6DNgX5MDlO4bJbHPrU4Xb+9Hs/zQp35jSTzWTGcVTrxLnlfJpsNAdiWmNOaAUO2A74oL
B7WrKlMcnvm28Psi9g9rAJPlVpu238RfoSbOLi62CHpa2eI4ScZcxB0mhosshEaa/TPR7aUxkUs5
axI+AKgdF9OxT9ttsYsFRXghzCdm94nh5/kRSm8fIBwZaAbgBHAn5SwMIeSWB/KXg7rbwi1khugt
jdHkvUQzUI+J64b5BQPI5+HOZpWlWV1jGX1emDXZXAuZ0QPBEoRvDNWayU0TEa+s4d4W+DtQYzPZ
KbGc5BtAEDdfacqz2pyJYOt/e41W7MPI/MQv3Yf9ybr/t24eeesuz7nWaKOaqGH8p/AsxCw3saLY
RACGVIj5ptTKopPnsX88Le+yHq0/jX0e3xscuOtUlb3RHr/dxE+oju68zQsbzkc7uJ7DdihlvTJx
njljcH6Sjjjv7QvuBwmuGduAT6CgbzjSvw8laQAVeHklnaSnvsDJeYD3gu6FgS6YzbpYUAntAQMf
fjSFcFx7mI8DjNWXaqAdogGchqpgY3VNKExTjm4UalLHyd6mECM8mFhngWf4+Q6EOOnyMFNkGPTL
OlrO6LeviKUxIgWhRYran4ujt7QoTq0RgCkflT5xm5vVacasH8KAkBaGnqzAkn8YStFC9RV7eGGm
jaaQYJQa2MabJojxX6cfFlVz+1YJzJ5pT8ykaEhvls6JMBSOas90WYxO8zn8DD76ZXyD0L+J/MmF
C7wAFL4Yolq/CrMdhZk+CT92lqp8p7vCJ8obdk0Z5Ys3Z5R9N8REWj0O9KoIoL3dmEKDfhphw1Es
MQnoWQzXXyLyT4fqg/MyqcorTX2M6TMM1F4ECka8wTl+LtKycOFsdSiyjJdoWK5JChzS1Y0wTxDf
qwj6+8lDIYlA9oa4SQpbpc4JTuO+HUl7Yf1w2m+NywHE0Af6YuGHCYB0de1mAMMjq4f9JqZV1+9D
tFjsf/ze1Sjohad+sW5r4f8lddvk85KxyhVOkDPM3HCPG1olWrrsIOvafnMx51i0nZUByo5tkLsF
LdD9btYIm12kcmqnhjCktSryhTD6mPPcN5Ye82LM0qVOgiRu2xLeU4hosDKULOGs/Oj6h2/VtWwJ
07JYSKeA+ywjgpgIO6a8ibzCk+4DYDVd+Jr2T7AciNVPA8f3t/ucceosXAEPTaowwK0FaEFqS19T
5QA81nruOgdVNfi083nd71CO4/KlCRPWePrMjtU9juECfRS9Hm91dFJEJLD0QJVlpektE2eapIjm
lEOnAhuPrfOVrVYh3gYGmNCzqtu5Sg+qIHdzd+u6v66GXu1tckvblYp9VgpvuBp/ZllNX+CG4SGx
VE+fv84VCtZWu84W1rOos/13dJACO7IyTqRZAP3aK9slptxSlN2CJWDziGePkrQXEO883e9pu2kd
ORv3uUSgatkg/D9CnyODwZ+lGAcdi9ZE4sXtLVAojX3MkK7+ERYPupzFB+PMf7m6K+ldMntx9aqD
FC2vYLgXpJvNwQcS2AFaGA44G9irg7Cm5F3ZroJqMoaFo7X+w4R5H6Hem77ihKOstr40BXoyfUxp
YW4/cZw+dK2lvkZ6QYNn3hBP5MoYDadXGSrCvsyvAhuPvPKWHY6dBCSIeyMW0ATP3EPE59uzoaH3
NW0rBfqzJse3zsxQ9Q3t7N2B3XxjpmVQ8jiVOmUg2nRjFp5uCl0/QQ80fuBFWzYLiiNc9zsGyEy6
4JYE0biVLt74/irQqNV7b8gqVsg+XTFX/q5q6pdxW5RrGtUpL5UPx1eNCyecN12Wmuj5WUQDAlYD
6Wc2EvCKR9NPKNy+bKYMb+6PFOOzY26xf6x0WlWOyjJmsfoQvlGso7cubrOlk4tNW6x8dn+o7Xei
UgvdWDkP8dht71zbkFmp3KQXggFKCdVUTWZ2HRZkguMjq9r8yrHcczmra0SoWo9q+rnAbm53QA4e
GmE3lPGRiiv6rRHzMb06eCniF82RJ/oMqsHWY7icA2qpy9o7o2s3cKwHqAo6gR72eJ61xgZ6Q9a5
20oVihGpE5lIlKYtDHsHhzzWiWjHL9hfm5JoR/XzBbjvcpJSZ2ZeF+BizkVtm2DnsJKedJHywkGl
mOu3i+fpPAi5g4HiIqqP/in6pe7h16JQHyCbmuLS4QzwFqUiBLPLvZE+oIIUW30Hklx1Kn8/Wen9
HZZdJhdSbs8YXDwRqRmAhxcGyC+2UmFtuiPs8hTYURfue8aiq8jbir6S9ZRvVQ6NB8Ueh53HYe0u
M/hWvibydUTOoHoSlduEf5dxPVq3MQDlzn46veQmCxg3l7B5XVN22u8VIT/WbY29Jpbm289Zz7nK
aCoxSn+8b+czKkKn0uqp1f+SmbDoHL46zcu7UNExYSm9dAFRGZInOjhADTH9fOBg+9aZWAlX4h1/
7z0+jNWVCAU6iGTIKoBp6DZqBt6tR+S87KSb5VMiBrsMZgZ7Y+iubV+fQP8XNCzrt8ktHeEYh00P
BLWC6L1o9rE2+tUhbdHwRjVAE+ASwqLWwO1kt2x05XY7nfBftErDvHCKnsWLYQ+uRNE7obS8Ct0w
QWryIjNYzAmVcUiLydnmr0KALF1tfzLFpJ4q/LbgJw+DPVz+VLsUUadBo03+J7E6gP9wEexD8BTF
jo8llOQLb5V+dfa+IxHx4hwjKeuTUZRgHaAXkDVeZYi2wOIcT8PtuYR7nE1UICqxKmzyrSUZwTpl
+hRoALlHRMADiYsf0VRwqMx3cuIcXW+52PqxwSb9P7wyubcRIQxps6ypoK0OhQO0W/hZD4cP8N9d
FGXdYoJL9ZlNJB/hvEHW0Lrft6L9NMvgNYKUEepqtX2KrZ28JKNt0wOXHkjmwitSZUG8qowcyBP8
XLfI2j2rzYlgEFuEK9dfFybqbVfOFq6ZiTGFWLvXOoCGBu2l0wqugj12BZXuyEOjAwMJdMUpkEqO
SsUjIPWZMg6eZsAvWVhQ+j64NPn2SjG3nEwuSlXD6cS7+zOQuP5m2XWmz0dpQINLvIlwIRc7RNaI
RxxzwUKiBJu8JT4m7lhmcycJesJATGca/QRFw2SiRpwFEZgkKgzenC5dSSmd+qsFnZ/i6RDztMt3
qnYUoEiHTexiKIxkVuzNvd4pviNFFynPfOBWoWjl8DI0/mEfzfcoCkB9aphaka9nB0p5ZDpLUYs+
CI2wIiJD+WB5zbR9JJvo7Mvf2CisbKJDY2QjUN9DTDl5vFsvejUgir7q8fnQ7B4KYjWqble3iBBw
Z3F2Lvr+V3DGJdNNWWnw76w9xWTNRZmHoVr+LElHzzuD/NdKyoJE4B8Mb/+nYLFAQb3nHqPh5Vkk
uR4MjSU2ohZBhSOLwXzFNH1jESHMcrmGzyPp8nf5tX9L4YAriu3V1iFd5zEK3/TzM98MhzuDSZj9
IeGgL5TefVj5PJR6iInG+no80P6rP4LqowCUTOuc+Gl0pWeqvekXmDsydubN4T4y6aRMx3whnpmn
Tt8jCvIJrFySREINWbGkKm+0Rj+6O44vChXcW61P1aovLLAxX1dT+82hHZ2efDKF7M2J1nr0ko9U
Z4vtXOD1tOYPlA+tYwAMS5ZAlREq6ljCCBXVylWdxIrtp2Jlb2OCnV4mK3Sr848qAoN0Ejwgvw/F
I/tZElhjupFsJAuq5OvBk5+Bw4wkQ//0VXor9/HGdyQLE0ScvCA5SmWx6L+IlfRXvXsvYh3vBeoT
HHXJdRCezpqQnAbq0T2eiuSKXjfBTaw9gh7hUJqACm6iSKIIAUvg+0CSKt8HPIGUha2vnTREFyVU
gAOsDTmPL8NuIZ/Suw7HRzTQ5XqSYNtivxKqZUlz1ENNXk8b1l0Jg+7kp/9Z96AtjDLVtAt3IKdV
2bvDl1KrtqGm/f+SNvom2YVV+/dYNLicMJhmtURVtuC8pcathSo2py3eo5QINiRUx1mC1C0/Sn1e
2oE6458soQZCcYSOQ2hv3+EI91BwmrZa+dbpA5Hvv72iWUug9JGxzlSm5ErhRDsjSxj90xY/7wEl
EaHApcu1SUTUAaACB1/xiab9arpbpWTejcZWH0VG3LRJBws+iy9atXTl0AP+w6l6AoBrV9wDVbWU
Nlp5Kx5LO/2E7FgT00n/p/QwRLkfl982zh6LdzFvbt3hPg+cddpx/dVtsozy84QOe3D4tXSRpSv2
pciCumR8ZxEegC8W1RFR4NjW44aOQJvkUoD/ZeSI18XXH+qM5uo39wUxoIIDMm3m2RIhOAHGTwvm
FRr2xspEzMk/FiIYovrBF8LrCSvZ1jXnKIfwMo0+IzL5mbLdoX4oEVAWH4zpEMKhsEua6rW+RmU2
t9Y67JSdHsazlDxN4f11twyxhA8DfFYQsFhkWiD4T+X9X2cm4SJEQ5RHbr1qt+TCk03upk7eGmIb
7QOWq68Kx0tH9LnzLiByBmqrkj4WI7lh7FU35BRvJJimTnMx/koZRGqbumPWEoSMGxeCxCVOm2Yt
EEpZ13r8vsefIP0MMRpzdTKwJoPORuWRV1jsM595Oz2Q3dHOUZYvYJGwqukv71sXX9EYMOYu9N7E
Aul5qcMIXtXabMTfBSNmdCMp+FlveWUhqz/1E70c3GP8Mx+8jMI2dNZ8XATxuNkPklmBtYuIsjGE
tqxigqMjeTg03vRz80yLO+gUyBPYeUkfgzAEAC1bZn9wbFgmdewHHuWMzXJM+UrWfrbQDwhr4AQQ
PmZlPTzSX2Fc9W+Y2xNNsL4R60nDplKtRUlTtyFPd+B5Fb9bDR4XXr89tiZK7uPztBUmvHwh89Kd
s91Jsa/GkUCurlzZuVc0Ofq8ofIqI+wlxcetuPQtFdqIJ65J4xZzDcl43fJ1thLVK0kys5moM+sf
sBJXN3spBkXox1MRLzheNXoT8wctyN3pIlCkOFY8V4giPBjSaaiOahzTQ3QevFLQZoFtFR0L4GST
DyIjo3yrJ0mND7mSOISk0TLn6kPL2ZXYECce+nFkMaUGmI7c/6Tqh8r17MFHFhgsvyRhB+cvRJVD
ARInWdvP+/41d8kDpOdgfSIM/B87Sx4GiCkoSLCdub8z6uOdWQzHg+xX5yBVTLFU4YIo9My2Hcls
m+3wjnhWy9zcECFL9TyaNcLRobIEx0bUY8ndZg+t8/ER4lWlJCcjfAacNp6HsUTLwLQrEa04cR0W
k/OURTPWqSiTFe6LUjt2EFVuhN0xYNB7phRGP1N8D7IKmD3UGT1nsR8q/EnGy5Da8OsbXv+aCOa3
6pRiRn3bcU6BdcwH5FkSH+ZMDCmcFNWL5SzHOW91AYI7WsVs5a5t3cbnNMthx5MjGiwPb0p6Cpp6
szJmyP7VYABmYiT448UMQpiRtQ1N+6IHkElevomg7SM905RtH/7Wbx5Uq4Hb8mWiYpAq7o1KLcQi
v5c4yr8kANb/nVVBFPLBbAIpvO8F+Tp0TnovpJvfOAZUOHx9oUzxNmEhgFtJT1jEHre0AqqM/I6H
fORnqE/7YmC0pl/ahxVjTlbPeQVjR1ji2XmPXvVFOXPCF8LuT3r7VkNSnzIZLD2m1vmX6Zg1kG6k
1Pvn2BeqUghUDRIkA8Dw7FvcrQqwiSJHal9LIKVeqm3hGygwalqzuTft2Ri5DJnixgqbB65FD28y
4TentgzSC5N0rAJIzgcLEbmmPyolMGRiRKZKuwNsH9PoMGKWPudGTdqxt2/6GBce4XbELggsZXgY
aTh6tZbTybZTU54DAqzhVFmPiCbCFbMZzKq4EWjxN9olZ63l40KUH7HxRjBZKcoi7x5kr5Pjn8nD
9ZYqMpzWOGu5rGRGCRPOMifyO24JfG6gGA/ki4LgmYWwaDWbgx48buDJHcgiaBJ2RbrzPRyx4cAZ
8y84rSSykNOtoOmXQRa2ebSD5CR2NwePF0WNDY8JVGsll2chGmjiAAweJ25JBX2AYbfUdv/g+0yN
/m9CMUFfu+qkIGt3XLdTFiTm48UdDaGb1jNcR9wM5t/dr8t7/4ls6weLV8yOCv8jfcZ3qEhYRJnp
QojqvmZMXYnouaIVahbfUwhiz0Fog06Ro+bZWtMLlCsWhqkOdj2icBA2Hy9NCy4yRNf+2stA411R
OqqongxdhsKAA17dhcK2vxUGMVfsE+rtZuje+FWQobDcPBaVT0howiwe23SRRIeeA15x78baIJl+
S1uQdiEJqWXNefTTUoFkKyrVhk/D1E+v+LcdRRTprjSMlv+C3LlBwZv1lvIMy+4nj3Ol0faT5+w6
B5xvj46i8U95lIhVPg2y35CnvrngW5MG04p35Gn7lGkvfhRnZ+Mouepi285HGJGP0Xn4lziny/bX
MJFW+hU6J9XVxAQJiGV9xZ2frPUhNIHLv4tsXoaBmmYNheyCe+9c4nSifKQJsZwrBlMV2j+P9Cam
TMg0/nvwZGNonckjWbis+74ulcGKrrfLYFQEW/NMobJp8iTvqKpZeOxrtX+DjB9rXLeei758WlwY
N3WoidZJ0N9u/zwHiaEl9MLgF+ds04rPl6QKRSfnsSmwAMQFFUW+rD4EL3J64MmwXewPD/zvIaAN
Yk75JW3wgc2S9/Xr6TWvhYEcEAFgbTMDxLYD0eI3PFY5/V5FVZl7MeeesdSxpQ3H2Ayh/O9XYPb9
Dzh5TBECjUWLT2RjfBT8rkTPB38WfwR3c5qyAtiNo9hp2HWt5LKEGLdG/BfXkJDPsfpTni1GZpRg
I+5NKcShgRoXxBuhTqXYpwPyID/s1Ft8LawV7AvwPX6WVRqdfO09ShEvGG1SEsuLjAIwlfuXXyaq
CGZkydfrJrbjz28WDfjcN8u3ZOuLgxbVaSZ7QjO/Sfe4M+mSkLW0W6rWNGl50nIte5kkWE4/VXcu
G+EpznZc17g4A2MIgWIQilznLrP3On/FzSEG1bxa/jktzx6MXgxccmWbu3kxdfuZRml72NWRH3zk
itcPtLYsoejAa/d/QT2MJUPQBbyWA1s70xGv8YsSAstb7y6JiusYRIdw+o4/+x6dW0UFw2HaKryL
E4l4JWya/C8+kZyFfbTp1LCBrsJBJxRuwqqhVewfNJQDb2D2bmAUZ+J/Tj0WSTADAdHD3bc8998s
WRB8QjQcN4VRfdsWDxhSWyJ2Dzq9OGcIY8LFoGAsAwpk9CObGJDCVfLrV3Oz7US5DDBz8XFl1GHt
Fm8ItQAVtZjIz/Xjb0QzAOQxXN8ooDFqkc8CXvKz4iA+WiEyQ5SIoNKx5QKDEahK6a1mkFjI3B4X
Eyp237/Urym2PjgcKd3m8jyI3tzFqIbnW2Ezc6boPPN0KNUz1TPZIYXaqfUpW9BYsXd2FdSruWCH
kA5N4+1RZSR7KbQ5nkY6lNlT3r8asEHcqLOTd/SxpqRWZHx4pWZ3q9CdwmmX2Q48c9++wCnFP2No
SaDNZyUDCPHwdZowwqsp/rUixNEZew1BGiPDPiV9BtNsO9T7M4Vxv4upe3pHRDy9b5fhWuFcWvVK
Rp7nj1PIy3hMMv6kamzklHOAgTnnmPMvdY7isBAZiDYAWpEzrPhCOyBVop8DtrzXOItnhNBWmGJ/
jnjglzNCmaJMm9lTsAeH2ZN8VuyjW4JhBS9SXJquWktG1npa2NzTOeQdq5QNHE2ryqz4Qs/vxhwI
XZRgDcfhYYZlT4RzBm2ag9hAAKFLPIWfqvtoZ8qK9CetYkREBtqTifcAHoTf8XxrhdjD5Fc4e9ls
D8afdE/GB6VYCDLh1MXZ8vBhImNdJR2LDe+Tj579htcVNjCp/f40hdR03Z+4jS3O4qH8a/PEaIoE
D+5KbLZYHP/BYb5/uYPu7CKVjM5jM3Y3Yt82FMXk7cZUroTE5aBbCS3uTvBhlwA6rJ/+3K2douFM
fhqSZzXRs8zGLrzxgs5eDvWPn7jTwuJVmIW6h07du9PQxdkLNkd4o+K8I7ZmOwGZc+zF4LNjQztr
rwLq79IaBFAs2jUpd6w9Rqc/aNf2B3U6ty7ERy0AxdAjMyn8FUo3Sb/8/JmCaB8Wt43R3gAb+j8H
k6WNc0/f76pbg1d4MSP274TQoSemA7+eTZGEXqh1Zj/PUZZ2hkiXUns6K2MnYS7nC2ax33oH583s
/UJ1FzMtQhYfIxWWrjd0tLwnOigBxINe6HeTFyMfVL/iSXUz5Y7v48JdPf2ut9aGqv6a1JpLBiaH
jtx/MYB409ntfltjoO6WoLfWMTTBDJ0uurANTcYxlN4aFa1TwQwWCrpQWo05CGijzTLvLYS90Odo
HKyeMGC2oJr2RQqC3JOhJMeJ5SR8Vy53Akmylp6lq/eu5u3msFeZZmND5fLcBWnJbM1K/o+Vivxu
UQmQjkk7m5vlxrpqc1RJZyMW45OUpBcSBXJ4FHj1n9JKx2t9JhzrBytfrv+KT8La7lhyELa9pirc
gWj0NVhOdKbSmx49WsHf9VxGV/m2owL/KO1fWei70mOeQe+Go6mrDtfmLNLcbtixhflxP4IjlTFe
Xk5bxV0egfuwruxV+0rFkX0VKX8YW6ZqjoRs2/2O9xPLYQ61zpGZhDLjeTJ/NU7fXDm8qoqxRX9I
z0TgCD0TnVnjpVdASYNSM2cm3MMT/dTSiXDY3WnZT0CHxxZbXogd7lJcqPvM4szkm1zSzehBc659
7KBRjfmUow11/UIHcJqGHw4XNZ2sLY+1ykBhGqg1YYL8G0j43/ZorktSrsNKHoYy3sGRrfonXOcK
IZeA9P1B/TD+REuH4EEAfUB/o2BG7zpqIryU1rzXkwgbOWQ4BTgWGEJPsrfkLsqU2Hks6w43GY1i
29gaSjB32Z2yOBsdEBBwJEhjfuS8DKzCnrYJ07YaKUUQWqsObUMXNVkZ96hWLWWBW4cCpVeLMrd6
0O7eYDwfOPGtU6YcaDVf/d9G4RAgcQE9ngz2GIU4u1CmphYbK5BRfk1MHvh63g2AyccFr9IBd7G/
nNYlDNzcpU8TW42u6pppUBCUh4GIKbshjGRykxIyZpO4b/l5MO3efJfipJ/47Sem5Hlp1sb0An/W
1/KKUvYMu1EwLkJUWjlvKr/FJq+UnyP23/+WHYRoJUu3gTcYtrBPB4nSJP9tiIsjqZFtpo+vXnoW
9/7uke4Llj4JawN1gViFewGpqpb8TyIHMuqjlT4BxgWNvu0DIFgvSMGZafm62XeD/DIhY4gR+jW7
8rby1AGSSSRAcR6BaNzkkBAAOMBKvKgH01EiQ+9dCnipwxUnoHCkeRHsvLq6TyW4aIH8gD/X77fe
DRAeXk141IhACpN0q1veMKr6z1OlLAxYHf9yb6iJe+s5lnQKrF5y6sNEctuBwC+y6eaMEY2S+A49
Zgb5SsDnacRPe9Q6aQE2qsvsElYi6LmmeHRhAjnnevGZ2sA/7t+3kv6WWrlW8XkOdy6kDxqOIa9n
jpTIzNjsPyZKKmU1eaU0emuQLfvZ+sNaTg69tf4LqepB0zTA3WFQ1VXQgPJUa+8CEMKuoi4IJGS8
+CxhtTGeKACP5eeLB93HTCd+akTyZNsaSAaghVmRgy63ck7xAS4sWuc68qoaaJapPgvFyvATgt12
pTn9RfcYzbTNNQBeh+b/BIJ9ZVW5oe5mOQXl1edxnq5cIPVXsphYg6FK9zVK+BxKbNH//J7kbuq7
60nvpJ14JWLNxbTGFe5QrbC8tzvf6YK5qI8OD6quROD8Ezh7mlZAVkKjndRPlsQv8CXGV22IZNK3
phcaB/DfXp5Fq1WOiw90/lTaBxZbd+kvThot2BRSrQToQa99N4stU8n9rAEcvjr2KEq0j5rNk05s
0PUVj1ZCw0Z67f7CDwoKT/PBQJ1tDvjsp2+6dx9lIoDPkwe4WvfuQV+k8ZKpytCe6Qpj9sj9BvNC
spQKi2bCFveILY9g/GhfuWpA7Tl3sVV8NY1flSduoeLRgr8WgXOHYQ7thYlZXDWFpLigk2Boq5fy
QgyJn2M1OyCNEHvHYFQlwst6UnV+lZsJvgvarbbkucAQ/0WP/K9TZafakZa/mgjzsYKzXm8w1NQ3
xh0pDgI9U4tXS7eAbswnjyagrxUjQIzBoJQnM88hBeLsrwpvKm9AnFDNWg8juyhYmGWFBDFj5GE7
yDc65b3lqSagsRcQ71qok0fNEYVQW3ucDqI8EmTtdQLNa2p/zWxb/7lzNWe3KQQmWGzmZDS84dm0
x1RvH9AY5bFR/V5bK8UPp/yG5rGfHqv+r7FcOy3U8bo1FgM4kZXrleWKgZUCCpOpTsL5WTrGqjKG
MXUGHfGD1wvOTMY2YYHqwMCUL8syah8cjH8N1BL0BFnWOtEimdQqjc5jWD45THGLbdLQM01uyAvo
j+x+ShmfAbGCs/uM/pXGpqnrfCfNUU79iOtmU+F3P1QGD0cn0paYPOysIm8kQuGk9UVypR5QyXub
73GnQUIQb4GgXSdgnuyXfW9qlZj5g0AO7aRpb5WkMwDYsepPMjtz2es93mw4C9r5tRZcouzRtlQt
y3Fn9FCD/UdRPeTagGEJmnGGMn7mH7xZvlAG8HbZ4SiWj/BDx3ocuDg9gBvU8huvsEWVaAcOPCDt
L/+Dg7jIcIcKndWNijmlDkuHKizpeJVEA/msomjeRHwwUMgzm++eHcqGRuzqIPAnk3prY79THP/r
NQlTNR3LBJ/ZhFz6UfsuW9ojDUBEQ5DwCwH1+rual34WhqMdBUU66AXAGuHY7HSjVHCzmedpZF8J
VJ4AQpPzkeqyELKihvwDWS6gfCF1eXOIRutbZ72qM6FCD+YYf0tj1Tb44m+N4Aer3q1wdwA+PHKV
KNnn/b+CGQvkpogGvGNq9AVRCihx1lXv91j9l5C61fA54dOh68O7h7JKl1MqCFQljGVz6VHiI+YY
S7JopW1IUSVD/5E0YxWFJDEg2o/NefFrooZ/T+hzqf5QruKDb73MjBxJab4aSpg9osS6vK/UjJfl
gLzmySulep5bkjtlAcJGrnmAiQuTmwnxBK/FZeTBZagEE0FvzAizsSyRt1KpgwXYnPek3mYbotH+
mUe6UjZQgZ4xH/fT5rVfFrAXh/oHFXdBYczAufZyiwUzgEEb5bkXjgm5gr6Wdj7ymTXWA9BeneJU
KcskLXRAmQunMhyYkYyH3EIBU5RHQkx+yrCzvP0kgb97YIu5K5r5MnBwB3Iex+0p+I0kDZ2BVbjC
3Dzh9CC6BvekXN/Ur57hIu2F7xIlI+jvtOmGjZ77BfSV9GRoNP4BODHq8qZm49I9KaDFF5WCR1Qc
gG9guHQE2ziq08IMLZlXslVCYn6/kh5gzWDHH6UsJMjKdtjZpA6mY0f55hVUFUPvamv14IxGx5m3
KmWnAuhRTxLrssGksAndBAaet8zJ9WHJd1Cfv3TEAW7p+mCgEGCgahrQK1Dumt+2yQG99lYGk/JJ
xHzBO03ElN2zNhH1fRsClMAPwcxtm6rrqv5VOkDWST8iyh1ZcAaAQdhnL3dNkjnNsvjL/XCLOpkx
LIRurjhgJBQ15dLdTVqIee3CZgaT7Q3CJPDx5P/7eslPY1y4+mVKKk4KRX75mJ7Nq8sVGp1YAWR1
2U5Y4g3tFsiJox8iqtu4llB8itM4cBjuQDmap5OK+FXjWgUNJMfpphA1msb8cGqELiT7oorNdd3d
dIL2PUZI+z8Z1zMPANHnPEkAVOYSDdS6KIMy9FzRKGV8EqNKJ68O87gL49jfsxDWyxWO3+zmYLe2
mr8oYRlIE4oVclhusCY3qKp4Rjd3+dD6yuM71tBwIqpJ8MqVZvGjyJj7g/CcIJ64FyiAKy2lAPA0
cilJJ+GinlcJMVL9MqlkcieT8zS/KU7qiKnIQ0Q8bDcO/JLbhMTFzo4NaF12vjkroqqwRScbCwI8
MOeHNiz6v1FoG1y34sH6BeUxW007xsI0JPVq4R9DLTXlgK/DpKcNQJ1g5pxMEHpf17zLFzR0kGpk
73qHZ8sJL2GzJATExLSlGD+g4l+/BHGgLgpiYwRai/35y6TukqydkC/Lsu5JVN7VcIDHU9KG5rtX
vm/brmePNIvKvnV5nMKs9Gm/65JM2fk2nVz+8gDcrqpD3IfptSmYvBklohyJ1POe5CMUafylkyQb
btO7pGM06DU+SfBDXqS6SCAXpPQf9Ku1xQWQXU+RIrDXk5dbTaZ8kQbL8PYRn4ZVi1izNI3UadXS
I9qHNqeeHGXbygAXJmKrjnReitxwOZWv7/7LBOeAgdsMQqY2hUVcmt1QcdqEYARu4Z9AICv6AUTM
orUJOE5Khuv4oh0mSNNIlnIiIVMZd9tS73dSpzXMiTstgn6mmJP7nVf+qltkszf3t9eb6mVSusn8
HEvaJf57lzgk6YgMaYBzydUoKVEly+qVR6S/MN31Gtg+4bE2oaDWAbZuYbFu0Y1M1xJK0t1yTo3V
t6r4ga70bYT4zrGmGlcN7Rwx55vdvnP4c5N3zJvJKD7SPfEPTI1wx9EB1cBcuWkjzUhu8MopsHuH
KmUClCogsiG9AH8BAQ8gic4MyGbjKPfaGZBES/AodcRHuZZWoEJXjfJZhI3+sryPv+2bZ8MBo4Nh
YlQZo3SrwGFNHcbuS6OmvouJDpWAKeZW2vohaaTRT74XcB8wdhLc5LxRJKLkkybCGRVCje2TMBaz
2ZfRFF+xPOiAP4/7Kdt4mspUevITZNL3kFLKHu2hqj0rWoFIz3jXxWklhVz2ifVG6wkCc+Fqibde
wecAI0Ancwp4pRK95v0nUYrhaTgBGpPGVOYQrulyb3h7PepIKtiGsCYoEXzyjIoq22gcpTlaQaYY
pMUOpyU+wM+Dco/BFxVg6AvlHvPEyTvGCmq6kQwDsZ4bRVoSqGlco+K059ZyxwpWl/Fk/1404TPw
LpFx98WRPNODH4V/H2qY7Qyo8BSV2gQAltGdajs2nX3aQzG6PKQl3HcSto5pcEOmDiSnM46eG5IX
du2fN9lmqcyhkbZgcIo1GGiNIFnXFtkRtmifRNAeNiAPsyu93ac7xvgdGwKsFLye3FZNGZEPOkxh
wduRwDu7BtN8GhWT8G9jbCtjxVapFy/+fVDhY9DsG+7Mhx+MmulKGh0jezOG1dt3NWmg0LqmF3f8
p7qre/bBGVcwCxIerFHycLdIggd31rZAefaFOLhdPQUzIkUkNqZu7m0BaUjV1reTdx8LvnLS/DkJ
SpmB3/btFiav6S9ztbwtvR212XebqXM5XkdHt0jSR6CYcPa9VN9LQTV4NDODg4CxZFZcDWlWiYzI
ZelLTfNUlBiaj4iJTUx3Bp9JTQMvPqwKcUFVDa6c3ZIPZjQnFxXVdrFsbqwpDZ0yLEbutsb+8Odm
ICwiO5xiF+8RVtGNFzny5ZRZFKGl758KLBv3SjZeTszbaakykkQGp9d3hWx1V3MJx7TDoTAwx6TV
ic3EVgkiFsMEztVpqFjl8puljTnwI3Lw/x1i1iTec5slLMdinK4Z+REqVW8jn/Eh3iBxV5YoGmGf
i5slDRNuSVCWJEkTH8j7yAN6zfhhg4Y6FidV9LJnEPbgpSUTc8PsMPTrpz60QH9FnJeetkJC2AqM
ni4Li0C89l6aCazZ2/bSWwhCv6e4mXW0VlkFGnrUnOMvistySWrUR0s8Ia6dkAsIZGSkB6LkLij5
XULGLpJUOFCJA9Fz/t+XBKxRuT9VRp23laU4h73iemSR+YVKw2QfMgu16h64UpNSz82YXYpba1z3
LtgfMY897tLvR0k1UGuOmoeCSFdm3ZD+1idm5mLihtM7fGEK4nuPgO7bvEa9Mo8qkbbONzm5DbcJ
U+/SR/bmO5Jba4jELzdeNmRSjrkJXuAscPgar9h7SsEOIy0nLuxHmXKwC5r4F6n1GZtCI1GLYNQD
cLxYqNaMeaNp9JJzKwxZha/tilksGOaUZDG6p7b+BhUkc1ggKXjPyfdlKXOrCeHF6Ila9ORraeIX
go/ZB5870lM4L/Ps0wSWwhgVI92VU61jtbwysDIGp5mmYp6zPTk1aiWXtxkwiVXqQT0FgrHy2pul
PKhTODledJDei2wYjkOwq/JAW8IUHlpaeFYS46oSVK92LG3/DyD9t7QOg6Lg7Se9tOCDXmfAfPxk
d60HHhs6LH3VzIME+6Qwb/Svwa1h0eLr6QKg/oH7ps5H0CbgtVv9TfvPWJwiPLfyAwRdwM6Ch/r4
ipqAMFPIL8yRVGbSPrCQ54ryG2ieVApb+9dukSS9KsIlemjo4rR/u8R9ZzhF/iG8i/3AHSyxaAlT
ZQULWxPOXnKlqYbj7QQVTQJ4D3MAdzcO88imK/1oXlxHiVp8KtXUQjhlLrH4op2CWl1z/8snD+07
2XJhXg3bSpI9W3SzPbjeM+DpbfgIdUs4P47i4OQ3RqD4wGr0t7s92gsmb0qoVYlmYqvamYo85RFA
afxOk32PKg0Id2wbU4jsg4PPCISw0JWdeGVwEGqAIudeer2cOAy1G+UstmbykKUtgKRmLnCwRXkn
6gZOHFpMr1KFGgRY0CoiaP+mZESUb508lXaotu7+rEJFousCfuISkiIdQDj2BXR/hDUf+sZPIwtK
LyaxqM2oEvqchhR39uJX8i6A8OVdGq/5S3YzAQNBPVBYU2t50Qd4Q6Q4sqyV3hx9ETISU6JtO+xf
CwMC1YQj8i1VFapteyJnAdsaDq3GIhqd/cIBL0SVIu8KUdIvg7PUlCpuPQlcSxhMEPnwnWgAIhwk
U7VM9Xa/SbaesErhZJkh1C6N1LFy6buAjOHDGUh9B6ZOcmH9R8KAIrwdFrrGS8o6LMVENACW7rcs
8hogbZ23piOFJ7lL+2N3dBuwD4aYnbHC7JPKD2jlv+8a9K3bDsoD6bmWCemJylqPgFCpol0lar8a
lJcq+kXYeO0TeEjVbIga8qs5cptsvHO+DX4IOHz1gT92n0y2yMPQgZHsY9elkOP1qantrjpv5xKC
vPCXogF/+S+Exct8OSGKHpIpUgjr9A+LuoNsBgs5TLTfU/xccOwBsHIjd/qQywuRR6VUePf+IBAQ
LKirqonP4PyMt1caDadwxuDD3b7Z7Kt373LOBcFF16GJ+PZG3JNeOWB1Eyr2BfSXgC/3vlpY+jG2
zwiniaXa0K6TXFuFLp9JuckAYmBFy+deeUt8HOt5JyoVbOu3l6nf/suya5QIkbp1Vn3aUk8+sPoW
sQNUU7LmnNS05Ckd3STdGxReLKwIgX+11AnI4rbPj8JTH1E9pOt0EmRL4wffCl7Fs3Bw3EHTBlQD
xmPbIuvOVmH/0CkI9iMuxeumaex5GGZD6xnRB+RzmlIDFVct701B+Nn1Sqk+Dw92byPEgonRBNKJ
k7CsSxttXCSXW65WVLaTnIV8JkZZ+KQIVJbYAc13xfDwdrSFgMNp+LXeflTqO7gwaqA5hN+u7Tr2
6vfOH4+7GcOa071Ij3fRZAVC+psgx0VhEpWhfTIphonzJFZ01gx5Fzc6ipBuPRU8uXPZXdbMg3Ab
RdACBYuCicDip0biB18XBWRALkX/8LYbpiQRwI/Y+CQTaSrF6fZyxxqpYVmqwrVgrP2AETRDonsb
6RCEIPjRkXF64OCDPx5h1HEUA7Q2vhWKLIakTZXJiEU7roOXJqh++HWAv8guSSWLNFih8y+Do2G7
887Aer83M5zHC4m4eV0+yy0cjR0TbiFU/eMMyvm+/WmpzFHqkuB20DSIf4N7wgLC5ge6oGqaZ8VA
wAekEGdfwWw1kpI49UrtXJOpsiin9jjIKbvIpSDjePwfQ5w6aqIDSquWqeNl/R7t6LfXUUxVGK+0
csmxhgk3NWDDbtFIGx+Uvsa+g2WIEJIcEigLDXY71UlnEbp/529u8s+kr/SfNboVG4RygX4SQilw
8nPsgFkaChu6+iBZmDLdTgNIp/EYVv6Eq9LzMucVh2JOoS8743ZjrPLod4iE8cSvL+Hw6qE27woQ
AAHgriv/BvWOaA4trzKV1+CiQZOyIXYhBnYRpFkPGF5kS+bBLhdJwR0y5J/A8lLN593EVpUoRjVj
PNZqdWgFo5Jm8fex/gKWFneqGahb7ApGlvWKygIKep5lTeHy0zQRpJjuYKf0wsZgtkxJeE9QKkeP
dW5vqdPy3RFz8ASONnXTGA8VPVjb4TO5Pf23MdiOVrK0T5jqNHV6yyRpvZnge2i8cpsl3SFJRp+J
LLu6jsV5MhEansVqU+R/BIw3E0VvyotQ7chkJNbRNAv6dQx66W3m8KqnUC7YP1gHMj4zBcj4CqQa
M/ZneV2KdyLis3waBpgiNu9iTbMo1sGfnefOCADWz4U3erpUJrOMgwpp3ah1U5KO2KnzifTcjtPW
0bL09xYaNsUHpjkWWad/ep3+ULEOFfrHpm0kvlk4mRHjhk1pe2jABRLRicoRg3IgPS0WVmbUg+K1
hXocTA8B6vvJpybaUTHzBDrFHGYkIHifdKnfB6/MtHqpXaIC3DT2+nRr0gNLFdRAAIkOGN4mKFL/
umyZJVTWWIQSGVm128CzkCRUTgpJBtwbSAGoWPNfEPVZOAOC3Bh0I1t2P5Q1WDM6iV7bS5c7lvjH
kDb9U/9rUqnMlTZq0ymPbu18tWNIaHcbp0hZCfGug+595Z5fmuBU8ALsggS0Z50nn7iLPGYNoN8h
KupsIyTXs2KBcdSgIoigonBruA47C7BhSFb3dH/RjU3zJNlMYiqD7H3O8Wm82IlD9rxXTbD6aCxa
l25vO3EOdIa9Q3odhfhtQBiSiw4mFL5YuefwMw6SECeOIwdJ5hUrdarkySF4luaO+qecf8ivSn4V
u/BaqUVC0xq5QerGCl1Ulqcw7J5JUzPHlc/U9YQA967FIYrbnxKk0YpYHj2jaJL1Wp446KLttgbZ
Y1J6kA+E9nUZ4xEZ7+ReSV/ci0PbuydmaRsBG+Zzq39VAIl1UkKvFJyaoOUBIc+qO1kJjK/qwRh0
xm/+/V7qdxE1ZOLTqE7YxrIhw5WQmp8gmlpd2MHBEPHLJmkbuTGZl9+WiJLbmeZy6CISoIAyP/Cp
UUZJOTHIl9G/QSF6ADkNkUw7KW45r4765ZXnXpPuca34a5bI2As/cc2X6lKVmVvuauvMXOImxTZ5
OZjfvmKTM7IkQa1zzo/iakjhQxsdGxkh8yXKDeivUpD+f3zXIlGay9E2SH+1yHXB4eInF4HdxHDi
KqpKddnxbQT6x0dtzR/UcMQOELEE4rWoNyfLtau4I7AVUPaH2Ie/uQFCdf2zQXoscNxenTvhVNgw
2072hUb4z1Qci2gFah8hfhMvwZkWOQcZelSK3tUi+hE9yi5weelPZ59rpFaX/E+REf9OJ/YWMIWZ
Fjjd6hKtvEaTkeueD8tbkmAwDCXVG/53OYhtjnBI6A3lvqmAz1UH452X+nNENHkTaD0W25d61gHA
9A4RNYrqLwQmJ4zWBfDTbtvVjcPe7loJl7jI8URTDTsghEnlhNHj3y+QFUZkMZXf25Ucd9OqDqsH
jLcTvnGtSEfbNRzhhoWXDINUa23odujP/ldlD5IdrikHA3+WBvt5bH7oxkOGBqR7hFlG3Q9pbtD8
DPZbKfoRXR05qhVoNIYTpP7P/J+/V3ALkRZD89xi7darb1PPh3lpS4nuSiiiRiXsb72NFcvyFfCf
r3K8C3m8Od3Uind9jA5RFuG00GaZD9q7tZri3F23YmabQVBUc0Nx8KzjZ1X3EUPkGrDcCwfs2myq
Ql50cPCzruAiH07fTkPZzvUkqCfXkyfPMx87geWvNVpGGw7YCnLv9jJ1NqLBg39w5ewCmlSpJnXE
P3nyiTs8SZOo42ya6WjNPrOTcpFFG5C47qtHn2Uc2U2cdLgWXCrsr6U7Bge2BN/9PqxUd89aAwa6
m3bAOLdbLtwi78S04nC+mn98SFgcmGPKcwvs2i6zFES+heFKATKaTWTcZxTqV/wTpc+0YokI5jLx
Y60fXV7rx4kOvSAZiZLJa665FeLMaJ+Ub7ojdMzurr3QnPZJI1ibn8rFNxfL6KyK/+fNP5mcEw/S
N81UR+zKynbs55YMZ38jre+Y0nGJTlsh2SD8/QnU9UV4oiq4ii4kNXS7UO173eNn5fFGxHSjWSzz
5V9JMcTXVtp+J6urZlaZLq8oYaXzY0EusFaOS/QVvYOJPusjoeE3TChP5IK72bhRcch8wG3QWtJ+
lOQ6e33I3SqTASmaWlZXcYrlZhCbUVqV70WQKZ+VTAc2javfBuQd2W5U/bpQv5Q8ORRi9jufyUwY
s17ZqzOy1S5UWvUHiI2BXHGZsneq3xsmy+WhGfPnMfGYkC1D7yIosoktcqms8DKUvCj0VSG+ofwT
W8Ya1MZ2myBVw+YKhpeAdavUmN/YY3y4h32lwYxqnXXoK+ozCGv2irEJqkODHcx/RXbjpbFh+0SS
xTWf/yosbHltYzy808UdtSxYzIHiyTrZzrCv980lPxKgCfxcUtDRp+7Y9wHb1em7OTFCuBX9cRNd
S5P0ESrCrslk9CV56V/JS98U47rsyOd2uAWRqRqeRy2H6iFkDzn6/HFuBc+xS1JGZ7VgOLaZqVxV
hkFWoeoPrVmZMpvjDzYVn4PDwJ4fJ4Fc8MaTsx+nY3yW7blysE2a7yFk/vogJWtrAtU5920O+chk
6rdt8emNDSZG7vqoYk3kZRE3ZQ6TKhwdCNa9xeCEyUYAafFwIk422xgqoc5PwgDD7DQOjGTVR2wK
iYINFdhMc4wUmRDCLASZOeIl1ISdLEaJD1o91m5iS1q5cI7NxY/Q859D4Kke4wkSbYo69PDcI7bU
D5J/1jJBzgPt2IZkufVXqoLQth0LipDl/rSwAvVemR124YLy31Tb3JoTDupcz+8ZhsO1bzGXLPfL
rfbjGA77CRHxWXn3kHYZmJl4Ui6tyxWn+y46rUyNABrKLgvpgfFFTph1TCZJWJh58O1FL2FaOP0z
6iCf/BLqAABgRjvdoWjtVa6dCPsPcFTlLFQ1tVcoPWFKZNWW2v5uvySf3tIhdg37MlhD6mGtB6QY
KN6pqtdOe+6qGoPYOMmpriD7XRk+XEd/cj5I0kwCICckM2hH38K3HKgV2EAIIlPEPtVE4xXkes0I
ia95wMdsHprFPEiojiB/+I1zaO6d7WI45bKmrlYFb/Ut+F6hw6kNxdu+ktjLb/Lc2qM0lfOXJxRt
yC23YqCy/CLwNYdep1kXEyvvvB+v0sotGaFjGNjBdq3ebph+mcnaxKM10VhSgCWwto8V/Cmt7fWK
Mqqdlz7p9fvMJXX++p6J91Hnord+rXVyx+Dz8Qly+1CvRbKyK4KUhZ0hx+A38aInwmIvIi8b3wto
+rhRVCWERsBIW5a0YbUDLDamqRg7gb3lAs6ae1pY3eUO2UBfo47TD6eJe7QZc4rWNZUW+lwbECeq
DEiDffsxU20uyhpZF9e9V7EstuQPZ+4DAa+aKqD+fvNay1lOjVgxxrM/uP01o1u+4yINq2eA5oCC
j1PL+Eouru7zfHpSOe/ZWYKCx0Lctq689GffLG5gwHjQ7qNF27w1QAgAtTdzu+9nT5kcRHoKtfTR
tH2bT/I+NEJGvTB+5EB5lAn2njWl9UIcQnVxHx5pLj5Ce+hgngXS1Z1UR7B7zY8uDwEHVfGJ4qcH
Iula64mz/7qIVE7st5jqYGr3xrzhMU9acGPrh8PZoVC5bfaoeQHMX48jfVM5t66p0ZbzkUSSytkC
FlWhe9Kg3K3j8oBHufhrXLY2LJRBfyHpDmbLrW7FEQNJ886ZsIhd+nF9+PWxRdGRP9QOzgBMzobh
8FzbUdosGP6CidEC3Xiz+BM/rebhJKJyMI/5cBrdUVbTo3F+zkYDo9NLT7+CbtmSehoaadErawDB
q44DaUrlTCWJWCs0DEixJNg6vcxuwQYnWBdDM2+r9KDtVnVg92cGFFo/CjRSnjxavjRgCEzeHW4R
5valSzS1y3mT+DKQCDE8wWvLWge/yEk9UU121ap2Fh7bm19Wa7gBxE8yy28wCZCQKFcqZ+gq+RSd
ZIjHQ1Hvmismq8y++JUMEaj1nQf0fLs9GjmlAnw3LYczsCKcWrVWoy1SG5WvjPhqvY2r/3tpE1lV
a/l0/geIX3cnBOIuOFZ5TMftQ0DK7Gar/d0yhbjfq0JyFYAg7zPVOo2KsPphCIY2ji1cPguoikbD
AhVLn8jDd/WrGvKdGt+r9wUR5t94IYYuCoLMNs2qLnFyi6y7q40/lLIYZi6ws32iXq2u8ygxE54C
Ie0cBhhHj8S57+hdnuRZZz20WAyGMJo7bG0IkwGKFEBnWt+WaIr4WtkxlJOBuQ/6yAveU98onLQn
MzKaOc7XkkHQNc1FUEnHwbDSj6I0oCFtVV4NBrTtxVkIATiFOYhoLQhPoZQ5GfeopDd2kDhIplmE
dfVTIHcAmS68tMcQJKhUmFkNKbhEBSBAJws3ceidagKRBljXSp/WjZfI9L4reQSUQwJ5XdEnlpfO
62A+cREFBI85lE55ZYU9gsiY/62m6Ofd5iRKMQ1NSv9yAcXq2UIqekSFrM13IYqAjD7xeE0hV+Kv
9TnaT00bf07lCuP6BfeGzqm8P380pzHVaA3g20SW5ypqKPLb0Skt/Q5q/R+cpDpMO14AJH8Ait5v
gHXyWtNHBAMRwkcO4bRQoHUYpMBb0heBqOd2aBkWMeURXSh3fNKr6D0w9g3EGh1BBpVpwc3LCvbP
Hnuv3atU4eMI2Igpo26RdAXGbff6cXK4mzMPJRA9zeH/3OBn174eUPSpJoUO4arPHyIFwzGkazjB
+lD6uq+1W4x0VJWvI/SMNH0SBWbwnTe5Woj4tcSDZjuVu4BoDXYZYpAzxBhBBEfE2U8BQKqS24Hf
8uTU3xQNwhkEH84DR3penAh28OZSiTMy424U6qmnW556xWIU4LXX0Lun1N/3bnWWJ9lRY10zvCFm
fzlaDUOOiCGCHW4vsVX4WGSAqCMEBKfk3rF6Up+YVt6jRr2KRbLr+G3JohIXobMFvPu8uMKFMg5k
jXt5F1a6PnZoc+MCZxGw79DCyScbhMkbE3t+beqQvu5d+QJCUHHj1+JmM30Akg12jA9x69f8NXDy
vZ/s4il510T3PxoFrPUoU9RWmxi2mFRabyTUler0Fib9Oci+YIFXIiZ7XDEbC3MVvyRFvk/H8qcF
Y82gExpeCkJg3fKsT1moQ6sB0uKLXgR8lHWJGT0aG9VeB4Cs/eAf0MKUr7vxgWZyS+dC3bJ5cOzm
1JJX9xINhzxNeedBqkH7b0u0c4iwI/6l4m5pcei7ZmeSLVXQqJFAAIgeqI8d8pVZgPVC0Mjvhr3n
MnLgQOw0k8pvdITzRCubZyOuD3jq2qZlmgCspIH3+IO+i71U38jGb3I9ziS+YOHuvSUCVJzr1Ewa
JveI5/e/+xfZmHG6QEY8LjLzFMUPegiR/t9iCkJDbbweJHZJZl9O8W6fsVJgK5h8SIRAiu9+8iYz
Ps/VpaJYc6+MnO4ttXKEGHDukhtxIauZqua139AkE8y/Vjim/1txzqWQc3OByQUbpoPFi2yUaOWX
3IriBSpdiTxPek6yz8zkERvtR0t4y4LFuCeqdTtU1tz7pGa2oC8+KcJJ07I4ysYhrn/oJPysyTHg
QhLBcCYB12UbINIxPS3BWTjF2mTbqaO9vTRqg4CimGAJ3rrdyen8lBaupc0pIZXqDhrNsT8YFjwh
vakD5P4LZaRfDO+P4Bp2GcAfpYd5opD2rNaT47zJJiXgn7I2ZphWg+ksaf+nsE/YGL6+5MCQrLrI
n8ZvoTYhA+w157Z5VNuwQ81N+45a4nVPrqndrqh2vCyjW75PrYsz8bsBezFTGO41UoOZ2GGXTYG4
+lcXD3Qz2WORyJMklPS8uw05hF2TNIIv+PmVVRWVGOs+S5LeSwUrL/2MDnWl7W4+ovXDRVshFPyl
lWyTVjTYvGeaMxs057VOjWNyONxswK5/wtieJn92sHr7liihg9cJSaoEf9d6FUrSHc28fl5fmME1
XX21cng8fV6xALkfNGAAXc6tccFT150WVBWRZCmh63Szeoqu3+n75/GVkxd8QiT4R8QCwOItI0C9
nhTmc/+j4JfNuWBzn11fOHR2NxpeNHTueBJ62jLxBvZGZwSYCj5NyKHTotkaJeyLg/NJSltlsyNU
UXCC3FvaGPBwGHARcGyhaRaMH8yjpsRx3LATuIflsVCPvJnVPKvPdUEpJbfCuABK4YIoBNsVT0WB
oN/GKk87NRTEt78fmBuZY+uCiUn9WB6SG5m6FdNu7syurlMgR5DI4FC903ze7Va+e4gwwLLVh4/V
JAOvlxREaRx5rVSlH9n/2sR16uh1E8zJ+7zsB5/YWrcUTWUB/kYMVJprLacZSLkoIRvmrC+I1nL3
tUgm7iY1Ehc4UlUBJCLc31VWeqGoEqmzLsxL67tKFkGQ9Zbxwdy7mHz86tPy3m7YOWQ2cVLpCbJ1
L91rTf22cVVTlEtka/XCJb/C0wOgH6BHvt507AiWnDnjfOwdiZtqNjIRT0UIH7mLkBXmrDBafqR4
5e8tt2eaMPABL3P3Lm+u24nKvDobYjHk3U9zbTQn+aC6psC73QjodlmiUFVFZYoa1y8Usll9gogX
IECA2oihtn5ZDV1xQM0fk77b9FEQ4CdgY5qHGA9eCmKDDiAxHnRuKbWoOF6DOwm3552sY0kGIoLp
s17mTfLw50aIB7urnOUU5Vb9lu1PR9Kz18sBtO8XppRXs2cj4i4W1Rp5SYSTsHDhywGI5lBOGU8g
NSAdSMk2GFqk4d4SBV0tZI7gKo+e0Q429re77MObZdwto4rGQlDQg+q/5VkkHnqJnpxaG5dLvFV1
x/PwJbVAUO7hlzfWoN92BXT+W1hPAhCYrlPYFaXVkPYW/ZQXtrvhpvY3DLnsIyeYuauFdps3OvaM
sHoS2rgirJwr9jzSsK62vAKpc080d3KmBen9A2SLnwbikSl9NoVWUr1EuxXLCsMISJnvAZhMi2cx
8NRibiqus9O8LGrkDz7I0bbfPI8EIfQRzbhvCTzPS9GgZnGS0yvadBmZ4LT/Ui/ibCXqhmxuu+lA
k+EW92gfTfgPD6bk2Kj5Zkol0FYPsOGRPzOEoaR3d7Rs65oLR5Pq/6HoouMJILczFbHU9rid0kUR
eu+skoI8voX1tzv3xBqbanEzxXM1xV24ja94XM9tJtBNcJPiWxWDUwvCj8VhDJvpaVIGkDJZWVIQ
ir5/XqqedMadmUJUHuRPX1g2wVFJOhjAfqHzENWdjMaEdGUSWZPSSiOWMo8G2Qb3J4RdqsWikq9f
bkclPlQc+yweT5ANRfyBsCKNm0UvgHs6go3GhXO154I95bVGIX2oweEZRRGBKTJcftTrv4n8U99s
gwaCeDsqyAryX8muZvClsQF4XO+zDaEckRrwmaAUM+h/+YEIUQAYvDabtquGwDe6yH8DFNKpyw5J
hYyGdSU/fkkBsDowhQio8Amy6NSxpc3Aea9Jfg8vMPpCZNxNlDwOJ6vUZprpPqCV1E1iKlTh5knJ
YLRRy/j4kk+usrwSMvuVNvy3Zyd5PsijY09oxzUMoHQJrMkCfK4BfUYF6R40axCXAPZ3cFTMdjIr
cdi76AGy3sbfcoe0v64gqZ71uLLrs2/FVPVC2QKFEXBxKjAndzIvKfx5IVjDBxIZPXmbLqRaTe9D
Ruvw/PxnhuaXnC40I84hHnYmvH6bXeNiJJt/p1hQRNdy9BiPj9u4YFbNXLeBeuXW8EwY2b1H08Sx
x5QhpCjgLAN52VrWAWGIxFonRm0sMuUzoF6kQXlgQYZgPbZJIFUDwr4d1tbbeVnmYPZL26Sxlplb
sHRxRRmjQluIzU+yoQa9IJzGvyU6R5EggZgOr04NYUkFdripWrEeePHBjzzW/2XykPA9/6TsulOg
xpk6EEAjrnMmORjhCn82UILFwMexmGQN1d191VVFtAtogiYvOI+SHwc4aluihWMws1FqzVv/muiM
cPbNkn13N1HLsYBrEpbnUnEC8DYtGLeLRQQOBJK/3nTk0H99sdgSNCAc/WOh8qe7LS7p6MojaA3l
oNy99ZDcO6lGvGHQd8K9oSbOOkhWDomT8BprqkkszmiLoqh3nKlyslUsibZGNQ8jyWzbLHvRzECO
pJMR57vLmz46lqfsJYSGI/LizTjL84De1Qd1ruhzO0/nMKi7SMSfNPwXHYBYYN3hb3ow5djR1+yp
jUVpcX9YKyX+B14KooiiJioJkDsa27bcuFsGeC8HsCicQl3+NTMh7F2zz/59lIoNGLf7ZueuEQui
rbtD9DZEcc3zbhICy3CaOgxJeBLBaDWHXktdH9N6t21SfYpoz/d/OjQiuEqxsk/6ES7ycTgWxJXE
ezz2Ur/bcgAXecUa6uCQ0ELleIOfJSVKTCUwg4bJ+KRMLRz/+d/H41ZVl+/2Az1CbxN9YKUfRpiY
e0t6IhsOVIwArNFvZhLaedKIwZUwc6zTVO4XnuvANTLD2dIPBrvOW4ntxerzMAPFq0grPud1wyN7
8/pzndUcSy/hsUQ5oEwkS+Ww0Enlv5Y55b0/kdeLr1yaslrDoL/7N8aXQc+WnX9J8cZmtCEH7dPJ
HWPAov4nnpJvYHZQXtVURCWNw/menTH+mqAFUGFlNPrzPLOfFMs3XrIXAblO5HscHGO4WttQ8Tgw
m7RDqZtgoJjCWIC+vL5wfe8fFr2co17doeNWFevRKh/WLqmkiZ0gpDoHFY/5/KscObMJDmGAZvzh
PjY46EBPULfNtMBlv6HUUdo4AgrJyAnUtLV1sJPZd2ar0gJ9q9oUHtA1Le98ILMqAJ7pnWIBZUcp
upby3bqNQhBO6yEXC8cyf6cUL2oGMbGLIQ++3N+qfWf+RTVuqW2dxdikLb0rOmnooMBq7eF5qVkI
7I10ZSFTU6EjQXwv1WlVszUbt9OsFOnlfQPK6XAAAKkaf5s4puwqdzwqMr3k3+VCQ4cvoJQkCiJl
Iqr74sac7OZAt++zS5eSYmDJ78iDP1IeA/NnzhFkZLUqLtTLmY87u2FYU+GxzqZBRctBiVvppb1B
ZzWUH8pts3oSAlEhsuwKGZHAh0xTWMX8ir2YeX3r2N4CcfOceLfUbF89n6jVmfXBVYj4VBo37W0O
oyU+7tuIuVcWMFuJTjsfdTWHFmLmTePyzwF+EkAKpaHEofE5m6SK+OtbU5dN/rKEqyxDqmf8GXKm
hZbSFccP40YIVtCACpC2Xf1ueTFKWop4U20F4y79Ny1w93zABePhq5d2tja/sTyqOONx9gKgQ+AJ
j1kYVbkoKIG/AgHWfnJ5SsiDAEiFB1p7Lmr671j4fzlo8Jnxo77a+tBSnD8W72YC3D3YUQtfyUoh
QKoCxsiWD9Tm5712Qdqb9sSlrNy4a/f1lLMEDL4X1KRvfkLa/O4qoAaIdfOvT5dbfAIPDBJXFOFV
Mh1/dXzbZABXyuhQJ/K9m/FLAa6NwBqbqJjgPEkvydKy3SBiQU/b5aTyY7/PCnb3b2Ss0tJx+FwE
u/G+MEZqJphJZmgZX6WHz2NkLkx3Nc3Bbi1BoPBsyjslo9+rKlOMEnWKt2AqdTZPxkJ0wDBNGLQ5
m5K5JlaG3sxG53lOJyAMencR/c2MNQaZV8BLq8fmsYiOPadOz/vGUKel55uZeRa6BlIUeosjM+a6
GdEi7GKLPnDHyoBBS8pws/8qB5/G38Y+dD3FGWF9mXSgvSVa2/UVpErwDfgprDfJMyIqEvUM2eZT
cOs4zesSpQHxl3VjfZLG93pMahizk16JxrkjrR5aFLyWpMXJ8quo2UIi3Dj5PigXBm/+SL9qQn3a
wrNIvk4vokKx39QbdaKyEO0YTuOh+DB74I8d2aDt+BYjvYmNRg0HmrOKhqg6e3l8bhvKgrppp+wd
xL+8Kmre7phUsfHgGpoGAo0SMO6Hl3Wuk1mwiJgPcmPlHryqn5R3u+Z44X3CGUUa5yce7HR3ot47
s4aVIMmC/1Sg+UgA9wG2HGE21wWx7DnHKOeC9nHQm/EXW75B0Y/qBnZ6GPkxAHk38BytO3h/MEbP
ICMYXkyRFqwe4HkAEiU8jj67tJkEuagSxskHqZEgqIkhRMuGTHB820fcLIRKjPoyRctWmj3FLkMq
P4+q8F3zBfnvvca2/NGNDRzd6UvuAX3qPNSddj+IdJb/2v4q+jZak2ESfIqJ5mJ77vTi7y9GS0kA
sqCFuLvIcSnPgL7TyIW5h2G3RYFwmP4d13Xu5o/dOnQjLUjm+so/AKr3P9YjkAK2rXR+LfPs9i0F
g0mhGHC9OeHbRFZSGdpjgcCUg+ovEQsaUF/qIuM3oZ26xnGsK0Blx/EczlIFEOHWuxwbH3CPvnu9
s2N4xzTGzAHeJaeBeaKDdu7wBke8GNqsxTNS16nW1DUvBLp3hxASWhw5QENgev6Kta41fcFvdAkR
tAc2OG5xTA6lvvkZfXl1nRiDY7xN8ExqdtPaZM9SKrsLrY3hXIHM8zKuBR6M+JNeVA3hKo+fpV2E
h71AvxBeRV+19XlTZbrUY/cBb5PWwlnBIsdgoyO/LPJ7gsbOhluvIs0XgIPZMIURsHIL11VBm/0D
0GbhKSkkwzenIp50VUgqoKKhxZ2AbINiJbB4Iio5/FzW3ys+hRHlg2Gv7hgPB4tcQOt77TYY2JWU
cxA95pGYllEG9pk9qtB3TfGaP4gZzW55VbTAt56Qc4AiR0d5eFPiegUWH7HlnLgGgVxnEX4SuCch
H9CGRKXYzcSs1UTzRqIRLtDuHsCEyjuTJqLp7+kjpBQ97J+1tVIkKM3d8JqzfE/NCl6OYzr88YzU
mkDcVj8DTcQjQCpepBpCbEao1TWH1ngz+lSqwSAbvyMhmcq1oRF/qvtDc4HVASWp8mmaBLk3kVVv
0fGBP/bepnYE8plOGVoCb8YX3ilIzXnlkL5MMBuKM+HYYyGLJX9Nf+rlzT7BPYmYXA8JTy8K49JB
0JlcR0sZbQQ5tuyoQmglDGa5NrrerrNG1AHWAA6wMk/Wbu3ya8lq5y3wvqhUUjzMJMYmM+0rsalm
tZ3drhMU8zfGsFiSliOJwdYwtS3ss+dEu+yfdFYQzcw0S533HCwu9nr1nbgFantCmn0+TXMwbl1u
6rZbKtL4/uxSuRirJlfvKDQdzuBEieW6TwwFR2mLaUJ0jA28lM1ussM90lW0cAS5wwZ6FPeOMabK
HHdKA6efyUSfbyewQeVYhMxJwC+FQ6FzsqRZ+RGM/nQ4HHJzMM6tQJVFWz0ZoqVgo987usGsxHyb
CNHJaT+m9LPMh9SmwF49WJQp6dJG+feTz3/L4EI/eVQIk8P2aKPuSMzCJseC90g1+08TP7qxfW8e
EEaJEh0N078KIMdEI3h4+U51ugtkF3IfWXk4IedEa2fdsDayusapmFPV8sNUqMbfbmVaZL872Otp
s5SGm4UrffNRy3znmJmwHbBgzoYBYx6iz3/irrd9L1iTnN1qCyufBgOCeYCsB/ufohiyNQclFDbt
ISxl5RM+ej64umdHVSe5c3v8PLy52MX4K+v8mCRK50DWdO4l2ZjZyOuif5nYja1aGw58n1Xm6E/9
r+uzLTQaaXjDyEewcjz7+KsOJ6PXuej/Mttmht2d15ftYX0LwFJqB1AL0m3HPPlso68gnNRVHiMD
UtNwr2Q90I8cEAJGtq2JDDQRhxvvi6/lP/m6cosjxprgK2kixLQfjYLGgSnUt5Zs4CaXv/gvK3t7
nn+Atfgs5Vx6G4O8cGl9/ciTYomx6i+fTCsW2ZnAEUHV4IAJgLzlxBiLQj97cFyDIBp0Luzf4Gut
5XkrSUsRo9iAPR40CQlebW2zGx1x08eHk2RtAmZKiXigXa836q206iNTTC+OT7SMvB/A9Xn6isvB
SUWLZKAUUGGoWhh1ArGEYDc9rzlBIcv5i7sdYQjn3v3bZgDW2mddsSFFl6aEhUUm0IKEEaUBAij1
p/DZiRKaErjO/4/b9g62ZIdjTI1/M9k8I7s6stIYI8aCtZC3nhUaBcsFaeWDo7huMdNfDrBGprxW
WJ942W0PiYVb1yT/TJj8L1Nvz79KsZsioFVy7uME3Rqg0BXzk80xdWsV56MmGb5S/P0Cxs/2sN/r
mllLUWb0r1S1gfGn1t7kmTjXlRpMa4qsldozeHNhRp+uCil4BWh+lPQvuSC+3kosDqlxcTd5cLlW
WnaWtvrlBV/V0Oy25Xg4fWQzqEhTDB+3xaP8aO2uupQYFA/6n7kqC1O/iUiT77NSEG3R2+Hc0EGV
h+/Du2xx6Q5F76w2WmmYMwtcIUhw/8HvqozaBlHaO8iVLElbpb0c053tBlVkRD3+M5H8Jt5uc0u2
rdV+ez70ernEmlcOJyXpcNH+CLPp+pIdIsESF9hKJJxm5AbI7759PLit4xiSwuPQ2bfbuxMDyrnh
mgKm6JbfO4/NlFgnfEHkEflH6ozyFVnlu8GnzJhY0eUMfRcBgKu81vDUP3EVB6hlduL5+BdVcY3Y
NGzot8dyYJ5j3kJi1+t7lSrN5vLkhJ4lRYCFEzpMT65kcpIIMFaMWYHHkFof6XrV1mfMaI1afK7H
if/MlGwwp+1wDEQeGcGcvZhSWf9fxG/Bx4Hiig/bsEvm3iKrFB4cvU8C9KrDDvF8G3H5FH30n4Xe
/z6EGVxTkbgmHymCBs7S/AdvsC4hCgbY9naJORBNnRmKyRR0KaagCtgQORNB28WnR2lXUu0cSHPc
AZqcw+L4I0QjPeqrpe5ttXIsI5f56JIUxE4g1vfYeWvLlcZsN8ZnNhLAPpzwXyRLVxYDQbT+Fm/S
Md2U4de1bFvsKCH6feGmF8/44njZ5hbLimkHuEwzzXCyJiK+Xu0KTjuH5va4iheK/DDM2Uawm7u9
RljbtDRq9qIYKIuZZglDTkEBxcGoGZ/amRSSWMHhGSHKg+xjmzqkh2mlE9qXBanLoMePBRnH4IOp
fY0/KQDwj759dujW0in2OmOORlZx1aDsMOYxggP2q6QEUeJ/WxmU3qO5hUhvtdOtuLrDZrpce2KL
0Yd/pEvxdyj0Jxhx4U8QwlDr4+6G3l6Uaxx3VKUBvufDJMwYGKZE/AwDHkjO5qjqoUE3JWPZMcnK
erPHCEZviifflxNNlGmo97SMnKvyEZJ3pVktIrtZK5gTEHChPEON0k+BynJZt9GePnborRmfvfbF
J9/gp+cuHu7hPjHDPiuDn0ZQiGk1YgObo1FCy2U+N6NCJiQ3YlMkh6/G05jaSnK08f9TOrrvMaG0
4zZ2EcOZ1wWRgwYn5I2wmNrHDvYM2qyn8f2Edl/2fPtx6w1jGqomVQlMj0gYQfNsRL+FVVfOTLnU
sSnkj/hz/dcDmslwLYb0ZMGAmM/ZikASd2mBN9TkTe+o2Az2DOGL3z0pMT8qrx+KmjzH3/DuPcw6
l8v7akN1TDsk0MARcxm0Xf5dz1E6wlE6OjZDTzD5GkGMPb/qFNkUo3wkxOhuYbpS3ybHSpfPVSo+
EubQhGLe55BJV5DociDuTt+yk2700P/3EQGuCCwKgeFR6lMSvKT0iMMn5babJcLetFXiCAlKTDfw
A82VFTYA+6eG8vPvpG/351q79fU6+mXufzk3wjVNC/XMegWN/bZCwMIFLwYlxUEnESRv/MYZ1P6x
XW0+Ig8rj5Mux/KuLNm8ILEY4s87oJejpfUXVwRmQzLfIOvOTineVNg/36oSBobp8Zgcz8cquGKi
ZPu7pWXmlXOgrCMPZYpuzfOOrszpHsBjTt9mzoAHvXp9D6KyZJSmRe0kHuL/dQQv5Xdd652b31Wl
p9/WlVqswapLaGcychX01EmQ6fJ3RdU5+hZajcF1Cr0CvFr6YSdStEIF9SBYuIJK5Nuir8rk0PAl
la0c/4rz5MfbFLSwtwh4L4reA5qOWwPBkHPdxoJZrubI3KNq4tQ6ofENOFdaG78RLK273h+xlMz4
Ieiw6Vyrn2XM5e9ZaPL2v7pJ2NqUbHv6K6jY9O5RXJHVz9siaUIeL1Heh2Dwrye9dg0n1+d0z8n/
QSyLbQrj0lPkBbu9fUOYkeejxxJ3aV4RQJH+baHKQxprny68Y1GVS5a8g0ZdaPENGRjCoxzYgUsl
4no0RvWo0DxQxlRKPNx+RB8yYhwLPWyIvXYHgOtX2N3t0R2pItNqAlRL+UeOQqU/62QjprZAlGE8
aiLTDZuqkkDctLWaEW9dHqV5KMCchQlp9tuqGaNLG5RrkQkP6sAS13i4Hi4vTyjLqbXt1relsK5t
rJsdKvYpYRaWmuhAPs0Za9aacPaKMhJkmgMpizZWx9RpXupEIcYlATuo7X7QM6eAvZbNmlgFzuxc
FQyxV/HSZwVy+AXkKDA7JHMBAaWGN1uxRDLsZUBAwPET29npJXtVmsVQ8tCpoYlvlxmiws2tfjfu
3PAcOOIEFtaPXXtT5Ay8ktPzdzK6y7UtSn4E+0KorETGnpaDRmaAtssKwYnhtlhVECo2/QGyQBqa
4bh3geNjWeEDNGvnalqfFzQUM2XF31bPNPyzqD4tpPrZqG37EDNgyK5zXy07Zcq9vDpIqQwUZ3NH
fKvD//BlOEFU36BKvDu4ITDCLJzR+Z04pmcW6jw0+eiHCShyWGxIdMkjkQ+KbUX0WT6j00R8BsBh
JRYHshFpvzEbUcMsTJiGRJREosD7vtlV2mcCDwvCfEAmm9FlNWZ1RMYaBBgB3V9+zS9+9Tm1PKRv
Z8S3jxwdxeCqGCW4+0KZ766Ys0Rg/gxP1nS+drYOKaeEmChJZpFkFXN/1Pa4OgcD3N+K5S08O65X
m+Eaa7PchdzinspWkdfV5uZ0MWOoanxCESEYBNEmxTKcNzi0jz0EinGkKWgKOhgVWxmx7HPtvT/7
xFTteqdQuzZgVU6yLG4Md6uiF4iumk3tn+39DEVojWNOot9e7sP4WNks2IPGYcGGQj2eqDfalrJ+
bPF+fHSPLcdT/2mmCdonYDfZLOh5a665XhBujG4+hKgtIwFO/Sx8lb+KAxb1KSTv4xx7kggSaPml
GU3cisiyL1AdXKshji6w4vpImbQm45T/F3YGpmR8M8uSj8/Kt7H0mIKqAXrxtNLiMFhjTSc3Wpde
slRJKFA0pgl2FcMOMwiXmzinL95s/ZVVfyLy201V9ZmaaTsKV3DYdkJ1FvhhoaL1FSKIu7+VYAja
lIrYqmI0KL4SE8hzDPhNbOtwNUojL5iIH3GrPxlK5PaMSbP7w8iyyZgY8fIorWc1A1M6FB5aH8Y/
GiMQp/nvcJZGE04OKbF48cX6YY7fFVmwgzs52mR9+G7LyCcb7i6A5vJXrardqiGd7wwUNRAEoH2Y
x+1ARBN97PL6IJLPdlZKZXvte5WLZfAfDYjMrbfM2e850wSzobHjBVwcH09L87nkowssXYr8NOD2
Utt1PDxfNcRol+46I8WsKP+JXk2MWjV8pJCiIBJARTgmnsnlKOPKnwrXKApYLmVFj67DgZZPL6aQ
jDiJfVtvvZwEg4FXR1c5HPMKb7k0OsqlaMdq+6LII3x5nTGjEC3PhqUHykCT8N2XIl9fU8fccPuN
D+qNAkA5oAfAfTnjZRMYg5yQnCrRK9b8X2kaO5l2RQbZCUlTncn8a3KVQT65AP8Wrkhcur0x0o1H
8Gs55WyNH5AM54WxES8MqhdKtm9hXX7BDeRA6fRWbf5hx6HZt6onkFi19MpqKcsNkMOnlNyzLpOz
p/fOFUeLcGCV65trwyaaIiUbOCmYG/a3Snuc6Qjic2vmiGmxqZKL2sWBrioX4QtOEtVs+bh6SrSq
U3PEI/lr/y4E9dsRuNTtglBXAHa5u0QKngmY2qQPI6uNqPlOwJhPHFcfPmT+BBhfIVeC3/2Cznd5
Mmmnr52aQRAdVZ5VjdY6mx9sa6ukY0zNqfSHW02K+kXR3qzKGdjiKG8aKCv8VSc+QDH+x8017zVu
+x5AHDuoWT67so79pwHAqfF7resReNpZyrpvtX4nq15KaEY/QyCd+aTiFiQZFnh/nYoDLmCcD36/
qNTBdpX9ZBW2IY/hx7/QUVaiGJ+EX9Qw61VfiVKNcOZ9HykLdVU3/982pF2EQD/QMI309qKWBI9R
RNeY3lzWzTmPdUDCB7yc6rUVB1c/A3zSJK3/gRUCL0spFSErgzEATbx9tnssGTkNcSfq82csDJYc
EKBnK9sltCfiNFVtoYUDnoXQfuakXmUjzA22UhPP1mbTY/Uao+Q1C6gKCLSJ55OK+metWC5jeMCY
4yvYtHk7Ztv5dm8zxQCgYcvYZIb92nUVD2Ut8PrDMhL2h8inz70i6XCAChucIW19m6qigMwkUC8a
QaD81eUvQvSX8zd6sOLTKMpLAf8zlb4Ggt+QmsZQb0WIlsTK2uJtAnbKal8wDv0rdqvK7BwRFzc2
3AEPXx8CuzxHFuPBmoR8mPG+cH3UvqdjYfaWnWEB27fHqt2WzNngpM0cf7q72f/3CiT0GocstimV
TeH8liE/eYn58moyf3tEsiVvxTDS/nxPyk4DC3T1cRWhXAp8uZGXUp6CCM2WrXcEyuRLKNW6egcf
Hy0IcGqiNDpkuwkFTA1OHO4Vbs9g4WoP4Fh1tbiW5jICw8YMi9M0IX6jWHBkUOCY+Vuydc14PkYY
PzWkV+XRHaCU64lPnt0m0ic76w1Xb2BErco1BBV0Q5IklbNr2inJuYNqu1/MtWd+iBzyhon29w6Y
atFAmUA/kOPQpjiVF64SJPGUsq/sCPXmw0XZhOE6QTyu9eMwCacRBZZuPbeEZ5/rzAszvEXSB7Go
beJJWL+i2FCjcrgL00HeelViIydbnB14mOW56LrCBhP9nO1lD1tmEBT2Tc1tHs762w6Vr3hmvgqT
BCfoegMN2y7oVnjb+95/NWhMtIzd2Ef7g6fg08UHQp1bSMO+U2mzB4n6XeU3LrejXYnwFxVR77dH
veJJmDME5boCeIffGjvThk208SVs0GLqOK6Wtip52EhcSEqAIvl5UKYacl7V5cEjoPQb9RXC6Z0P
O7m/G/NEzWm2dQc0u3pRTcjySYZacedrhCOKZOWZ73L9yXSS6UXfKnbJdPGvsVVtVNjNhhobqhym
vOs6wh4FvC1WhU/ux6KqavVUCabLZ0iONaemwLNoMvorHkqA8kZtdK8UMypPa9taT8uqMsnWbtxJ
UU17+REJEo8g0hQSyc9hKs+7VFLHEgYHTjSlYAJEC6jXkFlHoneDhD4xyTfS+JzXCgxl/+wHkujj
6B0HOwv06CORID985shkfxx0xKubBZfH7lu3w/xShhYOprhiV9C8XDdAC7gbdE2eHc1Kmi/sP2gG
NTMMbAtbW6riDBSSZrJyoXaueFzE8aqUEMzWgOgPSenhnsLeCMor+Of95XkDfaTBA05+UwzTo27l
LsN5xBG/ijAdDFwLNt3acO3jXZD45+mcurafwzdGc+1N/u34ghWqGw/EKwdL6wyNscalMgsZro5F
7gVG9CzDJPHLwSJ+FPnfY5UkqyuJ3L6LHYzOJbKnkyFFMQiNzKSn1tzTYJ/i+aT1j6RdtGiuSW3C
E5YiijPPDgFN93MICZkrtNCsR/LJGHQnXCrJTb/qJ+05ri0KL5CAEPE/ZCamLROljF5nANRL4KpS
9P3NV9kUg1neE0L0JVrIN8daMF4lanMLRgO3wbMpYv76nWsXRbJNrMFKRgpUDF8k+/fGVERkxr+P
nSKq66eoIjFJAR8nozTJ+27MvZmjtIRpX9UMXQM+Bbu7lsU/kGacZ7j05fEXtGehEvQs8pEetqfD
j8qJW9i9e/acrE0DD8tQqcN5lGDPbWvEEKR8tecqfHDYiuSpOcc2IavEcH8Fqtm7KjKF69Fov0dK
YAiUaBJxF4yPt/v2rJKfBNNofBgNMlMzh4sCV3eqdKQQpVK8AXwe3i6gC8Uf7siyU3cbTXz62l0Y
uA7ROWBHnXTw41Ha40dxkv6TQ0cOPxmaOpuHg67OerUnJUNvHylx0EdC/cmhXlDjdYPBF0b5WZTM
LASy07d58xKa2OveGUHGh50ua9lCbsx63u0fCSDuxKkDHbcV9oziGCZnc89sXwKnxucrrJiPorO/
ZVz+5rsId2QtLpLiUcc8P4BlFIV4wom9sqCbhnSz92nwYxtPwPMXy4RxRkI0G3XWmvv0b4iaq2Cp
kUUJpjCIAD6PsnOiC5iIX666QFKQiY5baHUxt1couJx2gODzVbP/lEm9jNwgFmky1h0FQD3VKimy
yRRHhm3FwfBPxoIssIrRsA+5cF3CXXDuOieRfpAg00P+13XCFm9SzeYbqWaEz6yhqEGVRPUiYodR
LQ3pwYc3vwfyCtmQrgZS3rgVOYxsCYOo7jAvRHZYi621mmfXl/ddxs3cBij5uMDUmWRNCweYPjV2
QqPuShuyu8q1JhU/fWEcES4lC4oCq+2IOUGgX/tuqYuMA3CWXGq50qQJaJIFM5fyfZlDsF4jP6e4
Al7RMgFVhZ0hxjBKdEqp8SlsGHiwSYx2A9zIqVnK4N919aw4ehlU8mW1NKr19EB2gv/Sx+M/enal
kLu9I7hqIwyg6m3GPSw0FKkd85kj8tUprAFaBcjK6GtyTHTgpfXANM3xga6VIq7AfCzzOusUoyWi
qgzia/StIMTxkP3cMFbrCG3DHaDyAxnyvQjxFTjyO8EUMcRfT1/4YvLo32VTVIXilkOHog0sAY34
qe9s/F2dO94BJ9zYUYGJsDI10e63tYNPnUUhZ5ZHQ//CrOa2YitUpv3si9yCesCSk+lreN4nj1y3
tj8oDvJcaQwL7968igOJF7f5aFZYk+MlctLRoLqJlVvqa2Nth48Ea9mzgexUoEhoQDXA1e24wz3g
8817s/PSSrssyxh3n1XtmGoRW2OtagYzpIyak5W19LmoLm/dHetp0rGu1WKA/C7BYfvaX4GjV/lX
LSH3bg8gGZY9owlvLl9sgU9UA/1IoNQZ1yiwmDFmhjjI8uWoyGqoS+YSxZ3/A6mgGLTDJaFFRcNl
38ODTH6Xy0VnIJWn/oJ06cqmak47ypJ8UKjUye8fyfWe5BtbLCOQQBZaSSVmcyCtOHnJBxsdYbZ3
BiEo73yddivDCJT0iOAF2e51f55Io3nTM5xfS2TCnCL9o5tz5RvOaQean/ND1M87kvykUcKnB4Ei
lifwzaJjxPDM1nFanMXgK0nzy89eY2Won0y6n6Je8UhmA6+sHcFkp8HoJLzr+282zJ+59hDHVzC8
keJz8QhOTMK0zOnB99M9rF9GKaSfvV6YztY/4rcAsLl7pytb0+OKwPgyygr0t14yrbK6wJBv/TR9
ZoIJZxcNRninH9HZ2hsXI1RiruUqwsDlMhLNaUYEdZPd2LctVhsMTpLMEmoUD84wrG8rxbDWoujT
mi+nUC0ZxQ88DjGLJyanohrgRSo7rr5FA/BHtPapRuoEJUvHHonaa9+llJ7qfAZ6enO6El31v3i4
yZQcvcB1FXUWw0qbspMShnSI3KY3wIj+eXGJAbE28siE/Pa4wDNLqfpzKjOh92EEBnbrbeVzLLRf
RusnSp4ykWkxBVqKCS38YC7lDCmzs7uMTCK5ibpuwdnwa6YY4KYKm4UzRtybAD8oFMBkQ9v4KMtT
GE71fyPlFDlTuot3mfBEBk+uCi9m5NtAZCqqhxTetVMxlsoNTUEhZ4Yfuu6MBLEtz+5FPoWueTUT
h0N24NPVlSE2ZwhtQb65mzyV/6+H0F96L1WqxNo1YKuBxFluv5UnRbz0/XWU2zzySS3n8C+Ht3QK
VSlS0MyTAYlox1SrqbqdKy+ycT1PGe2S9zLUTRouRKBCzpTyqXyX8TGnFYjKT4/nqdrCBN+c5T/8
LP5CQtt4/UMek0WcOTt0xHMJShjT8bDyCPYuwXmXkiUHOEUovq2cs4HvzS7zzDME/AO9dxGYCKBV
eedckosmfd5/Gwv9fltE0Y6ixM9w4aVvs5XYfGkuWmqMlmwt9tzx+KfpoN2v4mA4hKntlkhXbpxw
KHqQPb/3yIkNc9hdDpon/q06+2RK+iiMeEgUnxPuQ/gUvtrRuPoHa93q/Mj8kjg7KUuAwJOVGm4I
Aczx88GX4S/YcNmqFYEfoXGMevk71hsqgY+v2eZm+g2H3x3lNtK1wdkHMiLRjD+5SxGUdWhMjjHy
rHogdC1/TISY3+K2fcnUKxbVcImb0u/DU2LwJbGAtzjtLQ3ZJTtxidpK/2QZqwBsB+YPCS60YQoU
LN4KKS92JQXrJqOqAYtJtN78DgO7QCu8ifaZq/BuAuiJ4jmypmPsjKSmVwB7d8l+fC9mlQhCTqDn
83hi8nlS5TM88LKtI4XACTolxma78coE6Y1Yh/jiJkE5WkMWF38/+c2mjIOYF9PAi1RTgkj7bPnk
sRntbtdPnueHQOJKo79imIHGpO534uDZCLgXxM0wP25kLGaVTBhpnwcvhW+hlrI0/pcitf52ExNv
AYLMEZ/aE1RaA6l0gyfZ5XRohCN4hm4iqBA1Qoqv90FEH+fENh3mxCqNoIu8M7Fc30Bpl0Tgnv/U
pE8VO8sronTiy1NYbNzF2g2K0dVY/0KziAI0L0vYLJjlItKzgtc++sSxDV7OFiMlkdq2CczZ/GAp
OTrvdUZex/mv/rCsWa3XQXr4IsQmF6IO/t4zpKRy4M60e1+Vcmr5JY7JN8ZYqKFz/C76owjjTrMV
JTtk6faor9ZQ9Ls2i/wMapHCK2Xb77F+hC8AkzWkUZfKGGHdbktSXQ4cu4+K/Ug+dxHjXhsCkCb1
kl4bzDfMy6BFbcr0qMEffgP46HX7nj0JW6DaNj2hOOA0HapYlMiVEPfYau7UErsPUdAg8dUnLI5F
dpi4uGxkEUTKK6EKKt8mz3PHdhlgbCI7Vh2DQ+6lSJbaKSs9li4Yvm0FJCE4EzOJ/4w1aKTx8zvh
WMTGKUVOCliC+w9IbEIsyjeaXPIs83pxxQRrPWrhGPSqZp533sr1Zea5nLH2c1Ia6pN551KlTT7Y
EnrYrH56L/Njd9hP+AVx6YkQuHm8giK29oqLl+Nehois06ZPVjdO5s3c4c7ibOncJRRY57qvEeh3
uwgRv9tLC/ldA5qEA18fSFutWjJQfY3TbGs6oCQTRTopAYjONftG+Sx3S3qsa0X+eb059SJpsfaa
Btl0ueLtDsd6/ncfie9WWz+fx2uX0r9ojNDdMPNkLqPiPWQ6hoB4nQu+9ROJGx7Wy7frwP0oe0QU
yhGpGuKmi961h9Pp/ps2z9VzyxeMOf9OsatwVJ5g0KqEWAhG1Tal0xF2AEQ6y0G5qA0llwk7GmMP
zIC1q+Z7Bmdyk0aitDo1Re11swCHatVlyzhCyGs0aTbREv03Gvk56IofIGte6c02Gs7f5sFDFTqP
lPOdfM4okrQdO2BUJJqIa/uAj7Yr6Vw9Y+YEW0wyL6w993CX5MKK511uZWLkoohlO0Ws65pRGE6X
OMkAYkAtDRCVRjvaW/fjL0cN9GnTishwpchAFfFIcakUxqmh931NtAlb/k0ZDePBOxzgpKwPH0Nt
FwaZo7aRNADxz8GODR0Hq1SPV5VLLcVeRdmSBFjscpdyVZ2x/L90s5o5vaYxzAVXN7tZiG/7PUSB
esigADn4+YpQ5pV2eBd1H5UivCs54C6UK0sayfDaXGkQxzDSA+dNOgzFfYw35ZJUGQMPjrUWd2Q8
zznDJqZRs08JSr3V+bm+Pa9P6lK0nC6O2XqJ9x0uMr0lHLJutZlSF7js8O5K+V5clUVO1OaDjPua
GAwFFxj+dIuaxPDOuBGAKjscKyu6r54Losi0RfZXbeU8/px1aAvr/5SQDlg/tyzlbc6QM1ATp61h
btiqtC7JD7sme8bOWqntfgAYCN3CBCJBOtz0qTYeCAn8RxmFbyeOkxgYaLjLTBNd7+a/Cslske52
lUTZlyZsSgzdbE4RWbvBat3eAdbDFSoD9qRHKM3/0uWqcji5yJ6XN0exk7ieSjjpgn//amGoOZxj
UFErSe8jn37EQPqFbOZwcGOLZd+5VCHw7sM8X0jx5vjBbCj+Cm4ngWhyw+PL3Lj0E6gx13qhOIEC
qycvKzwgx97MWBkf+YvnLYLuPzphAJEgLltyIlJd6gDGDchJ4phFF5dGmzQWuIMC/9GxCA0K44QA
ZOOm4DyIefM+LATEMY2QHgqhPLA1wb/OaG0+CuCfQkvOI7YCpjNT5+dV9/LPytcWRkkQUy+Ta7TV
pb70GO6zdTUlL522eQPrsKrLOB8SQbCT9JEuGUYEsDr0mzP4k6kScEHwpbOt13K6/KDa8MLNx2Wc
vB6EUbGfWWyd/qcueL4+o0ANtL/uLXbKzunFfD36bT8nJiUUVOZjugEkXfbE+9vrc5ZqlTkdgCIM
MxH0T248LctfYQ1W5EOE2keEeDUrnq3QhWtHUFqrgn8GPwtTb/QUuC8d3p1ZQrG1XP6CLw699Fw8
OQohrxyy1LoLqPwQsIRtRST7lUZpAtO8gd9dKZ8DJeDeTZiTdp/Ce4g6ieohBYNMyXNjmfO/X1jC
/ynxQ6+AGzTo4BzhNLXwrUJJjkg9ERG8zEfsSr+NbeZcBWTeAn2QZYiWw0vArw/Jgg2dGLbz7lOl
AWMVVQ9OobsYacM4KGHzQw6EHvDkfLBrrrvcbqNkROdnH/kS6wikHDk6aE7KENO/FWkn0R9+nAoh
qUNVL789Ns2wAjl0ZFtCtdx8RBHXip51jAtme3buDbJoJ2ovWv643+OnMZ4pQD1wlnGDiBE+XQyn
D7dUAU2dytZiALOpTcl7yXwMxOiAg4wt75VrkbSbdkLoblI2tYDmHlJmAnuHuNbpT+dv0raZS6lY
eQAlA81qKjPm+ro8z/n06RXUEV3HisKKVvM9uyayOKBG9eGQbhckC/s2TsOyWwlrJC/v3cu4+DNe
6+45tY2ZXixZGpTOfJK0ROYWT51Ain/QfVXXadjs5it4hhSN8eAAP180H/Fie3nTZPudHhY65qOr
G+FviJWK2K298OW4uGnCaw6Ps4YZUedRbA3S6iSVje0gX67oAHRzkAkLe2EYkQthdetRsM4U2q1v
xQ+IKUEAj66qMTj/hFBr986ts8GF+cvBw1rlI7yrMwJnDvJaExrE/IBoIEk3KVhE98stDQtMpIss
uznhtHdBTMXNmrjqjP8z8cM7KCvm4lagAjKFkpTwRhP0nsPcD/2SRAk9FmzHxH+H1+I5HDj/B4JO
QpWb6olRHV62RJiqhuZAj3vIwkZ2wtYdqQnr/baOhBJpkAon6Gv2qe6O9e3Nbpt2fpZHNsgjR0Os
x21v8Olinwsh6SMaa+DEKUq6JpMAH2Igippr8DCXLFRqll283aROLPjkVeI429v5nfnQs3hkUrED
jQbCjKQLBXTQu3PM8EHP1qOjwhnI9V09YJocw/2nq2tnGrjW71KCQ0ag4+wR+uzu5TonVM1pyKJd
FqBWmciaWRyxX5QSTjCHVXbwt7vLk0/RcDA3W0fPcfOPHNLrFI1r24XoufMHpbRXovZaHev6DcGE
psFNVv+oK6FZaI1jYkHhj3GEoQc9NHxN51jww+5kPbH0zcV7aIs1C4BJF+TUXL4VOFhLoCkSKt7K
rWAea9J3rxQEPL1QruIDfpOdukNJTHuZrjDwfhpF7YpkxKihsJpqPGnPRll5KswGD5UxmMVdYIkx
3PvedA4FYBnuujTykLXVgccJSeOkE5XEh8O8GZJZHywD92DThLEl1b5928/Id3KlpI03yjlpe0QT
m8Ggusu5e34BUPVayHDdL844T4IFRH7gu8EgmhcOd2rbH2aEfF3A2t+3A7xpfDUylcCQiUWPOlRK
vZ+DfUk05mrEyOPiRLE5HEyJQGJIfuhN7uHc/w9DVXe9GibuIRvpPcDt9+oT0BqE9uWPuzyz7Jgd
ex6cS0Jaww+/WgXaaD6OnJm4JAvky9KvVGsqh5F79Sra6E6utTzJq4DZHtxTXrMCD/eP4qGpRrYO
hWo4IuyD4O/Y2bTGaXd2ppnLiN17S4SOXzlKmzyppLMJC+EV+vwWU4Cd3F0x9sJ8HVZ1XOYP9rGr
SB32aq5mLmr4/zsUo1Ab3tI+1LgdDsBs/T0Bn6d5S4BJuIq7KSLSiViczHjecxAWJZHgvTlDSlIC
AAwVueddj+CPuc/dxOgN0YxtgR5lRD0jRFQl6Rf88g63a1AmH8Yi0/bQee6K4qQIBBruGEltZkeX
+O4qxTEAkwIXcjqHsoHGMg8/36eMQZUq8vxapnNXmNyV6pOiZCpdD2YGSF3PR8wf/vp2Rzqan5E6
p3Y7hJ/2TKU8unjDgSvLzhESd3mj1A8lvqOllpuueNW7PTTqcDd/TaFl8NvVbRBie3Vf+/DG6fsr
hj3cTz7vKEjWPf8dhmGj7eDE1JSim7doeL4ngKm+WDQ0VqHXzlg6YpTVQngCwCzHR1Q91osD72C0
ssuJLNdNgsjQXLIa3uXSjbnAZ0hI8sEeDNdfaneuXqd90xSJNyPp8rdWxb0ttnnBxbe79ftNqOd4
MEhJ75J3v82pLUzd4Eohf9DnBOx/iy5Nh204Pg6WAJsjef0iQHqv4e/0Pan0/2F3VeHpjpa11coa
xFN0ZDlL8/936hThGdTQH/6FKbF+WxXi6sHF29k+pwK6ZyTcsc9hkQK2UN4uG2n8+HZGKIZr3vvk
jruWl1wDpbPTdowd8TMvpmpeZOpmNEdL6xZ6d+jCi0XM2Q7rMpAQEjaPzYCERO1P/m5NGE9fVFio
3+3So+ymUqZmV59pLE6D9U2I2r4vCndRQRox77KezoJ/s/5XKlyaPQ4kpKcEPklhKHwog38PeM9T
92FqTDq/B34QTR3S0wsfFHzNr8Ghnuh/EK8k6oO4IZiJN7SzwOiAXlZAhoO58izzViTzuaEbRpEa
aY49OxVN3RgGTr4ozeKBppN+kyK6U8LQBJBEu14zNjPBE8qvmMU8pNXAFR9caMOj5TE0lr10MkYM
ZXAFQuGbHUIxizhgZ/AKN58hcnJx4/LXH4UMtxS4f47Rox+ZuVT0rZUitUSTQel/56VacX7QWTGJ
QP1xeOqBoD62PKQPDzvsxfApepS2SFWQvld6laZwBriB1hBAISjFUBhlMXeufk4NmtPKFuwjAThh
KBC/b85BbSkK7ey7okx9RdCWGKaUbk/WNfmofT6ovE8sR5EMSbaUHjyrUS+ESnpCTDPY/6B1ObkH
bngLAIU5d+w/AVkrC9OSoKlEVuXHlkh+/ty8hxY0DSCWdX9ZaLpooBRsgo1OXlWt1is53gM1aS+W
bOs7oV4fYIq2sni175Y6CTzQueK+qVefUmJ5drgOqtiSRPIZrrDMfmys9UdGX+l1RkhGDcMSHY79
wtxbhi8Aodj7DiMxfGK92M53B7uK6kPXhGhOqzNivt8OhOyD+Nc63TGMPJPv038guLRI5eJ6GBdw
ETNv2BWqnHQ5hY6Vrc7GEZISxL0iWUAUSLU7cycnLBGMsLBuUarRQ6HVKWRBS+vPMtMgI+9G5dMH
3+kAdKG0T0E4IDwne0yfGelxGvpSxcHaR2b6fPBnJ5R83Gooz8tYGwhZxoIYg9Ieh9meQ3xC/DJ8
1eaY+T6BZBCcKSB/AN//T988kE+sxh3WfRDSO9nEy1qiLzpo4mPGGrsK6lepQ5RYr0CnJfxl8I0l
H2EQbNpoYZuPoII28/SB0ZiU97xSzbvqqRs9Rfw148r5uyjtmNeMqqNGeZ9fWtebYi3ttNJ1KhDT
Lo6rLpsu7oMl+DXoiYDMB/KlzJlKhXqhIDQj4koTJmjyW2rMFm1aVEQnSCMop2jzLkOr4zKAXj2j
I7B1ro13wET2mCKqTMVwJyFh5jZBQz66TCxAWOgGrmXip6g8O0ujGr35M6vleyEr2w8eCisUlXNW
oS3z7oeiMIrmLma7Qv12daDYPApP+wXTc23ZmGHsQQsI4y8/XyLYoTjF0yCSApAQWkv23Q5rVGG0
GV6N88USogHFzdWH5aV4y/lKKz0Bn1xODPIQErVT2n8ASgXp8CmekmLAj4dPRROzvYuJE8xwE96/
EQax43d1VXVhMw4/UVDWlaXUO7PSpsbWaalsP413FTqtB4W9VyhaROmTy4EddUjDFGRKRiLeNyn/
HALDbsvYJP4uyU+Fn70QaN22N0ez/8q/pfH4zZ6CrX2JXIYhRUbab/V3yPZQxSeGDW+Q2e1cUIzX
G9hffQuXQSOc7dwSCwzYQOgu68WJm9DRKXlTPfj9be8T/5+Mt1mS2ajQsML08exmsgSsSsyxqISH
vBoz9NQPrF7Zr1yDCyMhHCikxZuOh+miKE4RAA/m+xadVUWMQwmYZ1wxvL2/dVo1VGqHllDDhl5S
tScxvW6GnpnFrUJ60Zw6q5h9kgQ0PGUfEr+ufDNN49mIerBg1eYcoNKzhZn7MKYEjGagkvqqTK/O
EGKT1qNihJuo+oFWSDB92+k07S7zz22hzSPhxWjHKbqk0y+0x0XkpcdrP0OU0IluyhICHNJ6kK7k
Gyzu+OZhA20ZrGBXmwopOADs6+u1vUXwiBNxTUNCpxYBWLpM8NIn7ZjqjCvVObzd1MLtgvtKoUiJ
3almoflH9NNEmm+nnNq3nxcgEQe4+pIiUwJQ8r4UcKAjtET8vfkT1e3n4hXzloN/Q1K9O9EoNzhL
R473hDhKSFQiNMJ6+P/v+RN2fiVqV9NQ72GH5XDcNp+hv3zC1rrq/lPv0sjCEqmU9r0HPLWgr4Y5
oWZ+lK41QbRjKqcq0GVCIzaM8ZthLbalnu2Hcy2KdSI7FKWwdNSkcsCAxH1XtuapaAMMGGqWVoIv
igmKwv+2KB6z0XugG96ygnYqMw+iSS6R/PUY1GQAkNFIbYTyW+LKFxIW5kS6JZ/p6ud5CCHgmbMi
d+S9yKfamUBJj1SeYRYlZ0fj8112rUsN7/tijuTY2u4hTy8Fd8VNaSEH03Rdo8fA+UfXR5belmrP
jWljrdOjEhZflaRCbVlK7XywvS4CHc440cXHn1bz/IN+GXiEEJaCcYOpFFRysRtr3sIAaUABrMs6
j9UwbsF4eGMJp0kErS7FKzK6T7wyVVV4cV0CZpPm+HrwPJ6uEwxz7V87adclzKPB0j9He0W74REH
79dPSiorvkJInPgxubATQt6PFZm+iScrvT07ITE5KUmp+ShVkrA72etKzMABkRWQiaIEDY8m8N4x
HJ7SO6zt12numruBkB99AHUHMdJqR6ScUabf8sF+ArXUfOqtjCMmOgBhlZResStL+SaLNcPqGokX
dqPSuInURVtqJt9ubt68SXJen+q76S/b0fapipqCoaWI3aSiibBEL8PtBZGzLsnYj6wgVJq78yIK
yoMJVT+8S5j2wyM15TZ2kS15GF3wH4KF8xM0i5A9rGnG7QI2jwrBB4VcCA4q3QHK5Z9gIhJknzN4
fHRzdIZZZYS1nUsDvzXbzdJVKVmafJI3JfzEJPF8eyIRCsfSNWHbgv+K8Sx0kMDf8YB2dxHvRcVm
01H84khJsGDOXCttrTunSzZw0S6wSZTj7Pmn7XPJSVuPrxb8mlETZe7unTcyst9aSU5YUyUd8Eht
ZwcSRH7W2598dmJWGPvfqneIT8aRfmrAqLN5ZROVsdW+P/1ZbUcuwqVw0053zIPK3Tbhutg+Y9u/
XtAe6osV7FtR1AXHQCh6Njl4vzyRSU8+2gBNnij0EJYvU6w6MxXjv3loILnCBWOtO6ld4izf6BhF
EQN7ahI5r/vhO8wZcmoqsBeObjfO5KIkZ+uAr5asP6gMiHVG1AFYYYZmyXCL/tPVJRpcHOd0uXAf
jQKA76vOosFRcAs2HtX8gKMVXzsSfP0wCyBw4BBz3TPiFndAIBv1AZUU4N6YTL8JeOlu/JCtgkxO
At/GtJ7LeozhraDCrAT8R4L4mGTpPCP5mZXElPyTXKYxJ0jy03JBqATQpeH+CChM9YQB1ZN+izpn
TZQMM+AaQkfhG3FR7TtKb/w5u2bGqL0rscCAHvH4NTS1FynqtqT51zpd89LAdxxRZ88cmQCiEFPz
BsWdkMn40tQxcqAVw1KhhgFbdJ94r8Tkf9eNbVf/Ir4ZqsQIt2vNcuiR2b0UJA2z3JTPxhbqNZ6T
PLX7/iYVjAJh9UBkFPeuo1BOoFYyhuJgrf9P/ov8QoE65MsPdDhJovuBidX6V6SFrsjuFFqXFFXw
XIrryeIVc36zxH63rxXHFqSpRs61B34fspfsAsErEMDi+/uxc68ki2jA0RrwDIhr933t0IUeoaHn
8/7VbYOS2gT0Cz5+rUgZ1BzGGKNM/p79qu97dzu9bmfev55NXE3xXz0Yr/owTd9sq2H/i+xHo8n8
klTnuqbstj0fB162zK0xsEltGlEkM/Q3nkhQdSHA+3dPG3cm/ND6VLOI83SIwafHALh7Bxj4CjJi
gPn/GR2XTaoolwMsOkAxj4wR4udeWdfyVW5tmEPt3O2S2DMPotsqpwu0baL2uVubLBctfDH1A/65
0MEEm7x3PPzn8Zca0G4Wa9RW1gPXOvIGY52JOJ2Al8XAK7X6JQMeKP5nZULbcjohN0LbhKFts82H
6uR1kQO0pSHKaoqJY74GXC63/gZEzo9S/Vqhn5Z1RxizR4+135Z05Slvcq56S+hRQpfsfVMCkvzG
gd6Y0NpRrgKjlmhn6cmse/boDYPp2v/V6W1Y5WAaFDAidTTjlFWP/vcmQO5KGEPQjCuOFLyqy4e8
3kevZn3mbd9vWmFIij9c3SlLaZhdxbSSkVtsgqwU+TnPnty5Wd35vx4ZvAdiyeLV1T+LkZ07128X
d2+/ysc34/wfhtdZc3dmjpelmIySDju0hlAtkmhX5wcM4pesb7HgOdY6yZou6r1Z/ewamHhYPHOs
9xTSoJRwEqM/2NZ39FbO3D2/FoEmXdq32eoOtFg/SI5xGt7U97ESMOQ8CkM/H+y2PET9VK3L2kNA
bie1EgU+dcq/ZmPSeqyVzMBZuvjOBnCtf+QjoIwExV68i5n6laPw97yZ89NVfsV5Z/eBbVu2d4Ei
u7nlWQjfT75CPAJUQqalwv3ITUJeT36E1fqqh/Zi95hX0bFvbg9LlRJYkAcMvCCEL9lXHiipk1T+
96vh0HyT6Pdd4ULL/nkKC3aNtsBvdJoh+5babnDJm3JjPTYrPZxjdzUFBzjPL01V6uFiD8wufcVZ
cJFmtVXQttgb2h1gpO35CmammtNNZala/ohmDSEcqKB804eS01dU+0zRWHK2uffI7NGlGiyZCRim
Pxtw8seXpqHuORE7Z5k7NZwpuSxvvR0pv9/MH9RNQzkVtqauLwK/9STuRoxsOTaMmfL3wywh0YiX
TlvkcVEcyQQjHUVENSYlPgMYlmJGkImElteTYAGOUNWd+BusYfKpNDaYo83rQKE4RY3YwiknPRhX
QHphPHG43lehIiVi0ob0FsTpOhJrMGYnBAT2C3Ore+3UFG6Cdz5gcRzSJvxYmjJD7eZbdAd9wGVU
/I7nCAeox8JWt1cxLrIyFwP9t/A1OHJDmr4KqJ/IPI45yvcRqdYd20ySuDfDQIZRZQmNKOFM6KqD
obSe/ISiKJ9oFNw0OciRWLLpNZ6ldq3SJYDCNGH38G5Nze4SyU+eVbJvhKnMdtBYNLN4CLenFRZL
vOzsaayKigfcCw4OtIBEsCYC22qhfCEO6wW6pNaakuMVm81hOHVGbbbKgtHlTRss+K2r6fBh6DSg
KJt1iEBFtgL2oxbtNTpuHPAm0o700qIHtOoxH6Zaf/hwUSrpRBD6hxi/392AROPN2TC66vwnJUgF
8Mde7UzDJ6egIHbX3/qY/D8Wvh5YXwt1hG8G8fo3eOY7OckVF4pYvOi9emxarCYK6X/wRnycOxQ+
QM2i65EbTHFjrvsMQc+AMGabPH7D5VdArDYh0mNE/jjHkQfCutZbpfJR5O8ESfdr5benl5v+CM8t
gpdY4ORoFEtSYisPGXE4uQzlqj7sbm0LCvlsijnH2Fz43d4WUuFdbK+vvDZi8Ny0QMUxmcohXDW+
nQL9kQEVKAQZKpl1DE0aYBZmCdzy3aah/HJl/jgDWsF3fhS2V3n8BDMk/edexdMOEcEgzDvAZ/HZ
9dCYZErI8ju42ymBcx8WZny2N6nYoQZsPzuv7UQnhHlXDpuuw18GrPciCThQ/B/hK557hQSFS8rV
d+yj9jRGQJbWYlngs8SR97sYiXdzzz5dxUnEBWBI4LtgMc/Swi47MVi5nzkASNCKRJOWBfVecRpZ
4RsAryPVDSsfH1feAF3XBD0zq4txG26vIWipwZdO38w4h8EOWsAtwwGWTypKKlI8hdS/WxpNMDrf
v53LdizSbj84+119NrZyGnDhfD6d5kEPRBMavYYxk/DyGVz/fLXJVz09wtj9Ck9yX5PahNlldaji
/AalNZ7vtmQhewgPvcdPCotOtUDEMm/2yjJprb4ghXr9eVt23ip0wYpu/PL9inrannSQwo0PjEt+
/X1r77Hj0rfzM5f/nCQRpPWJ3977wLPngLivGdgl5ihxp4bpxNphIYw2mOlz3DVJ0nCskNR+EHrM
1S0CWMz6+rwhaxy1+DieazFi+SpJbkgTibuXBib9y4224OjrbNAAal3lTLImObZvkl/y6veC42Ua
563D5Qa/sOm+LH6SOkcMO9XdX6bJPc1D+aX7xyPzIbwexQbyHUX3DVMx/eHJ4UI1KQP2Sd0hEOYY
0NIYTTyje/8ve9hAeX1VpazYsn7obgFfxMn3ueCXLvbYZDy42wYy+ec3kyUIbgwe3SP8aEHDWG/M
51MOUOL8Fp2Ssxly8oSufkmTOvkhH9/RnarGThuN6RhidE+9RJjv/WgHxu1iA/i69BcLcZkyk/aJ
sbiXValBw6Y43Ob8mTu+lLBpGb+Ol7qcMBsB0UPwGDKA+kpsAOMed1yDYjKlT29Zw+88lsr2zWiP
ZkJbV7jIw5XwQ3nwNitOdAW9M4+7Shp/R1gT39OzEKwPFAWJ2THBvE2v91HYXUKMjjkeo1GhPgBH
ah2vDVGZ9+BtMGj8uJ22XQ3AaVBH/CKXb2azLa+LZJ1b6hCIovdkZV9Kko9WzMnYj5gpLRFRPmoS
Yq28DEKdGmDldhGA+NN9Z3ugm3xfVq9TzNcv/ijG9wVNjTyHb+BRL1siZnijZS9uSZ8M+x8LvMCp
Wa9x4zHYM2m+QsXV9mYIpJe9jJISaA2hsvxJ9gku7Giec+gFCiwJHwAs9ALanqoPLQx/dGMdDZH3
uxmiyk9nO0BR0KYqCoW+AHrtqBbQ0i3bOfPkMgSO5fNmgy5F+lxOCbq8qCquYOPbrh0l6pBcCAeB
7XutUTztC1oHHDzD8n+9CyKNMpEQf+KJmcn0CAkPr7T5yaF+7aJZGaw6LsIFZAUOKm6Cl8NnjBtt
ctHkoeXwIXsDUwdSMHBZQYDMW4csxTyC+A9skgmzc0C7iPc7ppsvlQTC6/2D1eXvZrDqGd0Wda8w
InfaPTypZWvqPLEb+2JZuV3dP+V52mAlDpnuj1rjuQmfDEJV/dkIwk3I94py5cwtZktmJ7hBqkrR
wEEC9daVgzi/4f+dqN8QQLHQ/6snZRuk1u0FX91cxZ0BF37mK5Ed1MlIxcrZNnafhp7qfr5ROBm2
H22wMWEq62yCdXddMHe8d9P4EEzTGIs2cEEv325AkYboyj5XvdQ17juv9rut23tdAzq74KA1Nbdk
kM4sTC9nc70aquPWyMBTPUgvlb8K6WLZieTn4dKbMa5RvPk7R0C7TgPV00ESKOZGZ4AlTKrWtIBH
2PxAoX4M3EITh5ujLv+s+IXfhje+zHD5kZn8Ve/D/iIQBEC52Pbk41/It8Ks6twdqxc4tOOSGdCs
ha5gSjJKFuKxEwq5Epg5Dg1ZRRrrjr+kvGfRLoJZEChwfV9UH2igXgP6UDoKOHqTxKu/fILiNE6q
WwmAI16EuU94KRxmnjpe7Mb7ozcudj5fvKS31bv/sJAxJyYbi/Di85SGR6QVDnXi4c/2Kl7hOM1Q
t+LKegZlWKI+Tx1mYbdVboFlDh4Yzi5xIH+uoeSeExZiqsnCY2b/eVtklcexxa6HyrSD5DYEmdz0
Pmk5c+xHBR4k2RcDfuJfWpLMmo/cEgLpjxM7Eg0EsNpUKbc4gMmKBISCmwCT06eUyAPXiHgljYwN
1LRa4WhOWD5aa/kimoy/xwhVhNV63jwEqz18qSd548pYUswVbm4dgncTwbvGrJQMa3ux1O9y8lCz
9hxFvAhUF7guzoAMkt2KvXN5NvI4zdCNQnu4VbbGFKpyETxlAsaqp6LqktoKkl7+WokmUDQ1U0ao
5nDua9iSZ5v+4Tt+z0REx/iPnAJRZvq1ZkTFsTxCPjujU2THvA5mPRjRvvQfIDp4jPmQC8KzE2pn
febBJDkR/3c6UEmlQ397hN2n43TsjyNNaYfPMa3teKkk+EMakS4rQq93Yty0pBnYGOxYmda32+IE
9H0qesV8wXlHAPHRBDM7iRP8xZYHAXSW0RFUZdF0JjBKdyAGAwA22TRwBN6j2pRRXb4SAZLmEM4O
aGKCCg8qS7lDoGLhMQz6DCATvA/Rnwjxw6GrbGMECI6huMMwGmd3xDL+LIbUWodcEUUs0y2Fh31D
+ajp3TtBzXGenVsU7sQvfib03fB8q3TNc0PoZ1L8rIyJxcGSaTaLKsRzu40CKNU6X5C6h213ou+/
5wFizWbt2Wt0T+guocVuPsPeihS8a7UtJyoEBPtIHrZY80BG0SCdux1aPhR3gpzLzYMVlRdFUyk3
+a43wRppx0DAJlYpn4kpVOIV48YjUg+U40jgUWUvyhfvFXvq4YC40dEKWjKtmEUPOEsHZpqjmZMl
cePDsMEgMNjc71CIcxZFNDsBwCNUNrk8OtUQo/7CC8fZfPhjVSe9FzrBAD3YhA3CfeSyn/Sjiv1a
8GIGHeb27kXYgppcWBWZG8xDcNa3rMenHndx580NHOekiKsk+EjwDZafe3hK3wMoc6zmk9WCNZFY
cWlUU5FOlkJ6cFZ3BaUcrcYrlaN9W1mDVSwKCKNuXJLbwiBkbMm7XMRBVorcticK429FLPw3KE4N
zBGVbD17r4MFoFHL9aARXW+3DLe99e9jFQ5kxa7Rnvr0hPaFCrMuFD951PFac+G9ipmJbYqoWRFB
mY72anvCJClaSjM/RifqxTo6nU7H3wiEsyfH/A51kzpnHWquUy/lxz6EB4MXBeHWIlmqhYZgAHpA
EVeLAqYurT4dsdKpcnulkx/M6yUmOOgYAtBpigpypgGhmT/3LOG9AzAWg8f944v8vzKeCmQgCOvW
bNOXPqMaQO5b+z7zS7/4ymRVdFeD6MXzYLqlKsNk8lmgI9HyBeA7LJ1OZLWiKULCCk21KbNYKrzy
5rcRFkbCThWgJ4TW+Ncz2zn5Ssv2yHfZPy6r1NLM2ySaYJ6zV7jbd+kZShItxTJot2qzZUTPgi8l
kCT1tNyRD/+6fJQN9MlsnNg7mnSsAAWet9s9h/GNHkKoekOg7bYt+LHsm/1YFNt5yH/8xmw09zXt
JG/OAT79fIBi+DnqDH1XDmXEnOQC2nKGzmiH0gAF9nhPGu7j1nTrD6vpfYmdT2Jv+jtUrFPjBU7u
sJDH5JDkUA7mjnZYzjd6n5fi3jslKnBNEO+uSBW4FCv+chlCPmqgH3YfQ5qfqbKygz9PcoInhHm6
sjO+IE4KMn8S03PrEUOyg80nS1g9WbDxYXTXBEfvr2s2+0UlYvDqmMqNMg+U+2YSaqllIkZrcQa3
WhLRnOn5jx3bKeRFbCN3Y93KGKeh/zcQxEkATyFstuHAWyFBlU9N0q2Q2BQZLNFcno7iI/qqG06O
RqIIiulnxYpxdvy60fMHXT72WSxW7IOvTwW1qSYEemGdAajoXBrclrIV2Uvoo3zRODcezGoR4mfw
+wCdbQeljnLdY/Lpt01q3078WLRWu6ZM0nJEdQoLz5NyTlbT0TtPpDfMsh96AsKGOZRUdfIjY/0y
T20Fc93apQXLktGhtKzuT2ql5M4/b4l1DTnB1/bOiJI3fYHkel7AkcsxHhzE2bYE/A3U6L4nwZgK
eeEl1rijHhkLg/Bzr2B2MxekDYXpTLNVpDswClWAW0NQ0SOBsTz81qDytFuU1feJ1hcCkbTxGksx
Zl5+0TwGCp45iyA5GgA9uIAero8equ23uzoR2DkIPJO8hswRHD6Q+kO0WJKr+eBpHIyVci8YQswK
0q8jALbLmPrutNqFDBfTSEms+c+AycuEs7X+hz4jPGcX42Dn8UpSywSUW3RJEa+SduAltkkttHAc
gm/P+XxjU0nfEoqlDaDQvTgq5f4We2IwdupKttB20vmFFZHWzr2cn4S3iiSQJqTFDUCPHPjUB4Do
Lj3PZWuMeoqvWj7GDqpH/AdAB0RUzhJCnk4YvADG1rcbWnUXbMUbSQ7AOs7S25t7nre7LeBP0egW
/IpGyk4e1saBEcAMESWKrb2e2J2wOqQo7JS3/X+tuivGqbJTuOrJhoxRKVEmwLujn37TXUyMd6fK
pzqA4UNc6fHKe5d5du25nsmoBXNq9B9o8rPTeWPo47pVX74A0RYVscu9PruEFnxae131q+QDEAZ2
VP8HL3bvVkPIxrWVM0/wfWyq0yiV4wLEZSNcHXupXNU0xjCKRwjZuv6mr89AweRgR1dkAB/fBQCZ
Af33D3qwmLA0hrySqHeykdgGS3Q0sHdn0Ed6dwMTBYIfVv/0bzTEK/+yQKudeUllynCXnXn2iOmI
QFmQ7eMqjUqMXlvXCMVSuBdD1Z/gUIvyA/Gc27RMi0NzlyN8CH1oF9NWuhXIDdDmnUbgbPj0mlzD
VV992BWERQulsTEN7Kzy/Ds5KqRINfwVwU12Bfl40FPVdOVoKBjp2UeiVz4fd+BwMiNWQKXmhaqm
4PGXxPvqA4C+W4LoGUVCNUDzEe93vU37EC4eheKON1sJXLtoRvmhW/2AQaIh5po9lOJpOg2TD2Jn
Jw2+dXCivEbADo73fpa67jibsLzXp3RP/CkuCZ+vSoZlO551lJm1MmbdQJEneY/eo+g+RlAfYfjB
Ka7FN2fJp4GtaR9d02FVgjzbGe+cREgwW3/hKnFJ2pjgGSl9Ohk4bbVc1TAiOYDvkJpwQTXp3hCR
jXbeprv0lRyrV+yrcRtXH3taN1jTshBq6DfYfy47+Pfc7ltTgeCn9hisGsPCwKF7615oTJCYx0cT
WK/k6nEkPQbPEQM4JHDDC+9pWpIEEV1hckYCkpfs8kR+FIb3JrV1d635kQbh9e3JOFyKzzEgcA5Y
giMZwHF0u8SGcFzHOTTbh6jsZdGkJi2DuS1So2+0YPiyNhw7oOw4oiH6Df2bG8MYxpg3kaXjWInU
GOUZX/UoNKapsv70uxuXGbwcH4moPqEPaeAqfotSWhbMhsuZdU/UQ9i1NYAYdzh1Oeoqt6fe/ocI
L/xd7AwkNq5r1GRZpgXFXNrRDEAL00KwbvbQXpYmB0F9VnBsEP22eRH+x6nwNtnAmJklwnnDPVAN
4E/as93NmrovVRG66Aq8jdJQ7IZTmm6YKxr2KA5WJqzNvU3RTrU2ik1eTtLAerqyPJbnSvcEtwTt
8ItU2CPRN/JpXW5+Lf/UeTfkAtBQf6WR36ikoVbKKvnN51yZ1H2YwFn1UVqPuxwNL2qsdZDKCzCc
VK1YX7kPgntLyDoMNY1uWGwYcPUtupSe5zZ41cvjEt2wqh0yGHfuuBNxPbaCWAC4zjSzMjP98Vf1
5OHU83HyvwuvB5zAV3MjA/pHbdoWUOzJzf5M/0HfotkEXe3/+haw0P+/g+HaK1wqdKSDIsekaoQZ
y3GKdwrh7wLc69LLpLBqcwyzc0NWkXd1M4NjxJC2haQWh4Bmva8pxBCC/9/aP1qVtXLhgP+QjseA
bQwYP5PryeN6XvC5KtY94GdCSSGbygs4ClZ12jGww2gIdh2c+vFSc6EqDyTq6E15XRj/KTYvQzqB
OZdJc67PBCVkzBGrkShwxehxIXlbOnWL0Q97oEcAsAnwGdSuCYDyVSG7ck+nhjrmZTeX4doHyuTU
OKl7UJxaXBpRHbmtwaX3qCxZa4qqeEX7zS2HeXFl44RQD2Gr2hgnMSL8UU/TBDVL/tdErpAopIb/
0cYkYgdSGSPCHeVBA6UAviRoKQKvGS/JBlvXEZs6PMVFxHk2Pd/FnT4wt8PmG3Inkpv+bJ4Pcw8U
v4OPMXC4PsMKgVG14t4G5Y8mKsja7B/SAKW+QspMBJEiq8Jgis4k2UEKECU+FptXxnWttANMl5FG
ud1bJ2dcCmNzSfSDg+9jgk/7JTPe7W9KGjw7yes5Alj5QZcf93/diCCzuRFe8TDin3Ueg1iF/YV7
RS6TQKpEqsWHBRP9Gj0gV0k8jMXu9bE7DTbeiMs/NxIcBCc0PonhP2neUZAXXjgypaj7X4BN3qpw
RiEBjQckclbCqhuz3y7wD8xBX4FIWZmx/Tp2jfaaRgJ5/7dAENuylMqAEKIbT+FSwz6sGKcLsy5y
yhaUbpZjeQkqwiCL0rC/qVo46Hm9ADWW9vwPufT5a6HYyUpEXwdlcuBPVcJNpLgf8bp3mHjgymTU
UNM018t03oXsJOQpbscH7G7L5+fQczK6miLfuw6Cr3bTonM/8O4K9NVldz5KPMLViYkWYo6cMyTx
KzVu22SsuweS4zukK4gpQxQlAQGn1/mj0tLeVvu4WeYwYVekAv1w6MAGailnkpXqvkWhJSNQUh/E
aKZxrhOooHi/IhQHhynbb9YAE5nzYvELd41wujr5xRXp2+yGtWhxnsVUQ8AiuonZT9r8mV783421
SWA0WQDhvslMlvcXkrFrMf49bhbfrNYblIK0kH+CkaBA3740/ZtlDl5NRwpBBWI2r/jqdJn1gP5k
dtXsTcEa7hIYy2QGzD6APQgYlhm4AuVIiRg02Dxcdj3BNdO9UBZHX12q6yPuUxAtKMAigntTdkAe
kqJ8btFKeaRBG4UtW3JjsqJKzQ3LPj2DscID8RMKuWvYuq/pwFk/9Ey7wNs1EL1qUh1HrVqYL/x3
KjHwGDNigPSiSYEhPcOwMCuqPLEzkqRpb65uJ4k2tWQBFzy4Yh5+ObNH8Dtl5V30dJOXiCN09+9k
dIr3Ld2qUEeU6RKKXVb4+rP4rrnHGeNmbq5aCCcZKiI7VjhGplFeH4q/fYp2f0G8I6OMLU6Q9MEO
+dELtlr99oVTfmWZ4iG2PuKty7WkyMk6ZNinwoCuj9IF9M8ar1RW4FkoNm8YX7yDxsw2Eq9+PF4C
Ex4HGtGnfJmXZtukOOd5FkZ4wBxtITXU74RjA8QT7/fWWJN/7bHDD+9FXq9VvuwGGst843SvPH05
yUsNE1RqfZRmq0Z6810Ux0UJt1n+JMsdunzPTSJwy8Os9vITqZgOEyhmtkp93+I8ajEEiMw4Ge7T
UA6rEzug/9F24wS416wcbQKDqzjCjEMig9iWdnmI7demTnBxQJqAPNGvEhUFy+Fl2jpP5tUsHBWN
hFMvJRhcvaA9EjQd8v/+YmcLO1v6IlHcn1XMR6fUtAOOitgYnjq9Gc6qL0ahNKHBez/4tL2fxFE2
W+/L4Jc1NSMV/ukuBncGleXRecn2FXllJPpRsEFXW7/0i6bvHOL+nTXjOC3o9JowLnpsIGPUtKsx
6dt65HQ1njtPEdXUeb3zrzw64X3JVjG6V5dcfiQFeZ+kBLNYQ0CODkgu+dLwf/7hG6oU+5QbIt3r
erWIYsLpQ/sJG3jMgAZYWZ1Jg0UQNgWRLf6qFi98obf4lfUGDRhmFs9Q9uqgwYcyqXFpQjYjg8hU
Me22L1dIAkXAYRXlOjW7ZR1ZwVManxpjjSAVUYWpNfbgIFzG3fprHSNP0VPSiyLy2iCoKv8/00em
iQqsd32m3LxlIcZoo9+m4CSIRikGKTQ4/R+cNJuj/iWeDgByoIM2GHDauqHMbXBDl7gpTmvrcEZN
VA+t/sDm9M4rF2OAMQ+sNcJILXIXyofCFkIi1LTfb/61f2zCqwIVEwrCYbeGzv2nympwwRZHEveY
IfHv1tW+vMz8o1JBURQ0hn7gv/jvzpdIZHJ1Q8+Xnb46WVTmP1og/UFBX/zHHD2Wy1GXsQ/K/FYL
GQodcNXHzOSrNe3ubJDFsDmC9PzrOBDzYdwuU/d8U2qIwk5JNrYDXUyDj3YnktUMijcJUVSiq0GK
4PwBX4P7RRB/RbVzxZAFadCWNYZt2lRe1KOy9zXjFh1ohlyuKvs8i+eNuYH5LZs25/fnyEM3vJJn
vTfCy8HrgTLast/k8jyw2HvmkGff46vRnwkpRSn98f1miVCBt8hbC6A8sWH/fddK07BOr0+8GlHF
t6ND0vgnc8f+vRiTYZ7ACF9PRqwI2dRWvwID3QvSMTKEuNcUIQj1Bpfyy8LVMiKwFYdP64XMpGlW
WrGgnCxEHIAfyf5aKXE/Oyh+UZkMUpkHMjkvB4b+hKYwBvskXKS9By8KaetXAoJPkjaH7HH0nCS+
2Xo9/WVmXXBlUqJS+jkWqyGtRy+ztHmbRzPwSwy3XKvgDeSfHdp9i+qN3BEMXXzrnJ+3xV7rchIy
3/Nmp6DwWT6H/XAhylMoRLoFZ/l++8BLOcRZWz8FwG2SC4dnU41Hj+piilky/vekJ1i+1iu6WLEs
KVgygN8H1pgGPxMwsolq6TmrnsqtJ+HI+drU2MOmKx7gSLZA0Oze/N9pJUoRIwpsuN1tM31s63HH
nZ28DguP+bTVoC81/L+kziQ4cDAISFmbj90pGEOqKMtxFez0i0o/cdPMSmMgLfPMoFeHo0W2JoBc
1SoI47TUF1ZdWruVkRSu/y0F2VPRwMPY8PB4E7jvuYv8DF/5eUcBR9D5+67jXJoBUjkd0YBerk3F
hxbPXz7+R7MQjawhmRXIbKAl12mIqWVZ7viO458cIZvfwGg98iob+KfG/RIsUK7Q7iNRh6IFLBo3
dColcrc6kMCEN6s90vN58nh+SGqycEeSGEuY+pNGYtUXTFgUKqgobXeSh99Dlgi1T6XNg1Iq/GC0
F3VVI+NzhHrXssMIfJvUcEjrrYPM0dGVaKjpUIg03z4TA413VHqzjSxuGHmAP9hnznlmJXzdWqBa
3X/X9F9ZHV1FID/95Amr6mqnfiY0p524mBCRzB+lYQ0tbiADEtNkTezJ4EOxNz/gsZI3pfaWmKLn
wBCbTLwd+9BAwE5GwvtS2wRmSgFCfCAPmo6qvau7QDofHbol4LCJoL8trufvg+Du0Zh6oxAY0e4f
r2TyKM9ltdaDpDbTdIwONTV2tPOOeNpENaZmoXeTAZxEOQgLSdlNXuJmOIq8S6FUtfPg1ORxFDVS
Eg6LrbIipSwqHEN4Ik+6Q4lvYK50ds0REYGjo5f0hAVEEQRAjZkH9pWXX6LOkUZs/a3nurfbX6Cy
30sLqqcQq7Qy3smmyl1Nl/I70AVahpAi62W2awPhR+aovFkhygjH+8dDGeGkvao6CqZtaAuVqST0
PWMGEEB0F7/B3S4vLA6z8injUhZ0XCFUV6GjzozHkUJnyWqbWd4YTUVLYbNw3W+qNpvbWk6sAgyP
Z6jhJdU2hhjd6K9zSAOIw168C/iCDrTnvE/asiQNWfScVImecMTxglqE3WDphj2ZRY2DOMPsrl8U
EH/0kbaTHpJq+mAgWKwnbdYuq3XMhH5FKHMwOYCVHv5EUBAdt50Fakhvr26x9f2zTJPEnln1tCXK
udp/HDXVbWsyuCrG4u7yRfzEQIT1Z0S1evYHHVPQl7AmVugmvavmzXNJjToGFrMd+LYDThFlPyK6
TCJs4QBYzCiJrvoxMscvOBK+j+HT/3RvMimOm+2IZxQoV4wDxCjHwDNWwQLRw/bua+/bQJ7RSFWd
9MqwRQD3ja0NX0HcU6xqYAjT//p2xm3hQyHGlAsz+LWonzqq5Edldi1ZInKdwEFNoVWjkQUGuGwt
wkKIYrgP/JSPmnfm10n7P6sE1Cg2phxKVmEtzZaZ3swDIf0FrcG/xDQJUvKcMv6UfmYeF+yPOAZA
H+QQWESSahlHkh/rMZmJmG1dtPqiJOxP6RJViMOtiUl6Buh34Jbp5snFe08yAxu2Hr8rjC5DU97r
eANxGhNiBTRzp0kS2uZTu62XApO9iXYJBVMzDo95jvkzTT8TlF+glJp6okCTVFOwMQz+799PHQW+
RyzPIBM0ZZVBT0Xz0qOKuw9srX38zGuHsc+ezZVHy107qr12agac0Ia+npyD+HcutJinuCBmm2G+
YkBQ0U+/HnqFefmQ21uuopNndl1s9+cv5oly932fbSBfoGJ/5D/r0yorws88GT4wF9s+J0vuQB8t
BcqrDqvY+gFMUIAgdL+YBVyyZ3lna+LgDZs+ZVNOj99npadpm1TQ4Jw3q9T/M9QdZ2Mf5jUcBPhk
GArGNnW5N1XvCWz71RXlnJMvOGLJBqQ8Z5FxP02Nbn97YmutTa1A3sJQJW/F/QgKnsiSQmS/2IQU
cZoLYozFnf4Nr0ChWeXAZDLtAakibOvlgq1dV/HQpeTuVNS2WZZyNCLkSjiMYRCrfZ+h1uZbDlpl
zmI5Ew1hrkLvXxC9r9OusAD6QLXCAEoXi+AZlybkmTil1/9oFaNPAjbSPbZoSNTUIh1WFJ2QWk3/
zqnOu/td4hy6bsq4j1vTzL4Or3EBDzIgGgBe0X/DcZpvp7HdsLZ+7/zIKZikLXnRMUKGnOQxb/0N
ws+VZUSsebpXJqVbKWe3wj87vfJ3nn6MAxbySWnHqo03E2ikdocdrIX1OeZxdbaE4ZRTEJdCPdyB
fMDVx3/r/DGY7tiqRpo3VnoWTc1apKEwXJYz78Ql5cDDBALUJQpJk8uFu3pNvFuIA0xjnNNpcJ9J
4RKIswweX5/rMzzy7HUyJocjgNsh4e3ZX0qvG4aE1oTEr4YuYxH+v0qNMdotSztOjdyhFAa8gLtW
H/yirOZU5BvcYjLUJOtQUxJbbZcLY1wDMTMGMpoo6Fv35DGkSpZQYpoSoT+9cxcph7/R/H3Xr2xE
oX8hzgAtzYAXSOWY4XZKgrhcwwu82KM9ZdvVPNh6kR6VzuqV1gzkdQAQs31hXagO7PIktaBLUM2c
VCuOs9ctBxYNWlZsZQYUbFUxZVQi2zhZATc+krR4YLh/MnbgqWKL60o3yEc7DoGOZbodOlZvAeS5
l4XQ8dzQGZb6KDmJqH0wGeH1Vw3K54ZuC8fQrZq52zPQA34lFcxqbZ3hqquqPbfEKXjzCAryUN36
I/2LyEiDgOTquQFc7gpTK8wTEwF6NWuyTPtbkDLYqhYzvgtCsWMamdNGdky2bsaHg64T02Wm0cIC
C0R0/Dh9ZivjK4RDKiFNdkAhhj7V9rjjOhb81D7/84FkNMrFfhcX1n0BlRBJB5sBfHQnu5G4VVod
4MsfBPPvEAzE7Wy+wZZocAtkl0/P99ZjDLNT7l3Bj71ulUbPyFQlzdoRy8WiyKWTytM03Na8c5lQ
553/ExWt+PCdNGu3q3NvmIL6qlDZs0l1DPZ2bkUOrLd8z2ciUbOfHf+sWrtDs+GoDT0bbdzdy4ny
Eks8zvxL4p6WcWHDz1mnaEiF6qM6c5cO0zJNm93MQfEbSMYmJPVdtHwnrR6H0ihf2akkKqMLIf7d
1FMgqSE0DPGj9D8iuBOjEmXgpSvMqIUvybGXJBDTzg4n7EzBBWdo9VMj0IU9SEy0nlOeLDSyLE3N
iFh+UYUj9PMc8x4KiVL6W3x4X5QMapwtCWwgKH3zzh46w7W27juyPowCeyyFUtHK8mz61AYxsbjd
rRoAfQ9FUUOhxQbyskm8FwPz5r9JS8FicRN8mPg98a9kj+LPMFtvUxLzc/F5q3GZ8N9LABUuct46
thLuribC5mJdcspSe5BnuhBlxY/PMFxFTrtZA3YKWuDXN956NxjebTL7xaMA0Zer7cwTUwBLqtEn
94WjRqbtcMrNFLKvEgI2zEvCYoYVXSVJUCscYZQWqFontGX3CZ/FydP7ZR/a7AwV+iVxNHWaFlas
/dpEioz+/ndFUAUKYKsMt0yJbTqmfZBXDWXcWhvpDAkKFUgQdWEzf9Y2ikilTAEDi6o6dh820b3T
tCKQ6MKo158Yh982ROozCreNqXQPorKPVSBGbFLw8bwWhhxWMZLYZLFTREwteKU4aT4kp/SPOU+F
KZFY6Bx5AdTzyvzYh407kM6N/6noomFNSu2uw5gGXFOWh05DG7pLqQU6sUk5poZZjfyO2xGpVpmB
HSdmGjMJkI6iZEWRvAE1/hLPqJkW9i/n4Y3ZcLGff+UwEPJ4Bxz0l2g2sLoDx+f/0nAoadmdX+4j
uyLKhcAqo71gViVnII+CaOgUSh3jpqsg36CIryTjqzMNsWKB+W4uj4ilGATd9+Wj1wQXamotb82b
/U1SrEnrZzRvaILNs46Kvql7H/n6BmV2ATQhPy2kGAQL57ECT8QjosgQYZOkCtxUPTd9gipIYa6C
QIyNC39xVcN3SKaysl64j2Tw8hu9j/HZG95mrc/TDRyaF5WCerTcv8Mc+z9CaYkeMitJ3hiHZ9id
EM1OrZG31YdECljl2+u2h0TKzxhRNUGimGsj66V+2X9pDfCpg0Tzfx1u0+xZlwcCsHFsv4V9mnf6
yh5bD1w0nkX+4uec0SEZ5cQ2GnP0cYpT5Fc90UgpGo92ajgkbMec/5ltb0ZJZmFXONnm4VBYsu9M
Z4FhVP1fzd2bZ+ypGAnOey6H/X2oyFZFmshnGhSSpRb5r9LY+dC6H9bFBFf9Xnpaa1zSM3KBZduj
In/QJZ1uOF+F0fsBm7A0WjCCsDY44y8fU7PcjdTbc3BoVwWKHcIESe4Xpz8qcDmVYTtFk1HEnpeL
+F66o2LCriQpcBvWGLuaKdu3sLToqMfAQ2yO4n3Z5QkuOC4CdrjnSX8BPirA5bx6mN/Q3abIQQ+K
BsVHSGXb3Z4Nik9pd7+Z4jo8yX+VbZCAKp6mgKOzaKbT/tWvL3rz/BwW32wqVK2dMaY51XVQe16X
3TsrmXabszC4BG2e2G5AUJCJncfEbsEXKuIySDEDWnqU//mt/73TqoefaOnzpUouo8b+0w921KYe
hYcUrBwKN9k1O4K9WcjXlKUg8pnFcPlb/2mbp2oHpO+zFZ0CQ5yBA5WgYbD75dgPpEtjGRFT5+kA
vADDa0ib2DO23AMItR/OiEidJLuZqfaaHwBb7G2/EHonE8r41Z+3O9acjx5jDdcTQwgztcWyZzdl
eXYQLsSMSvO1E0BvYw2BeWzh+jiIeYyrGy8yAXGiDZpfSBWIsSU7Gb4BaknNFkraE/4Rz9rSocsy
AMyPyPZtJ4EmuoFqoy0VwrVeujVASzKkHS6yGqGN0dgTDozvvNlvaiX51OUrNQjRaaFK+gsLwPTG
REyN+UFr8rB7UN7FQh6LFxjZkZVfTLktr6sk5GekNkMu82p1bj00wwv0NwIWyrwnO8ndEzOrkGUg
QNfZK+P1jwun4EZWRCXiABsTWSfKPEJLTijIs9pqF08XFjeMUo9Vzj/s85VgHbGPTURmNauWvyH5
9uFXCjgsaetPDCRzIR+aYjJP9FBxMldIUE3fdUNRJCQli8Q6CK7UlG94h6lZGD57EefJuNIbYxlY
cRq0e254BTcUgBaODjdW+dheI8Q61DZksd8nLI8e/x1XsiCDFgtNZCvNVOSDmIkloxEbc9eszl7G
m+Jck9xpJ00AOCFGFbsBrH3iQeZGYYrFpDkZHuGwTqV29iXXrcABaiGDe/EyheTajDK8vzdfqiae
82MElBTpxf0C1wZ8s8rozDsAFdHzaY/0mDEtpxkeGnJhBK1/kt0xrkDrNK2/B6qSTlB/CdUfsO9G
El1UzU9MxOwlNx8LxSTa3WdyMZK2Y2dmR4xkaM5ClDWQp2bQGdw+nPp/x7XX4LVEyg158nC1ey7r
ZyGyo+Oo7Iu/99cqR0POQ/1v28iOlX5ZkTJ7iWp3Bz/LVBcEthq7U5opoSTqt5uiIeoPuwfTy9o4
rTE48Pmbij1hO9nm+eNxY5Oa9d7DBjC+SYVYwbMIouKBlxSX8Fz7QpJmjRRisauiIKEXmLTn2bxr
GjiL6BvfpEorfFCcYQb9hNwXQBoVGTJ1eHCQvGYoTYbqlJk+zMAsPZm6kqdqgbIKKLARe9Lg3emK
AFRK/Fdky4YSwo3cmvmNhfDAf5kKLyxUCGkfmgxfOukIqqkvcqQToo14ETScfXfN0r7v5cNeLsn7
Uo+i0z7AT0dC7csEcMSlfs/BoU4iqLT6+Qczgf3Z4Tmw65I4oqKS/iB1saCRCl0oM6rJHKRVEJt0
IHpTjHd9YmWZgJU25RQipmYVuXIUgmV5bGZKegLJVlOXDOmmeUwWwINhB/vop0NQha9FzZ8mq+eO
ve/n6jKd8EZ8KWveLkmZBEtH7uaAXfEQCn9JGBTXpIijwq7OyVmDypYEKjMtBRSl9W8fh43FZJhc
3kz3i+gCL4ln3rmgJH5VdlFTz5JQpa/eU9SzYLBRj49Bq2QaoC66FjgReTe4Paz9QCUbnmlZk9Ur
W+gF1TNo4gnzW2gZIPNVmTOoYGrEuyi9YMeFo6qCFzL49xK2fb34vChT9xopeKJfLrnL31y5gH/E
gdZnJFhQxoO9TUzSdkeLZos5KOdS5Xbf/Zr93IRDVIM4m+bTIi6wPytmoFVvGdM/XMF4MPsCx6sg
c7vJD7uZ1eZNfan00hlSUR0B8LJ7CaBTNRuL0mEZukiB5+npP+OxE7FoJDmRwmJ/1E1o+vtKdgBg
toIoqjrEHbx/AEgqHmPAUkZcVBeB5nDw/7QcoHwyB/mTKQSZw4rf6e+LakIXhBOT4k1QwE6gYUNF
b7qr7ohDqGbwmceUlrXGE2rBo6MSw1EI2xQTNGWoZNz+c5QWp6QGsO0AOjxVKwc5tcUJ733BHyX9
ovPNAWzorJiRD4lAS6orDtQscGt9HYssD2QRWHRtatAAvNnxQrb6qn7KcHcNdvl9jrF/l3o3hp/V
dM4bs+IYeJNQ91Ja5hOOcuiZ2MMrp8lapxlKtNMlzxashGMsekUJIpN+PzgHy1LhMrPAzBPjWGki
SpalW22hqt6NtVHtapsSUaur7VUHbSPZl7fbUG//7RgL1PsJdpROKnptZ8x48qn7AXJlEgh6ONng
HMsrSAQd7FXhyXGpvRErwTwGjJ0Auj6MrG0tAAMn/g203OjrwzWHLGfWIU19ygGawPJqCU3fLE5C
+Gd9rQB2fqcM39NXOACrP1kLY5MhxbgwSC0ck7ML41hdmSNtoq865vkwStneqvbDTvlqjbVB1BaM
PLi0V6KHQ2Zao5y/0q1HvqnMXf4n2860KK4qUmxHgdbknyWfi3QpYjYTGuxl60rU1B6GjCIrRaaS
jpmM1qWrcOKvhBi7vSim1tYFvTHHETCcyTSSGgYJ8gVoga8jhOqcFUi3IxqCBRHK9Juo5ZLhBmVb
tsbhNv2worcfk3EFBtthSkBXqXpMLTlwcaZInLIMXC/nX6MGx0q2ZhEfYlzhot00qtvRUUPd2ng7
+qT6SXho/ntZUCtS87mIGHhtEZ4sEqMJRth3i73CSrtCwjIP3Pe9Gn+HdjqlPojeHNOmDb9NSccu
i85btxaWR9Vjz0jl8XGW1iT5jOhChdB2uBqaUQRape1d+BxO985UJ51gFBlLR3FFX0EmGKPW4sI7
pNREL4f7K6Jy/wq20Eu3/G2zzLsckkFstytfDMx6ArA+AVxFGRQACM9iPK6iKJBgSqqy/6RQcVod
N/6NkKFq/iHDLydT3lSyR2qSy/jgM896KlcysQO2aIPgz7V1TcabDf92Y4d5xc9vfrgDh4iTwoXL
YSG7ckp9fm0yG4V9//Cgp5t6ZQY1TXkvSR05e+gVaKIa+r2P7yrjiRfMR54fAgymLc13QwTlYhGk
NoO2nqDJ/AXAxjPUeLBhJL6Q9GbNuxqAY+vI7OJSSFgK8MHDvnFBhMLQ6GF07ilnPEDpAVp5UqXu
ESP3ntRXW2JntKS50Q9GLb9Q49kr1D6QDn7eXB7MLRikMXdXnI9gie4nPd+6abyVZ5VCjXvCfnLW
rCu6InJsfIsxP3jlnc8KHgHZEEajw7ETvwfi+6mDMIwB88JyrvIyEQk2dVy3rKlnuGNraTSqQ057
CpZUr8FqZri1aGPoebezc2mufpomEObI4cfe/oD/zlbVTm2JUxQPFr9I3/xz3i56AoUgKNH9+bla
6Bb3lYrcFyyj0hAX30i/mSALrlGjEIKgqBB599QmosvCPF95SIxRh6G8gHo9Y+XbPvzWKw5ZAsR4
mjrN98ranLCYIv/xWob2If4CUZq300buwPdr7h3Y3J6mThLWZwiuj5+0Hr4ZvKLzg8n9c9c+eh25
j37f0+a8qDjkJKDwcVpJkQd0BQSaZRE/W+jYnhvjPHo0EHgq8LZB+wDjtWgoAEGttip/wBw66Oh7
3n6ePC+KXeRPWYctcJrhCA4ijWKZ0dF9k00hjQw715D4StPBn3BNjF5Qi1sL51X/YLzVN3nKkXyS
zlhTP4OVcCnn8+p2b8tXBzXi8rA+j9Od/pJSJFVnw0VGxuuQhLuX4ZRs4TadFjvrisrO/gTTBUPn
LqTzoKdW/zAO3BiEaX+EGHacDN27kUncYOLDvcKe/tHgyJFERnjUEpZ8i+ym4q7k4PlECA+Kyz7i
Qvyc0ZialNMP+70aGA8+aEpY34z8tggf2cff37rDd0HmZbVAIAhHMg7U5X0g6l/eUrCgOCKx8/1+
DIeMYqVGbIgaZTrZ/yvho5EgL+6xSoqQI2R2LTlHO0LaHfdSK9jofzGs6Cg2ioX1T5UZcO+JZkuA
PJJJhZmMDP94teL7YAnd29EnFi9SJpi6q8QR1OvZkmiIFc/HAfBP12ZejX5WdIYzw0nNqU7y0fbw
vsTfE04qbjO7Smp0DBeRw01J865SqoYZSS/6xzaR8IW9je5EroeueGvDbQAY2UUztvNPYkkch3S5
3dEJMGCKYG0dAWFVrlMFYKDPc7vynIDcS8PdUeD0Jn6A9ByY3rQPgTr6S2M0lKiC8NwuyGFfwM+E
MI1NF7InMqsFUIdsgy1fLY70Dg/aFv7tswIUCBWk8+NKjAUgrylV9qn8G74UnWq0yX8rrakyahsG
6vdUDSLnm4+Aodyp7panwtGitgaaHjx7moIf2tcIo+zsLYoRJ6NnOxRN7Jrn3p3wThWio3tLXgjm
m0PMtFOTlyQ8VOvDtoDA6f5NKFXRoE6lLFdXyk0V8Y4lauwxtgzBGTKLPfU5pjGBAoRinkcAOBa9
p6B6Hg6cVpqa7dVPQq59FIgE6ZKtEz4GC/JaxWjCZ1uLa2X8GCM/jCv4mH/Dlenls3ephUmCmLmz
xI0hAXthUUQYpUggVtvTx4Fx3zqRzossECEuakJxQTIyBuCN7rGl2Sn9iKXXCDrL57GpHNoQ5MXn
f+QHdVLsKnIR49NGeI6DhcSvrP1DRWgcxNH8krmo8hHrXv6N6jRY0808FQiW7AK1OX2tg4ZEWEeA
Nzk+P5m3eZnPKg6ssaltSMOqGnGv/4p813tP2nYaKuECGsLw0cGl1L6Y/bpT/Rco590veJfoxczz
9yBUINa+R4/enDLsIfaZWMOeLYJB0Bht4rolROwB4L9Yt4fyPVhOONr1fj1TnMpcIHa4Aym6czhN
Pw2WfJ4HHp1b97qVqHFTYxUu1GluR6vGgUdoUBVaa39nOmZ+MCLUEAxSNS5yNZSuhD0mrtA+IaQe
LiX4aApbkgjZEqebsjvhtQs5SpcIrunzxzkNlvziSpnDY0H3hxgjhfRNsjt7jirDIZSQ2ui8rvBe
Yj+wKX5VKI9BarTYY0XWY+ck00odMR+U30etTckiwCLzpfIsWQAFx1rM3fVPPtKPWYaHmHXAD2oF
65/RzfHVigIoZMXTEUstJzQcL9iwV1ZRKB7zkDCxYfyfr3jz/nKbP91h3EEBcnUw1zNHzFHoheDk
9iPDCtSvoZ+BC2Qatp6k6OPv3TLDXjPO/f52wtrBbyv207aiw3FVcezja/S3J6xhPogF0cjFz2XH
zlnLnWVLsmVvQiBlSNOM5nsKvpyFPfW+zP0lSHXTZGUzdjV+7/CAWKCQQweUHVjMZfNpzprKx6/m
I4FDC97InW6aTgWekZFpHXGDj5UGhcQKmfPDA3Re78eF8AwuSnDvxKzB/D8vbOr1R2zJUkijY7Dd
Q7V4Zt4GFlXUx6SdcoZ4fMQaiFBdFT4uj7pjUncLTKhSRv65byl7WDw/klNCbR4nmIp3HriiiYtF
Ee/OHzlowRyOLjMHYnXGp4FfDLscWV3WRiB4p7iX7t3401dejj8KlqAuRBn3UJm8X90EsmK02d5E
2ek3dfAWKgT2Z0KUZpV3TqqNs6Nf3SsrULO12Dath/To9WZIX3TpxlliqGRHuMJgsABHTMi1UBTE
l/GxiefErGIjY3BeVpTVi6FHaJ0cF4g0OtOnBV5P2UeK+lYvoal8yOfj3CTFhmLssGsVLpWGNJmj
JH7BX9xbvQtAQSe+9cMfVDOzasyv7bJ/FOEMGFjFzEtnj+zUH3Uqh7xy+M6be6eAQucmmefQZa9v
QHLDy9RwO01WbtRAr9j/kOiA9gVDuJfFGc/h8uJvf8ZFoJmT67tSOX6dROxxYUtBXfMHkWIhapB8
w+UOOydknkCYI7oSv6LSJ6GlbldVUXUdv1gdQn3TRb+V8IiztfFFGEpLoL3P8BXjOi/PYp8QW1d8
DgJlItzt893BGo7Z9DFSlEFDxm9twhRJA78haGPrk3+L5+Ao2bZxoWeinRAkYmnpuHb4hr9jtGWv
WRmAKEMHpV6NHr+U+fMJlCqyprEn+qceY2qjs96i3/QMnpvOqOXPacwIHtOusNssfNbBPiiik8Fp
X6qMMK5XUmVmLvX68RVEuO/ql0A8xdVh/5S3/dkhW03D2lUZZV+gnoU9m2gOD+eJ2IszmUD4nkSW
wSd0tPYxDjlytfSBcLeJjB0/SkR1539f5BolcpMWfxTI+s1wXqfavlKxaEug73rynDq+pYxZgGS3
XSGcEJgi5zuYfGHxVo+7MqSNSAl9s7tmcuIoqfrx199eLRApBx//C7bVmpoi0hzAg4v/sU+Ndt0F
pazTNxx6iKpYThkVY2nnsCQYkSDgSRUiOEvU9PWObmGgk6QgDQQylWVQ/D6lZKcuXvYyo8oloCK1
8a4CItWjJ/RANCc/8Y7Meoa43kadwO+oa6S9Fa+hCdlpP5KjyORBC+gXs3crYPX/lmHn+0gOfk9W
yPyDBT6Ft+4zcyrKSB1iqA40ksfWNUYChmMkQ2ZuQ4CLETDHOdKrJgSmZJr1lQ3Ob4DRVyMgkqQC
HdGpyuAWwWBlAu3c20xYsYN3eL3F33vvUCnyL1wE7nDjzijp+qFvBT6hveIYlFb6/kPBqjqvMrCx
kFjky2TlzJ0mZ096Mwn2M2n0kKa2J5C+H7xpjKqGx/cN2FiiiPWaMcjpWD4bqDrezAUIokkc03+b
B/puJ+EjkPG2hvU0RDgYFKXjQKgZYJkpfixsagmRMrizbWI347S3wWeh04AgCICTWf1o7XJ49FMm
brLluwHxeaD9KtJOvxsBmhCS1ohDBgxezn1dBJ2Q0lVHC9fJdiSRF+GAxxHoF1gOKwa0TGuLuFXf
2sZ1GbmCvxtolHct8iScpqKsWtqCiPwDsfN8T8zyLnukgvgCYYvdEER1PzbEkprAsrX5veJU61oR
mb1evLwbcru3tCWH1bT8YJLgk5CK+HfxlLWNf44sBqdbaHTx0yhPHtDzVxjteaU+ev4MUYfB1MLS
8+NH26thsL00UtHDqgdkVpQMCuOQqz27lzWS5DAhuyIX6dmQzVlp3qXTOMYqcpZetNQeUOUu7U3X
m161GaA50UDJhb9UmV1twEzJMEpy2lEfsJ29o0AN6bDVqDHcEBgBb8Q3aLdhnQ7sGcDb9PyRWCD/
G7HcfpNtIBdac6q5l37a4CZdyrfHWzU4GmitX3lKH+N3zaS0NlFSPVOOyB5j6y3reYyvuBsx3TX4
Jdwozq1pAZNOcrk2XZRAN/RUhc5WcGyxWLTqv2xWoXqQxpRvdiJFaWUWSMxLSesXHjbpdbJesn7i
VFwQoUlaeQO1X/yQXYdOtx1468se7arj25EcOaB1v6RAikRqSJ7HRzby89Gx8nXGrXuFGhvMzoUq
QHk3ZWBoWxwR75i7p36tDzUgG3/Viwp9VqnswIYqynSOsBq7ToV9tz1hTe4LWFTeiQJ1agbKSCuI
NonmaaSH8xWcGxMz9oixOR31Clu50D3rllPkhNfSoWlznIhU7y66bvnuQROe9QQQ7SbIWqa4U5qP
jgoOBVg3vsWKmR4McKNiYqiwh4zI4iCayJBR7OozAo50jqnAK4agO4eXZJwnr17oG0T9YDSpcCmx
35XXF1k81kE+nEVb8PWvK3Lv+X9hGGeDNzdzjoRqj6f1chL2tgnDnSgpeZyK9ucyea6JVyph+iSZ
PyBNYHHoTiWoEE5wGOi5vuUWhMb1BcZ9WIowZuR3zxvvZy1lrX5jsqY98eouYbpl33bmMFvEL//0
ZyRrM3JILpRtKg4+OP9xBhqJYK7ox6v4NZTkijaa2hMP6bcbtjygkUuGxtWr745j9iw1eAihxhQy
A94hFsZs8nmnWaxPKHpoZ1fkP+OcB0jIvqC+nT7F+EfpCoh/8oZ5XMpZ/zWJyLipGlT7bSQxDN6G
7W83hTLvAroRXmDxDOZXLaW45vXfnTln34Pm3bVUxa9R6SKBTldJXSiQM0Tj+pm+ksPRn3rsE6GW
Ir95V+O4H7V4245x2dNR/kggDPAdtt+z648plqnaSvGYVAKOXfTQTu9hkQ24li6Xoh3TPmDelIcp
XEreA+tvjGBgxkS4XQ6OD5PKRMZObFH2E5rMsebO6Ay1HtkNKIGMvMp4ioQniBVyU+XtrHkdByUB
T7S6p67u3Ty/PfI2p8zn1gTLp4WXcipodOWyhSdueJ3EFWEoczKsuiZj4u5DcrJJTHP5SpqvLAca
tUKZeqEA882x+pESKLY/wacIWTenCk30rSTkv4bKEV21pcWcBHQzItQV+yRQjfZrOOuwWmht7mmc
yOQBfAd9pLJWJ/Nao9qrtIyKdTxCS1iAqY3OVwf6GInKMx6L6KI0gV8hCGsFxuvwZ3W2rNKKYZ2U
/oZhgNWdxNGE/jyEpImt4N0VpRdALrfrpPsD5yycWE32ExwwjqzPHSgJinCJG86y93TNu71bNJwW
jeZxIp8H18WzGpzpqLynwCinxd9PPYkOyRQIHrFXiZqZG06kJo6LcpAVxyPqajbJ44iboWC6hoAB
/0D9BjpAlYW8kIW6ISlX4k9o2RNnO3rKMSnlUxlrjYSjXRC/xGg1L7RCOzhbkb45SbgC8+SCX2p7
WvCVMik9P5XH8frvx2v8U2pFfmQ2TXxJCpgDg+6UAq55R2fsdrfLjWrz9NyR2wOy6azR3qect3ce
VF3ME52KzgKiTZJhP9/Tuiq7r2dR1wm2JAL29Z382nzXAwo77xE3A8QGb014Paob7mXi2STDa+To
Oa/6lYnefrtk5b+4aWCz59kAlWtWxwgSJnDmHZw1imTXrxuLibmJym7ZYjCXnbNIzkbz/cMrOxtT
/JU05rAHxdyVZrFadVKWOR+ruCXmmHGOdwgKqApqzQLFS3P1vFRk4D4/XWx8tn6Oedww96eF+ULX
0ZqXSYW7AwvhNK0EQ8RxpsllVXA1uwLEjVxUKcWlRFDCuKbu56PC0ScZe52KKN27vh4DNAeNYrjC
mTZEbwGatPJmPr2Nfl20pU/N3dFveA4MNSwjZeRSObUH1JbcJAia1Efk0dpqxwWLr6wTnoqt6F30
kKtwpxHQ1TPOv7/oB1dFxeKyOY1kjlGx1vNRoznSgMYGJ2SdxsQ1czQCe5FrtJdSNcRBooyNqADJ
eOtTcCYyVaqH1nW40hnIvXWw8wRTQihrMGst9sp1V3weKR9UtnSprlVeKQqGK7AP3FBPVRpNEmUT
cyhjxyWRXnH9C2A0HeihA4IIz7Ze+cHnSOO6zUtuOwtBWvzCTVzW9GwqOmnKtPsBFy2s5fGlolPx
8z8Sr3G81uFZVFoatObYWF4b1j3eBnK9zWm6eA0iXrrAmNFR3oeUFl7ZfQyDJ+W03O7XnzJrbPD3
1/GOAsT1R1rntFI+7w9Fs8yMTLWsvl/bWqPQlLiTy/jmsz3Lzk/5VG51N3cssOn/CHenkr+5IAJk
aatZerfhYkKzZwtECSkkn6CHZGK8FeB6A/xWeBQ1OPXeRHskmQLI5hr1AFdFjp+MTorj+ThAg5PN
yZjMqS6dVZF950inY1xIrY0UPnZ/nWnrzAdg+P8BgNBjrky4vkfoZragpB0whinVTWCvxlGGK553
c2z8aDqStnGhA+rEPor6C3bHHSnvCStCOtzFJIsXkdcx5MYe7V6/NQLBiUnknUbJ85GjZqtQakAM
l3Gb3dpmk9SHFHq1xht9EfG1BfFbEwCF+byWuSsNXj6+xo7JPWXo43gQG/5V9/bViGui/ZFG7az+
Kl/w89OlCnVaoS2yTzcorrf9CZRu9gNzi4sQBzH1skyim4edDE6HdlYns8mNzBRiZco9z1g1zSo+
vjTz4K1oXLq6VFu3ZsFATYMZqt+I4W5N4aED3fA0Qr8IwlBA1547lfk+asZMgWknEmllTAWSrO05
vYGvjzxtI0w0b78flHg94SLnbJjgLGZe02Po27KMttotQjZbP7nCmM0ID7A34avzRJCfSPd0kMsD
HiiH9YqkoxRubAvc7Iorb/icZey+qeTkuJ2yIOlmOIkjSZympcfxIfKFAQLuaN25NVdkDnn53Fcd
wPp/0bZRSxWafFtnJl5wvHlnNbkmHr3SpRaV2Ptwql2qXzD6U06xdW7I7KlarHUL53vIhoweKPjA
QOToTCP0JUASmX4ttCyfQzmjnEWqgqdZhywTfMQWoFQ+adSeycErji8BwBWJzgAzCfsrPNMKq3Eo
oo7bqeEzSQPzbCrae3tQVCdlId0EI17fiG6HHXYZ9+2Iwd9TNszUv7dMLe2n+tJ309r/u1wcxwGX
6S6EvKCbW+cqRc3StQaR1gC+0H9yicLbDxmYrvf6hLJLxubuvhMejY5+4yQ+UhK4WvZ/kwNjSBAM
lxkIHbkw3EJ4x/FZGwAmg/J3J0mjmOLGXVkLku7jYrQGyxIaI3YOeoaGwlqFdbpZAsgdbuLygFci
7dxzrHFl5003+3zMMESGBz5cU55h569uproemHdCyxRmwsRJoQ8qptosspoe7p2wDmEvLT0Fd4Gk
Xfb/gU8/BTnWmlFTsy1/6dckWSB7O3+/t8UZcMEqKF5JJxO/eQJtafQgluDEc/7gEPHkaFHTjy35
NVOmXkg87p0ND8QOEH2HQwUO1Syd3VSeynNjgSC102fhHnkk66VD44xSz2PvwQRFyOJ8ScldjRwY
Zo3f40YXYDZOmd85IvMeo5CB5cTD3cIrpZ0zEDRhyvpaBSn6IouqYYDWZGNNQnEhaFFn5o+icfcu
zj6r/bMFieIOWy5n2pIKIbB+6HRDS1WwasgK4RANFVYaZqWWnoOGP69+9MO43K2QiE6QzNPg9Cf1
SHEeMT8uul/mefEN4Fadmdmu6F3MzEDLB8y6Roarzr7l+NdNarcwXqx1/cjUIVLI2NymMiXYdp0Z
Btd0lgan3pC1hkdwOi5Np6aDkH1J/gFSnl896bNZaHqvXPgSzMAV0IpTftaWLa040+tY2368uJyW
7rBUabkJ/KOA1wnx+hX14+13YBM/NDZzADW9yWCqBXjV6ojjZ1f+RYQd4dbl4AtNizGMeJkU85gd
zXwoWL8gOV4+wyXSrEjoZnstxHYPzvIN1AEnFu7NX/sC0TW+TepMk69EINLcsZsG8urOLHxoaAt9
1CumyrwWGY6oqBTKx1/juwYaTrJXfEk2i2gge4SueAD8OoqbotG5hKbZ+BYjfHryrYYDoId2hBAR
yWsT28tkZSYs0UIqBhI3U8xfHktipfRl5oWCReFQWqnUiGS29vfdOYsBc4dUoyoFEKA95F0JqgMm
/ryYqoBQsAM7VIXh49z2OdwfZweIGISd69pe4poEcp+YevZsTQSWH33lCbMikKm2WMKFf3C9cOvd
lIUgZlgMgjN7ni+uPeN7y+XxBURNbIMrScFZTD83QZbtn5FKOOyQW/NygTVJnHF6DZL9QfaT9kD8
ue9S2bD9CZAnOrcD2w4FKeSuI54LrA0ZyssjVkzk37jg9EP7tEfGvUSBilD4MiW4DPdhEXU5u70h
4uNOJvyjfJE1UWB1L6y63KcA+jCKlz1SnKiW2BeCKdS7aFYhu7y/Vp/NGuRM0/NLt3QZFz2sMuVH
MWL8wYxlSyRDWRWcl2t+Ajdnqw5Nt6m/Jw95oPgixssUKQqjfK6jtagRnqqIEJ8vaRUGWbRKgxxM
vpRfPHHBX/9n4O2vuFwPZB/3Z5C2xb2+c7KC5z8ep4FSkmBH+KD2niE40Y+ggrx5n/NX1acmTjFc
/3ALFqHwFxtBTLl/KbMgIN2MGg9f2KJo3mvHgSS6cBuvf4y9A7J8SZr4rOYea/8zgmo1zE1EWfJY
NZ/M6EJX+xuHcuQp7h+u2GmpazkuW5M5iFxYOX1f9qP7zy6D8QVcCsFu4XFJRL0hgWjpMFp3+pB2
TMVlQwFL8tMpsZ8I7tq1/Ac/fEYH8T15Ml7Zsz4pAy/dyQuH7uTYd2BzDrd0ztrmSvtUHAUyztFr
9wu5HavXgdJDx77ARrMcERmed+iOoMVyelWQ4CJ7RX5XA5vDmonF88S9Njm2yKrfgo6c3vuNJfkh
y9kz3agS9Pw912Z84hFy5ZVAL/MEVWcgEwsF09yGYDnAL3R7T0b+SV2fZnSbgHQbCHevKj1ZNIEZ
tG7snLmMz7V6ecEkHen9AeodNdReGwIxH/FMFHVLRSin3OhoPYmkyQbYkjAvH4yx5RXqRSD62hT7
nECQeH04C3cVnY6V1uRiSNJiIUaack7cZx1E/HWYGQmL55KwGKbKXugJ/cDvsqoV686BqttM9vXN
NfMVqAsUnryEHT0Qmp4hokEIwG+NlGfnEcf/SgbpuEX7SKOzJtLlx+sy6hJz73OGSv6oLyO2cb/B
KnjHSYDMKtUohBAEv6sx5c3T7NikWTXx/Yn1cG+wx7KM+Y7+T25oF4jaqfooccqt6hsQWrLk/pxb
kBsIu6HUXoj6sU1PTG/UFA87OthajeKlDk2vRf6/zqZNvkn/QWjjinLXQrLUXqWY9a+Rhq4c2m/M
TjwdrwU+cqQI9sIoAvijZ7wr4pf+LCxCdVBJFL81G4nsc+HOacAGurDj2QuKijQD1FLtVrh220m3
w2KY8DYFxu/sq55DbMW+4yelnnU/bUFjkoVNfCb7+uXbtYvsRf5+0WPnDeq+S5vXmwdSY31tCBJc
q7a4E7Wc/Wbj4VbToQW9WnlYmjz4b/1FzknU4e5GzxfsWQ4UH2brtx2YvEGv1IdmSgh1uK5c74sg
UKoQ3MXP4Jq+DUDDAKxydXb5EijxTTN7sibtLbTw4b599cbKJRRzmpHmZdT+4zxzgW69/oFWKp24
hjo6zMrL9tyOEwyP1qukKqkvk7JtGrMGrX2+fHd30f3MIXukvJoxiTyDuF3KJbMWs8dez2Du+zrS
56grR7pODH+qeZFmNW+S8ObLolz6fHyJu88j9WHVHFkMguGTuWKMXSkc6/v6TdmbUHbJDHLAzabZ
EUy0OxhWNKQyFsDlgBCVds4q7kKLZNBOWUl6f97qinPRqKM5XymQqax9JxEMP7LY+Q//qPsVPYcA
XyKh5hmjAfEoa1zufxsi5kTvB/2g8nkNeQKLdiFxc/zOSAd/XHON804R+JivfIAo+yfN1URU1AFU
UEdDMgwhHbh7gDMI4YFpri/+yyHnUZPQOXTMw6ldVcua1qrPmawrWZ3U7v9i6J2CPBN0uGpk9eEZ
M2HHVNmZnS5cT0Yrl+6SrF0C4E9/T5ucchxqX61L67l6WKPmVxWFGQ2GHC89wkraWPI+Fvg8rtdV
4RkAkahS4+bK1kedDwqGb85IiqctVKta6ojfvpcBT9N6q0fz3fj4NVTzCIPY/ERtkTuZT02Csvps
iERd3RkyHuxb+SOXgHqNO+ZtESuW497qSeKGSOO18tSIEXvdcU1YXs6EhbXse6aqyMyhdnIUc7LD
/jYFkEES1NISHbDJWlh5mVGzQZq+QJCVJ41mYqkrMoyueNZlT1mCZ2YZoVfzuNhtH1IynKE6mNAq
+Z6YwmwXt4x0DZDPbkLmGCXrR5IhmN4V2yPsMhQnvr+S2DlZpIbbkx3MllW/nuuNyXH5ZP1iP1LU
JnOh+sXYP3okTuohrvq6kJLwxsT+cuuXKrN78FNmnFcWsTfvovHHR6Pq+ZPLNQR8pqGlm4UEecZd
dsK1ueCCwN24FsuyDXKbV1yGta3Y7iSqR0Ih+Ay2XtZwO73v9OTNMIheD4a8hd9HdkdppNfBTbQx
kMN6GGZ3rQTJhbX9wy2Dy5JzWNk8RCzAzHNf5zaLHqMTkAyTubMSmINL5P04AVf131Mjt7AXB9Ia
qfnfwSZI7V7HxRmFQE8VKEEpct/DkUDca/2V/sscLiBejtYohDrjNAZ8Wnh/4v3CRKi4p4FgLP0/
FoLlZHL/aPIpONpDbVNdiM9GEMx8b4H2QNQ/Fa576i16Vr+DOw/4XdCQdV80jBcf5h8hSUWmR9W+
g0vkVr9ppBKEeOvIxmva2VHzMcLC7tWB9DVIyoZ+9/fqLr+tjjRW8c62HWl2wjbiMPzmhSe4/RO1
yWRIL018jH8kuH2IpMGJ0eh65EDDu/CyBZgRgsJEhQSDnh/gs/rIkTuUkVRxWR3NBQAXAiXLeEpA
mYg4sYip/7aOdPPS6YvFE48VwrEF6OAX7ZHeTFeMqJ3hJBLdFHet8EEK/PizmMoQLrRYStLw6KxC
xQCrDiOkg8HNd7c6mL9ef7GuElZJ2awQAqijMICXQczO09c6gY1SnfzXKZrBSadunIpo1Hcz5FrF
RldfUYiPjeNLaR5z8Ueu2p9N6CgnVD6WY54KsZxi7/WXEHczPpHV/RogjsYn2EsySK6W3Wb6myjS
n4Ixcbtdb4NQh1gJB737gnYHWtDBjPhxICsFnPpPRoUv06MkMaHjmWLuaeuxSN6QajD7GMHYpRqI
CpM0vbzmd69HEJ68g4abBNZVCHZxpqR5sSaSUTQwrZpo95tukBlPhPZpbDxBGec+ooXaRChDx6oF
YtWKLzUe16SBnX2tPV4DLTwPwhft++bumB94FZ8LlFiaNKSlf6ETOAvtfRoLNlEooVmWC0T/80v2
VZZVJQqvFgLilpW3TVX+u74U6ldemtoVhT63/3+n9VYHfJ29eoVRt2U3rT4/bZcz+IV+s/XDpMgd
Awp5WpOJTOy2EE4nsdHDlml/rHocENyLFlDJ1R7CM7njW1jkU2wUnv4o+tLhQDXvmLMNwAWkNLC5
4U2UCEvnB5yoYvHaFCz/V1Ro3YdRa7ULo9ti21bt+E1pvFTgQHQwxT5THPHcFtfixs05SojO+gSi
FBEnagRbyCWnHZdsDt2bieDSlJMMWAlu6QNpg+QF6JN+YPib1JIVCvyDrZiFR6iNtAt+8YpWGvNS
Pt8EaBXVsVPgKYDNO8BPGu4BPch0pFUfPkwbgZtDHoW8qfVHaGuUh9XbvglyqlOSxNLGfH0Gnd0A
YpBcD1+BCZq7LKQmKgi96qv58Jrilzfi8faHxbE5fTVO4dDfkvU5GqVE/RCXeyuJVkLoJd7gJVbu
gOPp3K0HCEOTjhLaaRN5P2k1Sr8SF1LJ4JKq4K3oOuC4jMGi389RySdxjvcXdnVOBgirCu8VNqu5
ppQM//8yXZ1UWU+9rrxwEh9v2PT14UYToOca5Ca/ebvcMhuGSiBkW+UMm5SA9uznzMoy0Ho69bc3
07j5eKHsCEKXSEyvFEaBsHZckW7XgVFcALPqGLi7s4w7N8qMCmMbL63IUTeo6cfRi/bnWJLKoqbK
s5Q82L/WVdksmJwl7zVnikIw2K0u8bEvApCguCiExR3pVpocbWBUGOciSlENjKrgWBjRFgGxYBuY
k5U6bFpSi5o+KtkbuZ3RaOjzqgOKlDBypqzRmLMhTza/Yr138NHi4bQ7aysfBrk15NYKGqlLH6g5
Ke4VlEB1CE+T3TJ84A/+2RMq5Eh3G4vpVQ+b9SRn4WsxtPjRZGCPfXccWgEEhqHxumv2pgpJhFFD
WIrXpALggYW0wTsEH0BCrB4kwN9ASuGOv4BsXZMml8QrN0XD1bdlKG5rATxz6jtVDxHycaAbwNHm
jJH27BmvrtnXYyS4Hn12nL0h43AuelWHJY1BSAvMt2WmMT5RrZqtn5wicK1DHozJWWDxaNtkxIJ6
wQo/JkDFEnu7kDdmqRI5Jk0CnNmToUUG/6qJTvEo6+a8Ybq2vZ3W4/YaRDIlyKg1j0SCK0I77BuN
2SzC3dJoW2quI6XbBQQZkHPFt5WO93csz2ayLXkeiK69FhujDcf6UbpAVnYWzsdEaNHP5EiGwAUF
FIHC46xCOrTM3SwTtjqnq+INeqUomrAbk1UKSeOXf0YgcUPKB2NM4+FaZxoj9ptJ69Etkxgfkmg4
/9hIcTEV8rrEHh+HYqIbEJ8N0YwSKdMujnrh5ENhvEerHhA+YWvDKoBfZH3/MeHUaByWch4pPsFa
MOxvW+4rp/qAvwKXQzPz/OVV2syeXjnscv4F4GXCPjQ2zRzrOe/xtSloJm+qi+PhQN3DCm/CRCgi
rwFrmuOkMqh3g0cYfEGQtHL3+qMQ1KOHHnahW+WbElOB8T/eJgnNncwuzb5o9zOd/LEY3Sbjh3Mz
nIzERlRvXVTXb4Cw/BnnKmIhJWPawzL74lSmQstieBfOAQ3645K/Iq4hIDO4xjNtalxrBjGtMuen
A+62n2RZsHA0YsTUVjhqIikaMdYOA4aSJ6GXcsKU8adyPjpECjVyQ5heJur/vg5QEMOusd5LzQK0
0Zyd7Hg/xFiTkN0BU/B1L9jDzsIFfHF9gWDlP4lxjp96yb3aetAu9ynewv5YM65pmpjw7AIrgAiS
oHzXAe5KJUDStkt3kDSY7SP0c1V5WrRxHasj5Y5XVdMBWtkmlaskD0tjRadPZePF57v6lWSJoykR
Cs/zGaegNcS8DsSkomjmzI+oazN+qSY1sBx7vXF+kaDwPZVQroSROvfXK5wKKItvOfbXS4KWtL7A
79J+OwIObxmCKFfSS0oAAcHay+w0XBhe8xkUtLFSeao+6dSYggKbXhAQUILPgMDB/I867Izte7rN
6652dfefiQooDgrOwMWmjPVCZnVKU4RdNSDzIPcrw7qsTAMBeaV/xrjrftbOl4WzTVMO/N05m6l4
c23EbY8yHcRCzBg1MCaMNrTWZASe8xM+8l4WGMZnniM8Cfw5n50CgH3YRbiahogc/wRGLvMKQuQI
QvRaXVlqzltNG1jviEswFbqJA8DXV39nQXcnkk+O32OP0zdGoO8Lr9w88iSoLSJcyHnum+P0Mbsk
oSbjy8bzMPcbshgYYFZ2+sPjCPJimJ6H56MCv+GYyhpaohb2IWJT0LuxqTFtJ7PwvTOTjjPxYhR/
XO+nx8DtFg5xJ212AJLiHnKqFFey3vABthJ2hDxmq5j668YJWPlKRIKdjKyHi4HFpZmAj/wk67aj
/eWsHyftztkOD3t2X30d7ZWCirfgBnQuVlwiCm3oLWLuNpBvgKINNeReLEB9p+CSX5A+PKG0N7hL
ODnMiUi+uaVM70U+b5m2PrKA4BqetjfZn05p+Z0aFD997g+h3/lTlbH+GWBctDx+q2aEpahhjnjH
G0fdXKJIuakXrqQHQh7j6t/lkmZAFVOG8dmzh08WORRH05mw5YL0UOqbkkL4fJNvpkSY/ag/3hfH
bQ7dfN/Sc4yMkaSx4uqO2ZiVvdp1JM23B/J/uq1fOnNxJ3L4GlAg6bxFQozxhYSWK0d36HYfITmG
hZpDnBWXdELwNZ7O+AM+wIJW+s3198P+XCQx77t1Q3nUIyP+NrvpMquted1xYzx7ix8Dif+FYOM4
Ued06OiqnN2bR1sA4E6Aou8IVdCuspn4n0LvtcuJHwakdWOMT/u7sFoNL/z80kSTfGi9yQXXQqot
3r315EPo4E4TznVCTw67dwEH1TDQKHIalYqO99aBuzcSU+cd2koazj40Di4NgfGRyuP8NJBZHAHG
aie6Kjle/NdNgUh1VgV7nLSD3lTkNPxKylz82HQA4KnFrX4gVipIM0BricnWlXoykt81zwSG9utS
bH5vUR+dURvLX70WDLJKuoxe+eIF/cD0xhinhI8L4JRZs2JfMRO/I4Ci/91j8g33ybJfQKIm8lG9
8pdf7SWrzDUrC0jvEh+66liJtr6yOV66OSLEx4EgHPRmouv9Tin7b4ZKGZRa/GyOotbg/UZeM85J
GBZSDDFa1ey4KUtFD8qWjSF8OqKcrKecLcRvFnXQ8LMNRsYp77wBnkU6BzV98pOPezPpBdOJh0/I
mgzJp1Ysj0qUAIXJPWg6ogtqCoz1N2EH+42nyep+dD+iwKWF0RxEznsZzE+8zHtDAmwvImvv2p+C
EvUGP+ZsqMtcX6/sqZsVJttXFWV4vni0/PTzZlorR95OX7oTaXO6xKGbpOeKbe1PTGeOsROlQAvV
ytnBcV3Melb0wmeRGBsUHxIl4e2IGuG1XkCKY74hv484JMEyOc+MGuNM93+H9F6ha4xZLR95+ote
fc08rNZlLBaoeo5eVRc4rfv+tIl8SUiW4UM6PgImua1F8XpYpOmLQ0W5yKWxr3lcYwUPNZzCsXqu
WU/nWOAmh89EGujiWtWbUfsxc1ezPzOXBZh7GWk7Q8EOQhZqo0+bT7oAyWMHbeiBuevlcZ/7LRQe
//AkqoawaBbbTM93jGkYddf6dpAIthKcYGtHdyoi8mJLJRTaT2zAU5ZZBxe3LiOWSXP76TWLuR46
3Y1nqiqiPBQrzafMaUsgFHqoNMyT1IZNN+OXal6GQQulULeDnYs6DXiL3EMT+Ik3Q0eUKgq+xdg7
jJyUAGn3kt6G7R4HRkY2GnBiJJnEq1L2wu+FoPMrSEemRKQuc/sBTk2xF8+n2FwBClc7IBJXtN2w
oz31lTBax517+2NbZli71CjSLbZOgiQFTjPF+6dJF5epBtjVn1T70O9lVesITjuu3MEWOZO32Ft0
r9b4fFmrNQ05GVMFvkPj95j72Zx+HgYm2mUkvFXeKEyR2LAPRHtZuU8RmPstmcddy9p++seCnHm+
Cqaa49orlTThgcNTH/Rw2V0CmdzheL06GT3JS1+d8X1ZsSoqB/CQxo5T1vf7qvwaikHXnxTqm8mJ
btiNOIUSRDnpsU5CeJIhRPnaDzw3fHQ7z4laFpGUlewWcFJ2y8JbdolRwZv+r8wkFJB7pIjEOkwD
mWvB1Cgyv/R8qb+gCHF1fDof19QdaYmlZJ06k9hil0QdXT9yCJZVFmhTF/jJ6MCF/8ca2Bkr4EtO
9Y6KsM6xBfaZdXU0aC3ZOY2IMRPnuuZGXEApwGEY34cuNbx8M3e3sDo39LJ4Ci/6Bqz5JrPp/MpQ
fqNjpv/k5u0swTRn3W/WIeqwZD5PtoRx8JAs7ZVCxQRnkWyVaIEUE0JHK0auK3da4GXqghTYqLQc
Z4jnhTQVzwrIFYO7vmZcOW3+iJRuLk34zgoMKYAiQ8tDY1AjnDHZ5FOLFSwV3CBQ8QUYMyrEy7ue
gm7ybmWKop5qGVH16KxjWF2YBKi4bQIs3viyLVf6wRhz1UCjAbrVcnycMLwn+aEHzvAKy1oNMOjZ
OCvn9waoQd9MzchLyoHCoB8dbm0km/e0RJSymSMeg+1Fiv5Q7bWRm/5ay0DzH+hf48BOd5y4Qy9C
24gqKO2msPREqPSONz4GSb6O01r8ek32uFzAvt26RRxgDI3EF010BgnO9GfEEMYhGUG5KVAzlQVp
/weSba8VRKoGm6z/fkFrd2VyR5/eYbSrg61jhRDMjidzP0a7qE9kin9MY0N9IsgAtFmW2vigH0f1
+Z/ZFC0MVA/XPi2XVnEjPtkN/HBaufmH3B3vFYhJpI7PYA7gwQqA/4kOB7oXRXVa7m80CeJQvsch
sYmxb04NPxljfGVjq8n/+WVQY8n/l7pBg+e4SpiT/GCbQF8gMAFiT9V2HSavrZq6Fx7CTY8Wikl9
LkRmGTgQAmxuEBaQ9x2FRazwEOWdTvSz8Ci8uAvKCRGKxu6xYiACwM7PvdMGoxMW/0r27S7ym36F
nm/cbY5U0lKzu5vDbw9/FDik2UCw2Varyv5jGFY1LSuNdJGcsE86u+65pmCr2bpyItKQpAKghwIP
7UM1474SanV2PxfTd9SksvkPJ6ZRog9gs6+z1OwGWr3GPmuHDHKKQo0gCYYGTXg7FBcAKCVylvDx
+q3JEHNb39QgXYWDN/4V60Y0MFiMQLSV5ojjM6MwxnMWPK34U4S3dE52RXti3sLLmYiMRc7dsd9l
VGiok210bofaJbJZQzcyjCMIMxYfaf/9PBx0os+Lw1VK9fiNTrmGTHzvksSCqbdsY7NLWzQoj6TJ
XgvtLALdSx8f/mpJEMKE8AbhrLElqVB62+YYIUq1dhIZ6f0RKvBJwCAvUc7/MDP2TAh+idL3WPmJ
VI/Wq5fEn1TeG5uOuc6R/7rn8ITduIjN4aKiMFkSuo0pfg8OmBpNWVf/0thf7DMsCht/hCGA1622
NDYwfvkuApYL454OxUjIYiW1z9IEAL/cK6iH/djVcQB1FumGdlzdoER5PQv8lZEafT+nj0B7ibZ9
HZbl+2napOuqWwBn+GKnF/EIOFl8nl880XGmbuK57VgfAcmO/WlWhfX+3KyNJ/TQ3Zk8zQQxNEXY
uVPz4F5tw77YFj56MnlMpkRDjuqpviUvXAytC5wfhkNsyBOpPpWAh91c0L/gk2dzLS1353As13Et
DwdgIB81eb6aOFqz7Ubus3+FGeDjmQRUBgcToNmCDA1iixxZH39KG58aubYQaGKuAIQcXMTfdue6
LQD6cPD3NXSuoNfdLx3ilr3ErByi7OHK78qSudki8FVGshyiAxfU4uy21rYkx2Dia7omKNLJOoTo
6Po5SusaZ68qxEXvXK7wGoVe1ajXMsvBTwazB4ef6pD5qPoPQ+XSIaUsK2cS5SJwvoMAXPcr8imT
6Im3QL+vNnkM+cwRvgjR+j9zw0CEf6PcF0e3mAJKdg3uqb59oQUt5roFIybWgNGkSi2Xh9gg0eqK
CX747j0qoCKzAgy9Ac7i7Op9h6wZdIL1xyTg1ZUw4Jo+iZ0cVfu5KkD7v8pylp5ie6ZG4b1AB5ev
tci2wZwYl8CP3E2USV9qnGzTy2XkPrq1voWT/npzM/WsNDu3nwhchPzyV5MCN5DrrN+ltdclHqcm
rBkyvCrXWHCD99asA4mqsOrWPaIx676BEfGKti1Dp/JW5oMRipKk+AQi9VbSIh7rpTC/4VNxtXTx
CukWs8idedY7Ly0CXp9pxjlrUJiWUARh34/hbZBdmPfzoDC1PVns6A8sjZ3OETiMb9nPHDl85Etc
rqFkwgBLUTEVdZRP5RwkAxc1kazh3osfS7JGT+bXEKQUwfxTEjroc8+XSYlN53/srPfLxaaoBeKB
nWrWe5aZlgzXYcFk8zm92MCO+A/rULTdTge4zRirWfBmXcRXkMEjsjxrcofV2ESe3QLkTraFsUEO
7XU5k8jEU2XJyR2UgukhX9jL4kUo3kEujfdyUPx6J/ZhP/gV9L3OjFJt8/9OLyIIzPa1ZNQsWFU6
RhMmhHGUeqTcagMTVAMkj92w1l3jfd+tYzdpt84aSCY8o+Yv0+rtG7bLS7EGijyvxl2vFLNQxsPU
Gr/rvUf3A41Km/EVMsRzMp5ppsNsT1BYF/WW0oxrux6IKBhXZmRrAf8tr3QDS1NqIYfy0Qz8NmWd
fKBzUZ1vGTDNtO9uo3Mcwrm5FhiFdBVr7ikPQuMQ/mJe4zxODGuH8tYSSyFkjcqtfZwHv04vVsa2
o07G6VMtPjRwMpaqUhJQhdVBpY0FQsfSZW95VKZp903AFyo3lpOoOjXJ3XwvVrVbvD96H5l0i24y
/KFdY0wgne5o4M4tIzXrwkwIisYOPs6PtyDmTXxEYz2LJe9WQvFce7z1s4NKE360MW2LAHFdPmGl
Sv3s2E+0MwzoTAFF3+9PYt0Jg2f4kjRToulXido+XJvx3JVuI6BBVu3B9t4UzucMqi8pkjzVFXeN
MIHEgl1/yQbELFKwHVCePatAtVG3+C48kVjGkJcMgaBUMa/rwVpc8dMRp5fQB1qumEQK1IfKaQPf
rKU89IodiKoMmcH7VpsKsF4kZvteFFDXM2IlQA86i689rCChBMdT2p1phakT10wo8eImg//ZoQOx
fUFc/KX54Mo0iAufZgiE0fTPF/RWyyWKOWNzombe9RQv9ehVY224IDrjfv2AOueIWVakU02GT20B
b7UP+1b1DWZF/B6wfS8tIxpTmRyA1kQNlgisM4A1CrNDDkcIKjIbIfwDBmX3etV8+v23U7oys2OL
yqeXd15i6SQKDqTd1QeeZG9EVfy9+nJrfp43Qdgl/Fb2bwYHcaJKcuBLxAxa2ve3twMPOqWHRaYI
MYlgbTpNi7WuZIPERzWFvCE9SePqykbGOg13hbanOoTS6cY5TzKIWUF8hBQPC9AnnhUZyFAEJtTz
ZZu7A6QedW4cqWHoxxaOIcCsT1EfFhv2iswsGGiOl8IzG2Mgf0TmSe+A6T7GCBjoeEr7JVXk0I5m
EJOB+Y9vg8kMEJR2QtX0wCuT9cW1MFMk+Sf1VQTe2rOObvVTqNKaw7SPgBISDiaJXC0ywDQFo6T8
InvnL8w7kuyLfMAr6oAdPLy/JZHEZao4JpKLm/qXBI3tMdcnyCxg5K9k/K2sInqbpl5skwtLNQyc
jcNnmmnrcJLVY2kSXtaPO7Cbg2hgixY0rACmRFEgdowWtDqQfZ1qqKfhNwwtSGrWU+qdHUDqzdto
KYAP6XDSAbWfNUBWU/kniACb/XkiAVpWUY8HqHapInY609J3hZ5HkfJ4horbljoL5w227BJG4ABR
130bYp2c+umYncKzDWBf38H+VwJQOJ7xNyfiuBLrlI2LciNvs65Lvljg4IZtmXldTJ1VYGvH7+Of
TQ8ncHObsRXmuDfi8LzgcYb4Fn0LSM1vzMVudK+OfY5uRf4rr2lnKBK2iOjDunI9oGt/GaIBEwTS
dJ35pHrNMvV9YO8BNnyU9/SWYVwCA+t3grAMdZisSWMI7dLk/3ty1qICdzrhZ0PnHbGLEMjPmv/L
74uhnAiR0EZZH1z7z6RoIKx9Z9Yn4yAkkeTKGs8Bjkb1L4CuQzEaOFNQA8ao5TahZRWO1vo4s8In
k7mYiucXe6g0c/6jF6TLIYPEQ6Gytlcg2LzhMTCTej8uzeUwNNe4GstOLUxT3qL9bYV77iLhjhzy
tKsu+pzR5wTWhRTnq0DUXioaEqyNXNlZAVUFyyynMsLGMRGCtVq9FwpnlcgmjP2x8fr7KltE07bB
RCS8JbaXmZMnxjde/lDRsfjrM204w7MC5qU9bTfXm8G3rIq1P3mTFk2g5GQeidpwo05ASdRr5kt4
veCZWCPbq/Yz3uvxxGpi1FN1jvMpVa1/h+c5OKtjlN+KfmXVZG0mTueW3EjW/FVKnXN3wp45A2Fd
S4w9klti1yTZCK9z8dcr4o3+Ize7KzpUFJxuSOpQ9m5gJ23gLQREazXCk0J5FUadgU1FOX+vNaNY
1Wns5t9Q/8PJUfcS68xEDAZIm+FPPq4maj6+pw9f28YyioOeidxAxGdrzUwpn1oQfwv7z/dpJCzl
od/RaIwF1YKecyTsKmVWVJuvWC6+US0f5U+cd03W/tRsPGRxfrwu7fSezqmXycFWw2gNjozKEDh/
VwZrKT1/f1SIOBPfk6zf9Bg6wEFXC27h3gOspVuBmoJt9ATYzOIYcX1mmEXUKEFWbjHKr9cxKf3r
G++lwOUOOWWCV8CAKw8otTNfhFzvphZLijhqJV7+ppbPHyHZro/yQQv/uh7lEBRkyXOliWWpNAXX
uvqrbG6kFpOQPIPHIP/kx6tdbIbncZVXkedWwTj1KbriuJ4zA4dTmOFdekdKxuGqbY1lBwnfc5Rb
JEVGwtlOk/o9jaXSR4eHhIPoB6PhAM+eadPOCuxc1Nnpq+UaaW2daguQYZUGLJjglSixKli6ZZFY
NHmt7zA5GvlJDM8NrlZzorxlqvlfKFC5QcF9F6R+y7T/O3pCXb2SjlIFGjhpLxtTecGbYQ45jKSi
3uHZfs1c2rJGHkV/NgScFe19SuWxP4TjXtHeBQ0hW1Dk6JVZlBiNLNA0hEYy/OKn95IDxUVaFRzv
qnfBTbb0Bo+LrrOJ3NFxQNAye3j3u/0Nsoo2Ro3u04upz99QhQrx6DSiEXESdCMCyO4JblwhmG4D
ZzuRy5ZmlE9O6vbi3uX1kgmglZgGaayY5/7NbPdGv8oVgD0azqO7862KzzGOAvkEetvZ8n64tBjm
g3EEJ7UUYtrQIAtJQ5t8u/N2I3TjfwBbweUdsHlE48/Vkw7rHNBJbbUGh+A3rjPzJkfs8NaK4oP7
YWT5GBhWEo6RgsqJNMrQtyXX8uL86ymyaEV9Dgh8STGH5Uc+byt7vXQde8T1iDmXKUsckh8ZezOs
EiKMrspMfV7v7DPo2uZt570t/he39e7udTy10h49XjrswoNLfZVkEnOKa18xlN8DYjz0x/MYrHMb
QYn5mgCxi1UnmkKyupUF3b5Z/tnnWpGQNzzghWaWSxrE2gtiBq9tgbLSsTUUSfl8uEOGb2JlM5rh
Gx7VLDvNe9/N9hKqNXvgHhAWbTCdIrkIWleB5sM450V01z7Z+IRYCDl51YzWwHOaaQuwMoS6Xb5F
Ad9fMMba+IhSxsPe0cm5dADKA1d+l3s+5zwotRV/t4naj2yRnlNCkd3KhMYGb7TVUf5rmqCE48TL
EBhXCaqDVVB5ePjyhYcEudjPwjTA0+jAurgi55jJOYKBxrtgoiOKgejygVwqllWzjgSQmSDvxDYA
ZpedNY4ZaQwO1aIBxMcQnCwwg/1waB9YfnLkds87nGnmoKgpgUlQvkSHBVzqPaMa/nUOx5B85Icu
2RbA01WbmPs2v8CLvnk2XNFFGbQDvtm5f1IvX60LSVYk764qFgXJ5l6y0vUns8vfRRljBAe3gnRU
DL51bvkcjkk7Z2D2j+NzLefsf24+XkSHnyRWVQ2mnPwYHnYhFOYUbxZCilZA1dQSB51pyMA4UIiP
RY2Mrt0sm1ILKIUuSdWf1l/L4tauol0AHH7fRQk6QDr41m1QRl+UUG/KRM8Muq79i8SGWH4YCkXi
jH/icBG3SxJgaOojW/dekY69QQpqxIHQy8rCViWlng2dJrUJWUoB6Ane4r0PcnwoAvevfLKFP2mL
kBazwjo4QgbCuj1X0Y1QhRcwothQyRvU1XF6Uo6Ak0JM47CNE+NHOkTzexjJwWGzQFxk8rZ6FYGU
X8xHZGUmFLHJRpD96cY2bwq0rfqJc4lm8IJLfm8koZk2Nw+2tMQKC+E/j1Yd2hMcKo+sm/wMlVNo
VGkL63vXiMTyfClW2njKNItJOffUbhwuRg4ICAfNxWzDnU0SmeqRDqZJVeR6A9sp1nwoDnCUbzfi
dVLrHql3v+eatmycBZtCzB3lAZ6ZTqt1PWxM08yfOdMA5xEjwdZL1NEt4yTthPemZwgwyEwUhGcc
3VeghgXg5bfJ8n7fy8WNsuLFIZPeKi9Ub0sz/ZIMFTgnR+Of5tHJ4m/XYK7pEvtQdPv5bXnwGAfi
J/GWZisSAd8v2DpLokckbPa7d3miUePjFPpfdqixI5YGbEdpKap+Hmm0Fukhu3p36xWCRJO7puX3
OfWOPuFlMI2jOzHc0n+0G521cQs2c3VSMpsh6SGDrN+qG01BM4bhqdDLlSqSX2NRKZrcG5tA2tW7
ytj8ikNz90XxbMLbjOh+MlRgmVYaW4MumLrlgKyk2+Sa/SZvYwTxEV2cEbk3mmdB31UQGeA9VRSq
/QZ5yy0qImXidKjn9DdsgtkwnIhpZU57ibOI+49xgd8dOiEmkzEyeJom5G2Nsdhil6VtrFvwPr1E
jVvOvR6y8S+dOk1XBIdiWJ+5EY8Zt3gXzuUr0gYvQdIZb5npKpuAEGeJyJsGIRxfvvdv4B4YJwe7
U8a4nU7oEcez5dzrPWZnWyXsriMGV2pWvPNyH8j8urdVeD3z3dY+ARyHM8kwz1C2i0WkCK1cXjyK
9vsICmslZCgrCXXRFatCZRnPIUFyjzQPKYGH/MGOU/YrXIl4mWFytky3I8c4/zop0472qpSC+5yp
ICwIyjC+5218k68c+J9o96kuwHArLB0XX7hCMCNC1pCTzb35Txnj7RyEEGSRXnKzZsEBD0GTAHnv
8Mhoh24Hp+z1kUGDpwWNtjUSVIBPFWJxISS2qFohcnr2VA6Vnraqw++VdypN1d047uMyTpL83k1H
1hP29Z3kUxSoAI/W94kV559GhCf0q+VwFboSzlosLRHC7yin4HolkTQ67fAfAwXImwDcHZoqAO8m
6nAOzXM64xEBrxjdKIz8byZ8V0Cd850gaod2gV4hCgXCFj0Ebbkc1MGp5rG5uzMK6eCfcxuta92n
wj/nVcACEb6fV+ulo23iSP/NgdQ7eaHOGOmZSbXdSoHHMAqYS9Yj9i8oWnNrqm82MJr/00nQuI98
Re4MGkTNbOkaJc0U63ibzbm9fyYOCsGjTbU8PWugExyZuBKnzyfAcMkGhTQERTOYRGVs37/rVQzq
CIDtJ7rtfWM6YvMEnY/dGB0TTq9PteL+fLxO4ylrlRFS4bl+OTHksqt9o1xYnVQIUMH0cBpMKf30
jS+ggd/2AnUudWam50TPBv/T4cEeWEvjbIQ+5/Ct15srGfQLWBS/U50twpAcn2Fz3UW/QuMyiOv8
Vhi04zBrSTDrO4xLlOEeV545RJkZuIZM33SQJVnhlqAT0dHtigSShiLOOdP+gXFsmJxrJTuecTIC
3pLqzWzd4k1ZgdsElHMU0bTcLO5a5aQGegO7EKkZsZ5SRNOCfbJNpnGPCPXiBgDbdDArpG7uNBo5
633i/pkZAwnNxgrRDUg3nJlz9KZF2PqwLUrk92BmzZrSfDaZ/LDsh8anY+faW2raY9ubg55HIWAf
bdg5Em/zmSMuOo0ujup5Ai8prdf8IgvAhAerGQB6Zg4QF1G1nIaW37vF20VEyEphkUGK1IiwiOJN
l7+5rhLoGjB1h3Kh4tpp43NbOb0tcN1YGklUe0EjZSQczoepX1eatMAikbhl6AQyNyhLB/3EoacS
a0yTwxLCk89rQ4WykX57Ms0EQqo6fEOI1plsTJLhciTa43/OQaNQprAsVLIzOu0l4ywQMVRDofYp
3Uir1s1lzThaUXs2ZKULWsmI7SffN3naxvueDR24nPasTOOtKsy/3IkhBSnXf/54mtz586j8Rvk5
axi9qzOyCYsY6L3Df9LxcI05HvReFX/WWIPHZoeCnwIedNHHMQap3HBGBW28+Niwah2QUMd1ivyv
QjGtZutmsKR2/fMTaPNHmnn0VfSG3tQciO4W6zagoTOm5mNLpQ22vG5Cko9as139SAYz4+pPsu/M
41ZnrMwgBwJnCupyY6BXsoYIoNrqljmrqo6YkX9ccD9Vp+3ai7lWsLkNmXThKJvg9BdFB3JaL3lK
uxsO4TEEccydrP2lsT95MstwASCVUZ1wxYwi+MoQGGdH52OIDUA7nQWr6mDlB17VKt58hQrZBQct
iQf0MCwrfkIhOTmTFqVfGLepFQ9ZtZckZvadQsW3GETXDPgCo0AQLKUOGc7Y4IlWR0BtjJhFqS3f
EiTWkkuiBD9UfgrCG75hGyjB31p1mJFbmUCQqoFtMGRgCqnQN2RMfgJ6YOCGirVTM+YHzIIotcr0
bXOXO4p1C4kYLT3kTkFSzBiXrahDZsqTwVQivMhbamoPBwlg7p8TUsoM76WDXy5Moor/efKG2c5+
AC1jyEdMPYfOE9wwg/VMjYOknYwfCsUPGLSKVooY7BI7Wl7twBLeFe8rSk8Sh5ikXjgcsgbjnUkT
LtzspdetZjI86+ZEr0xJ8JfedkmokQ8mRNEpDH1KGBcC4Ut7TQ41Vp0/km5R5Aa4VfCP+yS58XHQ
dOzD+zVd5BP8GkC3VmdcLErczZ2h6gmEckC0CENDM+GJohHq//vHCwXEMCDEWjbJ/BpHMC6bpDXr
rLU/oEmg5dlCGvfv0iggGBB+x8yOApGlpazxqrO6uJ7xorybFOo1bDBZabvmbGN67q4Sw/rJA0LB
Vten46Q8tA27K0O3aKVNfJKk8d9PzyEwLaKVCkx4CdUIRKEivTLmIUaNH6F2+EqdZQjaGEwINj/3
n+qC9B5NHt47wfTKBYMRwGWxZ1ez0PA0YQNQO16Bx4BA10JePfnsc6oY8/hK9tZ3Fw/Xmjv+HZsE
/Ds0q+xg3yVt7yiqwX9GLZdyOWlj1J+dX/JwU6cpGNKF4vAOceF9yEu/cDtqOtTzEmiumMsu6k94
lBc5rBwaBrXtEXZ6kkJj9iCHQ7zaPoFewvZr+NhRyBfqnQqR514HH3EDK76T+c/aPBT6O69vnG/X
EF3WW2d50WC0zi1gMSzl0yPE+g6hEI42/FW30dhpp0tJl3NFmpEjVnWUurWh7LQ5wMiVDqzmBYDH
YmlxygWki/7GRZlxJwKXaQlGUYYbjfBA/Bq6Y4ORdo87LhkNw0IUOq/GPodbZ0HyUPEahanaBFHf
47oHUrZYFJSQZVwgspGNIg62cX3pZ9YAmlq9QxBqKcS44Qi1dnXcfV5YtJnYblneaL3WPHJC0W20
+xfJA6tyFygG7+7+p3ENYVi2tDi0QEjxd1oYHPhiRlLiVj5+5PGF7zqX697Vc8PkPzU+b7FJojIR
oyHLGxV/IKRWwDtE4sAxvuGJ8FF5GWoW8UXE211BBWOxlhmbkRe2ngn+m2qhgnO4ukbe8JJB09k3
adaWgLBpx7afgh/ZiVJ7rMkoCqDeflWT4xONuuHyo2KeVdUKGiTgIqBub2lxJ2IC8VPcKeRnL6sH
TaJeGksdQ4IL9wf9kpQ6ml/0/QOOKzs9Wen9MxhieN9fqMZ16Uq1ZMkXKiHIJU3o31DFCdAHkJod
5z9i7M+h/X17DVPV8TX+LAqJzZf/p0B0vpyFgtiPjvZ8ZtCjop3ds+mRo6Ivxswg3k5lcvXL6773
T2qKv2RtT7e6c8zsjtAa9Ivt6ELWjSpsy4PxZg3Bxp4eyY6LPQKsqVZgH3S0Z1Oi9kwpWgiwOT/v
SYCMGuWeDwXP86Ups83ETYvR2M/1NGS2BXDEJOj1f1R08OdWv9yxZF//ekF9wSrVClw82wW4b8Hh
YJx8VKS7in9/uYKPm8x+UY4/wY3RQKpvSUHVnRt2My1M/dI4kY2zNvL5wf43ZpIT6iN8oKrKMtUB
/zvfwfFMwCsQKDKu22Hz7QR0h2o1j5B1QNH0XRK1Ffzf+MsfNJPTrYxoeUp2ytemCol+hVm91+i+
OV4sqsIgKptl488cBcjoHUTRlLQSNOGhfghPv4zh0XUR1uqHUiI0Pnfyngfs5Wwpd7WoeThWR7p8
kA3Au6R1poW4PR0I1WDuZalpBHWU4UMS3Kun5Xw9nENh3NxWyA5wilvkTNzmdBaswZ8FP3SnTaTL
wXUbzciOFxsBtQ+RTl0GfLBPZDLQSqswwF1k9BVhkkos9D696uNzyaVByBhjwgWOctt+RCOG8nVr
U7xWoIb9f1F4M4R9Uo8sEJGQTVEb8Vt/SAFTFLVVucBVyJX7XrwMNFk9cw9Dddmo74kTPaYlp5To
sy8tWeTI+idnUiRLbNsSIZfkZbbAdu0icC7fXQ81U4S+Q3z4xabYZpkFXdAV2QGzd25XCe3H+Ypa
NkUI4CAQyP7r+UUy12nvm8nNWt7YB26RpmkxCwO8huGwiA6nhrB0vXPI9hqQH99Q1QEIbSDvs9Pd
s20u/wsqnnaOTQ2J2uwWnWIi/T+c+5nctVxAEOYaeL+o5rM6hODQ4iFx0b95q1HX9QN4w13s6HIM
jJ7d7XhogDJIe0FaO8V0NZvYHjGRdgmUyjTfS4F2/uR//AaAJUeJtTpKhLnHjmhJcuRLpUXS9spj
RaOgSs8WhmU/nmxaRSypsuNTEAWkXXEyWRhqNt981iiNGM/d/Zc4aS3RB7JyzzI/FxAeuJAe7OPc
6Ony4eeTqeYO2VZF0hQBtW/tsvYv3nsTlr6DeR+DwA8/+3bvzffw5J9NkYcmIcfwtEF5b3sv8xN+
RpQWEBXuo1t6UYwM7JmYo+QZcErOah8zHmxiEIRQoYwJSYJrQp82dLobciSmIW7HHHV0DeJNuOic
n1M3OqRVUH6FaS2Gkb+IqT0pRdxhbhQHvdgJOal2NHwNjPLcC43K17JTf+/YR9uMOAbg6roh0q2T
RdQDvOb2DL8nistd7Nf2eqKDwyRez4le0z9xQFrqo9GnFFvdTC6jRgtA/p32LQza0nBrF25ymvbK
k9egQKdUz6hmajDgi0yHd5jG1utT3XVUhP5vexyORZc8ju0JwaoQrsaDEayO3OyYJ1FxPjwPCkKa
RQacpBZ8zF0DReYSVcqRanvRyonCbdC6qRUvW8q717JFAHaVQvsSgZg5n4TuWlewE0sTygtrO0UN
49TsHYw+kHJHYU7IadZpeuG5LUhdP3fTGT6Lbh5xw7ylOOAB64nYOfXaCqFK9DdbM5Y1EbR8cXwt
Bnp0zVpDRP01h8gG5773izwSDL6RQ726LzPGcZt4lBDdFSEdjV4lwCzDCzgMMUu8f5Wj/n8pbz3W
TNzY8GiVsgSor/drdqccYOqhPzSTNg6HMWwEZekD1EyrzX6XiayxHPPWQ5wD7+/+YXkYJdYdSmCW
YmjafQUJECZn7y1Z+qMaQYMtJ6IM7+q1YJwyn6kGmZpSpyRTCDNNBavgswIRYlg8CmnQY70ykJtK
gxIXjb4wErBkOHmtrCftDdjW8J11u0YTXKCtOpQ5r+F3VGxPuibWaWNrZO4cN90MryplLDioQm1q
shpxuW5hOVRXCHR5lKhjO/ikiQWaCyuSvwM26/5ZOsz0nXHDhnpqtaa5uMra2B0rjkQP9n4Twmz0
wOf9XeNJqV95LPdLiBFqyi/UJSHz2JscxcgDzfrkbDZI/Dtu89JXWm15zA7gS+xA2sxI0IyWOWU2
33Env9toOzXO3MOfkG7jpIpGrZEiW8cp3FxvcmceeW/epODFZQntdDLBItK0ba944pYxnSRxOjCU
8n8ocNPJxhwZ1cWCDihcWcX6dQWJurfhcdaMj27/UdKpkkAbxRvH+9LpN/9WjjX8EbTV1qj4qI+Z
ts7nbUx6yKvqRSQgiwRj9pTneHRWUBG/5QjuUGu75GGWP5CXIB3gZB/cy10YE2iMAJ9PqfHyXFTr
w3uE0eYIssYfa2CeUTIY7txhEGcl85hBgDlLU0Qp+USALGSusiRQczp4oA1oQ0lW+RK1ZjAdZieV
2h9IR9eBwP857FjKRdip0I0ZgibZtOLuAhAVS4/qmGoE/w9c1TtRaRYac52DHhKYrjO70cf31dY2
kcO5hQOCl7P5w/G67B/CbaLx9IZ4xBWSSo6rqk1jkmGxUQQaf1EkYIxzdmGPKppBlF8idsA85jED
+xxC8EcErMy6ikTmEVLTR1/8huy6LBdiwhBmSScZUNEUOc8yi/Ac886F9kk5SfhPfVzcpiJgW0je
5o2A8nGKKViWozHfgjp2WsNKM+yE1PBrqLTIqBQOKUSVpxcTiypRlMlbTt+QDCnEnfNdnlzWDMur
SaSoPRhx58/w+4M5ALCx1I9Kxptacrug1eZ/jFieCHwsq/cCAZ2RS+FXpVLHuny7Y9hbw9m7mls9
faI4ShOYUtagjc1MI6EMVM+Wqv2nOcJAHcP2QOnlKsUj4+qyCE57VB2LWDR3Tpxpxjk5SmcoN2pA
mSQoixpnh0icZMCV5y5Y55CpnFunDbv8EnKbZ1bth4ikrAjcw8NxIoUQ3m6XFG6KhCE8PKY6nl8d
cO2faBXDoKHXDmfyHuD17S42CQrBLudL9FCVNuFqtfGKfjVIpR3C7bEQfB3A2zvK/BnK9VaOtLhL
g/ji90tsmRaiin+LZhK5DNnBaKIy1a/6sm1vErTSyI1fz8xvl7Jy2buBwksV4iEKqicfS1E3Gd5p
yyMYVOaEpmry51TYpOGQ3hZzwubKB7VEsIofXKbIB8iqdDQrG9uf+oj7BsFGoZzubSnl1xCZwlyL
59x5UKvRPDwfDf0de5uqSRiQE9AfgY1gBpT0GDIQ6qme8ojqh2/8WvLRcJM/A3ZXGAHjZJaC8Wt4
xDZhQ/IUXtswaXX8AAU3t256wWu0kMn7lY0dz/7FpojGADJ3HqAWMKU9G6vboBPQMqQGhW1MxkrY
vi11Jq0w+M5Fw42RFg/Paayuk20iYkhSG4EXpsIvMOdHJkaaPrGkK/2McUYPf7FnfGrQxEcI12gZ
+SKrzR5/AphHSrsHJF1qasX9xcLlliL6dGcpcnh7wVDK0HF2cOShrdPSb4WnGBrujb3XWpYg+5Iw
cbTWB/SfIMT6S0xev+VQN6BXbbZXsLqWj9IoO7GY5ofxb0d456/DkkXKxuF4mx4L6pixa+dhZqSz
VhKJSFas/yU6a3MaSXTQO+VfO0PrAg/fpV69+ypLcjJcovjBWbY5zb5OhF3fTu1qZ1GN38N0rCmp
FJEVV4SjiulFEOy4EFlXCdgJ6nwVMpqdvQXSTvKeXaJxmSm4IkjHAj6j3ae1zicVj+Cd1DUodiVA
B0/CB2STPGMe/tyVEg1OQDV++zw74vFWI24EPuagk7hTjBE5V2tdrmNRsB9UAbBhAI1f/tpQG++x
L97asS7TwDjqrP2iKxLRKTTXpTpfPnEI7VRHk5evbqSwGszjKmkeCx8szXxnJcjN1F3q7CIj7a+z
RjvaayxxUl5OmceCPhlAgzEyxBRQkqJcL0n0kVICO3+/RxwdPI3r4UJM/uEdYRr/3UqrIsKsgacT
GUviL3YtQZt9IQarWRj+lyqVVjeyayyk/E6iVAfGz2RiCFdDV0j1X7synbs/zNmpNbIUCSwaPWcU
avSwpYurw1dn4UhqEbHk0Z/N9iy1FPeu5wTTb2Cl2/W2aLJNY+tke4y1+AA8k6f2xpaOK3mIggzC
/2lyltBK8OtLSBh+ZLEL0gFV22lJCWX1hVeMTfFvYqd9vnfivtykzZQOTSMiOdtu8RF6ets1iDrj
F4WP/sA4/+SszsOj4NlLAizBdWn6SGEy0W0+0LDDP1ukOiErZemQrt0d5BBGzaZIZvNe1hWQBHah
3IpgMWaxnPw754+GKYOtJ5ScTDQWGzssq1vGvcG0L/OjTf3Hgi2Uh798Qd34W71BjYXaHoCDIqx6
c65O2WIKXu8J3kc57ANyv047PwDfmyDLmDeW59Dc0Lc7ZkSxNH75KGVMMDkRAyOv5E6lX1ZzVsTJ
TDwEHqsAgtQL5f+x7WmCLBuRvV7hNfx+ZAgFTsnmSVqhJbAd4pGKZ7nZ6xLXgaUlicPQt9kNUx7G
KI39Hpl5CNF8XV02IJsdiD7RP4taM0C9rtLLdc61ayQB2ddrm9OyZU/dxEdmNhOCcvR3vL0a0L7R
vZmeu4cpOLMwTThiUTaYiU41yw2M1aulatYPIKHYA1nDKXaKWgRqH3BGVxEXvTDEQor3I/ZD9jFZ
2dYo1rRmgwekJZ3pz6Iyy4qw2JUBHfcF8/xYn9gXQDFDri37LukSvjX78Z0tXNHcDRaz2GwG6wYz
1r58ikQYBk3at3KzIt+34a+Itz2n/dgOyBYKwOUTSQ4XNn4aVtJ55Yvkshak6+dBg/1YVd2QKYOX
yjEBIm+wowsGZBTiwbFzvf/rZzcYQLbYXQOAZJxjLsvIqhHL+tcqlptxG5ap6HNES7qp9R75FUWm
8oXCWCYcFr/OJkWA+eHSjkAqLquqD5ONW2FAmFUepUyOCPXNQ0HzuPsRqmBH+ZezKx7dUsCkoU9+
Lv1UWfFXWkWl1RDW7+0zKesXU7HvW3DNI+dixmBkblmH5Y9O1gX9tFjtzBY9PpmOy6JyebC+f+39
3qGg9+EOBMuZyOODduayk1SDLDl6Y3GZA/0bG7eolrUk3b1DmY/k+d+bp3rZDTqasMe1CPws79DA
skD4w1r+ZMdgbnCfHeveHSTCg0FV7RRRYH9/lwtdO6rNH+HSzRgf0C7FKeWc+wYQ8LvPpvuxTouD
Z4sOoKRGg9iIC+X6/zx5hVtqjlmHdxpPGKl1r+j5YIz5j/PcnuSQ3pUsr6ZfoQZ5LmYMmNykzPFl
5LsNuTLbQWAFJS9iDKD1tC/GNUd8tEqw8HkDGH/vjrGBELLjXtCV3+XKp/Z0rcDFqxyUXXlUFwdA
8SnLb9NbNz55c2/VCOwnjoL91X8/sygG9be6AMpDkHIlzBQwVUd3+qK8cR9d9xhluTTrCfgUY+NJ
iwsNRbe/GjFhGZRSDsc5ZUi42iNwk4Nnk8zTCyt332YKFmemcHH23LdT+8eKBt7Z3tAJ5fZ0pyid
SPad+LQAfguxfUffkaXNGxkJpCRR2iPyA4GOX6z4uWhChwCzglFurOKcKF+aO30/xwDqM1HD2t2f
CoS68tOjJEZFQDVGnpmGryPgRdVL7puacgrCilbqTGkFcinr7ZEG9VJneACOntRFGQaFfXh/fVaB
rJFR2yxr7FA2WZyFA0P0rB4ASp6SuikwVH8LJ2Caz1aZhlMCfMnBf5OV5hQG83Jt86F7T7vyeI7e
Q3i8XX3kX+xmOxJu3yVWXDyL4U7oTb/Grq/uus1ySfPKX1aoC0zuBLbI68SWN3uiJAZtZ2nJ5vIG
3pSZvFMWkAPCnnzPzTtssoBvVgqRnw7fYV5p4CigBLmdbalh6p00OPis4lr9hRc7lqb1Bsxq/kg1
IEx7Su+GiJtSvVzYBHI3ql6g4BUZ5KFKyxSW/s0ho9cIIm2TOfaXCwBspMF9eN/rk4WiWGguImz3
7gPiVnxUINVoI10MTR/dvUqzgtv3tkp3KezbY9lhiD6fGtcw4jDQWlfxfr0oQkmX7Jh+78B/CXu9
4reIje3klEa55XWpAeQ8KB7uSHeJAwm/S861WcSVzFKn2X7lqSCPLJq38DC1KrcxZkzMsiwbbMuO
lRc9FRM7i5GBVpHgNuaQuJIIWNMJGWMCpN7BRTpT3+RtW4mU/k6CcFr1jiyqU0vCt/t71blCoTol
cc2EgScCWRNqGC40myeOgmDbpyB7INP+jzdRgH7ETrmYLbwismPoKUiFAJxfrB6d+kqvOa96+5IT
n5DUv/CJ+EtHn3aEGRVV89kO6DVwi7UlTxriWM0oRMMJJakuWo/+KP/mnWzz4mU7VgElClwa38c0
NSwdrSxXENPtVgq1mnUhlmWqXBmFBwihNfig0QQFyrPXuvxv+CyWaBufYpBr7Cz+W0T+5yveZ6Nc
drykD84Aa0Omf3bBL6whxTuiIlvfuRMg8rVTjDAesO8iSWzs3tpHmsqBsVnwvVvLbo1DCM52DKOz
XnXj61eI2Mo0sHHHYv/LTiQBeBWCL4pVSuKZOifHFTnJ8owK9lIfh5RPWyd/ZPMnt4eux3aA1Mx+
bMEp3ESGrKsSdfAfLrCaQ+OaYR0dlUuTDnVKUOqZrbaCEflOk3kr9OkSAteVJofx4TPZN1n73BDH
9zRWZNtmdUz0wlmdeVGZTOd5DjrIxdooTWqy7/+0B3OH/jeu5JJ71r9Mvt7BhinGDbFAwvFk9q1u
X3V8IuBKmLQRDRa5Jnm/fMUJSOz+szauzjVUULHcSfgkbqp9PpD730TmfuryMq+/64X+xVAHYDut
N9N0fT5CPk79T9JbNkLfGgUgzPYUFVB67SD3BR+cHqgmvb6xBh2/rCJynnyF3Qn0RdGv6JvQsdbe
T8reweSLcGJU5Oxd5+Cqj7Kc9EW8xSSbZI6wfRHsFN6KzgP6c0gAfB72kiAe1yfKy0YEqp7U+5OS
3hbaioSsOt7h+tGKrrRljvVRID5xrYFfXqPJdeio4/0gvoYEmjK2eeIwKSql3X0QAg77y16QsXs/
NKnrOK73nUqoB7VyClPDCHGf1FmFU5BnmAp6VKJV3n3r+xVhVWBBlayRnvG9zctumuFIUf3aVoxw
3MGV0bttdYmHOGoC5FJ9tT+PkUa8NAajyaDgT0P2esyQFnD8fZf2k5SitSRCadQzRtO4VDhl9F89
xpU7fHQ7WGPs97kaYxp35w16L28UEO+gUuVWE1pj9534Bx+xW7fqgF7OrcmGt0WGelrOV0MjUFBQ
0PKmaNE5DxlsL780e2y2wHf1xwN7ify6LjVok07swVsUZzCCKCxJOnDmfIn+GVAU8tBX/E6dLC5A
uPeZLxmWJzQh4aUYq4q5ahgstQvo8qc59dy4NoORNIkUUIIMwDdXioYrAeAygwxTkuNx2EdOgQ4f
NC0/flI12Tyb6aYVVijhs4JzK9Axwftq1RcgtaePhwsgLOIcWOsBrMQSFCARUgIb9XNffkZMGVRV
2HiOCXXeLl3GZvh6MUeZxIHAQQ2iXlY1EYKN6pN1l1xYnUCjO/4BAy8+HwFaIxHUR/2rDOa/ugkm
cLPeilkSJPy6KXjJRmohE8j2FeTFlZatljb6rRDuJo1T840lVJIXIl1y1dHcWtM555jTGO3f41yo
NTLPPtcZNfeQsgMmPnCboM4cuRlEIEBrkHV8W82xE5vZQkABnBdbhKGJzTHu+U9hLtonnHEj42Vi
DHR3GWqoWXdFXgk9+RLjRCXS7OWEcOp70C8U9qLBecE6vq3/1CCuLplTmLEAzBG47ihlOQAWUnBi
N1qwLvcKzpOzrj7ZuZftD5PApGJ5/6BPdXbg67RDjcYVHyLOIYzo65WIpFItNxwlFm1UVknsoAsw
105DpoM5s5X0Je3GOeDJrO7yJxvN8pB/wz8XBZFQgTa+3d7bhfMljD5kX+bPp8g/HT9Hf232LLY0
oLB2AqSI7F7gRVMNwne5VZcLfkdyShYuwylM+rGTpMuLwgiN1p9H1fXb2cOU3u9Qu3TopJOlOHQl
zFge/NY/nJgq8vn5ZC5Y6HacguAERqaPrC+RdES4K342Bo5zitmc/BHC32G9mjlsDEOnmdg7sQPV
YrfG2u4ssR64wM4XlhLFbbxUwPmXnt9kEqGJewkKqgHIYlawsBJLb7GzGm6L3SbrEd0nMHpMgfFW
t9c4q9ntVz8GNnZZXt0HT2XvdfsKphGpUinJCMYYuKezlwHWadZd60I6Jfk95WIm+37EUa2+UmnG
mNgzTX+VzPSzh9MR5ED+dC18RcJEsD/2K/e3BfeRgZ3smdL7gz3KKVa5cFfGlNOafscFgz5v1pvc
WQVICG1qM6o4y8ohIEiIN+6ixujmb+7OBAyMrdZRd0qJDTLIuGEFV79Rjj4amsUCGPTk0Wm3rC5P
E+fiGElFXOZWds4FxC2F6qAc2h8edq1PKT8+yf8QB/ARzq85TBlJc28oGgoTjPAb0XLh6s8Wvf2U
MqM/OepNUa+MgAFdu1Hh250ELSqZKmGBWpotuLYiuiIQ/loPA7cTbqOkCD+eCm1Hr0fz66VbJLPM
sr02GHkQP3ZhdrJtuSu3aSRX10gm/7/KDufI6+qOHoM3Hp2gyOZ5VdLUGin62bpDCw6UCch4ZfFY
QG2oCjE9M435LxybIzrmhL2+eh5SqyULCll1lztFziArxiIZkZXLaZZAcCYkaqEsFaFx+pjwYTQA
8tdMdgzwTpXwqeqJ6KB1H8T1y9ttOJsagSZX7+C1lB9VP57QtprKyloPHGmF4nHAmFAng9sB/Nwe
X81ZZ8kb9/fWH3dzTQbq9A9OhgUT0SX0SDoU7pgBSNlIQcMMF4Y5W5YAc85JwtvXEjRAwgjPekVn
8eNDnYQbAw79u+ZlEYdvmR14c0yAhlmtWvCp4QsOlqE1XPXCHqTFhpgypV1wsFC6Bqkim/buuhU0
k7uDCcKXQsCywvaR2EJ7Glg6v/98dzxM5HI7M8bmYUFRfHLWyDepqfLo37sjiSAqfjWsiKNTIePU
UV4tRhXSPftLyhqBoRCKS2nI/BL6qR7c+uoxA5tRAi7J8pbV1+667pTX2bJIHqsCjhL0VHeNSsJY
9WJ4Cn4J9otwDcqe8LGGKrUupKP/P5+P+jEyNzS1JzXTTAhSHyMk5o3T/H0gLu89aEACVPuE+sLR
NCZ3R3+DDdCEF7CvlTe/2wYXl5rM77jnRxblKU80ZJ3uI2VMEWiAppNJ3eBVgGFom6NIP2YAfqwy
AoWRui1gLJjElDyZK2N80Xouz/zv2rsLyZSy/i+Dz5WUMayZUniAm1O14iy904wLZEoKkKr+fbYO
7g7/8hQWKuIcFtmkvXQlDICEahqhd9ua9Sb/PACtIMfc2X0razJKafTevWYd24vgVDETW8arhaHl
WbfFNtpOIdvpC2W1N/7FMoLV7w8kq1OPIUPq0K1ckR0i3C7CiLlC0pF77Id6plCw50nNPA62SqFH
2IW5ARLJbbon2leBktlY55syEHHnMRdjVanM2P+kkXb1LHZQnqHSK/viQIyzvwSVk/L7I5MKpLzu
AmPVuJl9tvq+LuBzMnUKtjM+9Lgf8/Eoq0LP7Laxg+IaEPzBXSLmuLmGHfR+f+3KwtYu2qi+NUIl
OXHbkSx2KE3YxpacMwnD4YW72R4vH/aCQcuWgTgLz+d8g6WimCr6Lm5a2HIYTkH42HPF0eRMNxcU
0/mGicH5ATP1wjAXo3yMpgf4LRcybD2AOWT1xpzhIusSHlU98MsritSPsN10Acaam5HVWacGQx8N
mnzl2VQrsOhDGTCOSCiOTQ/7okGSnnCW/lIfS8BQpHyBH/VYeFl3Mh7AePAy1863olDWbU1bfB7Y
sKDTNhl4O4yAtEMt7KNwnALj11vQ4/HG2nlH+zNSXn/FI8lZUsBjWSfLyt7L7dcZGS8OYWlXBQWu
xcsJoaCp1tvk/v19b66M0YCqZ/5XbKzYw7+63y4cw0lDJ9OIKROa5mmoWeI50UaasXN5M3PTydbu
JX+E0S00LrTd91y9RkifOKn4o+JAEI9c/QMRJElI7DW84RA31EujNhYxD2Qo+AB1JND3IHBx9eZ/
VBtFfEXhbr0hV/l+9J3kD3AYMAhemyci+oTyuj+tvJJf4ux7qZbmeEVQ9bTlX/ltj9mZrKSHbmXV
gFZdT8daCDQWRTZkeKPjxYfbGnQCXosrLkRnmt+Ir1393ffJbvYM2gwRvN55ZHb8Hc1s0MDNw6Ld
VNrdDtwYo69p9hlbHM68nJGU/DY82IJQL5H4R4oVQXf37wJPL7oS7MS6ebE61MznMskNZvcguK7u
o/uWvAHBRjKY02qGqhd4xA+igT2Ib4zvACJmWFZSTKrlzaKG8217dkfQbz3kqoIFYybdfd9Bv9MZ
VxUCsBcFRu6e11zCv4nXUFFWuhvNDVcBZai1M42i462wRdqA97a9q6l1dr+RT8Xw/JRDPF+sF8xI
lsyGf/3lL4xOZcAvr+DFORYiBx2OxxeCluXNy+7DrBBToSk+NxW1KuLCqdT6CTNBBFXDTJq6o6m6
YEVGXWgNxIUUXzYPvm5A6qQW3+M2WASrtHHj6iSvN/qkVev9dcjDBKCDJDpcjg5eS8hZjmn3AT+D
XCStct8GokHT3IX3teXAtvIlJz2OlXxBV46863P/qlY3LKhhIjzvpow7uFlBb/Pbuq1hnaz0iTwm
sVnBcH0ubmpkl7VoJQT8pE2Cfxav8G7U9nzYVCXi3G2dkyk7Qq/8+Mfzsi0roJthwpSGOxLOubWe
QFC8CsUkbF5lHnzJGoKt/EJu4t613ea4OwysbkiMEya8hS+VrpC7018IVFtni9utVDFlB5UPN7te
V62irsHDyLy+e4CTjcRvt+8xl2BqTrmbGaIBlyiq0RzJsWGILxzRNCIVL5y2g7BOof3F1jiW2uXz
YSRqMxf9u4Mn+zY3qBkMvPnHSNPCRtxb7GF0Bjqnln/zRLyO/4XmMbiL2DXkqhhXA66wr9dL1fpK
iZ3CqiTEcH4FSKIPQnQpYS1z4+IxVsKB81CYy1csRqgSh5ojeUhiiQGDq0ZaClcbOLvT+aV9kAQf
TJs1TWnfK3dnUaQ2QpF3TycALmXzLTw99DKWM8vRCLYlCHP4BxeDilRC+Im/zX7XeafOf6lEy239
HDBrL6JJZoSGtxqtS9hSuqDWij2zkRejhO/W+NzdoNncGeocAQNuWvN0Q+Gu53REtP0Z8SCWrDSu
7nUt+2s6U16aLfP7yne6bofEa39XL0IoiZq+FwRPYim6Kp0vtDWCwssTQYbaxc3elK2G7sXgPaUt
bVpm/Jqn01g2FiIqV+2Jn2MS1Fl9X/zCtrxb4+be3EL0xP8QgGxVnCUqHMIfnPvLQlf03V1nW0Lz
0W3LAbK0B6Nqxc/zHl4hUj84I7hWf4D0DudJOx47pfVsSCYZknJt/16jq0QK8Gd6WWAJr9/LQ3Y1
QKioRbE8Ks7JcE4RxwA7+fHPZ5jB8DTd/Ie5uKRbFZ4B9UTg7TIr753qOGr+WbkHyHk4S44SHgMM
2BTbfsSHWXqzW68TU8JCVOkCDp1slb+WFd19FVUtvzUGUI4J7PgXOtwXDlGcDBFVQFme4KGRUMEE
mcyX4BKMmoNkN8xBdqFqC26vBGSdR120T3Va2/X3lhHK8cgayr5hNEMLEkB8F6lRHrtCuLEKJF2G
8YylS+4V4kqEw3j+bVoj+Up1An3TmEvzOd/sF3VO93bNRTKHFbHMkHQ/y/UpNQy8e2cSoKnihoge
fTA3ckXfic5c14lzbU+YPGCdxYUYj3PnCPGXqgCK/WT+ExlTvkiT4tIfJMES9gmTBUb1S8b/rJj7
7nTmTz46O5LeMBchkrkVXlgfo8g8LBsfm4uc4wy8GPdZrvVxEOuhXSAlwHH4KsnZ9MzoR+o8cIJk
QCOdDE33RDcLQPShasnCGdM6vBi8Bo7XubR2TbzqGsuFyy8OIXWtSe0Z4jgKr+4Nn4E0/xlVT8E4
ET0eS6L2VRsbAqDxBodvbI2l+mmN8SYsEX4J0Ys7o61U71bAoHMn6Q2EM+oaQfXY8x0MrNwg/9i+
vfxRZ9gelp01SyQeLsAuy0fL8nECaCAMlmDWkMd6lBgtT9G6rBTi8Lp01Vm5r7ZnYw5pQ90DuoZH
IXM8/hnGQDhq3nzeO2HuYjYPUiPYc/ck6Hb0ZjCBzL8InSeRcvxo8G4k9pYePU/clVKKCsEmOX7K
dqx6VDFDdELEqkyw0aJu5BufLo9JqK1jH2P0BlS8qGamJGPTTaNkPlML7mP2lB2/SXXBqhyL4Gro
uF+wTmzb+OunuVsfPeYBp2LEd9L6JDPWNIA4/Xmx1s/ACbcDyw1M3XVXEED+us/h55IPahQyaay6
O3eRpmIvi8kkEIJ+RIU/0cvpOq6z42ouzn5YsRRIVHvtEPhCLxmQ16D3SvgK8+TAH6Sk7SO3Y/Rm
PDqAvwjnlWwy2tCYqG2QebfktCYltijqKUsboZA3muc4hXjrQETLm8rBuZkorYTR1HlMApApCtR1
DkxwkBkycj/tqBxbOqpVBtJ94O9Jgk0z3xdm7dZlNqVGlK+u7ZDnt5h8V1yLPg05Rs9KuKDpMpk3
LaKIFlbmu2VK6CwltYXJHXo5xSNxd/v4grGnkn+rLsABkelavtSRuw0/iEUNCS+pokGMPMKB1qaE
sej5Dn6UTuO113qPvcE1Tbpetq9XLvzGCsmGpKkb0zIaQG1QoSq1rQTi4PBfdyOyBqU1AhzHldaO
8C42EXjhUEg/mT1ZhgoDFeRo+XtXHkr7dP3/MevCJKAFmdSrjqVq3yKsdFiLIqbSa7PBjmwQDMBB
65eLtcZWJ5igfDh60Xzhq1ts+0Xz0M74WZXOgh/nsKt2KTIFEhynOvQLIUX9oyzyUVy3oMqUxURo
YaTyU9hPchn8sASBapW0/H96tuYD3YFXcPaxW9jzdD5i8ghvDVYqrFTdMUcsb4rqYcletQX3t75G
is+dlubVJMGTnH0aqYYz4VeN6lOMTx79h6Q3FYMT0bb2CLzriALKvLsoUGtXOhRgYXERWvq5zli+
unMvqVhfQhqCsftnGDiQX27ZHGcC0iKPCW/Jds/z6NYuJF1cWNDyKinuild27VGp/965YSsXeUc4
SpBkpiP7d6WR0erbTRzrYrY0xtwe4HoC5IfYa0t8gwqXs/hezASCE8fmDSkrOXiNoB3Lb8KIN3Gn
UuTvi1oiC1plXuueAFVb8oCUgRB4qttZV4y/YDVoT5Z6hR3jGyglrrOciXyL25MqtYPCn64HtIv1
DyI1f4aHcUypVOmLwZTZO66vPKPre+/XIIijO+Hc3MPMjN8/7WVzABSMEc/ySfC1Ir1lBdqZqMlM
p+QTqXw53sd/p1zTlDlR5f98Pv7WGzNsnedktzuLBl5zcbsP5M6Z1YYFRhFetlPqcsd7qMK/UviC
480IeeifN6NOl+rUcEk2bGD4n3iJwJnfLBNnSNjx3cd3APAJJMtNYFzFTzFoNRJdBRP1s5XYTtNL
EOJSvCGV2jFbM7OkCPctV37NZ1I7pRqu291ZikK8ZxibdZLGjs7uteh+gtU+Ca4geccarASqrjPH
SYnfWxX6X0vSuosf3Q2lzEmsAj8mbmIKuvpYGHMVxaL/ZrqM3Wjrq6wn0YJEY2yRhTL+6XvBN1KJ
iQpzTjRnBjngYGBnRycBFOEBVLR/mHTP5xgZ3j6Hl2AL+JueoSx3C+hr04vw8C0Gt1lPDjpmd62Q
7w/j2bHUpRJZgWfTRll7dBu67iFH+UuArQ9ze97u/Doh3pEvIDH/YN/+gyTRfQyOKUTOhb0a7khN
XPIXTV8LFbDMJbGRPukuPTvlGHkUtAM1c09REIVbmlL5/W6ic2K1jK3bSdqIeZwV7E6w/ABdJ2wt
GIuGHrAm3l41/otqiy4OTAgvwqxeiIHdbyjTUc7y8P5SdHUG/kakEHTKdXyz05Efzfrersu5HpCj
imUC2JoYXV0Y8wRJZ79xtrSpXQtmT7F0B/zDSljSQpx5lQV7AVp2XWF4GJuGNKcfl6NhacEUz/lk
JMSXPDcsaV3uq9TLPlXDSNZm4oNGKrw7QMozuMzGsY3lODFp+hFLLFkleF51tkFmDb03nOwXry4D
aOfbSvZsTIIkcFN+gdiMlMy9YmM1Hv5ehBfwAtr6EFsUFdZl65NVLGdiD2bT//1SJo5EkFUSi+2f
SWqVpMRsbIUN2Td50a43yZ8gpSAabEyZVnlWdIV3M7t7pp4rn9n+tE5VDFkue91zE2E6S6CJ/sDy
j2IEORjB/FCa3hx0nQqx3+mZI72ByD56dyD7JD6PyAg5rQoGeyoz1BsgjOgZZFusH+iqebn2cszI
kO35t+SKzMZfw+woJeTDkn2doxlgOA/VJoxHYEjlDoNPhZUrDhqz4fktk1HBw/jxvO/RDCnrYtgs
OEGqREgXYzFkcL8FMYbTxiksFJsibVISi5wguMs3q7FZJ/E4IDic5YlxU050KFf+x0aisEb+9irP
RO4D6QKyS5NbdUaPOoVTgmBeVu6UHkdMzLM3i1rkb0U8W4Jsk+kpgt5ThkjB5ExfLTpIlNny//1k
4AuDxktHSkMbPKTqiddaQO7hb3pE3CChNiT1GouQ1RvK9GqrZkUSHZCFpqNxLsd3rjD1VTwbaQUJ
VxFgIQKW6LyZ4mgEccnR3bD+QsEMMPAp3spwhXUICwzXFgpw6usAHh3yoeG9j/zozxwj1DFQNfsN
Tr4Gvl7/GZ5ZoA1ofxg2vn8J95NRshGk8+iuH19enXvovfJrZyvw/Gg9Fqepm3jdtkMLIFfNWG1a
11fOYIL63SBNr0w0GXQvVAuB8EXD/9EnPre2doPWgizL6k3O1w0oLM4Bfe9PkVSXtLSDOaRm9rlW
wIVvNZNqn2DKeF2uCjzdRp7Ev+H0tlSbui0IZtzzHUnzplV+lAKW1rLMqyUXpNORc06cBigBShLH
NRqMdSNzQ7t72hZJcbyRqymk3VrUS2ytcncYqCGwz0LEAqyaKlcF6IPjEoyal/QRF1xXmXUNaAsZ
MSMr9uXXBYCJD22ecwzkIn1lFuQThNvzxkC6YNCVzvbKfM//3/5ZCmghdm7YLaqGmq7jexKAWdRM
+WJVhKLHBNGFW4OCZQwy2Pl0e8RJWz3uXcdno8mfPK+SP5+p/SfnGZEion0A8sbTnOdQYnXAz2Qs
VRZvF1jrQFKpLpQD7UqL2zXy6SZfJwAJtWF3VSKdAtzD5zF8npAPw4mtF4eiM1yh7vQhdGpPd5AE
jjxIWSQ/f7ejAwcdX1aoUzwuR+cpa+TWvJ8Rv+IiiWkYglPE2LjZ0sL3VWT7mkzDa9oneKugG6vG
Km4R5cE+6G57MLdudqnOjBjWR/Bnt5YhXI4esmay6/LyzBMIo/Gq1rqWhvPs76Yr5Vr4nqolQVYw
ZsYU4U2AV2hfh8T+Gbvb0dVLpjOBpHq5pEdnR4+x7VrSm+3IfH0+0B514MDSQJNloji6tA5tR8Fy
qRGFchzoSjQAAUWcinzGL+csUKfVJayKxqGraSVNVs/i29pNZlPk0GjGn+OEX3w/su4mJ4g3hdcT
fp7X47QMxbb8loPZ3uMzp+B+55bxCu1r8KVo0z/ExPgi2OtkeegeqYhsXl4FNL/psGX6ksugwR/t
9VAMyZ13ohdf5eAFSZSc90ZZ1dXM5ALSjbTpk/EfCn/kB1x9MkvgHyQgH2M6+lBS1tEYpuWsLWwu
TqlIv+HDF5MxevH8Fu4YoEQddZkIQ8W0iTRCn1BrBxHiTMcN/VqHoln1K7C04Qlks7UkCTnN42Db
edPyXTjroze18eQ/drFiqjyXJAou4leLJfw6DqycbT/fL7skQAVNedCWjRJtZ/zol/sLr0ZREAFr
OK5jLZvEZ8LiW16CSAfJGrLZhy/5bFVMccnMbmncTFxQ5MC7zrC2ncRrD3Iwqyfcw7CaGEIdI9rm
7d1pCprT+3R+66vlf2m9Y0/ytEMA5ipWT5yHBNqeh1i+t4qi/1/ShDah4JCEbREbzU7cRT+f/iID
8zLJaunBZgq0fghcMNrAct2i3QBBgSBSRmGEl+CyqtCG5CGKR9GKppoa0Q2baUs6geDReYm+KWCQ
hs+AiBsYNzRemnm7clXYmouFw7/3Jbo3ETuBB6dgcO+9SMOx+fmmgukC4SFfq2xuC0KlC/ErZ0Hr
ml+AX7d94n8BTA3Q/wzKDlaXa//QEyzcXz77sxUAwbISbaddx5OS2yVSG3i+ajtPifDsSiW4ipH9
MdEQhO3R2nWyMhU5K8zEGPyPaHmXB5fSl/fidHL27mgkO01OYE3tBUaJM1H80+tYsQJpkovrQhtK
JDn/KkufGfGyfatUQVBSzrI4zJTep/edlp0Kkpr4YBBtaXx63IUnm8J9/PAzTYjfxH/ZV4nofu3M
hJiUqJVNYLch4pJ4Pg4wwmd39I/FtELp1Uvc86ASfwGN2jVf9Sdw4GrN1Bk09YGkumxgHVzHLJDD
JcjFPdHhPf1BvIGXXg4WHPetU9Zeu23+DJ85PgARTx5jXe9pnWm+od18zVuetNHI0hOwJpyjcisW
KjolcsB//TNUv9hkExitlF8RaQhjm+tAmjc30/u4yWqy+izV/RJ8l3L39R0OEvtt+IQbdl/1O9FI
GtTxZuFwjQKDGRB1LRXvT8vZj7e8KOkODrPZlXJshJdAGSB2Rr0AU6MxNaRANFdJk7lsaJ9YQxz8
sz8yNzlywUr681eWyoMlDVkp+6tJUgDTWdubmcGjFR/JsUZkG6ETpBfsrMOwMO58Hum0ZP4NrzpZ
ZXYUx5vpRspA7t8Gim/eejqwVBZYza+0AqrVaiAVGlm9/lfpzmhzLTAAU3C4m/jCjxcJVp7us1nl
htIrDLuKG4jXuF4M65FKFGsjJNPqFvK1/bN/nQTueVzArf/+CSFfRnENkamj8eWmc6Mz0bEmjX62
ojHBMIS2w+11mOqaIFbT005YXGEAVgSp6jK9Sf0rF9HfzVxHqedbSzGWgRfQ1TuFxvu+BsduN5be
kJ7CjbXbbzXberkrww6XgdKKvyIkssupJqVp8bwlzfCSoayV4uhQwELrOaVDXoZnp4o4KykMDDwS
dBsl2y1p1Qpil+q6EPTaKEahQXdMKf/+PMB66DmmSxM5tmReqwuEP0e4Q4Hea1C/9bdYSbo1Uwto
/OiCn/a31bXL6RxBzf2CvqJKg76YjEKcu/ljLyndb9hitVTIn4N6dFCBLBsspbR5TthYIzNABwEE
pnWxSGjtSK5x46VI1cXTBOMrmCW7jbbb0942Vn46g00d6b6UixQTajJimddKYxtrLdURfQZPt5tS
2UcL7IavUUHkx0yvo9WTsu8EErCXqthAspJQHLuBJNzgz1l/tejNwJE677e2K7PaYg8IfFH1oCpE
MIvE6lnnjmSSgKwA0qbMSF13fYcfiKv7QGrKU90BQo+OUC7GPoQ05ywvi0AdNljmqXzklXizqkEx
WYQK0vZ8SxnSDQFpxNxAAupCjwJwnSHr0rIr68G7Ats+IXZzfEf/JMtWG+O25YKdqX3M8WMs8qqG
Mq9+wBkb6RzMgKSUzmKJaxZs6KUBiaI385cc3N7Owenv0pl9YJZtdprHwFHGLeQb0K3Px+6Xuovw
G+c2sOp6ih7LlJD8cMOVV9c7Lgwj3n4MVbLx66Hpzd7la8s7d4HmJORR6a3J+J6HJF3q+n+nspg6
DLdp9cTY92Z9TvAFK/5wkQu6xPdA3S3LOG1fuH76g9YO8X8XXQf+gxwhsPdPdCWx23FTj7fTwNi+
xsuLijVyH7EuSTAlQBHEjY20pl3t02N7L378eMBk9/RUxKjTv0bYNB371r/jFRWo+YfdAoCWa8iI
LJADAwA6B5lKorbp24Vu+v33Yg70hzg80JI9nVHg7vwQAj3+KqN7SzOe4Yo4nmDsVMzE37yW7KdR
fx6wBsyG0qeiuyV4FbeJj63jHoQEyNZsmfBu/zxVdY2JS4mHkGVC7WLUxroZeHH4qbeqzWcEgkPu
GVT3AGOruShaoGIi5pvDhmHZa6QSM87vdu6jeqWPUQt/c4idLhDLVHLv/Q4y/pvCh0u8mb7q0jpp
1NYxRnjhpRMg48qn5A16vQHwPTQwkPUmKfO+xGxBIoaJlRPd11pMtBwCvGaoMrKZHwLBgfgGLppd
a09wOZzpWmD6NpcGYkFqQ3kQXc0e2SjU7VRJC7XhIkvZm8YWgJd5gps08OjiEyVbLzo18NowwG4E
H/cECS1iMaaLUd2EW7Q2tTQqiocfQ1x5v45JpPUMqT5CLhbIx/G8uI/2PXemjSr+pia1Vv3LZWCU
6SpF6x8MReFK1RZY9dSLt4/ZsT/1DE5s0nsxL7etdpAg0ZmUkB84GSw+Iq/9H7mYJgFY6WQMkgmj
dCHJh9TP7jitsiraY8TZfogYGt9JYDCdjls0M18wcPVshxlOdwxPWTHV4JGdSoMqp1STHGHCe+bg
2bHdAY7iwfl+8qaWcC3iYXC7HkZYlD9Mq1rE+ZEGjPNKzHMSeVq1eGtcQZ0ovJDEO2QorgiBGs0L
vIZ7uFARkwTdpxpD5UnsTXaJn/due54cNYY8WRspOkFYKk9+Orurx6arNUNICb9G/U4DHHcUmz8j
uG2NgwNq6GZqHaTIR04cfugrk1MeEKNkr/o6E0tovqxW6DInpMrIqohEHCbc4xdhDFdY+34xgPsV
AgXfbZkEH6DyNE9KSqjf5DChyAPtjudAARp0KfqaD8ZpKWhYuRYJO3mL7cNcaJ2xiCQh4GOxlJAT
Pcuz/piLVD7UpvH98GLp0pJGNIEwzz1w78UXl859TQSlBe+OBbVURgl7pld4q09qoWCMfFonW6ou
IXfRA0KSuA+XaYOQR5kzOuTTHb+CMRlrUhqfDccLLiBXwGpScUj3L86UOJEwSq2DrQeBLAr5sSs7
+5g28X6w88uh7ElkTrODQZKZTjPuP4AvVkui/6FgIgCFzGNTuueq3kceEWk7vNesjR937RY4flLa
bS2pn8CXG/QdO9hQ6PKiM9J7eolxQ9K74eYsYi9MFcmPsLoZV15AuGaqNSnSw9uKitE8DvMFSDnK
+Tg8hFef+iDC/qGa2OksnXpv+KZKaSi397WvcWdmiHcztJJzLIPKLgCJQSFN5fYgOQg4UBmibxlm
DkX5B7xyYEApVxhif+CzlEObhWoeYR9zWYwyGEs+fTaW5BjVgY9v6V8dMi2zNmMi2zCcNqWluTYg
jHFiLqLwAawEuGpajMzUeN+ANZSBNcC6tZmVJZ2caljU18F3/O4RcsVxJrTwZP6mA0y1K8eMrXNw
DvNkZP/4ALPKoJo34usWrsCP1qPSP+d2/j0Au9/knPapb8mYcH33putPHYP9uM8qo2fKNQOlFzBa
cPFJCPylD+UArzuUT0lcb0n3VGnxkTngUIEJmXn3fBxJ3z208p6Yr+xn/XKfBaCcjUk0TXRxBe09
2QO61wuq5C+e723g1lAtGm1XlcNUKEGlCMa6XtFnzbillx6eocTozMXCTqj666Uhp0BWDs1nQAX1
KjUDGmDj9IRcOSCbz6nCDAjf9pDxpyIK2PdIeCNltXOUEAfEa4WM157rJks8a/R0O8ERBiCQ0Nn6
CCo/dt58imnFGL0YVY1lOX8QAqzJ4Utill5EBwNC7ap0zwvJh8YAQz2kyzxQyhK56sF6HSQgYjkr
yn5I57TGC4ADz4C9Qxcq67ts4mnIIUF8KdOjVGUpm1CHISAUVSpsIO/4bHGtymERaha93eWYaqUm
czFkZSVgaZOzC09ikpmlhCXzViAms4896z0CLXdL3PHg59ODVqMXNELFLVAnNBM6r4nKogwtIbIo
QwAr19eJVo31o6eF0nMQ3alWBb+ABlA8S/hnlJYbg0g1bdq940hmuH/sipkhqEcUbZd2EgoQpv3J
oHozvICga9XM9mpEwK+TLFBro2AmWD/mcOtrhjovW91evciaVKSQrIl3VDNRanUGqQhnzX4gpFVh
fpDyYmVndZ7OeBZeQT46+GUEXXz0Lf0uagOcnQN8PbW0+dMZPv+2th4PcEMaY7cOQUTochcp1WQR
Yyva2IMDtOebfetQ67XYEr16Y4Ik1KawfQtLWhkDauqTLidUW1MHbD4CWrASOIfJA9tSCVXVOWyl
4xzbKkxzBZdnrrjeI7tohcO+7tNk0+PMzfcfTmR2BKZAMfM0zZjsCVKzYdcPgZR99IBsgg0J4S6P
c8ndUm1VO5+18bM6GmLESqK/UmcmDdZtO4AFmeceUUYERxuD3SjHtEFRDlOk+AkM0xiMXdC8Ilrm
VKyCLUKBBUV8vWqv6NeTiumhz/4TBZqjZQw+S9cLnH5LbJ+uxcob/mcSoQ/3kWkPailIy8VxCQiI
5bLwzDtzeoD4LLEOVwzZDWeLTS78yqfOx4OFb7ArR3EhTqKYAg8J7MVDqsfRoyUPTgEEgG7eM6cY
z84FD8l2k1rVHQIWtMZWHskAO9tlZ3LHW8JYJeVwpRC8kcvK4kdGt059E7B1j1RsYCYOof0eV2xZ
LEFj3TipXF9oPQwjA1+RMlnxnaDDpbrW0CWcy3lPOKPuYb45pX6/Su7PZ+QuVkLCOq9CfjSzOWqu
RuWod8E/x4vbK++hmDuWuYitAk3t5DNkC9mmfKZMhUYAebIQ/UYe4SXmIme3yKLQlncC9jjSd8KA
zMVXahUdkBynqXsQHyM7wVn5YXbpvCpleElS0QZB2MqN8cIfeiwFIMiCuHspInn79kSqcU/Vj6rq
y4U0hEgPJv6WFg8gKPsGjQ5TBYmATFvuhjbGNIq/Wr//kITj0+eDD6F0z3kq3/uxRma0YaoDxrqx
PHOaNkbC08ClWQ/uI1cMaIcJOJ5iacHD2EzCkTOeYdBb9cOhjLurc3bECl3XkJIHc5Wn6tLmI7Eb
KZU6edJ31P1ogoqcX4NYS2zv/TnCrQ+soi6spZOt7vDC3aCIDMSXCC5RqwYFqGAh1KanYCRH/Byt
ohopD3U7OWTQ5K5bCy/1YhhqjafydTWCcOTLOj29tSjvER7fqvGxE2TD3YMxLynDvUOGfbMOfGPb
isI3m19tpa76Eux4ZRxkPr3At09tHGhXeOumIEt/ZOum5IXQ9HZJIS1X/EnzJsPTIohJ5JYtG8pn
4b5zpaEoQ2CRh1f+Hxkz3cKNugEaPQV+Cd3FElxxV45Gu+HWff4jJQyC3JyUnpgOpwVwe7hqKu57
ozRNTJ47I9DF3QMLJZ04hWX4+aY3EhP5bDRb9JYwof2efl36IpB8/FZxel41dzil0c3tbbKe0X/0
boL77fn/oRdf6LcWyjgr7ZYKN2PKvatfnbZ80DZI9Gv4eKDkUZHTElJsx/IcX5NyW60Woe/5twsl
PrUDQx/ppAB5oRJzoG7M5g2N68QZxo5CBNu+FHkfAlo21Yuq2hT/Sdn7RLj2VoPoA/nppLob8V9X
Vw6W7MCZgIsWfbd5Ee8b+QydMIDYvW9J7ehFvSTn5cQiqgVl1tHCq8IWwvaF63bPgQvi4mGVNiVO
gZwe4CXx9tFS/vzlGPML1Jkq8T11Bldxli8xSZAXrCB4Yo7o/3uzmhujhmB+d9NEs3P2r03cacNH
H7UxTPvQPdHpygQKKLIEbIPwO80VQH0EKHgri5VfAAwNJaBcAvViDNpxOmOGpw/nbFA0MkTIwy3V
or9p5TCMQ5Nw0fp8qpk7u9+X4XSyBVNHqWsuc8yE49ytLP0bOwNHZokrXAx6pDPlWSuSwNArSBtT
8VShcOQoKy4qmT+v1lnQS852vJGcgP+qGYqatkKCfJdM3CFI4WM1gP+q6GGlzamoZcvD5+sGZy6x
hJT/v/GNpMDdI3CwKLrcr7JkguWbLCg0xuNUx7HuzMRtRfnHuq/wH14I7S4B9Y05gm/zZSBdryf2
UOwR62s6zAoLg25c7StlV44GZ7+/O46TDdnR2oEUxrMyKVXlGblI32p0jD7/CFKVXkK2W+wdNSPF
FxnSEl4tYUs9o8YdW9WNTPe6BYHBN4m7rbTRVVeKrPYhmvWkz4ssh8P+OS8noaBZ4WLm/w1pcL9M
eH5dALhTYKH9oefGaV0U9V4MeiDnm9ypAmR0uNLuTW6h9kCgkIelbb3Y6lK4WpWjy8YbzuhJfNnf
uxTLwHvr4IYxQ3SSIFb5NDGs/d/2qfzQUN1FKrcj3OFCVmZIwR/hwaiU3po/GXZR7GXYUfRrt5Rz
NIRqJzNu3/0qzNTcz72GfX7Qq5AFslQJD57Fvj8NCXAGA9GjA5fG85ilogURGEb6dCYkaw6niNl6
kAHYAokg067R5BksqgEzjFTKZKT3SnlPctEHUcyAoQLNTxTYFfuOvE2dXkIJhfSr0d01u0uFMpmN
hw2etEVyZrsoS9qG4XL479riPl77PQHB2OVKn4trPceYjRgwJJR3DwFXMVM6mfn7GPN3zxJAAxpp
gn21UEJxqMzVrvZdFkY88UCsRhNtCVZgjrpckIAhWMkky/rhDS0J2dCKQotM5PxCXubrhH1n9BQK
eOGAvGpIvbiwpXmRIzM02wosnoqPL6t/ldWJ3gI3fICzCGvj9wMG+xh+vm05i28s/SegopCPbVf5
vXKF/RHUjVT0Wkl2xpjg6Z2be6IUwRgOg2gciaix9wZXckZyRIoyuznzl4+zrIXe/jgCHNZGTsL5
q9hOOrSfAZaygeXYpRb7eDM26ze8nb1wE6ZEuyKI6RSuuYSTl/R/XGKyEx63eDSmiLoNv5P6Mn23
7RBCakN6njnRSKmQqjI74yIKHbuP3h7JNdk22x6aptrQP027j2wlrJrIEklBk7qnEhf0KPOpbrig
xkdhtXbrjzJKXJPt4jZe3Duyq5oDMmWvbV9orFSOhhLrL0EGVZ1xMqy4kXMKuo2Mp1mjXH7cV61P
wPudxR/6ZpFqAiSlBOjMJDtEc3zgkHCSB19sYD7fUMpwh+LXkrugzjpTq40a8gIhxm2pBOh213z9
cEoGRAVjSocl+r5GBttOs02IJYfd1yEeyXIk0Bsdq3dScxHH5lyTpWPp5CpkO1CFnukGPMvinQ23
gSNqJwpKjEn5PBswZkXlyzsh4erb+ogkn4nT4VdPvjztQw6g5HhRwB89WNKILYe93+gh4ocX/7zZ
1lJV1uJU7wUBpgDrP8cGNMP4DNnh5t0p1325R/IHJ/xzUa+tBqhCTpXxA7NJoBkvWkj+Zf54r1bY
c4gedcZ5NjTK4Y8qLwvT1sPopLLdUiPwlPI1AZP/veGaImfoGq2zWTg9biUMO+X5Re9bVAGRqnlT
8v0uY540bqTu2rJUFI7NWkct50HappEVN4YacV3dXr/qvEhCmADT+q4HMvV4De5AHiol0l6HbsyR
x4JpN+igy2eZglVeWqA6D2w6n27nTQKo4dZZsYFjFySrjxRf8Vg2GKeZyQfRxdn375uOXe/t3xAN
Z4EuU8LinUZ4mxE0uC1HxiNyegjEyGQ0CJiyU6N9vcRmYT6JQWIOqLfg20fcLJDdpw8/v1Ubpsc2
71ZbxbR1Z62apGuWo8VezYTsOpBQlUnNJHGsw3aujKVuSIpXpPE9cq4a1Twxn8xXyKT4y7ucrKVm
hpE9zVqNIJiEmBOZcDcwvmd/jvXjbOV240MZFSV81CP394j1Csv/AjwWKNilwx+SgVaj5ORR+STM
YRhiaYHemkazNSncAMyA2rkvXlih9kgyfgLkUXK/y/naPFyACXgx70fkb8EgZ27ZmYg1lLTowQVu
SzjK/9GIP7M2o5mx5Fywnlh1N4dzdSeT43hyYmRtOv3znqkctzr78a9b4gtXI0J2m5yrJor5A1zG
xH3PH2IfXJvtRQZTLNuLNZjQrR2pwENd9qpLw/PQl5FIYPq6UqkjvqZra99L4OMr0gdyMX1vbZHY
0UvZxgZBoLUPfUrx5Skvhvl1SgwJxCxXvfEZRWWpOwjjsWMLf2EYbEFXOhhXZFAmJGKwL97HByzz
CQihhuHKq2IlctglchhwfJTzNw0AP5lIqS6VvxG5e1Eymqg7bgu3eU6gvUym0nfs3tvElq6iFTtz
Ly/BHHmhQUpq0Fj2k/KEnSQ9EO5wmr4BPgRAT4z/mB6xlpkpB1wZ84eLt7BHF5gy8XpgeIWKwjEF
idWo8WlUNLn0FkEHeqWA7ueDYZpibeNC7NonVRk86rg5FYGUOf347T43xbN4BNn74A2PzR0pwIXP
TeoL8UTMu6o07tHUt42VlTfXDtHwHNHgGK6RN6dbtrmzpX3lW7iIxJOfTSYLlsLK9r410oVqhMM5
PWqahsG14uzSYhs2oKKmGbRiY4AG4sMu25RdquymmWLQv5ql1qqZQkibjsJjvoOwsViWdZZ672lv
sHGHNpgQjzu4k9N+6wA1Rx+4UTH+nRB4F7JO0wQh/OcYeTYW9ENdJkw0bhmban/GseBTMJE1kKlH
1VtNayNT2TDAM7fWGymcqUVPNw3Z5VjFgsSDaaZ7kuvsB9EwVSYK0XE0UMQVBWfGLl2K93MoTinC
4sKsUtSpw3SeilTAGv6y586TIA/QMuSRxqnzlmtx0cZQa0YxMPIqQ6Ud3c+9Pe1YAM7pmtouQjPX
oP0hFFOjaAxr1/fHVqp0ooLP5oDA//Fh3KjD3e3ohHYupqD0EERw/KiNlSk2s3xzTzqZGXDZ9Nb0
rEyxSDLQMoEdO6OdLXxpzGyIFkWxjPPIl5xeRJCAIiA2hxDo6fvV3RrIRrj+zszY/ufiZ7th3gqf
EoIKcjI4jgJoIk6/9wi63KR1bMNiH5dgQYMQsy7eHOxC1qKG2zYjzFSmp5kYVqBv9U5C/xTRPIaE
lgoY9OW0fyL4/GQDg9Qy1OzB1pYMz8FJ5Dst/qiJCFFIunlesw3krf/MJ9nSzh7KrhiEU3YlnZtW
EP0H9KZg7W9D89jS/2cOVP7/NwQbSSj1U/Y/9mO1bHzghHt2RcCdHPlfNwDEaCXa04k+/Hd3pVJO
wRIOIBV/aByJ7RlcOuquwxJQLlVUBJ0hiyOMoIXhg/i/WyzxJDTm4PUfWHeUba8oTqDsLUkAkPJU
dUvUqQiZihekwFCAa4HehKKKa7I+CQcxD4/LLAdp9zIxu3tgrIQgWbYIBD0Q16gARCO+MUCH4Jun
mfSc8JrfOROpXu0IKYMiNV9yW5YLXlhmzDI3JDjlER/FSBoA1OUq2o1l/pOEuRrwgGOVSh4Hfla/
4v9MZ6Lva3d3h7Y/pNdPa2xj62dxe9WSZbnXvaJj6GZJx4oXe7zepA9QdTCTG3bEAhlUxDP6CWnk
V+tzu469S4AnLAcDCA2MVINH4gyyEg9+rIIWA/u94EdWSOCrSOz6d1zanXuLG2sKGoOG1uaMuJ17
s0dh6w8BViQgHPFDbx8QrVFoOTnQkrVbAXHrhH5ORBW4TumcijY+Gi06FShhKCi8s4AKOSSVtRRO
vBMtl94aQ5ST+cOEWB5MZlV2cIDDaOjgxRU2nke47l2vg2swrWvAmnLhaiN1p9DkeLZFOViw5Jxi
cFF1Cnb+Q+7C+cAVEHgz0ko8yYDNyRAFrnOg5553N2BKokn8lwFaiTvPG+apg67ouMxc8Op/MNP+
vRFs/bgmOTfqOaJU3rFBWhha7uHgT+9J6cFVm+SiM8MjxW/qpKOTpQ5iSqEjDX22hMQCHzMp8pOI
Sf5DLcUn4ab1qP/0TuuJH7gL9n2qZRCKeG6gmLJzaklnAQlm1USv6nLo+01ywAKqvA6HYlfxcd4r
lZYM3EmJKqA97EHETssFh2/Sp/HhQ9Lfp7t72ECR8b6g0MM8itvTzu7E13iSe/JYKGAwpwt/xk78
gUdXWQmeneXBDptq7LocdT424XYDfs1KyPzBjdgrArGco+ijFfaHpBB7hoExLSMRueAW//d/Mzwx
xM64qJOm3cKQoO/cZr73s2Kl9f7nln0r2WWdDwcBpq95GiOCZSaYlBH2KsZ0uDr6JN/c5j7K6qRb
mInekEUAoNX9/zjn8QoWejkbl7eChXFxLfbXj0tbMVOb1yEH7e8HimUrN/fEGZtEDmEz/dAtei5d
D0ftStMYTvuOXd9Eh8lDpr1z5tQUYrPwCHDu/kLLeM1FViEvIZVw2AgS9B+n8z3A/YJRuWkhj6Ka
nIQAE3RoOQlviQgd/aXywXJas0lGBt4bdVmTuPN+qnBL2KA4Pa5WFxMpBIvIzNV8gQCAz5AbIOQX
wGRuVqefgyklb7TsFOkExcZYTU5+loaKXqWsnj79WmApXx6zeb7EhULqC+5f+w00X+rjUhk+z/pY
SoJrBaw2xJlU5G/d6bWqSn26l4JI21iCMIk+mv7ORyZ1z12n+GYq2vNdlGCiMah9CwaQzT5HkuWP
y8dSnAnSOgSyi0JekOlXviwRbfHqm6c7NQy954tRJBrlag1Dm/wX0drxi92WFfLmPuM7dg4FfNRe
LOcvczlIBAjbzMbsqLGATeLqNwTMHiFlCBom95WIMyFE4bQyOyxtFpqLrs7utg+6kXmAwxcZQdRd
Lwt3JcYMXHqG3yssMk78OzVfa05PUF+6lCsqYBctiEzGiduTIuIXWJOFrboVn8ZKqLZuIC94gIN4
tHeC5KbteWg1EXe7mbVFoBHHBf064CsccGhHiMFTFNASVrn4ENiWv+SSNRghwVAaKIieOhqxaDVX
QZ4hIRNIHtOqLAAgiinpUtWvoCta7i/q/+zTHcd9k8/0D6zZv4ckj5wV6qUKCi0jVaQndQs5WbWv
i04s6wGcbVhMPET12KN8jowel26u8tTT/rQD8PbKnrmhEo6HNV7ydCOgIrXFrs09PcpE4zsJlBdY
X4VQu82OPe/Syb82+WtYAbjzYgcP4uYfGK3iUbIaihuXiZzBMR2rNATvGvcFn/eJWa131Wx9s9yn
En+t9262e4GKGCEa3hdz0b7HRaGbNp5Us5koAV2Iu8uIpWDk2DBWd8DMTnQ8JtciHNIRqoFewTpD
7FPbYAq2W7/jTx7+Cn+AQACcuT/1u4IZX+R3n+n98NnMvBfHmcTiGl8FuOEciPVhpyZzCYwRf0EK
Q9o5w76OdKnudIZztGzOxYAjFa5VzYTkE6uZhkVWqAAVSGbhR8THEaMNugKWGa0i8oVheVTDi1oO
MTzND0Hq084f35IoCh6MHaN5KOchsDrpUs9UfxS/iPAvKj35oX9S8m7+wV5J+6EOqlFlA7BKxnlk
CYHdnMOJgeDN5JdxbHl97V8a/fbNvumJWRTMFuncihNqNZX5nhCWnox1mrMYNSqaqUqHmw7iKbHO
cpa850p9KYq/RBhE0bJyvTtKkphIty3dNTnA9P47IOIBaTAmHM9Q3U+fbp0+PmSm/Byp3chpwLHO
6IKUEDnI6I7ujXEiVM0tNL3hoN20NXOZdenVR0GFyHhVlwTzcc7zZwDfGLARqvSjuakcmuw/IlxK
knKpNaLP5nCikzy+gsEr23l0venT2o4Ue4gmvpPINljcppw6F8jeE/3gBDNJWEEag3vaBJZi2PmE
HTIQQmv73Tl9xvLYx8bqwOUo6V8E/trr4WFrVDqVeMpyn9snT9EYynnc+BIlYWOld6Xt8n2kiYi4
RPb5dImxdLjYk1R6LzUlQARIsHBXJ2J2+TfaknjEo21zFnw1KSt9tQU71lT0RbStwQ/Mg8nDXMRN
DGKRUfvM3NRxGOx9VB4fCnNLQinf2a/SV+NGxqvAmCXtF1G9nz802ZT0wUI9p1i9/xbcV7tKrzkd
TcMHv+hHzzpM5XW0uTmUx4pC7zr8VsYXfYkyazEaRAON/Bt36bKP0j9JTfPfsrp6uMk4cjZF+Ay4
ekGtHqvBzQsKxNdjp7zDml3zqa+cip0LOKDQQNqqNAKuNyQWAfi6s5HI9JeBXDaA8eyKV5DKcQTt
Cj4m+DmF5kXzNiyBYhcfxiRdnxX0O7GAKVUmyHsWcIFW3DnQSdS88Irc3CInKpmX6WKDLMrE6CsK
tURHRiH5Jsrt4sQJrBUV/TywgTfeclixQfbIBR953IOgncNn0dqK/QSf1Vhb7BALsIFFwZQx9F9m
N6bidFZOdKxA2NvmwAQnefCST9fakWcGFxgtQT0a00tZ7Yh7FyT5DcGTVOe96EvVOfFhHBo5Lt3K
zAseyuBAUwhINBPu2foQd4hnClZM5fWOfhwiCOcN4UtsEaKhuYzyMaM0hhO/QecyXuySsScQcvpy
11PQPx8v2ZTMDeG7yI0lXEsaowAKNR6gdZH5/vZRf2gba+sEY7O3VIZ2PJKOPfxf3hcxvW+1btY7
V9M7ORhrpocuyoru21ii7VTE2kjxONuyeKvJruf3KWVsDocQuzhUzb2wo/1ZtdQAtwtmaGWOC+ld
OIKIZAAUrwzUOYIXNMACnwuiuGkI9QblNxijRhRmY2lPv6XT8MjN1FhcIMkiDsfKUGmCpMgbn6ke
RSfRQ4JD9liPOmTi+JAw9MW573AOEWPUlAJE91K5KgswZG+UixMZeALEVlCCtI8IQDwHjm1BIZ+o
MZnAAApmoLmMhSJdpxNzgPeFo0dMnwEwAls9tl5gNg229Hn/BPtG61/Xnp9+RlRQmFiAN/1z1p90
chdtWxky1LN14M4Os4v7m51vEmwEe7nIcOSNdtzQsAz340A6x8D+Ot5tswGnzo8ralF/DYKJM9mj
ovfYS/7CHojPBzMDQuwl14mJLuzSYpnyKiwH8qvW0htak8l8I7dvwp/46n1Lq8vbA2y9jDhp3rz/
6yNrQ23pOGGGH5C6ucfJn1p+PhYeg7vnZZiuLrXXVzSfHd6nQXHVNH2kGb0k8RUQnrawgbZxBKdD
COOT4ENPcTNbh+Oebm1JvxJCH48Kv66BNAkgjplCDCzwH18pG2l55LI9NP3mChBNZQyKwYRMfjRI
iApcyGkfoAVG28CsLcaCC85qBi2Nf+MTSddnam2YNAutEnoUqzr5SXZKfDR9RIcFg2ePYJKjMnDT
OwEuDmot9VBCiea8s+3Pq4rQ0q6apqJfcfpH9yo4HMJTnHBiSy39vEdERU2SlZajoxLzdHlIDHri
aB2Djkovqfd7r5v4sjgmOdkQgArCKkLByTuNWmgxwJmKQBf+MFzxrv6YbwDfgsLyxY1GDRQ74Qy+
1cIM0KkrceRZWNq/twQxR1fm5Km0L/ksdAgE4G/ZI3p+7bTAnfxxvDEOd6aDgoS9qOmDEk8C4mhe
gw6cjnafWV3CyKH/fksxo7uDzZGucvyKTk3oo+nN8M5vXnZkByT/5BOEvsBcxXDtnSjRzhma24v8
5CiKzZElAeQnFCrIJkdQcHdrhmaa0Zab0rUghdIGPTMPpyZxSA+o0ilq6Dl3wVDmMl3f5l+RM3rD
1wf730S9AOlkqrOhLrI2+Pwgzq7wXbAKog5TEQDRMwYytcxtux8FTMr7lsMgPLCr+aC6Hh6Du+dM
uk+H6ffJGEkqXFEEtekisJoLXUxvCT5dZseOWzC0oipb+IKkw9qQc9tNWTgVH4F6/ckwA3dHdybX
/wkqd6Xf9jJhz0vnMVovKrmqhAQN5s0ixxLm2e+5nsTdQil6XL8+cLEuncWJvQOweXqeuC/eRne0
kJHeHoZrU2+ekWSmfT+nbkPCk7bAdCvLWqG8Xnknp7qP1ZL0lG69Bz7OcOslNmOf7dYffTHOjnTC
dJMND9+PhVcA4+SA1THRHg99zo7HL/FY6jdZoCpnPQiTg8nacmOwd/GiawBPpc/p9N3DacyLg/Ya
7D2L3Zb3N9ZP+jf8FtbzYciG0JApvgDvmhcuQrCSO0lO5tW6FT3oSyWyzzdqpth8vOhnpo6O1/ZF
t0n24IiP4RJcy3XAiWl4K9rR6Xa5HIDaKaL44J5G7OGUPYcHKCwg2+8O1khjNgAt5Hk8fqu33FgG
GAV2M0ubzPkLF8zVM2k7LaVy9p761e9FDdUKBlC0X9yOtt9TKIAl4WsaoOwu/k1jGiNJhf/mVV0r
pmgZ9MuS/JKlAOFLbiB8tb9eA4WIa/RXpq1bENSrSxvNlrhnU8WTzo26ogCH7w4FT7kW+Pg2WJcm
EbUWSI5RX5UVlB8V3X2wk/3q7E7zaJcIvcAwXhZQKy2YSUxRj/yC0U4pZiiAp8/XKXtihPhbyrGm
JbdNmvlF3ieFqvffaopScYnA5/NTnC3OCjInqZEI62hVCQB+zZMiJA24ALnX6o6nA4VAMKp8+RGC
ptm9TJcQnZzAB/lHpbVvDcTxU2ns8WvQD4wdBRuS5y7o4r9jWtepiYPvuHw2D9BFiEFFfiKFe3oX
+EnQqo9XrU5IN60qcxrMyx9a/zQrfmbLqKiFhk9/wO00ctag2/cDbfCFJfRQfzwhP7M2u5mKC/Di
SShq2jfgYKrd/OqgiEfUPicVF9HWvx/7NtZcwIdit3fAoDNLJyCQFKCkSC245fIJiAAcjHzwA2vi
Pwf3lNu1FlsUCKS5gdTSbss2T497EdFCQXoXei7ek/fFtuKQSIA3gw/+AGoI3WBXbH+3bk185aIX
j8YeE9UE53kIms0hIEfo/0kdMhqT4ztYOeWr9X3MqIv3K3Uub3kPQgrEX98W3MUdGuWzZqXCA97v
fGHwBW4hGUiK9a7swfphA/aHD7Ir/nn8drT0Ji9pgBCCnd+4COX3ZdNU4abfWuzaj5TVVkBIy/DU
XelqubIoBCyWebtP3YGszPWpUnEPVdVNJn7ycrBBWY3KlBjb0H5Qaxq6IghMZmJ6IUY3UNS1e46/
VQzffoYlGEB0v49Nbu52E4BmyH5pcgPEBM7D+DH/ea7mUv7VNyo7Ax3gRFvF/RxamLV/E8CPrldq
SYSRHJeA5j6jlGTkPGiqXHJWSTLmUjkBmnKddblTa3/Ep8APIFJoVZPRKryaT1fdkBorMiq8wREq
nkqsmfeqpqepj0r4kXbc6yKPE5gvTbuuFZD2NyanIJYJ116dNAlXA/o3yoO/MCc1hujrTGs5FrU2
NHPW0KdlnmXAXzmMWowiIk4keOsE+9GH/PS11Nxf8UtEubQ/gv1C1gFpmVvMcLAR2sSWym9/tLNf
CPYteYLoqSTZWd/Ow3uwr26T5OeVegb9lK1crDCIBERjI9jCbE/pvF8Wz/inE/RDNAcd4g/z5YGk
1izvScVYAbtruezyQbeML+xgy0j2mkzJNq/8kArdlA6hx/TURC3jnk54AYjY2m3n6vFhOoFNnT+X
PbUl51JUWJrqon60fZyLPqmNIFH2iavRlC9actp4rMu8i2ZLL2WK1dz6OhyzaCS+asAX2+reFlNH
jKLa5Tf4WLP6W/JqTsbStAX6qCz0raoi1uC12C4KPiQSWTfAsojv+Twk1rUYt/6/DURk6S0DSZMB
NQRU1ZMuqb/S7UGehs96LnQ3F6izoCsbm99I5mey5lBpypq2itu1V7rbtgkyl9VsHjyHL6/91KUj
jHtI2+YQu58hUAnYKQJrUU8JeU35yr8IcfX7mXm+CyVBEL5M/C2uTLpPBLrry2cCOL+S6KR8MmlP
/FViFi/ILfCef1moJm8p6Ta7cl31XOBWAc+rh51TI5d5JQhOTSsKdwdwGbQgh6n6Mlf8YmBPM5Do
UG0ZQchGI+qpbh7b8xIX9Tq2LBlhKQoZ/qmeik16YtnICcpFxXnwmRdUR4KS0DcOb006WqEiiHs+
0GfbOWrBnIWndIxaKBmucZgQ4iQfntjB+sz+tkhKBNCnPXZ142eQEPIE8myMoOlWraPm2dapDh7f
alLPR1hbVoCdYtPddw5azjVo96BmB7st0bzxV2YSWSKq8U93jki29Yi4mhLvEJC13/GmhazB4y3B
+XH1SXCOHGMgb0L2Cdf56PpclGz/d0d72ewHB0v9caqZeb0Wh6bKdyyvlA0xKUbdzZA4tuE2O843
4sI3qUzXaE2OEKCHPwtDsNY4gTBwVEz0/lXlue/IjcXELKqTUl9CpHLK2PuANSotaZhAYN8hPk7+
m411m/oFhd/fQbAVXGo5ohBzS+l6w1R4ebts5+OCJU03R9FQlBh4jxh5xa/sBIcLfTLaKPmQ3nkr
6GFMXd7bHGFHejxKUwyZEY3R8zLntXDMMMjfIElHIDJVag4fMiXjre7nfIZ5belnGd7OK2YCci66
Xf7MqOt4kXFYbGkjioluu3XTkjhlBbkXYmic2WucH/KvQE76JTd5+nJ09kd9wc+SY9n9yM3QbpFf
OwK5bZKMq3NqL3uTE3Tnku5KM9l+IndTv4RV9Qgcn26V2oITslnKu4Zjg++e8qC/m80hnlcs1CX2
TCWolJlLd8D19zuiFYKB1WcApdQmzDYs2wxVM6XLfCnCLyX4lrBVo4WuTf/4RCxB2LrvoLUN6RAi
XJn7t9/oMFveN0xX1YOw/XTqPdIHm22ehMsz3glmwSmOMa49IOMfYxzd9RbUfQ4FDtidkYd6whon
kur+hjyTEQkJO9ZaJBLI9704p2bemAx5glBeXJIckSmyFWFyq1f3eIf2j5jG4Yx8czsffIS7dTB2
1LFJjPOHgUw90pds/4JksSEHshG2kip5QFmwUKfHmPnwVtoJ0IYY9rjuCnA/wxUm1g9aPskx19VP
sQDuliIctzGwtXi4hfRjrl+6XSGNDhobfcCF6SxaFx885KnxD3aQlkRDzi+BTu3l2vK3PLbocL6F
Qz/wPGWO6g+/0jWVkMDPJzdxnM7LFfC3gFBw/bcr6fKqauGyHPHc56LKchAkYBoD52fQ5ORb94Z/
kjraAbrDv2BQ27Z0M23D8b1Xs8cjO8NDmx+3/Yz4GcxYJU0ijAqWjqBZv0niZFEBvmySUMBpDoQZ
k6IwoEtQ/s5G/BYJQJ+Pt3D0F5U94LO0pz3CqYePlgCxETiUycKSw+Q4AJLayE2PPGE5PtO6q1tb
UXceE6usXHLQ+usAi8cZRNo1tZG/EBtJH1EElcJslWNkI0Dv1gqJXzGw6M7NoEy9ZMsxGUSkQ+Cc
wcWxLM5eKxWg1K6OT14FdrzCJXIKflJN0PmySr3uaVQkISEq3W4SoZSanOtl9gvxq37MAMfGyxJE
VTJNCgr9FgbnTRH6PYmEN6RRnWNDIJSMAkjUuyMZGfo0/EUMzN7ureoHKoE9a44V7HBBIbOuJKRK
LUDI4BMvehqE2k3mX4iztViEIOH4QDG5S0VMTTFgee+G1Q+i4TLGJIu58iLnojYJIVaJBHTwM4dg
sdKCm86fUqnF4k7ogmmW1w/zr46TJEEhGWt8lu735G/u/g+3m8LYy3IcYp8tVcllh7rrA+pr8ACM
t67oWhcnli5+YRXXRfZWV7363cjL8SPPG1VfHOQ1tufoXUb7hcIB7A2tFwceg+7rBI20xa13Eka6
WNct7QXWX4a6c0eaNk2XQYR7weAITHGh+tslsT1bC6Xqb2dhFT+OTYbd7dteqQx8KktfF/E67rrr
iZlFZqB/fO9bTgNxECuopTLApW0Rly4TNCLNvQK9QhoRchpQF6Xtd9GdH1Bfqhj5ClUZiu6QrKub
s2OVRkxfqXkFahsC6AaZhbzCiHu7/8Lo2F0oSe1B6UYr12icD11rNVqy0ZxvEZYtT+DDXdnzdhFz
4lFkfB8doOa0cW2UZJaVDgnxWoyGGKt7g71B0kDmQ2fgxrrTm2CKe7OB0d5kDZ7KsY3H4H8jJl/4
cUmGp4C46urahDz/bUqIC1TElHg36zqqu4wTE9Dh2Y4KHeFofQ3U50A8F08cX1Y/gGi+XOSijXvG
nqqEB7hDEftXzECU7l0aeMCT8eSxcmRRHQWHlJTFAMNpb6pV41L7dDG7IY7pTyQnL/N4Kn+Jekn3
RC8add+jt+MEjF5dDslPRmI1pFYvNrxlVSkJ/luSyL8PUct+kKq7mHBSSwWgkKcVu1r2tfwa6MU0
O2uxr14jqQ62ow33BOTdWRZhYj/RS4NWhgtpmoGHDpDIqXx3drUkvNpXZD33sFb132PCwb8Sn+We
ojnTEEztr/N4ehnGBa1qsCl8ymISSnFeLlt9yR/o0gAKPFppytLJqv3yE1oV+cl9m30rn2Ffe4tO
BihmWrTe9PfaCvXkoU81xt5I3EULLtW63/cXO11XzeQa7l4EplPArpxHcpwPeb0aKQrVoP4Ig1YB
/bNYC1WnmyCTqKcw2kuH8ucPFuxy7xFw85MkLHUhjaL0fyK1qug9G9Mcoz4PRZZinKhr25SOLwHQ
8HkDcw9OQFyRElPdUV+cW1kiZU3R4GAwJfTE0MLb2lpnIUeJ2nRo0/zwgEo2Husy1IWi8+iDMiCc
lXT8/fOkxtJN0Gz51km7aU/iQ8YRmRqF0p73yd70A9LUfhyTIui0OEMPF9Cwr+AjAhGDX+x4fV0l
oxRIGirORDWQVTOmeNiimc5kk1v6YY38JKkp+koivtzApPY3rQ8boMKHjj8d1QRdVn3S8aGgQI20
dX5+zr47/CQohTug1AE03u39rIvFNIyr3s2512Fg8dxxqh64hYY19QLpRj0yQrrCWFj9kevf0oJd
ZuzyftyfKa2VwyPNsWpLJHsF4zT2DhWrUO0hCmgz1A1cGWEY1WAkQeuQrAwCpXKfZEttuXkHzqfr
R4lASsnr8nbT+Dhje8pXddZmlivinw1EY+Hng2UQIiq7O716m67JmsAdBZlB3nhTB9D90ABSexHY
9vA/SPO78NCB4wQI2X65bg5BMaVggz/SuXh9MKxmxA1lR1JTBaq3L7XZtHVksmmY8SjFM7DCcXwE
Em85jNB952r2B98FQaY3393bsWiidZMGFTpL/f1hqHUCKdO3aQ/+o9gaY0zZEW42LwjuhhYzWWeT
uFnRybAViK7Oai5HKf8OHeRmMvGqqwsexB6mmLRP/aQJ9ghszkEc1C/LVQWdBqUhnwceBpD/kvbz
PpvLw7CGiDA+Bae45hdGOQWqilgpFS2wL2VaxQFnQ9QHW8N+K5clWeRTjk5QZoasMnqA3stDRc4q
y7GS5R0D0qYF2akNts+ruXE10Ci/+FsHGbkVWWk6KmpZwn2OG3i11cNdl0P8wj+gUxZOXAzD5Cn0
oBvVkUjsqLbXA+Ye/U5NeTUfMz5W3X+4kcimS/EB2uBZ1e/9AS1ri2/+49D/kLGvgEs3qWRYSsnZ
wv9r3VUkh+I0yhoTMo7UpEOJka5eHjAk7yfgS382jRQKXcj2D1sdtk1HDy0dtaoQZZg9tGENO7D/
MocMu3y8TDOz2DONYG2xpf4CE9YXEmgcoaXlgM7CVn8lEgsYlhrNWwLKmIG63UpbRoD1cPuA6vDR
Hgy43Nnb/jvPw/78PTSUYcpDkMmJ3qwPJuEXEwYAsB/6LJ1+xg56SDSn1CwQolZYQ3RJbzCjE4SG
bUzjIn+2gQr8djViWwISFRtJvGZC9vX3LDfGIO5+xqV7HCSCARV9/gqr5mAHidwr5gNAgFkDQk6i
gUbjU+yP35vDVO0p5vl84zuuCviWDrSSL+mR6oFdnuIZNHRe1ilLbjSQShaQ3GQq/S3pfvn1J6yK
GfFeKHT0ImMFn8+oNWFMjA3SL4ZWYPusx8BEdwOqrULydO5L2QN1pvv2oNTaDoCrcM07VHSHpyKQ
c5QCALssniPhW4RWeT7EzGaGlsrHYOvDnt2F/QszIIcSMwLl5D0IpAjydPa9IcpOQ50vNZtO+iwQ
Lslv3ETupai0/eLo5GtprjpSZ6kDccFeDx5amFHn1nKSi03aFD7aWWEvxACOTzDWte0WymE7EBHh
Iz6S9h/5MlfcJGwcr0A2VX7oi7pJLEodwdv1AauVBKyUj6a/EiHn40dD8rM0pORMj9QYAy/nWtMN
p0jcwtpN1G6p0fYVliqSOXRhvcxSZd9XaNnSrSz6GJlU2IzMoG3xQQN1+ThQIiTsSbkDVYs2aR4W
6DJQqsESCX7yAaW++5NRI2B6ZKTeSHo18v0d08HY8DGf0+KgI1kTCmQOS6EK8yoy/kcvZpFUICNP
wtu8pNFkmhTWSQda9wuUTzaxOV7BXVhXmKY7yOYUB+rAesdpJ1XLBzfwb6qK2C5dkiYKq0H2RLsa
VNSyCwbbqzjndSVVGqmdbrhmovb8cEQNS5ogvqEQa5RSWbSTRdMdr18wo7q6gtJVY4tpBQWghrym
hDYoOyQ6L2RqnE62igQsdCgDkbRuCgYQPPsnYRWYrqxzI5MCx1EoCol4762040vvFVh4u69XrOXH
B78Gnaxrfk9O6XroYU8oyj5MWb/b+a8pvrm+Cs+Oi3HbipmEprQsZubfUZKQvEltUnF2RI2hhC5x
hhHokVs8EZ6Zx/fJmGcIwdscT6gqmDSjiZd6a43Ci1BmQqIFuUTl1LgcIjgSho0XU98Bonl2lTNq
+0Dwgm5Q7olQAjfAod4b6nL54gtVwWnElyJaxXuMTGzgC5hptS/V/+7jeSncHIlpnxV9HD9wk13C
xmVE7bjAHIpmp62tV/TeoBXjhL4BWZkmubOBUkjWqZ+wu3ZqQxtbpAh7QL/a8Wu1X/BpRUx46WCI
+jz6iZccE8hbecC3p7t6+Z3/k67aBrM4Rn+UNd5hE9xtuGYGcxxwvCewwXINrHSMaYSrdwvipz6N
N0W0BMJivwfLiK/xVbPdoYjBG+7NkxycDvDMuMybvZ3bPV85VGFbnf4gfqMx3df6+b6wHlbI3aWb
gRkOZ/NLK/tTRboIYNCTJrx6sU+s/ENrLmcwY67AnzDT48u1Vfjl/QqJ41Qio5f5rwRMjsf8bAF1
2X0VsF2BJ1as5F6ceFfsCTBI058KoI1aKsZWINdJYTwp7kDSCVGH64u0X6R6wri896EWvBUEx4LM
GHD/Mf4r68gt401Hf5CKss9kmGnzC3uYjiSuioWuUhA9dL/5pwrKyF5VVoXTd+EJ2QRA7hnhR+l/
KCsOHQYmtlwp8hYebuZyxyKRl+fyntIm0S32pjVe6raCq+gLZjbuA+9io+2lH0tv0OSiMerCc6w0
QDAZqFIBgBL/5c+NpM0xazoXlIT2c7O7dy+YStw0en2eno01I4AonuEy/LTeUSnqUrys7YuoB2MM
aDQg5eloEndTtCPMsx04/k2hzr7ujDX3Gu9JYLCt5zQUF5ojT14vK8/Uo25psZjeGiWOWIoWCRAr
yGmzrAaZcWFTJlCbs84OSTkM/1nebWQJ1NfmHhuu28lpF9bjak4+ehgQrh7qVFrTZYhOL5nZJgz3
kx4n0laVLH0pMY3HvnleiDxOPAK3VpwMTYrr7ausv70DAST29BfCQUBVhII2vDSnTDlzz4EFrsEC
unBLeAAsN7wqtgFeawo/+Vy78I+j6U4mGi+hp/7+Ep4r2ghfpGK+gx+AsFQoWpTZEQLJTpMLJ9Mz
CatDIXFoeC+e/owfqYccEbu1QaB99fp0lLUpe/hRRLhG0eUJ2eYRmCA9/hXkC2+FA7ttIUV9DsEt
owX5L4b7mf9GLmDvr4FIA2W//4ON8LQaLBc3baWmb8CzRcOi/wF8s52md7dXDlLg60zcuk9bmenI
2WUxsPTelh7dwoKdvhKBjH91miEfI36ACfzucj+9TthDi9skfLaN7e8l1Hu/Pl3o40IfaU9Vv+qY
dOooaY3QbefJgPAxVHpxV6+21PlnzD3/bXzsqwz7eKBplG3SXMsTcANO753YxPRp29LTeTLx14yz
ApQYW09/ML2Xt3IZ4JMsY5hAWoekWYkTFDWcZ5azI7pr22c/2ATylUUKnFdpvBE7x4+oHVb6IoWD
LsjGnXcK39aVIQbOhW4vjrGdFMZvoOfgMykIX4Sa8YFRSfTq+qnxaOuYl+kB9vOWgMD+wuGVhW1t
ftqCePYDqgVHiNVBC4cu53I3r6OriY5a+9LxeweX5mhlzHvgR8FbsP5ms/5BBBCRc970y4ZNZKEm
zSb4DJ+ijAQ8bCJYNLdp/ebj0uRNa/ObtQq12CLAAhfhcuM4gp8t32LUhHnlLN9Kqax/wbyFjgm6
aUonvpXQnW6nMtxV4/1GYoiqxHf1wDiRG1fPa40+2eE7+d58JdAFYP9bFF/ObwcooRHSTbTQfr4y
Dym3O6MSz5lUnIO2Rn0G4HIz9V1SJQaWmpW32tnypF50C7ijsQhlk4usxDQt8555SGjR6uLuedum
CdNo3TfNDyGRBhZK5V0ufmgueTIZk++DmcsXJ4IgbVz68Zyq1no9tdFEIkgen/iWaWrqPO6iUbeL
/p41jnmI2AO24mAtXbTOSZKjhFVfoZIsYwLtljDrK8z25+Bz25JA4GKDE8WD7cD9oo0GJI+U0jQG
Yiuqv7uWesLXGebtaoSQdA3cwxxIC2IEBsy9k/dK+ohlD7jP/3TiFLrEGV/0BcB25uTVkT9pYzmn
kafbO7nKRKu95eXSkhySuVMlIjdE1k8d39UPE16KBhmc5kjTL2xvPH6VSFhDeGXgqzWEDwDjnkk1
t38/bryugXEJpVU/m3LmTMsASzKnqhOVD4Ts2mekjy/Kwnl1w8urOY1a3UUCOTcZ+fFvB9C46x/G
HKOjRFL1RBYrKaazBhVqG/j79WKTbMJmyawaMhm3ZbijQc6LU39O9FplR5ykpBYBIiR3vLDrUkWV
Y/5z+p5NeheBJo/NehMjLl1jkZ+GAl1xcShWB/vOEHOYB6FZo/8D1Fl1F7lgm9534F83NMslmw9G
uDWaHh3JN0ULDCuQ2pxrPN3FBZJRfmnKzkm150Nq4Qurkqc8NJ4EFWtmcy36BWLl4YY+fVm3w6nY
Gz004EcwbID5PO5uB0DQxbHdIXHEI0ZOpp3s6Vrlm7JphdIrtDISwS8bn5+Xvg5fc1TWFqbAs3R/
70wiBSfV2MKFXOTmj0Rb6koR0CelEj5OloVtEV88tvDu7EX7gpeIf8kDWj8YuVWY51hR02PptkNi
PQMLF44o7Z3B7Lh6uWs4lC7O5NoSlcmCAWvJkc4ercGZkps5Zn+kYQkbyFYeWS4ngAdLSVTlrcqE
4tondTI5Th6aK5sH9V80CleilwoiIxMbH6BH2o1nkWS4gqdD6G5dXhucFzBI8CIKWoTD9NAgRXsl
BMbjhWk5iB8gc1nIoQk3nxkC4BivhabRGFC+frValH29o5hzwnm4txQ9H0W6CTbMl3DsbhUqCfLz
EN/HPVD+f1J/EWBe2BhnIAQg3v/oMIrOU1Fl2rSpqBYAUHoUpIRMMm+WSA/1Tv/9p7oJGQTlH4EZ
E/Qny3lOvvQrvHvu8yiUaZAeMDfYAMRZA7I30iEmlUI2FhX/EVRG2OJvKX6kSPRkRlRRzgeVx5Uq
LuF7CAnDHOiNOHQUxhnqtViq2Yfj/DDj/fIMwM2A+wDpJBgo9sMMcy9GeQYWMEUIiOuoJUAPEXHM
RNnvlQDqnRcNIR99mVmYvnyOcdmLNkvW3T6jSbRR8EqCP3O3PxW71C3Ai9L8JYMbMGM7wcMCZgOX
C0nlLBZcUcQSYRXWcREFDOISerHWA+AmecO5rwkjCqlX20jfG8wmNilH7GFYy+DkX+vMOs4tWUk1
lq9vtf9u3Hdpp7bx4cKbDJXbEAzvLBlerSXy/Z7n8VpRbpmQmB9+T11XrTb6qXf25Wy0Q/2690rn
noDyIBv2t2jPQrlFiJjQK4F7vyWaSR//h1IdontzyAyD2G/1iujCiNEwqM2IGhdI5UmHkYhfaQri
ucy16vhK/tKAUyb60oGcCjGG6LsJBCQ89CiwjyJ9KISJtFKxdGb/dUMLCFTEvjVz2VGF28x/UTcI
vq4A8LGr1QLJf8OeKEnxPFao+AKzSY2UdhcL609FIKO7QBEYKuqeo31/7RwFZqWpF8qt2jfdC/kL
GCyHoNxKQyagtJ+eLSuUfD5jb3nG/juUYAnKzKesX7b7i4nLsPtRN8gdsPdDe3FtUg5GiomLlhgq
iiPDfntX0jy5pVfP/4qphbhh4EVxtWsikLLQMiyHbe5UfbKcWW4omiCyKOqLXtMLr81IJfaJTTei
YBZvP6Gbo0ABu7HD6Uo52OHbnp0Tz5iHKtyjjTmEh7GQPJQXb0Q6FUNt0GWkG9vIR10RGr7RtX4t
YfIwHMwCCzp/cGlqdrXj99a6IEoJSQ8NkrOP8ktDUuXWc97kiTgapIl3OzPMgX4XbDVGfF4GiUJa
f1fL8KCNnpKEIhZGUFgxBVqFtyXfl7LpfQ8hhtn1xE1PeCrynlA80Dd9qoDcNics/YrDy7fgxkQV
CtIluMOQsxbe5IQlOTMRiRNvslMKbMYarDAxru90wYpAhOVSryzY1p/sugAJzHo4KyROefa3ZIno
Jw5j8mktSL62t3JeK4fqr7PfEtGZb5mklE2TtX4Vxq2B0GkF3o74Z4jTBX6SC/AhuXkAeT8C5tCq
0G1UpNwLzbJz1HN4mz/tmFUNotXfYHPoMQCwREGNIPHhi3R7e9YPD1xgxzxYdiBtLUFGhegCTUS6
Sioz32YKXUS2NuwD/g1cAw/3hd6+QOSsu2G+wQApr2VAIRLg1K0ijLL7OqFm6hFw0j4YhnnZNhrS
GeTUaPbrBZDZw+1zPySUa1CjrWA+18WKTLx9DC5S8UHvOIZqPUYsGSgBq10igtphYd3aNWUa2yxa
Sj1+PIJn9BPjKi7GZLsHcWFWezfE2xxQribWg8bi8QxePFQ/YIxjm5r8NTHI8QU+3PWPHir/hN4M
9cJ96lQJ8qOqK8f1T1cC0X828GMYcjgk24WRV7uq6LAR6QGtieIqbKMDFw5GJCAdCDxmig7olTGP
fhZ7ghxtbSO7zBJgUV/WnarbJAr/QvaH6h0+lgSC/CdXjDFfKD6bkvc40bHPNvSiDZgDnQ2tQ2rm
8I+PWeHjyWiofK12/HyGu4MOGFYpIqSYXZI071UnPBJfNUXgA0w3RFIW50lBUHqflrBBRcgfp+BT
XWJ16oKa+N3P/YPuUQDWBN6aPU1I0gd05DaWFMptnG3ZWS+ocCoaPiP1cK8E7xxVeHzzB3vK5eGA
B/l4HoIf/nt6tqF2eA3lrHxaeAYm8WuzEjSDMflrkNFVJqcey5TbXq3XLKnIXQITyCTFsFn3wWbZ
WddJ6jk5bp5qmPh2g/ac9e6ZFcZA1Q2UWmnoI63Wz4tyVykGSYAqeFFLG610y71U2DVdodGLRxif
84eQb/Tmer/xDfWig3MPqRh4RIrMFTzIcwlf+0zX80QuHCoVJODTveNV6eF6rMaVK+1XY65HKnJR
9PAQJQL0c6XJraJ31wE0ebt1jW+jVzPillkNfSqObOMuotMHfqLxormzk7g231j2bEkUaEsE4Xz3
CVHREOeLFQqllDv3ETO6ZkmQKc2uKoe9gbjsmDAG81WXF+rD127CyaZT4nf3h8XVK1Gn9I4bfPII
jSg/Py68sLYQNzly4QlsRzcmWtcINoat37W7e/TsKAGnmx1gIcKcmwoMY/Ex5O6v1gmGehAcmfTv
bsHMCTzc45+sc0e26JKuqy4RmxkphK3KaZiVjJeZM1G1ATxfaWbXSGbwPvDq98o11RK4nnTU3zHV
WxgzP1Hcxon7eL520vBHAMUbF33ZrJMDTuSaR+q+81ICOLZBTdTRsIf4Ge+LHh9LBujaC64fHYrN
+8zIhRSCmVkXOlzrL2IUZkOjN0CfgREtCLZro7smUav2CvuYn6vGdq9it7slQgQsW2wg40k8ngbZ
iIAlPxInMSVthAQPcLiQb5fXG/CLim+MDPzzO3P/wFc+ObTD/ttAhZnhOOqg4xYeJeSQ/q4Ae69d
4U9VIIo1p21rtzMUc2YvHaR8oQZjJTMme7zyQJlMspHUCD+PZOafMqSAOtGU0bsHfxb7QEujSeoa
xbORYpsTDAV1sFxS4M047pOcaTin0fPCcpN/bkV9j7SdGzaYDOoR6gIn0GnYlMe2s2wb7nOQQXQH
yJ2AwJQZgc+M7io7W4tFjhTC8ncSftgilnMxC/lN6ErhAYvlsjlC2N2NMSL91CSFOz/o9/SNDFtx
YmnHgfYOPwvmOKjcCjwgpYSgc2pYhfWE87+UBOfEI+pDIsdWkaXPW7kj38f/gGEwNMVTWF3/UaOG
qxnySEvhSMw1ulz0VOYhhuKZ8aZ3hpi+Rxj/n5YUvakocwicPkl7qDSB3pqc4Tu0wHs/XuaPNjpO
D3QDy2SBJdHUYTGYH+I+6yoU2amkkQmOvwilnYujtDgJPzkh61mqJK0rihWV7dhhiKaH05AbT2xg
3PdnU+hftjwWra0NKjysKI/0tiTz0VkfaUSPA0ZWo4MnWHeg7T3cE9/fuxSCpAF31tkItHmrhQFD
Xm0BkfoLLGIIxakKIlyIr8qK4v9q/i0IFVccW3B/zC/7/gHyHDyfOp5qmHSpyEj2f0yEPY9BGDl/
tO6XuJIOi+1IWBHzbBrUONfkfdSUHYXXk/Z6fLqDSwn1n+RO5FF6qaETmmK/1d9SvlWzOkEpCHTZ
9u4g53pWBujShwfecSd3qThTVomFIKWw6eno6gkPBS/Eb6YKDCq+4ZTzU5pkcXOvRyXDhPMyjOc5
EW6gA953yVwwGMbH0kpzNPwjnEdyi1Qp9NKa3ykrQ7RxZN2GYR+cHHnonaWqP6gzsrHCPm+41Mcr
vJ1OAO4zjMCGdvShavL4sZdImohSGbWyfSATom9kZYK0eUqsJTimMBgkGShMu5bkidObEgK5mYKU
W1f0kKnY0zccwnC5IgdRFAUBWVMI5OqkuM4Ya74tE8rxPS5zY9pUvys5rWn1LOM5zu86OIJTROTD
p/rKLUxGgO04M+kuf2M1VY1KFez9sf0JkR9PvSVgx9sAI3tGnX082xbi+KDiVURvG92xxtP8Er2A
QTx0F+cHcKu/epQOsP75D7hXNjsQ5hR5uZBP/jhs98dFap+jG3DP/fs92ihCNJeVD7/BAXl+P5Ql
R0ytb5d7agCbiCyqMrBqvXEl2+rTP7Dg7MymQorQFWX33fSViWwvJwImF9p3iR/Ke8xDyu9LdowL
iT2DFz5AGaCwUbE1O6HpigFImPuk73ptUcQryEWrge23k1cA3jtNrV23VvpyO15YjJAiW9bRKgEa
lVvgqGfl5VOmu1V9RSRAjDLOhgHhr5q9DJ9TjukA2jRRZBf+/Vkgo5pw9/wy65BZIfsEsDfF/H0W
gVY3/9DE4+4nComIVDsLtj9EOgK9lJg+i1GTF+eKc3AtC/KCxKw+nzr3GqIRneB3bil0WtspAGdk
eRSfvLHQFZNguhWvEMWcLcJa9xgLb8g+wHn0AUytuYteAqbljpzNLgrNAaoR8/ZKvH7lhSFkOU5t
gB1XQM1dO/+h6rO7dkra4xmS7Nuur3KvhQ+NFZHA0F1TDxKaB70WNKS+wAvF/ILT9dgCY2S0ByPf
nod3dRqxDVX/1jWxCkmeY5Gaa6DRYezEnaV6p4liQEfDw111P64jfQMYtYiuDQ+bpQlSODnWXqqv
sw/6Yn7TeTtok1tnmYrU3BIfgYXENal4VwPJTs50O68oAXOlorV0kq+qI03AhrJZ8V2xUiEvR34r
TBpUW4Hzlifj9fjBIw4zh+nCRIOL78KWjHz45JqkB+r38akeZBD3n/dOQpJRY5OwtwvwhC0hWtPi
/CVpie4u8he1BSb5eh+uMBv1lmVbCm4Hl8PVcX56GELjO6gKdF7O7W9pKcdIWoSAnXAPaBizeTCI
yDL/HwtBLK01XSpnQ6tBqtWYPQT+82aOqu2H19Oq0jAGVwwdBfXXhwi56kSTeaqaieClUFA+WXSv
m4uqn25jIivvA7bc1XOUKOHU6bM+4Bsh/bNma0x5tovld1YFZevBNXl3oBXor81U7bxOx0DGPDol
fdiJzZuHp9k851Rk+KHoRWndYZNxv36AbAr5n3g1/qRvXWKgo/mbb7Ho4X9NjP924TPZwZ4eUSHE
bARFGZQWT7X+lsfMHb5BHjirFvVzHLlxhrVw1g2bGzG9fwBLVsyPXIOQK96vnrTIJzBnvoa9Kemw
yyMdG/SRiB8lj0/fo8zcfB+b60hGOfyHneDKhACarY99XdBWlkFMKCrM82q/KSHZ7crhniekAVwC
s6kmyBnr0rBHAzbnrx0i3BnYiXKf9jZxKoBGOZRUFiU/+xB9OVUPE/tNct7YsMmj3NzWItqA+0aG
gui0EZPsy9FGkIVP3oXtb9ieX5mrn4kOQ/seFB+kjmAjDFM4KExyla4Xzq3xFtwWL8R29mhGJcrt
pICw6g6PSdUM48PAc2ahAkK+YZ5+yARXnvw9nxak3VI5Su8KqbSYtGzzdaU4QUlp3fNQlpwlf2mW
bXq0rw8PCq+mt7jY0pQzBOcV94zonzxMHQhsfGzSokSjFBL9dyfcLYQNaJOEGEUX3jWAm91DaY7h
1yVbr5MzL5Oa57U9yjpuLdHhg1BOKUmXyXcsuM79epXjrJQBEojGcBgOx+pZ8cuS3B0C0yyaCVi7
spr2qRmecmrxSCWiRyHnLFCxnLEOumluN8ZnzkMI8QpH+J537mt5FBjCpFtvU16R6LXRMOzZBNig
YHvvtGn0/+c625JOIXNACpE32QicRiBYrJCzR922bMdaj+kgkRVU+C6hmMrLLy1oTImfwQaabH+9
OnZEkMH9hbk2oSsUQQNGo7QBV700fj63OGmMKfXrGVe0eQJ0D0PDPvGKwsxheXYXrPihJ04Ponqt
PWm2SgI8gWfXbgd/Wgmm2/VWpeuBIbqiO+jJn1AFsAq2XrxjcrWc3JmfHTIhvgsBgMmobYewAgmA
QYef0qeoZx5OAakaTOVeiL5fF+SGvcAMaxS4Ckp/LeZicDSUA94/PPPJ0472mtvMcltzMJIuUx6L
ZEqIPWdwg1p6fuSLxm4eFN+j/Z2ow5p6uXwV0E67FxiAFYleEaNGcEbcNosbajDddJ7AbjQW25/5
F0rZ3TK7lvXSz2xhDKVBP5MqhT4tNAJDZ/Y/H6NuE+Wsc4itXiY9koCBSSEwlypsojjZEwjkPIzh
DCjCZmmMmcPPTb1BTohCgy6gUM9SLdAlB1AqNKhAzk/b9oMFrZDmc0rtCZQk9/VKzrIfag4dps/r
631HU6X+NVhXDV0ZrVYBjIuYGOwKkmN82eNXKQXhWBhGW2aADMWwhlL/9uM8P8+fUZ0vfWMsSeaM
J1JnJG3+B8boLYRQdrFmh+nLXGUQFjDl3lxOlkc0GMPVRA8U/aGuTGP8D1iVjINpl2lptHDcpsX+
a5EQZwDpOugN46R1uGfrwjMikTb574XTkjI0HLIoYKJ1fvaD/ngp6jQi3xDkIp1IuKiPduEo24LO
NWwILj7+QJ1ITZ0VY+BjTDaUu0UECNK0+TaxWhydMk0e9UBV7uyIepoVffMf/RLpGWJU1x3F7fL/
EGvS+oTnIfQy4klwUvnbvHJDRYzf0CGNnCMwkYhfFKeeS/19VznY3zFwHniKAFB6Tvv6Khrna/fF
lQBKdZO2kTId74fpdc22JL64rfSkU7nphyzkMAQjUnW/S/EGt2fVoL518EXozXfulFVHukOPRHhk
c5iAnWOY/31UJfd3v4fZjbbHFXB9APHC3fAeCFVUwdaNikN+/r5nINORpNlbjzE+Q51Kd0APbku6
ZJdjeautDOFBJWj0is4JEZQg0H3sFQjQdNGshYWeWNBPRdhWGuVBXV65VYV0cgiSiPAxaO6Li9Uu
SqwWnn7xYvfb3M+8SoKHRhWwimbvwIPNhJO9i07o1qQfYKexXLV7wCqlUwMareCZYWJ6gx/RGM/0
6eMAJp9XcPTecymoFn6F0aB7h4Y1K/b6OAKrryFsbzkQlST8M2vxtGUeob2rf12OBsQKmDAQ50vU
rkGsPwdoqcUchGz3l/KakahyfRiLdHbsVAE32/9tUCzElnB77aNJ71DBibxIbujRHeERTdf9o8kf
eytr+Al1hyqIPp/Nj+S+sMKpZ0g1sbZQvkGHTn+9NVm94TuVBwfp/lV2Hx/+T9uFsiSxSrPgCx/Q
t2BGOvjvY5tTsi2wIFj7Eto+vQlKhWkM0P4FijBeATp7KbOj5CLXhZ7lZzxZOVGkN/zamWWW9Ma/
zDHMbNyA/HOb3ppviOTYq1q+tagB3QvHPyN45nDS8NN1JpwU8/ta9T8RKsgm0tEwH2DW2C35mWfb
YeJjagIfNrX8rYfO2eKWgfiXA2r29efdPBKYZzxQ39vdW+72swtg4utBKxTCWv6c3LHvIfWRft+u
23abmGYuBMSTgBQ06FFgVpzUspkrWy7MNZHbhynXJHJvdJwJ+QLFUAJPuBL3rPzLdcNbOQIDg493
HoRQeA4Z3NlSvM4bN7Bb7MgAYzc1xXSzkuRc8BZ+5Ip07ehtSyVoUfGU2rZlrNNgOtxcDtcMpRXv
MWIB1511AYCxQ8HCK159zFZiZoQHJ+rHNHmcpCr4mkZANhN2gOtJSg+XWYZDyglExRas4DpHV5+E
lQrQMHprN5XlLhK1ERM5QOAF3IZ5VhQrreER+kINXh7RUiBARNY6iFqQM58EJ3els6Nv2SFz2Kt/
Wq6o5ER1FIxpY7aOYLziL6qKCEOt++FMM3xKSYAGDUwhoIAC0Vyb8aDuZ9rODaBgT8GqE285eBKX
cJWZJYyPNCY/PfXujKzk5LSNmXdd1fLP6ps7FpsgtEvMVxiCsy5tL10jGrAe49jbVJzpp9aMzplD
/pv93pBFbXsNIBOsQU1G0NF9HP9IunaHxsj0fp8fj0JvFvPTaM2lQdR2JuJVrhtCWYaNHYeYOpbL
NffFI1NxQss5hSubSbgwx4xEGGF2+xMnsb1YpOeoArOePzYzGZy7dqnGaorgk0tEy0mmRVKN7gl1
tfI8K+6Ua8JN2pXzU4jw5vTHkP2nFb4ZPc6yHpxhQHXD82qYSyC0P00nEuO3YR3n4raDnYjMD3eh
JgLdyOFRXuBoS1MSPcI8h4+vgReT/mbUyXVrmo1SCZLnq83SE/x+UDAOvbVbMQhRPpeJ1zy6P8R7
+1uPz+ToNADPPZzMOF0CKDsTingXFk5Fz6wxs9K+YvOf7BDTc2X36RC+qyYZPr3YaGiM+9V4INs5
fzNTCCDfYtCNiUq3EWHagOMNaXNoHVRIr8bExXspHUzupiGPz8D1fJgpeXcs/mZidksGb135ENsh
ikyUA7WZbJKmFugb4nkhSA0OCuVZBOnYYorp7NE94TSfJE7ikedmsk9PQtdgJvKSZNPz/jnxuBif
CYXbh5fjOCY8kDQwnm9rBVLez3WUYg3mWOLUtjTtFuCEfgBv0kKGJoPo7gpmMpCBef+kdheOrCeI
L/tia7qeNnTGSxFvnQU2Ug0NdP0AuNlcWmhGB6HYxcM6L5xi42kUBTVIODBlxQXyBXjzM3sn6SdY
5tHqM1Sbt+JoaBsxFGrsD8ZNCJYVGAWKEcp+6T4kzp1oD9zO4SswsjZ6iUrS/7/2VUEPL0/2yHbR
Pf636sSisagKSmpcNKXm3aksBy2Wg9g775ZWrteEjF7L+5ViSkqoamLhdXNN6mRi4JGYpZ5bub/3
GOFMm+lrpt2Ua7oGlDoz396a1+qkb4bpagaI96KRGc2bzEZ25dIxpwU4O0rf12xFdoe86XUVuhH1
S851ph1d1C216Tr5IYWdXXvJ8AgkLxSlBc8ghMT9m2Frr4teeecycbn09jeP4IOmScnMUKMJoDLy
/BPTQEfZjYlS+qdXDLjWG8GstXORqEdaKqtyNKj6piBTZlvdyFrQ7u0IwEEaE0oIJp7oCIHh3FvM
EujjVh5pkp6DCnDTxCXeP216tFgHjEzRUB4pDmyTNGpdMP7gyAefdlxzPl/VgQ9nOd1Z4PNAG2an
ncFKsJ30ZIjqWdf22i42smg91O4Z3qnOR0Esrc2M4VG15PfMnw4gUQJfYzdf1+86VLgFYWJRQm8G
dKUe/Z3YA1QmHOOC1ju8poVQ/8gaQh5dhg6LlIO+MyFajBpsWP5+1XBS+nH4GXKrEGo9tbUP+AIQ
qYURf2fO1TFFZL++/eitgzmWbAW71Q0rO4FfVSEJxVLA0w/FfAIXGaYgwcDZJAK15Yn9cZERrYGQ
SsidLJ+5V9ZofbHRPpNy0wQVHLyzY63OaNWDXLJ1vbGFm1q17VEYl6p4A1U7ZVKEOVQRutKCnuUA
Dsem1hSWTGMcUVbLCzaMwCR4m1JCIaer5n7LBtYcS8DGLkK4s6VTEVYGZXCghhxEPDOfFpSr8ibl
ZGzUm/MQKXPNXI/Sk2rv0r5glY0w0at1rJd9Iz1Jm/Y0JfxR2UwzCG1jHUCXxVkZbt5b319LaORx
OHZo8JdqZjEFJezJ3xfLCWG27atXQlTTVjzzuyeKGjATwz01/Lfx1Gfaxhk/3f8hMM4O0XoX4ved
jPqS40w0bVpsqhsoSEwjz/xNxKF016uQGxlmGdViAlfj1/Gsl3BLF7LnGvjqR/zd8USUV4Pp/rED
V+CEe1Cx9cZ9i3SGJBvareDKdRJfLZpAvbW4RzOkGv9ZmFzU5gLHRO78WLt0WITs0gTjxebA1yMh
JfRNyg49AWBjlYgRoabxhrXhYMKoELiBJgsCcTityTWcoljtgCoJnwDiRkA22aaPF3R9hV7ju8j6
ezBkYsXYW3HFMfpQIFfHQlbAU2k0emPbit0IBtYlCCSbtF0PTDuDa66CaEroofSxMbcCVD+dOIEM
EK/QBzPKqz7h+WiNCzCJCafEz7MjFHX16911vQ+/UsFw09PGjaaxvodjsYkGsbyfwd12iLa1z0b+
vBrK1NprahFjUoWWgOsFIgd22OYoHkICw4Lbqhw9u3JFXl1Pt8KSZ9/Or+rQjm53c552kss2o/cj
L3WzYbJMLIBHl6TZTtC9MWvRWEXUfsnxDdNHrO8CXJ57j9GKQC9WwlPum+kEJyCxBIuwergNuCFa
oX1FsgzXDczFRuEGfUo9F2yxKGS+KbACzuT8RbaBwK6MaiL/ygdw1TB9n/qw4kcnAn1a9IuVwZjc
p+ER5W3yAC0MEcJhXAmSQoqJSRPsvvkuMPTai+KNwEC/eCBJIdLgffEFZznaRGVtUj10jbkVMq7+
pB6aWmZMjsafvKanDCVnTchJnZE/uQLc1eeXbqjMhRUMCwD1Ki/TPzKZJCwZEmxE8Zt8mzUmQSHt
Oz1nIqPLfpuoCxCzTBmrayNbOls8Wbp3wIp7Da6EiU23OzBmH8WeHtwZ9dcDdrL9EdVZCbuKjEkg
+lX/lZEp/JX4vUHAvu6wPQFDKCfBdKWrdJu+cxhMUpV0sX/Vt/CUMCE4qBRPM0mKo5zGD8lAeARj
wCE3yhvHORUc1enC5+cvQvzbD4tYWkyhBSF8cxyqTPlqliYl1gh3Izju9sujwAMFeiK0bEYThHTr
AmCdbOQSWjBK1lVL7tb0A8maJMdG7SD24N5n3ywoiNwB8QCUsLhx1rTOzyN+Dolt/k8lfctDvywZ
V3eMzZlFV9GuNeBvrjK2Cv8MtPKaZFFz32QWIoUQxR+HWfN+RUIthJETPFUD4nFX1CBhyZmJzyaM
oMYlt7Z4oEno/zA6MMHXWX3XPo5y5nActZZ8Gzwm37aTqAia0/PiZxYPiaMAUMxlpsIFrlVBV40+
OWrSCkGEK/TkWMb8Qa+MiIcdguAsiihPKgqE6VEsbmLxG9eC8fjxOxhnq+i7Zq/U6RSshxYCEYFT
oCLzAD+lOEWDYKIobBcsT7GLMnk37h8HF6W2RJ1dhSA4hc7S3dkOSZvsfZG7qPGXT8cs1ToWeDnx
4mKzjtSu6/8JU4M1nj74g40zjjK6oDNtKgq5ReirJauGqm9B4+f3dSK5SgWRz2xn9mSwNzPLcMnf
RtzD38YGN4Z+btFJ7YAaRfSapTD7FrYVzehOUuBDpgFvF4MDd+ioaejZ6VssrkT8R8d0UFgOjTjR
i7ukRUq3RfiGkw6MFZfFsL6Gxm4zDdUfw5YqjHv4GcdtsfW2eUma7p5WQXBvIanpYhDwLgjwsU9L
ki2osjwIQm5GeDb3AYFqtx7q+a8LNiI3+urazSLWmemkdn2+pRv1iTS1gE5E9tckTyOfyJYlahEN
vo6uZKFb39aR5E2bRufVTVvVYBcTS2/0d6NMuPxCLS7GSjrhsnSwkHXVuf5xH4YfiOKC69V+VyEK
gX7fqDhb8pDJT4oQxupMhnDj6Tb136JsPCMC01An+On+xvmd8GIGppCsFsMEQ+xpSApJAnYZlqtU
6zgVPpA/LUB3sAZ92ROCdS9u8hQ0f6XybHSM/XJQrdpDqoG2AjWJ8w+1RTJ5z++aK2CRLEXrOjON
UiTbL2RpK3alRpVr/7Wn4GKlqAh1VNAiwz2WGfOukgu45pi0Wix6LO+N0CqhIQadWcIKzRRf0p90
i7FeUAnM5Z/xsaVlepxKIgN96rG+HC+MY/mmjqChhKII/x/Pi3VdoItMjZUbYEmOsv55JO6xz0wp
l52tbM0iD9LXydRCoReOwQERCtX1khvvVO54kF1A0j+RcxBwXTtbUV5zFTC1IQQYQd358w2DJ6/s
E9q3ec+ChBEcAcC314Ijsrby8M16pKJl7tnbO/5ea3mofakNexxdupC9bxNGwdJCrCgA81/qRij6
fl0+v46bC8BL7wBQMNtAyFAri+I62Xq6ywtq/1xGxcClAgbN3SPJztpmfQEITBiXW+pns1E9++mZ
83gktDltWqN91+C9iD2fvSrtAeUe0v1xg7cdx1xXkX2j+Q6DyIFVx6dwZQd4HkmOoB1O1o9WLV0A
kAkQfXusOkWtsqFMkDoozqLcldnJTiCOuaU+aG4y7fNGhtJIoFqU0vgNLYiECM9zzhvUf8it17Hd
SQzD/pG7sRapj3xBa3ne9qlzhMbMIQoNGik6drrgJDDKbwwqxX851AVuHqKmK55tRWYMpk27FrOZ
Xv2bSkHwdUp0k0FawjNsdDMpRCfg6aFb0j+bi0AOg+63frfFYRJ6U/N7XYNpfvcoV9xdHI8mL0+j
xnxTz0JHa2nikAKE2Q5n/9bsRQkfrrYsnOEi62xzhpxiTBL/9M8U1yQDkI3+fM0tdB2WSHPMUFuI
8z8ELWx5TfikfbmckalDWkudreSdpAh+PwVNk+DG8eL+M0Oa1mdqh8ziJOzOF3YIbqzA3QUM8C9w
jfwAQlVlDfjDNxekntQ4fMeGm1hXOZGpIV1M9ZA6LSjt24XY0Toxgcaj+XDj7Ekou3LC+NqoT19/
RGRxT9UCEN6CAIqB8Pdd7ci9fJLg5O1En0oShQtzkmhaAHLYYr0KZ9Vi+XJUKpKHDUQjMuardHjS
FIknm+jvStxH+bW1iuhxyI6QIPSSh1ti+66pd3WQ3G1lfSA5H0CQZ9BUQ1ecVquPIRzsL8605YLv
ykGl0NgjJdld/uJnPaMC6ZHZR/xKXW4bP+ZAUC2nAq3MoB5p9fuiZm03kyH8ioF8ZXCUPS8rKHZM
3Sjg4NcPrxQgf0KY3jo4kWowkog5fmpkvMBh6oRGpYTQrfWG1f1Fz/a6/+Qj1ph6bCkZfL5mvie5
YZgsUSYeEHWkQigqpj5XGozzQUcovm6xm2wPdEquboB4B8BxpHkQmDTTvjhkDFVIdaZH2GNMCpPK
gU4UjAu9VaIy5GZuVlFQ5hh3QcJGvUXMSALc6IRQaujVOexGH7T91kwZJsYV5dJ/0Kqy+lbR+0Cz
xV+3bkTuZfLJ/AeeHO5wEZ4HDQqdbDpoPleit0jEUbCuPOHyTKs3N6XEp7GqGFsuqi7z7BJX7g+X
+4M9v1BQdzxka7DUrdj0bhM8BdAKepcF7K15pFj+8O3fLVMBt/46qeS1lnGr9nXQ+tG3hlS/IED8
kOCUobbD97HbXWXQpTfoOXqWfF9mdn0jFO0osLaQT8ZB+LDW2+u8K2KNUzgy5QPuba/CJ1OJ//FT
bJW/JYU6GPrM2TYlCCo+bCCK9ZSyuL06RjyDrijfNQbSxiLZVHaSV0EQTB+MtsQmXnmo2vzPgTp9
Nuxr4VGpymc6rwMBTKyo2+r4dC2njyRQX8CsYu6zWbaDZy/36YvIFbQvWtDQLAJOvWxiuUO/gHkg
x18qweb9XxGc8pEkgdInxpRTUlNWLBedw6XZjAcEjMl+ackov8ulEOSAgqTgCREfuYHLAbj/wC85
sBaQ+454cj7yjMOIogocn+bi4e7PM+ksLAVJrdUlwPSdDXEmdYdy7ChhEz7CwKevfOUaH7yXhTI8
5EhN2DTVd5u0IoVywny7mPOG2u1fUWyOq6UkBQv1kdEfim9rTiHs7RDtGmiEYmg8NOVlN3hnk4Xd
O9xSXxJPIHzwJgrn8ExBqqWukfSFa94l3yv3Re/D++4fIMc2o49fegAdbeeJyhp92GznYn0MhTHs
LE0e4F96gyOId/su6fpLw171f0SD/HcJqHXcSFbbzEUFmZMIPvdEOYUsEogwR8Ija/ZgSO6I1DAp
KkunVxb01NeL2Byk2JuZLq6V5PjlI70a3MEYBcNYPVIHfeaXpo2Kt9fgs4h1YaCKiL8pntKhwpuf
xkr4pL2Dc/ozpk3wz2ZN6dEYgNJcqbDHbiXJWtkAD/EmcTrUJVDPdaYXh3ic22i0WlaHFOy/lXEn
TRtHkRBKBAYyTTvtnyBU4FH7YionbL7bILhJBLKCypotwikFh4BZyMGeZPeB8RHFcn5QiJK2L07c
L3yQbAu6IES3nanlF6M7uJtY/aX5TnnPLAFVo5KnG7wIMA/dB6MSZ5B9T9CrYQS1fg3RPX51VI0d
+DU8AhfONyIOdntESYZR+oBDv4FN5bPKvFQwmj7dw0bK0Akjt4G5euAQT4yv5endKzIlUA23DfSY
geXDEYfRg87sUCq45jNc97uqqdCToYDP5hmqAPWoaqJS7lIqPwrpYVCHAAG/TJ0u0nSP/ITkJW8l
/8G/me3T/URFOKsb4BnXwmcrSDavsyDtKfuyu5KrwZUjblan9YsWNn4W/ekHA4pkhIbG6H5FzpLY
ZWzR/S3BOe/znGcJ8xeFwK9fhOXmP4080f/KsEfrPiHeWcxxoYQwE8nlhQsIYFdUWKQN60w4js4d
q04kuwOV6rlQ46yy4xIw+a7AqFpu1ftmRx5XYmw/gPFMJBl1Elxfl1w91XVjC0sjLHL1bWqTtWqp
McDPewlg7qUXX0uQwxHkIc7+qhdv/Xo+xccRuVJozwFOL9ZfcTMPYuQCnWufQmM0kKTSFt4kDupo
rAneg+CkDZPDfmphrQ29t/yDKFEhuH7ph6WdFXBGweQbqFI55LWlIX/MxIsejvfCVnAps4zZ8tnr
oVhf7R0pWwQwltKq0fqsc0Ad38VDETfPR2xRndi7hdoFZ00NSreN7iPpVNiLbXY3wmvMM2zNMw+h
6RD6UMXdZhO8n0XKYLBIcw3DjgWiBe+K7FNDrL0LmbOGa6IXeSBjIWg2xFk2c/3bbxNJm503ItyK
K0KQspVb5XgCPP+hTBxtp6jMH6B1iFiOZFB01mLNlbLdmd3FpoOAeElqqkkNvrEF003UNxu/drFG
ApAZtGwGSWi16RpijbcKMuTMy+iCBU0P9vvdOp4VwrU7oxZiWyx4ssdL2UqX5BgXskEF9wuOho/p
VidyTmVHeU07gAHuj1lEoy9oDUnLQoTHCcxds1XHeilv8qvcpLf4TkUy5Coz+z/HNV5m22N/MIpS
o2vhzJd64tQ4vkXzUrySsVJOSdwuFxxAunUzG3BIi2JQCsGihiQoHQa52StQnZwnbtNtguxaAr1A
OX2rUjBWbLRyC+HzM8tg6k+yiglQ/dd3OhNXTlw/TRkvMiIHxhMzQu4nxAK+JkA1e06OiXEgqawV
8Is/qQSi+cdrOtn4kzh8c9x4wmvhnV+CjhpLLJg9l2FZoKsayBkaf+OcGSh4JFl9nXgNfpScqAy6
FLXkQJL9ZF3HUxtPxMIY0oAA8EIjnNYQTl3cKQIy9FTjESEWgo3oR1b8PEP583qdNpedIR2XUoMu
IIXzG9eOPdF6QyrIZcSMih+ob/W4eq/FQzX/hbzj7eHZloZ76Avg9pDeMqBNrRhlctbHpqVN7i5k
sgDTYOYBrDmdVA3NfSWn+dRoYobsBow4MJtXHyfcRuQs/64fMuCGqzpiC/M3esx0MEuaaDRmqSzl
QdQjMXyziCJuLjdk7tJ4qzM4zyGkAJ+2CeV3PQI4YumBkbpdUyWNwpVqEtypMOw2mzxw4/xDvAe1
DL4z9TB3iJeBUbnG98caO+Zj5qP4ubqFYz0ETkEjZ67aa2ojUb2n16fL9JDh+Cz5UkAiuyoCOx/V
hLAUJzRz6zuKSrh/yrXRTq7/xyuPEjaydAZNqw0knDiZPeVJmXhpqjnlaH2zT52e7WILO39oOVJi
y5BbWMhUbQ1BGVbIp81hAxLVwGDQA+64+uoX8tiQfjPIYka6Q/Ozxv4iXG5Cy3zk+FM1GgwnpXWI
/jdxy2s8TcJmTkBtdmo8ni3ZC0I1KHVw13kL+gSZgxCz5CiKvCRWMRzw/kEz/xazteCPA219V3dC
Yr+M8BUZsbVpjYpMOoBUA6NG84Po4tfWjuYKFwbL2D748/YL3FNouMCZv++IId7X+hRlcrMUHqWP
2HG9+d/0+v5DqZ1jeEfTRy8CxXOS0lWpDHZYP6E1ynz4kbpdknV+QqQZ2vUupT1uhYU/XXMX6hjs
IiOrzcGJTeiBHp8bzwDhiE3IfP+exKjyRhBTprrROHxR0OVnBt0UdgzqQvhsr/Tqm7kYAu54nRA8
Kf5FbRlsZXdgDAahqSGHpKW1FCX+AhdeqATxHIyJNN7VGv8D1JhIwAQAIrnhWJUy6o5DPFskdu9k
BGzlXnY5lqPmoXwx4KLxhG6qPmhJIctACz5bMs7vpeJ8+XWd5X3Y2fAXGJDrc50ohDyvWGchGrNk
/4WNui5sFN0HytBPgQr+aUrQdRpkMPmzq7bri8TvIynXkz7Fl/aXpSqXCRp5d8xFk5QEeDgCrC5u
mGhNwoPWr7/SgSYo/mvN8Ca6vUSFm3z5rJ98Bzc7ZOnugKjzIsJ/itzWywWG9AOZwJy8RztSOUe2
FNcPgrPafTVQbW1yUbLrqJ3+Qu825CFD4fwqf8PQvW7yQ4eYS8vRtAbvM9us66jgidiGKeOoCIkW
GBN6spWOx3vvsL6AhxZTcJkUj6ZzFvSrjigAHktgWVC+62sPjmGQWozz3SMRVUFns/JHziuKFQZW
9hBPCAQAOTYcZoarfL9Wesn2MxApqmAR9tPaSgLrGm0f+LviLjw/akEHRX4MfTjEzinxAIeVL9gE
zOrhTmc+ilPZflbdwbD85yyTx5UHmJMZjFyYZgYbJxTHwwRhDwvCuq2ixNLmlG19kwPp9e/ufS33
EZ5sg2abaNBdjnlzGnnOiqyJtRu8cMMzq5x/DmcftPU74TXpVk2Ei3kr5rvvG/cbWWJNHr+t4527
QrkcwWsW7L4BojzxReSIJWyGJ8VLwBd9MhWxoHZMwJWFZFyxIpylWsz4NpIYvcQHlHe8oPdk23j3
iIC0SUiiMfjfEb3r1NOwd8nFWlpsXtDBYbYgLCs9ZxXpiwzwcULTxIy61Qqdpsr6HVqgNmP6marc
oGZLiE3btk7+RGlVTHhcE86Tx7d79EmkYivMZbeS24ehGT0gI/pN7YuiJTclifatkAJISgUni8No
wzcpN6ymu5u1gG301Yt4Bw4AuBTFGxwoqPd4/Tfjro5G/LwnRHc5jkmOrBIVStpu+ngFq95jZT0N
NqFSu6NQEYajbN6emi604ehaKpgYMGqMuxnELKSSZCmmJXQYdgGWMQ2Irr9f8mqmLwtV0FdJeUIz
Xo6T6SuocB2J+L5eneoLCvXzTJ968ZnnRPxGt5CfqBg1Ra5JAoXRUiV8F+yWG1pQ8oV4ZrVOYHa0
qUvCrK4M2AT8uoslNKHo6RnuTn6yBHCduPVjV9tccjkmIk9MYbiAnoPew4aOb+pvyYCyx8RCqd60
DVj/6KBlrr4yOVExhYhChCdhDzUJKOfvpIwPCxhWdCm0b8GAqotg7u/onpvSXnhJk7eWgdoauYIv
5ik0ZqkskFYMv7vAfzLVJYP5pTSPdvAGbGQW35p6o8JkYU+WmcJ8hRoT6PninRD4yVimEFch3fQY
ROMR3YMPN3nAnpVrpJ6099f9EjNu+CqIvTKl2FO/zwXsB5KSnJiaQMr7/Y0UvREpc5cobdX2Brku
hb/37I5VfguHDrS0TKVxoEWmO4dCWsYjxkw2dhoqUsG7iIN4ih5dcmFcFigcskw/XVLnpmtt8BCT
/MJRd619/2tOsMN2sLJY7WlJKJTVzLE34T/HpTLOu1o4R497SYjovrx6j+JQtSpaJ0myGvGra1U0
FstawGFKJLfPA/oBwiB6p1Cj+s/cv6wv5DQ+dMfYbJ43UcZrsNfCa/JvleaSGWa8YFzUP8wGLqTM
W/a3TE/QW5dkOUK0XkvsdeN6YPqfczi+bCN3ODS8suSPDZUiMLpot3awx9N/wHw3HUupQDBSemWQ
nc+G7EnRjuD6+VYEixUEVoMQQ7OuDctIFwVAr5TaRRv83t+JaxCi35aKJnUNjz1u+p8SkPLn011S
P1WsZSSUYnEy7AZ+FvUlYZ3VfC9puHrcetHHndqoqxM0j8WOnbdfWyZi7BB3ZkfgcxW0IaZE8nFP
9alDVg/8U2faHz0GS4OtGTKSz+RPFcPw8BPISo86NLhhJYEoNjHo2ysJSFkYVYcuFWGulAAKbA0C
kH+S1VNllOePMU0EpWLWD3Ehf1q6GeyCyQmUInf3I/1zDz4va5OQdDNoQ93npheShxo3QkbHVxSS
1E5+/CuvQv9BwudQWXsf7Dkc9kzN1w+UmdGxpW7M6IXEZhk59Ihzhik5RA0InUTcTDwQT4uMpngk
HJ1Zn3aYW7JqjyJ6hbYyz4Q4BgEnQ5GlXu+sGmyFPBxmnkYSn/DMMsNDMZzBophK3KSJepkeF1fv
w/JPsV4aBmN0t04+t11cWV4Zvi/wS1NAndC2L/BNaX6KXNPRs/Opo4+8+Zxcy1ZmPm6dFQDUbazj
d+YzTo3Z2eULf2cx5oV/nxRbUiCQjfrvRXI61ZggycaIRU52zQ54PCvRF4HwOp31zeB0L0L+GTja
PkyctW5IUWja83C+uTX8wxexEbCV1V8Mn1KTPY1vvvBb6Odc++Nfk+afGj8eWPO+lM4HXgQ3WSxI
cYKe6VCqWtljE+RMFoHeqLIPoRqY4MyMli+erVFOuYhAHzKaAdu8cZjcFmiHSeTVqHTYhhwPg20C
k5YXq9BYeVJrrO42hOGef30ctGRB+jozoGzeqpbcJS9kgWaSmvQSWT+JxNR84+sUM9/zkAjomnXk
bWbhh/UBBIfKHAlsPTJS/7FBfIoKR9RFLJrPOw/RMoHig0ONVojYied+3ECoKkJyWMsst+C/c9ML
TnovYwI7dAVChG2l2N1X31Wa38JeB/PZl1XaXRnOPccbydZw55Nt3LPZOxHqCMLiLnJPwCBlhEZ3
29Dg83PpoJj4QdV+Muib4mkmVShNRubS1tyGQ2IE5A89Hy/12setESnosFowkH0euChjjKVlEj4t
HU4wDkMI2nfJlJkmTCTifhiudw+x/74MDwWsOgu4HuudIfEeN+myS/qq0r95cg/I+kiQkKOq+2P/
KRBZz3uqeaoyjov7Z3Xu4T784nGFfx0qnaFy/kuzm3Y3AQFy1H3kbPZBulRzFqp16Eo0RC2HAv49
iJeyha35uIOYArUZgz+cfbnsbYi/6smDJ33qLIoaPUmTY+ALhSid9zfCuZiCJIZXMliNnCF+IsJk
n61n+sx2eemv0TM2EUQDu8yAOKh53ha8sDexLbe6oPayVxUaDFHDYP9CVEJBlI9MGlz6elAmWqUc
Ur6jJkh8Q2LYkTU/BSg1slQs/ZRvGv2yDuwC2Ax1um03qGCosDhTDW26JtX2708TvvCdHN4gZTx9
TdXlhsdvgEv8VcG0TfGmm3FeG0vph6EueT8qr+kEMKaoVnDISPU0uOZ4AUU7+FO8OYffdauJ1DJR
mMoHyHgp2HUOTad/D7ADeGH2bQil3WBUz9ItA2LHr284wTFqqO3WLA8CcbV4pxLjizJ7wjgg5fPs
jqcDfHkWf9xliLhudAdbBrlCjkFcL+fxjMnVgTLe53tqm+JGhJD7BYMIFQh3cu+swa/cmptxjWpm
IZlenaEYTwRXKfbNZmezTb0QnsINE6GY+Sb1RecJyxonD3gt9Ley3QV42RERfEB8dvUTKy+Bwtg2
Is+c7b8tB17YMIyPHuKtQ0fST688mtRHHGyE9E9tlau4vh2gGQBuZUpoKd5nSsjdfP/VwXn7f55b
Zu4Ou7XeeH0/V+k6DiOY8jWVmgFz4Vl8DrQUdcLOs28q4qJQcyOELjKHKIj84H6b3qddOhtrKkSM
4IaWRnYe8awjeFojMIoy6//gTVlYE0f9UsZlfymgqnHLnaKrljlDE7VpQqf5oIyTgY1Ak8Ih6iKz
/NlYmkdh3ZsBEvGEgWR6Cq3b+8+FjLgA63HDPzjsKqHUIWFdEyASL+rCQkzsaGl2d83ZClM/V4Kk
Qyfn9kJ13S0x8lLfkEbm5+lbN7iQw6ZPBKk4UOjbRorrfDxBCaUW6VGOvvMVwvKHwzzzgSUlGLDd
rp4dL/omrQ6LY7snHFCftTNKpFBFEEGPGdj7wMvLWSEvAOcKTwGHJWY7fB0GMgOS4QXLKBHIOImT
POfk5vRJx8xPVjYvcgWwhf1fqHCt13FYhE/0S1IgEQLWUf7IefGk/0Jp7qAzRqpayln84qGly45n
W3VnTC1E6fSdNd0Y4SQ5m2PTwTqIwB8uAmN24vc7r9rSilFqVbMlQjLQ6ay3Z+LqIWxCw+wkTwBV
zvuRHOBe5tPYA5nphb9L+bQ/cvurve0ivgC1q6QzQogzAiH9WxkFsDEmG/0YKNickXyIP8xUKPbb
aZCjDagjMrnQ/INSVA/cjT5Qv0Ri8bW/0E+P47FKsEW6Y/AvwdJHaZgQZidL8Xy+CkHRdJoYCqdt
BeAuliMm3YgE2WSm5dzztBryh7zOHYxm3K38hQdS+XLvetZaY9Cr8PI/JxsyZTvfBtDio9j8ZTZr
nKaZmFeRhKl3+Ewp9bTkddJrKQMjr1rphjAbWl3P2A7Q8WTlZOTemeL6hLEDTTSLg3JBOnHr11fN
xb7ox7H3MJ0ZHx31UwnQaSbNwxuctW27gR8rPPyfOL2xFsSeE81y0AZa0Z5hXmMg0y8Ztr7d3/7d
Z5ornUsTS/uLV/UjydNJ7qwJ352m8kFh4nLeRGVDzUr+k6WqxS2fTQBgEPxlFmOGLk6T4W4O7Ehy
Av2957r8lChMYfAd/iaegKSazE83q4MIwOuslST/8fRv3v1a7BcJBAh6kSH3VYgd6i3rOLE0OCHi
zKyKZi+s7zNNgRDRIoCZmTuZVOpj5N9kWaQWyATdPvggMTlMp4kbUaa3y5fHywDDf8SgA5UrIWVv
NzaEqkZDPAi4Y+xdWGI6+8RgIlSQ+l+VR5u6bX0K2O1Bb3GGIg7RowpldyhKKX/FshxANPyqlmnD
jqv2kFAG+4Gt2ys2z00+pTUcHapKRk7NWJevJV68v8RVk7MAOYX6JT9N+BvCe2485R6A5C1TsReg
NwOAikwhndQZa1kjchSfixoAIQhW4oyXl7duiOED/C64GmN6NUVQDzgZscXGe3cSCnNfL6b6Qu3n
NGgfODgewWz38vGupVBapWzzKyEfxGQQpEr/fI+z0fJkRCkTyB6VfYmeNfPKFjNpQ13nTzw6oMSD
jEiwTBVRbrJjy/yoPaU/Oe+J6lklgdwKyiPEzxiRgVSTLx6ECjU/2bsa+bX38QNn/pr9m+VgsrRL
CCPCdmkgn2gbBRtAjLn6hywySVbJrrLdRZr6086nY3ok0zvTt9lXESUB55fZi6dQOFZPDRfpYSil
PHRCz7pKHhQRBfixJ91e5VsdzxZlpW5+SCSPMzaOr/uN/63YoyfwH8tiexOumTmEm6sO88LrDoxx
7nGRC7PMjBeKPwN845qG7H/rhWx7lq/tl/yFbjwt20YO3D3YCCFevQUIpHf78zY2pRu74dhZeY2L
+Q77ONZHwiOeeXjkg85f4OMtR0l/ULt6MX4gQvjVEIxtchNbi+R6JpSLW6qyFOw1PxTslsriOILP
2TgCCEyZ2SINVdjCR2fzhy1opXf270R0ooTuIG2nIiAMIFX+oYKJtnzB4+FuMtl8YNF1vHQyI/wa
La6pqfV3fjhNeGErwI4upFPu0oI+yOBsUb/xryFWH+eB22JuE3dxky4uED0wqENP+XHm5+4qfxmh
vAMsaqEadd6RrNGcPJq8FEy7WUTIZiTx4uXAgEd1t/sDdANSTR9h4XnebgEnkZmShCqC+oWy6U+l
YMnm+zgkPTTDyhU8pD8m7e9hJlgpT5d4lIJwzMzJ77IHWhlU6FN5YVgYaKzmA6kzPWKJJ4Ly0qgR
nx3BFC9zyWVgZ+m4ktaMhZ6HeESEBAcc5kGyHiu9r1f4rxokMIKjA+qyUwzInBTA6ksNDNe0J3cB
6PWhKc0gzsZVG1i1B+epc+7IG+jE2iNU76Eeq7ktMMVOV66+6Chk0rzEpVGN8DoNsTO7cP99QdV7
KvE/u+ovzHws4TxXvHzrK257Y7d4iv6BLJXLKuJx1KTdEtXkEouZBFKCZ1tkriv6nGQUS4PL0/N8
VKP4UGgk2i5taZAfYSvqVcwBsvVwCwP+v1GudSpM5MtZ7sjwaNSGFRKCRmRYi2M0mYZG0qRr1M6p
frgPJ6yzEERSP/8/hHp+DtTyz2A0Lr6BzhLXLPlhnwWUCaVlamN/xByg5UBAGtABOu9ly/ddB4U8
yD3PJ4UQIGyGwlVRqdOCGDqlhEjNcUlchSHHYbRZ59E1rKzwsxFccclHmlAxJaDB3cNN3npTI5RF
XySuIjnhZcMbt59AXQBLzhQOSse5QlQahTo9ykf5zn+iCv0Lf8FXkgnOGhbczLDIWA0o63OSCwbe
xUvZO+Z7Fft4sB5AbAxWw7YZ4gv3JL1hRv5qImsAG94SgFBwry/UokJuch2GmaxXgdFJfoU25qBs
6/G859URbAZ5E2bUGOiFQJ8UYX755F6suiLMcBYExk5uGoeD1HT9RDXbI2l4QDI05mkLy8rR0bWc
l5Cj2TCixHJkbe+y4WjwzYHUzJfSiDfvlEPDr+5ggYNUG5TKjeUaR3tR+q11S1mKJj0CovL98JSP
hmO8GtAr9ZmX0cWutLLA/+aoejWnW6GX3yVWmVGuH9CfKNWUFPehqJBP5GH9zKUbrOqXNqpVuY7e
wwtLDRNIMoNvoEYgSaoqNizQd0mdh1okV5Zun+RR243hx5pavMQlyNqk3130VrG1pVw4Y9iCGoYS
OsymLrDb6ip8XpXPxZeX+jZ1qwtbldcLNsZai/SrBqeDy1grR0gXEzFD0eNaav7l701ruQf3iTAs
MxNu1VxwH+kkNcaNQOE9h5G435G/J77G6Z7Gx3J8/aQ/ZrkrMOoxMp85ugwtqTeaVux/nI4JWlK0
J0nloIEZ5zte/Homa26vIHoBKgQDeZ3+hJzlWpeq907FZwnW/ZZoxfdsqExty3D2ToyafeEo+qrj
zQbKpKiEZ2GI2q7Saw3iD66X2rbIDtmFv3xbglIoMNHxX15SpiwyObPOPA/xv7emgdXFiL+DDdEW
X3kfNQe15MrOKbJZKa4VjPq3GXT3P0ZlPYmzojTi/asQD6XkH/CDhowI+g9BuzCbXXfKTEudq1ay
e/8DG+ag7oQB3rruhiuDZti5pP9EXxsRURX2pnxJ7UI5GoobKE0UIOpxlRlXjyq0oh35d6ZEaiEq
+UozbjCQuyHOjSBEWctFHRd59Ndc8A6eX0aenjj/omIaPNUbOTHKu4rlEIgkoVRipwChcA32iGJQ
xiMObvIRmx4DqOC0jSY6OgEgWKrPFIeeQxh7+T5zVv5qzTy4dqVcuMedHY5AF8UHcUSJtmcPjdDC
18LJtf9NwzdvVeg/tPjB76j5QmOj2OYKecfa+mwp8FABoe45jmTFd1JkD8YouOUp3iYTzfeiOxzc
BFVV5xQa+VWmiSkr9iMq2PNP+/06zA+dDL8ISBPkgsek6NaHdJU6EE1iPt2bciD8F08+wRnbcjBR
3nHE1fNARdt4YoFOVSKKnn0BafjtohkxXkjG03iB4Ah9JXxFtAJb6W1R2xR28dQtKLaaQbMiHdig
lLUG3OHJLmpD9/Nlli0IAJZxpmMZA5idPOEHWAQLdlQTc84OmnOEGtWRL6EHhkorasWGv2nc34Bm
xqjyFdoTV+yWJeRC7d6hvzXZ9XgQsMqnBuz/woVLPCobXHcIRVsWEiSoBhQR0uyuUi1RUC8+INRs
Cm9IhiP5cf1XNz6bhvxv/tnB0opHIUAvi8cjideM+cJ9TCbbTV35rkc5bx8gGTisWsaujXcFi/o4
LrRSMvDtC7LCXlQglc3Ruf2vXAd9oN7aSwRnjpjFeT3tIYWYtSStqG1+zEB/DbRSbLXW8wCf25bg
xwLIlSi8X5dmQNZBr3IJtuyv9/qACAbn5q4PlzSu171eekMkUrTfh1ib5ih5DpEWScYY+Ai4b3wa
9zDJjAoMmHqbJWfSa1DEqCn9ZTsE6Br5R5AJYvJJxbPNT7R/HSs34OLciv99gHkxFfxljPMGD9ZM
/R4ZoFvkmqMXprJOQSDty346SWAfVxtXaU7HhM8ELEjhlToSF2LV0Btc5kQK8E3d9b3AfrbPkHCj
lAUfTQKRsQHHVh5W7hofiVSCK5OybpEPwbDENaBMD9T6ZXobx9dEoGURixNNUxLwMIaz8L6YUbze
Tp0v9xnaDcg6UxX58M+Srh0JmYMG70uJkr47S5fsXf9IpKOtijaU8Gh7mmEL9UjZsXAi2HtEToxQ
zfUdfTAaCbAmrPjNxMyFrIl2f9OqI0ZfEXcRrkQXKjLcBJCeIl2pAqOWyRSjHYj9M8DgPublpAkh
cMIq069xJdzbRdp2xxG17v7axErZVM3y727VJ1uHHqfL/E7M7XSam+V4cWvxGCyZjJoLgqCpVxJf
dhkFk4KumhUP0R8tnbQ8v0rMqtxDb3+uAE0aSwxj4c4qR73QY0fij6oM/gOdBSbgsSTUOWVYXf1H
LGJ6cId3efhCY1snkh9Hr2JhX0T27hdSJLoVLVtpSDa4bCbAL6oWge2VKkSX6W8iRCTBd1igXmYZ
OXbsRnhO1t01LT2wCs5pDxJLlRZ4nFQBFT29UsqUZstscM7ZHwp5fiAJ5ZDJgKZx6JoXcJQpkI52
tUsuf77w8ytS1nM4tVpUkZyTyKcuDVzzGlgyMNrAqkdKqZ181WEacZtmczBvELgVBothTqDsPVrr
WnrOY3iX7JqoRznUdLAirMBA9SzsqaXgUWpoeH9Mc03gJl8QHzfFmeUI25bkbiAAn0CusvmRvVFv
3S+QRDcQfUpwUQ635ubR+omIrdi+s86UcZ+oRyjc7FfAtej2arzOHizwPz8B/LxWB3cZBQrmEFga
1vxqCx9lJaVRd8cgB4PdoT27w9+i8XD7Qkdio6l54EpPBBDV8ooo5pEsREh6MAMP78RT1rWYF0Nm
HcbPhJsaFzxmnpMJIIqnDXGcth1/Wo5Ud2f2jGuYpGbGxPUdTpyhG+4vvp2jm7yHaQu44DzAvS+B
tIR9BKutLa62TeXIZcoJERohasKghaNBV8MfbCXiivx2XJTWGHOeDYgcp5wuipkpOP1TlY1A/BPE
FbYilyN6ersj/iDZrNQws0zSe7Oue4dDT+kv+2dWtGX0RKR/aW5lHyEpXDavMpqaO73XH0d8011t
BBFK2XH6mopkiwfAYY2wsHfOb6MzeiEu9wO5uhP4ZzonDQwKPRJA6zjXAXEbm2zMeuFjRZroD27x
38q4dWzUGlvy3n/lHrSsBqydMmwPYpODLJnJZe21lvfcHwAKINukWIdphtEH2T08A473E75c+6u4
MdbdrAWwzGk1WFmDwbhKLK4VkPNNBCjut9qc4HXdx0tSq8HggA9JD2Hn2fO6qqK6mbxGNvjyoddg
WW2gwmZa8g9c8KyM9C8QK1DdRu9xDxqR3bmBi6aiSkGHmJNB8b44jupHyqDLhjPFa51eI6JgpZuZ
4uQu3qAl6sdeQZ3vOo9I+oSGc5E1+Be6FiSEm9qnrqezLF2QwW/wT9/tJ4G1DTOfBsj6kRlp9a5G
fVrZGjXbsRUaInPlwFc7Fif/51f7hET/ioEChvcvj3ZQfoQ0UwxR+JI0bb9dMFqqXKeyxR57yXmX
V8FguLArhtpfZSFWWBPe2Bj0gn+lVmb3r3y2pyXl4SrpT7n9nW132YTxnogFzax9Vbd7IX8PnvSo
485uJ3vLCt2hsNeB22y22EEKE1LvQCPvxIofczG6T5oaWz50MuqdQJoMOcbA9WH5mZ+NthkdnJhm
83CKx9cf6fx79Iq+wnXVexVPPBoMQFSqiux1driO1hIN+7q4v6AyXyCr+0cmT2cvUD4t9QAyoE6p
X0XFFhAPBMFZc/pZwBQKHQyj6vOrqHfRCOzMR56vF/Sml8rIHPOEICW5cZOQsMx2fXBInH77Livu
kANjmcKW1aX7Na3mZacDGgad/vxLbhSp5DoH9kDXmP8DiBUFknOkFy/wTagWXo2IjHim6TVzdk7x
mYrtJB4uq74gPXA07NYlr6+96xFBzLK2KbzjN5GmelkCDGD2ICPJAMrXvda7LElvpeErlVeDAP2S
BOFC4OiE3Jj9y3B2HsJRFE/vW/82w+AC/sP6oQJNCmQob21pcUXcZVDLkkUKWzWMSal1PgeZ+x3R
row1PbnTvaxyknXVC6mh0ZvCrM3HO1ZIupjG3fS6SAgDZI5yHzHdHIgleyhWaMAiZgoHYW5e3N0D
3UuRshlTRr1F/bTTI/Z6M4+i8erga1NM31gSw9s70LwAQiOsSW5c0Alzq1HeBnOQ9SsSCdQoQVBi
c8WFvvmvS18ctyTkLlkqmSFaXZgqt7KbnfMmas+ycPUWwL3JNTR2zmItMX+SS9T9F0s0tjKCmxkJ
4FsMG6ag6wsYyh8wUxzmrQK1eiJz+25SJNPR45ULENEqksjquVlNDO9uhAYMRUMUHa9IzH+gVmb4
iy9sZsKnb0h2D79mwawliF0okEbqUh1kHOmwpqfKaCm1KIRyWdQq4YuT8Oro6xAgogiscKtLEP0g
I+0/tHFuvnlsmNPe3Y8GotFcpiFozM/HKzLy8Pu/L2DfGAVRK230NfijntekEvOJoHtptYKcQqMf
SB4EskM26R8vN4A8MWrWOGTQ28KT+AdzMDw7Mpi7MKcnMkEbGM2zr84LWu0LiApVu7gMDEZ5fwJr
wG94qR+dNJ2yepHrb2qXASeUSq1nQzAsSQ3Nx/25DU5U9C+oIhNEvbiJ0TK2QZcjJYQ4Uu/JSgWE
lQaOl5DfycfZBs+O6RKzn+dap7XV/vcBY80kKGexDRDHtAvRPHWN5L/Pe1ZHTxSvNvaqDlloj3UC
qj7iA4zAFCfvwtsfTUxW24No9qKduQuEVIYdcr+rr3P5NDWc9klfcAjuiXpedPCoScIyhDujPNOC
T0ZbJrJo/yB8T/g+wv48j6eZSf15rmOMsxOn4BauKeOFlRTKxq1D4O4wF5fTIRpqLg11T1Yhh1V/
9deLFQVd6lV/kt5jw5wHxJw38IoonAUsqHj8s/JPAWIpNHyK3hnWFcCatxBpOWNbw6stPaLpq1vX
F4N0YTy93lUUNXYxWgXawuj4K2g7cxaN3SWGbhpnL07xWpbOdhrQPraq2ZnofmGZMMSfmV4c3Ntq
fMZZIjxMt6jLBirHOb38yhO1ZywxH6zRH1nZ/nQol8vKf9qM5Eh1e1qpk7JV+qaPmk19bcBoX2S6
XxzJ4wo1c4dPAyzBcQ64RZdYDVwm33KpmBTSSxq3MrkhqKb+9GunOeSxNjas+Y3a6xavIRRXM5Lw
gsB6hH3PDNg5fwM29GegX82PSaU2cspPQjawYEacfktJgleubR8sQIZat0vVPfwWWiTXY6B4bWXM
IEGMkneCME+Pje1RYgT4jjS8nmuVpe4hoxAXSvl7nwrkKYOP0y7xm2BemoIiYP9oX9zYcaM89AgS
Cro+nOfcfdJ1L6pp/5pGOMpZFG8uuDF0u368LHhERPEA1KJCmAtbXrDFu3kR1Qtu59MkNLx3bkNf
QeKVGbPTVhODg9FeDHDatEB6+SK4uk00R7e1K9eY2IXIXX8Ycmu9uwUDZYZg1I5GSx1VWsHVjMhG
vXWCVP6Apcxt9mNXogipz/eXumfGHHnX1SOKpSG+zwG3IPAMCJLhjlG4+wzne4zLc63mrzxGAhXB
bn0LVfAjs7By6h2YDM3Hoz8UgHFLPQp5Jz7ZZ8DuosfkpQ73iG4CfLAyU0tN8f8cnHyJjk8KIHIy
x3wleVYeWgd3+zEskOoJPuBRd2/BNXL5yphxItnMADZ0fI0fWz4gHP8I19N5USIpn/FKDsHxAOXI
BoMsR81kegNgUx9YWQZZvS9MrdAoZ1m2A9DpWxxtRKnWe+TNMVimNca2R+MzgaYG7n932WilLVQS
ahkX1Yv60v2SEQu2Xw3B3jmRCrc4eLp1FIDuq8h2Q7a2uChUty3ZIuZ2sZeAujMUxlySH+1FhiJ6
z4hHmOWu+V+LhpdowRL/SDZsIQnS/ELtNKJCtefRHIoTlKfq6eWbFp6wYcvocjcg5iwJNKga2D0L
9WUILzNXkNYGMIXYd0BGwtHLOnHCfIXNtLqQq8zLovtua/yoAUci6ntNqaH8RhXbRjI6VB8ndwEM
e3M7ACGNfBdfq0pcr2jA2MAIbt+omxFUIOjU0d/cjwYPV03HpOycoWBi2l4Mwo9LaWy/sOUyP5u9
b4BRQvVtFbBPg41bjFw9tPSYpoUx5qmZpNuo9PBHkt+ttHHRsR4KDNc76oYGOJ4959M0tnuTHLZz
gvOnylZdMFmHKJLEah+7hhlPxG1yXQVVz+qAoKvuz8iScVnzkdy1fO59y9BxBYSsPO+7OSD4ip14
TkMIdj4iCDJLgChstfEeNZ+g/4pxQIBwIdJW6pxOADAK3V5GZWAzCDx0ZwnCpwMfcb7U+yZMzAKA
2UIdCAlwfKnscd+UQzlW1Er5leiC86d9tWQK6xfV9xKWAvI4rCxkYTnnBYEA9YnqLqWSCxUzZ6qQ
yazYiJGF7ipuLawHtks2g9xw87bKPItLB8rHVNgpS9jci3X0upPJg2hrB1BoO6T8otnwJhP6A1cy
Jppf8LBe7eLD5vWBOKEHZo6xbDBZcZZ636VMwaJbI03VYbhuUYRKNg8S2Y0OWE9z0rBn2hMyDjHJ
TMFkVIX2Mbiwe3GBd4oDQpeOnsGs13jwq+LORC7t7RZ+McsY6S9M9jA4rOv9AqN7Ldmu0OCHp2u0
FrQ+23fBV0dLtuIoFPVqoC03gkU1VnUBv1/NkHVyDDqX3dpjpWzp04+m4a71fbwUWDsMxDACChLX
8ozIxZrzDtYsxGLAs2mRniG9Ug7fn00oKE0Q1L61ydaQVRbSQagrrm0d3Q4bnDNRAXAgxb4wUZOi
KslSxizIYvFdmHX696PSbooG7IzkSMRvJRV67EQ25cPP7id1NpxWiqgWiTOd0uYLf1pDYxK5PhFd
fiKnyqA9xbvCGHEYJxuXde6hPl8De4JTujzarWpnnsVtR96PoyNjgvCKGH9rauuIBDvVrUCoWouY
T0oTGdadPihXuyV+Fsyw78klYfV9TCsMlGe1TCnOqKZ+KnA/PcWyBy2Vf+z94XipkvPTHqIiRPO/
SsE8Z73i/XKu83FaXXvPl0/IqRkC+qXXrzpJDbQM6J+FntS7b5Jy4w9BiiGitW2bFX/x38s06B7K
65Mz66PcIQ2BiMTYT6eFzWiMBoMJPP/snxDczIf0izEK1YGcAsSAaqZPMzXJhzcITdjrbm8ksDsd
lTIq3FrjOxc764tWoJHmB8jO1A3oWykjgmamxmsXJNQ8t/uRd7nl1x9G3fwb/AJooBEpcYld4ZPn
9m00U8kOOgu0EMo5XncC0RNcUEyQvbTnHeaVVKK8j6Ht3fdq11x8QbS9HIioxfkXft+JtRjTWE6e
LRoXcRl+jKkDGeInyF5CaI4dAOk+CxUq3PiMVaaD4dKuiFX6gFvf+hL1nDpF78CMrt0SNuHoSewi
8Z70Z9mciBWWpy9Ez5Iofb9iC7cJ3TcdLtDdzUsXSIQ68y7U61pz5h5Tx7bU9QCIMCWjcarpIFsD
zuk0wEdXqTzdk14xGqdWzlrB2VHq1cIS1UYDCM3i1Uo/XsRCyvdLpO9luWPba4QBsCsiRqwOZXfS
E5fvdQcSoDxmSxhy7e6qBhPqpTeuH0ZPi7AfWcKgSItxF9iSV8LzpZT2vEn8ZFksL9KIvXyqJbHY
4asT+fehxD4F3Fo8Fi2rHkFCG2r5hES0wJ6j6SkBDNlmPfO7IPUfjQ5/VICKQeMdVIwTmJpHbgqi
HVhD3RdrpAZV0OcmBGnYb38b54XYiK7M6Y9xarZrUcXcaGWQmQS0V9XUXQRnBaxij2auO73rfYZ3
S2Qqnh75SBt0LNtsoK8fGu3FYGJOW6lQqfd1JH8Z8DpY5tla9ZSJus+Sd+SVYoulMHKrcLRcjsg9
6jHCf6JcCC3F/ZxBeL6w5Eh2Rsmt1rsoCYZD7z3RrwLKDkxz7qj3RFkk10NAk8rsApk1U2bQHOql
KY2gDI8SCxMKDGWPvjkv4J+uZosakNCcshXMue86Ll8BFwU+B7lkkH5AzBCAxkWdmgmoaemT76xy
c/HO4aUQXs+v4oVporP/JduXtYIYVtyxgACflVKihth9cbzJxWBI9qQAqKo8+9dHOKHf0AMpYLNw
uqGZb/FMfogSzeYZuMnwP34+rYt099vpTS81m7HLbIhISsqCr8MNgHUE0/ZyLc2OOR9L4K2DRhsB
/N+J5wNFnA1qHc4d1MqF4FEm1w1rMErTaMxg+yxy2kGrOyGWfUDWfpUUI4IHCYHoC3CrrMVX4VNn
S/ISqftKILQZKC70UMe2q40LxdU0xqj5Fkvu4mkAVXRbN23ACgCQDOrcIearTcgghpNgFoHy8szl
OFMb5NRovaQUItuz6pqbfOrogI6xzUozGMG5fdjB8SXN3eWkVh/0e3mzNZskcPrzYLqzCnl9E+Xj
Fy2J1P/KtP7eEcCRyuYTc3f4Ptsi7pGgpSJaHMcGM45uZ7TiEpqf/goi3oINIn2RGv751M47L9tG
ovXfTyTsaxByECIqIKDSA9jbtUOq9K962HlEdGlm75ff8DsZdlJ0U0LeOXe4BC8wLpUpCvW5Fojr
2JSNYgzxQQ8odR+jW1Dsb0+x9uoPLxb6eK8ZrsyJlvABSnjrvwUKGl+KJsJ2tG0tLWTO3w/PA8PN
CEkreVzBOuKkSFNJx16OdD03VKxZ17FrUG2me6m3FQNU5JqXI4aky8mAwD4/Vh8FXJJ6rLNziTle
o0Em1wPGN+7acs8WwG+SEiTzxznKxTgAmFJtDfMO7SsFFx4Z0S0dmDnBoOeN0oOQF/VPil09p3T3
2gXwvNc+aSg0dQ6o9sdrBNqeuCigyvaNfLoIqH+K3FzJNWDY8GaZHSOVHgfXo4Q6S8VYTUrQqZ6G
XU94KN1ZUlUVV757L0fSrDiD6l378LDOepBJwHEzB//uA1e6EuAblxo5aRxOfSppWHhaFMVGuajf
hEnufqdMZnc5ki3QplQFl4DoIUi3+TBr9+w9JOjhPZzpLCwUNkGxX4186roCRswmNfVoEbbgFa92
rb0rhM2zt4ogg1hK6gAeqEyUU+56fCjxexlWavEBeBWJ/MiNpnja+3bMMtpmIlvVXlhtyKKNOQLc
CmQSsmLrPuJX9/71R5WWLMXgjDJQPDbhC1kqC95WHlqeABMc1sey/U1bjZkNxldE98QpQxqNPcU3
A7RYmCqhBOXQDITq3P6SQirGMvox4/xckPkjdQCAX1oFgylf0ys80z/0PxrKBJf5EORnLHLevqM4
1LgPhZuk+62O+5TWnx9cGGBnsvpdtz8RqjyOmxy0GWpBMMJS7YQInkhooeAw4JH6shx+cepJ0d9y
UXIJHNjBnPhNcPNVagcTRc7Z0Pyr7MoYJxRVNC6R2D46c6hMjtYLHHtq8dyLYJqMY8J/CYMtWFSx
eA5KPo7cKpYMQdy/cSsx24aJMuhI9cKrmuWW8Y7UBhTzByVDGn++D2Ab+zHXfvMjck2T5YMHep2A
JK3d06nHoq00puNNXSiJ+okc7jd+1MQKjFj7IsB3etIM4x2wJNgwfYyQ0RtaWqlZakQHpf6/i2Ku
HYlU9qMfE6pxF9MQlVLmS4aw3yf6CtbUxWr4IEjoCan9lvG4VTTpcnFd1+ygYWGuzznNKzBWSMdt
WcOV+c7B2u9N2ewa92QqIUj9ly5V5cVDEzjEVk2HKsK5Cl6AqwfWLjXhM1IDodX+VWSXMEYEPply
Vo3gw6NQXFxeWLsUR/rWmgJbYyRRibGJ9tQajI/vSwwcRx8AD5Th5dgpitI/01Z58Fi2ZfLPVD+d
8N1qCYGkTrwbMNxYSj8fbyhWOHV7qQ6yNYGCJ7Jmtag5WDKxj9sx1s2lHLfHJirRU192LLhrjmdS
/j46Ng1/dHZ42q5CN5GiJMY2138AmSYf94WQExjC/OXLtGUdfIrgJKE4rR1NAEZfqs6W4VcwxhQn
LsO4XtwA4ujCgvcjMuiV8yaH8MoJSCTVfZkZQB/XREgq/i5uJ3+vIe47MLFl0cj2rS6au0EB+F8e
Ac1JQlso8hklnZ67ilsKdlBSQV2ybXEmCQaTk8bOm0Lvv21xOxaZhQh8fQLrmYirNHgIV7eBfUjb
zwHXgKYD/ZldnovCgLAavy0n81WBfCDFqZ9p2GZiWZM5b7bEIenJQdAkFmUXkrAFF92QlCttnFNB
EWFDIbQfdQ1jOZkV+OsebrfPUek9ufK/gGSylCN5gFnVRXNxeH2oTUdzC/UO9PtfMiqRwxCLLT/e
1dyNlk+AYdcbyiszF0VCW8myC3gd/eKhiR3Xq4HNYCRFRzbUq90+1kt8/FuH4uvWFGLFXweYYH6v
5vZXocPIOKn7eJg2jgsz//kqg8ezHyqkdgCcxmJIBq0eAn9nyvCluqHMYTfQ8YAyctx5jXj1YRuo
YhaPQsL4Yf02r2fz0La8NLab0EHpn18pTasWbdTTVInGEZH2sz9gpWqD2X4+HPSVzLpIAgux3//n
O3vv8wMZbG552vCBjXPwXxBHGN0TbG+ANhi6RMyY7946fF065NewSixrqEL1VrZlCZX9jZ1WT/u/
/T7ut6QeHExlRcjcReGbl/QIi7hv7pTRJKYyxlSM2QOs9YxSr5fqUJdlGb6m5llpwusZfr31Yax7
8dn3ZHnk5imD7yqM/vqACmWYRRIi6KBhqvt/JgltP24iNqMvb/N07mRJCFO5xlWgRwfEbm+a+yt/
vhbljsuFlDkOrQAcNOdxA0NAcUJuluxpAYZcNfOPy0PAHTuanPzXOXwTG3brivj1JsiGKfZPRxhF
xJTOO7dl8Bwy8OZy9v4n9FMNf1D3dxqFzGtqMGrBCoX8WrYaBPYt8aphA27GvFQV5g4O5j+x5hqZ
CBpJMLkNGggVYmxglj0jkqmL9u/Jea9njsY+OtOPMRN0zPS7wfg9SQGYkea7CrOfBWcxXnuYsCgv
RB1moJRCAgSZyhyaFegxbpOFVFlkcu6DGpETdcpjQ6hpNrHI6CPrcYAfn6zWKqf+B02SxGXbp+xC
0tHVH4xFJ7sORwAmW0OwbcvVjb5PjBPk5Qh5+XA4vybPF8DkdlDF1QVqinInTaqfG5eWklJ3yPR7
otAR2DqI7Q9khmqGUPOpJ7qLmDSReq3GEmS2K5MIQc7jVlliRFPeW4VYROZcZiP1p81HVO0Qhz4R
bus+4eoNh8y5sLFVWhPTUDAvMjc9cJTtlbehdSSAzBmELG5eSlys5Z3gC3kq3gJ256jFvxWjH2qm
0jxOqi/8Gjd0jUOpc1AM/WpDv+dIOj/EXgv9+1Ptr7uqb39va3/kIUYQuZnY+QMWasAU9dnGWQoE
b/2fduPEsKY1F3zg8M88+pe5t1Np/FBPOCCDoyrO8GIQhEwDE8dD9IM9BtDAauGQCioThdLkKG/o
j/z+qHpwIcydst+6m3lCT7bQYg4379wOUYFUiBlsj6K5lNGXKVZoOjQSVv2C3gW1ahG9jJ4ugD9f
BRJkcMWwG/JeUqBUGA2pmq1bfi82ojFAEcJpqJjTJ3GdmkEvHbGH1dTyXB9UPB8RadTITxwfY6TK
iPaZ9ZInd0ae/DxU47/zA+7xITl9C9ucmsMeJbp0UTzlrOUwfMf3nZJtIF+LnF6719XZndmIqnpa
z+Fo/tUyw7zrY1p5rRt1XP3mQu4W8Y8NpfyjQiCt4BHPlPZNprOWuoDYEoCAx5Miei/9OiOQkpz4
RK1q9TIYi3xqMVh4Athb4bxCuaSGEnZnQDYVMWAAsgPD1l+xTiYBgqIEWjg9czqFE1KFNOZsMBsA
wlsWOKbmrxBfnz19egrLClIK8QuvPQXFkYEBMT/N+y/wsBchUi4CI7uI0uGaMGGxmmydaJu/9RTz
JqTkD8ddfcg0YCdbYgHAeqXmmGxC1CHsZLpJ/Wc+wltzQ2ihHUCnM8ihOfVNoQ7eevOERul8Amll
fyq2KFw3b/BBTVngdu5ohH1AoWzJpD6KKrAJH7lTnQbOJpUDfxAEq4EvGbgY80ZCxfdBY1I5Hson
/mZ4JiTR0opaLy25ZtlnTLwRfoXs+tEWg7xDVUsslTmNx9MnUm3HPBpsRxfXf701m1JGZiw7X5DK
TQn10sWhIZcPCqY41jhXMOYrWdVvScxMyWRlSsLzBkd7+ZQa0XIxMAQ5hus30HMyUfvM+HBg/nUU
Z2bpjgvoXrslYf4NoDSjEQeutwJjctbItSyljfw8FKKkXL5aSa/bTwMYs7D0/oEm43j4vGDpjBZ6
ajgu0rl0swEhY1U0lxr3b14gOe6CXRo0UihFjaO5UjiS/5OJ6W1TU+FUoRpUBcBUZy0muqPGXM+Y
lv19USzLToIrTrJBowr2LThzHEHM5tFbYRZL7QpRsTJDTLe8a7LxM0+oLPeXPrz8COF5TSAC3kng
djTefbhAp9vG5tap4znPCgLoyXfiBqLigLjjbcX0cp49sNEX+Y/nyxuCFhX2+KRGu63dUgwbBoGn
lbR7D3uFt2d9fkvyIyOqiRyZbU0x8bYVcRVW61azGaDzRyQS+bi9QPnXGvjbgtSFtJfPUN2gtoxw
X2SY2oFnXLjZj2hS57X700xEBhMkow9HK68YXQkXJT3bgv69pG1PNSkzCLx8tXdFNnqCmHTo3cQR
57/S5HIoxU92EUyNLBOOs5UAVYf8nV0HHRtXB7oZZO9Fxygi6tL5+y2r48MTt9UyhF+pA7Ij+NVw
uJIMNcyEX+jSHGgzjn3sVZsM+sD+VvRdIkbcHLZFXduWIxRinGgXJEjUL6KDYjpK0oao1hlS5AfV
FRCttTWIAXa11cAAqcYBFQlRucOnCbVScBbjbpmPLpb8En3S4eAo6pwTKNCxJnuobo1asJaN09nT
PaMmU5FYGPrOTNhKWZhfIp7UwKDtD5F7XoBhXSCqgRn8MGnTrLPg7RCzOj6NOnEsZcKh82sy653X
ljIZsXUGn0X6mvw7zz+QgQQr4Msn8OuQddqljyURxp4VOmmitzrvmnLG+pe2H5OBEMPKnBYsVHPv
5qVJP8VZEhRZGzb0amS7OhecUTweYiw5Qv+GSPP2iN9k1aOKzxkmGjVZ6HpHSN22AFpoaSPbgjQm
4iNhZZ5EOipBiNbWBK7J28QZ+ETiErJtRyPi7zj4vhrQO/u5AILt6eek8sUDLFYcJH++R6KbK8nn
UubtQFSSDXef1GPVruVSKrd4KcJyyTPQUsWAGnjjQ92acSd+OrGxN41y5XBPEivzKIbCQklhikIS
6ZNi31YWY+IwWqzGqTl50PXnPq8qJ3CO7inanUOeP/9gjPW4VMTHDhDHwS2BfFRTlUIHCANzauR8
5zKynIwxQx7FDf23eZfGLuNbZ0Er5gH1cv80EVP/+YiU0qlmfDlt6JSjjLm4NJQTW5fKk0PKJnUp
E3WG9gImnEWPmSKSs4ULViZx1akhg7CTfYgWlcnVYRon68XoW0w7FF0Ivxjyufv12pZdVXKtHts8
QROiDjwDyYbyQmVpuVG7Y3kU4WwNINvoP5Sj12tmkWj5R+bZKIcXu/emKfunM/xcA7PZCNrlMiQi
882tkiva2MoHl2Ry7HyxIIumlZEO1U3NNHhdacFzuDgStAp2mk1KLyQC9gRG1FoQ74LobvCJ4n6D
9xfMuljpVt3OQzYwUHI9cYIQwcDTrA7AMiYjjr1LU1poGDZm/Xrr4hTB/FOMQfSieifoKslXy98R
JPhzjSqq9Ak8DG0OxczAyI4DKWOr5NGnOlc4KZwYC3/l0qcWktFlmr60CYxR4hmBgp+s9l54kovv
ayiDvYhJhHIqBqf/TYfP1rIjTJNrjGePYAJd+Mc/xMcYHWQPg/XPXWIWRVstQly87DGn+vK2GXWe
JnJGlDE66sTYtcyh+Nyu53AntehoU896/9hgauVXS6aBKDbFVq6S0sqsa1CoA60ra72Sdojj3cCv
ewWq6791LvajdxvqQzsqYSze7xdSTWqw7f5xUrLtGfVgcjmu4vXQUlYcr/Qux+jYlAFTHujWTQfF
gp3WXKMZGHPQ6Gn0pSWnITvEe+8NHM7Fr+k0aH1qz0IasZpsgrMAAF2BM5eYY+PArXzYmCxpPoGv
a+V7vFI0NsW9G7jhd968rbEoYF4WlD+3Z5qw284XFHtYx7GL343gEbbk6diOnRNc6/P+Sj5/XfH5
ZjqICyBVk7nW1URqYsLuuNb5p9b/6isHcR2PZM9raqZUZVLh7U1klbf7LYzq2j5ZObUmELe9HofX
8fVK+3vl+XSjJWc1yPlDWmvbm713jUI0ZiYtKb1uaiS7cBIDdq8X5V5VWL/DhafJWBOmEORPP0V9
GqozeWGNhRG6S/gZ3zPZeahyWZlmyEphf+T+5LseijylS2cNGyJSEyQgY1bF76wvsMWNUTl0o53G
QqnbAUGopcGchOou6yF5zXYzL9acTrwF83Pue55v0bVRYz035dMukMOu0rBuDoDqCwCxMTyFS/de
zrEYzXLhIXLupOR45ArIbu191N7F3aiVC4ECT1ZfRhP/B1RdVm0on3LcMyaB8/h8n1Qit6hAiNl2
gZVzqkgaV6Wn9m1JniwpFb8LlZPlhopmt378l7uOgeZrJvCV2UyIQir5Pf/URdqYD83A9FXa8eqJ
VaErk6nG2n7CAZY2+45jOl+0003jJf3u0zq8/+WTBVPusqS27j80APd9nZD+OIKAoDmotmqn95Wh
iaV5aREEVr4TKzROfgziw5QfxMALetEyu3YrRwr/ZHPHTXNwMmGA/BrzmKxkJRAhsw+h6FJR+3yP
DISVmbB6GoGPpsGdEomvyMJSYsQEJUVsOVS66zsdMvqXrKdlcvF6mivIdbXrsg6wLtAixXP2Zw3Z
xj2xrLJg8rQERFDzdl4hvm6f16kQxwjWiUglt+N6TdgD0OcYNDUl0HCuzgEX1AW4Nd5xRl7go53e
XWcBv7SSx8gX46/fgpGXSabMWgELRKMlnfVChKBWPKg3YLV1ufSzOmL2+t7bv7K8jSuDEHXyQ4+S
B3dZwQWSe0UXkyP0HDlql8uwaWgWGbyQlvzSc2R57GJ2OpKIVqVuis9ERUt60fcccMrQHODinNLx
CbRJMMuJ1+M+zId+zyiVvgRFZBef7Jszc8HNkGdGh2gb2EZDDLmABvtZaMWi8HJe43z3hOZr891L
udbWuVyRv6k49grIGbAiD7bkc/ZQ0Hak9CKSnQaAKoq1VcNXuy7V1yWXVVUNQc6WUrE2NPbvtBBa
nC6M11GrC1sjYIONx0bcFWIlWdGlYyW7ZAQezuPsRWPHRwg0HSvnbBeKlEtX17YjDkjTx7L/CdG+
lvqkgD8FhX/cYMdCDkt8UaraHv+nXjRzaMPUFs0JkbG3U4Xob1STZqT4HPoxcNU3tpyXAa96ayZj
qhADM4BZ0H0QdYocfaaoa8osEVM0XhNfP9t9lYay4P5tgfVazxUPrO1ayzNAILaZt9wO/QtFUi/o
G39mSmQ5IBfU4zEkZIoSPMBoPAgrYJHEGyWV1RIzxnIYxqric+iQ9MAvKBh6E7iqE8jacNEedNrN
p6rDBbOBm0watf7UUtRBiy7u1zsqi9SsCj9fmPywbqm0rj7s4kHrzuEjO3kFx7k6888VHTTAjlL8
Pi/K+6jlNlo6ax6tCAZC+R5toBZOQvbnhIdI1uj3eGZrpQ6LzRjs5HYiyl7vP16wHicYm0xXyFXO
pmzrpWjmy85xf30HZhSq3zXsT2diDajPQ85sDDlN0X3RqxXy8JAhzQnvfOnpMMDTkIGxHUOvMzJg
R2teVPQmHeNWQV8vu/VPYkVao9l2YliFS8qApSUpWJ1dW6KuA6gkZ74OojP1ZydNro7nt5QR7GS5
Gp2+Apw2dHRnxZ2R9ePEuxT+AKirRlMDvbgmjZCSLEWzUcgYtp6zJ5IGrVbVo2XSXsUy4oz5yMPn
tLMPP6qXam1p+D8qhzVpNAnkxA1Tmz+tJUGOpOPlFAsLkq+Iq5eZhrTDK7YGzJOHFfg/B+lqKnKN
s4XHSDZ6a0lMRWxTxUi1Utmf5FT4oQNw07/Qb3fbQlBQPEPhH1odQQHDTRz5XqCuc2QJMZLDcfVT
A9b6DOFQPH7IN8PADdBNTtekzxaVD5mzBRbXpjVTvChjR0okbBre5fsZx20eLtHHRtDFNsbMr841
jieEYBOhUAyK/aJWeQKdM11Snasvn6LbY9XvkXVSObO+ebj7rvs9U2jLO825OelSXwSdIJoXZ+TJ
0LTcftEN8xdlMIusZj93INpnY6R2kIUYd1AdQDvIoi9toGiIv+Z5nhplvIemkQJB7mDlnnto6AHj
h2/Bbmw8/kAQPnR3n/gsMHfVc8FM8hrAPv6K9ZYEgXDarumHmncrt+wUtmhF7QqpIYQe9rYMCneg
xe7qPZnr/dxVSkOtPDy4b7F0c3lybfLpkHWqP6dUsu6z8DEZYG1TfCPZ75JWcw1Xc5I2BYS3fCJq
e46OFJD0/PrSzFKUoR4J27w9jEykoqvzM7vNzUduExM+zO3lr5s9l2Zd8taBGyMvYv1qhIQVD7Jg
fqJ2FnObdDNB7R9Lz9yD2JKSm2GfU5LrLndTGQQO8D/NCxaoK7Cv3sCen0njCg8TOPrgquHDd3le
I6Ffqj+WXwOqVXnGgOZrLsvcyVCF3OLyxJeWURgvyZnVsyudEzcBcTYefSVbMei+wFJwbErpjpM8
aVvBiykSAfXbY/l3u4g6j04D2z+3HtOA0gryAaRXVZ83QHVB5/iNZAqtWcfgKyWHJbB47gNjMi7+
dJvXAe0F2P+40hP1y0E95zVDaYCBXABqNKMHGNnCffIwOoG/SoFget2BGZJzp8oBo/dXFVtxkGYp
Qafg9ejQwzs9SejQqS7H0IVIL4Rs4n9gD0wSk5uPwgdfW0DsX6ZLnYJDG/i7m2LgV7L+VLRNc4rq
+WLlsI+EwCk8RR4hyBSIwKIwLGBlVgUKsRYNz6EgURMOLE29hV/EobpeBEtiMYirfNsSnyj//KZ6
f+LKdxkfZB9OA2oL25z/gf+iaoXLoBTdLz/zCO0dm7P9rN6GuKFfvN08dvyw/IoZQuWKxjzXU+pf
Qswv94hpHPkKmplBwgYgDLDImwfZuKJgID63E5VD/qGOk2CrZqM1ErPm+OK6DXr3NU0GFNJtr6ud
veC0WOmoNBlYCrg5t1PI6Lz5bNCMCkTJTt0ehPmTSgZQbt302HI100rQpiemSRG5kZkkTCindzd0
9Xpkk00+chz2gq9wJcZpPdxNzswLDpiifJEVaFkapqpHKNgJ2vBApODgxp0yDmjX1WXjeg06zeea
ehyDmR3gdXCNmEPw3vWdfsv1IYxY27+Jaqwb5kSSWFf/hCiZXRzU5fEo3ln1ecdYodcFToMoxAj2
oU9kn+1H8JJ+I6irnUzgL+5zeTC1VbGfojIk739YQCxzCtNKHXuWu4iN/wN3ZDzdIF+kmTajiedj
7aLeqCJTko1RVokhSHpM/Ok0kHnkk4rWPZLEFi3hGJl2tmpCtMpYeSJcs+vMmmxMNk5osOi4jO0E
+cu4ik+aWPWDAfp9IU/D2zMOBAgREaYzgxBQzrXdI6LyoVtFLW3JPaW6mtj1ZPD3yz0aQe3oj/7x
i65GDY/YbxAz8Xc1Gqchner8a2ltGX/FCP9VrPJqc2sJru6sqwSI67vgEjKsknA/1jAke7y3AZbQ
dZTSQz6LAGayKVwXOL2tTEo0AcBkS4JIaoQQ9jczF7O+oY/ByZRQpQrmWJGXjkOr6+iBaRzMKUKe
vsn3ZzR51j/9HSAf3AoyLIoNyTIg43+S1/oTyCvsw+i9DpTgCbyKNECe6wRbOIiwruc15SofQaoT
VVr7F1Zgcpf4oCjRNiueAm6MceIOptq8oHRIAR4G/vyNEI/yHgZ7VUyvPRhznhMmVr5NtJrvm92W
6HASy1mLR2OaeGXOlU3BkcqS7cmNL1uj66KVn4zmz5Mq67kdAuEYAMoPeA8HM3uBkjbCdyKHT1r8
IXhJsmpdUagHppSTa4j3WmEHsPIKziO/20WY8GD23Llkv5HiduNh3ZiQzE/8XHLGi/edwqYp4dAQ
G/kzyW6JNazpyVYuxopmS5BmADF0PNlZuYFNCXLQxyjAxWmhrQdu+sUMyHHEsEf2vSeOpBQ6Anhj
lztZC4HlXeVEc5l4jkGvfwHRidniNf2h35b2ZbGxNpFwod//PBzLbQgH4MZXOyrRuusdJPvuA5YN
1m0FV5Lxow3uiduM3p5zpgAuBniEnM39E8Hs8aN0GIhPqhXKj6PAqUcXfONX9r4eAuwUIrNEKLno
Ey06ovbrgeQ0iCx8JaAPkn+XVjeJpwNbLIl53XhdwW15uVhDk4LWevlljHKjQEtPMKS7Kf9T+88o
ak0V1SmTGGzQeSDeqFGsZzubSwohq8H8plB8qFMvqKnc3A18FUawI/PPQ80M5jFulP5HuJ8oi9s4
cgXUI1OLoZUqMdXZYPaVKEeY5Od96rkHeA0p9bJafwkhVD6V7uptIyLmHcNJkf5Fhd15uHYaY1Yp
lMaET4c+HvBV6NRmjdZ6+cOACJnwNQX3pkpK0eXYPuahj5Jj19YkKI1acY121uaT4aVDCeROZZnF
j79/vAhqcyNC5M1WFeH9Jpt86JNMScciViSocy13+M0AbFYjEXPIQLHqgwUcP25uMarcoF0m1p5M
mk7h1+rhmhD0DZTdDPhuFV28GgJNtpnBWGvG5+IRrbIYH+k6dj3n/blx1A0wGtUHzDj/05NiMRWZ
H7B00onPYCs1UYa4WNX4be/DOxcugMieWZo+Uptk5Jf/YVKg0blPc5PTW3BfByl2OKIP0AbsLkdL
eA2SpnVBXkGo4t0RrydshOCQIiZHCxJpjkv+WhlxcBM7plGHGv1K8zITiQlQ8jr3lM1B58uOxgFR
VVYB/qz0hCvEQnq8L7jO7Hq5cvUKn2K12HLYKUu4pZzK6usVU856Q14J+MZ1+WvLUIWqV84bvI9h
rD9qcTJaWClhCUoIEUMkclcWqeNWquKY50iPDWnp2SKHCab4YaUD/TafLPuNkCq+t4PlmvDloRr7
eeXQ7aFQkvkXRW41Rbq2LAzMeV2nVZwLvK2l1rC1t952dyJ5mJGOZdhxL/6NoCIIoH44YAQQFWKU
pL2KL/PmPabHdtxeUY/nRVeixeW0n+YjHgocDoAEaEKncOC1eYVT+wI77wvZSTZ8nXMqryq49Vxb
e7m8Wf+rZlmB4fJicYJ5DNPAudibjDUA1egNRP+sROw/xQBOfvgfj+s3DYGuK30rvs8i5IMhBWYt
InYOD3CS5bgkp8fL5A2JgOqVz64gn23AeG+Lf0+gN/sCJPh1moN3MqGYJNS3sfuddUaWthvWmQqj
YY0Hjx9W9d9w7SuWDShZ4J28lNnfpNXBT9SJdX0ypwfrPHHx+407Bq92H0loXsBmHQBrweQDszYs
ojjg1DIMWvACHNBRkHB8+PgHgxXqKkHR767A7jXmc6POu9G7+TWWaQR/IhtYfh9llUBgbT20J3Wo
m2hSIGVXn3OvNrQwi76byNlsW8XqEOKl+r6lwoLgR+RbSDScoxjvY7JH9jSu0wwa+xXYQpQwFxkz
hUhb0jFPwL4JiD2Kx1paCZgN4nZ4L5f9uOrox3JTpeY9c8gBSb1qRZAYIYVgqz2A9II/GEseYRAX
YUQ/6ORAnVgrv43nRy+zZoETHLWTzaJWtyRWT7NaDpPwY1DEcII7FE6Qxc5CkvDhyeynHaj+zPiI
fC7GIFvEmFwRFj5utgcEePmpw8UJFosaECEsM6v0NTNn57I2e22feBOJz3EKPSV3z2Bq1pPxwX+O
a/yl8KG7tC+io7U0qTNDuFzRFO/cz9mC6vj7pvJvEdM/WNbBPuJNeiK0GqW9AWHZOqlDu93lLkNe
5ZgG0Vc0AedTphemuHLpZWUtPGyI8C5agMCg1evRj+ru93hfEf7ox/eFGeV2N0O2o3xLyZIzLN3i
p8c+4jKFqfgr534dmId/4fiSUlhM63siBZFDKSCWRqirZmRSE/an05UK9CoXiI0bZabFcqgdOYvy
UMGl85HAp4vE0F+UZh47p1zM/EW4jXvR2DQk88sh6BrXtAQ1TENmOXiBb+MMpGz5yS+zSXUJKMzd
oSnPusHrxduiR7OOWLM5WMvcnekyqnJw6zUelShqPp1mBG/AKkP3AKXzLZljoPhwYMvx9tMEKjVi
2h1/WGUmBi/ore9B2rdNG5LmR4SxQS7UBlV2hqHQx6jw3nNygeqJAwe4Ckm8W1oro4hFrvKxit3t
gGRMfiCu81+ul8bZQK1o7bOsEWKopVbmkVApV99aSPEUO52iE2yHEY8LHd+EUN8OhRKXSQesHcfM
rZKq8jI1j5r/RBmQ/rFvsvz2tYM3n4Eht7zElE43Q7h3nCcHuQ7onBIS3HYQrhuLg6AZaLiWyrSi
NNndxqi8Acl5FZDsLWovAnlGWkgPnmIyiTjoUzZRKWcoaVSlc0Ok9Ic3uJ3LrzQb9xeLOjX7s2tL
+NBK0ZIMXfidHAPXZqnoUIsgjTOmjCtdMLQ1h7wbB8BiGxkEFrzwDpQ2l8sLEjEEclloNRXDYLgB
i7AlbQp5b2pRfT1++k/k0b1XNTuEsWdzcT1pnmlTXzQ9GlZ4l3M9/LqIOC5n/Ya65HPzgCQzQFmR
T4H71LOJotDJaxPigmbsf6fyzZFJLX3cMAH6RtUz0xkfInNrgBEMMWuCfjhVdgSEvsrWryg/IQF0
oLSRnBBpw4yNqHVXG+K/jX+FSFbQdObxTtXkFRRveBEOWPpJJm9ZrzUTQsWQJVU2Ly1yXQjnNX8g
cimvIMFF8NnD3S3/BVcFWfr187XA+Ek7QSa72CB1AZkTQVfsW0cTQ0p/R2SPzqJWRxkJnOqWcZ3k
mqV+BKivfmr0UTml0w51cVoOY/djo6ALJvOKCApdObVKjLedpPIDSHHwurSWEfQ7TnvwbdJWt+zh
pQko1EPd7rRCrvFvMZvBNGyOTySTCF071is1b84/aKXoMac2STPCoWfcuiL4IejqioRbf+T3nDy1
gdUq0q8R8heVGExPdruN7U3aA4AuoSeVVgt1JEfzWZWcH0VYFgj5Hg51bHYPpisHm6L8dFXJ8A8X
OAftKk8/5wIigkWvu8AprWhPW2pQmjClV3e67mg/2TBfVMpNuMBluyKwr+W5adUQaOrGrmtVibPU
uru9CqMTREapAWwV4rOOLUalKblt67zyV0faH9b9qHXAWyPDEaaO1YGDBsM9gvolqKP1xHxPRPGJ
WSWWggVRs212U0mEAv+ncVnl5tCWJOLLsQ6WEY2RdeuzjGSLqXj0C2njyhT3KG63BJWTsUq6TNzj
ieiD1Q/4cpW+3chFy0eofhJbwWoYLjOzLRq+XyfX24G2M0a3nxuBCr2rAhEKsRVdCY3NMhJrY8MY
P8uJd5GF7yws+PpzbJb4NuKc0VgHIrx0vCRSWvL1DeKdssl7ouPjH1tAXWqKCnnHh86wHPmQkwPq
PcCHcpDVz5P530pIxfLyHczxa/3i5tgxZfAJy25kaSD8UClnGkMF8+/GlxbNArwKrQZJrrHt/T26
p6uFKqMwpPJ5wjjbJ6miOYNcIhyIUaWEltncVMxrX1xKUPsyKZCWXqdg7iK/jZc9xKgTZN3Uz0Cq
2AogzFjjtPk/ciRVhZcZLLjiZLNWpQ89yFvRpm7+egct1DU4ljJfgCTDWIzas+6v3lpiiVvCxiF3
KoEF3k9DXzcFRPZ9GNfdeOG3Eux2juCIrI1ISPlU3YYU2Go+mfteaU2wNJFSuvRgWi1FJq0arxkR
9qGHSfLjReasjyA4irkCh5cOUvw1eAF/A6+Uq/LuLzr1wzI4nmcxuyfdg5CeKw8cebSgohNN6KRV
Yl7r1zIH9wQ/uBpbaRVQKKV47ZS5YfPULtsECCe4Ceollc2ENJ0QLMB+04NGS26m+p1V+PaMV4T4
9bWiujcAIhx3BqizrI+KFD62yNuyOcPq5Zxm0c/AbzIq6UfYevItK5qD7OF/ZKjto8rk0AgmcK8l
wKnQBe1MMJt61lwB/qYE9tLiezMuuXBHZ2weOo35G3qvj8/FY1jizVIzQUWr9dxUi+gjQj1j0j0y
+E+ZJd1yMgs7duFTmpDtQkyg7M/h/XMlS+RtIUp4q3Ja1UKzFFcPddTDrEGX6cfpT7rhIlC4rdP9
UKXJp/y/Nd1NxE8vrMilKXyswgxo43EP3dy1au4SPfM3A5PZ7lGfI25OyjuYKdLkCq/gW12J/hTU
Avbj3sSYyMyWPW190rkHSU4bVX2KvE784SUIdI6+v7jObI8coeUymyM2LzoYzm7KNiN5I5ghnltV
bqusb2tgvfImVam3qFSCyGYgi0jka8rhpDaHuX9gglHfMztdQQa98auK8aEgar+ZSjAJg/c3tNmU
fbizW/3WQ4IbaRMP4E+ptBAhDgPlwGlxOazVjt8SnMGc0hq4sLEjRmTWP2rU99DzOBca7LAgAgS9
qeTk/lMYfK0P/Yl0KYkFqJT4Ko60xNIpZVpowbFn6O0AhhC1tzk2/8V0Fv2FPwVF195aUrNFEyRn
/m8ZzTCWF5z3m4hbjMEkvXabXYJHONd7piQudp2639qYV6eJG8L/F//lezY4KHMQ1uoKGtnSCJ/M
ugeZ/J9/Nn94JG1+Vj2HeI19ZcPVwDmYjS0FyypLTErSH2uTePV+xVWCw6lcD5f1HjLv5LbPzCUl
NDC5DCbwRHBfgeuIdGxl3pOROzViy6gymI2KpftArulDwF8ERd+GBcQm55i8u9O1p+lJ3tCFc0w5
A8iwTv7O/nUD6jQVjOrJa5kLsU6+sXM4HqchpiAXlWfkZ8DfffMsIaszUBxJis7GH+n/EXBkRPHy
JrixygEO/s9sRu3RGAMrJyRFHzLKpu8TcU7zPmRyhCgxHHatp6bqVp4RxOcL6NtBBKbCzMaGRjJn
fiHwhIs+gjeNwpsW4HQgyFOahngLXqGs09URDjFju95TRZoUlxCPevgTnLN4gRb6wuAdTIgkWmTy
GA7JDoBcKrqOPKhoEVZkSAR3Z15YFOMVJYIgmEhwf9Lm8WFVJ9pQjhcumzLyQp5RkEnaUFQL5eSO
dlBnl0qDtQjqcVEeKHqYLTjaXtBIfbnwbX7lkbuMHEyl98Qe9XyouIc9q6VVK9JPyhfCb/pkTgn1
ip6wvFA93AjDVU+4sqF782NqoX/z6d4E/61QKUyKfnSioqZxQ+oBbDtXDmDmjjiI/lKem8KfVorm
gueWjCBEPCxDH0tUhxrfFp/1P/ewl/UekOPeIIqPJiV2Fb3bMM3LshILjWnw/anyL19SnluDLLMs
Dk1/yZaMUESiv7d223XkO7MiuewJAmfMJsWrqnDENTjAMtSkMZhKEgYYec2/H5fT/f5EXoEmSQRo
4YzEA8Ajb12EN8jVxGyiimhZe3T3sJLmOXvPPofvqHxHX6V0K0cWK2EYCS0PApS5agveDMhkFCfR
RcUbNuyqSqiY/xFiqZrlE5mDksRsJy1eZM53d7KKWjJoEBKTigTKjiZB6+fraROR+Fs3GKjupuZT
4DMnxK6TZUIjHGNad0USfIPRXTgjDs0vMymiMaD8fEF9pXJOW/itrqT5pn6s/rwwq8H+/a7IcIsz
zYE3DpzxI6ifVNWDvOIwNLERhGXmUHjLg5Q2XFSDoyuZWbkim9024OCF2XjOpFtk1Z0WpED/L92g
ftZf/0fFT3VDo3XLGA+ika5pX3vKLs9X4OEr13z0LtGrphWOwsLKyMG3QNKfCSd/Ee5FjXwJi1lV
b+2/gIC2ln0OVlMgNmi77MVr2IeuqCQnRmmkvTDglmaMNygX5ZwVEepEIqpR9SGwlQe7Gwg4LTvy
A2mKyDoUnQBiPK3S5do7JgRBDn4Kn8uZCCL+GlbnJWNQ/dJ6HkFWXqd8T3cowlZEphGO7mtUlkD4
TZfBHe4fvnGRoufjs8WlzfpFC5+QRw3fMECnYRok1cipLwQLYCoGOq4zhr/YhJognNLZCSCEVaq9
lIZ/4A89krpbyajvf14b6PmRitBULeUKs0nZazB3pYslFkzZFmmbfzy+MYbl5Iqob2vsfYHRksve
mPMtJVyqs921B16nx0zvLJCeQxb0gCbU/MRCsFErGEsflnLvFRMmOuypGybs6OgH6GYODVIPXd/M
hnLS73mupVzlVYryqeJZkPPcgfvqi9vy7Gx4kTPiiIK0AzFJDYhtFNOoG/Aq2+rLwGQGbA04iTB7
lZFqx/lu9x5nQhCn0OkX5CLBVyAYEkBHY3zlE2yGfGWDrfU+nsDVPQdXKrmvamXEb7WhZZ8iWnNK
H5hzRe0zaEIzggkoRsg4vF8iq9a6py7PxRujG5VSO1JqmmMeg1s1MmYMiG6+s02s4wAPd4fftDZ3
vV5LhNVtxMxGYfJNs+f07bqrGo58JwqkOudra1E0xrJ7mcSEZKo/Xy8+a5ymIKHCAB0FNAbMoD5F
VpFI3ULd1iqIEffFyb1p7bLq1/fnBwy13+lWNXwTtSUqP/YEYxpZrKboU51qOxomo/Secfs8r8j/
+32c6Q+sHyBHEsSH1eZue66Flsk8nNT/APXD2JNe4PJ0CIgR+syb7v9T3JCTX+oJCqVU6W3vnSl+
R/jlTtRdwrs+J7haLte0mdElWL4kvXLhjbR7OrddqLYcvcKOM9H/Rq9fMZOeDap19uixKLat0i0R
/g9XU4cEOQ9gahx0r7dIZ4qfu/6o9PKhJ9ryxDsMzBGt4Ze41lHtxrrXlATEoKRhk11Tw0nMEjiF
uPN/NckjuzJWvnkHo+v8ROgCUIivOomgBkXNMQbovffMOkbUu30X5Qg+mit2g8BFU0a7HuuKZf9O
soR0WZtBM+KjkZlzpjrTRAA/umoItN3QfPQxy+ezdM4B2UY4fQXvpntutz63hjNdNQqAPQjOW15q
/w3lK6odIBEPVf+yYJEEcWWGhCFvm/vanga80p1Pyl+htl2FNY+IHwT8UM/hJmT1xxBISjSoGeqc
DezKEvfwX2ZfQP75zihJI3GG+cRQk3KxWrrbzvAguMg+/XexV7iiIsgnQ91CA4i1ClViaYbaY+SP
yfnRcVXn790tYeDU5AyQ8PKvJ/nMkQJm9ylaJBXiiC1lxxgeaa8c7lWabinUhbfr8bC18d67BcKi
P59AZAPP7Z6rMpu/DMw1mFlkx9TVaSPm1NG2o4wSIIZRmcPTJPJ7eTPE8m4G7m2tbvUg5+0Q7VXB
NThtRrwZxH8N9q1FpzAafoc0VoE2JkuadPz7ai8sjVg6APkgG8gvtz3fxXAb3zhRbKB1eQuBd/ni
mG23NtVXpw3FV5IUrWwCRsvBlkxBm1KmAbBjzpL1UDRwspmVQWUnAMGP3cbxDiavpcOd+Vm/LUlq
ki0WSOj40X90yKFt3zoNHS0KFHTcEnmkH/R6GT5sWzOSuQ1B5Kpi32cdQILdi4rF0GMjPyFhynIT
xB2P5liNFCczQ7jaM+4WQYlc9zJp+Vemq6RvXPXeODDuDVoYcJzVCA55kKrlNIua+E4BoBqt7EGc
EUUNtAyAm+StIaQEKMKN5D6i1lQc1A86dEgLoAHVQuTeWEAaI1XclSJf8qZjeOvw5K5MwA1+dwdT
3pYT/SEdzZYeFu7A9caJ5WY+BWAqgMYqA2q2589N03HI56TAJGMnQ8uEEj8j6jOrqodr83zdsg1J
KkeDsr5bEyVHk44S7GBywX0hF8hQ3Z2DdVoqW1wfO+v76XPFmyVLRGtGywiko44o05uKcIBCT3c0
8qyZ3G2Yi8sBW5JvTQiVr3zzx6rj3uVA525+H+XIZrYPRCaYWwoamXY5RO5hMoSvRdihowsTFIsS
4AJ1uZ4bdfS/V6DLAK0YRr/LAbs7TQCSsiU/c6DMaeIhN3wmg+fckIVtSaDl3CNt8sRru4m6vhaS
mKsXy8wUhfQ55KCilG3+2l4R+zGxZr8/J3PNAp67lfByxwhPUre7tuKHN7Nd9qNKQBilr9AIfZkk
6snFLTqZeUCZHDLYPcd0gk3mpx0GvlggzCkEjmezjw9sQR39D1J08Nc6dDZgKIh8wFr5ULt5clds
0Un89ErTgmPnEaJ54nGc2ImKyPccRmTh8DxJQam8oK60LNGzso/m5MIlf+JAkQQCzGfyauaoa/Lf
SYZEAvnSF1Tt9Fb9fkA7gQ8tQLxyx/8aT/5U18ipgp2cQlH00awZ/ncHCB7IrOw+yeqwyC1ydL1u
/vpU83J05+k/Lp6JrPyZ7cYJWD8li1JyWvBO1sQLcwwKhsE7OaohW+/L04cE3DqHUIiiDVdo6Bph
wZhMXRoVrvCvxQycIsruf9zfRH/5rk9GOlbBQtD4I3Ewl0flf9VnUuudEXAhR4FDiSQ4td5mEEYw
9OdZwrdlJlJup/7kJZrtfLA0XYg0rSo/4qwq1mzVSw7F+3j9UXGLNYWHFyWuvMnERLTLOYJjnT1d
IeOYTMpmA0q5GY4ibRadmm7ERImZBKoeyST+GDAup9PFv08uhw/HM7Gq/UTsQgNgULN0ha19qKnO
hW1sTgGpIZ0ePRGRmR68CgDKfvUy/p55GNqZCdwO3K1s951H8uIcxsa6c0VYpvVnSjwMCGtpqOUx
uhcmK/edSDkndZ/nSRmSIFUmNggTx8TIg8Nuianq2J3DybjPkbJ4uGpsEKxNsBXHS1ESmdhH85Lm
DypBGCaTgInIRASONaOY1/rxFtm8mAWICJ4dZFeL2Y4+ZAMDG0Lje8vxApynlIw0nw2OYOull7Cl
tnop2idG7CXREbkyyX0HuX4Bz20v6hmv63dU/Jp9w791QpcyxoxV1rhLnwnX4zBbUONkv/4ZyoTm
IhA+BhfAPyOqf3IA/me1XJ2PNMeR/cNkVQzvn5SB8oj6NR1DFKRf8ZsQCxzesqHpc5wsRg2Yx/mJ
TQhaqoEohLzJqNCEAxfXzfKMxFAzb4rTqMhFUZI4wPmq1vnOLDC8Put4Ir08HlRnS5rpquYqk6xB
TS4Q12/M47w9RKhjQllZjdmg1Q017c1Z5QKX/VRP99PtX3jACA+kVTMo+Jsi6isZWjPU2Pxd228S
qPXubZ9uZMfN4cwpmphWa/SnLLVkwJs0Ol/Ei0OBPiGUlgxQkn8aD1So/pICJNutbj2aAXWpzrIr
Vk7Go2S+FkAW7WtTxTKwFPmlXgB6i7o49U4SS698LjfVOnvq1N/6kUhyUPoWWQxZWVKKOUHJBZDq
9pwrIP1pANWxrbk0xmElmi9s5W0Asn3ij/brR6GYqtKvgdRcANOO/oo7zSHog4gvonnUYk5JKmdb
qRL79Vmygg9ziKXs3x/wYfCAzy3B98A9LTeOKFECsUqTzb0tkq+J4tU039ctRkmWcUc62fMAAqtc
lUq9nBbEhSVNXJXBsmvbrTMpMo8EjIqLDb2rZXJTOAqSp7bs9oQ2NJqJYtLzv3oPqnu6TzR5GMDW
KpyQUjl0onik9HyDyUn/+T3bery3Gxd0OJ05aqaAzrdG41NfhVreobcPSAuYN387GUzhDDNWG3S0
wRgyfupx+M2smoIo8REi9C0T4lQDfB1M06aIe0THKX/awPfrB8zSqff2QV7WSXhykCRHfwRl2i2C
TQWvkuemPGvHEU2xav/1SUK9MyPiT58rh/bYEorO0518NSXbwDEDhsRi/+TLhv8o7PLcUhOlSrBi
oGH1lhIjU0oDeU3y8kd4o+Ej9ftqRYH4LLW+Mg/Uz21H+DPx42f448eYP0Vqq3TaRXf1wXXG1hC9
JYkA2FB/4PLbG4LwW8xDnEBLF7mzrXxE9Rg6mOUzwMpUXlB3NLb9lL4C0kGe9idYtWWKgCxnl5GI
j6M0+EkFDUQAVcYh5owLEg6lfm6MewGfNnH+qBNgjBmqGXbsz39VN4ZQdUYOHEG96khc1OqiFleV
7EBTn2NOKyF43liYEhW69uvZYzipqvQ69TP4sF3JxNQRvwq+0t1FIZO4gSW8rh/uFSXUu6Iyz4NE
00QaKOX52DSvfRXK9Xoe06QXVTM2Axg2FH9xaTf2JoKEwsXlJ7q6CioHyjFiKsa/BHkMczjQeL8H
U74TnTa2UegFe7lDQYUL3R+2NJ9sSpzVsq+tnl0MbIGHHsW8qr3mkrdCyiQYalHv1Z7e97OTYhXO
Cj33cV6lXpCRlgGiQabYdiCogISF7ZwyapYysEl5HNYimzuwmvtTiEU9Uaa5N+xram0trvzpz30Z
QJqH8oPt4CVGvjya3bADTDXyQkX5nZJTq1CNjClXmnC6UJdKr/3u7SWC8Ts+deXMpq37n8+mlqy4
Jkz+kFwMIJQEhXmWIkrdE7t7a5GmLR5kL30YO0xym4CN/AioxDkPZTdUO7nh69j4BRBrROgikshX
g7tS3sHA/xYNhhBzt0Vbel3GWmfVPyTXxsljZ6r1Y3spx3gfJz1XStw0ZEokiH/eoLHnOWsTToVU
HAoPqM9NHlPhRdvkWclJ6h+2CGbOZViVHVNM2FLFVYXfrTs9yZIokuzxkbBelrHuyPeHu6MCbS4u
lv07lS8PIdPJrUPcmgTuH8Rmla5gMIoCPZw9iUC94s/jYWkXFBsjozQsyUu6CKLQAV9Z2XCkZgzF
TZ4XNxftBUInROQjNtXryuZRVEaPQlFqvgzkeKCJ8ri45iAGdVacnblLANqFE1TsKl+OSeEkeub3
I8JOJksgcy3OTyVeUDYWwGtlv9nKto7zFGCd8N6bnwHX6yl5gJXMy1pu+wgSxt2iWRD27qjT4h8J
ZPWWU+9y6fuGynELftGAddoyVGzTa9b/6TCLY5LAoK6cb3cQccwCsKMeJ1qafflVG7+JOl9izE5h
oEYMnRc8wLWjqcFsfKz2P/mvhNBc5AwBSnPthDiS6Yb5WQYt5zhVTgQt2O/rMdovSWtn9bWMcmUx
LTKso08fUGkZVKnG2Wa/5yfgA8/EuE/9de4uYJ57/iNCMRwaBpOVZ2WNHyZ8B8Zr/0/sTWSazusk
gbyRkvmrjN432Xk2LHrLaNXLZ+gXy0VYD6NHa9jWkonBt8x6LOriH6e/6L9IxyMY++QRLuGsGMvt
TLUeuNGfEw8dS7nhVMaR6aQyaMqB+sN86ncxdjJOrNOpyL9HxvpCKwQZ3nzFF1aK5eQ9GaRwTA6b
pUsWOQA4a286+zYaFDZN7VIsCtqtVqZl0adhfrUmxuEKPTx4dnwPDKi+mARmOe2/MNQYoMWqwuES
AMkTgxBI9Xjbf7imUQMCVTermBUTLmucxhp0unHmzerzv7zvDimhLpHKZblgENNwy4WjD4A+mBFm
Oztk8T0Vm0VIH6zXJgaecwySqscDwmX2JstkDdc/03H86NU5qfF02FVTnl0s0Of9S9fVC9zmXGnx
ZxprZ7pDG2dTKRguCjEZbHWAg7KE7EnxLGEI0C8OgY6tarm8jRdtxb9yfz7V3GNJZgwPuIjOWiRI
alC7IcDk/nY3WLUgo3VHAjttblZ2Qsf5M/Zo3OAaAOwtjCA3qKfhtOR2Lnvdbot4QX7zo4GTKPoY
lPg7gvtSYjq/YR+9rqEN746WHwu/A7hmIJbq72fWdw3ThWcf5vUhe7VX7CNGsYi56PBIvpGWFvAB
HkSd3U3ubAdBJ/IWz93j+WVUzrQC4zi2t6cb6+YctNQMNpg5tG7q1Kh02FJ0pdqcIpHgsgdfTRBS
KW0UcwjyXbDxRdQWpsTOe3B9mT3fQOOU9+WwzniGCOQxqrTr+exOn+HrcbP1bMtAvuiYjVbFvw0Y
sdEZCBSfgzrskyqyopqYNRdsRcOGbE95jKuTemBApmd91Qf4uRKwcSXAkwZGrqhXrjP5pT9hY7lF
PWlyfCQOzCZAOWbPpUeouTDiB0WcaS1HIjO4GJDecEs+eIDkBtoA4czhd3JW9/gm5r6U08bcucbs
yXRrXABMDvBUBTULQ/egCJ6U/QdLUO2ngiZeApIK/l//vjDWn41Z1AG8d6FaXAA5I6DWp5Mv4jy0
rsmKORLkJ900uLhWwtCl5bAbIXCg8xWm/06HhAvCUrV1x50WT8GWHMdo4t53pSZEPJ3A+6lSE/dt
hp9utF3/WrxDw3Z/rh3hMVhFY/1J7OvUnYhNnzQNww8/fhY9i4zyMVQzrrXVNU71Relsj+7rM1I/
H/NAOP2bEAvjyERpGJvIuYUpN9CjD0yo1iG5rMrQCIXuatlYIWkzjnti4oC2uOdXifj9zXYMBqeW
thqEJ5W86jH86QDh5arKt1EUbGQgK7148Uv7EZGHYdwT/E6rP3nW30JP/d1Dsmq3Tt78zN4zGabK
vMfJXcfjlcC6bEa3QPy8WJu0xi3lULF/Az5KTevirH/1rG9DhbzuNbCX1ZMAhhqOtjLeZr0TQE+B
7Zp5/MsfZeRFDZbGoIKrrG8h1GHG3Nhu9XrzH8WpT6fw8DYdPfCZZT0bXeZDOhDojnvejQmNe6Aj
YZxFGt3qmbtYc0ifcN99q2rEXreSR3qRjNpSvLsjs0NeXc9fBhWEi4jrDlNreO9Xst0U1jxF1JqS
0d3mviSrbR/O7N0keYKfzHPsogsf9iJ/nxzdrAm1SQsQ5Tsqnt1zpMW2oNN0ADZ3tqYvBHWJvMvA
a/I3EZgywa39uK867dHWx8piKRJGOPjXFotAeV3SiwXHiCrMcJzuyZMytleTZ+wWck4jWV9mAsGa
IBsDhAS04Qo1sdXS9Oh340Sr7FlO1eaIZ9PaGKYUTb0b0YJWpl/dMx/uk1MlWXXAqAiayexNijGI
6OuHc91ek7F87TFo88g/ptXcoCa4TyJRpcBTVVkXaa9V7mHKWierIb0Q8i8IY+tQQaXnbzwAoR7j
gWRpszOJ0Egr4+/kPFJLPYNoRMcXPHfv30XrssauFo2qfpPcdBAjoq7QAhm591gROlLxU+0K1+UJ
JGSYNRiWIJ3VEkriu5wZFUpXpW6joO2t9X2AbTHdVmEUMwwQtQCIYSRiy6ZDfBWclwkrR+LvgSAO
xI+qWeebPreDQDKDDTSZKZ/ooYWOopdbEZh8irEfEZM8gAlJkvhvLIHc4GXmhNV2dGKWn1gMu5vt
eZ7iPsBPpr/vm3aWG9xpAm3frElHiuzbnPJOgEJ2Pf3uMj0FNYNgc7hkiMGWPTA0GhvVmYe24YIT
lAmT0Dg7N/QpnslIlM7QU4PNwNOULifKlPTBD87D6OAmlTe5J3gh5m6gnnBsiGT4dz0/iNTNvTJW
icZ56MTqQj4kbpRu67G0Hns+YiTEu/NIv8+lILP+qwHHbLIzwyxOwYIkcWEAMg6rLYiNRzfLXYEz
MnK83iSDu+sMcHwOK8LdHnamN1j2ogdWgfAOh0LTUL88Gi47/Tlm5W22gPhUoSjxylq3wtfm+I3y
oKAil4xUqEjuHYSYH2TQ/dnlVCqF2Mln1nnFuwXsujimZVW+96Gc4hGA1lIu/qXTx+73mefkEtgo
8n318JRSV7d3Dd1I3YqUEK/Qo17JooPqMS0p84EVf7U2eHqbg4KGTekNeuxc12oQxbM6zVDIvCH4
XqMo9McRRgVDFCGVHnHzj2E6UGth0MYalJTwguFd2kxKLuhA+oqriWhuBwFVJ1IRwpvpi4VS34IE
zh/4RPB4KHUASS6DzMzvsFxRPAd/EYSQd8l/xrLK/oUOfhn2IkR4geffGP1/hoYh0yFPiOwqbpHA
1pgyzAuEMsPedD887g30z5bcezAMaRWqXXlxj8SqxNhklRvFOdM7I23j9F4GCiRfMsFeVT7rnYLj
BUcX+9wYpcNNm11pIY5iXUgOIYSMDt41QjlyYJWHEyaK9iLUcfeaXr/hfa9aTrgsoebI6oADnd5g
Pcm3ghlg+OhR70mjVJRaH4nuK+58viczuDj2IU2i+v5ulR40NNivoGYjLE3o0annNBPlsewpi987
jEyTATcCLMr5PHTvPiykHDpI755aLZmNRrZzyKC59mulxgpuriNQu3YEBQXTdRbC3CmMm8y9bo8b
DBiPRbG6/mNguSJPrH0faEjA58i/G7GwvE+vVdt+gAyd7TCO6d3OUdFGOi4Qe0jApOFID+B+Xvha
K5Inah3LrnO5mLreouBcBFjRU6lUDuWHNDzzedkI4hV3n/xvrsQThPdaqP3HREkf1kH3uAlNGDv5
PjIHLKOG04PM/j4ZdQ14dJwrj4PLUw2dh9tYuQ7vjcnosKHnQb+nofNgSV9KiuNtNMdrsYsojw62
QJJzMDuYgWkg0ppfPRJ/eFVR5Q9T9l069GSJH92Nt0AdC0XWi5w48Anm4xUFNJTG/xzbZWin7jPd
X2XkAnVPb2mt4dFt4eLvEjFydzLEXS9sKoZruP878leZPKBskecLQdGGzUf3vNdQYbQ4bVClIYHb
gCRBkMukuWaKZlXCUM+WKejTPK2JoMlqVNzgyveNqbF4eDxcph8/94h1Sc6GJWIVvyMFidlYZNBO
86R9Dltpc/SrrAn9UsYGYNyV9y3jqwbE5F+Oh/VjvEPcHWxGex1fGMgRpLpqN6boDfhTlrS2FpEN
SHzKGnpXI+bnydzEAdvv6ilV8EM9+dId2YrJEH/sTzDLJUQDPLoQcqYP/Wot1b3jZj9L2shd0vXb
O5Xs19u4Uqxtt6738XN34lc1WIzGl9DrEg5dj8cvd+9QdjVlPDAa+EdwczBgBhfWEektlJOx6XVE
QxyED6mOSZqBcJy4fv0Ny3scgTvjE3+0zCWKe7MZy12lf/jbU8ADNcrVUJzX4VsWUFSN9j876k+j
D7Fq3OC/8+O99r25kU/faEY1ERI4RJy6tjS9OBnmwh8ZGT09r74nbsjo2Y5qnOcZV1YR1ki8NYaJ
j8xZKxb2J7F9ldN3dW5N7sYMmuCkqZM6VZxsCb3wwbPFK6u7CZ7+/TL4+efriISR7VTiOdKM9SS9
iF18UfCc8iKpsVSDZMxSQFtvQEJnWhCLaGpWLG4/fWCdZKQYPGON3AJEO1qggoRmYS4BVhAhJzSc
qwRXY71hlvIFwRFj1iBFuKuD1oM1EC/j0mLX6unCoevWlp48MI9Nn/jHxOUZNcat8VODJhzl42uH
WY37LS2ORzLXAk7tMwSj4vUndCDSWVKot4bGMf97b6OZeUF2foUzsOP2LahpYcfMomAMbHXeF8ds
GQ0BynNrQcsQ06ki3f/X4Qx4QE9HB/OQfwq1yuy2y48NYuSfMR/ZYwfzszH6XojRuDrLC8RCORw5
Y1iOdWjR9ptd8QfQtCjpbu/BLWvHkHn89RpdAaTv73rvkj3J788KhPtSBJKfEj+HmGABIz8kS6CO
lLicjdOTc36gwF6sMoskpz7l8P+j/+qx5j+rLwZPuRyUJYQiJGmb2xk2/bIDRkCOIenN7bDULHgj
FckRaEpFkeeDnLHwtIAaKDjD56Wo5pn1SLxdGhFO2kDbv4BVJVfSmTalFrzvzUKtu7SUVlLqQMXU
EvHWp8ntZE+VnBgsMtEZJkStwg50+uBqWc7cFpZ1gXtokgbwQQpCl+zUwKiAc8hywh21vc3WtPBq
yBilbzCFHrY+oVIOkKe+q7/Ax5dTLc9ntrlU2YpeTAxW6Bt6WbBwgAyaKXM7HYMTw/j1Mnd9iosE
2OA5tZ7wJUROMjV/7H0t/PJZumD1319h7k+m0kN8PGrw1Eem7tENgT74v5v2sLjLzLkJ8UesusRK
5+k+wGI0ZV8xDGLtHlVWT7tm3/FBEKUKpYw8BzZHWJ2rJugltg4biMH1oshQVXcN68LqsfqjzBSg
tUzcMyNtQIiazfV0LreZV2HBVrccng6ZZJH1EioEb5xNZzOF5Vcelm2idrmslk/jJc4IHWCxPWQm
MSTKFPlyywcobbzOnXo/WjyTt3Xy53CpXbJS/vnPZzxxNlUjnyTR5tsgYbsPbgvah0VMJytcAqPR
eLJ08DVLLnlgDruGMQsMT4ptgUGh0riq2sYl4s06l4tXp28Ld3sEqGqVImUMRFMV8wN1KF2EvDxT
5rxgVFBw8kOqOMdIO24ZWa34KFAXVWaBFxQ40aeLXH8OzwReXcjxWFcRT0j+42ET3WTV2ZYolto/
G3DtLBYC1+p+6yTg/fax38O1/Q7OZGKlOB4DXCIFQh3/29kVwnZ70eIafntKcBQrBZkfn4kevAus
yiEbiKug8TjXnikzANUKj4yGgXP0AkaO3MHlxwIX+BVsqa2do/MJkGBpJq8h37LBvzXRXxcjezHw
qTcu0qC22gQvbxUbRlfnNgYUegpEqMGbdiK0kx9M3SbevHDfcY5rzbikZ8r70LsI+iYym6ije/OR
/4Gao27eXUGmV9Cu5p4zAZ8R6X0vY4nV3f/LXDZRcsAhZJUTNcqSOxx9VWlOme5jciZTTB+Hmwu9
qvoSI5Kwmx+qeml1lLu18uh3TMSybI7/FYPQH03v7yQH6SqyW1WoEqZYnY0YDgth4tdTiIJE0ufZ
YV4hNRi09Djj8nEMFVHLpuYUU+qZKnqILuzbF1MnIsOyCZvReCsDOLPjcgV/C6rVO1iTZa6FUk1h
2rabYRYL8ypV9UdyyFmoaT8pChFuTZl1Qw2y+yTW1+o7rKuZXMS/I+v5+JPhIeGg8jgZ9muPMEtS
+bmh50ZluJEt2piKvcPn6AOAio21AOSP4tq+9FYK5LfGQnsFz4/vothq/9my4q7E13LNwl2M5VRR
cJla5AK38C3hnoRc7FT2754qbVApNxeC5EqKUgl7iiLoEzJAikihaMsv57spKXzgGHcObyYXPmiU
/89kfQqVl2wevNG1mZoFUSwtCQ2QdNXIiu5EwrVyqBft0PAxOy6s94qKlpHqmcIxA3QbQSc19r+y
JWjexS+SvfbzDMkKhHdv5OfmBM70JvyR/vMw22/ho4v9aSNo4z427xU8QBEu0bdcCsrLQTZeVd/h
ujMp11IT4Mj/8/9O4RgomCOmGfLrqqpvxNp5xj2lBCPgz+xmpARmSXG2/LXHkmvGu+nNN9ze+Ucd
blj6YnWm+RZNTfP/s9Kw7+aaLEWBuGWmZMmiRQaekaEQDTrRBeZsJOF5EzRzsbGmTwtX3oDoY6uz
rZ1PIzzDTSkWqKMN3ir7EjE9W0gVPakc17qz/XWMb1WKXj+5P9zTfQgEPO47Y5zasqlzVvmPmhDs
djHMvIZiJVQY/8+jPMvmzfVCvR/syKUNLw7xO6uGHf7s0xi64P7ZNolJIrPcOaVhUQtbR2KvTvh4
2swjqLtdUjOJfoYSEv9GLusZeY1YFW4j7WNPBnOGqiB23nRJ6R7rJAbcKDYTzlkyIvIlSTx3LM7j
O55ZMIpVo+Sqq7zRcND3TxAqylRMlGlaRk0mDy8k8YgR8RoryJqWKf55yoa32nZnGLn57xsN2/+J
uU2R+FkcZONDGZlaP3Soap5cNMTOSql5VcB86OUS4A2Fb+/URUw6A4EHPaGoskb1ZLFNSdkgRceK
HZuG+3X2k20M/xbKpqpMrVeJ9HyUFPaKal/MrER/nWb0IN3OtVo2v/pK2nnYzZzs1nAeYZbrCmee
30xNW78iJPIMto8V4nBO7a6yP1/AVe3HD3TBCiERrhTzg0P70F0sSm86hzBgF/lU8hQFyCZfZUTL
w5b+hdiudcsK8vETSCklqbnxnv+vGFqXGgejp5g+p3UsW49+vj4cQMEHJ9/5myP6HOcGX4Pu/n2t
jBEn7dIcnU7diTc4h7753ndLte405lFgq7t2CBJwMdg50mw5Ei0DF61wXfKiLIV5jW5E/zSSQpKW
ViyFGESjxsLNPGOKXPzT8pkLdaNXB6H8tDH+yua9HxM0TltaLbIJjNBiZ5wxNI6lQEXN2LBg6SOj
ogMRCuucR1RimVBFl7l/da0/NuC+fmTAYn5WXCegwMVug/QiSLA/Wt04RrNeMypvOGhMqcP0EAIs
p/uHxbItPGVIRvrQSvKuhWg4Z0+x/38+iCFQzzWPcfRTDI3Ow7kzEuvU35UpAFRneCv1nknkaKkH
wLHmXnKbIB357K3XzMVgeXQNibrfKZJFxSL8SWUPjGIua3PQwxPeuki6up+fQsGGMv5KKrynmZTR
bQeoIjmbi8WopAQx3XOq3yJE8dhvlNa77NfZxxvfajNyPGJcUEdvCUOspDFI+anRoY/Lkq0jOigY
NCF3U+uHpAHKPPmDhdFTdkrRBKoA/kXewpG/43mBe1hprIhO1vT/JbiS124eJ0Q4jIyju/Y2MuOS
D96wQHqFEV6QIpofsLJbvU5+LpBUnL/rU450CEkGOMeiGnfrYsA0MmRIZzMLbCEMgMFqw5DYbMWK
FdFLWlLrBthG57WACiwg6bjdN4PsF6ZVo/vMA804vizGqdlKmNY8vc9ka2uhMpJzqkA+DUagNgAQ
LW9GeB2cD9M+d9nYcmS+ygWlkzsz35BnqovZrVaDHiUP/mLhhOrwDQIDKLIiC6Q/wjZHRMIFvNZ6
LxlkjS7zEvqJbm8rrMPoSeT+CpsXXFRRbDBhjq+0cUh/EWlMhcBGpMlNC8rLVKfFmwaB3PNb87I2
FlONuxTQ0CkdyFCJcbOqKhab+H1EbsFaaGjUomsyWYVPAIhfMUbas5jNyoIneoj2YfnSX9wpjSWF
JOuc0R2SdP5xp8LIH63t9jxNpS318T1ZVBRy8cUIPI5pTD9lnNeAoBi5LyX59lqdgckBoTMwE2/Z
l/glSsYI3EtZaAghBVSdbXcqwiMMlpyi6sA9swQLzrkiTijAdypXJT0rtKdQfqMnTI8LMq16yRSB
ufDB1lc9HpexRJMaitWgTPjdbPR0OnbU583gmXcLUKkBkGTD1ynFpgEtdgSSHPzfrYVUDmZfVWil
uZrCo78Yrv4H+2j3jA8JJKeu9Eex8zq9ZaCJagAEcqEN4PbnJPBHxZ/JEdtDlrgOwSOAuTqSP182
b7nIpVLHN7B7eOOKe3JT3U7sseQTkO3z8STdwD77UndD5qJjxh1JaCnW1svKgs82nqqjYAkJqmZo
PgvaUyvqcazgcXJeS+s4opFD3dk8h7/T8KX7qLMr7RSBy8UkoLbay+6oanoE1bGSVJEJmJc3lZ7W
WwJsogEPK62b5zBNoLiPGvB4VB6/u//gbC3UNuYZPYBdJbvY2+y3WlABMxu2kWl3nUB+oiLIszac
ZmYkUqBIaWX1x9iYFpmK4nHjVxLwYLw8OIe8wwXau8Rl9R5mIL6VVJn95a0QJj1/3MAvOlQcMpED
QzZx/xER/dm+9ppE+E3WScy2WS9iDCP42EsrEurRNIA3Dl4WGCSET1mSwda8Swa+tPakgRcjXgDp
xhnhREqqdtMThENHAL54CT0nUZvNV5bCyOIRwc6Gaq/dLPePQzfDl99dn+CAOkTZDFBMaTUJY7M0
vPWFtlhL5u7ZMQmLCXsKOinLfclN3o/luQKMBXagLlv81pdIsp1R32BH62ZKfg+s/XytuLmjt3Xg
vNG2LYDwAuyJdF/VR6/M/gUTC03je0wFj+z3TKsvUDJfJ25QsjiijtRBdCAbIRXaj83yUijXQwVR
Epk/fFZ0wOy2guxXwfF/ajQuT6m1bd5aMmqrqveh66+dpsmyKXIrpF+b1/1t1k1L4qgWW/E8pQfO
jCpPMVtuseKVGGvyv+ptScd5u/Yv6gJnHNP1uMSzJPuaT8PoBFMaAQWR/Ffhl6njD4k6vgIHYrCI
dUIA9OCA4jQ9Td27Kd17bmlPXSyPCM5YMJAlH/uqW0aKb7b88y4OUttvtnKoGdsz1dXvj6LTs9y+
xdITGIo0kJ89UY3kefuwIGRihrmOvGxXRu1dYxKYZ4XP0LmehmB7ck4kJ0jMirsIGDephOq478tj
3QoHBaZAZ2tSz3DaHSyJcoARyJbsMDyUAs21Fak3Ttwaq4W0D02QERYA8eT4srRODnx1fF5bNSKD
5mm5dPXlMc/a77sPKMMZJlDj3+0m6bFaioG9fYXJQT77gpZHb9QJJ7a+2URI16sXeFk3XlSNhBWM
66rv1ufgzS8/Pwx0Nu1FjS/W+dBH8L+VqNPExvMbQupLHhvDZRiSI/QF2QPuU5qohtPx2NkMCIUd
JxsKwlklpRBKf7I60sKpvtHo1jUtzWp/4vd1ViiM85jxphRqYPiaQpl72BvYB8CIjGPVEdM57Yqr
wwSeQna5DhkwhRr/OX+ZEU6ovr0ghjbzgaN60MU22MK+98umXQbZOqK9uQ+XjcJYiHtmh9XT06c+
Q2YYP0pYEBcJJUmjoegAt8uY4TGxot0cVxGhLdTC66so4ldIMo/psy/sZpHfXsLPoPaqX26fhHQV
CwRY89izx/9kDiQ1HVpFVoxjHHxbUHWhwGLQ4aOciq8vlhpaWBxTHAibnx1A6ue7jYXAmGdbSUJH
KiQM5diePaeexSJq+DjcsYJ2Pjxp2LYBF//cjC+3OdwjIGj302JN7YYX/QMDTyKxk4EYJvned7Nu
PTg3vJGjAr/cnntbn+QzZmMGnbbChUXIZTYzKMSqFhHWLvdonf7Clu6a43+tQUk1F3Jc5+nc1duz
nirxSGjfInMnf4AEQa+/4B4ALmo2M0EjfUq4yfA8lPCwpdaNgzJomIwmi2JiFjgeMz2Wo8jkyWBf
uTWV3B8FR6ln8ZxuXvnR+cKVqXuDef268vJksvzYxqz+JlTpGKibcZ7EE2OUt2/aMoCc05IItPam
Ihzbi8w/hW1681ey17LyBpUTNopcc0nZl5O9Zm5mG7SGhPqnPXkBNYzWOT3NF32yXTOXzA4BbUiX
gQG1wiFP+55j6O/Jam+bX4b/TX9DhoufsDXbbGo23wk+s9bHe9icgNx8FbYpvvG0+LnYmPaEInru
+1PNztXVMQpQ6cUg5QH39JhXgr3Azfd/D/xs56yt++AUHbhkpE7QNwrBCiTt8e00B1BjB1Bm1eA0
BE1GXRqJCJBSEyML1klS0MlehSbIqGS+I2NxSCOCXWtU9JxFy5QC1ieVfznnR9w+OYSSPryTHcts
moarxVzeH8VsCaa2PinkafGjj99nsTShhdvMSfWMElq3Aew24JAdV8QjQQlAzUtdt1va3zGsM6GN
oJdYWFwkEcpV0aqNcw63cXwnaProJbqwL2DAA8a/gsFPGm8icYIhK1UbS/aUfUPD55Sz3bsDDVd2
0xTWIuiouqr4CmDrNFCc9h6V+bFDr6ItvCwDZJ3bJk1SK2S8LcqUAw49Uw8lbxdo8gUILC1ivEpY
X6MuZG7MpHzJB6S7p7yv8U/MHUE6wgr4eImxEj3hC6WO6KqFV2H7MNjDwtJI30iJBi2jtkvFTo4t
EQXDi6WHyTh0hsOzWu4jgC272AwBH4alH/VGDml04tTycrU7yohuShkaMdm8vZpb763nYewHD4JD
TrYvf2uKDG420adiWv5m+C1Z5oGNTSx0w+wE90xbf+cmGQrXlLnmfFNPBK5bnI0Db9X7hoBXopUG
AJJZAG54f3MbZZnfH5h3fL6e1WYMxTM3xg9RlUoq8L0E6e8d66BW4q2MfzjrVRVR3LUsxk9P+6Y4
2+45GWnmJMmWdLAO/RYfN/svwrj+LzXfGpGjOoh5oX2ELvyoR8C2TwEmJSWXekbORe9KHcNh3omA
Z3jGDwMKzeqnPRhh5jpULgSGwwZbt4p0e4/gagEzvE7qNv3Bl3CcTypFxo2MQJj6YWM0XnVL6FLQ
wdIgO9rRWKYzqkm+bo/2ATiLtUI2iS+lu6ALx2CQe6ztKFt+JBcFyh4xaIMTM9j48uMtsKDFfbu6
uwd9PfJGMxUdILrdC3hf/cqUQkI1Ih23ng0qBpRfE9j/+UB1KXOm2rqtibZFtY80wBvKuPYbIkCI
Kj8HYdeQfZwHIs3d6YPphnC5cvSUmxsnkHJfsCCeqwBnioIMKHKF5Co6fjA2LTF87xuxeSAtRHA0
X3ZBz8KdLZQmxR5rT43f4lz0crFnbAuGFlpvcHVsxx3uwARLrCTkVeFc4K1gQ1CydeRHfTAD0W9c
DQ3tli/zILYL6szxyfnZajcLo+FBqj3ToSgDBm6B98ts2TqR+uNL9Z8MI6f1Pm66dsOOtLhz/VaK
2WnqLtrel9qvPijcVkXEklmDNwsWqv+ewdvDnKGXkkkYcWgdaeEq2ncrgNM+u1iUJpeskzvF6Df8
oX4dvY6UIdcfY4YP0PBZYbs5KjxWC7bacDNqNRowlNqKCuHFGv1+monMZ34InfhwWDVF7hqrXBY3
WziHbLPYBNu+bZm/5Cm+c8TMl1ggbkAgGnmRIBJzmbHsysZUSI313M47tsL+tJHS5x0qMd3oP11S
b9RKJx1kwgM7wPzfuh8k2htFAdZ/Rd/gxlD1HNgvv/BaN70iqGPIYFH0fXEoFxpYY1eRKO5vBVq4
3mz3n/FLpMV0bYuuTxwg4Vfby1bb5+kwkyZAUHHhq7gkt8hXJilKfQS/RnY61/XZ1wrhvfmNlCNc
47YlgylpSbxIDXXHYHxAEaofcslfq2rqfZrma0AEZr85sUN36KGOhRRkgGwZbSplbkQUN0fOoDvf
hYqhL0EiUvjKhikh4G+oYlTbO2AZ4LMgPr2Pcw9S97KzVClJY9R63ABMT4TzQ0D5YmkanILBy2Rc
tvLEzhwhuBIIpJfjN+R+qI398K0YKT1HuCf9Dir0G1TY31eremDI0Tf7+QdaD0fbRc4CyYtqGy73
ijAojdnmz5gv1V2enxRgo76T+KFGY0WTezPjcK0UCz5plr5gpnK4BpLoTYp/WlnKwQTC7Wy1osZE
AVsthzGu5V08gk4wgTuArHXhWvwgQ75pkf/35NwcJgZSUfasxB/A9WGztBAWAWG3AAUWXqo6AcRB
lKUekjGqXV61Fh2MKVD5aUopct9PZ4aZI1sfrx4X7iybHnCkvq6q+1MHN/AdsSgrYRxS+IxK7bIr
Ev8fvBkfxn1yZMtZCffDNSxa4arB66jJbKY415pXZA9dlZv8mDKlxbIvszzmG/9iMthoEVcF37Nb
2IXrKC/pWJmGSCty9GoNlemruXJCzgSc3opqrdtxP8Ps7fgxA949+hqQagoKdbVsHqE5Lr2H20/v
tEZV0fLNqv0Vqmd2CZqwTPbnATjXm3D+u0bmjmjIVpv/7QdIU/GmW92WchQIGUY0mxWDIqtJeTwK
BF5CDALFRHhO4EHI43MdApMMWyxH5lYdVE1KwyPP/SqEX/PAZSlMklsJgh/EFtSTmz2PFIFmLvS/
w+ig9r1efy+8guDK01GThDOYUpTOGono1iMb1HIBKUK64dbkFjettdk7XOWaVyjEud1wtkxaDG3g
bHJNuYV7aWCubF/JUevAIhF5R9sWsHJ86/lRIbfnhuIz+d5cSIuHttbYUqgi2HofZlwwQw2/O5En
0Erk0QhL9LbCQq+y9D7eBXYIzSQn61+YsfB4988C6out2+befOdGARJmDuiCZsLQfnTpRGt6KfnU
+JMOAZHcSlxcNuap51birqj9h/WNyN4j8KkN3CtzBJMd1310260wfEB7pDDvSKqN0J0wLE1eAiOX
7fHYM24RT8V8nXxvxzoM2B0DFbBlLZLsyW0hyE3sk4C3i/CtV9ICxboburghcZ5VJUAo8SAvzei7
0Eiq/KR0xc93sJROAIaeUUHFbUbbHbYz3LgzjpVVPzvPdImoE8xxTMejrhE9wkz0M6rGjFBLW7cM
BYEq0s5LRjTZWWUIAuI1BgI7HmOuMe5WOfzA9lcWCm3Yj3N7R3XEdpo2ztEs2bPy7pptxr3oveeF
/95DrUjI2cQ1MjUpSbeCxnv8OzQchNR5bKEcTu+gsTW1CBhOUWAG6JfbGKDfbHrXNh7qOxfA4IZx
3UWUqq4Y+AXOC3mAEBERw18xxzEXaRbuCpscHN/vSgESihwb/vZdNl1NQt9Y5D2hY4u1Ej36Zlsj
5cWZjntj0iI/yHdnAuIx08HwHT9Xgf4++2R3W/6Y92gzzSnI824bAYYM7BIMUBFFsy9aNx/fe+XX
aok/+gQyLXYs/BefM51DPPjKh7ZtiouWfGQQDRukRhuzsawfnocRgZjg1KiV+WKyj4NQxIYjdv6h
h8H2WHN4eXYDRNDadggsCI9PAUYMD9h9cBSNY/LO0CIgIdSJvbwgfCdFOxXgfMa/FNndI6XjVzgh
Hvvo31EA0S8LYD5zy4VRa4DWGMieqkXLeHQz4eYNaKQ3vBgUVfjE1qCEuRAXXLLKe9tEt1/GA2G1
p7WgtjPT+kNXUfnuk1AldttO1J01wsL8WgXfDxGPg4G2ucbnVBni4yNGmGzqEeeSKtOwZKK91Ah6
vzMNcLZFo1f1yZslzIYsG3LW3wqAQqO/54K74wUvyK+G+poHXVUcJI3DMmSd8cJYB2akN6cvWAMZ
3BbOwyu8OU4FEf6mWVcV/AJ3nFdWsLQGISGkYjoSDAeijU/z8fwI5QZtlya27bJ1lT7eOQxycZoJ
FRK8F0JUmFU3PaDSuQ+Bm+XvvOTNhVojzVGK2piMUzp/U+4ubYrVdmTRUwDBVvtuDAG+ghIdDXzs
0rBubQ3GY4rZ8hyxzwx3vlXrd0z7aDfIgVQZGqud9DiX0R++wxxRL9ucOWndeAiL1Gx/3qRNEPnD
2YYWch7S2LWMVRbD8nK8cKZHQv0c4eEhMbYQM5Ye2wk8Uja/PoPa/DhyVF6IB1K+DaNBHQa6sUdj
WBtUGKUUXH2ZiD7q9vDwNNN6paJzxTd4ivK3nTgtJoq/RvIjBN62ZlowwOrXt1DKekO3m1yB+Gjh
/Fya9EAAwx1TT/xGvsVl403Q2DulaCm27sFjHD6tHBvMbr1RjaCOvv9gm8Ube83IP4t+fRXwqqaj
mOx3/SrG+I7T0JqBTfGZ40liEzFUcM2u2qbF1a+wEkmp4ocCes1RnSXx0Lebu9gC+/J3ieR6NYuw
NsaWZl11ZH+KiJ+DJ0Bt6pumHlWIKEzugj1VJ1W1aOB+RpztRi7YlPiCGwfVVKv2Rpkg7osRe3O2
9MLV+Pt2UpXGsMIA3XtLDDMQqoAcv9/3BPWP0WdLwJ/DdogRlyATh4Pcm9agW6EU2Bqut6QB4F94
FR9Mm0LqU7DCkYGUT93M9j7OWf6+84RJINUqQVxmddFxYmz5d1gE9OHFios9wvRPI/KSt0lciR9R
0VA05ITkKhI2H00fwmf0x00+HHFPFyXHrL8ujEhUzzUcSwbZvDobfVQ6NsggPTgLl2atroOHwEHC
55XAz2dvfLS8nwAGkfxI3xgPGYQBQSBPg+WOppC1BiTrKFRJSSxsx6u70psSNZiqyS5RWwAoXwJN
kcWXTm9qhn3AN/iYvUuG7qOO6gW8QgzXXpes7VKbNm3kCguIS86/0R9QUEYWJNKZ74/Y1Uua6VMt
shoNG8hGilMj8R1SSGUlG4+gdYpm1mS66WMZJkrGk0lvhMub24Zg5VLUe4r80bH93yZta434XcBV
Ryp6jKvoTewoDL/UDwkDtG2U2wEwha7J55PWuEIzLWfbi/tzW/9e9lkK+beduNFd9Mof8Upy3q4W
buy2AyMIvNpFP1iwINi+5XozjEaAYstkTlYOUaztHjYubq8OqKyjjmV05P+ei8M8hkgEbFhwHQX/
kyMFNG/+h5sAzkQOy5qOY6Vu2tWJlhdfg/Wo/fQdMbKPjtrwsPNAD98JD13OHD74SWyV91udmMd+
zQnm/dbtrYPYtn9eIRUYPPU/M1HKfU3MveiwNfz0JATewQPa5tgYho6KWo4CAf3EBPxdFN9suYDg
vJs+WrTpxpVTLwP6YqEqBgCH7Vg6WH5uI7QGLtFJrL2zAmNvx29blPd83c/dMaJE7pvmzo10fZmY
CeEQAccV97ocbLMAYOpDwizNL5It4EeTmgnDPpGRJ2xMSXQVGre8/KXYctVLb5Hs7fc0Mcftzp3R
V4fEBP/vPO41Ys7MdBM+eTyPTYI787cuo3jzfj6wIV112Vv3CkOpziiTLC4S0kRVOoHtYGFDtHkJ
iWaR2XGu0tpwQP9uZYnl+WjYWIuXGXJR3VYnLHogab0yUTUl0NtkYoIDK8Kmenb7rzmYvCrFQ0r+
L5P7uB5ImWS0f2eYxcmQmJVdRDq1LLWlWp4uTt8dP0HgVlNjwJ+AOz4K1EPJ4CQbRFPMeoZsn9r5
8CQ5R8hKv7tvjpgxMS0GwKkC5579aIHisLhP2/DvjOsmGCrPpYYZwW9nUtskTnDilmKvAkuyJVTI
W7dc3nlSMLr0gyevhMIziPP4WXtFr/ToGonGGuBcGUbPsOJ/9kegDp9AYYfGpvON5Nzk+xA/IwuC
htps6t9u+erEIqSTZatI6MZ8bP31jL46tiHkAkS03cBGf1yamYUaL2deXTMJRgPdgm+9cw4qpBCP
o+6EH1ctgfSXI53l6j6kyWg2wwa6c7+/Bb+7t0tFFg+7fr/ZtO4ypPPJ8W8wCIac/SpUDVG/LCQI
I9Nrrxnc1fUquryFi9FpoUCA0aB/CZBpNJN1EhHO4+oYFGx+2TFKbRqQf8V4n5Rr6EXONxnSW/Fv
SfQJAbXfws6ePT2I/soc8WDZwlWYeYh0L8mUVeq2dK02TWQlMRfYx2vjCbBZ/W5wLalnfP0mPY2k
jDMURGt8x5kYM0VywaSrVb3zQV+rc1YvYivCFMKuMJHkTM3l0bP5AlQ+OhsrBR1tqsvtdA5rcnyC
RfNaxhPgYspJ4rDK/bhZjYzXOJFj//wVVuT+JdCdhb9QkIEzes88PD/WVS3CabvUC25YF8cIcjUl
0c36ytmmpbxGHtz3cTI50w15zVFSk5wqwMr6eBdD8xOY3TB7IoTEI5cSQ77HTtKikjPRYT8ZVdaT
N2MPIXY8N5AjfCdMD+c32pWoeTB9kV7zshiJ6QU4QjEylmwIylTIGb9BrgkLxaLA9A6OSWbkzvpY
AyCytARTdUnqHrmhYeY47kNHvXd+uZG9CGh4pUANLAKXe3DJ3aNVWZyX0zRXlie0hny1xOLevoR5
0CfnrN9s47uegE++a35Yi5G9b2Mtpz575Wv2Txz9abBA9lnE5T93CfIYBX4OHapv0+E3E0ylCXtA
9ofUmL7qmX9OPnGCIrAjM2JJmmSJFr7X2+5GTYsk2u43rt38pYgt1je5VeiQkvP6s0mrWwUqx9lf
jdbV3iHgPpPHpW69enSMSlRsvn0UqvdWdOa36f7lD2NEP3clIHcQmDNL+ZPm3eeozGqIlMQsVb8d
19W5yg93twZgPaekTWC6TUp5q6EF2B+Hm45ZoaHzDi151ifJa1XuiQJWueYI5JN9B2KELj/sjyTs
ZW6wilm+gsQTXqoojLp4ZbObSPCD0nJfVPQVUp3+O9W84wOdOEwhZ5amvmXxIHlS0wHUHSDMPoqY
KPjXCdX5jmVpMmdgv32WwZGCaehi0sjVmu1hlXF3b0GEUZAvxxlx3UNt+S3LlO1VEMJ13EL/w7pk
8rCVahP6JUJ+W0zHWmTSV3LeOLKuTnPuv++ss7vEllL3JqkBSa6guj6vCVeLQk8sGSIRoeUCp2lG
1rmbvYAdi/q1SFz4qcwBOWq4Owl5yGEYCY2tRplDkzSFirA9Nc0X0bs35eIHOlB0Oaa9LxJYvxBi
kffXj6bPZsbgrvTF9N6Oo7kM8d1XylxQ6ZkjoPFeNbQjj1trqVVjad8Tq7Q4vgOHAmvW0zBSG2WU
cSn2UPBmZZyEtNvDlh10L83lzKsFRvAZJd4kfqeWrYsOP/lpU/TdujbWOXJPQhKe4mpC8onY0gNY
PoUrnaqatiQG6gRj0FlYZGrVcwoIcRKFGh8KlH0cy0kXKMF0hJs7lLHoPPS8Okm8QwjwzqnFe+0a
DLdIhQWPHe4Mv0Bhx5xLcXevs9J/SEs96KIRN7o79IrniLTTrtAL9t5fbTuje3DK+6SOdOnyi3fj
qXuEcwT9oMcZNuiJb4xbLVuk9ldhU0/pdBDaB5ymtgDOTT8GyPX1vUC1Y+mbD+nvSM8v41VkvMex
DcD32S1o5Q7PLSphrHRCtEjpFvo5Te1peUh/EN7U9+4K0ppxhY1CIb5qV4Vw2oybyjD8jSm1qjeq
dAnvugiKuZb7eZglQX5AmeKQGOJXqSnb9pZh8CjmvQGS7U1MuVMdhJoDs3xDyhLfGdud5veIDCXq
wCxzY8GMsPJSMY/cWoV5OFg0bcYMIwwEmiGsYiR00xa6tHR6pljBYL5usU2LiYtV3fQYnK22y//H
CJf48DIPU6NG+p7TGLzC/dRV1gWgL4l8KdNbVYdjYCuT5pk8s+nF0vIn5/0I1PCN54cfPma2IDR5
k5AwPNSxNPRr+qW0WKoaBl0176/XWu2rNJzB+/+KuAbBrr7G19E8cWwh0p08YAj+as0/4BQKIRx7
OJXvmUL/LfyBGk7Ef5YyUNyLItE/j4/eoSBsm9022XSeteQPest7Za5L/6IdWvlEFuQvQKC+fMOL
Egk6qiBTP3PDEksb/vijw5tmlFC7cGhmbHcjqPA9bxfsqKcsZnT3oBPLk/B9THJerQQ/QuI+lYxA
AZAE7tVjviiAe1qk01TmTiv8E1LJNtitFl8NwJnid2t3PG/+Ae3K29RXxxQBPf3BGgmz26E/8J4A
wMOh8ZCO/M9FqwtL86Gb3v/fh1/0t5MkfEHr0d7EQu7V2nWUrSORW6nt/x2ZtKvxLGirf6RGzF0x
1EprsCjX4XudVEo1d9dvTLplO8FZXIi1SDIBeeI33L2HlPWSr5Y586G2VHnw7/tc7nJ95LaC+U5z
ef28tKw6Y8y9GdVo9lDBzrwNV8A8B7vMg6v9SCSm14Zv1gPtYjSls7R+ozcwfUbDBqmRAl0N8aOj
jE5puNMPi6JOYLfi/A0GuXXGSaEAyHgM4PxKdZ13BnDiLCAKIzHZvwAcu6+L4OW/5WmMufu7K0dA
a87oZDDSxWsjkofPjzWIQv1M2muYv1xea+iFuQKOeUkYcmuglndCBVwQQw+hfkhuj/P/ZXObNOwL
+WS1BDCrPc6QHNvTPERH3ZCw4ibnh6aIBqmj2GsJt8qOu53UpkB7jKZ3DoA7G0a3fO8h1YEbB68X
reyuxgEK8TZVAVUIjeDzgCkpOwPIT35fodUUu4CVV2laWoDP/XN77M7eWiUEsN/RIyewfWibCf5v
cJfzes4TWhPTHA+hOJJwOShAn5Y8ibkgl/K8alNIXOgsJ39W1FAm16Rv/FJm/sDyVsrx/DFyOBeV
ECmVWMCRnewb3xux/XcxNtuX1BKHaW84h/sFCi81Melorm4/N9WZ9UseoO050tyZjjOLG9pfZT2f
0qd/eoT276znWYqQ9z3PWxG3M/NDaxJGmJZ5GfopWtEHH9yaTzcPqgvGdjUNAoNr4NAaTtDYQHj0
dR1onTdRARJQOvkaRCrire/yfZ8NKgPP4SOuK3MXnfEZn8cYyn7Y1nSRuyUY1R8KLhhfKzazcDRq
jtjPy5CzsLoHiGoFGeuZdscDQVtBCAzdd/tkPxbI3Ym4hx1X4yzVWZk3Uas+EI9crMoDBY/r+Z4Q
Ld/qEoYkfDaQyBv4Vqf/6pDd06ZLXF0s2BwKxDH16P2ju61RhA/QdXaHfB1beQKMGDYLxLnnvBaV
qgSbx5uo9lhxehQpm63/fLEsvqKl9snuPO4Zr4zoMltFrzED5x3bmk7PQzv+6UzvZqGev8o5wdz2
aDmrpcZi9plyNB/SdNU+uev/6HfeKs8K2Ir5xKBT3JnIktE11MLDSJzoVMW2kmbYH7UwD1WCzUNw
qXUGMYM+UEQsV3TOrYUHiXtHU6C37z/X2lweSxmfs5oUUOiOTIa/FXmi3Oq6BUCGo1IPpDGjQLdx
qUD0YPTKhusgsx/DXSoFR7PcUhR3Zb1THhfBr6dAk2sj7q7SZhPCwXQWU/KrPfHFmsJhLhodh05v
kRb5oAhYFS1q5byDAEvOyK+QTs7FAcz3GoA9I7kC/skxFmjBbcWR3HSYIbtbx7UTt4VRKpC6H/8f
7QlPGeBYZqYIlvSX1m9rzEOobdAhQyubLOkffe6VPkUB9kTXjbyytocW3+LjR/YfG2WTqbw3A9mS
4u5tlXYoDljzyEw3BUT9+sWe5DjQkYZlMKq241CGOnkhWLetgZwl1wh4rSdB4/ijU53q+5VhUhSk
PYtYfgJIJotq+l61elmYVlyUqYo49dmJ6HysUAeO0WpEmEUQiRsZKJcNRoiDX/rONgCrfjsqR6mi
vBZ2STzTpANZOmSdX2JYduTp6kMIkuz1guhBeZLZrycM0u1rg2N+PDimb5BXOMysCuscYVmbNh6A
VTzLMrUDP7ApEL70nHY31uZ2SbHExBPODBPcmTBXtRzx3ZszJFdMQzX76pONgqIEpM+TGunwBF40
Y3MyJW5KiBiJn8J4gStHJCucy1zbRrTJy8a2ayn6deCgF1Twol2qIchtjFsvgcnItb2yM+6t0g6k
gK2+V4PM1TrsLSza+AWNjMkftZQLUS+lFdxLRmwK4I6G+QbYw93yhbe5pxPWERjVLK/olXzbJ19X
Syk2J+z8VnWExXwbubbURf0/UIs24FNAGbnS6mvLqWzcO8+DTy2BP5SkNHHFvIeBAz6j7FkwEbQB
w6db9ILpUwtKeAaUTBTTq0JzDmhw3ZgKVIdQg5JNkWL1QS3U2zhA4EQVV4ERNbpebSdx1er54y5N
kXVVF6zhT44pG2Zh65xi5KT6jkJTktUVnJ+nfXJl5mGvYi/68aGkxxxIO4xGSbBKwwp4co+GsF98
Sef271TYEE+mFCCmgBoE8hTzw0ccABikENQsm6wa8FfAs60ka4cPzeskJ6fGVRn7qGhQZXnFRCP9
UpouAEr0pC6bHzSe6KD9oy8tFPG7Sgd7lkH7qfhWRtXXRT/hCMLt4Urep7Hg9T9Juge5Hrv60bHV
ciS6GU24mckWLS5msCvvXvrasBa/baZDdtJO4c6PPxPR2+MlN808t3YPOWPQHGPk98MIKFGga8hK
aaWlQ4MzstPaouTadmOoo7kCT/uG1intTuKQNZG+/rwcgtZ3FMyRlZKl7tom56uhFRG7a/X2HXjU
PeV1esfc+bAwmAS2xGXLjvLZ0adbCLb4rwI4MLkEob39VVhu4wMFE19A4xSj/w7jCjTkz06kq+2J
GeiTIKvQFYnjjiG1xnkOXjtx3bpq5dmba2I7+mphHUdz4d/GpUSNVFn4onhUUe92uChp6NIexGTz
f8AnNswjKARREbZOc4kyw5AgvH0ljWRBNDlq+AoWts4tqoXIymHaAbJbRb55ZxtCGnu9bL5rJEQn
p04Th9e8+GrqYAZ9trHtwkS8Ajip+X7LneOua9VaaC+jjccBo9fc6/3jqgTJI7+ZXW945cA4KO7H
AN31D/wT7i9+Z3aQHlhrzw5v26qyXx/JDJwdHsY09mC4guUimIr/2EO57NO75vZL8ln0CyhWK1OC
tuMdb0aLr/MRVBhjAZlevIr/HmM7o+lpE6vRui6XVTETFsQK+lkWYCG2x91pIkA+xX68T2YmhzC2
czr0o6F9bpivBU0gsMFJLYf3OO9fyG3O0ywmHjTByFY12HVgl25QU0UpEsrJgroxaakcwht+gBbj
Mmeu09uC96q759TLEj5iCpvix/zeCXaON4Ior9SwRRriuNQPebn/U4gcy2lfulGltmPq3JjNcUTR
3NCeQAoQwlzHcFY6JYIOip0Q96er3QwWORTzj+yGVEbbvGES1Iy1rTVjHOuOkv38PQW5kaxoHhqY
U2IOYlzVUwLXSLHdPI+rcJmilkPJXQsdAAKvDDmNX3kVK3agkVoWM/YGH1Bd/Oy7z+WiXc/hvFie
ifwSFoJCd4M1AWsblPyl8U6yied2gdZgojZZvl/g5rHi128icTJQgQb/cr4P4sics11G64GDbo8K
bKvcL2Iw/wJebh6ZInnnzeVJGJLPGfXz9+E32mAYLUF1+BPe1UHgCXp2YHiamIyYQHOfr0Z7xx9v
jmDry49Zne4eHvkqyX+EhSJRNv2OdTmrBTjxj52PS9gEnv03c71ZKjqGn7H3hNPR8GjUom5kOHFE
VNBdstiiLviRejgdaFTnXuQzcB9KxruHU/lBQRm8G7YcQF3Csq0iCI3yA8582L+9pWivlCPaF4MU
ojwBTAZoHYZf2QSoTxykUjN0+5k7FOl/Pb6aDg0aBZvVzycxAf7SKHRupFD916rvs4d1fdSFd0Ch
wuRWBGEJ/TtrhTNqAA89WfVMfLF4sobgB9plFXH640BaFRqnpXwvD+U1x6yPPZt80zI928TP8TYe
ZIr8S4LGly52+dc9sLGsnSo+rttEHCZw802i9huMz46Px2TAa8Nm66Z6RGahWIsgFpaHiyQL+CW1
3jFmzHItUWF1VANqdaelWSjKbNxVkGm11ecw8lB3saYtLZkdmlze+1B/d8JKylRv1frWsAm0IkW4
NEj1U/8W0LFj5lmXM4lyxKIB9RpC4WQtn/nP0WFO97oM0UVQX87tUsbFIYXrjDhWdHi6e39/Rw3A
HHEsPi0pJqa0Ic/pCcOgMjUeKkDBU93c0cypeZdlkmOSlIxPTwRplgqCdBIDnT5g5EIWXzxx/POb
ZW8Z5tq2Fw61ICbA9TdZDMVHws5X0ej7YecQ4VZiUUso3fBUkTeBZQS6XJ1l4lJ2HSGBiBnON3px
bHDCcixInd4iterVI6+B/TOkUsZ55QxG+PqDPiStPj0iF1N/XieVr3ckqhDS0tk1fxwwjeUIfGCi
+NWyC9wZQdukBkJfdhJH3fm8I0MBBYPKfWDIkSojHCV2IE1m713HvNM5DdfNYllrVamYlrsHA4LC
dIDMvcQWFmFVxlRROHkaDCcYeDbB2yOnVb/77L1wuLEBJwcNjCqHodQm6n2rcRiI3NLiPPP2L/3T
SLKNgDI+nbLxbPfK5vtuQTk+cKF86gdHQ9+NhlXBAY87TNXGk/Vx25sTuWoAdlSaSjdfEh6ta9Y0
B1ENQAfxVt0/XEjockdavcFzTMCBSUWYEinXww0Vude/v4io5QYowVvRrqhBGxOxqBnsv2FL1piV
7mC5fSXWjf3Q1hdOxINh5ad7ctsPt+vNbhS1SmiyqdnHvu0hYSMekVUwkZS7omQ8tVr+k+r84VT7
kozvnM+C0co6grS2CoVwGDrze8FgJ625f+h7qBms368gs4INP34BfU/QcqCfpjq0f1Swqfte0fyj
/WALV3NfTnI+lhfyG+kq8uwdAhOEfqvQ7VCsgC19jOaA8MZ3cJnueeJAiOA7Hlq6Ak7t/nh5rkGA
Bb515o7XMs8r932Jia2mgInZYJ2bAk34Dt1hUkWWLYdX7twe9gmlBQ0bRfZblXC43etufNBQedG/
xa+t97c9akpBnBFPMEUOUXvhW+isNl6IJ5nqKkIdVOKIl6z4OrUpDOlKYJczM9aG5tzm/vC05PsZ
mS3h8CmKjb1Wd18iweGgAzb9R8DxhelqouBV1S+F2SnLaD0o7xCWEhmCwGz5gra+2xZ8bdxGKX4E
avFL5MkwB7ytTHQ8QPPtGItGQ+N07dK/U9IWl0sWw8JKp18J2LdMbfgwWVZKHGw2sAzHBhCq37R8
I6nsPkiRbo+uTO2psd8VFcYLk3F1tqF1kNtga61zXKnodO1iZW06g6Z6GKINopPfkO0UJIXEvLx7
vWa2NfLRacgD5J1S9Ojhyr6m24v62kRb6kHr3RxvW7UODAL2li7/SmqLiPksQ8DWhfoU+2b7dVu5
NEk0+fsKDiLvOF/dWszs28tF/RydRO4njCTH0Mu3x4/wN3zi4et0JUz7P3D8AwEXiOloFpaBIcG8
apbwbHqh0zfsHhduoQx6ubHYE6+h1vIueXosV+WRYCzAGh9dQ+kPFds21yyRWGQiEN/BvPX9eLZL
X/wTIyCt1eNGdPUVUkvu6UHetPnHIi616a+7f8pyVfVHcD9KHOUYLLoPLRAhc0/rc/53boBCKgN2
8ors5KeB+XVC0rXej5YS5BgJKV/MB8T0uwH9orz+ITEh0BQl8ht8agdLWmwg6Rruu1QkU0Izgfs+
sojSzU4p3heChL148D0QH3f1kiA2ejuXmAWCZl7QLQ5BeTs1j6jAniAdRYbg8npXKWe6msSHTAFQ
Ievlnf5kRezWhR3G0Y0Ze2VzVyHKv9zURN3tibjahuYWVCsb7nS68mnTCPOgDLaYLNqBSn2qQJXj
9++pb1K/U+IbU2I36QOhF6VTt9njx5jyWAuX1QVTyKD/84nFqiIi/MeuvLfV9SjQnEOa7mqZgiMU
r9AOFLq+VZJY+cyyu8zw2gVb/QtiG4RisHuhUYl89vq5eHJTyC7u5UblDHSK6AGhoOGnwNFYUxue
gWBL+QBWg5VXjjTZLabASq0dlulLjKXLw8pqJXqBZUXXCIdUjOAlvJWKaULrS0UaTLfaZNTbpKUa
d6rthW4P2WXtZRQ+ACLXGHaMh2HT3vzLf2uVzC942Yblr7rOylNwXiZyynQS6UGPt033KBK38OA3
xXa+KAci3MFMbA+dmveUWwu9+Y7ww0Pi+Dxq+FkFUzjJfDQ7UxgBd3aCt3FLJELUpcoUUY2gvQr+
DkH6AklnHZiRvzkyx51mZN5B6u8d/GpzoIxucP6oqKy0Y98q/BwHA74KM8Yu1fXCVK2LFGL1miG5
mOjpZhWBrFn8Ovt9NvURpIp+IbZyyyUtZDDwHcskufS/LFhWyZ/7qCqoYjg1NE8OMMV6YKDAlA/f
s0fg1VALbui0Ik0Rf+XBzjlIewCfpdpIymxaDZgcQIKeA7nu1GtUvrcVd4DH2cLyZeTYEg0pQ7rp
Jv+OL4sGtpX3jAtbnwV2I23ztVOp7IRGf9pMdboZRkHuIfiimsp6+Kw74QIKjbvBP4PDmm90TqdY
j+tJCp8H0MvXSCfXBQyqezza/9ro9hsHg1fn1axo7mXDZpKSKzGbcnv/gMXHGsk6L2cEMBnNfsxL
LZBW4OabrLc2yhcyHNEIvX2v6wNA4cE9kV//mtl8d2WIfJwxQFf4Ci6U1AVNU7KvsQ6pMXhSGIQJ
gkSvXtqVw3550bQP/4mmhi5eR/YFYR53gtsM1+0lvDZZN8PPpg99yLlED5d1L1XlbJaqrRAvfTyt
pbC0N2wTAV+YDz+hmDSZdKFySSdk9koqMic+BO+NYcuATFzlVZ4OJtXISPK4XUbAgm50inDkCvUO
/HzJuFHyQ7zaiSoglkj2oNR1J06ew2V+/eDpAQgThAjKgD/H+dJxRuHv2McEimX76B5lFVJ+SsWs
s/eb9mNtnI4OefjOMD3oSWBVcScipWNH1CA5z3bV0EnanmlJtw1W/zGpOhcRPFYnfgOyPljXVztR
4j3SqSXN2FymhundkWQp94cjG9lok2qcLy7b5/Rmjkh9wDdbKxABfuOqX6tiQgKWKk9w/OrOu6Za
+s9hzDPuMMuRHpkc1tgmoViZF853jNa7cUA/rcMpMND8Z2G4SoTpPMKsnnGtY+/V7hgzf3UzXTtQ
wA0tlG3Lg4+tWUQC3hpxhy/0MESh0uz20w+IqjrLKaG61gGT1CkG6Mb4ubCyFCTHwTiDf0QhKCwz
c2q1VIFSgnDqVLm9teSqSHA7RqsIyHL01+vChC1Cfa9Ydu4+pni6lNKxzLcaf1n6DhAx7hSDr7Jw
oTaeT9CkjBzUFiMEdqrbPq9efJsU0cSDUiK2VlyXGzUk6NEyg28rsz++weWZR1eI03SAbAHBWCNI
bydYJQ8OLJpF7AJ8cx6d2ueE4NJq5fBke+GXzQ/pd2lha8+dodPjlnQji1C+ZncjhlI1kSaDmCa7
r3dLyy0/B92M0PoMKn+ZoUQMOBSTenRooN3vKni+cCPuD0HXPYd1+xy/92A/xMx92/mI3DCsxl0l
mdEmtzG3OkL3YAL5p5zmnxtjy9Szt6Ky0xprvC13S8Ox1rmOcgHShRQO8yyrPMlOs7MYHLQjKY8W
KueAJHJHISSO+eTaq2CW3wR7NoKOvhe2OEZRgbjE6ou0icNqRD4N0WQGABFn9KvLQnaXbOBs8Mv2
Aq4zXsoyVJY9UnO2AChoef2ebU6IoJQ8V0fMsqrSVWJudQ35oPHUDvBLF/O+G3v4ftiPQBfy1Rn2
UAOt4ix/iTF1GglDiqEJTXNLC1Xd42vYQKUReQ1j7mCqIjFDFBR3rJ6ogZO0cvE9q9LG7R+xZBYf
g3Xcii4A+3XDWA1u5XGQ/KL/tLoQDiP9BCU90j0CtmAjxa9SXVMFgR43CUcfU530MYo5GEZ1ShFT
kb8VPtENv5AUq1EYO3/o8z3Kcf25NAO+d2uYYtU14HjPjn3KD8oeQpOsNK0qe2Km79waNxN6LHgQ
+v8ZT4VNEXO/VfxjEqpvBRZ19ySLUfcSuW6Rum3NfvTbzGfW3jbisOVH/vCn7Nge0w0TVvqs3deZ
uAmOQ42Rvo0QiSkRP1xAPIOCjfmYn80ZP7hL/olIvPq+9zz4537wrpYz0yyQ1VFCcRqVcVtLxSuo
24+NSxw7ywiCASfDnh13EnhIehb31/GVjghnsSwV1H9LLVrz4h8gyLyN3Bl5TmyewanTHg7RfW94
lku7Kl6F9EC3mAMjZw2keFAtFHyEbor9DvbIJbHRVIL0AjPKq3r0ZR159cf2wIegO/bQMe/iO452
zbig8ULlo8Xr1N8Y1aVsrPCV8SQsFq2Ln2pfaXJ/AMNU+xFgIrEm2HKs6mdzuu43pI/HWdzlRbDH
neI+NIO1/lb0pmz9HWotbDU8Yhn7Tyec4Xn/y+rd3mAR2t6ea30dXRKTktTfFREfTOcJ5iqoRXFf
5BIqRyRQOKrtyUuSkJwqC+HphPjkGIE9SPmbu2JaGKp88jqZk4HBCnCcTeSg7u5AfYbpNhM8xGWs
J0hE2KPCP/LJzlf5W0QoYmKVQzTlNV2K0Hk82KUEatfFIZJN7cIGj5BVhFMnbnc6SsM2kbs/mdPU
khzM3RNGqkz6RRq41tWDOG2L0IXXav6j1b4vkqUINCNpENSMVGe5LHYsw5SGuxt0JmeXfSxFcCGR
jO6+N5jZUYwOb3shyQHREUuTw59lHFzkGGfuFINLV7q6iY4SYSLGuo+y3H3EioIq4R+TWneuBNzj
bSbvhcHvH5v7LTVfgjou8pqPLxoEEF3irSM0Ij/9AjzJaVbstv9bAWNAV1TtwDh/EKd0eJxqNxce
eKeQ5SeCtVG6bWUT2lDd99G2x7ggzh7SgQRw6iFJ4K0Ic2EO+qfC2fp/hL95bXSoxZC/t04+/yv1
SzXRNDIsMfSp303YsU3TNRkXdzG3m1V1aJx4gcx8kKwjLEOCwCXFoxinrKkk9mKR+AAgscASurMh
aTmk3b4s/NShYHGdrvzxGbN7Zo4Q+ltztgbTho60z+ZM0SnlM8+va4XA8ptwLwCdwZLkzITewQwJ
lPcVQxd4g+DVGmMTYTy+Z7h+kyrlsIS8YCqxC8o0Kl/dJ7JCEVfvbDk4qhQjzXqwMoRXKcR8ylGx
L4z44ZrTvTLkhzKZDKo9w4ZfRrqZp/oJRQds1ypMeMY+Bp0RiJn5IUsNWMfRIfEVY1/V9AxMxQKo
zFSfQTfecZiPjpVauCnpn1ZMflnTux2Dxqudu4vcpysIsJmThpS+BEuFIAluRltUZYPINi6b7JU3
8EgSw2+Tx95DYoUwD819c43ECR9MM/YMiurM+nThyUKhcu5V0HdRJiEme7v3n+nOiupTkjisX22N
tONBXID0cms8XOHIQGe9JeQSmBe89LvZDFtT8aJYR9yRwiUi7dMwe2xiF4cJP1DrK5GjKogHINMI
d2BKyA10PNJYr5PFuHECIpwTsJ+2lVOLDR2Wi4Aoxgs2MiiRKSTVOUWoRMvRWRBl/9h7W3/l/0fD
LZy3cS4/JusqERa+CCJ7s4tGYogTsa5v9ICMpLGcnhMc0N1hm6rUnjkffycHVynqSvJXFFL2v+sC
sdZiV9livJd69DFGItYFSIPBjmVQ7HxVvAcPxtVZlN/taHyau/85cUdJWL7KSqP2BhR6mOTNkmBm
D3gfILNSqPQlsKfOKwukR0StnhACSZHiZRCbMeqFOnRuuC8N32uRN0JuyGbgtiqqPVgLIdrwKJy3
RZfGlwFfRCIRizYGyH3XdoqPa92cNlXjMzpAA8DehCG8+K1WmMUcjn86s0vhX3/FHLYA2xj1wc1q
jORBOBWykd8/5mHXS5MCiYKj9j77VE4gPQD/jprdj1OqLaC8TPQnxYoK/OaV5cCr0etC61Sq7UQJ
z9fC6iu1/MyyhCziidXrV062sI5FL9Llcue1ODhu39sR0KlmpBvg+OWVcCQMD+3UmV66PXZ3IrvN
nbNxSqokBawO/jkQL6+PmBkCXovTOhia0MW1hYG7zuf/3GKpdFVz7EYY46tWrQS2bme+Pb23tvJL
6adgBCty/7txMz+SaxVUIPxEKRQ3GOzpvu7vCaUJSdh/Gzo9ujIK54L7m0cw7Wo7ECQ+U0fStq+d
s5hLzSt2+GIykxlEqKDI8KabzyVxvkwwdOXT8YAUxMjFlwU4feoaBBfQLdlX0wBdfRFGLzSE7IXx
rCltcFsT/UdTEwo2oGJjae3yKMyyxSpVNXUOCb4VR4BEi2OcuJwCannc/YOarJGdKEG4D3zdTe3S
H3p0j7aYSv5xl9OJMHiH1hqme01h5KAhZCoe21wi6GYTq0LQkn+N/p7vb4/DS6s7rzFVSuVCfS4d
9XePRLWQY0RX/diUfuoVBK34/NXldVMFKYGRaMwUsbLj8AkTA8IdIzuSRDZA5mmJVyHZfwVQhPKo
oUEWycfBr0f9MW3MNpw8oVbWKqLMYjkk8duZBU+2aj+D7XUwM0qW2HMaUrwJV91wTZWaXRD5ZGVZ
NRyyxEi61rkFVCpJ6o3bkmZ0xnxSmXIu0M4DAwohn28GsemVG42tnrl4CrNRZVWsV0mDEr6Qh6gI
5snbtb0Z8GvPzUniCXiWRNULdsgxp6lupCl1BVsVMoQMGTxsr5D81I11prgIypvQBgXBY2rtPJQz
GzGs60fkikU0eSFmWFfzOTldKWyS9yDMnTm8GLF9FJ3M6aNQCy4/MnezLPOLhB3zrdUdfKXbECO3
rroQNSCpZsmJxydoh4om6XfkLP89vdPYJRHBgRL1lOtUVqv9phEoV9lvExKete2JoeDPy1P24EdI
fNbU/4mJ0M86I63vA+qqo2MmqN6IIwipFiFgj6u56sC5JV7R25oLi+QAbhZ159EZRoVxn92f4VMX
mvAeffblxQ/2+QjQ1JWpBwIiJ9uz+8ith2CAphb4rP0jEenUNBu22TwElGOdyrkyAyNCuevJHRD9
t9I3M+mAAyeQPBKGet2TGE5Ps4Sagyzj+eJW6CVeQd55z7Crl9h+26ZHgDcgtK+TgxoCzGLOpovi
2FZwcpT4fxBua5U3HS9zMRStNkRwN1r40ar65ciXEQhWRT4+WFrJ0fXHIUPwqMGArnwQ+BV6bIR3
j0Kj8out6T4X+qoHYGL6EvcpIVHu62Q7zm3BYVIdhqDppKtYnrPLZzOm8oBbPIePHEvKJV0q+kWD
Khr+ykjo0/l/BBVGGzXwIplD5CuKAJN8kDgxVDKCeMKnPmQVEGuPnVIv0TLpKsplTw0FqSVcOXPF
yHz09SOHb1nSF97dydifaQoFtjHlgWiC3zIex0sEBw0INKyabLJp+lTA6hOFuUKaVDOLKi7wYv2A
Jnwa69qxcR/oXOI9UZf+/tl5HegClf7K3Tsby7zjhPuhQiqp0beyYpGZIRxNkNluSXpuer2JzHly
WTAdPXUTFXnf8zojyyTw3I5kRkX+NUYJC++T1Ubr8uaeVAd6UqBYMZhflfAWpn3Ceofj3wiSc25J
y82ykU03FL8JXR80v1iCCO0d9mwawVpQGOj0p+TqoJPGI5ypObF0Jnqk48sGzHkpdjyYLlfKXo22
f9NFgr1yQCKz7zKOnR7+AnXZlX0HCHtxXeL/zjmK0bsj7ZP4dw8glIh1yXDc2alfmZ620kmnJREW
AYKvy8BWA/efuFRzdJODcYzNv+gjFVkwKVgDypQtjPXUA+ar4EOE/SHwjOXP6thTKokkDX1jx5hA
xQE8hnO7M76ZUk5tmqSrW/smVLV/iqomyA8RSXqp2AZ3HsZuSkgiY6VQS3zct/oY1INvb07Oukn5
OBY5pthfAFXf+1DO9cqdJmbrHMaqdsbJCmD0Xad5VUs3Njh5z++RPWUYDBJOx5OA47vsjyYdptta
owCf7eQkc+POBaYYon7BGkxgBfVAdJMYPBDX3y9I+kP2Sfrs3iPpBDKqON4MQ6dEd+MeFJnMb0HF
j6aKzREf40LHZLlfT95xtkFDbNjj5vImVy0BBvs70vcGe6CipMFxcGdupIaP/vb++4aOUD5rdM+Q
zbpUlXhoCdr5cQ9JIbC+V0YxxQtjyLFInrvoX6v14IRNuLLkbVVEt8SJ17qWHv/UXSiq+22FIQ7J
LpCms7ePBQ2m4yLnIbirGDQtRYm/zG5KdOjOkHeGJEfoTO992lWJ+Epm0D5EV5PIe0F0Lat/g5QJ
/bJRMfkGLiwMuhOw9PQPQgLk7M5R18jIPL9hp9a+iTh6qzuidyew8XATl1jZ1wJ0NpxrNjcNEMeu
fvDtgz3jurpelrGom3QOkZVUwMz/Y+ZLi49GGdBHS1QNIG53yWTBVv13FWkXnpUQchUUiZroxner
pd+aoFCCGmUynsyBY9j9ZB+Ogq5PuUwLueOOBjBuRGESZpdAjY0b3q0woj/UdlSQiQq8tq/z0DNi
tDOqDVl80jfzxRZdGiU9tcQz3Z3AeDEZusqoGCnfMnA7p0ZCg+wtaQSokr5Fr+xqZTHr8a6Y1kAH
+4j+z1Pemr3IhT8/1Bt3xRh7cPY25SFXrfRK7p+3VRKssO5ylVzfU9XlfT5m6sskvg7jwJXa9Hoj
3ERVfXWItGXM7B9gAdV52Zcl/Uo373cmxI7S7JtdF6e8Z5E3aYPjhccw+5CIAaOA2Tom9ylNwYYO
EUXXZgG5vuTSynQttcAZgB3P9h0PBxP0JUYfXiuDL37zKRpZaL51VHj5DDiixGoXy5sh3vAFzmGy
mOHgecYjloXGLq1e30fK79FQ8FTX6Yxd+TJf6ykJvuEj88DCLy+oK/UcIwTBuoSbQgtTqYMXDQlP
SkLAFIRwPkD6dxW0kwXTMJORxet3zfVUzUJOu6RcM9aZskNL/CvJp7DtdCoBwTPgHQfO3ZQSR4RO
rUznOAHvuTkvleRnS1pETr4tS/tALX9vxmzqt04kJ9PTfDy1zRPbH9hlhIOZIIBNUoZaX/RcZEsk
xdztoJ6t4jsBTiC/Tz0l1NLjvoyyHZOmZbW/fyUwmMNJALbt1fNIRCN+7bCSZ4VRCmcRSjlmA1Fo
sVigHx1g+DUa9EVVfJvAdW+By7B711UnLS0ppePKpjuRgU4ddqGQzAgbg29AM5FBU/m6CoIRpa5L
medt70UlxoEcA0PioafSjYn9jL/c3Qt6TCPWGhybZiBnI2HMK8nS92/1AqP4SBzpj6FGYqzfj+Qh
4coFxX3fVwH7+pg09QFLefPYm8V1h8VQUPu6MWNPAuTk0IVUdvX1BgRLGjsPzwGnFVBcZj2r+3KO
yzogS77GlY1VpjmjA7srdiogV9ZwCuM3R1lXxALnNf3UToTRIPr50ZjPjMaaffpCkaMBq0vfIkIF
4aVnNI0n4fjNFpSsPa1+BX8C+o7/HEtPCQ+W5aHVj+iU8B38+UNKk8EcFKDEwWMGBSpHhwzoQoPW
bCHpaRkov1TmxiAZrTMCIP/YXoWW81VZ8vnD2NAE2foRaV1EfkiY/w/Ikw99aoMCS8sRh0mziQcP
e7fZvTlx/xlo805hXXrqk/9U+slBZiDI4zmc2CDI0RsMvqVeFecKS1F/T1dI8VMK6gGA9TpFDX/h
xuY5yRk9bZqwp8YSx3G4o2g+2qdmCj4fDMap/EoVbymICCBT3Kw/BbTsz8fIzeTEy8fjGfGDl16f
OQLzfANNclWnEw9hjnUMHm0hIeCr+bL+6/fl8N1w/eyJDNGiCbEGSRYNDvfAYRQVuvIcXDkedJjx
cSb/H10G7QlitLRYPRfYTW5gcmQPtxhWzucXvRFLsSWJKG6d+CVoTg1XMW17SbiSHKEcAQ2eDQuG
8jbzfTBjIBjYOS9t8DD23Dcj4B5oG8o+4lFYs+tGUPn1hDoyfd2IZXwWUAOB1heKWIx6EpvQZ1Cd
cF2CzIdotgPGc9Va7ZgOwH/AmOn+z8msQBZZ5mfZ2ijXzHNhg1uqEsOCxIq0e+EHgx+3iQyWdyl9
wJme1vKYO6scpScOiJiE8AEZ8yXOUr7y5D1VfIkFiJu0dT8REKZ8hMB+rCeblWKtbCC1gmIconZU
ZoL7VCqVgZIu/sw5j8Xpo6IJ+O72/dQrxUFqdZI6x3La+ZrUS052R0VsmJOE1rmRdcTYRZDWS0Kh
A298rgpDk0L/sGHLSOYvd2yfSs2hipR25xnoGlqEB8/WF+Niko4GMSg70b7iosXKuN4VHSrmuoLO
bU703pYYKigCG9NRlyrpXptdGPH0PhaGiLx89iJC4ooIDz2me4I0hQdTjaZCGoaNJJ6UZWZgFxVR
Kxq8RaI3WU6jeae7Ihh+IagdwXBEieMFWkbcXyuvERbKJ3c2zx5ahJPTVuSd31aHQNhBreJpMSDG
mo5OPJ1Ck5FLBczX7wq8L/5UytyL7O4BBBEB3/dlWe2gVy8aDj2J6BOJTOWbA4MZi8YH6E60CAI3
EgyipF9+uLHyKAYe/f8O7kyorDSmxlqAHdCTuiRd6givE+/LjZDxkHeRx4aUwNsS8T1Be9CA17nA
11fT3idz2zzPqXc4v7ZhuRmdVII8yswz6WtGJlUDztDK18NJ/c8LJBKn9//ZxP/sEQYGYoZUDYOi
9uq7kLVQXw4782SrT2I7ple12I4V2tpJEAzdpLJL0HftmwM6CIzOL4FVo1IpDGmupVwxn+z1FOr8
ugtJAfd/ROUcqHOX4I1/xZJHJ9Rt/rkFW0OvH0gv/EIS9U4tkWlGZY2XPqI5HhbCQGS1c8AWbtE6
c9Jeu5IoTzqD6jqPJzzPlHRzb+fVDk93nGHe3tkJdw0O5i9stMe+YLAPQbP3aOOqRW8Z0xPg5bkU
zvVzE3jHP3IGOnaZ/+XBMasNOGZeT6/CW1qSFgDkRYZpkk8NffeneGZl+c6FpMlcfDsRvgwr5suw
Ls44KaQtqp3CLRrG+5ZcmFu+V8OLtfZULR8MNC9/3ehtXHLMTWSaj3i20NNLaCMdg1PAukkcbpVK
5bO+ox0op90ToYcm6Oco4DQvHkb2s67vz8ZC9stCgLYmkd/rxNe9v4ttU2F9KpDpTYjyEVDyfkPE
t0JxQgw7ER9eX/eDtess1AEM41ZDrji1AC3aOXKHgso1qSF0ZJyPkuF7d7IocJwA36W5FJ4ffPWg
sIkl0Cgn3D/HzgNK0Y9wmCL5XxqLSVwLctfLCxryP6gDtfKCSo6f8XqSmCbu48y7SeF0CTLoFYSO
3EbmyP6LHA/32jj6IdGerMTBe1e206MUeTatioS0NbHrUoyvaI3o/DLlra8yqtVwF29nw8alGyTY
mCFKwzhJM70B//d8i6+TK9fUKPMaUF4Tt7yhyM1aMZzGSFwwtiqjlDlcfNHSkWGMm7aT6Qtde6WQ
oMxaz/YHUzM6Rz4O5sCivDEKBdUK+OYDmbW/XtQ4q3dtTVIC73GnYnYhZddwUHUnMLYly96/i6Pp
HT7/uWZVOOwudb8tXP0W0gbFGVMZizmh7Ji74qmV4Eaq+t9VMxLHBeNuAIfkUE2ZW7CP3nmlinnm
jUQllNG97IAXxFjN2T1h0qJ5LfvMNp9bS5pZ3IK3EpABV5WWdQiV3drq8Ojbxdn3syXV4IHaSVa+
iNQjEu+lu0gCG16EzHkxQq6Yuku74PhsGsHf0S6ARGjscv/AaxByC6Ufa+f2vEfEhMDIazCPMy3U
xza4hyZRlO6WA20+fwR7PTWgl2/bYB0hclHz47YEjCkghiwLTLvDz5tlK0McLkvXX/iMcAVghPr5
7lI3NF7hPizr96mtx43DGbMZHX+c9g+PpjGZLFC8cHS7MbsBDdC/lNmUpmpkrIrCvdATANp/Fg9q
0yRD0nxwvouL4WVoAn4l9IdZJ7qVPAxBDpDPmYTsmiN1zeF6hECRAp1G6bS9omgoCq8zNW/0r0W2
oeXb9NH1E/AczpnLBR0HICmkIc/cu8GlG7goYdVS7MVIdnptunozMQLCyR+q1mpBRPJk35JyZ8RX
Ip4UKdy0WeRwnNmVUSYT4jYUPopr90kxqY7yK6P0FL0BhRXwjOkP/AqGjIvP0JcMTnhvLd4M2TDA
ZvIUNzbxYPhBmg7MBsq3ZrYdLjrsfLrgST77WXNddBP+8v991bGfMgV+95sjcwu9jp7DISsKWQgB
e0axdRlIU7+y+zBhSAr/mjyKnuk1hWvjZn/dxoMY0VdVaWUYP13EU7Zp05ASjRFva5zRCECzxtZg
s+cePYCE0wA0A0cO5C5d/2xmNqWjD1gmV9rgxS7aQ3+3YAw4aESx04VdR5acvPDx66CdM8Htz7jw
APD0msoyMF0tzORT+2rrN8SRgS3gIaO0PdzEYYRFPXLFMrOE8k8PY8nwdpfw57Unron7dtx2qzdq
cLluZgRwezJ3/tB5n5RjEzbaSmFaJX39HX25C73kamjhk7H3jaxHL0NoqvU0ahJ4or1zvHGZ+ZLI
/JzBVHtk9BfvLMsTNVOfY7OMesdbcqYJDU+zrgeqH/LVJj4XVhN/I9vK3yGa4k8lZGP6C0x0nU9l
ALB65tEQ+Rbm2fKUOKfjqs+xsBlPuSF3/Ub4ESCdNLXtEa2kfkQPLFk5sa/skIbJ9j5PNfNXUGlo
2AxoEO1kfMYksR6w69WbX+IgqJAFp8IAC6xiTcM7+ulOSQ+bYr1nDR83mzsK1IxNfKCPypzh7NQs
RkuXGYXsbs8c5BWQzXfXjiP/YyAe5m8SSjjCMvJYXYT3NzNMRKfVZv/N8MEb4R7w1U7gXh6CXAHx
l3kb7uZgT32PyIWDuE0bG7UMJnfbnoipl70HjFBsD10oSlcOicG/bVbBEffX/JTe4jEErYPh/w4I
M0Ks3hqrMZyb6xCp9JMmeQ9Q1qUbx5ZV/rbGNq2WUlGq8sSy8nnBk6+fsCoXPMXY6JxgPF+mI5pP
0i2qpR6o+0JPoJ5eU66IwvOFFrqP3nNCila/lP2mbZNiC4SU/YdGtzrPCmuGaF9ktZuXwFha5G4B
5nCoG2tdb17ksgh06aDmwP7LHV6U/1CvHaG6zXY2+pS7aJYadf0ZH3vks6vGcfHwgf1ju+5wup3Y
wFfLgChy9yWIIh+evEbqOc+mOAdDAHnBA7KiAC6O/pei1oLrDf37k3NUHIwlwtUuxPcZnzVar0cf
H3iTcIieqYW9ZYGFExq+SRJ9MpvNIIRxn5joxazB/9SNU3azTyPAvdLR5Y2WaqKxrmGViozrc/vp
h+QDQdjnHfZpPAISfDMn3CXoxi8q6nx9IJiS3l2E0dv4DyfBxkLeVVxM7+DpEwVz1focxG/1W5QI
F81RWqQ73NqpNCnAfo6bzdhMmhg2eY3xy8n9zoETUaG0+5Lo6Lw7rcRLPUofz+3Mm0OT3XQ9TRJC
5hHWtANEx4racXViz4WTcXVi0VrX6gXSCLdRDxrPmtiw4F8fXKXrONVsJYOGJIjy0dXPZNQ2ndbR
evl9ppH6IE+zmehWhboMbuKrHbmqLfLJbW7ZIyK1W32y8oTDDEYZWraiaCfDe1JE54tKXUhRPQg9
8weqbz+sp/NI8X6qynyEAMzSBEM0c/6Zmuy99p2JAfCgSr7vZJsaxrHnAIcYAXSBqaxku5FTfFs9
74jXnWSjzt2P/upvsTI5nM5E+bni7eTsOuuf1Ym/5FXxPBZYembQwuSNAfE1aOezsNuuxRa08SCB
88KIuka5kcMwxQdx7ihjt+tvmVbXXJW81qCzady3X8ZJ58ipU+8I44ErsCK3AxhbIGHZNKFtlh/k
m1/IdKu8qztPs9LEQfgJW9UzRedrLHKr1qBqIepvZEnSJJ0N3sflLyTdDD1UebHrct1MQ0Sq3BwM
t9BJeckFjTQ/lAMk1PEqw8lgfaD/DxBp8MqJfTW1y526qikTEnUZZzYLgv4LCoQvnZGriR1rm7v7
4Q/HE5dn55Oo+zyS97WIfFSmJCHeH6calp3jC7JYrB7QQchVNAF7wh/ir5/Xvt9+H6nEggpr1tY+
oVZQAFBf4FywWbcGGpWAJiRdZlbyvqnpe4+XoWXQVWMLTK5H63k1tnwc3IoOOU077+FlDb7AQS7H
rUmH+UIUGAxE5owYHZDnuoAXnGxl4PrbT9drYFYcAUB0hE7VmTKEMHq0qM+ZCrax+jjSTGwOa35I
/CNkkxwuPn3vOyv3XNxdnZk0Cv+u07LcH8Upu8JiIy0A6rbMReJEw5T1w25/eyQ/G9Zd9yZFIeXI
+x9gS6AOM9JJQn9oY2Ew8Fqk/aZ/oUz9cZS+E/a9bOPTSqyRo3stwd8N3lqc8+DUywvfWZ7EgRnY
aWZpT1Otb1l64F/Z2GBlEd1gB2kM2fyRhpr6N4fm7YLp72r7xGPLpBj7aPhd98BkKAD8oY778DRv
iSWcL33or6Dc+ANIyW4oBflg+wdJahOaATJGpYsjlwvCuEj58S8yjPJLcX7kyn3Ox0VWAawH3yX4
u6ENqgMM9TSH5hvhA99GsmMKsEvlD4kVEVR7Omn++4tznFCLuf7hInbZdxo5rQ6XVuHw0zwhHO+E
gW5YuXUidJB0zv8bJI1BQxW6p1N1I8pbN7MR5PENVrHZSJ+x6HU8jWWzzdwyzw0fBoDGUv+DovF/
6yENiE0CuY7lSh4kGD9AZkWQnSwmb7F/CjVmBkucj8utAM94Wo+Ab20xlvIPCxlk6WlMBajKPXq1
6AIEKyrkmJv349WgBCjBF+mI7gDg93mq2tEXzO46XuuuPM5nmRHmbtkuArcIilQ7sYZ+hiPOI3DH
2lxrsEFC/sZDA862KXEkVN5uQfpyoI/k2fmuBPREleB/PR0hWZfGXFHiOHUVFV3RQgQ+mLxECZXY
T8RALAvTxKN69X3Da9tuG5NjoFNSIdhmCsguhVjlJ1I0sHg9F3w6oQVZEEVb0bZJ6hGlFyrJbmDU
AR5I6lofT7VXkkGShUe7vJOCxiMI9nEeOH7+TY/kRwxYYlZU4eN8ip3GndNRL6w2ykQ5n77xZeSE
p8wCmD7UX4nkofK9DPNi15B0bfTi4q41ub7eEdoDNQcELnVqSyRYwYX8p+tbJsSRn3EayBTsmrar
2Iar8qBEmbDFl90bDB8lSqIf15w5j8OlVq9hOzDspINNrodP5DRN+8NkxY8IQ2dGR28TyBj1MTGD
e7e9FWDzkjoSdnUQlgSKXUWYgd++d6TdpQTpA+0pC6WQxrCtm5CwsRMVu9NDCZbs1DwC2QEJ+Wbp
g4EBfFBvSFahi2jfHO9nKXkUnFttHHJtVibnZ44QhcRhim6nb7H4eAOOVaBSBv+xZcz8gD33ql1T
dBcdYmnr6NN7Hox6UBQcMMmKzLcFuxND/nIzhP/+dGmwQJOVxBCmD42fO8znXkrYpxWgncrCNyLA
yxTB6UfKAm5NBYWRqV7LSwg/kodRJoWsuF167TceRdbEY7c8VXHlGNML/kISboG2sKKR0XWrOS5v
+W+bjKVEbS3rdYu83FtA9E7wnJBaI5x7IQ7M5h0HMsri8N8bcobMW/+JpibWk6m11bD9dQsAD3lO
CEsgxuA08OBZwzUqPF7F6JNAI460DiYOeE378zLQZZ2SeAo6cCW62Wu8gPVLb57/yflqa4mF7noH
DIG6CgJJy6bNC4LT3YzkHDblsec+0+anMCPVIfaPyWVmyIyHhQi+iR/gHb/Asq3mDxQ57EsF1P8A
twa2AOEb2QUp9C+m76yLvZLKRN3Urn0PCjN7XISBLIAx0cXcourx4Sxa8IDrFeICeNMyXyejLDH2
Zp3WOKkxC3lb/78iVJXyfn+z7iwnygzHVnQPKb2ZeH4sG4RnNWs6fmnQB0tsDNxMg5J4DDcff8bR
alXAJ6JAw20sYybfMPBKQcswcqUxtLse39C0aOFg9kORBsL1ZYXLwRQeKRxr0BHe0EYUx3+8DU58
hxVwFY1et1+ACzRkzxb4XBD6zbb3yRJ2x4Yf6Py+AlFA+idhvqrMdHd9YCb+pgV/Ihk+9P+qVIrf
JajLLEXOQvDeKA0twA8d7cSWkxlBoUBPOBpZRJBROwMQ1ei9PRMqH+0VHNbYcDc0HkjaSmQMnJm4
IvBaSlKfAogToKJ41u+tRhymMDSulZk3HOq1RjvMzjbnJ/CT9x+ZDt6c2nt+yLhfP2BukougE76J
aXk+5hl8f1IvvG84aAIySP80KsC7VY+SALKF+cmqZvIOF3WpRS5LzdY2xludo1LZh9UWb8ZMbuUF
5xG38rrIIR2TJbhNlsHTZH3EJtOWkEuTbttrf5ft/uJRrZ2WPDRlEpirDn0s8uYiJ9wUkwvFcfeM
pikoqZTe+1zSY+3QVhKdCMD+KCINiahiyfTCPJ2cSfdAF7WBGwlo8AiWf/5+ftPma3OAZFsjgqer
d3J6VHYKqhQ/qsDzsZJAIywMNZ8GwHjYs/k/e9Ob1I3/d2Fh5r2lXTjYZKt7e3rMZO5FvhX+/Wwp
ABObV9ne+UnW9a0wYrkHsQQemF+yF8Ng/4zmhBFFpKyIcZzW7YkxVyefqPowH83iQl6AjDiex51V
zDHjkIYuDQOO+uVEuIYiwr6S+DCGiemHp2t9Ijo5bJ+sx0jww+vshbDBTBFfkcCMACBXrbVFPCyn
DYTch5X7pAX07OWtA+vyKIPtdStr9WJrV0n0e2O3qPW2nL5QelB0TRkKwsDoaq25WuAuIn9c6bhA
8CP/6+cQHSx9LNIuIFa/aw+w0gDKgbb9jjKWKIUrgdJUYJbly6OCC/Wyo29+bR5kctGvzxVlwpk0
bvvWrgF6wYlLwJW1iHn3H/HTJnu4a8QmHCsg22RPQLMICTl4Vqum0QyCAAGmqVgYb24OSjXEc2sJ
KzLf/3PNnmLzRpcWKNdN0pRS+o8Sr9noyhuyZjPYltmMG5dts/sg0jPaN7nZZ3X26YaliHFhGpJU
9n/gjRAS4ibrbQsPjz5Q8qaqJbwyFlQPSkMVCXsy6Hmp3oaR1bAb7fbhYYc/bPbYKmVjAkSjjBL2
kTqey+GL6vCYn22unFYSbxbIKEHp4olKCGQH0B3jLOvs4Xn81/jBVpWfistpQ3eZNL67jxxzvaCP
PpFe3joTKz+u+uG+ZsvGfGfbK+vKkW5YdyhytbBW066jOtlYvt0pIzIml8UkfLo6nNBPwBl272iM
/YfIvhyyA+fCUBmQgx/3OZPJaS9NMdCcV8at33QG4j2wwKRkhoHvDsy3XwBjuy3j2Kj0lK6587mc
g3aabmaopN6GhkkGnW+vj12zapCPFoPT6zsjNJafUT5wiRj1KS9gFnCHDC36lG2HAdN0NwEg3lUX
OE0707U9WX2iztZZo/YpMrtGfnKzTZ3MUzrcLcI0khLNY+wVDrRV8YtpTCr1sc3CuTotLx+wWMb4
NN3rln6WesUmMPvyU8ZGMZj6M/jHfHoOflfI2+hRCnO6ro2atr6tRTJmRfYOvWcdnt/3duhdQe9G
eLmKCPm/PYwPo9dKGmwgnOgq+SqHjpgVWBnVJ6njdkbTxhWMWLtSkeH0lI6X/OHmd9QtwM5d1s99
IpNGAKJyuiYk6/f9sJOK2oMeJuJtswWrf/FqzTHVbKhVGY2eHTapo7mcq7due+mmK/ztqGpwgtu/
23CEmAk7cv4FzrPoKB6+s6NB7s4CjvdLkBhDPkKmgXZzmyx2xoeuPCRgImMAVJjURa9KcjLOipKO
y33RI0252/ElvWio9h7tetX5Cy+BLd16LHAECtPyzuS68SXMMtxZGN2Fgbv4YZG+HhYvEtNVmhLq
MqWJko2j2DI+zuaAN34SDvI8jkcCIN6eIUA6ZcAR2DV7ceKWP2YTEFzz171WlMakD5y+t/gZ6zCS
Duk79XX8rG73wH0h0TIzcs5b/ESunkZ5MqtElqQpqn05kfDN8bkvPIX2lZGeFQEmwMoJfozJET0i
+7LP6e5Ncm6l26khPEYHJfUJpZKOr17410nvPNHSLTbn4AfE5kjWqEzaWi3/AP8yeJ1y7Lvo467G
Xzk2f1AVQXX21rlQgV6/nlZV4WUIDWESts3EIeksr/G7GZn6eK4UNrW1+SpKK58r7aDs7UREqnBd
c2Dk9XEspPyd97bBSQWhhib+gNoKqUlJ2nc8BhDCanvSm4r9cRHs+SPq06BI1vnkGIllLIaEgHKn
JBx75BUZPaDyKvrx/nHc1rM2SR/4I0Sh+cynsdtPr6DV0mft65M0xgQWgET/QHHZrRK12Pb71J58
nojUuZinkfBMjmWgVcD8/mxberXRjYlI8bc5A8Wsb9OINvK3K/Y2s85eOTtS4r/KgObeq4qm8q4H
Xqg47n3eJWmntfW9kzpCNOeBndH9Ia7rHfT7ea6aSZOteMNF47vesjxyyaAh+FyAyAejZoHg1SpU
VrrFwEA9H4A4DqFQ5jUeFqVv/VrBvhknNHliexrwsgLKXgx2U33Zz0zaAGdrZkbCFk5rJdRtTLd2
bn/hEe0hzspOCbaHOHtTChb53IK2+iWy95T0uPkW8PytLVCaued+gzkEV4ZlcFCSC3FlVIv2K7r/
XCvm1NdBplirt0p0bXg0NdQZXzJ5J5bOwpBzOT7Fb0O1KeACy+6dVrTEG5H81vQ9DCJCowlyjrSf
MGaBm/uT2yABdsIbX7QdSev93NbLBIbQh3SDPBNUrflAAD4jFwKesolfCAoWu2dVxBY2rr1HbOF6
sVxGhYPqHADxzmsPV1YSdv888nKK0higM5ALre3193ERC2oz9I29+6RAkJlDNT+KmXFt1x0RMwnw
crvvG3bsgBMyn8px/HomOQQTSjZLq/pEJfeoTJcXTjVtg9oco4Cxj1Xr5YL8NeYKCuNN8v2/pA9+
/F7hrBrGv+FMS77ooyguHYI19piFtIHQYd+4zjDOaaU9QZshLF4YUmJg3sVg6AsbAy7PLWbBXxC5
oTCY6IsLDc2IQKdiaSHk8+TbsFz2Ng0opP2/cf1jgnDu1kOFWkKRRJaauVvjtTHrQHkShZuUTBpF
RL4LxsqKRYkzbR2dbbu0FFHLkfWi/YTJ/Rx4tgv6AOPmWWkvvJ2YM29PK2VBcPcwqIBEepLsIuHs
06rykSssy0jz8BmklshdkbBZjYTS4AV7bfsgzacN3iR7bWtWRpsJNfGQPQnyfBqDVxwnIE1Xmlm2
XKXfDpQfnTVoLQ52DqFmZy//C1B+IpAvuAOKrkIGIWWjs4ESCNGEQTXNIMp7RIjwXhOYFfmxCi/5
cDlLP2W8xEBhEY17vKidimJA9D2hrVwPEI8x+dPDkEVDEIr5FJcWh33y67AtjpYvutXMZhSFvnrX
KqChymmCh6U33OQZo12utLECl0I2ovO2wr9iPr+/b2gg05in0bYwtZGTCobvcxBDuBz8Fkf0hnXC
S96fvcdcSGZBtuh8waPMVzlsqTHg68V4C/32WHM4V0lIRMNmPr1dhweJxI23uFmcAdvcKxeF11MD
th2xcux/xWAYzje1hoUIYaOnqooAVlkBurXwZffcd1+b76wrQUskxICEJxvnoRIVaMi39oY1yDzt
gUOMjK9XUKzIGHWGaWCTuP8UlkQPFhwtRtEe58IeKT2vd+s9HOqo1SHtyH5pgZK50pxcb1jnmthv
4weVDh18ntHsX0Vqx5ZCQTG2Y3xzGLs1fA7AjipIWMOKCtrHQAu+MsR5cY4xdzGQJTSPNWKrpnug
TshfX+FSQJo8Vxzdhi+YVNj7IUttoRF1po2v+5o80pSAX4tYRDA4KipARdp7DB/JoZj8IMxJ0T/+
XbQHdlBT11u2/Jh5r4JDWw5AE/Ay34PW0zet6Z91NMmkhwb893dsjiW7iRjrjfUvd+tO9X7smQJR
0QXgqCMGwdfec1XkSKTzbUVJI4Js4Y/kMSGzAQuAuE85j7RrOp+as8TjutGbnQNr+/tFMACHk+hK
wbkv0Ho/0IWjRLe92G1mGVTAVPXbtllyVqmXZiU7+BiZhLxi4hQlJDl86UBFu+4+Ow4bljQr5se6
wzYMi+YkDSkZN4AOuWG9Rn7a58+PPt+lm8n1QCKZdmIapuJkJaEetlME3Urd3vGdoTsLJ4ScTgLE
BaINioh78mKT8nQSADhjwwHMCJRWhds5gWoVNJiugfR3MmadgH8DG27aZYBL0cXPTaVE9hXfcou1
5SoShz6bYRv/0Pax5BmJMCD/ZyrFaCInbpqJFfrCc86Rrdqt8iZniL3MD6Xfr7hFjZd0TpzNqX41
1iOGZGgxgGrVGQ7Bl/nZckmfzYR2hHXC496NNviW3amTTHyIDc4d+oJxaetpKXlAm55zIzQx/jqr
oMCF1AScSZwWzTnMsL+viwoojdYvIr7msMx5PgCfDIWBeaW1AwTaH3jnICT0eAVu66gXqM3KhI+n
Z2+R/2DlsLkIroMHJxowNxl7jqGPnLsF1es3HHepAfMxLKT0/EzJ8MDOocKMkTKsC0X3yT/M3/i6
z9pSE42Wz0unCd6uR2zRz30wFR5zZdjRJwqciY7TcT1ujLeS829zAKN1/srsRywzUjOlMhwfRe4l
5v2yW6jifZLP8FVwq57sEdDqBv+GqdN4qqcPJWLLSXLmd1S2ipfNUA1QR2EVW32oJkjtBvt5w34a
mY56Bp9RLQtLUMvbxpR0ZpxBwz5PJ8jhStkPlYb3HUW3JI4kcd40Z2P0VcXbZ9juI7CPw8waYDEn
GQnnPmEybR2AzMntrwGMjAKjZQOuiwj+9immNNVzRdsR4zs3MVyudiMPx+0Dg5ZsbMfcD/M4IBEP
YfU6O60gcY/zSuQXImlU7VdbPZfilrMurPXTw8NAyHGfZyo+yLMkNf4PQkMy8+ejcEHqR7ItoaXn
h75cQN18htkxIn+cJ728vokJ8vw5itVmnkcgtm08CPFj+gSDL456qmbtbw0i5Z22HO9G/XDD+7y6
5NMJZ+Z0csnG4TF2UNQd8EZbjOS1JgR8pTNNrVJ9BpfB351gi7tNxSlGYIVp+5xGAAa3o/FLeUjQ
AbawZ8dy5Ts5MS8bvQBz73N9/KJJ0vqa9tyhGD3yXfFvG7oxJ9b2+PW7arUSuNLjiNOqAnqtpQQj
IyB6ZSKq+9cCFldCTBCD66I6Rko5RO1JGPAKxB+tSfcKmeA5mCrZ0pALlQFUBzjvyr1FuUd4+I7Y
tDkF/FwR53STOfotj2vCH50hS2LDK0+0XRUIoSTQvXqwU+tJrkU4l7FMdCNfAMBtEXK67K7PtJ4o
pQMKm6Jo7KTnlYjrYMoSKWOhwVrYogT+vdWLbbvpUpXCFF5+PbnI4gqsAusU6zE1g1ydXGWNrOcN
y8sXEdDSfKWh1yp4ZZejw9gNPHUNPFU/QpbZGn/afoq3RZBncJMepLPnkmthl5Ohno8NIFNVbruq
fo1VT99h86bQ6HeMfL4NxNY+t97rA9QANqqwMtGLxR1okSfDkmxDN9ZAqb/xI27g8mbUpEmWO6z1
hVv4umqB5G7xu/XZLTDBvMiNfWF4PoWFgBtfgLtdnYM3/Fd1+BiiIK9ocp+thssONnI1w2rSJADr
VHgc8CZGsnuFoze6WqIrDdWg62oa/fsd685DzYLWe9D2ARy2xhFqYTF6Bd31SIn5PmgSg8Z+s9vy
1m97TgvTWjSnzFNnIZHriH9E9Dbed9WA3rtVbek2YirfNw010JAH37aw46SaNCTRgbNGQ+xsqNlW
sdALY2t/ltMNkR1pUSCHfy+VuMs63F0tHNRpRhVSPpBKgHOhFbAOA2JN3VDTVj8Ls5W8Rg67DZg4
kVy5RLAgp+T/23s2cY2xWK5VzXGuTa3325M/qAOh+BzmHIawuIkuYy/6dMst4FfHw/vRQX049naG
edMi0MFd0VmnxMTRcj744KhjSBTpKukYE04ClRFAGVZvTW31WVP7X2WfbHiiDQBryolPq85nTvqB
WgZ0TKV1rj1s4kIFo5l+/5vjCHCO32JpAjvlda2tG5Lip0THvBEiFTcgf3UXwqlFkZCniEna/3+m
d1P0Yv2PiTyhAstsyFEd/9ADFesMzjAk/2X8yauRTO2vvZp3JSeJBfMQ73TxzEB8gubSUchELJMb
BF8fbpdLCvRiw5niC0tZ7GANW0x/p36zxoI2cL4tOHwtMKM2HUPBaYIoO0RACzZjtk7MXMsMCf1h
cp0YASfJ40FNA7l38FoslgBhberSpKRlQijJdLnppab6nC1F5t/LXHH5Qc1KQmUb0NNKuIyiHHJC
qurbJiuhFV2vkhKmajO7BrouU6wBZRiuht+mKe51flhFc1WBE4qt7VIuET09vjSmFmdvFrPFhWLf
CDKqhGJO8JGdo+9qOdWfO0XYD1Hg0qdPQuusoWxCfjR+/RlAOL6j+8ksMVQiuRRE0gpyJd+xmK7k
jkuOziXyZslf08Dll6v+SVxvaBtS8XW7rdEN3nVjMN9V8bihl9I3zii6uVB/8bItkHGds9fZDG1p
d6wIaNb7Nmf0CwnqGgJnoWOBjzHTahmI3WKpZYkSQu6X8HqL42trwd8MJlnMuRFTB+G17+WZRwCn
z1Z/dUG5wEzaXLeIF1yaaR+zva6RYRIa9RNyYmtdn6UBoSzEdZ2/PwxEBscm/Q8Lg/TB47Y4hixO
lW+PPeAwfCcxNDbFWgzh8edABQrQZpmTEf6hJTasgoKgpOM8N96vRZQwk21q2ead3Mm2tDZHQHIk
EnMydOt25YwMw6IzSLhN9bQht8W0TyDWBE222oCfrGUM0wA++YJmmkDrQo7z/CNmqyQcMxV2TJJj
dhuZoW7Hyqvq3l1MwWfD1kVyJm/D4XR6cBsE6XjKHeb0QN3kRWrdrJi+mYROxZNDseMcDWS0NXUg
6Y+4AQRQwhBlVqMiavdb8S3J4hFY15d3YZF66d0Y/NX0RWt2udYlUtIaeKr3n+tgFOSfvzOyLjQB
OEOXNTZ6Zm2BojFo40O7Eh9xHDPXn6zjXBhzAAJPnKlzCi3ED732kyLTgipkmiXw8WOSaFVe/gcA
aTakb3KFljh3J+OCbEYHT/kWkwvh/4GGsmLK3tlO4lQKFNKktz/IwcdvDL+z5nTZLSO3Uw03Mk+j
Jtgw6YHnMBlrW4wP+G+BO5sTErxsn9IMm3bdnc49++h4I/KYfDY+S8MMDoa/kuPECL9Ci4j/Dne0
s61m7Y8MrOIlLVtpcixLgDNEJddJE6FrsF2N031+KbpXjg9OlZw+oOs2N3GPqjYSbI1+OB1m0fXH
dNPbmN4qBP2i8pw2paTfbhDg6X2okxU+Z3OuBRauhmtRHvGCB8tArfHTBO0oidwCOA1R2xdM3ZTw
E35kcN91kf3Ymrcj7U4f7grkyxJixL85axnRXPUTHfew+0GZ6Uvxr6DVmlAqQC30nK63e7y2Z9iJ
P/hcutzhNOig9bTwqb4ShxeP3rxexGtP1Jrvgj/PtyFN0j3wevAV0tnZQHD/zKCPgddw6q2T6EXr
p13RxVz8sNYQV25hermHBoRCZyvFMp156xAmV50U5o5EPpSZrErW1BYe1itHOH3a1h1X+IY6kuSo
ZGhydr4QsLUBleZXVHcSIL9MmGJC+OKhTfIuE6avkmvVha3Jah0nZS3vGRjtIm2Qui9kIvjrA9Fk
/4z6F8Xj8Y+p6ZsNZwwLJMJSKflBFmWmM0twsuyOd5AcQ0fYMF03gRXyXY5Aus/VIjuajBPvPXF8
eCNDtL/WCltde2wPA1bEGqPkyzPQ+KI2CcCaoo6MLTpxRrk4bDmHKkHUvn6YkOhbk2r/1/Lw+NKL
RRdu9BJ7LUkSFx7UJk83MZTFG5+FdWDBz7G0luzzMZLNdV/TrPhUamJWA2jfK44B1I/8epeCz986
gWO/c1NH3GJcNtFZ57blYA84JJqOLQptce8xgc5osMfvPQRploVcbqdqm7Gl2Jfk+xg8LytCQJfj
oA/HXLiX67JchYBUsEAE+HjuxbjuJYQ47HEcHfJduvgDa2EAquZUu56CGV0eo7shsoEAe7CQfDEs
91Jj4lH9Nb49917eMmb8KiRxdpDwjrDJ+nL6i/sfvtffk0dDhNY+ZYLvvrFcgawQIRlJ3kKdY0bg
TQWhOJopvPa4/naDPzqrirbFB41QuT9cbotR91i5zJbVWJr3lFBxGwvVAHdsCjFpNal8bzG2J6lm
i/b01N8kewKVeQUsiwCs6fyHx9jgqk9oztWCiBYOTdw5BO6r5HAuj/7wfBRu6viOvRT9mg+UcF55
77kLJ5YXt8xzhNuBOG6yTjI/28gmPVEEPQrfkOB7SckheyUTMRCq6+Mao7TZzwwumpFlpKE7dpYP
eLnjmjumv3A7KGbNzekUsXFqwK/2RN++2vux0RwK2kltDtFGaEcmNKhWz3Qj03FR+CtulysFCOyH
Wn2mCY/t+5PTlY1yKlwxDU7Zm4L5eAg+18Ov+3BBqPhMtHneC3xFbBsnBuV+HuFzVXeWB0iG3OM4
/sgMTZL+FcPIm55TntLjkKC6Rzeua/A7SJ9rrOvj0EIteGoocusNr8imqtL+A2n+iFSdfifTjuUi
iUdDoK9yubRd57TGImmNn133cgmVD+xMv47DetX5WliQ9ThIYpiOkRpyxIHI2DlcXUf8+uYQHAor
ajkGrlrg4dTlsukqEvjkZaSQDhRPUp3ATk9ihhIVoaspA2DZ1tx29dJ+Z5OA7KTMpdxlLjA4qUtS
lBN9ekCnUOVlvRqltfk8bqbikQ16Q1W6VpelZecTdBLXRKE8Vrxqb8m9eIg3ifAYhgjly7GdbdAO
bzKBgP8QB/UhKjQRT1IK+VxbCUas7UUAUEa3o7OorYLF8vJXA5etcd7nYew++/r9Fyl5Rq1FLn86
rFFRDmbB8Nvs6wvCzP2XhMeLUM4BEvf5DoVWLBLoEVYx0L9vVhC+QONCo5Vr5PLxlevQRWB7qVUU
ZU87HFxFYt4tbWRmihILLiWPtoMkutCzSzJpo8TrHwioY+JOCugFviIQsZQABlYoPezgDvw8vx2c
nFJcC49/cnfo6CUEF+Y6eNuJB1cfGxJB2baDfKcVDjK5mtYfgT3H6nmpIkIujfnwH9qdHNCgVqSc
zk2nNEF+xMcZuXFhOVvBNFc4S2wnwi6MWyyECZd3YN7virwtSkPtREJ6H5QB3J+uvyoCPQh/JQua
A/G3NNVlUeB5ZKl3xLxj/fftrxTDKl0fXmiW3l4daNeAYqWHvCFr97TZ60V3W4s67bs/ttDLRNU5
wD51ctX1kiMvPsDnPqxtJwmJ7Pqh89VPCKjjT+ETtSpZB71qEv5s1A/iXcTTbP6Ob0xYfwMBygKG
53kLnDPKG9UrxmXuoBFKdRkROweRpHPjNKayI1l9V/ORaIO+N3ZvQ3GLMv1j1VjJffbanccVaIvW
jVPjnMOBdyOvf8FjUsnJ6t9xB7DrsQ7LYEt2VvlcQn5d39enDUSnyOm3DwjhbzedPv47kxZv9k3s
31pP1o2xbK9NhUDbO1YYEfaS5/i5O/wCNsNJPCecBXW//Ijf0Iia40ZTP6if3g+3zFcLy4fkVoU6
f/TFmzP3vMR0zAXDGtjJ/3pzuoxiJmgCm1XyyAJA4LurLB8VevJ/J4rZLtzwEERhB2p6n9X99Joh
9cqEq7oULPck6EFsz4pelh24KKQeXfD5/LZzJJ9KTsdjYnJmozsf9xlqDH4ewquVsv5Q3sJicJva
61VRRtloNd4jxlfpzSibCL+meIcvSBLaA0Lh0AoAw7tGXyvUp6msiMDJCGjUdo7O1fjRMCvzFVdD
bpe0TnmV/piJ/r19m4ZlldiJLRmVP24v6njzWryOK22pDyZDWxxucEAsHcQPAwmN/gDpTLIsG5y7
DknEWAzqAbwC2JXNb5j44TXHLw4KwFm61rOna4Z2qcr6DSjda0mH+XyLnMXr5S5dXrV9ctANtmSi
DqhiO6YnHRc/t0BbYSlOt6ZuM0dQFjcn0JmBjUnjdno1KZmpIJ5zJPccP7G/1lwq4jnmLIGw2wtj
bN0PLJCQi8O/jbuFBlT3W5rwLjWFVB8oZrF8UoIISib6VJf0mHjuN99tHEMYQurVahypMFjIabKG
N6O13NQb3/FlxcOCvcdnikOweEatFyUq1dKojrVOYTtcmoh/Bhpwuujn8qADlOlV+sdjE1zSlcFK
dgAVBbec5QwE3xm276vvVsjf08DjcnB7ZCZF5t7vpLr/0pvz3QbhO4VLhIwTe3ZDdCh3Do/22H68
pv7WXOnMa0BDjqrHHp05t3NyGenfHfFeqPRxqfkJFZ+mor1MB9+g/UNkZzrssQwJR1eQpYDLUF8C
Pkj3auL9ryNUdfMFg/kPCkoyxYgVsOdtfOX6s9UmrwPxQQB63RW3sXFEyXRFWPvAAM5SVGfFSoMy
5hJBheUXy3PH2N3qiP0ku15Up429x/JPK7Nngrh8fCA0AXgTJd9e7ZCSMqto9bWG/n6yVFnw21Ij
594x8aDB4oYOaVcUhE0tyjJMIjveP0ZdryBEMc8qS7C3cNAf5BgqSOikr970cxjVF5o1SmWLqSav
kQkLR9a+4AmX2Lvsxv2UmdlJ1mvUhpg8noG+mObXFaxoZOjKdgs5cs4TJb/CPlfU8YcAKqAh0ow4
NETGm8VZJwEYcsRJMtHOPAM3U9NuI8HNCh1VolRX7Uqmky6O9oNiz5X9LMX0i3a76yZRmo88rG5G
sUngsipoULcxqTBjQ0Igh76yff6YoJkEYVf8XMsmIzxpgivbo4ZyMlDZtGTw3A0J180gHaZYhwya
U6h0ilQI6nkp3//DPc6e5OY4PyLXLRMRO6fa3AblfV3nEV9EP0odNjfQfYzaC3eqwje8cSABtLEE
qOdecDMx9cWgaaQYcxavZPTSEKdYmbu0n5h8EeL8OFiEO0RG0gfitINGwTqmHtLaChXYH2SIBccw
f5UcO+PjlEco9q9WTO1vN2srXf5LACYWBhsFo2Qdk7o2NrLyd2LC/ZTWMxvoErpybEdcchI7Tamb
S3+5O1fL5edrx34CZH28JldrUsHfSShyT83fvq2sLbtY+fsLJCtodwY5sntTC2Bg5gue8+85nfU6
XuOHYuiswVyYBfvtUMcSv+/w13xgi0TjmbawTnv8IF1WudjmpG8ZcmLBbD5PNuBFp8bbULdHgmpL
We++4pISBJqUA/Y1QfXvaskS/ZhaFJIsw6nEpkR3jhAk951FGKirJ3MaxcQnWicRZ2vmtkaVVr7H
4HqOfQLFDdCWBXISyQWB0YdS2I3gMfE16cSzczEq9+pQqRQSC+AJRGQL+IRrXL7jABwIyXbmIEo0
KR7hyYvhB6C3tZWND7jd0pTyC8m3c0QRgJ0q4DOoAzJAQ/XVA+OZfl7t18Dcwp0WFWQzxqWI1Nig
u5tgOkFfjIiAn4fNmiM5Omj9poMMz+s0M7hDEqWGaMairtSgE/YzFfJ1A27mxduo3AZbA2OcspQb
+tF8ke8VgE7vbeKbK2jqM2TzLCoTHRKHBZaEQgGKAXNxoIzpNQwBCTUarsWiJpUaMEkfVSXVuCkm
k9Q4MNkxiakl33xEAGkCiovT600F/rEOSxxRwx+6b95RQmXV0Hi3P/WZsS6DRFUhxLd7WkpnkWep
9UEi+vkxIMpzLwtKA61/zjVCQbApFn5CT15Wk0W/5Yh64E3An2KBQ2AJ5A2MeXz0VBHNg5vTuaFk
aHWZApbn5Iv/q3OyLbelLXoDIJuaBNVf0CH2R4j9/tJ0IAeIm/IMAvtgF3/6YG7XMrKeS9BXC1i3
WaH7wQGJv5FQ/fphLhUqvdqXzZ+6yaTI68kTm+N0tLMyHuQDFwTGWbAubCkqDWmqqaIx9Fqo0uv+
2KRwrtgBWjRyZhWiLLQdbuVrSAQb14HiIEtlDjabL/aeLvpUrw5v8OQyNVCngn00LsNJe3ZjUWZU
odb++yGAdTLvNAOGHSywN5TfujpPwlt2mPwlYIPfAcmkPqLWqUT/PxW2dZ31GbGhPo942aN04kYI
YxpiXVtqjp4uf3si3DJYm9770fubJ9djy8RgyprHovJcWHIXqW126DWo+0IH17K6aI0rb2s8eh4z
+/mmrp2bt4ThJdsvgDQPdG7OD2aVTR/YDdWPNao06ts8jhDxjyODUNpDw4MGiiiFA2Hs+2YRbQFX
znGN7w48Ft7WyecjuNvZ6TCI/hMAdwmshhFx1zvvxnN//xe1iCKx6czXHDt+h7RduktTIbz0+Zjj
iMeHxdM2xbriobb8JNJBvVz5FOMCgfdU9Uzs9SXFS06yX6LtECziposSF9sHCOFZLA2uxuhP01t4
O+kE7r8WSJMhc1jOIbqhm0tVoWv8VvtFrhlSc6pzzXa4DbMES3Btp53lX8FdzORsy/UtTwNrZynU
NaIEidKerRO/bqC97ied7fAYyN/RRi4rmCWDcbJ5Hi3CkGK0NkC9iGrQifHke4CfyM5EcPSNruvm
Hiq2ujjWypqiGkchD7XgANH3FFhZXUWIqWCozft1ILar/lJ952OpZhQ5F+AOeHDbGZr7EcVLX+7t
8s6FvWJvZ4slr4KmU6ZQG6w3sSv5PqonVEMbfAbQteQAgeSLLrmeyeygqKAcGRkhJ6rSRCs8uyTk
+MBl5N7E/0SnnL87Ce2urrEICG2+WgU7mtmOrEIYk2KZIQHrkDHvTGbddW6nSuxQQJ6pxgIcWzVB
ShtX/HmNT2MpMLQEmJBLiWTv6hIn8qbbJln8bjoeIsVrCm/n3+vXoh6cQp1gkBaJY6SZ9qwSoFV9
Y950BFaBOyr+ErGvCXtGaXfnlabNNiYJBxm1wDyLegYgqn/2CHDPd4xVNeeMHv+mhW4fq2S1hovw
kpbZgk/PFNMRbZeQmFNxjEn1rHBINEzLf9pEFL09Uun8sMQAT0Ie+f1TnLL7quY2+smrSByu4wyR
RTEnwuWv0QgincP0nCU3UMHnwZtlAtXGEG2kI3xqPtt4JzYVnAB319brlShcXtrmvoysDVphleH0
QgJ9xmJ4VhpGjirkEM9LoUHArXuOYga5f2fIZFTlvO5icPepwnCHd3JATnxi355a1P70Ad4mtoVw
AigY1oQ0dmlThxh4PPBi6jwzr38LcGyrf1D7bP5tZAZqFvQ9bgzkqwFaZoUE63NzokDEYwjHPm5A
FadWZDpkgkg+x+wlzVD+LUuPbOtL/Lh/JUuONgP4lY1R1mrEGU5F4OQgpnC5cFBzNB9P1iOX4bAQ
2i5VNfBi/JTry4WtseWeK9LrEDTfpQT4nwXz5GyvRbDpKVhwEkC8PxWSsAmTSZ4FUQ58Za6huPeZ
wuWng4PWZ6KfvKu0Dp7hZKDFvyI6mXliUVbxiWPZk+pcSi58+aIWEz2WgGqZzDbcZRVpDirwyIfc
tmUOzCFTQVmnql1eFLt1a9y5sLdqfFl4lcewS0vO/3S2z7cymt1WXokvDxxC9TpU5s3cY9MP1xBM
I0Z8YVCH5T6XdwBvuLlGSNpRMMJL1Q56Sb3gkPKD3ONY56gxBoLz81n7iyWJJMbKtf0+HCWIYWpC
lGlkTOejxb14f1ddqf7BMWw7KXHDjDIdfby6fqi3ipBVUs8ONopl2FmFTF1T7KzYWsn3EVPGZH2D
bgR+9BSQfZGVOBx0gIvmzuuZ8tKkw6h8b4FU0Am3M/CgAfZjsKGnw6Y7pfZS/j9g27SpjW204bzP
1Oz++IG/k8gTv89sRLYk8Y9NezugERmaQw70I4Gll/AE8s3ss8fYF9F5obB8KzonfY6HpF8WBnXS
iYyiKkj+4LL0SSpXSB6vw71ykWtvcGhIfrSE7ryySnesysEtZQiDJD7TWUDY/0B0XNnli7KfPvbO
w9Wc6qKwzLpd4+1N7y7wRnBKAyYc3roIL41gvC7+cr1g8px+J1Gz+9ACfqwf3diJdB/ckSmT63jz
p/e/77bE0h4x9D+oDTUb1luP7h9QB/prUS9sBUbOjlDZjFmBmExSvy+Li4K9OKhoRpi2vpKGh+/g
kcSFemaH5gIWYH6KCOdoYCQ505VoDX5FwE813ax0pIlU/QfqCZwTvwNte8vStV9IRS/mhMuwVb0Z
yAPcekAnykw9WNU8xFa3/BpbHDsUlIJMu7vZrqUi5ZNQm7SRB5lIFu6/D6K1PqWlu+hdU3QuaVOL
PxqM4ZY3vqpTCp0UDgfaWswvkvX5zT7baeoUrhvKiRoiofvn4VY+MtTwbd2T49sTfbstCEGsdVZX
DNFLwkn6ppQVmA8pEttk7Ee28dAfgyXL+uShsRSoI1s1f9tNWlSIy35Jo8VceHP+MaQwSWcD3htZ
IhE4GuqjIVTRE4V+xJNybrQu7Jn0xAoZ4AIR9hACi7BjU6GkWH8+2jZYprOKp9J9wJniA/X/aD9A
BwhZlnskbBCgIq+xjnCpFl+11yUROSCZo9SwA4VoCnXermJR5lrNAXhoBpk1vHqS7u0XxJRD4G7Z
/7F9nfXFGq8M27QZkGCkAIwCvR+AfUgUs19/zcZ1nvTg9FkDNqhfLNOxT8lFZZl5XiUAOsgFU+40
06ixBs/gBd72FxViGgoPWsfPdgklLa0+APR73RuRFsr8tHq8PSLebCjNZ3+rLBxjID6xexM7NQOF
VUXlDJvDKSiBgMbHjHKxTl1txUYVdVcoqDgBiz29KGP1MsIfZrLYj08IJ3hZWGQBSm048Ifq2Som
AtsAxLTdjTdsVdkGtEq3eFF1YMSfrb1QrSHwn/e/laNw3zI9mrgOjvYmprQ3J/jS8axXSBZSQBgX
y6fJftOJXyxsByYHAVrgOcdBQyhARYzLOTdpAInSdhks7K/YUk8pO0YFwG7Kvaycu4yqc951HmXm
4mU3jtx3I2Tf6TbcwzG7aTKfwEgiiDk4bRw4u/+UR/bVjq479FqVUsBlDEQN/+UTrsd0XkOzoXr8
NTi4BKcYd+DEsyEfTA3yj22G7ycR6hyly7liAUHcyxwl8hIBSjTzpd+00x+o6fmVZ/mT81rYZ88F
8yYzPqX7mpnl3eXUgMNt7fDOEopCwIJiVzgBmaTlcUNcVnYvG/AmQaptUEoS8Rt8oiF27XINEqyg
uzhWifFghNG6jrXqzU2vqDe9JITpyJU66yq+ux7CubFTFnj/BGcq9ueWLNDjmon/sFXq7LT7Qs8E
y/D+YelP0n2OQDGsXCBDrzTsE5ffEMWuixd5NZOf4vfOm1qWFip6TInp9OJaLDjvUX8LwRGAGAB9
x6IW72bvCptKYCVb0eTsT6XYw3wfD4qLYUBnL8nlu4uTVK8QnVC56C5QX+Vi2vtKQC6NPOLww2Gs
pjuuyM+Evoonx2YvHp+mV2NXdFSNmxqaAWRuJiS7vqL5ax42l4kCrqxQqQKgp5EQ1t598PnYb1T0
qxx5FOup3nsO1Z/hOAQ7mIh6Ij13iON5MyMFgPojck5jB/AtUAPFknrd9SWY6z/3MWDN8BCK8MgR
BBXkpF4NF9nvXPmWMpBhhr97J0PB381g1rPrBzJt+7M4ipqc4o9bRubU6EFhRiMGpGlK8C2j+1zX
v/ttWVQAPE1FkBw3Wb1llXvm0O10H0nEwSHxNcmPstgHWXzjMpyzZpY8vXXRyavz1H5X+SxiJRkS
TR7SD6LwYv/BOFN581D7a1aB7w2FOQ4A+ErJtjr+97FMmTwaJcAgcKlFIm10lf1zd9NvJ9HdhFUu
rdCYxX3IZM8fSieM2IVOxITgK9RqLBWj2gKQJ72TTLRCFaNSYkullO+6kSHNijR6/klR0Ywnr9BE
Jp4Lqf2xmCpXFi8JFQFhkUFnyL4kmveq9xtXR4c3w/E/ch/RONRCafbVh88vnB9tEq2iXrbUuQXq
a/P+52QtM2xpbMTx/ONf2qAAc8Ak+VMQox3FMR8S+WiKnTpNibSBHww2LT5RzkqTL/VMXFlacWlE
ZX9vePnqyL/246l4Y+Jele7CdoJ19bjRRcKlvbH9/LAv1oQ/mlHlRiT3zpHasDsvD/30lS+SFBt3
IxH7sPzv27M///Q55WofdbG6vtZ0bQwq8zFZoVeyK2DHesqbLhkbHVynoSJrvkCoLOJwrqx8KdYr
qxdhHK2mnY8zjaq21A7sfRDJ5Ac8O2DNkl94s7lkLiXMhtTMCEdOdZdSMN69SCco7x7VJRo7RgSP
HTJn8uXetjHNjxbjxM8W/Gijgjf2JN/edgPlM+KQga/+ZTEW9Oj4bVB0K7McGYoFwNAXeFpO8LrC
cZiBf3gktiJuKbw11RAL2L1k+wwkv1A4wQeuW6iPSBRp3k7ZQf5+kl3Z7falyXyIp66L3jWw9TJN
UDibnTu6FaHn/uIbji9R2iMb9dAUhTE+Y9EedqpWi7+5nhNkLcTxC41+my7FQEIwP3/9TLq0A/Ow
ic0WedK1dynKmKpiOL5pVfDj1SG0zLBugVnK64YNkeDTVtYhwxZ1ZpMBQc2HDqx0lJrEO2559J0f
JMNrolO0iG29zOWNdCbSendu7WuyIzfVKPCjTCowwroz6I8Omr0SubnPOEi0qAncnxSi4IYNaiTt
JftdJBQqmBD+vbKXqkh2eaDFnK0BW48TfCNuQ7CbockjbwN9t14ZDJeO+wPfdfwx/NYnZelJmS9H
+GAGrw8BG5ovBfFWrq8Gi/tzFHyNulBRC899Mehfyyavx+h/NEaL0TzlybkMNcu9az/Ov/2ynoKH
awp73J7fJN/Nw/3sofA2cVPbDxX0W1ImGZaKHX2t1PPZBfzHhsDHskdyaf/SbfyYM1g+FPJGAuLa
ThTXqS2esJtbkz9xPpqDq4lTQlUCb1HaOjN9FAMNmC9YJuWWOUMjLJr01kqPW7l0c+OgoqSsAzat
oldXX6pevsLOL/syqwbBE+m/aQHn++7/PpUbJ6GdSWhTT0jDakXhSoqTe5w6dT847lAmtdS4/l00
cj+eEbNAQarfLOyjr4U0PKdQxjVYil1sMBkUgLA5nF/PBGKXR0SFkjk06EkO9hosai9D2v2Gkj3H
l1wrxcGswq9LzrahLSiM8U+syLZ4tGjC9sE9xqIXzfSB9EQFpUFWRTi4rhTKNUK4tCZUWb9w6pfK
+xr5Ybl6E88nII9YScXkpLbJZ75+Ra279gZtDTs/rtlXwW3blw0tzo5wB3uHC6HmdNd6Y9K+oDM6
Yas+gNFHE4fgboqbslqyBSsoymXfzDnxbw1ZE++JZipnWqwfFt60QE3/Dmep5WUVtaDhDKHpszfW
Dpw6REfMv7FPGX0HZMzP4tWem8a28q77Q6rGAf7gfeoo3jzgKwEswSeuJbX1dSpQXVDy2HzAy0A5
wVUwR6iv3FCAfyAq2L1dpoQEkgKMTvtMGb0piALsyzsSTmpNCyKdVl4MEe/uWI0XxyoC0X3Qnrwg
p/FzXFQa0GQA2Dy7UEwGr7F3F2vCOfNkBpPnWzgst6m08WbOSrzz20Ex19o/r0qrkcRLm0F/pym9
iEwZdYFiHpa8wqE21F+dRj7v8QC5JOvFdeQ4RPXEqj91WBOBDIO1izmZowJ6sOh7Ev99ontrtGWw
VDjKWHPYrORmpfXhP51S0TtW63KNaWPlKKHlMfhaR3nXWFF8ovUmNWPoNPMR1/VkO9Db2tsf3VAV
aYen1pKiu7NkngpJloSb7K9p6o24LB7UQqwhtnRLZZTWes4mljU1xG+uIN2dekb2l3IDzpm/3Tq3
EjPBGOZjAoRVg5X8J+XG3VZkg3xidx1hemZ/9RlcGmU2Fv4524EwEg+cZMCfaxSyjCQVwEbOzUnx
bQuYdFXyzw3RCgHSV9RUM7QhZ0OG8fuTWwM9dcwbVA2Xh+Wo7RzU8vqXM7HtHwpyG05215Y3mnXr
mbr88KNLcrvm5MTPp6vzbT0tHXb8PpApYqsws6RH30YGZwF43ixmthqc8vA3PyEt3hoET2Wc4woC
dHYPla/HmDaFLRpaOUdcvuM0fZ6+DaCndGVZhFbWI7X7a9n0VMyen8wSuvNk8ok9cl6wkfdJegIH
JtBh9Alz2z9cSjCBxrmrDtmvDSUyGPFtYVMgrzvvAoJ13H9IsoFXsMWbPYl/MpUS5RdRpVXKEcls
vEh9XZtECfI1zy3m7QP9LqHMqxPPrz3AK+4xSMbfXxpG/bGHL6Ur4e6wNwAH//ixiBTaandk2M76
7/6wTO9ADKIZPhWgQOtkEhHp9Z29fFcaX8BvIlld6ff+wSXX2xffj9iuZT6jbKQZaqXUv/1NLO0a
mTFNeSzUyAuTewAsC7+HFcN2n4NSaftJtLF9Tet0yze9zwNsshgiA775qNyLyKs4gavCi6XoZLIO
nw6gJSBzSSp0Dv2tJd66H3c91FuJA0DZuDpwo3t+Ks+mkPQdenqzSY2gh+BcHDYScyYxIPe8ewl8
oGtREqsvuO8NwIduPdXzGsBCokTNMhyKUA98VkMZ3y2sA8x9ot9HICkiMizz48Acl23tNmszhiHu
a/YFDFZnxK2zIJaunu1M+eKzlRys6CmtDZ+FJte5ih3zlUDBJ/WN84CUngWrifpK6JvG1iWbiCn3
iBb9NxGtfDmA4khUQNzcHoQf6bmMlW4+i5j0Iq2hesye3JDtzL/pxYTf3FoZcXbXpVskaUsApcod
0/odkiKIksT2YFVTyFGgly644fRgiY2wcN8cVa8V66xYjxGehsegX2ISEKXR+quwqfBb6zFiDHKo
HEX5ubhXBgNG8u9qUxKUIzz4nlNMF8qfoNeJftC78Zth0yUHxr9QqG80BB8qFUu0lzYLLomPNBgS
0ivgEoeiMBcFv4bfs6eU4AkpDh/bCkSY+B73IRQsMwQvfKO8tFbNByFvXsaVzJHLIoBe6eLvBgvW
khQTshFQ9DLNAqb/A/M+jRRzJ2s8aDEc2Wk83HD5aasUnvKXAgSwpvhyrvPLmJ8WIJy9gk7rsbO5
P8JoL/laBDfrc3WTX3+8gCR9acAtvsTDzQUTHueVjv2OYd4A/ari5jpG8Lcyuz0JhdEzsCCMaueY
U981JAlP70MnsMrLoxWjeJNXAQxzpCE+VESigVN4BlQJ3wP0iw8kx+ABpCC+OmiMuqViVoyomlGF
R2OfvHe6EbDpA+ViPcaTZpyI/XD1MpFBZKgeNw0uSAfmobQbm8Cnz9/T7AdsAGDiwOmRUlNnpJTk
FZKNZMzLcVsqlmOq5tgRdZrlV4lK/rVH8aAHOBU8XLAVdi+h3NTnxiS4mQMdK8VLWZj7sZvECtqc
2jHINPzwQLXWNwGZeFZuLZY7jXmXbkCdk2FRllZpXgLjLD28f/ZWf5gOiItZ2f3RzSl/4HOWfMCN
aHQ03P2aJmV/B6bqvj1pGc/i7Ut23L/KQHfYuT/526yuVqcFQQHudn+cvN6SiXB4jqyn2O2UBnO0
J5xowGsq7FoqeMiSWEiinVNeqPfwrnXZHeO/E5Lb/0xyGEhYFT2ssIddRL0R2v3g1e+YgW/wcQu+
G70sJgI9runpSP+7NG6vJsbt5zNGfI7psR4aHg3tMw6SjHERBCLcIjTZ0dHiFR8sQA2J31pLzPHc
Y2Ub/95EI0tUw21AAbLi6Fhp/gx96BrFjjwPQuXV4CcjOgBXz/lBSXF7qmJcQaVtbMHfkcusDx/o
ofVA2TEGkG6qgoeQ9fqkGc4z1Tn5vxbvW4MnRzmCfoMx1R4v5NeRyRpFNWtX3aP5/8r8iwKRG4S7
BptZ8Fjwiuk72EARuL2ti/ne0boll5uwqueDlYMieQ4GPwO2rU7O1lU6NemQFdyP+97dnj9vSh16
bLfEtAyPBLcUWAl82WfkqZsd28boG77cvd7HOead0vUYfv8fYyNGjIyMMk+HCsGXdjPaeb1jyjTp
MCRSBlxORmjArxwD/0QNNHQWqPOQR7RThoNgAQ4cztVfFlOAWZfJ9LtEdQ3Sf9unSF/exL/Bd/hh
EG/xxe+Mi9h3gM7zERBJ+aYPO1HdOoMnLGlpxCtN3anwgXPxRlaUPFFkzOnlIoYaWb7OkCFjX7UE
V+ZPCtPYVm8qt9qdLrqTdgU9T9v5VGfdgft25/w7T8VQ8AitB4Qfevfr9U73umuuULw9C02NyK9a
BiQae0ZyFYAEvcA/oNzVBUNSOFYnep1afcsYnhT0uv7PcMuKSEWzgpr4p63DPmw7L2K0boCvsx0C
+ICqp91G3iKMlkRPi+r0A+jJhJWGq6VlzFE8g/jJVfx/h3laKiwyD706XteG7tDCUh0qRT431FP8
g0VdfU1+7UoSerGiXHusUCsNafzP3slB+/NghTJixnLvHJ1wRaBHNGhXhDoEssPr8KmX8EU8qYoY
fHJF/J1SFnR95xwvt3OG8M7TR9yHLs/XxMlyErFPaRmvBwv7X497fez4kLWEad+HkfPyd2s6aXv8
D/VNTXBEX/i5hwFu7IdCBI+1K2zbFDOMwUAOLFxN5/ejNW7doPv+E6sxBQD/+ZTdAKc4biGr/owK
XQh3bxG/H/3faXieoAt4DEhLR8hzxpViBe3yfibH6oemnBzR/whvW3zoaqNRg2s1+oMDCYOsn2Dc
mxdhsKkfBUloZVpyXp3wQ8j8fXArhnrm4o3sCo7lrguMNxon9nUj7b/CRCKSlRYlFvpPNSykltNT
0lnlL7BdG3hwu82/D4uj1BsM6NTYASmpR3FpCIg0H8cXYT+SzgRjZMYpiMhCMm5YAuGUG7GDjfPE
+gtW4SqZzi9kDMKyfVGOW7p79uBfLNR//yvmnf2PKbg9dQOw8YF1OoHJ7cd+PEo0yj/ZaxPXXUUs
SDtMtmsN1YXPYDTd5Yxntk9+f1k7/BfqjpWWy5mnGhhVKjqEKV7iISuIhpGOi/KOdbF+G8LiQcqG
uiixoySQX1t39ojZ9WGcrgWbjHrjgq15tVP9n5ytoUyXqrpQ+Gr83XvR4KI83SZN50d9S6Q98Jw4
XEUu22mNY/WL7fAYbJukXEswwjOfp7ThjW68OBknPY64HvaNt+UQI1zskTonzvOoSuzA+xO8thZk
FTWYDrEKSJzvyAIUNk3ESTHy8s3YGx3Z627zD8qRRdkiaR/BK0PiVNtskB1SrEXunx263BawYatB
I0DZdqpwlbDvzZUKNgxlrj8IPt+ADf4yXzdppVbbwlgLmNzYeRYQ/qdV8/Jf9qm889GAloS11HF5
x8wLaWCZOcs4VJswHiUwjBAMlYpGPrSw39p54BYlqycCdjik2nFhHVQFBvZgrdiXYwOp91eKyxRD
64hk2IySMf60+VsYy/R2BTRgRt96pZTdIQgPpLLf352O/x24EN7hIO3tKbPHCCYo7X8U+AaKn63F
kOukp2s1TfZ0+tShQBY+W+BkBCV82E7I6GifjHBDaXVfJX3/1xepUUvG+lfHRAJP6fKJtxMC//Y/
D6c3ebsg2kyWCD592j2dcdko3fEvndc2e0nr1SlO0CnFbj/4n+oM0/3aZcQl3NnjJ6RROJmCfKTR
uCFpH6po7rrUFPQHW6D2+HyEnQcrb1x1vCNnYRTgR3xs38Lg2Hq8KyFYvP/IRZzw/8sBjgGScYW0
j5KDHI1cTVdPYklyHvoiLoEdeo5XwtcnYJNg09cehlY4GHiwBhJz1CoAKQzLJwxQQXCZCG6IaGzJ
ecv+wVfTZdOlYTlktpbofbmJs6yU5gmeMyCMM4B2DY3k6YaqLU8k5u57y28uZe3/hsiPbidOdHaz
9+z8tqrWdRJ8yXB+zhmjxytzUcAQ2OSIqtoMcgeTR7vsxMwNekoKr5xMS9XgiQ9WIw9W+9qFzVq+
y/BHbNuy54l/y7MNobvEZaO7OLtOHbDOfEFcGWHlnfhn4ji1uNPr46HnDC0nDxlbV13Xx477liQm
O2tAtjzIoYiwZ67ZhrR5s3PDO4u+UTnAGI79JQfxur68WqNrjyYvgvfeNgOcDXfTg7yxhUo3iXGw
XlKO8WBZkaAdcrpIh/nSM1YBY0X3bOGpx58PjpqmR4USEiFnYc81XAudSqyRcRLCh2XnEK7GEK85
4LqoxkhHm/YgQ68i3LrZzIyRFSb0GV3LC9gr0FXh4H8myeaem2wUoFKVLMIVVLeKsFeD+rOlIeyX
NfZrwRy3MN1gK2XyJAFrRiK7TDkg7VcH19Tm0DGaL0LgOS93mabM0E/HySnPUHK4IPLnIrhdqRcM
v0chj4XEj0yhFo551MKC4/frN6i22qOfeHel7w3FqUexXfXOfEo/P6U+HjAe1lJ7dVyJ2LmovUUt
cg9tzJddMViKaF95yC1RKAieWHq/gH4qL4Z1l+nYM0NXjsumkLZIE9uqDZ1TdrBCL9uEPLrslQ/T
oxh1tBbHJtelvUaek0Yyi2/M6Nvjrvq6CUjxkLT+jFYrB7vaUqhN2GutsmvnE2Q/6G7vMdmxzyJd
DMBxTbyMnlbhvR1DpUtdnd6oZTMjdoUAF8c0JhBHxIWAYKeO1Kwm6qW6qvGszGJTcFhXyKkH4Z64
hb8rIFxoTns8U8m+rxvlb5W7BYopy0PfvXhZrvlJA91j20lK9kPom6SQE11Wg7e3NZPubzSzRZnq
pSx/nG8oWzRfdV/BW6iKJ9dec76BVPk0CLvxwdtFwCERgq0mEtk4AuJPiYKwU5w5bWYV4X13wIN4
7464tgI6CIEGuN3k0OT8PaHpiCWe/kPQmxlKdcyaqycRUAuMZNPtca+8hUVo0KeBhJajnxfpTNkl
y8TEmB7rujnxhtUD65ZPJFpqBuY0mV74awFw2JBRiqrxsujZraoWYQNpSKCFfLoaOZzZG4yv4k2F
uOn+ER5newAaJyeyug+ynfR3kLdh0lMAlnpG/GgRz2dvVfS3Yn3M/vAgh4MHX7lVfFUZEqKv/JiL
oZhtopWlc00HQugR83L5f26B0fQpTq4VAJ9bN/Z32f3daLL3V0XlkQReIOl46FtXcQferQzIEwrX
jxCvjQnjSxs5z4mR+YXW+giXgiTmaH0s1f8Yb2xpcXDzkm72e1VgzDLwhkYyMOtB/2MJKKGLLosI
cuSvnt281zeutt4BvAb4ZkIhUZY/7zeaFJyIB3L9ZvH+xskblgjS5damu9OmwXKbDihOJhucnT8n
7C38SORZoIQ1eFyyR/Wg/L02xwLgXPjl223e/uHJcHlbdWPbCDTzX/Vnq1r08ZncG1BKzWVP329l
P0sYV5cqgTuikle4eM6eS+TntS4UX2g+/LbtIRaEvxQGhIGtk6wb8aGVGMyi8fKhi+Vk6MaIPj9Q
tlildO2J8d/cixhUjKXSgsBf5jKUL1a3fGAW+rNyi9Yv4n2pDPNuEZTCms7xgCvDokwaTTRPNpcZ
0dZ/FJG6qmeIo/zlG2RJBQ2mMXO18GuOci1UdjuRnyEPtkTi9LAf3RekTUC1d2v7gAPmOfw8usDX
RUF7GyGRI2gG40LgJ8GCZ9pjopyryr6xPw8ShFNHEX+18l0iqcIxgJNE5LKx1KKC9sbeXv+rmjX/
a3PlQFL59gsMSvT3xBM9wXMimlBAl6jdCmaMU2IogXQN06E6AqsS5ivncuGREWrX5fRr+fYtibAK
o9QioodhWR0ythH/Wh/YF+CeAQZEdXvxhO0owJT86AomR0JNbA1rbQ+udP0kv/CGnKFP8115PveO
VAnbT5AR9mgPbiupSq34p6IEP9oKzLHMG4okAKz1uO7/MOSHnVxr7rbPH/Nn6TzDopgiiW1WaCAo
3K9yQK0HFcBVOCEV/YeQFv0NCW0kfQnp9tNWYRjWRJJJXGxHs1bjAJiKpx0Xek+RPTRhjU6OZDNI
XPsBLjWrOPGGvmOn+pNHMUwfLPJlCc+/Oht1cJHiln1T61es+ZbPgtmTxVOmdbDcphpkUoFB3ZAY
JaAc6OqlzOqa+wMVVyQWGIqS6bzanBfQH4+uiuZSmYTm7+av61LxuCWDQKVUgtv6BlHzfORNmNnj
fLnmg1D2r0muUiB4Q4CERGm1a0fE4Mf5//eHgsypeVpaCx05iL86Pm4YMFQl9Dt869LRyUa97sie
G+hh9lazsuQhPEhM5YUpDYfq6lqUcde6k+NQDIZIs0urHlrbXWIvubB8J67GnGi3mvuyYWlcqkSu
SjBFnZRdn5HUZ2PnUkGD9IPzm/rRiYRVXjDeWNnifVE+fTA7n2Rc9873N6F9t7a0k32Vk+kJYHs4
MkCzatTYzhUpu2F1fveE6Yseo+hkDfp0TcO1fQ2bYoUD+Y1w8aUyz/IAfE1btBjqcCFLFPMCdrZF
liyX+dyR380ZlCfLSJMpOk30nM9NuA7+nBT+d4U6jCBCaqES2ZRdJY5A8g8d8iN4E7jh+js5XB9R
Xp0Xq120iTIxgDoAWf1zRddyAjh1TF7zqLdxT8C2khmxW2hn1yHB40jXmptivSTuxa6+V9VWSlKR
rHtqBXSV/o9U41PLxTjsmdc63Fcypccc9NZb/2mkI/rqbh8K/BwZXZ/Ex8nMxa5ycawbDwrHY/Fm
o5NpaYUZY6FMusMDde0rr00ZUMLq4u0PdeK5EZQXNfZcTytp/PfEt8E9o8V/deh+D0kDVOra3Y+D
gu3UtRFc4+bvPDUAdPeU12zxtIBldiXGrxTBRWtbPQ0nPtcgvtIIo8bAKX1+WlbetxyWZwIA78hN
spH9oGmgOMB6bhiulYYrXzCXUX8U3rk+AnfVmFJQxXSj2ARzrBehx+MwT59zIjV/xsCqrkfyAmfK
851c76oMYxvR9oovvXoT/mXZUkunqB9BGGx8nZ0mxCURjJGa2Qjxhj9gv0/BokWOQ9el6WNCpC93
S1AMyAvlhASmWxIa6oqWrdKYDeJvUT6R1spIO2DlvoPQU8FBZAJ9jIzVClxcDtp6LkWc8A5JCxqM
d/iOEdHMYaDYIUi0/BVN71NG7Q5nY7RZPGfasAkMEuWLx2Cu7Cz0SPBBr++gma0+TWkn+kO++3JQ
Y8UIIsNijkH1VTB/0DsI8o15+Pypv/2OKvahcXB+JjeTCxkXeZI+MzdZI0SQVfbcuoqMxfAiHbOF
Q7Y6P6c0ERCc+gXMPBWeArHgcjwk++lNmwPe022/NQPBAIiv3OtQPIzngdLhMcORtm3TuiUEUK4w
3g3smhPu35p4WQcQRcgYTq06r9gY4rLao2Rbtw5sfTFHDC+eJnbzY2xCuef8L4wrRiSO2NoHSKW6
anQg+grui1x+ZBF1eq2196ufj94Okczq885ea8F06YwAmizB1qFAhaU9QHx/bF6uN86O3L1S+fFQ
mqaMoaE/srpNDjW2Sl58M99H+S3Yy4Ggv/kWzComZOClrwd98ouwTSdStld8zdJXKlvcCcXCtouS
kuMNCcjHKeN5+TOV66HuX1guDhAmSrC2r7jNkZ6GhDTXZl2YmTWkoGSXDPl3WUpHlf3ZzKB2xZrO
HbkSyj3NG7nioS5eZvCC3hzbCzvQQzWvzeL/dxvkg/4L+mvZN+PQaE32fzY+CF5GzdqHKq1gAeXX
Cu2D7Sg8iV/hs1jwiDlOclOpIYugU0loPm/8mXXIciT3OjMf0r3bNAS+ZWWEaR1CFb/pGm9fKIF3
ykDZ658Cc8MU5CoGHeCYskUy7F5carOf1ojD1BqIJQBtWeJC1XOC2cy8/nL+5m6aLuFIKvlDVynB
05az+gMJCY5OlTgqeH2HbBBPnk4cakuQoKZ44iWEpymQg4oJcCp4H/uNMZdtIiKJ6Mbk6upVowcq
T78QZEYDKEDjwsSJ8PASbSjbBIx8Zk7Xjks8sBZy3rNeMUJJBnGOg45/p31XdO2TeVKWqL35yfio
ueLRFMlyiS3OEPjCMCqS7VptLt3lYclDoElwefLIbEaYG4YtMjPVTaxT/O3K5WDI2A96TwPow1JK
A6NV77OOdztZll1A4Y/ezoFxtR7/3bWWdxNCRBtNgfRxU01G88oQk5sifgwknyNmpdZf3cRmCdN8
R18LFHlMuTdd6G9slB0IPd8slVJuLXO+/ucEOzXvp/hxlg7MHNScNYUQyRZH+YFoyZkmylHfsMOA
QZbCN83uJR+ZbiQ9L5Mtjdq9mEb0ODoXqA0/b9GTk/XKlFUxZqwWiUC5dXdNUMZJCd6JTi+94/yV
hNpUAyeaJInQB0HX7NlKpiejrHNYs6/xihUJ2sfIIDij41jGHkbujlM2HQk9iH3jeOIAVciiTLXh
Ql8sYNFGwh8pQJDYAg1SwXDtBX0sRZHT7kVw7LPPL1DWBIq9nz0tUG/dDQcVkl0GNcFW+N83nA+w
kTW5x98AZeCn1y2xXoBSJowZQxlMeSq7pC1BFFA8O0O5wXHM3+65oaibJ3YVPzoBjJjxeS2tPX4e
yJrkqrVKsimCSE8DNIaS/er/TyClNhEK7r2vIEzlPX/zv04rVbRVd7uTLWcLmEOC9zOhSB+tX0CH
/zmVmOrlGqkJr497H21R02Pe5iZultmDfP60n2/KCXYXYyQGN9Jb6RA4MSYPdqhHiE2EAxk11IDB
LOC5kIt9OU7ms2HIvXFlENw6kCgepFh7wp7C94xGUD62J48xf77Ekk/XV7wWrZY1Veklj4kc2HET
HQDUlESoQHvZs2LCUMXUo0lEmB+cugQgXhwzw2aCjnoq4CHatTtQ3WWu27RxmyB3pf3Q0Ewuu/Ex
6VWpLbPucUkPaZUiFZvETOvjpXux+jvUw1HywyAayBgd/ud33woIP51fwDrohF+1fdB1Vvy24Kcv
Od71MPApxklMooVr4nlpL1RdSomfHDTLIVz4zYHKTaVt+4jIC7RfXle24Cg6ap+BcyvqRb13/pTK
ZA4UqYUlHRabaGBClTEIk4zz4yG3ZqtxTxMzqjbEg0Nk4hqAspvrg8UMCtkClmkDwB9E0ScBNKwc
Y7iHarHAnzBAZ845AQrbMxLYhp7AdBCh6vPM4QPdw76x/1bW3S5scStezW7J5J/Pw2CRiJt1zJsL
sRbob1yG5DJ3m/xjLnrn5VZlKwy0+N6kIQGGSdgh0VgiOE5IxcgqpKbAX3rYDj7IIL+M/8eUQKZ5
g3Zytcur+IIHefYYh/RNdt56y3SVj70zCTOGadvg8y7oFaAOtS8Klw2+E1Gt5qTa8tGRa1/ldE86
YSOL7BRGVEZfFCzNk8lno8TKOSR2s/9ef4WFxQiKZdNcx7AMk2UUHvSQ9HlywQyKfD5ZyUQKWiUk
uW+i3a6Hj6WVOXzuYh52KALtQBgfQ0TI8TCiW5u1WBb4ALI+MJzMCpUn0i1j6FdmWiTnclt5Zw+c
uiOgqaBMoHyoUTR1O3J7/tE12mmc8glCDmyC0euzVJUFvJ91eamty0XtnPDT9HwBjU+JO4AIpwzR
/R7lB92DIybW1OnQQDj1ocK5OXsRN015ALWcLgXuR5LbimDwzv6S8l4XPKDZWa9eM8Jv3fTnAMaQ
Je3U+OygXsg6jMd2ijox0StEzqX2uGw8LzIOT/8uyV8vzOH4CGhDdRkOBep96O3ou9Mg8dmjbOSl
JXuO0mv52Q7PlNq7qA54kWNUGAZ0rqNGArWMjtU9cdqVFzHlvAdwNi3YkfwfeRyJzOrjDy9stOHA
AIjbKKA1ieLvQB0QrKGitJDph14GEHH3RvfwDtTbEV2MhukVN72/QF3Jwefn2iAeoSSI/kXLKnoi
pDjuUHWz/9LP2uCurxFZRObct3MnHe6SzOwKmHOHYUb0llqsaPLTL4HteXIzbudknF+Jey59duD0
Pm9UHeHSJty1cssa+k+OaurBpw9bJ1lfxucfbbH2QHVXQk/0aVWXT9QAY+9D6l5dK0vM1LijKhQc
0Aj0bVY6z0uhO1Jvz2htql5O6bkFZ9lAZI3BkOngNf2VAaQpoKQb3SJWNMs4M8HfXeYrO8zDrYa7
JyfNpck1Wx91/gEwkygSdKUMUOZHMNYLqKrnkSfM42oMfl5ByG7h/3ymDns8apSwUd7NVA7Rj/55
mXR0YlF5MOoDT8jt/3e2GQSOklbZX47l/xPycyRSE/8Gk72hmkQleip5KpsF743uW2kqFGowdw8B
B2n/9wJS0G1u6bXPlylz7usN9KR/lQ7GgIej1Lq/ohlY2bCYxwOQKs0KPUQWzWnctkMl8tjkrQDj
f8yoQwfL9UrjUs5zaAv7fP8XV0FjuDQptXuPr8MnkZAunYn780JEy7PiVHRPAUL3+KTpbkpyBdWS
LvTVvJRXtL335Psp2+1XN0J0GqFaF4q4z8vC8QeONEn0Gxgboc4HDnvMyYAvYcdPY1UpwZ1SqMQx
IibRm7LOqU4QCV5u6iRc45mG8MXCIqIRg19rXvJGrYXKThxv77NnNlKf1TX1IpWzFpVCEiTQZms6
ky6YJ3ddXAnFxWRyrkwt23VvdFF1k1AkgPy3sGX1HLkGpni0UZE9U1AUGeIWH4OUa2R9IgapEPcj
YvD+qqIUpuXTfZ+ESaS5JEUFZWTERabVRfPAVtR6rncpKgvhee6qWGqD5ggNTKdElQitI7X6BalN
oqtTj67/EJL/30oItA4Oqw6upZrre5WN84xrVDWhcc1hUa7Hr3bk2Q1Cg8Nk2AWpOcx5t4/paS/d
y/do9sSS8R7l+A399MPIIQtZcBaYhWi5PBgwrGCNDmtybdVKV1EbpRuvf5ugdcmMD9kuU00m/Z0e
9xnr0lHw8yfyyYUiwo4yErgn6GCqZACaLgz6hLCOoekJ7yXoCJh54MXlSr/Iw4JKuU+qNV15RghV
6eP4FXK9m2XaclZCdr2xrKveO6VK7dzVFR+e4U2FNc6TSC7/xzA+lJJKweeIatqk2+MkhOlxkfSO
yFV40vog9RkXzwEI2h6p3H++YxhuRkw2lJ5rtHRsRM87A51ZJAqbS0Oj3EDPSOy4Fsckf8wj3qQT
VL+TCia5prAnHIqOl9b1BN6ipTsr35lmFEsLS8xyTXehJWSRVmf5570hcZYwOtAj1kf+VM6eu4lM
cZYa+dOx3xscHQhUHGWxICpcCZTedeCZkFOaUMT45zZN2b7+BdF2FOvxqPstd81qxUWUAOe2Od09
ya3zpXOJSD2bh8M2263+Is5zcOYPbzbfvY7QrF7F11m/O0NMFALCMDj1j8jXTQf7wadnAO7utO9E
UOA7N/Ff6BlAkS7mES+hMn5Ew/J60S9zwIGzv1oETbzcFIRpRP2lt0hhjtb1YTYDAuw94jVwv21i
l3Bz5OhO3JbYJsCMZx8cJzum1AJ7nxuGpEoYYmbyVMneMsQLfuRqi7RvWHdMFHIgUSFzHh72gqMq
ZYWPDR8wW3S/r69HVwk2vKTTr1/fsCmYjH6WnP56otuSJN+Ocz3nOEirO1JC7bBSwESV0ssPDmml
6B9w8yxPNKHe6OONunbb9zeoNBzivaS6f/SR7NtHaQdNQF9CWkTVS6eYnypK93iuW+0maGG5Cwh9
/r+MkgNTtdmSDII6OrZO7apTrjbMq/SXZNDIKOgA4YR6S0UxXUzhst/mYnZagBZ9vpdtzGs7sbjS
iPZaFD3NjoUnLjaATWsmUnPAvtsLTLBdmLYpffYyeW93Cu64zzRMGLkxmSAboEcIRIlEaKagiRPA
DhoVypvSlkeCHAjRv2Y3WRmx8FEGC+GsVCAmhiIh6KYeAHycko9tN/C0S0WBy0Or0gOv1iOY4ive
vde//FX2t3reMf7wlGTYby+KZhtostikZXBwscDD0d3KlLdRBp9NZOr2rrTU/RATrv92xQZymnet
cpWMAhydPPfa+M9by8HmEwmAAvUJk9RdZecXbYvWdER+dCAGlTE++25PwLRpVORTKvpqwgsK18c9
DRve6V0Ewg8H8kij6qJTORUOOPfNWYE0OpJJL/LzSbDvrdTGAsRnV6MVDF4aXXsE+nKWY+97OENs
GU1Y1oJ0s4n7dktVVwlcVrIVCe16h8/tS7qceK9+/UTlDC75D37YhIPYn/2mTAFpc1E5/9EFm+WO
5tBLYePAbKT7/Vvw4osCxazc/kGp/4Xd9j/nK5KRsoL/6b1YIvW7hwzAntVmM3Qn8IAt61FHUaY6
c3/mGdsqA0hQxTfjSdHAPPqUzWXITTPPTt63j4pz/klS/GyxizD5ipjbRn0qpeOGWwwsHHVS3bhp
zZLPIhGu2K/fHsL8FUbGx/ByIFR37L5JfuisEgLxmuLwY3+Nxc7Tu93X/GK2KGFB2x6oKVKnWx1G
6/+Yw/SadUjCsOI6sySpnZNBc6wZtxOLdyYD1tprH0mP+TceEvp3VjFlRYtVHfx9ZfgPgdJ6O2+8
EzXwu5iRB6XJpTwQLUCb68p6O8/Fttc3V3UgaRynW0uhlLFrVBK3HsopvUaSGMSWo4PRz14hKrCy
LaMl8GoF7CeQQN8w3Hu9J4PKe+nS9w6CucquXi20SmQDoSQwUGnPOc3bGqlncdc/yPHkTJMPuNQZ
I7aFSMJt3jSZGuwVL7ecZXttN5B6R+rirUFFkF2HV2O98DR4LMmTpT88b9VD1e1951VKGtRzBt1A
f1ENxpveyZg00ugPUyb/O2nQRKEGCUTkTDtg5mMi6qNAD3ODgpx5GMC24ux7jC0DXwAZD5zZmMlk
tJQJy5d0J/Ox6fUC3X8mL+3gQAw7EAovS5x9vS6lGV+rdsjgB7IkS41eZ80WOdnI5vK174Btx3CH
b8y15Cf2nGBad51WbWVsmM+kOZclxVGlXqx46x90dTc79du7D8HiX4EgPBRXpMHvDwBCsvHeCPzc
Mt1Tt3T7Gh+xnRFUikZdGmndo8UngcY6gif6rgj8U1Ijs0jcEeOKfR/YHuy+N3pmoe5+UdCOz358
RBK25j197TtsbWZuLrHNfVw55lggAiG2eY11Dxn4piAYpi0irdJCm7ZFDGe/t4lKxB10SjHGPzYl
Id6MG3x5MQtKL0N0X0Nakw9fialCS52U21n+wWVfmFA8Pr7XhLinA5Jy3wH7KfjKxTr9zc462KlM
cm+JbCA+MzEAbop3FsETczhkGP8cU4o5trXGBMTVQc3LamWEvqVIis4iRRgXU47aKaY9UElDMNAp
K5ILeWGu0cvv9L5dnCOfafEy10sDZpLKvItEAn89GVMcDjmupmy2BRxFD8JWp8epE97wa7kDXMAZ
F4ixM8DBen12gok5etmPni3eqXBqYzQxEFJnKAEDShwUBd9uXbPZd/zPlp1F01O6H5Khbzdtx4Fd
nhDMBoZ8mrKrUn3XY/zD8EbbOKKMEVcTADGlQJN0TVcO9b9DNGD/dLuckbIZRCniHgettb9PCaOV
59vbAJoUsqAR3/fsmkZt3wfLuhBFJmKncvSHNINIsk1xns087qXauqJhg6RURHQ1smBIzFvYPwpi
qijhgXxJ6UoOssyxTIHSeFptcQn/SgmmR70UzlPuOsGrPElGmKxqbyL6GiVp0K8J+wtvG22MiXud
9q4JLKOLA5EmHHjFo4yezDoAQXige95TOIYrKamn/6i9X8CEeWAPuzQ/lIYKMoOl0c1oj5yaPQ3p
tBoelw0woG8p3Seq2Q5k3l3WjrnIs2Dn+LipZoP4BXlpwi1PiW+ZvTtaQXWAJgA6V07PrS8bH166
96GToWlIq1u+AFvnRTMNHtqHoCBxI3I56raaX2+aeGDCRjtX7hmz7dYKCHKbBiw+x2dBb95nLU2u
3dR78cCuf8NeQs+RzYYbWupwBZfxXlLYECru9WLJZjEQBTjCG1ZXza506NG200piGA6z0HKcGNHN
YFYwPQg28vW1DbIs1b2xrGoXnxf/TWGIdCz4yaM/fIHEmV5i9/pvAM3wZHOmPZnDfsuVP9HahI7w
fJu5mpLK8m+R2LZYxrfib0CDm2d2WkqUZv/1m3nTmm2dhYmQiNWxilOkYEuspRKKRBhhnaaURAFP
9dzBu+p0fVZwluA9qUU2TF6m9Kq48Qprmvt5TRwMA9SyKDZhTp/ENOVFEAMpB6gb2b6JMrjfiTAl
5xc9mUAcl+sqF9/c6zos1nEcs3KsK/sMviMHNSAMPiPGnkdraWH347/nK6050A5xORva9j6xUvf8
suyeVeXodM5PCTSQPIsewBao3iqiK96drhmDGNX59H0nm82iGAVS66al0p9iJzDbmsDOZb7hBLZV
kqWDnxQ/VlxbWOTHfnXIhQp8xf4WqVY+Ech3rraza0JCBvw6De4oUl2+OMhXrZVGLLXDWUP7v9PR
dnn66RXDpZ5f6H0Qj4M41zylYssjSWqLZZtWhxHTYgc5w/uKIlY2iTqRoAYN1YcgDFmAOUv/UWzg
mpbA6f2rWtYVkffxuy/kxcFHgJELr/qsDeFjhlHyTHdPWQKYZBxwWqNfzMS+Hs1sMFzESuxZQ6Vu
JPnZKGPpyeX8DHQQBnHugVOAni+34a451Uf0QQGKJtYgnFC/I9cP0GT6+FbUJBCDYXgAUWf+FqXB
SkkhF/+T5TuOlS9z0P4lXVjxVI2TRRSAQzDlXWJ8GC90Kka5QyIFXRQ5dRd9A7g0X594pYRYNgqF
xvoRBUaXQ7rFIcvSbkQ6NHVewmDjDqgT5564/4JtOoAcp4grwkwzpqC7QidsaEFsuLh+AE5y6jnW
LDJyqdO8IXiiXsJuBNAjo4nxRA+aT81CVt9S+BkSpEXmZ758hiRBfoHlvEdzbjW+wCZbc62AsiAo
d+gBgwsR+YkRSq7qlH7gveC49HdkyFfAp0Pg+CWl3i6iKS9zrXWu8IAaiIJdQZv9rNluaq594e/E
1KOjbEFEGAq0GQWbg086VF8Mg08+oYeL3TlaKZa03Z3ewF2XstlZKDbQtzonn8bIiOe3JBiit00v
rVoMm0W7ro0wftQY1wmq4QDNaIfokpxzf0gHhZWhrh04n9EgKDZsBwaLkjamCFfEjcJxzFhLgxYI
abKACiMXQe0/oDXcCoNhVvuy2oqBUi0sia2TCMgwfKWVaD0vTLQv/Q9AwOtV4k2PgC1GxApaDvz5
yAFaT6F4ULlvLOS/+M4MB5IUUEl8J7VpJFMv2TzlQN4l9n1yFgXJ4YBYv4AmWeA+3Lb+qPfZkSzJ
tiXy6SbIOrmAkMVB7VR6AU1XhbzfwZHE9dctlidcn81MnNYXrpRs22nkbEszT+hZ1ujjMtldvhh/
sY8IA5/xuQpOWuhY2v+EpYqMO7dqN8mhSz3P8CDRKFcfZcL8J8RtnirPvSy1dyxgazTGmR1Wbyd6
aOotm9Y5AVUyrZO5y2iWYrCuYfbPkQoKXdGXNrJDNCj+ag8gXH/NSRfsweoeei72erlQntJSirRa
HqbddSQHvKBQyNfUqb6MybSnWfWZ0sdf/GXY1dss82jpSLYNIADBw6KYXB2d64/0OsFisior67iH
KbepUnMMuIQ4yss2o7DYHW4TKvwftM7kpfZ+2MsLenAPmUJhKWlMfpd4KG+9v/c38hDWpMI+uN+0
3QPGrHoCzAvrM3l7oSiimw5uhDMQeD3TAyHfFKyy9kb9UHXSMuMwd8ovNigT/4hKu/91LpfgQvGs
zerC7t/Nr7GlVzE2n/9s8rxfSKxXoV0X7xFYKUA5zIAx981zd6M4/mwhKUJomJU2iplEXj+XBhff
UN2BHlJ8vDHtXG9TapQRvkR2Vkg4NPGnYvA7iBxEwZiFU7Oum/3ZOWbNQ+b0alfc+/XPDnBs45fm
T3AcNDKEnXn8TK9p1NzXH3EYjDs3pTsxm3VNRH6TxgA9gEf+3aVVyrIaVKqUnRQ9eEhbr3psTQ77
1svLb0o9kxTSOdOo51HO+h5m/dxHrrALhz3ed5zrxOH9xH7vdrTC+WlFCojG6u9e26reRksm0A/t
U3n5EetHvexLnMz4nSPwXuFd45EQSwrkMdkr20V9f3PPosRdGBWrku3hA3EMSu87el9zKEKcz908
VSZsQiZWpRE8snDsBHTkS6GYuHekd4CaBalQU4NaYXJuaqzgZftVJ3Z2JvjWel2AnZtfejCLxzb8
PFl8hernuzhVug4r6nzC+uJKmylDVDqSWVAw1cinLJRbVL9nBTbViU0qU3pR5RlDzpDaJKIkAAx/
8ZoVAiiVFAILTelJ6s6KDY2d4GS8a8HXYgdPahKD+cId6pyDuCD4zjwEc8HcL0EKRdzG1YgJ55xF
Tu4VqoEHLqTGjagzruer4eQhMqa5TxaoDGBANHwLLSIN5jrr6Rj+Z5Zr8SVfcOZJrLkb4zqkOTgK
pXM+adoHrJVp8wNLwSFH0s3B7RJpMthC8x9DU4WFpt356mvZDSBWedcx0+E6H1h1bWj4NhQF4LLM
Rjfmd4xve3RFHwxTd6XFREIPgAVQ/byqvve7+7kixf6LB1vxkFXD5d5RsUWcflZdxS7QoLoiNq2J
nVPrepFaB1WVTp42+l4PTaMI+qRuFouU+0M/IUvvChlk58uUo1LO9EkPhJ7Z3wEidy4qV2SaHIU5
q1fbR7VSzOzMzRZoJ8bb2G/nnhxdPtEY5XDm3Odo0OMuMFqpXJ1WghSlzssATS4uJ7cbyXH5hWDv
YR52fG4Zr49e2wnUZojtGkCevjQyqtTqdrUlEhgU42uGaNqIvWkZkurr1DdC3aMnVtouYgSuzQEz
09njW3jF87E1MvYg1Z5RH5i5ZceEtkFmNfCg7pJau05OlVJes4J1MLtUBd7pcO/IlVEx6FDKGaQU
kj+FKg4aAO6PYXkgZH5mfi1S4llXqasHB+u9uQO9aiTbCQxWCRqIDQ4yRhq94CpbEpYep0Li2pvf
KpiAkQBWBTyaZbptNN2u1vSW550v0j2b/KUhWZvv8EreifhwaKxHMZusSVdNu3oKoeI6EQvAPfMU
LATHtjRGO3SFdLZ8AE7PjYoURfIxLO6Lst19lCrrVWWNHwP1IzLG98xsxjhCMznP/nuD1x6noTLI
tfr4BI//JPPOtUvKu8t4UqleCWgRUvtIhqlT90enVR+025obh8Oy7VaKbFkcGXJdRM92Ma8g2tv3
nO8h5WmkyZ7ukoSy6NCnVFnz2k8P1jcBuELek0J/k1XXeTmwLI+q0kjvA0uaBdU0pRDvxMdsj5mB
sdWdgj9hH06sMoWWR9d5AOgSR14Y57DlFA5tGzJ7KZsug+T22fvo50rCfTRIFewwRI1/rD+sXn/K
62vxZIPoPs/BY9FIMVrveue9+1gU/JsiJncrbTmBDb8LiScHDw4VEnubi2Hg6O/6sdWRhphmgHtd
V/V3Z5kht75Ofxv28kQ1wXn9mMObgHtLyOipdw57PC8SXQc5Ax3ct02G+yUNpuOY8ngBC3N12egC
oFzKnbCcKRZP2Zn/9r998QQlHdYiZZUP2DTku/4hV6j3z1xnswHtIvLAfBwMdTY3j4iMBAwBG49z
Dh57fRvPeTx2+8VevhVEc3eKKfX/UOl1zq+hefvx6DuMXXrtACUIZpqyy4VAFfS+ttrmghZTHOuu
jBQ1kA4aW7Ga8IG2j+nua2X3VJSWRVEgzObYTY4JoPRnT6mk1XWZPODnqKPf7AR6JmNnzItP830n
1vlG51NmaNS2gU1nOdbt1TmUQBbE97ZlpE461+bxY3hq1fLaEjMsZlMoodnihIR/etT48kICwtnd
c2oKsv2MYxhC+7dzqFgwDXl++8q+hvlCsBsOchuPvE24ZlomJsRCToylYHfoAQ/PseeB2+MlkZwO
sLI4gM5OTLpN0OeGid1eGJdPCoH74JzR3pjSfhksnz/BzwAiZdoJWv7fHuWgVaKPpmBc40QrrdTa
1s8U+3iKlxhi4Qb9yDyTRkecifSj0bIH/XnCNETM2s30wIvuYFL2ga/e8rb4AMqUMVNHPdPu+7D3
OXOFJjLjGYGDhPcooDbCo25xLC2pOG1IfcLO2jIg9qsXeZpJnMUKZoeJCgtQ+/Fdq83hIkCacf3u
smw29X2CD4pXw7Zuti+lVxeXIyPDrS7YNgzgK+ypC7078yrt7mue78OaW+1Viv6qeSB8NL6XCfAz
3HeisZ30zivnkEu/v8te4Vt6Th0yOxxPQqvijb9gkZmW2hcyX0wTp4o43I0Qdth3o/KrzaHvNLIy
E4Eb50PCZ/Wu4dFfrZXfFmoPJ4R2vPsysLtem7T5Pd+Nu9Y8fbvqQVWQ9O1x/41FVfHRSM4DtEwh
Kz42EJJugbUQdk5aS1n50oaCn8QahFFLz6Ldzh3ViCE6yP+AV7qxDzSpyJsK6EPosqBd41rI/vLG
RfV7/FNKWXEeLW6uW9wGb0I9pFR+VGEwTt3mDnyAJrezVNb71JZFvPDGKETPaQ2tUEHBPfx12/yn
uWabC3H7fLlG36Ug+bQiJdLa0wz1JrOhR3ezQ8ide/t2MwWFji/A97lNMG4BffmP6tMVgtEBZaxh
BlLV7W+Zs/QAh2v3E9cmN/RKk0vEXy5u2wwdwHwfixAW2QqOKRPr5MOiH4H7D+wQe82NxCueOVoo
suSo4lr8K3R9bffQUTEIrC1aiqetP8DZ6Q0k/FQq3pBLD5mWvHKkEnmCR7NqRXnGqGVHBb929QP6
xMY8GKHb9pdNR4WE59/EOP88QGRpXd1j/5d/wHTccZpD9z6z1KQ98AHPD6mmi+Uqo2iz0Giv9T+Y
/McPHB4OT/MFCapvv3hHoKCTW1EnhhSWA+OWJz/Z2tfxbfXPvUicSu6RW39UnzeYqL9ElJPSClw4
qThWYHZEni7IaN1oVLFZLcVSZ7WaoKlE94Ss3R2v2uKz2Z6FJsMir3/1lhsEulsuYQCJcQMe34iw
tkCEY94EPmrpJn8orbCJyXrxOwTfJDdUbcg8VDYnQGCyXHvWEAFtUXCFRL7zHe0+vjLFPRcM/wnM
P1sxr0udx1K1MK6bfYWcvlCYj8m3FNO/xveig0zmglJWkpgZVpVmY8pw2kKY/SBFkWxyTf1/sgpf
DL9WZDKWmCr2bdJqcQiFRwvkkxYvxiRc9qUCpPxUx9KqZtzGslNY4ivaZ3954oQzIY9160Ieelnm
nTGumKDI53jXXU31Hu3LHoANJXtxO8DxvYmYr+1ptIf2X1dcnYEAipxk8KDHvTc0NnQLuD9N/ZoY
Z0ts2EGRo+eUBt78vKii/OHexrmPJEbXnCfWcmdiWEb1fDRhmveXzXxvhtRmsKm5SQLm0M0rcjqs
lICAzb/ipBTKVUohxOpQhEt10zGeTOYHjtwOb/xy5sDYovdbyhZYVM4EH5lsgG05e97rDaP6a1l/
Jr4jNYt30b/OeCazlzNshbe+We58wrZmQXLia7BNE0HlcNUKlAQrjUPW0Shd2+y3UCyX2r9r4JgI
MH4DwQIQRgRrMkIuyMSkWW++paAjK7TxtLCLYYSGmi114NYEkPf97nAjT9DPi+bNxZLpjaoKoVUO
RXncG8C6nNQB9LBvprVQJR3n20fyk/azKHpoUhghKld8FYDHIY4xoL2PWsxnbiK+REpOKUouoe7o
0HV30JrzYj4V1Z/ioqyVUagPyF0MePrUIq+iZ44/PUu0nIUKwy3O6G23iStEoK/QSV/r0P57uJ0x
DSUPrWO2+hr9rxf+M5/iAWgPMshNA79xyGgJN1JDOydjmC6PmcnSLN0zulOdwy3zgc7CAFQBMAJr
C8ipaotvt005ugVgyjMkMAKmY8vLc8mlyQvC2L+VJrRBmd7uWno25LHP/oq2tFbqlphQ2kBoagv3
61f7qTRCBk4BdSOca+WCJA2Ion1eo82KJp3IkJ4eH4629i/TYvgUJLCCX+EhieMF0dKLCAcDlT6T
CebqfrcVCLsSudqkSO7dwIrcEORyNPe1BWg5UdTPHQBxFgzfZTFveU0hB8zNcvNyVNmu/RnIg/mU
zNwfRm7pai5Es+FDAZfSmX9W4cwMg49r7fnCPQmKLoYoc99jGd4X60iNBR6vUBc3YAxGLy7P69aL
+yo7UT9TAQrN/mdfoGNh5QAIvl86rjSAwyeU9yVH1tbMME8kMScTGeKfFfgJ60anhlMPTYiq7MkA
tohHOGnfdP0MjCPwcg9GSYPEEgAhqexj/chM1D22m73uCbqNikpSu5mAxhh+dkVfAdwj8TZ59DCm
A1LUOhNr70/7kbFjDjgrL+M+aqcgFRkgzo+IuKyaNMElVFlROblDuO4/naiiFyH+l4fUFLBZXVz1
6Ly6muUQahSYplPxA5sPn0AJpT/AjcaJa7nUpstF3TVh8ZCtoOJl6QdkTDMq4F7TIBWBBghQj8S9
s1vgjnM6swP41wlN5TQ2f1fHJMj6fSpcRSYmc8+BNIQ2Oyo6U+O+uJeijSO34uF4OZd7mqptREIm
qoOhyjIcSNny3s9Ckf352jtpwg2vGEBLAQg6OYg+h7akkf7txxkRkbEfvpZik1vm8IbEpxylnv1A
CGm6v0Ju2l8WUno9IDj3co2rwJZ38vQvdMacCKiXBzIjv0amvEqmJyyw6nP9mM0lh0jY8AUYvP6e
i3n/jWECd+alYvQgz2T97mk2T269szGsDkZUfK2RlIuNh3R3GPdMfzn2wW+hKXeoHZ0dVDPIN/yk
SzMZkXroyTNdaRsWwWVbtDSbvx5VS7xbVPWp9Yy7ooWkT9hamViHsTtey/4ruHvFGvDy8Bd0rPag
MPxQZ3yaVY72JrWyYvYJYUpSG1MI21OEvTkZsJY60XEiKuX9m0xHbLJFcjNv9XT329UV+l2/ZahH
2ki5fKXxZilK8J84qsd2WygtqVrZscoP7TlgHxDVMY67roS6hdvLr9QBu7fQ9d4WAY1l6wHXTYez
zUVwHK+RR4UaRXEkwUaF/0OkBUWMB1gyv6KJo4UuYBcbJ+nXgw2OFIECxTcyXWMdNBYKYIGJp1Hs
YH97GfDQQ8KPD1WUjKrFtjDDH4VmNTFeCNOkVrzmvDO+rC3q4Dh7gjfyWE3UY2/bbk6bzkuavEM6
utM27aB+/eWJV1EH3EWI5UKL1S5HccbUl5wZvhlnL8UfGfs0/PTybEAq19y/so2UzGZGbyZIxmzt
BikJEOlzkaJgzJgE3s1OkfUoHhdBt2Wb0mWi9IDD1noMI+DzujdKZXozx1lqtCnn4boxCmk82KRD
0aJui3kb+lTnn20N91L8bZzCouS0+LYTahWNbyGyXdI7nflsAMd2FY5OwZwoS6ycC1v+dz/YuMTJ
lUJyFhmA0kzVBlKdHlsjr+YJC7ObEoVDatVO3xr7jXGkRhG3G2/MZ7CcYdlmJtm6YNiH8DtOB94F
MaaqKD6iqhlD3IvFzuEaMWvvxu9zRt1mlIWavwG+B+UzZ+YqOCro8oXnG36yj07MoHmVayEeWXG6
+drEr6GSLdj021AkVIFBqyubuixGsdkmHTDVJjDMxGTa5oEypmVlPZiGFVADrgHJKhvSjr99+Vw+
w9SLCkGPVhcZjBgXMKKgyRSnfO7yE47sZKjluAec/F/FV573RlAbmPQ/s+qgvrpdLwSP4VXJalFb
oTf9FBNiweQcIIJimy69qcuRVre0sS8IOEpQlpY6pF5WraFgecjVarFiZcWHogClqFmR+ZNUw8Ba
LkzZ5XFm82RKfD2Gp7pSFWcgF4Jh2q36xuR4w1+zWOwcO73tvXUx6ajUA3GTID+Z3gDYdMeeha30
Tl8htPolz32O8+i4P7DlYRpbi49LOX/LdJvs49sevAIw5PPMfwyznIP14emeaMHPTQkmtEqM1J7l
cnHkEPaaKKWwgLYIVYIFokG4y5m5X3loq0Se0Fzzx2dKUuNR+HjXR7x+IH3HpE7dTilv6f2hcm7B
pXgYd7epwp3x/SoNmvIvQaNLTDRE1N6Da8TN35pmJ/lrlflCydudUdSxeodbKF0GckPgOWub7I+7
Pzu5EeWYZb5WOBTxRwhHVS4SPN9k13GzgqeWG84A4bJEeTw3d1Jzj466Au/QUtq1vsB1GE/dL6+c
aBA8lm5dVK++ux0bKrixZ8XOb8lWVBpBXKE1wrfxNzV/hZRdO8XPOpkHlpmPWWy89ZLtM75zPkBO
kW3HNWgm+rBtz/adlq8cqhiJfQ8N+ww1LSZK3rtprdOdCZ8em3bpYRnT+w/LwET0xBty6zHPyL0k
Yjh0FxaoTWF96vBUXYisSlLr55NCPlW0Q6owA87jzRvlWTkQY4eDG9eGSktyAsKkC/NdJStLDH+u
QDdrWHnF0+P9XGG5Nz7aT8IhHqt1R7C3b7ZkVrTX5OxXi8rKXUm4o2YFGTdh6TP7UMFweSbyhTz0
JHQzcpAdoThGYzmRlKPokJsxARMiRiivcdUAv2yeACE1rl0LkRwyimP/J55B9gCOIvw6/yO0pq2X
oovfWYvWfxBcExsk5oz2XNuVB96smpR3fc1GRlaL6YcvTlmy0qjg+6FFu9U3vSZ1E9KQKoYSKigB
2gibhz01KW52CmSX1diZhAT13tmTpz21aIMM7cxERgD59rqq4rzeYXTSEyBDqhrHatlhLNDDatLu
qZTTabjG+AwJgMM/mrqioHHmk+xSX+MVfTWJ+247BR1GVYrx2Cr0vVtAA8tnuxhLApjLt3hUmIPq
ZDbjo+3yNih8A9Cc96V7zmJY54DEm8+buBcgvOJXaORyBeElsjciM4+358+nAXnQELkR20mE4d9F
LbVRlEJbLS+uMvYusL2BSlIdKu52BJVutBQ9GMH8F1AnqEEfd14gE5uJkbWHCKBKpttgp3tol1rD
kfgR/M07ChQ+z0T9bgKxGNG3Bsnw4iblwVHK2O9lyFaueX7mWtrrejE6+Q9ML4Do5OKglGW/jGlj
rkicm6sNI5BNVXoiRWXDPAzQ4I4odE7mGuw28Qj9u1NzfKJV/N4oIXaCK29FqnznsI0I1OqSFYpF
ssUJURYnkZAaICW6ZdlUv01dJ4UZcHd+SbDa8GT6OnEYxo4Ld1PgXnxThomE94H31hxs1/3tlmeR
RlmGTq4jtG6fvufnrql+OqQ43zgR62Xy3cA6/dJrk2a1f3kOd+sFAc/MDGMGnUHlvUNiXDaOAfOu
vHlMCvZwV0kw841AE2PQmoiLYDLPQ/OBX+6/ICY1ReTfYaEaO+5uuBDuMEGvfbDcZSb18EvJvNmJ
++juSpywQVc9+52NVEKNhsKVUaDSo1aAjsEGfEstzIX72ky/OGoZ5siA+9BAjQUbpCOwnbsWEsQl
RMtKmE27KXIAx6UvZGfW01asUsBdOuNiSnmkZbAylYYeqXJY56W8fCPEQT4mq8oFa+T512SWp24C
vpOwymF42jdK3VkVmiFdcUX327Lp8+eDQQoOD/jRs3yvezQJRkD7GJ+RAUuOEVAjQXOKiapDKYcH
ae/0z+gN8VtKKXkwznBHlQ3iCuYIgGJnB1/OHt8z9pbcoHNTm5APbURGIF3c6Gz73mO7L+4otQUA
MalP/dMpBq2PS/P0WdhsivnF9DkZPw4+fqh+yQ40picGfyc1Ou03+n/1vMhHH9gLoXaHol3EQMJq
Mzap0L31BVMV8FuItCph5fJEIKiUSK2Y5mUtbHMjbvj8Avtiz9d5C5nJPpvJh7UjaKbxQYjlsqg0
GuvBZqZqh28kj8OUw31ub/b1FJFkGarP5UDCT5lIB9RUdTgMC1i+GZwliiUySjp669yd48k9PBem
3sz8Lsu4KR+N+bMcvKoyPMx/qXxDu7sZCB23j8rhlJt/JHlhb/oXBFjpiZgZhh3wlvYd+swYkQ/I
ihrwrKf8+tuWo1gxfhJ3OPBbL4kr1QZDcwn57kwShxzUPV1ICxZEzhrj5YCqLOCdJlJiJIRmzgn5
6byyEmSK5OTZnnb6d1G7RQdatkkgKVKsF5DyZwqf5CSeubjks5D6db3L0cZyfe8QO8c3UnqkgPLb
K9zA2Tn94itQEzb06w5kcM/yeY0+bpmyURuyq2Gk45R7ut/9mYmyKhKZUFikxqwOt6hjMCydqQKy
w+dVRcc4puFqYoKGxrF1KGsn9jsqKiZDb8hDUclVL8pOAv0Nir5sUK85QbtCmhnXaXVpIOd7Eo9L
i76g938DHOHAyp6NmDtAHROa2fjbhSx2dGt4gpvwQIFOTyqx8Fb1VxtOQI33sXbqwed/TSOxYf2V
ZWd3d4gqsDStcFFZdVrCfI7FS0gUJmB/0RO+o9F6u6tyERhIj4+b/AYD41uxIq2VeYx5HAQoqtIS
w6TWMYKbOL1EM2xrxf9iYhJOQry7B9JPImn7qxJgqThOsFeXS8ho6obhCkkMNU7gvrKsGZKOCOal
UxOYXc3eIKvZNOUoqdGReqYqkSTT7yiV3C/rS46qmZdOdVHPeMkLcRmrLrunTCyAFw7DLHPJDT+B
UqfZvzCjQsOQMMhH8Mee5qh5vwmDgOyTKrzpIot1t/2NSKQcvTEqZh0sYcnt3Js5c0SwnbjDLd86
g7jVAkCUzoDcLOgtZkuj7xN+A1Jn3tWEITQJ8le/O+5ZSMDk8/Y/+3Avvd573BAQ30KL81TMxH2e
BrzegqrlBFOJyW8PrMC/uskVj+0yVe5dt7qpb2JaxPoUsJ87mw4tV1ddIZwncPTTCcoIhWBTRL68
4NZsV9FHgDQl4LbP/dOqKhm7yHVUhUACQPl5LxNSbyuFY8KL89/BN9jq5d0xxOXWqFZfDhbbIRzC
oKeC5M3G03m0Z/jUG2YidKUP1bgM1YuaUb4ct1kPFLZFD9kPfglRJa8Co3pqB/aYKxaOrLQLPkV6
beXmbzlweEi1JP9WgmqH8/HZTO4M1mpBSqqi6g9Y031adxrmzPwAX37NqQRh1SVZWldA50Iny11B
0Xc+0bDfN56YA6iZGXHpLhzGY9n6CPo5zMfwJQhMU87G7tPSdIUqpDI8+j5SsvbB/XyaOKWiCgaX
H12XJw3/JGDp28VANkwoaxBX4GTQFuzdzjDsE/f0ZZWjcjEQ0zmeWNW0qOzpBR/MybmnY+hjVGsC
RfZup9c3t1Wx0/Sp11ZwGSwdcG+yfjUX18/LAPCA7vf9LbfkSl7wPxiCJNFEJ5tYaJMe4enDVl0D
AKMIDHid7d7bkq0nIyalVfsAs5GctdHmn+QHhsH8+UL/Td4gBhUGmq2R7SKevIqKJQPK92U6mo9r
LYTshraiB1ZQxIxjwJWdt++c0ADgw8IPTVpmkrViYpSchV+N/kFI/vtprVAgjREVUFXnmdtKPdel
XvF4y6dP2v7tSwoseveEiTY+zXRhNQGVZbn9cI8HY69r4eVXlfPX+yYx7uNiJvspt2Dy6DpLvjiX
6AGA12xb4sQmjdDMJRMUHg/zvBgaq64ZfdjwuCu6BJaqd8DDMQqaom2hKhERCtr3KoidluaMofwP
2RgmuY3FTVNyqRmCAc7zTw9LZA9vmONgmj9kAEljc88lxpGVX3BSehVZLr/D0DhyBKOzQpRi7Sun
GukAnhdQQBoyRsrzYoYnNCXnO6WKS8y/WK8RjAKgatwaeEagNv7iElp5cq7m7ja/+nGlDa+nJAPA
Zo3TIWgU8D8NvZl68FTdsJO/Te1+2jbyNpU5Lxoj1dlSQ3HWqOw6z+JJfIrCiQU/r0gsycAitZk4
KUcNEm2dC1jMcXxxVBQxRZbxr6CAa9e4m840e2gcz+UNdgMJx9ZpcbHatXZE05BxcLFt2D9mOw35
tS6Ar2sHT1uAUVKAPD/r2GpiS22zu773AXUeTL2nuHAxngJ/YRJCwYgno/KyG/9IO5Iv4fzsdUWb
/BE1N75JmFmXy5m0xl0FuPxORlVQWQ4DKNvqKFQf96RAtH6/QGGF32oFVQmdhg5bCKrffx1R5nLn
KgM5EnOse7k+DCWy42KwIvLq7TLC2Enm02Tj1CW7AM9u54TYcU/2PwMU8Vrky79UWLfhT3l7yOT1
3Zabgs2X/WXvSxwGNUkkvVS9mVC88F6z8QvFyhb3dFWPYrDBK3L1++uzCfLL8B1mpf8lmIL4YK43
NfHq+D1BPjecKlcQ13EReFzv4qAZzzptzn9m81R09iijyMnZMKhIkwZPv4g+J4p00c0dMDJ3lvAm
susLraIYIIRHGjG+1cG+06NZ9AGf9mVoogf9lil9RZguK135L2YNLL7m9L8DCXHE/vkpnATp4iXO
Z0DBMFXSlzAzkGVsUo9HPO78HA00ki6jiZ0dpPHjffvbWR/EgWfv8ymiatYuewQWNGGLPPmSJWcn
L63qwvwtPbx6cNVIbE5Ck4c2diN2HyXo0qwzUyqY7nD6tID7W9aYsqVsqmjB+OgOY3APIrigXqD2
5KKtIfBWV9HFALTv1OflCJXE5p+eZOblDMDVlcshMuns9XCWq9XiMjJVLvQFVY2cYeEW5CoNPiwI
gZiwd6BjX55jFfQ6PfTjNwI+rw31NV4XuX5dSeNn1Lg5OIjqjXA6rJYBxX9+YIjProYw0p81U+BC
ZbEK2DqVn0LOvhgjv3k0i2LVr4SAhnfnp3QWb9dqucjFSj2p229tVHQiabkTFFCjEnuU8PjFnR9O
4VkIvkbSYbN0CAn9h+Xz8yBswWwcFqJIA+fB1bdj2H2DmwmNSomK3xYOy8e/O0/0Hw/UrBEN25Q9
ww1J6RK3wKvEr//rYa1yU7ri6w37OUuDw9fsD28ZOBFShc1IkJVHGPKGSaPrjB3KYZsTxJUDHSSt
gefPdJPvAyGBlxB0COAZPJzTKAtg6fTR7fSxg1SWz/PHjF4LH1Amwnq4vJ/cHkZDnfFO0Pwpp90A
3TBQtIFMgXDoEYMXZjNsyvcAPNajvUUu2BrVLJ1uSQL8P5DYw6H8FMZMUyUSl2oViyjT/ZamuIlo
5J5HIoHHjwNQD3Uhr+gINdQ7BQB6zqw6pZ9zW0eMuHokWndbeCrJqkrUGLlG0f6D+kByh0wUjMzF
d/hunKCN2PuSGV/gIxjYrWrIWFZBcJlt2U/lJi6y2hLv/y1//6L0aFAhSZepC0jI5aqFY9fT21Mm
xJH4Pi9FtU9i8ZbEy/G7z6bU/DHwO7UFtUhPtVUifkUTvgBqUkJclhwS5tifBNzmzn161KEGGTEl
pVKQXKM6lwx0tBDhGdXiWiacaulIxH3xfk74wbQtodYgjgZtZZBRrsyQ5YSuC2/7hwn8M0+yIXes
71gNNdsqhCRUNu/C+emb7yTJxlEG0Jd8tTn5wCQzLdv/r1bVuT71XlLFpy/4XeRD3Y3S+qz2/ZLD
rbdc8sXnjtm3n9XzjpST4M4HxblMPoZ4Q/NzJYSWcW6QpFTCD7JHRb3wzUyGGQWAiTa9Jo1ZpDuJ
xhGc0SZALCM3cfhEZFFGVAeQOPjquQjTzmCKQuO0T8kFNf1qypn9yVmxq4qoC6KeUu3W4JFFcZqB
IKSEUEi1QiFDVpKxTogGNQBDv2teoCE4CBdELf0zyG92I53JmQk9qH7nhLihnxCUQ7cVhvlYAVfN
WbeCIeduCcM6RF9+9ZV2rU8NJfpXoDRm2pSGlkbBVMtYG+4t/KLR+xRVGCY3YM3KFzkUJ0Xhj7E0
/qMfkP1UTinY3kguIgik/53hAJ5R3DDooykNFHAtVc8E5x5G1BYG4sM4vhkEpvSEhXDo+nB19pFg
P4Q2Mn+E5VkA3nWhJ0BMBWTICuipBM2mmp3YXn4ZbydvtDEFHNfVmqF3ZFQoKDMrYISo+je0qaN0
mkMtNgqtRp6ZDHJfGPTjyZ+LqvHVzWYEI6Iejf5RZAxSrWCCKwximdVruIv9+xakr1ARrpJgH1kz
Yl0mEAes+eTwcuae5aBt1CL8zPksF8T3rB2wFUr2EjNONWXqSXEbAPYB07irUcN/lHub55XPnzOM
Ex1JppzjSf9C2TxeraJKOuzMNDsWhCoRhWVBnAgFn0fNqYHIdebv0xTtPQl11BgN1uonscSRlQ8U
nOZOlDAg002N259eh56JQdifpK0fp2kb+8k7vwnl82Gc77YvsSpQl5+S5GxjIK7YKa0e597iY6lw
S6Aidv4rGXne3gBuDaslsHlmds6O8beflZQxf/t6YQJ7v42QUTrlSjXOUq7Y5A6a1D9rgtd13Tt9
Kr5qhD73D65iH7qjxLMeYaEvvfhfeeFm7Db9L9HJlbV1aLfODvNlp+DzpF1PfiaprtyNFoRvYMF6
rZ4FBUf+K2aGDIZBXwCSZ3wylmFk7AOPfPOWECCOupXrwSKO5uhDE/zs1Gixu7MfYPxiG/uJsYIx
/cwEloMwao0axjI1lufc9/hmxSa+Cx/MAk1B2FDZuAuhLwAjyhibkRc3+ytFjVlQ54m0myoRhHnF
a2g3klujWixBoMRKkTFkbMPdqSlj+qwnkFzTGrMqD8MM6SPNMnunGKSNiz9VCbK2utVsLB5Ugk/o
kBDC1iVTOzCB5KvsdBq3yb3DzAUXFj/GSjWbURWVZtjM4pCn8ZrlUN5Rw8Gf0bhoTWE3WF6MYod3
UTUXD5H5rTsLMDuCQPca3j7zxTXlirzoeJnTva+JIFV/drX5KWc21O0kMyv1CqMbvuDLGeirwvFY
yhrlNS5lWYrzpmw1ENdAkTdVqw3PlBJ8iroMcXMRBIDT7gF6pBe1WNZhq35sxOgYtg5T1SG1Fi1u
c+FiCkM8+8hZEtztITd/xGa9zeSGT2rOy9WjHIRUFUD0oAnP4581FggYQ/bUdZYZjLvn266GJ6M4
CL1IbdNzvDb60yNmr0BWmEJU4tZFg0A/wKy8VzVoWEwcupI1Gl9WGsoNvMzFZbkQ8u4/zVVLjnKo
ponFp9H/PlPzrQbOUgO/ZjCGHlrQuIp6qVJvY8iWY91hOX8tqVftmTCVRnF4zYasBuJoVraKtqa5
rpyK8cHtsbKdYPbICvwmt1pojxOzTUfw33lqC64eEtzldqxhGnFJpRkyVoTTtZPk8DFLQIJ0ajIj
IXqrXAynpS2B10ROWhQUJZ20DKz6cUSbpXJFx3BchQsCPB8eMHvi2GggXYt1fXHENQtapt1vIluN
7ziUluM0nsnolMz3nVgTAPaocVRqsAoLjzzs9MqGKGFEUaDx5ns2mqdDNQnNNGwAyW7Glxxeu8m5
7SF/JSsvpOCN484PEbufudCxHEF5djWjKQuutOch1NLl/KO1bJU0HEAjE+uRtMJ0G/7jIBaF/nft
ZRq/FTgU5hGmjxQ2MuRaOEENzCOqAk/rFsbqaqj+KQa+yPjbUqg6gnB13LZyWZ+zJCTai4muUImP
2txR6cxhvHaj5tMiVW+cEt40aLjoMknrnKv+rl2lOfAJhIzLMtikoqCumRUbzn4kN4po/9XT3l6N
LBvHJ3zlVvG52bgowSc2UohVu7eQRsQgCwpoKYx16qznCq7dWNGi8qwXyjyomB57Y2vhC1Zy95Ls
YgfTewYRtkeabmlolKBZwwfCQ9MoHjfPvdc8JBPNA3mLzXa3WJsEnTLzEfLAb4u5d4OOHVM0X3ty
Y6qv00cln4zUEJsm8X/gYRH9HL7ySQC6XFyMDeAz5tt2utEkrKgG8/F4qvHCRUO6Ima6dLJmCcPR
UxqD6yYEQ1AJlNuzKSn15Txt5JrutON0CQ5CfiknUPLU/h2YJNEQXNaYlQhrmQjCXu3qNTG5dZS+
uqIm2N+rAfaVoxb066nPFQWsjuACvO9raZrUNyqppVij0LFAoRVq+fWJSSTbOzlm4kX0CNJ+6DBU
BB2mkNaC4qZnOE2a4kQF7jAthnYLyqz1Qgnvqm1O0i1UEwFRBG1lugEAKQGUluXiuDFTPSSDRiU6
6vG5XZ7Sy3XcZ46k2Pt4vzEdgMA04CpXiaOihC9DhObLnMcC4471Zd/stX7SF1QcA6eQFbj/fPSN
XG4sqb/ZZS6UI7UHuAbrIFV4ZDtyvRGo6CtRjEAOd+ZC4DL+ZpQQF9gxto+U4xKZHLw23hirFnSK
SG3fDM7JxDdJmuRtCFzGM/oSWKuz0G93zEHBEsnFOxnQQRoDsKUgHpMhkzbcRH41Nd+pbpZdknBB
FNluzuBr4qw/4bFRbqScELvL/av9+uPGV4okIQp46z/W+RK7m8i7z7a5UGuPl7Tz8VHJ3X0bX9yy
e9NkSOf5IrEtJYnO3KwX1dMyiPsqDnlU2Ce8qkz1E1/mJavFEfNKkqNFNbFEyVLCFQpbvgg50wk0
+ypH0eOAwrGcUoE5qfxXartNJiUjJdVduYPjtaw7rlO2VI7oVd3ZRBlex0mDy514u90grXQFex5l
B4XGjMmVAsbqq/8MAsDwPjgUYqxkdBpuiP5wo6SxY/j/Cn9TZLO7nPoT1jJIBsrH13BoPS1LqSPB
oztQ0XpQaNep8psXJcxqjDXZQOU1NhKGIE0IOhJr40WfysSZze+uHf9gr7oeVJ2IW55rDg/o6TqD
D0WmT+n64rZdqFZ2pAG5U5jR1RN/QTYI3o1bu1Hx0UhMREnAmWLZaD0LWb6zrwFCJ/D6x1c/QIQR
q/F7hM+2pSqLYRctf6GFWyZsON5ntwu7g66ThOSNr3d6EiIJksilMtypQTEbWJjG/kD35121Dr6o
s1PMFLSYuuo/e12ZqJzCyjSuqTBgE88+l6XRYrB2gKLa+UH2VCPYUtWhNsZGYdfttn9ZRROYCCyp
i+ufyUwaxqtytHZl2Idm4L+1THkypIkmHLxF9LfjdyHwYhipP8qKA+//U2QY7F2t+whzJSWgAGKp
aRNnTsmpVJDOn9nqtHXOwXjUJGszDzzJfpZA0kMdJEAtlP0kL0/rXvSO839krmcqbOvZUdqZZdon
mbPCri9qUFEDkyFDee+SEpHj9bFHMa3QzeElBUJK4H6wmTlv3BoCWPE6ARmNhxeS30XiNOPuOl8R
blflgkJXbZdt5QyxDcBtLRbjjKRhJv6jB7YydtlACvWOQHuFUCr87ypRzRTRe07GhF6QKaf9QlbN
3+BCC4hb9zc3kO9lx/JhqgEkob+KHYjUwesSZhxYdzaAbr2SiQIjB6it454dlxoGShwmxwwEJCpi
dWiG92CBFkM7o9YdvM1pj070OTZXMvKKRsX77TP6sCesoKebYNzvCEMlMx+Xch9eKEiXG/ulhDLy
/7yZu74+LDEBBDhoIdo2ARXHcyh7F+GXMhBgvjVZ+n1YePDIU5i3X87G//ivcWpU5WdggOuKK22n
7BhXVY8J0qKZxbJmePhmiePsWje0D4ebDM4daU/3

`protect end_protected

