------------------------------------------------------------------------
----
---- This file has been generated the 2021/11/22 - 15:46:18.
---- This file can be used with modelsim tools.
---- This file is not synthesizable and does not target any FPGAs.
---- DRM HDK VERSION 7.0.0.0.
---- DRM VERSION 7.0.0.
----
------------------------------------------------------------------------

`protect begin_protected
`protect version=1
`protect encrypt_agent="Synplify encryptP1735.pl"
`protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`protect encoding=(enctype="base64", line_length=76, bytes=128)
`protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`protect key_block
aLKGtZxiX/VvUy208eCy/Pt4frYR9JKaXargrPm8+BMkw8KeiYFKM6iYRotbplYKHbQjOaAVsSNj
Zf5KxZXU1udfNBHaEmjbWuPe37/P3ygfaZKcNS4rjwCpZ1XWHVheKQJ5w2EGLq2euj/IXl2YJ+uj
vNn2WircMn/I5eSRfpo=

`protect encoding=(enctype="base64", line_length=76, bytes=869984)
`protect data_method="aes128-cbc"
`protect data_block
RBQ43laTZQI9h9jdKDQblsCHQSTDP72+EMf28wi9LB+1F5wvX0yV8aKo4meAeatOrrhIfzsOy8iv
RNV/QAbhZyoK0mwGJiX/WITZCgZWtvLpcT44k+kbfe2r8EEzn0We5Ndm3StsOqyynGeIsdGXemI0
/TXHfXX9O8cV/41zqAUjXxyX/6rCc3Ko3pD7cZ6wdJHE+5cp+aJXwyKLILgGVq9WwIN9+Wp7sgxu
Pzk3JTmU75UYpgvThFeAnRC7XiKwuRKMbI2lL59OtfzyYCSgzD6kFo9qZnnPp7GMad+WYNWklEXy
esgVM7m5duPMgv9juaCcg0yGBLPvxdIouT5Qe36VnXBsojfDObaVEEQr0pqZ/mP6UDqrF4C83bbf
YmKBAkxEOsJFY4XtCQ8fB4s7JGjxZ+6MgVWqz5jrV1FZPALiIqi1MNqnmTkwbitTRE3JZYO44TEi
Ge8TiwMDVkkU91aVt7gDl1Vs4ar7st00785WKwIiBFadLkaos9hr0QhnDqZayE7cg5bp+mT8LCyf
goGBmAl47malqzrb2DP1VsI0vWezLQcRt3rBxBtOD4GFBO+jWMJNlYZX5azYcY/BnOwyKti9HgqX
ELZf3Q+wnamxkUP8hAhkRHHa6SefA1555PWiRJ/VykkBnYk+I0DwfBgzN86yg77iMYLblT0BmmWb
sw5+3jLxmtjOsbbnFamYR6kLU6JZtOvYH6S964KzfGIpQS4aduvzvdok8yAE+nJ16XJXwHBQLDKp
WXdo21A38IKAIydJNXHiLa0rhKSnwLtRLnwX3xxtH+GVoSvRq8erlGBL3avhuCaxi2UnV+8bQvjn
0wwP+nDfJ2jG4TTISCbdrglKdIjG25gd/Nz7SAh/LV3HzWFAK4snADEbZMFvbw3EhirAuxaURPmV
o29ETU+392jbeauqIAv4iarI+k5+gXeyWBKPV/gryhzuh/RQF2YaXgHAf5UPfQSUmQ9dfJ1qW+qc
+EDXzZMMBPBv6GPWCJbtrNIcpie9PiFaAhAxi1P2tNNAlUaFcIRLfmWP3Z+ycie60HkFS/mQpAQe
FPL4MLfCERl8TFJ+/Jb8qY8XmCo3kDed3Kf+fPOGyDk5Lu/1u6qwxHhKvIOxP6WbLcEbYbJEoXmA
mz0rsfkyhsClfPCyShFovQ3oFuQ4ilPaiN91RGFVLw/gWc2/xwSUWbOoBi2JTQIiIvYbB6j1+KBC
HEf3QwWmJRZpe/wgwzKbjeKQLaMGv1iq1zeq7VNv33Amn9FLXAAg5ELcONUxEJYc1DbWBlZrgtmB
p5fx6jc256EnxBuEpHz/jFuK4yn9GYLqGNNUolYerddBFn5lg6v0CGirzkTfTKSFbBg8JpeNkkOT
WDSW8Jg49vRfNmVbt/hzdD89Nyi9ys4ZA2/TUI2gqvt5l/HH05gp1lhk+4JhY2DqKHaVX8J3sJ2h
YJ4nj9IfVWsy9vVaX3BuNUfyxUlDZ3Ecvnrm5fpyufNCnrTbWmqz+AujWd8nSSwB8Y6PQK34Az37
lomQPj+h8JNYzPYoJrMkJ34vrxsXGWSIp9s9jr2M/Dy53/e2lHKW7EDqGbM+m2/kxILo3kbJ4nQi
M9tNtHWXCDQ+6hmFOAuvxaX1DSmXXiihxVMdmpFYxZzvf+hI9rcp/ft8KvW5vhVn08fm58npOMLa
6cNQTZUq1ZsO2wCmbaCW1x/+dnrvX5fDW1avzyh660wpyqCkvXWpI4KTVYk1m5+D/wlRFRx/+Pfv
NDQMIjvOw/dlFcqBkTpIaSPQrL2JPOt8a7zZyEKibhBh3ro0Uj9DEaFW6+wOQZZsz50pb2M+uZv0
QlG6xVd/i5179dkwm92kT2tatVLt/FFv7adglpDFPsyawX/ACu5gBzDY78gbO1ge5eXxRFHkSZf0
NJhx8uDqth6nK4wotFyYf+uBJ320iLDuYAIblydWZkT//43UeGet8WHLF5b50cl3NyLuEZuFaK6L
HBkTI9A8u4teqHJn24YOXaYJNNTL7030V72alJF+H2KevEyl+Ly0QALGa+W344Mk8LKAhiDuprgi
Cx4zUFK3wqJBoz4to0s8GbOasPJ+msMZaHf+J0oCbT9IgGRLOj6fylE9nhMbdJ91v4l0WtyYEOfG
MBHjYqX05ngvFJ+pbEeCM8CCDSdVsvKTw/IjNhNs9P7Gk4J13aizniB7p3XQLNPNT2/0/WDtonVq
IcIkzgRW1RixQlhrG+T9yYMme9T0THOwbrgyfiNGxjkgRke5hlKqlglNmi8GMF6bsvUj/fm9XLVx
zE1c0hDAgRkkdIbaByhqq+tc4lREhQlqdrNxLiYnBCnCY29EnkzeRd7hn8b8fQLLEb1SaGVB6jst
A5UGS31vpv3LVd1Gbed206PVyw92rRCcs5FeKPfm0XRSXRDhr7OMhuJD+g/HhiDsoX6WVgKXaZgL
oNlS/hqxTpZ7jgbcjsfLnspc5s9uxWzfe/W+LaaQFs0Xe1Oyuw6p5spVT1itVzNPibmRvsBGmVxI
G+Va9knAmQAGl02WJzjErhufHVTPAMa087cuaBhPPQU3rre9RggkyZ5VFDf2gmtXdilldMmlwLEw
RIpFwFriPHTGdL/8lj9pz4o0/FTkYmCSg/RK7QQK3Je6k/j8M1L2ghpNlyXehQxHbao/MUE1cod1
xB/vj4NYSwopPKiPq9n2BnPOM+TG97IHAlq9ueJHfeGrPqRVqG95S+h6/p6lUyRUmrN+Y+B+js1N
gnwUc4XuZoHn3NNvTu8KhPiisPnj1wGQtG9N/hVtE/4d7nn56o7jflALZr+88tSDn1DACL0/I25/
IK/3a3qaIAl1z4XDTkiHKCjrpcoxy0Jzf2vWYG+G5bue3tlv0FxK5/KW4TKlHFKkH7GXY2PQhJhz
78jsA5XOyq4TTxoILz27nZlaznVnZccGZ0Q08UNjU6wWM7WrhKWT5nNIg6csfjW8xwEXHx4er5vS
PDssB+aHMYBrQNZHgAMfXpR2/eQehxk8CdyU86/BFoup14JzVFYT3ucJiA6YgVkXgg+2TaDabgKy
a5vhhrCvy58jNY7ISsTj9go+hZ1pX9zyIpS/mSnbnV75C34Pw0iUzNhqCc3ghFEj88u2Jvc+1L++
1tQwpW3p0Co7XfhlW6sGg/b+DxpV8K3ZVAbB5UriBEZMtGYcqAjPV8l3STwwqWk9eZNkbai2jUI2
M7sFgcObkA2sl2oGYuQ7Ze0jOHYGmMmgtPmJHyG7kEkpWtKc9RwQvRsSWOHwKdcPE/v9SlpLR9Un
oc/y/gJq8Aymk8jQqYxyKrI62u1qixYz0+SZUlm+KN7LxSCvBuB1Smmz4Ac+QKeceg5GiLDsSJEy
382skFHvdlFsMAeOa+o+rIxJ72FraX4uyE9I72EMEFhfIPyATJxvqSUELHDnDGSxz8zOqw6St5mk
+/EnywHI+KSOjrk3PS2qG4zDxxzTjV8IZPZi2jHPCFfZOfdJJyUx0jFqqKlVOHVvJK8a+opOuk9k
hEQXk8b73/zzGC8CtD8tRCu+hoqOiBuu3fevkux9XOosjjTXHZiyz17edzuQ7mQqkAXEGwGMJhMm
myT7l7gkJ921OoSGFgTCqD0Ria06MWZ2VEH0WMeS/pjdFqm3wGMAMu53mhC6HAdPbvSewSpoCp4l
EZnc1mDipIcwhmj/Iz8BJ49dz2WT1u44c98rgK4bcDTQ3xP9d1lZXBGwDfsHsro9VXInwUdpI4DD
KIBNd1g8TxWX1xUNWKNjP956efOohHOOMhbuGCecGs3OJzcn3BI3KcEMaZ+vrrCyI228ksg7GdM3
v+U7QKQFmdQfavuvrPTddjeFzYHWil5R/gw+cYgwXJy20QTxR5zAv87WhNw4u/DKSpXyqXzCOBDd
aC+/RhI7JgyoYQn/6lhnv63NkL8tdQ9ki7UIB0NlAyIsRI8Iu1ELEWhMYI24q/ItU+ThJobufS4N
SmMXvpdernfGjRrrfQm7lNMNLTLcsyfAcBEVJja79nxP4QzOIysWHYcMLm/kXpTTPglyaaQ7B+GC
W0hIgbZos7IbUvOaUf4CQxjH+qWoje60ciwJ0N0Z3Qx3+4vjdkAirgjKXR9tBbiqUNM/Z8ZwKtqJ
aHdhWesfQ97+iE1K4vwwg1NppME5u0KBGsOFUVkwkScQo+LNPGy3dzn7nEZMlX4nO/gujZaoJm5s
S1D1/Y8ZrPRmEHgg21m06oK51264Q8qdsLCIMTR/kjHxYvKM5d5WJJQuGkAu9/gt+2IVNXj449dh
juz4DPJOr4FXV6WOjae6sI5IweqigsVonk9txvdIn/O8Zfow56gl3algf9WeTw3w+SROOdVHawed
9yi8VL98oGrZYhDLBE1e35MuAmlMMgE8h+AL0l2+/cM3KAOEmTPJlz1Y/H53N8q1Yta3f0XJ3nQy
ZZdCSmiPv2WFmw7bLXu7Omx/oDDi8lrhHwquGe6p8nXur8J9wqiHZjXa6gtegeALLygtN/4mh88Q
aH2xsLR2I10Zk/Skbk3FqHPM2qAllTunlWDdGcLorrZI2Wk8lWpp2OK++zZ2ZS+qmk5sh6L4n6Z1
tSAStDiAFUc0Cndgh3S45Vm6pe7/o95HIzB0hiMzgY5bgxyk9lIsx6r/sD3CvKrf1BaSM36a7r9r
kXWYvBqoF0WVLGA0ineo1lJG1CaIqGlytQimkIOx4tV8Pr5sCKBJtQJK92f5KLrRH6fM9k41omwa
ntInZLvQ6vui1O6hvbQUNl8Netmi+j+Y9KnJvs5KyhcImzeZZkprMYj+uDby2Pf1ZkXTMfJk1BgY
2VPF7YNvglisgdVZ9WKkKy3UMndUrxZjZS7bwmdDmsBokHyx1zrniqL4ohOIQbWPC0kZIZrrM28j
CVVaGsE2ZC2PJm/KEMFTQrDSeKBkio417ri2RWtTSUbnyuknD8WdjJG6MdfgQmr2KQJm/5CZuqZq
21VX1gUb4e5GGV+nWn+4zPgdzK7kRAoDCV8GRdsYBA8j2kaPmddlfOsBrB6s1nGEFo9n/MaE8TUT
PMJetKip/kPYsq4PbFN6YAfuRR8q4TcwDmFDRccsQRk9dkrQ9UOI3fcXSFacHyLX7PvWw030sNDW
pW5U34MAzH0e4ESGlZECKz9ue7rP9LX+fd9fyqryzFwwzlJQo8Gr0Ta03CkZSRIVrLCf+7tjvHsM
fjsvEaVp/PnCdNAu7Pa2ryzE4k27y4dMNgycJt/Ka4Cakeh5thbib2SvlyRiXOMqDtLDXYpqu0oQ
4tfcKxgdDob8tfNJm3se909Mh9cARBdvmcdGXM7wZbAtrnUhDwd7hi1AuIGhO10aVX0V1h2k0r5f
DvnqWbvwRJucxVjzk5nmRV4WxejgKLZvGd2xzqNMKPMV7fCAiW4PGZn1k8i39NRe9Y6lx6QEfuxr
vC3FYxwMAOcduSwNtY458alE+ouVfkbDCkM/Sy8wa6aGWUxIZR0gjX9+YV++cnEZRlFfMriRznmm
/HHNZlxiw87Hem09MaD+JuyKDxCtdG1Ha3PgRJFk3FacV+nWFvecZO48TLq0RMGDFwltVNhmoypx
rzzc9FqEnw+ZTUVCQ+mg2KzH+EFY/Jze6WtkrrvGnUKZvcwCHdim2vNhb51qJVmHJe4U4EuPlBBp
eTlJ/jcTSS6jP/GsAiRDJkUuSQqP2nTAjf5Ku3rN3dkpdSWk5pmXq0XJnJpQc1uh5fulA81y1+zm
ITzlRn+k2WT7uv2iY1psQtJx8Mn0e4CFMMg4FXi8inPa11tAgjMF5YHW64aASivdSfgpGB/a12Rh
b5YJNFX20hY4DiHyzHLIkvtmDbHqTjcAibGF9D8qOguLOYOzxeYfJQgGZES+YEUG20gFMaqj2LAb
9tbQXVnIMneL0MDP87ANpoWfaTWdUFD7xn0huXxlZf+WPntCPmx1lQxQo9clRDo3kdu+ZWDELLwA
WnSSlNV3jDSpdIfmkmRLahLChh0ei4q18rW44Pjb9DDxxs0mEBPqq+rDqujhn/Cbs3wE1KcYC+Ac
KaaNUuZON2YVURxp5tRKOCDr7b7Av6kgphmJuDt5QjhoK8/1ff6zLgAkuo+R4Nx6uwkvBMPuP6OO
6GIcK3mbOaPTjtfkVCrgjA1Bfm41fzL0nWST58zuSK8xDa/fbkFn7tr4biSnxrAhUi/AtnqIw/pt
KDWNR6xBV8Fjf9vhSp/g0E0Isto+bo4cwqTCEkQ3QaqE/7fMPuTU4ypAbbmY2UQmUrb8x6CAQnn8
ri6yj/SzZYshRPXqkZMenUK5JxaY73wKK6rdP/jOlCbedr//uHfvx8h2E/FnjrLpm2QDpPSBnMhn
zXQmtGLtFSzUhclPJibKDg29qJyGXWcsaH5HiM9o4dunr9onfhjoly4MA4S24oScLh6gaxbLAGjG
QZyyCQuBRh+4x3RLy3T+aNDOcwkh5QVH/8xVJJDeqMCsLLt2j5kj5Y+smRxoPjb2ywTgO1JKgoNk
VOAhoJCjDDSbU7Bl44ViCWKEdXQoOwLqEuvwD8nZUvcKk3TXNpfPJqKy32q1Mvau/CgwlK7glvHY
HzPNCGwLLQl7szH/lm5Z9Ol5UXRW/Tqw76viWVD2aYe94JvknLyhXRpGXpdZt8tUhCcksNtM9Vo2
ToPb0KhrojebVjIF8k/B+xYJg4M2PpuXXMSPyzx0F6jLEA7HU8Ku0V69mwvuQU3rQyPngx6+SBho
I6lhYbqaWNGumbUbvOKY+uleaEGwoe3MKlt3AR/NvxFMYjeNPqGiuZmg2nu3UXYI5aa3fasXx4ZM
LNEGxcQb+1R+pUDc6pweZgtjHFEKruxPhxS1e2B9U13kISyorz9Bzt589NabajBjaI/4cF+HjkPn
YpG04F3UiLAqmUPVSKm8d6u7ksVN0ClsvqNLfd12gvZXHJ7q2El+me1F9U2AqRiH2w4id1L/nNNJ
UMOLxV0a5GXX+hDnFCGEOPtX7KiqUqp5eCbmU2TKjZu3UX0EmNeHGhZ+1Ve4nloGDzUL874++8S4
y/uVxnTMxVjs6jJsjXuhYJa5r5QdtynqNnIcrtdBc6rNhriwF4KAL2Lt9h9Scoh4j5YpddsYBFxs
WnETNHgxExh5Z7ORKRFKjumZcy+ibJx6qlK21TPIAnu7c/iYfPkEC8xyKWYHyys3syLxtkFB28sP
PoSImV9i+PE9BTodOhtS56sgmGWuMjuhasmNNjE/f+Cx5oe2iOM+Dt6osxVYz6mntpoa0FD42zUJ
ifrUDgRSNHg5hSnmmXWhiZX7DNwJ6/g0sYYmwc0svXy+SJYbi3JECDgiWuoyIt1sxGCxIqUoHFrW
D7tJEwx3yNarbbo9ohx/9qhDV3aUI3Mebf3t82WdZFXjcHZNo8FcnKY87LchCSH9zcDEphPwjZXl
BrWhYKuNluAnL/H0r364JtGrptIYc0G1eFMuJI0gu+la3dMGNIsz968EErFs4vbyX2iKL35h8peU
U8/vbz8sAZq4efg3P90jJOpQ47MNMJXSxSZNoP/YBrzJGyk6Xm2Ydhd5ptU0BcDxlPU0CA1odtJK
mD/aMqWqODcvPcthyVOx9uNQnmpkMuGNai7IzBSeEqu/n+M0XKQV2NHDpK8tSKUxxWNVCcq1Jz/K
6naEMYuoXKTGiVgDvIMcfkbZKZg4MgJPsyRMVTJdSYL376NUjBq1mLc785iR5o1eiiYcqUd1NdBB
KWVzox4WNiKYajtlKVV+ijIA5d4cenGOwy5CLJ+MFZ5cIqTSPEk6hVsgN38H0S42hZ2VoSleGkRT
7iBVA8QxWhbB6IG/c1fmCnTeTeIJLaytgzZ30FJkYE4ThrWc+mGRIbwDd6s7W3nBFcFvspaJW2Bs
Tf9Tt5/r7IuaGWU5tKCR/DBpibpExU+JIsNAnwkwWn0TQE3pFu9Jz8zVya/p6zkIMbh6QpbrNgb+
fV6a/e0XxEyVqObEc1vv+lVH8jxFy6pn014K3PqjWYd85yXEblVTEXayUNg6PGnOgFbNI9CpzvJR
t7+t9HbDtwsOrc13IGZ9nwNm+Y3lV19anheXxTl389X0Ahk14b1YChQuXShMImw9E37+HXRQ5R82
gyBhgkeeiJHq//WWFSdYxDM8Xh6KQSX7yu/BhqW8RaE0z+8KG8ebDVhEcRpGIRuxtHeSa4ePCC9p
llUT2v/cYL6LZRmHMCu2hzNboc6cS/BBAARVJogpXBWNMpa5ChCgNyNOQsWJsXB7/a/SpKFRjLE2
aqplS5/19JQeSEpsCzkxACgHQ+b3UQlBaKzOce7Iu1Q9C1gr3OnQMA8QOFKTjGOaVoZIN5p2eVTu
ETwoFfk5JKeMq6Jt5nz/V8Sl2vlB+diknXERGunrNFUasIc7JLX5dJ3CF89nNKZW1GLkjjciwhao
l+sNf3go4rgW3opMpxbftGbu5Ds4YxMDU9y3cm5r0f8cc25zMKSMwnwrUYDNZrIm8tTOg/azIHiT
wN4YOJITsW2blJb4VrNYvdvpJTvH1rII320VALva8ZZmx8J084z0omC38xINk1LIcAYPWDM87rOY
q5FwQVQmR2yy1tndpGo8+mM4VzDW/rQ2kU/VphTKbRD7mPfwuToZjaoWmdtJ9s+Nv9FHjfFOi71+
LOP7An4XCEryiWcLUBcFjAk4KU9w5b6jVK3V+QQPErZZlRBPqH59fH8FGyvuqeh2aaTOyqKQsKN1
oqwKlPiLfd4iFx4Cj0MNDTmQcOXXGFvWCfzTAvgNWWOPwQ9uvr9NeI7ku3dHLz0Axn6AaO+d1iZM
Xt0Ugu0s3l17dnGFQp4fYqJlwdyYcUgpgKZfucji4nf8g0arHN65E2Itl/EftVuLcv1YF/Ylrle/
Cb/Ox3sygBeEIi7HxqO3veIg5W8WMLxM+xZDup0pyPZnEbHYiPSmTJF09GhdiXjVdfNFSZJVwI/W
T4y4gg52gb1KBNPV375K+NAsOUmHYH49Nh4IoAgVffEVB9zrXqYo7RFifigCbAAMUMqwWostCaYj
LW4K6g1hCkD6ghJNUFiSM76Pyl/H0xZobK8KYk9ahGlqmYQx7OK5/TBXQ+w8FBqMAsQ6+YTPfI/J
RClyKUfjOueB+3xBWV5EmF7tvH6imN+HPKGNVIdDV9TByHHfg5wH/XAVp9808SYjVkKxsUQv/xAp
9ez0rYAc7fvoAib638ymzLf+JA9l4fHB+6k8Wu8FplhhgOsFN0At0jumq6uMgZgfMRBD8pr/o1n6
dvBNTBY0/wFq+btC/iLk/ZDJoYLz2Fhaq0gaKjThZ/gwlc7ukWsIXzlkupfjKXx/0ZRpHHnEtAnT
xz8ve9+eIZIhiUtnFjw3HBRnMJHbKHeYjszIOek5XrcXPs4UaTuIOMDNyuCxBgNsYp0zktrJk1IX
Yace5lPyVo0fcIfXo2SDJez20iGBRwAEEZZviP8WCwqSgMUxNF3KsZviNDPw8YEkHhQSKO9UOCZB
+9aYKY06az8xbH8AqOonP4DKvzFLbC4ee7/e6ajaBnE8jJrkhX8z4MV1XEnaQbKqjGpawire9dJg
nrs+o0O9R/tTxIs8zN8C7ws4+3V5on2AIznEZ9VHQhCP7gTq92fOEU9njObOv/2UZXZY7x4glgLv
cgnTgpJCQku8GH6rWUDFIs/SfGJ4u8fnRO9AKtAy8BrCjHMrQiTWXFwlzfDwLRy9i2l/5HJlb9AH
91DkP2Bk4NYen/IhHJqlIQ4PG5PHxUt6fQmQQ1MJH7gumzC5EPjUW/WprzOo6/inVff1lIMm8WfB
CSAh5kD9+yj7AKi1rzzwGT2YPShREMu1d7AKLLfecOX+tlUlHbpLA5U5760/DhZAYEkacAS9rOnd
6Quq+nm3/f3N5TUDhWag7fqMVbBeCwoBE0UqUgYzhbcDsaNl2uQ8Z+w2j2LZz0gUqqBeYRerD2ZF
7xex0v3TcYYtSRmjsiYBu3An9G39pX6qQhVyUBhRZ2ji2U+fKm9T0o6zjR3/DEH6ydwXTgEbmskK
LllIcZ7EiASNws40nXcCg3N3jALfJnQOgidtu/ocIXDyvRZpU8x4GZzUCLQqA9yzq57VF7BGkDaf
tlipAg5eJZmYnfB5Gs1qDoS4ZCZZIYye7Ieh4s/sXCyVvupAIvPVp5Lg9Tuxfx5bzg4setKjswOk
yP+4zwXO8GWA0c5JZ2Ro1sf6yuxTptcmxwnE6YS5/e/Jd0tFxQBYBOkcQz3UOtj3ADXnl6VrXBGF
UazqEgMAMs96dGDg21+ZlTiUvCksIoqB1zTQXIVonGe5Im8l52oqAS6lUfSzb5YjwUa+TfNeikY+
Uso7FFNGbWMQHYtdTts0bBMXwq1hnE9AAjg9gyTxhuAWNdbkLqpF6hzAxvnW7bcewRTpbEkOeroR
jeBQPxhj1y2Ma2t9y9EBZKPgrD7P1In6Ngu2rr5ZRHob+QzL0vkEzd9yc5UbRdg5PDvM26QNOLqC
4c14nGfHsHfZFIKykpbK0YigKbig24YvhLPqojS4waYLY80+SPQdrC8qXA90qZ+WWxN9FiNjDw0J
LhdWNNg2lVE5FQ99KQXNPuHuwvZprd79SwogxaFnbmouSLfize+GZ0tejoLyTBDZyvpk26AWCWk6
B4BPP4Rj1cuLhG8eT9gp4EmsFx1mXI6p562AkrwaB+nZIYOymrfwzkK2wFfzQbsxHwFgbzfJzrin
l2gEz+QhQAN88YXs+iMAWG/t9wxUtz5W4xTgOVwIaa6wjj+fS/sAVePfgjUTmnPntyoJD0kxWez1
Ol8ZSQ1ShVJnVeGIna5+S4Mvq9MBEt1Ec11bFUsIYDGLRdUiq3Ek3X2WUH5pmXNgz5KixkQj5Pqd
NyKcd2jr+RmABxCw0eAwAdK39tvFaGb1jtRzZgxp+yj+pbcTzGJyJ2H+8cfDGiA1OfUDqbMT46db
lKlkUw9Ike1WYVgse7KmacgDvq1/j2k42KPKHU8IR628HzEfcrDkCLB+xmmaZ90Py0Wh/rfXz/1s
wQmoKHRuhWxIXX1CZJEBipJ8UPZSumIYUOdTo5KA91cHW0OQLQIvpXFITa5Klq+QJwOg0MwZym60
G+I3oxk5H6c2pAfv5XSZR5EqfSV7o/taNFDQelbJQ5fgv9hCxoe0cP6Gv7za5JB4t3S7Pd66kbQV
ubRKMluuncEwLmGsggFm5APIjpjMTsHghWj80UewrXOHQt1mvre27tYDSPMVQfPTR2J16p+nmJtz
1dIBiuLS1N59IRrm1sBy77n/1RPFxvLt+roapqleYC9ZhlTPsZYIoY0oIj0c81pAplDUNJYHTTun
ZF0jeVousbICGSKBzETndreZbGHtBv5X4kB6kHWAw3ZgN/cyd5P7hpfcPeKek7ZQQ7vaDo5fVFUl
GxbN8Y/X6YqRGLibEXL71yhDxQhFc4uWzvbquNk6II0Scbls4shTBxFgh0IlDADoz+gt2k5Mw2Q1
Bsos8Evs5KBbguBhqFL7nn5rQXoI48IU+Al2MmS2k54J19DQi7PoeotK94YOzhGD/gKGn1RELiRo
AV/JQDiyYBnjxdeWuSazqDzrp+i4GzRHq95SJASl43rlIBPVBM92vvJaUQS9SDnHepzxgULejfXa
uWRzjoS+ODnyL9PJYwqICxDv+l5gCW0IKM6H1bMVV4BFVk4y2LmcsvHBLRysz51C4dx4PLTXJ/Tq
jG8ArrVn2splB0QLpSMxFZ66Sl7977uqV5w11MeBIDXQuivI5bTjtc3Euj6WCIoFI8cNTYafTxt+
hSO+5EmPpnsD/CR2mOFKi3OAuR82Y4sqTUr3i5N1u/b+P8R7UL3Y+lGjH/cnV6Q/2ZtfiPfCsr/b
8NyA4sO7pcUgVb4A0t+2o39AMoWo/axA9MQQ1RO5TLIE+x3RDslnMUvcmlwSx7lvAkOq6tyY+Bt2
vu+aa+D4hlRSdSslzbknVckfiYnYSpvkuBN9NkmS2yR+3JA8N3gegCGQSDNIEc3AC97cJUeIY9Cn
zM3OzDk/jJgbQqraRmlgz00N3HGiNlPFyfZUVNAooUTvTINUdSO9Aj5PD5+XP1qNiYDgIP9BMBel
jNVLfKmUNIN6UJ3bkyI9A6jOMx/6Q3cdAVhdmJUNhajSytHHjtpnT/2G0xj6nrPPxUaSHQ5dnCQb
drS9HMpVD1ElimVVSC7k0jvSmWmfrzhMh0EunyrxbVy7s8lE5brEUu+Z+IOkRhzye74qmwOmUrLh
6fworVtCjsgaOSiFxArb14gqleRhAXG0dyTdVydwgGSsBCxu8C12Euwei6cUA8d7zJMbH0L6jxvO
z3ZTOOePQM4RMtPIPxmtNnQ114T92lCpglOrPlBqMqCrs6pzkzr+0rrOyhjZQfAUOpW58aJK7w8Z
+n7xcPxmpnpROmy0v6lNsT2s+ZrwbRwS49dDKn5FoOdyB5E5PCioES0Yc/4H9fVUInnxPYfg4SPo
wT8xWTa1jMopRap7f/81mmHH370Tp0G7YoKzkPF9tzlyJ4BAt503Hjrxs2DrR9shA2aSOaJmpuaj
KX3y6UHpg97moAU/Ol7ipi8+4NlT0g+LnkrTkOzKrLZsvmCu8funpcyIuHcInxc/0AQCGvw6XMiD
LHRjIUpGh+52xnNWlPDyL8ZI8A62cBgkDuR+9Z8hjdHfjGDu85ps9MMom1eKyJYHzxk07Xu6ndGp
+BWgmVaKhz9fE0YyqUv0jw49upIPIllTZIqRS4cRYbK7BTYYq0OT/G1l8RpOMG6wqJ/hJqhmLXAh
pKlQU0ARSnzRBqbY1vBqGSZ4lNDP1XODCjz7u7ZKgeaBYhyibgZuu2prB1CrmigCHZDBGXGmhx5l
2iBiHjP6Xk7WpR3/x1ee6oCbIRa/W2TZmF7F4B8GecjXLX7TO6+jJD17GZFHNGVylzgdDmJMpstV
5CONNaai6ADjhfs0U1lDvyaOsCAOqNzCfP8pMplRwTG5h4s3CWkCMQK1xwz46KMytKO+rp/N+4M8
U17JoyoP94AfCUc0+Zdh1vfWGou0NCRbAzDokrQCj+cmvikrfmEyOkOweExKl9npiobYQab93Wym
BQKyj2vRckFqWSg/WPqNZy9QFhYuis8h8U24Wd+2HBmnIeRQTkBwB/lPJtT0FuY239HrgGqhp4DH
uKKcEb/v0NqK3UAqPjqQMiOkNneVOVsWCjY1FbUBsiNhq6xpj2dCFdYBPol32qz/cWodrNkvSSgm
yoo+F4/gKHwEDeApTsNBj143HT17FiwcgQUW+ECJr+d4MlNTN8jurezgLAcV/nmYDngcG6pUWskr
ToZcESW/2JfHntbGVNAQhOhmCc3SLDybEXxigMwWYkpW1obHa/B4/cpAoDRrQRngtqkGVVdlGRxE
+o7Sjo/thjobPM4TnrgKTtMMPG+1MH4v7pJPGJw24ZDO4mhjYQBjL0pInEWc+cPbVOQun2LQNVu1
p3Ps24lsfC/cU47m6NM2LodK1fuvUwscBEo8BhUkRRkJy1P8PLJws6o/epMudFkSn8GTmAofi7fv
WrXj0BXaC4joyED27cr5Pd6c5wiWxWW+SdVB78dtFEm2JXd6CYD1TMvwqaYSvt8gIsn05AcjjnEN
RYuTlLB5PKjU7P2ROFq5tFJmpzN9dqEWOy5DwCGlw0gYygHHAoGwpDsIlCGN8Pdsw3jlbfrUDk+5
jkvdEh41hP2TjPY52yn01cbWiAtQ40Ue40DhyCIgaM6d7fSa5SeZEsS4BtR///JrZUsPh4+HYqPY
z9Z5lzu4VbCT41z2Awj7aElMDDjzLdjAXn+QptI6+wkoZh8Sso35UcVXdOJwNGfZ1Ht7heHQg6hV
NUgDg4hlrcYegCUEVsTTfwptfbZzPEArHjYH7hapbGsMhmHUQtbGB5g8/Vun8a5lcihVp1C/mUaq
c4QlhGCNWcbLHYRaMUtZNaLTdVhru7+hYAKm06df90cX+abE8cvRRQQQ4QPKkJzobL+bWG4J9d86
NCNg/fGUWny9VhY/4RH7K+1Ewovxhz8vdMfMFuDxHc+fqtzecdGIwsuoqzOdwK9w2xrlZ/AGQxI+
KHRA/+HPA90CXaIBi9xbyc2ZSP29e5/4d624eXsIXFno0gDUkDVI6WcIghiZWmHw4Wj65n2A+fCB
LlbgnDa/XHoBWRdwgrr61VZXabqjLshFdsvdc3WoSIx64fq9yMbFzCCWBPAgEbfKcgTmSEVmAm2K
uTpV9z2ZlP0sUIw8eAJ65SePz3ZtCNyzr/UnpJCL4mcyxtAY4WEt7VATI7Ug+QIu1BuPW93azsFV
PRXmfnzT0XuVgeuHaTNm2Vd3oWXb4EFPu2aM2/fpRPwClw4mdrY9/5grqf8xKGznxGP9o3j3hnFk
97hzqfPPruUebqaxsoZfpZa23w1GK+9GEY32f4oarcVUYL83RS0H1ZXt3CTvVPjq6ed2vC/1ZsVC
NSunCpCkwYUIYunrZ8nRoaoVRY7OhG5qSuy2VaARhzVmU1q2Uu3eIE1GIgyMorhaERn7trFFmJRq
vylv12Ephq4ZlLUOwEK4jZmciGrbWW64GTcXvAF51tCswsqE2XhXh5Hq50QE7WmUdM327I/lZX5C
JQQv8YKWJ7zWuHL1rhaWoMWu06ApVYkkzKpCSo3NKbomkeiliwHCiZLEF/QyNU1ofG4wlFIatLb1
eJ2rlHevB+cJMiWM82I3mochXaox5ceDXv5KjQZllFkbVHHx9rop8UgOnCe1Iztojd8s5EknT0cD
4NTYPNaxjLbpKtTBur/IbbqBV2GSv1mEfnFHEA1Q5Woy+1umjdxMbYDsM8g3k1f6hEJ7CHmfxVYO
x8TNh+BWpVvTpglZNhUpIEi7vSqAo85PLzvHPuLRrfg5H5H6j/OawOJ3V3LKD04FsrZSdygA3jKG
kP0r3IoaAZ+ntAAAarbfDB0Jrgx2gf6zeErwh/7Eab8JDY5PnN/4xc0lj3+OZyiTd5SQaajiSu9x
w4NlR6+nTmSIHJTAnX/S9cNfmrc1/8YyFcsOVNEReXvwoeM+3xaHzGKLuw2+PrezbR5qAz3ANHLl
51ZJdwBGTTiFOR952NS7TCKGOS1t4qjE/Q6NYEiW4pOvBwkSbYiY1NMLY1Oh2/R1Po5tT94tZr7c
i6RedPJQDzn+Ht5wVmjtgAF43Y+BPkrkYWFlZmky6ZREgcX3HoSmqAN/ECT1XbMPGTyZgqZ5x0Hg
Zuk1cAf6ZWKnsSnOfOixTgRRovdb8kB6ciBN3AVmOKlSzmpQmyd0MqJoTheauowVSBA2rdIF6PvG
9UMg3liZfn4t8LA/E8guhMEMU0WCnlAqkyuRYhNyLb1Qd/+3APzyEYJwBXw9yt1Nu29EXwtG3DO0
mg/UxGzbP+h9ziyt3UOn6+K1xskeRJUrQJgTaA2SOfw4NjnXZYPCEEzv4HGZ8OL1ap+addlb+IF6
LxKbdDPTk9ZtSc6OESwt79mcnscRqsEfuPMdYIMF8bJxnHqtGZGeLziAPC5sKYT6R1nDDdPXEhfF
t7baDldbRhK2gh9+FaudW77ufciCHRfMM9Qt459UTpoAe2TaKqYZXfMqlfilZ4/sTchIGJHCdir4
a7LwWCf17n2RZZqO/H4Q207glAQu3djaTKNJHGLlQyYafNkNrlmGSKyu2edoJXreTgbyU88Delk4
rHNvF+i67miliiDlg8pYQsWoCELX31h++c3jHQY+lygIzsanGuu17yKvsr35orzEbS69vW3ssR/N
IjqjJdVgwr/ixjpjV2BQm1t623hpbD50jKVdoflDN4UkEKGbzmXIGXczKfpTrf06fpK9qEBpzf4g
ZpRi5dFz26vTAE2Uy12Cg3qAN/TI5y1ca8zYJRn/0az92R/tztZ77Cq0n61gfvw8ssV52cvwUzp4
fs42V05hhc3NeEffRCepJp2r2TjIRKnUKpn+WDEmknSEOyL0gRpu3kGw9Emk3L1dsHNvVYCP0AEF
4scZxUwPt1bdMX4yOPF1sICEyG6ttOK5DnBGjiEXeKe6ABS+ZCmbl9jVIkeyJY083p69wWRKna8c
TU9Q/6oIc0w4psYB4kPlrV5c54np5qwxTpAV4TUzno7TvPyJRUqwOeOyTEOBVmm+fDGMcSGqFOia
30rsujDhJ5H8DqZRVGpAw06IbnOm2Uu7D5F4+WlFtkdUiYAFlypoUnPzut1psYDDAL54azhAyQYa
JVe25Agu4RxI6r0JN7Nh2TMcnnGWugdGoYDtBDGP2KX4l2Q7TrmLYw2fSepvTCFosJDf/gRiizAq
fErIsqPdE4Q1zkgnu2cjHgaY/epNTg2xX/ycdrUvHFS6MC0Pr0LN8GmXeNHHDyv6StxA17+WPWNU
zziglFeZW2yGCdHHP3fijfuFCv1wBW6G+r+A57XWJuKkSMuavEnk1zTliovRX4eAdKf4x8zAcOdy
LNDrPAEXW4onSzyjGg/Qo4E2sqTCfH2uDlPnA9HZP2p9dt6u3VfA/QNqw6djMc0UChspQQZ8Pllo
h0FYw9QoA0l+TOQdWduj0jP/RszjkgArxYSssp02FjdQrl5Faa390XxAvJ36GMhODGuDfE7D0yGP
xn08jjGaTyPRKdLymKcbPyS/h85IgmWQNTp/zrRJhoSuwKGvWgDcDxWyTWtu2eLO5KQzpeibBxV+
+Jrss9bmcPAd8p+/pPeYM+6FJQnypyZCiBEjDPgRAjoOq2lYFuX769g4RQ2TG40UDLg74x9Ky4Id
yiOIhZnYo2nDxgEJxqCip0JnB2/yfZg7UBc1h/y2T0d18ymmGFCY4L2zKcNTApeTtgrQcU6zOuIj
6L3Rqt1VLWxCnlr+3XckFscVfhbnxttEAVSYgZjrePgy0q+bo/aUMNftzY2vxXClC0W4qWC55Iy9
VOMq9Bk0hhqO3JPioqE8LvIr3ULIk3FOisv7gIogKuienOXDbVz1E4qTv7QQO0t+zoiZUHMswBQD
YNkyf/iF3Dy4fy58LWPh3Bp8T2NPf+2aZJxBJANCRO6aHoyBQmCakE59nkKCUmd48ouQfMr4gitd
+F+/cOgCRPL6UKs9GV6oT5XQG13jda8sJvUMow8t6IrZ96iMH7nSYG109+fuA8whf1Yv7fAnrw0M
4hyRzCCIk59Ns9iWTdOsiONXj9BhI8Dc5O53eiaO0cUo6/TAqT5thHZrfM8W059ke84W4Y/QGOPb
R5Hfz3QsEla42ng/ELtwNDYpo/it10/12xA4QE4Kh2wuEmL2d6UMw/9cNRQgptZd+ZkoeGJh7CkW
8buRKlW0VE8wpadRo5ACC3ls8Zhx6txXTccpANIlbMXDxPrMtYk8Z/IoGlD/QApnvl7P/4FbYTvi
FOJKe09SRY1emH+QLN/0j05BxS2AzrhQEX4xyJE5qxLFiZmz2Zisp+uqT4yat51pctHAaYX/ha7H
kSetbNSmyvfJUsvZz3xTLNX98RZ9Xc1GkNdjdmtFjoH1f5t7ia7eOrIlOFOx99bfRSWJoJbBfkCQ
ubHa7v+MTCF33M6y/8iBfciYYgCLRhPf8LR4MmxS5zWl5sdGjVDSNoBLgyDDH0lht4B9Xl+wggPy
EEOFvp739LlOO8MLoQtBLZhziPFKKRi7M8kN+/lCHui7GLKlDwr87evtnnLZF96Z3afALd+yJ1Gz
vrqd+F5PF6/egbtuC1Q9zPubiwSXDrgny+i+22xb3Ru+x33ydQc/DMKtmqpKFYAkZPB9EJHaU1x3
SNFM9klyzvRAbdEEsFc4fYT/H0zMmWr7Ub6av1OlnkQJYilRDSgy2cZ1dzknZk/R4mIHTugo1WhW
JWCfos3S/KG8UaLwy0nOCZEyXyVDKfYOjaCOuA+GW7UGYyK9Ey7n74zjqFHnANjjkdFxRP6JCiIR
iiTCIURDF42qQdq77oNLwkzCLWAsduXG57Y1NL4aJ6QvHrmvbaJXcU+1G4yWnbxUPDZeZXArnzMB
I2WKnUM0vpvuaOXU8S5BBIbDoAak22AQU9JlxsVL5e7J7k8WiC9wgZ9EO3cT+u5Pfu3pATvZVv9T
Sy+eMSkEtvISyFXOCzyHH+eecZl/YhnQW6USqqFLXrPcruUOQtfzHoqbgatE1MZxrzW6peVaF8G8
I0e5+LZUct3e2x4uRwphf05j2uPWsTmQjB3SQu3PTP8RnOy/KdQZZUPhoBBeDSNwr38u3ygr9BsA
UE5uIPd2eL08l8JDRAmtlXTe7UpDbNmvxOg8EB5rW3rPzLdrTZ2XlAbLwnt+DISw5tWLous46kIW
kYVSw/LghSNCeEMYjatFks+ntxBydEHGd4/TVJhFoPusT4Y4pILndh2kIrEt5ujLtYmHvCY8T5eB
s+Lv2AR7vLHPWznVtfaX/aRtIaC9XkYDnpe3IurqU5OW6w5JC4Dt5xRGC0sB24vXgc7voaXppUMQ
JUT/j4XrZgpYcK6pxaQtLpzN3JrbWnnCMhSAcnKZ6fsD0Xly/Lh5j5oiS291Pzdu6Pzf9XMY9r65
8bItNshMLfAkOof3cgBw2VoLwaYen492k3B5OwgINmRd+01XoNE1PFe+O/pZLxAwQJBezRkoKXTb
iq8JbDd/2KYbutZiOzR8y95Tn+mZLN+wkbbIgrmb020WD2k9muqENV4iFWmOm/9j5c1tZogvGMmt
HxJkuQTrHSzhvHoQOToemIzJfrQG9hqRwPqanOyL4uiaf1syF7HmpGKNE23/WD8sxmA357CdMZO8
O/ccOlCdAAaVumVQX+mhWcxVMzsjZDTusY9IJJqFsQ31eERcN5W9CMK2OeWRMy5gzwGgujun77jM
l2vro1PXrZ1Gx9e7Phoe+k3FWj2ZYwI6JJxKceC5mM+vWBLE3tO1/liSVQiYeO1En9WA+fCXhVA6
rdgHEZo3rN2VjbU0ZNcWOo9g2n+k4clEFB2oOGQOMtWbBZ0n+mPrCJGgeZ8M6ywJwZwI85i4mURW
NRMgEEyKBunyG4C9i3atJmjKfVfscmSV9eVrsTvNzh+vUveNBpM4qCzndCxk79H0UZ0aNOX50vdQ
XmJhK8421thAj/kYPAR96EacfUVFVYBdw/035i/iUowGbAjNTWJohH9lSeznpnrbRV7x1Gh3QP5n
gy/IemfEIbK7lRaH5Mgo4JcUvHOM150dhe5RhOj3aaEW5qPsBFtfIypayVYBeGuf55v3kkAQbxEN
8j0UrNXP7zVmrduvQmaT7O5DSqUmzqNeGWBdiwW95dyOT6u8IC+lk8hz4w7rqttXU7yvzWHvV9kB
c0QYLalBKYAUTAwm+TRRE1bvqkhio3RexTpxYilSCN1KxB9cmFJcVGrbeniQd8KHvgATF2jDIzVO
cW/GGr3rkQGDGOAV2dKwyhK8MxCzzt0jwSZw/xOncBc2kW6JP8g6fnGEGCwxhLJfYJl+5bBWJH1V
YsVNQvIzTD68rYOMwqmNjgZA9EzR9LvY6K6Wc5DSWn46Yt4jmHaAJLPmVlNFRHlf7VqfP/iOwJgo
Sn5xyaTh+bYQ7ZEQpQyUoQxXlCVNC6ZGKeBZmZ1WwMfLAZPyfgvTcnUqpK5gQ0IqlNHe3vShrx6b
7Gdv17k+puUIJAt6ayStHmXDdCDbx6qcUhyiK4mWkm8dIkjBRVmkL0iXkPJx3tbCoSj4pRoeYU4i
GHJCtIuj97aouSn3u7yzqk42PoMOubuWGZeXU1A0dK/cmRsdtRIXwuS44F6lxEX31ad9ig4zPIXA
S6xZvXxz2PqpI5/XwpViBdJRR+UErK7U55CGUiiFbc6MOxNGg1KiCFX8LjISdhvl+E42dhn4pNo9
RgKjaDSnsGhQ+mDF9xBQJA/afpBg+CK+PW8kqNX3wvCqLNwawqP3/OpWij8TT2AHmqSL9HrJPZ2K
VieqmCFW9bpVfXFzADXAtpdZaK85kU5EiaV4wyenY3RgiZNp4AwYNpVpBlf3SYHnPiFy5fDp2Xf6
HyuVFkG7loffi9O8KGcRJIoVy3c4kr9NJNw/JCzur+XAcHW7yx8Oe3tm0/BDqLx4Q66FsHkWAAUi
58HIQe9VMtO9QBrUyjX4dTbqBfsd3iANBQdbrRp8XwR5n0jNqb3dKSh6BXZEpCJAseKh5FOw+xPz
qtDRvIVH+5HH8Nb6hr5xnmYvZ/LFwwy7bM92uwbgPBSnqTZOCbQW3aQyCfBINqFj212GtA650tRk
gOMael65TN6UidCafO/KAQ7EKw2KKQYMvY6yOce3m5EUNWZ1usDmoOTSx2ME+o2PM7St1ufGcIcq
WCwvaTrPdZff5j9gzkE7uEyltS7S8AM2WrWCW3fSaY2nRZhU5pLts2BY8qN90jiRoaCnPgFvwI4Z
EkobFfzbvUr/QqggfnBqaYOUNUFd3JACVt82Fx0uYaxrueY6vUKwBo8zxP7ttopnP3McphmC+1Gh
s8KFVSlJp7jRuGcDji6aOkZrquZ1B+iHxULJJut7K5TqgufcDpSBL5k94i/yr/n4Hiq+RGmluSJw
L6jVhY1vt1Nvghdq0s1WKzI9R9CjNUuNducdUSQcFEB3V8s8tfMleOMDQ7HNcjeP6ZFstDTDs4+d
sWUwJ2lH4miMOiG2TxYtD9vKA6f48XBRuEsBVFvc4VwnG+FqoK4h/HmwpEvsvnML3XyGew/9kHZF
QhZe7ICKqtRkw1pQadZ1fJDVSG1ytKjlDTsDOOYed0eHZGCbLtx1pqoPujubHCOonlXHX/TH6ywd
EmEUc+r4+9ExvqrToVD4Itue+DgSEX+wwsDTPs56flFm5CXMdaOwLQVuqLq3FDC/fMvyN8uAK/uA
fjJKgLbbBPaIHkA7b8SM8hcabSFzFW1F5iv03E4dt1SEMfadMVmnRHscexc3hqhlScKEIiJmlB6j
q2cJYdPtPe00GxoGqXT8n3O8asQatnZdj8gmtmxsWXACg91QifmLqyPp8zz62y28sL88+AKQ9eKc
7jqJHsZzzy6e7CMvhrT6knKGxksptGgrw/OfWSgDFq4VVkPGRTttP0QvxFiIDFXgep0DVc+36ijm
NkfJO/lDPMEcePiguyAYrtFw8npOpcHWz0VDP5T+n5/UwPXpSRGNZv+iDsJTJqfbhJzk14HXgCRg
ZNaShf+8ZeOrQhTq8b68Lqj+6e2tTUf6ph75l/SE5aihRhgjxYVBPs3ebVgwWTLAnIeQ1IzvTL2D
d0+5jxMweCNnFCC0KAIOfu63U+t/ebPAO3SpOAlXueZq6EUE9/pAvUd42B09T+CUdtl5a/Aja2PM
1sEn6xOAa1QTZKXH8I/DrW+ganQcsGw/hIcAsV2WXy1ufVlNNJterLMzWBALTvGBjEYGm1KU1Un9
9VVgvWj581gpS7TCwlwOmFXalsvmE0WzzHnRVDfUg4YhNqtDPEFUxa1HmpF3k2V3LjDFAJMxtWDD
eVF3wsA1EdFgrtbvNXZ3IFVbOVkLGfsIuvj8ySP904phNMiR7O/SWPkTnRHgAtFiYP0Imgzo7S0C
FPx5Mw+Crq7Pr2z6fMienttCslNRqXrqFZnAAQUJbaAvO4KpJJ/Sfwd/hVO5bkPLh1cnM1xHKeMm
9X0kjn7jeaC2nvcPo10A2uYZspdsyjfB3g/47obLzeLMBCO+zCBbeyqqlA0z+XBcSGtNZjUaAAon
o7ylxUUsp9PA32GUnZui1MHVRkmmFPWpxPBXPzisrmRCo6iPikhBltLAtnNzEkdVVok1y245QRbC
1eCGDd17Q3lFOjiRXzTkR4JjjUcxOaHUWWn2Yhdxf+MZjWr0gJn9+bMwcrALC7vdbIFPNwJmpn/r
UfrZMF1yuDDNqzhatkZzSKfl30LK2ZPbBSbaeLEUFJ4Dhw+h6LrOLnufwoTVIj9fab9rM+5VTJ9O
G3oH/copXuQMIc8Pka5Cft66SCy9gFuCzGwGpwzea4o887bxF1E6rT1lYmB+0Ieiw2Z+j0SJNBcb
2Go66fXzRRXl05ynNf7eBwlLjRbXxbWAKFTmmAh4YOqRPkhxOixsiVCuzrulFbRCCWUnkQHfEonw
2jXyLrq/+St9m4VUNY2WN8UmMFbrgyj/kHrIE47lIS1eB+zz8SNkr1YVK8UfFfJDZRQ2dOdk4CMH
1M6rRo86+Cqw5wt+LFcz5Lox9ilzPP0jeH80DDCW7hQg3DLM0AeUQapcnof+oeRqYDW4p8Y16NXY
GJYWXux5aZNs//0qSvEC9DBzOsMKtCYEZPVZ6ZphWG9yfuuEy7rE2ZCa+I/6UhUgVnDTGPMWXQdr
A/1rEHBDXJ2KGjfMeJ+kct64eK8zVm73c1KzakT5psxlRM221BccnrnO6lkExKA0zhS1xYgwOI04
rP52NvI2ZhGPlEPo5AA3B3zr0Rj76t/d1CKZsZev2Vkv8rjX65iDiZs9PwRcRQj6dO6MVpGMd3dJ
gphX2shhX9EuHOOZMhAagKJT0zUZzFch19otoF+x4/v6a5MfFNHlLjKqAPOCJGpV1r0ypWYHZ0ph
MXEGqHpW9Z5ZKRnVv3iD+f04aAHOqWsUUewRJXoZqAdJyZnBNVn4pIwmCtkDo8LTv6KfSmJFQYJm
k08iPk78JmoryqJcq4++xuziKQCY5IfvXIkdY8y55xiZU07VSZtImga3qULGKkVyqckmju6DUexA
uZFH/Y+1RD4Cn30psno2RyRrexlLWpXJDoSvVwWCsv84xnkMEnOKfNUvXK8Iv/PvhJoFZoX/wI98
dZYPFL1HtHdqNmqv1AyfSpWbMDErAt5WO3OE9MzIHsT2gXNYOLNTBfZPFtQk5ForIkNgjzXRn1dB
d655CZyNu1+ENP9WV9oNSEXIJueXEpQPAdBvOwXdK76qxh5T1swhgWlu6XtWB8MR+9CyeimJS7/a
QvB3o6XOWUJjTdryVt9Nq3R1PotE2PQDrCJ4ONMFpkfHBoZ7yF9CNirSOCERkMZCtfD0tMSaCVHH
mzdtZ4gvg2oq+/74g0cXvkJxiI/XSZOPnLasdepcT7asFezsR7Ko6wEOhdDN9oFDGNT/Pd3mV+vy
syJDZzxErhnrvxcWv71RyLqT6xE/oGyjrmSojusPW8pVj355OI8JQ6Vx215xNxLgxXSakXRp6LLA
1TQA5JoXWPKkvofUTHhC6XtRJVyBhac/qFwE5ejKQyQv8opWBxzII7/qCOXa/ycugaMVItMG8wh4
miUNfKSEUXn3VqgyfSetO1eEaPVuWHOiixDXX5gU35r0BFpSSZRRXsoHxcFE4eEsVDnzSu3A4htk
mo3uvtv1bY9uTgJ9fQQqmU+iczwYMgXjtdK3DkDpKB5Tu2c31LcbWjAJQyp+Aof1dVkpXV9esdTI
szqaAghtqZUOkMjfbRpE+1um3GoPH4rSmt4BedYc3nG5ED2KymhT0DrH67opIuFy6X8u9sqrv48C
+iWmAnAVqKajiwqEn7/qWnmJBn/7sOD7yBrwcIL7Hdwi5lIVzl97B8L0OG9LzGYTgNQBFIcxaeQL
GULprxhYT1cv6kAtzmaUBHb1Y9OTdRy6HvqigmPx0d9iI16F4Od77VsBCTvJjuY42uxBy2UnxYF1
1s8/cdfVNIUpPyuEGpXXuTCxTmLfR4pxdbgk7lm98UyMMrQBO4JcUMiqwBRqWe3P7LTgnmFLGskO
MlIZJXhDAl2wIaF44OzDe/32v6YWVdL3cJp2pKhQSN1DfJ2TflIIqaBvXq6dwCBqskj1wI1MlkKP
NDqXhj6nvo7eckB11zBQ5zyrg7JpusdBU6AES7IslRIYtosy3FGG4XE6rvmyGha4Z7u+5r6ZAr/I
v+z/fug0mHKu1BpiItD+m2GuZ4rxOCbUN/q6kOV8t+gXBM8lERhOGaWI3OV4RNXTYMUYJzDcCDu1
FL/u52DKASxJQl9LuwQNQKhGxIqbZ9EUHc9fRNl5lk4XVUxE93Z7B3oaOVcc4O+Rd0XC6CVshwZo
8T1WORCAW2QxhloLvAlkyfKpGpg4FxK0gGRF96cybzDTAMvGubJTajSmjWsjZTVf0uzsHhQ9TMvI
TWhO25tF9SszfhQZov/XBEvyMjcPce66dyGw6vxOuWSqq860fCO68EV9mFlL+695ds4RRE93+H6F
8bSD4Z6wCWeqfebBx/Tk0+9D5ROBXe8+mOXQrZp6wBhgrYwUHEDPcSKzuQU8Mr2SGVETsjtiNOLF
9R6/IpyeRLoVAAp2sC4twYFCZr14LJBejDDQoXYOmSHXE5UOXpzFbZJLjqZKq84CXTrfAHzS+cYY
kw0qv8+LyWq4ZMVW6gtBq5CM8kLOZbPw7mpGkq/xYH6cAtflcasEGetDMZuUOWAZY555Up5Ts7LV
vVW0EREW+FfuoEOPRAUcQVKIWNMoSlPR6VeLAZ4QkonLDIrS+itfhPLkqBEyjuAI2Zq04AuD1beK
AMkM032FXkGOjwbvgDJb2BT5POEVS3ApZupHoxMmCh42SvgHLPsrKUBKc9+RsLHjzuVncKuQsVYR
o6pfh/vJa5x1uL2xYn3jbqMUtUzrOQssotahxGD8/6gAfsgxIthNr2bSgPKpDr57BzOtVTUZ9nli
kIFUrJb9F9Eyq2BB/2z1VITKM04duZ3XOZki5mGXUJgxk+34RuuachzCC5ycket5O6OySCh7a4eu
e3iP3T3z+3DHyEjDDNMyphKha6ImP5C+Ab/VhpKZC7fO7rTHFDNErmFQFVKgxZN46cmkyQNSE8Wd
U/3fU0y6IsbRmi3UTB0Dwkn27HbuOSMxhhONgs/9F5opQichEv7vaJmdJUX5tb/vM5hm9CB1LnRm
Ipe8C5usEaTpi5cMc9S1dY43UzfDVVQdvymZujntgCaM8kNQNlCO5QPNv9ot4nTY7ebs3PMbUQ/z
ud/CT/Juq/12ySN658wQGG49AyUEnVAumg+zQ4zxNo1OqidEJ+5Tq6MOuseKJ+A51pVsG+xzsGQ+
aFXLI3R8ixATwBjHG9+aIxJDi6egqzUOiR3m9fR/NFp9ASRS14Hqa/q8aktEZ9xsK1NxAH9cDcDz
0u7ksyt6A8pOHbBO3ojmAvcb+ezDAwAuQZ+EjqNIzGa7uSjuy0tGIWrr+qZpcT5OMb+xBRa9QVHt
tqikl4Aqk4Sl51VlVuBQSyzR7oB5FT0Hi5+ifFsJrl6Ulrz6iTWrfFeL9VBw9nWjnkV/F1OtQ1NF
8TCa49Bl8oHKmQClJoMt3WihEnibcrU1/HRzWPwG65hf5rqFx+32hej0R9mB53oG8PW/rZWEAVb+
xVX0ZIzY5E9S3CMMkqgwf++XYouBMaZq2SDc0HSyYl1AnjKXUwmxPkjjYSFdqr5isKe2D2oVp2q+
8uEkNwi3qgIrk9kFL1QGNLRgUjHfPw6T858rWzblRW0R2TAa24yUpS2U1ohEDFfmM6Jpr9UaW09C
hF12JOIsk2mYj91Imupo2tx/UnJVzuYqfFZysjDdOZCi6/5g3asKoOFk99kC8rO41TDMViNIig9n
/ozqQhmd3wFTGP38YR92iMZaX05poi8Cfe1mQ74I6ZW/IeLOKPH1bW+Y6/iGWdQO7MjVdwJoaljf
tgDuma3oiZN9OpKjeM2g3DpcjzgOaaIbe/sAkWZfTHyCjOHsgbt0brNG4Rvp6FEm4ri6BrJOAjKF
sIesLLpx3tb++pP2y30j1+1CTR5Hs0/57T49NGCZgCT2fmP/NpXpfxDgFLUTPXVBwIhOHjfDvYnQ
RpcWm0OPwsA9GVZnPvG/6NY+3nD9bgfifJqyx3D5U1GjqNXaGbOlWK+kxjgI6BKV2LZwo3dgeSWl
x6e0JmPg2DNEJsvBNNq+BfEirqmhX0MRzFuUU6vgby6Z9Enxaq7MpflrvO/dF3IwvcVuFtNXur2N
qy4shRfCn+Yzq9mRrwkm4iKwhB5JvCTNq1Rwum0lqsDqeOPZ/UZY1ta4Z0afAsBcjW/Lbkk5W+wW
+pwWE0fq9QC+m9Vq99XCJZyjaBZg5HYxH7zkJbaTirFrtAj0qsAlvyK3wtKA5QffZeJe2rF87taY
bhmMCK1dvaJY6YfRWjecEcz7WD5LQuMXbgPZgy9Z8uxrq1zFp/GuV3RoFRxBCfwTy5uvbLcC00tI
GN8I41ja4Lg+reLG2doYITL6EbHhQhTsSzSJhdzeoD5FfD2Y4PTfws1nA8n98aOBkDWK9Psp9vta
6rHke7pLo6C+H1IFkp51hx3L+p++Sy12nDmplpi2p0ApVe7jJ+blrC1Ih8XsyQbFpoGcbeHJUl6f
oi6bSyCqxqIQlqe/GB8MwiFtYf5nRzdp3b+N7JCA4yEc4LMtb5/yPeKbynU5TqgElMHjlkVmTnq8
DJ7H4XQSOWVsvQT0RKZd7yPuZ3VceK4REEBlvFnb6EI1IG+kI3Rmzbqa5OrFWdclkfOMHMD2IoYx
l1SbzgNKoJ6XqktBswrCd34YVnILTksdVlHCUy7Jl1AwN68D9Jo/Wlnb4S73s5H95UHfzJLBMq7K
XUKrXMAeIxbloTD/lZEq2zzk5gU6VJyPNTmhsgXjxfn0ptWo7yUHLi7ee4bsj6iOGsX9DYGqnKmJ
Kw3suDFbbsr+QX8O6asgLsHdLpQC16FNJUa7UWEOP7wgxvDTWUqmv5sbHwVYY8bJWlj27Kg6vfXo
ixN6r1pjmYFNrXRTm+4LqU3AV7rCXGsCt7MvZDEBoaer6xtz5PFoRvbV1oTJu1fmmeNBxRLm46x2
H9GFbJxPwQBIaKti9kxQ133DUP1617iaiejzef1/EAGmlc4lrWHQqR6q0HmRNLPKrIhR9WNz90bD
upFpj+UZ8/dxgkZVZBOniTV/Fww2LFAx1nGUcX3/pYSu5zshhbTwxmvH0Cx1QgR2r6rGcaj4kTwY
dyJxfCoyByBxbyb1GkL10g96+z6IOL2r2Aief+m1asYVhX3MFiTTO6laz6ru1BLXpDl7RD5HeA8R
1AqD8z8SsNI6Qr2/maDAbXAq2MjNIxXi3zRHpmRwJhQ9MQN/tJnMhdqCM6zL9R02IlQDdPb8FrJe
GVppRnVzE5L1iA2Q5gxPeVc4uK/pZshkCe2fap9J+AI2fJUIulPN4RY5WxbqxKwMs/brRBuUhYuZ
5MZAHfJi4uTAis5I1do193KreL8DQRwP0v+jt6O/Sjc+0sW8TcKnbbdKpzyYWENp8VO1lGGAeeVe
XIh2xIppADidtYMwBmrG4Q7//T4r0/AlH7FsWTVdCAjcGKfUqKoQ7TcyyckaAsaI9RHorAofTMyF
NDLoC5jATZ+HXcJAT+EDQXDHYu+f/Z3+NQxMvpmlULQIsBv2CMVFu3X+F0HyKqLH1rqGkBOPQ+IU
21qrvZXVbm4HlU4HQvdkDK19dXlQxgVDeBFek7aBIdz6l3J9kz2OVruF4d5WGn55sK92nD4f0VpF
S380/FJxRZ94BpQ1m2qAlm9osM0qSOIRe8ZOGmkJ+yQ4MmHlD3uSHu1NVDEpBRn+MhA3Fm0Yh3Ir
ZpQ9R5tPVo7etw4G2t5cFaAOnxIF+qiBodDCmW6qRgMDPIgP6NtuxwANSIM09y1UPAS0xJfew1uB
WuDXbCvOV47NX/teJNadN2RiJIY3fPkjZxteE+zulLuLd6cPNDM32Se+McfurIeHUG1R+ZikTdKY
4/LQwkBxOY+J7ydLgN6I2tQwOJaUYf9H7O0JRGG6MtgFDYxXIIT7svouvloSAXVPP2ky1KM6YqSF
ht+FkITXcWHDFESZfgCFHlCvB5zYNzHTecHe6xvnnyIvlo/aFxOSIfw0KAOnNFOO4kOLjEqy2uvL
bIEliq+Y542Fzh2yagjZvZR/qPZt2ZXvvdo/tDg9XO+S7ckSNoudppMXBphGdrobdLh+Dq+bsND9
aG/Bws/+UI7S1XLMMv8uWgMr+Ayj88UlyYXl5dv99LmmsO+kfi4mN5883D/AQutWtdNYRsP90/Kz
4MSlM4nKne7Fi4c41qwR+J+8sFzoqDkgr0KLd9UOmWeBG5TmJsxhruNSJGF9qT3l53s5iD2nAHOu
KGJRSub6LOOJJUmPpVNipYN/hlRSlLbPI9gEaIQK8Hp7F5bn4sJiyuPPyS4SZIxfLR7ceFJbHie5
smyBRtToJs5kjMGlOCxXDjIT2XKDFgCNxGXLJfxZjOvOSdp9vQDQTFINa471BWK8MAJ8tooyfdc0
UrjYeWr6gyuwUawY+hnTrkr8wn3K6KPPdrP2WmAXmbB8veJgc/2rA1NMnTdUWvmatmm2+3p5zA1K
q7jv4lgI+A1YAK2Cdht6K/Fz+yrf+zNDrzqODOcbxZu3fiy/RK2o5nQwR+jICaBGA+f9KDIuzp11
Qq4OHT1trb4y1VWAna9OBjXLmkZ4sUaiwl/1nQnQlRUSVKtpXSXh1j/fTUkUImTB9pLP0JcmLRZd
wvXRnarj4LJ1/r7f9XQa7QhyEc7hVXIXryGbx3egHxRULX5c9HvNkwRdesPako31ZYoiKpLSUS5p
XDI04cOxwJhVWrqOPLDuaH4yHjUpHD7rVNsUJv0UAMDoq7kLqGx6+Vv7pfOJyYllxtRs7f5iCwEU
qd/HKQSAyNWfabkxMPxKh4g3K8c02xaeuQSOPjFXuE9iUrzx1NohuA8IvlhS/M3RFwLSs95FrZ3z
1xk1Z1OF0nX2ylUYwyEwdNmn/B22hBjxTAurSu2iNS8RBkmj8Yd/L3iZYcVdiptI9Yst1syx3SFa
S2/MVu7TqLsO2uee+DweP9bRnUymsc8QJWVNNiP49aTudhLLn5gsIKO0ZHzZ4dCXiQqjwJuKGfiM
Ro3yLDxRZ+oR7RS443xwbpMlHpGW2vzyQhaRW8n1yI7ffwjNi+u3+738hM/NburZtsYSHhG9WBNU
o1OknYH7ZBF5xe7mpgaxeNhSw2iAKrD7xVFkbtDl9iAxl7UM5dOkUfzVxHLm1dZOsnlh8fyeZg72
XY3rD8s22IDXbokuDWAcp5d8RneSPlpdMdW86JMQLbZWEeD36VLFH66t7EI9KiRXCDdOmRwJPCX8
Ksxgg11Pxo+L983q4JRZk4Wx2R63E1vshgVS5Mu8BHQo44tEy5/a3RxzKJ+cakI4jYHT+TOFyuMr
AAu2ciuO6zOk6HOHJp4Gia6u0DkX1ymv7JlI/yRTga1GgNK5w3iWmMlKRKtkPSW5NT8/H8DEF1xo
7iZNXW7k6G9yu3vhr31FanvrHi20Bpo/k2br4IkCKGKXyiZsu15ZaRmnQUiNLld/JlUhp/CafQ5t
stp5+tkx1xtp7XmWP/ZbekUe13wsKlhVodP2GrSG/Si939EhCAySpT4ciMF4OjkYkeaNnUk0v9eY
lJ2hJSjam4BX8Ns9TltrhBy1NNHSvfGHompzt2GOqPmBFb2tCSDY2fEXTNz3OLBMgXiRBCkriMzG
4BxG37cmi7bG3LrOm71fTiz+j7yh7T2q2eJKi6Q5sOEtA8D3qlG13r2CrLJ9Jhf3qfKA95cG+cxS
/kvIynwaGGDY/xgaFRGmxMXxogB/6lhP2xTF3Y2LnRc+6wxmf9Bm519ukAeR6cKdMsDKLaUAAm3O
4aMAK0C2/AHmVKYCOofVwgkh6VTwOgVvKDp37rhGYGghO5/0Qw12CZ+XloI2IB8clvEJOx7PXa2A
ww2CIaJab1CMHZrFQf5BLdb3QCDh6Ktz+Kw/1ebzkhXKme1kjkeGmBZUrQ4vQxdj/NkssprqyC/1
ixzjVTTAz8QCRCyY58qc8iuMHjlygvp632FhG8vS9rPeC7wTOJaHTpmZDtfAWphPI2BD57Gnyu30
BxlN8nF2NaT1P05hZiVkE/LEDPVn/Gh3x37+c8eFDgr6PMI93RjH//Up0+FVIbf4m52CTOh36P0c
oKsPcI2x9Vz/sBRdvEkv1Tz1CCct9fst/WEcSeIerruMPuy40qhkzwTIvGwFLzPEa6cyHyGArF3y
qWtWEk4PLaXEzVAqg6Kl7xuOjHYfDBVuoMPjt0OQjZUl6D2sy5nAzCK0cW0CZzkzRk87cbIl6eGs
kI8XGqhzIxjUMHQAuQvyQ7oEklM6wi6LVSVUNUdaOZViDXS8MsNkWDbFfCYhQNzJtTr7A9q0h6TJ
dL8lFYw6BEMuFZC7hPBGzF0KGl1z2nYTMT0C1JGnSmELbJbVzCrgEc6zGHYfFfEe68wAuSSok6p7
PrtF/r1+mridbhziLCGRJuxZhtevDIbF1QP5kgGH4HPMfdor+OTx6ioQrczXDtpKEd2WEgj4PLWg
J9bXTYxocS969g34trACYaDM6suFDCDI8pJzJyjycT9VuKdwb4f+qiZVdJOEuQuCnDD94B39QJHQ
XBUyMreYIY8WtZC+o6cBUeKmZ18NLsXkw9RE5zyCuSQ8fo+9VVNRFqaGTR5N+ZW5UsHm+0Wc1yrv
16f+VDKKon6qYbzSAIrzOez1PaWqRm0IqnlRb388xzeS+veEm+JozLJxeN6J7YN5/hVuZJjFMhgp
34iHPhjWjvca7g8Qrm3Xm54C78l2PGFRJ6PGi3pFoX11XOrKmpdBIgLKYdP3GrpXzeqzLQcm0UwT
aqlk8RyTB4rvfGiPQDkF3nHhqqBzv+oNjBkr9B/Be7IolGq4oU8n07IUwDZALSF6mUp4zFTArYqS
XGjvENO4ecK4RyW6RBSvlwJ58XTIdVEnAAWbzV+HKfbmzD3u+r5BvmpkSBeBLD322eGhZXGWuaIa
IotlKI3hy8TefJ/MjH5bmdfOAbbuZciG873mQUUtV447aJqVLdZlr1SBlOV8iei1wRQ5JFModmgO
6Xy6/itsWoh/9ZTA6pwjtme9HayE9KqxLPRtJxzxOBqt7JB9NmpjqB7C1zQKNSnTNuWiHAOg+bf6
qh9C8DQ/5TBlCBRUsZiWmSm1mBqImRIn/NBojLEVv4g2ZTSKsDXInz/BLB7uPSqYfIyaNwbuexNh
4a5eeQ5CS1fa/H4Ju9s9Nhq3MuM6mS7230Zbi5aGbhqIxXqTYncLFmdM/UQVXsN7rF9HpXVevdGb
JLRa5lQUgKJOvzuB1qmqMB2uq/E0OoXxffGauSqo0GCcIn6+GB3ZG7VWRfAOIi3Wtanm+x1x1QXU
iiob0eQXKXGru3LeemPBT/zwhNNKJGZm2lvUZTFU598PSZHk41obVu0HS9rO3epnZb2c1uR92U8n
nqd9NZ3YZQ0Uvx2tCFlrvRQX1OwEXJdfthuSF6nham7H4fsssWWY2DIdYkkxonXu0FwH3UIVdbD+
ml0jZyxQLb1XZcWVD9EAv9IbiJ7cH3RjVGT+Fkk4vBYYm00U1OPeZ7kUo8yyTPpr9GiQ5UkiDvgW
/Lmrgs9cAYRCQki66MjkwoGHIr6tgyUgP9DEk6rI5UJujhfhtusxY1Fq0MRiYoxC4qvfifMP4eC7
XnmfM8eeTgtvuP2bik+WkrsjeqHs/6CUUjXUXmKeVs1MdTASNIGJsGVBy8Uo19tVM1G6pepxo3D6
7i3uZmG4CXqDPQNmvgU2XxprVi8+yM0PeKvXjygJgEKe/x9tdbZ9/gqGKKxri2zdtmal+7TQGELV
iI9mWPFzOKj5y7f/GVXabtgOibqg73BqZFi4FE9Gl74DhkbSSiQtsNYfzGK8rDWP21zXskAISvRt
2HM+z0R5Fpa59QgdUgdPJpdXl1ch/qnG1uGIvmi3LFPMM0KmmfgzKsDZAriYOsfOszbV/LCRrIxY
1ifamsIj8HMWvSCj8Y6NuPyRfDErAmTg46J7haCtVuRw6CKKwF+/t+Wt+YSLtOGpMomGiDYB9RmU
L5bAlON7A8y73CGdbaeXptV5oos13WFKE5IMuAyegZnvlrPoa6Ah5EB97sIvkrCep3wz/G06mmej
6Ykn8j+F6TQNmfe1yqPIkoCgGAM+JnI663I6V+oLYoRm7AJyZRQ1neLQ8yF628WwGKxoY1GSStfe
utXeVO4Gsy9PLeK4tbPRuNx+RHMBtovIQjhw/9V2wv/JsolEOPqsahEKhf7J0ND4mWRmvSVeGEQ/
vv8ULg7vY6DQkAc76pY+TYUU4+4Llphu6X6+Si9i5nYZCVQRV8hrbh/+I9arMJnm0pSHuFhoKjhn
aCvxsOqBA9/9vDSG9VepOUuX5Y9Uorls+OdeIMFkyETdJAWmuRCxwldC3beAOI6NH4Hvfk5TTdzm
g8hfNr69ODzJ9j+wvRIhtD3gcsajO6BeKXgFxCe6UZMaTg89QmypyQIhZMkJpdcsIEKktAP9wHHK
2IDOyCWN5MhJG/+RivkHauBn9fzEK3ESgt8BQChVdb/vyylLVV+88Ipp2Le1yo5GAW9z8q0LzZcO
23y/aoBWZl3N2r/Rkba1LgQAXUyXiL8GfiGx9phTEw7WGPPQxj5pOSmWiBZkUbV15S9fgdim7wzQ
pd9HG3hBebEXVH0Z6wnRIecmgGPEAg1fQQ1+Domc30VKALZ6f772BDd3PR3scOWlWiTOHL0HYzaq
K/vup1tyQTtDoTxKkNK8enNAe9/uJ13pC43DDr4DrdLsAh4CiZvKY7K0hhH5RUcZEkzN3e9iesAu
5oG0bodaQYVnMa8ZbPJjNCXOfeIl705njQZsg3MPAagsixRrpr+6th+4VyZRKfyjumaOXaVhshX8
UtatzqfZb8dgLNb1yqSm/C4uQLjlj648e8xgtOGx/EzVjHEveYTtFLSokXjzPYt6JXhtZOBVlYQ3
+03Uy9y8pzItNMnYY8YzwWasa+5VjoEvbkUQYyzgSQ9KwFOPonnc57kJV7GuYpDVX5KkYJ7QZjPA
vAFV1w+lJuiRK+1idy7teF7iI/5SvshbqOsiH/tNCL46cYE7e9o8akcKr30CaAReixMaC+fkiAcW
FNmXmxT6PRyC9z0/HlMtuAfbqNnbCD+L21ICoXC3fmO/RI2FcTnHk61NyTuTtpJQMIqHHyAVv9v/
UgetMXd/wuxK45NcEvc24k/KkzvdlHyYqa7rsbH3iSyoaNXCQVoK7RnfutLXFO/ElZyh+P/Vm5x8
CEEYm6OSJngUsDXVay/1b1bz+op7NzHSIG2PM15pcupJxZy7dev01zwdxV70raGCXJCBqeDP1dYw
8fhL9f+eJJXHqt4s9znnXU2mF0KTODU54Dq1X5le0kolkcSKKjs9aSJgJRjMJEry41IudDWlAK6+
WeXFzXsby+F7TXpPDhUejM/WYSh0SVbfwmcr+36SNcFJMKH3C4BhVX+hUh2qbafSK3DHsORp67H2
nz2d+uluqSKQHdag2xPTNAD6ExQ3V3dQbGh7lF9pNG2nbC5G6i1eWuLyIMG4p6MA+mzpq3JpmaUU
dfwUbYpjt6JyqGXgxwixYNHjkOZqVb+AkNjzj4wr5li5+tP+raaBJb+c3XKkIWjX7RE0SxDAJ+D9
khfunKz+1Z3kmCwrv0IZ9wqtU8/6sH/QHat6BvzcloPDLX8CPNZsQpxycvpXSNBKM2yMgRYr/GZE
Fp3DnBS73iQaM4mI5ZkuJx3Jb5bnQkXe5RInEeUv52EM9E2IsbU8QsuokMO9n0Ba8Wn795PxtRWS
jJn3KhDk0IAuhGAYD6ApHp+P1WCl4vTZVbe6mWMTCwmYeJv5teTu/q1TzpVrMWfT+lgLPg7JoqG8
vHYC6VOCSgEouB35QWuYMdjBjkFQA4ksKQt0D+PSenSeMUfQDyaXuc9j1AFxtxWEiceGFwchMrG1
UNQfv9s80G5ikSS1GtsijANKB1oMmHujkFHcikVv7fPWET1SckBUGJI5JO0UhQMvmeTv87SehvwL
x7yOvV+2TAAw0IzdjCfoTLe2yKcE2wyxafYADpn8SIroGgdw2MwrzIArKJSzxWf1SUZ2ceeXP9YS
Hj9x8ARZ5kNuHCfnomUeJi4vAzT371csBf0LgSR16SC3yhFxmRUawJNvR0v/6PVJFmQ9HGUN7IfK
iKp7vnixJzQf80NwbNl2LOxCq1xYrI73inO89xSZER+k/zQlNzsI/3z5eEAkw1GsGsueTRMjzi7o
XszjO3pFRdzOBfBAK1ptnrjkf9OEmgXOtz5H8xsfxPwto8jmaaOR/b9yrY28D66kmPyVFMjLS4bQ
DnQec3e3l7Xxa6tc/f6PMYPKWiYDGU7cSdAYDrY2OHXSQ/+K7o14xbQqwiqgGmebaCY9cZ0Yr20P
0s9PqXz+RbouKNKdk9Swh7IcfiqKBgcSJadwQ5sz8caJxo5pK7xLx5nBbAfpW0cWTdL4MgNHhyab
s1FCHFgJ3TakKUj3w6Ok7yLZXk5nQdw4FOR7ShMDJOyXXV9qzdid2x54ett+pDgnGapNzYLPQepc
guS2vIA8o69fev7wpEqZaS5taS2RWI4LTHBE40EoAT5qde2gpRm7LBmL+S0O2E5aUbNdyzfjO2zx
jK6l4ck/EuoLwvtCMtyxnaQrUMfYYd4hSbI+6ZjTwrF7lk9pTSSSmqqYn/GGlhUy1yUCKsF8A8SC
MV1row7wfMYWxIvDn2PzBDd6wVGvFTOE403OOujLjBSjmOXslAbrM/WG34ybmdlSFhgjuaeutDc5
vcSixttSmHmui8Bn4cSZocVJkN8nsg/RzkOlHZWdMZM3LeskL/+2xyOQpbnnNOEkITl5sDB4HNS+
T7UV6fredm4Hkq6JUiq40sYMkS1UCjd4Rn4ySLBVtzEZqylrr3gT+4zkC4HZp+OOSbnB3K9Vk6Vv
B14IMeLnNFFqdWMgyGGvCN6pP0icmIwfAzoXtwHmjejzHmfKduAc4ACktkQaX+wuOSuDIamP/6Lu
xwDjODI7EkhhbXzb/wgI/Itx1sTEj3ZzE6toIuQQRWExT1MHIcxqekRGC2KGnG6FmboeH1yK1NwF
KJnJHRbbPaCial0/5q4GiFHP+PZJzLH1l6BE89kaUoDxccnk5xcflhXgFBdsgIRyGwnXlBG+oFsC
dNnGnI/MtNeomgea5adpJvfEqFRNWAWjC7sTcX6wJvj2ghJqBAcGcu0IY1yIYVlTiTjMgRLGufH6
9s1+XkaCInVND8HfR/TFb3juKQNijf0FqkTbbgZymQor2s6SmjNBtWMXgQgU0cpHapujn1Re9JDP
cVQszXUbstYGUyWf4s6AkNUdu63X/wH/WfGbQci7DkmqGuB3HMuPkXbLARpW351ErD7HDvQXbCcM
PL4OyBPEdRIT3mOegCLBy94xYEBDgpeuCawP3Omuttjbb9VjPVW2D3xyr9OJhv7q/sKnieoxFvZR
I6tLob96zzZGichGfjj8PwtOn49gstEjYgR5xjSER+6lLjFrRPI9hhp65uBeqCrT9OljS86aed4Q
Sq2kwgSbAYOJ6txnUUT3k6hes1auRNPDLFRO87/AP1PGbifp34JIdflAlLE37axsqMetC5s80H19
d7lUDa9pOcBSJ0MzecDdwZtEDX22rmu/wjIHzerOBLikEYO/xQN2Mrvpcc7UJUeF0S5k9VwkBFRt
+r+pZJ/ZUWILivhaP4lAao16JJoBsZlPFxSBDz4OjG0lkRezdxNXHLymESCOCqdn8i2ybw3TsC3G
4f4qsqlIqHLTH5pBFDTVgKOC11xwsWZ0a3EmCRxQqboNTpP2mjgAuiZ7hgcTRsWvrnLgerz8x8MN
Rsn68tNwenjR57ULWrOdB8VXJpd5On0LHXW9arQF4bRqyYPcGEdu0mSA0umVcoNTqyU08wSHLD2P
+IvxfcaJ9cqa75+YqE33BZK80bBXQJ81Ve2amn0vbFbmPsZY1zjpxsv/Mh+cRT7iRwUPD6x25c4T
0MbI68XCZPxgOrIVDe1LjDCWtsoVxvKMg0vco1nkrz0EtZLhCT1SP8jzxZtIqwgZ1UrGEk6N4t/J
HJ08e+cTxemBmakxZxoXdRLVDvzcgPqpi7HQtRFWerS9K3Z3n5lf+j5YmzzNG4vZstfm8SOfZYF9
HNdCTm7woVPFSa/3w+FwdybLpusBLRAxRgEw4b7z4DHTggMq9CnKy0SeTnThXvPl5HWhcE58zeoq
bO80qw0ov4awVlxttnsn2n1X69GSVj+/lMTNKFkKHJvZXmmDLjkcn1yPx8Bx0fhP1ch5chwAY2vv
ewUo4qNk9MywJlMI1GMyoI9pUmSRItOprQLbA1CLLOW0LsOWNLOlG00bKtoyVrWQcFCt7aGIVvCH
h7YVPHgsRv/+fvqoo30iRAM7sSrW+3xg3AeD1m21Y2Nrsb2f7CvDS/lZ11vIoieCfcNpJ/cZDgvb
0jpla2K1jn4tg8v52iMFUnqJDcR4otXhMxztNb8QvKtg3CU9VlNlUgQPw1661cT7ZRgfqLnYHLPa
COd72wplapNAdJHcQPHUPDvKzYHjV3JqaAaTHp4B/gRO3+sI3GVYG0ZYxblKxYqv/hXA5GryGapu
I354eX/AH15me+YYJKdlIld9hRuBDhnzyzD8y4RTn0wH+xIEyh9Y7RXHvq0wFHQWC71qTApLYrUg
EDUx3ntj5aAgfDiPtyZSTwXjs/D/ErDpfQgqqmDIAHbtTnqfTo/vs2slwhWUjdXdIpSTdC2GOBD3
5NGtwG01ywm6a8UAeIzaYY4lcoS0hqaUO2fsFmQiPQGDfza+vzLZNpdScr1JmYcIxFADIrZvvNqd
0dNenBCEHiUV10Qqq2D8T0EUZTX6cV9mLXyJV6gM37rfUhyCtGQrzQhd4+SlAbGtUB5Dlvy8YYFQ
y+EIa6qzdwuXm0Wx/kUp/eMU7ty4fr7464Gia36X1epWqDKQ3nz0at9IZ+Nc1F6Fdb1evOm+fyHD
JrQKIA1AvytP2nGELARvRnZAKOLZ6rhT7q7T+LXzmnXhuuBs1f/qLHmI9nll6lZ0EwQH6OlFOG0Q
GFE+a+tm4jVoReZmBsA9UqKjd+4Ymuie5IyuBfruDnJc4MsAqavVERdiMgpZhWnTMvUEC1FfcKNv
eqykqxOiSIU0F8sbkewFsE0knHPSPzc9CwahPSBSlo2sPutUGALL6i61C83Di/aG6sKOlBswVbFK
Ig7e4tEoEQVL4TL7s603GC24of+9muZrtXtK7klEbaep17L4xL75THIIb3WPzQDk2oTPDcq9SwsV
wZepu9OalNu2p5Zina4Y1CtgTFKUFviNTeuriRdsXtxGZNthBw4EE3kqvy27NL28x1dxIrR2q/gW
lYMvdZGhrExNjiSP4zz4TewBuTRoeE5cU63hgza4ciKQ8DRVdmK51wWFWALt2Nn+ntQ/tTvvNaWH
o05qtTUYo/7VViq5J6xcu96UX5/C1d3KOJYQR9ifMAC0u5p376+CQdzxrlN4Cly6FkHYqK8zIj6A
t+bvTj9lZpaPC/Z1EfVeBtHCoNwRjTdzooFC9vTXsY9eNar/Yiu81/+5YYRnayz77c2iSukbX5eR
dGTdZfmWrxOzP6nChMOIJSrYk7WCRMFeO2AC5n3hX5U63zvpALNGrIM2brugyeCtOTj5pi01aftZ
Wtn5fPu7KFru4tjiXHoBUBFR60G5f7YegNxmsP4nO81lGEjyNNLKZsj6OSivWUjqVEW/pWaB54uF
6onlrCmfW6xjIJ2VkJ4HABnMfKIHq6aT39CKlmJlupl3rW2gN8W2GDknopgwIM+9hrbuwzSnqmB4
2pRdjHTRonRi/cXw3N7omGfkB8PYhRtwr9x1um95T+Gvy9i22kJEy/SS2tXm9pziEDPiqiMwKwpI
tgsqF9ZKRKURb68OWmCs95B1CerSYwE+Mt+VxM49EfBBxPb844aswjhVawbuus26R7CzNU1UuKAs
k9RmeFmsS5HyTeTeU2kwb4fVRPlVVlwNHQEos4LkcHViM02pYPbl5PgDjhydL/AA0ybl9izHv+oJ
sctw8PNco0Fit3zDlX6rvbfDBL5OUm9OJwJuPhVckFxNXXMVvWm0B6knik5FQKH63M5YHaPfPkWp
8vf3sstKfDRtAU1iONFFJGuzEWSXidXaPPnPxTuo4J9KDVOwP3GGeE/obwOwL27+bVx8F6bAsdia
Voe/fbD1zoCIlsaD3KcXmGh4jPBOSJaOL9aXfRP2LVQEZh4UHaZJ8Mb3oGMdmxM126uoz/5xe8cY
A+lsWckDe7JWBkBvoOq3G2qX4+Cubh52F5eYXdpfuBaoFKaHGZ6MjQWzwv1Tduf96PVNsD1khQ4O
Jy6eURn+6GeU3IqiyyZvOExzxWBuIHWASPCZWgwCkbBtIoCv4uhszzLL1g9isI2AuToRXR2wkrP3
ObroPlu0IxDhO6vmVeA0ehPIpebpMOEPL8hijFMxDWXXTZqVQEIz+/AYpanRUV06S9jTrlUz7Dgf
kYuvtFmbBXCgoXnv+X8//zF4qDTzNn/CZdgKgNnVoJ2u9yTzENvMa2dOjo/cwybMAdgwTs/vw++v
AYsErvalZPdeZWMZhANV1Y9gslMDEbKSbuG7cPo3p/RmVCHDqqYk7mojdwjVzA8fCeIhzq/5GFI8
XZBIGDVdPYeTKpZN9/8UF9Q62ZJeZHPllmb05FrSFq/Hr2obGCSz0GXUsFp8bYfrYm/PFqONFTUB
vKLOZeMxGSF3AGvVVd3oSb8E8y4VQ4PRV5cMQWl0ijl5D9/tUqm+vVln0vkRE+QM0Oie9/GUC303
Ypv3KOHI829nR/38zP/270zh9Pb5GpRwpsZNmXCToiExP3EWTj3pZ3oEiAp3N+2fMzXFIP4+vose
wyXA34+/a4r0Q+1rV9+Zu50raZFE7rjgkkz7B9cKogOsfz+qqQCBduReqJbS/PsK2lJnn2RMeFMo
JeKezhlI75Mf6va66TF9GSEd9R5j2/2SZfCTjdyqf4pE87hDWkrc/wVGg3gL70zDPgY3CozIEr1L
t4dvroB2zOztuCn6NTo6UlS7Rtm0MFZ7Xg4VubQmhebYcu2Z02C1RuvQxd10k1OGITQQi7n9m395
GTF8DA2m6Hvvi8pTOujpeJIMKNZsM68inFa6eyBw4va5b0OJE++borW2wbe9tCfiohlXC4Cosbmt
gjAr9EvzABwOraWg9eWwsa3e1qClwXWfevi/tcmfbfL0wV7OBWF16VaaGijVha6s/mdIGPKHXMEF
2/diPhO8tmmnRUZ7ZUU7iL8FAvf9j/D+0uOLoSIPbuBDWhn+ApdvS2CD/nz6vm0Z5g6hset7/40c
F+OO5xSsDwBElQNsyrnRYJMfEviTxEtNzK6/CmwfXLVsfhToUxRHcaVIPgumgSV8s0YvAfTv6g69
mMIw/PeUP9bb1f4ifaWv7XF9GSDJxkMGDg/84Z6yoh4o4rO6PykC4NxJUI65YC7zz82DMTrmF+MD
ZwFSJ6Or1R12BZd75ktqpKTVziRtS+Z8C3f0UvpxZD4YmLY79ymyZelIBwhGtiN/7IoMyIgOEPfq
lpdaj7S3gFmN5WjmAjWAUEJYfiRgs0ndsdsjyIy6QsFTDJb0M/EFEjDFtZnYVSDIZDJsgQ8C0dL6
mqNZpQe5dcwH6tV4hoOMQ8a1xoGgHUiVo6rE1XY99sEA8HrFcjZdlqYx5kDl0g19FNcWc18YdKAz
ayFFcDFH67wyXE2U9fotpfiRUYnnF2bPJDIsOzlMN6+HVJALy7wA8wZbKEcu7A1buq38dBp3K8n2
ZbhkhLB1BT0gk4/3ck7QUVcRBnFpMdPR0tfDYWSLR/oQ5HxiPVZ9FI8lKTBIw+1lnqSSXHdQGGmX
C51gIWS46U+pmnGrllkXzMIxinwfOFsGtH3aluJ5uXEK5OYxE4sQX3nvZmBaSpXCLaFa6txF0lUL
5f0QT5Fq0fdao/gWLAZ6dxKoziwa5ebBgpiPgGJPHYoRpZhyQjNMZiA7IueWJUfTwf7v4GgoiF5B
Z10BQIiVfvk2dN+NDP3CIGaNgsUY1JuPo3dLuNI3QuPSsxULdtWlAMcYzUXGbagC9S4f41F99FWd
TPkX43MMRBgHW3Yi7fNVC/++dOKHvjvhu20vydnnAQEQQNWvjNxxz6si6M6NKEY7PrripLA3B7EK
6i0pFL0W0ykVSFlr/wyMCOl9YMi7sm+NZuK/zonvbK+hEoP8E+VVzlqdrW5nsUbDbtzY53MAqmaf
KGWVBhDjY7MdZcs7u9MgAAW5js4LNG4MKB+xLCzpd1rrj2oVnthuqIQt9zm7HMNoyd8elZOpaHWl
WkZhcjIqhyns4I6aqTZ1poWy1PHnYOzgAjYDTRB0NY+9ozdXFb/ki3mpVVk29sruKeeXW8JpTiJ0
lG/8ZvTgHinq4Wno1YU8B0Oo/RKT5OsQQgYgIPKLHR0xF/1EDcnLzEoTj9i57FQDU/rPCwMM81Ui
8jjlWd7lv/5QWhSpEY8qZ20+5Fsd79n7gtAdvP8hOptMkTq8LQg/Ix1HYzyA4fNd5vg8HA/XBTUM
HqrkwSHeaajIT25KSjclcKfHp3vDxgF49Gc7jtn69usyPZFenAhX0AR/XyMcuOxtDfM+ObtaqQae
yGBVh7dOHrbqiQulOShJoBi/uJulFi8ySG1GsD0F6tb13xjQTNLFj33CyO1IbiHBjZlpCBBP+0c1
2PdOqjwHYZao4TjyRXRDyRtWA7WbbIAAF+314uh02bLkXhccvrIJD8P2hV1sXLf7Jsv1pI5mEYVb
s9/JqYYmUe3A/zZrXZraoUpeOeatjm0QmdLTP2uCQ1EZ5d//O4p+l+yqOyxF+Gy0fQsZ/+/ce0fL
sfopNIXxgPyQAS/pr3ulpCczeEJdNO0dNF/toz6v23ijRRGLjhFG5uTuaTHhkmetg+B0qUHwmlVS
HURBiOa4kCsyIrIFPBHFvyFJHPMUR4/W1FsOw7tCgFaDZ2biDfuzTiZoGLqEBzfE81zIiK4cAz+p
lrpaVoTLIqtENxKHwW9ZjZK14JE8tKxZhDETW/3gtyi9oZd2aL7BZQa5c7/9oK7o706OR8AMCE6g
PtgDWDIfHwDTtg7lsiABcx3AjjvAy4RfA7E2a8dxJ0Fn+t/9QoAzakAXFZbo/0kxAvRDeXNQqCPF
EnsogTwOqAAGPIvWe86/IM7dOGYr40WVVoeJ6S5e/Em15KmsjF9AeDwkBZgd1lWv0/lA/E+tnu0x
VpPoo0p0knlcgdovm0TFSjwFVlvTeIqS8FoH7ymCNYFBeOvahqkSHInSRCQvwmtwCL3Co2sUdeJI
sF70z4/do1tvdfpW8OkxW22hbK5Whb3zveSvko4Cs93k+aSEniT6DhKweBNLJwAv/k7rVkg8Jxyi
6yvBWwpwGxJd6y0ggyQlqKevLInAzdmmaPT0htKKlWstlqw1S5JEEYD0PjPcX6SbB80VTvamCKKJ
Y21FPHkDOPzx1vdCV7Wi4JMwEfQUDfp/kdrWCD8pbX/b3oT6pTZguAM4hfXCwk5DfM6W6TFFidVz
fJ2Twi3mMAeuAg8Sr1P+WrVTbs+Y9ScDatCCztPZmTmlgcHCccm2LZnrVRiGQatngXOou/Zmj+D4
/vKCuL9waCxdPQZSEZ8koqRn/yUxdFwXNSORGOxOc2IKXRGsJ/wpYuMNJULRhMg6oVDeXA0S56Yi
PXrOkxQutILsI8Wt8Agb4EOvZpFD5IhZz6ojwVhTo+sMsXFghcIWoeJPPklhIE65vlkIdq43AwH7
hayJrEXO7Qm525XSQ9zMHjcz3RJtdwAxj+mtoklsntt/bI9otvvSHxISq0ULsKOtVkL10gZy9Lt3
fGx5H+1B/ajP+IIKelh1+rGCnTT01GExiHRJ+UDigAeuhSUMeViLjqkv5hEdhKvc2oftdo56E/q1
dOrVLF83zTV8bsEWm0QvXXavReskypWzI8iey39LM/k+mv3I0eGN0ZYnM6LMNImvB2ZhYMakTmQg
5HLWS6mKdkIZPQ73IZ//mhxJK19Xp98rtd+NKW0DoXXvwrbRd1fcsLRAhWJ3X/Xi45Bg5Htv+MVL
ozEdq3wgKOCIRNfpgYU5SXokPd0lG30R+TFcaMfcUlawe+yFzLG4V08m/s64F/ZDONLvyAm1IAkk
LI5pUaoPHy/6gtwoVFGIranUy2ZeO8mjuCOD3Znzm2MrSkvVgf4WWqT22TSTCvX1hfw/oYkpqjvX
jtJIrtmqovCWRI2rZP8zS336LMeMSKbs/WXT1/OHaBs6H0Nsy9nMMuTwOtn9jzlsF7ujlWi3zMGC
4E/9p3i+UKNrszqudHbTE4fOnJPsF6Vhg1WfCZoR6iHDSbg2ZbfrMeyriBV2j9d4qFhICeu42VnA
z7aNmKBs6gdbCLh0WyEJnI/2D83jyvaOXM81sDeDzKTexYYjwvhZ4947j/N+2E+qtm6ngwBebkL3
BK9lmVg9rlhjJhYBbcg7Y667J8wmGYwZiosvpLwTXhZdi77lXFoPsWYm5yZ4hR4LL1bJOB5rsHLO
UEqPk2lkmfkPyOziHgkDzv0rNTZBfq9aFjdX5K6iR8zizENDf4LiJbhIMhs8bBXK/5jhgwELXpkO
Pz9H4NnuoirRPKz6HizgF6x1a1hUIJ0U3JKHfeVYZ4RgNnEtK2dmL7A+iZRWOGRe1sB+navYPSqh
S8ADa3aWjENtO1xHy5Gx0u/xEqVlgJUnhWbxv7eP7JAd4IO2Agj9KlKNRx31B8VDHB9azD/LpFgY
6NbLeCU07hq7enKJNOBxBWLj5KZ+o8CtxB1db3c5g9k+yhW2baLAmtzAuTJLQLGviztGUu7S4CWJ
TxFi5l2pFqyAmsemW5ofj0aysRNuG5tm0njeGRA4Yf09A7Sv13wmxvVXZekL892A0zwLFZnxzt9s
FpWBBFBUSZtzclzb9Q9xps5h6Kgt77AkdLaBkD5Ql7+uZFUGyRHiR/XWKURXcE/yI+mrHlXlLAwc
5fXZy9kStwtL0GwBMlAEPiwWw7c8AuoS2OO3/OcpxGJA9mVn8pu1d1bfoFRYI5eYsOXdVe/72GNM
7KMBraMAEJX0hpNcLXO8CLFffFShIrMOhd0dHCWwUcydPkf1G5LwMDL2dGh3Yda0xeOUB0uPtF4Q
8IQbJizuy+jP2BAvcpwkrf42KGpoaXWCKDJ3vL1z966v3omymVdQAP7yTX7yxTZ/N9P1mLUZUR0i
xtKEcQh03o0oipjsohqiuMif48y6xK/Q9p9YK3kbJ2uQDkLKgOlbFjOWXtgzz8DDUjPjK+z8GDS7
L8M3KGF7jgtFZgpvlex/S5s3b1VvJ7GjqFOf/ZIjxGJd3c9KrZLjU1z6zQ7W2ayflRh+0JO167Uz
4Pxd3kssQBhYf8i4140+cVeeG7pe+TKW+aTstVvaAQsKgMZRKWmJtcCrhApDUzstnd2xj6wyFCqp
0AXt36Z3OO97jrzlEFsmrVx1M6MnjOL6ehyKTkcDFCsTJqUs2qIFoYLkBhWRCFIlKdgpOXAif4rL
9cy+pMjC+QxaAP4OWEPEsXObSP6GBKsBei4wafrKDMaTTjEB+G1TiTpoR56ZyJHDDEmc2+zLNn7N
PwOM/lAeHhOVmDRHMYdeIONdxmD7khFJYhUXSRsmTIuOp35mWOz4/KVHpCmg7Gzyr/vE4c8pY3lV
xW3BZB15A2CfjpHHj0bp+mUVUruFyfppJ8F9u/sv34vXzBnfQXbGRKbK5kSIpJtNLu9Wrb0zvpzZ
wcS0idpI1I7BbtnmHnamsrHSQvzZ++o1+6zhPHFQNKWKWqxuFaF1vEGG1bo025fNdwtsSjNjxNGY
Jr6Z7hEX08tEz+RH/3teYawVrm8FNiYdDyfF0YDszhmn03PEm8BPQLm74fTFhzZf+gRLDcmnqEkO
4iKxJu4ny8WsjnRpAQVVYtD11bvPqYkJSSqPkaN1/EhCOcpbM3qYge6rHZiR2F+3mDhPxCpIf9b3
/aoR/9pZp7zv6SML7y5rfFLpEFUgB+RUAA43QE9DoiJUve+7DmkkwdyYVLtkVSlJRQ7O6igqEZB3
Y+E1eurk3cYX7nW7i3vI9UZM40r6f2OeAFdPwk8IzAc+KsI+NlgtJNAekMRo8gebcAhEj47sCLzD
0xR2gUmg98C57TUcMBay/bQuwHGSWeElae3d8ta1QyRRgBHY6tQZO4SnkYj7f0kbaHF+RGwmZ9/p
soVQ8ZmLdvsqvFzurn+Wa+2H+jl3n2fXOWT6AL0YwS0fl7KdkEKBwjqCt7tMS5G+Zo4UaUZOkAOJ
Fo/zWfyb5zybAM4elR9Hg5ImB01450RBV5LlXr5KdcuuGAmAc0+cC/Hs18goawuDNnyaAWx4QUSk
WHNXYnRw77oxXYSlmK6l3DwpHgrmXENU0cBOEMiCSRhcgjjdue5HJuMZHSlD76rvodXmkxumIhnD
nUt7/Jyk+uDn6cWZzufDYLgE/fPPU5P4Htq3YMgGMeaye6pv+hab0B2OuJtg0PbsBQoAiGlthdw5
5I21K1nXrMQdHsGNVrYRs87HElCWTO9xVPrTv0RoGanuuWkPPNhoVoG8RMcw1HDiMkHoK3CePldL
9VquonrdQSIPdabKmLaYAJ8X1fsXALyOOKIF0wrI2eve6nsDeWIs+4O7ApLrYDO81kRXaTE3BdjD
cBOoLGTMjp9Jq2RS3S4ZPpX+sX1IldNmqr+Ntq7DdrpJmgMdV4ReNkyhJyPfh9+fFoVAL3LFpTzz
R3S1QaIdEAT5Mptv2yLNoglnFQXahmnTEJbrXxeY8YTPNrqWPpsU/7vN2r18Ua3JXGxTlPh6Kpsu
fAc7EfCcUG1N72ptbG7nNnEBnZlwjDYPUkEggaNbiEEWRr2GUF7atqZX9okg1YovxUvL7jY80uka
HUuRSNAQdDu55b5CbHc0/rV6a7dplrFp6J6t0gOlUu50H5xfxlAdTQYN87q5dakAu/lYAskG3eG3
Eu4OhAZlo4csqXhNqCoJ9hAwCQ9TbDviedOrZF0C4ANI1wjx3cWUgOUIOpD+YgIY7aaGjbcnvx8B
5qo/3qL5KDrB8px6gfLuXb+TQBRsoJDmeIX34vdrUOO13WY9SCQQlpHhP9ztSGcrC/uV0ysZpdu5
w7y6bjeUyeZMaVXDEeUSzNOLzmLTZCVcyWmcSxxdUiOH2o7cdp9J0Eq/+pKnwAQCnFeUzULiowmz
IJqNedOojFkJyPaRgpXH6oN1EVbXaw7OZ8wFr/S1zQStoqA9RCH5jlv15AdyvNH3i8GdWr7e1jO1
f+ssEcUnfRFdEySAZQI8TyZH3pXjXs8LM3to65Srdo3wMXSLtM1oUczH8JFdSuv5w44doKL2QbGg
ykdPDKZWF0reSpi3tI9dKJxp641dWPWt3WXYlsojr1ZvBu13froTvLSyutl5fOBfKu6104FSHv3W
hI19OP73r+Gbdrl2o02q09ZdTR9AqP0KQMjP6BCWeYpzC8A71ZfoaFah3V2mRcioYo90CzhyZ0bb
0HROpNzKNepqeH70CqVyxWdgzdET8J86TxIYE7ysJLcCy6lQ1LjglQLMdjYH9F4+IcYax3NwwvFc
5faDgOG5ETnCHUsaVZMAWe1offdZKJiaDe6JnTEbPTElstiS2r9pUiNCZTI5nKGGlT0lyvvyZEFq
5ltc6v83qFqp0UH9IyuKG9PKWqakR493zZMMUKWkPIq56bVxBkxqnm1uLfsaWVwvIvCrXwWITtS8
juZl/zSDy9FYzMXMowNlLMqwZ8OrWtBHPo9+2L52Y7ZL2kXfMkqxcuoUzGicjZ4rnevUFrw2Fxly
5k0xXPchuwF+gw5zrawwbk97X9a8/E4++KDRG+4Tc2H+d+XMiCGEONKuK8m6DVWFuFxzD21gVqSW
Q+HdhXWqRdyMeOvFYUO2EYrFQbFW4WAhRDDn8VziDgssgQjDYCHPqeFpFk9kzJjqXOv+NJ73V0y+
nr9ndor1ftWPW9Xc6DVr+qoEDSgohIisv/nuHXO4a62FyEf3PD4Sdbbt+3d5/lsgb7uHbVlHAWyI
btt3vHIeGpgqMAaLAdo228YLjng6WMI087v0YCKc0ebUsBIdS3m+/gOVmClasgVTVRPVE5GDf92Y
3VZDYJ/kbOHFZPlaglt2JetyxHNQB5yTazWwBd6R11n0/oU7kbvOj6BobkDBXJhqLCuKfG0zZaYw
utl7/MwFZRsR6m3tXKZyA1eT4bgM2qZTICewJ4ufKOOh+tYSj4K/kfV5XySygKz2ldu0/KPGx3U/
AKeVNcfag/y5ErODrpWMJQ1OqVSs9jHdy8z/D6YOyYqkfGUwEHzLq0RjsuMemh6ylpyST924850w
d03qB9UEeGpYZMBRUvaVy47BfsPVO11mE+3N7MBriPqdL5ezDL98UX93ZVcFJvAmePOH3m9C0C7q
Huzk7LVkvIDV1sUfHzhAyyqxBLAqRo5mwWGrqUm6snurf/yom358YP5cRCn2o0M8YaBTxszpfDH0
CYfWpHUfSi6m2pOs8lbwHOHSh5t9BSyFwiONvv17Qb9zDa5BIZw7MFLarQWVQGRL9V7ipJAEiaU1
pRGP0+S9HZNhPxW40Q5eRnXCSRy4D8zJSVH5PhUFPOU0feqwyslOBlUpzgGEgXznbMbtLmbeo3F6
8fBokIOAkG72cVtzZU7JME0z4XNE8ECJuA2IoBIQDX/YnNbHWoEb3c+NjZCpryB2ck0onO9BEfd1
UTWJL+GA2WQqyPZkIwJCZO4qGuBvXF+wvKVA61XPTu5ZfZhr7zict7x81njhijy4RZu0bgGkmYCi
on2/giFzNDtBe9CEf0NjNKquNFo2cAK+Z7QsvzGJJf8RuKF+9fAEObU2KJnnL/rkdZMRw6jteIwM
0MV8ICQIVApQmccIL/Ql67dPKh6hTZrSRPaFTb4ZlUJq5MEcyULwam0nQL/R1B8BItF58aB5nuHc
/dvyPP53AgvvoEotR3U5mVOIyTZmGgBrEP0BoVNXnRn1A3DoLALuhEqyNuchkfJbJPNvIM9mpaun
HRqtV/6QBe2xHh5cLeZVT62fIE2C3nwpU4pO/21nFHH7VyMBtZcogHkPRmebANVl7JaPkm7H6rla
g5NK2QwKEk4w4rq4R/ZA6vwDFYcgZ0K4BrIUkOrWeEI2c1qlS71LA7G5+G7T/bUMJmhxAeyqXhxu
qZiSv6ve9mDKBG4tenzn+3EkF7uIRBLxRGEH4VjUw1KLiJGMcSlkjO8Z8kE/4ZNlWP1Deh3VZiOc
z/Gb6urrnlQ9tm4sp7yK1ywHHjHLpJqOIq94Q+/a1zsK0sBLevARfMBnwi+va0sP58GKU/rcX8Ub
2JLf9e067SLGPy8RfuoWHKftE1I6Svh1aTcJWItn8x8pHNlfEjyO/QC7dsKMLof5HdVBrHvt0hp1
O5Bu7V1DleGYTzgUzayCfiBv8dKgMbrwIKfx6KF9idehagQpNYgRj+CoZarI8WNG60s9cb7BNn5T
2F/3zmZatCqN0o2/8NteUusNEODlrFGT13oEngZoHyn8olhlkfPCII1qo9sCWQX8IdguWrxB3ZIy
ogkZyC3SEyXt8UIJ9oPbkuMBSZIWksovN1LOx59GLi647PjpQg92Dcqt9rWAZW5zA6sAQ7hG1wMR
WySQZs5qUMaL8SYu9XjekklivKnwpl+i+2ya50V5sLplBbE43QrejXtL4ZNxA6UyQgJTAPZkg3Yn
9djJyQS+N0VcwI02uq453RA6+SM9MS0LsPcxSqAhjnmpoVrCMoW+bDpDe3tE8iw7w6LaN6Dv0iNx
p32PdmHCQdl3ojCi5ccxir1dLO3KWx/zyeaYKHBD0nWqIhKN9vfmXIZj+KCDUlYblbWCBocga4Cf
COXpG3UaV6eY1M1n4nDTHBG0GMap0kDsaWcrlpB9UpU+3uV6HGuArzVlJhXkmQ+6AUATfPb7g98k
yr2Pbm1/gTnbd1owLclXNi+Kg39qwuA84JwpSkKNnPByM68vi5q7M40Jm1+s9YHhwKIiS5XcVVrA
l196UfuqPU/GnNdKr4X0vyFZh3RCpNzzKiTkbGaTameTok8hN4gWDxWaER9Iwpd4m9yoqpx9e853
yt+JawPGcYwauU1zLDgQxF0RCcTlQmygyKRrzQ38TIQEI1rITBGAPiEyU02AnerztxJNSLvKIyd1
hK95m2N2vH+1WlWfKXYjlf/OAQ/7P8OxHj/whhQMZP6mJdrc+Sxvy+5+panQlaVfr3Dcndmlkp41
Gg0bAnk7wIHsj3mkMWLBxNrrKyQUTJiJnE8QN1p8R0C0FQWHoquzK/1ytqSCvtB360c/j4i+SKZ7
/CpFFhz6bfvHsqL7nB52sb3zodu120ycAGpFpK2LnbLq7otHt0rvKDE+d838tQhmHrgvkLXcj4te
gtQhw+2DLJ7LhLocs2I2pslJ5tetuAmb9MCfz8je4RkvV0H9hCaexzfZE1U8aQI0xdUnZ87ZhGTE
Yl2sjDithcJWoMPnSxeZiUJYCsT/gQkh+OebC6Fkigde+L8kAjB5LvFRZScxOFYBMVJywqtSO1uJ
Qrfk9P9CJOd/bWdY893JLA4QOBGnT4tLLc4uYAKa1WMjdgXwJYSQz7Y6mljJUtmlg8piDOaIgfz+
7ugf5uzfN985beUbxNEcA/jqwZU58sFsGiCRiDO6gGSUJ+fe0sF+cjQi6IhHQblU5FkCtUrN06v/
BuD18sM3Luu/DLBuhGu73f7NqoNeNsPZRNxJ9oghHChDwBHzriU0Lv6hMJvyHTtJ+hQaN8go/xGu
kSuA3Z2C6CiWEDNKbJHbgRTO6/z1j5R0BIimJTRA7QTxL6zXusUvexHwEh5QdMlTAXV5r4dSbtD2
ereg4GFJvWaxDUQYyW2ZZrYHymRgVJSb+a37w7jFsWpWEptHJOyE3Ts1gGMiUsrULMgErL1ySRJJ
A02m8TBc1jmDAfsQUYRs3QaqD7b6SC9RMCTzKEvBoiyQV7Syfr6/m+XFl2WcyT61JnIRgfrWq2F4
VjHCk4CHcWS+nXYP69LnhoPflH4DdHrthtEE9LerYaSO9XgKveVPtOo8LvoWW6VVxHC1IF/CXcJY
5YtwCa/Px6O3/AN23H20/hwT0dvNIvAgGgpOhEFZD78VhLo7VyfqeJQ6lxwR+Q9NNePB9j/uKR6S
di65fd3NI+UVSuGS4gNwPYsfPJQZNUVB0tn3fKbkORV0OPp5gIfqWSTsgshM0heBxCWUcsFsa1aM
JcoLNzHnyyFFJgWdAhYhp6Kgsa6FVHIoo2oq1UdoZ0ekb8C3C/RgkBZN+jQX60SxSIDrapE1lhCl
kyBQyVfrSG/rpfDskG1lGS0M17jfIRIe2pvzsppIUWzucrQ5xJBMu8IzQ2GYpL+8R7uwiPGfKHd7
NIatW4cd91y3J8Nu4iKv/vm2iXmI3VNBCZIKsFK++47AagVJFmpnldsVVGkMj/MoEG+qrcOpoZ5/
S/JRE5+foPqhz8iU6jRXvt9fUEI9dPdyedALR9JewV2mwtkGfnVT1T8/m8voy6pIyOWR+dlhDNXL
C5ZeiiJDFFq7vSLiru6RDN4MObyzMvSTNZ5jwK5iXbT0TkhggsvObIh45qwYH7vvZmHLhXDia270
zmFXAAOHnnWGxsj8RzBJCNANOm9IM7mcfGMPtsw9no6Iz+3h6Lfiz6NrUvSSKo2jXNRkAWZOGS4f
tqQJlEnIArUmz/hkVwt09qEaapFsnibtmHENE761a5NSa2as864482BN1+ZPe6zrv/srHrZAh00m
FAfnBvF2X4CO8chw9gZUeMzpMbaTvB9qOXL5QzfBnOOaPF1nZ/DU4nwLvVx2dR+SUToyLQW+0HMZ
zKq3TvM1jOkH1rNMvctmOz1T3x97BCnelHpAyrBb6e4iLeoRV2LIefYlWXJKtYBpPNhk7uWXAHo9
18HMCpsthFN1O75k0pll7Td4BRjMb/CAEUymkhLy6sHXSp0qi35olIvmR5EUVa3tt7mc42HTgDh5
tunsyBbL46iJDH5QeZCZVUkiiBcRIuOYbmEPSR5qK4YX6XF9SF6KLaSEI3nvzJMvfKriefOHMNtI
SRAMMmnU00gG4lkCofjZqs9c8pwKpLY+fcOIyvcgxxse0SI805Dn8bOWrnLIOaSLm9MZ8J4LS9Cx
joLDD9sSLSmjyB4AghiFX3z1zz8H8jJKtT9icGaC8/t1JLty7H6oIR0LFO0UAW7rOTuRNfth4uu7
hMsMuLHObYoHJWRyISlSZBQcc1XezUyCYtKrARy0YZ9ocoF30PocI5GDKYcDuGB07hE0et3jGQHE
mUm7/edBdBDJI9gJkAV7rQs+DnvWmZfhoyaOFprK0I9elUt66PhSCx8icE0hjH1if2iukERp8wHE
L8u6orCqLwlV2Dp0EDfiaD4VYHS6VX2c4pI7Kz0AexGmGeQi+jYAFPz/RoGaFxn1qJjl1UVP+6j7
A1EQND5GpOZTz9Hrif27nZ+7oSsJDJij96rW+Td009XSPhPYexe+aO693IStJ+KnoMhdDiY21Ejj
Mnm4X0gZpXwd6QhSSNKObbw4i7oLxu8yZM5CvSD3qfxmdhtO+xEK3O7CrxZzVvvKz7QLyirBA8Wf
5kpXzMySYa1iQONgS4wchBGBB+68uJO+ZXkwvmJ+1J3CytqVSr7oU8CfPQ2S/Q5xcWHg6GE0e+qS
2vfzWqCiHOASDgckw7WyX660Yd/l+77Ze3La4maagsMAu92i+PIjhvMBdh842wlsisTLh2rU2TR4
zLJNQntJVMkFuxvfAIZm1Cxee7+bOQZdTTba7TbiMwO1QUZA4WEKJb0pThBjApvjtHX0WkbkHmlC
3lQO/I3OU1QxVfsYUBH3kMvELBjJuVs7rFXYrQezIv8N/pcaDwDE8dWaxMGGQBDXyCcI7aCeI5gf
Hpj2SBN3FOlsofm1fZU5h0t3pfd5HlmzHdogCpdULcSl0tspZGYs+YqBOUFNxuROQMPpTFBuAkhQ
98kr8zgTKc9Q4nl2P7Be+0We/A7d9+RPET0abxX+xlV1e2WPKlXmic4QHmYXgHBtybBfLcA9gfep
3BaBT7V9oY7jU9X5SIT8oLGY3p+wSAUW2GjFp4RgcnJ5/JYvuACThgQstJK0hol9rb7HcDPd/t2P
4bwORm8swF5nKNE6O5uZ403/OKjY3ZWJrrT+b04IvnS5yzH6PfWSwsHQdO+3/dkYIaHL30y8a2ZN
H98xi2ZGJIxMVKUVKECGNnkJNIacnyBsN3d1x1yowN6P7SF1JsQBYFatVGlauZioAt27aH3e0kmY
ykTcLxEO/Y5D48CNOPMYPy+EJDFl/H1xzTcazkjzmZOm8v7tlY0IE+yF+jmH02t9fJAetm/fi2+V
AKuGDBECRr+8FiTHyQ8CcHj/3Y5r0Uz5K0J6tFu+LxmI/GKnh4tsQhHb1y+r+Zt4LHR5CzaFIw2c
xPX9cTP9eiBYgup5Go5HAIvDwsSyZfDvsu5VlUt5jJk29g4YDudEX6A9Lfn5ok2rQBZQesHXC5vp
otB3iPoCf7O/zEhOrb9JdHn03RhWypkS/21lfgceX+XBQP2xOl3Xji6JXyxcPeNkXV/raOvJ8PH7
ium2CXmw0qvlXKFLe+jbCUe1p6KzqRZ9AxjkC10uKXJHpBvLHEBpTTHQFpC1Gu9id8e2QG6J8kGh
ulsvwO7DGqmu9JcuezFhZlPpYPRI2K3UBB7Vr4Ce5iDkIaB2xBEXgFcHtfeMoAYot15x75PrDqHK
nNH5hbzesD48c7uFStnsp0Btw1lzcIitxBANUpXuz9hOT6iyKRuQLnYbuYi0BBbslpqVPuJHtO+C
bpg9ezveoES05wdt3VRaAP2jXaqIpbOGvPW0KvF0O35wcJjxs0vRU2Mstl3IgCb0ENrutL5yFV8n
EELpVT6ej+elZSX7qUN4Vo2c1gUkwm6BDz+AVVbYyfBYHOTNp0mrUjhPzaLpvxZoLfKMah7Zkn7y
4LYVTftOY5iHafciamMkGA4rJ+M8gGsTKMjrvq47J5JXkxfGZR4ugCjwm+o48r67kTZlkhreljz4
1rwrSE25a9ZpnjQ3PDhFs0zqtQnPJ7i/tEe+PquubQ8B9gAZXv60S5cYBtEZ80EFUhGBs9yVH43T
eoFQLDLLXu+dx8QKXLwiRyPkjR16GS0+sF9gY2PpkT1Yi2pUdNBPH8i08n96/gj+NAunQDwUwVs3
Xi4SwQcgemgAiRVJKU+7UI5UzUuZbScWGXpUWFCOTXCb//iuAJ8adxYyYwtYQcIbypcWrmVgV6/j
naQW28urn0O6E6hLQtrvh/rQtyF1HwyVzUDIhU/ybWnHtlKbIS3ThynbJeXQEinCjTAMhURdl1PA
R1WtSk1X5f0gu57cAKNP1xQy+kzfP0X+6Ftx/C7tIuUqYO7+gSb/OCZVRkBaxZY0PuE1M2Js25G/
MmhnU6hu5a+0mfo/Vkxcwxjk1M1DEakisX7YuDjiSTj/YNBJE8iozM1zCMNYajrnUYGLV+Vs1xBz
UKM8VfOfZnb/GidFfrJFAPqDHdHWU8Ctxi8JHfv07kZq1jtSHFi9zBE+FDpHadSlnjyK8jj1eWiq
axwHr4Q801lxl3Zf5NRubLzPSzjeyjYOhD+U2eFvLJiXa4bHNAHefW7PXJqL147etvS6WNjCkn9+
MlJ7ckhvMoWwJ61xSCnjSuto1HdGdd5wzC604/QfkLZrbyGr/FONAhGcqLaLwVx/YBzjQMCZT2/t
Dw2T30HHHTuFZUyQP5sohHi0GCjLGlpm487Sy0+sxxCJ/QKk9vu8sLBYWRSz2BNkI5vU+7L3yzTN
Hj3Boa5lbICZxH0SU5aqd2/ZeIpxyY60uA71wJ5QaKXuPN29bAYdh8+TYGuKgNkChlhbcqFQ9cO+
Ex3hTC9SBkxpcAfBdMpDrxHP1OW3Zv0eE7LY4XEqn0FShipooY37Wi/i5msKcDwe1qVw8oemBttX
FPxBP0oLzQg9Zg+2+in7EHZEZf0+ojYJb+V6SczdNFhuGThcW/frFym8FC53T9VZD5y8zG5uwvYL
BIYI64ULIjGMsLxTLeriX/R8KRfJG1JUB+T3nZeYQfS4wda2SgVkuue2AHP7INl1TS4PIpLPLE1j
7xcYLJlTaD5KITNcPGYaLBn98t6yR1Q5/gOf7x8WJcxqNO5gaEEbv0NusqyPTA+MU6SilQsXNrsT
w6u3nAL0rW2mBX7Po9LDxbp4ODwZl8MqWDi/c4DbcvCD0QfLq/km13JBTLgDUSTSQfrz/YkaI/Wy
kETb+ipynWGf5rkLshnK/SpudJko2xq/5/rzHKOf7wb88HIodjbDQNyHw1KCYU/Wzzz8PNr4KPx8
3Rt2M3pE2/2OZh039W/o6FTy7o4viYC1wH/viN8Afw019Xp1DbVM1DrajwhQps/1tmemfUTXF62j
l1eV+HebGUPtBsDcDSPL8d7XfWUJhUGWEn5lbf6yNM6KGq6SpZuiSBhM5lwyMZSQQmJCiR8bKBON
mlnNFpGiJMnNswxWg7+/mOvlZbcUlTVTMBoqhCvIFJ0L8ToYP0iiH5J9Eqa/8zP22rLSLrik7iR+
TwVlq6LnPVMoalCFTIoZ4Ud8ERi6VfIm2LqXxzv3J7yyJC6KtTRo+3QWWOJA5hahNhQM4UnlTXKu
xRy1z3cqVu8nGqqaWwrNrBkwK6jahrY7w9H3rX3jRXhh8mQTvgQAVnC1oxgZFCbVzGYKQ0yP+ggs
apYeUz6XjFMMTHPJ6/Q8mSgzaGgjcZTjWbkG32whVsVhQgjHpN6y5UoHLPUW9+FlSM3s0FBXjZ8V
/2GWOtPYij62sD3z2GME5VkclLTgjyNzbKYMcs45XSW9XUnUy6/AHiFOejLM9p5ZUrNP8D+ZNyvl
cf+cLfr6be062x5UzLSQeZcIZFT9IIT+viYd9YyZ+aTi8zf6giuxF2nLVr42yAr7aEROlt5RKdmh
6gOxYyIZIRuIJ7CGIry3J+1GR47Eqve299NBRyEGXyYLAFvkr+YkKiNTaWxqw9HERt8/0fsD/3+R
9iTpXSlsDWLfLu4tWJoS7+Z2NMfoEQbimGwFctiT871Tl6tb4caMiNGA6AA5zS8Dw6F5NLPp/H0X
lq3Q9oVZ7Hz6B+gabpVEfsCAl/MrjSUKLz2crmGkndBjDmv1Qo8nl4qlixQXWOYr85gS/+xa0rwk
nV7GChcm5mDWLA9ZuYPBRkstT+0ruSl48FBiuT6WzoFdjv49JGyXRbjvYaYPKniWpMZJY2McixUg
/2DO/4NuF7kyOc/POQfrbxCLa7E/GrvE2UiTiWAQrrotGOwl26eeQejGL3vNf+kW3rikMuvV/tWE
c2GycplneBMRGhsngbkZqTcklzgtOr5DUMhNNIPOIDkqt2eZ0PZx0rdQ+akGqSld+m+RqPLAfSRq
3Wlfhe7+RkQ8NZOTc4DDL5jbEXLjlN1opcUAQYfkZu1qR3P9Z2w1jBKW7zzBwGsyNy6McxngmjVl
IZEqbnfQwDA6XPTKbp1APt4jVt0HKLj06zhrIpl01U9Q5rwXYhmnwagLO1o9MnksHs2AQjAkkzqa
nqYjJw4yX8K77hfkMMyTtsb1niA1tuyZpUTTgroI4GxpwPUXPuLj+ed3fV/wy71q5BPUyHHOIR1l
KzmHP2jxDWV5n5DSzmFKwY84j//bKY8Gn04EWD8VuCv4a3bvLrCgfrrCNlfrrxFCNVs6LM4mBB6O
GnXC8nxg/MjhGZzb1fSZJxOkqk5ZSWu6nTbbk+fJN/PZCA0qGQkHhou8H2GBhaCr7R0KGJ0CUtYP
X8dzX2EI3WYVaxxGtMBSe5Wva/ZNAHntYM7HWurcgZqDYPHKf/G5KQ5MVV/0jRUNpAboAlJ3KFMh
zO+bOGWIrBFi+RrllCFz1Kst0FDvTCEihvR1ldj5qpS8/tey9yaOC+8OgHBmRGsQlF6e0rYxDN/Z
r9R27w3lrtwGeYdPmQNVCgl9alPGSlJsMmO05QJLZ98t44ZrLct/JAXih97izJ9tLwVeZxxHOwGk
sZTQVtyMttwSRvkhgOKvH9eLnCfVdWDZS7e1almX4AgrcHY0QIoasXJKdZC8ST0RnxzsPIcgP0zj
6MwKTmpTH5qjmVb0Rv1VaxW/XmX7R099HbPaoWZMWsnHNxzbNI+1cipj+1swl9MF1KO0VaW7nVG6
EcQch7T4Ej8jX6opQkKLPFgSxIQWqIHCq9dau+vTMPHeFXzOqCW9gKou2Q2ihJ83UqFl9tTIT/kh
kug0CUnKz6fhuh0Q5VI4+25Re7IgzHYb2kqIk4JTxmrOZrP+kIuJQsXLldWOoAfd1YPyQqTamhKJ
lLNqw+BA8jY2u5ZKMVZu56Lk7RLKPTuHsCf2O9z2qPRkafRGylewusEphSlv8UjsTFmAjqTajk8b
VusE7GvJ27SXNY8SZiVXcLhVT4yoi5tAgkLaEmIXrkrAgoy5/+cOYie5Xb59NAfiupa/9i0ZL1ED
M9O1EM+NEppvIi0eyRnsbcLJeufkkBxI949Vsdg5e/LfiP9wzmIDEzrl8nigIhcWfmYYiH9u24WO
554X2EFNWrIt0CWOL2iCMxF76SSiPzYR1QZ9HmKxLm3eKafrJ6Gckls0kVrrxbjdNDs94LxhOFSi
S9yQehzv/XTz6HHdqlXs2Nro6xMVGARglmIUm9vwWVPY2Rp6zc9U8KnR97Bps1uO6FpUr2wK/942
H4QFyi9DRHMw0jQ4Q8vYAfExtgOCSrGpgWm/pzB7wz2SfPVVdK2XjOa8gL/sulVyeujrctybOcWj
MTp1/iOvxKpVdkIKS56nVSXdCjTStE67qY+O+gY5/bsmm9bPavEMPLdvSDuFgp9/VQMc+iPUeP/a
NWGSL15SEiZuORQudJB/AH5AXF6waFa8ax64Vf6hPx/JaO2EHN65OELsCBf0+zv4K/XWHtKPe5LB
jqkCd5V0az69r0w/B+rGqWm0musNHlHqjBWEfveZ9Y346I8HPixm0UOaTMcbqA4SflJ7xifc9i93
gmvGVssGpJgTF+b6ED2xSdT79KXhjdf1nVHgV3N7ksknrNi7BxW6ghOjV5VK8LAPS/5drY6JeFMZ
q6VencUJ6Bq7VrAm6iDu2auPd8oSUtMApOeMpWWMJ3VBjKSp8ZEWPCNI7oFFlHgOmj2yG/UVO2Fz
bHWPN3mITq66+SxxsPKTxM4iMOueMq2BUXLqlVPC9BBkZhHvywWOTLwvXFdwyOeH6PCT/gaTkCQi
bEv/20i4QJgo2mrCKO9KQ5tkodPNLC68Snwe67eBDWUg6LF62UkY9PVV6MfUoH0wIhAinWzsgDhT
c8L0wvAeySFP463mqssaUK79QiuhzAEwTTO2d9DHOYARNDoS56YCa4PFMVBpIvGc9yBSX+mYNLOs
Wg4bRpzitaTnLnf846oe4E0NHl1xCt4WcLdWaQe5SP1emKa5TuaCvZUBhCPcQLilcTfiobPEo+s3
9uwaKs4KZ2rsZle3LfI/VCxmNyVZZaRy/tNFHNm7IsNUZnVkZeu7xeyRKPkt0jd9bmjfijh9rIEW
mLyB7ZvBpqlhPvMZqqTe2m8pI41a+uf6t4/BraulQ5e7KuIerVNTYA8WkNrjgH6AEuvQV4mCqFGh
fxNQXe0QVRiqUm7FK4+HVEGgFqeGtMiANekG+xxoS2g1BGuotPn2Rca5dMHFMhkGjs1Qmdt8zpyK
H5YotX7mjR9dotD0wDMS/y8d9LGGnNa6L+LGwPVFTS4lptw/Ba+hu6e3FR2ljI8DqQSPhZCwcr0M
EOe5oi+EkkApivwFGPJgSCfevgi9aKEiAng+ZyrYNXIz2PJiC/CHxwk8U0nGGn/IfqdPjvbR+NiX
hY5cq0kVLSP4UjKYl7U1gdTg+aSl/TivnNY6A5+p1F2KNqrCpbs/x/fcB3k1IhO+qBkMrVTR3xR5
iOp9z1VgQiZjHadtpOWXVoPda8+WwSuC1rA01DCFjYqG0DMe47EPh46/SJQHKHQgNaIcI29Q7LDy
PjKEvRzWAmXlc7JJTTHSRFoV2I3hmeGaKz+4ZitgDqvNh0QIgN//SFWyQq+dYvpsnJki/zPoUOuy
REWZqIUq7bH184K025ZqpPNShKWqbibbfphywCGfYztFqPF6EI9qIwFXN5ySmNIQI6Fzi38mjyiy
6rrO4wuwYCnbNON0/rW/dgvpzwCEmYegKiPBaJLb+6GjTrns7e6L+rh8Cqj/X+BDo7QcDYjxij7H
w0FNaFa6t11Fjkx70IJwxYbD+9FweGQaNYT7defxZQSXAJgQfc1NxEBjxUl+5CT65TRwoArLFwtc
HoaCkaQcvl7SdgMFteWCRK0ha4i6VznBNY45gyl+Hc+0+MgxLzAl19cEbu/pQuBJJeu0wSDE2iNW
FHknJJZxpchNFMNN4LYpbv/CIAIXln5SJTmqvqPv15bw+38dA8bl/mvdUNcJWOnZsvbhdfCO5Ihl
ioyQxQmtnnBofXzYPthR83h3Vdn9p+W8lzgSVaeazhI/EQ+KGX7X+klZiKK3+cQ+chy/9BMMBO5E
7lIPgzIoeHIAV577dvRg8mivFClgcdnQIdi1ZgDEUiP33vXXhkYGuPHgJuAuX1pLzqnCWkgOW0bI
lUAZnDpwT1dQY75OZh79EPvfaDYh+Tk6euTJqQw07py98SSk6kgak//gaJn0zMn/Z9wkuPAOZCuc
wxc8sqVheFGJJhEcp/cSVuth9+DyxAqOE/AnlT5D/E2nPgrRP03MYRVLAtdN34G4Q4U+W8XkVhHN
b8znwdhD9WItUoW4w+HFryRl0RueStMN0LK2P7WWlM8iRkHQ5OEDMj+6qkZMd/bGypcWdkp7FIcH
vNWsyxCj3XorkJt/qecPaiahi6DEHkC0Bb2tueOG+kpXEajSU/2ZY+KICxxBDqEj3e8CtyED73U9
1xFWkqVpvYa4yWMML1cSdB/1alVLtpMXtU67kgjO6EV0aSLwivEywpnMYZRf3JrA5/uupb0s6i9K
syOnsdAe7ESEK95z8Oko2ydpq3eNQjhmsNWR3jS2E5UXVecQnlhMNOjht4sxMXj+UaaTX9NwC9sw
zp+QQVmniRaLf6rYzxt1rqQY68LbcRvORlsDZ3oy8rh1f+iSeYJs3hfLQRQOLYbFfOWJy8j2A88h
kwYzbD9WEhuGjP5icuJFPzWKN2qMz8F1iGxDing8SlMkSrwN6cTyJmlY37s5/h33+5f7PoCsdzWh
Kcja2h2VEVKGt4tZ6PO+Yvs5fri1EqtBQZA2vOjnmpS0ffioxIRZoXNm9Jgjc3AoCROf9jvmElqC
FDZmtJMLlRU1qVhtzVv5GCWF7B8b36/XlaFusjCch/Yk+GYjfvl2b8Gnx/JwGiSrePU3MGcPoC1P
xQrmRSUjOdoC7JVxVJ150FdMTo9FMlxemY7TJclyOff2FIDNnk5QTAZtpDgkAeGZefdPtMYYkKX7
mN3sGquIX7JMryO/rRenvjZoXLEq4MdsaMAH3jV+bpPPhwrgpNeat06yhZjR+T/OlW3yco3HjXKO
x9fPaXr4vl3VyuqaBmzGEmtTQajZyntx6zwX5WrrC+j7zwTm59y8YFXFowd7Tobmmo3gn4OZN6j6
gCjJwcVELug19yBgySKR8PvoGJdaMATQDAn/3pvv4Q9gm3mih9tO+WirEsosc0vVGSSYwQe4vjhX
8jA5/5OhV2tHSa2icbS2mgYjNiruDZgUKjPTl1awLF99MbkblWmvJF4Cx1WbUdMqcr2iUxQq9Y+l
pSC9hpayraAer1Qt75HbPCypCCTSYkjDXRgyH7f0HN0mZZHr+bMA9T4S6bae8ohXIlP525KumzjS
nYXTb0lPU0BSp4RrhcWnn6uVoPOlTVRpXCusEE84FYO853DOlbhBj3cDP8jibDil/JDZ+dCyp/DW
uE4X4Sgtz/rDOP1XGy69E7BHMrWu174oIAe7LJbfQo42cq3YTokF5sRwbUapZpekRRo1X7ODRxbJ
H84p0SyEK8OcjRyZguFG839uyna7MwWxx/T61biz8bFwgYIVA081r1LA9uq3HTZq3GfVRAUzLDJb
AxZzX7NQnC1hAc13RW7EOqX0L92DItzgkxEsBj5qqIPVFjWciBawd0uKUDYLKjE/R20gI5VzvHCQ
/oTcY2PI8mDqZn0GuAyVWmxhZRZvYes3vYvnvUMCTyXj49ZN/KiTB9wivJo8Eecw39ACotDTtFv2
NC2qnKHbXtR5dsbu5Ujq/YshCMAnuiDMWTX9sVT5NkZVGC2ldYr6j04AQOXv7VvVyrwvNZDA/58z
PZkF3m2la8bEYCgYtDdi6t5NDeDyWJTLxY2frd76C8c8I1V+mxEQhN1QoFMCBv60ZpwrnqjXROVh
EXt3o1rKi3oIwqe9FtQsmxw48Rh/JowcHXqEZcXkkh4lz4oPjSEnM87TRTtQBq8JAGL6vcUw+9I7
ZoHdSxrCUF8lERaYvhdmg6GljCgSGPIPk1ju4ZYv97DWhkS89rUD6o0Tv7Aosgn9LKqlbDKgxvpg
d/l20HZDp/Yl+CPQTmrOsqkdmYvfUrVvjKrAuS5/V32GpiST2wythH8vzE4RZvIv2y9vDpl0/Ggg
L/ncp6e4L6EHXxmkKmUFWsKvcrY1Dg2qInIkI/vn1m96IEFGxBj8hhGHSv1RgmXwQUvkaTh633Cc
y8iA0bUYL4HkmJQQLcGeasBCPSbWOJF8GpFvZVVE8jKW1jUOPtw89XfsmJH5Xk+k8qLJzgaHeSBz
G0ZxdS16RgkkxulO9kWZIzOmdXQnQwF2iZ0P7AIFQJ4Ftn25ePsLPQUpbsyzN7bEIS4Gm2TMdQqg
QWIZfqsRdzodNT9SfUPKVt/+bsXtEpUW8TTlNFpLtH3Ok4gXstDSned8DCM1VxwBxYJLSGRL2nDt
4t6gZZO3UtvuNaFkDYz3L7Hbpi8k/bAc0mpQ6zbAVC9Ip+w2OcvRaEYkYMw3w1w8AJNMPwIUhT4F
+ALDTINPdV1NVt1DFJT48P4nU/b5hXg1qPhLUBjDfMKZg10+NNq8TwgV/zk8phoFH9LhYbP/NWzi
VeErA/K01b0/Q5IYhM3Dw0IBEPqN2KEaU39Xmz3bfifXXvn4O8qP16mSRMEmyCfjxWc90S4y8vpE
UcEB7J08J4kOEErM5vY6/FAEX0wWPQSXGs6Ji8VoHXMQoBXjKcewB7rhfSflktvevFJ9RM8aBCn3
e7SOvcr2U7QnpymIezGobMQKlWTt1YDV1JOWnxRF5jKbufVUT1+4W0vSIUjhn0sTGU43YycUprfk
dJU94+C+/xKTsX1DzqdEnh7kzpL4/xIQ58JdExLiS9v4C0w+mO9DBiK9ab+whOhtOs7dFCbnPXun
1o6uMVxW2B3OoEgr4JnGnd2RTQGeplspHFhnRID2pU/iuWIcwJ9XS6+hfgPTDZB8E7Xb4bOPi6VY
EOVw76u7jxq/IkMeFmo7MGTA2E1e01IU4fip17T+rSPk74K9ZiASBJMVb0eMePQyz5ZqJOjxONTc
Ix77Y5nwgtut54eYc2A6kfJtNvFCCZbuxyEGSUulK5aBDEDGcuHm1lJjzxKHmNhJ3wcoaaC9G/o1
XzUDWAasnQfo8+jiUofJ6F+aCdOBUrDa7f8QV7WMfEBizAVdkSn+c5ZnYNSjcQknU/aYNC8jFvjg
v6YSo2umey6V78tpayqPYX9Rx8eX4mCck0YwhhFivKeY3MDFcKxgNGjBAteYIFT1jxv4KX9SLGeM
2oyE3vMr7bAY3tCCWX1BHsJcwwFhARugbYGAtoWBlAv081T9P7GEKJ+hO319w0C+WpTHf/XPVzFj
I6lvaXPC1sH89hq4DH+d6VfFqL7qQIvs2+5nKXU59c1bqyHY7SyZ/mvXLCiGp2+Zhd1gnaa7wkJ7
Ndg9fns0CZbvCBoFXVh4XpN4KpNGArkwEpkmH+JOIY7WnHncbmZBbLb5FhSTfVjffR7PHvwxKs54
X2qbjidxVr7OMIFgmk+jFNcIRV8PmyFrJR8Fckpn2zexnwJxqPX/gjkisBtxAlz0jPX5iZJDQXY6
9n2Y/StS95XhX6s1f2to542MnJTYdiFqV1N+O88yf5yiuGYkAVs5yrbFJ/HmbhJtAWiDbvP8A5us
T7duop4qtOzAVzplYBZKFuY6iwbKka1eKtS7oZ1jxS3OhCfVfcMeaKC7sJTahvR6pdWldgDfEOha
UK7fz4Z7vfRdPf40/Ti1YurGDS61swBjDPFUt9dV3dsF2z/BUvAfKlIqEmipQqKdmjlhRcvZTzP0
5FVEOVB7Xx0ly87Mv5B7h8v2oHlh4jo5GFwPykrHhXbQA5ZuAVuDz3/yXRGNlv/Qm5UJqrEd57ag
aZ17dVvFeYyqf6gop/QdLWyoRw+UXqluggf2NVjXJTQxyElTq13qe0MW3EPC51h31m5nmOyY8MlJ
fVNiTTVuZGkAJyEMkl4tzJVdJ55ypsnNWeWNgl8go/5cLjbJj9ZiZNDb38H22u4T1Jr7BmQF+zGN
XnRdIlgJZ0e8r4gIm8gVooU2BQAfZDKDJNlNmwifu55h43ov4hwPHtkGjhuxVuLdLKIauQiBTq5s
ypnUUq+sSSDCx6+eu0Di3x+g10vAFQgMiwJnqCsKysXSL0sTcI4HDL+fl3SRiWVS4aSwzcsLs+Fi
fLki54CbHEsAYABhcAq1aB3U9oKnxpTM8kpIuaa1YB+rquEjVvOG9Go8PFzu2ycP69hbBwmXqlOf
O1X7DiCOnho0Z7qTnW6gTI5y98Rzynxu517qzIXkIzqLdK/imnzsi0nCzTv58yhCl/WsuDDxZSL7
HFgzxJ+PZGN0a+7tcBqMRMQrPIvHliA8sv0f5BeoJyUzO7ajeYVff4blVEkt7Gbv49AP2Cv4yTlR
hxR8N51co/LGvkndj7gTNhRHWhg9i8h6uQFzhCqITAOA1nbFEOFNE4tCzudcQmjMIHUOvcWzIKIA
8ChXzNje8Oqe87jtjywi7izvGx7Qgnfn6MVmWUolwcasccM7YcAM3lEXMa4pUIvIh8/mRF2+Kq8c
1RiTx3k1EI4A0Ys/rg+LwxL58zWOHjC3oOqpi90S/2+Uqoxyag8l4hA0V2SgFO7wlNk48fvRQsHf
+Qta6dhfZICX1f3aqCo41YyEoK5EzD025YNp0fJX796/5bWFUH37Qy76PgaaKYQ8/bh11olw7cR+
4GmouDJco2C/VZJ1Jz9avhbxZJzPRBIqN8CGhs+xI4ur5zHLDN0JuwGiS+ceDE9juvBmquPj53wJ
I9MB7eWc5Q4BjztmnNoscA9MLdO1Myl8PaydhDqF50JAsxhvalRolSInE+oF8JvRKiIKQNXIznGy
BzLKTnvFJC4sw42aVDCSaxNU4LjCzYiDqn40b+G4aoauSLlx1IVJ6HniKBBjjwvLBMHAfsO783JG
lRQcjJg7A77haRi6ydxa7H4b7GsCMf4sZYzTpUvqK5M8+fnJz3Lh21sceBoOAg+ou7WzblEIsWz+
si2jGz8HFOtBAeAvuem7btzzLzHi3XF343AucxyGhqmxFUHMN0qfiqxCTkyZrYDVaFTty5q0TnLH
RcwZHSziC2c+1ncr5eAR7cE0O1A0WZ6/po227DD5kc9Gv+jYyToxyJizlXIAyyme/xiqUhn1zSiR
fl8CI7ss2oz20LEQWJVXfNTzkXBV4R226vF+D4po+31ILBBjra7iDaluMj1j4Z9BSIermoCnuMGh
bM4Y9B2yGjJNn7IJQ/mRxFi9C4+YdEGBTuAuBoUSQdKyG+L2W4OQ1ue5pClir9XlWJOuyJ1uxqD1
dFlcVglF08jn3cwWcT1Yc8OG3Yk5Dd68vC4mW+0Ij8sjfoR4DO8leZ0j6ZEx7aBC10afldUWuAGO
9MxAuA+6khKLGwapZ6TJ3Jfg9gtXfghO/LJON9/HQM+0TyKsrSX7jxtdsZI8JCWQb1NZ/v1NXkEx
j7t7vTqesFnO/oySd41y7zzIG+QAGPK8TCInR+uJhddQmmAJvKHrOr1T0rKNiljvQrPkLHmrH0vP
wkqvOUB9xfid4+hyao3pQSP5cXe+nXoV4e+9HAd2UMpStAokbYn2ikBZr4B9q7jyBjVJmrxH0coA
2GSvOWuBFY4Z9hUB0LSMkTnPkzTtAQBYirQ/yLiD9Vb7vbdQqbzbxS1FN14FlBY73/MA2V7xQsl6
Tk54jhtkFuuj6TotvMvdaYt3v8EWgLWOAkcziUCY9aCYBynD/sdLbAseTysPtEiUdAZQ2qw8Ric6
3jeOzoBgFH1gL1/X0M5vj4cyst1b6TQnLzH0MhDvzm9UHVzL3f3YzJ4o1afrHsJ+Z3gADsKsCsF5
8oFJCjT0/WcmbXQEiKGQ6GIadKnYdKZnilhGiDcKX7ihUIFarn2XdbW/MBW4QXSaP6dyfdFsOmd9
UFEpgSt1yb7GsdqoSX8KSG/I3Y+Z9zfKdi9NWe3lion0GW+guF1cGQ6LFnIS5IMRulk5bInWPauJ
WwFtcNycDvIdxplyYF2aJ5YY3vgl8DSS8p08NT/2s+YFervuHiqHDm4ZcTucu41pht1yRWG6Qz2/
EMxF6d7Uzf8Vm4KJ4XmVONfLhJs7asiFd8tmp113P4eNwm2SyB887bnxiKhu8LZsxrMlbZJ2BqZY
Y3fkmypEFOnECBOaQ6rLujWVmZukLHXhdYN7m5vP2zB1EpjrDoyS6wzklqM2CNIhzOsEgAO61eyV
21FUgngso3BNo+knpqHqBRjtnF6q3MsIaLI4afQIB58CvJO5/mk1jqj3TeH3QrezcRlDW0koT9Jy
cGkTN2s127ZU39Tpk/sZ+7urVBCoyuMCSWWJIevEQCCyXQnqqMPKBAr3cyA+3DoF232zs9C4WoNK
/4qZu1v9lrOcA2Pv5Jt+WcG5r5BSnod5annNGYL7x8MmzalJKSBuiNUIJjmprX4pZ2AVNzpHMBmz
cU0KIDkr1OUbI4NPWE8wty24oAngUzmqYcRMZWlYLZIa/Ix1tukuQz9nL2WJxzPiuG5vLKJCMspq
jiI/O9yrcA6F/oBlfuSb4OopioWAFQHXq/MebwsCVfMxEQmiP7tQ8suhKrBHgib8Fm0jEgvYr9vu
pOp91zI/CwcE9KPZ6ieLdfldMIhk+lPC5AhZKapC05uFd6UPAWeE2buEsXOTVNqW9CGvHl+3a9lJ
BvLWithQPBHu+UWg5OqpNie/37FGtWGuVaSkDjLCi1q1ei6quwY/BYnA+PycjJkPo8qjqFcXK7aD
Tqlx1fotqsmCJAbaXCvvi0ArP7Yr5elpIAAFPsU394fggVEo0tUXW9K1pcHIMrz7x2NQkE2j+k9T
BusNMgJLBsvGlk3rjIOJJsZmhKPBmOQ9NXuAdGXLmBX8bIl7wjVH/cZaCW1h4nZrcRoCX33byOb0
MextVFjp8bNsq81MSZ9qSDgn58ugALLnTZUM1u0UpsfWC/sGi/tCt4Vu1SiDiy7rMe0Dkmc57/SA
OvocYNKmdLftNups5ye/lYmkMxQuqrK4BIUt3tOEk/Ur8Ihf4iKOsZv2KZ5fvmyJUQC1XRlIZGKb
GK85uJEf+tegyEN86/nLr9pE1z5TLdAYCedqva9bdur2ujhrcv5f/DNfbGal1ceVW+UEDhZ6vUsz
G8QuZlhL40gaY9VavBZ4n5w2SoetvVlugATzL6FMz4drgYYoq4aP5PNHTGmOvJulaVAVKdp4+24u
E2q/YcU6z7fQFES2M8PpspF0o8cVz6o0BX24j8AMG3NS0WYYw9FtHN+rdEbWbVcCnIMT3h/jawoo
OKfJSHbNNBFdvHJ77b6uRs7lPa/wtL1hhqqjjckWZf35nEbrCwbkrKljwj4hf7tMOPoDfpTy45gD
5QvhkWrh6QywWISncn/DkBczml66P3RyN9gT68KHe3zupYv6kr3dUF1tIi6SIdD48IGYlFaK44hy
en/vehlSsJT6TNaPa/PdjwQPxRl9Z2HdaQ/4dSHV+b0oq60x7QxpL2AI073b7W277UNik+Iuzhu4
XnVhauI3HJxUw0UxkLZzWNSQW9q+zmSl1lYkhlUN0fbIjMvM02N13JJ2aoTIvfm0fcGWwweqQkJs
aT9wSFGKMRcMaeM9qv0woCaWb0T2kKmgpM++VspAyLNMZxi8Zy8knXU5B/HNF6oOkAFTHgz834tm
H4zmsEggyFrN2p2mHyCMRVxDmlyA31iSF+KpMC+CYYlDzKx63IdIbiVF3RJ+dp/iEAlNAHc1iIO0
ThcOGlFbmSqIkq34ycJ1xDL+qZaHEkKXfhyVSaLsrJbECxsxhpOwG+mBgdYy5jOhqk/28bFjIBl7
ZH7wbryzcrZjp962fSqAedEJp+lBE1tygcQoyV+7+32ZMujuDOBdozP3zJ3F1oisixiydd4JFdnb
krAy6NDuI8kEMV2pTJYaJ1SukGZ3N71v5wvVJUVZWKHJgXmEU0/jfligeGXDwQHjoYf52LD6tpZB
v24Ia91tF2TaaFr4UEPNdTzQDzsjf401fFgRxK4AtgqC41h9+NVAt7Zzb/STcJoaV4jfzS1l2F5u
qjKbSjaqJkGBkGMC8DNtEiSTvgIHy/rigW3z8HCt0RwkMtOrMLgyCD3S1XLQRFOchKatMgiKJzhH
PzEK/t+1NXUIazTjS68spl9vm4isuz8iohW86PQQ4sZZ+z1L23inc5+2Bp7zRDCwBj3Aneyaz0Z+
y2t8b0rZKpJkEL47NK13hus0+aqtgSX99gxAJNSmSmdLncT/M0NdvZkt/YGjR4w9RCTEIvk+2wPu
H3nxhayay+ZCjQjnax3eCP2MoM7qCinJHQNpwEUloBOsab1+yceyVRlPbGL5+zNQTq5+lnEX2G9o
B9k0IuN924bIQCOQzq3lb0PPlrTN01ZLwzgKOisi+nWGZLoV4urwk0EzDAO/aC6LDKDomJ2gqHIT
HMYwL4eDZGkM1JQAff/rcC7MaFSk5Fv9OgJqZPrHEsoIT3dJrwGafxviiAioq/hLv88yGmV49p5o
t7TdBEsNvjlatSo+H3dUee2zytjV0p7A73Q683R8BG/m4IjwbZRp5+VIbCy0MDR8ItYaY+d6XA3E
/nK+kuXDTHuz9OkwcLB2tCJW/kv9/9usmJWLo5194yRxkcRNqUT3joJ0Z8zwV+GKqEMvbhHadI1b
gh4c7PsLt429TojtJ7iltrdg8OandjEvCRFW3HgtcKQXYLfha2wlPnVdIdFjNC49sJFuHNfof4Ue
la+6U0GnpJwcG/WhPKP9Ea5RFk8XNwbOlaRSw8RSlWOqKS3cS2vqTGzwEjj+wQXJN4iNWjZ14W1I
1qkvRQLx0rWaFVRaKpVYdg+nbyT+oTDaS25Tf0RemKfuL1TQfSBbbX/MWm1e6rzttzaTINmziZEw
QXLq2jGslLxko/lYy1HXCD8JnuloSWQWoT/ScT1coogUJVnq7FLNKDymcy3DetsOTa3Am0f3P7E1
4TnBcEZnNaIpb0nTrQ5t8MjuSUhx390UkJhMlLAzyIyRxMUzHRNelwRzGgy12W0oF3tSw1dq5qS6
+Vay5FKo+ZCnASSc98glKlntqQ4goz9iy8nKapOGC3BFVUrxb9KKwU3Ae8FKEJI71CkWJXn9iJwA
2pP6ViAoEAvhsdiPTfcYJtCPjUmmi7hobuWwCJFwB3oJCFmQLdj+ommHtuculY6kDGrx+n3Y1odf
DVSfrgMkXRoi01axqWxROl9724ThHOKDcQI50WLhu6tCh2/+R1uaShv1oDay395FPZvSZJFLpWqL
/ZlHzC13H8Xim2RxBPQFsidVM0Qleul0lAKjo/8kwjUcQhynDX0aahnJBEUQQXTm89IuetG5ejFC
azAsJBW7HBfTU/ot+8tLxZ6+wQnXBpIeM+2hBUld3XT4zul3LbzV+D0PWC71tN92an9gweSllFoD
a/6kjWL7T42UEhqyHgr7P+MA+Xs857mSUB5gta/cSZxY4ere+Hq5MpA8BBlujI7iJTXG+olfjv/C
UBBdi99kdDriK9h/pz195ASG6ifZTvyjKvhUSAveaNg2yvvlIcLkPIU8/yMI3tlouMQrJ3NKCEKa
pqYCGo478KC7WZfM4/s1wSH9EZWx6TuMDFdDLYVoLLEDcLS6mMNnuR5cppTEsGMMhsfs9qd/uOE4
to0X7OMGJSba336eWYQ3CeBMZLKQe/vp7OD9fbslka2uapjRg9DB0jQJszmL3XETXbfhhApgokgl
M4xRnQOeKGtaRMKvWiI3gJnGfT25GQv/jTgxPcpYtM4rakGLkfVbpDo4q1r0hgSx7fCIoC42HrwJ
7v32vwm5QhEA99e5TwbNfeY9bON86ftx27CEYfqL4SQhY0OzIRWYEZylZfG5mIrsRca7HlCwN0T/
YFp26WvzqaHVe7LA4XRpoW0Nkcjz26dPuTwIHfRv38KWiWgHQd5iFtvtQy2ljpTJJQnvfOAXMvsl
f74WjE4yIwFvtZmiwwfdmUkHmrFShzC+uDFxnS/DZrY6LPt/dlg5x3P75Rp6AJyvuFjGZ4NZdLb2
MOx9ZtyAy9QUeBkb2umhgydd/ryx4ZNxsRkPy04rwa6YXmL1NgdBPX6NbZdkkOMCAhV7O3yYEb/8
A2IP8lmOxtj+SSX5lrWxcM3K7DZVpMqLKFrs3QjSQPE+s3UoWQuiCcskbilViiOMWUgJjuHfe4am
A7MihGY+OSKTSPoWlQmPYHV5wdA6gYmlCK7CbYm2OoQGGre7P6YwiWMxQKVru04/pxrn6LBp/6ZZ
k3cYZ8fO7Fz3q8Raef8zjlAIhg34Pkc43Hj9M7z0hStTZXAh33PULwV8gZIDhJpI4O/GLDS0ae+L
+pyM3HxuCDZDrUOMuQWhj78pjUWOXOggEw/sG/lns8C7wMXpJbUKe5hQwoHHUHon+/WaJxwvKXKt
46jKC8iw6Iej9FH15uLOF/OBGMW3Ov2dQ/YaQE4gfhHWetkukT3WY15093Hckb51FNG48odWwVlT
TAfms2K7zog1EcXi2xyM5/IAq6/twiM/ju1HCt4vVPlYaiIy70Af5BnPWvk0l4kGKYE2Lv12Oy9B
XJFzjsoDeF7ZBFMNrt2AroxdPoL0ZWCEqoFL4duooJEMhXLSgooBezjJZJki6fpKuoiH6U3uTeaY
C2OHA2jmOoY1yFN5KCHTb8s3R2jrusLsP06eQqcOvmzwG9AmJ8prwHw65rfoaVQHs9A6h5qedyVY
Y+Dq9iPr07qhqsFMpjg6ePB1Nqty25SCTxj/v4L/AtTEzjE+2yH+3ruKwttD2cm/EaS8Srth5iOj
GqzQwM9k73iUi5omXRSr1bDRyQ35z68t4LSXxkkyPaQ3v7JEdrS5iAq0FT3GvXIfm845Vklts9ml
CiU9sNDT3gy5TW0nNu60SB2F9Xaecv/WD0aoZCnCqfMJ430YoUBh/GC6KfkqvG/9ywPHmvVQQRty
Rm/MTrKKFWXRSxtJPWs2cvO5nbJqz0C1k7MfKQr3t4Yw2T5o4ftHnNCa7TAnh4uPWXQ3kbLCENrX
fj1q3syl+mz/S6n7Lqx2I7JXsXxJnrn5Y/cTFLihxP6y/QYg0lGJY8jdrgwyRRVhUsoAk0wn8lYt
/3hAPjd0iA+DAMYb4BRQ1EP+7Aua/uxO/Uqv6bXqJDvHHlvTgjcW2fNBW45QTiWV/M6P9BziHq7h
tKH6KYCUriI3IR4jObSYvvSlJLVqoK0k9PqXCtH8BecV7IOFtd4gFD9ycWjdySR6C3z104DiCGR8
6CsdbuiDZWIGkLyut00SkAGsnUJVVpq8AgB9dk5sUWu6F+wJM26zZY3Kd+u76PE+A/F8zSSFHgaG
74oJim3S1eplja7pxaPBIaUPOa49q3l53Nf7hZjgk9ggS06VVK+j40yeTFA1lSyGsNfaJRg4+Avb
gBiV42oXUeMZZ9r6mZKgC/qKZiaVu3PD3b5E7Fb0ClNKNS88RE+eVFAJ0c4L1AkZBDF8zs35/2Ls
WDCXWHaZ2yLN7kc17bGP8hMJGs26MzHSoFdANVkA03Ub2JcpYuA5icx+v3Dl3RApPLWJKqyTDPEX
hoztjw6UFRG+rMYe3eIaKnU8xo6R9m+X4OTvJvJPIUTdpMQlaJQgIkta869Hu7zPy+j0bZ0tw6NZ
xG34sfc2s02N/a5sZyHLwZPwbRlwr7IODbf8XEAywQIgPgoPYUjgNHMOjX95+3X0IUZClue3GFp7
q+3Izl2zSyoI4RvzRWSPhXezyixTE2pibVZb2v1LJQo9AB6k7OLfyIH5uMEIceGu4tc70KkdL7DL
1H7yfLNRmIm2ENeDHse+Q+0mgmam0KHUqyMX/hXaeUWgggqtcmT9fK6ax/b7NglE7czxPyGqCaj+
u7GSKWjEJujnceAILiMimht3ifN2YLpcfosEIJo5uCdtj1mhrssY0t3lzJHS6ndpexRsfvRtAQgd
NfjnGoRS8P0nv4dzmosL3v5RU0f1ct8ZhKD0Niz8FkDwXRs8stP5bQz/RnuZ4DJJ7zJNGb4itc0p
4t4KRQoTQDzYE13ky+qpPzGGNBi0bSl13mzaiohARGvvUGTDHPAtuL9uQkgHJEF5q1ywcLcReWEb
9N4+GcuRwcUaw23iN0PvVa77YpNA5tYeV5G7RG0rwEeHCtMmYzyOw7mymE75X10SBk1+ak83lHwi
9RyV3KL8XWmckNmnq6RPU6LqtF6A9iAx8xWbnAhzFJsuZzmFenvY5aB6+JdXbwuMTkVQSvQAawOL
9GZ5xwD8J2uDTf/V2zJQZnrj79KLSMHVD42elr2QVj4ygpiy/kx4FVievY9qKzLZh1ouS1pF5gZI
b8AS6ePDnOlLXWnXxsQ/g1DULQEgKg3os4c2P6TQ317vtJjOJFedD1KoKuw5Wz9TbDII/YajBIGR
ByPcIg5sXrRcYzQ1M8vw7xKXQRhOF6mXNiUMrJMCWKHJCdJ1R14xBHPHDCmFDopQ165OzMp7K1om
tBTHf372rquj2uJBX7hmw22pVnrx/GaqtUQGY6OOzfmsYictPZh1oLluivhUrJDYvY9yATiUJX/F
8sG/J8PxQCDvJ7yoaSTX9UZVLrin/uwN2cplRg0hEIsh5BPZCmLDL9rdYVvA85klFX4JHKKlpCfI
kLtLqhh1izfe9DOhly8Vp2wOddDlZZGLgfzgLNZlG/j6xMTQth9TzhIWTV49E7LDoOGg6v9rolIg
tNvAvp69Ei7UfTV23Vnk+RIXmhEBvwnGHaiNQw5wqvuOqHVWOkOnS5ZtGMgD9+HpJ0fuuCVxsru1
oatinN47l/vEgUWdMvlA+AcC089Bvu7p27NG2XD0D72fyLXgsYKYQrXgOSfOsyX5p5sgZdrW19jJ
8Km24Jpk2mXcJOhVwa6HGLPNAXUnFMA6wymwQlOcWx52XVu09Ww0HK+DrTODgvocp0u3VdzaWhiT
AcpyIlY5fMIy4dDIdgzglrGUPqzKD37LamnYiNK5usimm/prGPdF9WT19Nk1fkOgLYnaHRTXS70l
3uwzJbafvym9gE9FiggqQmEzCqsuroVv45CO8Vp1AyTVNSFdMQB8lmsy4NCBhwtFfTIC2uXJMrsA
iaBN3a8STeZnkiXI86yPLRznlpk6o412v+RFG/LWtOefY60WzXk09dM+hf6L3V9lPr0i9AQxU02+
szLdjZh6n6ooHzecPtNTESbyJZ+deXO0UzKfZJlxFTvv44h/FuzuGMZ1Nx/b/zeV0qPMKyCWwh+b
jutlgyxSJb6Lvt9fspNalMwhWm/bHkW8XSidikp07M4ceCO5yqqdVw0jyTAdB+Htecu6ji9Mbrqv
ifjkGsjsbKRt/mqyJs25OS4gVuAWaVejJshQW/xGnpdUxj7ZP21rdQlaasCwY9p2kX1FMy4MglvO
MaFyZgGpMHBXkRisEfkqt0iaV7bUSXLouaB3PBmcxEl5bvqp6PVJv1zYyNaiV+iLF18uUTlfRYs+
KGdqCEjaGDZToL8OcJviDaNuHGk0Xt6ausdRcYnpK+BQJXobihSFRCk4kN3/gVV1GBXIwKOXoQNV
N3Foj1QOWXqWrTasAIKvZMMCjbHHJiUO9IsHk2ayhxdPXWxtQAzBg+4DnJ9/aO48YXC5FA3n5/kN
XH7i95m+gI4HZg3BWJ2NRXl6rd04GntwS/LXzC5r0B+Ep1WD3CXjGeyfmZLs4QiDyiebfxldTk5A
6T89DCLxPfdbE8U6dMiXIqd1EpL6yHCGTL+Jmn8kmaaeubcovODCmEOR6pDM73y0i0A87ewQOHRW
yiZhl2b2jG9mUcJ51/lUFQbb1GdXmKAFI20JZe4ra66YOC1GMWix5ugmJJd40nglu/Od0P45OExv
+T0Yp720/FzaRUfkLyTX1IAO/gT/Wdjm3nYBrBA/PoCZwYytLUGiQ7EoPY6QHlfiR2UKcYgyNE3Q
BPt5e2Lo76Tom+SKYCKL2RVP057nLzBdQSnRdiwuNwYt/0HzdNCc1KogmPVJIm+IWweLxnaXRQHc
rnFrP7AEhUJACRd1FwHy8NdNuCMvkqQTYsg1METE5lEBwQVUMXdvm9/V+Et4Ivd4Mra/6zv9o9da
5X4r7jjQGh1+ytGvOZq8xDsgs7BBCzCqRDbwCVDfLXOMthDno6y2bKzqcH0WeanYMrsW+kAsWs1+
7MbRiaUOHYr3aRC3yqIYceLuee3L7RNmcrwttnejQlAHkK+swduETXMHMVDj0m+GhKmP4Ym7EN1/
MsIizwxFY7pNkoiaIrSyLLyqy5zwuTptEpwlXNaBEUeZ4asUMy+Qbe0x5ma9VaPGuDjOUpYP+5Tq
/YYu5xtcULoTPVZVl09vvkKX52j7jogABQXaat//cHbPA/50XMSPbpoBc+VV+62XU4sobTBziOZr
jzwlhK8/6L6DJ77WqMgHNg62MKWjOmT/yIJMI+8tQa5kikx8PUWh86q2dzC2mdwEZuIt/F3s+S/m
7p/pqri6EE4ZjiLDvSdZOZD2iFcZLjF6hWbJDd5PEm42LB2AMDoji4p3almRKuECLE707VoWWmi7
BRb3R/HogN83ryJr20IOiZJ4/gtbxPODtXm92AL5IMKZ7nJTi6y6UGrsPNPK4L7T6mSaoPSV5xa/
RXFxRA0RjuCfBAtUrQu9V/11h2q4yaboJPUTkmI7oSaTfOMF+a8I8dRaexlXwOiryCNQ95w9Q5NQ
bNA33tSjnogkSzoMOokSVttDFkhdTbnVHjp9d0Hu5hQMl1rt62CLrKTycIGpMq4zkpwMAF6lQdNr
qO/BaTfY0qzluZ4PSqHqGsK+/J5a91vYdlh0MKilQD9VB5etIjYob6cX0xQOF03jBT36pMayM0C0
qnaVCvZo13Jz+xPIgoOcG4NgcBCYVkl4FnGbIIJ674BdIA449hko6novgZoEd3+ypyXXbdLnO7x0
bmQuspbTiMhOLbA6YOSupGiVA+Ltb54gc38wu0NIcbcH05AF4DbOv33Ah2AB+q+vgi4a7d3WRAtX
YYJZFfdCWi+eIqWG5GtE873qvLTcdI5eh3W5UGFAhdptC8H2syLXuHSGIgExctfplEFv9uVJWjev
MppCJqCYEWBSyEdAiNcSDNd2tyrL1FQ8LQi6+l/yDCFtOx0U+uJUy9rlf7oVB0iQYHDlQ5l3yM+C
7fmhKRzNT4QCquQMPUASN5HM06jb5Nwk1rIsikpt3/zVaZTLpMuMtSzgSTmHIy3zX6TLxKgvCCTt
PWWeFi/1UIRkGpTrVlGrszzjLxlMM9XJNjcDoWfpA+QK+Jba+VP0smAZbVc2LFQfiHRG2mwwv/Z6
s8cBtAxz18CK/WIhlkwYdnhH8ptTzBWMuMy+qHS4ODrGoG4AJTvPgb/4mt8QAFNDm1kPIWrRED8+
ugVtPvj+184yrbXvJfoU1Vksu8cl61YeoagkVQsbV4Zznex9q3E1M6/e5chJJ/7jsBV4W0NeEp3+
eVkrSis9/D7CbdC5a1sv+Mv0q112jrNkiNmIiYb+lp9WH3vPp3HalXem7keZpL7dKWPAsmc8FiQv
RNDR1Ks1u/IXS0gyx58gebG/naNrcpT615PaC32hC9wBlf1ImLnQXbm3eWFXHvOdF4Bl1UHh+RTA
ViX4YXtZKlwgxe9SKnHmgoIOSKyg3AqkyMi0764sayInNnBHTJQ2FbcYeC+WEow3dlS3BOAWdIpP
O7wlUcbt+VRoUpU4jAo/83djzX80D9W/vg9/p2xCwf4csBeDI0XEYcBeaRc1x5e2zQqyHY81MgRm
Qr7f8IsKd33WCzmDWgHQzeOJSoYg3zO2T6078qdGn6D3GqQPFGxdwvDbpUo06u1Ntj6VQBW/QBIW
SYHAAHo+6qUIl137HtJ4if9QDM1KgqX4Scic7fnOJb6Dx4QXG+FW19oZz8PzDPMzppGxOdJXLz1U
8+hO3damL3CLCDmLLaxidyJ3FkLqIvoj/BCdw3qumXOYVN5PT7Wx8pIbUdN4ZwssmT/keV1bObNJ
q1s3imYTwXsgIiAtT46qYdvI9gDFucX41pd297/W4gc7iS+eMgDyZ44aH0PGgFnxErb1RKn4CQj5
m9pLtgmU/SKz1Ua0PjM7EUxx4tqmP1L4L8zY0H92KVFz7AtuhenHlEhE8iDYkP2bqJua1j6oGnq/
EPDfvqcMT6hocXWIA44eu8U8r9zsVEfXkh8dGQ5AWV79BgaJyi9Gt3SdEcT6c7D8W8w/tffP7cG7
ZLizKQ0ik/nOwPRgJNdvlgHWo6bIpnDjtGY8qoylQtetkaV4v6uAh5GH2fJd4FSIuo1nfkh/D+8a
T15/VVMNqmT68r9FkSIOHwQLA+PPiuSIsBJhWfhtrKv+t3ZAfrGGm0ojF+PxqtZJDnAPH+cqGiME
S7t9+0KQYBs5t/qKJpRcDowGvlmQIaThm0LAysTby+JFJPp/7nC9oSQmqY6okzIhPrD0gBq9umGu
zh6w9EiTh6U2xNrGMX6ntWQHIW1x0+1KCXRKTasolJGuj9Jj4t2qvO+uexjJS01X7NiRLKH7rGD3
JGdqbnAZIO4pawZ50zP3H2nRBUubNE80uUg9NU8GQ89yOnhOsn4KjI7f2/f9P4kKvs4qSb0c4zOs
MjwUba2lTiEVa1UeakGLqYcnStfY9wVXdUUpjEotcdP/m3mQJ0K1sBSP4dVOnzTM2GQ5vk38EjNf
8kNMVt71q1rAgLOIupDJkQTw4+uMcSSksthMTdZSuBXIDkgtTYc9WsDMpI3qHwzv6x6PLe9uFWQ9
uNcRUZCXDGxpBTOJdKCzqmgA4O2b5AdfhCHZSp8//iTUS2oEpn31C5n4579obI9SO46Tfqtntd3O
VyqBdVsPRxZWx4TKjwVwMohn8nA52ht1VPaMRta3c61gJZD2joDjv5YieOMLrmEwFnx3yn8DHxxv
sa6/1DplPIZ+fHhT9WSUuYddo4msPfdbh3GEBlXAqK53Gya0NGamMJ0fnGQeDUBbnYaDE2Wv4rbS
l0Z0NIdJTTfvnv8rjNMHOqfKctFuxabpPsiveH230HFdPKn+ZAs7K7qQFLnZsdisdFoZfzhvvWiy
Mm4xR6WuTmeiKtDUszA0nHYf0lYf0RBfZDi7Fo6esNaQ0QRz891PqyFSmsiGcFB0fsIYqK0yBHf7
Brx2e/nzSehhxT/gIEr9p2HEM60LXaT8iyDR2EcuQ28aV6s0EJkkgxatckxgFge5z+tkqnBEgtMK
GMDHbuMChFgjif1OlAGdfgSL3Dh+PoIZGPw2WsrqYTuf4J1blXBkIxV+PuZWuvS78erxjeq+aWPg
d3q2SRnUDHjGjEK1ZiSjAbEbLq5uA1df2pU0SLGtbV3sojwRmNMu0hrqoblJ+EznlJA/t8Y59y1q
lZqg+Cu0j4kCgnU3sCiTbMKc3s64QIYY/J45QyQG7X7S0J/29AABtz9kqJ1pldhfJV9GLUH2ldDo
2hOelBqPaaDVJ64GJgqLEQ4fr37Dsycujy4wlaMHGNx4jBFpWb9179zKfG14PvxLSkFlCj8pI9r6
IXhBKv5N1oSKJwiC9Je1oW2jQFvcZ1CIgdAhgteEbOawFi/Ix9j9VVc6wXYQSDelo9d/OAyyFIti
aqT9FesYpHPoh4+p6CZ7H35VH0MLV99GgxcebotFa4VJkXis4XoW7zNThe1axCotGaGitoe0TQLM
2Kg/mEFfte6uK5UUs8/ENrzFqForSNx1jE4TwzR96RXVghzimrhv1yKe8xKwn3X33Yx9GU5RfzFK
s/6SCpxplM5edjDGB/FIfhycVf0KJvNAFn7eO0nP9jLBTM0/IE0E9g2ThU0OpHg9CHwEXIpkuarU
UqMUy54L+Yo507kzzFuIfAh6v8/PY+ockzGxajejCKniW+OuFvjfd3LrUG2fawX57iWsgS8MtwHj
FktWF1y/zLBk4vMhU8fx6+xEm7vPo5km0HWA4QKCoDpP2CG65Nb0Wh7E8gmnu7QlR+3fbVfyYLFi
enpYpqimkN5kLI6vI0gHNErCV/liiOmFPthPutiV/vrwSLyaSuTy4gaTLPV8fC7tdixlrtCOgWb1
/T99L71XYX+Q5O+wbnnuZ0fjv987zwREAQoOClfECB6FU7csvBVgycDtxyOJ/u3DEp4mY66YEMKH
5ywxxx/uVEQ9HAaEvWP6cLewIkG4EuoRAatwvNXepk4tqB4ToNGgELziTz/x6fWXZmiCI3ay5ItX
5RQBGDcbaivCu9MpRlWj++zzFGJlOERFErJSIlPiLIwd4yNzUoM2raP1aAhmAVPA+BDKeKFndJDC
tvZ6A7pHvB4tkGHUbVH+uMrVd+Y3JnNaRL7mo34u5Lrsxo8lvdIaruQJ/X4wa7foehLa1bEgbc/v
IG22HDlkbLHVpBKkZ+NOAb1YOqO81QatgrQdxAITeEMPr0URs5X8zS9ehHzni5//MiLyHxThjqrF
fLOME2AABUp3O6vQIJuEzgfAE1n8TmRk8mVUnm9MTbclUyHKx1ovh2MG+JuAnN7h8KRH58uutmIm
MDAr5mUrTtBuG7CYcKJlSfRXjgi/5r9EX0SDIkEgP7nrspSBAI0/FlzXMF4+8k+p53iAZt/+Swpa
UJrUHEx35+y/Xc4gJmfwr4epIUUBoJWRiJ3zxAjX8oK44veTg6h/FnYmW/ay31ntOn0iPJlDEd6Y
/FMgQ/RpPARWdJtOQOSTfpB6mpAgZVEm3/S4wX5RfrHCRxMRR7sitj7YtLRBEtlyvYtkAJBWFCCP
HJ2royUJdBfMErEnGMbcqAHPUu8w5cRCmlon0qq/pYt9fVIptIy8mDFI5xuyj2fcvXCNC9e4MO9n
SwLtxPHyS14AGURjEkHSK18a0LtVuQqSKAw+/G88t8OqoWo87ZR/Y/FxYKibgI3MoxTQDuLkUutj
XjHf6WtqXBjIJgN8sDDOdXAsErbde/Z1tHibQ5LMHASpyGkoPW3tkqa3QE1zu5mzhPJj+e5DaZPd
unPK4onvij8eOEGdmyyefNxdXpWPM3F/T3FGZYN1ShPe+mm5VdyNaCKy7vy9sDhnukZYOl/M1nF9
FVepd5mAMQh1d82Tcd2Be3Qu432EPMmNL6bQyaUKNP9vG7bz7rGObVDNmb7QjaCmHgH9Vd83xWlt
hp4OLXy/W65koZxEhzy1H/c5NF3UaDLp9t1H5XhIFAZrzKLYQ92gOYJWetddTmT56wXGRx/DhVu+
1xKE4jyBGX4FOXGOU1iMb7gfBnGZvlFI5eie5YlMyIxLdZJR1P4Bt4R+srGe+eLbBydchtQo1sct
eOkVEAfhKe1qiQdZxqMqHLwb9L5N5NDb53XpBqsHZBFidroph2VNaf0omHeDGnwT3fJBGmFfFfBl
C8w67qgUGDUUAjwOEqmH2QwCjFuvAklc3hec2J2YVuQux6QgqLeGXdxaLrHLxwRvan7AMNTu+2sG
8u7hxjqAOqoAGqP7/FHL0Kj2bmkaqmRM8MG6gd9TR98uOrcyepEZOqpPOEfo8HiA+fgA4QIf1eZL
3c78Ez6KwEOAKZhjQtHcI0b0q6Tufqahlk2gkLxqRkOTjfkOumaxyS0nQCW+RDFytveugUBq6kmh
TcNkjUDnMNvNWrSRDx6dvLeyGP4FWP9XBCgRoW3b9nbQH0CLGJXzJHCkOLySpNz6ju5jr+zjyoy/
/GhSL3jFNeyVoXO4jpLSV9dbsRlkUgcUJPNcqmVR4I8Vb7Mi3dXMHw0PlOd3+9ncuKJ0bKkZTBUA
dQNCOtaqdOhk6/1XVdA/fIeURaW1hM1HjNAYpODGzhCF0KjuNteuenea+f+we5jQKr22iEWFNHZx
R91ZiPAMSPOmyW/5tpKX04AC0pMC24pWxCI6sPIQV179jOMFngW7WQCBLaVAlCqItqFnK+nVnCKN
6lo4GmhD1/mq/FSduiAovQBlgVfNEtm2JowwdnuhqARYQsF2Uyv2VKaKqTCjv0nP3wcSVn6ktygh
sdXSIfqnAOAxoVpOoA99P5uO7HLL87+nfriANvXmrH7wMARH2REx7MbgBnnVPulW7+E2LV6qWjQb
OHCNfbD30qgYXzUqRt3dphKmkf2xjGBGdIKcro0DrdtTZ5hXLl9vNxPdDRXj2t+9FIKCq2VwzUG6
rNmmJCYfCShFh+3m9g4qiYIVdZ/40rfxX1gVfSQsRP2rDEIujyBam1kNy3Fr01/IgOeC/vVs0ike
yo35lvI9fpL10QFiI3k1a6myJ9Q/ZDtcDv8mmRT7iTsTHvAarPHFTKgIt+zdVgjV0IEfM43Ic3U5
cY/tnyiAnAQd9gX7CuHUm4p/kxhfyRmWKqRDueHE+IYi5sdy9g5O5JAiHxWFzJv3wpZwcl/qVjjN
3oR7EBR/hQysrFH57sigzZCwD/Vemc5cLkamZugdiZuNDy2jD1ho+VNy3wbvv/bioV/txatJNcA6
Nug101K6GLyptAZelQyd8gq8juUX0TXmNhTYZ48fh0SpDTAMpJ4F+FFYwlg1ir3OODqrSzsxa7BP
2/gKmnD2mtw51T2/BAb93a3G810VoQPRk2nWKZBvRP4P48Sl6xRK7mDTZ1ELI2wP8N/b6WI5XOED
bpawTztfYO9JPvlfrhESIBod5QtkBKcVQq+F5bKsS7SLvfONsVNt7btnRoL/UHlJj+/40e2MY1iE
EiA6GlKll2EMadpVYebj3BqhYN1V3oH69h5MaEsG1rbmMAYZMf3jtkpJB97ADqw7A8NmrRMpG0sv
it8zgliF3aRVh3mT65+dZMDlfey+DKeY5xt8qw7aHqbrvJ7+8HYdehbm3Fy5d4+rwVGjz5GRdDC4
CsWmVIXiC/JHPBw1wFWLFaewsjwU6oTAUf/FS1M0S3+1j3eNgPs/1qVKusqWeBysSUkHhZOPktxw
Y1w1un2lQMqwjytOl0Naf0TM0nDR1de7rXXHa1lk7gkRq0W9MIutGvrz6Dr8OLOaiKuXHkzfMrKv
66sK/FEk3QV5X+56glF1XmT76Jg1qnYqutWHYqtfbvdwBnmV2pang/y7ZuNlttNsjw5zOrG5IHWD
3RslKGb6qi3szZcRKvduHKFxuH4elx64mnCJlqfpYyC3GLMODXI7oYiS0d1TWdCt5+hmtHr9RPRU
WvpmGmZ+uiZsh814/cKZtMkdW4xONo4nht9WYHVg+4tycsmjsJHVMNEdx+bvAndW841F2aqdpPmj
jRgbWCwnt7SqS7QodkPk10IWxVGCD3WnIm+vCqg3FjfLq5Es6T7y1eUWwZ6Kk2CVJ/p5p3p3Tk7u
TvfomisyaqA2B6YO9ghcMp3A1/lloOrFGIzQbNI0EQs+H+ej+X8BA7PjbVS1EcUcdv3iy4Ny0y4j
Y21WbZV7jqcK/ebHH0tmPtNrKBK+P78bBqcGcOV3x/qODC8zzGk7/H/JKjRcDeBC6msq3rb4rUYT
V+LVBjak8njfPihddlvGHjPGbm62fLsLWPBAFIxHozy1vxwAEcZCrZykXkkP4eXdgVe8qqUEFkLY
QQeOdnsuj8uCnVK7o2LP90rz7pAuwQziCyTaJMpsu6mIiuyEh/wKuEVXcrmcS+pjnGRpv0EbI1mL
BE7neDcIrECVenq3kGKeD0DGGOoceuwlhGcPpYCSF8oKHjS912pa97An6j7bRLQos58HCH3P5scA
OaXePKEBlk4SOuWT+FwdDgR71ACjfj1HbC9GTgJu08tpfqKnaXmpxgZgpeEtrM/gxFlWzu9Ijwz+
PdWdiDLpLSwluuujSFrgigj8GAriuwTWtQWz9fLyfyFhGupn8/eHN4/Fo5JqPvmMiEVnP1pCAXce
tGFOaH6IxrLo0c/yg1o5MiZC20+ojsHxgWFt73CwH6kG6jkH5GUHmtDwAifq1Rs3maGoOfXVJOJ8
mXpl3wUg5qIcJM0TKVjymycYJyEtVp/EnJ10EftrMlkUTBDVGOEyY+5gcLfw+c21KN6J7QSrBbSE
A4D6zlU628vuHNtHIsXb6m6CZbukaZcJ2Q65kDxmfhIcT+53c+EHDXDy/Qy0BvbT5yG2cJ3g09eN
Ixy/iGH1kOIHXcmJ1NZSskFSD0B3By18uDu+a660D2hm1gtol/xOj4EhHvnAgddzg0pQgSuuQcTx
1jqDtGbdkxFoVPVDrc2H0Fkt03naz5ahWwzfok3M9J3gQFhrzqBnKgoL5S4bHlSDFMb8sMKU4F4d
rmFtllU5abIw4Ta1C40mot6yP+xhhE1LslEu+UBap2ZPqp5hc1VPbLKKIETY1T7Fs/X0rWYE49Wg
DFTCdIub2audecg4YlRbOSNgb1EO80BxfQeyx+ollk7cTDM+f9ITYjINtxKXothIYSRI5SKGhRiD
mEg0jVdBwgJCUy6lTfBQAuj5Zb3w+SvOwi3vZik+KbmugQ5/3Bb2Dpbbpkg7k7ztovAVccePpn+R
PPpwIqiyFX4zD9DB5jgSww9AEANaqDHUIyhD8Q+/tMWzeLXq2uZq/PL2dvtbk82QsDIvT5dFtkqk
rb/lI6j2/u0R/+LVbjkoqDIrWasog8Ta7Z3cPwLrcXloiL5+z+sz8roTqECM6BJea0x3C23nLIjT
AKS7Rt7VWW1LLtj69SLdk7FtbZG36wy3B3vKZJ6SIsSmNsfIzlZ4D7FtxwO2Gr4U/wTZwuKwZJh8
1ZujREdWsMueotOQ6Qbz1FxD0JR5kzW8chGwudghed//ZWXhMRVB41mGu/FHUQtGGRpqvhbVmQXW
dX5UagjOrJ0KQBzWNw0FnVY7N7joERDqYEtkV7gHxPAJ1gBA+3CMDqbnJp3+eckYvt/ozePQ9W9L
H6LN+Z2QjtkHtcUZE4IVse2nYvgp9giBmkiFHCtjIWg5V1CMaJjG/1obZLbjhakuoK0+c9Qkuzeb
kneFzOXZihD1NNpum92enE58yz8GDAo4A4LJsKt5k0TQhK+DksRTK8Ve52HAldtFoJ2CtDqT7sHo
sDdlsgOZBtINcQpM89va8UA5d8iwSJr3dHLVcSHtbb4eQE3N7Of1Qv5nJxFhTJed7mEih/YKcNgb
TPTmNUbcMwC/p63jjFj9BBCKqWL/PmP5weLWD1qjlAcjn6M0JlfIVEhrBaxuB3oOTQzakzYtfUGp
ydL9Z5B0EaYaWju/S4b78dXoe2iVZC+2VQTIfZ+bfmGal+JyDBNkfr1ccal7XiK0mltJ/m4hST5G
CNb02LGODEI6AWcNCmQwbQUnthkmsbVfHQJpCOI/V+LpfsIjCp6Fxph+aKiEHlWYM8afKtiwlaWN
WHvT2ySl+M6U+fzVp3mG8twqPsiREK7WPvGP2xPtFK9o+nP8YG6y0QpdxxNdvmOtQawNuusHnhOy
0dIP8OTDYZ1roacANOh9BCNV8W62Y17ssV1ToeFQfxaWzNS9m1K2y+CP/6OeZcnh891Ym9YUexQ+
l0ddxWYr+xBeJrL2LasG+ICIgMKksLjsK9oYNPPIcMOhzICithXhsaDwTthyF8wR5nRpSnl3Bqs3
wWEKF49V0nucBwT+RXcgclqOj7lzV17AhgspkyOvwfVEtt+7n9kt8ntanCpPWltfZF0NfKl7mwcx
tH0oXyljHwuFRDGX9SgR6mO59NC/KtkCrsZJQzbvhCXK/1bc4pp7IsNsZiYRJYF+E7csmf24gD9g
mswBVPCgzZm3O2U6rJv48PrYsvdqeyQtIcMOT4z05iMkWoMm11rcGG/7cuaUBdoB949EnI+Jau0i
7sOQTdSUFxL4A+UsKlGbHqH8YF5O0HQlFoaJi9/lBQrENU0qDHRFRD2XTEJhZIVSJzh2WvOmpL5B
ww4303JWRQZMiJh6A2RpUdi4c3HyhgK3Yld4RPf/0jy0FYw8b4VKtdIZ9wGpGXLZzVAdBKIcAVZH
K5+FfZX+reWZfR/CAMd19piNssqPLW3eCet0O7Kpo9YKAIiAqxnINUxvKWzqlAwWiSEjZve2yzKG
GRIjiAT1wVL1uYD4oeyknKstwh4PY86YVGUcIWp+UX+iylympHItJKN6CMaTBz0uwmc5g6djHLE+
yeI+b9FM/aFe+zoCzK/MJD125brAR3jqAmmAgvqMJOzvcIl/6wVjDoTcmePicHNaAB7c9aMS9IJO
svSV5RZvATIAQGpAeYSnAcKcQ3fk4NdYg5AGEUN3uL3aRWZvB9tuHTF9uI6JDk59YmSZd0HJQSFU
3lsaI2zhFt7oCBtbsIH0UXaECW9s7i2/s+IHGsiB73J/+iUQVJJj5dzW3FE/LuOJM9Q5CUNsL4wE
XVtR9TzvrOoVsruvUPTZfC26Zdfybs9BXEbxBzDgPn1xwBp3OJUK/i/1Ctv+FPlWjhL27vnMkkpR
dOMJ/K/PT8WrGOKQly/QBv9cZdbw44khIXxsqNHdu/TfIGkCJxuaC7lWGVzVk9/hCxEkbNEXSr5s
4Iakj4ecDB7WSO8/Z1YfvJjv2j89iq41DK8VQt6Qne+Xs+gnPdL6PDFt/0bq46GYrE6tpxVzNSXU
76xLuhQtFAp4q22PSmD0L78L4yx0u2CsM4YXAk1plBp63lgN4ZAG+W0R0LI0rle4g3d7ksZcw6dS
KRg0pONFEzLzcDxM5HFvZGI3RH1TjE7Qxm3116WVQGAF8Bif//CspIRRlGh2krKynWFVvwRelx+2
6uH5Oz3A1iCbgajONntI+GMir2Rpt8BQhxQZg6TFOLgDIAbztGNVntS18KfLSMY3gbNe2tjLsmVn
UpZW4+5uL0ML7Or/OXEgQKHmPfJA1rxegpBDPkLqa5t7Mumbt/go+f5xn30tnBNXJggK2T8p+q0R
Bzf0DcZHd3foEZKIGPgraRMGjFXhynJ1uXI0bCUFOyIfyf09351dhfFoQRo6AWZB37hpHSuB7W/4
+X8XU00a8QsMRG6It95OcoXzc2A3CT5fcu/bim6IM6TUsAuEGa0CMJWl/hU50lzYG9orN4Wn/Nn7
BXxns7KV7pEjpPLg0hGxGJaWfqUn24ZsfhZbopsv3buTT4rB+0DZAhLwttqjbOJjCrDjc55sujoW
lXZz4lqHHbhIToopiaLXHdXNkdBnRE53PrFHAQSb9aiZ/xY1Je6+d71SESwLjGnW9kHuy3Pve1N8
FUzYO3AnLwulwtPBWFaNcCdK4p96bc9HrL4DWFXl3TpnXqpNs6Mhfx/TJIQY1/ydaJwYAukHmxtq
sSxm5ZLgi15SzJXOuOZf+5wzqvjrOmL71Scg+fv5JrWDuGkyfnMr3O9urNMQkKhiSXV0Sxi8FYqZ
9qN16JNPDLqBVGQjF50FqlE2s4PDZVR1aeHE9932KjSUWfo9spvxBeIvl9PtrX26it0KGI0D9zOQ
fR1giwAYbXZ5ln3DgpELxvEP3H8mRAqzzVYs2/sOEAVOuG/AZvlFyB8d1EqXR2o6uzj/uY+n2i9U
qlzq3v+jYHmW0T7ewK96hLCxwAI5vU0fb2QBnnvF22dLhaCpcxMrrqQSzFivij2SzpG2GyQk/vpb
fInS+d//4aGqTeZCAjqY6wbnc2HnUPtzbd3UGt37YU0BOLKCN0uO9ro3sOgCfciJhurmNumQVUBf
sLGq5OFr19bk1f1qJq9F+NeHfOh3v3kwp7nl/lL/Hbo/A9wLv2g8VDxiT1+N06KuHjgPFLhFu9BK
9kGz9hDjQQVRxsuwOCnDNdNt3oNaSGanxJ2JgxnIe+xtcamFFTr1c9PadNvunSJlJntUI9Yz7pAz
LtgfeWkTUKHTKkSUxhUrDJZzeKZdJvoyNLKs9cSxH42KVT5u1HhMopK2LiBLgOEiFCQNdlogJ++o
s6NVfgPKs8iLn8fiqi0UP9XDPe3Sdf+91QR/Mu2pGrNROjXwyCIwi8/JSd5jPCiUItj/aoUF5fpb
QJcHgAMsHPwi192khI/Uk3NC1CzD88c/5ZMnIvUYQlmJ5djoHgLPB4TIjzZsN0S/3+d7j+ThGDfZ
Ohz9C8op4NxLrXyKJMsz57zXPXlcWzwB6E1XHuZVnnnnPjiRlJCPq85+i1VFigpfit7hyYBw5hJY
U+GG4/6xrkJ+ThpEg9mqTrwE7GQ54MmauoU0lFDRBkVXMrz/deG5z3mvyUxbiZnjIkMyxYKZYtmM
3HqgkXNPJQiBpxgtKAfb0+FD4cdIzJVXAXRyJLXqWids1hHd4S5t94FQdSyUSh5OqBKcl6U+44GK
X95kptV5yWHpTXThnH+EG9pztzXzynIHhzlMtWMCiYql9l3llLJK5VkMC7nLjTNUxa4XwjoqX2R/
nDsd4yjP5tu4x1Aw9GnydZU0ev8fXjOV/cSHjWx7zy2mjKT3DWSBAQsCAmTbMxWwrLZfyBxb1aNx
0PCtYHJjxHnJyR+0WaDOQb3AMpYx7Optvmvwxe9kUF6gkUD0pS5PWX0BfG0bHv5l+KOwauCulcGk
rGvUfkMU0eMujjSJjcTYv57PNuoiJ9PWY5cQrrRD/ZMvZgh3Lw4OQF8boBJ8kDw2dzYW73RChdEh
1rPm3LLrpLYwaH4glY6yL9RACbTN974GPJczF/CgvFtU/fVLAKZp9a6e65Tl9Sj30k26a3f4yexT
TzOEYkGc2p+conT3LmAug48f68gpS8rm0YhodkqNZI4N5yNGhd7XrvxKe0pgK4jaqpf2dPnjnVFk
+dtxuw3y8PZaruJVMhergGRbtsls4GkW3+stgpTRiZSglx93yh77s4AOUKfQMAcsD8RnUzF8WA0J
fP8Yr1Q9xunE4H04pOhUIsdEkVnXHA/Rgi/fJJmAG/1Rr+7qZ1kZDbWJjcIvZ3kjTVeVYYJU5GP0
FIZt1QPmP+XXFMDHWu3SU1mbVeYZ375VsGlyfB+tySzfIwEUPhJV/16vCvDAKDilMq/mjWZ+RT6c
8cl+YEMZ1pJeyvpgZ7BHMJw5zWk/YJVg8d69Hqv+L1jd8hItUfAJz8nyt2Osn34DRQLUgCLg52G6
Rwpxp8Lypb3q1hebyKONfvoVueDBjPxhuhANqERhrXyow0YePNieIhsfe9Nyl7fv/6Ia6YQdFoVo
oIpM/uUbfFY2egWvhpcHKLmnZbblh6fXdieTmCHcQamRKiTnxyACVP4//P+P0hpLk8PecHPO/oYS
f2n4+rNmLZ1aYZD7muVg0/ylUVApQDvOifGdyhIZzXcbYw3REt21fcPM4VKRt/2pg3NzeoM/ZJo3
kYRzXEHLaI5qFFrFFO8w8I2i3TS0NAo+sIWMMwIZBsQBs1Ul8G++1d7YaJBH+4nZT6TC+7yzr+XP
ntpBIJyi2xiroDzLzH95+86rTPYeIXKG3YgqJhonDksVwSPPysRm4RDXP3Pd1B0Nfu862PU417l0
kEGXwPlH5Qu0doLmAlVdTPA9iYzpF+jlpwpkD8PK7r+kJB7ewusEyVJ/hr0tYLZxZsRa0+ae5n3D
xrCAtsuFJTzjj1OkxtzUiNXWH5852ZuPZndvsF9Wq6HSHTcrOZXCqFmf9gihwW10CIGO49zZtTiF
l4QDhEIFlSvuy1RDKsCaDPnZXH6wmd8kWW/usCc4aS/tDvpqd8u+SW6mtYDSpdvCaVZbgUnXGX72
NYV3USIkC7zX8as3ldUOnUWdsBOQcUK9n02ybLtYVvPgBFQnNe77ATqlXkxFD3CGFL0tFrrwAr/Z
lKS6HQjt+3gG699fJRwTny56NCQCEOAQCwgzHv72TIjvJwJr38k1vN3HD7J4DYZ8NmD3McJpqM5Y
asmKxGcQU713ukLeSmZwkEmOFNlRUilIg2lc8mdDFDXxj0ca2TUuCYwTB+TK2HPPSsmgaIzKt+36
Y+RiAheaFg9LJRvdsPEGMtcAfv4qyc4T2Gsi3UvMBdX20VTTWADdu6+5Tnua/6YOzPbMRhk2n+Ts
wQsZup3Vlon9XBwhnbb+G8XPa1I596laJFrBPMioQOrnx07+qYsQeMSPIjnqz95GSDNDzEM2sAbc
O8o8ujL/nVUs4itR9rhWcyK01vFLzVhLIvvquh/poP3u2H81XPkfEohx3SQ8gyY+fOAxSUho3IKx
b2/O6OyR9+AdAI6NloJFZOSsoUW5Zdh+WIj8JX1eUx77GbbPl2nVQYY9vwkXEY1lTmogcXQHWkKu
Qz+mTHJp8f1mT1AgLM9L+kpZjORkl/Vdcn7tEVbg1CrF+cMMnKiocyJMxdcpjof81g37rTEvqXN4
1nOivQwI0hhoCk8rz9acg5yLvTN9Xo8Me64ljeb133KxrhcLTU0pa9XI3MrdTgwgeVJJ+uvI9kCC
9PmXmEDx9kBf9FE6PMoZ2KFZtJOHr9ndPxKUXpX9DuibP7W6U67TCNgA3ou4gS83nvkwK4UU9Itz
Syss4L3TRl0IFhVyVvEC7zYCamIUtzkHnuiEc21TvZNGcR/E5EbsgVhbdon1pXlMy6itGnsU9sUB
7QSL3hDr6I4Un+d87XKeHcptHogR0TrXsATaF7vwveJ0PBa6wuUJ1xLDi6u2tT6Z1vx/4M0/TT/i
0ut9AS+LwvcaXHEuH3OxE6FoyzOvA4V9X6XZk1Bmqgl7CQ2UjtUpVJBnKvFR8W1ZN6G6K8wiSA4K
1JxOglMOsnOVNm8EJlCzialKL5ONEJlqz3kr//wvBMqcmWBqto74hw2SIWmRHPNhz88h71CtBuVO
QmefbqIzT+a8U+kzB2kpEXT02L9Q/EBBfIJx77VCxer9j8bY/kE2TofLKf6GdNonAMpXkkz7Tkho
Fvi6nrGUSfCcKrr7/bSG5/SiL/cqnFGSrwohuKpCxsEQTG+rcvqQE3BBsh9V+4zCaMOEahc2xITp
tGlyEps4JDbFKTCZ81GL14TEY2FO/jqMykhNdwiXvimQpOupPLz+FJdRIfXLdGS1rM8/GrmIKI59
gG3LvNKbO87c1OtmigR2rSL/b9pvdHCxiX3N1YuvqooFk/I71dpiS3APr3q2lkpY6NC+/dF93HeZ
RPxiQuRrwUe7kplcOihK2aos4ODXTvwToqLuLOphfFyn5HWNC3Ll6hXYyQC60hMSdCTlvLljnu/0
b6uNDAdZvgxaKZVWzaULbAfUD8kTxa5gI4Hc2wHY8RkPfaOHo6j/fpW0k1tgbq+2rTgzSXaEfDnl
TMHcGWvl9hOlKdvKV1KSt2IYgy8t7Oy4WSMYdBNcopLt0ZST38qrZ0AsYv36oP1KtSmI+wEdqLVd
oRqirbl4ra98QiAMDLK3w0gqrdZznL/O1qVVG4grrA/Nc9UGiQ6KiSVPLmZfBabk+l329GTMIdap
VS+YpC8TV9II37IvnoB7i2obVuf+Cpwu8yIVc0V0eCjrWfuO3CuYpYY1WSdG+NnSnL/bQxyhXXeO
B2zWCsiZZ2wfXDj07SZ/gKNvA+RaqWr+nuNUrZjXT4+pE1My90ITZ6Jm4g0jfzF6fNb2o8AAwgro
SRFJGHlkeX42y8Obp+iEQbTHc001sjpRmNGHViEAhx1S2ZYp7jCBIjMAQzgVLpC6fCCDeuUiRi2S
2BRwKlHd2K0amZynCikt0XnGEiV1vZ0Ahy+XTDlrPJFiQcgewxkXjJVOdCSQT1+zDjhf3+aWRwww
BEV3wodsQGDdeNdSgf0FfqMgeh0l3coh++xsKi6wgKZqX2SZ6r9BYN+0yjzY1BjWeP7fGM1B1gAa
TqbJ31sJtis8fGDm0K7+2RERQ0+SVWTAo+SNDQYlNB2wOvU9l67X5+H34jNiIyYeaaxVlTA2rP5b
lce4yXTxstS000UF99lxwmBnTskm66n80zbpN4usGYW0jvKIjlSCL8UWeE4Qe1BBdQC3Gbs7hs/W
SnkRidSl79iBdGDCghXfU1f6t5joV74xpPbJhBj/BqMbSwvxBML0oqBQU8bcxT8g4jkJJznabL0D
nHbgN3od1b/YS1RxQZEzYJGhG4vGaeSz8HPnWlMascbsWcZsQiWLFxKe10leqAM35w7LWqjDvcd9
7vZLEGQgRX3LA4ZYQKATxjMc8+iiiTq2So8oqsaveKsrSY1DtVZp16fHcFczFZfujFWjagNqsSuL
2IpXjo0WaNONakva6XFr2mf1rEogLVOdIJTghrltd6VJ3bDHCNBptkFKpAH2O8CDT0l9Mk410GM4
fptdg8xy01S/cZQ05Wv5hXjoj1Yer5E8XxuPt6PXFvWdj1cYuNqHS/PYEAY96ubrpg1UHXqrkWh7
FBFoEzfAQ58dsMfZpcjFqMvggBVsAQk5E2AkWrOZSK/fOiSSX/t+HOshW0POIxs5nk9fOuIqMsyj
Sx4LHIE9q8O37wgNBmd01nHrCm6/SXdas13gLr8mDW74m0tX+bxVUSdm22K9O19LEQewuZy6iSpY
1ljo0b6vXRYb9HIow16hczRFHZes8Yv5mrHIc11bZz4NUOEP8eQHfIGAYb10pMQ0ln0Fd5FKUU54
TYwkK/b/d/MDLtRqA3ZX1zUBXaRpgP68pSYl2rRhS3r2pY1+gF4cCWc3rD1oA5cE+tS48eLazpds
tZodG+4zTOZm9ZCTF8lDCyycV+HWcBrqy3Mfr72DBOEABfjrmxrXGUxbI6ep5O5+af35aCDviE0h
7CJacIvvgozJEQNlRdkPwS/ISLzsyJW/qW1nzLFsip/J5bPIJAKiXpj//xQfyHyf/KCaEdp5/EMJ
LTukr6sexp3ew81EFFpcFC+6U3TMR8gaGLZ+Qu54Gv5lKD0DNYO17qzJDrGXBtsAw9YOmYI1Y+dd
5dxt8bEhY1Y1WI0nqCHCsYL9ZrU5OfV0frbceyj3ygi9A+xPUtVXEoZkivOW+x6PBvlU73M2ex02
A5nZTqQJxKfCNEDExrtFSjipnCZd2nYO0VqRf0p9IK4lk0nbXaWaVNjE4Rj0vMrdkeO4P98KfZ61
Jzcd5J/FMBbRsO4eeowjp5KwbLNFWf6n53y5p2AHxYvqLY0Jw5GDr0pCoOIBzfa53Qys/D3DbhCE
Mt22U8vYN3LVgGrypPJy7DFpEvjTqZODJ8TKcI2rJiZThT2h5a9QYYvHe+ypeIWyAu2rfg771eGA
L2KYwn4VunZZtYiIuSE5H27PMyR1GITIE/uiw6djwInO5R8vM79NbE8EcUYMuZE1qlPwrkP2r3YH
bnGSECqm6g3pVKRnxRvJ1Y9XfCsj5dTVchzZfnBc2+RYE4ZQ5pTWArr4K7TpmsXOcuFesBbep42b
MY5tYsN2Z4145ZPKr4sw5h4xAkemXtyMpm6Fy0Ghd8O27L4eWFa6UVXSGZjtXFptWWgvriqeLuFP
EMhVHBLxYSn6vzmcPjpJKGIok3E7AErqztnXmDj5IXHit6WDRsySwuEFtg7mn0tIiY6cY4ywGD18
/K5znZlDmxI+eishFzTEl2OUL0Jo+TWhA6kiJhcAKm5qlEscyySWR+5/vAgUKJNosQJo1e2j10iK
cMNyWFFOF5a1/PqQ93+Ln9bhZjzooS0pEiqkgVLbTJt5q6X9tp48eYMw8yuMpD+CXnvw18u+JxWz
ptQtz7Qeg+0m5+9qAHRWuly15rH0vbPOKRNJb/4x/zvnUNC/OmgGGaEatJ12BNzhQjX5IcPXxQuG
2LRoWDVPGoWqyRq7XXVg8S4JJiRt2wftOGUPSebFwUyJBCecb4FZ09DMypZ2KDl3z8Y83KKaCQTp
e9W1Vu8aX3BNQbODhNAD3vNXAU4ZwdRv3FS7BnqdLVTVlJOB40KQUEJODgyj2Q1fAytPqaehyH4N
5pFxZOgFlclkwLONhG+C0kNnxfRjznSBar2fIYMtkTRCkLo+ODvsORc44lCG5uiwfBAi3Unyqjz4
zCnGFDNfpjkZsPLlONtr5GduU7NL8rQgn9mq2lrltK0XBye07AQxpuI24ZstjrJe9HLEpOT9EoyN
DNtKCWuAsXWP/fQYOwg05trGL2OkVOdi4UbZVLmUK1pnpA2lIid9QXejThCvy1r1NtIusqraXGQT
zPsfUO0BVIPjoqrDQzqLgnf6k5z+3SDFcsTNbYRPVGeaYMheMXN4SHVQK/t32S0tZCL0BXOe7sGH
2EzW03oJJvzO3HOki+Z2TMfsTlOEx+HzjV5ZD6WODKVjGdGc6nAny2On5IPJbXQZ13oHMsKpu3Us
YMRFdP9KcRy1Wl9W9C17R6jdrQwlzhhQvKxgvYnYQzT58FQ0lQOBcvPiJoCvP0s0QYRuLepvIm9M
8ajLi+312oaTMp7euOlA4BxE2trJ+yxMi/rnhXdOzLTD7cCG7CSDQSsQDweFFxyraUW2Z6WltRkO
qM9HXMStIKSZkKNXlt7t+LjlMJ71wvvnCRkTlxWFd3GJdQs1leVzh09pVvGjW1umvkuKR6JlN//e
O3Vlkwl3DXh0tqPKoG6KHajstHgJ/Fq8TL81YHbXgqKMfwH+ch6RA1o5Kzr/6WnEIicYDphiGWwH
2fE6G1pbU4L2XxQvtEjbH38w3e+KxECeu+wOttPhdIYh3hA5JRt3uNf6mSjd2vHKWO7I/AhIi/hK
6tv1iPz1tWOnXONCsoBPEQ8b3uaG6nIzuurHvChVdlsXWy65Z0n3HoZd/4Qmj/SnhKK5hHWVZKYz
gqiTHuyFRHOgowRrXRkSHDJB2sLkTfXE0KWNToKmYJSgDJjY3SeSrIFkDLyCPu7sF2L3ru21G7jA
ZLCKWXY95wMF8saSqt1xKk1gXPoQ1Msq/9bV6JcaC2MaJttAbZlslQQ5eWTIRz1sPmgAzT2pRcMR
T6Dp5w902UNmyoHhHjLGKwmRfY45gxj1KJLoGsFOFV9a+OtnupSi9DtxZl0h7R06JYErv0bdjeiS
N8G6I6q0lfeclkyURWJHW3oj4BAdtyT1kegvF6CbucH0EXyIpCCVLaWXuxIP7ps4W0EAz0diVvIW
VP7M9GLM0zvvUMUInhduX0KHMuzOs880OqubyfGGUf4FUi1qSUjPvttCbryfuZOxl7ZJoXqiFQG6
oY8NzqyiidMlyTVYx19rBwo18utzsFFghrDCaS4DFBMGq6fnAslcT1poWuvp77lY5PekaA01Y6Cd
xrdQ90m7g0CuLx05Dh5SLwuEvTSHJluWzQ5cEI7YtZAgr4hNHThO3jq9K/ar5qXxWvuIxrACb98h
FoUTAarCFONV2PSmUr+H6WSLRloDQhZpXXb+DtdxYYCup6f6LwKT0u60iT6aOUJiWkMHlpJ5+FWU
sBwHYTF3xdUTHPTHAS+rkk8seNtIevPg0UzASqQyti+YKOUSqHQuO56ZrIKx7Fcha586c9miQ+Iw
JOba5tE8+Kq89nBRb6ik53g7GkK7GueURKJlpCcCR/5tREVu/RrDHwEFdgH8Ngd7IkpJvPyd2RqQ
occ8Dhz3XuO8qPKMFInP/snYlDsPpl6pXRFwoKUTEcHgxcU+b7StXJ/FdToEUxoW9bDheJAALNLe
tKZBHysh7AyvsePE2t3yx9BP8+NQxP7ztwEWFtzEl09MErX1hBCekF28CnppYfEAe1oAAMYCbp3G
KRXET0SOD7d7eBJWbOeIvwUKEaVw/khCJ8FOEjzIJMnOe3j0ddpl39+8Mp2KT/gdvz65had0qlJ6
KpfQB8mvHNgmshADIITFLbTaXJ8Olk+rCPJMoKUG58YhzRTZi8/xRF+Ws0fejEF6hLRhybCXfCrh
co0oUziWIP+IY9aWBDtP3yJ43D+6VOYgk1BJNh76TVZG2jWNC4byMJvO1tjITL1ljUaA8+vIpTVd
PtetUfyTtxvOPGniWlq3fe1x/WmrR3VIQjPoH3RUhluwiDs4179v2y9VQ1tquKzNPa9Vy+0O0iex
0frgYdqrbK0xmz4WosvjP2D1jkNY8/09d3cnTFQ2tj2ziQKgr1EVGsskTFERHguVjuiGi7j2tdt7
mo4SKtX47CslnC0B4ujIj4KJF3YF1SviL/ViTX3fdAjSkSbhFW8/loF77+qKFZ080gwId+nzDP6h
0xNvd9qyAmX7r9rz4Um2X/tPl0vCUD4vSV5JMKpkh3ZhpcSzopvaJ/ZV9fklW1Jp+FYWn0ClpZMh
7rSmUOh/WJlXw19aqo1MnebvRAXP4Iu4Z4cljkz/ew3SuXy4gJPLziRJih7WbekFh3mSS7ZJQmJM
GFj0irrzUncG+3cQnxv+286r/o3Gm5JAifF++apmcHxik33npgu9ym1qEIsCIZ54fdq8VrMUmbix
BqcX39uTqHH0B1E/2VVQR6jMrn1QkVq2mFkkMZhv7xBqb+ju1KCXolGX+SiwNARaXsTV7vTk1ehq
aw+Q7xwdP/8ReAUDJLYezhl95+XK4xggmfam+HRckCAGtgC9GZiwpADNyg7Kv+xBGujFZnV6MZ6C
5xJQveleG3Ym+WroDk+yAXACAn54dtF9wLWgxhSDM6QIItVnf+FydzYupm7MX39/eTk+fF6sxX+D
Cun1sJHma0QHBOAW/s+vaSAhIiZQ1H1PqaGuAAefrQFI5KI7tySwIfjuTKPNAEJ07ChHt4+G6gO3
MRXobGQ+j7c90kBubBKnNPSXnzz0csKD5H94BFiMMD0tf4jqbdMRUpHEQ/HBKFJxDivS8oQT0cZN
Ezbt01yRmFO9Ti8TtLnYuCGgDHmCbDRK00OHKlDqaJv2Vf8fBrgkcMKzCoVisTTi9JgiZGNOC8Kp
XcD+rwvJic79ndVFPG4aDKkwHbWfbx3m8lCX2QcALPmt/CXbwZ2/uHdg07QD4paaIb1L0ChqaDoI
YmVf4+O3Z/krSWLMdsHXm8SbzRXsrcoFqE+iAv8L4q6uP8EyfI/S6n4JUzmkgQGe750YP9Zec8DV
YO6XCvTl9Juq/UdcwWqTVI9n94VU7wXH6kGc3zwj+QtQ3F0cU2itEtbj1UvuU/6eTEgx26BK4AHc
1HDJzbG7gkqqVsc4gpkq/09XuVFou+JETVM9R0WMjwuyhoOMZQu087t7LRfp+VXRHZuZZB0H5z7q
S9FwSRCi/Tu38Z/GV7J0tXVPUYO067eGHGX+Xg3mxX7IFrGNW24d0ProWg3syDmu9xOgM75fuzsZ
CoVleS70O99ynMMG2QxvUdxZUfjjza6aiI/hCWYY5ZZyq+cdeI6gAHrekrPngxkAr1IGszsegmDX
WPo1DcFkSckVfKqDIbbZRXlpgqpE0w/Ii28kyjUbusncQGBmT4/WpVtLtstP+DzvN4QKkWaEp8ST
8yicSNijYJMdsgA6kG9n6JV+f9saxa7BZI+LzKxGS2xBB8fZUhs18lWzoORB6amp0oX6hleGuner
sK2IAWZQsaNuwssk+W3U8vbMfBcC7PLK5+W5HsXdL4rps5YvDzg97csR4xB74cGjWAA1d3YM+9os
iHt0TZscpRzf0NlngLQt03FspvQiF8YOqATEjiPv2D7teXLpvVasU6e8begOmtHQTXB/mp1P1WEp
B62WHphLQrRidsCzPDr6fb49OcENiglzOjJv7VvRMMGHL5gLlZ5d9Ixei5LEgjXdvvw5FKYwKwGf
XtLxLMN3QBnKwEDZFgHdozuLHqnjEj5h7qw9MdMlMydA9tM3H+koldjmlorDy7gDWdePxPl+zqtf
xrAspje5MP8kxjKe09+UWx173l2Z7SloLIPQrevXXAz7kc1nTB1doCUz3vH2okzzD2mFBRDEVXFi
0ZgQySIObmbqGYf+Yc8OVLRYvUmllbUWgKqJA4csoGg7iYGX0fKgktHpfzK6leTbv/a3QIAmO0KG
W+JKLhW+BYn7AXYqyh1aEkEiVDHEwYFV+5VqB4EqsyaWeraTKqq6ErUw54QShbNgA/OT337wGzlo
fThQfkXWDrB/PIVd0DvfkWNkDUh3L8ClmX2JviVkU+HdBgwDSDboqJijVh5qfQU6cReiQ69RK02A
IkNpymARTWeEyGjZPGEHZnq7MqEx87JYPURJySPhvK7WxPZATNjCLbZHhTeaz43LWrh7p6kzH11H
pTAr4bAcSZmIrfpMnSWR5fsaMnFh9aSbP9jPwy4KW+p8GEjkdf56PSRfW+kosr9zIO0UnAj2NoQs
ByIbPlYXtCWSSx5hJkuW1tTK1bYNufJwWYnEG1iVrxOq2tvHayoJOse1PQcW6vJX9d01lpaiFhgh
u5Nbju+f+YQ8bfUHv9WVlfrSsd6TZtLMF+Ft+XljhHO6AC2Za9Z3RQgw9N/4sxobIe8ZM/eJwBbS
CmE/BR0gltWm13C/h+yLisXRoHqcwO7HXcqIKEx/mmaWnzQm5OxMqhUfvWn9MHwupJXEDsjEsLcv
Eco9QOHWceRDKQrWMeP6wODxVc6NBHekKj+66w6bECLgt/ZJhLLqhS0ElqY3gShdP9ZxWd6zfcvX
+QFc4/KhU7aCjULJNOM1079mW/YajkJp5Wsx2mTiLhl6MvQuwi9I1kpwxZ7APUQECIkLWBTw8qdl
LsqsZDTp5CCaha8uex2N2mO3iAI1YMRPP/iIXtDEtbM545+9SmKjp+kcEHDfCF/3BAsdyaWgMIt/
5u2soH6ctcycCZ1HSblVM2QV2L0EEZW1Gah3/mQptGJdijkLM18u3hARvdkPvN/GcH4zaLrU7AS0
SnjOkyp6hOOPqnvD4R0bkdoSWZPqUNwkscqymzgjJi5e7Pot/QPz/a+woE49Ll2Z2cq+uCH0qw0U
8R4tAVb3GFjRycDdqV/iqptQIF0LO2tclxa+RJlwsqpm8F67FO0TdjljHmYPUzlwxDewCEZ4pMxi
zydhL3fyJb7Owja2pOSUqtujM3NEggEh3aDKnyRPl1QXBIxqEgh/hXnOK1q6YcsbmxHHDzfGgNCT
iVwdFiNby/E0knZ/NR+VsNFA58Y8/QyqZiyEO7g/XEEWKGb5BzG9OQ/8J4vLlxzNeKjYXT6kJlv8
nyS9G2fNXYxdA2orrT/4MQLdFZJWp8W9FGHG4x/ngiLu0f6r6KxqKtNw7gK1bp5VKfNUcC1uZ5nf
KcbC3k6pPJFnQA3ZJD4tgN2mkcu2T6mZ37+mFkVLbakeUu+i6+F1sFTovTgc1EEMMcf6HGUDL7vl
Qg6COMX8m8GrMC5fJ1zC1pGgzG4SOvliEfRnPktmdk5ZevfMJFMvJ1W3DhfXEXU0ypxdHHBN1djp
PPWIX9s3Nu+uoubP9Rfe8xw8spcU2YutWJeYzWGrFwJ/wvykM2QLmTkBpWSe+IEG34zx6uBzsIIv
N+BDxxZNa3xiPCHYwixgKYiOANYLTEaRLYdWz89jUHwx8whmoCXjun1gWU98icvNM9kCzJmbf9VP
P6GIG2UG3eqqluJaJnXAFThCOWsAEOfTpiWCcAlJlFTdylQcAbRteuZ/D0i8N05u3IU3Ftv6Ynhq
L+qhVWU7wc0Ko5mLInrtd9kXJBSnuQwLjgtiYXEtyeER9w/w1JS/m66J25Pp0Z5QRanh4ShZnE0J
Yp/XWRt51sPyWNQy43GVrH/cWvqwR3VZZnPg7gyDShWwWmzPgSizUIdvVtMyw9aK7wlyHo5kzEpj
//+K4LljyHJQg4aNp+qXSJuxAenn9ABfzNLZycWUp+Xop4NiP1O1S5GFoJcpitbP+AenmgtqlZzT
Eujt4ethso8BNZVrM5pqGpm/MjT/5aGRTo5PW+vtNu3caNKNlVL6TYnYxQtOWm0sbcGSCaLMGtLz
4/ePzMs37dOj11zqOQ93ajgzZ0lMQ+2r8L9u8GSZz8pjoiZEYkkm+Nzzy1Pagb/CJoJpRnvkcRkk
P/Y548bWAdE2dx2T6hf8Jeoe9f0ULfCFbnVlw+kykShkyJ3W21Ep1e7OZAujFT+UBKjWGI0JXmop
PL3II106ct0/Sp/hA9ZPRhcCX0f13Cer+Jxb9QJZ9q78KYCPhKobRPpzv3RwwJa23f/lN8GX+AKy
mwsRWWU1NdYfllVHTrWhiL5FIuOppJ4GPWAKESqKlu4J78RgeOUfVwaBMIocJ1YM6uppmaKc1R6z
3QV+LJ/B/f91JGktD9lvIHTQyRSs0ZpZlMIVTdh8R8kSXhlvIUhmeXaN1ZmFXKPnYFGhHb3YPg4I
vyrVOvCzVDj4yyZ6yKReso4Bgza1PcyjOvR7Ckr5DwsIrGC46eOU6hurIIo86WCawMR18y36F/yn
fgrg/NG9SiSRyn/WzwM2ZzZln0rPwnammCUn+HuH3h3MbZlZ9wv98CmxnPpLGX2y4/0wR849txs4
6mSJLqYOMU+MoRA9xp0Ac71gIM079wXjoYtiAMbGXFGK+Pc9l0xyR1BwKRL3wMuisN152jPQFx83
gIyClce5g8aWtJXjOYUsstD2kABm4XxGw4ZZTQ5uYQZ/gqgCNW/Lpj2Bi8RLvoXsmj4lpCOWgXhG
B6yqseI7q/LzX9ZrPX/lWpZEWvbFR6w4+b+nwHdQ/FuF6QS75uoTRDhTyKe3heXmrqH2ZvZDxkoe
ZmFIXA9qt1FWpDX79DUWRYqZPiEiyzddMWEjpBTVifzxMT4bKSipzbwF4DFg8a2Iu70pgo8rORkH
u+LuYflcW5v7iDe+xXyUqRpWtW0y+w+Mt5QGWGMdZWU3jU45TOYWnFiTQ+k9jGIieEcSqPh4qmFl
fhNE7Zwfo1ALsQ82dOckTbw6Y2Uf8/61poDYHiE/EN3HQf68sL63zWjgkQ6oGuqBezWWRiGyAmST
fZ1DUHnX+Hb6q/iWLYQhoC2Gpxf4qOyVPgdZnLAHAMVa5ybDI3d82WQx7E7s5M/v9/lOWPyQ879Q
Q76sh5PL58ZFdH6tt1EDfPt05HUvxfXkzMipqBinklK0MmIIFeVyNYNz2FhHdpraqSIT2IKrn9hl
DjUJVsaprdH6nUF/X39HOf1L9dqWilpSy9+14BxLRbhcdvh0r32dh+tvI1bIFNbQJ+nX5JkrNOHk
fCTxUuFi/ox83AdtZN2pYa5/ST7QN+jeg7L2zAeif24+JVffK1+cLH5hV8ZE37YDi4mIUzE0XOfg
6sEAz+Uk91kxkNafUZiZ7JlMW0mW2P/hh7UNsQZ/rLIcp2hOaFIb+vb/bMJ9zJ/yHupcnrLu9+JV
TdZ0/gz+02ljV/F5ZKOG8zIHoepvylRTXChtm/qxIg8ZLU6kccOKeShwf1UbYZQpDwrUWKiWiJ1X
MiXnq/kv7q4oeHDDJkN2/nd/NPSYXmmXfbdYC/mEa804Yxy+Z3HshKEs72HyGwaPZWu/CXmByzwX
6Q+Mj+ZabELwh8KcJxKhWc2TrJMljKjQsmYQtKdAFbh09vxPANTODbJHZXx4o2cNCYrKLVTb7+jl
GZsrPyZU4tSVVuqi03eP0aLPLLdgm3HvOFhZWuxjmupnpbTZVW7xWRjbyGLT7aHa3y9AiOxsHfhT
VqyayoYypOrShF8/rF8hpI+QH+60YE7Lx+jaufPXn0cJyvPNqV3xNepv3alUnsNZ5ay2DS1IunjW
992xbBXQTS0wkUDClZiU0VUk+ZA1ZO5L9b8CEN7oSp83NK4edQ9Sj9stSYc2iy848VDqAct76Yp6
WqQQqTgK+ugThG5/P6gk4/CBvERZsOfH4F2ah87rwpCB4Det5Ulua9tF1wP/LyhYhxDC4i3rJacq
rD0x+fHQl8I5EkthDEqRyBT41TETmzuOsH5jU29lJd3rkbQSEAoE9Kpljd2dZr9i2XmEFJPjW4J2
457QbKBxS7niQsDAbbd1bU3TjZRPJVD2eB8FLgL3w/znEJnTNhNeC5OVD/ub+Nn1MuOtdwszdTxx
kKc9GbAp7lJbOq6LDg0TtEE5wbCDQuqEchD7MMcoTWnIe7Phy4N/McU2iV7pDDkvNcr/u/PPQPQe
PwwYsn2tTpOvJEH1Kyw0jwmBwOSsmqUOwFMQPFFDENT9fCmWctIG914KDEqRNQTItFZanVaj2CyN
Q02SnWJBoSgo8aeQWaX+ihZ4Jon+47jrTL/itzUjxfSvM5njnDs28/2hN1WpJ3hSZwOZqDAJV/p4
2UCyBclJVGrbrKTXD99FjIvI1StDv8lVSe4xVus0/7gxUh2J1f5NmZYIedeUwGgOmuqEWS0wBkNX
5kL1npW0DAb11AQ3fi6yvzyX09ufbjaa/X6KjVvou+8XvIHl8YCfKiXs8N5Z9MW8DJM+OWbKdT+k
bOR/S7tLMjSRqfHm7HPIgHTnxTflDQlwu77uWXRmPi48SUkgtN6elIY+b650apJlKVgUciXMCUqT
neZWXI06WrRU6n+kiPGB9bYnlDFaznXK1BOR1OOkdc6mm8cTh8OQ7LIz1/BMNMEa8F/CShNL5nGW
7XjrsGrrpjERq0f1UVoXYmMzKNLoCDmxk1dPO/oist6mcKL/YYhdcHuGS8prmTNQcey6o9oP2QJs
1yjteJ2/xugIwQ0MIwSyyEJlwz/BEMYeRHvi8lEOkGxKwrbxZfX/Gc14pS9yLXDOiFW7c+Yo3Fg3
aScWAgKNGFsWYnk8HerfI0DeGOno0Br1dWrsBRYiH6A3IdTEHEikWyjrr2CzS9T+UFfLR5dqdkrW
t1jSwMbhVCorT9FnBSe/7LKRajsAvcZmEJihhpAJnFnNNKgVAYKcpDBG9kpSyu7QKK0AtQ7entgR
UuVZNF9pjl6v1GWT8yZArc2fcgmZQK4DtKoxDNWJ/UgHQM41zCBrjQqpHqBYww2ye6rQbQwc0vGl
VY0XWvZvU8TYr65yYEv8nW5F9bqN1kSsqywlqTv9hpeAjVN2gdvxxGh8rbZYWPUBNdBavPoj5nGf
7EzGbGExdHRwAjWHcBUVRpgTKAB+hbTM5ClMnmy2akIO8VwMiUCc7HhmwYXpVkswV/ad3+AmSQpb
zs/yPvNf9aNI3CybtHnfVPD5V1pQy+Xh/1pjbgJjJwrRnnhOzLc5EoIoSlhKz7vOM+HZMqdq1Jm4
Q3wT7sFdYb7qcGUpZPLAUplzoJo+A7eO1XF2g7aMX40S4FclI2XxqnEgn9graDaTsLRly4/0SvQ5
CTOyHG4XPsgk1O1b0zHKpxJ9ZyXQHoBx9UvVavOiGBEAEDdpaHDV0T64ubOJXr+01nFe0chXxSpr
NhgbBEp2vyK+MVIo1P8k2u/4SwkrRHx7RDtZTH0aJEYYgGhnvimurjhln6n1ZHk4Lno6+Sdf24yr
jgaxQKgw8z+/LVEGQ8NrJp3GaYZb3+sEiRiUnNqDB8vafWMbZqOpkxinBeCMJ9xzUXW26oekRC4U
uxRVtZiLn3mS2nQLwGC8EE1Nk12gL2CFJTjXHGygeMgQYEi+AU435CjPNDYyphKEpRo2etRpKU1h
pCRb+Bt3VlBpkUqV9C6/1B1tYQjv6KbBkKYEDaqv+Mcu+NU5zrPoXyYxb+l/81m8mhHWXPBJxC6p
8w4o/CMpYDFPPMnSfZ9EaVHj4vbf3FM/mp9wSjnfiv2/ndI6bSlkM4BTPsPkIJgp6q062o5hlQb4
PTOlsTpg5XhsnPDlFU2//+XHCRBUDpHfW9Ki6GlHzHe1ViMQuY6V5zMvKg7g+3YFAWuBpjhePnMu
Y4CY1eu4XYO1oIerEfnhTmd6OpjX0/3SDzFJRYNoZUOxGBwUmno0tNF2lx5A31yom9yrOJWkW75L
yh+N6aoYkodiPREDrgneGbqScdktnivB+e4aJuscGb1SjH2njrGHUoF2bvYmQkEzaDn9SYrbK5mi
fXcsaOu5CWIfuElOYL7QkMa/aMxzCJjMZVriuuTF5Wo4a1XUviAgqL4Uh378CWbBCYVdnbltHmEe
ndsOXAEs2QGyZoYlJXxxf/RIV07EsI+RbU3+MAUVE3BRBpJbtBuXGdsYpryTFIsPrd2eLIfOOI1A
hSmngEgnkZPm5D4RBxEI2hDv6Wf0QCXFbNeQXOVkaDxu2NPRnF0gr0Xw2/CFFMaHTX+QrA4FAzYT
XN/ZvvTriQyXRbwTIuT8gAM3BxBpsnd+2j+EvPkQwZf9CTaL972Fb1tyg7c/Bc565pLOV4H+7B9c
/51UqupXtZoJZUdf1tYUBGLethYZd+8yuQtULVTYJhHS5gNQZpxxM4N5btbU8899XIOp6jRXt9nY
WwAQCwxnjkHFiVrgc2mlQz/cCO9cyPTc7KUclZKo8D3YQ2HHZnyIZ0HkEfVSMhWlmDDlbp7KBYbp
bEXSfShYVOa8XFOLjCRybOr2r9ypKD37mazsBFxS7vKhQyT24BgCBm+wgQlZmw8Y+N/Kb7jv0dBC
BB0iLW2pbAtzD8LV3QzIKobxqZRSEHygNZnV0N97jowbInUDUaZHwI66cU9tAKijwDNegUZztxcl
eddI6ZOeREsDJmM90YXvuSZsq7azrWX8sBFqxZ/QJZ2qOQ2iQPwLhSqyZJX+gALnI+PkVwPb1z39
olrcDygrJfjWNYSjvp8UdkV4gjFjMTRQ0vp2XiaWPaUouItlOfySpDnAbwi8f6toKEpSq4xcVoO7
hFP+TmIHnLg1uJktHewPEwThaQyuaIxbMKF2vYfr/Q3L/P0EmVO3XJ1kJkLMri/t24Zr0UjYlWny
b/5sjbhSbDafMVFUitKhUJar552swzOyMnZy7fYpOO+iGmGRhb2TgVwK3Gv+feqtMBGFtDM3hR28
WF8t3XtSvPS+FREGgcknL5yRHAVJJoNvEwBsVznOjBaGn+erWdvIhJ244NtIcDD5UvzwzUn5TyJR
JCJeaGGpax8zD/8cGNbh2yuZXXI5ILnm6mTNkfyXCecAKwWMUZxEQ2KNvC6E6Xcm8FceG/tu+b1e
zw2dpPEHLqXYPyEEM7K1/lRtJ+1Ih9pHJAnvmhTLaR9ux/NFuq4rAdQP6nMTKE4+IobbDvZtwykB
PLA6/8ZOjCYPpUjrdxuvV131LD7agfFJZoAk5wzTmeirX/eqgb4jLoUY6W7BHZUD7yyfDPUc8LD0
xP4IATRTP+/cC5Iat1aUyNCUHCURb7xAZRUl5kGPsj+cr/OmlK2oH75J58TgDtnOf2eh99FiLxuj
plggRtdkZjSK3KJgARWofylR9D+lCIkXuLsT1qeJ23nB7MugRUIhfq63nSFLgTdAiQNSsqZ0LUEi
6sGxTbn07LqMo9u//X1Yl3UJUla5YXmtEbkeXAuQP+l8WA9X3TjcDJiMMkGgEdqcdOD8pj2TIXsl
BmdvLcbEI9tww7pY9tfgOnhFk2IjAHV0bj+/4Uds3lOoMjQIYmCVnEyAMYvGS4cVYp5sRRAa3KJO
pX30OUUZ+DTZMhcBLLRGwSyCQnEcxRZnpM6Urq0ukBf4QBf/RrZ5tg4Vz+FVlCqvn1iR7XX9f4ta
kFCBFY73B3pA5okZkGbk/vZJG7t+BPPQoTt8tSqW1B4Cml0ocsY6YVYJq2F8RDpn1DppRplvAHQ/
R80S05L8cXF7ne9TAZ9RVZbWow8bHnfAqFEQgOZQ6zix8taRGL38MUJ05l3zBeBw6jkNj3T99C1E
W/C7+35PuMo/CM3p35ULGNiIKX8mIyqqEdZT0PaC9id0J4BGHsvInghsCwNnS/uR9RbLIKptNJAz
ch+Xt20DngFR+uBYFce9GoBzC2wc+85X8tBZaWN+3DpPdzP2l++GOgp1VVGETyypkkryrEjvXwIl
1K6aMX47FVzUaFbAZ8KODooiO+WqDLFOFL+h+VmJ84mhVNNCodho4A0lWXLBR9WtMC4dr0y0UONY
Yjmprkun4qaQbP1jfe8rO6O81xDwhT+Ygmn1qvAoDksAnTzKEdJH6Dg/q1CN7safVQBcg9FignL5
maSIlfJ2T1/EpYzlusz/RvCrI8aX7x8pHFmQqRIeJesgqoLzwqDDhQ7bDsHXt+FoF8rkI6Sb7X7R
rIzi7jHtv5NzLPITU5hK3Xa7k+L0r38GCuzLO9aMEecX5Z/qK+oo/h4IFQ6OqYcKNeHwuqWDNSED
obJZeGSaHiQ3b7Aph5IE081Hc1QZik3yiWqYCwtJWNzpMI6GsVKYhfwKE2FVonDAzTU3aV/foJ3f
UJceP2n0TmpoxEk545B7jXdyP9CovP3Yv7hnchYKr0j2qm8qe/tNVJ6edAfbGuXjsSQNIRnh2Jz7
9YYauYy95QQx7U3pTCW39L1uScPfs1aZfD2c1V59n4GAKM3V5C1ZSLveePe54ZeENQvbT3W2N3+l
XmdFY1esVpt9pLmQAPIVWGHDHqIbsBY/JRzUDWUogykDTcqFFPCwBC21HEUhMsU0McxY9NhmQnoL
UPgcRq7jJtnKlk2l9f8eKz8vDO3qthz/IZI4dz5Sg17jpki6wAVhKoMY4ZPWrsFgLutJi4DDRMNs
YWFezPS9CELYfphZT4DbWLCID9A9C7V1r0BXU9Dhs8CAeWKB4vIP3cwEl5ljR5eHHX0TBi2IdF92
Tv0rXWIWWwZT2Okt2wadiSb8TH+UFYvn+ZOYgq2xqsRDG3pRvGcGRpPFPRZRVJHLHqAbnu5OgngJ
iBx0sPSngvvp2iMNeX2YnvYAPCVnEmfcQtPREVNnGPZiIjXgP4/BDQ27jYDmfSlS+wvjqY1r28Wv
qA/klQPuhRzwMDXZ+xkJCoikwTrIRfbSmblNi7DAbOXEX/DKmrDI+jXF4aE3g2oCjmJezGEYVFUm
YbLxv+YmInSQiYjzLMYvbN4t8YWm7bSYjFJtni4IIXFYnx7Wnu2ofUl7XmJZe5I2ohuOfxePRFGh
uvnLzJzmnqmTZza7bmjnOrCjEwLuaeTZlCHt+v0ulyCESv87bIZB617dCKc+2fEWAa7PHUIR6GiO
OiM5p1RPCVE8BCQSgA5gNlp1oydpi2s51jblOL1zGKfPUrGY0CAxNK/LQtGnA5aD6GBHNGPJRw++
fk6OxwpBEx+47FaFr4w9XbMpwz44u09MP8f+jzIQ8F7t8SXHVji/T+GlCA+kFOP/Pww7DEW7Ne82
R8RR8sDNMxUe/RLqKKOz02FtXrf99aWFPF2xj81Inlqw7vxBU2wphP5nTdXb7QtqhfseHuEQiopd
Rn2ITl8q4wpi3AOGtvSax94+lGm9hfKKv2tdA2Mc7jMaa5gXCZVxnlR30IOJINkqTiS253yDQ9l4
+eAQAYEa4bsr5N7MLAm8RixdVPnKPPLrhyDlZWmcaiIE356kMw8+WxjGmo3n/t7Q+I05y7D50ULF
b6V5q2Je57SsYKsXKaPXX02fNePx/1YF/9yGWJv5uWzXQGpdSsykkGkCeENs8i+tU9U4QKLzhLTG
3Bgqrmpyb/2D5EyZSDy/VgISsBafGnQQvF3oqDKs8ZiiWG0j1h1TXUgWsHeusGaNK/WkMZ0w6Tux
ibwuTFi9/Qqc5XdbHVkszWGKtqcV4O3bcNvWQpSWJh+dwrf+82Fg9gvzht4kDfQGF5OeUYzOYi9O
IsyOEpH+B1ulmQ9322CVVpA2Z4ft7U9/fO3oy5qqMCTSzs4+w75F/JTSJxBhhtUw/6HaOI05ypwn
lI347/EPTQrMAS1qPonA3GL45gjZRU/Ae7sUNB5OVTumOAKrYiW9tKEXEfEYRg3SRIbZR5NCN1k2
UaJO3vKD+BhMCMclikuBqkH9dgjXqWDXlR197uv8X95ww4ORuBeWIsry4AXv42E2AZ7EgjWcyVGY
Hw3TtCZ1GZnWMdItAsR+mKSp/6hIzxCinNbbPdcgSt5Ill3CJ5AVGgntHZosnsTuL9VAoq+MYtVL
ZcEL63zsP0fuzGbfPE7YvDmpzjJE+9wV8rdgC6vnBkIkAOSp/VO3CWomJglITSDviFPO/lZOWQ6S
uLM/leb/OCwnVwfMXrBngUAes12f7c6y9QzP+t0PHV4tnHY+is0bXWnPBpPTVABRUaUER0wRsxQK
jHosFAWTQbdawLX88p0AuhrD3W3yYArp8GJVhqHQRXaFwdOoMI+F5KlMM9DvfFF8drIKcj082qcO
+WlSGAT0NUyO585pZ+RodMcbrIz9EIXi2ypdOnyD34bfXBopgmx7ZM9RvGn4VL+Izxr4Z6/EoN+o
pgGsX8R7muyETgPCargpyRhmXIQEmilDzUsnpGXPRgV73K6IJbHTdCpRlyfqfFvwnirPnn3r0HjJ
y4p82xCLAFcSL16EedII6WLCrqOKE+4R7BMUhG1U6QjG8Ka21jNrnaDpqKZ5Ve4RTIhHYc2rbEj9
v/qNpUNoPRS9TWzALofUj4JtUMJS7NIODugYX6v4o5bKw7Fha+Z8i930J8xZvIoUR9HyojCUnbPA
Sci07yMBu0H2cA+ts/rF3QBBLcVNQ6Fjy0PNzBLd1AolOSuYbRYh3FafU1a/psOWFURBB8uUHAsp
nhA1X/l1LwGiheiq4plvhYl/WWvWSLzt3bCJLdBp+9epEptvZDGkGPi0bvWDzP9ZyEelv1F/ufpR
hzRrsMtjHm0l45D0nukD/1gQsi8JOA0NemzoZoISYwUz8LyegEXT6IbYrOVKM9NMNQU4zH+semw6
UeFRarqQxQ6GGsi2Cz6agJ28caMHx8B8o359OD5vWhVddVxL6JMRXjjhRJh4japTeT+97WWYAaed
3KGwEZSk1XhclR0iifaZtndcnU1Mn3qPSVIUGpPHEVoEDDbOZs0bcQyQv7EQ6pzrZIFxrVD6tHm+
GmAOpjglc2rA8CTuLZBXa1DOP+n0jazl02YRAZFWE16LpIUAkWFCYnFxsQSupcemKNSd+wzSIO7p
eckj+0Y7U/30Tykw0NE6OHCSKPR3Ekbv3NRLE+xLsKwycXdHby1r+TG0Eo43Vvl1rEFz5Sg9fjYB
QY0ghbqznIa51KXUeH5q7GluNy6eqiI/ry918cIEcUNIbqDgnAMcnRfHjBJA/yVWCUubOjh9IPCx
nkajfMxepoMUixSKJ0bB/uswYf3mbc9lMQ9eWTVVjTBA5fA1EWNLtGlBtjNNJ9T5QnQ0I7gH0xI8
wc38fWL9Eli4aGRumDxtVr8n517bRFjOgptI4hBWeKchBC9fINcFgRyzKrxvIlKv06Jy8EQ0vrRs
iJ7zJXleYUXZP1C3laaIyEZr6HuLc0R7q2kWDm3br08xLtIY7+h6PREFF9iTvXqp4NMG1D7BCeXr
YYOjy/wgDdK68Tzqtmme4efJ/kbI6QKLE7Ou7MpYC5xnts81IvxVvL/AWOoTPbGSrtIwgCoWGMS0
1C7vYIZMjH802BJKAbq8mJt7ObBtpTi2uZdd1apT00IBSwtDidvBHjngAD1NFgGDxxduORVOsU9w
0J/CiiRdv/iFsQvU4WmZKmUp+2Grte2uClQH60GCWGRbGS48wfjC3OBm3ga192CKeqvwJ9aXRovD
f9lwbi8lRS7NC1nS/90c4TwDqBMbzB0BHJcJfHwrW5v5nCvad+WMyAYlvKgNeRMOCryqswC4FcKV
EVXz/ntRoIGUDq0ArVk7oUgRlfIGGuyWxbUWZ79KKwxvsOqSZmsFH6UrDBGGHlVZmnbZMjLKOe9B
USjGd4b0s491FiHTne17fUOwCK50kJ3ilTpGEHjEA8OwRP31oUWIrxb+FYe/cnE9lN+95iQJfGTo
Ho3bj5KS7FqURUlhQ+noJBGlLQvTmeMYQTQlTpy+PN3aq6Qj2HH498Go8vkde/fOf8oAGzYACl03
1WRNvOF48OEFNpACPkV3jxzAI9tfJC63nPaQID5tSowJYyGoOwp6KWI8anWt9w1bhU/XoXC6aEeP
flFxb/YRQjZnvUUgIYx5F429aVx+y1s4t8JGpkTLvAiQjfGCw4zjYEgu4OWqL1ALsxzWqVSvAMX7
VvKQTdICS2wEInbDq0L/BW8ynip9BYGwe3NscBGrUo3SVnYJjw6qgnE1ED4CTDIU0Ij/Xs1moM+v
JUlhc0nY/NOKvJvlp/2saUzMI8I291LteW0AoX3sxBEZ2vO34iiZ4cwIVyiDH18ErEyQLlyzdlbn
LtPoeijHLRyM+OSNhsIqv2gW3pczUKs7pzEeLvxBlUQB3R9kkdzZjLHu81WcxlFblyI97PUPaCBP
bDgAbKSMOdTvSSGtABc++L8BwwSKq6jhdAaN+KTB8D/IA7BbPTYh8Z6PLdFgXoJ6MSg5ezEZQGQx
apKL70h82UTjKlRDMIkd2IPNMqiLM8rtzzWgWtjfoSl0ZldBHHB2ECLAZJxPGPIQKbLdoCkFqyuq
NVVi0YTN3jD5FhXYvcGeuHkvvNufzRvwYWtMtEMcdCthRpFgv2NTkr4HI8ogxRaPSHwrEWufcP4P
41Jko49xEtLb5b3zrICygIV/Kde+8aHQkau6kNIERFiXrkjWJLxLiJ9OKx7G0mm+M8KYltqTvycb
EHuwEQk7D2NfN2lQMECWam/w+gu4mU2jdA5fnYUhQhuZxL/uI8YHaVT0SvfBfOaWWWHsWg0RmJVF
t/350g+nkRM3874iUL47fmxQTanHU4tBTf6iKoskmdJh0Bu934pwZR41nhbjlTQTgJT0rKvzx3z3
fTp2AJ8g7fjFzEGnRrefRCQ8I6vu+bKPejPKRNcPL+Inuv9ajz6ltcNLqAtONMdc0cEsnYvA/Ix+
vNy+2NIxsQyFcbd2JgLDCMRhSwwwL9ecPbah44WTVMCg8AlhB9iI1owycT708BIGFy9Dqwg+15Yb
CyuanD67G8LSZexHyieaV6njiN1fz0nV+Pvzr4/pIOk6Fl3MJ5DlLTtX2IYq7kPe1a3GFDSlpMU/
JHA7o59qlRl1HiBzoI1sFhzkZ/x8AmC12SDNHQMoBZQUMAU3WRRP6LXKKWlSGmydWB7n90tPKUGu
e3nngkwFr9p7b1zkQAwXw8I5L92a66/KakeruKNEte6VWG5senqpEi3dAPO5RgDpO7lwQrs0hPTD
7xeBJHwGvBHr0Oe6jC8pYY4FRnhxXOSY76+lxJ7EPz8x33jE/pDns/YJfSwj38Z5rppKh/RtkhLh
nIAqZArxwaDkHb0BYcJN+goYxMHx9Uvg+0HQxKwSOmFogfYMRdB6sZ4rXrJnZn3OUq4vxj9hLy7a
cKggDb+KqhJOL+Zh5VPsjQoOHw6rLa5C9hFDBx+Q3MM5EWqGUTKK5IeWdBQgRzN28ClyLgJ7GSEv
aLdRzlwMfNQiccVY6sKwwoLoSRvxoShtYAnBucMEsY1iIlvkt/Uag4F6/45LLiUILz5OAYGCbYLo
gBk6U0PZPs7AxTgHPIdKAolcFLMnppJauFHSgHxDAT17aTtYKRgn0jpTsFzrhxUKz8oNsjzkZILg
Gwe9dvvBTJU8DS5Ci0vYBGRtbzUonZJr8ro0YSvZnXugTmad398zmVRdIQ1YWqU9NYoq64U1YWUp
vVG6JnxExg110jeFzIh3AfQS4sWG1bJdn15jDuVZrAWYjCUUbcEnqNgsMWn+ICZepsBChhwikV96
M1+XfZwit9N8YCwsh13eWiktJsv0YjnsYtSzU+PYVsnDx+w+2RcjzEBGDDJme3RynslvJf6SdxUH
kyYTqWChSD1Kh9T3fgrvpiXWhnh6Xd8Jpqps4rJco+/SE7JGsLL61Jt5M8cnEW2A3SZ4dLIkQ/1d
Zv99cMmZeuMVzoJh35Ge5m8gLHBwnLHEU4Ilj7XIc/YeaXUio7jSoILSI0+1Af1nCyUCeJewG1f/
vmwk76nYMF7yNZFfp7zcC3iHHlkwDeL7690GR0t+P8a9Q+mN9pNBRUOhRFgL2zSRL2Ah8wUxE5iB
a/0Wc2tbdh16E3G5rJ0yzAGY60TQU5L4UqYtzLiAb4O4CKiRIMVbwv/deMECh6yjhrbFYi1UU2ki
NdJ65tcUQ8MOvWPv/EGAMTqBAFEK0epazUMlPLTBsBjaehf2WZgfMfoZy8RFTlozdueLN1fiSUBj
xK+MgmNEzmONnZIEuNJ5T5GKMdd7cqUR49F46Qi5d3TWQFfRvYXF2YSjNG/xhcQ3h9hhOD4ui35N
bR6JY9pxom+YcXY9H3qLsmq7job2EmWzuE76Tklj3pFzRRGCjgY4CGq6t1wN6r5FrKDAVbKtrYWF
oqzkYntcvJXk+sShBZbTkyKSMrxVGX2ykRt9LE5ccTpLofDowQxMU4uhLpQD/e0d25+uFD/LzT+y
EcZEZt7pA/2TYpsnNNET/VamW7zz+xYrSO74OJ43gtGIuYfHzs5McbzdomAdh5Js8j7j7Om780Zy
t7OUkcQUjFJTh96yq88oD07g+BajuJ93IttIIL3OaEdGgr5EMgzjh+JjXSqRcoqB1OCBdM9IJDuw
U+4tqHYPI9QWppkOYSsd7XvvyHfBFa2sWoXGqlCsbkh6EDgC2fijHDU0bkLuN+J25ijH6gCx12Ns
hd7TXVMx/L6EQEllbjJpeFda8GTW5ZnCZ1a5tnD1t4XKp8dwXx+dDLB7xCdce92Pa7TbypBteDZx
Ry468fQfmQD7XjkXMfpQ8k1sEPBQlg4Kn99hdz5I53FCKyHsXjk6MChpCwgvCk/oyVcak6CLUcSG
f9mRCPZqoYaXfU8C6WJQXtej4B04yOcc6H8Wtb9FqZkKx2xxTz9D9r3iFcxK20FJsJG/4rZ6dIhK
T5YvsyoPxpJ+qFzY2EBcw3OAk16+t5pvtk0fbLRsIJjLa48SonQNw5dknBJS8VDLfVGccC9sjKyX
oc0QA4euCIf+c4PbtIiNgjdtl/hsNUWrwDt3DGO51NUGzcdQil35RlfnrP6Od5e4SJzWmqKosPna
gNklWcyCtPKnFuK2j+Arg7YkWMQXau/klYjgA/ySx2ZMxrPnqlX552hDqXqB20mncfDPo1y38XDZ
afYnzcUaQVOsYbeycrpZHou61pfZ7435n0hts174Ck7xAHmXXVuFraaG2qwj5VLE7HRGMTSGLAGN
sYXvMRFgWRuWJz/FYy/Afbbp3E2oP7Zz6WKrhHOtL9VYZcjibJPYJnxCUehGsgBaSqnlmmCyHkiR
H02LePfjrzUsFPbb6x5Rxu6k3X7cnToY9I9WKDD5792AjlirDIleq+7zaNLh/u4GtY1hQYVO1v4E
upLER0+h7a/LNKhFwZ3RltTAvYf+mFat8Z+arh0K29zSwhOrtkaEI1ARnrpPfF6POhAsx1zQwamt
OfmLU6jfOVkS5ix8USA9DlNq1HUntItOMQ8RzE3EuQ+DozS67NTNBS2s8HpHWz3GvJCg1vi7472G
w6cz9GKLBhQys/e93txYgAAQiWVM+5UeQkRVbqOD5PkGgtGAF1vpV9b5dShgz/rz56FJWTkeJx4l
ja8Rz2E2oMwzIxmnWEp+WwCUuPVQUVWnA/5xZXEwEUX+eWfy86SykrFIstZIoZTWHsfDABTUsOMW
XF3VhhWciIGEO8PGRx6IX+bj8/QHd08S6BBY2hWsZLGGo43uHbcVVqhxLBlXyTtSRyezcXEFfZql
/tctXfB0/ZEkyoCVbdcxmk8OrVIr+4Xb3ajhQhYWIgSv+Xllos2DhznS4Wq/WDvh8pkk54kNGRCa
TR4OmOHoWiH6KBMe3K3p56UXCR8NDb/M+Iy0xiE8YWBI1oUqrkI1WoMt/Q6QU5mUXjDO+EOox5iu
ZmYKJOTCgIAL90mOSV5GhUJGlsu8JwTDu9ziB2HESX5UBD/3Izn3LQWlAcfSPS3ujcEWif+wQBi2
3QM8KB521YJ3eGJ3+8oMpL8ZnZrKmmRMx/Vex8QN1qAZqgWC6k2KAJb8mJUTWMTM0ZlWKtja7K6L
FWzXDf670Ep8orbR35wyaAHSbECVxiwiGMqmPi9e641e4dvxqX9DTgSvOPRKv6Byz3/igRJZBXZg
H6HIPA7QGDCgjThAtCnbs8rMlpJqgc3kIOJPskIxiIgh62EC7NXO/RXV4iDOMvilfnCDWBNCw6Iu
HgEKWyboOyEZDAUBg5fzqJtjwByaH504R5UmHSW54WVbsBP+gaICS9AYrkoS9MJTOUGqexzlDOI6
Ou+qgbC4h20VqrDWPJ09wOxVBt0Nw8+a8gIbd2sARvw8Ojg5dbKD07wd/0mPHY2spxwPAeJW2RuY
IAT2xNfg7sUKlvEpA8iTRb7ErEYT2e0fKYfaibgcHkFcfewPK0gL3jZCzjwdzQ+XRyKYfSZqTZ9E
EIqoMfcBqXPivC6H6KaXGZMbQkiFGmEN8S8T6LbHftMwEJamPluIjK/3WmZJbaOdmiTx7OAipEnu
l0sfxCXPI0HG6SZT3VeUcj1AdIq0AJSN8w3pyNDOlo1y5Reri69NgUZmmxiktiGVzaSj5naA/c6O
Tf8NMSYkoBDOqG+o4UCiptYFVEcHPBU9RmJxdwdJk1nCso/vEalzhYG3Dqp5h81lCY9ucR3Wtttz
mvIj0Mh66YS+P3xIZvtOV5FxCcaWM9lQ9+QbEnU0j9LeQgredoCzLub6TnvW82iVyZ+Bd+FSIbe/
Qr+iQX1l9SMfd2Za8lEMwwX8I3BZjwhNmQkATxMRu2v2/WSRzDle0Y2Xr9qxA57RdNAmex4dS8U/
QF3Yt0oD6diIaOybcDUvjLVAOLfIy3rH3JZULcFLL3/2ZSLd6TU6o31XWZ7Br18DVscELfh8YRPR
d31kMQ4P6CUBm43CTXytUoqPzzi/CYbpkIZKx4NehyLe99boIPuxjevI4i5tLap3/5KmleXcsDMH
iCuA9iUroNiQMza9/hs8yIxfMk6UqDr8JhQFXY5UMfa8sNPtcljIyS3jJN0Xq27s0NPoAQz194yi
J+aSVj/2rdSt96czBivhMv0wJ/7xSrla8yMulI32pP9SiX0+pQmvT+h3kemqDYF2b/Iixwtts6F2
o5DDpnJiP/ggMK0vjWZqHoBoxeFhoBKcPq7QtZWmThVYXzrBZocM7o5s/Cqf6nqw1d6Q1S3TK6sx
x4z/NFb9KTqxrJl0gd1RrANks25wUTxQAawbs7HFmGqm8WDOnDNu1TH1lhJHunnl98qCzmsTHWVU
axYa3Iw3YTU7ViYK8LaXl0TJrE8eutWRVjXkah1ADedTRfnU+0as1ypQm0iirfiFm7L+2cgcsfr0
LuklM714mJOF0h2xUfJYo/FSTDVCoOoeSouNhB1HPmTe42s8cqlyMHMOrz8nSE+xzbF1+wLZ6oRH
rJRLzjFM6WuCX3BfbEB8RRbz+X0+kLTFMuRkJAPDLK6eqEQ2Tivtp3Fq7lXbtThj2PR6CihGpJ8Y
jzievoLUaXXJb7UM37JhJLDiHE9YHGN2fOL6P4yV6nrObNcf/aZIVSK+Pqpo6Y+Nt8b6IBf+bvzz
7uezgmpBgikiCqEbVm8s9JTU6NQ06Q2eyuNru8025BGH2FnquvyzOtdrgl9jRNNOy1WwQNzuH4Fm
UR1qnPCdsA7Hz5TKda/i7MhQ2C8MrBrx9DJt59dI4fBgKJS1KJJpNp+CiR+a1CTwfP/f61IeR8tQ
Fg3ZH/onngbXMr4TLO+sHAqLq1STf0Saqj3s2y8MTwrJj6IJGWMnHRaf/NEJsxRx9ZCqduHL1K8Q
SOMUuMfPqUVfwivCnrqkNxjU8aEg7hyTiRcNujNury2gF6EgoFb8eKUa97DoTWMI69q66E4GQBPO
qOjIQa0UG+buLiU7KbACMIcnE/hbT9VogAMzmcJsbBv4KDgohUgylWYlzkF++VkXdBEQEMvyEAXr
5kX81Jp9ydvNesJUYnOj0EjL15QLw/FT7UC4Zk8tFAFIxgfehSSFGzyNYPPLcpcAVVff6CBiB9LJ
V95ZaJBsrZbS9K80HsOFrplIsWsk383bbnsksnnoLvgHQVMBjAGpe1+QcCmEKAF+kB4LH/HEvcpW
asfBWBPT/39geUfoXPDeK84fz60lWhGZFOsr6HSKpDznU/Rs1B4GQGlByJV/6L2ZDerkDiKPzhQw
7+NyVRuGaYAokEZtD6c5CP+j1yXuRsZlO1E2EQc8FxlIDUnfQrpRLO3ghCivNlfTbC8mndAYnPtM
FguP/g0Z26yJQe2Bdt1LWDx1t1x9hgrJgY5yByTNpC6PJdkdte+Cn4DZuydnLg7xIG0UD2/cQRs+
Gazn4LkOBTBN+G96QhO7rxAihGntk3E7HXEEGYU6lvjHLPvXpgNLcsvi7W2Ncu0Bry1KlUMrw0LP
V3it0ueoi/EwyL05VO9SG9Oy0TrnQRjvMuVFflsQmSfziJJf9mHpSL/MpzZ5L7dPnnGrWeITgZkT
erV1yrlXssnrYbOYtDi6+XK9q2ZIi4JC7cb+mC+MDVOYgeoscstmr6JQCY23//A8BLdQt72gaEJI
RvyUNM+zkUfOHBZ1IT6Qs522av/axdVHApOlmAJEYaVaJmG5tgno5vOta0ufq40zRrlpJcAhHF2W
HntrnBQyPhd0lDCrx3gxQ5gs2zG7et8YjIZeHfqdhaztuuf8fR/zGpVWlfFs3xIB/gsbpbFZiPfI
S5wfCaQEjaK7q3GpA3bXkBqs7mmU6gfV0zBF5q5+7ZXjPO3g88xJL88JlM6jjaP5oTP0Joluq9gC
GstVziXh6z3ogWlpqHC9KR0QlnIEyhQ1aqzzlUqSi5Yr4qRDfYOGsljcs7xyhv9OyESQOEfEj5zC
zl05qBBi/CCIv9VvCZPce5P0zG5ZcuPxzWakAI0l1a0qHMjRTghbF6niZ0HKpHYGEzcvSXJBUGJK
I1GAk5A1luxemNrlck1G8zsdOvfEH1NuUW7ujGfADGOtc4DFWqxqNJr4AlzqB0HSPyTKXyygxXaU
CbhmQcJIY//sVTckcWglJmc5FFzeUkLo+xG67009MMnKlVYklvKpIndqwT9v6O41aZmq4jgLv/MF
VJ/VdFtxBsmBXphj0/JIV+1rF1C9r59bSSaX3jC5VBMBUZ5/K1eNAuYGLRuLtsDHc6Ib0T7frnpV
AJ37xHpnOTOoZ20sr693p9aYjxDYFr32GEfnXQqzbWYcAVokC0uf5zeJjk76Bae5m5M399rd17lA
ZmbciVhrW4fDdbGRAPMQx0IIMoDza4Iw+4rsmhG+VXgTV6BHyD7xiotqAT5LkKGwedZzypmM4mkC
64iyESHH3VN6joDpB1UoFVu4sxUaQty55QnoQxZqRKYy8UUuGOrBuohAPdQiAUyTegxdN9sEedd9
K5lrGtCnpQDaApVXJKtSZOym7+Mb8jrNmYTsfGREdJfpQIWfGHyjzZpMOcG7heSzuK8vlV12M1Xk
Vqck6UteC+f6p0C6geMF6a46XGQj18O9LJRxZ33bAocVfwd2iV0OnXW9+z5JFDzTTNJAPRVxdpdQ
tUXihsr4keju3Tk9UyoggfnLaWl8v1Ahj0Ak/CRSZqBoEmk7RUJm8SXQzKtbbeYJQ5gTSwq5ktLn
gBgZR4NzswqT2ExHb7T70g9XNPI6N8oOKcyD4h/GM7r+fotj1eG7kk913y7DIGUjejPTHNJ0kW89
VOH70lgAXyJw7Iz3osEYqMxa/dFVsZPS/l6Ld/N6iGEwkLt3KLeSEjhdjuXmhpT8eHchfi4eLH9c
6Wyzx7H5g+wmWab/Xw5xRkG/jyhEmEq4/VfIT6Csg/T0m0Ldo+65hfEZ83TogVxyyVi2brx5sEKP
N5yQr6MCEeKWi3tq/Cwc/+rCKbLZf4AATJZ1Tj4Khill8GsUskOiQt1B8jfZg9rIcQlHdUVx3X50
bTE92BUcimZ5gGGbN6j8/6tAKiUOYfR/CdbaeL1F/7v4s6Mh492/xBs8SuFTiNGr2f78IBmoH21t
xatSh0r0uKP/QYptIYGuumsUT9cncsMcTCV1bpwBGZ6nOgUZyHvAeG8b2oCS1GduXcQWo4SBmury
x8uAB/+9X/tycklWQXSqqp8v8SDTQyaxWXabGlPabOvC+Z/2EaaX6/1b53Km27JpwD3+F29SP/fr
UwpCJ/+q7gtTw/u13/L6lXgSrhVRCGfgMlK3LQffGFSdTa91zNrvAlbmkJDn8zo5m27Cgcc9bSzC
Y4cwMYgm1b2OaB+UsnFyfe6N3mdnRT3zXRRNisfjLUvvhByrS3gXkFhtK7qN3op5Hd+xZ37LT1XJ
ecwFHw9P9gwLr8kqnnyBd/XWW1YFTFgQWWZdJLhrjTrFYYng4l0BEpzmhm+IE44mZ7HYmzg7rFB5
8ene7pQIGnBf28fbUDntsjQw0vSxX3usjnUzyNCLY2lfn+bUucaghLFXt1+0QR4MsJZYddrI5EZt
03+gGJHayHXm4p/AAOriPcIdBQZsG+i6gQQPX2B+cpfSgda12/rcSfKcGq2FKL9Iv7ATNT5CFqW/
7SREEyK3t0zEuRfu398LylZzJV9a/P91m4LHR5Q8ylzyNKjkNR9Z3dvXFrzyV3AKQQIFxkps65uZ
wZbUSYR6w6cZdLrauLI5+aPQtChdMvDory0DlEzXsLvGGPQIgsM9y2m0CQwPGFGiY8tSm6FtYx8X
lEchWWkagAzonvkqZX/WX5/ES7Yonr0OT/TN35qBsA5xpbIW8LivABayjGftSyJhhAZhEmS/Wnw5
1uHRGtZndcb5x0Xc9+7XGYySYpGEmOjutxIitSGNnuKIRGc3UMSOeEocDc5JpCtWLuJMw6Nb6sE1
d12q/xCYJTJIPAxMExGuRi34XIE+Zj1X5oj+Pd/5TNnylRCGqEv1dWMPZmt4YlyEu1DXb3V6N3ZS
gyDXUnGzKFVRrThemFQRCqlGEHLGX7rt5KoQJBkiHC0OEAe1X6Th/x+CFOPXvUrQxGCgFwNEFstW
8awQ4KaDsz0W+iSNtPQeVqTVqIDCubrU3xP11//OskuQOv6dZgEp2t3/5qCKBlqugSbYuWW6cXSw
ezIh/k6dtnDi/O9C4e3iT79HTS7v2zbLUGhybFsy2Chzn/ULkh8WL7aRJ1eWdo6JAzt66ThX70vz
rpx0PHQW/J/v6YDm1rCv40Tju9iA5SUB6IZo/6SJpQsS4hQG/UV0TKlVmiz/fbQwD9i3Ofd2fG8D
DipgJmqGOkgyfqqmSS8QJ2mCngc2MSh695MlP2XvU5SmgkErUJOUGyNxobCkpzPTbkp1kYgerU2G
pne5y8ed4DM9WRHImztmSldSToX/otEZYKzjCDiFgCciKfd7fNsx+ji/Zq03sM4BIONQi6dXnkSv
BInHFlh8vGdAPyFbvgLDfrAVhOyX25JItsfeYaWe155qSC/zJpeImKBV71Dzuer3G3kpQEW2IiWb
bCvs/SnsL9ieH5KlVjU8VLxtuv3j5g1WmcRxqKYMsmh4lx3JUoQu2DwVRYq5dNozsmWTfeKdv2lr
Jn0tnNO8wxoZRhksrKERbcbjz9XwFtcUj/iYQombnX1XFvPi5MB2DZrFm/vv49IZHAbUsS/5mGMI
zAXYuFUDckYYziaNltj1kJBQ10sKBEUXMdupHajBhpStxxwP6Rd5oxoJwRk5vfyhEDtJ8tgiT+yz
JZNQJ8BvoZzp+xv1N0PnfmWbLEVODg3LZufpIaaekk87J3gSfTZ5c/z3JFdq6F64dmPj+EDwd6R3
JnXIQ3TFetrni+AaMUGaujYAhg8SmFGAiVlHqnlPQqQBlVRxzjK46gPjWrn0QWkykmD2QuJxBig0
RS/TEEfhRz0Ripep82xTK/c9ficDsU1z7VM1k0W4OtjZRBucTEM3xqFHpFu7Ru4gQlZSoK8wSkbH
DrFDKTE+Nnpb4xFPYjJeR0Ue0rgPK15owi2zOLZHaUoZiwz2O45qSGOalk+LNheYkSkLNbOx8Dv6
ceT4XHiO7KIxPIeych5HcqXJYet/2QRIw1C7WdiOD/0tKSoxdtVbi0ScP5wm90uIB0wkU/2EYVF3
R2DiFHqgwXa8HqPtT/EO/7hvB2TW3y0V0Thdk2SSPmLt1iEhFCwvVuz0uX8aRFZM9Wfzb8QcQ9VE
cTXHJNdoqItJ/5dn/8tUcqvjjf/ugWHh1VaDjz2cWe/luxvBGuXg5v8qvY4lTFr2C4whSc2Bteyt
KZhRut5MWas6252xudWvz6oKwZ2uCdTErZQHrCfPpPdU5UnBqy16kCfncDkKysMbG/ZHLQscuPFP
hjaVgVMQGNj8AyM9Id3w01vFNe6UIiAT2C92E25k9OmCNNnFAP7s/35rwPp8aQLDzpbxMKlkC3rm
CUu4bV2nuOqz82Cy6TkiHHl92sujahyOjLcbPVnP6qJVvdoDcSLyeMSu8W25GRsQRIqoxis/BBE9
o1UddTjn1UySq1slT6Yg2FcCfASE5L7aP35SkhKcmxSVC6X4pKFaWggw3Q0ZLMVU4OUo7SwPGETb
bYZJpvxzYkXRkOyamA9ojit7ltA9K81gnedyue0Q1GnXThAZ+mOQ6QMsztWP8c5bXOeQuhhBxGdM
Sygps+NOoFpHVtOzyM9dKL7FZqM5+KwFeA90x1AMNcu0GFGL45TrqTcpJQO7rQa6wwathW6t+KSI
C/jstmROtxRF4ORNUM594M8QetRNK4C+wcpsHJgtrIQa8heNbanqJv+uf6ApyE1MG8rii0UZHdcv
vRaqrmEcZQoZPJZrFb72GTNQF2u5IfDN6TlD0w4n8xorp7pqcaIRSOQa6oXc76Bic0tu6wEVvI9R
YRQuzb7vJy+cUyWbp0/Lq0I8SLpSWqlFpbN0+YE8GcnuULjr4dce0pivPMHoG8cX5bIZloczBhjh
4RGIlJL8i88MY3O/sX8lYQG5tSdjKi5NYM/bM+BymjZ86/csctrYgMHZ3qm3UxvSEENfbhMKEWyZ
A9w7Z5VtV75UgPBs6BG8BLuDvnQopuQC2xDd+zIez/XpwjThOtMhhz+uLK+YpTMdAjMbamqkkYQv
rbUbFsYDtPeVK/2xLAD7rRyWmHutl+clZcOEGnlX6e7v6wOQ1/K8hQwzr2E8ttCpSL84TpRUAycE
G7uN2/LTDsyLxoVl35DAPLLgSTR37YnCPmqYkBy/rBupFEur8xdBpTBfmrbIM3MW/xmjfu+SJg7K
j/Cj6252t0T07HaxmN63uu5Z6bRHDBmVssct9Dax9ea6/ZNgxWzw1EHrKkhV9Sua1DaeWXgQpZtb
wHqe6tDS85ca1Q6SvaRTR9ll65+FBvmJOwWaobxa9wzS0Yihii4ePpY1c4R1lJ8C/1AF4uPFFepr
YXR/+vD7wkdB/RididK+BjvldZnyrOqC2ORGN1SDHuCVejq/lrm2Z2EHyMdYVfH2/dYUYUZjaXWl
Z9SIBUafx4zLejbhyOASrYTUu9VpCXtOonTlXZDADsP1FcH1Z+48oXfjcHDtUjQH9eK7wN8cEVCf
8KcknjBvlD4kK6b/M6qvXH40iwsXhSdAV+ZlvmmsRivABiR4SGI4CFqh1eltIfuVqczS3UqqrLJe
IinSLnArvYvoovGzJA3zf/I+AQBLkVIRTINQuUsq90h6S9bl+mm+BLIaii6sUrYpN4aPYb34rMwZ
p5odjaeBrRb43C8U7xp59BaOGBqjRVL/EuXNecfZHw+1J2ZAkgiP2w+afNsBSJtOlqifh2TlvD7r
Y3aMixXMC1j6sbxWw54ACEnFmZ8kK0GF6+pFHMj0Um3envlb1EMaoIisGDI8KSRc+FAU3meMt02S
+kXb2XWu5eoGISnYiWXYldINatpPlEZuFBgZRRPKUbnRQRUNuM3+74pe5cgK/4tBNLkHmg1eOo7U
p1jZAkmKhZFT9JAAs2FGRarBJEIwj01pj7ozpIrbvSzabptuHNCLYjDIfF4XISHOCz1PJSQc5DbH
eDAnQCqPcM+hqaCXXYdseqAFMmbRfcOL3phXPVJgPAuiYTn6iZpV58UBVWbDR180r5zyTDgEY1YO
xnsBjj8zAUdxIxx3eZuV2Se20L4WDnRAR2UkZY5ouLNzcXEhXD57PsWpP6SdyTLQRXlEOnTJJ5o4
isF0P2f8j1w2aXtaeNGSt8iiIzagEr8UE/IoErSKLiIBhcWQeNLwFBK/KKvpR5s/P3iCU7wAd/J1
dMl6TG1I/gV1YeMhcYz+sXIk4oXkVLA2jjiRWbQYS4fx16IMDWUDuXp3TIQP5Q5fqjdovmcYYwR6
J7CKsUisE8MfNCr0M93iDBQBoYtRtIyTuqQKyW8UTM2TXpq71V4SR4gkPnC0E2RNs+OpbVfJ44Z0
2deutardAf7PF49F8+iDZgyEyiSEocghNwP8K9qIZ+MmDrOJHi7ZHxkXVXho9GwJ8MyFLP2b6Slq
Y8r3pNT8Z+3rcMQp5B2pyRiQFJAkQg6kfn9U3clx3abpZjVcinsh3jc284Lk7Qv0dFNMUsOv1NMa
4wJkRVSVy3LH4neUrIt+nJGQyTNg2UzCmg/z45impnQyCYdmOpb5wtOkpjoRMKH18YX422lfc2bN
1Ex1p7SbserbSNSQKSLofqZbf1e7d8qwao3TXgWQuJGU+OvfB2aTFwReTOVsV/EHpazokBRe/k2n
VWg1EtuQ1QZ8PT/HtpAb/KgEXMv+59/ImLXjs3R5Tikd9+6GyS/iBTswzJAUqlCr513BQ9aEqcsD
xFshUYo/m/tbSRLMrAlrHci3tEKdQNVdbnfHQfzsDfe8Z4c212oGkg6CT1CLoMjJH+DVoyDI6glM
PCF5vg7/FjK9CVQ5IXVMbTaaxsfkXNegRQsKjJoWpy4KudRkFpl1w9o7cqDahladZf4iPci4lUvf
I6j1OluV9hdZlR+eMjVcm3+nDha5kKj96ct9nrm/Gik3kSEHhyCK0BsamJsDHMoKNshSwRel7cao
NShUgyTYgotzg8INS2dZM0udFmxvVdKWYLIJkN4ExyJUD61zYP+WG/4JzqjAPZ13UtBCyTJxhFJM
RE50EzT31kAGc4j3Qts1VodfYjDlFC9eBVAQFLkm0e614xM4C1b+Ox5X/XEJQkQJo57zaMDSEHLT
fhgzEdfLF9j+/7KSb82b42+d6R8EADNz7lfieQIEW5UAS2+KQzVYGdlbCiBQFWdKq+M6irl1vIx5
7kgCDIH/fIFRj5xSy7LtxQf+sgnt+iR4R+cXiA5KvX/LX7unM0UPjsO5W6KvarhTJAsjKiDGYnHm
GF8Z6Qf0ZWOwfbFWNj0oH9DwY0PaEqo+Cx/BkktOCTsMd47X8a7bOjj0BpXQeA2MwEq5fp3Gm+7o
d5iLxQR9Fd/OBSJhYHpS7Kl1PY0dWVpraFFGSdosBIo6pabNeHOuRuCx/8y9Y1r+V48BYTjL+GqJ
lBQHPUUuOMX0mi4/jgFHV8v7WDzqPuBwnmETLxCoLynTpYf0qwOwj+4Vp8qINqbmITMc9+wVWlNY
8A8/XmVOiOacm34gAsgBbFq29e9Nlr0oLteru1MXnUlq8vWpm1rRcjaZBrimpUpE9/8YBhweSqC4
SjkSUrTAm8opu0qKHt3LBY4ADMTqd/FO+FIkxIShsJ8c84tQGvD/d8tFK4LktCALQEkUwK2oq2Zm
y4eY3O3Ftmw9DfLroSum2D3sRdVWdR80CwArPe4V6feIpgayEjTkA5SEoysFbXfll0+gq7JI6z9o
vGVJGRY21vj4US3jkvBuMKyVzZZ6eA4Axpcy1NM7X3ttGVxDrLOvoyNUHvh1N1M0lOvTfzqXACgE
RUARc4YdiXIiwi2t3j4jpxprK7zidYVcbCS9J9uiWBkeolLL9UZAtUrlXwig6Kcna+SaD99UciSu
tPj+FjbNZvdnIBx8lMn3rw7kKbHYV6fR/LTP/M+e4US1/lMq6Uddnlv4Sj4kSvAsdT1hZ9b49l96
sGja4oKJqcTUZZLOOPTeVl1yWTQtqxJeoRKD6NNiCtBRsnuwkvSBVLoE+c/+fVM23y3Vn7r3TIXn
E5E/lw9vFp12emv1jkoSH7QpH/4GhcoJISGoW+Vt10sdWOtw1kuu7TpIa8jIc1Xgb9aXJUKyUnkw
oULGXXYKFPiJcMznhhDGeWX7391Rc5QzJsK7QP6+vXnbCOHfwVJSw15xq8hX9JCY/kXhZHoEpb4d
vUDXEnkFekcNnKfBxXH2jckcHNsEZRTWGxIvxcK1BxIIu9dqHCi0aF7C9Y2YOUG3TX0SiDsMLuoK
kO/6PcUzKXT7uuLsTUtXf/taORrzupHt9rJRLq3oz90PsD1xMcbvzpWviaOrFlxgKn3VdWxg1KG+
zDr2aPz4EiLm5qEAsYKXrSUoUCY9QXWcCj3bDF8iRFrEXfAlznRUYfFaej6ap6qHrWOlwINRti7i
Rs27r6ByBSYkT887T0eMvpKh5jqc4eEh4R+k32k3ct+kffazAkXHA8gDuNdfmNJI5SaW0pLFuisT
1/09JIwcgEDyz0fQ9a+/xqTacXaUHY8hOTSIMKIuu3j9rCcPKgeX6xmTi5nx75/VQsBW+Rl/UdET
3A97hfwBVTfk0Stl9P/6TS1ByBP//qgbd0B2qmWBxSGcYf7YYW7/IJDdnaIZJp9d4wf5wePO8zT0
MVxgz0MzGxm51rftJGLgUBk7QHJouHCb+6NgLFd9HaNtp/BMwX12c7RFQKKqmIrYmrD0vnpkYKvf
3rNC5SOWNA+EE/0h/LKIjrhdiJ9kpcIXtvGBG/7VkJqzGkI2fdYqRkrHXH0N5PihCFuuIpih8Ppe
WGVRY9Xknyc5ss5a/9PkdSdiqvYUKAKuPDzHND6luS/IHcAn0yT20RB699aOSMAjZBYkgHU8ayEe
mXYTlnj8zhdQse4iEh8CoClrNyZfKba0NVaNl4e2sK7IHiIKO1/WzeMIn2TSYoS5o01QZ43zG54z
vL5XP9gGuiSmMEU9/6iOaPMI01R4RXXDZVcBzwjnfTcizRIqusCFoL9iwkF0pN3XK3VOjDV8jLAl
LnUdoxXCcUeVzh2jcXVGBXXyYVLadjwUScA0VXI9/JqZe87riXQyicthWTIpvdcjrNDCAOHU0pVd
4W60wWdd8jbESxm25eaPjMwv//CZmszgzDapKEPsiatAVmgWUq0VbuA8ulP6MHvERz8NDRlPcEkP
HBDTvjiYF4JmDG9v2IKg8U060PxP/a6vjU23azbEA/EGQDBY0WssGsuqUJGizd+lzpROBSKXcIeb
t0MhhAmnAAP101mB5uabBCRKr9S0dLDoDwaFTCPKHEJ0iU1skJlIjOZyU/OahKuP9oUlaNIIHzP8
udnD7R7O2IsMvUQ1V3ij1S7jnmzJaAU+bpdvEE+wC0M56htu1yUllGopMhN7Wn8OpAqgl/CE/eG+
Lp9Xk0D8dqO/ULe0JkphB0eLhEXGHIVpcvHmnTAIzW4MS0ckpm1E4CqqY+QJRZQdniUoZxmC19jo
gOpi5NxVOPSZP4EBzcqJWdsHmSBE7XZwe7G+WDqXNAU+3YWyjz8Oi6/b672z/xVytiB4FdPQf7tb
8cWyxMXaFjOhRa/3X232o7IJuzNf7cONsZhjZAXf22H1egIdQGmn8rvia56THWhNCTKvVXfcK8Ix
ArwwBk2OVMVcd0XpxQeHQCI6dlLACiaqqrVCbtzgjJ6oGtT7SWQ6u2hWwXlwPgc1JGo2YQlET3pn
CYMUnJ85xBPHTCMBrRSQu55TD/bjbHL/8li1DuiHtxttCohjp2g917qUuYWUl4MANyszvkjXRgIe
eUzzL7Yo8CC0hlY8DcEtEB97fMcmJHncjg7Qjt3KNso7nghQGszrMIC8iCtYkx+1ZnyEr0yt0SD0
mCcbnnrxYyLNPj67appeQXw6Jpn4uA9HgVzLNruGroJsdJAQaQCav/6p8K3+El+GBhidpv546zqS
9bFYn05x2RU5xHeM2dmaBAUU4/NtLbh8sQgrYoNUXOreyyDx/xuUofe++Nxji6SBW8ACy9mClm6f
QiBeMx7zS6sZf+wGT+gvlzoOqxf07iWmWB9s0/vPPd0bB3DoF2cgYeyrVD+p6cY1FzmZol6vZVPw
I36QkhztQK4q403b+uHfL7ffGJjd3ZgGLQJm1tlLKOEDAJrkUIkHE9K+Uwfp6cOpQbcwjXEzFhtx
CBupmuq0A9q5rFkTUjMoa8KeZO0GAd6fLjMXqrCmjhLs5cPJKLIHkLuph6d5ccQpGjFARsIINuK5
Z3vREK8Z/dcM0qe+mSj14OfV2fUC/qpV+Jrdj0bXrVPv13P/yxeYxyqM9fe18q6I+iU2AdW7RTXH
veqocxab9qnzlgNTMrDUjTcp4vGAAhtITnzHvf/qTlz/oMYultlazD/jE7YqHDzGpr0S9Pa9WK+2
mz86ZqpJQR8RyeC8K8deLjyjKHArN75IcQ7m3Ful/soiMjT5AjbzowvIDxOED4KqoeqTXWwvfM5E
l7dD+28MhLg9Ck9YiLLdORVhzRTIO2mbWXrspo4IgbaDcd5Xk3jzfA8NSaLvcFSx91fNGv3HBt9t
/HnsB649xkR+ZAGoDShbiWLsbWporCh8uGRw9qW1j2ja/SUJR/meWO4lhEsNCWCVsvD+RhKtkyNf
a8oDqhaDdE0+IMTcoR57rJP+1v4bZY1VMbJH9NeB+ZHTeMI2IxtVIwMimPu4fcPAyYqwvXd/zsUd
Qv0r5bu348y/gQtZz6zU9WpjXeGgfDIv4DfXPt84Sn7pQ+MbRIstXSjQMnbZgivnmcln7fJaEByi
F0pPZzRRCQNbOkgLO4KtX9aKs7adrexodMJN2TwoAkg59iShIv4M/bDvhUsOdFTNjyEX32Dvk303
zqBu12ayy5O7L4kkt9mR9h/rf4t+l7D0GWBDuWx4tEY8wIN2BxWq14pfltmISmMNi4vFTu1N77yu
t212P6Egbov4m7Bez6jnGYPzsQD4NXIXIRRWelQMA42xGwOQcF6LnpfIllJz2N48HNSTMFbWvyXo
CFUdKt5+fthNfEeGvehjGqFVuVt3wUk4V9ChTMB2IVRiBfWb2weME+7jTVX5i3QKXtbRTvgzfSVQ
4/nNE5i2UfhXukb8lAT0BW4W3UVUpgiPkoSvA5xrawkItRcsqfNBB4Rw+/G0rhp30JbTFMq6K8er
0aNHWOcnIGTip30d4igHv8+9xrJnmMAjihzXce707ekSf3OK4/BW+d+mDb21qGCpZe2OeEdj6ICA
7vXQqgabj/f1xUjDZsQpZf4HRHXKWi/4idt0j5aa+y3hMLZfkFAOwkgSsbr0wIeyQi26vWJ+LEel
7VfMEraoUTFWjdKM/Um7A2nWuuzb6Y9oLXt75XeAir9LFbPgIkngXdGFICt8DLeliFrY3YMa2lPK
xKFntP5EybR7eR5cR3ieoHWOkmKhR1nbs1bvvF4x0HCooWPX1Q1MoG+xi6+vykDIXvEwnHeEP3Oo
K/FXC2M4kkjGga11fBzeK9K2CJK4sSBZt2t7OucdABZCIWtzOsDDTNUrCjiSof0CM9G5iaj7YTLw
6rZxIjcCQaCuuefh1fezcW7NsN0Saaqawk5qRX46Bc1kBtQN/Qqgj8f4blgCYR9MqF/7LNawOlLc
0sWa4zMZaI6JdAqp/Ykgk1+Z+VT+8CS+GZRuxT6t/hUTgXT8GYnW/9ZB5UUuCNpziZt117vo7YBb
kSn/6CMefOkO1nYL8f1L7YUOkBqDoBgpoxmXyVUOeiYx0OJgPFAnSATF2QuQk0SChe2gjxV8VTrF
ZpvEmpr8jMolQdSNe23cbhIoN5taoCJQqehBdYc9+j3LNNUHQZgCy1mePyoZxMmqGE/iQ2Rf+4wk
9pApniwuEtJ4BCoGBLt1OevJIlxe1Bs9FCdqkj6fo4p1eHk2EhmqvLQI4BRkDE07OSJageTkCVW0
Dhds6+cMC5KASlhH3BBAfqFCQdOSiO3Z97mMoaNICI7VtEYMmXGuyExNIEcGH35FqLNmn4JIofwn
O0hhjCow56cjfYGYLncZivGBjmX4tpj6LFH1jqi7rzP/8Fp+C/VTqhS2X5XtG8XUkEHg9opcI0z1
/JG7VbhUYM9nSi7ef8mSf8u9ClcjrSt2zteQx0BWPjmoZ829hHJNJ32CS9aANfjys/OFslbhCQTv
HtHd2uKpW7IczvTovObmVvNbV/s2eXXj9f4r25iUM8zKnBeMpdlSy11NlGjrRCu7IwFgMn2qjKb7
D2rWonGQYblfmGEWz1JSCW8a9qRPUvkbF17V4w94mg10Um+DXHZ25xj/VT7VLIbicm33R6onrnW3
ib3IRaKxftTl6n0Cxs10GU08yCYJU+PIu1VZoQReasI/1GrRmZzM4WLQKJDTAsco5fQC3EUxX9W8
5l2J8RW4viL0eSGbkrFo5OGXkAr+bCc5tOUnJtJoGXxn2gs8hFRnI4CEmmqNz3Tv7YadyoQgzy9n
pw9+94uHaHkT8NKE83muBBw9fBNG9WD5NeG5QYadmm5hsL1agdMYIqLdkUqK4LPH61B2LwnSiwgR
6DaLX0TQdcuo1A0gHNGn72DxzZmcdyQGvUpMLfwg44hlqkBJegDUAZKr65dzbGpkCWcrc3lrDtYz
7IBh0avZ4MflUEEwwenJMPWYDNRLlBcwXQ8wuAZAnzi1UT8Ai4K+OG3i7xQHk8IRrg8WFvrSFXgr
a2M0Re/6rbLiDuzwLgwNFFL5THg0T9QyeVho0oYL5YX0fykcgFP+tuDkoc04kVZHh/QTPv/Is45H
O6x6bXayp1BZyv+YgoOWeiySnbOnc+CdtcWHbhWNbXy9Ce3nGlzkZS6/1amuSjT3SJC72ttVwmfJ
ChsEksusbcYaa3HfGaB+HuCHqihb4H3J2gUBQ96gIfHtB1neXg5cq4mpUEvFub5T0AAbxkpqNH4Q
s2heBJ/If5kL8DsISWcX51kJrBy/i+bWVgx25xQ346mQFVyHOnVGFMN8siHPBniT4PMuritUQqra
epOTSZzataK4H9FpfDWWXKKheV6Z7Rl+T3mwQOtPS+bBOmJ+FtnVu/ZLn5bcnroW9KPXKUvnqVqQ
Q7j6h18pSZGLi6ow7nqqTuxjtsFWWIqL1FIvCJi4096mX52VGWBfBVwmrntsPuw5cwzCIW4XSNOC
KjRrGS4UzpgQ+mJJTwnP8kXfPduaZZXC5KNoa1zrz8yLwB/N2jzz4JgdxtVFr6g681icFZsbwh2r
6uNj4WttYsSd2P3EYoIKbuYBV34096MmjLp+Z8FR0z2opsWioBqH1u0Nq4CDzJs4/pqWDORRq8a6
VffSuCACkm9CI6WzEXea39U+0xxojmIWoXdKzINgchDS0A3iu6f+jXiOSI+ScR+Wh1mpwi2TXiED
gSfY7JDWC6ifYGc79XMscACZwYS7MLJ2ui15jVglb8iqXoEMQ48AEzcpvCKFmGn/A2lvQ8zVrlDi
aSU7Z7zZNVgHD6joO23w3Gl+xmy1d/Op9+cHfdPajzo8FZdt60MicV1Pl0X7byJ8/R5Lfc5ERzNZ
v58so9u+1bSMDXWD5miRmffqZg4flBFuYyv71yhUd9S4bXatvVv1imazBII+OzBj1VxVnnz3f3mT
eykNKTHdHm1029XpVyN3l/JptdkgP6sjuiP70jRJDvoJDBZY0Z0+duGLdhaLRGLcZj2jVlZ4ylFi
/2H0zbBccrAuQI97pltKOB4hJkVN01DT2/wNd6aS/x7TyAau0UQLkPONQ+KdIxzQ+KGBS6yj3Fj4
ckWlMqYbh/RZ7YG462uj06fX0d9pbP9L08mhbKIG0Qhc3xHF2qrt5U02KYztDrZzmW1V0FJPBVZB
h4+IVk+5EJ4BBL5RqVzFED6XiOxJ6U7LWjDtsDbG+WIQ6K9tPa9P4uC/eHTNCCAMRw8Vu+Fxu3EL
Cvnv9wLyBwrAdtlSql29J8nEuqNVweKuZwFeUzpKAxl7ZTutpckm6+8OaQQxw2QpO469SYntkwXM
Yd3fOs3o/YCs1UzBbmBaAQoi9roGCEfMW5IwZMZfQaKWLd7navZn3K6wQGPi6QMb63qas5adolW2
CrLPoEI2N3z6vsznrXF6VHHBZl4+cr4BcrC1KsCizgStUE6fBIO+u5CYB1A+1LrMXqQ9ZM96Lig/
1mVluINQSJk7AZMgzx/pfePVSPtUjka2/BVwemS1puYSdEEdzca8EfAic0vYUZsRd+cJtdu9NGGH
QevRKcGoZwvuWgscMr77OnU4ZfpYeFDsEkx+PasmXb59ZQi2+SQwpZGOnn35CId7JKVaWuSyplnk
Zf4G0mou9CGV+xR4YjihFbF5HdS9XSED4rvz94VKzy8NghRnI90iZjrNR4rDx7T6XA77NrSBILkc
0elFNFnDOVBQl8ncxBYJr0slsoiLywPeWzJIFupp6q1hu5dahwuTLAk9e8adz7Wc6PqkEJN60Zw2
DE19GKEy1wTBivGHvtVdU+d19fUIopoyTYZzZSrG0l/D+t4AjFKufodoZFaIgpMWaiEZnidSzEsR
bCTNTmJCv8TYIgvs0onsBaJo+rtKdlypb5m8PyBLMrpmML6yMsAr4PqQm5+DXTkSv7Zi8ysVpCLs
GOapEkUTTZW16ZGlkO9Vjru4bVGXDZumRpuFCvfbNZhKvAsZmnY5syMKdKpUCdXJQxo3LsnoIUIe
fWb6JeKnlr9Es6CmR6VGHE8Qbq4MVaE0hRrdDP82FgWMfT5293uveDrQban1dhqRSKch7SlRTc+r
BVIasBAOyDfoffjKs4Fx0/lUqe0S3fHdJkuS2N/1BgVXboZS5x5UgH5xlnifQNpE0nvGkzrn/NoD
U+g5RRWKWpWADNFsCbByEUbT3OvO0Z3atRYEmqZ2ae7lmkiy7gXniwpTuHmjXVBImTWv3lLCPuP4
CeN/srszm1NAy13oeCKo8JlQ7Kv1LKb/46+KeNOu/lLzvDWKC2dekfWfMy1SFtGwl9kkE9dCZATR
WdUmX48sFbvGBO2Htkoo9FRfr+iE8kt6a/JxXq37CV5CfZp8A0kUREbbTA7nhU+GJFttQmd7Vqa0
jJLMvg/LlfRIG5quZK/me4dfbbmx6iYOE4CghOA9HNUoNWzh8cKzi3QqR6A3m8V3PvwW8o6bweFe
R3D74kOXyPjPphTrusJ+NyEdipRON4d+E6DHUwRxwQgRJlwP/NwvCyJJZMscRP8r+atflNlh3Ws2
+VXWdpr0BuzMEGnIyVRCv9FSW8fPstNJNnp2CGVErEcVmTeAzVM8tvIjW0BfPLszVL/q4MLkv69S
Jwv3K7U42zhwaLIEl7OYor648Ru9HKoPBmIYNwgaqn+IV4z5HNgx4upe1o4oIZFoE+XKAdbAVFjZ
yfVxViPc40iMKJaa6pJC02WQ80eNmFv/anGh4icPwqePI7RBPbldVP0Cw2C0wk6ty9FHQK+bjtMa
xm58nDyc2Dc/xPADoXVypZUYVWeiAUglOWD7YbdaEeEH3JpHcq88csB814Tq4m81wpzS31jOrU2Y
UjA50C2S1ETJe3DD4XJE6H1cXkcfeWu8ANDa0Tb7A9AQludK8k8c1F4nkDsvYSrHqhApHh4t5seW
ts/s4+yYr2XvQzCKzDVD2Kp3YzPQ+8iBSJVlrSn78UGk7iuDfKLCQlmQob/iniJTJXDr3FGSbYBR
n2JWCGV6CXyxCt5/hopMELJ4RctEM3pI8itvokJBjt43iEVbESamCaNYeaFbrxZZo5FWL/0PkFRa
be84oIGepF3DpObVTKbnY10CMkO5dCkBqGc30n2RxF3oeMfA5vuq+6z0RELBvFgC/wiNMZJnho1e
mGGKNB9AD8uGZ07d2U8hTFdWeRGA3ojLjcgbO2tLAJDH/RQJOQe23NqA8Tzm12+TPJ5p/XweuO3O
I222bC8ELm4PoIob/Z5p+l8vNcvNrVH9nD+fy+ZBIRiR0heNt0MqIQW3IJn1D5w6ptv41LnHo4Sm
eBc8u/c3YhC3xVIsKEJqYGzhQ4fPm1ZZkXJNOCpHMOT7nhUY8RmkaSURZRg5bfa3yfe8N3GFgMPv
uExPZCIddM1Hv98S2c4KbUV0RAp56T1Rf3sOQCiSJnAe2ZExrdGtgUcGsw3anohv3EG+bejIVSBq
tiWEw1obgSk7bbb1KraSomTqq4PJVbmbYoLz9IKa8LJ0sLw94O5bJLZuMWPSEdLaSQo/pfBwh/ng
HJF40hSizhLcnR1RUgoFfuT2p4p/ix7j2U6OfxYVt7CwXkskb+W2GmNunrz0Q5AVoE3Fd6tDD8TV
cil+nrziluEQojnyeDu5c2G0/8i/0eMc4MAJTVrBFuWLWR/LSLnl4Q7zqAwfgJKcxsn2P3u9h5OI
MFoKmv0u9GHJPGnSUm/elAzexburlY3fewW30e2n8tPxvTU3yjDxJaIHy+JjZDUrexhlf+1ihxRY
6rs4TT0qhZfqYJ/V8eM9aRGPaLaQl+qx+rNdf82HrqgdZ6F/lziL8SXAe5Cc+OnNrbrfgJXTVVrS
1syRk9Xw1yKhdUuVrIY0ZMdBWaq6o9LFPPnu22MKoBpbeIooCVq1kq3EvlSeLvoAH49rWL65Z2Zq
+eghGUXHC1m0ZQ3z1446ex5c84ItvXxWL/bXaf2/Nj8Y9sRE4CugM91hSz4rxa0513KLfPrTAXAn
+CPCYxnoY+VOD1pOmrkptF9UWQw1LEkeEI5MAzsvzlVJU47iVaXiKAZPaNWNPCRBHXIQaoTGf4PG
to75caGB1fa2AwPDMosZ0BoOtpCwo7q8ESka0MawyU1d0djizEInAukdbx9LRN/846cMWM6BQHpO
azDiYbMMZJxb/yE1OQFRI8z131jELu4aCZiebE/FpwnFUU8R0a6adodk706ivHErShojiuvzv0V3
/evwhd9tonob9l5bl+J5sP0/gr57leWG+YEeboB1RWHEZjvOxtZyJq9D/f0T7zefTjtQAKvw2Zad
ueDR/ZjlRLWuaCW03Wm/99YxZAakXyuH0Kkr5Z2YJxjdt6m7yqP63DyzJXjPVlSwSGdzJKd3vqhN
FpQ8zW7oIRgJ4jaAudtUJqVsDc7oSF/UKcKG6gEszVlVr/pd/e7PB/3F1GOBNSvkK4R5eLc1YL5j
dp/qVTzEe1tYHVgt6U+AG2M8HzYjUTFkrNfQ+GTq99eEm9xee2/CeeJLbpxJ09iOMfjqlaoxzHRq
xjLsDBlv4qjzTAmKCD7tFgLmT7pRSyN2/SQHFRDnMauZEWtBQQe32y/4GOGrgXksWbrGzH+5Lndc
EwCh6TDBBDD2pnmG/t73i8AUX4UxPyebR7q7RjrTnqMDo8vqVV3O3a/9LuJyRED3XawLrm0rAzM0
xyUuhv7wY/RMwLg3Z9W8xKg6cNiV72XXLlzKh8kcyxZZsbL1YWHcON5K+UTC6UMwIoelwdLeaUgk
+PFaowpo2Zs5EfcBSlkQCUqJyGBZ5domHd+0DomR0Krnw9lKQK5expKN5DjMCUnARqNK7kh4XtaH
5E5lSsp9MF1/CkXkAO1VGAa/FY1krRYTGWIiuwGCzQY3mSu3bma/WqdyOQX7+xBnMr31KVYHflv/
4IS8p7YR7AVOB97ma/yzPduqy7Zj0/HCDfUENGAP6nz9p92nCbut29jUA07TV5m7MQKAPsUyNjQ1
PdPg5AjvuxUaTaETzsknsSUkLNYDLQ+Y71OgpwfbMG+cwDRLL9+0yP4SwapDGRpLmHZXZI+5Rs78
QbsQWGYTGz9sgO5aMYx8uXAss/Mg3FduoTuurxljemPvWT9UUykFjjB4LcxvFvv2xACSGUpWdjaj
haFNdvzoaO+Sig3+II1Qaam/F33i38tv7OsQ7fQSnlIwNpEQteuALvObDDCfMmIzKdvuy9jzw3Iu
dOpz14po3F/mfhvhvFSdpSKXA2rOYrCFsUnbBkjrGikgilDeJrJcoCdu3llSJ8Iw++EtpUU1Cj5u
96Uc5+lES69LgziNs84tqXPQs7wkvPMKxqvgGI3Qc1k6wBTl94J/KJaS3wpC9J1ov24mdOg87XvR
Zn57qDM7wDMDordg+5AI4bFujAwt9VRaWN+aj7UTwf6lzirz2BJ3KedUs17WYxuXVrdnmzd8qwwX
3wwJVT1C/hHmybjEo22LM4pLg6w4qVnqKvWL4Hysl+aEUhkWS4oq4cNbvTJaqCbpZ+lJjTLkdaII
DrHJgnJzRm20sMG8PQrLYNdftIgXNGKWLZ8QMd/R4EME/Tb1Ngt0YyduGS+WhLKyoevM14wzHOr4
f5Ne3z52Qgnrv4nwYjfWlLRKZxSwz5L1WZgO1V6EqlbVglR44RU4jxEwAVCrW3gCg4Xv/VyG0/f5
Yy++bW/RfiAFHYvlceFXo7lKgNDLWO0LnG1nKvJG6e2d9n+iJFPkrFvUkW2LEot+McTjWMvah2pm
RPcn+iH/eF1Jp2StnomdLMB0tUlL7CveOkwQ9Qinm9kZ8F8Fc12PUlkXHW2bQ0SolCBrnShUlrZ8
aUTEbK87lsRGVOwArxzL2BKEA9iVPIJyyoFba+pq55aQXjqvghUdsB8ssVXk/ggWbsWBPutuY0/t
WX0pB2ma7tqaRXhEqFhkaq9EWDXW4pNJeqL968oJp6FNelUVICgblU+uwNmdlMAFzCcxWbf9X1m5
QdKjCvFOS4YEIC4XNlM+V7wr23h3jiaJv/vknpiyNr1HDdhX3B7N4UuuF6KYuNrt2LkraOzogW1S
4hzTeXfquNG+vgiWmahm5SMcD8I9NIxK3OOPiUQa+tA39mu8iX62gSoRZA0zFLgkHZBtKeWfNOJY
znnQdvinWWOBC2H90BET3qoJGmXhq1w/I2OmrkRgYsXY6pdgJdX+nq5uvH78jiHIFujIF1PTwbUe
85rZFO4VpgExidgmd5I8PoPjtsOld7GK6gr+IbGak14e8pBtyO0sBm96DdYboeudPpShrYP4qFmv
051hZOp/JPMpxv2JDgodcxUslSLwcBpZtyCFU91KKqy6bty69iU7yiHs8hvJ3xSgQM4m3m/u0cr8
yVOMUvItbr+q47Jk+KWof2RKM+IcbBkguElqqdcrvNqZsp8rqOdLkIxBblvTlBb2EtoJH40HWKyA
ZiXGq7ACFbM6oWa6REpRLL+gEreLrg65WZL1ypFvUZbwlVkA0bHUCtbjqkjHaStWcqjpHyCp9Hj6
ZvgFdNzDUaIbfGF2HQFsmiPki6YRMYxJPYzg6oFtBBIGVqtDlbXHnQagtPwJjAL1mm8P64+r3k89
ZCpXCGkIr1bHBZROkYnVnFHRkdc+FluSwuo7eyAvIOSPonhPqwemBk+4e3pR5YUD5w9/FWKWOPO4
8dMtOUd+5pTHxzDKRok14jUAfy130+ay6dLa6Sf5MIp7UsFyKlT+6XrsRICD69FBMRvAYMEO8bhL
MnVpeqHuZEo0aIqfM8p1qPhVxM1Rs8mgL5cOrIkk5LkUP80YUHwi9qKht+SzVKSuR3UdN5OP68xA
9kSPVoJt/4HgNQWyF3pB5y7IKIG9ljBdCbqOASfvHbK5fpnec3Ai3Id+YuUuiBUBZNi3Egy8+yKn
OIzoMRb+C7xjH/ZoBRjSg6Ni+eOdoXR2JbaHGcUisUwEom8wEa8LvFwfgyEs8M0/Y6+crEQ1ASy1
wqmFVKpsvZxLIyBjW0Lo8aT6ioEC6UeqcDYjHXt4NoB5pfdpAO0Vn5yIElse62o0CYoRoAJzJmWC
sE9USO9TwdVeRgwNlimtKysd7JIVX05rsje792ZZAmlxRcyNEVTlW5fYfNuqtNpkzV0OLnZRshXv
Ioitp6WZA3Sq8H5GGtNLlUuDvOTyxF4ei5QLE4OHH2igR0l4RV0GA10hgLrkE5lMru8rwyIkihvv
LmdIqY/pliL11EOJGHYIDGzjSKJ4VWqvjp/jbUlUMFn1xd3MwK5fioih5rPDGnUwGb00vHU3y3fZ
kg2wPjLLxf7LcY8vFSPwITYjOBmnW4ZxxZM4Sj0QySzwKd9hchlpE/C0lg/yNc08hmCpbIy2d+Bz
8+u/TIpyjs0sNFS4CGbR8uNa8r/dGAXuw/S9JxbQAOnVGvwtEtpN5CaqeKUootat/yguSx5NGQ7e
4GBHywhr87oltL+OAYSbkWi0vhkLVDA9ou4B+RSLC6SsrZm1vviX9bwhzDzU1t0TMwUi6vhSgrE+
0lDuuqA0Iu0X8ilLocgLmmftHHq/+HJKVQfGF6OYjsPjRJ9YzxcytOI0bQ9ZFFQsjrOPum87s5W9
AODMCngfMh6cEEuhlNWOtKcdbRTf/gtEHj+rnolBEBTrRvlqSFyAv61Y5l+szk7sPSHeiTYAkxEr
6VTl8GAt4kWFetzkcTQ16neNxsyq2QxjYx2O4y284EUj2P3h+TkL5l2qrQhaafnp5EBvpLqySD7D
IhFJma6hQxAIuur6BwJyd/o2Q8j8uV3d05lPpAwjkUcztzcJhAR8HEoCyc4gwC0w8XZw/J3F3b2/
PsKyfTQTqkKvkbeYTWhOlPAugSpXTn2Qi+lDADTSUw5iX21BLUzwPlXNP6VJsFl+ZhMl0rv1AanL
nWw1MksmugeAR1pqZtEua2q08pMZIHkl+XAjzv1DUFucuXCdXUAQGle25bjEJC5DkRfGYtQqlP8H
vabAJFJwS0S3EsqoVDGB725QsSofbS3K8ugruW/U3t71GyqR4jgf4SIRF4dWmeYn4lI0zMnEodlI
npk/LEKRgV5SOMv1OElosrNXSwoWbOcXdVJFm5tGSYNEDHBz7rx9tT8Bpwva68GvWIUcWjVPmQ//
n3I+8vxlqWLe64mSlCw1/Vy60jXj9FdddCLz2G025vOImDn/HRXFl/5SSrDz3rI9XE9840ax+fnv
VV/dmC/LSA5rDbRgfrfqML1RA5pPUDaTkkzYg93RUBIbLhIlzTGzLN9Tx9OwSN6EkGMZcnZPlEEe
uclEf8SCh7LWxN4tGHr5YzlPhCDdBTIZ1y/WkMBip94SiRAXkKA8ak4+g28qbhv4pLyOSkJ06bLQ
kRYw3NvbFevcvpPCl/V9EqcP+cnd/xLmOmVcP7yEQUptPBe9CKathT+tb8KJ+LD6tFvd8Lm7zZ7R
4QoDwGUQyT0VFVksBAFRptDWOJy/jePkrzgEAsnEnqA8FNV/BrPLSk98RPetvDT0FJmxZW/t9UXA
s2ocsV6Ea+ijA9c6fkBLA1zCA07P6Xk104V3LVM3UtdPsRuj8Vy7ZcXWZujsHJonZXcJJEyZX6KY
JEuEA6WkVhMIPV2ZonzHqwj0+A7tEKQQHszYj907pAD2oLwSpDKdGKWaL4ctQBk4aqDBSHxPVUTp
YSFlB+kDgYKV/rkgiSAYmeRreAKFUzgaRK4kM+LxQHnzsKnUIPgf96KOnvzJj6Ndd4yHkeDnM9HU
bkcbzWFqzPLU+L3bQCW6F9UPlhKQU5yls5Gu7QPawAiP1dKRf38CE3V4ppqgerdr5cYL8/kJIdcF
swZcv7xAi6NW1JAsoEX6U9EjJb7/z2WMrjojABHDOSPPDDueSNaAxLkUvo6ZONlod1rZmR+Mco9f
wLSwNRsYUZIETSrYv272UnNE4meawv6odErLqCfSLqHdVbJOO1epZVIGS1WCZQS3q2NQRQTbgy2a
zFfbHr9vlDnKQlXgtz+eV70Ey37bgAHjUHXuZzh/g7hoTvVQXzC6J1Ed8TzUl2IAEdbb/BzcW43Z
DTFdtgIgCsQCwPG3jHLPJa9r3KFOK9pEUGqsQXG/q6ekv28VmShOgN535+1Kj4ezUDEMfZWk3cke
R1DmsS1HbOKSesta9fa7GfTvjRkYDN6vFnIhiYVMVASLBOfFrR461VzSEwijT4Wod2G0Ns1KEjYQ
kfE9uYYhWoQMQQrRcBdySgf3TFfZC86PsA+D8eUmq/rzVRKo79BtJ8qat+ZcYNh+NLWyX5f6VgIa
vh32M5y8JPpngmyWFEIylTdgaEKIrO72uvh5+fNMD5Nh+D4aKHq1Jt6SXiUPlZ5NH2la5WQv0bUJ
rnBuR9ej/95E3QljUeI20MSuJentzGfuAKzw2ALADm6xiDFavT+DUGxYKUm4OgFuHMBDTpTZf9/6
KKGo+iMgQFJ4oYy0oDQpLLkLFozQjgD5GcEaqgdhil0jGi1jzikMiWoKAFveVeTUO/ExJqFPWPJM
uFD1u+Tld/FOK5jq0uKNy/UB0JxNHkSmoPkBncoT7iJ7og1C7hQokLpwHb3J0QuyYhHxiHAQD7Uq
X1ZJEyeOehH2ECsMlV0Kse2H/+vdBxxWAdffOFinHyUU4s/WKcAGbPVR6F51kmgQDzoA/v09AP1H
eTxDZamfhBbHjG0Um9jr2e7j9unVD5eV89x5aJjAA3J5Dg79uSHB5969kaHN4w1USeI3Qwfvcbc7
czd+Qn5JHK734vlvgMRvjIdt2PisR5VZDEE8gFCnHVkwMY7yHCijaSwYs35nlLN+r2g2WeR7jUDV
ylL3KD2+SSbOwwA0MMZ11cbdc/6qqCRNox5uihlQco70dhB8aiukdP9ZbplH0Rlu5bpokiE+3ESq
e/rptnbH9jF8XNAxrBXw7OGRm8BMpEtFIK77hqAj3hoENl/M14x8ONEAd4XYmafBzUh8tPfOQt8A
ZnJHFxIxtkc/x/87t1kaKI7L6TwrCfEtBhLOHI0V4ILSoQdycg1712DClpZkGu9gxGQGFdqPYsqO
ywkpig6JBn42dHdg9SnugxYH77UMAi1bFrf5c/nGndsoZ63CUgRJmtlPr/nbnNCjj9ePQXVEtHHy
jvZB3ViO+BEqMXanoT9onw1hJY3g2HhEXqSsLW/Na7X7SGat3wXwGzQl/0U62wTQqPXWq8pi4R3T
dOz6DY3o5uLPDYp9QRcIdosmPQtl++E9SqZ6cRh8K2ePE0Ibm9qMOFJu3i0Sgol/oPo3tTTRfXHh
l71LCVY31W5QHfcuXOHRjZzirRlfIWDU1E7qwlH5DdEy98CnPhLD/AtOLUMvdSQ/JX7zDdN7AFW3
FDamBL9XZga4aK47XFTGmqmtSIVtylNkW7BPSAagoyjWgUroRkdypOiZ+Nd1lx1l5Ej+7IJfXa1J
QiMMrsFm4pSPw8kDyyscwoPxu+kHxLzWGW7rTMr2kqTomXrVw1DOnL+UhHIWEPQOq5Cbc/wIej+7
Og/YiZFWPJcOM1U53idU6fwVBnIDlA2ceEDT+aeV6WSOK5GfUnDRqaX8R24HCN40KkmBXgx8Rpcu
k6V+PFMn8HrQ4QLvKsiwdMOSSmecqRVEkt3yBf9nSwLRPvgth7nqPNzadqBppExMj3ZgMFoCaDxx
qPuW2hzAMhT3NM5AADDHgvLC5AELQqS/BBePOX0qOrM6KrIllDZH60egtSjUlAbdHBVYK0XKpITP
xZKnwC+VF2WG/dOUo4oqkwdJDF37jp40eu2yzns7UxNQeMJlWAGKO9ibMb0BN3aXSYNr7vl8CcRs
il8GxXjgaTCsyP/oLEJD7OsF8AgNdTOzOPCkiAlOH10u39vxOdaI/XLP8T2defkxJpn2Bt72bNiv
7X/0F+R8TNmHt+rvmTQg053qeaAJ8In54uTWLXViykUPng/NJzuGHf3doxAMhiB7/bsLGaqbRhTi
5PzOqDECVDKydPD2dGGVLejAAPMAdgsr0aip+eB/aar9Gqwq5PwinEEuxlvhQs5ePOSCx15mYxFL
qMAalhImayST9D5z4uTiO73OEepOJTE7gWe1YMamcwDL+kol7Wbp9pSFat2M88pW+eDdUmpgsMIw
JuuJTXkoZ/xcOXyXlOT7sPWOwOTGk2m82ARD/9rm+NMx3xmEZ74wSoiB/f9Pkr9eULkrslGm8c5X
kgISU/1DtHepM3fQFAngHRg8mzV4oE527egEIfMTEl+6pczHkECGTwxLoAQS2vTIxJOhTheDTdRy
V4+Je6FPhVFkTHuZQrLm7Ry2TVOLtnKJiLy5mJTme6F3hCl3j0+2Ocra4obGMsrj7hQD8sp3DcKC
mND4ApusAM2F1EXkel0bs28VcdA7uae9wQ6YTrQxriwAHSy/8rheYHsHzVaNzHtgTOyaCYhkEITy
TDTrxKlnsvNNbmM6xyjkEoiwFAcdoCuDs+RIvDJnLEaEvMmhbxy03VEfvnfeD4RP5OB8wuhRc+Q7
24UPwotoQsA+lLwVSMh5eXjDRMT5S9nsB2hWzr2PpnpkVxBODn47j0G5NT/8Zbb9N4A2Xe27+iIO
lEo7xRb9+Yu/4EB9T+Fxb4DhUyL8LyzvlYbJpV1kmBZKvcwo1MvTWipCKCUS2gAU2hJ1ib16YxgA
0ngDw+y1hF0UySWHyfLC9Ldl0o1h+MHCKP3Wk9udiWyAyIyGDpvdMc5oVu+bx41tjwSuTXFCHUos
zKClSEITzC64d0GK7gqQv0DbNSg0e4D7JcRWr2FqRp9r+s3cytcL0avQgR7WH9W/sU1iGX4NFn0m
CowzJVu6YADgdk6i9n56+OWKdqhJNRKM4X++v0fRMKchJ3WaSD/ZQb7vWbDw1yMFE0sRTsNlpf3W
m5tnb30ab5R8AiQ8l/aZWgsc8CKhMzdSHoyNJHC6yVym1Olz6+GYcARzKEUUmXJ2n4zp5RGt8MsB
RNgFjmo2u9zBJedA+zWYUIEYDSwGob9nBgLuETJgUWULhVsgkAGfSUsIeqL1QAqXmQRuWTcdSsKR
ABd6nJCd+HDKIYDb8YpG+WPzoH+Qp6gqKk6qKaEn+zzGZrfyfcK+Pc1O4R9xjBs8lnERPnFbph+j
1KCox6xIA3XbrcaQQ/5vJjaFoSffDVA8AsLKSHVR77SzMu8OieDbGyqPs8sPuS+y4hHpsLLUxA5s
T4VamGuARJfLYrWr78FeG8eiEwOOxvG25ddQeBoNMMErye3QgWQrEgDAknlvlqTzKKjpBa4ESRJe
8obUn8t62nc2OS2/ORGEjjm+LNDpbatG63NE8sZW06OL3+QpDQ01t5kJbkfHggco/eNWzEkH/ptg
fuvKpsrHMYIsjIw5+wauVjzIxR0gFZteo4PPLwjG2+dSN/q/dItj7La8r9mGku6EOKHBTDnMs04/
7hR+z3yIWffaveWaZaYZOCbboIoEnw1Ym9YTBa+u2oBHojf1V2arEEdy4ymy1S2emMKrI4JamErn
UEh71+3oTy7Fz1sauaUJhQdv2rvnvuHzvlSLLD5vJbM7r369P1TnwbnbX8f/fl/ZZsN5QA6Cau2U
b/JoCBRikGNKWfQPxgI8RrqnFd00JamL/OJzXqUGkGnjCtpjZR3rUf6roKSux8K+/qNAP/BH7DnL
9bVo7Y0QsCUF9Tja/Y+/y9QBHZE8Tk+6tlkVCnupQO7BaNsSrQy9x++VnzkahXA+MnPXgrNavQZP
JscQbbV3yc90Qsgg2RzqJwCVVfSJRPhbOl7QGu6Bm2qyZo4Y/rz67W8J3odx0qNLqi9h5Uj51xdR
xtO2lQUQcJka/+Mk4TSWdN410lfpAjdVCDOyErOWEa0FtT/4pm1uyWEu8RtwQaahMGCb8INJTs8l
g3CA2pUifsjQPHLXYNvUfQp7pLDKOOQNMvTUBiTIuw3lZDpdH3GI8UFdnaitpXMl1Iozamp6LOj2
xOPK0aP9XF20+VUs8PBEtyvvPiSYIiJh3w3qe6v8xzdiZNdGUg7QcwA4v58VkINTfC0yr1+eKHs/
BLLMIN3MWo7wJbwIpYQblnToHQXjcOQ8cjdjsVqHq4Dyyit2vS0vXD/xAxEcfKMYmuCOPKZIdG8M
cy+EPEsdpI4Hx9fvAN0awZ3D8Vqt6wqGHnLRs9kYwCwOaP59z0IWdu1sXgUOzGn7Y2eGH+qiJa/1
T9PSS65fLnL7Nm/l5Za7hV4IFeLWcCQhmM67JnIMkm750JNs9jVx0Kz8fwEjKH1byEc6aEVm9LUx
KnNhJjDVYjs0nsWSk03X/Mgpki74qj9OleieyCxKfdmEsA9O0mS+tgdNzwOArsjDadQHLYd8hhTv
Ow4HIvX3DUto8gBHtIcfQ2DjZSIDSrM1mN8b2C0QSOjLoD9hWVo/P5T/dhgktDzu394jVn5caym/
9ZKRvI/G+A90eSpbHsRGwJdZgTGv6EaK/V/QY4vONoKl3CPg2Fj+vCEV0oxhiS5CI9V4U0XPxivq
0xTSLTvYwzGu8XZ0puca942YsbbxHz3UiOjIhOQFOdPVASzsID7c26wC2cbDqgF1WYYImCy4mI+W
3wEWaX1M8EfyBlEy4dOUKi+8cJXQblMjGwxv1bCsVoXlFFPrkcO/8mpRVeq271jr/mqFrkP/NcuU
uxWpJ+vk946Y0vtJ+a8rQrLbuyTUuQ8Kx23Dr9cPKO0T2htZ6nu2AaNmnF/c8XWsxeV+LFs8Zi66
jXYBWsZ2FNXcqyVteYz95/Emb1zxblRxH6yWtAqmLvirr7lmAaJRhxaB/OGDv03N8blIgiegjeNl
b5WwlMQiLj+S56DTFQuIyW6ZoBGIpLjtDSrMCR+hcvlLMBfZpreoRvw0AdKh4EH6aMOpMuQxHhyB
0TPHPQgM4pb/vqRehQ1TzRKUxiWVoAzDQ9HHISl67SLM/jBqXJTmxwj5P4UusnaYiTmEU/Q0Rrgp
PrDyyc4yG/qjgi4XKzCLdEGJXPaWBYPv6NHAy1ZXPECLGhqCVx8UnDEd8m5TZtx79R9iaP6j0ZkU
5MbPE0Foz/guuUaP1s19f829Yz9HjlQhBtx2WWDw0JeRZb/8s60lRfiDNZ1wP3iKs7UDtacwDSfy
iKSEvvowfWiCtnqauwI15g1jcfhol+Zj5JhWVMe7wdTTdLop1S+bNz8PfAuSFq9Pm9+uuYZoQ7Am
E5fWkxw4Krxe8ogOZ7lxBjN0aLKo/WUJCs3bFipVnk0bQu74BujXI/wJY1x9GpBXWx779sw7H+9A
qOpiFGmOdowmt9zJ3UmCyMRU/sPZdtyaryIWBrmlqNoq06cBTmGNALuYx9tlHfClLiqbub64rhbC
41bnRllr9YDGWKlUyoPluVY1iC6+faH16yP+jmQpBf/JBsD2r3PLR/X0onvZTX5691wncEGHMsGt
W8uH6BJpZq6afIs6D570cCbBY/CSTCoZnouapwi2Z9h6TflvY+zWOaoagdxpFee5xNSLAEJRfRcD
A+HERQIPynkAuYkuG8n8hw10y3CgQfOtF6qw2H4mrNEATaUERMeu+SavDORvvSrtS5mLgXmwj7ZD
xiligwtdxqXYZrfwt2Je4dY7vOXrfvqINkSn+E8+PEm1R7B8oQFDH1hN92Iq9pkYMwLKjpCriMoh
mMRTMKixCz72QuznJvyxKBAA2hb2uhzJqqp/LiTMhYwUsfVu9hAJOjOCcnaQv0D5CF4D+bxAyO4m
cx++6lgY1HalRvgNy+QEKBmM2f6BuQsivwbMeK1En6JAN5YMY6YXMWRnZ7FEl27s61nE4myrHwuK
g7yOeXo3IkRefsv4HMHHtKM2xd+BgKK+F2coRM9IE5AIb63uL+j6ivri2uVqQkvML4JJS1CqBlx5
ZpI6DPQfwfTRv7uOxb20c26DDZzcSpEZInuzIlka7ZP48jMQ5ap8SroknkgM4yeIdVStXSq5FTgP
QTkfoVJukK9ebqz0g76/sMCqgIHTNhZoXL8GY/72qYhnkJIkgtkQK9jLWFpc/l4GRW9XeLhYrRgb
ieV+8mDNBaa4JQl7wA20Vd1L8ABVAZNQ06YK/vlA6/eKMxz0BKWSYnYn316KgA3LmYFH/Q+pmElv
Rd8FX/cULnFQJ37OdE+5Wdv5IoJH4K20ZeDwmgAARgKZ7TVnoQNnnhv5NV1fWc4QiY3Zgc/A9AKu
dmXazr0q2UDyHuecRKVmohs3ehMY0tRSRDiUc08De/4n/f59nMDEkTp6Od7z+19VqPwTGGgLY1ej
855jfvAr6b20ZKsfrehoEX/W90/9AgHT3toxDOxKcwyzczaASQpNv3Q7AxApPWR6TIFkf4mn+UjH
FGzuWAmaJcSGyzIhdhm1VxjAY2ZK6ADQQ9dkM1VKpnMwePy7ci8azDfU1q36CfDFeUrpFjjMbQwp
raSAdtUJIkLv/BbiRKE8a7HgG0ksb7k6FMf/jVvJADeN3rLr5OSIE+igPZ8GskWR34h795Tr9G0n
EdVmpvYJuAUayBELKUxvOHJsvb6iMbfgICItWL3BSOwv0MZbhSbnWCeuDPwlRKj7DMdRs4L3MwKj
acvEQkIZuGRpU63MsIxfWua2vm3y0d/VfnqF4gxjxCHWhswwsn1djXMj8BV7IThcz+EC/p762mba
W2q5QJVH8hYWrSU+5tPi1MCkI2gdFsB0piiZQ+tZ6CDPYEXdOiO8KKRMkIG/PUJpwoFFnnjdU74H
XH3PFy/Z6fNdPhpNbv+6zJAGqu6id0yB7fwa6QR+amp+oUV0Jp1Db0MZfJOlmy9yKrN+zT67JImp
PN96Xr6Smg6gleJboqvNlbtsKYtn29aMzB42Jr/mqSpxB7sndhb+9Pj1r1WKjimCdTC17ZUdk5VI
VpDghWudeZ1b2CrNLFrmOcJX4jJrkqD+SBP54BnK+0oX4VwhR4EZoNDbCGR/zME3+L3SSCkEJ5YT
++F5V20S9MFMUjyS/GOuav6+X9ZmAi6gNJ+abIBm/UmCWXAyd2IkpNvpOf9wTMcUV8RB6A5vkMQs
O3GJv7H+RX3O+V3s6qj7f3k9L2Q98czBX4dmhEPyN5CCwg3P8RVmdALWFz4XlF9Rj1y1rrm9UdGQ
/4NRTgeBg385wZw0bBtIraLE0m0rJI7zmdkQ3yUmkRyDDhoMX6KOR/Bg2Rf0tS8aXMHP56n0KGXB
0Trlz1ojax802fEco+9nONJkTR0R2T3XDjh2U7u9SoF5MypJszyH6DkgLoTRj21I4G3NQcMphS5f
IPv5CX5AfqG6urtBQKGABS36DklseLMyzDytODFgMveQ32McFktOkN5P5UWN+dhUDIK+MoV5BbYI
PY4Wq613aROFgHHFcNRQkUBL7d4cUIN39xwMqW43dbf2nKqbo/j0YlYmx5R+AHO9kat8tJ5Uhuic
rB9DjUgZo0+Nr9s7bCHs/QVIHy1JK0kSyJztOMtnsMvaSeNRdEl/lcRMK1GRo+LbOCnxCW5POS15
WB/eq7CltO+sOJZU08rbV5MHDShWBZQR6auaU6gC6yHP0cIzPwgh4StZh6HG9asqNG7kgm2tHexJ
fHVqw+hWpArBLy2afNc9oMvFDStFB54+/ufnJSpGHeffZpQwNAW/+att8/UvrQfgcq5NpBInCsQb
K4oFTTzMdHiq24j33w4SylNnCCRQpzrmiMorDXRhaNHAQZNA2cMe7V9/ZGJrxsEmsBJqNYIXKiXh
bH+61M47Ozx+nrlhLnqNLaGllGJBe9R/Fp5yWSWKYEsVopvNDNZwxYw/wrIx2CC4TM2BSiWfvk2S
IO+qG0l51hBca4VV+oKdbkONhd+ROBFqC0qkM7Beq83msWSea7k1UitnJZSRfOpwt7EoBMX/6Mkf
z6RInbt58MZsHQu1kQwOKAyNB/YlxanrWvfS2Nfe+Suzs89vUmSQoHuTFwO4smLJCPRHShIhb8kJ
FgSlwQ71vvDP1hdRgTInw88jBlWCZIMdIkapisCraJkcVcxA72zeJVqTSsdi4VbctxPYUeNDshlc
ISqG3LZvkWZVtlKiNC5v1v1mCVELr2QHTs3kgCGmCKojctrVzyFvIhVo7Fo2dCR9ISJeblKBvcNS
i7bsrO9zwcpja5tgix1dfTDtepGb/Amfayy+1DBBlqtsvVP6G8Yzgzv09DG0zVDXO6/7++P5i6TY
KkPkz6nBiEOWfelf7rC5FcMZ+r1ZEIzoIp8oSBhyaoOFv9gYLo9K67+871KbogKVP0VbBOMJkia9
/DSaYKtHQMVsBSHX0pxSyLKk4I0Mzf4A3V0gb7/lynox6oXp13DrxUlM9nMFRvbQHlQA3FkcTc5q
LCz8GAUeHSp69UbOWytZ9+1rO/3PpqOPn2lzZoNF6TXAnleGiDDQVOLbNfAfm92RCntkBttrBLNp
LKN701M546XyOezvQRHabs+yUPxXD1uOuau2GjO4jcTlTnEw3ImWIzv3El/neLCe9cUf6y1S1Ozx
0brEQXh4wdw9TNbRZ+U1PobPnLXWy635rapMAW94m/sc4qxHt9VHX29jELouqutiShGmnzWh5YBn
i9A4FXMhYP5/jKbsitJ7HHSOAUOv7Bx67rlzUcsLwSI38+WkRxEKIJtW8g74c8eyhEItIbC+oPlc
wRAqMMjGgsQ8ecg7a/Ve5R7e5Pgdf/iZfqs8jHcpU22EexHOeNyEjMmf8ooX27993a1tQU4JTbwt
uzYZUQyCswqdY1pTScuF5zVTIuceMNMpo5a8rTnQnwLCLNWVj0BsE7+YkYGR+lmq08rEuA84kvnI
FfpoR6kblQPKPnRY6qqF8NsHJZGRjyK4rQ88o8wkIQCN7cuOwiyAQJkM4xCAkYmQBQNxBPdYdpWn
fA+zADia0JbCyPYMPL9d4BUUOw6qz/4d8hkarIGqY71DXUHNtwaZTRQVn0WVAOxUAqF0tUiLjh9p
ctPCb9v3aN0jkLjUEBu9FNwaaZ5qForw9W4Waej68YtfWeIJymyp0uJaJ+rI334HYbN9F3pw9qOO
OuLfpxgnY7LKJ+iKzZRFBUpLxq0RlEy4OWQSBn6PoGCE7wgtTGoM8BYEOOcql0NgYNNYB/+rYFHs
wyVOXhwQCiHKwSNq6msfNbqQbHbiEqWG1Qy6eYVb1TwPdGhg9r8rFQlEesSPc2BBn1Ueepl89DpK
tR3L+x6yF/K34vfgi0egoS2Z6uhrTCPzcI9wbltZsrNP7NszCSkx7Mj/DU5zTWYiUrOJVKynmDLv
FChMgUe+5ekKYemmW3OB+FkxtCP1+uIMousyAsk0QmW+/Yk0oaIMuWUnookUD0A2+zcdxuKlNWGw
/SV+APOgrOt95/6+WrOr85jvjWfAYBWTUftl/yDMKsOrUmYVz64eKffN4zHKjvhufds9xcsWE2bA
2nDRBtCeYx9jpbJ1Tb7DgZBAFo1EcUq1EP4sho6M01AOO2KWh4XSjhU682yMctiuUpeDo6V62ZIr
XCDRWLclSZACJJA1jyBcItHooTJdBAUlBvOe4BqcmH0wg/9hahnwE5gbPr/qSVTZjNrK56eA2LeW
3Ep/CGpgQqc7qf9NBdpEr82kyX6/vQDHQY3V8YGuihdIbhbSW72bKpfADixiYsFVp/SQowejdpQl
RrmLkHyECBm2m/guWEbPpTt8b7NL+WW/8DFgDN+UYC0d5P7CVCtZFIsSenBU7r0lQeGroIWQ7ePT
N5VpJOh6AtB3LLSHQhBwMdxH1eGtQME6h+oiCB2eEN4tbQC+kjEYBDVJZz4B8DthC/REDr/xvLM1
dvQk/+1zM1cJCezuF5O6yVCI+/Cp4vZT1EyZzGsXXAn6ZiRKTJJs79QET8niYNoMgLJlgZpXnII1
E+vU/h2Yf9GmdKJR+BzyN+aM3y+jpzJZMW/EiqWV84srADsGjILXy5II94o0r3DizM3UMmD0wOGc
0lwmCkVQRj9C3J16zUtcb3XALmq1lS+ff8RUzdnAQS5b1zr0LPMQw10t0sz6zX7k/g0zDPobgon5
FUR9LRyT/+hPGxaryjTiFFO5yB/xANPN+zM6FOrSdg32+XoTHtK25LKezYCRNdynzs7VOQwFxaYw
no4VV/nPsmOrvs0WFKFbgQKmzNBw2SFvKC7oSjrYUJGlMeGDrxRh/6SZT0BQ9k3XB/97tFMNN6Pf
Xk2VU9onQDvaxDvGJRsZ0oVPeYqdhz9YODh0WgI479ULm72w8wHqst7ENtefi/JlXv7lS4U2UkMg
CkLq2rexe6BEHW/FMDzSdoQn0hDLKXPfUSe0O2U2JHfX7tbESgSmkFc220M5+/yqBNR4A3h/TMx0
qwux7zp/TJbFP7J1JbJg+ykrOBCQZouVeSbD7XWGQK9miB1IfNssHE8wd45Voel6GzlYGxHZx8dN
hMeDJGzeoBKXj513OYgQl6eQcMwskNYPGq1uu/JCASijDg+aYzoqqo0pTF+zWYi7kRJUrAyVPKSI
Rj7Run7QJ4as/D8+OXfEQFZDy6p337enXHuV9pz1hGDf0CJE+xpLRMs8CuyNnqNbkr9RWchWjlgp
80wYI/ZNhHq0eGJmaVS4gAkdnowHUtQDOhqnav6zZ9sNa12pbu2Y+JCnyFMRfHON+6RpIMGSgJJh
UwfuvMdUoFmRubXLLI/amOzvcun1/L0EsghjsWY5ja6jczObGxwuFIyut01P825lWfNJqVEOvZ9x
sUNH8yHGwzmmP74yIgbqbsUAWdkQibmq3CnUO9LD4NBoOkJSyByH78/tWyXknzBtROJNCHHTs7lm
Iv2t9pVXVnKH+6mmgZGcWnLpEhE/pyOv/e4XYmMRMKN3zLd4VIJTk5I0MKRdm6pxb9/hQHkZTgKP
R++YkWBeb6vxR0eYlWIEkVo2vlObSel6UEbPdviTBaI9gnvj+DK0ndPKuWWzUm4/SrAE/CfAswtg
Pp+VKesomPHiHUGC8RgM3NACvt2d7ZkM0CCpga4oFF9FxSC1hQ3aiOjp5hOAX/0cjb28DufCmNfh
feZbupJL+WTogP1GZJa8DgWahbJeRAuk0DktfexWoSiyBQJfRT9kHJVUs4tUg6HcWwnvadwj6QO2
fNR3yW9MIcX6+/aCCc3oAmqUVz4paX3/xAYu+BP/8ogs1/fpN628yb+Q80uCjN4m7U7C7GIXkZMC
fPy/tDFTwJviIPR8yvP7KayC/3a2HstDG/rhwiL+2hDBPg/PPM2/f1WSGt9wIB3sr23pj5ElA60S
xfsDBfg0dXUVCmv97E1bf7Z3j16OQ8XROtqccF3tUEYB+rpFfKb85L/95XygDnd6pNXBfO7JJBSk
r8tbRIM27EjFwdZ6EoBXH5geQ2Qmww5D1o9q0z8CbB7F1D6ghrGtzIhWPSjbQUMMkrwE1MfTPuML
PIKtm5qw8ne0SEL5/+gQmW6KvHUp7rRRCaJMpwMu6qpQOY4WTrdJidwVTy8tQKJCWjnlmaWPTuX9
Zh3CK4ILrXYj9euv/EcMUEoennfUNazS9pydYTkv/fmn2OeiRfDhAuOSg9Bdw/TcvqgRabSaxESu
bYu8a3lNeWB6YdK0j3vmnW5cC5JR0LDaHtiit/vCIc2OPebz0vcVYvjS87DtLkyG/NenICcIriKj
SIbk1PEcfxHZR6FnMv5uSa2egRjblqbSs3DKhh9Bf520SfCUcnuW4yLH1n5VzllWj86ItKDZWOFb
yAIOEgkx0tMdMT85Ie7nYsXL6/r3LJF5oc785Mp1yyCJWmsQfKm2cQEh8hVnhbujSl8CQFoVKfzg
bc0CaQyiSy2Hw+B2NiTkX9uBxS8h98AL71OuD56WpEWxdIMnNOsw34+ArsqhGExa4rHOTv5TuEgF
4/CrSpmA8fWGXRzIBWSY0+dR4IxUQwUkkdofvvNmggP+B2Ks6s1SvpE9nueN0csv2OMZYDscYbz6
pJ/iFxil2ntTzUG84hpx6abXjBw4FEfg+iRVi0v3z7G6M/j8z0DAbjA3P5VyWqrNpOtHXQhkgXoj
8c3GyHduQ21756ZLGuGWARC91/TYLBCnNZvVZ4KTiGhO8jlVGQP4k+zY6uvhUwEbS8y9UcDWGVma
sKVn97eQA54g9vamDtD6yIbeEBCVaU2mt11yh67XtHdocxnsD7+m/hH0KPqZoUV1STOIi/xLQ/nz
dfrzps1uuaTsHkhbRa4G7HYGU6nRhBVvZLzCCIMutsrDWF3ECXtn3QPTo/LWchUpav4mW9fwDsEM
Msr0JqP6Ce7a8ybl0ua88m10N8S0L6WpTp0UXYUJZpiWuYrx7DzOadOpJ9fBey3Oe6DPY/k/h4bx
fjH4NgOExswbQ9vYkTh2YjAeUk9m7f6Peom4TRvxmwOR+isKtD8/oLKITAQ6jk7ZXN8TEorhc1O8
NpXrsEuaqGlO0CNNN+hZHP4tIte40hmxHg5saGN1oh3XjS8LIrp3RHpF+/wEMCvz5ncijHrGx/dW
Tcedw32ZIkUE+YgN7W69VU6tgzFzrwI1I79KxFRQ76RrNaMnPGq+m9iOp64wmuayF402BOAWEwBJ
o7For0/Ht2d6TiuakRx7Ex80m+bUJOV5KsBadC0JH1pOCeu0uW+KremeZTIEJguXuaC6YjfuqfUU
ctquZUmdCpFBadgNwvC3fk3URMnC9FlIW4mFy2z7JIMvlCNtBFfDeD+n4+YjuBpmMB0LlM0+Hog+
q7wmWKe9JCLFWGaBsU1oM8mGxz+XKipVnT0+qVPzsSkhlwPbFDVPueRfBWYfZyjI1O31uD1ltscD
yzxLvMQiBN+jpT+U5c3Vd67JzbSsHPVT5FRKS9ajw53NADOBUfJvoNqxAAzEOGtnNmuN+HJukFNH
ZjsFceY9NgU+TqVzE25BVZexHlSFyhNRhRb3VCeYS4yJMqvO1J1FeUoVnd/Zz55TW57OHrhWGR8Z
dKAqfKQ1P1+/c7n+jXxwU8BgDo201e26GU3zWRNbPCRw6elJSl6SoZeGw03YyQzalXJvzdNjXV2X
u+qaCbdABTT1JUqwD4A5OhgAz6xEPdVR1ZFiAae9FddHv8f05iYSLo/DWQa0GM9BfkFJ8h/0Cc9+
HsHQSgz18SQ5gjItMT1fmIlXJ2eqpLhGWW9BXrGPxlUr2ZN83nXOk36hMeattTUihJxxd1KDwFU+
+eFT4GOEX3ai7vzdJNPSVq6TdR/5bZZvRo/W70JFmL2jKEveGX8xyU/g6uJUXmHyTqgFWd2KifKY
86kvPeSHu8XVrquVe8ohHFG6HefRZY3y8G8RfmU4oArcdk2aRZvsbyWLG02HPxqwmumUSYN9Rk06
MsdIh/4EPOKURi2pfYf5o4CI+vPYTqNsA9gDR4rHOwtYn8LMcIEKuNjquczn+IXH6MNtgQ+b0rBs
38jPICCjUIOTPtahlxO5oYqirELGElnjYy+fZS9jGbjEPr/H8CxGRHDTqfxGmclGrKskqqWAKRD/
WfjAeEpkLBm3bzqL3q/v0bwHSKAqDJz8BJHQD8d2gOKlHrNei3cGrAoUH2l6GoqHjqBQfo8KhgzB
WZLskqF2gcr2lSukIOk3AA2wdlFu/ZWhjswflmisQfW7oLilfDN8QSpHLak/gSDi71c2wuKKQaJm
l89X4wWR+rfnS9uvmC4BBnYq48u89YYFl5Ra2vGLwEMdStyDmdVyQFqXpR/L97lJFVxxdjbKY0h7
56GXlBqIs/Hl0Plau2UVjOiw4wjBatxI2I830aPiirtMcKrzsCtqBNrTxd+SqDWNUsgxkrvee8FE
3Zk1TxDzszFt0nX0tF2nRilCJkLZVHJsw1H9PkSWGpuXf+stIdZchLdJ1FWDEHL/A9Ur4jCp53Q+
1+zSIMAeQp9Zl4nq1pl7kZCq6zYnfn7srde1dChp1q029Y79jYfnHQKfTpG+FQhkT+Rndpj75i2p
WgV9Dm8b8hqiOcT/8NmHjOE9JW1DRJh1eZhFfyKF0RqU+fCh61ccDo/xf2Ud4aow9BGy8feI65ww
FWYCqsTA1+ebYcrwNstlQJ4lSagrNRoVBK2bSHHpl26ixBYz0SifBqGyrW8VQ39BmPjGTn4VW5qa
RMsiK7kZgHdi7p8OaLG5Qex/LWpNU7nF2nAOP/Il6puJ0Qh24TmvFVQSi1w4fm6COEBJE0iIlsrX
DE3vQElAQ2BeEqLmZux372JkG5EpKjckouYHkJ5GMCk8ieW7uwmWJgkxSEXJq/C2LGqsXCV7QQr/
u3EIjpWrWOtLMHsquhgWdpzHWaHJACqlUmRQd+w3O/wK3ZUll4pgi9djbFi6Tul6bkLmvnGSqb9y
J9AIvrG0iXj8Vp7s69HJYB+Qvp2YOzYHaDkMG7MbgrxwngzCwQeNfq+WQ+9HMqpfnweSELrZKSDo
ssn1vHbWOgdoQkl4QXNF92VC2lG3oHz96iQiaU+SLzAZNeSsJ765lPclq1uYU3eQPhS+yIuT/1bl
vwtE0srGgriONZsy4X2142cCEL/LFepZZ7wb4jj//Um7n571PRdGOtkzXqVX2yYZvcwm4G51Iad6
B3wqSfbjOSby9gazD7gyUoPltchMXZFjyL6PqlAu6bnVuXy7W4yeF4qQ813qvEApf8E34Bi5hFFY
cDwBj5C/l8JYVEJbvhpX4ygQpObiZVNlfu1iHlN7C3eyDJGM5mkJPsNOH6Ke9FbvGI9YQqKjBVnz
fcSQPaRqsN47hf4yf9d8qlNEk3dLmNpohMZKTtdjTuR9YLiPtwlEvNYcGjGvf3B4HHmPS/IkSJZb
wvXubyAKAGXveQ/pq/Ae648UPd56ky19KxTPqE4Y2Ja+FsNUJYKwz4NfL7gx8sedp7TmgkIDxRUr
pPcPeyZsb9W62uekKC52MZH46Rh+7iqo4uegcMqSwiMKhjMNfJskeEuJO6OTeIB5fZgWyhDDuMnW
d/YfYtXXz9JWgjoDOCemgMaAAKdHVpgH5qIY+Nqq1fhwgVPIBVjfnfD5c+JjhZCvTROz1Aqasbuw
JjQ6qQzEJm3ZKyGPb9j8cUj7PFcGiCKhQl6d8Gbnv/oOQFdCbOvm+rYFl/mjB/JRE8YP+S3GN08u
ierqkMfuwLOiQNvLuio7gCcLnSc/2WnvCu0S1atJEMM2CpDWUutHkI5ttIawl2J3Sa4Ygd/htuQG
hEPzRFpLRYhzjUbww3pJUwV13N1r/JJH6mvPeeJ+gqnnt+ZA+xje9dpN2jo5CflKRXWf++H7L11D
IVe6apcTWCsVrY4+kwUkOqpffJ89CTi3eSnuXmEVn+sxlaaaaguhLCbIqyPSiV7vC4wDjk3//sUE
wpkgZwUlyqoOMRHxmWM9+oSKvB5KympGQckMrLM0oETST7zJevCx/f/L2b1b3JhbipVx1RKY4OMW
ul6P7wavkpnzrndd/MO3b2NJZVZuLo5yBkYLBXvKfydkXQlxSmJr0BnoKAmISNpq6H6OAaEvpfJw
bQtFZH4AQqx73SFCTzIc2Yeibmqz16tLLfAHsQptVFlfSy3seBXlKFfQgExffltGnzpgeKmoGNpf
+0Fr0Ap7yMugQvLdrl5IbgQw4fBHVXNvjgvtHa6T8dVs/hZ2ONZJKrtYl1/ADSc/sBleh+IaiWWE
wwP+yw+DbsvN/aRzopm9u9Hgusz2UpDFILcPC7wJMMxWrjBG1puihXW/iBdLCxRb3/pCltlwUcVv
TfYD6no2O8tXNYI5AzT60KnLcYF2EJuOz5m39NDaDgY6uSKNYcT4rNX5r1wxQ6+htu8Qa0dYr/+B
AG9vNMoaR93p3/2wCKk2Nre6oNcZa5ehGOMtVywv5SrDsFYA5jS8Au/aYZaRgokjDGYrhd+YuK4D
Wj2Cj1O0uFHZ2twy7ryLtytN9S3ISSIb9P4hoSfz7PvZISqcAOxtMzRx2OIVRxhloOtNS6v8UMCO
pWl+W+3954uvRPDd6+f5j/3O2E1aFX+1WX9Qw7lgkeTnCd4r1Qfzlrygy6mkp9RO2f/6bjyUT4/L
ljcMrrb9vi6LkQkmnDa2JyW9xoa+6Op54yc6y9V2tgzb23OW1R5ju2T3vjTayiSiPKDoPQjEpVu1
5Y2SXBW632fJXN7iDHcjpt+pCAVrjwH5huypmcDzx/fUrLtZ/B+AvkMSaUfwQiqK6KCla063aBPK
/wdePIQ9Sj3UNr5RZVOYKgz0mlmpze64lH2nGiZSNFfG+gvEbPwYHnRmWRZP0VFzuJ7Pc3RO45zD
zAZ8YChWrmGAgN7n+H794RttacUoC1DJzN592kpL4/eo9f3BFTQaWPE0/wnULSQcMmTW9nq911Sa
o98fA3Q8R7ti0XQSHPSWK7F22DmDr6Ef+ie0WE3oMDPgCowQqpJMk/U9AZpY3Bsz2pLPWQKdh9Jq
neWTW2WkOV+33ehoVX4e8j3owMgSwfvXYNbEiJ43PsJvcUXmhVn82iGitPenB93hpBnnbaccYIS4
/GXRRm2nhqA0esRbi8R81jpqSdzS+8zOKlVftwxhJC5SAt8fujGS1iFNyGbAcP9W9dUuvwVjqmf7
S5EgJieYzg7aLqbUfD48JTZnT+Nlx6tSuCj609zO742/0MsBvP80iuM/nzcz9uKi7xavuFZ1NuAg
eH3BxrhwQcf5cidaOHlAQN/7QN8MHat7aqyxW1ydiV+VdPDM+rpZdkOp2NmEGvywlx+UfRGqwFXD
KzMWMJ41awPKncKVwr3KySg3oVMuqnUZ3Rm/7uHPSPHP6kGunxIJgCqLE9++DR9+lhZhrHZPjqRJ
0GW7R+pmEPVwMGEKhinlhvDdwb7IntZZruo6z/clUQwkb4GdTxez+VKcd3uixF7DnXiF0RYSGRG/
k6Yf2dASZDINSsPzYSmI+PaHVu1IL/fiGHoq9tKErva20FTpm5KUJWfy9/SGKkE9iE5y4QenYK+6
SWDSrf/urPk+HuVKGjvR7JXT024TOfatI7CUybTKIywU97uUxXOaJPDjIYF4XtNN55nNjCs4LJNa
NeBqKizIvVfWXeoVRwCtYAgAQL64fQbtOlYktAP2eWTODFjCocavWh6emVlytkUHBO+B8IU0rxAl
m/VEKES0SjIKtP0LP6G3nr+mofLFFZd1Hjot06KvWiDd1cM5Nwr6eRqSbeDZdhotPGKYCCKMU/rh
QJQCla4SMxlwNl5Rrd1xTzkki4tk/XXa+8eHVL/uyNkmzgtqT0tLXL/hSDW/SNRrbCJBncnwOzgm
9JkpWjqF63/LE3BAgODY3+psd2I5kxeg9UghF3QG2s5Mn2dnHyXoBHaA0+XPKia9Ylo+w2isOcQU
bxwQVkTpN34eWiLV9ovPg7JvsccBhEHvhMT/7651r45GFPuoB4d6+5olGRneVZiju4aP/y8a22Uz
szOwRKwhELKbQ2m0OqWtghvCP1+XesJkxT9iLMtbKM3qHzBe+N9NjV5p+xhm6S96ZalH8FTSY6uw
Sow9H1VrgbgTFp5Qy4uLvgXjIbtm+U3YO3CNY7xARo02KYUasXPvt3kSKiFWDU0VlSxvpzoo2onv
C25tUzpzGakW2P/KlTVE5u3xG/Lwlp4AxwOBjm0DZhQ07YLKRQkjbazVc8/JZdggyxZ8Q05xe+r5
K0ysIG2rKTEkjCAuhJOclI39CCGv9HUvoab5yKPftM7laKTxeL7uUPkPxcYz3+7ZRKW3HR1Xjujo
CdWdV5PnEh5ikEbKxqVAO3q6aUNpzaGjkAaNZEdoLyWzDr7gEgwMVXJoWMUs5i2AnKUc+D82tGNq
WTNnYpN9pmnz3xzIhwUiLBM6AmK+J0eTXqqaFyoRpTIwra4oJcGGYyZOc/HIZ3DiuofswIJxOlAh
ZwI+proZCpZnSZvJ39rvj2FUIwZgmD8/vSRcoSRBRCvLNAa1LNT8u4iCx9Y45L/jf7bRzT1AGeG5
jvdAUB053Ps5S9eSpAhlcJTR9Rujby8Fto7TJqSnH6rdFyT4Q9lK09dOgkop43QOLQwPI2V1K/my
d07c5Qx8qaku3z7JvIupljU5/YeWvTTVyWN5HCC+sjmEcRYyPWhDfpQV+19Z2DZ2wS0cGxFGiXJH
IgOZh8cX2vEYAOIqs4QihCd4kPb1apDoibQTbdKj0ZG4HKsVTrMCcZ87Su8N6vg4E3p6iSiIihwY
h9Ljxhg89J4BBvTcWQ7m+R0izQ3FE/3MtheffUlpc6lbEMBH7qmwfDLJb/57hh+ikM9N6igJrLpV
19gKvLeT6BEOXqJXHsTvZbpN4frNul2H6t/9eiQVd6ye5jKVM82BIZqhTOXVWKrgx9dn/u84C2da
KEceS0btsnBwKb6sodEvnHkEshNwg5U5ArK0Ywa2caFv4yzAq+OIHfw0IOtPYGFJaE/D542BrSPf
U16FuY1nzteA5WY/CYC90Y/mTZwTu0j8asKfgEmQAkbaIn2ZsIkJft0LAMvOgKEIAmJz+XjfTR1v
t5VyOEKVD5yK5DAzIggxXXtovvt+CjF5OsYXQfEHPHz3Lj7K41/G5bIFerj3YGuIUveGUHzajaQ8
dGAC2uNoGvbKWFATwp0hR70Zd0XC0BJxFEJJmQ6RlqQpogIUXy+IE39l5CI62sxJtRto0nL47L5K
vkeRR6rvLXsiTOidRyEVCM9Ouxteb3H54lc1SD/lSoB8a7j97CDTPfR/e4CxKpLwApVAh/L2AuWw
mnKZ32z0J+6UzoqF6lIgtjTYxy76mzE71MolIx4r3M1nWnDPUhkmwj8gucxSUXYpQbDz886X5SNc
L8E+PZytVA+0wunBw8zJ6yHu8FQ/MlxUMK+is8V86cj2Tr9JoYlneDnh3gaOl/yVbn1gbOJLzpeT
DgCyvbZ6uS4zqTVHHnR2Janv3ADeEJ5DXELv499wDTWYTiTmzELzR21oc53si4Ju9pEhJGzQBxOj
iMrROkfLk2EppClw5RStp8veko5yPxBQWLOAK5teSj2f4TGaxhldwtA6yWe1RvQeK+A45/2Xls4u
qC6gy+wV5IY7xPQTpEl4oRLfelURqVMyZRGTwzj0azyEYWgOBABcUag4rLkEKRZHWvc8e30odlPR
UyK8w57CnIo/oFmRDk6OzguMlLNxgWWRwQCzhEGtoiBNcZ+qf82//tmkWqFXXgkqu5u+/EvX98eO
CtYDbFcKwv6UIjyEAqMPPKXDwEP9N4ZXWabTEef9gi4fKEbzTwos6ybih5XL2xfrS/SJDHD28syA
X2dGxdmSYVxAZOdiakPpw2gxuZU2sLW+I/bd0XcqvjjhG+EC0WXvV9+pA3k7xJxhz9fJLjlh8Miy
rakPwDyTooOaRI1GftYFdeigL2xqR0BO+Y+MbxiD5sCVlsOausa9zQ1uvGIb7WIisLznNLkKGIGd
jEkByOOHHBTQDKMSPNfY8IpfSjYqYSf9COBt/ErRhjjbs/fI9rlrhZX5nb9Q21FBcLIcDsAGifxN
g08GBbd96c57htOj/VeZsTdpsgK9GYUOR9ClCl2PWdzNe4iDMwgikVd1l13XlIeFOeOtP1xqHQ5D
0YY4GLZZp0Xv+xMWp5D6WrW9n2EphJmSfxXp0FooNZpK9islnThh3JyXwTqTfR2Io7L6arZCPCKf
t2qeLjhzrUcIaUZWRbIDMssPYOwKUi7gR8BcB+k/tZwUg2HT3SxEo/zxgtugdvRLbUk/D6uN9+03
kuOUW4BAaAlZ4wOYGkTyQZnzgWhPJAnNCizNtx6oiqRO0ujCwR5Uow7S4NPOhmmmVTacXlkRno9e
6Wjz+NWUT7tCUn03xxe47hQiyyeqmsax51LZo2xdcXQos3Vv8ZCftgaNlMh+9ce4eEIBFN0gt4Od
8B9O3rtP6eQjBxEcxWtHZ4YaFsYGdcR3GL+a0gF/QYnTwNkvMhbGqntc0ZEy9Tm6H1HWyXLnaBMl
qJc+g5QdvpIO7z9FacNuBxxDMraPY97PuxyqNL7lEk5fUtOeUb7nasz8OdGhuLN09I2y5ohO30zR
bQIPBfKSJ+MCWx7ueyquvs9Qfwu4i/irE1skxaxEaMucDEKOJNrGXYoUqsNw7gxWErS6R1aYtGfV
FBrJ4F5O0wDpcm1UOixrGmCek6tb27hqJtfjEA9LpD1MEbPDmJGOfMQN8CTOC6y52V5n6PBNcnFZ
618b44k90CUOINu4vVOtzs2o65EJA0C3EdTf8atF4yCv36rKPKDM8M0Cy+Rufdmx0pP9M2whubyM
ec2TwazJapF0pvIKHkc43VuGI1zRWJ8XHLM7g3RCKlEFHu2uJVjQqKwP/EjYAxJE1SM5u13xPGa+
sfJyPYlYW2FFhHOf5VSEC6WM9WdzIhkCIQl1K0D4Usv0eGaE4D8muV4kYhpfRXolk5ReIKkMNVql
nXB5FzpHdy+7Ie4OXtokkNbWc9JtEV6Mj/qAU07GM9l50m1lDTyVj6fV09TC5u+xyLDfIhUjhWRZ
Z6/U0KL6f1SuQUoLf9VS3HO1IINLVeONNPKY89gvj+wRGI62KV5GhtDcoWuD2HYOyEkIbEtpw2wi
MxabLt2pcrqshYk3SMapBGs9ctOtklmpKhBApKc5/Pl4rM2RW96RN1mb3CFiJ31BMLaxLHB9NMok
FCSq+qxOgPnK6LvabOSvkiMmuw/cVDLvvamleIMIzddUjyyfNaS2uMdTp5Sgjm9rivcwVfcXW2fX
vusUp9XzMeN6nvmVO25OAJgO3VehiakaBrkewC+xS3f2uQW0blm9D2KT6U3nls8NaVV9yUMOQern
iLonNh14pXR9Ue8VQkKBAwIha4dZ8tAzZm8ZrjgGVw0Pcd+cPnva7oZ2YWhPOQiPhVVP6gX7wlum
iQ1QkzQ2ZoaBmZdpOEpFdaRfaewPqnQu7u36xt1iLn1BvABf/7/Ngl7xaNFPfsx7Yiq/xS/a1NEL
TTv4CKMQWRGSF98QOj8n0sG4yAh9gx7xkavCe++MQlikFrvcullyG4uh+2/kjlVZbrGpxLOS9rqD
kXI81gjsR07fNbeF1KK/MUKz25iLGZAPhKNUpOEAaWkUc0ZMjsO9aSXqIa6o65ELp6wHtCEDeIZq
uAK/hrFV4rzOVMY5q720gT3I0f0MCfwF47ENWJHsK/I235dyQpjX+6NAmk8WtVEpijdLQ/zFbJl/
LLntEVQTB28G+eIRQRyY32tmxFd8jofzdWWyPD5JEeNB6Mx7SmjAEOSE8TcxbtrFNdWzUWV7gahI
e9qOEvo+xky+lnxBBf3Sum/HCp+f+KHWKLoRS0yGPS21vFg5pu3TpbwNCkgOfp5gddknaEHhZ/hA
oTAs5ePQx/hJN1ARNpzfxLIZ0apPZg7GZnezkm697lWjZ32My/o1e2LzY3DOBdIYlvKPXBb7mMT4
SP6/BZHuivKD2gXVfmGWCfhBYprjQMucR3t2Whvwxmg1e1sBzcLhpfAqnRxteZrWfpvbF1vBRuaw
TROXxTknBVJe5/gQRWE9HdIfDLds/j2B6gEoCN3dH7oT8oxtcE7sIERK92kDdYfWgw7F9825a5P0
qYsttWSBZfhTAvfuIIqzhARr65GBXVpdRjOScZwUz8npHgKVPvTlSXMhQ+FTzAaAiJsnEa3FY8qc
2k4eFT1cQt9m8DvLBWjvVUiF//u7zhKS7xix2FYvFfDLXrANRD6GVndqGeKmkkCVZRGB/OGMsreo
xxM32Y7kY0eMcp5zGuZA9QWw5w6La0gMK9hRNkSBJgVMMFNcrLOuhKH/BXPHU1mRvCqC074VBAUg
z13QhNtF2sWIloaqJqBlc3ICwU/QCIS7npvjAgqWyYxLEzVGPfs+F9r4TihoNaC/+uk9H+cHNcky
IIBIiLfwnqMG4kOgtEB0YfqFpnPn4I7mVpdW6smZJY5tYlYZLq/8Fs160Kl3w48aSMCWHB78u4XB
d9EXcpwd8AduF6fBmrMlyFxgZpoUblYULkeTNKVb2KfHptgjKVcJllFLokht8EUduo2xihdNyLN1
pImRB+XItcs9aMPRzfR1kl+AaUL9mk5UjtnfyUCmpZ4pBkGFRziLdAOSnIRNCyaz3JZzxnJN5NGB
nLNpe4eHH+ztDgJV3R+Hld5QMalbRiLJYdvnKGuBhAXTUS1J/FaVcScg6GGsR7GkAjCHKPiL9oFu
I+dI+xMwAn25C7W2WE475+DND5HhwbAeEmeaxLvvwX0qvT9KD8AGOj1x/gv0eb7y1BWoTf+YM8VU
QNsU3ykO6YZzVrFSeY7hM7knjwPJUEfQrY9RWXdji12NWO3HeVSCLWqNWenbzAUatQ3Heu1qXRFB
3dur2HpKwaLqW9RrMPTNSAeq7Hfld7KwohCtl3c9Piee6aeGsktaNsoaIWNz83n24QUtU7tz+eBA
ofb9rIbd4Dq8Fj5z8wYn1LXYyB80WXF7iUJ82+7LQchFs+ubdJ4+HNNJZ7KunJFUfyP3OVl1z1Xi
mOHghsRJ6uE+9GVSU4dmdbAiaxkwQh68L6ilLsMHu8xVjg5Pbon9ihEHmEPjWWOAfxqCp0KyUR9y
2U3dsGQ5l2wnc2pk+Zl4JDYNqLe7GpL76r+gHQNJ16G8j1/iB+7kzaaoxx5jcD0ETX0aq7ki118o
LLO63b3r8Cf2sywTye8Fzo/jhZdOfDLPC4ThBQBuEdwkvAxG9FltGyiszHfPP0GZVSfLZHA0dooL
SwadwXKuu0F+bUJtQTUOheVG1/1cQmwHhStfst4OfmBEYnXL6XmLmuokPP2PS3JHnhf4NWfP1EPu
QOak4mpefk4nh75q5v2xxh6GOBpmK4MVQtCd4NmmOptW9b7oXAuKjHN3QgfHUBr/eUqzJH5+qXO2
ALfvjjbvNtNxpP7JThY3VYYtD12eogD8dmtw4sjafDUQG0C7aG9KkymUOjHF24SIDvzUnw0Kwt2f
YjQCkLze3EVJeoFiV1MW2kHYZrxbWX+8ch05QtN+S0hYLsWg0LeoFad54ikbJDIafGKCXqEgFoU8
t5sktJ2hogu1B2CfQpdOpbpqBbnhH2WI/fJcafYiGX32FOLHNO+xcfM8Zvlp3pPTKonjxPEwN9ax
njxMsJDiUTmF9/3XIJzmCzhu261TYM4i0iCzkTy9/539sA7vxjcYDHJkwivQxn6jKdbVSdH2Yuqu
R53LCYI+vJKqvxOXVm27EzUyMSP4kNibKzHmuTa8ZaquWyC7wCKsJ5XiN03+AwHp8jwVaKT/Y4DV
7sdyIHEYJUdgIgsmwZU3D7kNj16tMYyOGooMiFbM+oJlqIsEJAYmz9DvYA1WqHDPnmO+AQWxUyl6
wSfyNUJt7C/RZZVklHumRGMNi9Zye7ouza3NFAK8LGXG2s2Vcd+WHLsYw5WP3WF8U7gykUe4Lr47
r/zQl9Zh9WRsmpuIwn8X17wPohC/uYP7OhzziN0fPQnBREACpZ2bHkBKl4ZhjyKwtmZj+66vBzbM
GogKAyA3OMgFzTtYhHcTX3kxZ91cfwQoXHUWUNXpOE8m7Vt2sno2XCIXljAyoQrDLfkLXNAFDMq9
oB3sXPKT3SmTDN9u+Uw7ZB4U9RutV6TWOsSSpeOsq2QqMiBD806NRaZp5ivA1/M/J28NEINEc53u
34qV/9CKSXIQaQCM2I5UQB0ao+PrGKp2FIYVjJA8oHCaTbcKjqqsArkDWtsx9yTB2xwX+JQKX7Gy
ac5Tra5iJjC6RE3x/O/frmOmxk35eNW4yqhD/i7m4Xhas+lF7jCy/Y3JlQFzRJHbRdx0dpeNuOHP
LBkvrCQ6n20X6imsCjs60glogmiqe/T7pF9hOEt6oQB+iXCnDDsuxLFkOmSkj1RZn5nmFXXesuWw
KcjGbhHLvSmzQwodbMSsgV9QpJPY/w4Yxje3m/x9b5dtDaIanA1u1Xqm7KoYiW2D+gmqvPZJq+If
HDvpIguWTGUuWcs4fWDe8lMDg3NZYVYMdh452IvST8o4EiJ8Yj3PXXM8A7N1rEQMO1buYL3fMQOi
sb1H1Cg//GLFCqzpxE1Z8aPSvqs3Vub9mQ55/NSXXbxX5TXc9rQ/PPBxTrJOG1rVF3O8y1CnocGC
ja7I0BGBpPhanOyJSgx8Utiean2dMWp/FTFZrF+SZgqyRgmG6zPlO4dF7bSWstcm1RQoujsVIP6J
Q215GEd9mvh6UwV7Hs38/GKTUyo6Hj+MlDmrQqEdWyUiF6kYk11dlqK6/CvEiaj4+QVT6a1yZ0on
6hNJDY80leB+PYakc0DwKS7YJTbA0o3oMjYkJDfiJty5CQP20OCTxYqFOUwXEhatEO9mh9HeZ/32
Lkx/4m+y94CnbkqLEEAY7YMwGsvgaB9tHD/hoC5IrebJ0bEp6c6xlYhqmqrIPJ6dBlpVOgdf5Ckv
koVjIqieU6vQ5V+NNefbkwvXElfT7nfdhfXjkMbu8nZmFI0QIfEbrb0XpVdcz2BvB1db5X5Mxm9z
MejkTlF831kqrrwfFal7tX5CbGv+2VsAPRjE3SDq+aGZ7NreQ7YPf7aA6SvP25QtIN50OziJ/YDt
TPDN486N6Vfuqs6Tmk02jj7TMqu06xcRZRnef+BL2uOtS0jeGczBa7F1LCDNl51lvuCawL0GOv6i
YI+QyeBXAdETylz3buALyFN3fC4nEWUa2QanHemLhxj1NPU+kE5eqhnnDdH1aWPTlKMdEXFu/htP
Eg6DF1T9bE7f72ZCJYgQTJomFCwQzH+cIQw/ub8hqK2WDPUVr9c4v3yQI6PNfiogOLGpp6dHLDpY
O8066a8LvGxktXaHIqvki/LTc7l0ItVlCwNURidcmaD0v19QZIyC2X4Wb4aLtDmfOOuvdKki2pYf
ewsjpyTw1q+UVmx51anKAaf4+qwN0P+t6bEP0nfkV+gkAvtTspk7ZcKhIm1uqCIAMy/rDibgra4e
f8PDr4bJtePMuOlu0eDwsmFq3TCd/QvQ5dpapCZTChnHzRrlYSELZCdfnK6pn5LvBEqdb4L661QF
DHyGS3yMGwEB6By4B3aA6kiKCPS1+vYll/5kCfd3e89ix5FBRT3YHawP3C5Nnhyn1IQHEji0iAVR
xTwBuvz3P8mNob1lgixZcYv87Hl6WPLjKt2ryoHyXaXMdJQyfv20ts5gWyXW43v1dITOV8ytW8C5
Hoa5DqIPQcxv4x/2OBmK89AaAAUEfcb+Ymlzr51K1aMNQcqXjZ+LZOR29CxA10G9zB0d3RCzjoms
4YF9Kb2gMyFVWlC2jAumx5HLhrRweO6o+ArvoiZ0UKxPq5h7NI44sqFDljDJCam5a6O67k7WH8YI
M8JOM3lQLIW5bVQ9cTFgL3ktp8CwovY+OjGLjr6VNqHmN04iyBccm+xyCT4jbWO775NeqNiWL4GK
7BwhdODExHj2cNh15MV7EM1dhkdLEcGYAEP6GSlAr5mnu7i127aRLsGKnv9GPLcBC7u6Jgye1E03
VzIU7ALgeETJmk9caemKftLeBGuf6owIak5sAuY4NJz8kTkwOHF6saBxob8ihKLxr/Pmjupllxbo
iT+e4sWSHTKW0ufmPHyALz0PXftecFUC7AUq32UmzPKK5SfIkKk7P9Y2HMBMfaWNIs/T1GNBWMKZ
X73bNN2+JguKN30ND9GGd1dVAbSoRxiusVFhDrKf4+aePpmT+r0++C9bH2auZkPr30YBs/q2GfD/
zYsbRuA+Gi09+0fPi0kxA8/VuDWEgO7ICaUoKMD4BdmmMSa5h5eqknexbmy2/jLyo71r8HE7qiBw
kPZe8F6EOSAIFDE4+IOUW0z9eCTWj8nOZy80JT2LZxxXePwKA3c/mpc5ffVsGUXg+pYlwhqGBqNr
Y0hrgkI4V26sHDIvdasmc6EIKLBFKaHc7wXaacDCn1W+qjNylUvBUloMC3ClC9MPhfxzklvkcb81
IwXjdMMZxZoetQnKG2YO4xHxq5UWa3K3Kphhnp3GPT+u5Xv6twzWBg/YaSv2nTMp7uXaoGF/8ItZ
Mio1W/k8Du6ggn90k0bGqeoslXcbd7lqTJviWNWGeBpnNNAxZMjRB0ZnJxZK5LeVhjQdTLVVxNAz
d63XoUn/Tjx3OpiQers2EOE68CZ4ZgOdw35Qt+fmDzJTG6DNxPK9402Qt30aDERKVSYsqKInt9Fd
ZozvkRPNjv285bhPoSLpJM6pNWSz8kNDAFRl4P1f5O5bxPhlImMsoqIa43etHAeZU7Mka1zTTB3o
siDzxMHvCJ3s3egUceWzr9KbZ7GjhGydYx9OYpFcYtJ6BsZzFA62y2ihaJi79RoKkFCn2zjPUOhh
26aCvxUjJ2GJ22Npjpou82//b/uejvnsIAmsLxHHX3sf/V/K6ouJZcQXZIADFd6aK1ZHWWpgChcL
maxzx3mUmhywaMWbn8Yfp1nm8cvQQ/0sOVWqDC39IOp5tuY1zVnc89rkwejHtw1glYDd5Nw0NzsS
pA76Gqo3OowWC38H8Mo5f6805GlMLK1HU6H1fmsLrat9CaobcQ1FVyg5M18TxA2is/XTlWUQyAH0
W880ifMuSL+80V9+4q6g2aw8xPFGYe7LyT7XprFifkqL138dsqtwgrFfciZikRUwdal7Stp8R/g5
xdQte3CC0tSxD8PYzew8vIH5GTUR52POLcQSwH5TnUm8KHLs3kAMyua8zXY4knI1RhnR/ubCUmeX
BYSsXVaeDLWokBUVRVoKE4YRjV1JVTZ63Z3THjVMOefYEDz6qSHsyjjjq/20c2pg7Z1/X55r9zsq
myV5Evf6j/uO5R+AKwHOU92EHsbDzP2hguWcPsrmiqHcjXpPOaJV8Gvzq6YwfPJpnx/XB4qo+Upt
EYFmL4Ycnrs036FU+CuQyxXsiKEdGhz09HM3QmwP8JTeTozuVvlIwihvtFW5szdxaXn1kaZNMylE
VuN/K8wgLkQEmfSzuSPvPvB9/SR2gQE/WsfJCsFmRGgae+mTfdvrz3QJNFgDKGsUX9xPQys+Tbms
d1+gv7JQJf766VDAPyH5zmRkJIVmVP7kZfuNeil36bnQ8fsqycELH3NzYgjfu40qX2GZc/FyEJNt
z6FHqoJ6U5ZrH6TYEFkkI0setfl8IP4SnQW74+15hdEc37YRfMNitJMUllQFjlFVjtTtV1TQOUNw
MBBGbC9QOms8fktz03kWqu45kHKhtFMD4rWL/TDxx5TDQLyRT3MEaQShtXTeIrndpSbrtRIwlLqj
tedqQ8Sh9+2+TBcWHdYZ0xvl6MlqCv58cDQOJEuvDnpYqiSw+xlAjYBQsuEAPoiuIoO3GfyHvrtE
SZIpKqk+qOvIMFdRXfkDhnUphJapUaDZQb+0137mqLOXqJHxWS0XoNF80FzglZbzCSoV42sTd4Oz
PtfQb7PVogLwWf6P2sprNngTYE9899o2zbQRPyIIGVcQfBAAPufHMSBitA3RsC/QaQLS4ysue2oG
O7cG8pBHRBcuCjzasp6TjFdCYX3X3RG5ax8gAlYNVXNDbiOqnEE7VrzqwEgb2cSKFQa+BdUa01nX
2MWe25k3bwRoaTD2/leIW4zWfTcJQjnhipH9Wh4nuFZoG6S6nLn7rAWWxORzWL+R5sA0+ad6QobB
9yO9960CfdQRXFH39jH19TUy33T9OalIt0utDzfiMeC9hL6fjIcqVINukY3jLfO4h3Mf7kMl9ETg
jNyKFXwLERFBqs6jmqB6jM8ZEekZ2Nz9ty5Evi/nnc7XmK5jUNZS+y/EMdra/cNKVXiUAtEYRfqP
CTUsrgjt8oTCNDt5+ccuvAh7YP9OqHe3tDE/Xks1tuY/9sUTPRwZ+XZo3HwYXBvKIGOUoggTJRWf
baDutimmnEPNFsLCK6eXC6rjGhodICRcsdCIiPSa2P0izKfY4eTsBmPmgNLGvFOpJCgEaujYjEnS
JqtjTGhKJaq9XQypSSNWCqEBp8wWeqJgZ6y5ZlcuW7c3vx7Wdpv3itKazPeqtNPb4hDvoGxKVn1w
NK85BeeimQWfFMJVcTBTDddje/tGqS11JCvAse74xJY/GlWTvgoH75rFMrM6RnWlpBci3kzQY3rP
RD+g5BbrcpGuS2MAL6Fdm9/VjcN5I4liY8cPE0O4UacooH2dZGkkNONaUxcBF2DTh61D9oLaHDqR
CWhWxUN+Qvz4OLPJhpEu6nOjZHyB/DLEhiInBRRKsYI3mRepNc3vkmxmZtqRsNiHEsvlB2H5IJee
K5X9x+XDN4Skn5pSChOA08UGwC48jyQmYdlf3OPCCZvRQnnMDEWj0QTWf6wtrkWpPRccqKOnI5Ki
HF/1yKRiXKB7qAVJQbrzmjhWgNEYthR8ikk5m7i5VIKw7QEerIKp9WkCjU2XHxBjz+wL/w2L1+Y6
TYGtHx9hKr6kCB4DHROxMIEhkchvjZcwvyZnaFltkQciJsrvovjkBIk+BNH5I+AATRI9JVgraIKI
BnEsIY3Th4+ofFic/D0ONuvPKdcvA6iGQbllAXzUQxjTWXrxP7l05IyuUDw+Ilk/R3zv+m48aq5d
wsxtmxDLQyFW9d/YznlwtrkKiP6P5GEjVPadrpSG7s6/0YHF6hAEAz5cntXFXmzVvnC9MJEozueD
8O8Il/a1NXizLPi9Atn1dfqzlUG1Uer05zpPWd0vi4LzJm++GTV8FsvbsKOghLQ4930ZgHGCgLSn
aW/hgIHXfKp3CJZbn7nohtUOmEiqHnkvAy002ioTgtXWwOXRbFGH2GpIV8thTwImvEndCMfM99JW
dXAEyj/0OUAx7eXHpxAue0uvWnF68+fitcQseC6EV1Tgu0kD1WUf0eg2ZE7fB9M8VbN5CjsQ9yCb
Q5SM/u+dcCBo0TsSd3V6xsReOC61hQPYxhe269bXIdGz5ylpuub5NEx9dZ/5VQymdiF4YK+G9eYw
wSsr7Rde475hBi2Xq33MAuYzo7ndBx75O8XEQyvKDp/wjDIlHa1srr8YeyKIAUBg9reT1IPHo+Re
poSvWU1zRz18HOYp6SlO1bBOFYaRnUnFvEw2FrhJgJsfQAV5qA8ial1fwCR+053vvwlejcYA84tR
ZS93GN7HU5+5mAGMvBldez4kJJn3NDeyj20+mvfo6UfsUZDr3UkgjvqcBTYktYVndVtF2FMo+7mu
sHe+Kt7qd4zCbgiqhEjbMQ+BSYyp8QsHyGEOK/Zy7EC6E3IJ1Ilu5CX88Wo1jU/zEn6J1ubt9WWC
PJgqjYZhkfqbr6I+l3A69sxfkjWpmyBA30eI9q8Qu/0ELYkJuqxDL/pzultjatToaYKwgwFNZyW2
e/eUcpULthrI7VoNJBXPwb0Kw9fFuyHi98o5sMHRQofoXDc9I1siHV7wL6hWl0iCkS1qLflVFpg6
RTpRmJFiCm/s+uY6ueVgsDQq3ozwOKy1ALoAJKg/mrAnZfGE5XvZ4RzOxJb+4CkEVyEK3aNQuOhq
Pu0fmN+xglqGRYwQwBnEbdHXkrr2OaE1Icu+377hyE6CUJw2zvQzJ40oQEc4Y/yzL/cIP+q7F/mo
pPcrrdSuJ3EW7oskBbmcAMRuGYwsY/4j8YC2I4k99lI3eHuw6YFVXcM/wDchhQJrtRWfp3cdB1QQ
212VhVrupIW2FZHsyf6ABquu3YR1ehT9LGS/Z3T5QIsyPkbiaNdf49v9K2RSy3p74ZGCp4KfNslg
L+eRxinnFRDDMgK3h05LRRd+31R5mgwXVi+4nPUpAgFGuitCLTv35y/cuEAHDLv0SuQAGoZjunZr
BLrLB2zRtbNoCf4XKUH8S81WK54/AKbtQADEJyM3tpXaH2og9ztSfSb8oP1YnUGOWgFYnmTdcfq7
JxNCk3qH7OdeRG688A8vdbG1CFqvPC4XLcouVWkc+rrtp41kvUpKt7KpwSzJbp4TCdy0gyOMAkoF
URAC4Yzl+BnicUkVUx6vTbW0C+3il+dK7jXThlJKsqbykrAyO3ZbxDt9voIYABNvA5tUvZfxImE8
qEh44QT+4KiM6P1IlXTqhAL2QQxqelxtuDrmBVZKAGjhC8SxCI6RskVqpk2Qi7QxiiA9vyGgTMF9
odvgDHH1qBDttpzz/pt37TKXi/fWKyf0VQcB80MGzU/J4bSb9q/S5lQNbwjRfqDigClDcwih7jQz
hQkQ2r+NGf1bbikwx4g3CNri7vKdpGupE9v1uY1r6ScJaNyhXqX8I14jTTLBcKL05QACK62EJZ4t
QkTA2ydlWOSGbsEeKGSBZv+5A4oJqY956Gc9xPLGRiOyc1TOukWE1r+3KT2IAfKE38baJUII3qoq
Oweb6wepoIm8YzKmHj1DxriHpr4Gzi73l8EySONWsaPeD0J3nz4tlLoSoDu6wVfOlh2G1sBsLBej
oIfj0QZ3NrnA14Sj0HxfpBXjMB8eDWDiBcVJ5Rum54qgdjYMmfOzohSU6L2nzmc0hQVYP16MHwtg
seE+nPh8TC/UjHw/YP/FM4gZPBCHEvBnUx2csswxOgCtQtwqDWjWe/qlBRyCHyQlgMg2TBDfks63
5ndFd7hHkl4hVBEh7LPZpsWSwElJHuLxy2+Tl77pmDGLb814bWI6C36lL3Z+hkJSeNi/iYsmOPcz
ksfXMSWYmv9hmoks52EsLRT6zKd2oeF7rXYm14pLNrysttFfjR6ErvMC8VU+qa+7nCHWKCDv9GrP
1q+k8S/+VUWXM+oDqeW4/XI+Ru847XWaM8TqaHjjd0E2nh+oW/ON46XaYm5X3CwXNDqrMuDSYLkG
TfcCCYo69EmCBKoEDi6yRO57ss3t90eZI4GGqrAg9EV7zc5cjxZMx1L5q1/MrSdldRXPV3j3ZUnJ
L5gPQTz6zuh4RqZbZSGNp07esgCZb7bYvB7m20qFdQVQuJ+vtRNj1XMq9xpP9SU5kAPgGjMjescA
u5kEaDpYn/oYDXL4tTwb26STGylP49XTl7lC3yfS/6wU6ADBJi4UEBuOc4qeyBDaNPb+1XYVRtC9
daQ0HpBP3iEtgLj1E/a82IZLTIYWKpC4FxCvYtnip2umC7JxWrvgvPFrzWh7lGncvnKddwe/uUR5
JNuWHiAwXZnVeGJ2Xwab2RX5kNartp7MPOuRm/Y+cOYOlNEi/VO4b2gX5lH/zRg61Q4MhYTzZxTX
Knt25lZE0n+huE30Gv4U67yK51nQc8lIg+Dbmcd2emYhNxKoXJLt8BqMieOt4B6JRxOCHbo1Hhxu
PaCWO6yHbDlC+Q+h9yFvDih2nELekPOBfXg7MuwSQTNE1R9Bx1vgFG6f4GzFsONxsL+1BcvRjKQ1
pwvqqfQfAxS9Wiu/PY2HJ7ksp3BPqgk9crHSSGgGr9qnu44uRBJ99Ybt+TTQGmV1zvt6mSk1uocu
EWNknMPSHfZm8CNsoWviojp3FfItzbrGVCdIwO59PwG4ye5gbBlmO0QNQH4af5C+RGbxw/HP61Xj
4u20ZS57wnpPktKfJYr61SNTptEbT9fubiVLpbpXTE0UTp+AMsZ3WukvynINOxMB8MTCPvdhJlb6
8uI1ol+rSy40CpZKkxcO+vnwvy/dA1eDSeXAVilqecc3u1hH9OioUAUPz/4hChoLS47/b3RNELTv
G8JKH7GmQW4XyBDBkQtFSTUN4q+J2Pkt6xS5gPtIYhBs+pwEQp0krGAMAoPPKnnwkcyUQDLEtQQC
7i+ymFuB3SmqSiYwnKOMn0Om+d7n8oa18Z5G/k6flEhJW9HLUpkwj0ANR+J3T8XQ1c7Q+76LYA5E
yxcsstlZZtveLFTpYduvDuBw1gdvW/2uxlTIc6CKOrKAzxcDCQDvJ6Pu9Pd8sYb15Vg/KX392Mvy
Ct0yjAIl6srzHp93/HH4uD5g6Z4T8NYSSj/7trd40akTSwFIvQ/mJcFN9ejRastVopCOzdcmMQbn
I2MIH7iOe64YSJwUeG7tGcoa5YkO9PcGeGScoqP/aS7Gu25H0hgpuZO+CRzL8Ap51u6TbQkpU1+b
O/GwYcxDTJweSQV5y2CDO6EiRlUh3G64Dhe04VoqX9Dpw8ruVSrszqPXDz1cUw4mV2/kTew9iFox
IGEpUBhJs27pB36ap3ub0LTEJZV2v1OG9it+zmtbeCUc/wRhfeGxtDZkQBJiY0POhjRuzoRPPIw3
FXzI4HAdY4muNbV9HNBJjPDck4jDyhkxyoUxgKkfSFHu0ZR48OdKAgqNhTXKLSsjK+oXeAoIL9gP
6Whk7Ff4vlcTIYnzmXBjh2cipCpMwBjB3mhq0YRH4VLSpQvUa8y2Lhi0+kGNnYeAALHk+PK3yr9o
pyzAMoLyt9oq45xesrfKsNwPpH370jt94Zc03HMclTePwL4R5NOqiMHIhvjgER1P251JCzztM2Fw
Kb+SIsB/nN0Z+MvWEnGMw1Oj30/r9t2FVmL9Rmr9fAN9FpjXMVX83TDNyTCVvsGrMr+GFLYAfixC
TNG1txuDCcnQS905pYzNGE+lGMcIwC/9NJ40Pu5jvSx7QHaiGyiwln2PAqt5Gjgqjf+NLKerwIRH
EiMpWKgsY50JmT0PlA6nBB7zACs0IgXQzqfasHaXOc+pHIqcnkjkg6jRTqr0dt6g1U4p4SnYjQRo
2UJVTZ9itXSEw5BJ74iUOKvMrRs2kD0wr3j6eUw7Z2sM0A+xuXJeXxxf5aJ4O/8k89l3WFoetGK7
CcPvVZP0sfARVsm7EAQhM7JQjm1PDG/VtgakymFIV06Dwz53YEw9wNb68I3PVPfvwdudpfaEBXfR
GXaLGx5Re986TFk31RkXxYZ8VaHyCQ0+O6MECUm2Y4lcgLhdhgom3yP/hiH7JB7QQd7uIjZSBQtZ
OrdhCVqNpCbVcnVDjgq4JPf+GQTmcacjlNY4+FDA6T4zVA+2T4F0WrvxO7ygHY0K1a1GCRwB9Iap
WcKAJle+1es0ZMghkfshpopU6B7EHAsbPy/s/pVRd0z5xj/OnGQwGGpVJx9K317eBwdYjcGFT9It
AYN8y+NnA7dCIqB4LNFYj50SRLPtHqOHr+TFyRJyfhwYOp8YX3bJ9gAq1//djAwxD4nm+ilTsOZ7
JLqOuLtgtFKDM0XM4EFBuZlclceAOge+sVJytZGkXkZK8j1C8PNZMTtHoq7hjSHZ2roUEyxxQmdQ
Ni5lBjwi50K2/XnvomcrY4f5ifgaUtUswJ+XOdOugmFdowZUhXfAJFYUfgHwtiJrS4t3evjhoPCN
Q4BfVJMxjEDRi8Bdbo+Ppz3AUtoqY8mO6qGwvEPj0bcnX5/shH05lRv+2TMCRm6ShaWNNkzgOVeX
H2mn2bhXlcHsDYdwZhh7ldd/iBFV0FxK0sfggSDKo7nKOTQpyiqFp5xeZoAOw92S+97gIL/K1T71
FFbbVOrBQbIVzOPgy0h1xAHC0ee87A9DtxK1iSg6++kxgJz5lTyria1yA3ba/j9cROVZy6jrI/Lf
Rf+/3hqz/zEyI5M766SYCGfXUHzGPFUsO4Vwuv54B73cMAF18/dn3q4V2TSYJlmlMrS4RHMjL3NQ
H3yewsS0iiw7xAdY8h1v+i/rDXqWrq6OHVYDLkGL1bNfL7O030Trv/GtuT9CMhDkgyWtGXoWQBL3
pXD6Rt0jw6vx0dU5lJJizhL/8bqpWqV3ritLZ1XP1yGjtl8WY8P6GxTwvMMmt75CXRS+mtc8M6ms
G2w+R9wBZRmgTwmPaMv/HjHCNt7is0BUQKZgLB59P2h3KA/38Sm8evINq+f1yw79bnQJhNB97nZf
TYbiOitipL/MdhhNiu7mRuPewxNWrsbeva+ywzjMXezFZheLjSfircaK1n21wPf4JzQ8nbQUj8T/
Azf5iX2NTOusUAHrXWWWNL4Rw38gSjsN0iTN/pxanaty4DqJkQt25nmoZMp3kS0sE5DgJuBW7fzd
jTGPdMLFYd/XzStMYgCUr6aiUQmGl7ZaDEOKQoB+Dwn1vjfvQR1PDNeW80453Twi8Zy7i79KZMFp
nsLqwtAXH2z6a1VtwfoAOBNwEaKtKLVSgjgMIHhoDTdiRnOGtotIFN70OAATZ7m4sglWiLQtQ28t
Adbho6agzgfcdCra2B1P3xRZR5Am1waUCR1eJpvAAW5iTwt2pn5vPq7hvyKzL+SD9y+9KZM+tRdL
ebl79iyhp2TdAAjC9YjCLRMFTGhjfW1jUk0ZeQzBj/sAlHkGx2FFqfAZ+1OzgbVpjYkXAK+e5YT5
W6q3Wb8NR28x7oBdx6iQI3WIma3nCZJdiKPGObfDT2bRMP7NpuEsWYNGL22wzKL+RI59rr/4qGhf
aEeNyqDFyTJTaQFiklvPYrhei+HMorhc4aHLqgOpvcBX71DBEr9+Lj3lYqNxq0XrzR0a6R50zDYm
akgRvDzIwqhJQ7AZuffUXneTs4qGPZPOWKGVfjI3ZgxXA7hnzU3ji0W1a+PGPkoyj8mrQ2ot2mtd
qf6YmrMEAbsJCQK7XHDtw4Mch9j6gMVL2P6qCDoOGISNW6fitgc150pUr00wH421nK3hGO+dSh2A
zYMBtMhM+Zvf3Q7L12edPFnNtQ4HADk2kGwGDOIywPy56fzjow9LTGn9mIB22rc1wyT6qSf3nuDX
5eLCkjpE5wQ83MRyFtVWcAe9XkJUscKC/uMVCEvAe3QhDqnC3BMYSRhjNzpLWXshfr5oDEjL3/BU
EJmvbSI+BsZpAmylSpJ6C76bhQudggEOr+RQS03dd1oRcWaRoHYetClwuo/PrYE7iyxnX2QnYHvP
2o4FplTYiMpumT8dZkZ7KdCyutVFb0icwBZ2WPGwKAKVQdok67Zx7fQUP+4RRdW0cV0OmahrH2sw
+n+JSq3yqD54qoqtN6DiTeOADhvxQI814693CCoI09uV5UFQnPCmqYp6IqARyhowWpGX/8KTEwFV
jiMA2F3LN9mm2mgtKQzwmG/ANWWTmXpKGnBac5Ff4/ZZ6pa6mhZ6Q6fBZUwvuLta6WXNBxj6lX8A
vtq45loWQFIQoyg835SSpmnmjp1EoalsN/Nf+KNF8q9GQoIPLScbQJIRCfiu8Gwo29TzFxX86p+H
PJvHdLzvbJd9XbZhn/p6w8CCn64Har/Z1W7StSc3Yvin6pReSPaXZJFCNWBkgxqSFUuxRTDSZeRT
a1Lx/OsI0Avpo31EanwwVxCQy5ZYU3zi1QZvaOWAEPwNX15/cs2Vgs18tilHoxicvwp2rwh2JUY3
o9AQ0tBhfZjxyPv5lrU5jkh58RPWUDisgmbLQ/X4A3+4V0d3XQVl5H4nqiv9zU3NR0u3o8tMKNHV
jlHWRE4gDgM8ur2i8Lc4FYlNh6s9h16wvqSYtnbgp8ZuZweMZrMxH5fO2/8T+AldK/dovmtD7VGu
FlGatqfyo7iu7UZ3f+eczSOQJpFzr8snFOur4zaDF1DYa3taitaAdeBgTrVWgMCP0QlOU70AjfQ/
OFwI8JKx+QNS12xY+0+z7nGvSvqJrV3TLLOzehIDE462oTFzxU93tRyO8k2muE9BOM8r/fgfx9us
f1SfdLZafw9NmUfRYxzCPcljQQiGMFwHi9kt9tLOt4Yzp3KydJZHnvcSWA2G1Dr/XaVHcampbzcC
qVK39ZNzf6C/fYlW7+dLihpKOte7veWZF67Nl3kyRC+wM9smK9dh4kx6CujTHs2waBeZ2HBbh8eV
KQ3grxFcatOrEC64evAFm5+MEIISGC09doTeO78J+Cv11Q3kMu45/2DgIlimi5LkdPiPSOFeoNm+
fNaI0YPb9otP1SzD3f6QfdiPBjw891FcWlm45UgBzfnj+w6JqSTQi1R0eVHdt0KOj9cQ+euvSUfV
gZOPIS7fF0/WI8yUBj45vlbOS9lxPkfmFlSyDOacCd209+KxkoFNak7oC8qQz20PXYEL5BOC37Ko
1o72Or6TSHUKYHvL3knLyzjkB7tt2H8AHvtvMc7P5nR9HHQB9xFbtk4wthP2lSP8kq3lOAbcIvq7
jQHHECr/wS1R3eQGVJD7NSJAe0tjFVAbSxpATZjnd6vLSfcQNycTEdGrVRLJ3Gqah7dyDvaC9x12
W3JX+RL8NQ4DyumT7MH5lmDyZT1DwlYTqzGxuI+1pWMHyl6H7KhYZBrDt0nqS4WtY5TKZKz+lJmt
QMX5zp7CTj9tbGDcuB731wxrRMrRw3cuw1KQjzda72B3ymy/CinSmsoKNa+XUiMihpsMyzn+89Pt
rh+xEbeNXmd3sUIzZf25NIWos//e18+SWmi35+On+lBdC9w2A6bam1X69a2KYIwagfwZyl1MMHi8
fOBVwiUYRHHdiuOpT7NQs6sCadRAFLth/+X7Grt+brjO1FBBpwQu4/fj5pyK5ywGq4tliaRSnLQ3
wwT+hGeuzt884WylZ5MLhXVv9TFpsuAp+Dvg6czIK0tj0yojtPAQhI7K5bZTzAPGRHOTKF2InzFB
iVi3zJBAE0+alSqwlbxUEQB2suVEfwtFoul7XXXk2LYYOUeo3DW0lpA3axWxZGYr5wwg3oBj/Q95
GUCIpm5jj3ph1EoJcimZMTzzp9EA5/6zH95VsWJO3PhQ+vYdNN2Xg2EpiP2re3TVMVj1Yglz9umP
zrhfLX3IshZVI7pgUE8E97ZyVZZxM7C97u4RiJYkGhoTmS4iBz2FKQPwhLuh4zPKarAyZwcnKsqi
svrs6Gjy1vYyihhHx3eLaBH91RQ98v5bl6ict91Z68/y1RoAjoZP953/UD6BBy4KsiIYuF/bccay
pimu5jY8fKKbhiaVlKGUu7Xzrm66FyftYejRoCdqRDcFUJ0cnR7y2rWsGCNWiKvxZAKaroo0US+R
K4YEAgrUBm2zEtHzgBzIXtGZE5wbWlF7Ulk3wR45r50K+/L3uGgxPXZLveVSOkgDZYvDXMMr4/b+
EuG6MDSf0S6V02obS95PCoKeZi+gup/w1lXTg6DOCUizg/vjr4vw4loSqXIzah29uITKJyzVkllB
Y8FwwSUavyuIOwe+6Awx2E5flnJ5rooi9LqTr+syt8ia79io8KOSrt7nvcf9ngcnydfdWOb7ZDkX
1mHrtZHM43O/qmQ2NcQIwiO/YOt8YDe+UWZe//eGUvOEuryJd2fRjsT/deP8l3LGm311yuQOXNMt
GwjW/tvwdXVh5PiV3A05nQZjdabXlX6wX8HE2+cTW68yyom3828nZcDtkbjgI7iEXxFbTcCm9OFW
maoXmmn4FxgVLLcdw+uRlLr5bC+EevQtHlzbvJ1i9vfGLMJVX/wjd2+oqH7N8apZc6p2XH+nUGnU
dW7AKrMq+LOEuu0gF5wi1hhEKpAFG9gtInJF78r7tG/7ML5JXTh8IdOZdILpgYHUqWLPMeK4km92
sB6I0vVjkE0GIO4vA1/BgGl+6atcdrbDPV5BYhPI9tIzGQ8qScyLuoH5VhgXOzCHprcWVvmkNxWD
6XdklPXCDo5pCAdlcz7rexIeJkV0FwrILSahIHmPAtkaALyUoNaCmtnUlzDQSS2MfdfHIUEBG3ou
tdl9DcIpcSiDTUiYw7S7qFDkwdnrkAvc7h9NviksaTiZA/B0bqyMn4EitxpqJbM4yGnP+oTyjCdl
3an/WxD13q8YWm+SCwDZfrEGzNrD05XuzjQ1maj5w5Ud4M3JP1fHnZcqJaUSOcyZvlzdra+oCdDI
XguqpWXXtSbN4OeKdG/jGfU3KBodOnnyKHXrGibVY2gNTAz6eOwoyXOc9xCj/qWjPN7l2qN/igIi
OKCgB2dOTlolv7z9esup3ZTfaRn6k6WZuE7z/GCeagfH2IYCEZj8KYW6VUP0wF7GRoevtRuwUMUP
sFQSDh+6bfvhAHFISj2ice91m9KPYJ/LmDqf3IbsiQGEe4wAsiQ0+Uv6Jkc1s5wgExtttivTSnn+
qqXt2DdECgNX6Bzpkn8tl/A53jNa3kHDxD80v9p3OJbZHmU149h7g0BIWFE1+AHVW2KjrhHPfmRs
BjlJ07WONBvSDU8x1BU2qCuY/DAJr/ISLL71ZGU7VpPDCj9Hyst9LaQax4vBSO2SMTacMQnTQXp6
EnZW4P4famuSBELM779YvqUjhKhH39+gsisFWIkNznDshv8jeOa1z50Hqh9mKUL5vr6YgffuqDdb
dtdDUHOGHwV49RkTSgK65aRJuXE3uX85f1FjEWXm13b3MF9nFsVrMWVUbBtqI/zQpCjrdERt13b1
NmuQOuBTMHE4uff3aqur7yGe4tMLMDv8nrvxNAIMrjPRIuctf0ZDR33g8TpCQpzJ5j9BXxJ6aKCt
IASOnFQ4Ab/m8l/vFsG5KsoTHsx7E0LEU8dmU2M1WXt0hDxqofyyL2Menex/Owa+eaotdcDkZAxO
Vvwe1PddsSPXK1GXUgN1idoIKd7iFM+BmyIA9NI7bgdNkM6xZfhdLYd3nN1kvgblNxr1XO9FRA4L
py3Bb/JEWF3yHc4HMnXPqa+OZbLUuXTFBNgLeNbA3C3a4dpCva5+X4XpujkUX/owVH1UaS56dQGe
dESUAXo2iqznZKTebQgbRSUACA3XJztlR8EvtgWQ69e2Ln1dqDcCxSRipB3rm9gPhVwxWvrOBCn0
A1Ons/kI1oY2QpzdArX08JEhQ73B/vEHRGVuIMvTbK0nRge+l4GtASUvZKjnoMlzJ2gZcm/Bdqc5
VGjz+V0MNwkdr0+YiTr3tnHv6dfFM/rbFfa0eeapRwJrPOoK62HTMaHcoPy9/NQlykOjYVGocQTV
eC3HaX86+m+DBahF6X9dvhj6cqH36aaRT2COyDaUa5oDg3FIb5IlrjWeeVdnKaiE79FOCdchMBGV
sIxOSvRo9LyHm4sM60k7Qzcc8t4yeUTY/4mqne0RyNhBPg/M2a0suALolmPDIdj/22R6wIDmI7Rw
mxsb/Ee4+86LWWe9thktWjpMLUG05AzwflZajNhB6kR+UwigSeTugDZ+3RyoehChVi+TmsRWXeOy
BPFo48Rn3AUBJf+fqEJmuGFVDzlIxU7FlNSxjkg2Hpumm+4H0eYeqiarCAg/FSlpdjOTUFse9Viq
rvaQfFF58gRRLncQbqnBJobx5XPDpdgh2VuzcpkkdbeN9WHxWjIHB9o4imhFiGPnVhDCD45p9TdA
ZlVRlsCr3IH6otMc9L2eqfg9yW/6aJhrnDInPADKd/CGeTTL7o7T2prx/VTj+0znbtizYnTQflgo
QZs9mg0Q0DNP6gmGnMJEhp3nr8FoQW1xuYsTAF5PiSUFaMineBcNw5o2ZqH2Tfc1GuPOBabjOiM5
6CAmNPksqefzlBd5y+7DmAb1ZSbN4FOi+NDJL8SClD7AzWWU6EQUeCcx93CLSgsWT0DwBTsmKlkh
hemjOrmXVsUo99D1mBnriKcWX4hTVv1b7uGZul9Xv9AUOJsnKYgAE4R6stMjHCqJgXoXE7ByKm74
+QLiAnfcPqP9c/bl9NU5KyS5jS2DKhhREqfHD1C0uJ0eY7huG9ip/QqfTTFhfvWRr3LOdHKEB6KZ
8gFn2PpuMekHvlTIx0ON01q/xhkSiPA5T2WfwrOrGToGFPqVHfe4Lu17g89nzbK0Poq1CmgDVCIp
BWw4O1e116piIRN8tM9D5uCeYAcHpDDwiHCabLf8KZoUbwvl8KZalpph1Quj7FRR2zAZMMoPjlv8
/enRHGOE3Swc7hetJR5580z/FleDBlk67EbUqJqut0dir4mhTyRrTFqnU3djE9SJu37d7vfN32wO
bXxy/4cewhArQkTRbqzUAYhq0Ym6VCMK+iBGUP16yGf+ILJlmG7mCs5kW3xzSSuvvNx8zeEVv9aJ
+5qH3hZECIlomOB9nPGD8n7TCMcXhsipeYkBZeu3zWX2nd5+bTmF7c42/PD6ySEjPFe0pJGcjzxj
742Uohp0ZSf5oWPVvcnud6qePMGHnJJmFwbzp1iK1RJZSavEC5MSEBcqYX/6IMW8dOzC7JZzegfN
m0Qv7ItDGctPJRaGOhujDQ74EQTyCPLD6FXvkWrmRCS882gbAAHXa6oGpTce2H+r1mUfKHoj9HeW
nMssduEOpqVDiprJWsF4J3yC2LRbU2vfpKKWI++DQlOUbWVgc1tHcAWJ2SFn/7QvervjCKuv+WKh
QytVAwBX3SpoyxAbJD1CHV3/dfSak+RMdCEMB1IwpfLR/DnqRBh69YVnebKwb6zbBsp08H8qhohv
CUTVXI9ZAtD7MHn+QhIPqm2k5vHT4UsEvYiV/1TBidEWMyirajKirrET1bolpSc0/ALcVX4HredD
uxEcNJ6da93QsqhwAgmCnwBSWc0mQmw5smsCR2m1xC6tj7OCQBsBsFtrLrEAb8EBfvxHpG0MojDd
zebbG0zj9v9lDzq9inU3YM8yAW9xkQdA1MjyDiqQNpZtNcYkn2KLTBaa75BlW2sE9R4WHZn59y7c
zJSwDWj2LPNKsH7EqEGr8Gjoy9yMbwnvlJG1+maKw+BrDIxBfMoq9y1+nx/Q5veBw7vd+G6YnaI4
0kXp0F05IbP4oq+Bth3Hu240y1d7jKUloa4OjFfaKY8pj7oi5Vjh/EbLxuamlTzn5BHhF/xE169x
9JqeJC8bf+5xetttZQExw8mUPIzhY1XoBfyhVFfrcaZkmqt9+wYj7lIPd6vf1ZLBkZa4nwHC8deD
0JjrJfenEeUAZfb3NGr1TsBoyAHeopWictvGLEWYszAW2p4vlgz6jxZB2bBsc11c3HplaqePJAcH
cKriFr71hxXi7ci8jpr2Ug5K5uBN9vfsaTtkdFVAg+2nKMTrLDETLq7+T5+Oblc3IRV1SE7GKdMW
SV9YgvWucB7s1MnJzeP2uGyRzbQw7qRj7oWXushvb2zGnvf5QjqV7ZAXwnJ/YrJplh3FNtbAM9PA
eIU6/Rg5+m2b8VMQZWgCKiHvqb8ZzD17FE4wYAqLLdTHmQr6YSGJxa8nc3V29uk8MdKbW5UnNQnu
7SNTcOxG8F338pThf7HRqcTmmPD7uoYdadBbGLTXj5KAA8f0PjG099caB+RNvILR4t5u5TLRqW24
sErCLXPxHAluudtZSOVHcldiuJm75UTEtXSzpCp8yO3w5fQPCg/0NqBxu09jLfEAsmPUC4ZEQsFp
9TOMgahfDSOHBVmJ2GnOkWqHQSnvewNa0v3NXWEU139NYUmCG48MBFql70pBELN660Rj5w0cxIa1
shPuLV/iAsQDPQmTd0uAmDb0dg9o0HgCynMv+9/5FSyZUsy+rQ4UafuqcYd/xxlWaenpY0B1R8VQ
gLYadl9+Z52I5xi5GZrB+1r7uJoGv1cdsEE/iyQC4zf7GDTXt17NFkcOxvsYPwqNuvjt0gTMC133
ZGRdGFEq21rzUlI3d6zXRgQWTd+pUMeQhNqzQG/meu/l3omU4ZPTYu3Aldg7LC9fgcJSFpOBG6JL
Elcfz+hnEeqRHNFTQPbyvm1l4u53Cv9Oau/eUgTDnD8eg2aoCKiH7c7MqizzlEdi9uPbB6LQi8Ql
43UBlW89G2cvHVRVw9baxdHNlHyOW36HhZ7hwN23TYHOQ48ANCNlg1Ld+khfhILpggT67hsStM7t
sfskMYUnZCuEdjDq2gBtOMDIFP86YAcLYwyQl6IxNtMok3GBOCKqNoFoP0bQuiAhvUEsQq95EMoA
+S9ioQl7fVvq67gpbHOsfL5hXH5SHjqZqfdq7aNhF6lsOHMSoYEAWypbnR26Y5jFfGZlOIzrCuAm
967rXtb1RcBHwK6pCT+qEQT0pG/OZlHfND+pCE3KuWnbQvk9KtxqL6JASsgtK2Zb73R80iim0t+3
mBbVGiXnjbpS9LMWXCTu3xF5aZWHQLlt4j8/lPuMIAkdopYEFftQoQLlKBN8AL0TJNNhobhJnse3
bICuRX9Zoe+rXcmIRFrp39UXNKojdoRFfA1yN3YgPYBShYJgW6w4MA3ieWHE21GZjzHagL/8TygU
w2rc+oDU/Zx8K8oTNcsgpKctinDDXUit49Mp4N5lgNqbaMOkv0DVrMyin6eIUnK0/qGviwpDnksN
J+1k7zdyzLMlAp0NWxEPV6Q/zIDPlI8UGl2JH2jqfbFgoPM8SXgP8+1oOeBnCb4xJKMXr8TkmOBr
xEP5qR1E+XIC/Nxs467/VHicjKSu6p64pn02tilQ1tRgWPBibdYnpyHHZcQ77hz2EGGzSsn0Q9Y7
6s9mZxlfTnRC8Qui7+HY0/Fqz+CY0iTmOij4qMgW2Rqidh6HkUTOTg/D9ssYUUJQgdtfkudHZDX+
kQZwNEq4zFHJNWvap00tIVHNSaaBY3tOVy5/KBpErQlPwv80jn56dkiL7RnX/g3tPvpztRt2n7Ay
8PZO+RpTjelSh1lWH080y9OF5SMTVp4gw5zvp8dNMj2zWr4rClYT/q6r4Nqcnq/8IDraccMoqejK
LtYYmzZP/KStdZGbVGAgVC2jNOHgfXZHTWaAaMC+uZQ4Tbd3juySRK7gkEGMn4zRl3gEuPteDL2P
aQn9lVZol4YoJObQsV/hki8uGdcJqKxaL580gitge0VSaBGuwA2/EpOS8TrmULFbi7FZYkFK9PWX
5DUH2i2ngh6QY+t9Y2YkCYmVshEQ0tenP0hDiEX9Zq/nsGVFotyCnvbDhhYRCdK95Kq3kSUaeyyD
MLDGK5tnZEgtPuhY7JaMfSG8PQnAusK2LfuIis8tifPRARwT+AN6aJbxVt5PeWphOuzo2ovw+1io
wx+Udqn1Dtv9HVHm80I5qqoOmOSDpOuezxZLkkEuZ5DPZFJsi9h6oZe4llQ9GYR0vMRK74rY1mFB
2MV+1C8mA0oxzzkPSuVamo5P5o7pV0bq/55YbUy7SDeoQqmvvbpMc4NvykODUQ8ETlgY5bA2Vwuz
Be9O0kqq2Wmr2+cQHMnG6zmzEoD9IW2rSMoR1UDgz3O99BSdShgwTPVbi/EJw0i8G3wRprY4q2ZW
+0YgIFbuqlN3PZUjpR0XaCcAyB9OaPCe7zGtKRTGPHrqSLGqxFtAzF0XDCorVMCf1j53+RAJubh4
J9gtY9tgMfqqeVBvxmhqaA8c2PcLcrMhFF8du7FA2vWUGb3rEBjqMfzeHE6+l0ATu09fhnxgqQKi
Rtf+F3awjkX3NKiBUchyLmgBSvKIDeIUGcdzQb3qua3ux1DxzxgOlWW+lF7qsxLzz7OEoa1oBF1S
mkpBr7gXub/YRk/VgyQTmHwxlZ1C302snkk83/xoWwBRbgnk8HL1yeH5RAIjof233Rb8YBUxXY7D
Pc1tc7g8zYCk2T8fxmPFyMunlSS1bu1E2KPPYuJB6IPaHAZG7uVnAhdTvVGuLenxaRdpicstCnkk
Q1JK/v9PlfOADvmGQt16VvqLqLpP/NaKwguU6kksmQDByT8EI6dPrpRzIpcbSO+W/HrNPWOPFit8
I4LwZKdLrfLTr0bozv4AZ27nqkm1JctM9TKdLGlbGDcfL5hc0h6zpDG0fZKcSJ5YuZwqZE0UZrzP
R43nnswMov40CRjqFDfAZdX0xvsPg03r13Pj126IDdmIuTD4KJ1c5XR9qlmg7a2T7Zl1eMfnnunc
FmPVM+JN9GApgH9E2Zr6am34tAMoAfp69s7urw+eDTvZkHpoE5ul163HdfUChjFvcjpiMZzmu4LH
9ZArRYAe5KLJgDhFJCKy+O+6jzX/RqHtSlENkO5w+0vNjJerxxQo5zYsiyQ0p/QJ0UXqKrAnAhuP
4rpHvDxp2mqHSdfqgLjknH0UnT1av7NsxLhulUIcpFmgcPd+QtMcxuLGdSm3Tfz3nXk7MtiemDwk
DKQ1qoDvd8gy8E7EHZuDOdldr7tFwM5ArkMHl8D5lLKO7mCCrE4P8mWo+gj/2JNzZD6tqB2I07nY
5wSgjm6WF9/e754cTeY9M6xVaq1GKXJyFlz95MWwbu/6l4/XXlb1y/1uvonJgSHdQ/v4U/OXx20y
f6IlovB85bKHaY27AK/Lv/JmpZsky9aFvRfWA3qHWgHfPhmfwyd/uWMZLEdpuTM5mrxcmNuWdOBj
0wP0ogi1REYfA/xUWf6e2i9rFwiOoPYPN87JkhEv/rgeREhJmBbLp7vtk74pfJw6d9nZctpnvCtY
E9vYgCprSH+B+tYtn04KEfyeBeh/roIxouVZfXRD+RYJw2H2GdVq2HEwfwOtBLodo240cUkR/MxY
bjYGyysAdmW4U0zyNJ/KYCaHhoAbr9XDbtrfIT6SNFipXlqrEUYRJvPJdewEkC/u+3G6Pmatf/P7
tmlBbQBsk0g52Tt1Aw27iLZtcNoD3DN7qY7OpwkvbqIcCJSHP5caTbBH2t0zjbCGsPgYNJqTzXuW
yVJaXM/M1MqG7Sh1FTo/t37QiBt6fQTUQoHbtTNR2akAzS6DZYDUJnLfbFdqoix7ReyCn3HCLFsb
5561Fv49DMzxh0RaMFJ8B9ouSu/IaaB1E1ZO45YmbxKvaRqhiOqaTIndQujUYpi5OVtuQrCxW/Bm
hu4+iO8RCCB/Z5tp/aSZygvNKhKetJrHHUtFIvyzzmXkvNrhNwL9xykoxhzeSjwgsBqj04ewXfu/
ss6b2g+ql0EY0u0lpZi2qwPxlq4Ibf2p0ADjozTrX1JqfJ0g0I7yX29KBnDRhjND+9r36Ny2hIyB
Q4ZqZGY2pon1jk+/K6rlH0YjTRrJHv8lykMEVnNnXfnidTIdisArWu73wE/aCmae6oHGOTsDdMND
Q2FJdzBS2wNnX0+jdcr5xyRqRzJVM4R6fNIwD3phB5u1Os9a3pmo+O+pV1c6FIEqn37rhcLPvbWV
Uq2ymV0lxbB7F/Jz7J8CFwTB0UxXeGcowEkiN+lhQwrXHoWd06sFVxjq8yEOCmPvwfAvPm0dMbue
8TpSnY4msQM2gM7HhJg9DgEdDS3Kme2my9Y3El+1rm/DrpkBpf0Jvvh/Y91+Q92BlkWDC4iNv/Xn
I9Myel/uKzH4hSV2DO/ko03D94gkzEVc8GFV1ujQ8e0vjIDgHV+cgFyl3f0YfDMLy5xbpVafASdF
IbTlqlIa9knJtFPlWKt2+kI6quztI6eRebOXoe/8IfwpXHettKeh2II30x84CAscnVkM8X4G+0Lg
QvBb3c6TOPMQrErelUheoDv2gAg4DFPI2Jb3PpX/NYDhDIBPnRzojJh+7r6l9mVkHPwIp/dRNPVn
v5GnPuQlhtuhrzd56nbg0F2lpI1NNerUkE4PBRxggGH/YllQnJ6S6bvXgKZQ3898wh9xNQW5DG2y
qCWi0TCECxZJyVp2BHb8azy/Ea2aKdwSvDHm02CrejEpS8hNra9ARi1/dNBX9oMo2nbbL9V7xEmX
vBQwgG6PFFLAPgjbO2iGJjmfIN/kzgmKSgUffcNZOWiKZVlAtjPkDAfqsQEucWw2nMfUurjHkxdG
Y/uvgvyTVudFmmzGRnNOM9sQjDjNmohbyscBwypV957opg9shY38q/gHXPmQDkj0TkHNQF6S+GJQ
HL2D2QsPiRkmg9CyjeOGadC1ASOv62nyM+Sc7FdtoXA9a+qo2MvegpbPTwKfLaOXJ2MQcF5GdO/j
FuXtqfxqnf/+P87CsQYaed9orFjcGsy/e+lf8v0V9CtTqm1ljPW1ky6K85NWUEiULPxMPzYPqA5x
qYRaSDkEIy1FN2ik8Xj2jOMAYoICea8nmv4NNNtffqTUReLRLI9sMhVmvgpkiKMCzvTDWKnHB+ve
Or9uCHHYERkhoASevhCqM9q5CWzgfYna/+1x49u3XKpuXJUS9NBzo6jJDpm7nEdoZQvsz2TGhJ+w
yzY6S+y95lSlNPakgj7S/lK4Ly2TV32f37ZTURX+4klAB0HQwKjjY2JP06HrgfYhtHIrVQay/fmz
CgT4ERSMCS5HrQNG6aOJwjuIPDMKFO8XM+W7xaXGYda7TunPLbPlO8KZgkH6/O4Mf7vbgHEcRaUf
LrQzz7hTlAap/NTeYLHXDlJ236WYeGZpz4ynkZOHfjSe/wAAFtimxoSmHgOQq6HNwoiyU6/ka2Xs
v2xVcFS2e9bAtNdUT1o78MM3x/ApV/TUVHc/IUevmRskIITEzI/kUYP/1WnN1mNYM3STUBwfMOEV
RWF5wvbE8ucmBMWkzYu+XZ74Rlxa7ZEmObLm7Qq/bzwTZLAXxZBVbyx+0VebntUC5giRzvZBFRZJ
WbDxl/KnXHx38M5tolcP/mIA28cl+hwh8mOPS/SArBplnOuaBsEUZdXGsmhuULfvWdnp9xYqYVA3
74lNvFmNhlLYzlNzfK3hMEC+FQ0VVvqDuuIsfFH4z20X815ATSCVYDr2R5mvsiOgMM9fWrHQUs/d
UXdF7kgy1fHUlfCdiuRpwMoEtmTkJnfbA9cd2SDgcExc/s022LbSTihgmu8ZvWbePLupMdRsWvsE
nxRww/+cI5PSuSJZXGtF3dznD6rNPJJY81JyZKR08o+UePeg9mk37S2HpXS5e13D31DpMxWAyLgr
FaXHNDWGwG7GgwZpVqXuHCWPzMwqQZXCRpnvJEtU6cInOKcKN3GbmP2C0KDqlQJFwic8cpOr9W7X
DAa8c6s4AG0BKSRLNlKZOTTML9f6pk4AkTbRJ34m4PQ2eRsEtOTrA6x2+S9TikB1ojQsqRfJr25l
A4oKvvsB9x9nKyxchS7kw7MsNMr2Tsx3icqyZHXigqPTkK4G85En7kFnaG/iJTmpDBuHLf+bVG/5
PZoyoIeeuL2wqEBNzjiPIh6irmJCKa58g/D2qdLPjw3dGBqT+Q7TXkpSlKbXCW0dhF6fj4EESsh3
sn+7Gy4Uspuk/RtNtmVNHUTd5bQeHoVtFEEcWmxWYD1GeQ3uV/4MDfHhTdfzM/NRI/mgaOsTzwYa
OG/x9nQIckSsUah5zGW58jqIjtJX9QGWACJZwWaqCiTWzSssMULUeBQPTDNja2WhG527neqFZK75
XHRfQa+Dk1wC/mdG6JdmKWCJAy0QzXbou6CiuAtMHtFv4yByFWSbCiXB2eLSPnB70H/cYi7xoCcR
RBqqykwe9hyK/0ua13gulALs7WGOtQ6R7LVEJ3Hkp87q3ZuXlMAScWkKBctHps5JgPg6r64H0V04
LpsI7ypwn9YdOXvO35cK2mWNnbRzLbLmJ0+uJesG7AyYP5InmA0D9VFiB9hevYKcmuVSVj23TUSL
14FgRlyb0LSe2T54AyXPIG63MTDUOu0WqIpOWEEfHr/KMuk8KHsHv79UjrM9QewlP2fE0f4OCAws
rlNfIRrCp3yV3QohjGiS/KtYp2R4SN4DrB0TxoUb6WwwtdfW8YNhiZR1CufcEJ3hvztx+7mGw2eO
K1fQ6KteVRbwuWXOakeaFfVTu/7GVdt6H/AMT/gd3KH264iFc/levQvYZcdV2tYgex5p4F0wYf9a
MsJMd2Y/QYhhwPm79xE3aM2fRq/BNP967DrFNnWtYTVLiBYO9r1KA5tObRJ43N+08VUvX7jejRVl
3aMoIfb1+4E4akDe+iN5okopWxO37Cwn5OD7mhnsIkD1/0F5VvhSzgo8t03fucymNN0QDInd5Pc4
MLzwjVr/pewVVgKXGZGouJx037pmfyAkP9m5sWcEtsHFnmni2IOKh7/YZBYN6ZTdtEY3fLqvg8FJ
NZR1vHHfZXCN1mZGSuMnksSZX/8cY6ve55DlLXQ+CRxi3EHxP5iyQZzf3m75fWY/GczdXdoncdBG
/OmSRbC2++q7Z1oUqp3d2KJEf5kAj6W5mkGpFkOC09UVMZnU1r4jDpuzS2KhLMMT5oeGSzPdtPl6
Aw4tvV5xa303KyVzIVJ0cdA3rmGTtlHvdNKE3wkQqgAxi1XshkDusVnEG/i90bkEWJyOKC0QnOSy
vfWBp1hwP6mSqXcSIIoUnXztic+h7D43x2gNa57+sA/5AKo3J5XBs1qWbu4H6t9frdeTeZCScEyw
zzVvvQ+0+Adyb/2h5D4uGOtN6TlJp/BA7hhjcuhnv5VG2hR/veyPnO78tRWOHweZ/0ZwNiLVenTd
LQdEdsS9e7ejwHz+pbSMceiFW2ZhgLa6lWcCguTC6pSqXKZc7k8txqV7c9lYekNy8k0nANQwZcts
e85zDpYNQTdMGwYZ+xDT4VVnux1PnAYMu4vQ1nUG4Cf3yvNJopMrMYWqU6BoRFB2N/RSYIe0dNbC
GUNRIrwk7Vy3Bs4oDiUx483eau0FCi1mtkjT/JAubvCBUmPiX4MLyjPWnMXLI/LNWQProFYL4ynq
2YnwTU0GtkVdx5XNjo7wzo8+/1Q7SPqOjLiJlTrP/01y+u0J4kOlIEzrts+fZQ9IYhM2GtY1kizx
3eU1a3bcLwHSkMntfNvpTGIovAi80JyJCERx17I4TIQfcLElghKusbtY/VEJ5s2E2R7umc+cSz7v
vUSnoFhz+A11mrBV7v9FwldeMbOdi9v794fUUZFkEeqtfE/vTwCV+l7cRTyVlud11kDcmMLyyQbY
CwzPH1g+Bf+QwFO6/ATN7MM1gR10uHySaoB0153u2nqpRC97RsWzapOM9idzBCWy9Ji6FpdlgkHl
kvNy3V7nhVksdc+FzM/iRFaAw5eJchyfcAkrEPYGsB7wxSaXfhOdCx0ou9dn/z0nSmrUxgteB7uf
XfAIwCDALahZjGHvgKl1K33Hn/YwAglHZUDuG9pI55onDYcNKGN7BgblJ/MGdeVBlVu9xHHv4LO1
2+4T7+DNdRw0D4j6wEyWeolDyfZewkPjFgMAlQ4JF3Ul7Baw2QGcPl8UoR7nvxrLJgQFt3tU/0VE
MRhizrC6PRXBhbko3X6+R5j/5kG5A13UKQzt3bL0JrCyjMdzDVIYR8YcAdJRGJ+3/It6Dj/vP5m/
HjWEGhKoRdZWm+ZjaiUun1vF8Tdn+8Am/7e8D1fGpNH53NjoNk74M6wTmJ4O5f3Es5erT4cYlB0i
CYvzO3RWH88RACCndh4ms5Q5N4ZrllPsR70Gjh3h3vq4tJm5mf1DOjfOTDtqC5+jh7EfffBDjUAD
8XrPV1qLlODQGHHTxzuCILu5Dar9P/y5UqKkrBuU4uqsP9iuXeAdtK9HnKVhRmRu5Uhx9ts3ciFp
SFpfFomiYf5Wka3QY8nKUPopN80ooTOXCpyw60TvnheBiBpo/JL7SBK2Mg4Hu3KeWrMl4UTLu6UO
a7xwTgIR48r3Vv7Vzjad75NErPBWg//p2ckbHG7/3Vs0uClN/jcfvHjBqpmRPjV21Imt7TtumW+z
AN9vh7L48K1Iajdyr4DNFjf3N6HPujrHwL9NobPWm/MUKmSXdvGqweM4lDT+3BzHmD1+dIFH/7Ro
iiHEAsFJ88Olbnv8suBq2DI4/kjMCQiz81Cjk5KbpNU+7CJ3fI/HKBeZPQ1jQELaQuj3ihlKYA4n
6HO0RLmcj2TFDYzGf+HQ6nTTNL564VbC7GV+dvP7g+eevrstW+YdK6TCqQo/f8FHBcA6s0ANmzsy
KAOQN4sKFleHFoGjNm20FIqo9EcGiIcTBed2eCRVms3428pAHUdEocoMdreGDIPAFQaZOvkhFumb
5K8PqgFXAtEvZZvdcm9RU+6dGGzvDT4vjjDDD/p6csHkuWKlEoivMhX17c9S1e17CDWJQLQmiEo/
I4IWqZqebshE6L9S1G5s7qsGGBXPlm/PYdm8SECW5hlHpUPP6uUq8rQH2ILfbbQbfcWfwmoJsSlI
IOZeav1nMXAxt+T8xcdY2Gj1q0wkdDOt1HWpnLWM2xahmDx3JvQenZ6QepYJ901e2yB3nFpawNsy
wC588875PNSNtOWSZijLhEhLwqdDOOYwy8Qiv1+t7Q2tbYBUzStW/wN0zniVTPbD1J+UlUGSlS5K
72tP32PYc/phee/F1G3cYLmb0HsBFDhsVL/yIh56d8kHNxxd41YcndKhqGWixzJeuQDRKjv3OHZ7
lnyc+tOPtty5qiCtnw31SYYrnGBYKdD8My2wIejr2omzWPiN0D+u67DAsrEylkpeCo3UlZXQV3el
lSz18ebWfTmMqWw9YzeEElhCWGpnnf3/uj3SyMFnmfGLMAEZdqtJjc5khjygY0xzuuSvINsPSENy
tGW8VaMC5tuLge+1uHzqeV+V3Aa9b6BOhqW7Tf+pZlxuWspdmT5sCdsJHdygH76xomxnWInqflje
mwOv7l/2IQdFWiXmbwoHMxhsvxlVD3gd/1QHJEkzREC5MIuOblrjZBVV2oVjF5r6QyrbUEiD1/LS
y6VHIfmcpNlMJJiGknTM7kYf/vs7hF84VRQQCQuQxb4kqlndqPmJ0BbVa1/8iIyXdDhZYULGMDYZ
UYdO0+cJxE2agVJOpiX6SvYrvVWPEO+Q/X0WwRHa7K2RKQYRzEk4C/XH+M0bXg147ffn7UDo0gpZ
dpeKY6xNYLhyQhQOrA0qUCIcWaxbLzEuRACNuabCb5pHlEr7iYLHRROMAEUAa9CVgznaTqaR+1Ef
hFnmMSwUS34Q4J2EmgIENAb8wdA/apaLAEDTBbpI4QVvGGwNW9YC2Vtd62cCSrC8Dn9QQwdcWYLJ
hWdvf9NthFQ8QFH9de4rZfGWCDDw8At3fEgCR6OGfbADD+FbmQbF/xR2pPwKOhly11Q/6wAhIuty
W8WlJe4BCsOKu+KTZDXAFAxzDI19BpitB/sd0kclDtOe6j/oXB9mW+nRpv7ffT2JJonuQ/4Hwkv9
mC2DMBXyXxXQm9r13rlLP+dq59dR+4io+rjLMHaVwRQvC2zxSe9GtN0+cmHe+KK4Pj2MGmv8T2Ey
nPk6rg9z1UPQmppz4VlRFA33KgNtltDvoV57DWoA+sAZc/30yZ9N60l/cI1JighXI5uCs7lzk7bP
bAErN6TCTb3jfdArwdR/v3TCmXSEOiF39b1Yzx8OVqjTKayUOOfqfJ3HGrjd8s5Jgf9ivTpP9KfP
FJn6JS5o9/JV6GYerbfOZNOoRPwzQsCpQanAYs3dvGNUaLfJOlQ5PnT0FRVHKfdq9gLIY3GcVVys
xFGCNenh4oePX01FIB5EcELF9ty2dhBg0/74hSuVkJ7Zq3bg2QQW5LASg3rRSDNq+ZjgAvKuYNGf
uMJ/RzxtJxOdBQR2lxAIwdusdRebAqDPV3X8qqZYU3eoMnrxMaGTJIC9+JtaSqDxp0p39UeGnDmx
JArPeEm88gxv/9/7mU1imT3zgMlWjUi+LHkHXlh8cnHORCMvZNmo8rZwOfX085F88Be6hdY+IlAZ
q7AZF3T78ubUCTjl7rGC3A/OOmbHSTfX0DkaZ0IMl56AObtuAGX3btTDNYl3gZrXS5evGJoCArsr
O6PuEngyTCBP1PWI+xqVKNLUq/v38u9FC62Oy2GEeiAlQY/PlM1sfGR1WlhXpEfs2umJHtBCxC8B
3umsSCyKLM9xXIo0GCW40zy2fDkGuJivsXoifmsL/VCT+3nTh/fDEIwIVErl/7zi72XSlcHnFouo
seeahkop4HeTxlWNNPf8W17ScZsiRdAITM6KFHU12mQntoYkLYskQWZGz28K+pYAOAadtM+WPO4y
A+ebIBxqUKWHrs2zkx7SDQsRqhBtp4TG5Q2bxgsf9edOS459kev3gTZodxmX+J1Sg904K3H8cKRd
Nx5QyNyFtB25O+kQAAeRyJceQt3QaEX4VFScU61r3t6y2cV3SY+AsQVi/ImhgLTrZWaPYM+gKBBb
s8BxMrkaji3ZGCR9FiTxcW8FCoMkxoV4mHFo+DpNJcx6ZT9DSEZUQjJV17hbxMfoxpDTPBDQZr8r
MgZdqbOv0GurUtNjaIwc8GrGyDXWzo61sGSDanld2AsyGklc8ilGzbu8tcyV9+cpbgB06vtE5qyY
CVCTGM65T4GPNrFAimWsyEBM3glY4ZbeDclI2oKyjZFRxlRnvpRj0KC4ZW/EOB3+PcGdZKZqNY0z
5x/VyQ9IJp14pO7bo8iT28I8ITBOWypUux42YaI4C+Fop/nSjxlg8FGIH48lOvAPSWh6D/FrUSDu
3QQz+5F/3qybCCCXuHTrjmqYbZdTxfnCBvcJkJDi695JTmGVbMaILOy8t3vHAz4WEsPRgX4GrUHQ
kTRWawpGcYwfqOpDy4JkZR9WEWnUxz4ZRUwL5Nv+vc2BanukojHKbGG8oNyR126DfNwx3ujJ5YOE
kr2qb3tCMo3lXb+KJa4h5uXl50N72+g0vk1E4mUK5yTpLApFLmRbO6Jy6j1gQu9+YButaHoknF5u
RkmYlEaL+/9p4IRSlLFLj0t9Xg9YbyXC2AWZ6/YcYX2NnWCl/ufrasP38scmLGDckVv5qi4TX4ug
IvQe3NyfDXziqEZta9LitKaMYkRlzINjBvSJf4xaEhxvTX9uvVYEbAGgiDTyCm9nvHYkRD/xx+48
cvqbyfBtPxH9gVVUPXWU290A4x2U95nwM/LO0PP9Qst+8rUz9jMfjOl6MxEMjKHFoVuaxDUzY4s5
2xLU7MFnYkh/0QDnjyFgdev5CzJ8nRk4si4isA9CvSpZUmWkBP/h1HiqOQxDg27p4h1h98Q/1sYs
v810CjSrqgykafTSAO9BdNWLmBwCbaw06WYzKc1fHqIhZb6RuCnbjRENh4cZLTVXt+F39QAvTHL1
qXOsYFNBRsG5o9c3PYV2aC8MFB/LWkT/ipOmTOMG1ztpPW9TVVjNo/gXXbk5cmd7G2DmJu3SBkEJ
LtyfpRvH3htWXsSxI9iidPLVvfHuXwH0MBEmzhUVtW2Ftm6l8Wjs5apaetdH/A5grw3bag0EC2Vv
F6Wnj+KanScSQOx3PZoTPdS95PLImD7SuDjaLVNrv4TMIGdKdm3CXnxBhpRpa8gcrdkmgAnSp+vk
iRIj5h9r0r1nYtubdUvMMyuVfcvyUCn//8OfrGl4uFxLShimKixbsC+P+8sH1hGjD0nTxHxpqPmT
ORRhEcwKswUSejaVImlduwesmQiLVu/VvOPq1iXWWjqRpbJN/+QTP2r4iXMxrLxgOIR/tjDkCo0Q
NafAtTjuqDpTib5bKKGKgm8FB7n8B9iXnzzJ0fiUTiAFrXO/EfzGvNgExd8Hi14bT7TVadmj3s7u
pB/DB9gG4QBxTnzz+Bp5HQSDBCMzP+1t3CnEyPlSwDlN3fg0Ft2iFrrTXQ5onws1Ig0XeB9WggEE
Rwh/kfbzMM/rOD35rJqOlohTucF/ogdLAS0XKQ0J3JBwr21GCQHj7LqRDefhu5Lj9+FZbPGlgKM+
KfE2Cu3kVjfE8ooLwSpiQwNuyQFGJ8Q+RaXQxJXnw7zudUIRE1gzthpKc8ZRLyMk0ish+xGeLqDI
UZA7Yr91zGJHmmSINE1+SC33Gi2WPh4u7D+/SB4PgN3jN+U+BdBPb72M4lxupsCCS7sa4lhShkju
Kuo+jWJstrDgnVyqA4XcknCmk+xHk1I6KndAhJHU1yGWu2lkedav9WB8fyh1TuY8K3n0yEBk3L7r
HGDiDCWaNMqcDCVLUsz3OVJK6B2fvOL2G2ezgjUuXFe/lfAWWBsZzU22yBQ59Eo6ysLUjoVZnF/b
TXkEw3zNP9gTnJr9qHp+ZaIL4By7bpxDyvQu7X3UbeIy08i9YdB0NYKak7ZS2DAymTYTHlCk0I8M
1PKkAyCXkSnHD1j1W4KZHSMnJEGoyzbK+v/sasfb0f5M8iJgb6aO8Aju2sHqRu7kemrpFYDWh+a8
12bCzVs9+WgP/MCo6h4hZ0/4HTRB5MEBjyvbwhRTO3KaNQuKYTzrLJ7z1SDVeDXXHWl+ZIItY1mv
b5GwE6snVpHLjsTA0TTw4OVVIEvZzF7KAk0PnY09uYIESbHnNfENtvpg94+ggv37EtA2smDWvLln
T/wsLMWCHhId1smR7UQItdc/iKxsmy84MU1Qve/nXzPkxSbYC/A765LCr2XFdLGX65jZk9LGf761
rGVa8mM0sfwmUAVqoNnnSnxHaNtvcSRoeZvPSGJY/qbpgc0xtHAXuzLUGlxoLcolgJ60WjLCDEzG
vbVotb+TepjngrJyGN3N3H/xevi5kDKa5vZGngAN2vDRAemIGGi17+9h9B7+Rx4uUHN9bgE0iakp
s6xi4INq2ihAZgyZemYnjklvNxPTRg311XcTIawaLWMGBICWE+qxbhi8rOFHQFN24klZyAxupDnV
DlKE+DJvneZAoN0SXftmEiRGKcQbSoZ81X+Fo8sVFDoRD0nVOBwsuND3oz9NoKnTpU4zDhvW7+Mc
3kXY3qiIReKBFBkhK7ECYWjFSHQZXESttnbz4KIScTIW6aS4uToAAO8Nse56wUbVubmVFzSRLmL5
a2b+4sM+8Fp8U0Q2bTaYRnb7FVfBVyu7tjc0R4X/bEAtdiKMoMwPX/5PHB46CBSvkN4MZWA3UXoJ
xhIYY7IWIQtx6pn7o/vFWQwS4Ortzs1yh60Iizm5QQB1P+1RHbmdNgg06fxZqHBsuWRMNtsNxNMX
aH/Dda7+aGokVrcxiJ+ypIt31tdY8PMABBVoXRSepyu0x4IJG4zp2pq9A+ChRNLg2mURueDa1mPk
aGdyCPFhf968CfkYj7OwNuCdtNs5zEBHMLG4Iz721yk9sU2QV3CCROMrUXyD9ppsX2GKebT0dOrM
1WTMzSKCUEOsiPePMpjKYqRwvMnobYLXiXsnNbTeGawHTpcfzNoeL/ZtnGYaOsRDy6tCSy2HXWvK
Gos0dI0FjeXFsxhWTYHrVw5jORByo0SxHIw2R5NoYohVypmDMMl6PgfoKVYleyqpp77OdS2IC+Nf
YKs8QGm0uGr9+4oHeeiP0tiYj5ANOvGFjkJXnqyWodxKzkOyd8YvV3jZnuN0kUe+TADdhW91YgPu
xZvtYzyl/q+pZ8I/dIGIXMQrJw72HrXQnH8Ie3JfH3L+wpo4qH9AhWx9i9FRoYsZRMj6RDQQqZS8
83hn72R9D3AZgt5/RiPzJ8rEEza6/zR++Hdd4dYIpTWS+eWolG3HW0TuhtBEvNlyGK/JHq3Vrblh
vpl+iMIcicb+VTzTTB7OHf+wXXK1ZrKICBhl8mL6QzNt94Ql/K6adNhtEa0Hn7T5X4HJx4TEpgGX
pVebA7AgUoX1dnlabBQTp9T3sJ2eByMH8C2g2pKSIpEnB9a1DAk0caEY1nLQgUc4qzTG28wb7p8k
Em5Hj5pK4ybgKQT1S+SMhCOpXV3oLL9zpl2AZ5MKR7nnSXqp/s+akO5P70JNFu+W2oj2r8n1UQc9
n6cD9mCUk+UGiDV6huHwKCm+ZTdtN3z28b1AYaGay2p6/7eaJxQBndtS4R8z5xXl4jn3boM+Ty6C
Q4pzO+t+z+XgXHNmhgN9eHxe1NauXvGihT6lhq+ms5hr1BwEyGnZnN4td4XJY3Kfp06AOmmenn0V
DmQQDromhEcmKm2zqlzNSN4aMI5EoDS5pbrksHlkNYzB5R6mHEjtFHDtWkxqwZur9DwRD9MqwROp
OMaW9Ki5YGSIL4QzWQxZ3o2eTaZJfM79YmUsMRttlNpATjza5AAzvyNOZm/Knq1IfJp8bdj9Kq0Y
0lwICqhXHw6GLl9fnbcRCLW4VpXQ+gn3lpxEoMf+vQ5fcaFhY/CAgBs/Pf7H3uY2ffwu5qp6HUsc
FZHVshg9A65tXsxKB+EzDeGekYkt3hHcSMEClXKZLu29lOT/fAjiM5xaIRFkvvAcD/XSLuXsPISk
X5n2edMgPi0Ni+4zrR6m5H7IcY1abDDsSVwPjeBTRuK3T33OSDoxdla9UFWS1CjT1tByZPMQ6lS4
zklfld0nbkE5x+bpuepJQTE5QVZc/EXOPy9GcN5srWplQDOePyYbYSWMY6Xy5oktidEQ4TuxB3B6
OZBiJyRKcY1pGl+KBouPZpTudvRc0v4ca9BmFsQU6IkwHdWpNra7gmbmknPvP0e0p1nWZgWnCtbJ
w9rBn/2xdybLFcUB0+NYGx4D6pLswsUVrhyqTBjVyY/mQcDNaOusogfNHQHpXnQ9xBv2+gZZI92C
SMyQp+7cLPhH2WOMNFd0WwOU1awXIZaPKLQMpdki4CIsGc2gylfsH3/bZMP/zCB/iHYLshVzLzrG
5e2DZ2y9oEjV/spB8g9clq0EnAwGAWet7VTVlB0fz/8VHHNCvrf/rqRV/aeTzj85q+c71i+Tv7ud
ApaYM3KXwgVM6WZ0bbvMk1838lR13QpmHd9fiAVbW6wT+d3tkEIwNt+begMALiL5zyp9WiZLlrEl
pVu67iha6Hk3MJjKxY6MaLp3y8Fpv8Nz438V0+BQv97V0PSshU9G0sI3IahBQ2xPFiylDx+R9DsO
OZJTUeataJjd+uV0E/4HVXJoIoCe/zBPoNZOvFwT+W/tdBbDQpjmmnW3VSORPLGEeWPD8i9mCAIQ
5qLJMC3u0gVhKTRFmw+77m7Skk1l73XwB7SE9c6Ex+Kte8CbTXPrOmH92Y3ezFJPcVbGFoBdk5R/
Fkn78jEtsHOYK9h+WV1zh6ysNyLczgq3Kw8EQI+pYmDsguRgDm3+kVO/X3GVMpu7dsloV/bwVeOq
vBcaPNzd2QP3E9A1ISAoqyxxE1NAoshrGvyAbEOw0POABtZg+oAQQ+FvM+TV21D/4xVna86qL61G
OtdzG6I6GXvMsIjK95CGI5TCIaWn8UpBjeCZ+ep06F6Ot2S8SxL+81EOSWcLvYr/umO0ZuXS2PT/
DPuj9V81PDrcqJCzLhBqlcTZV5TbJnJHWcF77e5xgRviEaKO8O73SHR8Gtw8/oi50+kmRltOFUdv
RtCt2sygjcUSLBWJ9LstMqsm8vVg61GJZVVn+k8J6Z3yK8cAUWcZzaTPvY2hKyktHxRDP7b8cTAU
RqhlgcIbhTk+kOJJQ1zSuseDsDVQwE0LTahpUgJVXD7jDxhfhAOdB3sewEgx+zMZ/4wtEyd2hrqh
B6o1ciR4QSl7f14Uf1Q8OBvDwNCA3YXgyinWYWh56aiesuGD8kGrircgL0+dpccPM667UVGcsF6k
H7mcRdnSn3JvNtp/1xmde1hal+5d2kCpSyWxJ+qSFwXyC2gfojUG2jbgEoZqugp0Y1tZQpayeogK
gHgI3jEflk+aT5zinDnUKTN2Snk62S3nkcgO9AXEAB3jxrH9ClYHzIFWujrhyXG2tDffaGG3p9GR
CYGZJ6/zYRjh6soMW30XcbkwxQBXIFo9lnwKV3WKTgzs1Xfti51Rz/S6LXePkGePPgl7QZRsZxau
y+YSDDUIZejjsTHC8m6WrB7IuJaHUMjxILNhXgepbd4fVbVR7vZLfd2j9nK7wX9C3nZeglLz51jF
yFlweflmPbSCTDlrzTxX5Yj4Z5xI07Df43KtWvcDPIOUgKZIaF5QMKOMbLtXpr6X0enxVtWUtrjk
4SNs6siD112VwuXnVwbLYrKSvEWs8zlcN7homRlhlY85EEEIZ1UrZ20c0p2HAgwXpaZ99I8sNQEv
Kd2PKwW8cnhaLj7vQWAa7HgaeBGYqsKH1o/leYSUsvOhrb6lk4AWBtGjKW6PcHV85fMZ+v2Lrj6a
/B7e5mKsaLur3RyR86Xgu3MVVJVhMTM5tmThg0mmiTYPgfdFIAFyWRSCbMs7dk3qS/Aw4s/NbsmA
kcuAO5ch/upKXxs3HTDfOI6IQ8ZHV09HH+ARUxHddcddvj3SAN4pi+RvnnzaVPzRjPgFofyVh7Vi
n5CyXKC9rX+SJuBU3/qKE9ma+z3vd8MrsRaBYu32o5Wk09wEGxQNkbQYzau962cRA5+BUEGEPEmY
o1qaTJgcuzBYpKMBgILb/o3laEiFki3LZS4WqRfhZbJwdCqACo7nilSbTitmAF3tWWZ4mXqiTK6l
tSiPYI8Xo8jGBKlizRK0RojiALcWTLL2s+z4SjROM1+oNq4lwzgdaY8oJKGwwj37ZrCOjL8bIfA5
WCVxmez7UKXebWZ65DfAgzrFR9OdaP+tJsN/Ix7WlvytGOrShA2uGhQqpQlbNYwxz5MNlcBRcaE9
BCw03XFw3TTQrNJbN3YvQ9dCWoL4UeAcOZjhavVJ7qfKkP7eTKwEm2cMRzhPQu69camo85TgzCSg
CkLyqF58SMSRDLNpCadeTXXXvkottqmBmIxPKrqoRl0fIkeXn2yEgoqg5kjvVJPzfr6HisfN0+Nn
2R7UgI45drQitgDf9WqR3+dNgGhLkU5HKCiUnFOzBCdHB+q691T6PuyDtgHF8gpCOg/bH9mhxvDq
NzozESTGrJCVSGceF6x2DMIp332Nc/OvYp2x1niURiHW+MLyv2QpLObGB0RkxojlzadFFfrEa+xh
oXA6ggl+HU4Op9NaSTfPXnclsPrx+vMfxdonFEOQzkEbXGiRlTz2layHyQ7N0BfiZ70x/KCNgRnw
x7SAXJRQ+pN7AdtDQTWXQQlSynS+JjiGB8w3wyHf9Ux1eAYm1ClWuOs6Azn1a9ZO1Jljt0BmTrkr
6ra6MGCFPIk+y3hZNMd9j/GQZfCfWruR82xK4YSXYjtR2WuNwckVjiizallOzY4OIWK7KY7SbkkD
lPPqCmN1ICixknmGlUPE7BTd0f2yS6MRCJ2IbFbrF4W76+ArS1eJAqxR11/vhbPTTjSUv7Bf5pAl
8o+8pzttTphl10fqVF7yMAzEMgRVtj8wgEHdNM17p31BcaJkRN6VzscxAp5OY/JZf/YaR56Qgg9x
ewuG73ku87lISFPncZen14regPp6uXc6pEEdyrHhB+y6QCsPiCba/EaLF3gf9weMgiTwvQBj1WL3
Kz65Pc2iQfgvHf7fvmh3g0mMGvtGJVENMcb0a2uc594xyh88M27Rt7Cfd/lSULifQg5SrCcTtU1H
TywSNC1s7j8z9gEABD+TTv6wDK59xKKg6ov7lnGi8IPBzLshz4elZ+MFdRP2R0pFCoh+IiPAA374
Q5MAVm5AJTagDuTR20P1tWJSjVM5KKRaPW2frZEcIz7x0lIAuUkk+sjWffyo/p2hgpej7EPY6bY1
BARH+Xt0+2/nr4TlIktyJdnPCcOnsNZakiw5K11WfcttPTCGWR82O5vNw7eOiQkyjj2L2x8/M4B/
demow0/DthFRy0Uzdtq5aMXz0fn14Iy0R9x0SboyrjOGWHIphvyQ113H2oyoe4SUTLZ50nzyQp1i
Rv8n9/X5hLRAoVqs6O+T847M0hZIw83AdcBnzLMs35d4NmnH5TrNHAVcUySsNdkcXG1Y/UuGKeWT
mRNybHSt2CQNj1vUu/R4ag4vpH2K+R8zGmvADvJDl56p8sbOq16dFsqmUDxhZ1WzO249hqHbgx7U
J/ZE2uT5I0OWKQNuwPwQPQd0Q2+ZjxtlMVHVURXcmA1UHQFbR+1UDwDgE93okjrC2zzN+U9Hc5eg
5EcCviZRjkcm9cEmob6ZmKE03ULyjdH4VYbMg4pfSGo7qgnzDGbJiawcSuwRD4LURx+ofiBhCm4K
PULSw8mcCKBmwE6dRKqwokXOImfu5U88T73m23HJ68noiMrN5DQllJcqg6eFiTkog0Sa/rnVBjfl
emydBYLbAMynxZ0Zi3eofgEGmOeJkc8qrv9LEl4tlc4/wL1VZ6Waa92cchPjA1xGIhVeytJvLBn3
41YZQZLITMAKk6KIgcmnGFeLaT27ouhk6PBiv/2UDZ4Ddyr2SozVp0XjFg1v/SDwE/aS0jQKvjln
m06/GCYnDvqdXLe81I4nAm9RRyfDTW2tSiTUBuyF02LHkBoG4w/dhoxR66/ebRId4zL24HULHRPh
XChy7PcBToyPMhBMh65IB25x82fyOzC/N/BYV71ucl5c76PIjhnRGEEk0O5W+viaQPXkSqVmtM3H
Nw3+i7byfKPjC27bPN9GSEG0GRjzgr5EZQbyDLzNd7RngZ3u0iwCt4FPVAY0fGDjwPNUjUJQewJD
clsLHXEt7J1ZsENP2Z5XcOXnyuAqc/qCJZ6wxVA/eLB14sPWTrAxguHi1OUbCwsRPCtcI3On9VvK
ydbcpa/xSQede3irpFloSu706li21qhWcvw3EKMGUGsPGP6oOWO6Ip4B2Hz0dMspDWOiJmGlIc3n
3w9zTX8uXfN3pGVRVPhrYtE0LrVqfqkK1mCbH9DZf4IC7dcAAqTWxpIoSrNbygMNQjRxU/LFIq6o
BuiiLP/2AFnCv5eVuz6o1Hp6sj3txNvnkX5eeQ7DppU62DhABVQ+ztnVDH8w16lfr9jGsDYf9Ceg
PNul33SebNTGexI+yzDXuJM04M6Rdvr48jDjaSBSXtgi6rmdE0047yC/wHD57HK9SEBrXVhRjarw
L0FoQplvzAVCyDUObY8WMTeu/xukK5CGjlttpzSvRRE0zf6v22t9k7OeQGi84g6Q9kPvc1YQuihS
qMHpJ5E1OPD9CDOkeBGqJT/TE0460wlBJq9BLDHKfIL5/Y8+UMDzqlcTg8k+JNajPc2HbgRHQ3/X
/RT3QtrA4+5OEOzVlGVBya6YTtMKNhaTsxn9xpa8sZGCD54hTEC+V79P9t3Wzo5uF2eNkg4hMJNq
pOiHmREsBJ8FlNOxG/UIRnYMh7FZTq0OnoZLHRfatgLxyp86MrLkkrH9F/QidpuWMDTmaq4INtWT
gT5BUZw48Yu2fylfN3r2CmWC6f01ADwXKrKcyP1AS8TDcHrylKLhQ68dD9pP2ecrV6u0tCKwETg/
3TaDB40GKimjvJMCnxvgCIRYIu6p57EPU3mftuw5Fm9tMqvo45ldin5Gn6Bdl7YMHsQVehFhK4e+
2350jFeimoY7IwmT8KV0nAK/B7Ow1hNi4pLfrI++DsAw4Tkg+SK9pHRRi8X57IAYWy2SnboOVq9z
WGqlEqRzpL86qi76jZAAwW6z25sJVtd9Virt96dwntQWXGcARC2oqj/kQwxA1F5GljZN871zs1+6
LHOq6fxhcEEr3AlnVC8mlV6ibcNA63PZjQIsUjavK4GHbZufxUoYd4EbNpnv9C53PjEXpFt2h1bs
tWYWmS3AhkX+1gzNz15nElCmveUWsl0uOrlynzVhiFJT2Ek8+ETzwI5gQ/tW+FtA9sOcQ0Tz5yfe
3QSJ3hWOwtkgrMRVX3Osc+9VT2INcfVjqARpjahfk2qP4ijv0vh14dbmUwjZOzQ40tSLD3p4/YZN
kvPlRRPZcpVXD1ZgC/HxbQVOIIEcavw+USFEC3RdxOym9WbYpQEB+SpJAC1la9W98iCC+z3tnXIn
6HvORXWpWvkOMe5f1rq7aQVOYn4AVLLEjyXU/8uGMmDaZuuO4GqjuhLE223mqDyA28233nZRnNZ+
qt/E6D3LPfi+XdZWipnLeMEqvl96NFnBp8Tgod78ZXQ9/rjdyZjQgglFaD3+EGKqYbQuALY3/IXU
obzHN7zRodORCdd0gPxskg8U1Ft/9L+QWIQ0wdF2IabRxpOSE16EFAYhATdyGY3BO3wfRL6vUwus
R/QQz7D9GhmDISRgkttmVrEVET9GjzRHqhpsBBfkO+SvFkdFbqoqGLrODV3OBBuGdlvshZiF4FZj
Gisbm4YZOU/1WKulNAjKrjUjcJe8wxtny8jb5Q3MsRDLmEQvocF1c309qqvfXcUtbA0wTSSulME6
iTjuy8ad8jU8J+90MwMdGJ0aBLPXgpeXSkQfeBPN8ROhfR7tWajRO00e+kHrmyCbpvEfKBnNtS32
iy0qdHktpWQdMNDqYbnCPa7oXxfiGz9gjuDjeOCtbSio0vsvPaK3AvrHL5A+ZyvElKTxsJdefDHr
Mg2ToBkkJ+DBibA7Kh+QGtpsBvZzY1BXP3iguKpjLfgxbl8Cx9COOr8OtO+m4h/Vbttt3ni4v8dQ
9fRNgdGHAOwezX18DMV8eU2HDG5Bf6UU4Wz0QiBc9BO/HhOqT3TwuQQDKuiCCG4RoMXk/n2aSv+A
GLWx6X8kA0kEolkamgFz5OcyNFzzCssNoOMhMcGw+jts/L/7+Jrp/DImqMnPUr4uoweHfQICDNi4
QrcX6vaMUL5wnfULrwfVSemrIiUNrT9qSZr8QHsRGz808iByHutegGbbhAq+KqKldzS0aAk1AEfh
tllKYV7aKXsedbJiJS+qHm4bc7tl8XNmbwmj6gXS9zU50pbrkG4AX95q+e6Dqmgf2GEllwW5Ea//
3NdgI9zwU9IKbBogoX6vuxeTQZ4wKlOmjgWQ/tQj8dfNBHDNzQQ6Cvcdr47c2v5xSEn8isyvtZbX
d0hIyCLqnHdWcEQEjhFJUdsgjbYXdfsw+uCLJD+owo2r6420sKXZPnwyhxyVn2FXReXMnYfj+dwj
l77EK4S4EZqIR25UX917Jt7vYYEXLDfOh3l0CbusaSRuKLmKATshvrqJhDHtqGVRPxHBCxt88sT9
AYLJkNZtyKPLce9S9Xf1Rexumfjm9YgKVTNMhJ8LWXg7qhLPqygo08OeZcfnQlNiXfvDrA44JO55
vpl4SHNT17wisa1vMB8LWrkUB+zDTw0QH/wFqdKGfQeuVhOJwKGPfbxaS2efwuP96/t3wLU+ZpKA
fybpT21H+/l4oxQeLWpFpfWtHgVabw0hNoiaZtgNG/TrHCMLew7Z1lrReU7id4ITgGboQWzJFqfD
+Pd8yTNQyLmyulzB7PnnUY/8YqOxP8qe1Iy02k9XJZrCBL+gTXwSqMcpmW7k4qrKcBhASyYRpL7k
lyq0tjBaiJgTQCp2ncBzigNSiYTJnKF8h1zOAD/9muGRhFlR2LXjRGU22GV71hIa847rjLOe65nO
o0RedOkmQiaE3qjvSWjHvjyKf8yKj8QkPJ2CeKv1xlHR5tt8fcdDs/zhRw/o4XWZtWUMJuL4KpVj
wuxR9BkAE3RiCQhL2b8FUvGS/g9ioXaO0Wigxqikz08asnlDyHtaScqMla8OlmcxbYE7iw/MuYih
XD9+AwDEnqVRlqSUzRSi6uSUqK/y1bL+F3/7kb0KrVxk+AGeQWjoKi1I911O1pDuZNRvRcMvx53p
DuuvIqKCWco91tke5a99Cj0bbsLPB1PnEjN7yyJWkUgfJQDi/ycVmhjN4Qmttwe/+rIjnhtq90Jb
imOSHRN3wyVRA+QK7BDmCvcR/q+gaToVWHs9YxhWYWpD5GXD4aCPthfIzTy8kR7tklD9xv+R6JLr
6fCk6oJKgj8K4EtCPJFeBYhBhthl5RGySrHrPHi4dSFgfc89d/dghkU4iu8oP0cFXaootVk1raIY
dVxYuTEyYrPuOe+yrJr6P83Do4kxzeUyDex3/Oyc44GYinGy66O8dySBXqS4fT1grM5ntvxIPrYb
Rn1yBbDse/u+P9dwoAhPvavJBALs3ACFdCMvH0Vo1IgB1GJzG3Wc2MI3sstHJWtVhj3b5bzLLwz9
3o/PniEUDPy3CYmwzhh3XA7YFPhuXOWbvPHG/yHcMEqzgDFVKIc3zkPp9WLgWG8VsqtJbI88bWk5
6ZoXvFj5C5UIKcT0EhivBkNknfwl4tDTLKUqke6NZXsN7q5F3pBGKc5DLeVb9fUbY4AC8bq9/WNa
4FNQVfU24eX2iEDJdtpcpnU7mQ6x2H3pCH9pxmCrRFesZADE7VtocKOwNzJWRtfe21I7v7tu4P+3
nm9PVh1wujRIIl3MTziriAgC0K85e33hV/CmwTX/RMF5ufUE/mYbz+C5fI0cDqPGA+pOn256+W0h
C4AKpEVfxz2TX1Ytue5RkSkvvlxF57o6DIJzhCaaITT32cnTFVWYjsR+fKyGpQmVbEDV5jPIlN5B
XNkVZKPEj23rAch9x675MvpqNwIf7rQGzJufhhPdEtnb/Es6hx7omD3YhlYa1K0Uloqgy8NLYCxF
JIBccIR5oqAYPRroUrNMlmV+sL9FsnZtXK2oaQ9qyBH91PUYEdm4lJCdIYsDVFNrS/aymdjcHdUp
PlaonrlsXsc2V61w+iGSwOdyKa/brKUon+nwlsrH2dwuIBAGRzgP8QLmU7bBCDOnlQXJwCWPExc6
qRwqCo2o5iW+wyYD5MKnd074+3K3WTCJt8KwMssQk3hJ4Ehryj3T2f1hYwptJOkDZZYIuUCFfTR3
dVFqzyscqqylfzDqBklT+n5D/yOcAsX8ljckXKn4vS1g+N57Tt5EHski3yMWpRb4JBsuC1dlQiJ+
PIU53asGN8YWLzL3jMp19BWnffcOBXg5qJsrT0Ld/1sPii0JvoF/b3/TdVP7vIcmLlB92Xfj1evo
UyJCaGkx51ZDPf+bzXLf2QOio6kHcdV5l7Kp9Zajql5nB7rLhCVRmRR2gON4w984XDWemMQUsPLF
Ivpyvc3tZJw0WP40xGEmFjDeqFY7/Y44AgV1IKIAMSV4qOVqs/cmNLQDwykl0XyBGtJDmq+NgZ8g
h0F52yyL4EXS3BZJX7ZZt+dCl3Tr5y/0ZfLbnrQk1gGF6M2c45Ewm6Un9Pejl+3vrs4lO/iYTjxp
ldppr7OEmdMCTp9U53EN9hjgM5NKKsaBlDxkbvT608IKgFLwLHgg8RTq87zMByXg0LHyg4jefiiT
QRYr984byDEQJscI8qEN0+a6vq1zbbE6p/rubijrjYurccxKq4BBX+9EQrTvfkebII+5otH0Ijwa
VZRF/FQ/FLfDPqgFr/ThrF1Zd3eSxqtQgX6JOglYHyfQ6FZe+2OLjqoZ2UFroyaUXtiGhkI1OSMy
lJSOvHrSsvsiuFEz6kOsbV3w0ZFh768Kt2/YGBiLStVDJMe4VOmAKkcOps+6ahegR441tS9pLJYV
AtVq/ZSIMscLzpFkcmW2TbJbeLBc6e0VyqjUCW0vIRZmMn0MVxXS8SpguyOvhP0eUvRAh4WDbDzO
djTBoA8fMJp78McXq5z6j5UPAEa+6Mv+GOWPEcnjzA5gyztw5G7i02VgTDP1I9obpuL6whZEuOX6
uaX+70o21AtegdEUAz68TuVn/3uzRzqvMvvje31Nrgxd096mH/1KZHYY04bWGbsJzugJzdvTdNm8
ha8xsyuz9jvcrkYgkbJSlftEFJTgvMkM2ywiuSTxUeOCf4+854b8gytmb6SRHVOCmUMjHxgD31Hm
I8WIpa5jToo9HUz7roteJqQ44BRJwzwzhZ68yhw+2lb1R3mFuFBW2fz33wqfXAnFM5/Ji4dyLUAP
vAj2Hd5mtLNR6K6hAVWfda/56aZfE8M0NB/zcSg8sae9QFxRSbTZVGJVh6ZmJWbxqdCzW5K2NH9g
D+RYectrj3CAovkcZP/CznE+lFDGF0sopJ0P1uSHH7G6XDMl8sgCpVcrEyVmcbEfNFRGwCf8FMbL
ujTGNawCdztfQtOO7Uq0EGP3TB9CB9UEZRTcaQyVMDTIVDHnvUKAntzjzPw5cLqdCE8VVeR/zj/w
kwok++BoR/rtBKTYr82CbctQJadtmD3PexcPKp3ZqZPJ5w+Yo5inP7fkAipr2EI019E8+wlLcS+/
eUK+GMfOLYYz0rubcHQZnbhlKTp5gnkoKq9fDUwHO+pKk2R6+yfrRTlGUUZGS0TtRWV24nukF8f2
uImcYvIESibm70RxLlWV/6byfOP9HeqzjOlFbualzgevjpTR0orRQ/gQGaXvKuiEAwU6q17YIryp
BoEB3N8I3y2pWSxwFdwiFOy+vfj6LimviG6zgOURBCUErfkfkrLu8mXewFZ3SOrJjdV2grfN1ufd
REpe4Yn2seRZdg/x12eidwZfjpD8VyZktYNe2ugcF2AOWnnkVZplSJDoSyiF/bBQbPaB5oNzJxPj
pt323ug62H95Mwi2CizAw1miMMJMqIX2c04Bz6WfgpusY7JRFMy45zQr0du3YI2XUw1NHXpuSY48
RmIp1VYNITCAE/Sj+xN7HhpG1WhQH9WDuCYYAuDICTZwXIwslPlnIqeMbrsmefE3p1Xkuo7taXVB
bCKmCxe8egQmg63YftvAe6U7zn6MmxsC0kvkPYAVBDSAPcYDdX/vyGwt4lSbRtfah650IdVtPEsY
Y/+lhf3hb2fzIwGGEYUoQMNrBIkC9aWtuFK1qb22vjK5dLsXAIclycfovp5e1gD+XAqPGpBAoZCs
q8vb0+jhBBTbtxbCm6Q7iNMoIEqoSvxlWeQcU8wjCYXZLQn9GAt4g3SJNkWshxn2FZjkk8V/uYdI
3MRiY23U9uD/qgD0WB93zzxnXvmicUhSqYJnn8kP7REaW2EI/GCWjqHsruKIhO+ZaFv6TUzAYTGw
IH4uI14wtvj/XXi/j5fDp3toxSBwwEpgrIwg7XpJ5ZvyQ/KaDAc8OJaF/GPSW759HQ5dmt0QgB7s
Va7aC4djuFdpr3ccQFLfZdACMn4uCjEVuHUHopfnjgIz01vNoDUfoMgIb9e+CxRlXnafvvNqeHzJ
NLstLn+n61ddyVEh2LeHM0miVIyVWUNaFW+h+W0raCpqJWeSIxRJuOuAOgW+iKwzVfFxngln57Q1
czIHaFaDSLB/oNOtGAoL1z1Lx1rRTsE9L2GzSZEdJAqWw8MBcwpkqm9ouOIfljUmBTtMx0BpqIVY
lt5TmHTnYXZrWttODClUPdNshjSHmOSitk5DHvc08wk366u2Zur5IiVyADtVo6CIb7X6gPKiBjoD
snDI195jMKZSdZ9Yn48B0+V2dOmQG8Gd2qVBDqkINMasgS9YQ6eGuYvu8F0N8CYuA/QsPaOQwnpV
FrUhXU4wNXV8guU8ZYTUG0Wm8SJ2YNEA3mYyADPPz6+1HNIHtCgHrkZXxPxNBm7MaRao0IjG0rTr
8eQbCilXSrP3Co5kkwTSSi0iJq1kgvNxHT2ZRfEAGTSi4uJp5W6aozCcqe9rr+lcjboe7OhcSgRB
GqEgEQMkXZTQ0YX0h/sO2Ws5ISrSz/xgwpkBnZiC5GNl521VOlixuiREjQBrrQNJFReUsYU8RwDh
e4cRzzKhxe7mzhYQSFWJHtIu8NHnXmqWcaI/Pc80FZ3dazJhW1hnvYt1yZ4Z/tfdtb//qx+6+IBG
P76S7wlhaBpycAHPcmYJgyiaeBV0suTr9YgabPKAyeC0OrSb3AEsGq3udkc8WM3ae3tn27u0/CfM
ydCB7DGxfhW6DnwFwcyHx48WL+yrBvkqz2vBFRtORDG8g6YQYBA+1uhERD2KbO1rXgDwcoSvgDdA
wvJYLrAsWKiTtT70xr0KWssAR89dyUHV5qLYn463JIcj4HEvMlgSUJrX3wHgmN97J0UlVkR9UEjZ
bzcG9Em4QFGO8VZFh+ggeDXNqd8YHIRXi+6Mhx0X3z6bMIUhAhlWiHGtac81DpEq1tK1Mm/HMDXh
zNgfp9uGrHbyH3ZmDIHLQ+YiMZY+cXNcjpAQkY+tczoGjms717RpN3dEj/DfuSIxDX7HDyhFl168
Gut5eqpm0b2l8LXhBoApVUD1Qa+o4esbXxXig1N95RavKPmCr27km0ytBwhmKtpCtnwdi2dVJCPL
RotiRtCrMpx3kfaBkFAXC+JtssKuocrD0RXoQmh/Urfnx/BoBVyleJQUF9UTTD+NImLlJE3vAA4u
bEdvuLcmL14228ediGTbUZcjvD3QSHUyCkNIi8qGxtkKz/sZ07b9AQKltKriX4rtDhryw5gPaTvL
eQdVc5KVQLBmZ0uHQgsiFp4wcyfJFN/D0500LrCap2bCVyAyGMlsULQTMXzqdCdlfUg1V9ULUh8m
mKdvORP4MMyXbBgmnkP59gaUC10syqW37wKqoesCUIXfs/She6qZQLX5TKqVlm+Hs+L4LvPBshtj
QxLRBvBK5qs8XT2me9Xe9zvciUzcyrCXCh34RlEzZhpivJC4Dxx+Bk5U3OQsMKXmp8PV4hLcKSVG
HgamU8AR9Evf0xbwxTcftAMFrGoMfGXE6yes1EJymX0nXJrEX83Xxol/sH7IcAsUKzdbLk3Xp7ic
v19au3SRP2Q7Pb6H5e4qhrP7Jglx/ERuF3l7l9eEPE3huKbqQedORcvNMQV+Kk8Y+/M1W/h832fg
t4itbHAIILHl6lPVfa3GbQUdTsfaxg6g3RCS/CYlMljmu5Z4QVvx7f0d5W8YEPo+VcN4m9Q8B4Nb
vCEpD9/cg8MKw/mvKTgIlnwgxqRf5Mkr1/MdzQ3UKyk5ryaVWK29KwZRayvk+Ss/AfWZzXVGlhv/
EgaLYYssq7feBZzF6MCSy01B21IfSPu8QRvow2yo4i23Yj0FiHnFTEnSIqyhKjJHEYScmGmympSB
1Kfxe0O5KHODCZTCJts3aHl4VvWbu6Rov/21a3EKQV379nkEK0Vy/PY9KsivCPVbLd9Mr/CvZlLc
kdQrSNojHHptve7WMug1Bh85WEejZQDWx4j7Cty5SUGy8CuJzyDFR9UIs5meemMW+Sk3l9ZgocH4
0e41beoTPwNQ2bTIbHfhhpMsdLDAFCSpCJBdt8TxJm7OzwWvrz2MKpxierwVJNO1/wbNWmOUr7PI
vp29Z8wTXLub6nxGsWYuUyyqF7Ta9YyhS+A7veCbmLKav//4RAlNm/d62lSJHR6lTjVM9Jz8590f
Cb/hj8Qt3/xWyNVXugrupopsdMFcgRgh2ZuPsZ5LwEfv83KcrktGIUfmvPXIpdiOluUw8YbGqSV+
Ds9ke/XoAFienL7L9JvN9rWZKTutjaNSZLc+8oDJINaHbfUiGs/NLAvjcksnvtWb4hjNJyxcYaWv
eWOv1YpxBFa5ozz2NM38AHWzi3+IOZZj0f+ow1QEjD2zTlbf1YTeLcSIcguZLhCjrwcbiavOQhr5
MFLAkueda1QIdvDSJWNW70I6WJelpbisfWi3EPgb4aEyO2XlyWVG1VXwA13+uAc8xh+7j94xEoGy
+bu2EVP5yDXWJJqxFw96+ajpIDIIa3wmhTNmcFG88aO0GhrKqtsGaZvzIUDyL+ylD6pmMzAfd6xq
eAAFd8OKtey6aLV2alCSsIabZpmCFnYV8lVSb8rsOPYsky9FLDBIZ+2mm4wUNFOI/sKPdvudP6j4
wN0j8BAyEpEaVCCjLNaUnD/dx3KhA9kCyzjIGKtf5vOcCFKhGd+kMeEbDXBJRF/18Go8qza0k+z7
SEsjzXbE8QagQkggET5kyybPnI0NEUetzfpVcPa4uCQvRUGKX/VWd0rqhYp6HV4wajUiMsvt5DRz
Dek9zfB/mjMyJifzLNCdDgkSHf/IGsBNSTremPsrQ8NBdw47aceDq4SPcD8fB7KzBEgjOj44FvCM
n6hu++ZaHMszEpM/mTK8cvaflWImfSC37YnMlCTQKMDzlS0Iq3VZEeGcgEeUeZ636KVaoKQihpsT
4Rs0nioaJKP3YZ2dL+KHHyekGkiUgYG10Aopr9t9LBbFWNYGA5agviBmHitG7EToLED53zZPMBhD
utm1xge1wNW5Kn2NVKCZnt3f7Wj0UBc+bLKaP9YFQ7PxXmUFmImUFGWvRFG4OJpWFvW5w1ofZ8vZ
AfYm/6HziPLf0i/oeEVnjgQZ9cjcHFgQdzMpaRpeIcO77ucoZYCmjeHRlbmugWtUDuLeJvxznnp0
66ggC0CXrPUuMaNcYKZFSZZ3NaJtduYFLUHCAywVaX/XdjAkZUJU6SYk8LzMRzzaM/3MPKd57f4Y
+vikNP/l4WpmMlOlHeuEQxeM2bXvhwbF2ypgSbRGUAKTSfNEA9jQWljwpn6Gbefj/wIcjWrkD/+q
KOyBbOCxks53DCKcKbfJADAWW3QWd6a2EOK4JJuxVBhbUI0FJMXSqGk5tPAQHJ8TjP6ilySYvX4u
h/OxWkAXd3hugISoZUKd1pZx78EasLgbnnmK5/vNMRUWUN5a14rv0ojwk46tlkQ2YDfaUr1s6kib
zXDKKvcb5+h5v3VOxC1pK6AzFjAh7HprVGFAQU/a1nq3Z+GaJhj/VyYlkwsCPOl4Euw93pWKSgBB
YzApjR7KU0IrXkqlowMilBamTp9v3D8pHnHU/FxmlgjlJQP3q4xRm7j8wg4h7cbAQPhfVhj3ZhyL
zx0NeKG8JXQLAej4DFXWOPgUOaddBILjOOUWe5jVdTgBisMrAOqNGPw6f+pmF+mFr+eSy/wSiCbR
0TNIW4kOLnmZvNlhVgy01uiE4NnoWvlgGAf3ODcssyUOJRfSxmPr9fnKBFzCwPPviVGIXy6cnHP8
pxhqV0qSyIRVdI28s3PJLfyMV4ycDKzuPGpNlVnSnz6kYmR8bXzU4xFq89eQU3btEmSmr0t/uqew
v84vxTJONTUpgubF+Et4DC6A2W5PZdKwWfq70FO4ugQTzjJdoOr+YvYoFu/7mcd7RRCgeyq9v0pY
I08FAWCqGPs//ibozh85xUW9aJeILahu54CmtEQxVoxfdD0305gUpSdBYXifUnVzpWJw4IXf3mj5
zCb6FfdiX6h+taJK81KdMyy++Hvv6rkJo6dqHORHH+R6ipCF/N/9PpBrxGLvSoUKyUlTv4JcNnqJ
RNVVvBBeylSPVqNwkUHi+SGRP10b4kpc9Y1KPXM4SAYsa1NcsBjszfU3VDHSHIckbCsOz8TV0imh
k2yqrTR35mOF3QGBJ14MfLbwT89dhD1/EnpEL3btNxaYbjT/+Zve6gzARbJItWTkiTKoRzOcFXis
ny5wyLSCWze389waWUlPgwIUfBkrHxmHcfnwybz88Uco89MF6H+thWpFPOtnMc3B3goVY0gcoYgN
Q6CjBhethqQ+f1yK/UqYeK3KtXaXYt5hY6KizRDZp2jgQcTFBwJc/7HWSJczcaBhZJOhR4ClngCN
2Spt4auU5jWVtrESKup931po7ibzZ7wISTIsK2Tq3yLSCvHeExcJDy7EGypfSeZqIOA6kkKjx1ts
1PEKOP2aKtxSw0Vc2r0qzUn8NASnBoXOWui+uecDW6CB+NA1laGw96U2cQpRog71Sg+DR3k2WXcT
BblqMFA4yJwTg1hUvAhtYh6MdKC27R/O8cDJea30R2COsMrlQ3l5CCkB8ekLELO0PqFXSyMYbDnD
1aBqxbPrGih67nY3iBIuz0OqzI3HGqiCVwtx7ECJCzlZupaojMdDIGRxTQlQnQ0uMQJ7/UDhQBg3
Ite4uqA7seub89bWkXbXj0E4SvReP6UNQp6A+k13ZWKFmVz0Er6X/5klwRkyxfaMzIY3yCQNByDX
/OswtiaHOOysxMTjhxmc1uKnP5OLEyNPxp8ZySGgcL0l/2cpBx6sqFjOMqm0sB73A7+LoVMjKxpI
CDaZRqtU/XqcCuxqUo1sswjedCtaYxIiFWp8/YYz+tcQOxJI3wx3AtBLoQmem6/ag1B3s9MLeJ0C
DNiGfsv5nxn54rNNUqAtBuhGe6wna4t0Q2fsul1efK8dRy3Z9JlLEytD72qAcwEVsG/HTjW4FnKp
WzWuu0Cj/g/d4K1kOlIsi76kit0IV6N1id88QKR980ninFtS4lO0wJpqH9NykloQQGdDn/UMIiqD
jQBPlgccd+xnjVYIKJK7JDSDuuXpgiH/KdxUS065D2Qm/qUEo31/UjHx3wTPFY0iENGlb+eGjJXM
0LsPbaoE2OB/WM3j9FGf2M4CJ5paZIsh/N3op7poZaLFYd++VeWVkFpiHJnibqLEdtfmJFMr7Z2X
D8ETIftum4dt0rLGHkYPIwXgYgMmdGybae03L+UvUs0Zdnj7c7uebKq0F4XkNtx18B7tN7aXNSYJ
jHtFvWqfTwt4/SMCp/6AG/OmO867+xAHLmVmkC3UbvDuQhmZNn9bBfazHn9v6erkCOKwgasSoz5R
y+laHwYCTLT07SICG3lsaFFYrMM2M32FLpalF9/pNgfqWYkACgRCFusmnYojX8swk8rTopQNJ1FN
H4TX8lcFU4I6Fwaj5qlgG/ZYPFN+9155dM1Bset94TdqodYlZ/DYeOyUiOIiEkoOblhlBoxdmXYj
sFN/Difk2u6C6oHw3Mtws/k4kuAwv7gVkE8fD+r4L/9+BA0oaBmR6tjoq6EmDywS7NQDbh6UQvqo
hK2w/4znpKZ1VseVZgE09ce0zS2SjkV03dkLKN6uSbZJxIFS0JdihYy2axGofl75/xgRDTZf1tBR
IlRQar/t+/Zn3JZvuGioRebFfMgWWUZD9mKZcIg+a5Q3d+YRBJlwMMe9OYQnb95jBUgHpimmjxg4
5shLL5yLNcCbASoVa8oYlaFondHrEqE20xoL6+aEh7wdVglivS9VTz/+/0tXWDb7E4THDX8yjSA5
aChba5uLg0OMbskTHDcuGu/cg+AdkOY05d1tq+X+m0T4pCKEnJGo7UnSdhJBBWJM+HlfCgiSLSKm
9NaWLT2vSe8nqI1kqEMMTQ4key8KvaANn/0xyC9uAfJsOtWtqsd+JI8Poz4UuxEXQbpaw5bsX7fe
V+OgTwouymIKEnPWHlssFC3zxWP4krbV0if6VGxkXLZyjMqfM3SxmzIQt2sSE4MZQKk5j4pdFYVm
nZfkxsBCXXGynkdsHZrgSQJmRpFKrNx1gzakikeDxEDEf4jBX36WXW++oiadAO3sGBuR6Hzr1gPy
x7g2mKieADVeDRrawtp34cw7SVhsLXLNy3JtOmCjGg0ULz+ElqfDG4oW8IKdw6Fyp/StGp0dP5QO
96lAAICfVer7oljnIGHhpm3wGggkCZLi6RmHR/whJ+i8cT4uW7KbXgEy5kaAOqTPZjs8Y0x5kvi4
RlOIykpLPG5pRYVsHd8VOcI1QF6dUDNADNqMucLaAtsj5CqJdJ6hQnmT7hAzcjgwyntLZ8SkcIEw
57PPSuRCPZE2mhVGQFwbQiltroZ2YEHxt+PfV3dTOzfYNqJ2Eq5BHyievqcLbJPTy1gypoFgdWvR
IrXHDtwpD+6HbsFdKwMXaSVFvzIzYfMe/t6N90AGd+eabCvBe8lrCgFoNye7ncBo3TzrhYwrlHZT
8WmkxMKqhH2AMQC2rfRn7dqIeio4hegABtaVhoZNu8WP0eydixJ8k0BmmQVN4HOjaqYcJ+J9wriQ
NoY+eSTCNQ/+VNbHX6/ldCMpq06mm6gLay3b4idZMGoPZVCE17F3Hj0xCIVPq96RyQJQcL4BdgHR
WSjZCmXp8ILPvZhVE8LzrrpEVGCqfEvIdhXtDWBMRxQpGqCu9Pwwe6uVCTCbRx96YYmTAvlS45Ro
eXQgPWZBmMSioy5e+wV3bzrelnGW72AqS6hR5EoDx+vLDPByZaCHGPriwmf3D8/4XGKOeeFtAI5E
hgD+Qsohaxp3TsTlqukYf0uG7lEX5pf815EK3V1Zy48Csid9iZmZSKWH6PicDrG6tXlAq4HbiD9L
Bo0Wcvba4LbNwnZMubyxcsiN8QxicFjG8ONjO3/poahxArGJ2+41ruu21V5OpWjsMgtXhVgQ7jBD
vjVPwlyLOqZWvQYbX9j1+2HIE93/9/kXMfAykNnXAUsOALDv00U3Bxvclt9KlPAYTFfUpaTi8mWN
alsHQNrF4pKkTHuhvWuvjZtnSO5CwJrE9MZXMjc0t8mTlt0SIVrhPHC00Zl15WCSwIGMKZUznT1c
IJmFpBWgPzj5ky4NBG5sH4yDmuHZcTLe+gpQwjY+Vp1PJQuurRkdBoJ5QFtCn9q7uZB7iYn6NcVT
V1x3mFSrzLGbInhfm8CzR/G1d3GU+XkpXrt2nIidsokE/ISNHx6s6jl0sbXoH/Evt0CQOuSfOcus
bot7vKvTCcXGiNQbTFidlQfiTWcOIcRgwPmhvDAzrbmyl1QXfRKOYcxOXNYhXxopt+jK8UDyop/a
Im2lWJYAmhra3/f9bHvw3PM84s6a/BA/NCJ4urRzspB4UCxKpV8j/tPqe75/JmYH9tLrkhXUlZmM
wVkMxXhIkzTJ8z2EG0iEPqeKVDa9oj3CHTcXb6CTRZxBTZ94p8SwnpygqqNz7k74Uda7z5l8LUx1
S85uJvQebYsQc/CDhJ4GcihvtYGWv8ZTI9jytF5iy4ibcNgLcJEUCqVTvUIf8+XeJrvcy/W176oD
L33wHvMXKIkGF2XGe/fzB7EvRhWhcQylcQTWsan6Rhw6NdLgdhMZfyVlDzfWys8Dc+/MV28tOIRz
K+vr8J52OoVFc4Fta8QL94yF3uwPY8/4jwn5Xm6qbSdR8g3LXXlp/oXQOXL7eTsij6D6RXDpwyhY
B2SA6UVvkHRnNBNNdHibGpU/o/WCcHcj5DZzDgdjwSC9oj1u/0iuKhR9rQzmT/qIsVxkrdoLt6LW
hE9spr0654oHK522LuHK/ZL61AVotUgwNnak2e+H5ngYcjcsSs0M6yxP+ad8FitBvF8jMr+aE6iw
1RjUb1GR5UQVKOI/61EWxweUfX0SCeW2qPVEKeMIq/Y7bmxYH097q1wU5O+mRHMLZcMUVKWIUe+X
aO2Esj7t8dN1jg39y+XhpF8r+kaPCcfAAjCsPtYdk8SUBBcxzL+1638s7G3W3aHHFZDhVpZpZfXo
/fC/CHW9/vjdh7Rws9fDdan4ARdAr5yLyd0/TPlilZzpbB8SaroBoiQpq2xRl0mXxcWKAUaaR8c9
vT1U9h7OQkJQRwyVK2sfo+1TBLPtUWR4bfKBMIwtULCwskbBS7pyWpueYv0Gu0isMxBzvf9ugy0U
M4Skm4pj5hN3xyHN/wF5IvwXQmdWJOz4HDCzQKZz2fS1xAnWj8agMJhl5AwztjZIkqutfeOrsYCe
5qgQwq2fJwmToLv+mjO15ebDxW1PypcfrsTMNqXs2I1vInqO/yLkySR9FGR3XqeHaHpwZREED9O3
aZ9TN6iV56f2XzacfE6T7/aJA6Y2UuUz+QIzDvZhbK1R5vb+GVfjQgdRu/Qs0GF6WBGQC0GjrVTt
3/aKWwL+6pP1BlpRGf5PdqvEWTDK9AP95wc43iUA6u6ROsrsG94xB+Pc5LIYYW5Ck0PGVfLgAAL0
+RuHk5W7KEurTocR5Ehssp5el1WOA87H2yJGWi+9XO1gBJ+pLukoMh1oFcoEVV0QDvGCd/PxZ0wK
T59xBCMzXZm9ZgpRQL7C36oU41HLqCAzmUhFtNIeAMZgD7QaVV9kycNu5LeLk8Lq24VObHL5mhov
f1H4rYFBOYTLwYbu63YYHf6yAtz1628K1Yhpupq76vYuqMWeWyyx8A8XkVMHD11lX/1okp3p55Wq
31KwmSRGP183AhbeiyOzrxKJxVeWKp8hHWrfJnYP+Xgaq5OhlG6uC8HW53ex43UhoH1FJdUMnJp/
+PJZEemObGv4+Io+hAsnz6zQjvlBmHUrux8y/H7Ztl3oxJD/F95zXEdOC7ayT6PWCqzhHFjcqofA
XFQ8ZOAIbkZj+HLd8bHUKEKaG6MsfNAY7wkfFR/NG6urzZlgYSdEiRj486MS+BGCsAovkJaGcrSQ
CliNxvxi4oPJGwWLjZtxkYuY/NBZxcAOYllSsbu5y69Wqh+p7hjDa0LJ3dtgt8mypsdxIq2NX6xu
55RgzEd0kHggpbLIjaZywxFJA6eL+Mf9nz1BN0fYW3T/Mq1ZZj10dAS5L6dE6TDEwO+Bith6fI5O
TPo6i2+nEOlGhgr7hZN1kclPm+k9qNk/Qysfw/GPl7WWNmdi+fstfYkKnF6AmVE8ObBjKopu4fos
aRxycq52uxwOFrgcEB/NYKUxx4HtrY42SeHQp40Zr4MUBYAAij3Juf2pKEpOcpOuZiBkqg0+zcO9
PcWzws+bXldkbn0MwY7R+8e+cjGbFEmQ83BiAisWfdDpgHM4rLBg0nFBcCN1fdOHV7K3jOhsP8uS
Mabj9Cb9GBOSRL+h5ff2HkigQzTyi5UeLK9OE/xkvAiP7zZn8XjcQ8a37MDpXIwF2GfLxBCkaV8T
GQB4GH2EbxwD7PEbyeVd0j7LtMyvX7H9zy4T7LEhE4s7f/h4xCQiXgp5Uyyz49bqga2qP0TRwACb
Sl5pPWPfJeCg7swYmcTO8B3fT82ZFfXhyDjgjaZULHOLMZVan/rhFOM/b5BT5D1+bQ6AyFI0uPvg
Ew/A/8feKAz9k4nJvyWVOhU3+TRP/MUQqMnmCBZE3Tq1f9B6CIm9U02vybGhAzcyv4tbWi487/LJ
I8fueYbWRP5D5c1ANbb7OUTt01O4rsNwznHD1kytex8UOjSwKeD8jFyTYuGkSvgOeNXI/8otlc9R
4XzN56ZulIX2L7+zzzEguBoHMHrPrTf5p1mSnaGpb7AVuJ7HWwb4sH4+sp50BZSnjcTiJH32tvTX
JHSZ58HOkNCVcfpPiKYc1qrX7UOJfvEKg8YJAbxwVKgtQuW3bxjpuw7iWZ2BzsSuft7hRqEjn1gB
J8p3OoMgUXBUTBXR0URCNGZVhUiEPcBX7ZzfSSkIA3/dRlSCfxUIpD6ZGDXkBV2ddAwRNHuZ9gIY
vzexBwGJ1dBAyikkA3ZWxJXFMF409OJgoJ2uqDoGs6MOZvnizlKrTwEU4Dc4wGFSeYYrRE4K/GaO
xpLMf24eljGyCaBe3/ARZA082T+dwoLJb4USlAWRY+7TlIXbMP/8M2FMm1efC0KyCzDthwFGymB8
qUuHLCaEZfT1+AQ+utvgvFH3lsvOTdlbBoYOzd4AsZDaa0Ft9T4yvZ58hgP04zG6acZIS+MF7m09
IGx+ao53uF6/CAWvUTCs6DuVDJVFk/XWddtozS6hTSADTg3uZcFAoXG+BYF6F8rX8PyQpA6iv1zi
5x1QEDhX1cxVJ+ZW3dG9LuqA0bpDTANRMcT7B6rGc4uqGStJpf7jPD2HYbP82ul+qI/+mktRZcuY
UdelSenKyEwv/Nw/5TrHjWEXYLlD29TOFpJLECH4wmZJNmYG/sPHUW2RXpKmvpqJouqdvL2xrapW
PtSpiIyPZUz2X8I12vYrK/4PjoeH2WkXcYzC+5nh4IkF7Ht8xxk/LnS3PEMB7JM/MunaR3NQkIsQ
So/LMthf0QGT4T8UrF9bmIdrUUqcOW6By7+KmMp5UuzaCxnC9fim5Vmfe3oXXAYQKM/tA1awm6iK
JNX8daUlWJpOe3Ex0ZOXPwkn/pEvXax6bnFcjzQqxZpHxw0wJTC9a7RkSEzYe2yggzLnUJjrKgef
AM86EZSYwfq/+4Cb7Ll9HUQn8v1Z3CvN+EftjqMV4oamX5ZxFmMSB68ngUA0nK98ruuxQE1uB4cO
EA3fDI2u17zAGFAXsAB5j+f25+MCnuXGbTfITQ/kBmRKmGT4pmyEF7NJ/xiSmxw3/rGfg+/RgqPl
Nc2EWB+WXv6rxbNkuLEBX+BPxOWmPi7wM/qDXP0ZrPqGdCAdd0OYiz1L7NI06338fCK8Ba39W78f
js2aYG0liWfO8RCzmPyiDDL3VMfzONs12O5A9XJWnVrQiyCZ+r2IpuffG5LgKTvUjBJ9ENjKvZBM
X4Ym6XD+zCsisCNyEhYqrPcYzYr7L2jti1qqn8yXkMLpz7AcGAKTX7bXcXEWHDsPcrjT7monVC0p
I6M17KFluG8vaRrXAzIcFxE/+XxBmeO6yav1WcUr7IYrXM7wLXVXCIpQxTFjJitvcRlrNLWIUOkL
C7Ss5fniYA8oIaG4L3evveGzI5A959JyFy8CXTp1AMdq9PmOACbhdv48nJSmZVlB6xU7H1vdjyz/
SuRg8voR9/p/HpYtgG64ONMxAgFUuFMsBxOtabhlO3PXupaTA52SfiZ59VAXM/0o2EN+DP7JS/k/
TFQszJ+qbjy6BZc8LpAM7LLdd9j3ZFmKkudqIL6XLy6kFmy+l03vc1zX0L8osce3++pPpFcUWRCe
3F0QQREFJECbBrqAJE/5UDckRAst/HuqnuwOERMofj5IxNqCwJoL95OdM3VeV3Yob5dKtqlgUCKo
dLY3LRm+g16+SIeFR4kuwWXIaYVkKq7Kp8CRvUc78ukrc20/L1gphZmEgk2OBuLe4v7HYzEdTeF/
vjCLUq4VFbrZ7dkWEkc63rK8DaOnjFxt6WKPpXQ7agdQqJt2IPcqBpHmAHEmPU315/CRpzOcN025
qnO+3CTppjyN/XmJrJGvEJWv94ZdQxDUBeA5oIiQ6zlfrBkAdO2dhczz8iRwIZDs5o/Na2ldVS8D
PKjzKBDNC3gB7VaCOfnY2Ka1uyHPqIelEuuU/O0YZtKraMFbeE5b5xqFDFebtoIsRbYaY6cw5/u+
WoRwGqrMl5LoZU3YfoXERDGxl9Bzbr4ezKjhDeciyjOQB6nILK39LGTR1w9NRDs3k15X2EyP8UIx
uZgDALcLtJLSQmaDyn/fk+vidTzKGNvdiXePAceVMFvKhY7btXklPq+ZRWR+fnRPlEgRO0ho6KgQ
l12YPlCmtRo8Ytcjuf8Pe8so7MUizxEmpyKC1tsIy21GJXLIwBnaKBQ4AIz9jMdNCB0ApI4lDJ9z
a7v6YJBX9GF3ADRNa9YQTHdlB5zHJimGge/TN7j5xd5FCzUEiBlWOvo6sUduXw1v3Fx6Z8dH5cbV
6cH5K7q0x1XM1Nou7VlALv3/IoffJ0csTQyuObt8FCOHWg/pntxCnMRNMbUZD/49OgkbDO8LMxvk
G/dy9US/GOQHFupC2dKST5L4ClbrZ/n8PQepzmU5vGgcKFMxxsXiAazfu4ajbHD0OHHBMCj80zZ8
hhyqEflI8f73PXbLtHWQ0Wxe+V6zIKJia5GpYIZU8M0qXLr7/6jRgLNs0ExSQqGKGE8k6XXuT46g
ksCppg7fDDhQpBRdPzTkQUOyQ6ZHIbWiow2GsyoROVSbi6KHheGsk18t9B6BsTyIPWmi0ufMptKL
rD3OOQgZ3SVo2EH7bp8Cx7ojqAUYH7V+i2l8LUOGl2/1sfvkXjlVB/d7jBwZ2XA5qkABkSbkW2jW
4793xCU+yelMUqgXDUQTMX6Jhk/TiUdBEh+3mToSTEVzRqKgYvpyrL6TMz0zJBSWxHOYQtOmsdTq
R/PIgBfimXHqWCtzE7QNEldV545gw8jfna971N0FlDlSgdQKuuYdFSF9JG2RhrIMpydcr2RPWLi8
A+9xLZBqsQTq2WQF0EjKn+EgjrOiEKZNEhj8oKMocLXvIvf8TX910b0dDQP/Pi0dUWOzcgx5n4vi
UUmmB4kdWEkoqjLoLja8L9ppu2q32MqlUi5jp/fWj+F7TxugukQK/jnlR1tOaZ54cQmnqprshQj+
wmZUeqzB7WPWipx/FfU4wmCHiLJFAMM3q6YOj0BciMpA+7YgRpzxcGnLh1cK/cBysYMhMb+isDuS
nBI4g6PhFNOci2WSV83DOwspBDhUyWpDcX8NB78gOAWe3od0VBYnQvIMidQhOINutqw100/MF7Wz
9ikPldPksXNtn8vSl2oj6WDKHHsgc4FWr66H7FCCdedIdbovE45oZoJ/N4oj6CDKVjA2N7NkBf6F
jnjBWsvRLrUiBNDM7dJeFcV0nKnwVrsdaO4uifiSEHtHw6nZ2hwGCTaEnMW4mTrgsX49BE+dceTU
ffs0a0QSamVTKpXGHB3Yo4q3/Ufe+zE+51pedsWhThK2K9fgxAd++EfwRTgkI2vaJMInRIw3HNGX
sqMJ3ISobT7X6slL25Oy8QNsLlJpsE9F9TEIVNiLkpmgi7bGXcLHF1NsEmt48CdUDfoQgbVYYmhM
6NOvFfTwzdU6qVbf9LMnVrfsKSX+QoVEOXAMZFLOumrUcrdCRVilPafD0cruziUUHaur05p5wcEM
BltLydZc9LsGrMWFzfHtapy87Z1JVxUT4HgEHoCwV/zcx4Af1GLzfj/OkAStJfedWSaFV2sxMpq8
zoGMDAzOteWpm8XSZ6VDYYiQRj286xhf18t6O5kLA2A7bEBKtfnpHT6K0y5qho1xJJBpaN0jHATb
4LM4R738dPTkLlYiY2DfuveHVSmNoBu9p5Mdyv7d6B+OtbhnBHOMuRJ88NSX3gElOHKmFn8qMjQ7
rQkp+5wRAbLEMq2uickcFAOOkCKBr9/2HupS7/04K1DboQM8EwsORl2Y6oqVN5ACvjtR/LZSde1g
O6SDTjy0P6hSKFCUvjcFeAb8mSpJakx4sn611Vo2cEn0wfcR/BUXoQ+sJNyJy7i9MH795lPc3qTN
WPJ9A2twLtD4sJh65jzRzrPB9ocDQw7STPIcx99dTKHqMbLnb1Gpfmss6C54IDvqu9cm/5Q8IbQM
yANh3zUSD3tshTvNEg8wLjycplTmgslql8OvJlCPoHMNW69igy4Xt+ySuUQsvgEqxf495CSPStb1
7QIYM3DRHDvz6gzHlfrDKwtLEpSRhrlGRAyL0KGGtlkFfLsIO/j6W6sepJdlFdNt2gp561buKrWj
+0NOP84yeguCvOlioClnxAezzZ5teed6mzRW4T0ZOAPhprfdIgEQeHtqcJLJuHRkAOlbZYdneNFv
ypF0FEu/pmTw+y+LbjZVlwmp63Aue4RtcUGtWvrIf8g/hg97yhKmmBRYU1FXUcyktcuZ8xhaYTh7
iKHOt7dlFtcPz3RNYSK7CEyJOqSn63bpVXyCHCp11VejEFi/N1MASJpcAzL/ZfkXhJGBp2BGPAlE
zuWl8hsK+O9IP/KixnS+hPVfR+YTqxbUuv1ndzFPuPUdz+Ea9QTZ/HFhQI45Dxlen1+71rN5fPV6
HVmp0b/+b3YCLcq02qQhaQTHxUVFTzqxlWNXvMJTGk46BGgk7y17DoxgO97drmzKWKurY2ELNpTE
OZxUo2P+r2cKcg9jPkCDQ6CTycEZ6eUO6KI+BHwDMKvUlP3Qotj4otfOnB8uaJF8PZFQQxKW8t9F
N36m4ZJ+KNNbjUHM6YnK2l6PzmnJ+63NADRU3qyWpV5hHgrg5ihk6q2zQeWAyN42OEmv4GPr8gFA
CMh/2TkF18pui/xe5wQdt0RIMJGQlbka1cZGwD99SVJzJZji4SCoTl6DrWWnRX9CE7Lx0JhFkeE3
qP9UuTmzxcnHujf4LiIspe/i7/abT+eP6kgtVstOWUdCXTxGKUMMH9d3jY0ywniRRm3YJbgjUogN
jwTr1kGrbPQPeNvNxD50b5fKVdjY13Uw8ExBq9hdms2o87ht2xZENkSsW8P7ihKSRI44PASxf1Ay
PJsFVOX7nCqRfLC58hf1Vv++vIs0BZp0OHebA6Zl0TdoUR5GJw0AFl9lGEM8bh/zqL33QALcPNWz
/fRGmBoMHVXvrYGwPwco+eRdLaUj7fxomEHSqHXevuBVW7/pdUcN45xAD2MrmP+5N820kHh+guHq
iy2aSX+I5v2JkaguzaP0bW7145AmOaKw5cEtbwdnsvhCVtNcQstpikNMJbY0hoIkUKq7cS7ni7vv
vWFwufcCtWNxUhzYw5kZ41Wlmgt1s4JKH4YuRzb+8YT1Na8lHzpEToiw3kg5Svg/KiMb7vorMYSA
KG99qbHOgLiqhBU5k1V9DsfTJh16jRsycRaLTCKPIdI0S74B/ljtvCzqlDBCWiGP/oxIowcRFTXU
2FmPo9hj5XSDBsdKpDhf4alnXHD53Z/piGjCXAc37f3qrdHTgw8OEom9J8+WnpNHOBKzS2oMlJpB
fzybtkwxAnFHytPqpZ/uOh7e1K//TKB/3y9+1Uvp5DFlo41NJCBtXMFevc6Z0uxqg4bDkw9oRPnT
kh+5MBy70siXXovYq3gAyrJXVTaOZpcyrZ7uihaO1bTmYYtB7X8iDT0PvzGnMpykG5jgSdve6tD6
agDxwRnQV79sJXrRZ2NZXxeFrUd7PksHVQQ0zfhphzH/CpThtq6UNfh3+hUIw1h3kpCgllOlS/JT
wDYMmp0mhtlkLi5/i+d5ArDUTYBjMtEbWzOyHdusod2NIJaBy/U04dOwvGuT+Ssd5jg9hnbRIt+o
HVtW8LjuZVUbAXl/l7pn1OXi6/4AqCBJv5nCdjKaohJZO73mgd0uAYOy+TVOs/Eyq2ZFmUdheMQR
nHrhP0GLMdxdM5Y0lnPnlf9w3UN769dJmRwR5PMk28hyaQPEwZXhJYr6Rg8X7M3Yv9RSejJ1i+Xu
SvAZZVz4UWzZDknzRv38G1t+qMYGu2jLFuS1zfN5I/IJepv2+FVBE847INFpKFznmB9Yvts3LxCo
qQeTZKeQKOU2D2J84yeZANy1j0kGnxyUsv0Lozm0USq95ulMp3eEs4udPn1qrEJ/gt+HFZHaU/Sr
ZsoyzSoBoYKjoFfj1Y6BkKChZZMIGmptHi5PDn2wVeKyoeH/mG7hKDKkfvkp4RFjxnF4n9Q0WKT2
4XRgZ2eYzL9oiTjdKEw/59FAI0x9aT7m1Rbsn+PpYBCVU//znFpNBchaWb4Lvxj4BA8qcBXclKKE
cyfWn5WTiWHWGDvQHuQpDZlrTZ5/kYZai+gUMt05ejfkTTSgaFhd5E4yQuolHDJ/Gtg690pHFYKq
IhpLZLJYRk2Jxu0CFaxbOC8HbYZkGigPJljpojQ+5Y3feyMuWxsNQyFQhXtKWYsopKnD+zUPvbsR
0RD63ymEXHXwD1WWt2G/KrFJG/OkqXUkkxD/Nwg5xHAY3rL31L3cp347uiWSIqaQsBN4D8slk2qt
ItvvpTM9q39PqNVtOmvq7fkR4sW9YvLQESs8XirkjTcaFz3iS7W0/tYLZGbgILTd/yPnS/5Rl4cO
FQchA0EWgAFr6UHZCjPbBbnMEdQhHbmYJr0T1lvI8g/EdvzdYlf3yaMGJztkmBAIxURa68aJDCUp
1UVtHUg44YVUNp2IYgybXxxuzFTxB4Yn9E6ym6tqmleSU3KN9K/L0o3PuPWcbqbdT1wUsIXK9dUo
Pt7RjHjqEkPNV+W3J3q7Qe90Bpwg/5k2OuQg3sfxUIHe86moPph4Hr20WpG65x9npKEl78G/UCz6
r8E+u8wxMfSDzMr9j1LA+jTEjhChoYSqOhXSMLu5pMht78mPDnSlxTH6pA+M2qdRKD1zM8aPzAE1
lMDrLt9f7Egxps9DhtVgkiFgYLta1YIvg99yTTekmiKNlQJvPDOY51vIZGj1nynKiGOXPA8k1fGS
YTa6turuUtO5H8j9SMaV8WO9CPwIijzmz81FJyNLmUDZAL1eIY94X6andlDlVbGgj4FV2Eta8OAn
e6aRHjPLbQKEtuYuPo9W2fIeXLTX9lP7wd6AYmfXtkLUOCVtmUPuHSbI0GEcZCgtTGK3vUM0gKrI
lW8Vm+uyAUF2uR39bXztGYIcWdK2ZOFSdV6qGvuH7qWlq66UU7Aqc3jvVpDqqBQfd4u2XkGXmaO0
9J+ig+cmNEyVQkZwLrz1Moop9yB4bsko0dld9ZGve1ut5Ihjhk8VP24uexdFuBUCZGGBN40va0h7
CVPDgiz0MXTyOIyidPO7Krz5L3/gbU0FIUIKSayroBpoCIqCqUUb4m6GI6RFamA4uPVFgEqX8Gz1
vuART6NKyXTp4PLK/N8r9GFt8YEt6/ZZBI0S3xZ/Gd6DREnpIJRvAyvSDNo3xfcrBqR1MEXq9yJh
vBgGLORyTghcd8ZJNWOMbxjFncxR8v9O6yIh/PFcaU7clIGghiKYp5wQyqt63ghsk8CfRES1MghU
vb1T8vAqquU542/QgKl9eQy2wbwf7vxSYlZNGiZ345sfIV5o2vUOqbm4UVRR81Na5mdv4MpDQYcF
zLTToFpDBLnFn/gdaBsxhnNauyqLzUDculgf7Q4PZXPA01uncXPngYwi0PJm22neHh8fhQkM7baD
ny9f28pcwwhw2ZrLH/dsAyFftnDjQbb37h9vEK93OpGuZ0w4qnZRnr3nes4jhU17vvz9EO1Xsxkz
6WUXHT1yCBDc/q09XbASpNr/5DJnORp1/6dQUo9Hhdu5zKBaSO18olpyN20mbeWfGKrChq5UUsYi
KzKssh8TM7H0B3NbYJSWFPLC/xVG6L5AIP4zjNKeK49v+cvdZf4JuHkrZ/ebXHIc1igNSmX+RWMw
bOgDAiSV6/vEO4I23olMb88+A5iGzX08vB0qH1Ub4L9Ok+Q+tK/+fYc8Z4nSLNpbc/NY629hSWsf
rKdUilhALwL9OaQv1qWJk5fPboYn9c+Hjw14MUt99TcLxMS3H53MYCENNwBuuaJkeYscEMJkWfGY
xjDpigRtvMeiE86cBda7tmunOH5HqBgEgkkcAK/gX9EBXpB/OQ/0sA+ks+tXiWfnfJEGVeEjMwq7
/oNV62PB0NPeX4M/ehaSwtvadLzkBTSAFLP3eNkZHFO+31TflaRGxWSY8zinROmXx+kVazLwmKBv
zj6s3YDDtBVPz2n5XD8CiAP7IogYE/qScH40I+EHyY8uNMESaVrt0g7EmcG6dO0OHrOqtWJWYu3G
LAUvd9Yu3nL3F3bSlpzmTDKZOpYGEjWyXA8Xd8QD92pYJO+NJV4EL77ZQTKt8Y4/bzrlFshjtpMv
EWSOXArAtbbAOKaDWyKR1gmaZZAz2395wjh/lRpa1hcGcAWjjGunwPKbHHm7HumggZfo2X1J3dih
rdeCNioUl1Lpv5IouYsuDowoLHSHCBI5n+Ka6lzGb+3A87ZaO2A42X1ndKtXqaS6J1e5TZ5Rbryb
L+mgsSGHeELSHBnwBhfUmjTst7l8atNMakZvyj3+A4q1T5gnagvvFrQj1JNxzCSbv3KvHnbTfst7
XpCcBlwebWfj2W2UZ1NbpmycRoeXWtuQoBOxNkDv9sTJWP+ld3zLgD7K2fnGM+W/eLMaD8H/zwOT
wRwEHnj/rP92sd5+oCC4bSDjerrZkNhGxtKNtHgvOkRYGh2niqxBZqjnAIFSPFH/0/ce0Kwpgz6b
3QL5d27G1lD7nKlt7S2GuSa9tDpW97UH27bHdceJzgUiX98hQID0/4xMEhfk49u5D3DWKrVVBr/m
kdjyfzaJtuZ5IqnL8oF/cDKahYvlwds5uFQQ9wsO8FNbXbKYBS8+oxzTIaWLn+2WQxXG6OU7Es8c
GkdAG/uBpm8tkUpio3DCU5vRUIGU4Hy78tAo37p2r7r4xhMKf99YBRWZ5ZpfEe1t7FyzKc+XScz5
5qjUr9UZYsgJTkPtADdW0M0NLawR4zwTPv7EghpLB3XvxO2vworvTo/90TZ6+He3p8HA7DvGISjr
IuCtrKWEJuyAHoyBHtlitZ/YZ7FYl60xh9j4qY0sVOU4ecxSOWKMEeyRkQIPKwGDonDfBY+1KV5S
8r8T2+c35LsNfwYF1ZPKPP1slSS3yVn2GdN9FZxpB6iXOy1t3r04srKzz5MTetEmxKE6vyxD25Wx
YoVCk3btcjNOjONEDR9YU/87mWQOJnUOm/CverX9VT+hG1zcLcaOUA0qdIuRUbwlTqnmdmCA2i5l
ka6RaSFyRP+3dVlEZqjcIg2ow0DiWIAw4dkkrUkXEnPdOZZMLtqYSXnKNjrnYtpJL4d6sdgbClKe
3aY+3LBnmxifCJZb/AZKgWgkzmYaM5vI1FGDneJhynyoCUI2Rirp5rJfw605rSlllkmpkIx93Mgd
dVLQgOQHszMI8iL0tt4/exIhJqMjSgEzVjLwQ0uDiImj0onYRPfssdLj4ont2PQ5e0dkKpJAKgk4
/qC931vB3B/sSa0n43lLe3vOFA8szrbx2KaaOUcr2+Wz9QFUQT1+Zox0LrTGYGI92HGQ/Cai3qcq
5k05tudmy7/ipkAKDs0zQx3ozt2WIB/Rb7otWuO5Ajioi0Ixr1bGB11uhajSNyWO4a0+8FwktOyY
b3Uwden0oavcSItWV0JK9UC2sa2ACG33EVE/lcb2Gwtyl4ciHVGeXaXdMaGPfBS7VFf3HTZF7QbG
1JCrFftXpQ7JDqf7G1RXeISzftXzxnhacmvWK/cihyCCpgHbiU8J70ag4byYm/FoeodTjsIT56/v
+4uHC8vYKxat06+JV/s+2CfqqpiI6Z8KgEzPg+LfFLfPTIIz3K6nG8FwrejK3O1pky0LsZ3nqjgr
K19+6TOCL7PLUtAny1gBzEB2ivQp9fFEe10jQ7brBSh9uJSguzameA7R7uCA8gBT0nCTmM8L+/y8
62S/rq3VlSAYt0uXs6yY7km+sMEgd/0dKjEt4GVaYT5eOxuTJLLj2XxGf0FKjQ/qfeo16DZOLSC+
yvwJaFTKsLuEOjOkBZkR9ox5OUDFDDb+q3X4YlgFugoM3RzrrnWQUxTTAkVnsTc5cYLDQmhdRJH5
SuswFr8oIXrPRXR/WR4zyGn+avfJ2Eh26SOeIiTwhXDlg5Se69dqXlgUHcWmV8+m10uMNT0tOvrc
2CscgbU3dZG1/jFrQesBoSLMXIxU3dLO9PSf5enSxLaOYRm8mMyK4g8kFHoUtN3H3Emyt+ALVyND
50/GLXi51J2IIj2ZVw1vtD9grsIil8rdHTXv300Q+Vyx3u/m6My7F2sGmUbs3FxWctKVQ8ZcrwGD
OgWpeI7/sWEz3WO+VHM1YMZPSngT+z7IWMftXKKNUgCRuK/0OXBu653TQmMEZ5s613w8uSfBgbtB
/HJE7Wg/4tSIHl+ONjtSwB2U3DsNCue1LotkMQ065dwH8e3dT2k7XmJpodCu5nePZjnaLAAJM4ah
FzJv4I2/GYsIdSvhrHzCKh7yC669K8h1jtfq/pOJI+wDIe6qKjokxwn2OnzhM3wjk+7Mv/QH0bIp
6QCtD44Em1u4QzYUUmx3kBe3j5viiHXB6N937S2URGPOTXwtxg/NAOYayQT7XYaR9RDa8T/jqYLP
6VbgK/q6HhB05iw915K9PNBGgCvfAa+CnhhoXlIi9+Szg+e/nTLCD3KwrugvOyHsbLLFyuNLDg7l
lUyhKnju2OSZ8N6zSndLh0AZ9MmqGQLFnk/ns2Gc+4sICckFoSj3TmEFyCQnQb/tGKkP/LWtpT6H
PM9HVNZgm7IUwwrROuv4E+cB3kuBV4lswRjSkRI9AaP1Y0jE8P52KF7khMXTOhP8J1hdIgMBoU/m
e12AvWiMY3JrmscE0sbpuKHNDfa413YIJqoRUjUZRTpSjUwED90ut4HGmsKcvv9L7m229rVvNTFZ
qAWXh2fCvToeKNZHWLWLehqg/nS+LkD15veDcl5uCzB27wxzmJXn1LOK780lLcGn9xF6t0leDA8Y
DCeANREWIUFlg9xq/X4L+JHYNJut3dwhV3c2MahE+Om7MG8CJ9/xXidzPdRiB3KYWYtjshPJxHHd
cr5RYVebcna8HqWpWVY5nA8ciBODPI9wXfpRekhsQGyA9mX4dIxOaMKaAPhSfkGHqccVHOUsxX92
jSBLR9PFuLzaUgGneC2MR2lg3AI7okpbDzvBCJgBxH0l+XVEoXscynQidaQha3yafCxkO/w9qXAD
PdwjK4Xa6ayQ4XOwJ35PDOPWk8SgcWJ+LTmO8C7XY90q7vzC50IVc9Ab8Lh8c+WxP+1Nl4mlorV2
4L/dTC/uS89xQA2li9xRZSnKMug3T9CS12cU6Caw8OI8L65N44oCd/Qrdzh202XornOTucMhAcII
GNYEY9WK7WXjGFxJb/X2JkCGqDJiUEEZiGHal7OqOq8Tag3V5qpILG4V0eSBCuDdEAWoL7Z6/ggm
zOMlEXIK5RLvFwCcxnlQjzwP+Efx8qoYFFYuXkr9fUhaL83rejGrbWB89HV9WTBI7efJpYE6DWSb
vIGk+vLmrTGicq3yhNfthG21xNIej33uvSgWh/CfrHSfJAoC/4Kj58K6OVbW4e7zOJaPml2kOnYo
LehPBYsTAcnK6uNgMHynDATmSQ/Ezn0SCJ9xuIJLtENHpYojqGgfJ2bBpWxZxUSPj2eWibFQ44ZN
y08bXcBRTo2RptWytaSty7EdNh9/Vrw3hSM4W/0nmjxTIwgL1ZHxaGxbiBMmt3jlLUvThklFyq6z
I48y+6vorFsmisPA+U4tDyqzn3PmFWwyQ3UuuxpQKU+Wao+ZjNih1VSn1YMgmPZdiuGCbRiJ5Qn7
yHV3gshZ2VEDhd1pKPQn3HUsdCthxpXDDffi9YL8zlNucfmwNKUAfglaCLxa9HIwfSZvAKSTgWbD
y9ILe5F3uE6LWgNjhUy3wz1qgWwkbOz5bkkKyZWdsaYdbn3ASjMIg5x7rdkCQDgikWUm28ajbofN
gvb6+6GzQ8UP1uBs0MrQRSl9G9lwVqB3Q0aN3QaNDU6MGHiAAGmovy8AwCjLB2T1U4YDNoz8SnMV
+zfh27HSoyLUoVtezAdxUiIYkoDT0LlntCdCULwKsc/kSjJID7LtHNjD3w4XQx+wgHF7LULgsSO6
4R05mtFCNrd3ldKMGWX/LStRod04oo+NVXYjIFYjWUMeA3AHvn9i8E0jTh/hUfqVKGsVUEv8wXw4
oW8nl9mQ4Mjt3cqLqxFl2zD+36e02hJz9wvkO+0uxprZqPOKEKZUcF5GyP4mR8XgjDzRwR0rm7JH
++cCtHDo7r/fPu861lvgj1PsMqixkqhIl4FYmIvz5cj35iXBQsqyOiUDaX7NB9nghMVbzqiHPSj1
vvzwhCFWHYK17mSBEGeiykojWViGBx1gB33KzhZAsrqKiRN2PsvP2kCNudxagFpgKB8t1HoCXkO7
O/wtvrRssxX8ZjAkpHghyZC+uPVPpZMEDqjcVpJSBcDhpbPZzdBEN1o0Pd/3uvggzch8/e+drvOH
L+TtVHFX/F6axoL4Yd0s9LEUVXNNiZhQpPiCaZFUKq+qEp6IQUxkUrPup5GQprxkpiwEsMXMV0h4
dAKRq5ipgTACAX4b2GLnUt5pbGFyZ0capKoCIH8P+KMlbKcQ0v4hRCQLQX1l0w4WxMDM2OaAZvI3
mnXZwQURZXhvU+Vc/2TO7Hi9BtKbpSe5cfxzZPx78Bpg1wvs6/o6YnMuH7ZMqAY70K5UrQEDZ/sC
wCaie6H8X19Up6dtvJQcBCi6fHCQ0i5ncNSjSTV2z+URKn4cjFELEzX90GUu6JlTsrjYSWwucjGM
+WSTf6V895og2YjE+exrbxhFWVRTu04kmrLJ1KJrOt0UdURP6jnaUEASLAVWdd4IuY35YeTVdBT9
+blqXKSjEX4Xx/pVNK3/OVpr9WNZZDQV4bXhlfAHPGbGCI0MthIYc6KWlWx3W0TQYAwXxAOayq06
VhGVqqJ9tqenlB+lbq5D/Be2ZOAGND6aN3HrL8FsmZCxYq68LTR9SOe7eAzICF+fcVyCkjvF4QHy
ixClws3lPmKNEZlJ1zXcPr7AeuUvzDZ9apV5rCbj+FLH6PnrJkXzYsHKqjYy7yHmUEl9EpJwC27H
Kg2cgC1zq76UYikoZqQ/JE5ueEqCKJORtYATD1GDFRIY23E7Jcjyn5xiSNv0KkdgnpD3TbLsTxsi
PmDBPbKfaDIQ3m16z/oTInwTcizudZWdxBZkdGpCQGJnz9XQ4wVuHiLFeC4iMvJogzqEEtrM+6qM
hVhkRI8o37hd+dytmzLXhzHf5EJTUACGjNil834snxyInbQyFEHPxT+0eBmU4rCgb7smToysfkpk
DKfdu638L6CnuOJMjTVqPfeEOVZhj7F+K68PoCaTeLrZqdBehaP0NTA2khG4Zhxf4bxf8rJNumzY
Ldd7AQzCTrFBna2OzeG809OZvYTi3N7apyI3HtCXfKQQVlIQUWJyeKqydCVwp6yXpuOXZ4EBETDp
aRogmDMe3XnUmpA2SNeoeHIyNfhUYpHpws79ucTvgGqSFzGcaqQbThOUjd//spPpP6PDB/qwANog
TtO0QnUTBYaC7H41vmbI1+X/l/nbdOFEaxNKniXIL4J5H3D4qAjzo2xIagHcJKmhTozsFzKkas1z
NFyLs47K14do/SpXb3eS85pFHqzLU957Q3C0mhrIY0zKU3lUmyMJIkAugQJsHmG6TLZ1D3qodPYt
lIP2cPl8p2QkbU+g2aEBLhr1BlOw1mZBgKn5cH0xWO5OFSH5geXtlC/sDeTye5vCr/85ACG5m8KY
ux2xgBFlX8wwHAHx97jygTqg5qIOztvi63E2CScNbPapLDfu4w+9Av6cKmsxOIGnzWaRDP95cXMt
R4OK+vEA9pGQsyfWVFBBHDzxXbVM0izIzzD+qcXzf1kYInmG943w/03IhQ/m3y1wMhAZ9skXYfu/
jqVn4l1co9U+yfPlLMvPLwHcasCe3glmbHdFgBdugPUJhUy1/MPI2TJuiwu2Wai5fX/ZHenAa+fY
YhGjwRs61PBbwIly0CvCMf8xMbh2byPZoQJkZN/HmC3rkljh6s0F5J1cYBdRxYRqhg3Ooz7yN9yK
RysLt5sIEqlyAuVJ2elxsylIfAS+tEv9//ZWjeaoob+Fsyx5cG0SpS5zHz0LdLWKh0EFNenR2E2F
YCr4cOp07Ao+QiFDjlwQmf4EyCDMgWoW/PUIzfhpw+b3+xOCSuMrAbKxgoMN2YKL/jq9pzlgudxc
YgRkmiaSPxRmCG2huCPzSj58LAhsFw+MPd9cg6s1s+65qw8Mvs8VfqX+h2t2KKwfgkKlHazAn5jw
bOg+eICq5li8BpvfVIPITXD1zGcTH5A+OMzmAfYIvG87Q1WD8pvtTyTuZDATRI3wNTdDM1uIeIAj
Xx/31hOGavoMjL+9rCsZDOnBbgmgeWFTG/G2jIHwjB5jWfqU6r7A9OYaBpgDt05EzjLuREvx6c3g
4sQb8KWJ0W02Kn8QTup7Py7cHZL5luU1BLvgzsjK+o2nItY8Nd8ItSgw0aPxHV+auWO+TZvRb0pC
Ft+ELX9mgHQv1dDTmwLNTlEvhmTKTguBznbPphMIAMucGyv0tYAw5jAY2lFNPKWArVvCP4M4TovA
Aa5QFQ/NiMAdZ74/SkfmPOn2AShknttDnxnwwhAggXynuVJj2uUR5uS6V+yRsjccATbC82ilVlRF
LeFKC8wvamJPYtKcNSeE2zK+Ynncyof2gq6W46rdy8dKa9WAZ6iDp3ylp49P/Ok9YLwBNYSZphKw
ri7At18A2VzgLDK238WIivckN5x3F/2x3y+Dds75d2k9XeFoXpZ+sMl21YtpT92zB9YSDRpnR7kB
Utat5UxqjNSWkmb1RrZFquapRtWb4XRQmmAIjfuRSfWcAK38OmIyXTj5vT5b9qUiBCYNRFlw3do/
2kui+fXE6oUYAWkWTWJIGgBtP7n67OUVGfFXvsEbX/On0NSjJIMbXQ6duHUrfjcXGPgd3mHVsxC8
W6hgjI+I54aYvr3jP+CIGhim7UI98TqLE5C87IQUoupnm6ELOkv+ibK73A4DcU6bnWO0WaDWqDBP
3FlNSTQNgaRjAzBorNOKvWiDYTEW49chdimOUxQkPlPP0jnRHNkjVPXWG8nOZ38w1i9fsFIoEojk
xoIE1XEoOIT7Pj+v9O9eXZPWLN/iCabVXsJ50Lvf3Sn1w95PpUeRlHVA1POXnLcXM8gV10FmPH4s
yD1lsrRmFaRY6L9LFyiacMlL+wuz1lU0i+o5e6HnsGs8f1tQ6924z9L+Aqlu3eE6/GHfSTvKR85P
sUGvM706YJFwia+Q6tgRgP0fuAdmmHi1mwHWE/neXff2nloThPDI5hhfkBTqqxg9e3iXm4XLOWjX
CW5qOj9xSIlnoZTYVOjNbFY8rNnhfo5vQmr3oa1YNqsNl7KggkKhyvlKYtVCwCHzBIL9nSckp1zF
qXALpZlJqi69qak8tS3IQOnNrLJoUKi+a2QyQCp5TggyPxoWA562NtchtYYNs+/gmHEZur/XFdIc
0YJCKrxZ3KwfO6kFOK6+Od5FiCjlns59Oz6DU7D0UHQWNepl1Tefe53avS6IrLPhJGIEbWPpX3SN
OB3Jooo5DHZLrHrVG+13FoKDY4/1/aChCj9wiNfIZ2BxsjUiAuTH/MNj8qjCQFEEw47Zw6yr4DSZ
32pFRZPEuUW7eSetFXG+7NFhtMeORsVWB3QEzRic2WuUyWfy85P8Z9aI0+fWDhaVWBY7K0Yjhdqq
8Oap7MC7CMNTtF93vvHFlBUOkDcM5dhQDlTf6eBB+HFiSmub8RLDGgVMEwJkp3Mm68Hj9IxrBzwD
X7YVC/hV8SZO1+qm5bdqobESqE6MrnXikvzd4uTOnU8qJUN+Lr6632skmrkCbZHMXjt68kegyT3F
8vWROpvLwuOXLHeRcbHdgHGXP6SICXkTGMvLcumz7pWfAxXpchqQC2HC3pRwxU/ukUs5fvdhQfqe
YKqi4aEHaAiiWV+3g1FiCX6WKqCcnWXZtIlMtNkuYf+AqyklCqW+AE7WIixNP6dHqBySnlpvBQu8
RWDvYYv8Q0S2esyhECTV7VyJEeZVmLnJHPt4wRKYHw7Bw1Iq+ApmAyjbe3HEk+1A4VoQwLHrLswL
7mVZHj4OUdPUrtPcyP+EmAGVsoOrlYM0asMpMQwuZLR/sXft7i2ugK2ZcSx8TAFEoA19MB7rqk1O
6KNjn4AieB50al85Au/bbcu8dCl72kASjrD/43H4vsMwBWZTlCfmBuSXIToD9g5ImPTn5mf50zrW
TBJlK1MTMxLxQFFKFVgOZKXRRs9MrWMToeJjbwyJz5rRjrUfpjypG7WhiOtj/kWHg7LGDOuNl5/T
D1gxjgC5b1GVfd8fOBfjJfMH/aMtc9fx/eTxzza8ZFNn9S+k+nb0Q+43sSYj47GISP2hiOE5exy+
aWcXQ3JVPQc5IEJ82UeiRPcX/phqUPqmkxqq4VuTWIkXZHeq+kR4uLF4iya3qUmCjYimS4gdWt9P
kKcnMnVPqBkfsu5a+LFcMyN4OIfBpE5vgaVStK0FreUQ5uYqrJClpDyTd+rdWPM2yp5IEp8CqmxS
7P2CQVouDSjLA2hIjkb5pXOunMpJhEkz6BIrMjoDWTB8jrISjnPmobhBis66MRIop4w32pleX2sY
I5iCVi887lcXmuNS9PvivHEfEnzciW733faFKPv9ayYMM3GgBfDC6mFNpOpHPhJCHIII7SO7vgBF
bwID0zpjRUvpetcezIEQLIHcF+g8x04oRtQ95JGDhi3/FxERyOLPnKApvVgAdWYFUOg2iPc8q8Em
WHDp6ps0Urh1ubKV3FnLcr5ZOYdJxhCfHjlN3dJfi77oYYquiNj5ZovZNdeT7JsIlt68xrtCQM2g
ob+2gr2lBniNPGHefHqapvAoflWcMMhVOleTsnhc20ohqy7M1j2h9wQUePcATillYskEGj3co9jf
9hhVFfHA9RWY/u/VqJEpGKiFDRyzjjad5Wr4rg6GEnZhMpmirDEl61BI7lObKuKElLFgaUjw2JvX
+zIp7lG3hzPhYt8MHu7IGbcEUJpoSLMXGzSdTUm4GarTQIRfhZft/sesmsvMbcXNj2fydGHwHt0L
2WWTDJniaUue2uYhRWJ+5o5Ch148N9BBnk2v0TXaQ4F6uEhG4LU2acvORAlyo5/Kbks6726bb+sg
E5jxQ1dW3lE4A0Dp3llT0mZVuMt99MAaIxKvM1NXdYS28BXgJzffIev+Mf8qdStxaYHoZKMjWzhQ
SXh+MU5cRNqgLM0mlBWtD8lDG4Ji7VzshPO1pe61R8FH6Iz1P2miNJB2U+HYbtVUfehFc9fDMi3R
NL9XxQ4SlNcP1qBbT7rVZSORJYs4D5K6UcAC3eJZU0ZLdYt51mpFxBEKX9tAI8puY264Lrn56EOV
edFUn5JpD+FVwlAlQ63SRlaIgX1Zt2ahVejlTaImKEV4S8FVd4xD4TdtNM/CawTqOrEwKsfV+Z1d
2CvYelQlGRFcgp9ANUR4koYXuiKIrAKKxBl+wvldJ3EvwPJlv0hB1b7oooguXbxVAH1znlmKTkHa
uaIIU8TG1YS8iErVIQ1jIiLHd/VVeftMOrN7dSfIbkt3m4UxLNnwtm6myKy6NThoq0bWy2ZA34QI
mFSS8+4eazWr2kdcNgu04KC70FdoSDw/pYuZCc+oajtOCitn00ANMpNTgF9KD5/WS73brqF71XQT
ZCz86/vb00pJVBj1ZYgQsYWk8Zc/Pfs/hTpYaelM5c26lJnmuDrEeotwgt6Mqrmorx2PKMnoH0Ja
UAHYHUL1ubT2d8ZKq0YceLrxxadOi5ohXQmVvJMLsGzo2zBH+298LWWE4FKtG1am1Ym0ZI/pBMj8
3hr3lN58YLK/H6+5YQkBqqxecWuRSiJj/TO1oPRwFFzNfVDK0rUMzGBxuRlWGO+l3el3QVE006z/
g/2Zdc16SwpH8qpZbRzguN+TvibosM7OcW3OULFXd9MjcIlxV6q/wP5b+jABW4xct2GCSzVZLUNg
rI6qtJQA1Xh1kwBwMQPIUV5cKGBwIkjbKYXdiIOafvul2/zPiJaUVJpb1PQtRb5EWRe8OnKMJzTf
O2L95ixcfa8wu1apRWjyFtD7LW6I7rB8wEBY5+Iq5S0GZ5vQpPjdbbgIuUT/9ReHvrGSjcEI+ZG2
L96RhONPtrCd/1x/Cic+J3QEcS1pe6LnQv4sTvMnB0VgFeO0/Ungr0bLoDyUKi1nU7ybtZ0zSDA2
fQ0EwWu4edsb8gcXkHgj2OnA+l5eFCjIywbiU9aQr0VHmS5qlletIA0yT0gz/T+sjBsZWmQxd+Xt
YXpGM/r6bsrFOhH/8GC76NgPUJCSJ5tnYTua2arCui+8IOnZwxcpkEDljZd3sm+Ticp0+9Y1iEdo
usOBxKUrwCZtjnqQFjyWiR3cF/wLHDX6ecVtjIPELVWJU1VfdIBu8QVfhx77LRq5d0dSxURsQ2Qx
ZtS5nU13b3ZpqpHnH3uSro+dIRu9WczRhZwfofTIguervy/851AMH3yvdaa3luXQQn14m7XzEBAV
Ig6aiiZM9+/YmiuQE0BQlysVLPcdoKrhKBuB+KiR+Bv4A/mZC41nnSh1v6KyzTPGEyvrXBimGCy1
bXQ/NLR+I7z0pqwKMzEFyso7fYB6mxiJ+CGmaH7GnucQmpzcDRoFa9y6AbGHm0ifiEAVl70LTkWR
911A3LKVCAVzJIUuGM7sN+8Vv093NBK3u9aGQJcOiG3f46l71GnIql+asp9y0FqrSLnEQ0HjCYGl
TysJWvfBxyPKqCmuZdmfO7PPZ6cpxjrxgEr4KZzBf0mYeriThO7FEPsW/kXxtl4yZhEjmJpGHO1D
wchcLxYorUTQv0wqqX39v99z5/gpmTWy4GSETvO/GjUpg/U1qNNbWH/CU+OLaELwsDezzrqblGH8
0Sg6F0M5yOGUZNzwPlfUj61JPDPXTJUYLB07+qFqOBcaEEYtC60baDcOWhTrJ59VrsEDllymb/cF
5JuGtZnNQGYSSdfdtBKKMn7WXPlYiUKNaVnRVl9kYA8VY/HZYwhRSW8fEwUkxSFLsm4Ewg+TUjdx
4MmHGdyeTmuc7a0C0b9ZRYFClS6Hkt0HtMcnTihXGm/vNKPcEHbbbMIlMgh4VK3ayl4lJyNW7onq
3DyWVbsS6NB1uZPJPtQsge3NPyQSONFbV9tzZMWmypTu67j8ZTzyR59DyEKPIc5vz5UFUuTkxoO0
1mMTRVC7bpZHIj8aAih/b0yKLHoPaHPIymNINqjFDKiWmnrwe4RSg8Ga2tDistKSmd5BH+xD7qde
xzkKPpA/cw3fVaDjkspHnWdHTaM4i9SIE31OtQW+/I5p2V/OYVXMWNXlOtOQktjWd2LeosSptauW
E8fvlnWWnAEAfz+Vk1TDk3Z8B5PSpEgIPhHzo69wZB6rr/fOWvPPrmV+qaPyLwuY5PhI9KTixq0s
OJxHPXxwQmH5L3BkSRdVYuRhP96G7+260bPYVoGs/mxpA2EKJ8iOivA+IkUM1+gvfv4xsKwGyBHF
RHI3tEQWMaR3T8HGwS+BtlfDE3SWQ7j6L014u1frGaQwbf6NivlkYnoM1K8dJDYb787EPq+72k9E
yyL6FCimH6gZoZrffRY+1X2SitctJal/dgcr7XfMCdPZWLKU8eoXFK4VlOMqPDgmHU54vzlr2nZ1
M20DTVf5SNOFDABcylYzy33vaDbuPHyhE1Ml4hXJiP3YKC6sfy79d5FlW+sex6+/7vWFFdtUcQ0l
WDCGZY8MNEOFPyN3dUdPkqUAhXSpWVSBL8KIHGT1puged4lgFwo6op1DmX21J8XwiVXPVkzm2nLe
8PhfkJkmjWgSrusRkj8pj87a9Z/bDWJJR5IAh8JEAheU52573imV++RMT8E4UKx6WhBT82IAFNYH
LWYuigkqGDHIACzg4pCJBwrnJA0IXR+e8VNFHZ8pc1xd/Y4JWiU+6TvFg0iOZoyxZHazMFsuI75g
Si+dPzaoFwU/0ufUUx9jV3sPayPzaaRJCUhEfWJelGsglLLCvMblU3WHwOwjZpsVf03xKodcWaIg
Eo/g3CkdgVpwd2OmxJS5zSsZLdA/nCF8nFGoxH0DK07YW3GXypUg9pahnvNo8fbMOdkDxFdYnf7Q
31ZgRnNxC1uEzCKayVPXNaz7mMop2JpZLxZP7AyQDKK0nzweOJxjGC8RahdLTRY6UluRYA9K5LJj
kIMCAfJVwSrJOP30q5BX5IlLNMrw09sIyRjUWB82+4dHPTEDicvUF4SZE8kMBshaAjgnc+7Xp5px
AMrBA4kle0zZQWB2dLWYOrVsCIC0gwhYCsvEhcVFylMaYU866CRXAlLzrsb9AXIYR/bNhYeqctuV
E5RF+t6PQNIMnF3XN8T9ZuuGD0Th3tu1lcS3eY0988SisphKgpb2epzNZCw1yclc9GKbKWLm15aV
Nj48RMG2BsclkEYA+QVA5diOYwWdcZ4Oxu01lWebRwWtOOxfCl1Vd5QE8tgsCr+yisPFF33FrF1F
EWBGDs1Vpi5NKbmhQDToEOAZkifeXVwpUv8SocFa+a4Jx8JfIcUCFNwHZZ4aaLdosy69rlUpg3hb
iRg2N4Ky6ZQ1eyuzcm/OFsU5EZc7dzAjzrMn+zE2DvPbOjsVsFvFq8I31uIuzi89ZzyeyrNByg0r
JK1XfBfxiuMC97P21dpJRtHJTrzlnqMwhac2s2nvey9deArc/vmm70kFknoZQDvrhvTF5f8ENbMf
Hmnaz7/xICoqIWSMKfw5jpXGyR+ys4a/JGKudwXNQXOKMOALEObqp8cgKz9TTmVmI0/U4V+uUMPW
xRVXdb84SpiirD9oIJ5aFMoee74P1jEY/fSA4tMWNzGieZgkgM32Qsu3NeLuPcWpd6OQPcyLMlrD
s1PqU9YShoG0nlYBj0kAJHTTYOtFAp3qILtKl4+jXVZl7EGseuyeX1nzI3VmST9zG/77A4YqOgvo
r5AsV3crku3ShPllm2QhpBh3WdcoE0Qniee56MEey5jChjXyg9hcMTAFNNVOo5GJAZW0pDQ9SQ3K
2LVMWZ3kxJaqfmK2tcvQpUNlniQumQt8yC+hCjisRf8STi31Hr0rGw9dOp6Tx5t5I8q0UEHs/GCk
d4KPMOvAUGp/Seh8LuVwfEjdXqbaMpUEoAmrnTqUN4bdGguh0zvyxPiUqZO8QxY5sv9FBFy6Pf+/
LzsS272LC8tq8CZkO7N3z79CEojXC9cjvSEWTSRz2Oic5Zc1+s3NgB+hs7kP/Bkr/89jFXTFh0Tm
F8be8qNNKXo0n6R2g3XdADOQPLKd/pI1COayJGdhvRh40zE3iGq5gxo0oCrxWoPJ4mpae85q3VZB
w3hMoSgl4mUfAna/10zfmjscmOOAvW6xYWexwz7kddHJwKBiqd6s+PIzKkD1k8d+B1P8bkETT9nt
r1pKvgZN+MDL0lSMqO6xlH3nO9IEa+MhlLu4fwL7we5HsojuqnlQWkBvrGu10quSF1Z3ajRQNYWx
iiGz8hqyBnZKyNNra1aFKQ4tEvoIBR6IctcYtdR7E25+ad4YiVvxF2E1ny2lco29AC9mxyy2aQzq
Ln7exGm54VmODATipVLauOKGvYInvhZnGzM9V9joG52rYugx8c6aDBiTdE+a8DHgI0Qc/Ly4RObY
eYrMuE551rVcTkWnCpVegknIDn8l3+uCc8RxKqHnyhWxlK+k9Q/QSbfrIMAeXbXAiWo79BKAKoK3
MPjpVyj7gFdez7qoudF/XSOA5QCSnhvKen3AHMBIL1GC09m8ITC8l/FOCJSI6hLYfb4FY4OMT7tw
P50NnX2mh84Yh+Ad3bmNQLB1gv5RjoIX1tk7rQmxBegrYaUiW6MWRQByJ459QIEKQHqnYcYCZD1Q
hbiC8qePOCKDxyDbtm5w5Si7Hu34rBVFsO1QDsShTURhJ38Fgm12LBridpqk92xZmCU/LTt0yqXf
JGRjTh1ajxDdDr2zJ2By1WhxPrN+yBDZ2eeJ+ftoI+gEaK8mCIc6C/XX1gU1ex6kLa2DpEig1+cE
0LFXXNgtd7eqicspSuRZnrXxlcHaow2z0BKYDQPNaZrXI4mHoQ62aRAlIujUVEbxRP6PJj1Aclkn
mf1wwDItfearoXqTsSgyBSp8BEIlGHEeXKE+pZOxtSAVdbknoWhpszDzTQnFZ/Bjm3v/D6v04lzz
UigML/UyrPJBKKzuK4f36gMnRVrLY8JQSYkCIZHKGuIHTu9oRQPH6BaKT7Mrv7LjWKS+8cO0W3cI
DSJhIxoRGIYP5Pm/+8IbkhJB9O19oSAl9wVITYN1cDu0jU8+QhEX9vpSoF2PtNqz7EPxR44M/EE7
Ljvj7K6KMy3Lq2V6+nt+V90PR9QYp8TPcOO65XgJ0B3a7SXG4CfRoSUZchDh7PuPZb8aMN0khjSP
SFx9IO7Nnj2Ncg27bRvmjc0nfkyHoVC3U2Np69z7h/CbPlXA1CKiJ5HzCd2OnHeZgmomHq9IEBOd
A5Ibgtxwlo6n056lUIz96d1Q6xIs0KcjIXxB39Q0NSuhOgAqnW+KtpkfHVLqZbkM0c7JwEKtyiBX
pA5QctfIy8ggv1wV9F1ZVxZqXYJiwTPYGHLhFffFDVmO5Sc0LO5yiAcVWrY+txBCYpYNJuJ/qXvL
MDP9yzGS0vGn5rM8Q8H2kc+/s9yCAwje7BvF1zJAZ1Ll1bj/386ujt1wUFPmoBEkT1Ap0fADsiPz
RFlSzPEj/v17POE0JTVoS6mGkYRYLnmeog3yiMA3d+tHMoJ0tadjyl0fiyxayspFMSDDqo/yEi7l
s4LsrrLiLS6yNUzyMw0586dKCPysrlGQagmWeDPRuj7GnWPVr/wvp8af1C8lfeU0xZebdymK3O5V
8Dw7VidNTWfb3GFkzWQeNqG7EQsQkwhHe+zsXoEy2q22QqxBvF3ID2AczCWHYcIDzPKp/oLcbS0d
jYBo0KrkYlCDnIl7IJk99MUiZj/BCNLmYpO1f3GG/DKFsjSI1PQ7Li+WPe0glWRg8J4o7FBm8XSY
ktHN6dy65lF+3zKjogFZBZ8RfaQgXgvEq5mI4lZQA7sKlrblK+S9+HsU5w9YxL29xQLuXVgyeiMg
P3mUBjzzwY8Log1D3/Icr5VG1ho7L73cKF/y1RCpcF9J5s8ceGsJN+agl6SQqeUIeJCQXfWquf/c
2Tf65TzDpcAaejgT/dqZR8aO+t7PTwNSmcFSOqeXRnbaKUD+ousIsQbX/p2CtpN/UrBvm002Y6Jb
InXM+nLtWCg7OO4WfyTvhMf7sAoViufcf6zAQ46zZeQr9FUXYpkyrzy1j3GtaC4a1IpO2vks6QTs
fA01CXpuuAbSwrrBN9n508Xo4rRmgiepqkxLzGXQIPZhwJ1OtBuWDLKWRZt1euqil4zVSMSM6qiy
JpaDn7LTUVvSO01D1EmKYTs5xGESwcHq3eBQYYHbSDUF8NXsXKOBzBp6rL9Ruuq9Xv8TT0w5PPmL
NCJxVHGCvsROj+2g8x7mdxBUXNEcACw8yfXyrW3tgRNemtGz9c0oFUYQZaNSJS4aj6UcU+7fT1Q0
qhHs6ddzzyk7bE80R2QyIwbCLWCO++0/jBzMsKEHbbcjURQ6vR3xftRSVf/Zb1ei8Y5Q2C1pEPFi
iGB5a2XQfyhs7z/6bhmenX5gG1TnePdxipuRQM1VW/d+g/SKl+Psq1xz2vVFti9bSutL46Vi6kTm
yguO/5uhor3YX2TfWhemEEMpbJUo9u5A/lNmiK3zVsvLyXUDEJNw3VmlMwM6h8tZ819ryjniJDCb
/jsMbP5vtIGKegq68OXPiJHVD+TObNaGhVYYZyEylZ4cKXslj/pRIFTqENlbhSlrkuxxpZnwo+WN
h3+QBh5fNSqWJjtEdrc2gx7aEJ3gx3GZ7s/O2scyPKU/8qQNzBcJbyWFt5uMwWcwM4HpgY0SevMt
/Ove/A3ToxRwdINYmH4HV6KOkpxuOo9k0WVlMnHwjUD4IZrpciMkY60RTkmaVTAISGtYIg3zGCnS
7PKmqGtcUPs21eBszf71epAh+i3o+L8JWZ9tAiLhm/frps0V23K7ZjIAy5FXHcWmmMWhz04pdjSE
BrUSA2ZeBNQwJE2fn+JzxkxbloZdMeQHIfZhuhogW8oEAVszImQe2ZwhVukDerfPVEzhEB48b134
49X7VtjNqeWOSe9t10w68LVdKKRSrdYJk6IU7IQSZCw3UH9kKgcOwUpVxhHkDk257c5fQqWBQpbD
3YitMGvcRzId8yWXRl1hKU/zDJbVwic6QrsDYAE/wfXTYPG+N4alUT5uONQaHXV5DOl4Nnkh+rSG
ngN4gkBkajKnQDz5bZYsfGFKid20LfbA/nrBHzt6YwMIVQYpD5vVcnnZO+3L9scPe0w92SAAdHUd
7wgcbLBYXR+evBir5S7U0mCxQCcLNU0y+ltlaQyrVAi0SPKrsYKptRlHa/pZG5/wAFYJ3sBl/F7e
o0q5/q+vJSy33O8ss7aBwbUkl8rfr4EBCh/IqcLjKWapYkaTz6GZtJQ5ZGL+FKf0TnCh9lsh+ojz
rIhK65SlBHDoPKjbeG6doR3eejpknt/ZpRIOV2+rM4/5mjAcZRoRbFFiQD7lYvgpcZWWexZ8e7WV
WLCSwBHhVTXrG13xrVOFfKPp0Z8+6kVbbS9p2Va9B1zotdCJEgaxyMUFXqUkpJEt4nSuDufWqzeM
6wXBsso6MnboSVU6z4VdgEnD8FlMJtRSYzm1vr9NolTEJhzhhpnynosaNqcskqFwxkYMYNwP0vt+
U/B+301Agi8ikkffobh5C98Y/mcG5LrUr/SwERgQNmsXBd4f1Lm0d25Y7McR0Hc3MzFjXjkLKhdV
6QTOhFxIZd6/KcN7jr7l6o9HavCCj9rhjJfLjZ0Q3unFfpdokBfND0RJyaHBkhMkDQO/2S+AWpos
WUxCgGcYvYfvQR9bdk1FE75Oud/Y2+fwX9BumlCwmdJ9JDLw8NQgVFpf0oMouI98hr2QUyrQ40TS
UGXZeXlC0WyCQXDYBAaIkvXT3H0ofvRCKWaRrPcuqoRvKGd5PW5i7UX0ekoPRgF2vhMWIZl+wblM
1BKJ0i7Pql4MKEASxdiY0xXfmPzPHrII2ARsd/G4+C9X0ENphYdYnjqRmZAHXuhZtEjlu1zSRTd1
u+TOjmlo7AsO62XsaPFlcJVuhonNbGX++IlGtkETsQAPZTODYdODRDnY78u61yAhIT8RmKT2oj6Y
bPTyVjaD6QKFg38ZI3bFEGJqLDdI8MxMBTEIZTtdpInQDeUrHWXtoL/ygrbv5bUv3qUBgPPkkSmJ
egbRBLLCO0I+oFOyndpXy16/XYoNmskIiNPs4UHylbbBeeE7gJe7VDzkufhb5+8OAtVYUzJizISQ
SEnnDgIIOR2zyS/mTMXRA3kz9aC/3pL6p1rYTDrr6QOcyJsWd7zBsC8mGCz1x0kSZdJbl2cPMOkm
rP6tMWuK8rwtv/Sg+NpAJZyShbZfLbg3orjVMZEgjSqtQofSVp3/Sfs4pmhqBBy8LmwnjQD9egMV
i9WUJ1a3Oag4bzpOw/g4MdrJXsxUxFABFQElOQOzzWM8AIObkPdzH2t8yRNS1V/fZsXG8bhZQLsS
ivwwHC+lsx2TP5CAqXawp1gcFmw4dRLdDg0+QsNdvbBgRVnFjNmredBulB70TbTagzgWNutSns/O
/hoqRWUwyq1/L6GrydoZ4pf7RjziiG//bykXJiZoC8SvAd7F6Xrs9yLNSXyFOcCXojU30ONn89ax
cdroW0dj7BmoM1NzzOjcdoFomRKtwIha+V7xNB6MGf2rqHY++QC90B/rSGMmdV24lvH3ipcIbDLJ
B08kWY+tAl46UIerEeDvnkws70GstQdZIWnSTbkdRIeLVGbwv1l1KptbFfRXVHqc95MwXynBcKeW
1vMDGL79kJbZOKRHfKzNcogVrcW6ovibOgZgjIE/50P9b4bfWSQjoWcGu/zD2x7YtbwD6KTRhx6a
vxFP1ks4e338JVX4VpdO2v1nEw/ZIOzWuGsE+LcopeUclsES1v4X1ET3lcgpgAoTtIGkqXOrjJZO
PN1tZE9UkXPoxI6t/zCoASb5VQxv+MOEeHF6NT9Bp1xF6p66wv5sT7AI9iDn6hLJI3SWBm2oh98d
1wfD0if6dAih0W1heTGunWO8mJ/Yf5uP+bswQdfXJz6HKj/bRmLNkUsLxpIm7ULrdCDlN1yJOMuz
aX0ZhSGBeCbRAf17yaUXClMyLiovnqMRX2y4EVLbtMTfZWsBysUF4z2tu14P5wDpxD2y0X6VfmZl
yZUG2L31RHTxtaXD2HRl1h6+TDGZNWViq3MUFFKJO26GVr0mpV4CLWrGjkIdrbtvkZMMoeeRbion
RnONySX0s3OU2/WJohuAGfUjckONAKg0VmHNc0UtUcZXxwARENYNCOf0lplfqr3CfAMD2zSHxUom
wHHBkOIh4qiIkZi9FtEhdbyCyMubre/YvF67skO80I6imEYKzumRV1KSjy3yQrovCCg4UjAC4du/
22QTeieGQjKU4cjcU3pht9zwDEF7CFWzhcxHV1quRNXJUxXOr1m0mFb/xLr4iEYuhj96G2OBRMMt
2HFLK1y1YIj9ip8hzlWOuNZE7XFdxtqbFw0XkEBmPdPTTZlpmjA/0HIKBM8/+DouaGkB7/83t134
H5qhAa9WCb5OUk3u2VgoUtHv5Xe3TaqM9CGyiFGp8Dc0UrLFuOI7vVNfk5Gp879h9RCaZ8mEOkoK
3Gp6siLhR9HYTa0k/qqphLVT9KTn3fcbTCDcbbuU8PVaC5YnqdlWkAv4ZQUJVv5HXxUd8WahLJaX
qmtWL9f4PAcKHNBFiIRlDZamufDi0my4G5Zj/+UTX0hXlEFG5gbe12tyio/gx8BUBFMypjPGEnIs
d91PkqOB8NqHYw73nno4LxrydIFgIjb00mlLp7cT3V4JwN0v6BeuFdNLzf9S323zHnnyBwHoTVqn
EbCCD8qkEggC7d1mu52xf2GFle+JAakV/SQJVLuNmEpqEh2ab5AN0M+2bZNf84GAMfiSzHbNbpvA
qpll/NTPg8Mhp2GuphSBkOBCZTVLpXcc2ttpanj5kyyfyvD46R3IwO+HYT3MVGZc7tc+I90WUp4Z
uaFC1/79ThpFTSwuwkMVSSC8gpBBazStnBZLJDU4cgaZBQYJfbYQsuXiw8U7ILBlvjVNQHUyLefK
xEA7HaJQhCeJ2ML3Gsf6qqdtKQc8dkWtyUhSAsILRNcwN/jl59LYsv1lfDtkKdIFFBcjLNnUxhx7
C0T+KSB7ebv6TtA7EM1idW9Ga6V0PrGBtnyBgfnyXBOYPh0X9niUgGw/avMnSb5hSbaRJwugz1uU
2QulLgvK7RAUZAJxnf4lRQ76cHxfjebHfa2RaLpjDlgjIgYmZZOU/DJsthATUxoYypS56sEgNrxI
8fZafw8PCB6vsW/3KW1a/yboQc3aW0Ip3Hh+tTCvS0GvdwoR+5ywun8CTrHN6WWng3uhk8BNQFJG
fGlIHFYMDCrYCSsPVSUrquFZD5SNBRUGWwGgjMs0e2Er2Nkw/KG+VSjnYhgjK0HxCHbdgiYmyl+C
gGlH928BeijntT0Hqc0ieolAp3cZECU9/J6zBFy/+6SqNOH7AQaxXatHywHmxFuQYe0e7eYmJvKm
0gjpL8dfWZwmi+kVjjyme1mwdIB05y+GVtGp0mXPN3tY8IP1mGaSk+goCmq+t2rmCrWw2O/PJAyl
Loqo463lxJKp5nFidpmDh2egyRKILCTPyMZCevxAwuET5CD0ppONUewDa6ZNczXaFd4oxrH5yCey
sec2E38+0UrPA+TXkoCbjD0OFagZJ8Lri1o41v6l3ti1Daa0RHzAJLylJxeAsJEl2Cx9EinHLdvd
TR0FY1/CWJMXmjDEqAKVnSmRagnnOJFbmNOTkWxvOmYdWbwHuh1Je9VvaanmcEfQAQDXaQvJL+Sf
7AgmsjdKbEoLT4WQ2TjNIWisw7btHpi9L/6g3AYhsJRBIAw56eDej+JVUyhMgANvCUnFLcqRt3aD
PoeLyaG22s6ZwtQ9cnwmvXA9BvXIhxN2GXuxkNr9y6Xz4/3AwQr0SaxPz6s9nMMGbYSx9hPZovOF
OsTqXafy5xsM1uA188hWjglgDz3g06JIILAGgIHgmllCMZ/LC50rW7TU5IjqLt8SPgB/8Ajf3/7A
aU+0cLKINebVTZVoOCqWv4A+nI7uO6+JWiquTAprszmBeDuQXZuDSHpPy4ZBFL9xmfqeCF7UUaDu
p2nGkf9qwjQ4r2TCsjSrt5z6f3n3goi8jy+XCCNawvQ8NlSVzsKodx7++yxr5xvAD7t51eNxHX+p
/8clD9BKDtgT5ENXkYMAeL08zS8FzB6GHnCrjHTYoWilPsv/D2tLoPCSNA7dAGYcC8JuPMO6FlZk
QJinY4NDxj9ll8lLJPxIi5fMrWugrH7swYMzyXcTwNMyndMoE+pjrQHQhgmw+PQluGyo6mlWG3du
Jla0imF7CdOGFiskDz8Z3xhieYj2APaT07R/mfXTO0Wq8TlrkWMig4pzg9bk+35UAzQWjqsmMfUr
GmSCzzbkcSzvKKPo3gs2jwFyn4BolyR5Vtozzv3ivEjoA4rMBUlM4Oo+uko9RV0SoY77xcngjUjK
JXNL039mYaaXBkhFVmbgTBZ+MoldxNQ1YwId6qoKSU+uFqjmk0JKMM/1zz1dJpKsz0N1Cy1CWR12
7kfAsCRTWCl1ITTOfRgf7mdHkjgOMIoO24qY14LsvbfWOAGBvuDPlrs1cYzct6r/KjF6EcrQ2iEg
WqFg5d0sv55IDUUN0ksRt8jR+0LmCyryd4tkK/35ejg7wQYLhY5zRBl9CpoT3jT3rFzIJ0JaIxq5
ZoLbn9lPqD3TdKFbhqdIzARYtLI/GysTT8A9ArK5M3mhszyHN9+obcUlO55EVUtVwBpNOtJ4G1nf
OmL2VzpGQzwYHaDk8l/NN2t0Wuxzi/ExJDJ8vOp4pgNFUXT4Vu7QRGloaYY0WiNrC4rdtr17Bj+l
TQSUJ/QICDUQsJcjs0WLEM4sft4ud4QpLh2H/eDP/kROO4nISdYN3dXpjD8Se5EC4+9i5ciSUJ2q
s6EfSLkC0KK0sSE88FizbtPnEDr9/lLbNf8S5zrXzCizOF7WI5hazul/NqfcZ/qKHI8y0mkLIZnw
5Al2FO84jSkrFpCuBJemSDmUfduSSpNCZAlBm1kudDLWI0W4IeNcUYVixyuxJcgAffV1LcE8aL7J
p4MK1RiGhWbUQQURtF0Z6PA8n50twpK+I1ZTdpM7SQryT7I6cPci9VXh3kdiR9h+EVQQs86qQVnx
8dF+MYBSzpHUWD4m3v6/Wnl6e0EVFi6RZd65oszkjQnSwVCWGldVcBBR3eBf4qrJE2ajPT16wq0F
QMBB4F55wAwlOaywdWhrbch7mVi3AuJeEL3SIPcSAkmyetvHcU1R0XIZw0DeflmuapPAn0A5GTKp
FM61Ra0PY00SSZpOX47e5jzmi0rdxjO9e/pIAl5Ehdk/cWKQnShc5PbHXopB6tpqHxJvOCrkrFXz
4BtKeYiYwHACkil1wQZOy4XxY+xxr3TWNzsnGmvc/kvaStjxjxrghiSqldYLm/6xldOG03tI94jO
8JnLlCOq01tz8PMOmsAzc3J0HGXUcq8evuxkZNwi8Cp69GC8j8sdbYyK0RekjnOEBzj+/o6auecb
0ZURPpECU4Thtuk3MGX3WcKp22bL5T3PRJskLeMfUZKWWMI4hNQFl4o2/fP6d+fIbdkVlXk80oYj
jlideWHw+reqyxOt7oB/uasFYPJDAiIZ4W+naYRAJg8EbLJPS5lZd5Qcn37JPRn8r8s5xPlnVFeq
ZcJVreTmXR1eKKO+nalx6etsv4lnSJoQT2QviqbPjJv/aPMqnDKbuJGU78MSicp8O1dHgDtVNC28
qqOnbBEl7mlsfW4VvPiD0cOj3RrgjniFdwIgLSficZTzWWwPGtL8QC2D25jHOKtUvZSAYFbI0qfF
eXWbpFFxozL1w98LRoHnFHpoFtJb/TIhliwxIa4cXPnEx9pGjE1XIikvxZei/fLtrG0CIdODtjUk
93ennwMZEt6CBJaDFkK/4BtFsrsPtC/AmBtMvi2OZ2W3s1gaZYFgA+X+dfj+JaTIsBFYm/RGApQw
uqnkWxTbsuoJQCHXgGMx07ngRTluQds9qZ5FjmoZXDbQtH+2ix7TGy38Vv5+NW7MtUUvYg9ACuoi
EVMtr4nyx6U+QaR2AJkBf+f2RoGzh8AKYjG3BeZJGqPty9fgu50rlcvntnqFhfhLSe1vfraaWlGM
ftKrG/gn9Zw01wneTFe7XwRd9iTDS/8xAcP59pbEDG6R2XTBKN0pqyJb/ePyf9uGUcBMllK/w7Va
8V5D26Ey+ggA45onFa/lrCWtWVrpkSvfDFs2h1igfbvjeUWfijrF3aBqunfL7bwpntgDUPqxwMMR
hnrZ4rKtm2Q4KS6RmKpdyAtyXASrQXgmFG/C4G/ljBsRAYek3IRTgJ7YmdMb1i25DFyzpIS+tYfw
s2cH28F2mqtJHBoVZUhQnGYxZORm7/L7gy6sQf22xV92CJ0oSOfIjzVXCJjbvi/u/UPp2bS2h22c
LJ+jtJTIFLuLdOgUv8xIIk9SAYQpXO/SmOJlXyEvgd5EMecUjrQEWpkGTszIrkjA2OuXRCxZ0j1J
isBAE8XxumANL0m7b1Ht6Nnzo2IX5Z4+p3d8ws5e+GWidM3hhlxmxkH6s1nt/dHsfSh3iwu2kXM9
hpspdXYIazWrrBegCyOnYF16G3icwIIjwE0iDDzQwXeoxDG/gy8tEawORTPllN3T9rql8QJjadGu
0nm2KT5MmPvKCDpyyalFERiB/0Xy3AQndoQvpTptZlmpWEfOqUIT17oYps2nP/8O2wyyRVwlmOhp
j4hiE26uTT+GvKoNtRb5quCymOWFk5Bx1FO6/w84dD1w6j0XUwzwDKBlSuDWpw0eLCspRvvu1roD
n2rfsG0sdB2yBLQfNFwnTuOK11d7/PrGbu9uJAwczcVdq9Drs65g5dUoWCNi9MOm9CdMzPW736MK
UfJPv87cbo8kMMDXBbaDzNWjEWeWj+m87Cw3X8kzB6keBnrVUPOVLiMdQidAXVkmmtRWgJ1laPuX
nF/53czpTRENBg/uET1qNdGqIiUOPeLcx+quR069AqNK8jKD/g+O8PrtZUF7aregFIq92hikzu5p
PJbNumjq4E+P70YaKytVh9kno74bx9+GmefwJxqkiL2WAkNiB/I5A4ttVw8VEed4bU27bFQ5um/G
jmPpELwzVwYNhmRESRyvfXZg5h4ZIEYyTZ7NdhCMHammGl40YYqYsR15eM6SmsuWfdV0/DUNUlDT
KcmNItWmMmlmazsC+m28du0d8cjnvW0/zpBZyUV7kwNDyEluTzj5Peym0srvKQ0ToruhI8CMndOx
EPiAe8KP3cs7ibzmaONBy8j/SFoUJuN2TXcjC9QlWLHMQtMQBUdqAlT+sotzt2iHmgXPUiMgtm6T
87PygnNaCjbHRTiwlGVMFZ639HngbM3AabYWfS9jZ2CFbyUBG/0QBE2/oB1/VXoAa6u0YxprT8cE
dU2bKg7hnbWvlySW1BZbTzstpqQrOq1QsWGcHcf58B29h4cQugrsntK5OCKoWNeKaMJ7oe0ROYJv
jx2bm77j5O2fs1E69hIyZVwMo2T/QF8Wsim1MnF5v9z8o4bx+lYP3gC0sZf9p5SW8gEfb+h82LVx
AAGXmLv+Vuzhh1l17pQahVxQJp/hu40cT7qJNO6NCY7TypMdOVJfpvL+31GDsc4Rs1+VGR6hXeia
HLSpjjs7DeodG0ruTGmaIM6BmdiREdkgU0IhvryKcKSe7L5q15wdzAqLz+6iOi52DzjZ6a+Xt/1D
yv83bRcCCTo7jknhunolru/y4/CbjOLUNrkFeKEU+oOa36gQdX+dNsonO3/Ib9l5oRX9S7TUIL+Q
xq6oDwl3soHtoMiPuhxOzb8ISqgPzP6WGcEfCfMO75vr4Gz8KTU4lNLZnpQkNWi8AD9+8Adx9g93
tVmLSc8UjDnaf5/lUH3+zg9p6lDX+qkrioehjWh/HcbGpErq311UWZVBx8bPsiiRp+gbdv7Zcl8R
Zhj+pJrvYqBlnv14znNdiYXJsFLiRFg7+i1ARC7jwsR4hvS0qS4oMw/43CIT1B/fjO05T+IyitS0
rwjQqAHOwRX+hcB0bmWLtGDjUCmVj6/k6R79h3+9zpsbT0R8YlnN/XjfJWR2zApjoU8+O+E46Mo/
hAx9aoYBuelHu6UswluUSNeeVt4ZwHSSI+8KneRk38S+cvRRUADVhztOPb9lT1rUMUh+i9yLtEFc
dtmvtglB58s+DZ6bys4yG8sU/UiwXXLkRi8ev1ZzpUa9M67NcfrXrInAkREyeYiA9rJHkrjwpxvt
3WFDJz9r48Hfx56c+uIP1QyOTDC9yTMmPOxq+5q0sYFgaQe4v64z4if/kRKgSs21h+1piLe8QG6N
rf8/aVt8+Zo9zWA2JLuiosUJQ4OCQffKJoc2pV56mNkDm70fMBOK57w+7TH+doQ5bja1JlTVUbRv
ZheTOxCqpKj+qQY7o6mhmJ3Upk7aLpNe21sBHeYH6PfLehZKaLBmJvANABrY5cI/KlYf1r5j3X23
n/u1bhWbkojmZaMSlOulA1LkmvtpxORuZCNPtWVamEcCkKIuLPGG0ez3iFHCmp+ECMNk74vNr4yo
CygUHZpkzwFZJJf3z9M8AK5DlcAKbdU9zbxyyOuIbWPjLONtztlZpJlHzG3luJr8tWtKz5sLLMo+
NOK3i0uZPzy4x1oKgto4XLH942CBMWyBwwUEteAT38C61MNuSkcfBvuq5piYNon6e6e7zYYGj7yG
JbF6BZv27w9nT2tnuA9rlsLmrFK49V3O3PRqp9P9h3m9WxPBNitEN/vEl1RNtJogKqD8XS/EGEZY
CgrjZm/JHca+To+hBly5vvVccttRT45PLEWQ7a4Nyt8+2qrzgAa1xt5mrmkTXkyzh5LMVwSxMHKb
hlzhO3pxkyez3yVpamobWC69XsSpLRQJJF/6fIldJAdu+p3IxpmX4mf46q7sqmbHEyK6Ka2rmBsp
B5AFb0gPz8m+wNLjSyduMn0kKoSJbeAXKHdtvTdBm2Ug2tvQtYYUtFGyiPUyagGKcJM4nooCvWaW
i4YHRRfVg9ZLP1NzDDat4d7a7O4Fcz9J54IHerOcfMKn8BSXbx+gWeFpSSDWwZ1bo73PrQv1WVlp
LJ+cTXTCnxuwTwdoRGu6FmdpH59s39Dx2QdyAF3o4ZJLjbMCP9tSzw7ZIDJxqdIYfcjrYElsCIzO
VL+OhOGGSozzvKxhwuagkhIIYzSBQwLonvmCnnb3HtP/Rrj0X8WnSyv7kSUfCi8ayXd5IrhQaiq7
kQS6rN7vMhMPA2d9L/qPv+0r0P2os0fCMTuQkNcco18qYSWo8r1DW1Px/Bi5Isp+RH0D+hVE5f4d
wul3ccXB4Ryj/elut1U06GQv0ZMcYWkPDNVilRLpJzcRag6chflA88LuxCI+Xn/EL+88Ejp5X5Sx
Tt55r0LTRGVFQ7s/uI9DeJGlo6JdThIBziYycOtMOuUrh0IYF5GshKw2y3X4Gkal4UPhqnxdfZAU
uIgqSJt7zMHyGNSiPaIDef2nqC72l4rv4qacs22EtlKAA5ofKC+HTEu784JTDF0I2eFBid6rOrDi
FdMei3qMEQxHKgcOYyaOWLz4k7F+Z15m3NkIbczMlrnqFLNBZrNBgN+oA+tNU0L8CpPc5IwipiXE
1CRo5PHFd35Y8GeQOm19AhvJ8fYA2HcCyvPmnmNFluZjun/ctgHtp8hXYxtNUeQH4k5p+mGuosYb
PetkffErr7+ANDlxCBSY4lRhaILjr5Klt5dkll04Gn/qBebCaoKnbMme6dCAN01oE1SiOkiOzMU8
F7UNFJ0DZl+lrlCRq+Z2yhcZB4RDNzszp1Um4DwVKxxtoYXO3XK5AvW3l7R64iHhhc7hy0YntR+4
+/veS/gTYl84deJcVQEACgfOKadXFGeiqhFCKchvxJQ7lC5nZaVGprk4aClcmmtrjQNkgm7A/9Ta
xWbfoKMOfJUhw1ytenKB343mVZBIJvdxkrFZ3lNYFaoLiUx9w/5EsRZbG6r1WmuivEj4XzU9bTPO
Phh+PtMs2lOurDYeGnjVWDwx2fo+wKgzLBPQV/+06GRaoi8L1SPj0+OXCveQqNv80vPnP+tclg9s
BKK298hBCGz2CCFiRBP/2J+1W+uexmYlay3TWgfoGt49ZLu5GHfcnT8gvS1Q0G6U6/oKGQqNG2zW
ZjtR4aiAvHWVl7cxMCCZ6imI9mjDvZl2Os4+ng2Acn8gZR/pU/VtUjCCLahGC6i3jUc0hZqyJOyg
qf3jH14iMS34B/flXbKVkV/F7he2JZ4Y/d/uonrJqvLrCOVlja0FpAWn2PwmYVQG6cqGEGwkMGfx
gUwQI7/7mInmzDMPMUJqRQ337IqIgVXBLl2DCIZ9VWVCMT8AHPNStpBslsySaMUVDE/ueiEvKpVV
indh/kWPJPvEBWo+4lWrKF5nriKIrEs/D5HzYQ6eCwE4UTMblSMq2uUOJvwSNdSF5ZohZbej4l/R
sCj65yiKVy1Ykt4EzeIn7OBfbwj+wprlLvZQ+p1Jzf7TgosrGuRr/qaiZkrz96eC9PyW+++tY3P2
xjkM86EhM5EuU9koVK9VRXFSvlx8TlVFAaS1qtn8t6Qtjuo3PHZW3CIAwvcsGc/YW/P0GJBmbDZY
fvO34kaPQ1hUasfuURnEZ2oA/fIzDdeDE9Vi2QvAwJ9xdhNhzy3X92Xqjiq9CZFKPBzTkO4nSvet
OarSviTFYwwtOw4ugIaI1av6du2uZEVzZQM10zxBSy+JcI+qqMksXh/g3FcdAAmsIQph0kYqhbni
CrmhsHk1tRnRMRix0+mLDESwO8H+Fac+lQqNmRErFh7/zwqKiEosSVt56WychxILr49hk8BMER8H
PGNiGmvmfHFsEvqpzdBEDYgr+knRpTc7yen7XCoJ1EoM6iLNLkstMiZXM97um5qrJCuXTSY14uLn
6V9ychSeBDmGnY0+lcApktGDM8tuOrQ9Xwg6bfAcjkhxISX/iptER5e/jRZ4IQD1QvgoAHdLD4fO
3kM5PJaqwBFskyna0aK5h8LQPoaN4LD7aB6S87WIAGDBxqYp/Kz/pYsoaqQFpbsJk3iAdZQlMXWi
i7H2AtraXRBtPXIp9FkufYRQqmfvFwcCc64hZ5Ku9bYVRodT0o+5Ep8erdcq8fDhuktIf7QVsF0n
3/8eeWo61MjfVVzgws94dcd3HCP7JNRHwFGd/xcsDDJsMp3MQfyZUzr1s8XNpf5BN+KN7gxA/BfO
uAKk9eDVVlKF4FmN/acrugEbxkY8jQV5LMYSvSnpEBYkjYcpekXhRpwh3AAJB4KuYpzhCLNGIfe2
ph+JrNR/kqcB5syl6EIZLJSbuhOkXLs3I+4gFtBIauPShAeLYUQgotAK+oOOpgHFsJ20EXx/vUA8
h1u+c4u2osmOgMGlPTI+7mznbsngrdBT1gS+VCqu3g7afytVPxkFohNRFJ7HQj2GT1+y8NuKj6Fq
qKFXI1QxLZDbs408pZOnL/vkP1B2CtvydkdotZL7uawsrNjj4Hwy/Czp21lkPmH4sMNEDEo0ZQot
Bkyv4Lgx9zc9EQUHjLsuei+5dUCO5Uetyea0IwporaB6vnz9o4+3o2Ti2B2jmj1GwCFq46EHbSXj
80667/OQ7nzPtlKou5Jz5BqtcVeiIwKSaIrGAxsJFtgxEWXXpXH60GkkfvqGAUpaXgymA43P4XJT
b7I6kMki7KVkxFLvpqAXI0wgo/wsH4r4SrLsMUHYh4wguOPWPgottXezAwDCY4oVpzoiiyQUU0yi
HotyPCWJpElCUv1Qi1ry3cEfdgm7L833kWrZy/B4bpSXMKB/P++kwQdDJqrBpubEq80mBvyyUZTm
BpGJmDO2dGjPdeJZucxdhOJxO3Ui99GtdezcRSEUzzGlfpJ/PYLVxgjoBABrWpl9M1UosiLcGVkA
dB6ZVt5CuiUy7aSj/ST1xpvYXzuZvKTqt1ZZUW3EzDcZXYee7sNuc9Mv+gIj/lXjYa60V22ZTZIG
mHvFFMIO8lAUzF44UBTJ/OG3aQbMZO3NC+EseLCabZdtiZXVN/7Jv2oKcTa/PfRLGEa6+XzdXhwU
6cILlosMUVE/1TZgDQ7VNqmZzuTmiYd6bpD2ZfS1VMNwgRaZS5MfrzviKHQEpRum1SJzZR57iTzf
2Mdv9+4MEx5gp5FqyOoClurs8aCE6gPruNKfgschj74EBCLhRhQU31Ro72F8Fgf09riSxViMgCUa
17a27YOhCj664bmTsyQTcVWtSNd1gpF8NJQ97B/rWlFach6grBNGQI8LewBFlS3HEmvMI/T1wIDy
UijS7kyP/yw9e+5r6EFFOKajH4N8t/nNBpn5S8kmqxqPde0HRSZ92lcfFbSz+t8KB3LHoFr9xJI+
O/xCq374E4PBM5VyHDfOJ94pqnd16Q5u3JgABUnm6EedvpKGLz5JM0PRxiAs0MZehuEwVWAxsRYY
CKQjyuAOM8xaQFoCA7ka1h+tbjIY4iupGSfEMx+843+J5xmXxuK4cVgTosz0GzWR3MgamTKUyJ38
z2tCqPH+UAWWlvTabkwLYrKsxLznzmIfzaUCxVX3KOsItIa4GyGjVoKAszSWmupFJU2clkU2aSzJ
rXaOwLRWAvhbVCYX5/c2DQCOFBTfp1d4zxRirQ5lWZ7Peh5n9+UZJ/DJATVWcttz/AzLX1KC58AT
9IqeMF6k1+iEq5fU934x2MQa3X3qlg29Sk2QhJk7U7hC8q8gWxrdXyk+6kdyuA753Ywa3rxGZbwZ
HKMRSUeQkLtR5grJy7yayflEoDsYI7Di9541bRZB+3gGL4n1Cb/DvF4p4F+bFSWJ36Xqzhdkbk/M
237YnkPOpEVoBKup7LbynnQbTZYbxGAHIq/boBOVYnD/GiRb/DAjQR2DDwE2mGb9vRU9Zcn84mDY
vSP1Pn++4PXkX8GUCNAtGg2sfdrECn3XhSYzHI0PO4NN+ugxcym0nMf6MDDPsM1PiRdzyPbHgc3o
B++1T7xAZAfJbN72Ad+9UCz6XbtoWMcAyIVqamYUK6yWPOgS5z70Yp980jUJtYELxR64rDem3+e8
w6cOrJlP9XChjr//COERydiNBr7i+4f7NEihtlKc5LoeBQo/O5V2te+PGKSe3kDgMlDdylyz4MvV
4aHW9yL4iKNecjWum57eM/NU07j0PyYBnTN0oMV3fmyTku0rFewohp0uYwj1SyL1SDB9P6GRDXvO
N92MlcImgu4+IdXrfxVJEUj9sQPVT4uD9vzKkoZkJStdQVeX+BuV6Xr+peGMWiJNwPJbb75hFolP
NWMatHg6lVmkXh8AhV1ZmPaIpJx7u6dBN4JmkJRVfRYWjYUMXcN/7s0N4tvOroP/3mmEVp59Angn
Dr7bngjLF48UU8Kaqy5Z52wpy95WSfkGbDa5Zzu8S5QZmTHmgwXUIGXQJTlJY7SO4iDLr/x89HfL
KB4wVEcTuU78LTlY7ME4CNPzJlLG+FTRC7LPjzkZRbVmbb3bBtBvs7c37vli3uMxKjrkYSajIU+r
2FfrlcEZzsypgiC37EDtzoA9QA8ZIlebNHeG6BQ0Vgz1VKEuH0Lz5p9TaEzRKG4WOLRiMtXBf7G3
1fFGKlUDboK1LX/jCPK3JdPPGpkrXqx+OWKaIJqCqY/6WH5d8akRYq9K/NEc0qUlGC2UihvMyD4n
MaV5m+zbvCHCUdYO9xsOnVO3tPuOZxls2pO+CY02VtepY2LaYYFbBs0dygeQwBLV4wQNAgAV650k
ugQOmd57oSZy35tJg1lxCeB+5RoGYzdxr2M0dL6TqCSS7ghtCeAusL1/KhriUbbI6xVtiJYcb+RI
XlJHM2hsOB4RiLqmt+MgKnIlOonLfx/BmLrXcyAv3Az3OQAyw5fg9OVb3Yh5Gu9N/b451fBeb6Ky
JRBwBS5exZ2RJED/iwkWxVYATPWLniSvSgqX25891E8fRlAS4h4scZfsSrf5hAJ+xUIbibpVphtq
QK3JO7UDQg6HcnHXxRPdsov5TpMWDuRoK+UKdjryQ9wOsKz/k7o1lyYNYVueJv1jB0s6yZv8TIMz
px72ekvut58nguJIwz8+9sH5JtGjK3U/osLGq5aovHAY3Yf0ZjxTZpDC0i0wum/WOoSWt3CJ/g+x
zlQ8CG9wloiuXff7oDiHyaI3hbkHUpyhrnwY/3pxty9aATxfqCULJg0n0+WJVk61ZEQUczgB4mAo
hMfGRApK8tegbucxn20idBZ9EXsF2U0DPspg0jbFpceZUhGGWEewtY+dEE/3nQfK6C+lpiLgf0PO
Fjb0lUJcXn8IeLvNx3QHKZuV2oLiNxsVrECA/GOu2eJUn08aPnAeLKRYfj43C+YHQe/vLnfFAJCA
p0A3qea05rkKljxgTyNQi57nEiRHxmcKfaf9sM00ywgjH2sqyF537X2MP2mZuSixGklh2CU+nAlm
lMRRW7/kVBgNqlHoatnevNXop/RONYTxpuZ+4IvRlX9K8f8HuSoKjavCnEtEuKsHSEgvPfT6CToW
qmjc+35y0wqTAm1q+TLWcBdUt83OSrRU62c5oSZx5KoWlIZ5zgw7CUDASxEnyZfEaEw9hPw+qqNC
ikqxUGo+Ll0ksPMUbt1meCKHQXDO4eDi9jUFGJqwq6wixo5AZ8CVumuM6Qoi4clLyH0NwSoNAno6
RBnpZV0nO1fkDsOqAVyf6lEuHY5uZpVMjnnZvdCcWJ/HG8gBw2uKfM9WoT5/5GNXW1n2PL8iCAPt
oDKRDgmmCGPm4QKD1OTxmuTk06oRe9Gm1cfOiJHs8TpYwaUwR0pphbj9ygTEwH+Xd6EWw7DIgPuq
gUtKoavkDbeuByMdeUsIdXIFLrKqNR1V0+M29z+a0iTjAA9SFyX/osIORMoFYVIIwITqoZ6HsRjL
vLLetIw9e0Q7TwustakRn/Kq62FZah39t5VlYpjMUA5Eu4nq8LL4hrfhOgPWbFekIiWLD4/TgQ+w
6xjchjifIZWG8aW/RkUG2sRLGird1lOTMf+EZN4p4LKnWxEx/FPEVR3pnfcjBm/8qJcGV+MvnEi5
r5zta4o/J/Tic0Qg6wZaGR1mqUJOEqE7nonKHj/zOheAayLuiDv9t51vKdREP+EjLCo6SXntkhbJ
RbAdOrZDeTAOQVsM8GQolDuTgeEmy7gFg6KyHyfJa4mma2gDXDRkcokPB714EwopIWr8C/FbNcLC
r1YNhYGlpynzhQi8b3ZyPMRBY04HzrVntjbi0/nHD87N4KSgZsp71JzwM5q/X6LOFZ8bqVLprrec
l+BOyt5dgZdcbL/9Dd59UWR955AjMlb65y9dMhB4vq8NITRpy9x3hq3LFhpyQxBVsZYt+F5FSDTk
X/KXb0EV4k/GL7hV7gSaJh3cp5WybUXT9j0dwa8F7fJ3jIG+5OvSFnB0okI1f/33SMypmznVWniL
xVph+6VvxYVOFPzK7SyoksrgbVt9DK9IiaA0tVEDFZHVU04WtFqYcSzZJ5r/yV2542SfLZ2hCcC3
0F3jEDSuwRBi2qrNsPSSDRLudUuvgwmDY+F3l746P3NQeUfJ4n7/hRMG4JRomvofhYOQhH0pFEv3
t9zTDXY+ZnY5E0gDD5+NxC2KHRzX8+iwBzJX4T8iRxqw1e+YNu7Dj27yDpyHxXroi3dW9QZI3Zp5
ubtdW9qt5A1jTy7cmSXuHcA5lWw59OOcxfmNCIrQvBG6t769eb3Nyyo3SUCVghGqi5buIazMaWWi
GbiL0HsGsOJ1fz0rz7CNNOmTUCAdTjIE9Pclw/kCdbBmR9ogE4nTcj40oa6nIUmb4q+VxnCQ+ppf
+UNYl16bePLaXiZxPc72gsmb2/AdulnO4gphw5T8rsBWKoiQmUgWX44DCycaSof43tWf5Bqii1F+
XYzcMWtnaXtwLS78sh/AV19+KnHfA+XxGeXpNO6lQQYBDlIEC0+bA8Y5IKGHt5+U5khJlr4sS4sd
mjGXU36MsrSjOiO5+oA6qV1MW1rJDRyoIdy0anrQ7L5xNJZDatU7MIRi4y+p+t3iqT+oPOojClM6
2EOA2HeDEzpuNSGGZKpC64SAo3n7xfA2XamQjCNtxThNzjc1NLLJBIVu/vUnt+JSKPlruy2wyfkD
trkRkuMh2Dm8/WX6C0kxcTIqoMCH2a0lSQL/7plzXMsR5jgKpLgR0A0JjxFUcr7LfHMcPz/fIkBN
AqJ0zLJ8yVtBquYnZ1NBwmz4cGJuD01BzMBL7WLtA5ep5xaMi/b75TaqG836anwQ1WwD5oQCYfZ9
QI56CJ8SsCYkvnnUYTtbvcw3uysuVBX4rXtqYlyLN/QPxSAyJ9anuaN6ifWKZhqmieZTT8Ilp2re
VYe9QltUNM9WHw9mpe1mDGY2NUEJmLZvlcN3iM5vBKc7CyInM6dYO7blVwH65/DzPJU0ednY4ZZk
Ym473u53cjGlDBqH07JrhjjqGxk/eliv523KZh7Vq3exFhYBx6jtYoRnOZ9lw1Wx6R4KF37P7ocv
oTHNKIkXyjr7Sv6U77QwvooSa7mpAcl8JTxbbNzKFfqC7ebiynsCGARd7BjBqN0ulPYJa9gIi9g/
L/28qXZkZW8NdkcpKwMtSR6Vcpwwk+aiyir966Ub4IG7TmvsLCpi6PN3ySv7znrwkSGqPhrHBQyG
xGjjlnlAx92rODVjHQUvCzlEAkR8+EknjU3IPOax7Cc2RggKavM6ISSH/REQK/vuTmRGqWUCvEP6
EzSYJThO8NTvdXRzK1vkrknFKOHzvJoOb3dCFtKUxK59/XZcDTPx/NBAyWWuW6ccGBg/tz9Hb4J6
iIi+GSlQKfugWDC7ebo2YIDA5gYdRxvMVdaeQXAhLgv5MNTY6JNdiRfwgcTAceSsSNpIqi/uGwTw
wm3viQ9V3ho0bUerh/3IVTSjY/RItNX66bNkgWm5GjZxIATPS5WTWU1tJ8FwzdFrGBZEfwTb2/so
PeVaAeUKo8Zsei8CA4g+lAC4P3km3La5lMv30WRJ+X1NXn3PJM0+ifvi8texEe295SUM6FkJWd27
JzkInwh/9s4kZBQzcDADfvuVrQtVkltlYuWXy7oGseGxdU0YGNSYktphYI7XytnASqJUQ3ZaLITW
WLVrTOYeZ4KmF6p6PmXiHvw54NGEtgHSlO6KQC1W+ahn4msI+hYEpV0dPEvgt8TDnn8H+uqkCJ7u
UTSXKc8Ph1nLgkEf3XMVICils5Y7cO4E8wcNUvjha9WWOJXW+l00OMZU7XTM1VaT9MbsYZYIkMjG
rrwjlx5ogdzZnweUo5E1uRm9vmp+7MxirhSMlo0Zntykyo2cC/LtBsgwNhsQrhXJl3dipa4S6r9u
XV3kCQfQshlEdD7DcfPzh1lEjahPjs2FtPcGNcu8vR+KAKOa3umBhYSWhJdLcrplP5bX2iDz7CLW
QAGbVF8pcWvsDC7ea1HQ71RhW0x+t7HEieSg1vjdD+4/gJb2II8AgDj/HIMi0Yb5CkAk9bu+Cv2b
kEfYyPl9GtsgmTVHmuzXakJqK8X60qyi01eAdztQabMWlY/bKl91WGkjqOUOuUr/MnbWxIxftJE+
apwNmetDavGPEpbDbuOUuju7CwCyj8SrvtJa+gazBpTEPqfIN8ZuUEFXMyvVBVYfnDfImkbGJM1i
opWEQBP3FD0ldJunUH+7IAzEZaQCXjpMCO0/Xly+lx6UZkWvYTe2T33Z7mZdIeTnuRvcwTfKoGJn
9qEijj0d7ZOm4V0lKwJPncAAxiiHt04IVWDCdtXePEFyU61l+1vdHVrrwVAkuUNorhyYDYs6tCf7
Z+nzqQv4QY+oUgbnLIj0Brp9h+y+LYtsXyvk2TGnB2Z1aWS5sGKiJwywJJl7oEtF3Y+sVTTJQqaU
yrblASds9lRIM5Ke4MYHktVoxUAa4V1DcVcFGg9YBGCfoi2Uu70FkkOWfF/tFgkOqfwTNDA8+D5n
csLs8IDgCIAF53AocdSjNFg6zXkd6IhzE6KJa/Rkh/sUWlSVEZE/iN/0SpHhjaqtMYWc3EceUy/g
ZqnXkGot2mhTjfOivcwR0XTvc8HmM4zx93J7dCa9TSA/+htIkMuVNaSrUZi2MQnwmiInedTwhMkF
yE5iDHZeSZj9HGJui/3mxY8BB/VDfeywJGnBIYnlfsEaLowD7+F5c4NRj8cAzxlg9dEVS0NMoL2W
rl/d6t50/oX4Ie6lKHkFsHGSkmtaHL0eINNn81Xh5j5u8qLp68VCecoES0Ia/jGrUK8DOMRfl6Oc
czg55xeC9w8ydsXTRQh9/mvuCYf41GhxouyP4xzBuDdiuNYpHGRvzgGqYLHlg0dwh69anVrMLaQN
o4MsCD7roR2+TC25PgsTFHy8OpStPp0uS6Dp6nio+9+Z8F1yy9aA3psCXVcaaoidPpk1zgskz/cm
iNNkNrDKLyYzkokIbh59HM6MPD6oBVqE8B3UHbl9q/vBjqJIYCzWpsk4Znw025crTnmUCr3xOf7v
HyGadNJHwZAyQWSYqSlPIJRzO7upxle4mh4DVRsvop5MtTYrBMETDifpS7sHdTEOCvs4SvT4cnwm
sJFuR+TlM8E0bABfO91+vjASlgze3MGNf7S+Qv5UmeEWd5P6kT9wj5AVD5xmYcmdPsIgXyVZOwtd
lsG6H60pkmxEik7muip+2TZtWTlAFJZ/v0c8BI8ppwWpw7Upc4LTw1FO817uhKlUQ2hHfrTIbBWE
sqFvARKnZu2B+SkqsH+im9xur79pN1QuZfJgCvGfVnVmDN1UHpq3HfADMe4DliIBW5TJJNEvgZ3N
RlIrowr+e6mmVyssQWTgpDM6UKACQloCmSBhDVbBDhXlFI/B+Pyv7fHqJjgit4IxYfL1Gp+jMDI6
raI7jac8X4lbt17qvKvYT7Zt5yFYUITDXRyMPyX6XKGHpqu6WEU22LvthPOyG0C2xXJz7frUTAdC
TJF6FbxOQzLY369yg4qNxhfCD43fJgRe5y6+FUAHL2MvvOvr5LKi7kGsYJpszubeQ81MEMy71ZjW
/p3OQRIdvzP7B6D8mPM3aDooY6foH0lOD8S6UjhTsxpEYIdshdrQ2GAHqS+S53F3+h4lEu7uordH
ap6znLPkldaBo/jNDxFWgo+5EkDgppuGTKM2RyjW7oR/RX+TqsOcgJ201lkdlmLg5Z4IelYYdOx1
chd5xqJ4Mrew0+vAYsMgltca5kRo1dni5itjuCWYxdJozaT2bOdKryYiTWiofbuU6fjLLDOzBo/P
TRCGsqPqDhWCy3tK1vnsRJSpQa6LumQAg7XUnugcKi7YN3IMEtFQrK2uvm15CBSoC1Uj31L4ZE/O
HopYCYnOUWXKBjKc8iKu9HiS+1wwewXBeRhpyBZjZVQ/ReLwCHaZSmitCvUuWFNQjtT1QA9OwpJ0
TDF5IBtxu7De6eVjpA6FITda2rUlNb/NPuqjBGTg0Dp/RLP0CBREGakcRemDw1hmCJ1f4C7gYzh7
sIfAJXt2KzgVNG2d0jnbzG2MjDAVIlajx5wvR+zyGygI6NWFlpYV7Cj21CaYZvrp4iKA5MJ6WN/y
JyGdlXoNtvZOlInS+a3DifCclIMKUYgFNFnl0aGO4JMcqgNCgH7Ws7+PdEBMteljdBliKXdwcozG
Z1QMA0jXXb6KBZTQYqjaEnnszk3foC3TDQHoConIcfAB/aY9ywbUVU7gkXVUVRHrGDU9CMsZ9GSk
UTcefUg3JMf7sfh+/WCFlDysJQ6O4ZPLOr5LJ373Xzsqsf2f52sNnVQ4rU82YsLfJf1JLJ7cyqQU
QNpZoWXthwiWTZTf02vMkBVHjYOB0DwFytiaI0dvCV0WmhSZzJjfL2vDJqfkU9LZMcitAKpI2ScW
Zt31vf75HiXq6wF5vaEg6C7PxWIWpVOuRRPkC7leAiXKQDYFJRtMPwNsmftJ9KFmeCTaG0g9Vd5F
O3wTf6+YpZG/qgazMPI7W76g4QpPOMjOJ8G6tCdoBvbNyT8dqhGVi/5zXDgXxnHe5vbiQL+BDCS5
ciJ+FNixIvxOFkVAx0DQ6bUianOkuuoDQ9zCRxHNxsODuEyVqrdEHtcIQkNzTVxsv5MkItNd8wXs
TvwbU1GiEciW6XesN4fIBMjmqtoMTGexGr+F+flG638G2+gpdhpSZpTBQSUKeMlshYxPKZ6x1pqr
EOYljZ1FI4evzyq5uLvX1TGBxRaE2mD3FlHzIqmtH8V44RaXw5rTK4usPRI8QcxL1HfBeJAYeyU9
zeeFIfL4h2sMidINRm6FFLzTbb0XW5lU7Vkbiuu2zTdU400WA8s9uZqOQfakaV+91nmlg8PZdVZG
PoOnQUaHT3h7Ueho0R5pzB5hDBxgBn0mRRgBYrmdM329LY9PQObDi1dvsJmqWLN1k5DF2ZqU4m9W
Ogy3KitmzUlsmKwTmwfobbHvfPBqCl+bZZgipFEDcAgIS4V/V2kLg9PKGIQQcQVLk1bsqCyE30bB
dQQj9e1iufIfsl5FzRjWMJuzSAXc5a3tRqi2MbxW9F9eWr79muYfDXBjg9vXIWLSELudHyJndcFR
FRTAkVAcjYPwd2hCGko/UJLBad+XrnPghfuLyDIvpjNDPkKykb3BMlumZPslgRjmAt/WTngBc8QW
NhlcrSD4YxAXiueRiBxq3rsnJGVWg96+JS8xZ+ts/VwSySfc+z6OUew7ImxI9VRa4nGbzopMRlmB
nbqFCEf0Gszvq2KQr8cFJ7ti/vGW0toDjiobysTV03YHyCmDwpcPKLLRxM3Bg3OHe975zhMTUIi0
VBjaiEExVmqko5fnGvZ55pOIFe7JTuS4k/0xW2aFcxKFrjhx1pqvelm2GCghHVkI+TtAlx8LlV+e
xpkNnEYglLQxHlO7vvEpO1aaOK7rUcy2IrtdR+i3equIAdjwJwTXAgMmaOvqYTLKHoUdaUtPd8FL
4U1N2H1r+otlBK2qLqb2GOZLSIk0HvBaL7dDE62GW8Q75htD2owvtacscVEkSd0Bh1K6jpdZXfKg
4Du2y8gfeoE3BcYohBJZMlHYWPkAoJ/1bcluwc+cnN5qjiFoTuDucXRv4++VLKU+iNMMpc4MxLXu
dftZ0Ilu6mPJkfFsy+We916lDrcPHMsSdx6vCA95r+RV29hMQjKhCZ/R1qpdHhJowP2nClEXxb6N
kRbWNezqIZz4mpANn/boa0r9NPuX7xt6zQdNdCY0hdBLBetbBHpwmnfGl9NykWvP5z7xReg3Hz70
F29yLI6POi934eFRsIziCe8ZZ4C5qwvimCUKJOCDQx+/Tp5Z3VA3uy0ZloVPP+n05aads641f6Dl
7an1AdSzzKEnydMfH0FSy2AUUhOSE7lCEf8rk9nWXAia0LOwwO/R6wKQ0c9fOgBlOyGGDgp9pNYb
BSOMhG/GcIlqDkNBPAbPN0V+TZEx1RZPnUIPLQh3O5U/AEg1w5LbjDsMdo9yBX1uZcPhdCbkz9oh
HMJ3qCyeisdzngqfyisUtG3xa5HPKRX3smzo43W3m6Z0CZ3bm2oVVkLn+gP8mzeJKoO6hU93qr9S
Vv20fz3wZPpYIF2oGZ/7ptMldgXs+l/ZfFnZHerexeBihorrpoiR890Qt9rPULEGf+YHGL59OndD
vlnk//HojkzkN0ch17ggNrY/PWBOODubRemojOXFSRPMa+GI1ZhJweAWkSIISRwyeecyeNJmRVXF
2pB3/yawmS0CTD3UVB0oip3pahS/uD6Y1k7YPd6pCz2Bg27qZK+H3TB26cMsbIxFFFtd2sl1Yv6F
WBTj+pzbA1ML3pFyoDdU7DTSusG0/kJLcxEVbYTl7FqIkHsZ9AKxVax4o6ASUpn4pjCQRGlLjkvW
aj5HnQWLezs0uKcd8KGAJ1J0Tq5LUKGEYNuxHF6uSCGSr56R34HGDfmjEMXI45CO/v+mFBMhaHR9
nShSlJvxd3meAVNwxmlarPf7UVnDRKUAIpH6QHJ63yJdHkYNyi1LeOPuxlGKGoIvWFIEMU8E0cL3
tS3uqbe1ST8S81nfTwQFQIunWISBcc6z7Yu1I3JHA5GkwmOBftMlsF0JImipWx+yRQPokL4xm+rR
LwbV3oQ/EDUKrx2hXcE5gedfBlmOy0mpZltVlVrp0QuP0qQ8Pj37gdkweH5GnnZhl7QSZVbU+7EI
SNnytvrDeX1Ge52y2H4jVGP9bzhCTBSqWhy8JNJWpP3ihMMnH0paU8hFO0yTvio3i3XiSlOl2GfW
or59w4id71/2mDzUQ8cRD3HrhPfzBPubVIdiXD6OId4wQqHuw8j+uk5f+X/RE/4aODvK9qnEmpx/
1DuHulL19PttN1CzOI7ZELrvkBx73jf8bJ7oWAlzc9rjcjbRQY78ChDzzN40J1u6DX/scWaOlbdR
TShTkN1J+MVisyp28Xaq2qUmhpbzj3Vv+ar5i4VSzDo5FJ1TjRdmnkh/0bDoOjOWB+H3N2WJ0ht1
isvIiEDKZj3idgLbenNXETD5iIf0RBlTyG9hECoeUnmYBUiU4L/k9otXcvMDLUBcyyeEgtz1FGLn
NG/qayfCIt3LRDK9eDS31lUFyX8Kz9jiwsgceU4dCA2Uh+6YEDOulGzE/2P6GA6bVXJ3mOK044l5
grCntK2EtKX8mhfKy1e175l+klKWIuSEcARfxh6eSWtZEPKkGTyaEf6xvNEzo7ApsTMs/NenU7yp
V5g+VHUafZM6ifbp8tLyyVvPBpizJmsIfu/erS9c2E/0V8qXFjyWQrjRHM3KUWUhoTvE7aPziuYW
QGt+mQzfzaJ5GJpHVRK//seyIgOeNpuS2Rf2bWWB5Tv8EhFoqGWxBuqT1kv7y+xyFoIzonQ6rfCw
YF0yTcVyiyn6luzqZsr3GZHgaA9SXXrzEKgpk0vA1SnLnlNpwxRQGF0KkxOMIhnz0oKBwJceIU7X
IZTtN4SeESZnzF1jQPxmCTFYy4UUdg5il77F+kWmrgkXXeGn8a/hahyapwbfM0M/13CQAlIfDpLe
yfczJhNA1uoNcim0302+J1jwlKdzfOThaiiji97Zr8bbwMgunXu5OGBujPIeP4ZsAswhUAvEffJg
nYuB4C4WYZF2HnoYWy9xrzlf7m6iBsI8uWRh2YY6705Q4zTe+3YSfYEi6rfwmfNCLgTUvny7qWEk
Z9lR+sYpDg3NgFGkeHldWrzAQhwQ2J38PLFrRoinI8GmqgtaWY09lV6qnBD/GtqTD7m5kON0FNgk
QXfqkR8mj1lWedWJovpkw72Bxo/KynrWyz+x3w64tGl2lhbZC6smBcDDMf14tzNFNlGqg0NgWpo/
oxYj7FNL9ZbNzKNNRQZMFsXdOhGG0uupeIsANU7PifNGAffSfe2Sw5+xrzDIPCeAcEEIfxCYo/bg
WF4D4i9l/B6pil4kVOMzgqp1WKo7FLiRMDsO2IMXsj5P7lECQbKybeOIYJ8EBS0LtvpFpUPfQieo
xO3asjlCTr1IkxXJkj/AFiKlIfQ5GvtbGiIenrf+2ql4pXztGVKz2iW3jNpHTBivAxgMEZDhcvS9
AJHE7Ml6jD2ReCjVTLBVQNoDtxTnxbYGLT0vWyhU0QoazvpJjLPQT1V3daVr6btWyeCt10vGLwWF
ZvWC5uoR333nArPhKFzFuY44BkSfUayCJs8J0grsCJH46B9FGlhILweoc4AxHNZFoz4/loWV0gUo
sTpRlodSxKbRLgSxs1vZjAAKOdsh4ti4aor2/v50xaeJRRamQvvaStVG6Y6RSUCir7MAK6Ly/py1
UhyO5pg46SS9+9fyiWBHt6XzbvpGI8nxyuNzYmsQ397gweqofl9gK7WIslEg+Mx0WCIJA4EID4dQ
zmLfuEapyCPLNmcERTR/+S8Wk4vaVYVui3YmpGSQsKYClZykBJKgec1OTKsuCznD03T/oBecdLOw
dsPcxXOzdLwSicG1svvJC/XUx85ky08ZEcfa5So0ILNcry72g6Byp5NtpB6vYCHUL+cWalq58C/p
+mI37fe5iFQXcRcazro4ii5kOkEXZTFNc8LseTbxZfn0jDvI6Q3PG937L39CUKnstx2HUgZHtUTT
8YhMFDk3zm8OXGiLB275fq5N1E0EuoqYMeiFA2mhKdHGbyMuYPvZ23HqAymKRuasuUWDxBkBvNqF
1uS8N7imTPgRWWvoYjxwVejJ2uRQQ8kBkWKo16UnL+iHn9W6M71pYrLw38za8k7yfmHXCiDZJT0/
537+khLjn7CG7v9hJIlUnZSt75rLLCC0QliOBOBzUUfgHNZEB60ICa3EOj9V/gmAr6OaySYkVZsJ
hnuym9aHNvctdTddrTUZS4sBAedVvLUJzkvHnAXIOzcEhqJr3o8c5AZc198L2nbODeCS2QpOouQF
VLmFzjguHLzHtJf0quUiIyXM10rclgcjdx2oKoCR+wZiriRxaLzWoAyyMdEOkLjv8CWQgkn4v7Su
38v1g385v64Jbe7GxnKn0H0/MqjXD/ZQazBJT716c+jqe1Vjb+IsBHmfEDdkteUz0HiJdhjX2om9
1+1TTDt05+9R62bUgiMo3UA5BZAqlWsBRJt9Xf2SR6FXbUND7C/buAk+MOzbnhkubriii3Hi3RJt
+CMTm9S+lcgN7Q9CNuoz1j03SgKy6d3vxpaL4ZASA0T/dhIxDq6alKMxUdXTyrxT+DkKkrz6N/i+
SEHQbVUMC5x18Q7lN56o55Eb7efzlqsTno/WjEeev2SLvHR1IdINYJ+mTPBI+2gG4jKWIcttyAH1
q2ZP7RK99xwLmhxWCR+OKI84Udg5LMKEIzNWYuVkNeMWg+RKT9ya5WmS5z+1oxOEKid9fdovDNaT
LOAi0Ft/MXX4bYKia5hqr7MTp5mMqmGFkMzkHyjiPNxkfBbLEZLhb+DOUuOm89qsieqPTUWj3Vz8
uK8QMjxJg5Ehd9/VeHXG3vlnV8Ql0f3IKZ/GlknL2cSOdbYfjTcKSyC/y8knLEufWEz7Z9PIkn17
EogZYMQMVuuN4i8IMElRLqC3QEIJo++gw3CAIcPGvLX3g+BUxpYyep6c49uRD2S21O6MWoQ7o5mY
NNQL1Xc9GQwSBb9lkVVfEYcro/X9FIDTXVq5qWySfKgnmAp5TlHOaxerb8S1J3HnGOGBgxeqNDy5
4SdrAJ2WquW6uvfF0B19gyssfTphvHiMty8PoHHGLy3Cqvr8kCpjiue8YHMqEHv3jS5R6kbYqzkA
QN5smKdbRX1x/D2u0sqi0nqUrzYWfy1Cxu2dfQe03z5ZNg0tLqfNwLLBUR4Nmj90uHxcHR5z5k9q
muEftgjIaamS1v6yoRO7b4c1Dw7T0cp8exhr2fZ5m6GT80bZjSJLR8qPtWFoeQIePuFvgWE1opZg
S5wOqo+T+U0chYhW1c5y1SIeB+94iXT4qcobDb7+WD/UBj/Ly6LbgCiiDnad6dMMVkbMjoQDHI39
anFLc9KB6PiMcHNv/MXnHF4JEyNzYzzTF5DxMuu3M5v3wzNYXFJ1ZjHRBMBgOEGzmSVWmWADNxqd
Qz+/yF5z2Luhm1UWEeKlxCEd9ilovgpUIIQmuCv9ORjTzI/g7mO0KBazO8a+xZWT8MdTj9fOvOKW
HpkKCYCh+8bFC0S5TFG/9T2WXIqA8ZHoypwhYHHANUtrzsvCFOSZZ5eFGJie8GJkQHcY+fqXKzG2
fBBVhcAUFd4M7O6+rj/xAKXZ9DtY6AL5pIczd5adhfwWO2tryQoeTge91idw2K5DSOtNJqffoOz7
tmVscYTod3drxnVl7qW913Ulpc2zSHreBrqfCyIdDmXjoZ768CBW9CYoEdppxfVW4NjNZvgHqfpk
mzC/vGrVP3wkv8qCaIpbj0D/kWSXKUYPIyp1nbqkJKp7HyYW7iJVi5SdUYHWsh6mFYXLMdQLkw7x
lpSSp/vrV1/+BGlZrzG3x/RLBWr+wEawbzyBn6HyXGBVDtxDuKYi2/8Zo0buaNqOzxWqhXr5lnuG
j/MAdZYUedy45o10x5SEYIv2E+KjiF2DzWMRxGSrJJga0T21t7cgKW9vPtUuZcYxsQozbMekv+SQ
dOBLUjTR/EntJJKwTuwXYb3knNHGlZyBvZ86qZR7cjIREA4NVRjgtyBVkKGwBsnyiO5UAUOGbrJO
Xi1AhY1zc+YmmnVQMizCdaqyv9Znb7/pLVR9vUcdzxgdFH918f5+oZTPM+O06ugQnArDW0E27mbI
iL6QPW2xh0/G5gi30SMRWqlyvRgODd5csddriMQvEKb2GjTVlQTbBFQxOzq8/LqN9xxRfsx5+2JO
OAgcDfj94I1aRiyW2WFumyWeGjG6ohcZldobxuAvUupNYPuseWR7F4t/rfkqmslpiwasiaPyhoa+
SnkgWD+vEqGbkuQkTFEG+EwxpXBrZSHzWBEdlPtd19V/qzuBuxYH8ANvW33VXproKCCIdLYLDgdf
niREU/TelEGkG3q4/HGIlCKgsb4UnPxdCMiShyjjf7lAkaE0ngPe7e6osWer4xoZRimHVqf3xWIO
3GEa0sg56NBFCjTHZTAov+wVt0EDBN7tWWT6Gop64ws9WR+xVC7YJdYF8X4el5Wr7dQ1fBZmDC/F
IBId557guF6qppAjjncYxv3B08dPw+PzzyUOSiJNcBdIERtRLHkVHHZvyYsgK2elBdyqsDLzV0iC
/vZQuCcLrptXLZLMhfQOLfjfEx4/NlaUlE/L5192FRiE5MivmC8jSwEdzb+NFiXzfcEH7DQS3iwr
+lkrYYd0bcewO+V3yaWKjb9GX++1Zm/ZkBfSzWSqxnI++VJpnXAz+bXs8dqneGCbdZmYzgvfBEJW
qqT1Qep3DOYdW6KVEipmrPT3YBfZWPKo4ZNYIkeDp0Yn/lTIT+CbTSMaOIr1FZiG8dhNfjChwTIT
PPd0QZcRc0iFpeVAmqddVMNTftlW8fM8alHbbQ3ib8S69Rci2FeA3HyA+FYmGD5c3HZNTFsfvBhz
KLjA/Tr9EToSnj9kUaljGWgvql9ntg26UhV1t8xC0VOjaEOjXTc/rfot+oTey7HrXKrwh+5AkowS
GOk7WFjb20uDNCV2XuGUS2bDQbhoXfz5r7QPdvlgWzElr2peGiBh22BD6fO3NzFKB6YFEqD9u5IM
LDqAmgiJF9ofZL4tS4QVfISkzO+760m+/lqlxXDm4NzYkIicl4QY60IIPPvcdfzftAXIzFP+AWhO
VGgd3pYl3CDWwgEVKbhb5CdYrIj/chWJY8L1esuFqwrkHP1sUoRXDwF3bUTudPcZt5K3K2hWku/L
VqNQ9YGwb5Pe7K+75SHSSEEZAhsNtHUbC8VPlI/4NnuXDeTsVeABb5M39ZR3o6YzH4sGgP/yZka+
ANBPmyVmJuVMy/hVDC0CwEkZ1U+DrlejyFqPsb3zmWfJ13TrnNrLGfkdtN1ZPTYQlDAY5fTw4UaM
HCSAqGMdrDCKXz2p7j/UMUL+mMwD2gevn0P/2DsNi1BggrJSZriLCYXBQWEmK1UQJe/OF8UfFTIM
ZVfQBa7rWuM8sTFYBw/gREKCnmVzhC5dhpNbRQ6cz/1T4zj7fUzh5eBDaM50rQD00eOkkMT7Yw9L
k/rywIY9DnTjNVrMucMz/+xK1ObkuK9zIsUScy6Hqh1asDpHL5Ywxg8tVRQsY1iBYSB4BhJ68dAt
zFpK+iIAxv0kTHJNvBfnuFMaimm0mF4efh1MKjho0jWEdMMlLPctgvI2zAlN1LU0R2N+x74V1IHX
bzVZIaOe8w1bwwDN6somgu1tndzwVnjV9b2Y1oyKNXU8ByEC/Zd7WmlP2nEW6at14fzRwmEQDtKS
iuVPYUhAL7xo+0WhSGap6p5eJsdVAcPiRHYX7aiHCH3HJ89TNE2sDyRmg7M7GPmT3BXD0BhiDfJ0
NF/3CsrcVOUjlYBtNGMYUAi/riEnvyk4y3aA27Xcxhz1jCBi+BCCzamPxCB3aJJbxaCZ2CaC+VnB
IRO6qRt/QM54RQ3U6nDXN4ZvzJp6tlgFpdXb7ExZEQofRA4g8T9oVddyee3ZLa6QAJR1IV/hojuM
RA2sTiKlg6XuUB6cKvkzTmG2XAMoCbcxgt+o+PN4YbZ872ISz5BwUBKqcYjGEUFb1KC96LPl+a2F
XkWews6+DyVQAF/oy7Sry4QCBr+PFkx2KZE7JacaVi0IiI+wcdc8qabR7LbAxJmR0wZg0Yi+WXgx
g4sfiNFstohu5CLw4NEFggQnIDuVJ+OyT0V+qVuAonPCSDrwApyWhY63zcEzUeIKMu/G9+vgbfzL
uN/j2+635bL3JWK0lhiwPPOtKYhbLPlqN0azaXXSahENccfQcRb8rDcvP0r+3bvV+zOp00/47dbv
rO5E3Ygj640qRLUmqkqD5vYzVUnfgS6TkSKxAD3sAOhpL2X2P2wKG7V0QCyyd66tWBDkuERYeH8B
tWd7Y2GjNJRaJxeg8j83+qg3g9XZZOGc2lYjswg97Iu+VRuL1iGdpTuaLH2ztmDaAAmVdGfhqiNO
1aD7W9i0oqGGETp3ru11oc5Ep2Ae7JkpO7QI2X7tAH3eOSgzA8Nfnh9a4Io/jrh/fcaCqAE+f5m/
2/Z4KsClWYfhxA8rVLSajon8LOQc6jRlbin7LEFAq++/sfmU/xuE0VqJECNb2RF6b8wr5YShzpTk
k/LR+ldAe3lk31r7s47T/skZl5HcDueyzsbyZCd0OAVTDl2apxRuafgmCgAqyEhviAnUDQmUnhGn
qSwZPIihJIRnN2IcIez7G3vO3nkQaA/ALE9xNKQqlVVRubZdP5WpLjPpSmdzxa7JYroix7j6LhVv
ui410MeZIHRbQhMzj8dBVzg2PFu3X+ValwGP22TYnijE/dAU7+TVgRyEt1jMq7SUJppGptnWU1Ny
9h+Sj+yweRNPihWPBlxTxwmeALK0ncCTakqYuyfdKfDRE35rw1f9flJSrgswIHZIUOcxRmnf80En
YBBlPduc8ZW5y6wVUlISJOVgsLlObO5CwGg0UMDh4evojQtNF3w8MKMwFaA4Q45Hv8Wxv63IYLrb
ADHR3DduSYSmWTdkpMTavoHb1OTswPOZaaWhMwzKfoFZ6KrCAd//yda4WQBmhLCeONy8XPOXyhw/
xeH19sHeJniQMF4USOY6chRP0tHXQfnryULhTAKdbngm6VzsMXGr8fAkBbm6vCCvcTUrMbXY5rV2
qke/c+W3hLTnOSBkwYtsTs2hjJavMbb/C3BjX+nxAFalTIEOnM7nEzJDd6PJMCBSTJwPdzP4q5wu
Jy+p4IlJv5JiIhgysc1XStt72QLZQpW2i6AgdNo8aaxYLlV/BGO1jGV5cp4lROal1Judlug4Zfks
c22iWTnsSj0igBJDVoe0zybqSgK8vYzVs7rPztx5/nYhz4Zo5b9MhMfXwVq9/WbpCIgtOX+VwKbb
hvKikWaWscDotJuyVSwL5rBlw+EaEK52LFMc/k1q4ZceaPdw3PNftLlMqzhatcREK6/6jWjDaTco
Zxx7/P+RgfskxVeUi7GS8jfRyoFFKV/L4OP3rYRbQFSUZlFzopHrBCaLH8ISilS7Bgi7klzJyqmR
Nay8+d0ZHlGYEH5YNCQKsVWctk1Na+rdsrHHv40kEWQjVudYNLks1MEDMHk8iOnibns54VF3jawn
M6MjAmOCbB8TNWi5Q59ravxphvT2bzENGJQXfKsYpvR+HY26eueZVjoOyKNX2UjO/RYjJS1x1Wbf
zJpee074PXXNsXfDPru8h1mirTOVnKx3c/zUxAbj/RocemRoNFe55Mgpqg7TM7QFtwdfCz8UxUgs
BVecH15EtFwPLrJTIUOSQeBWOfIx7bRw5xqVlWA5HFROmsqoBNnsBqTr2R1vVpHSqMABWLnH+nOi
OFsDB9frLD3G4XxmuzY0gKnsYYl1PDS4/yCdkwccCfSRtdDq3gtNSFNMdpKn81OMoYnL7reNqkSb
1alTHgE+o9hpIe/c+LJP17STpbR6IEDZDprylgb240bwwrKxppWmiwmdPlu1bLoMuMaq6aCo+q0t
j+aYOu/EtTYdY8RbREY7KI9ebUxmE7TvU/id4HDdptJl0824+34CwsndwxbcxgO1byrYTbSkmGJK
T6ivlwX4PUtE9S4y05b2FuUOs3dbf+VXwiv2dqyfD5jtEe+q4xdpNVw32iDY2DRJxnhXBAK2RhTf
E6fQtfcY2NCBeTdtOVFZqq2WFMZBfAGSr9mi6hRb3i1FEavftjmELZe1J+vlF7Il+O251f/D0pNN
EDLsq0TVGEmmrSgrT64V3ZzkijAsntXRjaWn1SinVigGP9J3x6/ZnBxCZIPQG56025lcUVYSw0JL
TQwoLs1Y3sCF9AqSslciuJ1OhoEQsc/UdutBBaf1vQY7EwyxdUpRXgLCGW9l2oVBes31SEbbcR7U
kTMaNYcXGsd5NiXWr3zZ1cxVNKjjvFS3F5qEXMrnaM3GFvtSjXzz/j7TKX86Fu+/uYM8OcFZnfx/
ddpJlpHnijlAMEujyElZMI/+dUdTCUBi8Lz1vAtIxKymdFAjCbl033UOzD/syQasCv3+tf/vUF0v
mkIBCdX6ZOSuqdStrCS0c1DX7tZfJe9St44z9GfCrPCSfP35OxoNgw9sIpDHOGqSFwCI5RoQSjKN
wM+UDOIu+gHFYtuGpcNSpx/wcVL/siCXt6L883zRLI+f79akGynLmZAPmNkof7/bJCD9rCVLPnAP
Sf9NGgt5xrwgQmMPGbe0ndNiQc6mTHUTMR8pMB8uZ0r4EAS1uL9tHTMJRaFNPgrvfGEf5Xh/VQDQ
eroh/QPO7nl7RfLDkKDkLLr4psCr2mrFwkFbXgVrC2pl+h4pU5Wf7+M8m/487W0IXHuKKmkzqVQ3
d7/GBsW9DQ+DBxgQqf4LW1ddeJQzoGrAOhSRtKW1KW43ElovO6urk7MJ8GZxQnQxaDjU2F3auqBX
EwJGu25mNaGdeD6qUdaF1lqy/OOCUsE1YjFJZkno3g0Eh4cjhDztC2fmWUpfPsx5Xii7CEAS+L8K
8hdViVJYS7C8FjZkWBZ0ufnoSLs7T/33FOD48PuK++ror29hju7X51fXrrMlCdGsu7kRBFOHWzeZ
x99KSBtEgHONAfOgysD5/D6bSca3fe88CrBIqjpreHjVqqpz8Hq+oWUBEY5EZiSM36VGPWwheNFS
67I1L/Glo/q9MmhHOIysJ+Qz9oSx3/hQxRTFLfXyD7rm9GWFeY2KTHoXOzU4dHHpFSI3lLHg2zq3
l1RBB4+TDOwSBb2pArY6VXfReHij8wNUo80Fx6wA1dfqaIO0+xsxJhsCu1260iSVtnq+EzQ29VVh
jab1NYxI1bOLDDZsXFFtXcPDfcDxhUE6b6NpAekoRNQZafpDExcCES7J1kz0ju4WxANjVrE/5xcv
TOyZbgLiTDp+vKSZBVHyFBBPcsKIt6D7DEUZ2MknB/uFxpoVOaLS5/zQupQVj3z+c2WuyC351kyt
UthIJlIHZRr7ScJR2F+/cpLqA0RgYYhnNH39xa6q1M96c6YuFNuDB3KnS92ZogpqXh28BsycXVZv
Rz5aXhpS2cmLHUKDNBmZj5eYba1LcPsGWOAFgC3lXJ/zTxh9lUmoeY9y2qnorzBjRr0vM8SuvNfh
7o6LWm7ZUvNhrgXIYfR+lpDZiXBP0d4xPSDqXiy3UQhkA3Kvx7crfP5waQe/ulWWrbRiXWpwi2Du
bI7TYemXfv+sCMlU6T39yi5jLNm2F15EA9FwuiBYQ9IvTL5BsO6kernh7pTfQoFYMxft+WfxgkJV
zkQhGFmFmP0mBqraXpkB6m8Ioxi3I51WPJmoy+Q8lWGqADIM/aMra/ns4MqRORNNQt2r7UC1qKWT
SATke2xatlRrNW3+xuvxRDpjCEDxMG+Ee4e4BmDqZ6cJTDw30VbeYp+Sc+iIgSU517GJyn1l83MG
wyVb+ro6PjV5/yJein8K26GElkgSYlaB65JesDEAGx1M8zfzS/1idtGjj/YGjEwmP3/EqeJsWp8J
K0k1KGWfOjx/mSG0CeLRpS0M+ggZDYPYpHIx4pxC/X5qG+WITAzwVevPWSRbmNffjCumEKKYkfWH
/ocv4EwVKIHZOsq1KxrKTI7Bx5xXE7LZkESxSx9HgX8ZSELUEoDiZa6fMK1qvlXsZfmkPqf+c1dS
XvD4xN4dL4kduc4Ad9R8lt/X4S6Z1wk9mn4aNiAM4lAVc4PXjpo/NuSWjPLxmJdyFs6nZt1ZyeEi
dwNkRYrb+WkarhKv/9HKt7en5cY+XfqvdR1vTSnbCVkjFyUpWaoXbZXZTesHLPthrQzVpJKZyoHY
78IUVVYR7dB4Fc8cRQSHDLhnCD2eoV9lMRHpSy3aFQwTssXrPnU5ZbxB8mKX/zphn8q0d5OftbGx
kmM2EiYozgUVzAgIn/Id/lhfaxtkxAHdibQfOdRJTU+16Y9Euui71aJleKCEZlys6QqVTa/qimzQ
JNFHypzTc9S+hk2hSXBqjN9sRLfMaVf2jRKqpfYL42uyaMgoRQBN2nSgqcs6tk/beSmZuZIk63se
SFYXdq6lbr6/9hY85oe7XQGGLdabJaqHcDqoatEYhg11xypsz7nghgvDKJOs/2DyY7rRjPHQG46S
4/DvXieMqkIUdzgH5Ct/0pMxmFr6mqDuj30NRd14NXNOvhgvL2r6P00HOmQA01iiw/po79cRu4Ko
sgXjnbq6sdRbA7C3UI/c5R/m6JHiCEuJpEWXmuHxzUdIOW3EX6pnyxXzTUleBCH9TrFS8fKSTNiA
raqwyb7IZTS8jn0UmDgCt+PTlpFWy/iGSCyXbyzZs6mE19k7aFn44LYkJ18lT6mNhmiPH3Seev7G
l1uR0LRplLNdPrG5Kg1X/CzGeXht6Uohw5Xml9VqFo9OCMPRo7aX0K0B7Fvt3PN5UkF6yjpHkn8h
t02ypW94ggY9pYQO3bYF8h1zLBZYihrAzsUTD5BmIqlf9aRRLcq4cCbC+M0JlWhmzFEo1dyiSmEI
Stt8qiHVRGjZgut9vc5OIbW61iUiNZt7kCjWaITxXv0CJQ8pf0Lm6u2FCSsvtMNRsM+3TM3rEnY4
4ssvp1eRLaDlbVp4PYdsG0yjG8Tb7HTSzLrXvMHERuTHb3AfrhoN+pG8EOd4tj1F4BzIA4ZfWAuk
vODmaW73yHMJ/l7eKqUoSZxB6MLznUxCU2GfFJ6F1zzoZzWlGZ6Dh6xICwk5l4Oo7HFb1ZWB5UYy
TNa0YTqTntvv1AP0ESO6PrRIzFfWb7Hqu97PsEDADd5L0LcX/cWDjB7oekhrBE8X/rjc8928gkHa
LhS7EgiXzSF4R8+4G0ssWOwprOnOXmLsBJWWXwRk16DXpZeNaKho54TjlQRAvi1CRuBSqg5kuFqS
lDCIufQIVfY8w0I9gUEK3uBD6RWO9xUHdtf+3UEFIDJMUPXfnGmbx4Xd/bnXwVoiAxrgKft/FQZh
eIJELEHLAtI/dCQsPZGEKju+z3FYAZsaKLsz4IWqtGADTYakjGpV2DAEH/8VF7ynjFVdbNRqjkJK
BUNcwIyqwZQdcfzgxeyKpymiGnbiSTSKhq+qdpHBf8LqCDvoWrzVOiZsoCyP2FK+N+HtLGnbV3/f
Dq7l/lgIEC90VWsplTrBDqf2G8Es9ZshDOVH7+lpWqKgmm6OR/vfrofwumlHT46exID9XSDU4cMl
0wPLS3+boobu0sx40tVEm+OefBHZw0I6d6o9Pf6UxOhFE5W38KlUpfhhnu2NapmZe11Fz49nBRtQ
rLdJDg//YvAA2SyB8piZOlHjOJJQYCLAWPtcGIXjPO3l3ZYetPFA2qOp7nSE8jWsPrGSvNoRwcru
YKOh5dkY47AcoIm2xO/Rr52ZicDB6jBNEaA7yliyl2reFTuURtDLqRadDvEF0MTSKdXWTGnnXrXS
RYkQIv1oww7zdjs5/xftPME8zTQ56pfUEGym3ev0AiG8yk7a9/qg1XkWvV9rIbxcy3V/BhfxPc4/
klZKrzlNmwQLc/BzWYeCHWusz6fmVy2cpjbZ3LhqvAA1B07why4S7tNGhKvpZYvM4DpnKru+dBwv
fHIiPRMQgEiCZMLUMu9snfatT7moVjD4rSJTB08n7Ce15yiALBD9YVH6zbY3Qul056cHGpDK6tJ5
E8mVSf5w2SUNFKlaJXglCaVKjZ78JbSaonKsC62oAsPSHu+d2Qkwk6xyWUmK9+Ow09rv9xJEktkM
6XAkIpk3hcsu3802W71Xm68RDL3wuxjLlkm+dVrrTEV3b1CH7B7/btV/oYbzSqLEspPXxBqYkW0f
uk1r0ndlSR0F+qXsR2NxySO9H1QnJtW2iZBnPJYgDw9LncPCIk1rOqnCFW8I25vwueDaQKaE/PGt
UTLGesWKkHcV3RNZ1QeB4J1OuzD7bdWUex9OpnMJFNSlN5dwIpbWlivAvI/g2FVkRTA316ffXXVX
Pi57aI+Li44DKakqNDkAp9HbwzZPyCrRWAVWWpZxFZYBxw1XXBHKhBY8GqrAJltKusOF9cQrYZ3B
u9EeBpeNCNDFxtPMRMFYTRo7KesRky4zn1UOpTQH7mbRKPwTXf589mdUmqMAP4aPPt8LiMPyDVdn
JdgDqd2xAlSuMTcky3YEagENvtnkSsSUpEkRxtrfD5rB/qI54SJghmeAK1UBY4NoehNQMn05SeCn
Xv4N1VXHWI5GZsu2dUtVA1kvWgzNdmHggTwyr8g1vWUbx+rhGx/mRkiEThLUmrT2rllX3TJZpf2E
YHKt8SNyIR+eSCZDsOg5v7Jyf3D8fCxsB7ap74RrtvWeggwMGS6Q9EK1td0MUoGdNpuSby0488Mp
6V0UGtJfAre08PQgC0lUIqqSFiun1S1SHcWwtMtGShV74NTJ6ByG5LHPZy+wh2EqxlA2JZxHEKH3
mv2w5QDmHj8fL3OgpeVTYXb3qiyk8EneG2HOI62qFxO5pVaYD+wy6daxXE+7k2S2qCDNpXudi+Rb
D4XiAUNiXx1ZRlpSLFfW4F5gEy25YLt5rv9HE8BfdOCIvJajOzS7cwIVdhcGLJOgTYID7Mbxqs2R
DJaGEhwr9D1leTIyiEuqqm2uOVYSeXCGsHEuwyXNQ4YGfglKa7bfrj5BzlE2XSgbXdlInIz98v8Q
HGDlf9eqK6TBNXGucPdFfd5w/MTiPMWLCjufgH25lvVqps6HWooXWX5/SDT/zZm2y5l+PvmbM6k3
YStP/ZtEVBvNE+nr5ou8Z5PWo0g0K4IzFotvJOwmmBfiaSvrGsuHhejaVtkzqIib0D7wIz5sRq3W
0w9kdr9178ywDE3ARfn8FyT9hoL6xSUabbABiTkdH6qkGjxH85v05bvTk0wMqgqHmRT5fIJSIVzW
LnuIYdVRlFX9S3AWCEICOBU9prp/yBKDBLIw/g5qScrvaPRvVcd6KVXBn5cze2MDVVD9pj93ZmM7
KbXhvRDxSaGbaKkJsDBbPekEUKL3OAwDfKGR73Fdr803LAV5Yaxu4Tk72tcGevX1Jp/k+aVFgUls
FjqwzCVlFl5uW1A1CRz5D+H5DygeAgajpROGwqY8s7K/V1yaVOFeFSlbZVBAZuGYXjTeSgV8Whe5
dSxGcj8f2esUQ+XOFWRpU3Bzm5fwUpp91OrfaVNGY7E7APxVbvgsUjxLydcl5LIRPzTzgLs/1P2K
C/sQ/kG758YMbOTDt+mIaLpOJyg97AD922RvHmnHkQBKHcGzTiaHRGia03izqa+GsrrlwUDpZLFs
5FkEsYfQMV0+9UHf+HQN2GBIza967OmyC3tVM/OorGvFRF4iKfdPMdgftqfMDm2sjlWMRtnfAMjR
7o6IGKwfMuhgxa3nv6eHZf2fdVyNj08WGDzE5gMg2O9Ha1xSQKCYF00uCInDFUZ0sBu1BKlHVE8q
yCZX63lMvrvAKgDRaZNCBfHM9PrBrXUxddtNnUJB8LAH0H52d9pFfxadzOgiFcb3LVrGcOf8EJBH
QVWeM8XDl4YgUbrkq8Ae/+SRFFZ8CFTzlYr1qvdFCMStc6I6jfCW3zlEiST/TqCjY2SBuRcy89Ih
uQ8vMDucQNTASJ8r1lL0RRufCWJ9m8LcPU47FE2Qnpan748xD+IfeZzfX7KYF9NH+/6JtmWtsSch
gCtD3vuY+an3Q1qcMVcIZzLR3VnNZSsWdYRMnfOso3IMeICheI7KO1KEMmImbDugticdnXoMjWwa
VIKTn6SpkT62d6KCgX9jVb2Ed53A86Z14LQbtmIkyD+9fWpwc//40DqnAlLDOJ/v9n21K7lrrcDO
nBHuGpGomcZeZCVKMZmACcPsw0LCDR8pOIhDZhuT+Q5Ay84XfmVdJ87eX9jwzihiVNQ8gy3Gc42l
XOSkoYrRWAO6CggIDydJgZ0PvnmYy0cH0+vt59NDTx1Now5ciM08f39ReLHnXC/IrxF9vbMk4Ozm
EopWsT2RR7VkzvbjXHArMX3gNw5XskFfb0isC9nGeflW7RcLI30nwze1QOjVgBEOpTlPMZMKmXXB
bX0afTxnVJizSpNoz02lCk6EzLQURuF4oo8dpqEwjdPT70sgpt0HINq6tNZU5dSOwd9e1maCjbR0
v9hlb+jVWrzH45u5eUqdWbn34za/8P6gwVNh6koLafgybBawFhg33VdG1Za2z5J8hJTBNW9LQmc1
ps19c3Sn0nQYVJkX1BhO5z7RSOIQ//MfaF2E74lf3fTWZhjcDOwx2BTSDwjJwM/j3KhGg6QfHImx
qcM8dekSx8Wt5+SP7pPxaasck0qLvQ9T338PHB+KM0RHLYq+3IeiIrftfil2KYVquRXJWAkfYB2e
vTkVrweSSXD27SiZtsPoefQgjb9FRqXJWbsuNtIknzRZs33042sT4+N0uuwYQF3JxecW6Hnqt2xi
zoGHCacTi+izZfI/BL1hKtFX088DyxqbgIwIchUw6e0atjrwcCY7gQ9wv7cZeGYhzw3GW8U355oR
pDQMPYi+edvv3T1a5b+2wNpmJnJDEUTteJbEsUllXimqPCU1Bto+EsHuKxHKxmFRqUXhSwSwHqDI
zA1p6G9izQPorXfoPhUzKm5233C/HKQzgA2ifFayrxdM0nc+a+ROJ5SbydkZEeundWT8/DdjapaP
Yl9ols7pVayn8Yc0GPT8cbk60Ikmj2eRJ0R9FORLZu9XGEZMNg9p+5DdbBIf6ZW/zcl0TEiqh8QC
MIaOiMUQflSgO/pwxsH1NPY7exW+d7XPT1kWW7AUlLVwn3/8lnrxz8iT+02f0PPCNNaQh57x96hh
9zwhkRK74wP9jrz8ByjMO3I8+TGH1g0UOHyHX7UnEOJkPoNrzU5rDnLb4P2BaxYQfCQd1irONawO
FjSZeWFaxrjsAG/rIOUfHmBbxAhUBwj7rhm3JHaCX8crZjiT2w4yaRZQp0lYVXn7a/2feo2gFkM+
PbBgSvPtdReq5cyguCoaEwX50ZHm20fYvkGmgWlR+EH/6FPGn5UJyNG3sTV2FIOO1sJLvmohGgg6
tvG1AJi0m4DgAP/updNXCWXY3GI8NM/O7cP/6yExkks2uORjFkpgpJPvKK5DxoefxvRXUqYyS93Y
9TyXdtZCXYufo/QVNK90aFmC0DDlHFnMnm1EbC0el+j5u0kDg2nY08LGJnPOmP8Gve3pVAigndVU
c/Ra/S7IOof1GEGxnHN9strxFqvuSdvSJNPbacXTFXj8kjM0M/65twTNcVh7nX8lNR8SRZVfo+hy
aBF/BJRG0nkdRn0z+txA6rIuShK9reXWi/9C2ovYS5B03E4fCAhS3aFxeNucsZmUve18vs9frL3j
2cPG6ATCQ1NV5yGK8GguSAhj6qq/UkI8WIpMYpJwc89f33NVwdiJ9V6iqRE/Ae13nmkIzy1WPg6W
Yxujwd9OvJrBoYJFzA5hzi0vJBehuI8t6dcwjwrB1o8Aq+CEqvJ/0KvsQOz/fb951pT1CsLQDanh
uSrGK3sxgyebQvbysiPUeDpuMs8Y6AE7LrTpPnBN2nMzzc/ka3pBuK8XQdbdA5rY9Mp8vFKzmfBN
z8IlGE8gaRFkr0aMPu1KRBpfw4393aIpEkUcuvlXXEl6ZbW+InT4eltF7uFxLu2WmodcP7Iwhch0
aa6xhqxCjGO/iNMy+05xNXOOVpd4aYEU/EtuOLdsabeOd9PatsJyakheFbUw+YmpBvxtffZckNaE
GK5ZknYnJTHXO6pOHx72rEG05JqCwB/OwIJgWb73l3C9uOk/m2oiM2GiBtzanXyAoFBgC7VWZFGL
hSYZMvpXhbZtuDQHusU8Be3MhOrwM2G7Tgb4+H9tIN8V7M+S1jmgVb7MBSD8cK0SsmfHXEkGEWdF
yVOJpCMRd58bcuG9a0Z6XwA09KJ3QUZve/uS6DaPE5PCRsenArXkXSCTAALHlyUv4NqE3gju+6+m
d+UYr39ipEHK0FYgp2/QrehM910fyAdSUHJGOm26tElbUVYt1BnLUZmxyoot3NTBuVDGgsLgGauo
FHnj+MgflQrDiNytE1bsajAZ/lQRdZcFHdqez637KZb0KO5ynHE3+W0UXD3nnLgoDlv9tvp0Buqm
XYuMFHSiTZVRfSwBMiyunDq2cJ2ARA0/sfIGCLFv5XwNa79dCNFHG0UtGIF3r7oQ848dP3e94T1M
JfIBhU6BLUZW9c+7w/4R9RxBEHyCfFmoa8G7geRMJrubF1UWR6NW1LgQGwQsv842H23pCOJU/Kaa
79hC6q/7TLOJK7EoCjFaxgpscCefmc+4JJJBGyiI0U1hp2zjm7For8T3yyPH4sXCf5K6WdCYFHIv
QRmUeqa5X15TIyEUV4AFrd8p+cMZ++2zmEwP9KthT8R25ZiHzBDqEsRI2+EEJFky4dcdsf08gUdk
oRZaKjLdwo86p7jHledaxpqfQTCzHQ//sVNutkrYDurFUfeS8gU3ZRXVdnmtZh/PE3MxAK8A1f9K
2WJ9sBQqv+sdaQQZ446x3N31yCyixyK7c9LK3E4RpUORcf9g5fQk/fJJIMlQDhQf8ILGQgDj5j1t
Pxb4Ffp6zXx/+ngLcVe+X8avQSTfa0UdnIJc6DJiyWKu9xwMErCTojJ+rHNR2pzL9LHWuQXoi5c/
Pr6c+yoqWGlIXz8izmKdlsvyhxwD5mttXbJ2E9tmcBj0ZzwQvfJokQOVAG+bM9tv8q9Up1wIr2r7
Hern5is9XqmulZq4nzDsAdWZI7ddWMiE2NiSPqvqz3JNn9gzvomGEIkKdEXUpUoLT51XJLpx40en
nJ6niH3F6mc11jlYRKUpliSTzf5XDiiwuWeav1BbMj7TLhmPHQ0feIf4qDsow4A9xqLf8HArsqKf
CSqvr8U3W1VfxF4MrddD8Q9hKhOq5YaOHoTEFEd5YL4DNLt0ikDFGPDf7DVOws+DBQRnztA19Jro
FfWrQchN+wdcJYf2qKeo99AqqV2PLV8MMr2cI9v/0EaCfPpzemtkySX2JNblwkiD83JkMRlqzShr
R2RNgC4OaLg6/+erh1IupIzaO7O1j8qU5q3FiOyRmt/12Z+WP4zxhoxdhTeL5SJwKV01Y2PaXPUg
FKAIf8EYbE5qoTGsII8+rYS6sLP0OcgMl2RwlfC2YN3AvBasM6v082lkslUrUZuZDwUXuRr5WJNo
wG2qME45DCS+0PTrLHsHjK+p8iOwdsBS1v75nmcmQl/96hjQiuLeLAuFUIL1PxxeiNXuhehWhXdK
vk2iDbYLcmHoUMmvHB7c2/a+ZAxwkJF+gSgtLESirqognBHEtNSFcNer1rsPcZE+iNdwD7Ra3u7z
wH+KLA9fADoBUA3lswGHJQkiHSImhCR2evtRcJgz7jN4EVF40vXjjF3qQXOGuMqlMbsfGoN7EPNe
aACICGZYMIOYOzo5WoNqUEksFaKdSXNihmcCbA5rFzEWn0WqM1rARUAv9HvYPoivkVJZEwoWZ75S
h9W1Mlu7+/3fRX7RNyCmaqscIjwoZZJZ3Bg+Z1MhYE+lXRwHTNhLYkS73+Jm7cWa+Ps178+jm9Kq
ubSyfKJ7Oy9Bic5dNcd+UpDugPc2eB3zJAH1tYpdz1IrYb4VA5eti+UB5JskJ7py2KPcLOuERjKJ
wn2+as54JQMWoF5C3ua9Xipo2nFlCVV/VzwzwEHhaafYWu2QONKlvTJKDW7nmn9mxVuhkCKuWbgZ
ehu6n/7PxJX2AupkNhrynQylqC+cvwHP5pxzZqaN8DBfAlXZuz6A+/OjAZsXJYDYZ1TLZGKsLgoA
fux6t/0q5Tzl48MqDt4qNbx4Zf1tZKnRgMQxuyji/DyP7UlnnW1MAz7i7YSYXhLUYg60pUYxrgQb
lqZVahXxLjUAj7/NV1uEYZsYYsdu59NvMk0ogMOa3eZKNCvxpLgUGIn8XAUb4NaPwRoFP+mYq4yw
OI0UIpVUEnSb8q6Efu0W4dhlPNd1mgvt5CDfKuHZzroTVQ+wNwUZxnf8CJJstMPz6BCLtMVULYJ1
VlyRbtcxSPtierD6fdY3fZKXxdrRZoOPeB8ze/0yzIdToiiKuJ80sCv2hv3rvOaW9zDX0pGrStXO
tc4261aJLWv9JHTbav2X/XBGEUpS+cuiZt5SpMgUJYzTazLrESikaJsrVyNgWgX/XPTuMmBNVd1q
PGdWVAhZQK/32zQ/iKui1W5k3MU/rRc50n6osBTluTLy7MF4TQSz/jPziqX7EPmz/qnhktKiEPCF
JIwexSG+4OntOxat9mE6Gadk9uR2+P7tmmp8wKKmT1lGgymE1L26x3teWiPDx4+UCG0tm5JBWLcZ
SM0nmwHVemp6PLDErMYKtaWaD6V+6BQgTnJWLsAk0UvAZqD5fo2udxPhIPH33onmseJjPEIySry9
veaE0GpLuaB/B4TchT0dHY+mC4Zgv14+qUZgmZZ1Uqhk7tpl9ta23f5QmIvXBx3J1XrQBeKvGo9i
tJ4rCO9g8gQJovxu0Azv/KucvgRYKxMmZAGUFi3Ziz8tFHKpN0+WB9aJRsxjYp33ltfyEloPlJTy
n06AScS3Udpcn1RNLNn5UXnfVpuzLz9Fmy0wwVicQw/GsLHwEX3drvV29XSRWjLeT4GF/h9ciYS2
cVjxWeLyOlivrFzyGsPo5TIlaB6gHmBS5XUbDqpGBekaUrh+AY+phivdHlFc3y5d2AWxGvD5+XkY
okMATB+jC2dxB4XJ2JVYcivOmlyebpZm6Myy/tz4D1AuoQ0HXXvXRLAH01N/BzBb/RjF0+6qITd3
lAkCnDZdBoOA+gICezouAkxR9zSO9czBNf9uOlMIhLktlse5Iuvh99nf2WfC+a8htb1jhDtwfq0l
uOYWdmzxmhOTdxGasplTmI6rTxj8zobpUzqNxVMXbtV95Vp7Pmfkfw7rGQRo4sKdhXH2Qmph0WL5
8vttrcWUE+uEfs3cuTDf/og1N5+uERxnlVKCOjsu04Vxylhweu1U8ZhtrHb6PIPf14Q+TM11miB9
GuBEmWYeLhOSvB0vO5cZ/Rcg12V8MSbOhVwVZPNoBAHiRNMB9krHu15ywIyPpACFlIWIto2TfbDg
CcIjnCZBEBQmJThaCdZ2d9/oDszcDFv5tWPUmtlBe0eAC+m1GzLFlzC7rvu5dKRYoJUqme6XiiZM
Pjjzq3pW9ZC/KQKPijnqrlWNwuD8Ub5QRV6VwVFJkYasN4yc2vCss/30qC3WHNBh+s09O/dJbGb3
c29gTbEHuJ7rum+C62RB8/QOgmdaAvhopxbk5KdsB+6CCBi4SOZ1OER5w93XpbDMYeMTGohn5XRD
qkMvkYnViIltTqjZVOWny/AjBdjRJIxvXpflAa7WxK4cNgoyVz1Kfl6FMcweC9oE0S4wpKGVQqqL
HxMzEc0cJs+cbbVF2kPJFzAcz/e9OBRaWAoUhCqYbtYdpFzozzOMlEke3UPwXOoUI4cpR5ihky3v
rnIk7qH7d0q4CNk6+nM+t3ozQl9o2CYSBjRkxwCjSSjIiOV3d9MPP3t+nYpjNWAFHrUHsLpPMbZY
uXn8WLNFDSij3FQJSkec9IKMsrUBcfnVOrJsJlyuJpLi42icBBcjBqpRyyotHmA1vXzujMtXF8QJ
w+2OKouAXHdha+CQYnMO7fch66yILb6x03PlKkLr/XoZ79F1rcLNK06PAIo11tsqRyoVWCvm+rGB
45sHI3+5b0dfnpYJYJD0hYhEB/9hy4IZhMLIYf2RyE+2WnB/z5vPAhEt5jeEoKF+XNk0Ge5JXJ79
jxxuek2a6Wb0sJhM52siyXGgDkGGf8bXDoELLhAny15OeHTjFHvdUlJ0As5V4/FEBbskSC+lZsz+
fzL+rA99+jbGTz/FboDstcU/oYKaJETBF/m2MAMV/oyopQIbfw9yHhhPuBEnn0iTnGjHt5lpmEJP
1Q4AsTWUSkqvpZaFgvQziDhOa/sofJnUTW3o+OWOSSJZuZ0x4I8C1OOdjhGtkPCCgCTEAPECN/Wf
vt38XPoWmA1bSDMocoqp6Z/0ZcZGnJjEi1q0Yvtj3/nQZFB7u8l53p1Regjv6CjhjwPnRPipFNXd
2Ia0n83pEiQslEc7K/QjxjVhgISZXdcYR0JbYivzPAzw+/G65Zv22HIn7HbZ2kMT1kwTh//uDpiX
foxFpkJGc20vV8xPQWgjrXlHHtsW8hDzdGXcNb1vUYAwOGRX+um+mrClu8vzIQaO7mFEdexvrw6n
KGhhnP69S/IK0OfVeu7FrkQYgFFp441hM/1IVTyv7OZgekDizPfAfiidjCwGz+sGweB1HudfRBOo
Rk0WwhgXFRpPXs2Tus8+D+MeJC85bIu+vNqP+iOPKunLqhKvvjI0MCTX84ylMooBnv4HVv9DrJZ8
eWaufyzcc1zQqLpI18bUzbWY27XO9Gc2gJIFe18RlktvwHNdyydBXVSNPqGTn+jX3tL3RCek+ykl
qwf8YGY3jDuYxCzcQpnFdtli1X6oioZN0vX3AjuMDY+Shztr+vBRdX+uWehpDqfZ9Edvns5BhSgZ
eKXz78Nw7bQWzsfxVCKKuX8s/zHx1h4c/RqYhFRpjiQtochY77ijbBW3qQQggMAJBxR5Z6qDN/re
KO7LRwqMceQLhCWgLSmXTReRswmSRIdtUKyRH9Bi1hhzTkQIVI/jCrelxoAnAZs4qaU0lT3sf3UH
LhWqhzHPE9M0xdL4jlADnoJWeGYWY1kJdQWRuvYvnLRFhJPGV5PDXntx6jqpKHqPQtO00v+yCbT6
1LRc+KEPrTzW5HO1VH/Gdc1OYmPhbrX+6qik37DFgCzSyebhMWQsMQoKHSnwnqRzoqEmU9GaHV/r
+bmLPCFvDjZy5mVo+jL/Upf783kO4qUM5D/EFspa8A2x84k8zN2LATE/qACfSy6Kl+eiK9AIzSWN
umg3Pe/KzbfB7219wPYzGtO6m2bBsHWCRsqI+zdYSoiQydaBNfW+/rdYvOE8nXrt7w7eCRGG/umT
PkuMwAByycK0CRRMV+wEorrqzTm/ZvlsurwwolxQNDywx6trAerufSsffEEYbYZjpCYEFW+KgUQc
azJ0KCmKzTj6g/2ztK6WbPv9vm4s/wNC6Ou+L3V5h3Eq8OzF6eduUAzP13kqjImfm4HAWboPYuq/
uNUs0nBjYNDlFibFdJVU32zUx9I2x787a21NURsP8p2FdvmJwGPlIS2LJoT3N3E7CR+M/CI4AQG1
Ab22OXFt6LPZRrpoXDHSo0f7K1x8+mteDKs/ixunYdPMh9PLya7BKB2mSWgYy6axnI74qCs5nb5x
atT4Kub3hjs0kf4Zq90iA0VXaj1ZguaGiJUnMK0SOhm3fzsfzzM1BuHhmxpc2Q20LaDBGERmdf6H
FT/w7jwHhUySQntGuo/BxI8iLusW58znJT0IlVzI5x5prFZFYcp00i3jYUrOHf8ExzjKlMOukoJ3
fAyLQQs9ZxLNefprRDH4CV+4Z6yWSSAaPaqXUwF3h/c/cf35ibHoJoQY2g/AJ3NDW7pXgjrsjVXV
yHNAJ3+zM/WbJE2NCe5/rDU0hhMZK0npiP37gwXTfu7Uh1tCXw2VO4py04gy1wRyqQyzhAhmrvsu
sPP0V0wjkc0kHfV3Tm7P5at7T6lLv6/lg5eb3TeBnkeEs05bFGwBM0dpLNH1utb9uX2x9NzxJEi3
NFV7Z5UzY7Sn34kvRr1f0amDTdTxjxKq+x8ghfhE0cH1++JKePOD4eHwVDZvIgCZ7rfCmBy5d1cQ
7yDkAKx6nV9krSMhIvutT/y7hSbslk3icm+RTFUOefhdMShY+5WOfMWj/WKyoyOId0lqC4PYe3tv
9SmWSt3FEnbKlzdkdwistxtYCfjrIlnw3YE4UyDpFQLEBXvS+kp+KaHhl7g+ez2aagaSwci365rU
tBn8CSMxz2ppy9F0rDw8fshDesiZ5SJqs3BDwMtDOIuqc8GB6505GyxCBxLUg0/O3xpeQ2TJULzL
8haDibW0zXfUcXlyR/f3MSWaZUYfDmik48snQPd5B5NomwWY6DHsrsRwoRhH7w/MgNP1cw1EVa+W
J0xYb/ynOFIFO0Fg5Pib6tHcPSFRu2EQPCpIFjTqUUWP1vQ1wdv9dfaQ6QMrJwaVHAGbJh9bvvs2
pQNDxBLDd84XOVOmK1CyeQ9skfpqnZuIzRqrzrzYihPxhhmd2sHAqKlI6jy34aVpbHz2MXRsJkIM
ZXELbBT+WYe0O5NvvYybyFlH1koCxvd3HLGGgzpXbZhBQ6Mg1j4su4Axjd/8FsFe05f5X8jyBl1N
eDPrDS/ArGvZNk3OjAR5n833pPIU1F7y5ciaEE3JINhNZDcLWhvt3uHPyynZdRXzeEa/77ZKXC40
AWMN++C4nHVFC7dzqBayHLxlx1ytGSC5y9EgGGGg+DrwkFpy3e1GWQVgsV+0HCkuRg0Kf8jsVX4j
+WU4rCdjCcbUTALS1qSBFMKTafNG3429xON7rngOrNAuKYEhOqgcQP4hjZziX2r6yPyQ0klDWp0t
Pe+OLiPS6vFUdDnZjw9w9tBzooNOY8cde/9Kq4zUUe/UVgJU9rYRD93TkBLnwU3sc/wsEJh+G1uI
FueMCY4oOVfXvJPaJOreqzS9r1g9hFnmsTHxHhc48ydQHfH9tATB7b2EyUcoWW7fLWII7f/yhwC7
9lFkvJS+SFaLiDKHUMT/+twRtsvfFfnGp9cXxfZJvWKVXQN+ihj+IbSTMAQCNZJ7+seuCJNdgKpO
YdGgVn/8s71x/wmnewMT0zKaA+oHFYD9EODM/fhFQqSG0jFRTW3WnLBFC95VMWw3o0PGFxRLGeFz
Lr/SRX3HliZXC/pfoXyIG9rS1Fo1q4zwrWgqnpkSfbjHOJhsYMZca/mTf7jWRmxf2y6/URRLeY00
qhmftDr8GtHPKd3rYjK6/YnpgduWjGLRNdUWkcamRxnU6u1pYzHzGF0yBJdtOfMaWLQY3SshZma1
0XyN0q7Z568jxvZJEWD8ruigxq+UrIZqijjlMvYfG/NhIJfAFQQ2WNK+xo/jd01yowNhlZnd2NUO
v0GNRvS1tkzb7lfjzb1GZAvrYgUar6fSGbD4NKYoo+BiJGgpUosVBL/os5eDb/n9CSJbw2TXs6ww
wYCYE13/oJhoaKCH7Sh0RKo6x+FwfqSHCFzxfJTr4GQlG2pbjUUo8SKyKVmRBwtu04nzclsBuk/8
USPxqaQtwHaenxpW4amYcLW2t0UkKURYQT/myp1jdY4PEt9nyeEDaBpP/Tc3mNR68lbieQzgFD6E
C2rJzgQJTBrp6LPppppbH+luGdJTZ/3BMBrnJ2P/wAsKybJCUnf9PgEI4MP1FANTtL+GRGtIhT13
4uU/5A/LvIVLO6NuHyKjKmtlg7FlCaAZdTWfAEfCu1MPfamOB5lE1uKFIAKTfje2OlMQzaFDiEfj
yqPUn+DT1wOjlseR9PtRi6ZoCinX+ATAWPBgRPwQLXzommqSSXiJS7nG8G2z7ff2EEVE+8abRrS9
VHrW0EAl2we3xpYK9ZCirqY4YvtXMHwubg0+uqk5hSoySod4/KxIBgu0zWWtMR4u53/e4batZrVU
6uqnVxN1lSSpSzwflYsPaoJvuEcgcs+FBzGV+P4w0w9ym1fpm64m6YE+74B1VGbfwwk015h5hzmP
KlBepip/poy2L20j0NJ5ZRPYNStAW1he/adLuKE2lkhylZFTp1aZ8L3ZuU6srvs4IMh5JHc2JGKK
qRTvNOt+dMTsqE4EW2kCaIzrDOLOYzfzWV/xvQOUS1RtU2GYFXKvErD2XGfV09gaSauakCTufzPk
r0mpIOHmqHtNz/Do3nUJDPZOpjNAD8BS8o+euyUp97r6R1cNL+rtbR/wEKuo5Q8tqv1UlTya7X8k
VykB6VYAtBrmT2B87SPA9grJFgpvety+Yy+lY1LNzkWs1FJTacEsoqpCqAHjSbAi08n6VnWkhA9O
gH6zws9C+0+B48hMe/6AM6NwkjNr4IHxEkyROtfNgGxSp0FipHb4CSIG6mgLxNNfxXdh01vJO1nH
ZZs9sap2/FzseJqXBvGn1PNX8Q348DdQpxGf6mORCL4QR8ZxyV9yF4ndhwNVi89rKpXhkHHSe8kX
sAz6FePTMJZtg6KoQ2z1ov/ObI59YwICP8HXYw+4zaUSRsRnKt6R7utw1J/3ijULLHL/vOTWJxTq
FnnFOIsWqY2UM1Mi0eYZ7JcJjyk6PyDUhwzCoTQlLRXlw/mKzB4iTGwZc6chZQgXWMrIvP37SuHV
+BxKgeSAobdcqKElAkfZKub9sQawFfcWodX5gMcbcT8h31Vj4Cc/UfwObtSXdkTAgVZ063hKBAo0
dwl286orxQxShCU3NWK3cx5f38bgnf4E3eC+YEVjYpAOAekWUdcNZGzgF5UbvQQqbHNLHQHiZgyb
5YCDW9IOGNBaok6x1cVTIsyIdMcoNfP+HyUDhqEGTLqaTtcwrm9E6fbB4TIVxMjJVRD3P4AoXXHA
LhNt/KSXE1e3G2IaPNTIlr0P+IK8P32/oEPvOpdFBIEElHhOUM6u+BybS59DpDogzTasbz9hujkc
broudi7IZ/w9BGBhnmEdcebh5RRLFcALvXIJVyMxq2nDyIYk+AMLj8ybNPVa98hU5Ytii7qzWz2B
F1MuysOEvojKNrn9ehGzBgEZQaRxFT1bvVZO1CQJD5vdNYEOWhKqAiAIC5Vzzjm688e/JPw+TroI
8d0cCjxBQGTp5CM/pzEzP6Tf/m+FZXVaU4rMktL1kebZPOCoxjlUYNoMrFKSeXE2A5XyM+1sNSYw
KBdg3HmrGof3RaZVqRwdhLROTCDLypahbkjJxlFxjT6aNX1jSGHv2HLu7illVHCbmzCPRNRhGE+T
VNXvRnsRzTBfNLc+dTLDPMD85AdSY2lFakspfzrdAZrzH/0mg6/B8VmTQwrRkWZKT3ZlUFYkvbXA
D5Ye5z/a8jLrU9sviOy/0llf2t2mBaohUT7a6RFkSjYTbz60RdoBvviUnzPWvQuRw2pJ9LNzboh/
63JKb86xepQ4JBp7MboGNS3PI34ADswu5cv/LMZr/lL3ApZp/+7YyhaZ0CBmYufbRAlck1Nlv1s/
Nz+v7NXzFdHsf0Wv/1X4BNjndAfg+OIbrdWJOFO8cXD42OFagl8pvk5AMYnKMIdPGGbgxHNzf+4m
3+Z+x7BxwgKUPGchZD2xM6R+vXFfITH87Vn/x7hi4xE7rNw5NF+7I9dg3MsK6n0bLlJ84hvPLvgY
vbfiGtBKhJgO23Gc5f1SAxFHd+b1ffdrQECJi+I5qUQrnwdGb6HIguhI1QZeXNi+73YOFDk48AKP
+NFYI06yCQDNQuaL1glOMhpkvEZDyG/y0B+rfn6AAsRqNVrRGxd083x+XRZTsFmgIJ5iwnk1uRwG
wOXgzv6zC1sFR0XvVbswoqstgLEq06JbWWqmBvtxyBxb9VFoLv6rxnZpyU+3m3y419L3xJX5gfp0
VjCeyLmKksz2lNgqZPaPT4PiAoo98GEKf+lqlOxPjOkPcWGgj4yo+YnoZRfKAU34LF/cskYLc3G3
bqiVtmcHf567Iw5XaA+UO7S1jWeUStQSuHAcrvdVMTSMwSQ6OxyH/ehrScMNirAIOKqXAcQFZujD
XZyYKAPKEFEIq2DzQhuBbTLa2on9b57HI7LeqlaJkDpfAtwYQoJpGZvK0LGqcNswQnRxM9c3NHs0
TH02ZPT5h8so4tiyJsBuqlkUR1aIymtzbX8kBTTonMuIVt6eRwdgk5csBOI3q7ELWFbgd99oFPO2
uf2XWhHlDOPFdBuH5Yf2n19aD9LJa5Qhd5brg+Ge81kzKI99PfJBt4QypGQ3oVvv7eF71EmmkN5J
DfyBGYgEo17YVzXPlXgQLsphO9kmg7aFwwN9GASS8vlyad2Gua+k+Ta14rCwTL84UR8b38N1vKMz
7Xo26vUU+IOEvf+paGCglmA1B9/1FErlpUf+qyu3TwhaPi01kOrbtz+mouhAjYFOaobEEeO5WJn8
A7LK56sVLwEouXTbxmuAtCpOFj41pEAA4U5jmIPk9nF1eAgaaAvEDcb37ZB8yLO6BcdE3ij7EEw1
ncJcKjNDy+iol6XYJehZo1348F5dWutbCIzToSxIfreG2o5SCldUMfwUweKdr29pJzHNvn8e3aP1
F6H5s8zHe5J2OpCeqp03J/1zduRUfhdVG/BaGaxXGhXj4qNsdB3TNiXqpjVp0gO2zr5k/GvOzXA5
cvHqR5O9y6NwlTeR7VZlYDmdYZ/ERlZv7QemHDVvsPjRfax/dIWjMS8l7KKAcYG0wtV0Ay3Z/RCP
YoIkFcMFAkBa8bnW+GhjKGIUUPO5BgPzI3mgEFaEolkXW0VJjII3LB9D4N5K1dPomzl+SJALkhyI
1H58J5wR/KyL4tf91KY9BNU11Wes8gtsmpDsIAwe6XorG7XZTdTK2NKw8Dz2QtRCq4gZrEtbDF6l
m9665U0Tuhwse/Op6KRvqMeRcqapU3EvSC9mXIPB5MoqgM8JkATAxVL+gkMcd6VhvnUMDVBIQGvC
RqtJ4uyXmCNeQuzsbLY0Li7KPMXUBu/QNHKP4frgbLawKNaiMQ5S+2UoFk7HDIg/EUtVF76/xbF5
WqCPsQtkF6I7s7i5O8RxhNnamr9gMd6H9tahRSn2mPML9KMlg4WAkJ03QJkpQI76y6EbYcNb1po2
9GiAaTwOiqBq8iGYzWlEfQ3ap2rHVMsTU1G6jc9pzzGQbtqFGRo9ZyTD5pnqHHBFi31Ypfs7Oqwu
FVf6DnhCp11Nr3OGC78LWGz5xdHjpp76AfJvOzKqfOFXacWqVM5EFQg/Z4Z2dyBnifeXR2UXKnUb
UEbQ0MO4z6giwMKKi/CVflrOBfXYZ1cFtzRey5nYfYygHhzCB8vW44HwVJC7uxyPeIqmbbOi3xDs
vpM+rTQs1y9kjlPGdzq9vWeQ+W2H16krehafWaiD0S3yi1Nu8fSeazDDHcaBGeAU319FiC88oUem
tal5eihi7qImko4d62HxPVrnEPxLQePiVb8dqFwunIaM2DL4XnxZppbvwDPhZMbtiTh18VBZK/12
D53sIpCH7Ph5tCHbDVdBW+gRU9h2Ob+yQW3EG9tmw/CaaxpjU/o/7SU+gjB3YPPUjQHjdXsL8gVx
/Y7plM7RCFbF1OGigI/IoKn2hyzm2j+yGkRNWYAXCcoS1je8olNbulslrI8TLaWvdW497VF3yCOr
fH3ElNnoyJC1Z2VfLNdBE2ssksdXVXXojtd7R1S/5rhSTCWvh0QKpcIRGHlNetIHfsjgca2oSdN9
Byp6acXDOSwnqJ+/EFrQty6rAOXpUvGJkzaMJfvwhmgsbWQKyesUOWKkwigME7Pch0z3uFXLMzfn
RoHDxmjpzuhW1L9+CnLckbbfNWY0FtfhoYA4yFQz23XGANyEnTOa+L/WyGdrqgGKZiJEG2gPWJmY
JDXRX0txIl8kApgx9ldKOplYwwugHAn/Gf/wDuCcXp5GBkUtGASpe/VvlXQKl2QbmZ80fVkuBAqk
xUyYYdiawUattw+t/ej/qEb+m1mXUFFnzPFyhSxWXTSmuHCoVJlkpilzd/nZBH2psMkpKWZ9hfbm
UsluMxJW3Q2Psu1hqg12VVdh65M8XxUCbWX0btyRh6Oy54r/4plIC2SqKHgcSxgP0zyyHFej9RhJ
x0CX0ptIooQLsvcvenxSc37wfAAELWb1gFSUY4DKnIWKQIBQsYEcJf8RUQQR1sa9DdeZuT2tVu8I
S8oXg+M2b2mVdm8RCTIXf4XJw3KNrzzkM435fV6JT9LcVVePWDz5o3Z+FsH/fZ9Wf4AXG7xQetIg
7L6ayB0ahQM18m+Abm2qVgucTYDg/p8GePCj/E4XyqGpz6ajwdUGtRmPnlJSWrL4/sbt6gzyJoZG
txVYtrnOmuhywQAO/J1xmRcH5blqjua5j6tgd8UUq7/rJJy2SBYTNeKupRxgFRB10tSO3g01v0TA
cIQiIAlBj5CzpbOsqlU703DQj46VykZe2Chyr36/gLoNy3A6pshbx/BgnztwD54oBJFkr63x+YuG
mDrgd3FsBJwQNvdDIAEWpvUZ2q4zY+2zyXGhd+pTMQv6YAJNgcy5NzQWC2jyl6lynA2ifeI5ZCnu
eLu5lov/bFyoxTVU5UZE7DHZRTPw/yQR1qx95VSnt+JlFno3kBC2WHN0ZT1qId9Ojiu3upJI21Fx
3AbOFA99ASrAv2pmZnomROgmT/hJKklOFxgFDrCPkQekSbG10HHASlvIhE1Sh8O69/cS48yF7VUI
AxHiYgzo5iJBAFuAg1oi5TJtm/1hlE2g70UCFe9j6YQ+klHZ3jY/ZFvyI2/oT9P4CIi6gYFFrB6J
hg+NFwGGh+/ZC1XuyNeWkkgn+OTqU1TxUkWSb/tnc/sQy7sb+iOkuHaB8DRY2uZ1qMk9NCVvBjV0
YM+cpqHgefN3jTrPdz0Fxd/KMa7vSevchLro+dxAjaSx6EqUNlvk/0rqvwSL7B/+RgwAtZR9l700
5MAu8KTqYH30UXATEl1lFvXptHtMTe0XDdAxD/xXT61pCeJHBNgA7oUkNRmd9gQtZSGhz6FPX3Yv
GH6dKxMo7NFuV5Duz2pfVtExuQkD5J5sdezi1UoJCPiIT0ZpuAPgZ9iSbZ5pyTvDhT0p8ZipTTPc
XzEuE5/fR/+0gDZzOxvG0efVf4+MSiEO4P0eiCbYGSumu9pSGGSEO+fTaiT9I10qbxZskEr9+qXP
pXeOHM+WDmlMasIs2kIVYMoQiNZ0ae9npQu53iTF/iswEvuiodt80uxDdeTaElF0mbOKXn+BRhWt
LEmbvu1jTQ6VT00L75YtPzPKxitcV05eGGgeSNYRK7r6rktyl+Kc0mBoigDgzqcs7RZ33zQvo4M+
DBn46eDVJVG+rzuk/UPSVNEVUr0dmHmwrEz4QHSLBvpD1bqEZX2G4FDzbhX3lZJSCFjeageD3VEg
plaPqZrnCC71XlJ4wXZnuq0cMo5gcA7HBYBxSnO4s5WadSA9DIQqceWW8citcczlc9HHSImNPJK0
yxB6lMSS2bYDeSZaLQTLVy+K3Cn9skGP1trlVjinDSyC5kh8L2rtTy/bGDTjlqJXMhddeOdW6HSm
hLBOIzeOj4pPxFBy6NBRVFDJ3x+/vGMMht2s9aE6oHiYe+3l8XwZzSEmPGVQNPlZ9WpJv8JkHsVD
r4p+llOZTBtcorKO/RcCpo/brftqseuzppahiFg6JfWygNmEC92FU/fAb4yqeVASBKbApw0boYYi
0DW2dhHRti00SYmmbSYhWBOIMq7bfcsyNPK030k1SRpSbV2DW3xyI6M4YJaq/IvV8KZH4aFLlNAJ
euLqLMFOrM0Uo0oc/3F9PbfyY7JweD8+jYscysy8xDFVo5W3RG8GtX8Cmsz1gl3T3QaghNaRCOqa
uTo08/65MgAZr8z6Guu7+W0NS4DqNV4bwYAIC1xYHZj5FTzDLe0pz4GVIAkTFPX8/SPGDKDB+yGK
1wNyJWWhL1xTlKJ6hcl2KfxFym0MVHjf6LS617kH+bWmu1GlZ/DD6wHBxqB+HfAJ51yBxf140Bfu
H9+YHhBrSqiCtJiyEi6MwKEkv1q46FgWJlpMjLMS0+mDOSDUkVATccjOxZHvnNF87IBfQjh+RHju
EXtgtEYVzyhnGA/2oklvYxhg/g7qa7A6l7kP/ReX0JbDhr999ZaomuGfEK5TvLBOsAAyeSBl9wn1
Is9KQ+785PgG8vMmfssbRKezkpsmB/tiLyc5aZQ82k5eD4T2PinQ2uQ9Hy1pNTbNum+tvZljM3cF
hVxdUELIXS0746hatzi+c2NP2z8UICLHoTikWP+Sfu2d/sTweSxYLmJb9zbT6s2N1i51LguqzSo+
gQZp4v54As6eZkdPIoZXAgHeS8jS3+htyIDtgoq2nC/FN2aUPWctK+fAq0wrnD0xtJ7NQlFXRbsR
tUV82pHoxintut/BP3OAOaVc3KVbv3Q0BDtCqX1ueFz2g7eeMhs8dNVLIlKBH+OkCeDvrR1Qs12N
uNMGT/uMCSonFWYKmobgQF0CNTkAmz/5DkWC+ByMGqL9jw/fq4KkL4lKRZb/CwpPqFr+K/W1zuoG
3ioeRN49ysSSY6GpVeTOGHgIuQHpA1KKH/7L9f4EDk8vzjd/2qHU3La0AtGtmKwOSHPdQzZ0Bp0v
L6mxB+UAo0UmFZeQ1rmPv0/YAiVJc1KH7Ejuy9S5MzSiKFXGd8eNFOFt06Ku6qiMebVCwso54HSs
gwfZxPC77/b1uatdH9th8CkI4nML7Rtigbi0BHq3a2OHPioR7YyD8+QwARkP9yo6aWpGU7M3Czp8
L9V7+LJqYJ++c+IMrrs0DC7nWy7NMvv9N+ki8CiyQBGnI1A1Cpi3R5iHYYRujgRqJkjX5+6sPTP3
tyaabQ3nZizRbkYP/ugtn0TeVVgIAH3SSv3tlschywzF8whCZWeM9uSBIaeMoJ/Vuj96AXkgr9pm
NROmB1lFQyQQOMhuXD/2qbiEw/X4fsPZmMD/TxJqLdGF3CVOHOoeOZnSNtkkghgCxupwSUQkKlLL
UYK29Hc/A08wzamslGf1+sWw6E4XFPMenmh5eS07qPS9+5DV/hClY9Fi1Q9MKcW+VmoWnaTSpkAd
PuEw/KOQax3uVbFMhFG0jXw/X9kUsSL2yuKGaj4pu1EvT7MERBWBF0CGo5aPKuYjKR1Y0vJiTFwF
/fOmu1505gfc6Ke9BO25i4e/ie01jxCuP6AdGV2dFdWIvZWel4FPaav7ZO27nG9bvcZnguh4C90p
vyO/mASDNCVUWS9N3kWCe8QAWxu4TI0PMhrxeBTO24N8ULE2dVhfFUn/roh/MTSqgRZGqeJgPji5
TcIrjDCLpN3aDtXvCyMUySmICdfpb4T+XJKE4IU7LmSQae7IQYOKlS+R//54Tm11mOHu2+16QTnp
InMNt3VomvtC+u4Fvmp5/1Ubgv8qsC0BaqR4tElAamlKGsxO+l7bPZ2TVxGb3M3HgsTbrt97uUeh
AiCqKg0LoDL8AKqGmMDaXT2NtKPeokjMfVlcBYWwklT4l9uEllgKjuHx/XBZHf8u5lMuT+Cus450
kUCuPNpuBkewJLCUgWhtfS6AX9cJrXledcH/JGpnxUIqarX09elUuxNGB+ZoomTGwywkpa5sf29g
BAfq5LizIhg7YG97dd71IM3CyGwz1ycrLP/l0KAwtlPXlV6U7s3bOVAc/jx5zSmPVFbe4gjtgPg/
gX7AhZzEzm1aV+X9DMsle5HA3FeApClwAJayYF81YY2kUJ/lvFlTW1Uv53wCJlyI6Mw2HEdyoR4v
4z5PLJB5+DpLAdvzdk0PmPBPsatF92cy9SCNHFzHJgiP6tzwjSjetI5fFbLerbVNEEPxGKyWLnzp
T5cJi3fBCjI0eRhN2JDuXw6mEJhtbwYzfzZGsXSaAXihnQ/PcHTIhpAXlDMqK2XTnzyYSo6tVzX+
GOc0T5VLPaGT04KuLcHIVEpISJTjK/kCbGClhs8TpHBtD988GR4yLdh2Qt8Ht9AcurznezGAGCcy
zqNbMdWdB9Lj9rrHE73wYr42o/AnbNo4HOpHuJifHj0N2uHZLTLv9+A1AUNzRsTZPiAigd2EUp4a
YFt/WsVTihU3BS+po5sI6wsMkiGG/J0+Vlmapvl+b+6dAX7voBVniYkdnn5JBIEitYkhBQGZ89zG
1I0GD4cugBdqIHdowSlcLg1DXWSwhYLLnNOcX28sxbTWMOKn6aQ6XPvAdN7zBnAf8K/HoxpLfkNR
14D+YWJalClsLaiNwwxJTYD+IAHCRkwdkp9BCrrwHpGgT/MrJy8DMRd0phS8oZdnTrxOzQmqjqdC
p7a4uMBKXl+Yb2Tiao0gT22waNhhQnJjAUO0P+regbSyT62NBqJfPgU6wMHJaJvnaPOvPCV9gh1x
QnvYMEr2Qo4/9H8ZKGkFXjY/AHUzgI7z4ljEMMLbF/erBQaZKop+Ox/9zDI+TkuJzpW5vfIoF+MK
UxjnHDTqfSNSLkAEoOd4KW44G1Dqbvam76xBPRtOga57hOdeDuZ6YtQFOt0ZYmdCqnRx2VFNGZJ+
dbLs2tmMgZfFbNp3T2W86NsMJjrhBW65g4jHcITfIXTe509FG6S5RiKO+tc5yztsjFc/RT24YYhz
1IuLXTGjupqfm21xr/92AAuDBrQlgJavhK6i++4GQU7AHWdPfPuuGS4FZUR5E/ft/Oxn/4kmyLyq
Y2zS8vNTICWaTgafYvtAPRxZy7iaI7Rpp0Lee5li2Jq2gZ5QQDoCXx6exdbENXKeX0sySGhLPzT4
dDECiSmUYnpQ/ubNlVnn3HrteRU2ZftfDcnroDufG2L0MwaDrgkMmbBOX2PuwMGGAgFGk7LE6KtR
mZSy90lmP9/ge/t5YC3NlHSbpMPd8QJeuUa6xKYctIcQB7FGVC09U3s9bC9Afu3PBt1pxBkZagFw
19rB2+VIfRQUazyMcpJ2W+KLAmLq4RD0aFFlA5XWH+ZMoRyJGGaGu1O/VOgYCmw6m6qwjM3MoHLx
59PVNzB1Wd1+VGRZBbUTCPZOUL6vvrFD0o9qs8gFvgO9TQxeM61xQT0lUjGfGa767aogBmPEs1jw
2OenW4sA9z1Qr1taeTHaFDwbjrluzNrbUBGpCVsKCjVrQlubRRBjJHGDbRYAWvmdksxVHea9Bm+1
CtT4vBcTQt1Z0ZCLlABmC8l/8f24L+LJGX+EMw94HO7gAHVN+WegeukVqmD5nFtM3/jBnsNTNEnR
P07ZVGfUZJaywIlZDiAO/NLPCT4TxDm6DM3MZitpAGmH0THwzlRS9dSrrCuu9oGEUPNguNGKu4E0
iRY/EKuemaRssNlr2ZfOKz6rf0gYyra/aq/zhDm+DqrO7f6DYQS54OkDK8OZTlXNcG9R3v39+KB7
N4YVpB28j5VttjjHokhppRJcb/PwO4B+bnIIzV5NIluKNXoItOR8d3ZpU5TzAGSIfIu0u3LRCCd4
kac7iUg+oFKthzo5mUhxI7zPWe93jBBXu7Bu4QsjOSiYQwqXojeaRndMtwiPNOzmOni4TEi+9+n2
r67G8dq3lRe0LnZKzXPFBos76+DZQ8xcRydV5O4yoBeKyYAlbrlqzR35VBaCx1EQfLDgIhC4Woc5
FuPoUUx85LvYswPRIfHPTiD41Q+2hNvPvCQtqmmRul28enIawo29febppKoXfc8ALOk/UqWuCSoZ
UOYwmJD1nhsCoiqsgb10h8rTcd0fSQHNrhPhVmZ8b38MRuDC1JMXwP4HkCCjRSr4tWkJd8G9YEBG
kLVq7DV5xoof/eFwMw+cci2z4hC00k0QgqUU8IcZymM2H/Pdrioe5t9awBQ0jxCchcyLFZ7O5Asm
t+SI7s4nlx4KOvA7wKIBXEYN3fM3Ic5FK7FXZCIpwKBgA15EBlCjK9bVUR/zHzzDlhiyHDqDUwpS
3stnSWpSNHGebE3el/P4wiuPyNbfCTR24bB7P9VFZwKZzB9pS9annSwOjk/5FHt3FIwDVfJgeq/e
yTsDlBnt2k2HJmW0DeJud/Mc1XfuMT3/aciflfspfsZHEeGIL1H47s/UZehLLFhirz+8wbddOZNP
77ZbglFkH2gAQ9cKjYkpG7s579x1nTSirj3HoluTIxSzlq4ktVTXAhPAaYMcJk2qE16m2obmfDCh
5JKwSgeEQpikiwHc/fldIoaT5JamzMXcigci5h6Wx/WH4wxthXRD/HlgDZHWrfVzzSfMHkYEBrR3
+XTMUCpAXPIVlXyWjwc0qfsWY9fcudzXl+a7lGySVjrlRhfGRX1hwS7voLCIPq3jXgPYuV9r1s0a
+mCBzdl5YlIAErudY4KpwUXOnmX+1GtwgJI1rWEZ3EDc/cSLC7Cs06odQjh9DyVbiMHJWofSZnKH
dfHcshrNMMMndWRx2M/WFX3MP/4UU84DXm+LOoPURu4lOfQAUMo/3cCCynrUBeERNZrGIV+Jl/Uu
q/gOkevAqrkH2VyGSvhalTSf9ZhjhN+LKCHMEgHszZv+X64Q1qTQYwlCVPPBB68M4X2to9TL8XWa
zvQd+M/wmn19r9JEBdRSpf3RiZFYklintlUaA5qlYWm7fCBneB57vzrcnO4bIXRMyG0jwICv/giw
1rf7hk7WWSsrVdtuVoEmi+pnw9DKIkgl1RUiNA0dVVwkAp87s965RwrVE+5AxDfhmRvbVEDtPQ8S
d2HsuJs/dClJ3QqTNISFUGgcOm2dZ7/cznebC2J6lstHjqS85Xh2l5LbqAwm/c+6Ux0jLS/hVwMw
g/J1baFiOfFV/OuKnTbvE6yVNQ/PWvdOU93+5OA4o8cuboZztXAoBRiqWx6ayVlx2GAxlgaw11GY
AHJCDRwQmd7s6uEEfs+yeZRKmwMwwTfw1JsQN/hduoArbDwQT6a7J6vNfxi75mvepz0Dw104Kp3g
uhc/WRiaAp/EozhXOwjd6xubhO+aqhmkhwcc8nE5CcbxfvbVoBgTtxqZ6kpTGckDCKryi2gLkZNf
k3zr5lU6LnQaJz9NnmvKOUzCnV1JIF/A+F0c9SZp1aQsUNS+bKwlse9aEh53evfJ/0V5GOwCb2AW
qcHv4HRY0bxXvJRnbUZRgENgqfBDpmtT2sP1zdjPOCDqjdwe9ILY0Wy/1kGnYZ+VJnj3J9eLC5JB
B699jHhO2RCsJ4v20LTJNDgHs9pJlxphs4gKeT764j+q5tKuA8VDth8GitpwTDXtDnK95Mz8IYRG
4UkpcubXoJ+gh9L6hQAvq2IE3P/PboOQ5O7oBPJyskelooTzeL5rrUt+LFt0ON/sCyirV70rq31r
Cv7WDRZstm8a0gwbUEeONnmqnqw6uPCXo1C5nP7+ZAGjeEfOs2iTm3q94jEHDdsnV8d460EUu7VY
lF5tKAN5+8Marr1oSa4lwfQvRaAJvMbmTFItFHaaRq8yRJZDRzQprUkipYSl3hjwtuNyLD0Gi2VJ
79XXd1hcnk8zILW/SLTIniY89OXd9yt6M/1cy970wJ/zQ1X3GKZppvd7SbzTLmTswnbE3eA6B+HP
gJuJXxXhpeM5RfIb8nEjQYNDDEuVUd60FaC/dBuPMA59yr/sPJ6RJ48A7yHoKGpi6ZeVR53Az9U0
28Te/4d1YGJqTN38eSCNNHP8PCTnAlPBmfc9Ayc1AqeyiRjMGZrbgcV11zTZ5/pki2iGc9bt++zD
orZ32ctXZN7n+8mr2ZdWR4kVabSl/dA+z2pisaMgSNMP/fHt2UmF/Zt3MfEHjcRi9Y2ltdB0OEhr
VWO3eCKVLRxkBBCNKpGGRV/WpIOxiKgCBXq4xEjzHm5T9Y3iYiAlHBvilDDiDw/7BnjvTYQzPhK0
tO52GzZygWRrzYvN7CmtY8rGZCndrFYkoG6k3QwOOEZV2J/SQb6aT4lCb06pyttCzmmvvVzaQ7kI
4uRkaq+jrNEdTgmTWxXpM4/mwrbVq2O0uHUmShJfG499urTvudIp8gEiU3Higw0AOVJG8yLh6EAR
JUlSopZ5O48zj85v9M1id0IL4ZOPk5O8ZaddqODE7suVIcVl3hWVb8ST61MS2g+eVR2fyNOGe59/
jh3CZbsKaNmPe7tmPofMFYfUBRjPYlomei73bobW0/tHXS+ZI1GteN2tpLszO9aKlYQRr3vdmJlZ
1YOH4W3KBd1JhnoH1UUDTtYkumw/B2uIcn/WDkRuzbwP9CeXjybmfQj3DmhWDCge9brFIY/T9dT8
Ey6igdYCe2hhRTmPsYYFhvXkRWHhOuxsXqNXM/fVQbCkJrzKaTUX2OhGEmU1LJLi2TK6hYhT8YD7
dpz4CcEuPxlSTrzQ+MvCNCS+uf9ZMmJixGPT+2IVBuhvY1Uia+Drapdfgi5uSQnGSaVbHfVaNQeJ
+DvWuYZrlX82pO0+kSg1sGQTPrIpNW48hEP6YY94V5YWSjCKemHW96P/CZ36G6OGoe0DAhWXFG6p
TOkSaM0fQunT4HBZilrxGL+3Iubi8Y2lmpfGuKI124Bg9wUuDT5uAzFU7kY2f9NO+TGtvzcU5wUd
r0KYeY5pu1CKKfov0CJL0jSQhAqOMf8ssH7HdhZKcvGgTc29eEY+u1zoI7YaTF3cpc8FmBBETaFg
Q2xJcJes9L2WUoVvrcyQqZMYSsUSy9H/vodoNCr0OLEKMiWDR7a1w6Pl1wqSfsjtfvV3RDEG3vFD
AZbO4vJLwrNn38E0I/leGYuybbGRrDgZFenTZWiBOYDi7wNCBDODmigBKB8XZV9UmAZ7cc6RTT38
5/dqQi37Xq8tw2pKiHl/+6eK4EVmrEFn/jnMcj/09SBqyXs0FqBm/r3Pzx6p+2Q1Jp7CVOWO1Z3y
hROoZpgyW6fMT9OYjskGYW5mdzRrBEAD1RgUBkHbG5B4J5ZmsBBrB+b7gFVMe9fvoCHCEtHPgiR9
kpLWaz9lFwwcJAfATI48mT0qTjg051b8DOsM9qCuWVygsaOhzkPlvu7bVsB8qiRYJIOg3Vc2PyoX
ljWPv7UbNoMzZ71x4lxUBHXkU+Ghei8F8Y41W2+wtQo0XLBiqZLKnb+znzxwqzPt/HgNqTrAaVg+
zAyUFPmPMwPwMqtVw7oHCkcRDtu+wiOg2cHDcmy6MleyD3UWpaBlzUX+eoCyVeyGZx/88rQW7vos
6ZumijhXtNfLD5XqlrRObftzxWKQVMoJ/HQmH0VQi3H4Oo1GhZUs2eofIOL94L3yFGr1a/X14utu
9XQgRAYO/8LfOEmwsy4OhfShnlWUOqRQ8ncgvvmTlw3XE1G/h2eghcdnFEDyWxp5C4J0ggY24pBm
pnphPZ3U1T4ViUN9sL2Cii/CSXvCdi2+O/1q3RwpLGBxR8JrRm47rdSfYWMVZlzEzReKsW5EcaPA
nyXbH1to20v6vJ41BE4PIsFs2hl7n+mASyE3fN8CbEd4qb5cTDbDsEMjFrO2+5K0b0c1VuRnIpDy
FiCU/2NBVtdgZZBiK6CV4V+4yIR0Fcxw5+hHbWZNMHRMWvFhYBhNS9BvcZM7OjGgF2kf5xdZIESj
DZloBKDeRtlKLbMJELKXan+Y9g0KbIDBmvyKbvEZ6+mvZkQ+XjyIU2ig2sjxUaX/q106uYvd+okC
1RI5Vi3BC0XQrogP2HeGs/cBjQTritgy0hYc7RoxttpXfrlLGAZpG1qLRWfHWA2hIE8goYi1cKNT
+omqJZBqYnM3fuytJ0RWYSeCP217IM8D+fr1ZxcN+MwAYnwQm7M36q7TRhMV4X+bqd7UenEGQJ1H
xTY/cvjt0bgQY7hpFy8BhIj+tMBUH+YwJpGXDEBFTkG7c0n0P/sdissJsrPJacqzd5PIPtIC9NCC
FwLMHOHlPZ4cslfoGLw/8Zmvv80jgHBKwRtDrzRGUNZra6SuHT6rddFakDp9q5LZR9nklZAaHlFz
O47/7K1WAKUt/37UDk+AJ0YyI+gECR6oXLgrMUPIqBFZL4W2iqWnreVm0GGLkHK51qbxT0Ck0qYU
I4zYc/L4jvlaOOXfMf6+9X8+VStSAIl3IdCQeTc/4kNjO4ZEa2vzQdB05oxSlbvIurt7edizsX+8
+Xfl2Bt026truYd6X83KsjeyoB51e/WpYmAmgrIyT4u5JPQfUWO2n5ns1dx2A6MJn40pnXnaL9HD
UjtJTNTv5tYGXV5L1eXPVN+h+UArjScfS3lY3Z0jbu4wsoKT8gRdHxi2Ro3dvO+7lKGatbfnhh8u
v6UeG7m6pRe1pqTJTt7PYL5FQ2yh+v9d+8UgVdxi0z6MBkaOqd+PK+u4KFlQtnNJju/KV8dYhgYf
4vW/sFTGYJ9H1rodVVasyobqB/yzLZQLtCXF0p6NLckmKWBBssNFGo3Nh4VOlUmh0mQF1busy9xl
lL25ALXtcBEa68wuPTecVCXeM+ncsindjGAyaECKFbCa2kIYg2sMJm/b2giy6ugo0zYoVhFgPeKf
RIoiDBDHe5zATtoXL7rtWB1hE2i1uofagU2kaDvRv3d3zhz1KHHjeSJUBoap/Z17qnp/8su7pzrJ
TLVzKdRp/XKMYpJDmwddqEv/FgkOLmMcCQjC8yf4ZXZTauovZ6+gzXbjn2kAyM9wUtvIjeoKWMmm
u0hdeR+OBszWYie8ovYe5s5thaN2Ui1MK+Hvcu5v2/NwB057eyFp5xP4XyxtBlB1JxwD5zOTr1yL
G+GbVNv43YPSsk78EmeV8piYMMPOnWPgzrnvNIXvrkOjbGtWY508TYPfhKQIE/34idfOKfvM2LnD
ke1SaI6pPKp1XL4xeXPL7WLlgK8MYDTw/cgrjB+R3lKZrQtl3VHDjjho+sygMotgkVvSlIrF3CY3
8dEL7fHgSjE8zPxR4562vMLytLZaoZrbSehJtq2utPRaedbRqLh6nuA9vRoaGWHcS6O+PuMWmVCN
PsxOYTFpm6w4aeF1R/bZrWkkU0BYv+rT0xb4ArLZWKSVrYNpK7p6nIvK5Wm6xLAdG5Ad3jtZCtIr
LqIJwMT1DoCiOJTIW3bsxORB0grTetkYE18znHkK/cH7NduBdtj9Ms7wp2708a+24vvLvF49PGif
WZ7VWS7iHBAVf+f5/T5O6iXTR63uRueuTZmUlowHRas0lABWfr/xpI1EdAhx3pP79eQBVTYeIhi4
JkOe1MJAFIWXowp5WdodMxWce73VMa4fQanBoZg5LnGkVKXY6rf4Qa5IQpJo3k3AN5e19oSQv5cR
IVzmGXTdELULGEa3PGsyjexrKj1NMjhIT5+Af4mYN+qzgJDYgxZjHgOMjAV+JwYjJ5vSlUdZ0sGR
4hmn5qqLNtlmhxaVwD3ACB6GXRefKHCeEpAPWpmLf0VczjwIrzPgBkG8Lmc4QHjPeBbvaTLl+QO4
LLkJiacsaK7wGKiz600m9H6ZvD3iJL5XdOLNCfUkuZE2BbTrX2wnbCp5JeHwpXmB8/pNXEe3e4k1
e0FPp8kQb1P/mqtpY58C2Lk2ZB3Lafebouc3nKZGlmPXdTCvxsah0yn9w94uLpM7lx72Flo87xw+
xaXtxDLWq3VdzaS5fmXfiscckhW2dVwFQQ/24Hs/n65K6mcnJ1LvNxZlQGdryJzF+QktuJ0KWYFX
mKr/86TPnbEMD29I1OBwQWQiWe+mQLf5nzjAiUeqO9bFUAq+01H+p3QedmMdkpITA9xHL8+6ozv0
wEbEbYPUt2Oh/AXg8JnzCL8RjsBa6WpiH9tKSVnyjqdhXyFaa7SayR1rHgUGXHvgISyuWt6Gk8GF
Q/2ob3fmQDq2D2Tcz7n5vfrjBJgTKcZqKfQEH3RMJy1nI3yzQJHF4Z5F7N+VHKPGNfMPe1H+TVHO
dLLbkRKe5vIAXYkXJ2ue1Z1hmVDA176/M+cUHFpkV9zGC8i1J/iWJezXlHrplf+BJq6c5La5kTT/
KFx0i7MwIJzfkVfWHnkVmk08lATBbTkAfNAn0zSpaAGAPtPTNP04fL4ekgkPGI+ga7xm5ZmZJG/x
IKvculBZiOVT1JoevhQj2XgjlFJvisYdGtWP3qoCR62Sbktj2ucQeh+cv2J2RFGI7yNGXDTX/5Hk
2sVPM1TviM+zVt5POrM51jhCUrI8Y7wWWWXhTOfYCcIkf+NY+bo/AINlHF+5yf4YB1psmak8u8wf
noVGVSK/m7ELcHc/ZsamLUWhNWO6s/xiY7Ah4OkhF+GaSk3Go/MptjeljU+ZZy7+5vgvpgj/Mym+
gDoD8lcP5m7Q3lIcZmSF6YKvFCw/CbtqlE/7mEvmsit6mQa4UDYQ7TIo67V4BSo18/AJ2SMnlVuu
R7t+joCZyvtkBUTRzL2srtkUJuDQQounVQ/RC6ow5S9OgV3XiqloXMfRnuBDESrGNwh91zha7WuH
2oRNOzMOJypVzLYizWlOPgodHcYgG23Dblp/si50Z3cfqY8IZHbiMFSzH84RskjprXK1bIQM02k4
kuLkcpjdWblks3Bh/VG3WD1KPg5ABZipXPW8fuguY9IgoHj/pnXLW4UXI/KTksszJ5ZxHpT8vlAU
nKbkBVsxIK0jrmm4xd2xon0fH+0YywAV0opPMSEwNnsJ4XbYONUMNNn0dmqPBLzX+sYiP92N0sOW
+rfEYZJkXX6uCZ/BUh9hbwNkZzqNqcKyyWaOamQxqmHx5HzXjbY9WSc5cOEMuyG/yiwzR58MBzXx
WO8CKtfe/ZQJIx2IflQNBO8au14DCYmmzIfxNbdFSbLjvmzWb684vLTQLFBofgPEAyEIurXFsy0U
uzMj3Udg8bU+I0dJTnDHEw7ELp/hs8jj5Y0m7l1lRG0LZ1j4Iyh9eYA0GLZSHZe2nbCJgKZABbGs
dNnlEx2e9LclfIQMsX4DkgbmKS5M4GG0bibE0eMpWiKYiTBi6BxJZ2eGyl1eRo3z32ocpZgpDS6+
DAIHEK+/ucVooP5JI4JB7sxJ+YhtwCQsyWu5BTSxfCupMAoiipjPr3mzvCaAG68j2I4nD5vEnd54
bSoNEdXVdM5RPZ9opOE66WvIvUQlH7GHpuw1UShlsFy0dmB10EFqidRgg84z8PHPN/hpHWnqWAOK
A753rtAjupzQTS+AcckOcJOnftd0090Y1NjdWCzbckddHLdhKG72xwBtDWmJ53C1/qaFHzYN71e9
ONE5UOHTkZ3m4L50bY3K+siYnrvrp2eW+Wqi3XEkbrda14Q5oD6t8uKSzMnx22YFnY4Aa08GxF7A
0oFgJkHWVLK2BSYRdIYB0J1dygX+NZ7uigfVP8JQJAsTi9xN04Kt0YsiF9cc3x1M60Is/5jODQog
hkLuJbd1pdLaOCW0liWPCFNB3Cvk8BT8Jfltw6uHYwl1VXNioRt+i8efbhOv3ImRj4WWlZHcJ7Sx
9kN7dahuJ/Y73hfIadwJwG2NMInzmklP26RUeulw6o9iq1dPtt+OOO8km2qTL9VpF7pYtbv4kT5X
H7aTYEx8ph0fxcWZxC/EDxKBnDA37/PX7xgTNQNnKYLKjFXqBoLjcW8h+ErQVJbh5JF3U4yurOcu
rSx5gEIv8gWgBRtEAtYZkAGMDafwJUUnXEDhj74ZSsizOsbxFtVomWfslUQ26tKl/cOTeMzOxJE6
yqLVMFqbLhhgU6cbrTtwNuEH2akic2qXVQksVdFwUWtf1DNSq/YvkP1zPZ+FWdkb+SqjkKlqd0HS
/tID2BA1MTWsZizH7srBjAKQS0diD5lpnAfGOS7e6+YHos/iSflFFW9Na7f3HxcfDEvt4vzyPtUf
yTGi055QZN2av7U//EogFvVEQ00O398taWi+NXKOM+zjsXsYjYJ3AHRijnLowQLzB2+0JwMq8QAT
JKS6My8gLOWOpe14l8SJUuGTirM/my6HHadIR+FDhe4SBwBHl+3ZexibqEFg5RyRf8amoWbj9nA0
yT5aVvcssFb4W5QUUcaYMPxSgC6Zu+rbVHwQJ2rqwQHT3wlL2olIyOAfA3gcmBwWDGY6GCIYsoPn
HisjRuEYTzAkfkKM9Gafd2m5SdG5gKkzsYfNNFVpOl02h5oJJmy/3E4tSeW5GH+92cdXD6EGsuVZ
DaWpAlHeLudx5amcWRn9eTMpKkKML2J5PtDK2GFoIaIYQ1gNShwkQ9+fzoDTSFHS7UxuULYFvLt0
D5cKwg1D9ZyDeuIha8FwxfidpKRhq6y0si//mxvnftisBhqmTq7Rxp7EpQUcGF4TfSm6LaRHDAiP
enM6AXuF6eUBkq3Ou2xo7RGy+9CpZJvXpfeemknIp+/z17vYirvlFXLF5D8qzrM42mh+8CzIJ/od
pKBxbQ3hAtJEMt07tZidMS123OTGT9z8Om8HonuFaHznBukqR4/potCt5jlSwTl6AWU1TUy3bCz5
1muk26WEckSesGPnNmgxtbXV0OrHZ4UCngcVCuxwQNPg8Rh1ZTkSiGd2YTJ+XJTKjheOwGLgu+Bn
0IiGuqgzUxSxYJiOCEBP/4+laKFRgpABz4TyjRvA/xeJzdlUtQtL1NjxsDqi9IG5IvqggYRAbWGb
4skLK7H4TILrxDjyR1nb2jAGD8Ha/0oxjigPv8SMIN4FSym2ibjyqIRL3nXU0TwIXkixD4BQgv/m
O0r8ZbfUxdzaeZpcrJgieEWxIyjJM9sXv8rKtPy1mBAPEqn3LmRK6ptu7QlFQX8M3WLeGFy0U7O4
EPT785Buzq4Gv7V5lkejrHP9Lz52DMOnuXcehYHTNE8jHb8kCWhSTXa3vjVgXcqgRKcZjP0GPyq+
GRLhJ1K3/3wrGbT+GDsA0mOKbhwwh5UuXbiChgCXXBBLK2qYd1THZjy+JjGs566wxVFDYLZWrV9j
/I0rGfRSxpfDqSVr5x5/tBd+VW5k2QGTe53uB93tKdYYMOl2tuKAFd4/7wBEl3eePozzE9Ef3asg
rMh0zjy1g7hzC9Wq0V+IEmn9HVsCa8IvgWjurMSGCKo+fZ1HnRIwNGv63wR67mVEAUVxIYM4pw32
MVwNNQvcrpYseFHtEjJu2pZsv4EyXe/OZ7OU9CKM92t87Mw6lCjQGCIyHVK2pEZGvhq/whYk04Mh
vhVmRL2XcVZaM/KIn0wiVRNPYhJ5VEUp+jftmyNefKs6VfmxVkxgAhGtXVxOYs2bOGnoOROCkyew
cna6B18ciqO1gxxAUVLJUqcd7lEX7q32gIhowmDUJkbHix4mWomb6QT5ut4N1WA5+BmB2gNDdYCx
XGFaapNSjGVi4G6lCDkkDBKBM8d1ov7JZE7KQcjn6gg50XuW14VB4xn4RaSknr0VfAnpUXpsEXNQ
w3NzRsZmQuwKXIUfpjTaRZtauiUlFvCy73uT3YI3j0cFHu3WZUlhdrzTHpn2hX0fZRPhgtWurbqq
LT+AFLj0aM3Q9Up2XoGe0rFO7spXePYOUoZPzeEs5S2GfNLxzlq/bdrTULfgioxr16aIqK0WqwLr
0iHLXRmE40rKw7KMtOehq6NeA7YqB13HCw4Eko3KzaFpAgb/oX30c6s483XuV6eI42cz01nUvxhh
qkxJFPoTqONMv4Ggipk87C1N/FzWrQLbor3XSBcSFEMgiJ0vFaHjwfP52mu0KOqSETZRnQuS6fmR
iO4IMFwOb2ACnzBHos4r0J9bWErxxoyg5yuoNSdWsi2AaGOVWAQqKah7l+Q6KuZycJzSxZVpkBuu
gjBrG3x4rJZTg/2LQvf1NaQOJsReGCBJMyM9ZZSrnT2Dx5V8+h03Xz4PxqCDEIoUp6xAuqFq49vg
E3bCR3NM0vStvTDltU/ZeUTy9oUpmiN7uTSONWH/cPN9POYy6LLuPephavIsqW9U6wRiuy22DbkP
7bTa8ysrp0B48G8DZUw577hUqjbxAJF4wp4go/nVxbzpRrKLQQa9nZnXRPB4jsIoO3Q1/NHo45HQ
jGlIPPUroWhI3/Uy1l40Lbf8HHNr2ZIJt5DVRvsYeYvmMOM1FMcukZ1YfAIcdMBHS0/cEEys/srW
W32Kvm6Ft1t3BrTasoSbxmAX9W8IPlUFUN8KuenrUrak+Pv/K2JOpadqAIPK4pAXcHt9AN6WfcFi
I3cVkqNg7SVqnL7Jm58jm63zDe56UQiy4yO/cJUO0jkjujUVwF94+iToVF9Sb5fBaSEX2SxDoZ9l
D/XVchuvDDcz40YI7xdvXSrFdlBg7XlanIfuk2TAQNShYj5e4VOe45q2JLJ9zepEzwS8ctw0CBzj
7jycK++YXbEk1gaInVdKpw2CxYqZyMuPoy26+9eWea9gwZm3V6ejcWj4Kf/ITH92TIMvhwdMUXQn
Xw2rYGuiKIFINJ6yNJZ8bunTXhiVIK0j6XV/mgu73XdwyU4xadCftMItZJ81biWUkLteokcseaPQ
DXYGpZqhQx8SLmXrt6rHIh2cHSDEdFbotCKPvxOwZ93qFN4IjbmkITNFcmiTZQLdyY7OYuujgOIW
1/DRQbOwYz7cf4pD+D0AgoNLm/gvyAGVoTvoVaqxwhTGL140zawcs6d7dNywjl3cRDBdruy0U+Pm
bspXAEzonNNoiHSP0odNOVjTzX99fIo5E+q+9cGQ4kmAZjv9Y23gZ0M9LucBsyNK9dFclwkdpgcC
GuGwLMLFdUd1sSXJevmCFD1M2F5X7ys21imcVOttJz5rslmNFAbe3QS0pNdp0VAB40sYJbGDavel
XcVtLxM5/J7dHpIC4bC0kTUdOlOF9DYtOkx6pFMCxG/JzdZ7UgTbT8CBEywhaOp6S7m2vgdfGjfQ
FlahULjwikZWDevbY+ucakDfbS9GEPSPxjOzQziZpHRwpuU7+mGt35Y8v2bvIP1mx5Ppi6QNLwBZ
5xbEQ3zToE4JMGN3IeCEeXQWBk63578yyw49bayFwAgVLmiuag+kELyHlHeRLcnpypBfAnQXJBK2
szvbtC626TWGwKq+kgyPjubdWGno6HlEQ6/0n408HKA1b5S+w+4umyVkJZy59qQR5s5MUkn5vMn6
XLUCmXN/2LUfdQ6fERgDQR40s6Y2N8Zo+Qd208x5PIUyn6jnaRmA3/PBKT5pNtsatcAT32RS30WP
3nYvYRiHExtOKqjb/6aRn8yrJzsu8V1sRpPtO7sIIoN7FMzL6X65ArD/6HTl97yM5gdAsRCMDotd
zRRRWuUzxMKg4JTzwf4LoGyu0sU3JlGVegcD4FndWyZbF2PCq/qY5gxmPqdRX4VdCSTXkE6zDM9Y
J98TYrAxkY1kU3mWBHHgCGLNGLp+NdcuIuZepOl3JaLzcc8Ey1lQmvUiHHVybaS7a7qBHGX6buxz
oZmw/7ycU1ac6ILUHcNGEthcd6lr46kIHtFp608tZAudaUIWG8oEjXahy2IRlPO7tpOLsXh+y3K6
Gsttf+vCZGck+QyLX57la7ktSOAIAjIufbi9M7jEknhnbBB1IpqYbB3TF/tGJAK3zFzGnMNlZoxs
fF8BrESnRYz9N6zvXFa9RsG1frL+DXk+GP35abjijIJaQIY7oIPiAyQeTXhO88zBRsr1+GC5Y/VD
CRO4/7WaniCdn0O+pZlQ0Fo28eFRMK/YPXx6PlJu8tHDTB7dxUPITN5ymqYUCNy3pgWaAZQ1bNyf
3Z1zDMvLYDq0jSAQP9GV5mKlB+b96zjYPh6AijrA7Z110iqKX6lgf04QlJ0cdMPMsUJd0l5GHls5
6vKAjt7DIZaB3z05Krsap9Dhl3CDDSNix4xaunGVwSLKTJjUnnmDzsFcIQLb1hzUi/fL752PwxmU
uU3Xo6YO3imiCT29oig368VLxJfNpEE6VhS+zb2JxbxlxXLSxsSniuYHRuC+Ak52f11WLG/KMqmr
naOjaLFVV7mh01QzNqtZqr+/cew1DjGWc39nddTlBjjUX77pexFh/3Rxh0i2nClHX+BV35Nxig5Z
PY2/rA9aJC6NbwJAabGxGD+cWWt1NDI/iLNqB8RxhCS6dfzkUWpmkDGcgxcQL0Jk9630HA/tOpL2
Ca/o3yMvYxWDlEW/R6Q0cPv/gSL9DBmwsi8+Jh1WWluv+BR43YZ2Ybh3IuC2GdNZVLu9zVdrc9NG
PGrqKVW6geI3T6uM50sbHmwYNdMAQx5hDbnzX9dkIdP6oqsO6h2ilsy1GPvofOVHdyPLW7F6lacj
fCTg8dMlaulj67tg+aIxiPnxCsHN3OraW/oYunb/tkIh1QMe/vwslH4rwbF4g0Z18CMnaR/Gcpdp
pc0RgoIRBDq+YY7WQbkEgjNL2WZcsBXHH3SqDX9M3Ppq4ye+xShZIbh9OzOA3d6JuIaWf0xNS3R5
qmGKzaK95EyiqoIxvWG5YRPC7ziKOj/v6HRh8fshI/auFNn6Ro5AB6G1fNws5CVKUCyRdOUfyBi3
mP4v5WA/QXivtfH6s8hpPlYFDCdljtzBJWPGe7l/6qwojLlpnVsgk+BVosictI4ceh9sxcpN0cLn
eiIKqVtbd4MBUBY/APabV1kg7q5n6bhR1n2b1+0lk8xLeVCJXu5p9ooDKig0pDyHan6p7XFkupL6
g99cmbpu2eGHsUj30UmB1D/QZG+4xANCfa96uJrp/8FycnTBZT+kxd4oC5aV8jb9JSkD2ymY008s
Iv2B/R9BUsYoly8eiMEXxA9CrPdQxUPF3NepQhKt8n1uaZDJ4hz0Wlttk5SSSGVryeFN5o978k7m
eD73sROw83CUyGC7wWDy49iLhWqAYRyoQZ7w8rWxGV8o2afHOkfagED6g2yDg8L7NlXAGPkKOq66
016G4uPruqp/FiVA33qyr/63Ayz/IKFu5iWn2OSK7oyE4SV0Vy7lS4w94D8PrDt7SZ3ne1C5ab51
YJra83NYNznxyHjcd2gFNz2IrMAkRBlNrchJZEEmfbFKMgv7vBK51sRIx9656f1KcsabBUC9zwam
CaO1fBKUcJE6uXC+hOnjVT7E3RMzWnMd7JmuJGZSNmZgd5f+Bzbmtx8zGy5dwst+/hixNatIxnyx
U+StAwJH4eeaNurghSljYQ0L/Mps+BXhU+jBKlRpv2UPk2aboUal8wgQsL1IDEWr7rJRPWD4V3WY
RVHOXyPJV4MZqV5auvOJ/rzDP9smLZ2Jddm+ODNGNXMS4SwykRaEWnIP3B1EmeqMWIpdu4SpYfLl
s9GL281g/tJJNYfXs+DXutOiWp8hknT6Cjr99JHBVHZq+9Kdk11Xkegu5hhDl8k0r9hHapGItlAC
w1nIbVdQSONyVG6zKEbGKHNy8XXZmiHFyZLut4BbmXmSqPStnZl96CUQPnzcMhQ/ClmXYEhOBzVq
kLG3Ls2sC2Ti6NW7MsfuI6+EZOu15/taE/afBtuhQAZ5fulHjepdTub4fm3819PlcwdsgYokyIgW
w8r342qOQTlka6covFkfHfTVgNJAE/RdgySXmOf898k9XZzMVjLB9myE65dAWmem+0PvQIxHybly
c1SHK1qRwDD2pfQosE6yujbokBumVpSGus1vUdkXomaerSOSe/fF7IWXhQJ6C8fIF+LYw+o7c+Ft
kjpxQ7utQrtwSZ0rf2tag4yP6lLC/sQPduNAnWRW5MiVioXle5+p4RuKvV++DwnzOs3fmnZn2rQP
rEKcpkGEEt0PMCo/VoAE6VAecaon8encTVCc3vkpFV5P5hvAoViY9U5APyFcWrMtq3rQ0Uk6MvG5
t+ffxM1LQ8yzaCNuD0uipPN3rY4rI9KLs+r2Kncoi7xoSLmd3Sk48VtPSQVsYSB+xhxYK/008iiD
vgw1/Sva9fgxHn6i04SNV6EFNaBIwrRDfFypEazVQdvB+pZe8IkVLYcCOWd7+2YvYGkhTn9/1cz4
LzTQPSDRzN8IhiqfokFJPtigMt8pc2c+5ZHhfdeH18TE+QdGOrkv8T7hrBAuWfzKWIlp1dYqoRDD
K2N3/UXMAuiX899BvGdqg8VIGMxaXsSb8t+8ffd27LWrQMgi9YuojJUi3sT17bnUulJLg93zz907
jpo0s69jPo0ssYhvw4p0J/CR0ELZKzOYkQV8BR9ueonpgtzy3VLnqGWBNXnYQWPCBs0Vig4Hpgrc
4jCZIditgHuaVmokW7Ol6hcivsW65766cFdJuyDnE0holIqQEMvXVVd5SnZuwDgDmS5w9EXHiYHD
Dkxm4kBmP4uqLcIf1emriE4Q4DwtaeEnt8Wi3tYsj7WR1fN0IegbQ9MxSqQSD0m2TZahTnZwAXGz
f2lWKptffLKW0rZXHae0MPdTqwyuUGoN/mqutVPAmUE9w4a6kmrM031HCZt5nnIqYUpstcHmCpRC
HYO7RLCkBS9GDP69jd42zkrKD1AMJ43VYeSXDsl3XAoRsaemDiOcCMbDjtmoWyLPCMvSPJopgXkB
81VJyCreDaSQqDB00fgKjBF18l3Tv9u+StOlrtF6549jBCBVa0Ugwk0+t3e1d3Tg2lh4U7+J1PeH
P0Gcr3S5gorYUX4Ml67FELIRxVJ7YuyOdiz3KYuyGQMYBk5LvOF4wtMY5cCsmpO+Tn2qhQla5y7w
IHKNgSi5N5RgcHtDNr0ZRoTEh5xb/2ducRAdnTaFPn62XaLgjoC8sWe3qeCAYoJ5gID1zqRtL1CD
wpQhuKdx43cq1Zfi6ePRaIIgoOmEIwC6SMaze3NiAsLbivkJsw9lWh+GRatSkL/fn36NRHi5EOw0
w9KQu5LdtUxkxB+b+e1yEnCbz2RzlqXZg/tNfoXErStuJVpfeyEijv0bgcztQ0KFRiHmaTBPpyTr
GR7vg3k0e17Ym1jr0MvqjxKOpLJmg0MqY95G/XYji0nYm6pF0J2jhUFO8cpV72W4A9eHVyLAKZLn
DCeQiz8bS8LLwHVbseNAzrBvkd4dtozsimrJD/E2tmIQhqaLnhjZYUSuuzZ0I3y8W7WZv5N7YLvm
lZCG/XaDt+drI7k25TOctYBVQKcY7wQ6dTPjHXYx4vCr1zkBPZ2hd4MPleJfD0e6CEwicj+77qUZ
DpvLBJcWWwaDXMYS6tQ/1954KOtOiHu0U8i+sL6cJYtLnTfpbLSdXoasljc3LSeYUII7pKWK/b9Y
XnGc246iAaM+1hQf3k7foE2Cw6NQM/U0iAfRUoIsWZon4jEjJuV7hNzJ+M38aZK8K/heAMPS9mn5
3l2MarUqgT0iS3XyXAyR4gAB2DVsPyGtABxQrNP6et7Ep/9wYXb10o+c+UItUcbSpY7cLqw/yN8d
oTQUOsjiXEiyX+VyQr18k7S0KPNC8Ur9GTXuhKngD+cgU629ralQ1tly7jIvD/oJ9XfLl9TqPcKV
WX3z2QOpbj6vduxCQ3KZADRbbvcB8QzlbTxTVdnXHuuoXt45rpHwjPxQM5RUP5abG72ZzFQfSajf
uZ91qy0FG57vqIMdiJw8HOUb4uzArEW0CCLPqnBIIKveNOCqGCjT1coIK5USzQPSjybW3kpooXJb
+Fkw2kIq+i0J3XRe4M/KyKII9ww2FVJ/y8dHsH9NFhUeisn2XQUwgE6Ny07ucYUVCIZyuRNSvN1K
G97qEosndhSfovz3rZIntq/FKl2S1p+KGyQx8Ge1vdMxB8w/DyFza2ukd8vjR8A55cvGLG+UiiAg
GpEPsb70sLPRTCKEzLFXa7J+OAzl0NPqE9RPGouhWfMqZlFNwDSysgQKXeEx9YwEbc7aGALpMbS7
RyDgjoD7mp4Ub6mVaokczrevdcSTUnkOHexNmTMftnOHJnnfDQWu7d+4fhW9DgCwjlo5dRl13qxR
1TNIoZSfrJ4AfxbUzay8rJ5Kcvwp72JNRbpmD6X+FvhfWxwfHbAJR9gZbRlAmXyi8NNqo9qButGY
qCHmduOXmhgT8eK0Xn99A8naCZ3ZOdNtS4ykrKF7UTO3r+KKoGJgN+KkzadtjxU85V3LDDAVQ5B4
Q3Sqhe0YqQ1XFS29X/DP/KR8CYnw/MAuVEG24PfYY/Z3wGy6951uyfpM9aMS1Iq8lExWnjz1KH71
AtDnvgYthk52hZK3wv0/uG2lzGVI/qVeLaDcmtI94Mlp6D8reJavTiT4EC9jJ/6tMRqx2OOdikpi
fVyWbEKOxiCK3OCUj9ijq7xnGazebDsG2c5JjdkKBI4oSRAn9hxmQCFBHRHXQfK7wJrPQ4zD9nV0
WzVxu8zFP/8WLC4vNSbjhSqpAQB9RV7C/4Y3q/HeSSmhBSPdrDbEh+460PyXarq7BJRXqMcNS/Jp
VgdxwPZXEIMUD5m1wjjw1x8+xddUlcr4X2h4nJpPglR4QO9IJRPmNd+9ZI0IeCzfmlWrSuZKeW74
leRRpI+rppAA/8J0SXp6ujFAqUMIi4yH9kAfLImxtdf4nnqwN4BgHLT+iiy6TzFnjlcbkGNfd0Oz
Cfj8L8+zaJFObuHrNtSO3aji0NjI1fMYZr+eQ6XqdP/v49kUEMGdLsrVXc3GPSBBF4RgEkImV5Ec
vOjPsxkN+5Lpm9FocN9H0QOAueaZFWom3jqppQawjUiHw8U2fjMOxG/Hjllbn3Gox781jC2j3o5A
Wai9tw/JZOblogAAX1TbtEiXjPQ+XRtNsmfeHBiOErL3hresbG9S6rGGg1gjcVYohdWVAOSILTj1
I4mr8cstIrWxhDsMHUHEfqGwMNRDApq8Ep9FKUkjezIg0skitUHLjcQn6FCw+iCiUaEPzue89y2T
Pwk3OU8PRR0PHmj3AKXcSOZ9fH9B0g3aLMv6Zljg2iTEUPFQzoNhbSqeKmNQ5gRDFUHB5/NUzx8i
nHdatE+cdMnrj1gsDDB/cFVh6SKdeAr+J4TSHzvAKbbzMcugCtixmGN1YcVVQXe4Qd7eH4LdGY1c
rMAeFAfLMH0UmFGVHDKWWBRcMN/NtIVa3PsUgLmybZUN9vGt5vi22lqZyBshdOqYfMhD7dgefSkt
RYhSbKxTdS00SPhF3/fk46RkrR9K8Niql1WD1sK9saXHyfpobyC91wzVi/rZGaZk79CJEk0eEje4
CiPKiVGGmMUncQxziEjD6QHv5bhLwg9k+WEbd6dqCGPiF/N6H3eh6q2WL0WfLvQKxYN35aq0OPgn
80+UUlbmEul8lXLqj3vYPg/q/Qn/kAyzkSPUQSK71fFm6XPIXlY5x9/dlP9h+fNOjYG5sEmUoro2
whgPNIkjOXjpLvtVAyBuS1li/2Z//KIpaiFvvsRi0JhjVtd3QLiJIamtmZst/jDtiajkpe3oJreq
W8/FqN/Qe3jiTLjvzMZdFkY5BGJPZoIObltM+lzHOzGZGs+MA9wU8NphTrKItfor1US5TbpAYKfA
fc2w5pf7zU6gVBCRZItnAuzghHsRNjIDGx8+w/eSZmRI0sbAAWtIknBFSHhjZsu7T1h0I/nqGaKX
v8Z1YrJhvv+eUTOVTuqVjK539yhOlgNcZ+4ts8FuCGM76qY+5QLVRw1lgzSUCG2+j5KSnLJ2Bifg
12O9w1sTk1pq3Lb/rdyEivyQ9H86nxqW2r92+0tIe7s2SeOBoHdpLH2r+F3UiwhrCilSysi2/Sxq
JtZWR+o22nP9p0U/1TG493owHBvP1atSWwO5eIZRv14rx49aEH3JMH4zzpdb5/SDsHdz4yjRfn7S
3U9mVxoSNGUnoaApNlUggonW6fpPfBMTQux2tSxOljgscZRDgG+VYD098BGY5uTtxX5YWfXplGfj
yP0ejgDX8nPnWdibooipDEZr6idNtNCYDgcUzdbY18ruam/A2D8j/HitSKsnNIP8Th1JAk2796cB
pZ8hF/QkS9EU+6IFLfjgL9xKvK1cWvco4hi2+TVjFLAFPoEnynVquo/SgjdDc4WiF7wzKJkB99rW
Uf1CLDSK56acXiVhfJXXx9wD4IWHiv81jv7s0cEBVUoPUsQWOkurMDJbKUww1fNvdYWQ6dF/dtAo
6b1brBFTQ6VCFzDesm11dp9NdLf8KyodyRe6rVKlUYWiq2jR/83z3WhGCDOHXTJJOMXhc7DNeCxQ
TJMvJemAAtwH4/AHJ7mfg1w2oUIww1BJKBf8ZeMiMhKDNgsZnvo0NMBmSAyTrRYpjfikgKbv2ZTU
IQKXcsd8LTTE4DWU/Rmm8Eihc/gJGr6L3c19HNodqLI0NO/TaZFrQOqjuFyxy9t26Ak+E2ISXaSe
QCVNGM1ynphMYP3R2os0z3xdk3Y6pHfmTd6W+GD16Ij6DrhW0IKKRyDmKqJNqhAgAA444z/Xj92L
pyi3gGagtAKqU3rYXImDDboEPgdBuQMWXwRDjrBH/WJ3CKaHVQntaIyfpi/wsLTnidOI+5Gngc9L
yVnrfXcsZl8TEmwnQ5Q+mRG8raCfVPb/G7z5IJUyDhEUbnCgpEOV5cmS1cx2FPNtKUNxeO/6qXJH
56xddLvjB80W7i6KjFgJrtelYevS4Axs80BKuQFHwCVfpe1hVBFefnYu0iqewn57GyxNS1/VtIH7
17tS5xDw0yF5VjfFmsrhJ0XYD1S4i0DUr17iXdfaOWbY+7g/fO7sd/jcI4lnAqLeB/+D3gdK9K5W
oVzG9BOGD2txtVyt2PJwFQ5J3fqEU/0agvHEKqRHU8SugdjCVcdZb88iu/YCiMVh6aW3zrquPyOX
EoAD8tjUP9/YFsS5Hg9AZsceJrlw6qTjMNoAVwaRakkbiURNJLvgZ+HM7HxfPDJC3QZnae3VjC8O
dCL0U+aYVG2pTpp9DJODh+BLN/h536j+dE5eIaUgHQpd57rEr1h8E+6EEo1ZdZgDstUyiK5htiwB
ZE6HAHUn2iBYN9dCcWD7kvAEauKWXxToalz6q2pxwaEj0qX74jdhA9N7shSRHCY+C9Z78YXGP8Jo
WjgSCC0fF0POA7ck4KFmAwtwsA1+E1/2p3hyha+ft0VPYyhV1jFO3lZ/gkWNEPceFsDJl2vh0kHu
KHjYMgrlx2JkV1H9g+xLUpo2WXBzv1oy6Mt2v0CuVKm3o5uxwpdLaux/e5EnOnlbSh4Xxl1UwifA
wyz5jQzPQDQecvS+USj31Mwdca7y82AgwSKtyROaB6sb2oiIQ/Bx2X3/UZRu2xBCiMo+652qfxAA
lPe0YHeW7lsqhFWHMn26iEZbH8uZg3Et2psI3qjBv2bwbMM2acPWK6K6tWJqc8HlVfODLh9E+GgE
1dpLDptoL9bUPCjN+fES0kiSBjcU7LEB/FpZUE2mIT7LvfuJEGBtdDNFuuWacoUW9NpAhRKHTiCx
hN4Rirj6mM+unTTPb2zbKV4vaeKz+EibA+i2Re616tCfAGXg4sXy/gOb7+CeNucC7AxINXm8jTCy
7HujFtYAG5hRxZsVKdEsdNOCiFVa5Es56a9Bn7wSvtrrkS2REuB+UBIvTokSUOTKQo1Hh3v6m7P4
ZB1rkV1KsTFWkLb19u1dMwXPC1LgB/+nnopradEfO9ekEMKCVferWjyJNm58m2e1h3FLO0Km3ogG
xvPkduXJ48N0N3We2Q0t9zYDK8s/ATcpWvLad/fUInS2ZW2SPhDB2FiF0IEebyHUnMDFTL4R0Cbc
3mSD3eOEU0IWTtFLgD+TuqexY5AdgrXmnmdXvsOuo1AC/dM3O3Q9J/CpizvpDTlqGkQCbMBJ8Zg2
g/VV3djaEZNQ06dUO4WzCZ04cxk0XMA9OO5c4PiXt4s5HqLtuD7VSc4JcFNVu/ivaz5a5gdMDFbm
+Sv0hH++QyD9JIi2SvlPWhDODckmuiZXnhGp0w2UFvtpA6BT8w9nbs+Ft7ilP3/BoOeEg2T+fn4B
CF+ScL9IHEGhzYArW1UyDVm9UjgpRZRshkdkh4fZHvPQB6SbDzvcQGCzJKVANJ7bp6EuF4EAQrmE
QGbJBiLP6yTsLQmU2NY6bevRe5znzC3794m8MBBzpP59po1wrxA9nt45nVnVEpGVYcYwDWbdmHaO
fkTKd3iTrbJObjs1wJVznlYrLkJQVJ/BImHauIASmZEofcqUt3vGZfCFBed1I+PtW3xu5/hbL6AD
G+eMQvQQ64jwUsoSQHx6KGlP6bMuEmWJ5gDEHiArLpHZMWanjrqT+ThNiA4iuekKGYY+yaH9tuUB
6Uxlo8aKJLr8fsPv2qFjliCS6v4D8oxN0Q2VdO4sCHhjBWKK3zJoyPWiVBzpONRyFEaEgIWx/fqN
+8ljTSQAmf5vGT4jqb2q1nAaZRn23fxcLyLZ7mfZbJ86P2BfbT4RErL4mPJkUIN3Z7XgxpjpftZZ
3V6b8nY6/7UdV4Ca9O9Eh0DvxUzY7WmQ9/swfxLCTwj7wAkD5in/Nk3+eexB2jKjSh+L0+tVJHDw
jy9Hp6ZEL6hDeRhC/xIXO5uSR7Zi1zPTnZCTORexMGq2dXSkqP+RKuCa3lUWLWzZQ22xosu07fG6
nnmmlaxtra0JSlRp6XfGj2AX6gX+xfdXcVjmgtwDLcXkdMbpbsq/XdaQq7a6hYNzhqYvFftdR0oT
ItVfSFotTNpHtaT9NZQwI3V+VnZgBNp15/I0AMEMb2t81XXDuFzqiNQYMUk8wYxGQG0Zz+yGYJdv
SBNSTLeJx6+JBAQSbOg4s1O1qL9rAeAHD4Y4o2r7XHeN+CaowJUb2pFqhvkASs78W48JpWxybqME
yIBEcH0VCv7BXuwLy1cjIqLoyRL+rn19l0QyG1LYB0mbxtASIOB+kParR0UkK1rb8wnVE7aliabY
gU9XOtDO8dY7RO1zwCLloI/DCnhxzXAmNiU4eCSreuUwh4xym9Aj3JaVol9vAOb/F3poMmYy2CjY
QYXqW9bhNJdV5kH/j3glsTdkJ5QdcPKmRBX9nHveggU1KJR0cIYR1QXPfKKChkDLp3cqsYUURedk
MwX3/PkVge1qc1mSa70Sh9z7Vq1h+eYztx+FKV2dCZfFt4LM5akEuvFH22m2s7QHchbfwCYfgxaE
eh2rJpsUvF/jwHj7jFrMk8/8m6eC/xeSPwgCnC4l1nnWzWrw+te8UmsHn6sVNBwpgYYh5zdWbMiR
T/rbJ8DU/lNBcclZ9kV38LycA0v6zPpL3TtA/kpUjd1rZKQvfc4wOmYf2V+CqeLZDA+ecGz1yfNR
jsupO6ZTJEIfGccC7mkP7f1s/R08YQTDrpv44fHHBR2IkC3f9ldKxlx0RWscTj0eyd5QoZ3P6OTp
IvChJxoxjjTLU2INsiDlfz6ecmCyjgDZrB5ol2OaS1HviKaN3JTmy/AHZEl5ivOzR0hMrlDPuoGb
Qc5n6/pR7YA27MvlDVHRz7hyRQzmTneh/kjTjrPxDwsN1G3M9wS7gaUGVfwC2hTIfv+QXu4GQxx+
vsdm04MGtZ4drrKdbZIEVTts7G/tkW6a16FbHGP4MHe91fhxIFLU3UUDwC9Lluk9Hqpu6lR9f+eE
dGLCd/mEbF0RpyQPlIMbahHcHIDVgxEjAML3IuJJSPZF4RcJtlnllJeoWLDPJopsILkLugNPc27/
7oDRtI+97rE35nFRwI08awqqkpvfTEGbTpAx4a8VLvp10zQEJY6cWAb0uJAL2CdM8aXVwumVxVPv
u3uQRUzkRGvEhMBjM+8xOUer1I4+skAUEGBgeUT689rXmBQB8OH72Tuc/BnUMaFNFguE7FCi7ezA
CFWjanp9jtnzGrBAGMQR0GToqOJtw1NQHnvA2RfrJCwl863T7O7RnTC45AgZ0nOzVgWTfIM97LX/
ipLXfDhkqjPuxB/BGKFzobEIVap2u42hc1i8SHmwjuKjxt6WvILYYadt6wc3KcG/disxYF0w6yZS
4Pn3NEFO8MqIiYMw2PDwnSY+JWlWNo2psCimVAp9R60FgLnSxKDt48+BVT+rZJ4PmCKea5ser//H
YskIG0UO8cC/cFuvUl+emzSNd4GaROlUo7oTE2yI/Fl+49s3oCc47Fjsmd32g0Wv4rn9zBB0Sivu
j2nviVR+xem9Z4ZikgA17P+i9tdtkwjgd6jC6HOC5DGbPHNypTZi7N3RyTA96KgPz3kTJEpl0ucu
OdszoC2JJYjvSwH60V8xlwQ5vtK0ePqvG59cSdFQ73GXlbhR8HAhlhDTtGq7doo30YABijpfwxFw
rYqiQ+SqR7v/oT/nvuzPQYVyEk9QXSlsaWtwex5ORyMdx6reeVk7PKEnXtRMryVRbwGhIIABOb7o
rjZ0nvWSsoBUYLh9kU0TB7cdd4+ea1sOavqwHaQAc48dRsXFTKFaFsWWogmnpi2XgxUrCpNnnMpi
B/DjK8llhbLs9M/didnteEoP15/ln+mErD/DC4Vj/WvBKOPcLFDhIXFEi5PKIzzTax/3+JjXPrvV
kRjSerxeljVgAmpXghsxK7lWvPCATmNROrxlOcijSiv7zcoEbImtKOM9kTektKy4aoUZhPSXTo5+
1oFxdCIuOWgrlVpzPQ3uW9qVrHdemywCWHbi7E1cFNPMa/+SXT450hTO3coMywE0Iw5EHsnEcIFm
+rVXcgz8R4XmQbp2KICGMEz27oC6xC+dc5S4WLEQSxZsQDX0srdYADd5+ctTPe5BUTbaDvNVlWnN
j1lI6cdCMpw1S4CJPs5QlpaXGHxm7fibfpmzBswQ6mxWfPmDSgnE6zgL4gL2/uM4Ff/yVuqknQ24
TYsmHIpEE030YrMUJGL0gydy3yHmPLszFZSgjiaP2eZYueHv6yhkn4WDDx+MEsOZD5Wf4b8E99Il
zKifFf7VHiuuDvXVezPSFYgIfcs6Zw5oQSnex8a0XHrKyVb6LzBzKmsiciaVmxuK1PwuwNsW05rQ
3TqQ9Cs52XYrw4fmLHh09Dzbjy/4dBVjRMO6X4B/rZyf9tRLM2UpUMLTurJCxxZGpbDGvSwF9anA
kEsG+Tixmc5xV7POGewMMxbctKE5AwxyFmNqPdEhq04qVQoFRGyYTU3Le2496/jmp0fnyYEMUn4z
6NuxjxwMpQmuIli1Sgslah2vU8MhG6/StX9WI5T4SQ3m+TtfDOEOBfE6DfIq+qhXInbIH2eKZRC5
G7WL3n2ELQgoDzURa8LfphYZn5tgYHZrdCQKdxGxut8QahIRWqXhwC12wWGtjY8F547cvWZSqIxN
MzfWFTwr5bm7+SmYjyAlF0LwVQdywjSh25THIjcngp/MUBRLz7hczVBrXx0Pb0pm9emELKoJVvfu
zQpLNL0nhZ1K42pXM/PV0stcSiRvQvk7NoHbypU0rdGgVwtals9sFY/HPf4dGfZ/b9gfOD5FSEZ3
AzIPjjLKLyqZC3JQT4NMd5qmkHqkgWG21pqQw3fqUKw5ijOmyCKSjZnkXKnmASsCMmcmeU5/Y8wq
sUHhY7iJcE5Vqk0w6/DH0+kbxf4pcdDEV3tahPYLuyM3gdR7JmiPLxoXk3dnQZWAlnmV+3e3LFKe
UiShsa7oLBfNljGw+0IyKfe0GXjoGOp4mGq/H0msZNPg764L5AZrafMNuBRaz9hH5X12T2I5egxs
5Ri5ZYrGUtffiyJ+GlA3oBN0V/vftHXELmZ6qgJn5HpLRrEcE97gxsK3Sn6SdJep+yz/ZN3zK/Wf
Yq1c3fnmMpjr4NMDjBXD9PC0HOKlRUpqfLvzv4HdQyVajehXdoZtTnlyQuROZDXsfWnwlx8wfkMG
JT5Vc3ipta8pvQYKiXslP4JTsr1z4RwgUc/8QX2KIPSQYP6S6Zpsz39+SMpam/aL20blCV1DYEHM
N6zvjKFvP4N1ujZbgFgbH8aI8wEh+yID/Pfm7mHIgpEj3OWiykufsE264ENuvOY221V8EHIO7bbI
r62zdzjogzv+D/ZHjkFeed+fzxa5LkjFwpt8ubONwWX5qh0s3Mm5FLoOAe+iwegDwnq8QwJjU5Kp
wHPLYezbdCJv7U1svbFfjoiGZos8aGO98wJufyXU8ACM6kjJeAF0AooQ7OqGXaqQ7GycVCE1sDYM
bAdf3sHgSiYFXjDtBFDwWmsHUFHB9mB8LGk8tfAA/O7XRbuEzVSQZ1NIJhM/fSEJCLNGo3+pfnlL
JHWfVfKtuVKDcG/z1PelfWcHyO92u4mOFQHQ+gdC2zjZ4jOY0UpvPtujDDuZ1iZtB+JWn6y45oMv
1o4Oi26AsS2zx3s4WwyAN/dG/4+/CDO9V9v4mnDoiMzi9+QlPMkUuPxph5S5Mkhde5ARRf58W3L6
QkLEyDV28GgdWbkIbdqGN6xG55XHKckCCEZwbt+hCg/2FZcyZy1CQD0XZnxrMD9cxYlUnUDpv0Ej
67it7Rdhn6naQk0R+8AFeklcoSAanqCTh5kFqf4sCpRmL8P0ZhPnrxU0U8x/Uiei6yZVH7jra+pS
JmZZgTZbwyULf9/uThqAcZgSjN8HSMa3omYwA8vbxKg1gZk/9y8BkhqrFam60Bigu4hBRCG9JTIy
WGQe8/BTGxsrczExZ8f+cdYIQBkQEJwi4lgV8Ncl8wGrz17uC7Pa9g2XVlL8G9Uyfpej1Ss5dN2e
Bk9tpb7Oiyn5ccRbKCpDRdG4w6Epb6kFBbrVnxjKIFxx1dKKbavvixgSrCMdvAsmawv4bDxo8QTR
WgruBkwYAx6Atsy/S3sy02csKxIOU9sSP8OPMi72Zp9wjnMg+SmNtVqYVW8OZ+toVXwlEe6io5Vj
ki3O+n0UKVy0qbi0etVCAvSOvYPt7HjJBHk7WnkgKOMkCjVwP9wAzY8/ZktjKzxyctG/Vl/Kk7gh
cTI8/375LcwaSdMouukFmo4mgLQD/B/3MGGqR7NRQYuQryScBHlVflDOBikP7wddlTt/A/diIEAS
45REhFLi0FKkU6kbP+hHCOcKPEnC5iZXuWuiVfR7qUISloEi4d1DfZPWau7ot8HWOV8F7nN76FmF
Qru3T0SXqcrmlU/NcVWX+d+xJmlsrIO680/5yuLr2IBrhDgDwgJW2jCbY2FRZehhQxN9lBStBR0K
iQFXmyOhf4/BM2YDN5j74BBg0Da79hgT57/DZsg3kl5p1zrtgT+QWDYNUhixlNlzVg43BICl4hZm
Uj57wpZbKBpiIgk5El49XVLkFr3mDWTwXxet5eMzUeB+0/eubGJqaF77d8oMwdpMAo/kSFb4eXpk
qDyNQj09pgZaKHq+bPJroNilNe6Zucs0G37oRsTCXMbhwsSjMY8MLvV0HigrCutSQWeNvBdG/x8v
14eTX054/yVdcR/gsPBb3loq8Qz2pyXwrXY+wmMxA5ygqqh8/MIuf4GZPIYrhS6lFbKxzDYFwQRG
o2yVkJcaz4jRJFq5zIpVu6cAtR+EEEw6o/PFYcBBdLctb+W/joroPjWH56LcFlG2kDrYGj1h0oqb
NsHKjeL/Xt+bSn8n4zvb+HxORCHOHomS6vycK0fKSpH3LhA7UJd1BiKulYsCaaFksh1bot6dx2B7
95ODJI2vKJD0WgWwp3DleWcpT+3in6ZNYiHlY8CRKphfa+lwzM5oU9zFmCMqxw0M4ZtKXrUn4efG
4q/RrL65wV46ZwsyE9SwmMeNw0RDG5xlOdfDhpybDTm02I6HDnzDcmFK1D/2AsfcRS6k2jcpOL2y
FBHBSkA7ggHekJgNvOFSkv6a9NUD+aLfsziv7X72WqDbHmHj9Vi0Z/4EZ0AyWhVQWRURx+rLOK0m
Og13gb5rDY+hPXpgQWRAAQYG61+trDK6xFIv1n6zt2zdXxGmeCsziQQMq6h9Mfxd2Z+Ct1R5YCyP
0zhGRE+1lUAji9r5+n7xYvzrmduuQbpdfaFBHPbMY1BuqzplTXiqaqKXIu0tQXY+UcKwpzHBVN+P
RxAbG+qaM2/OQ+QhcPpyTqfQ9DcCXk0kSujH278hhMIz+Sh+8rYV370jwb95TEw9BVRQUfLtCFOQ
JdmMkYZ5RACqs0CA5vR88N3ts0uLm3mFsyiaWpqXGVCBwrgaGbbp1vR+8/sBjpsQ8jy0Miks0cUT
bVun0SdX8zMppkDppR9YmuxhZGS7HGIDBxUVNVphWlX8Ut6JB2Ve4ClIi+UQgGzrGH+4WSKUgQP3
9lkt0ZZiLIWdxl1QFTUqLJoE7X8xIljfxHKcr6R7ijE/14bKFglIdUb1Ocz+7ssHWwFkzTjkZjyy
Tj9T24qThm0HQOI4Uf3p18Wrs7LFdSHkPx/FCE5KYUNti1JUQ6k+gkIL+ayce0a1qODfb5Bv4Tkh
TX941kQJ7gM+phn2hlzfYebDvQLNuDbK3h/t05YWT1FmxYWkhh9lo1hY1K1vCgMRiyHO5KjDLjVP
DaGSg12LM8mHGEHpPAp5cc2s3OcPxKHOYyt1ellGw17bceYH8SDrZ45Zj24URdpAF7wP2tE4Q9pp
nPuH/fig56PrMYT0gc1boIqul/ZrsEjw/5QFYKCBsbVrX6LZIRlEHZD7JswFXSS4/LGX1Wo2gQSd
WyOh1RXti/iL/6rf69it9+lkqL3rcFYWLUzbVO1AhDkEFjY2GNpkOoKeegy/O2RTLkbfDl2YMHj5
HFl7aNf9jt0RcQKxr+iL6h123YNI2RROZupGJaOi6+R83fu1EZQQkLlhqMEEosZjugWWnhOG+ezZ
GOTbEu0t6MI1MRSXYKH/s3YNoLKuy9q0k0a60Jn5tci8w1KI4P/b7D1fSPhTNYd0hj82laMyTHMH
s7FmFUbjgNVTbJsCTVfvtizmz6ypv3m7m7RhfAvITHJxM+WXV9Rko7V992AZ2LFtHLw8qvDGqb9e
ghbWc9EHyJnOyaPfBWlg/1BQbOUDLXKldXhQcBcTjjWPyztb2oAqp4jXCCEofzW71K+EoQvsWZpM
PE4nvAlWNOTizgspcBoKCnF1uJgWPj7ctuh5b2z48DyovsGv6VeKEj6Y+9DTS+GUEuCUVUkBIGvM
cmzKgukAjg7WywYMFFSEBHX6KVTod518UlD5bsh09OjYRxM3TT/1evrLgL0+Ce6wC+0hESwF+0Vo
aRYVzTvmNjusT1xWdRf94G+v3uKVMKy3pg3pLKXOXE/Ab1KqYWlnoksjQoXOB27Iat5OnO6cB5Co
q/nP5NaVUoMywM5dag1YCLJRw/BDEvdPeoSid13adqSEmbjTTWCBt10vNA1oKzQU47Wz7ZbrE8L6
QqmCWPpxTya5nb//vQ9dvJC9moFj9u2SEUH1VfiS/Mh9PdXd3mteb9ad8RTo2t91hhZvLEK/HMRC
8bPGNoLTScut79UdZM17A67H1Y2Gm3ecJCtOX542MHrIaOlTmMJ4tVnWwtFUzGm7dDALxsYIRsXN
0VSzYHtRvC5UhBxpkiyQSuBbE3ek37R5PZ3ZJIJPeR1WMBUkHk6XZH/ncJpmBvamL4kMy4iPcrY+
a1cufMQBNRmSNUIw4cXa6N/bp0LaZDHMJAzHCgZh1LAptWcKzxSBBJROTs7CNhxFfVGUdsuzAnjs
QhaUMBjFysRp060MTB/F/PKTdYX/GvpOkUdrITVgAfamFk7tF5Egh/6gbRNkTL2gTY/dWEjpVEKf
eekFKn2fKr0rdwGc1ebulLBeM/N9omXQkclS6o2GD0Q6bly0OEaQxXxCL/8YwlujcQCydNBLOs0d
1Vc6HZ+iauTy0/42liaJIY4gGy1Lr3BXvbhimHT5ar6ZAM1n+zxPJI7Rmb4mzCsqQMt8o3qH0osC
yBn1g0jSL7PCFYMy31pvSDpL/tk4K9FV6xNBy+zTN/r3ChcDyZeZJ/rjlXctti+68XrSJNmJW5gh
0RCxrJ+29MM3t/DxGQeQYteBZ2rySNSiWwyr/68qdBathPshb/+XRSrWT78Sy+/pGL0QDF8mU+Yn
rIO91NoXdX+fc2ponMCKj2c04Ee33//Bva9cXX8Jo9L5/uC0qSOqCaJCqyLmUvKoEQ9rawi7NUJg
SR1x1Ovre3flKfvGLT+jWRRQOsbINA/b4riiREh9E/NByVleMaqeiBdCbDiKzO9sVEUsM6vdl0mM
UmVOcWrB4Bhk4PS3fEcATXBCXxyJyExxMEfF8Ne5cIt9k90HidF7UzCT+BXW3BrWHp5c5AFOTFby
YPYnVUHNsx1DK2dQT8lFg50RX38VFLEqXfzZijbdYp1TljS/W3s0s4LxN7WKIszM4iwBILbgHAme
NrlFQ9c/rocqLJRPByZ58G3DejAK6nwlLWxLWMsiNzHf5M6UEoQROBigomTDw+6DqNgR7PYndIN3
6ev3w/QxKmBMqM3HlFpRFqiZMeJ6EprM0AjGhtaLMH0SMwwVDHEQcXos2qv3prd0gEnWNZakKG3J
Dstga4GXmO6r/+MQyUhwKaPXEjc6dIYW3vCaUsx7kkgicMZI3Oc60up8QbOwHKRVi5nPoRVNcgl1
h8/icmzcetPTGyNu/yXyBpkDEnUoovpl9EXUQya4jVswgn59AbcyfApyJ8uhy8Smlb+7ooZ1g/5/
jbEHtEPtPrAVYUWBGUBgyAw1kyNQMQm3V1nDXp8BpBGEPma/3RoNt6XE15ogqIGbamnCt1OLzYAw
7q46jV+cRKGWvwH67/SzV8UBP4s3FVXo0pnektRgGrl/3pKQRPyE69bYj39ifvA6FsIp6f7kF0SK
/O2uFg9dvqkEi1/YKPDYK4BoO8UKzJgqmfqjYne64q0np0QgKRwQ3KPvDbZqaWg7bC1NmVIQPo23
JrxBjSMGMV7ZxT+cbD0maD3Tvh95Zcjiq5oIdsTO2pHy4wNlHzhzHG4ukMnYZExx5AsL9T+2zaYT
0VehnvBOBjIO3TwUjncDY9JhjuQJ9XN8u4ESYbnF4UuPdZzyPk8Ty2SQ72zEtrIt0uVkcPZ7oqJg
wCnHhxCvDgFJRMwptBoK2p3QUxxirImG034oK99A/mQlOXZHTDRy78Y35xHPHESIvsNngbPtcCmy
HFPAUoiaZH2OKvgexq+zL7EHs/ko2rn5UceJOFNkfpZrmBwE2D9dU+u2822yVO85zDaMjF6sJDSm
JJyn+3nS/O/NVoCNgikj8A7QL4jEp3wVSaaqWwpXalogFYq16O9yloSvqTw4AKLtXK9k69Rd+Z4Q
B+sU6dKmONBqkm15PpdpcK9FEHvGVxXT8VR8FOIkwLtLKilgsIqhJVTlzRT+f57YUCQuvqNOQTIX
vOt2suq7kzjwKanUfBAPP5NIFBR3uSWb9PeE/qfBQH2UV0eMNDMAk8yV1kjCYB0oRrGj5m10VSLH
K8dwmxiizCCicGPSqrKVlKBf632IE91m0mfTqCDDXczTaqf0NKryU/Eug8DZn9S+fxAuxwnx+XSv
gtJ31dm8daepI6MpyssCWCUIrfKSZX+2J8OcdlnlzfiyBZu/9czeNxGsEiv7l8TbJHZDqgjdmsAE
V0t8LSOUyoKnB4Z3K2ZRa4hrp/Y/yjE+CiKRBTSO6p8aOWN19UlQkkPFhibEefjjilKT93pE9lj3
uz1ZxMzz06Hl1xvI/s3lJKm4I6/IDmQUIwU+7jd90hS5wF2njlRkPOjmFbmJmGb8kZXIUNHp1sUi
7dWxugR3s9BiCzjtgH4edkc2ziWMV7A0PIAx/1/nVhlSG3E/C38NyX+E/wQB2q5jIeroJp0xcIwl
H3GdjC8+d5/MQkmTNMIh8nGsxMNjqjdkGy+WJDBI9mGdVQleVdl53rEby1GwZoqkdLYYET3wfWjP
OggUrNYbSToZCp/BO0mg/FbF4UOwHMv8mji58F7QR/iy8BrkXDbAoGSPjIhYFevqYlloZHwfLn8S
j2DYrUn7sWf1ugfmxhvDtdpYx3A0PIYhRxAWBsCIimFY6q4xnL2ggvORHiI+0lFF/Lu1TDEUGNtI
HFHoS4xiLE/tKXv7yDdFhaUIbWS2BN2fDVVEjJ9+kz6cWrZyxM1c1ZZsIQ8VNvvcZPp4E/3NZF5J
HzcD+du1K1YKaiqTxY5wS3Xcxxqv/cASn+XYasgCgSw8RaVQLYI607U0u6OFY5D1UzZdUkOxuuhI
sGkYSCOInXhj8L5quWd0PbBQ9426CD6nZIZ/yaCzQIe2VpgxHLBl5CqUNGM32lMWvSgjM8/tR2r+
uOsNCSJPysMZUFAsilVp3WswqP6E4+GJJRWkjMQGar4Pg2FHN4fHZLaej++2yybSMcIdC2ygvWA5
3qk9hRpy7PVxXY09DAarhRof0M1tRYoglXkdn0AFYzO2Dvf32SN2kxhvxCbin942JVHJ58z8zeWD
4KvYzpWx3pYOP7kurmagUFSEeEYLXoVPjj4ij3IdM0akSn3YxyDtkns84aqzMQd4fsJxzt2eDgVc
fZNUtgn/O6YVqdKYNr+ALpR3dZkJ2ufD4POv1yvUoXST461ifX3MAwbOlPr3t+1bjg83qVwYa1SW
6tr3B0U0uWMaHjnH5Y6+kwKkmFQx4qxwDNTkKj9iLvDUZHECcmmeuyp5b+M1gSq5vQawnaKY4Igz
ZWk+LdytiW69k1LNadrGtnE9HDaZByoUBxv2kLYhU6xLPWucGbB9sfTG54nMGE9aQ8+DewjYbptN
1tcqvJE4Q4+GnpYg9/I7Jf0gYZrylO67GP0JBqfcXIYwI7FEDGhBxOSwVCXx6sHIBjnVXT4Sa8/d
qA7QjmwD+mOr1xm+l3c9zlqz+dLJ7Dgi6P1EmS01KOEyba8vy0U3WhH7Wh/8/2mwQuFxK2FxSvhC
FD5frSpYx2c3unU4BN/kv6568de3CejcheIskoaXXOkj+ouorU7vn/Nb1re7zaSbzNHway24cUfb
K+Pgqf/juCKVzEOaHl45eyKsMat7vqthnHQ+N4TA9YyEauF40tUkE3C7DXu1QS/PvqaauGWEaQmX
6TYKvFLMwsBp4PoDsQRoF4fNUOjVunUrLpwZo+EEQ5T6PEeL7vWuo1C5d00GEQyuE9SrZjIeGL8G
sQL8LjTzBspUPdccdxIi20p4iUR0jkRP8iJei527GsN0GFDZqOU4TZ6FJZYyIlcaYwoNhwwt6evz
23UaKp24o7qkN/Fg3/ZmVD5WFyKPD8vHBSnOw6OEMSjrlgQoZGrQRf2ADbjnpNT/bD0sSjCVbR6f
UMP7XyXIB49lb/zmsR5F9yXr1PO0dvxm4267sHclvX0ObWqUsNekzZJVhYSaqJuPQkCBUV+Sl2zA
YOBsxecEvZcys9UtnxlPImCL+k16vIPn5pwQrgBYOM5UI46roam2MX3r4l12VmIaPuaesFbsq2FP
qAtKalvVhOKUO8/at6+mfVB0qiDsq623Qc6OOFdJFtQwygLBLGGoPzloS8GTYFl8zCD7nmVvzoc+
YCAO0bfVhTGUdmPbvc476ienEaQ6J48UcGcNtbeXhiiY99AwjsFW5PARNE5XU/9hFrfefyoS0Lk7
mDCVPbMPicKlN4dR9YuuGAoOJsQQ4Gk4wrbxhDDwpUP/F4NWJqi+q3Z+7rHJ92RSVoCvLu+iPyhW
RMyg1cVOYWtNPa323976+gCDk/fnp2XVEc3jBQCle5bdni47ah4aPqAOACtYzDZpgPHn5mAmUIPi
Ijk6BRhH/S7i4jBtgjDeAiy0I16o5c4rkMUtYuYyfeJLHR0XOwDtGUJQPKYgISKs1sqjFH1RDq0c
zxJXGv/mmfA/VX+ocBz7OwUVIR1wqhqpE3R0rTIGkTm/r+utS8Qcpv/+ZUXK93LFlV7FI7rTzsMD
BdeMsX3TSLpsKCKoT5XQ42vN5MU/GAxRzWOSMWHceBOzEm0Zihkl6mx/qGBoaygln2jLJAoz4e/h
Cc1/oiSFZd7/RYk8IY2JgjWM06lsjUbXCmhE/Bw25DrVxLHmKCE+Q5zcPDu9BJl6rxIXHkzO+kO8
eFuzg3gFY3Cwd+zLYhoMEfUll+JEwx4rHRRyxEm5nzel8+rIeW6d/n3iPMnq0gFXCyI+vtg7MdBY
Et1IkRgVtfddgPndBTfrCVbCONgOFE4J/jI6sauOmiMYdXrHHgIpfX00GSPqy5KsCErQr6P2jsjo
9zWvyIh5M0WmpJA/7xnpk0pmqu9UrD1ITVlrHZQwRwaSfbHq6coE3nP/x3hfiP3hd/nNSzApRiyt
Exlt7XfunprrrsaAOIREDwUXcmzODSXrgSa4JVe23GOHDA71k7qdtfMn2YQ+9YDA+KeGTgQSUJn9
iAX5akCPaiLuWqtqtGNuzeYuOrqTtXW43vmdbhtZb2LAUxeEYLEMJNM9Qi/u/3PRcbXXxyxIu8D6
dS3tvA/OD36BkCKUsk4amN11vBmVQbUWIxCR6BX3/pD+8fWrTt7Hd5uyBqRXLKDC7zxDd8VngRQy
VhGshxbuM19CQubvxG2FaaA/U0J4aE8qrlvDZ97MueGrlQ7F8a8ZbR+xVFdbZGlSr945H6pfvPX0
3v96JyCdc8B5JWjjbrJBilNfbum1uAkLnMsC9fMIkfsHdfT5d06FG0+OedoA+dHwJONkJdUcJiyi
6rA/yQz7Mg73sYWIw4y2qKAsCVUhGqVu5CZH/8u57kLaV1YiDP3GLhj6zy4FG1K5fJG/3hgzFC3k
6o8NOhXg6pYkXdh1PhHaWR5dF0JP/fXXY1oBcEMlrazaZ8oe6ACLhMmJ88+ZazA66ShW/DkSZa1R
kdKXnZR9u/KQ51qpz5SGgFi9aPqF8PPS0qmLv/wtrYilK1s6sZIteZ3G134tH1OI97G/SIaIRsJM
gObQY73VihR1lwxIKBd7VmBClBB6OlplFxfqdY+Dxko2i6bXC5Kc//aCr1UMkUubDcE/AdyuS6ZE
5DDsYRflQRt3c9DcT0ke6MLjy3tENdJ8nNREylLOvBMZQHc8jn7XMfTRfrnAG4cMo4NpUkKCoD3Q
DQke2VAMxXb/RAi2WwppIgqu81scTUoH6acMkTHbwbB55N7t1Wb+WqkwziY2fPsIvkX2xFRPIKxg
I3l8+fqCh9YqERogUp4t/dIrNneWtXuIr/Ii+z9eBlJV24B1ay2lXRb9mJY4nNCoS2PKd1WxIK+F
+yEkACrrZ+q+xSqjAecS/x6BGJKtUDfRA6U7AC+JZzjWdWS8gwfWtN3GC9OXQshNLeKavvG9bn0x
jqmJ8dMwaPN+EpEs2nJvw56q3++jC1EEIzZKs+r4Jh28T76yMLD5L92nX+OSiFblj+q2Rwluhhlo
ms9Ao/XGxmRTRpM/OLuazP3B+JMBOfcvc2WstPXghyMXsvPCaLLCAJiyCDARuN3mBb032OJCEDAb
cBtoCkkMfPTatH/DVzado2aO20DMn2eQ9k6s/BUbh3vZ1Z/doGwH3m0MJg5sQC8kbtBbzFTomdzB
IPKlKtfy6+uRc4rtX98KiZHUXHfNhst66449hdTSVILXKtw82b80CvArK40lQXFEBHoaJqopAMJm
wPqf+199VDNiAjw8RqRQ35H1MrDXKDWQYOONqP1yaAqySzn7uJL0zycW8T5POD+TEe3dzcbDvB9d
qGQBX1MYO6TWmdINhTNhN7zOfVcTFyP4evB4ZNPey/E38E+4gviffkXWzgKiR9z0tKwYmZrgh+LU
iHLPj6KW1P6x0BeXY+vKZXcLLdzreczFl1w3Yd5RtugYrvNp6UNjibaPcmRlniTfzDFY2VTe9vkb
dT4L3Ix08Q2U6yle+ipLzIvzRnb5LJML/hUvfrN4RigEeG0KpVhIVj/WXsQdAPjVMRr+bchwEKJF
0S61Xo+vIQ71amlT2U8ttqcgRI+UVOS7JsiJyqKPEJqUsS+azhBXj7EKg2hpQnKGWYACBSLcZr9B
KLKS2KYoOsKLgiorrKSNDDL5gFf/7i7mbeHb9P2mQZCdHOvzHazQDtzsw2ZBQZOxvP+uYHyyoygL
G2sPumVPvag/TqOvdVB9YleBF9+U9M+V1AKBJDra/78hnBs8/lB6LiFZGNGrVBg72K+JwE8wtQ/n
AATjel6oEjpv/LsiwrtQf5XvadAWjPe5meYLg9JnItAjHlYwDy3K+xd73jdcypxyluz7MayDoSLH
+g1q+8MNBVV4JMmplgtCepJY548NRq9Erw1lAaiNEOsqvsh5pdMbNIqgTow1Qj6/mjZ/dAPkw0Vb
9Hi557wmx10VVPXIhIurPCLw/hQP83W7HAdD0bM9AQOTMRIW0BdgEMpq9cVClgfY3O2mByXcP39l
mxpvfwtHZhbptYpHtAIuyNz5F3eZ0sw2BQjZ+Bwu3UDBa5TsAGe4W/IWbUoOMpbWwSl3zVj7Lp6u
RYhfObiSy2CNSf65IwVbj7viPrSQeJGahiUY+Ie6rfrQJ04LZyJn9UWKnaZS/WCAPuTY063qsC8K
H/OlJOccuylejeicbM3Tf9kfAjNGLTUFf8stkuUNjwmYgMrYIF2lGBW+hRJEG1UVEYl3eMhjOIv7
qbOvaARG7pZ29Nhjjww4ZmEgXImQXzU7Qo0ZDsfzcKKKRxVQvjr0ROtCJR4IJ7MLkuxN5Znvx/OI
a12oauY52xbLCWcx9yr5ZVcZe14Tlb5CnhlGms7X7D3QFQvsRZJ8U2atv6zylrcCK1SmI1Bi9KzK
C7eFlspbYhpsnutvmVlB+cXmQwF1D3VY2oqn7Dn6PMjqVO+9uhGVFBsI05o+IonMo22HOJQl1y/a
f3IQIBnxzXXlbtFEdt8FqTUiSJS3sHn3QJRLFPky5vhovnRvdKcSf11DR2wQsfv/K572txMpdmDg
k+Zlwm9KHrvQlRc6RZVDrr7eFn01lhq5HDJYFev3ZAJCPWV5jwd/jHcSl0fU72KgTvBuofSIvl8S
2bf556KUrGowfAjIt6eFhca/UKnr3DpvxGaUziN+5R3SvZg2G3/djT0W6iJTdKZTi9ZBV+tHI1nJ
ZnHSqsSErkExJuhpFC3K3mQ+Li38Kh/RA4E7XmOpJYGhRk0NeUELLoe4s2JQOilIhMAVa5Koke65
4sf1yHIlD7726MGDGqg4K6//oCATKkPUekHyC9RkhsHpM/doU2oVU2wDO3WwNP+md4Wmc7eq6kBY
O6GjbSi+dBsu1QgZ9Wa6WzhF2ckcZxbRXJ88IiOKbKCQ3CuQsWGfH953V2GXXbqsDFmCAgd6PM+b
v2Sy8e5ijFKrpt+VAX0DPXnoe9QZ04yWWK4V0bv5pSyrR+FwbTbbVfu50TAnL23gQXNOeE6ORxkb
/sCQFBhQzKFDEU7c9FDaCzhbcb8HtUaqrsQvtXjmb/Derf/qDVOBSwrgDLwCdh+UHdXysPfGAnyu
BzpBRbIiYqZ39u5obt3l1vDAvOgxcth5Vyf9ss0CFbydIS7S2X1Y0zGXSR1cIqJoWtazRv68Jbl6
JAL/OhmuimibUc/bxnD2zdXsueKropSIuWEml5QzSpIElwPLPe0LVviYYjXhIfvIrbcxKlNLBsq+
HWJU2tHFi4P5WT75ScW7l4W+N2UdH8KBUoD3ioWWTpOlXr9NC0mNCo9TJYhq6zAQyMdNp1KM55mx
b1vhi/rX7EePfNrzMYXSn+5DUWBUEzTIQaJh3E58wGyO4eE00EF+MjmW8I5iNa8GIB6rX+n98mId
L3E3tBy7b/p9qop8LgEjmLLhKXSI31JiJtHf+sa5SVdka0gGFJKYhGYLXOobMOTXQbEsy9WscHmP
X4+KuQ+Tjzd33qqSDT5mxuC4eI3hfakZE0D06QdO+uq5I+gE2UeHyjc9dJ/mA9cRPBAKLu9+NuvO
5iRVlqyqd4juMJmg+7xuO/W3sxJoJZZy1tqAU2t4is9v0u3CQ1sG/e3pSXJWenhvr75Ibnp/UD4+
FIoKLXec9wxACZ/dZDpiLczW+ihaN4PDw5VqbcfxNAq0smb8KvEuA8bmGGyFkO5nGz0dCsHflZFj
oj0lljzQ32z6HGBsZK4n/pKnsbGeGeERAZpH+ByUEXQRw+4iYjFS6Y2Vua8lxdmfhpcTYvwTKcsX
WlMAMlVwTX0kFJR8CrUdU1WmJcdanM0ZBuwiNCrtosxdOOUJuDrMckaCoMaVm03VhVqP8DJ1tbaA
aJOF8Jj9bvHBCBzLILnXhhmmD1RUeWAKkFusFirMmNPcLazSITv+KhCXGB5jHMHtdiqL0UwRQFYr
3LjdfJtKeYa0EXFaEIpZwzjNFI3rtQA4zetJws9IgRKrXrHy4OfB7NTIMNZ22TeBvUaoyjWFajF5
ynJ32+Q3ySiE4GEP41Up524yWgCOgFawFYLyHD4S3rGKyHaxeNJLQvaaqiVxCZoPYZKwrIseVBxi
W99cIkM4i45J/q8KYSQyNNd78YsbQB6YihNN/P2xZ3xSEzW5Te8K9nCTlNRQG/uLeGHRSaHgGElq
yVYXciprjYL29FnYAy7WUqgURTbUKtaj9JDkUFoIWJaNsS8at/rbEbftiS98KzsMDqAs1jagZ5hd
FA4ubhQ2/Lb6t2MrdMF3JFSqEZoC/vBQbU5OlzmgZ7287z60CgQFONpq+9NEgNO1nOADJCEZbmy4
1on+FcZlEDzScnLdWlRcEvwa7tbEGc9hvtjy3RDB+qs9dV/5+BV1X/3FVIZ31/pLS0rD9MwblyS4
O6DC9GiZkpzGm9gOxDyQzmPhK+rHWTwLE450Zw8zGQWSx8MXs8wOYKaZq6TG4F5EP8Le9kocWis2
JgYPJQDYF3nd2omBN39UKq0vpRRK1MaOFRWb2okE9MUsMq3d6DkIwpdYEhq3V5r5b0LBalMr00PY
1OJywpDC0Qs8QezGfO6SQdBeTcEQRIUSh9TBvbpUz0x/2rtDng/1zVsPNyS8h6LHxQcz9vaB5I/6
usd3oZdAqRdErbRPDI9geYsif9Fhs+BKfYyl0O3MHkaH92n6I6/IvbVbGFHUKkxrMkXxE954MSea
6MMX3uJX0Lrimk1fqqXb0pUT3x5zaiEOrkxKPSVh8uHIps8YnmZOBYuC14/xeFC5RRNVIv6Pg0Ey
43NYxXZNkQSu8HA//chphn6d2UzS9veX18NTY06hXgl6XAXOpRXOKO7ORfPvJGtz2KtDiwz6wyoy
FYn4FnHtyMMDvFvUY6Mb/iCDH+uD1++5zV1wMiXmwYP1LDQtSODga1u4CTb9TLbzIfs1tLcGu+lt
sh9QzwcStdkwhBfKOLG8TdhXdoG3l+zFoA2T6zLqKOUyHIMyjdPCAYHSYR0EjkPPpq6CwgFBtR11
q77r9vqr8dc1t0+Fv96AFccxZo/Bqfco84f6NWYgXyBAa0DyRZbaXFc+goEuOt42e4JAsyTyNXwG
qDkK41RC58q6G2nmzGOI+8zkzLBDKRFXA+KbQyudHmV8b44Xn0UY73K5exXtasluBiXn8iARqICd
2JWzoWLo6g+SWNi7MHwxfDJSDm5hom8kJ9Rv5pRo9ZKY0aK23iPfogrRRizKjX4EidzZnxdtB2Lt
/lqMImi+Tiz6DP9IzQT47/ydPc1bxPRQA5B6eEL7xiL29QHbVPM/WrEvQHtokZWBMfMub99s7d7q
A3zdLppmNXFHYlPG0bf9ZuTKsxSR1SuL8EcXY2ZYJpPlHdOZ1ZL1icgsA8uDWducthTeJuPuB+BF
AIc1yPAcVCGICALOAeXHq0PaXvnvoKv/rZnINaR1JiZWgfIzArHU+3JgO0xnIFiY+6wvEiakFJdW
NexpGv+5+iYqlEKLQCQLiH5kKMC0dunrN6aO9vsYRTqq37OYBV76jEmLIVVlIrWicuVrcQEkzh/J
j5cxK1X0e2jXhGeSonFxmzmUzy8p0aTaLcBwzvMi3bUuyaceCeSaujTsIt19q8xhOrn/HsTdbfdg
tdS/IBnINeXRjJQDEq1TcE1yxIe2e30rhRuscjy0j0Mx18ZhVuFXmrDWrWmz6dz/AP7Af7KMmrpu
EsOZ95/KO3UU68OClDA4iglxJbzqCGCUC3mjtQbwK5y8XQ87I1RIlFZOeGdwhceTK+2+CfBYWXEN
Xtk59ZA+vFeAEWbkUk2sAX0u1mBtFwfoxRzDxQw0vE3/1DMGd2/YfPKbfpjBCqQzr2wJm0gYoh6M
ZG9FuEbLdwkR53vxm8nUNrSC6R4d+RMpbMwRZGqm8uR0gTvmzlAgIgErlP6aWdJhzx/aGZNpcLfd
w6XMQhHqehXuIsbYTgb2kuOH2nuLZhkhDlWloksMQcCI2iMDMFBtmiezq+yWIBdZgKeDm1X8fgJ1
X2VvGMIbCxRfwU0FDuiYRUX3mjMTIotyiug1o9z+Xh6Rky0aSNVdL9UiBOItaibKxbAGD5zvUiHO
/yInxdniEbBL/0+Aod4RndUVaI49X8SgkZ8xAqj/dsFambiUaOjT254uDpMbPv3xQqlgUF4+UGYz
rSDZ5VjAcLcjuINaTg/EDFq96TSMF0uB99dHGqhmZtux+NU7MbaselsMlBrHy29AMvYtgR1ls9uQ
hHWrmE9yQ03Zl8uKvev+ZYJCm10AEehIcoOmmNhPQfN2RgSf+LcfRkHEzEP2bKbTocqf+xAsUOBv
a3Dx7WSmWmMwPZ9olEzjWeggdmR0jUbI2z0rF8YGQC1+2J7ptucjj/tLtT835BPo3+fQzso4BqIw
xyJi7gEPa36ukMOWIes+j5C/BGGu/SLh9hqrFR1OEvaeUSQZ0latN8Y3B24geEuJNoFS+yAfNF22
fO1Hf3y6jyiCefwttFNlTu5TRF9+bul0NNKWIhN10RDC9ZnqFgoXqyI4kPy1bDJBTPbf3F+ewgPn
R9dMSzXHILZ9EkC97QGOEtnOCx4znrYRXdppXVnal1LesYo4fSCpgY/ihFdlkINiomN6bn1gQgRm
iqMcxcK1MLiGJ38WpUXr4QbGmLorvU8GKP1x6fv3Z4qpl6yaGLDbmVDRAe0lddfArBFGjJZStMop
RYNULuS14G6lk8qoIM96FQnEo10XCJIPpD2VfqXGVDU63T++qj/eNDBshWMgDg6QVobPdUztekqN
v9N25ZSvLi2JSdDxzNWWGp1Z7lH+R+b3KtxEhV7NRh2YixC5D9lkIuBpzD9zvuE39UkT7TnCnTFa
FBxVjD/ZHmPvPMX8qdhoyOtYipcH+/WBSfCu+mA22zE7nfbNtkxvc3NnXtZFjjWqKbl+71aJ1cj+
yxmYU+6jTR70GBN3uWpMIaj9LUE0Ch/FAy8XdaXvf7EjCgvhnY4O4PmDlYmk+PsJgpmB5NMVRR2K
9mkX+zTi82eFzgOVpSaa9I7+u2kFzO4PZmERtybn6xevgU71O0KZACzpll0iI81gvw0QK2FXRgx5
klr7d3C7buWsN1JWYR09a42UvlO6rLai8zTCaG9u5gYQdlJGs0Ie1QREhfwKCJJUurPs3VJEpvkG
rv798GPO3UiyWsjZJULXZfwEXGWduJSmrBXZysDnnZS98J091Bb60tpduUBxKyz0/lDIlTSrQOcs
a3QTrCBZjx3rFUM9vIJJ2kGIINAKxv01DQVgDdQb2CgiOjrF/thQO+gYRfczabE7BnjBs4qC8tIZ
EgubYqf/3++s5+WbfA/8uK28cWXQNlEDPwb25kjAqm/PB+8UiEDVZ4xYOulout63WreYwWsOSlHd
nC8akSay3nm/GvNVGicXKJAj8VuS8JokqL/pXPYisXm0ukFkG9dFzbA4crSxKE7VSDQuDtREvtSG
HAil9LI4E9Nttu4r8vNj/Z0RmPGGERT7FzUcad7Cfu9yEuV/7auvqCzMxlq9DmPb4YAqxuvA9nyW
pRGI/w9e+wvtF3WyfowRgD1bzQjouiy1OVjQmmC+brSbs/OI0Kkdd7fIUY3uqXs53EzOqKXyWUi8
mgo/FU5Zi2cO6GBIOg7vUS+K3tOoDGAv6CnTVrXIMnBEh4gWTWmihPudVITDeVa1lTfheTjGEMhg
l/g1F89wQvz1SZMy3rbYF8pz2pDbZiRwwRPMWDe4TcLylxSxZLC3v4Ty/vjhMcvleSRAbESJCMrQ
AK6sT7Vlq2YjBJQ6KGdxLX/Qww58KNGREanvddGwR/WJgFFWDigAzMDJ2EogGTqVqF46ni5gmZC4
uTo+HTQs7qFoEf2l24XlsqMprM/1DLOI8E5KrhwBS+G3i3BxxMLDwgQsV5e00U5HlohFPiCP6fQk
KCIlOG1YuWQ5/nZxqBzu3bMUm20OibRgF9oA4ZbfcB80GqCOfvgMoYT1gMv8D9s4qubHaUqfEazp
MyUfrzbtRQBoo+uUMwZaePJi+kTtFDQOq0ytk0vdLn0fkCy1+91reeqJejdnY7mV7UrpN4m0yatx
ijUpW1jJniyPbKgTglj6zbQAxMJ416jRulEwuOu7Xetp14K+GlngzOrjlG2sWeLoRBMAS71YCnqp
J8VQekkAACabNH9BVhXNT5HHCbfue1JN2uqiLn66g5n1O6zb2iAqMjoBFLeg3deG3z/ETYVhMrYy
qAuN+CKF15Yphnebd57iPc03cF15w4Lpngf6M9GU1QCrPCeN82+q1kUu1lDJj4luW77ZJSLCUenc
E1SqUuev2vnnAFxDRAU24U1aRNd7jHHgAFwR27RLHsRLfpL33XjempkTLyHyu7OR72OtGnR3JxlF
oGJDqc699ZLTmDKcsiAEiUvf8jJfvTD3dw7PtVUGmATNdd1yUIciedxCquFdM930AszvIVg4ZzGa
wGMmg9XeBissqAmdb1IxXz2R8dTTcdzsx+8oP8fD0gR0D+lB+j/wOcAWM7ORjWH4ZRjKIobZ4QT/
fT4zvD/YRJlZByn8FSMzf8i2VPMWXMT9kle9rnDZ6sh14mTpH3vxLvHuwMTIYWz6E8kBa4VljpYJ
2tnQoHibB4s2t7Mffck3RMcm83eo57KrEBlOQhl4+EKJwpdgtV5FYt+wlKZ8+GU2h6N4jQ4NlN+e
JjuiCGRhOzAuNVCzx4WNR1I5FIvOKL12ku33SMVCB2ijKMG4HXowylN6Jav8IPm4dH78XnHvPNqa
7HGsxJxJuhd3E/L9voljILew8ixsGWHSbf54X/0Cf79H/tzZpV3Z5QQACRQ/ALRJV30WMcB+KIsH
UlwKlXWQ0tsG5Zmq6AgseJxIQGDUgvXPDASf/O9Rk/PFCI6qZTG/3cfhMH/xiGB9kS16FOsqUSoS
zvR9b8ccIUmkhVoslvLYWAC3fM+W/LbbA2vyqMj2qCl706oPd9MTwuntjC+YIGuddbY2vGXPhlpy
o8R80ZpN8m9Uv9646MGHEs39/OYWn21KwGYakrm2Agr57qV15cMsoWLbI5Hi9RcrT2ybIK06AwwY
xMjI/WSswBgsRW3pzG2O5FHhZbTwad+0q+7aXS9TdUsexDtuiKk5nYvAXnviZPkXmDM+AlPO0b2j
b5G8Doq4wJQXrrp+mon33NC453CucyXEPSIf7EKwS4BOFDPbB26XZ1HjT200uJjsQHgjRKU4YjCC
lOum0HzUi+TOHz5FUGtiM9lYVYuj2urOXN4CSUhDl3f3+hB0c6LCDKtyJV8AEr4F2YCPvT9tHg7H
3YcscyNvqAlPmDpF/O/zelwJNyvr1KF+26p0evP6iGv96LmW8XIN36o+9FeiWSaqjDRru2AIfcgJ
/TjJ31iVfKxXx0zNia4bu8iuyx4ICYEmlYInlnthxLo0gDYeylr2WhfpFoyrkl6K/LTRUwXhPbwa
OA8FKIoNumCa10grYLyS2QOBV6/upfmM55HwiiMEHNWQYsixq6Wm32fkkg9FIFMnZGNAZbpcGi4I
+C/7KBQEruOPYKzA67NuWCtEEbPnfsIywW78KTSFhZOmPLZD9nsOktuLuhPPig1mZ1UuMY5y5hhB
498HXca8jkm5GzFEcGJ/aQpYqxqPKsqeV9S+lTK0mrfHrcTUB4/94RyeQ72PZdRAVqGXWB5P0zQ+
drA1yQ5lIf8YvFNaMJ2AfbBt7jWNYUyjhYxMZU6szEyhGGIkTMb6ybA/rHMmwYwByYQtOrdpzC4Y
7mlqOvsO4MlFBC4YuxwgenpktkT6snVQ/Er58JYs6HXQMMc0DS/Bxr+7cuuvUYSDqXpE4NyWZ7vY
uDgSdL/kQRR+nrjI1o8TFDDQ00Qn63Oo4huKBIKn9YZn81SxiutLBtY4qhDQdxlXV+qV5+rFVGUy
q3GYwNTRN+qaKC/DSjetQgVqBUDsGZSQi30pK04TbQ/4ImoRzjrWcnARwjOkm02bvdkZWe1KnvE2
cxssuj0bhY4XWWFxRAZhIXXrfbqiZSrqcZWNa0dV2KVJSHPfYvfxIJvhY7LeHXOgpR7PU7cbE44r
XmsAd4lQJZuZzIRk4SdWDM5J7OUyCm4ewZgjoDez8gYNyvSlGbzrc0RIQrV4dk449b2CZTXe8zOT
hgrQe+87JeoxHD+UGQ4KNo1HoL426qldYGjEP++SSjVthtqmawSnviuKNAlvNYG6Js+2vlqOGWtg
SiKy0ig+NUPQAPPczRrhERO5eVRxweb81V0cxPm+f1AbBmD/b5kjM2hUnpp32Y/it7xE+jBMhQ1I
nkKnDnfpZKRq/XlJf9naShZ1h6TIn0K96Wd4NmYYEly3R2isS5KIE5Xm/MyKFSsf9DtYPHKa6G7B
dVcy6//wEdDeUkKWlqj9pZLEPrRom0IFL+rJbgn61Knf7b9K1vope7gpqWOHNaECeRTjeDE1mBA4
1XU4bo9btozGSUGCMco5IPZBLmnImZZ2POZTO1EXZueVlh5+UNmNjcPob5qCmcsbizuG4BpJlbMT
zFBqpyj4Jh4JoPEBTWSUGBwpDcI5Rb+mmbJERgwtUERSGuByYAYhbFhGTD/RgbHBAeq04pyi4DMn
B4G6z0eXPSsXwVIWlea+nQ9Xx2sdrgI/Trlg93MrGmR+9JPZtB9GYcra/HthxHKu92dhsClyncLl
pKJZ/LVRlzzvsWNEDN0Fu0pJmVWuzRv/ddDy+YVrqZe1aJqhnJDc25J9KIAF/U9Xmlm4ne8oQ4G6
xo2GRlQDCZRLrTZFo0vZXkqMlj5TY6hdtG4vr+zb+YqXn9i+b0vaiARGQimRjbWEseakGVWFZC2i
B7tuJ/P5cIVUxJkf9tGUhwLWfGHlF3ygJKvPJ6Xxd+JDnHr1BFGy4pVtPWRJiQEpedQhtYnzTIbk
oydJvJJIkepMVQt4ZA25grZXtp9fc4u1t9RqKO43iC9JhZK8Um+9WylVYbFLUOKHlDDlfwmbJvrx
anFTtkdvpHfvEV0SNnY1R/tvzGg/go9KLyBjf4/Xr6IF2zx51n2pmFBBGUvs0Q+bZVlDYdzcPtTo
6NaszO7bjWpt5LSYC6GD6f82mQQ1zCHyV7hcyilZ9iIcCB7OreNO1KsAOAolT0zf3LGr12Y7GNQD
m0ajsdABSBhYjMHlklxyelf6xAZseQN4EyUxXw5OxhttcSm2BBUFpEDm1hULioMiLtlKmR2c4w20
0SXxkzt0DngU8uN3dnVG/rSkPDaZ5kGWDMDLbLVnfl+6SWnjaovhVJcW5XcYN/YF0lOhnCXHU02U
bPLecRKkfC95LQwCotSqB3aLCsilcJT4tEdxdQVQQykM4rRxRYKj/CBVGgbYLiJp2MhMbyAHB7sj
yAjekKWwNllIjJCXYIm39knWz/Ix0SRLoj3z6Zj/dk2jsVYaEU3nXUeAhbmyNO/VinLZJd+DUKQ1
dwbMCaDHuHgrR+7IkIg2vGAosp1r49fT2XAKKJbn3DcrPruj6rca3rLeZqC1e5EIRrTvqHmyjSpL
lCSvrZ5tK0pbHtJoO3SwL9/tPjUYhHEEKYHXLcEROYssDDtG/JmQFBwmoTKxGBQGhsIyJR49hUSD
wsn7Exda9v8bZax9xIjDeJ+6vMGk+5AWEaSEOlhhurtHthSQEwqomvDKCt6okmo70Uolfbl6O6MV
73yCjxr0CKtbMv805IJjdJHyBQcLRoR8vQTdNhxcnPueO6ORM/b8a7mMU3KS5X2lSjDOnqeVRZ31
tI8dE6ZSdVPBIb/iqTvv60/kfLgZXhcm/x+ka8Lxuc7sPiEkaGN3FYkTi1nrrQJYZGYMKfDs/H65
my6DOjcllonr0Afl77SRPzSAad14pNLy1bVDJXKkEy8ZRX0EDjNw0mpcfNePaE2FXTKkqf4lyuFd
WPXFJSu0HdfkMK5JZBH0Sjy7uUfiidSqtN8BFIqDVQ/BbKL7ulC6cfz0uyFP7XueLw56wzCngueb
ZASJsVhckAbZRWzONsTwYGmiremx5sW7JWbkBcNVVTZFDqS2DM6v4vZBvfsQ3gGRqUUefrJ+yV3p
iJXZQZ5oAh4Dt4TFPyvqbehA0yMbZwub9brj7Q6fqWo1pJtZE8/HR8hxEVn6oT2a1lMG8qODCkQm
VCrdDsexD+WlKLgqCefAeRxT1qDhdw5x1o2fLoN6jtN62vKLnM6XfXxfNcrGzZAfhp07wtZNCCLh
VtfwBfHAhPRvRzBAlP/bAwVBBIsqATwG+YommL188Oa5cxfM/Euo/N0g0CTiMhWN7uEDfJ+SuDhp
5XADE+9ki2rhIrWmvlZwtHJkScvkIisf65Si4EEWTowv3L1py8M7hjNw1MAZJI+/ASydMuDCGsoB
2abFYRKt0xUOSREicowZGw3b+9bIrakxSaZVePp1hxzl8CiKlINOfKbtoUTiNzmvLzoLg+4z/Xzp
wZ0YtkrcBU+RpOEeAE98ZbKPlUJMPF+bkfUdqxpUUtwMN22MmjpErkX8C4ztGZQ7TtjvuKjYGm7o
7xjniZ/NEL6XuEH4PC4OFHFMZvRXlUwJOMvIeFrBbqc/6GJnD1bdL1ujy/6kBHKZqlbHp4xmLq8N
E3s+cxG6buh/GSMxYbQfPS8nPhBogA4Dc8h7wIDtgXu7L3Umip5TS80gTsQjRXI1c4NF2KDrmlv9
GIbpj4TIdw/3BxJo4zXaV+pJw9AvsdgNbFMfXk11WiYTWQgcK0RQpURaet7OMH6hlI57UlwXe+vP
hQGqIypnjucpa7/3qun5UU7J/7qt7km7ZLRlpaT5W7CpxwPTO/bU7CVUXb3/N4BBeR2ABQyfjrlD
eAS/ukWOF6oj/cjuMHOHN5dAc99s74pKiTR6Y8Kv7XMVPoNf0rBH3tAz1bCmV5ovzbx2Sfhu5W/y
4UPtwbUTkqdXkd4OdltsF5yHPpDv15Xd3mnnUjyvKpkClq1jzGeXjWwfg9zey+VUoDXWIwNXjRlP
XmH41v4qj2uJIlZuab5nBYB4v7KCP9/Tg2VZl8J0bFDN4dYg2S+BlVXeyxFUyZOS/pYonCGoKTtH
C2JkXv4xGh2ndtYgsgpkE6nYdDM3qYnGbudeXz24egMZ65f3v4ELLvVQPqHnDr5xtbuCMqu+w0IK
6RqXBYwgtP46kfQDt/NlzrRSIYj7GrliaiDiJM+R5nS4NpDWpOkjAiHfoT6pIHLewn31pKdhJJJs
/+lmMBaS2Fdx33n4dqUnWlrBa1ofS+J5ZLeu09uM+G9+jE0bsBAXWJM1fMdh+edEU2IqJoFfLh6F
twNWxTea7QvDajMv8RtQ2iZxzzvajGJ7Hw6x/nE8qdymk0p38pF9JdCHJ4R2QyyE4z6kJTPGsylw
iy3OpaI0lOoLPx70Xedzp5gJllMsPQVX/DhYGPyULAGKJyo/13/Mth20suaYWIYz9JTIKbYqofNR
46onhPERVoZJMVbPphzXguyxzBYg+82FwKdh6tJjSc7NUaI5MjmNF2byhcgbzJYanKpAl/NSQbdi
hXHpJ5PbLUQHR/EQ7IU5BlrRPRK4u3uoU97bFup+DUbH9oihoZQs3Vs88IZbmsNEyX3+filmoWwQ
1yufr57HFj1n9yfzby5odG4MEzZLuwEgpqvNp+LKbCfP/g0jrWuUQJnGIPHLYoFWKutyMU71BbLH
jgb5YMNwHCZg7k9ZCi7eESSP/LT/VeqX/g13S+t9j8WiHiY9Om4Rcu4w7CoeG72LvZV9DZzlgjle
gGK2Cw9fsArHSDWcXv/Bb7suVSJbbQo8ZgaHeuV4xPNxorgzsL1GqUtgKhaJKh3TNEWlVAXSiY03
Oms090PTvDaubhmyYO1lQtYd1UW/Kh5jLtgKUmGoLksOMyBf5UExU+p8R1ktXxj2UeqzmvdhpGIO
FOaS2HimFW0sIOEMcTVXLYdtswbuhwlKHdfKZobe2v/Ruetl4uMlASx/fYXQFn+99bEDgqdkCETo
3/Tb5eLLg7gagXbIMye35KQKt5yfryNxyX6tM1StXHPzyEIcUK4oeQpUhcWDzT0Gt64TqBh5Irfy
FBr0oGhd/UuJ6i4JEtKwAl8WXbh8USWGuhGm9TYXjlyhQ77ACRMsWZ5N1Z67TV+bD/k/EjfbWb0i
DJYgLYvOVGUYc/eE4hGXvfl7NXho4zj6EUqXnSa9Kp2jPPYm+n+y+rbVzZ9kd+WKoAO+2MfLna2y
uLP+Yl5GzDOiPj38gUIsjHqOpGLJcKnqdHR0AX9hg1zku1LdYXmnaWIhj8L21fBKGuqdRUmjhvYD
sSjGljEjxPTU4dApURyzMjI+Ikv9e//k4nA6bqdO6LLDg7XcXoTQXg1+Ei3asbnOfpvcS9HC/QUZ
Xshhbjwj3qaJVg0baNDxZoiKbL76aT6XymqqhJahFg9BPstdBpnoZL1T76+P7wzTFtmHqAJQKZCa
WcZI3sD/lpz2iRv4o09bPhPdxRKg2ctQmFKBLrrM3RhdPmjRcSzyarb/mKlUxDonLYQmDFx5qG4k
zWCIzCyc63mQh69toL3Ii22eJO9FuNeyieofTM33gva1qCkLaQY9L6k/PiaRsDJiX4Y0kfIUMcGW
koCzl0ip+Ssxh6muVv4DlbfAp8YVpXKFEfhGCvYBrK++oVe8TTIEY+WsSH79UpmETUxDbUPubMgX
x8EoD2lm/wdilnPrsvHGHpb9NBlYldCpxPEZuIXmos6jLxKNo04hE/+dSXh1otOpnUZst0Q9ms84
P9hjfLzyzhOOPa1rr2JGFv1sSCMVy1YzSBt4dSe5EjKzPfILPvEeC0QLdMuoBebeLN+xYYbT3RvX
KLLXtJJlIOUBow2OOeL4Hmb1c0+qiu9/1EoJOy1jFzH+aX/HWfECeECXduF4/o/Vw2ICL2o33O24
TpSNBjS5duM0uWCBGrOe1E+LpN/k3SuQrOhZIfBca5QPd4vTZVRONHYIi00yFnukSOOfGLTybrZi
agyjWluf+4uIF0jtSFCiZKsn+AQ8O5k86l0XXjoqC21mE1Htl7j8RyNwcRYMTt2vyTXJ4teDsMAf
8kKi/qf7qyx7e+XSM4f+CxiCQNkP97zALQmj5QhIOLAhgfwe6PYSST7VW5dibTXshx66qnENxZiZ
1tNkFR1S/2E/AV+N0qx/gCMFjeQ6o/SnD6rM4IXCdh7m8mZJqcF5CzXBKjbZxWySGJ0AD9AfjLu8
JjJXeLYHwgL4i+NVn+bK1WV0ML4a0BSDoiF/awD9HHlnQQXfY3/j+96keBkNlnWXMYpqLlM9sOkC
D7gfkC/TdyRxUynYicxdxgOTPW+N4Mctr2DT3VPGwiCbPP8nT922jid2GlT6bIN7CcqKTXAlpgJ0
Hik0jF1n8oDF5Gsvho7aCy/z1sRPzcisWHFom4jtHkBuvoZfk/sFLfOnb9QWHbtJbjvvczUpvYki
Fa9ZXlzNapO0/7kYXwGo34y+M2PlPLBFK+w1kltl0MIBMEvZ5N7iXJhzog81ENlTwFxsZumgdYwi
oiEa+M9TKjQAcr0HN1LInrrlKIRcYpdSAyX0y7daXne+JZuLXZUElMhpv1y5GjdwOZtBnotLnksc
zfzzljW7XCChrrPEWRIumHD/D8HfTJAaYi+g15mvdQlx2MJ6TMki9umm8cRWrDU5h05FlJ+9LPQf
Z/ebO8ASg72SrA9x+Du5aPB6Ow0KCWyH5rg09AZOyJHDROVs45i6lwugae+9NpJhfOHGWGW2mim7
4erUIY4mSKFxLow+ojBFRNiJbfI3qp1rVRUAtjPpBZ+piRW6BAQaewpAnjNBeS51d1mioCLCscoD
XT8jKXkYzK7752MvNGbqa85K+llledrAmttoJsc4+XnRhm5TMiSkAS+l/YD+HjRjz/fawPpFeotS
F0LlN34UXUoAPeVsv5kne3dUjBrsxIz1uKgvkSfC41WM0UI+ZpF6/NVk7v6Emobv7bVQSTnYJeJo
zw1LX5V9fexTxzcSn168bOoctJCGmcIdRc5bjpsgCRIR5AmA+NNvNrS3m26ch2iIOdIVJQemK88o
HM4PpGgN+IsxcUrC6Au/okgzk4l9MdbxEk5mBTa/3hBQMHDNmxHF5ohuZy72lFn9sYn5+sdoW47N
FXbxPSV8J7mlPjW/uMEtbf4FCge1INfntwWRleiVpGdwiqh0fwMsRuhDF+6w/dviIm7hSg0Bm3bc
QDxbpoIv8MKBWs9seORaWurDlZmUNrm2DpVImmNfcj26xedaBcmZk5XJpPcCt9dArYFRlOLQ4bDt
twRA4RitBW4t4HWNO+H6ycMseUr+eB6jzGq66ZTn1ALTJQKe45s1YwGN4qQrP1rIPUiW0p2h+noh
mdHUIg/uH0ukikbZqqP/qcJ+rnB5dQ8I5hHwMsdleXFPDXII7ct2joB0e9gosrtEePGr5M93SorK
rzCpxIaXufqVyTmm0swawMf2aNwYitdj9HruK9QaiY0RYGX42+AdFfpRZiRQlXOOeuA9bj4vSwHh
ZYMYvCQcvmCG0kyfeJLaciI96e1YtXXfHp8fWHtqhpmBdz4okkwIsBVZTJPzO2JmKqUfGg+/4qiA
MF8gHPowVkZwlzqJtxlOobHpl/mnRQEqg4gc8uCJIuA75W0VYCsDVAfgiRVds8Ub6vUE3/V2nF6Q
YScVda4wXGEWTFw1xEdO6dAzdtbrwif0CpED0+1iwWf+/QTuSbjGXZO7MW3MdSiNnP3VeiMcsNc3
2HoOecBxNnSW+uJ5OrId+eN1ZFiX3WXBLDP5jRWlB5iAqNWlpyyQvcAZ78X9+5cMBQATqVDMI3n3
8XvoTeU6QtktScnzo+Ns+9qUX92y8wsj2n9WBDZ+XLfWTocbujzPT0z4SESR8lcaki1Qd7DkoWOC
fnH9SptdWbk341lUpOQYgJxcNyEC2yOOtKgQ2FhrBpRMZ2YZlmywOXxLd7vLVmA9y53AT+/I5seJ
ojbLZktv7SVcYwdTDNpNGhfh51lovdXmhg8N7mpmSt5G63w8XyzvrUAYopg2nj9oBDOMpu8MenSo
LnZe3oZe/CXGIUXi0+HTBfQtqB4O1ilVK2OP0ifv4TvsQOZqThwJB4EgosEizHZxqR+dydCvB2XO
4j172tuvYf/wbYiJPrKOQR3GN3v65USfzHHFPnOXL8vrKWQTBk9AzYSikLa6qWTlodo65aOPJ676
cmivXkeIqE1rRy5NzkT3CSyEYOTcKCMa9JevrgCasZgkyu8kzadrbW7K8JkZE4misiKAsvAwy76Y
guNzuNRYK/dWneZ0EqRflGl2FXKsk5excvuNb4EhJNH/Ctc6bz/YoGLjAefqQQAsa5NcHUXcbFbd
C4LE5G/UlG1J/Q0/XTcMvCGKcscMKy70K9MvNpos129KVmQClhZ+6v29Tr/ssjG5YLl6cyefEO2U
br87VrTShTb+L29usSxyXp5KMXgrzhzhemIrt+H4Tczj7pGM8PJ2+H3h3p4XF/Nhx/jCAFbBhcWv
3B6NndzhOfH1X5gShgi/1KUV6+1DeCluXyxSgkeLcLBhyNiuU/UltrvRdwRDbLxEoPEajBC1jtP4
08pkNdyI3pPs8J2/4CLAHSG8dFF2ctv/qjuMwo7CKgloHiiQL/aoiM+dvI+ZXCJM/22d2CjXaJZ/
63+3cUPu/BhXwrB2VCbwGIz5/BnKB3MeX5G+nU74YxYsteOXeyIcDAbt+co2s/8GUJSTSTdvhVAh
xkNuYl9LcF4FrgEkFTSdfCFUWhxtqRLKsFs3ES/qvpyZIBt/0h9vFZySbJaVfn8Y3fxJ0eN/6csN
o6nvoPMzgFEUCNi9HHT1JjXiLGQ4Ptt7XGHBlyPRcoijzBPpUi2b8WnGiu9+qtxG/9az3OnLOM75
dVT5OYVRyJnFx6cHqYR2+/+mjhguiLJ71c2AXLfHRZGl/Df1RIhV6O4YnDE1wB5T3h3nWb3CAqb8
VOGD/IeH7JH1aqU07pme6X5qs9x11SXuwVVqOaAhCqgL1g15FqC2UBTDh7i7BU/v4P/HDTXcLZna
Rd3Rz9bYPn0eM8luAM+O/JFVqtQRkeSNNyCetp+S7Bqo2rNhk4OrbzAIoGkaIRR+RazPMm3NMuAu
lGK31QRvaF4HuPASqgxaMlRcKPcdEMiQaQ61M7369+pFSmkT6pDPDQXIyQ0JNenrQFMg9EaAs4w4
d2ztXwdNgpFbapaLGp+8Iz2PlI9IUZvJmeH4X7kQGO1Xv+vtk+AhVPPdkxNupqM8KbY41biktNE+
dpdqsYbJB2kXNEYh53T9/bs5ooaYdfZtzYhXMvjrCCRFjyzZLaLHLsNXhwlfg3Dp+ZSBjtEAZu33
iuoo/GZlAXl/2z5pB9F1d7fmm2ybsraqBS2sSirsMuPVVLk2Xpb4vVzbcB6v4dasgHDKBdHDS4SN
SwIHul9xehgyIzeHyL43syU2nfQ68pL4EjcGIwIKKg2XxloYg4+Z0qoVstE/z8fOlUWA51UtgY5G
8xLYUlEeMZun0E5P/rFs2z8SVOxmLKHSctLXCD6+/w9b+TtcOzMxjHOwno3zVx3DMLSn8rgZRdcb
Rz6wxy5YQK/WOt6GS6+QpTZ817LJApKMurEpZvxiEMW7wJYkgofS77zSkh1nUzQresArXynmWeM2
ep4QfKZOx8/0oFS6E5NkbRD/uKd31KErpqBdRx2rRcGljZipbw2yfXN2GSPJlYCX9O29PE3fmyM+
kq55KxvRyjpNmv7XbbUjjJsYMu6xluDD1gWs3EyykkPRXu11anUPlaG2+GQpU/jxO/qgmvMocsi0
KSc58/U9Hk+ScaJIpAw3OVXGc/auHn+KH4/lZUav2ZXF73a9JwkKjyv4pO733D1GgHoemoe2dgA7
VmzQhUepyMG0cA5ee/YbTc7G/7gJWyiOU3yKSB6Z5fOXNW1IeRByjFbo854odGvidc2x2RC79Opr
fjDX7hrZL/IZ7FVahaBiOMKajx70S8Nkbtib/WulL3ytedHD2raE5lEc43gg0QZi027zOZHQZ+5j
mkOr7C8/C7kwG8r9DRwl61NKDdRIBkxNgKrXk8WE6kqm/f1l3wLxz38s5VxKTVrQ4fqGEKiwNjcK
6lA6uPOTVQDot2cy/fhzT+b1fN7nWUSuB4tLGdBBxj6nJDDwhfjDLknD4k5HMY0ak504ZBoPE/FK
2XOo5MCwoRV7nFqLVvDfS5MSHIf/p9pMuK5SNCw0wbRwV5l7jY/rsIyz0bcFyWB+MGrMtEj74JRv
REYBgVEyoY8GT4YZD5kr2x0ez+xRL/LSjQ9sOTOQieviale2Q9bDUcgWHSmzwGUiGV1JweSGj4lk
zDCMh1qNlF7xbolaTubPX0i3s9t9c5bxIlmlThSJ8pyV27o95ts6MOk1jdpptvvWpaVcH+kPiCCB
fyO0uxoXXIamOZTclWTYzCMUGuVyHnV4ch+bnhfHVknuAKowgKazjJ7BqbqZJpHDuOxtPQKL93le
m8TIKm+GShuaxg4Tv0r7taMD5Pn7vfjUMl5l7JZlFl4vsG3XL18djz8NLsSfrdXI/ZH7WhIoHCFX
9WsXvOY44UJEYbiKkBzop6jkBDFG9SdKV4aiWP0GegKlYwyPJAXQ7QCacEhu5JCg/GyIuTOzAt4L
gMOfhRzmxQlcRj/6TIdhfHnMQs6X1H3xOO+c+EvjLrVKKLkXwWZM+ubswDWrPL+4Xa81EJhUpdaL
rlwsfWDJmpQyopenLYry/GBn2e71SiTrOL2QjeoUT1wZhHWeAvVxAyvdGLkPcGkHSiuqTATCq9VK
vfttjnIKbHo5l06Ya+64rZR4EIypwWlsZcSBJD5Tk6ALcS0Jnj4uHfG37uDUIiOSkJTgzA8soVq6
hf7RjZau8vqVQRy9D1XuXPOiQHRH1P2OpixWmT+LDVWskcXsy4QB0d9FBebYATwWjF4xT44RyOZY
jEp+1EmwkvHkFZ9TXo2n/zOTjjkYItXHJPnGhF/nU05U4Ad6W+khrVZ+8hJ9+Noav0eSX3JOO6fn
6fKAD+nAopdQ7hES6g8D3ZkGA3ORrWBHwmyz1IbwXQKbQUDWDXIcKcBFevwAcLrybgmXdgs3563I
1FAF99CpdIqi/tqzZJul+3KsLtcBEYvek7DNshg0migLO5/kaZt3OPhJuk7Fs0dLBgSR2yjY3/Rg
xL0htMXMra1I1JBryR1LeN97TurGWOj8vMqBL1tZ3QLEulnh3KXHg3tHsL+crnrZM6C4m9BYQ/u6
k2THNEy2idz8zd2YNK3EEizcb8sQjoLu2NNoSfzZ2EjFObY071sysQ+IxIPpwveZVzHgXnW5QK+M
dFILjyWkeCQCjkOCqOJR3987pMce/nNE9vQverf1NW/wF/WxoPiF87Gd1J6RibtwN/oYDYzXhvED
3bpvsEljRTc3vbr2TkTTSHhfoJnVYJpR1aO8DTXC+uECm1yaWCQvA/lx8qD1i9ZSlIETZR/yl5Vb
EaMJ0FuL+BC4/cLHEwMsPRXiwaIWpgPnvz2K5HeTcUZi4yc+GcmmT4u7zjykzw1UmkIy43bUXzE/
SZGsRdTXojWbV2Xl62JiopL38Pi+AnsRjwUulWsTnpGCRauMxJzANu6CHyOAJjs8VlMS8Cv681fy
WC6i5Iyaw+F5sgmZKPhAkE0KhNzu+Jd3Ae5qhcSQVzh1jPi0o0JTzGjCR/bo5lFb0V6L6DkugOpl
IsUdnZbJFDsUduk5rQlJMDYw0OqPsn6a8R/gE7bcMXAw25diK3NtEutf2vBrRJeb9ARePocRVvuB
dcByJQ47k11QQiLHXo8b3JjeFpeo9VHiwLr3+hP+rMHM27zJWSJwPybGJk0zQXxiyy3UJXNZhrzn
XLQYhE0B0M3gWDx8gP3sDi3XqNcGCrG+j/+hNZoex6ez+qk86Q62IV7ZOR+Y7L16yPwFrpQniYgA
e9NzpB+tma//nXTgj44V9UIulj35Y3LFiJ55d8nEgjTjncSqMu7eoaE+S0KoVCMJAY5WbozOX7W+
i/lhtw+CWxWhJwn0ssZ0GvQW28qoP61bkQ011w0Gh31lLsASjUTdki8pjhNv/QeueaVY39LtI81c
gWtEVwj3p8oJPLeXMCWRU939/KkWMaiL+Cykqyjy1txfNxuymcj9Lfo/nWVvV/dhZ7H/AZn9bdeq
QI6wf4eFXoAqn2Wjvv4EeLPfOjCZ8PJMXSppIPwxeWb9a84rzmWZEwg40/vOxhqyMtMlHdt3k4fj
njYJ8njKn8Fm0X2qrYPF1D+HM7NfnjCWEPsaFeWyJrojm00b8bG8rgwhyZZIQVIlibaIZsIz+huJ
HHnTtlAB4eVRvQn+RTaXSdVhZHj7HZ58ciDcqt0pHZTfIk3zMbrBcB1oNtjnu9SnqkBI8VlO1+89
UDrh5mykQP3p0pyf7mGp4/dLndH8W/QE8EP2DSlxIDMX3WuYKZ6QlYaB+rqrvyD5SGO8BejUgaXv
MMy13jPXPThT6UCe3zVRS7Yrn6+Vu0oYLdmtVEXZPCbQtFFNQBMNQRwZAaXfH5uwVMp27nWSvF2h
u2wHDJxE3odwRRx48Bh5UxEV6FstlNEk7kkMsCvNcw3hcdqSOkjR+5QT73lzWMvUU8uCoKToTcO+
UjRXC9ujMwGW7gE/cUu2jx4QWjPT4LsBQ72Nng4sb2ZWL+hnJKi8bXg1JtFkyXlJlQKKZl3nkASF
DaHm6PUtqJAnjljLIe+cprfxXUPI9JiXBY19WgFq3smWRztmAJpA3cAhX7AARs9VrpBtZZYxJQAD
PpFJg4gYpVdBQthjYwGy0fQLxx02yrLKKU57kijm5qANDNcI+V8j2puLjba0ADaUHZXTvfIpsG2d
G+RYtcr6oUUZAdLjfyP7RSG0lFoXqj5HzwlTjEDfTXMN2UXkGxiS7BGyiJoLE8QY0ZNr9FjoKXGM
gYutvjTEj/Ty77fyZ1S/qD6CBPguqSUbeZ5QknZEnR3FEuORkNT8fh5P/HS83c+axGDnhi2+8E6/
JIDgYWyYCBYOOOCmLZZS8K3xWhJvH3xhepvaDi83RRyd37FQO4cTivGvbPn/iBbHoUcEgjXvjBBY
TQXXoUBBDBzsESztHxYGKpNhN6FwfXQOHIkzIuN1jCFMqmdDXz+epCHY3h3f2uySlRRANr8fRvap
mv3meXSmfrpkuORxvV7Ulhrt4UPh0U+2NoRV5VyOIKcKK/6ViMAY3KRRYGov6WG+1vwd7XyaQlN2
W4slLCQM4iekF8zUcuY+2knjANWWv+V0p3dKHGKHlCGqgWMZZBC7SVH3raWmgY9WtlDic4Ewxcd8
HI+BKGX7ftEaPMLECvJbLAZSPg58o7CB8GDyHKdnitY/tx/NFxTG1eV38XO9oVy0AaHmqMSjq7u9
Gs9u3/80DDYAQJit9DAYQusPuW5nQLcFxRtDnC461sRqXcv0Bdm3L6YDAYgDqRI46FUFR0Jr7neC
Gyskm4keSx34A+EXp3BKbQh/tSNltb7g1UAtIWiRD71nEBC0rHHe778cA5bNFmhVjuLAi7ahmRi2
o6mM7wVITWvSYCOOLs3Gd2clOW//TjTTGJr6a+3EafPt8fohHToVhiTbnN0oyYN4eFeup90Zi0wP
E4f+VdTip7eHf8gSsMX3OVba7QySHK205WxIY32lrNBd2eUEGujDu/0OdAcMZGOFZgNjHz9lqMga
LLltbpME0JPP1O+5UmIlnk48esnk3AUuqaV6OYOfCFDjcuNqjlJDkyUDoNSBe9CFOSVSKlo1CCsS
PtlIurb8FTIrJGXCoABrtY9lDFgBHE3INsktisAKqh5TYysNadqn/RWc9s0sjnkj3PYLxVNDmG3L
tKLQr1BL0h4vfTWgxk+Vf7YxEbpp33m7UW+d99RZSBp44CLByzhCExW7CY8OI/mLUsMPWV678nmP
7UuqJEQP3hF2hNMDyUmhOA6/WG8h+55zbcR6nVSbh+Ah2C6lX88s9s1Ydbkth0dISdfUAGNB4SLe
8BwYF0hvBf+mdoYsBbSpPm3b9iz59Xbmlq3TzdP/A3ycHs02mmVa9k6uEyVc5y9rKoxT2QiqB3VP
veJFmfNWefAbXb1cXZNmbMnGCf2Z/epNGCztPMKwzUJ0SeGdUHscksEhReUusxNCj2EgHwWiYK3K
5iCXCQat4h7ZiViF0Utk7dazMyWGG1L4ggd+gsPCo1Owmn/E2Cu6WJmMIIRO2J1eAaXx/h33x+V+
Rov6tmJC2EzmVFgLo8k3AL8ZaWexklWzD6znWfkwW9LJhMmFN6CRIK+VPSGB5SiECXdFHAAJSwqr
BLd+OlJb5PxfRzDg3OgwibQAmOZXcZh24xS5NvjntV69fFYNjjeQEde7j0FcLZ9ZRWEUvkiJhOvL
C5AFFoLHYdPe4zZlSVO+USra03tMEOF5ijPrTOogbUDPfYZU88ieUUtbhlZgXOrRyg1kylDwr3aT
KU702JPJhbo3thDOWc59U5whH1Msozl9gNHFfso/XLeeTggMeOmjZAh2AwGg78mbDcbG2vYwrA3a
PezRYSPY1KqJUg4BUmbGuiHvCElPiEt8OhsCahhZ01nFSxxgw2SZWrerVh8roJChNKzOq07tlTFl
2GrW3KG5tc7ckP/Hc7SxPgYnJssTuS5N2coIcMh8QZtWy/mI/VwkxMNhyl7cK4+LfoLq6LqQ2mg4
6HRBCjgbsJC25BJWNtYLll9XOy1qfSpQoLn1wz1MmPxq6r+6A/cW8wEAm1/nNNCda9/6k7zqRLuK
pqu2qddHuTHIc2r19gkRO7NfGrJMLAZb0GKDV2HuDZ7q472qT1ZYD5irfXEwzmYEmtIC1ta1TsVa
8a6HdsNlKU5rlhl3qDb0wBwWTNwogtEVtDr5g57QKQaGnCpM0csnaX3wPdqNyIJtukNC03tUwpXF
I79QFv7faI6+8okjYqwnpDmRjE4f2tm+CHbDbIJpFVbexGrRV0Fno5PSzUb49EXZVun9vgIdMWXR
obb1ccZWlmSyc3WALn3/cLbRZ2QSulEHprbj230lc+RxgMnt0blH/05rZ7c41PFH8Uk31WfpVi2n
eKGLPeOT9hioZXd0DZTLt8QC2S/jVzde+FfPV4WrAexfUe+qeh8Ilr8ILJF8B2qaKG4hGd7gyxoC
mPIfHK9fcXoMIVMo6yiZAdzVMgJrIDtxcJlFqoJpayQHPqhS4N3w8Fih04X52Z1k2DPqG+sOMgIW
/z8LrixgpL3QMpeOCPFUGckk48neINZ94897i1MW08CwxddNFNAnz/QXHtkTqG9Z9GADN+efmP9A
GpRZt2DXwpTAYnsnGRFSFMuYyTLxXSYCHuo14YgMivwfOn7jx+SGr/e0FPbFh4nR+gihkwon0i1l
Je6es9pHoZ4QFYuqqJSRbnA+zKU3T52T5bB0DxLzs+wJhdfTxZDmZtXQk/d/YeA3mUErunQOWmjp
pjqLukPmjvnpxwI+dQflN6cZe+746iBlXMvuEunEq3h4hkNmB2XvQ528cUDV52jymcw70UynMrd7
RzjgI7naVuWNGloUFYOxG0KjF6sm6H1QErmZahtLGbpYSZUuNHjyWEwPi+AQXBWddEcT2a/igC3T
83cJKaBap+n02a/xGB0KgLWWpXEWvXdUMAIPN1chUnR1rO0hmpbZKP9f1ZnkSfQ2cco9gjV2UowR
BPZHLRLyN3EoNe92LGHdqO8eBd3At8puzbXE1Mn8jLt2b4HEqBuFJ51fbLd1L2O1nRDomvxAEVxi
WMDSIJbTa/vR/qRQcz/YWJfeZkOusGS/dAIEcZQb3mrnqkPkU1alAFQYfDZHqcyb2eeFZ+rWuYbj
Z1doslzJ4z0jPHlZdt7N3Y/VN7mgTZYPs0Uf4YnHLSYldeWnBjtG6963Xzbv60bCYwJZghM35QVA
I+5RqRDYlC9HdKY2uOf3UKbvk7yhMnpGbQkmM+BKC2/dsP3jLbBLNVwZ/mVGpWEntvd/0kfxuju/
o9nih2tYQvS0tBpVj94AOSrZDha7/mY6c9oiEhhX9038ZURU93DaHjoFQzmbw49y1FmWnkTNPoBd
dMOgz81eMDSdxGd1M39ImS5cndEBqe0PLy4WumoSHR/WsKDN6fCa/VfhRgflJMTG8TzunawYwnkX
fz49OSLcmTOcqGlEOc8/zXg9RL33WxtnvRT1xNZHZA4JmKZQ3p3+7GhlQh5qfGRhk9npoAgCjHbz
Bf02Imvy6vQ8iYlL7K9/6pE6eSmGotDS2+HujHEdAp2eDTF1+EZCqjASHKUyN16i96c9qrkEdBFu
JjGjM5yzWrtkbSE6lL+plSA5HcQI7K+PENcIK/sjt3Jpy4nnd96d+gRk+Bb1hpD2YAlYQ4uafOjT
uXfV2JIpNi3gmIqaXTEmKVxqdA6DYC/On7RC7dSXuRMxbFLLVLDu06ZArPWqlWFCZgEweCk9qdYz
MmbjZFmuCC1GxnQ7ytk5bqL1trTPdEz3i3FlGuz/PwW3QMfGd3dLN5trET0DIg8sLk5WHGrRNdQJ
CiGwNNkMBsKkKprWhmV97tHfcxmZW+nPfEzWDYeN/NfuVL2nSMzvLAi9mC+/2H+DERzEgZ4tgBE3
5oogApzO6NI5zTpbLzrKChPuvfAwsbwy07YMWQ/oQHq4eNmotvzJG3Erb1mQLcTOt6UiClEejYsA
YfhS2yv1Sh7jxRwnnQ2HctcRczecoMIqFwPR2+H2tPoujovpIiido99Ac+3FMxuXo87YwCb3/NwE
yjSuy/c2i6IY7bp3z0O7i9OhM00lUAEDNWrlmXHBCsFvgcLwe6sKbWrKQLaeSHpcgIg+L2QlZoGi
0KeIhxcrEeLyRlr7ftmdAEtYKm9AM9rqr9OixaeJO8X2jLP8osEDEezsz0iUiBd33WpEtDGe+nNx
fR6iyLqt/ifJCtKxiifkK4APtjY7+riDMx/PBOLdR4pllid2KKOMzJ9Q/CwTnzqYSnia2reN4sTj
KsO6sUj6xTRYplEtcvd8Kb7SwW0tESY/9hOiakjO1cV43AJxSiyC5BxFXHpwZdeGvyLr6Wiy2eTw
S8SQT8BbFyzos/aXjn8EMaNfKhflMQQU6Ecg0eUJndzIOeA2x4nB/xRL7Godxwmo56/VRFj+Zpqv
BPiLxsyLiPyJV8PZolHITIAolvs9dZfaFk6/oe4oRBz48bJgtpjJLPK5Xfm4/cKCDuxWZfKhR9l0
1TWrEszxYjfPPHHVK40mOiE4psWPdenTNO8J27qLcbYm1h9rXGaAiAtOCtKD4NqqsBEtmVb3Oloz
IUxDyEOZcFq1dFQoxM5FZFfMynjV68b3ZrfvH/IMbA3/Bqi88m0qduQlRKQT6fovVwFBIAM0EzQu
8g3LuaXVG41skNDWIrcD7mtBtkqxTyqgCiggc5nGuNOt3tG456s4E1H+silf6xc1nirZZsDU/m5y
ZTNCCmsGxEt4BPhThwmuhWYqGWgwdXCZd8k74anACwbb4khbSDIB1QMke3mVdgx549TSwoeQmrI3
fewRIQZQFm9VPGPRl55W13oAWKz6f+SZf5kKvYfcPVnE2le0OAuylCqrW9IitRMG+LtZoqYZhymU
GKFh7lOySCwM/3Ut+DWyw89ylZTMDNtoQae+M47fom9RuI/F9zCCQWuuKbwTSirlxqzZAKl9ZT45
OZeTyhV8i2dwVMvq/0sQY2Zly63wT/jcjR7dxCFZe6Lt/kU0otbd925jv96jtflpD563WQAIjuqx
OtPmkmHoDfrr1isVNaxj1oibcFAHcdnQcw8/F/JJtIPis7zfGU6Wg1oXlRA5b+odYGixRwG2JtBp
tzMwOomzvjCccImqc0I21H0MmCQX9HLodKVWUhN7M0AT7EPTmXkINRAm+w+SGgRcR1EEgNm/H+5r
3stF+oQz/vgyc5QSOCVu6nNYvDfSyY1//8RvkGaxqhAWPJSQ9N9hIPmrkk9Ml8gkQ4iK/IbxnwdN
4lrjOmbadAsl6EvKXC8u/b4duALnHd7ADqq/ZdWPGoMP+SUmOpEJA6HFWyrOZ3l5qjm42CLyZi3Q
2bTM1rJ3yBEn428qPNlMklxDjvgPnQ8Ze9Vx20sXFPYGfewUaDuzscJWhydv81oeDeiaFX+R9hJ8
SVJuzd4fV0RPM+dAh/l7OGIH/WH+cybGyijgo2WQ5AW8Ym0QkmuMS7lEJpL47x2a1ixZT6Wr24s0
l0f80fgT+2a6xDbVnKeVv1Qz2uLwWtJtv/M4gygq1QzGh8FaZiZvOsfTXqnWczxkrui7coTHNw2T
7iRg5Jjmgtxqktkt2BJt9AHG2UVQs7bNxNd9LhCsiB9xnz/HIIsfQA7ooXIcgDTG5dfWqKNyOXnJ
udgMItZ32ymSQhUNZbjm6YG6MkN8t62t3wXHySY8wtdHunB9fsKOOekaH5zRhlok4MT1ZOsSS39a
9JCCtB6F5LW8KT8sjid6fYZzW04jjZmzuu/h42iOu9IN6cup6tkDuGTuvoUwPQIbx7uWhiQBZs5e
LwY3U3bnBdMK3mR2Qqj8PoJyPqN8YPztYn6RvENWX7YjsuGwvyLi2hf88avau5xsb721as/KfHh9
urkY9oYwyYPv5QXicdTIN6pS+/psTlu9oqVUt9CnRITwCXh7JIO9VIVKbMWurgMr4DzhLDGK42nA
FSVd2N+svW6nr5cIgO3sDniTAQg9OhzFYeHGMfogPpoIYjevCufv8/aX/URwyErfJI++w6sg1nGM
hQ4e57LE8ozzIA71WHw03tG8eP9+rD61cjM0qU6HyPuKC9yqcLBZo71UM4bbG29U6XUbByToivJO
R9hEKLTONeu56fluTJhLgdEDe/IXc3OPe8caGCsEfNWJBYY4flO9o98sU8UfhQEdeznN8NGlC3Sy
QhBD+auSXF2slgxkfQCN8Yl73eEzcGJS8LxoHqw3NCffHJfEY6yf8NXN7GttV7PK/nOA5EnUucz2
X9bzb3zU1ksG9OlOS76iBiTX0ZXKOHirLNyVkRcnAkm/Ahs+HKlP4x2cFLIoiWM8QeEcihw5Llpk
FeSB1riu0Xa2ZYL3bSAIGiF8eiAsIUzXX8BZLph639t36TU+y5qg5RFkT18oHr2i2Ov2A/NzEASe
6PGCMUEHzVGcREVdht/Q/BEH5lsQfwFP5vZd0nqna2u52SAdGN4FE7K3Lx5M1YktYTTik+arg0ol
zMwsjNbigAcr9kCYkVHAMe+PeUxyFtaY3vtAVvVXfUlhxHLw1E25NKXsDMYsfGcoQyu1Z9WCZeKN
zFyzTq6zZSHQJzCIYuFavcuNGEaqf1pRUjc90d4Dz8f0etD7cFFIEZcPD84kim4AOf5WYBXKZuG9
x9N7enGSajier6+Qzu4Tdi7nJuGtbUYD0+Q/L+jQb3MICMaBQzP2MKZmYxdQ6CT03a2nZp8oz3FL
i7LqYr9d6ybCtNyeFIAr1rb8b3LTaT5yW1Xt/Emgfsktjxik/Tg7mfogEIjZ/FcfZHTUb87z17N5
L5slTOxucT4Jl5D80OiRugMQNn5BBZLswf5w+I7l/ejqqW81KPr+cqLSYoFbvRmqiL8i5mGmIiFb
bTUe2nelljULKibMEKiCIxqwapzBbvyR6202UiFVR22xzEAawuLj2yN8q1USGxVSUDlM+Q6lnbbs
JkfB0w5ddAkIfHG21TL8saYGNfvsRgv67xVhsMg0XXFLatBVhDdc8FtKwdXWqkR+L2YwG685Alvy
IHaXOgLAwXqUtoEqCTdR7zpA4P1vIj+IxUNU7HXWIJ1iJX9Lqme51n2GyG/g9hdPKjHZVbYs3MR4
hdjE9wqrhVmktwqGl2yaQmfVq9gdxv179tIPWIWdYHL24WkpmTre2RK3WpvlaUP4WZT2tzAloPyg
kaX7WGYtL1YgYMKg4NtQyRxCMYnDDhIrp5qbl1bgFdbZiQ5CCkGCI6c8fSbosI/w0X24T0FfWzz8
g9TSeqVapR1zNOUmx36rdwkRllLO4vEagC2AqQSW7mG2m5Ww8J974JQaJ9N6YL8Rx0EKuONr5mvw
f7+UfLTi5WQBCbs8HPl8BdF+gIViYQ4TwwDiYqHwTuo+hf4bC/lQBiIZWk9RLjj08HQUiYNWOIZP
Rz5ekkN1qZIr9WcJrG2hCingGsMr+uSrxPXfQeearppk5lAPi8QxC0wXxVoZeNRn+VPFF4fBXDqr
ZqmQGSFicSUo67hJ/hBNCoBRNjnKAVqu3lRPLtdtIsWcdbQy13xOrrlgLEqfip6+3YWuZhlJAS6+
4hub1JOJsZNWYO5nUkDWq3wZRuQP2GmuuMFL1Al/psGBbQGgbMP/9y2IfnQm4Nc5ynSHMZMI4ivM
qHbgt16jyzQce9gkKflUvcrrAn9+1X9V4FQlnhGqye+k1MZmDY6IFfKshZhpFa7lXq+dN65Hz5cM
RsMXo/Pky8rygWD9HhsX2wAr8k/5MDktpF5MG2xxRh6XNIDakl3YDQN2p8VreoE6CCWVc0y9XqZc
BnAkD1vxLlqpWttaPEDZwG2zN4m/DKE3UP1J5D8yCPAR0ISu+g1mGK5UyKV0Wpn+MSPw9ocjWUBl
jhwblEyUX3ErCVj8aDelzYv6A44wFPqT5U8bDPEsZd6dJ0frpkceNVnRwuiN79i8cSHjcg4xMaP6
GaEz2PDl1XyWp3/n8x3hluLKCWP1qiQvIJ45ri9T2e3XSqKJZK2NDqTCA2lphnTa7cRnNperUb3N
zPbSoOLJOloqDhyqe1HOLDPrE0oe+gZsEsSM+Tu+BwFwIGIvsztVLxp77iYKoN2bn1RetglZHqgw
B9GIp5aPt0zVy6sZdqScr4p4ARuHN6D9ZAjCaiWCurmXFgh7XpjZLJ5KO9iAIAPTiENI2zw5EieE
+a4HoHyypqJp+9GQq0J8Je0gFI+Rg09ll18Uny8aSMn3fKPYa3vFXW8NrkNA6ZFaiFUneNKQQj7O
mr9mYQ5jPpnxwE33XfBdtguTVwKPJg0PZKMbEEpMlaiJ90w//cVjQXm+vIpjsdHvn/7QkG0efkle
PvaWZZVHPTFqdssD36BjOZymL6FZXRoNWp5Y5QOwQW6lWADp+ZscvnIh63JHrySaCuMhvXHJFLQv
P/LP19vuqmHQ6QkmtpCzg3/dPUY8L64o3HYvzN+zsqQBoMJw6b2Yomms08I64YEubqgdFHb7KhuG
f8pNL2snJF3W44d1m/7wC5XH0d95x5Db6UnXbGHblr/Az0NrCymaTs/dnFXH9NARZ9zoNOVPbfyy
UqgayGRdqtWk/t6HsoQah8vDY7KxdqPHbX/JItgRbIh0t7p/UK3ZBSS66jV33hxs2nJfPIuzlETB
KG1GlwHE8ztWzuhK/J/FTaqn9QiiaNffVvTYWovyvAb7bL5baQNEFQPYKRtzGtpUpCYm79WXD72w
51kBsqwqAiCTlperzTD5G87jmi5KDwslrPBrRC+C8pS5YrKFBQAnh2wPwtkOYH4E3z6Dd7pORcTc
oixfdZ9mEnuelLr884AWrh2HEh/Cjl6eYfYfBB4RS25B4ASmScERs64f965PGNpDgaRURpnm2iBU
PP9xR3lWZwCz6U1PCHVTr+PR8ZShF+W9Kg6a0RsdcUJtkux7lfsiLHmn5zeCVnfi2B7qhAAQ9BFW
gHt6JGTkCuGyVxi6ldIX+t8pVPAs4B5Oy//rvaQMFCteI5T3KXfkeXMjS7h4QY/NeMsFGPK/pUaF
xM6J7CP7LkGW5RLmdN/L0BPRVUzixJ3XE8wRAwJvVVwxuaONM4pZ2NEGqprRYfOqhqZ+4vbOdjCb
lCMMxsDjfOyHShsNrfPZmvxgpJkDLeh++36yAjdG8P51+sNo1vWuxyoIov2uC74XNhpQAgn+NAMY
gMxICJpyU/wErXixGhtSTg/lW3kRiGlDVa0An7yVZUBjIKERm5e0VOP5LepxEMcD+kuVNu8ue//R
h3D4FQj7jgu3pbcfx7pZlFPOWFhSxa8335wq+Im0o0mlcgdrdmGyszARDb66eFz9BxlKiSoEe7II
fv1I6RzyqCcfWeCwvvy3I49d0j3GXlND9Q1EviVNLAQN0ot7K2HsgR+B5WS6wW4iLXKzp/KZ3Y25
ie620EuPvWtOiw1kYaBNE4orLRjISnS9udbKF1mztuOy1tagAszQQJ2mUUPrUsBDbwB1R6wJdzQz
gKTYEjRpqNRAMJaWeiE22FtuokHH53zH3aY09MHIU/DaucAxrFpgmegtO98/9IiQwPh5HPvMPU7a
kMU43vrt+B8fsINk2HD/vKRF7Jx3+5dEpellKJvqknfnKBT8Ixh1M89rISxMpn5BWVrhJ1sovVnN
jF/crPK/OVko9HY8OfXHN/V4qubWJUMwSDVC54AKKfYHbZo6P9OEZ46EqNVSYErOu5aVrML/xVGo
qp92vpGLmmQv4nZiiyaZqNW/07xVfoVlyBSj2s38niAe5MYvc2XghcNaUFG3uO2nJ+5TVAkYCQ2R
mfX661unibArmFYKAWtIKDRE/38u3uSagfD1jsoFXH01HHK2hhuMdwTsvObS7N6/om5EkJ0vZXnz
6ek5lmy2KSYx1DLnppoE4UQazjcc+rK7DCyCRKMVldbOed6G12ElhB6PO5XhHQSoGzumzps7AnAy
lvyiYWEgM21rz/IeDJGhPPT/S3sWEvZWaCdSSOHjqL4Srg/zZMMtAa8vJDqhssPOcjphlGOepfh7
ju3yTLTVjYtAMyF6z/6Kr2np7EECUOxwWyfAz4vbNTXEpJecajXtPUVQpinvZJwjp5ffAHG71n8B
A1j5fBhejM9B7rYHi5rma1AF3oZQhx+OZ0/pLqOA0vPE1zm/ePJesloSPTIrO/4km/UpcsP9uarM
jv/ceSrX5wHgyNfIoGNMS7Yks3S79Gv3wAUMlW9hyCuIF31CYcF3rryHm8/Nx32h7MdISGyUwVpz
0U6y30DygHotr3CUxsuWwSoNeU/uw6xGvbG+uvM7E4O1sNAj0cbQJZGUSxZzrDRuxZnRWBEFBeKF
94s+MyJjwTTWsvFOUbUBQmt4foI5jKgmkMGgf8QY94jjVmrwkDX6xB2SgOKHj1gUUwE3IkCmnCuw
TofIrhxQ+UCJpNHDcgemTbPLcSkV3pXktnOI0vBY7yDXq6vCAXmeVZRIu9edqCnvGx1rPodAiRe/
rpxlpGpNGwuUpLE50Vw7x6s1UhqYD1RUE2s9VlSvPpaAMvv4Knj+YMCvg1fJE0FNaCrAjWQ6iOlv
kMkHH4W7ev9KNkonCk6l+RccXK3fSwrxwAvvLjG/y1oerv3PKbp+FtLfRgiQPvoX/VvZjzkylioh
vO9TwRy8dFJRckkNbm3BRMZmLnu+cmVsfxfgV4UaJZkLo+lSpYzbJwLDPEvegsbEciqImuGcv3Hk
Bq3rMB/57gn54AYKTWFK3yS+Jq2MoM0dm8hbkDCsJzMGcnRWJzy7xdgtA0UhCeDDt6PQQxyie5I0
8H0kOfHS/RaSBUU+PUMqq6rmugUdq4UAAbDiyzN7jsTrtOnzIYsmyY++5H7Elw6pv5k2P9E0SUu9
oko0qWhF+TgHeFsPhr/0LO1wZYS2Gh8Nl2ZgsnxZxh1mIFi4H7d3xX4fMayx6zy7kb59GbAph6HN
SEBdbUGoCvLZ+Zo8TUpsCXwkB4J2fQa8S/2/kASxmOM86ug388cyrC1q06MdnBRJ7hP/K4Kkt1wy
TALPXfjMPocHgox1ecDvR/lOS9SouH+bFdSHK7+TBk7Pxnn7J+AGw0m2hqpqLIMftyDOPjpcGGg6
+V5oRqCrpOMvHH6ZTy67jr5irUVf9cRLh4fv6/12tIJTey7kFTKT6z5pq4g5heoySFJMcsUjm3zG
zgfqjlrH6Ghybd/4W4yuJdLw9iM6ql9Z220IE8zASBgJ3/osfyKlcjEUpHlj9rSn9F4gXMvYBf3T
DE/fZKiuZtq0JrvBDOPr3VGPpkhgoazx/jJEahbOTo0poBx9wPj2Cfg4oPOi9CdOb7XlSe/YdJyf
B6cuzCUBACs6V8ivKY2izaa2YZ+k6H/TDp2NliKbheK/Rd7WbRt/woZWkUKpJyPInt4h0Ew7gyN9
ZV9Vz9/b5dMfJzlsfHFP0FxMKMIj/UrmsMDc7Nl/mSp849DQ+WSkgZA6gow25izxbkQCdhyJHkJG
fy+pO1f5QgTPLzd9Fu29MI5AdsTHqV0zWmOneTp8llJX34qe4aO1OhVfejcR9Anc25z1XWq40cY7
5aS2uAVPLwehzuteNVhxw3GmKMUzfDqUvzZCV4hlHX2R1hqof9cu1yrf1sQR66M8hSu+lTYWp/2C
PEecWbDlmlWsFV+mnSiLKo+JDJTSPFolF2wGepii/yo/AstvYum18c/yGb6F1TFO9XRCuiCY34mO
HHD0PEM/a6Q6A1T5YiQ89dyZs0OGcQQ5taMSj9y8Z2xVoSNK+Wmy+LxKFGFJ5oyVuoxDi/LfNwrZ
L11NnFhcbKpVvt85IybC4pvXSbfm9BxLScDQd5tc8fFUseae8MwfFpIBgxA//PC/qX/4v0mGXe7j
OCvLr6ykZd9RuBqQGumjvfdr2B7Au/mWCn0DdNKm+cUhCIWLVujmmIApieYJK5v/R7rpgaLXdbEC
clPdbaFb0+CSPyvsmYzFVYmAGODuTIZM0VQUXY+J7gjToxZv+/ChqgzBtKi7OxVtZK76GNLeyOoc
OmqspseyPt1R7YTaJNMu301AFtBJVZxL011mYd4xFaNTeRrjL40goh+/6ptrSyWPHxAZApJu31L+
77AvavWJiXBIgTc/D/plM/o/G2OsuF5oHn1t5Bg3n7TbiZLLMHU6hcgk2mM8LQv2hxqxuOLA291w
R0rscIy/911bXmKxwwYkDsK52B8x4MLMb62cSm6SX5kF1Zhi/0mUXBvE9h98iCrrQX4XZhfPLwzo
qRzj/zGLa8jfZjACaNLtu7Yj7zVRGRSMdtrfyFFjo43M53WtQomS9LDxmn0fgWq9l890eB8dDFcF
Bq/C9lXGLAv26DVqSesa0eLBQVjUmc6/GCOLdbhJI3XN1r9xaBMfMDBCOWFH0B6kKEG41T/c4bOU
MgWYi3QlZFZ4CEHcnfxy5tjmcQ3EcL9S+l1GxSbtQxDmdWoDRksKTN7zmrHDzxyogxFU/ANSyAyK
/5xb2Spg8W3ujxjvluX7VYIGSjYY8oRyZwf9vbLB/M99NWcSztRqu2os+Av05yKbdetjyUEBfyFW
iIOYmjyiu+Ag2i4moXrjnTZ06DWOaXnWonjW7cxuxg9rwOwTEi6tJiJ+v1YqBUUG5HSLd1cr7ROV
IXOs0QwuqsnpdQ3CTy0AZO3IFrl68CQOuwB8yfSALxfpefab69mLZ4aKYjdx2G6DZSlFlNz36YIG
eKFvWhQTqpcrmsYBqMYPaPDMWjF5sP/uNMRtD4V2Lek8Aa+8zhC4zmbGbKpAtz0Vgja1ekuAi94G
bagpkLHgANWQCK8cZQk/3pwnDxu9FBgYDSFzmNTsmzls/xJ3cR+RvARnM3UNQPsObaFZbxKiihlr
Y0hWIJYKYm7mfhe9TQsKM1ysvDcIUxdydUsq76j28CM14bUI+u57Ep9JC3Ef2AoiwTbaJpd3bqf0
ueiuImNelLO3v95ETIv2Bq0R7mbMYD49djDvWt8A5PsSrSxHOvtP9YPM13uGlYlrTvxwJ6NhojnL
dplYYC4j0FYL6BeQtgzJBs6O1kJMnl00krhqa6O7EmphKRqs/j4m96noqCXxv/mCQylN0HbKNARc
0JxUsPsE8h6AKfXR78CuObvDV0w505MHhKfQN/bgSY/7yF8EpbGyXs3ICdgBTeGBxLVrv+ZNTzRB
dhY8wzWMrn+8ymrjnCqmaOxrUu8GWRKzbl+RPMQbpZhKwJPThK+KmxVyx3ZbbnY8SuPtu1iTxWFo
f40tMwL4kCFvgjRz3RDtbSd4SMGGXeOWr+OChFJntiP/+80flbrIIz/Ku8zooRv+WOl9/WbU2FO7
ExBklKAnohWgmN7gL0U9b8DdG8SbmDELyULMqWrn/YKxvNiH/wQpqaMpmOMwfbgOhJVMRSzmf/TL
UpFK12qjURtjxU7TuVh7iCw3aRBkQO6MbIBNFJ9b3xtDWgkyhBNB3afQh1a0O773BxhyQjXZp1hE
y+6L1cle6O9yD9pYpRq5A6vzLafPDT02Yn0R5PQWDqxuCnGfF6MPZLBqTb2SBGUb/flQmvxz+b97
NV9Q333UPT0IoYgbcklHzyvSj54qa8zBqdH4Jp5HXubBeKQuDm4uIkfz8wTfqesvJH+GH5nWMegZ
TWuX8i7LMjCwh3jrIbnTg31PBKyQO7chupzT4OQZMbWditW/c1Po55zCH7Jg7angUCfCN6+iDBcX
EXas6x1Gbb4VUlDrHkmixDdbAfvPueZWBmE8LHt227XGK5Pv3SyREW26nRs88M1vebiizDzb5fx/
656jMx5DlAHTxRqA6L7XpL0rNarGmvEX0FLAkEt80cOUeR5fw3v1Iwfeq+rXYqb7BsSbJ1/bw5Ba
zwhM4atNbuskNoK8pkAEWjAhS+o5IeShAdoApphjuZMumo1NC4Kz5Cpjm3mrT7gT/pwYhjsi76IK
Kuma2U6dfrIh1acQqZ4u+tL5jVStlu6IDKQiC95ZPSeJOqw4Jv1KBGhdQ8YhbFYoaNjg9IRU6TWb
MpRYBWMCnv1lU4W/H6W0Hqg6pRt/i0N+he0ZXD4ph33w5sBBccGFozZqF2XZiNtyhQDBygVDcK27
usPcJy9RJWyUbAZcLxBZQNw4N7AAxqPPs6e2rL1xQwqufKB+oCi6d1ahk0tuRSYjOviX2jMYBnve
C87h4s4pOl4wF+Hvky3lvIaHjxPybQpV3P3EaY2Cumdw8+I2xVU32/TEz3TkYqdc1lu1ikDUePYL
+Ok5m/tiAdS1dZfiMYhay0pJHrQRstVDnTxC1XtrjaHZzR7qiFlDmCauUOQmkHpT7UAyDT+h75Zg
c6vS36h2XaenYdYSEttgdp+AVrnINDBlMLCQ0Bj3hJ7x0VqqxZqjpkG9Kz7osce+LKRTKBx7ax1G
CC3tuxtI30UqQr9iVZidlrTsa9r8bcriDTvQu9wQyDwzcbP9+DU9nShUAKC1zu6kiCk71CFpVuI6
OvtVqs3M9Nhy7h5ReYkgKq0dy1pYpwtpz7w9e5jQ9VE3NDYut9gFhjBxjuFliegAhquyFw0k+BfP
VOfwrzddHOeHaroCfuKMEKGEo/pzlQAxtALhNfdSSc+87jR+I0ofW9B8NYWnKwjexNoRnaNlPC4G
fCJg2X1lhFxVWNJtyFovfrNy7s9BGLTnAOeWZEF9fliqxeZhH5qDnRwlGnVMZetOoMQF1FqT1hFn
X7B3gUSOQGwK2YM/qHybDeB9bWYErPOE36J6n1mg9wFZHXWVBIsDtfbhMFGcSt8holx3bjhvTyP2
dRmYQOLnezF+/c2D1weXrBwNksXy+9b6c0mPvFMCDEIDIjZw3kTlpNsmr3uaXwh3tvJ4zwpjmZu3
Qu4F7HEZHKUU6+AvS13xg3uuh/UuIUYRzAjjWgNZhJeJQ5Q7sP4mCBlwKHUSnx8zMB3tNcdOLHOx
K+8DXsTtBj+FNwhVynEuZwgyXhJEtpNTxcnu4JM8MRYxdVK3w1oOGJMYG/sUEA2//v4M799zd86l
aV7wtNnlVbD+d1ydZzqR3ygYpBhGalXb/VwyaQL65CpZCWX4Ud4J2qh3CPUX4Lh63zmTnby4sr+C
Df/1P1MvcTtMLyET0L0Jt2fcoXGt9mVYwiezoYvBBqrCKbo5NiJ6u02/pBpa46bNATVIsB7nkWpB
132Bvyl4lVIROEfCwTyEhC7y3M5NcLuEJnORH+5TwRv4iHA8EPYCCNGq5acK2Ltl0IU/PDITtvKT
8iiirGXKq3vX4GnyHX2hkhChovOfYYC35SBAvrEqOXRIIbIxrg497gBtft7yU/5VG5TGNnLTDDXq
/O9LmKXBQQoDv6J9SwkwM8124h5VVQRCrIAn3zCjjSepicERn6tdx1Z8dXIKABr1S2+7wWenEjJw
QkHzuYdRkzoTApUjw6ZO6SR5FTerel7cQZkJp0VD0oU2G5L0iz/9qkEk5JiQpkbnTqcv6a42H3kK
+t61ZCbS/FzVT/lbpyf6YcftfcpjQy4PUAlArOPRASHo5Wrsv7DVQD/d6IZ1JMJpzSKCcaNZ2JRq
i0SOXi5oagy7hLjtrLyWHreb0jDI0BcbxbPO+de3P8KrdhdG2Ch+k7Edlz0LuRB/de7fDQqsd6fu
UIEXsXps9EP2+9ex68YYqALDaU7utE1OCQgCe5F8WMEOl8YCV3m12dzWXyStYEldhD2zjt1Ez3Hw
836hhh1r+b9iJfIeJKpfCU2H+LGx8YkqXY5QaGZ/HBc0hwxL6U/6k14LTtlIwV7Oikp+6O40OHcC
IZefCcp0vQWZNjsFnFfYpBG5joqun372LxP041uIufmimZGLTCh6b71BVgoXPZ3MydiYkp44cwVF
zeXtjtSUo8qTAqC0Obg4LbYoPqtUXunQdaR6J6is5N2ghpVXMYq085wZht5pDEoJftyvzxCZS2BC
ChJ1rkP5ZrPRR0d5aG6JNWccjUy3XEMESMur+/Ja0duq/eyi5snC1xNcl7ui9BaOId6nXRMEfE2r
xMUJ7Ww2HD7zHhV13M50x0AiZ8iVtEerpwcwL0EmYFyEH1NVainU9V+0HzatS1wlf3zu3sDgRprO
zSnTmAsLhiMRpzR8+FLNCvGqwkW0ZYRc/KSCNsLJvubIdwNlJY/jtFbpF/vO2gVtvG4umElgC5lP
xdVvNLs9HwsZAPf3AZ0TqDMzMKtYiaPhIIWAB4m7Gnt24jyovwbzz/B1bEaqXSfZfBhYFEqOKdIG
Dvi4bbT94Gi0FleKi+he976SL++MFXx1hxh35bKlTYAmgLTYOd6LccleAcwVJ7RwXZDBOljHYwaF
ORelmKK5/qW/Qdne6fT+nHc+vsGfi+FG/J+Cw2ks9AvZrLJDM9XpE/PSXz549KuwCZBFQJqBU/n9
27GtvY8+sDdk9SEEDqgt9HrtchTAI33bJvuC1vkQExDM5ju6zQ9G18A8/BgArP3lr8DXrme+u4Ll
56lYSdZRBoIjAIQlrmZ7YPT0m4O2v/9zAkNMkxAtXZ5mPjdJeJZKU+DcfFC9PPVnw4p5rQRo0O/9
z1bn+5VVFLEwll0ABMLgkZr0WrDr0qffFfdd1Mh/hsBop7KjWEzB2pZimuVPBhQCJIVK8ApG5Aqg
/3EPXPfGGm8bvVCqx+GO6jErvSWfZ0xPMoJQiPK/0OvhY99VRUxSFiGrKZir7URuOEaH4rAyRbvD
o0IlY2gQ2qxRJ4LoQM+mOuwKl27GQcREctstwOJWXO+VbzvXv/Op1Ns4VLCMidEbPCmX0aQURloV
29f/4ruAFj0olOI3N+3WGysoeVH5SnZpfH/YIOvVWcVtdg7hUriFOCT5YsZextuEEBVfBi4fmL0F
xPQ+VRcJO8SamaxHe44HAPTAfUg1MhxrAgxYEyVTq0VtnPsuu9/WpQAn5GPqOOhEYA128nVRS//x
hI7NAnD0qnWaud9CkqNn4/h/Sas7vHUfHbNR44umkAEl5NaQ3FZMDe7OJq5ArDAyZAa/adp+z8TI
F8kbkfvT2LXl1TRAmLMN3MbGNmNqEcodxpzdmAx3SHC/4JuBUVKR64XP0OD7K2XuWzi/4TcVicvE
myFsyQUEWxOzvoB60GSigQfLLTyKC3v6sR62BJ8lOjfyG0qXDUcFZoY5gfijyvLLr/r5BRSXwVM9
qg686L3Z928YCQZq3L48vu5WVSr9euHXuudw7fX4XcZ93PZDb+TYL6x6/3QBuv8jTvNH3/TGRFz9
lUAk04xlqJha+eAgb/eWTrrJ6AortQ3BlY7VYmwSfS7b0PGkFblzazNWhZP6dt9lQuIMycjl993I
GH66cs5A3nTroV82t2FfqfbI9EndMAoBEY8KquzugMHBlFd28hXu3ZAq6huYDSEfyTbU14Q1xsBn
6f+Uw4luY7EBj1KbQ/dlBzHvpMV7z9qm3NlKIysAGmMZiRN7DW4FuKvdXE0lYMs8fJmedZAPwXw6
U1okALoZOgIJUBmP0yTaf5G0QYvDBQlniTkaxukCNIkXcF6oygiBaT60CqG2yqrJRcK1oXC37c2t
cG9OfuYz9NfiRR1IxwHES89r4iVbQbekaTSSxxmrqBG8fTf49jxLyqa85l/Zcq9VAxLv3Zf0065L
tg6M3NdqnKPofDMfv1QelY9ml8+Qowdwzw5iOG2sc2cKaBhpb68LZB0UjkVK8KqMnljQedr7O0zm
DPgMPQ2u9vuOGkY0g3b7QT9qldROTMBlrY8ZBm5vnsoZ7EJgLUGCL9JE9a5mOEtkvxxbnxjsZjXg
9LjfIZI7ILhEN0UOwWh5aLkxxLBr1e5gfHvjaKIqyrIPA++26ix36a7RdUDLNaZTu/z9N/8jBr54
01tOqc9HlsM+/aVdlf7TYihpZK7eQr5JhPi5WUhn8xmefsJOac2mW/tPc3cufePNbvMIE6mPzHpZ
EaOTBmIcyMsmJwp69nO6Vg5w+PchcuXkDsh1JQTAznCC87ovfQnMNNvojBO2mOBypi2eR84ZiFA3
9qFJdEPxb4lSeUJ6HBzmyhK2ohuP5rg+Db1POzXoFGAV1lstZypOA4v9CJ20vkvUdc4XpoyOYwFd
d3qi/p7XB0GXE97BcQrIMGXCP4otrnkFtBiSLfwErlsbA8Cy6RpmMgBGwIyn0YdJuszdtMBU9JgZ
hUYH/Hh8EAbNTHIjz4tNAV9HnIeIgXY2PDExV/rZqVbc2RWBwEl8b4cJL6Vn0ydySh2+7H0IuLgt
F45O8/hmLcZUDLrXboKoHRCQE+w9SNCyxutkUB/VMPM+fPI0JbkY4t3/f/id9cssZEyxK9YPx1Ib
xtz7roCsWkP+Z8/m9hExJZ1LoQUHV1kp13ofmB2ZV18t2M2So8GvU5/vSbLNubgd4OXCVdRdhquP
949HN3XBIAAEXcT0FD5r8N7cZMaxMwFdSNAnTwjdyXagHrCAV4fHPRHaX7ElkY99TWtzZpeviMX9
IFT8YpfIsnX2VzYfBm3G9/m1qfpt6aShqksRIHuPtJArZkvdS4SYl3hr81JbBXVtQ+eREKLUHWsU
uDmavIy8GZMXXZm0GFPpHbpym9B+VuHBg6lc0JDvdtJh+KC5RBGBtXQ/UE98xMPMEr3ylM+gzRM7
8VIKXTQjuqb9T57y7wYTCktsCMMDJDnnqrrYAo/9T6GGdykUgdNZJRUj7dKo3JiAzUof4nYZYxA+
+x7ZQL52Nr39Q/aSsv/tAgmzINJbWCCWL6yWDaKOVX/GRya81uFCn26oCBtecGjZyY+PPiopE46l
aTLrMb/m3vOycYuuBRdtX3+nPswbL7IMMFMaGpO87nNTSFLejll0sjkDNm0+WXgPdpy1oBoTqKbJ
IKcOdh1mAjiAZ9nwVCFO10tq9moOIiuqNAKa7yb5FGWz0ePvwPmoL3w8KKYTFuk9bVspDfjeAsz/
CLUgmbjlkTfnUbPJQNNsGZuUdeDOxOj1wyTYh3MZGklUiUKS3CQlZwifLPpPraHG7EfUzD0ekFMH
9YGg/WGIlL1t+urFCpf430pSxru2usUOZbHS6EG61KUUlJ51q1joWfhLSocyr7OcCPOPbDPzyEKP
/x6CrwfsXjhR46BBlqZ1lTp8hQWSBCWlkkW/lMTr6Kz6+D8e8n3AI/uULHDGNgw0lqIc1q3t50AC
kvUhf96+n3NjT4qiCsUwpL9xmlg1Oe/eJmfuRJpmEEmc7YbbOh3HKXcjpK2Y9IdEkC7rI3jYuE2+
09PDpl3BYHlAqwUeSxAcrKrUPvquIPfPXfkzqyEYK070T7n0/ZyZbokQ0aRSWlxTTza+FEFs8nNP
e0DyCUgJzLo6pYd4JZqTG9UIbYgeGw41jTWwikn4RfCaExUsWGo9YWMj3IEAww8tuRQ2GDTA5TOY
4vUkI7lF4tHH2GB1fh+yI8zkTHqTLhgmN35AKJw4zmjVm1X2zWycnojyNWg+HERYI54LRZ4XAvEE
1yfH9gcjD5JeIJllByu6Cc9muLopdh+BE++5Jw7qaz2M52GUu5Pk2S1WSWN9nXnh5C5rJMbJZZds
M280u8259XXCEAoPCzB4e4u8+o0PNP1zhpcT2K3nEyhkkaClTAfjQxFVaXvY5/ejawQyWYSWPUWp
THyP2U+rbAQrehM+3pCORYaJkVeTeFuL7Vck3UF5pLN4rsRGrTtGSz13lqZJZKAY3cetZg6p27u2
fs7hGF4C7jqNRprjj4VlW1pqNTdyagBbMJWNoiNqlYWOpE8MsmDQXbd1OjiTNvd55jJFvqPlnz9A
5FgUb/I98fJtw2IkGDC893gxvoKhPKp2lMTFs79tAyIbpnOMQfrUZpv9JRj/ENDuud5ASffaldDB
mLa9ZM/AsWuUiQx0bjQ2vwbGDBrgb1P9QMtTuDxorVw74rB9FXhzxGt4ejlI60ncD4FWjSMgqFD2
u7p5biaeCRFq9kC505j7S4KGeaiBF2Vw6q7IqQYVPJmjGmKS6m9jrMZY7xUyJWiVhrxJc/3XIUzS
wYAW1Eshro3CHr+0ZBrxBSdr+h88m37HnxtpWV/eB9AWCQ7yBGSyEIqe17M0vCBO8l+9vkKsFROq
fjTAZzbkM77Y5CyLBraCfWAdUD3jy4bLbLFHHA/EMOcfQQ8v6rlEeCl7jvX9175Rq5m+9j/1k7/V
rNr2JvVLAaNhG2bBFL/KSzgonRezABaYcDXvXncKXSQUddU+o4kDdFwkVLFV+KJ/ZvSLixH4QsR7
O42trA9tiqRuFj2D09n/GgRTqAh+ZRbhMNbc1Eu1B8/s+ep1eg8CuYh1kIVjM/yShFFcRU0nDPXj
JkLAHam8ne+nYi/fDD4aIjZrfe+/VSq6+lxyPe4dfYPyKbN8896DxeoW0t6iYCC/x97aP6vys5+0
4F6EFMkr8bfLo9EA4NFc32ZvqGTQxOMfCmwbgCtwOqHvw+9Zq9fcTjbIen8j46vJrFQCFnK/rwec
aS6ORz/ElVDW3WRnHDF1laVTq9JKIKoBrlLfnFSjPUV2K+b2qQ6pzRY/3C2Wf6k3U4j8PuzcNel9
wcMHbN7wiBOa/vivLJKLKjY0+9RWIPumk/AqMHzrErRz3qESQb/csKxWIeYAAyCMoqsWrK+C7BJy
DxYXG0dSeIIvZHPeJQqMWMLF4xBo9h4wUWt8VYnPX1CdUkWONeAj+vtkyB/ENWZHcnu5RSoEiWVG
ejNNH5saGfT8n1H0JMYmAed8jhFZ6crvQLgeiRhIDaRFTc3nx09EoqqZ5DxPP80FDQ8958wbPusw
OHZT2Wbfd/TDGvfH+yNVuZMqu+wB7apsFQSGwrTVMubzdNH13cSdK+sjxtBuOe8xLmpkLOF4Pzq7
pq/UJOIS3q5xMTTlvaPtXX5ULaUxzxjD9vNIOtisdJKwFZd8HOt5oxAYFDIQdNgB1ki6cvLDG3vA
XRrJM3tX+qhubyc220YqqzFYtpMXLxx1yssUuLMYtQzZTjT3Gt2IKTSJovAkmI6P1oLiGHMtVY3Z
uoaB+gtdqcC7Pj0bHpmDsnM6nIjND5tG08JfH+dPcqqW0B+QA1smz2xbU7hMXOmkkwE9VqkKNChQ
VCtUZe3H1bAfhMda9uzuu8lXmJjJv7QSJ3R7myVpdiTIBszyOSC0Fn4sFDgR1mTQ1XghLh1/XZj+
o1pnPDgoRs0PtVm/nyt4llqSeo1bJszHepYTXqqBYwBwEHjJVKM1YwOZX/Ym9TwzbPSBOwuJ0u5F
deTDVeJQ8WiF/vu1PSzUWSbEIomH90HmnpqItre34IysWFMiDpNYmmoB3p4XZCZnNQ9tjWuSijfh
D4sT/AXMkfkX0ocaT0W0DAEUf43giw8DmmTHNT+iWodwTlYRrA9a14VGb3pJIQqkwUiLMU7tqZ1O
0rSMOW+o8lXusYKjr7nCQCW8/iQuAVCEjSC78vMQgzZPM/kP/HoakDZzARB/fTs3c7B8Zzqx0Uow
MAaCA9Cpk3xljRVlm5f35AeHgs1PCvASIeLYg2adU24H4rJoCd/Y4qYzapxKr2k/CbFtTc2h5HEh
b4HrpN0/cWEAwVi7W3tOMgVD8BgPb0GW2NBvovTaJtBJ1+k9IpOxOUt7NNTXjhN+pl4bSFyXIykG
tp/2gOqGLvl0yCExDdCFCXgDlcU5+vinx5NTB4seP6vWI/lWuUvoUNdKzL30cY42cwd2N1lPSvOq
B5FGFnAWvte5rpizAXiVVwFH8wBEffzbFt/vcNgvDI0Iw+9xg/qTHn/UI4nZ4i9rJuSblC1bbudc
K4pY9CRCt/ZOPvLL8mHRga0LByuVqRzhAfHn44X0xZdWNEzP6qltDLKvGfw7HfZXa4oFVhlO0XJU
2wMUnC21O1EOTkePgIC5kgW4Go5MYHFw6M2yFq1syJ+h1vXksMONxKBH+5CQNxNV5XD4GOHL/QfC
z/fqAkjtWDwx/FazQoDWvDLFF7i/J54Q0tRCJkxU9ZM1QkxMPt9Pasv/ieQW2EcjL0Tn1n6PEnXn
sdlqvE/jUfyEGChd85tsg/hLWCqkOsqEfdbhkqb1+ZMmUIf9NQEWW1vcwrzpnFYJ4GTlEE6fvNyS
Ct5gLgL/24Tdu1sNvOW4f9fKYBrFEhvR2a2ztISNStBVqq6qw7+TO+jTQZkQ9ebTEKgAUeM5Zlsw
upzVF8A1SPvhCZaR82icDdCqonYl0Q8h+ykEoEkjoKFXE8qjS+5/z2TavJsGV1b0FiYZGefahkSj
2F4CcpQ/i7UceKvaKCJIkphEdvCRwXRmhxzkPm/YjuNod5COSJEVZGVII2GlIadXAgxwnWd00u3G
sxxSSWi5qRWb/gPmkPBcxRY7vQyQ9iU8kUYWV1qWZVIadlQ8x33JPwA7fvbOaEBNJIxGtSDvi6cz
MrZ8CXyHf9NEfkkHib6Lv3cMtbKncKTDHAjPbvawIlu/eHUUjuuGxN0SwxrwzTcmmalw4u0bSV5P
ToFRfDoCI6OABzJYFRraYgRBjc6DJp+mXJbQOq4Kxr2Ay4oYgQwcJ+uvx5vwT3bI2beHJNtfHPXA
Yv4caSp7us0pxMrFbMfDYtqHPIUK4IQHjcLGgDYjBi+UAs5O5Pfstruplc4fv+auZLz9+yJk5eiK
njxOL2mrvMagSfe3MUI+eaMXYDao7E9F0CxVsJ3UFzSdMnGh2RYuSVm2zNzwLNRn/nfkF04p0OuE
obpUwLHnjSMcPdO2ymh+iGIIB4eT8xymjbsHmcO9Twnv9w9/0204KOivD1uszNrHgFSxwJNe6YYV
+IDucarVX6X9tJA8OD5Q9WLqTji3XqvdsapQ77nCMcOTDtQGJ4MfNt0jbm30kBKiDXu37rou9UoX
UxKXzbXwwVU91k7rOC1F1NF7xhtwtPD9sWtNbRYfFxSeb0I9Kfo+6VcwfiRIx1rdm4izIuFVskeF
b7qiSpYYD90PocT7opIE78ZEXXepPeVzKTjsJf/4PJWCkx5lmxCw2X65q8EP/kFKsuZJGVZFcKNl
8d1fG13GySrWK5xMjFGd17I2AfwsQjIKwAuD5IU3IM6/EmSEU7pNPpjSPS25jfNBvu53kzGahHdU
pEE07ne+ICGxDGNsL5TnIkEz2beEvjuUGf+L0yjN28hlVpO7ytm0eanz4nsKes45xZCCik+Trg6i
JeJ0AZH6jpOpAdRIe+0b/XBLQJUhRSJqGAaPdBiLGvXGMHzRP7nhL3/jz5xlIUY4CehTOgT1YMgH
5spw3WY52EeNzJ5l4Ak2K+zIeCboGHnFeyLKK/a3KwlqYIZfiLAJLAcMZ/KbzC3fPgpYpnWfM1nF
aKdDFZD1GCU3YbxJXQmXfYzf/sAtTuQ7nk3CSiaeXhKcol/bbvltXiaQeZrv3mNNe+O1B3d2gA9s
5GgNRgvAl6ymZNTyZFf+/DUwrzZMrvYcqMbS+yDdl58+GTMeZoYWijkU2nOl847XDCLmAnTE5RKp
/Bkj4XWU5UDzcMOaj7LdOBqNmANiULBbvARr9g+jSFcgPMFmBQ/4/MvOFIgukPK/V2ThVrRgT1qN
nv162ymk2/5LmfZX2+ZJq7f1TY7/INJpzGDyVrL+wuFIysdMo9Y1R/2659tDqZFSRiw1+UPDsIbY
KnuMftyQyXGc51mMPVppoXShr9GzBce6YA1CYmfP/4i+frkg8trYL76m3Q1FIAtcg4Xns8ynxUwP
NlY4KBH2zUQ1O7PwVknTYKWU61tjZBarFtmPycFPlS0FvAjRfqbEPLsEieQUvaxq9wqyZoVrBILZ
E5llEyyEVLShQpIDu95C+JjvXzopJNDzIqvCkhgj7zJNN6GGlT/oYVfEZYL2Z9w8wXvCUQQtmoeA
hcqnbbY1Ot3zCQl75PZHLTS+IXqbT09FMasm7W5MmYmZS4Bx0qfWxxS72zIiPAi1jJmHLWfq3vED
Nmah8mL3spvBoIN2MAQxOs5TPravkCmSXIYULqB3dp7ivVoqYppuwqxkYq8J0/L1x8OEvL1ROTz9
6Qcy/00iKEco+HNvu+M4mXZLRK3Vtd/4y1c1IiL4WkFOpimH2og1dvh+QpgmqheBKEOiF+BnS3EB
Jl7dax45b3deDjcf2q75AVib8y36TFFnTSp0KBsUuHY4CyWeVON4Rrtlr0ib2Ra/RCI4f406YWac
cmy1kuKXRTyvHIdKL7VJTaVXQ9Rw18tViuKDE/hP3xWZSOvRl4c3Bahz3P7TgGeHYOCkyXOLitqp
kRpyx1kIvvTP4byF71DXDnez6halEn5Cj3fxugH3/qF4r2jyNPGHBTHvVj2axAraWPnkKW5h4Jf8
FVfCBY+Dbkb+xc11UIo/IiTbJklhBS6t8GBZLFcBw54KwISKD691T9MjcqByEgajQGRk5gZDSx5W
/BisWxR8O/Cv730YMjvR93I5+O7MpZvHdgXtzhy/iZjlHdHh+Mx94nfgUMwUj/2xgy75zf2gFs2Z
fJGq0z9kapkgx5PAFSKAQWnQ7DxVnWMTjzz14hM1mzZi//6nYHebDY2Nux1lvtoAq4M8G5ZV7sv8
MbtrAH3RgbKy36el3XeUj0eT3ztZVx2qsd6k2y+EszwTiIeBF+tssI123NoQr2y+aq2QaFtM+PBi
F+Y7ftivkR4MqPB2nT8ZXxxOomWqGA7dEJA3u/x5VauAMqJdVsQxN4D8alE/6pW/FnmzGdY/SrsQ
zD3thNjaZqf2rVygT2+3j5IV7yQN29ws9QMsdT0IkgYAoPalJ6T15fURXgfxrRvItgg3Y4UviiNy
3B93KCe7ygyQcCoM4ITNnbvFwGZeTfXY30FCcFMY0A6WqixTAJZ26JUN2tNEZ+A7LHjz3v7220PA
OeYzXeE/dg40Ro2fv3iZcou/IfwrPazsrDKANVEpDj4S5bbue5ZcTOjXdXjip/5QUGk74lhsYCAG
HdhvxcmVgMwqjLlgP6qEPDhlSsKyIGX5ReIpEbq2PinQ1So4/V8TWOcPZQ5qSe3H7QBksltVCvB/
kvIUH9kCF8Aow78OMzOZi/oERT3P4yKSHxn/8HcByXve6BligJIS5DMMIg9J/CqrkLt7/4X3FMhY
2f6QfiwcLN+X+GhJkqllucRo05j7LRjs7GUkefgsIBJ4PUOrkalLXn0YnusL4mhh0uVsrMH09MJr
1JWWzks3ldGrtiJy4X2Kg17ejTEPzFj2NKt1XnG16iDhkOhZ4s2wESqfL0dj7VtG1sQgxQkQx0uc
l36M+SZu0q9lGqthoLZb/GJt48RAhImaIaro5VutJSbGAG2TywqLgoaFquxeFyoJ81ltzXX2fhlr
QM7Pr3uN9atL+zMR5rVmJ8pvYxT20iMY+AUYrZfk9D3oRvEpgQUs4SXQ14i2C3ioGM1BihuWmgdB
BO2/gAyoppyiCNQe9TaWKaYQ+92XgdYB0CoZoYu1rjzEgeyamtUXRglPVNQDZeluKrQdQnQXHfCk
lxhDcH+lnMMhdUjifGdXcam089Glq1l2yLWO5RxwNML4Vbcgb5JzwoDOtrlIqR1N51I6pOax6eON
pGtw/jJfFgeOdPZC9mPljlRhrxPUpIUUHcK+6fqhNDUjioKzDFEmz2rr8PhBqSba6isKc5NX1+Sk
iUn2IszzNkoL4Njx1LbnMBgkZbXzXAWDhwuimtg/wn89rNmSMJLZs4adc9LQkY5CYT/OVQN+TjCS
Eq92BWvg8F3yZNA2o4s3Wp2XnO93VnY/SrmXO/Dni+qy4p0JxKAGfMjCE2izO5A6uO2BCM7jJgSC
d97r67qP1SkMeibJRlj9kv85h7QUAGDER32b1oY3x3RL/Nvd/YKN+RGI/EAVnYd4A6RyNe4hnj/s
tmGvrNtwL+Uu4YnNhTrO5peAsIPdfvVvoH6X8GGgtKKyS9h4dDHmVdcNnc05yCsi7Kr1b11Gr8eK
5cF99TRNThSrIP7TsXLtXbDvjrG/3+1yYwsTgB1asthsl8TwCfpZnr6ptu2LbahjRuHgDyxT1OfO
ZxaLrxIEnAOiN95EE6bINHvFBVhpFOKbVIcJSXUiXE72LZQ5sdtngFYV1yRgfDPLIHJpCUs0AdRw
58sYMUFQiGn3jn7qn/EfLBn+pYujBz0bbpeePjNe+2GAteovo+4nogDX67AGTzMv19CE6V8LOkkf
m04BPuaYBvkqvngdqOxH1ilgDqFALKcqAKQmo307XsijgwvoRFSyqiY3kuVRVV0OK+o8fJCp1oJ4
oQETMfnMzDDp6xVxt7hWUuYTV/EhT0VJSSMndwW3fC6KnhZ197YhI/zhsw8G8A5sHLUfpkZCmD5f
A9xZ1YC8APsRlaCVdd0Z/JfgLzwXk41NoQgAunCsumdlF8R2lMfS3R1eo3I/53qVybP+vHQHmRuN
cVAwoqkJdzY2wQGT+k34VHL6ybHXnwE/sUJ4ulKuHsYDiOUkeXGo7qKVvdbHulNT8i13y2yBisVp
95BWs1ApQB6cPkRZwIhXa9y13udS+pAEvl4n5SuYZF6axQ/2rowfneLRcxE4/PjSiDPJW0/6A60D
TH4jeAFajxlUc4suxOihlEGKf4fR93L7KCqawbsy7U5g9JzXE1lE20PJUkD5DmxZHZnGsYU3oyMb
egh9A0hrK68J2+jRLcODJqwbVwE/M5Jn67qITIOLxl0oZtBGB06cisqQNQOHO8eT1vE2jjqIs7BX
EKi9xgKmUhYwIYNlHD4PLeHUgrTEcSMLGna+FfuAzawzoT5zA/473+rmZJY47dY3iUhJjfFYJ+yD
kiFdjj0ggZ3NbkgHU6d9Xgt+hagRNdRKZ4VWjiZAczfd6XV4hcQZ84lOyQdYbZhTBKvGbpIk7omf
eufZgbu8QdPgC32XEwj845HJRsC2ZsvraorCiZRm6EWgxpg6vlueFPUwzNa0OV19jLfqL+ljd1Qe
BXKsfELEbrjkxmb+sWuM1lfehZLAPXqCpGOjE2VnmxN3DMPUPOEc5grNHxDnpEezaN7mlKLg6VtA
np+rQrzrUhtTZ5rUDR4Aa8uaitR9Y+Lb+c8IlMkbhOClqTptpLkizJideewJUSm7ub34tNPGAhYW
Bwmo1s0q5FtJromIbMqTAHjtxb+S1yEBwTg3vx1OGkvo0cgs/kIfJvdVxTmikUMoEozHL6J3wNnV
7O7wV9xLXOa+QzbQx6sB1+hEPamd+X2Wn4By2yJ7r/+Ft2UVM6i5h5HS0I0bpYRN+gfihyJCWIDc
u0zmF/+UeRQv7cPlwdjm5IKAZxhDZianjyHXwYXfsQ/TLMQ9aOMtkEr81TOd23zmvNbwsFsvm/q3
2qxhnaPyf33O4XDcVF+P0n2eNJ5sxsFtqaZZ1yXWYST6eFaXD3zJiTp51OSJrySwaVxXWyLIvoGG
KSZAbw90XRUvBjD/la3L99nDeRscUapyI7rUBrcFq4eiX7hJloKRIyOYcCk8jPurRBLJ58GHsCwu
OhSuNuYlCm2JB4MAg3jXn/QDnWNh5jDt9ioT04tfTktURZn9HBLbNaoT5qcBuNLreY5d2eMwusgn
GLn0W3veeBGxJSsQCSvGh1EE+z2yxR9PlfKSGN9H06kgjBV2z3MN8K9WXQQCyucKcMwbw7nrzwgP
+jlV/QgdRnEnNNOayzfpPhisOBESgeOgLzI2RLgu1URlYBskRRx7rGkRHGA5Gl7NF4AWPgvAssbu
Hb+Hr0pBv4S07TwwZ1J01uVrmf5EX3qpCxSvS5j3+xTgT5I7xW8RnRyqchx5culTU4wp+Id13/qV
u9EGH3Uz5VEncuXGPgk3knGWxsXgpRydW7dfvrBwSaZ7fz9n7v0BpnuxmnAqJgGSI6FY0kdJpSDJ
zt9AJbYHAxDUHT9ufmrFSKdqA/EU/FFJUCTF68SApMLCoQ6mH0ofKYayApfXkstR1W4CvjNNW5Cc
iYcR/uyH9qTtVdeuFe4Y3Ug0FIpMMhGAtXKGa2Gd+ttm3ahDfys+V/+z+qUayM2xriC1KbmF3eCZ
9Uh15UivpvSOI72TjZlldCtbxZF1eDp4N0/XfhQYUFz4RqAJI2xpzM87pMC1V9dAA4jN6uejtlD0
I2rV4eW7DBdXdjLGW1xx/K0grdkE6QaDPcHCsRsJVX5dFyzyTMvcikFF8V9YsQ9oGT8+CsFhFVCg
HfSd0LPCMHgTON1QETUy2EEaTuKgO0+PFzQI/QHXINFGLis4AxwHFofmyCpKXayF/vSzVJHMdWe3
U8T4PmD6vLOD0znxVbZFe97pvfMYitGxG2jIiCTehmkGy3LnoojQzBmh+PsFm+WD1DH+1do4TncK
5HgWXrJgDOavhZzFKqftmvPY5z3Evt3+uLk2rKafkvaHbBW7cdA/oAi881Sz/+e4ZqUsNpVloTwi
r1YfE4+RbtZIpVUY+st0C0OX4dbpIeaEzH5z/rh43aot9UI6piyeWwEUImoC5wyK9qHQIZTEjjHT
RHk8+q7+ukxmzZ/lW5kkG9Sf5evYuwIJ4qTn48FUl8LXm1Gr9yoQNARS+D2NFlI2DclO5NSVKBJe
bQWyGxJV4onMMo7IdfFAeM8E4h9hqso9H3j05ne+1Gn4JzMDY90eIwRYvHRb9m/cPbM0AphM6DBJ
rkBEUY8O4ITBsVwilVexx45Ildi/1nPqeVBQFGUXKFF/N1WcJb7dzNtIkpn1w7rcjcWg+eYZ9vN+
HI92TlQRTiCsJSS1QwZYkKJw0rqcwUX7rOp453AgW8c/FoYeLz0PD9SpE1Hkd/XbJQD92koi4O2n
SRjtikwTOWF/vWfrPXJDOTxunPXdHuL+GS0ijUj+sJEbMbu0Y8lLSK4aHp1o/twbCZIU7romz29v
zd++k1MaayYnnUNCH2QymAYUfcO8pGo8oO8F4ZYC6RutUuLxk1dLUuq4tZ8JKriRrplcLTOfr4jK
QJyg87/0f40K9U3t/aldFbQO2Ank4oEznWx24FCyfShHTixbD1HGEPt7W4RXtQQzxVY/mOo294dm
Kb3hrK58H2NchJGufch/XtEbMSlJbIVnc9yyARC52EKPYzxakIy0QDB0OZRROPJmfXi71qxuW0R+
Vj7aLTlLTMaaHy+lY7enocxLFTxc/yIt7GIAbXDrg/pHZkweI9qgdkQrkONjEkan95SgcAPUmemt
tG5muejt9CPhgYrf2UKmyDUQvUZhpelGpIHO8dNhSAiQEN4moVyTdohZ+AYSe617MpHYkfa8Kc6J
FRWmxu7F6K4P35tcDG8gIsqDIkkRXuSPd6Y2KTk9GkM3e8Uzvx8o9vtxnHzGQ/9TWv6wz6Jie0Gn
RGx01cvri+jw7PqR7CC/x8+n56J6HZOxQCdwLbcfMPlpl1fIJz7OElpmt5feUMxAaeJhHsNDBevD
m1vR4AQuX7zaK1F3shzAm4NvOfY3POc6H7ocQ7DMv0k77ErgUaWgaQ1kMHOK8vAmubmopMWsQz0Y
A0D73iv+vzU2stfd09W1AJ5S7EJU1FRpu+gmSq/xR3t9boV9zlJpZzK55I0XsIZzV35/NFiGjpE2
qXgVUEjOz5GF3H239xlQ/CiDa+CMXegJOgUYef2s6/d9vI2ftH333BELluRLnIdRmCt9zi8LTof7
0alKsTnYzIOCYP1XluU+hWJdlGbwm9uYXmERm/gRqAuIMgX814MdPHH+AiLGj1YUkzo2ZxQzkoK+
pgiBDdUaChjqi2vnetRiCGjnAz2DfSRB1WF4VUU3tUyn2hTCNnAtQgZlpsClDTLJdIEpBBqqgC1v
6s+4RQGIwrhsbCUzdnPVSnbYr8lHV4J2UcYS5zSNyBWegun8wVxAdfBhoB4FOYH/BJFOVUuVvymR
uGgytqfRd//HB7Ei1mlAwEC7iVnihLas1T0E1qXl/PhuGgvovEc8JSvZRnqH4J/8uK7j+HjcJLjb
t8/SPUbs+7wBBe96hUTXY0iHzqDNjHga+sLtfvtlU+jWbGBUT02JsdMJW9KH55+5eOaG/uQV98eD
ou33OBcpi1MfthQ/uQpR2Al/Wjrnwa0+hDq4K6QWDoq9+1jt9b78Gx+o1MsY/YJdc3/9xw/i434S
FpSXz7wsTjxEiZKaGMC55EGaYQd55Qx8b2jRFohi4NsutKdIwF1gVle4v/DVXoMPiHaTHXAwgcEl
ry+Pehhwz34VNFEgh+NhRhy8gv79gtfJBAREgWFNozDvZmDWLhnT46HqdaKG2MscF9mqJ7gbxW6T
i7xbEq6Ds/KTdPH9aScZ2vlyS4RO5BykqJYLZ3QVFQ5TbwF1sNH1R4ErGdMyRuI2Pxfz8dAgaypT
Ws3GngdFnOiUTkz0QXNQ+EccdhBgbaU0cp9WndQxbr2eInl/BRTVJMDKniCCoolQKQ9ilYlcONmR
Tb2vrArMPfH1M4x2ID1VmWr9gzQ1yBQ9hOoa1F5SPbW2RtIaua1LG+9Kd4a9aFzEnTDP6pOasH7f
6gQqQprnh792ycWfK2nNnCDo+2U5hzwmiakemNg40MX2UXNb68tFO+GJCYTPXdCCyAbZOvLSzNan
suOFyg1Pfw5goRcQPBwKZrG9nDD23LHns4ek+JraESK5xKsJ53W3d9/30dSc48WvrQ73mKXxxXvl
pQoG25S+5pwcbDS6VUuOl+gMmqe7BZ8abqhtvCwtKwYj6Y89ZfFps+5gVs6mE01oA87ysMMfogdQ
rQaLnmPautsvSpeEdhTgNhNt/b+vwTtCjX2SI7As+dRw5FLchwgTww2P+37RB605+7uQIQWS3ioq
FV1m4AqpsRprBGC1SAUD2qKX8LS7t6C1YoFPathhSeitjzmPV8RIdOMxmHCZ+TyRO9KXb9BXkQxG
V7HoDfx8fab4DMJN9om892ys+Fg7tc3JUIoJV4wL1bj1KiU+yO2TZ6dGN76S1eNFLOS1xRizj3Oe
m4/126+bPmHrOaEXfZetBYI4lTogYV6ekhQz38XJsmCD4EMynUp2W80238uEhTYvcqgqG+g96vfI
EA4dM4ZuP1jAPDd+8m4t+UpQQhYIDif417xD0vRmwUKJ2/9pKEbJg+v9mFns0mXexVjfo5F524of
uoS7nxbr7iIvsinWXR7IMDKSLZl1rrOJFWxxq0PmM0mW/spjzKKauH0Sg/O4TeQveTZUIRcG7WKR
izPYmHONvofec1JqVUI6CGdbXw6I7AOgk7HovfVhIBmbxeLmAhc0HdUrd9SiBhA73l2wSoqDwlfB
m1Pz/LSV0RE/uayEAJl+HxPKIe6rGAP9Kw8XWwTFZ0M15CINc3PAxQitPrDvGF3ppQHy7EvcCDVK
sLzhKxx/pSWu/GvMDYgEoEXWinVvJJg/lkrNSOBr3kiuEVLXDL4VtYfIbpekwHtZlTdUAUWoU8kP
ZXXhceiT/rzCLyKD+N7vwK5zwwj+CjhA32kuvUSSywig1ZIEo5NgEa86pPHpHiTXb3L7VNTk6kiU
wnQu/fqMU4yq9K5uGwYnESOIMIW3RjuSggxaMm4qdA9aUOzVYGJMq00fBq4TcYGtzXUMsItqjgap
hbNxWRbTFiOVD0g3ZCRXbeHODxm/84QBIi+fASqMu6rWSdkz8n9G4diI1EDkJ5q1FWmHcuEAEiyb
O06e0l2NbeD2hsCItdizXcA3ZtmyKYO/Y6oSyFmql9R40uWHkshQbOoaaSVDhK3ArYnanNwZ4FQG
C/b9i4OroXAP1syf9pjK2glyHXHtzkZGnb1VEYPD0dcUqILgOz/P5/LTGahEp+kQPRur+BNuOa9T
LS9hkRs5aSfHz3SvOSUMk97xIOaKK7hoqEBdiH+u6iD+Mp9iOy8keP2qhhKB8Ns3Ry/b8Tn9iJfB
w8F1sCBsVZGCXsX5UM7CgHXPm9q0uHluhOVe0wdufmEhxvmB8/I1S9rlOryaSczZjnaEv813NqDd
mb8U66cK/322UDDRBci4+FOZbWPj9bmlpzP9nDMkHYDC4FOSg8gu25CZE+mW/wqr8fgzjW0qKyzA
23Mi0L28ZCl4PYBZqAWNasLBdyqlyZq5mKbCWgoFkmeiK0/e5xgsheMmDaqNZ7OeVbUtgpULbn55
l5WWcGNsgBnNg02ezFQnjdFXMKtZ6fF6bKYcXVLeZ72S3yJLq1kAN5a5+ZSPsMiQMyXCDISv6jQO
2lTT10TPvwbC1sQ8qQlCdGbZcb/jkYybHhGCkx0wJuIMVKKIbwlr1d/QbtwqlV29oReAtd1UvuKT
YD/0TnbMqvY/oqT9QiSEZ8wSXOxoJslBd2igSyjbjxEo+TCk9zjh81Fk4eHVYdF7NhRcITBNOAv8
vSNkrdluipwhmUgJcdU2E45mOkFzWcrtEL6Xw/LSqdhFHt5cBVdyMd+hI52HfslQshyC9R/+bge6
AWLbWzXjGByUeC+5ev2umx4wiMJb/Ty4GOlmQqpCUc1GN7h4LJ9ChLZD3tR84VPu6FndEQpu4qHk
p3fOb9wqY6ZeBbdLjKmyvmx7ZX6Ufw5++li0ozsE39bGgl6mHL7h2jSuxec3Gt2iNjX7P/aKb21S
iPVrAHQkA1ZtIGa/YppBMF04K33MGv/u+z1anK8VVMDixcZyqBPqZMIeBQREHwifsYYF+yxB+h6u
7+5xQEZ1mOAAb2XTdiZ2pHqzvW79UC/Fa4x8lZAZMxF8GASBqY3W267I/qLjo16ZiQ6Xq3x/67fC
RgpkQT9swTLgO0ISvaJGBTJElQAFhPFF+uNkw0+LL5XA/Jh6PPiR3+WhP+YYuvqHdfQl5bWPIiMf
B4YwiasdoC5zmMCWTUvA5C1bYD9t5ttHWYqhHeJ/vaQGl8vBnBQpEWfKwBNYADkf6mirj8DDdxA3
4PikQdkFm2W3Tgw1tVKnG+810zmF4++V9saVnk/zJ15ZxSu2kHaoaHIIezK3gYZq5XgbQ3HqHJdh
+ERNvgErBMI1F4jLDAhVlKr6UUI2LC5E3vpypIZ8Y4RMB8ezOmPmJowypREehA8XJPulc807ZRMC
KqDuzyY/SLlHyl3wPVT/D/fsxMK1bXgjZpn5YkUfqNWxKlD1tBi+TFPf5BoXE0PPZUuYfNkPHuSv
JuGKR5NJQEALQzognGe9JPyfnV+jcPkiSp5C3Dr/3XGwVrDAfctAuPj/rlFF95dNzPST/uGRVs4r
OVDaRFcY3jfmS25IO0FpuT+DnVzdOONfNx4eQ1XUUAXjlWgsfDlIbUwZBygwuTGApbLIoz3LRYyD
2zOSMCIPuhyC4Z2ebkRIvrlZZnXZ41AIAPzfagz7DhcbWB44ZRkHlit8TUgpnCq6AhJmrf3hZLuu
q0XL9S5YPg502aOXJE67Gcu5t4g+j2iwyAyEwLTviC14hWgKFkp1F8gpfE74WD8nGmn7IQxGbxEo
9XtKnEH1AYeuJnM2SKvF/riYic/E+EoOgmYul+08wMrrNfkt2ro/p0FKNcBBxzlFzmPLc/ns7gJX
R1gviNnfvfgdNmWUeWTI8DkzQn1UXNYn+4zOVly5SuY7omMeVpmNl3usALh5tFcNn86qJLVcxP/l
Ocqc/J0nBhx+SIw9R8tqAS8uO1RHvfYW94b1V0WowH916RA2TKVxHdh37GiGdYEHHnEE0zpjePTa
9M1IUkSYQPeo+1dLRd6oCuNvvSraQEUmiVFZw4QsoON7CxuI5YDDj9n6mmTGfcUG78w1LsMLFJK7
NjV4q22limvEmXZ5HpLJWAr6AoQ7DOLuO6BbaituNh+Y0v/yXeX9BzraXKbYn6HVOOG5Fe/rRP+u
49rfhbaRa+klZ1Cb1c/8kSuv+jaa5tX/RZ3lyXb3lUlQA606DvTQyrMIUxxVJgKnsglohey/UKIm
/4aZjpvC/E+B1RycKFwgHGeYRJEaMLf5hh9e4a513epNEFMWX9oQAXDBAODgcFFe9qfyGfSUqSmC
rv2NY7zzmhB1eXwcJScngmxcl+D+WMn7xsbOcooxPprPf+uieMcBfRDG3pcXiyX5/g93l4enTV4M
iA7HWADUJJFXSE7XOWMuKBv4OlYxVDSVDX8rtal8dft+wK9X2vVVLtL/UpaU8xtdPYLQ5yhwSVKb
wigia+nLv2IwihRJjZZFwzLRaTBwepUL8YGuxcxVa0a9NKtJZCJobFlRefE+5npMdqdtlkoOavWe
Pg0I0M7YTIQcmWDcfMpA6iHqaEqUHvLe3LNDuyG3Q+wbNiKxlSOS8A2jDcysETMD80gHsr9+2zmB
mo3ZY0TTmLT+ytyEhlyubbiG5rR43Q2+yVwoCO3gvdDorz0ATG+K1Xq5YBtYN2DZvTAP871cIBqv
9W2FakaZcreeQMFbOZSMI+hyux4rtQFnsHQ4TUTs/3IxR3aYAFyz56nxRW01LtHSlb5zPFZRUx/y
cqnSXGhYoD7i+1fhyZMmCx7KCejO4xF6QKWefKBmQEWIALL1cZkAsIYrOTkCN4pgcCwTppwPolK0
Fj3400QmP58ZE8QbP7vj6UuFY4APLqpH+y9p65Vgwxn+j/3vMk6NISd4ZrYmyQU9+JU4F7at4xAW
gI1wqlYcZZmwMItiDepG3fIVQtJlhh/yu2whyDTqYvj0Puxx8w2q22atx1U9tNgAn/iPMPchvVEu
Z7PDtJRSFG7lk7obE0hI3hkjf0fjRcFCtsGykZckGwZZlnHInp1cZ5L2SIOLmlPvCi5/LsD3QOfJ
OfoZsuv4CR9koXRyCJRKVsHOgqGXnhNyIOFh3zbjrZBHc+oF+6vhgaHw5vBHKOwsbPpKEuEDiLGW
RXA+6VjHQ6YNqEdkjCQ8ST+as5YjoPKQWXE2juwSr/ysk35mB17RqSb/caVlQhYEqBCYZyPfA4Vd
rpqf/psDso3zWKuQ+wextDYE3BZS2slZy1eGcTFyLWnO7SlDGU+eT1uuXK833+JvgMvr45GnAyns
aEMOFj66b9LDsYE8BMZDzsVMouyQaU6aXRSEg/f3YDdVITKeE1Ooosc3p0z3+x15Ck+T13+PvaKK
ePiddLmO4PKvilvOKWlzyjyyU3rUo/eNaO2HpKjwKQnT04YNnFJsLAOyTv/vHtkzgMn/7qYwMAs7
5I0lOtn4h5X3ZBljiQnxfALbpuy6NflhImIb049hoRcArJt9L6czKNuL6dVvj2r8haLa2VMeEMF3
biM68yovhX9zGju18yxsxl8LXk00WVoYdiZTFYvJa5haSejinwf9JLF7+QkYrxjOXoVz0rkY7G2W
xbWFo+LmzSvjP+A2iGj8IHRQiyjsRAM+klGkF3vkwT3Q70RmLo1r/U1qnHciRpdVDGGY9qypRkPd
ymUWyiba9aYvl181WLlms33aUtxbtc+//pejZHsHs/SRXJ5tM7kFVbyWE6dRrCYedtiuQ+xn1aNt
uZ6bxeVLLosUE3YXEJiY0hhRrzECpPbPZtJxdv6WR7EKyoBPA8Rv/X4Gsb14w1UPorZzxvaS4lsw
ysaf6JNgTWEa7P5M1onSTtaaFdN7EqJsc5MnEtAVrckNPSjGoZnSzh5MSEvtGOvfx/sbwXEbHXe5
zyINAsqopeAPfmjGHwZ7DvdHgin7OnQACxoqitrLh4xbWbuT62GNsE50AEsrypp2W9HFSBUOIJdV
qcz5RhEthMh7YafkDFRWQt3bo35Cu3tRnTL+v83wg3NqRJuDGilKNoB5/+stZ3F+3D0nF+rYUoAX
IvYcUPDETuXtsIWqwSjMIBRZqcKiMlu1HpPvwC/MKBFq1Dee9Zh+Rlfu2bIj1GWGMcP545vwbZoW
mIqS45CaFEdexYBnB3tH+Kec6Ynn+cP03IpJlsM94anEFv3zziTLUuDzojS5UJRZgYbUth6BMhaS
gLkZDJA4qOV4fSyD5J4WeyPqIUtkZgdO98RPrTTE4VTEa2dQhwBfk5X+NQ7PR+ZzCt0zSixLpqGF
MfuZX1dQIAlb1GLSZOWuq04/8R5c3xMifp77QdLsRdRtYgrXJBMEH9iDx0yHpg/rKWa1aZgkSJ6t
e6v133cGNXNVawnBQkwQG6RPyGEcNbkwSoxzGvQfATclxmpetOr4pwwlWW22sdKQNExYrfy7z0CG
7g5WHJwwUpqI7uKpLvpXu2tpMJz5nsM98QNI17GmyNkVZyKpkHwJ/0rw1lKjM4DXP4hqYTjRgRoi
1hAtE3naCqaWkBeUs7sPOF57oQmRmagNAAV0ae1xBUo30+2STILZm4JLUiuObwCe5frQBCcHTnkU
nCURO/sNJo20nVAH8f9qxJDdtd4l50akZcFoiMxRD7SrxkMMFfOyeKggAcXBCcP1l7FuDATgT87Z
Vl6iav/iM7h6oJJaUUIWtOOU5gXmx+cQlSzwwoIMWhTUit8NIKRBaMYtS9/V5L2oCOJpLTc+Sgn3
SfQmMFJol99FJFfWCRspy4qsiQ79+IR59NNOf2dCMemkpVNLO9Np8NuaBvQSVIxP29b67eQBK8SY
FufIcXmTPTEh9oXdXKq3qhRfdO/gnQiAXkEMWXYLzlpxaPaj25wOWe4fP9CdZKt8Qj/+OySlERun
Pk5A4QXhdpGXgNMQ/NfTn4wpjEbqQiPXwWTHM7XwyeuqJJeVVqnCr9mXs2DScbD/Hrik3T8ofCQe
63JE4pkXS3scBpHKl92uGWbmSow3RDEWmzAxvfvto35sYG9bjD+i9WyacLScCV6L7CCBmdKNXNDE
pfasyqmdrkUjB1SlpNa7/l+R06O8KG0U1HUKJZ4GpaAyQrkoRjr1rf6QcH6Ak0FaPQZMnfPe/8Bc
T+81v0hUlUdWuCcLy3jEvkjJ0IVOLSWs0fHYpXRQZEZnVzzGwrD3vf+B4YVGbQIOdWE1kIAuYtNt
CRAXSrOsCO6G/Bljbb+t2/qhzXqNDpjPol2nYHWFRV9rVXio+/HZcbVqx1F0CNvN2NlA1sGR0z4K
2uUw9hc06bwohelSbmBSnvlxAVlYsD7ApwofxbmQWfbeNhO08+1S3PcYOSgULDDgm/i9wYXd282Y
J6PuBnHjCvKTngG2rIf2tMotTTjshBgrLajt7npbaqBMrDxZqKZmzJLWVQcWtm93nRBhTjgN3byS
iRVqoE4g5pIisv3GoJ81V1NoQ8tBDHlD0kQQK4hKUY5cuPPxkHo3sT8quSMZ1B2qv0v8SSY2s3MX
9njkuJ2T9XyEFxP7ihpJFWCmz89nTNzPXUu5JioGDYLoz8XZhScCkh2kZMkNbTiRPw1eHlw8kA/y
l8YW1Ff4VEHukh5FpD5aiw5pBxdDJBLsmSCHkjgvDthQb6zAbRR63QfwK2n7eXB0vVGbr0GeeVFY
G0wU3FXCy5Tw1Kb12Tzc7MVpnDeJzZ81JFYxC3BL7YFLsyNGF0nrVlJFUIii4awBNP05Kb3KCA2I
05wKZx3Fssxa3uoW347yo48cHmHh3q8kqje9QIm+7DDKCxbBIhp/eYq5LZLhso54IBzq78ECCrRQ
r2YNeybSsPKUyBNDsqvl7vKNaNgpOtOeROeOtf0ns0PDeJ/Tdm48s68KGQCOfhWOHl2dfwTIJlaf
T1uIMRdEyy3zUEYNegmQX72Kfay9ZIMMAxQOfiMtY2suSiw2Etjf+aCW1jVFo/1q+gUmOEDnHfG4
8kerpw4Wchfue/ICXYjjW536/zVhyecMaS+V9eAc8yJaYPgvmM2Oesjv3GoYYlTE1wAKJLoHtp1A
Ru9tJTTih0AFoUfRcZPEhuMrmhAAdbO734KmfeTTQOIaJeORxHdlu23lHeVNJPWM5fBguzePTcZi
EiA2ozDBSvBE+iFtMlg2z3Jpnaw5FFtLBnzOtw2H6MZrNibiXy0hzc3XHRoQ6hudl1w9e6qPLWEB
lhyPtBUbiGw2RXfobhx4oK55S/bNLmfbowY6IS1lbUMBlDvD9dm1Jhd9yD3Y9a8yN6l3C7QjSXSr
tTkAElbS+Mz21EWM6hn142NL4jgG1UUodcO1nZ32jghqCUwoQFO/ysda2Qa6TW2QjQrttag2xiYC
NX0KqyNK6pI3PO46HU8RIJHd+M0gX02L6cIBQ3TDTfpUmlISLJJ2cfHDkttWF9RhWxtsN7gFiPqe
MhchAA5OY6cTD/LXOL3vszkwqj7411Bu1PuXA834wZdU7MnWe8BD+OKgQfuGsEzSKuluuLZPh/ii
JQj3f5h9cwBjXGLqvAhBeVEOgvd14nR5qET9wWcLRFSBOjwLxL3NC72P48aar1N5h8YPhzI+SDa/
uZAXQvUBuQ1kYtzxP3OS4I56yMlx1GnQlGZwbupPVFqsBWRzXkE8kYZkf6cbzdDDWii6kHW9BO3z
dHBoI2Vt9gnnFuGc1IxrvUMep3ehG94kCzzzqlt4RwJvPqvDGAKB+lZePf8/B5Ub0dUNsvIOcsqN
VREqQQqIjH7KWjtxbXCEQSJ2tWdaQGwkhPcvv6v8laPBx2Wm/fn/53YvfXbGXUgzWu8PLVh5JtlA
jWD7G2JjPxxFFtUoEkuZJRm9dIqug1t7wv18nn97vvJ8JwjixgDGXKZGGXhMMTAPF0MMxY+wFqay
U79Lxh4UYjYVtGOllXckJit+VoLCgSACfrgbPs6Nje/6kaGCMqQsLzWH0uT3tskKk4DNAFnE2NIf
MAgD3IMTFd1G06vQA+yLTIhooxlxbnave9upb+uQFiuWTgBAu5YWuo4NoLB2H1mokohaW09evP6T
Cu1P/bmMvtgytZofelqKwLfc/KBMefFsmSNhLFa7lhN0Q+Ecgu82gjDzN2qBuFSJi0+pyTqB3W0m
Cc1wy63qohAQD42rhcxshbxEkWxG2547NFXshTwRDbofDrXKsO/wYDKSLpo80ICezS6bMQm9HYO+
yN2crAmxrn68wCDpHA8sny9YIRuHIK2xrDp+FgGGdtogXVNQslDGVCoYXVlrlhAKoKXapbZrGrKq
duCpq1nD7Gkq/5xHg1OYP6DSzBGi5UB3+k+1iyVlPhsK7PXoejeg71SJi5lrPhCQSQo7Z3YQ9g02
49ME6UZGc5ncIH6cSCi6y93NrgmIsaTrlqwv6J9j+cdKSW+dlsbDDCTUs2KGRLIqYTkBUq/RSRQV
c7vFd9OHv6H97Ah3EvOWIkxpZdsisVfHvb9hBnA+Ld6rE+DfLaKfYzZlQyAXxM8E9Bb185dzXRo7
YXt9wUJ21WqCZsqdz8sqdftFMk0Gw1/zXCLPMpch+nM3zLnnzMljuY6j88h7PxOH3x57fwrCwQwr
DVmHebQ68udvoidRGq/4zMMjWeXbQC3S2ieB1YGbSykFjDeqZ47VeQEIHkNo7r3GVVOA1Yd+SiyI
FIj9CCKNTEuEAj1UoSgZHZw9ODEBe30T89O7WavtGidV8SZSWwRpDBeugg6tmNdKcfbW9dDAZFkI
EmfOOr0rRVLGBhQBT5xYp3kMHI68/5oqDO3inqDnFoNUJgJgkklShQyqO8rYFulxbsJFPBhrXA7j
bL1Fv+dsBv9ATiMo1CO+WrQZevesaAM7qd6sNVTGOSShuIr02kYj0ZIa+3XuqCTngnBXxzS5vpCr
jiAoQeA0tLDd6lOmqT62iJaG1x6CUgHqe9/o5Oi3+ezLBZC8by6duWYIxx81wQbqlGJGmgrEGceX
GR6qRHxW3ETtgio4YuJJh3CUWK5eBi9l1CjHAjuIzUsOJ9xeKkw8QNYTo//x6eaMh5HZLA3+eBli
8IJ+pUJxqh1f970Z5Qpl5UOqOR1s/5qW6nXlsmA0cQpsw57GCOwVyGGA4HHMQrqbBTkYN08ET6OU
ZEmv0g4UpfBQ/3H4HXp4VVFsYyu0AckOz4zUsi8bGfiFsKhyY1Zi+NixBIRED2gWMCqKt2UndHCa
c5HLgUrsQ6sDspY5Sm8uURmL8s8sB3WS+1L6KCACM93rfOXrEdZGF4CdM+3DsWGn+/Ji5l1q6WdN
G4w4xuLLzKoZPD2MLFS8p7ZxNNZWptBGmkQL4DnjoeIAbNsBvUtuSluA4CGRRyriSCoXBihGWGd9
NSEX/enD3xT/MH828FfLDEoEFSRZC0+us3svVT4HZWm+h9C/cgGu9q02tlm2ASSy5LouPV5eNur6
W0Wlf4LK0vjJUiWMbSbhYVmKiWal78hSBhIZUsWLE7IY5zM2Gvg/mmhopmner6Gi0jY+wul9z4lj
KOM29XGXw+5elpxGGJTWt8kt2bxMO1qsoMCp2r0Db1c3XcQeHM7QNBA4zUltMl2ma50q6fcOWX/F
MVjd2qLZf9LwlDZeZ2RGZ1r7Ysm4pPjdLHjgqRIWMpb/6f6RgG75EF9CS7Iexw7h8blqioQoCg+k
eKHFU5hNBXrfkMhWTODGK4L/olof8IY+NKIx5QEfXjgq2ccJcc0oXaiuYzrast/z/x89lQedL2Fn
WiGmfYCPi9Z4khQvX1YIxzECqMv+FfhXVL9q3fE+haaJwFxr4G0JqRsF0hZtL1RsdBzD2P9GqIcW
qaCfzAv9hQ/ZBDerqzU/STiJwinU1EjS8i//7iQC0GF6qycyUW7vJxW05im1/bZ/WvD32URLEDE6
+xaTSChuQZCthnHuQ8ma7DVuXQHa/OymmyNw+Ia9uBOBlOZvY95vFSS21rf7PjjtcUtD1ojlSA8G
SJzGuXMQ1kJmoQaxFRfC1vx6wVQPcGe1OWr74FMy+LjrzX1diaf90tahv5QfuVx928lDH5w+RNDF
sue5t8gluy6N7hjr7wxS6SktGcD7CR9V6pis96tR14WxIx1QLG1HAWw22Xl3kvQpyyacJ3TZhaNl
nQpWweSyWSRBjC1Rb1sGOpNiEtaw16uCMsDm29hENAPriJwAnglr2Cx8b0D06d5HgxplnyDqiUSR
9xFJkkPLLgm9D7gFR/zq3EgKnUVw5ZZNQ2EKcQXzMiZpmfspX/XCbscl6vS4dWZwPYWskT3E+MDN
dBI9dQQSCWYiUQgnYDf8DrhtaWQYXzBsNNl5AnXD0+Wvl78qROHyjoNKJWViXCSl8WE1DLdnqFI7
7IGqNEPlK/o7GMKflTXIN5syyNGuVLR50Er1H2hNM8ObGzAI31QG7mrqZERRPPK4Xb8ulci/4NJK
nkfyPm1QMliniAEIQ2axnhqYupqowcUHNztGt1UF6rsNv0zm0NUE25iXKkJPvuEEcmwez9PGdeid
5VjmK7lsapDLivGCAuoYf3qzUnwdz2RR34XgnqbLvVT8fp+WnCCmFcildV3IsrsUQsckY5rIFJWk
PYGG4ig4mprlLVYZcuA2tDwp+bLNVR4jO7dNsse2ubekBYo5nD6Wq269tjVKv8/EymY8akRzaxrt
l9dGMvaWbFAYXNDzc/ilOiHAL7nvOM8q8IumfLPTDL3HS2/1dwQAFRdq4dwpoDCKZInB4I1ViGD1
S5eee7LlvbAhCZL+IUW2YMWk86oUE8AkZx7Jm8ZHhdWk0Ry7DgvOWMwxqGxBIBrr7w/eo/gzFPgi
ykA9iaDOfRgpmkQ1TpVqAAw10hUxQp8eKX+I26NsfVjMC0d66CHnOKjW/tUjGqcEvwB83fpzjtz4
lVJDrmCy5Z2xtnlw3VCayd2tFVOkhTgKmC8EdqL3bnp9NUOFJi5AkwH0XC80lgZIlvKyRgcux5jO
1d+LRptjS/qnd5GCnXf83xBQGocd9G54ty1L8TQy7XeqshbmqTqApjuVF3kCVGAljAEmFpnGitKi
EZj2XGVTU/EyuoN4xB+ZKKZR/6Ue4CNIiJxOBF6vCiCZL7D5CIAAd/uxCV/mf9yerOsTlhFnv3tj
JI56zu9PdB2odv5YQCI3jvvaD/Otl/HPlkeJLJRhoBhDv4QXd3hgD4X1YtMDSyDoFBNAAYWBbORe
CFIx38S1VDl5skh3D1KEZG9r2dwv1leHvBOeOpBYw8p24iyYxxEzbt3VR0PfFi/36gWqZrW23cJO
qAGnAjIr1Q9e14E0727ZvxuYrbWvafFZbdqC1k4p4TOSrTm6Hwfj1y9CKlrEiRMA/d3Ouxz22twh
UDFETXYlIrJUyRO5DyJJWKjvu3+8F6vl1ZKZA/o3aeNhAy803+hCd69M1qxzz1b/YG0AxASqWr5z
y9f7Fd2GCNvBpjThb6eG24nbTtWdCRsJ2rDtvbNI1rXuuektlNTEqOxKagElZsJanR3mj5QbjU4r
QN54Hs53AIi7SS6klxA7PM/L/60uOIW1rDlmx+On6xXM+Xjp6VSRjDVW2J4WooFe/IHfMX7MfF2Z
inFQ2xASZhf0OftKIn8Nv5Dto1/V212lj2zQZIaFwn9a4BQEK0zLXutJqD3T5KIV63LjrTawmqZG
xOVWuTN/zraw1uwnyi3a4u/21JCHaXSRxGC/K0+LS3PlkwG+6VCA4+kidEAfsD8gEFcUAMdIk+s1
uP3bzEHKnysWviQx2MWLF4G9cz85z1/aqc4kk+Fj98rR0HHWrtDSRtuxJiv/X3SyoqUIza8amRnd
leOH1U67IJZmjVrLYWAL7ax3RYUnNXDSN4DHAqfFGGRfzPGZfkC/AZGtR7L89FevU6ABgPDOfQ/F
Ez+Zy4b7VbVULnDiOntuot8MtervlYELihRPPRTjVcsyx2TpurOb7geyT4084Hfg5/HseqMIRuGV
LPIaewayT/9Or5JuQ7eiQxu3oVds6YbMLv6eeVVpH9df/8Y8DLWU1hYgQtZ9hnmDKAUhLbw3fEPb
iYIl6E6NBePX31FACYXeYPwdEkeWwM+wauXiWLyrclTGeDiXD6cdxhv0+vErK21jygJzaQNusXNT
Unjf06wURpbu+RWASe33/lg0pkNsaD3hiOLLZr769YOY5Uvz+SXeFFevYxYmDmZfjuDXhllIkqc4
hAkEjd/9CXRKH+9YVV7xRy7MBn6s3mJsEvCmc8W/Dq1LEIswRWWcfUDHhv+3R7l9oV5bTyAdbg3M
ZFX+i9E1YAiXPHPcQVMSeJ2oKNG12OGHJKy4NUfnxFyvWKCTqiaLbmQo4H6nxOVtcc9NlexSflnO
y5XY80R0jZSQJF7+iFfKxpjl4P3kONGZyHx4Yavewv7Wo/YVOrE//6BBUjc/KEP+4dE107Zm5jCr
50UWN0mR62R6QrKdYtcUkb+ZLKazXfELKGkViMRXjehl1VDIN7DHM4uxZwnDGfDXjM9SQ1oZ/mC5
TM0NGWybdbv7RdjxyE4E7YYWiDUwCXbPlFAZM9qklCy902L/q2BegECZCvL+sLJi4EREh3D0b1rx
veq5tMhokj2QN/fAq8BbyfLbutxL+asXgS10Rnf9cZ0MIyVPEqCS//tkrveB3duDCpVR2Qc8lMFm
4xPMVMgpIzXZYFC2e53q3lsxjw5ClDFuetYcJuKIlPNCU1jdYHutfre7f+yusxDHFvXFyLOAdhA6
KiCl1CU4PsCxMOx//VLljOMge1AMo2Xqs0FUVHggSSm1FyTf+GiqBNWqTkDPWD9i/ZtSHOLZIWbw
vJefTs41qifULahnl2Jb+yTVzrFZHyZ1VzGf1VkXfoedkTp+MoArEpV/YQRcEERJ85YYwNFicNXF
8cdwEu0dpVvcD793VU4jF5dqjtS1t2n3UKL2Nbbom/SMRGaEu+2HjMDEz2beb9sTvuXJZ0kI+HFN
UN6YjlAunlX5C0l3gb4WxilPlx7wXh/HOoGIml32G3SrYWktx0ZHwT96LHZVLIw7/KxViqMxdRaH
D9rYf9nAG49L+gAHoPCKcWxPP5f8rmeQ2nkbMLCMcr72wRvWMivKLbs9vxoNTxSznAqccen15WfI
ENkrESEOFEbfzc7t/wimjgWn6XiF9Nnszsn1vYE4dXON9Bj7KMBVbQ37Nh8eDi+SOImpvEVV/CIs
4r9EF4qfLDxlbaywMeRlZ+RqhCJDkxwnlQGzaTxRy4JWHrIyqsJoDQdYw678SXFEKIn7dcKO0+os
zNUvhxmqafUQWUD0vTfCJr4iOUipz5AnlieLJvBkunE9T+xIiycZGB67/ad9McPSujUwD7xO4vlE
sDNdFJ8DZTsjF7VGI58i4UXOe7r/V1hEXq5o5PPWoz1C8GiL1VE+92GdevDzRGkBfhuybniNmz4s
lP9DH85Es7lC65MEQBMMLsTWKdUnq1K1ng3e+rFGlABBh/9cnhrsqiCFsLErn2L+VtdqPpvr+AmI
FJACS9QP9GhPDef7MNJPGQWHda9KTxBGOy8L90hd9qmEvo+5LJ0eVfkSxpEDEs3Ncu5Tx8icx0kU
3zfqi6pHJmcYeRcVm9laFpbxfNqpB0CtZ1HHlto518m6SvZVvUoarQckQXUZZr9/Tfwsh5yzzPlx
Q7z5TqyLbvpQ0FMDcsf11v1JKrIiGl4HrZFvnR7Jtfvqg3gBbXsOaPGH5YenjrRADbsb9bES17lL
vU/kST9d/kQ1dManXFVB1rQp6Gbp8qx1je76WC0b0qXELaA28RAAHENR83tD8uYjjBHa3rGolGwf
Edr8WkMsj9UqitNHHVFlLIj3MbFUcVSCq2sBbB+mmSc2eVOlJOhN+W/lK45dWb/CNXXhPWwWJPFE
FNIB4e2oUQsgi0RTzB0pmcGLO94pUGS3DlFOSpKRdECmUfUhRvxRFQVTg7onUWVzmdFJbxWJ2llP
GIsWKrbyeevXx/YOMuKVbb+U4EwTK8RjFGS33CW+QMD45NXrVy3j+Bn285HJ+XHrbB7YYjJfBlx0
Iso2mPI12Z/1IzQhfQ7VIeL6BeAzO6PXHeLOQcLObfSrGvYzZR1LD8NsyimSU9QyE0HwtYQnrKbD
r7hrItlS+bII5M6bXyzwMNmMUKUx6+wYRlR47KhuFMrNJGSt+GjGKCc5Bu4ADk5v1Js5zl3EmXKj
Qq9jTBNbCgHMY/qfDizkxDH1WhqtWR91s7X6gcp2R31jEss+7nfEizG+0FmRpSM/j5ZmhQfzwO+Q
0MMkzwtv6LXG3jCM+8KTjd8zHnqXOIEWJRTcPLaHf9axOIfBijWPlppknAPaoPZzuk0KPHaULroG
ar4ze7uJMKhGA5DwO4p5RjuGU8CVdsIuzIcGYx4rxo36kwRLXKJ2dSyVYisIiiR6yCgUfdGrPagK
1qnHBDKpKIkjB1aEAQDP+BwCDkdxn0QzvcSb/IzZ/IF7SAr3BMPcE21ehFZJI0h83lXoYOJzc0c/
9aCeSYKa7txjb72PxttbM0A1TPGGXhQOPMLUfPdCMAp7VcdJ/7RwE7zmUVU+16XseQ752uI14KZF
DdNeagp9vNVEvM9fC3x+3aHW0wGSXoYiHopO8tTYiwz01A73Oa+Qy6XDPc0seZZ7BM4XewuOQGAf
wE3rALp7lLmXuu/4rOHKvxzx6SuHW75/XmfbCnjtGGE9GS9ro9LIIzaXLZjymw0zgy4kFW9l/k98
yDPCiuWAxCmWL13OeXDFKic9a9tpE2llJSn34cXaE5XdHODTENMbvgHVDHCe3gz1MZDmECx6AVpa
Yq3AR9/j0DOmf2cDwZrEPCkHhlwhYx/SzBrSDgAuJmKhVSMcRmH8EN6XJ+eBO3nXsKY80Id2Lv4g
vigGLYRNjf44nKAltxVswemC556GJuvzszYjxG6AtDQBI7uCT5BShdwFZJ61YMMUktH68ucHFIK4
s4HOBcDuX8I7omwyim1BwoecwizJ2ZUV9T5sZqdWKK81/iDB9OZgqIU4rEQuRyZUSEJFprijBeSM
qvqhEqkAiPiGpT7PeDyTc4+JWPt8LOgHzphk47TCzq5KEmazJQa4B6NSQMVm8dRp5O6bcNIEt6DI
yW8aQ9I7YNcjdsn+W/WbNFGZw5vkHvICACnWURhj0liZv6C7wqJlS396DiK1toN9w8ExijoDNvsE
X+TJmM7IiPeGd30EOVwmpxFSjnBBBH79LlAqTTLXUhVrwOtV0unuJaSKWqf2H25BzbW0NPTf/uFY
S3NndSUWpdFzmt0WfrE7qMvLnfRuKUZ3PFyc7oxRHhHjkGSNu1nSSzzzdbO4Lro57JZGjT4M9l59
O3JBGM55HoYSMRYRyFKx/Dq4IyPesk8ocg+ebM80wT4fhOFj9MjXEAOkKaoWE7ZqUUJlAdf2tkim
Pq6lJagBd+v51Q35gTdSh4502NO30+Naw6Z3FfwMp8mrIhA6ETM2j2XQtQUAlqlhFIVpK8b77lb5
SOQwxanYq6gZ8LdyKl5QJRzw5R3herl0yzWBBo6HBaZd1rv7GSWiazfgf4bg4mgRW4Lt5WiBtYFz
aQdRZRt26vo0Omb7ON3wq9wKxYXLVdrhEk5m7kpGEAJejGF+vpA4Z9B6UQazrl6CzEgMMZt0Rq6x
UXcSxUf1KZcjDX3r/g7RLlYas/UcOJw0S3SdjVGYUnnZ0xO2t53K051PpvDVDSTfXTYH0TRBL+4u
nE8KoqVjwCvwmJDhgRAf9vEJhrIjG50l/5+gyg/GU1zG/80mNYkUTOAZzFsAmQW0H+aFZOPvfSeW
LMOJwi+A+U7hOun19v3sD6fJZPBLxZG5x7xvmnshb8cEqDlzBxtiCAZBA0mb6cfgv7B9C9tfufbT
rN1Vfy3cP5BD99DIbLDUOmEPV6uTtCFVTl2RyDAxXUGZKTIFJsIqqlYQR5m0sPiI7eK0OP9Iw2G9
rENMSabP+bY/kjh2J4NZ7N64oG1A+KzLRKN1vN3sfiV8sOe44aduhAUY8FWhc4hTGj0Jm71a5+QX
cyfmw9KN9t0racqZraRSoug2Y6QWnSeJfffR1uXX6OxEBOtGc6Fn+pF821lwVi9XVa7BC0oyX37K
oLjuP9lSgfpIWaRT2cGy+AXEk6HSZNfRsta60MIoMDBaLPR966ed/52rWI7hvpQRZC9k9AkhPEs6
7u8AGQKv8nPcvKbTus1T1jVIYvsjgOLI+527QAkJSRZhrq6aIoDZASc1bVZFnCBJf5i4O9joBA1G
VLK3oFV2LplrPCyL18mfe3+/PjbLGkpYBSAsAnm0HIhkgO/HHW2eu5V802kTWRDTtwZaY9nRleDy
e//NTBnc7R1QDXRHu1BkA/eUVnzN/HnBfMl+cyy8ls2WB9vv6IC0yzkOrd9ekq5W7nKhWfT3zNox
sXejfTSFa1Biw3GuATcvFpfFOrLy62tt+D/hSID3kGAfZoRQ6zYunlDSJ55dn22FHRYurPZCwKKz
LqjFViGp0Wr8bBaNKZXnZHxcs9rpl+lBAPXuMDbzSnsdZqG09JzQJHwRWlN9JQpoJRKdtHfGiIkp
4OzGaxHViE0B63fgs7UGvXSG8JkuqD1rnOTvuS8pAZYM/H/kKivQiBLDuCsdtSIQzf0CTwJq6y1Q
JlTk8umvjJcim1mBeL06HoFg0vxvKq4T2gCCEd9D1UyjEsBBTAiVzmgI2OuE2FrNX45gNo2qjTC7
OWSG9L8YEdAfFT3Vp6/tzHOyXbcO69dqs5mbdW2ASLEt3BsxGy7UGBCPvqAxlmgC5OLZBuIoqSpf
nOKHDmvOlRfXZ8VNjwNlk12ZOMEJhWKy2v8RW9Zu3fUXherwMsRzhPbih5T6rj6tpRCtBNd8B8qU
ucwQnFMMznf0w6NAo4ffk+BBuJiIDAtdC5sLovPSVG05Lwy2oLhLJ6EV2rqOdiYdRtrZ8Cvd74X/
aF/J5Ejlwwzzk/JYNlvnLoTKdRitAxC5y7KaNyjMP0UtHaZyDrmgh2vHxTPdkawDsBec65yK8+XZ
vZK9xqonECfoqP/KAEKxIsRktmsij2Z/Cqz0LjfzHYdpsXDkTyc0OyD+ne9aBbR0o9xuIb36VFyJ
GdRRV2/KUC0XCdDE1vl8GokNffKev7HiJrg9kw0mXFd6MRHCdN6zvHxWlFCLN2Zb1wUPvm6NagOK
NDN/h1OP3nTw7xdKnuj2GCIhhhHwRVLSofA8kSx1Rqbej4L2LefsUsvHBqCuzHyplCphTSTyfiIo
v0OHw8N3whN5JJJdMR+Kfgh04khkT2ZnRVYIK0+8oXqP3wN9kJ1ZBl/8eeKPFTtcIcIFJSnr/yB8
EqZz+GvGXY/xqjsMuG1pec5bIE5ctkuhwxZo9aFkWx/2LdrbujcXEtC9hrbWMuK5A/B1EWmxcbxG
IBNLjP3Ukez88cgoV0vSPisMu7FUVCO4SaL8TTqC4QZ/oD95N+p99h+4M+gO+AFfr2pPBPE9tpYM
kN7hYuRy2HLbCVUd6GgBMjwmi3CUixHZJ9+BnVtgt3+3zW5S/FpZGiczoGavZn1lx6ogQjZs3GQo
8yHhSi1CYvRMGSyAZpzIyke28/3H1F/lGeb6wOzKuHpND3RuLSIaj7G+T9bkKeTDxngXW+l3EQT3
Az4xv52G9C59JHdWd9KAgrPftItcxqe9arPl9d10m5vBlIy3MsiKXC9+JIR931/HbeiPZNeJVSuR
fQU5yYOO2U7gZ/oAGf8dLEcDSechMrPwR4ZV7hc6W7v45jSA5kb/uNAj9E4eXuIw2x4QQ0nw/gU3
Z5l11eIdYyKHxxrE23IO4hNPxZpseohQxNnQ0PDFhMIydvRGziYTuikrNuJx9b0c1W92x90u3dGc
FfZ3O7Yyl88L9j3M/X5vVTlWhVJliGOo7nT+CyvhS4DCMrrfqcYnwPodWHbeZjlTi2fBaL0YpBeZ
BlZJD38yoTPLyIjaXrS1/xNtwUjtyt9OHApCVnxkZ47owG0aSqPM+zmPatGyZrznu6UDWe0fviaH
lStmJSd/vT3L1cYTr8Y5QbJvaErk/DZVgLlse0BdJkj0DriWmm49FA+U20s9tDjDByUzFn0GNkf6
A6KyOJy4pD57hhKuWLokA+vABGEhlNba6NKbR0lNMg6z1aVSZPCzBYCq/F0aKUEX78Amd2in+4nV
kxpvH71AOAN6f/z5jtPrRVjyybqE9OFYqMYYhcwX6q9NmqylHHcD+Km7S17Z6Ew6GF+beqyPQuBo
Sbd+qrs6/G3orWOFfN2cdlX71sEokCEkd4v58oXBgLsE3kYQXnx6leAeWYvYOf+BP7PXInill+0H
VsFjEyQ/vNbScTsVGNFqRixY/JlDSa+QlTdLkwXxU7IAfPMmelYBTJGloplzpb8aELjH6/Xhpm0k
ZNi23uJilY3o8+jKm8db3Mjaw4OtcUCM4NCQupCsnjDNV1q6029XyWjPpZ6fgFUG1yOvXjSwcsDj
3wtAOuqfJuR1W+TPxKeD7LufKG6sbFzWC+sVCBLWkfWTr77G6soy8Q73q7pEQDFYfJCUISzcdfH6
NR8ea9xJakuX0/Bbh1dTx27IlbpMtpFri3jNMeTBmEbcNvK0zzofr6cosR/TgtzqAgu9EqswGLco
sBqwx7FJ5JFXzn6lp2j+FulMbrOKC9bSkZfKTNx6UwOCuA3zQB7DKRcPAgxVUXkj0ssedjYN2G1K
+JxPvBNG05swZ47Vk+choLMesAWEsS7L768fDKKjMDhAn21h0fnEPDoKBHutcs8GEA3xM1Olf4cN
O4YCYQ211FgErp/FRgFFaVuIRIWOGvBbis7LxN75vV4jKz1NERI1xrvpMzK2UxukzFIAUc1s8CDu
ZeVwIKtkUBpEiKM+RbcSuwRfZU0BoOnYzYp1LPnBcLaeM/Jg0iskb01nquR8bxtHN6ZIqf/Rm4LH
fPZi6ye7IoIH4RjroMbMRpmpizOmbSkwmuZQp5uirJS+BXY4eHa0n1HKl7h/WQnedMo6N+rGk8o9
dsrQXLLY6w6+d4MrK4w87Ibz9sCiJ1GyVDmUd6ADs3Y1Cl9KjnJOvGJ2ajLBKg5oT0v2kYu0JFaH
DlFnuptxKcDSiR/gHp/TuLP0wxFVduuowwZ8zgN3ZmQnw+tET69nta0zTINt2fbwLsQ2uO9odtgY
Wfc6+Bm3Mu5KUiTSw6Rk+V9XVpT1x9ewauSD6IzMPD94kKFfj/9/y4mpAqUwd7IR8/VPHk3KzCX5
bML4a5unTYLzOWxShVFskH4ZPzWo2u+fD/tPgkxCq2yO9BEV5/aYvecAUk6j4JceP2EC+KPOpVIE
tyOpw05bv4NiXn2CDB0JFfvadBYovJsoy3dC27uofRGoJ5+gpfJi6ACBHgNeIwsVPlGu3dnONiRh
Bx832lqrPnv+J+wFEaOrzpTtf+8caFn8OE0UI4POEzRuLHYn+LnQfZd0RnN757pFK3gBau+R28sU
L79SLZm/lWZ4Sio+svYvF5g6yNiU/jIsbPGiBIg8NLpFdwnL8GBjqgD/34Iidh1zKpk1J3IJ1Oeq
S0OxAJzjdRe27PqaQ9oxEhuTl0rzBRWvSndESnS88caalqZQrAhBhl+tfzQZThjxyNGTcpk+RXxv
qxC7mSDN5eMS3g9S2tUGQlxAO12eCU7lFKPLSg/gV4AatxxN2rnl2XoBV60Oy6lh945K+aaL+/0j
OZ7d8E9wyCymx9VCLh+8pWqPvVwWTLJtU52CqIFvfwnw6UcQ5i5QarOMp97J8bVsomLl+77Zjj6b
c9UeZ35VwAoSuAwJKKwLB/+UCo4aLSzsYke+kE7UP3PN4cIITQHOvk8YOBubyb/eTLaQ0xYqyHDL
cbC49j5SsB40dcb/beoTn6VNk/blpFZWAEB7UFxhqRUHeOSttOOv1sS5zasj+FXsrBOWh7tgcUd8
lTm7hOsx6W8+NADqBK+7H7lwJQWaOPracEctB7MzKbtABQHzYjxPcIZGPgPf7v/lgKlmPvkvL3lw
qcN4B827brAARTjzwBeJAdyYZZfe6YAzp1YMAGcmrLSaCId+gZnghgwbnd23Sp3HV/h6c0+iqtqs
KX6TE1uzl5RGKIsrtNUS4dvQmXUwXyZa6pi4dbxZuNUWi3vZxI0ZTCXofRlr2z7ePg6dKfXV0/Ei
raWQUVdXenctwYVUUkZADbU079tRs4ToPHbH3Oau4hAq31m/t0K3oWI7qDoAuz/vtbgmBtktKpRN
Pj8Z5oOh8vL7aW1xP8258RJOWUS76Kq3c9xChktiDtN4/8yIulP7WInYHa2UXRy8ZDwc8cYI7pVb
hELuZBM2wQ+MGzy9TTQY/DukpVwHzhgwv8Q2yj2nrJ7Zw8zRvkj2FruGPFnyR1Kx3T/4EzUMT8qi
w9Gh1btuUAnL6Mzyg0G5I5UaY80Jc3Hx355VAfu2h4l5U5doaotT8s7ot31oU8DnLq7TfUYSbsgf
jDlzKz1Tji1sP1kS0C8MNtiimTY4910xE3O1K9W41vRg6hXCstbC+OZYON6R2O+5NIoCPlh0grwa
jnZqqPVIjayciGyHCo3NMjK23wmvvjVLu5wBAtF/hK1QeKO13y+iFPghMZBd771ntLb7R9N/Kdmk
GzkCWWRfl85eRk+kO7NCA9sX02zlSuyMoDkeaQSajXbXSs/ZdN/VR6hiy+sQk4PIFPqzsRDKe4Da
7pn0OOg9OWhvJcA/d5OtRAyNCpum7ZrOiXeVv+SmlPySoX0+1vApShg0crtddPtNFCRy876rtN+P
hcmAndH7cu4jA1Jffoa9o+eJbL0dX3MXBcZx6JoDV+s7hdbTrscgzKl0rgSyj+CRTsBznczbDRNH
TjnnbOZSzUAr08JYFBG3m4l50uctvF4jURQySaMC/vF6zweXr5HJwoQZxfSrktIov4Uw6aLjRdFl
4Kr7kTv5etnq04KxfG3dNW34dXGDhYMsdzVMHlHQkqLp7iUpptAMl4PeUZ9t/u2+C7MAawGvWT4f
s4X7+SQRKYtmOvW97k43UbwJAt5xxRk+O+bknvhreIjjF+V+md3dVTal2uKOlGMm5NTi86cKzph7
n6uuoQ4WhuTLyVGhTL2Jb3ohiIBEPusf8xXz6KAHuGvQUafrrEiEICBwswyd3W8Eo6t9FcgVZuiw
jm2UV56x2K6AY13D0tdb2BqsrBcDjYocshocwKhP/4F54BOyiuExVty59j21/U7fF/1fJa5ExQgZ
4lv5Gouw8jmOllloWaq50KXxQSIj1CEcVX4VZjlb6UVLgX1RNW0ZZErFAyf4ChQC88I4rZtqBYxt
M15Yq5z0m83JF6v2RtcK/m9DykJL0Sk9cWBcYZauO7YjFmOGzJeiFidXt4dP7yNsNLj5jQu+5Bvp
q1/0hQgNu7bpgGmeBXs6zcpRw54ybAJvR37THcE65mjbUUmV3B1Suf3sOYLMAM3wrZhVZAVX0p2L
M8AL+5d0syzmVbdt5ENIoBmTvBzGv1Z70efkQKRKMoIbXjDL9qL+yP/jfrKswwTwnolS+Zv5gcrB
l/zU27uDB6ystiZ1yxfG6nvd/yeCnwoabL4bWO/JnvDcwgrGJ6/lcEiAHf11iMcX8tlQmmBGFDle
IYbmf+R/8Lg0Jtk5gyu5V1YQOCrX2RY/TJV3Qt7g1BR4oyx+nVZaXqDig2X6E5eQtiPeUg+xLApX
/veleUV1XDO42CjPqzfOoa9BAi4HNHe7Yoxy57pQKWage4KI2aW1P6o28qYqXvDgrFzJjXo4J6mO
fvuFF+JefTNujcLbukWnFCTXL2z9gJu+R2ykhwGcqY2SiMdL0U27Ou9XhVVrtI9ofKRNaN9tborn
GNocuP4OQu7IEZdcsdkSbEqi32Kwx2gMahV5PDnfMVOgtddc4r2W81Sttbm+F1qc4FxYp5sTxYLz
JWqfwRDF0b4fBHN1R2gjQLn0hSrAlc3BgVc/IMRcfFfiH10gni4HVXO9DBactLNMZJeu3Q0VLA9R
SymP/YsAdtWeANbchJu1uUX5B6OJy7x9nd9soCjexk4Szq4oRgt7RBXtwrRKXokJmDKnrZpOKkW1
lXLjg1J1MiDq9GWdg1+qesqNLTx3z/sa809I0PZtqLFxig0ScSywfDBx7Zuz2MbK6/d0LPdXEcn+
aF4x38RrgIS8gyDAIynMbN5Mw30JBUxhX4oY9GhdhJzS7+izf+gvfkTLOFqxC+fO7LMJ7r5HrkgE
Q3RxyXnf7vjdQIYYcqjILdGC25pey6x2uyGHxXLPrUtkbifeSAFpBBvaab5fswPIYZrgVXGky4Hn
NmRxTGLXAKGzqamINgEaJU2lYksy1Zy7LoNd2WAFx1Sdd79kQeGJqLK/hCtjueITmnGAmmeqUqFT
YHgRXh9lFihW4REdolgN69sUCzIuJAoAj9BotaY9G7aEqW9ly06BeamtvaOhjB9oD07JVP+PZ1Ey
1eqig2oE+A2GlreaIdH1x2HTfnQnpQxJfYCDbSjldABfoqrs8ZCGm5XjxHnZcVos0JNXaQHXN7NE
xErXaUghm3eTrPrnGF5G+YYNTIahmNTEIV/w+4axcXJW3v4CMrkaY0dpcLJWssu6sRfMovQ4rnFv
s+DW7f13BjqUl8kNbtrlojxP7545LMiL4kqVgqCXGykLQN+trMoIn6oCYqTXQI7vcq4YAhOvvmXH
Qmt6Aa/PUXxOSWyqgDRWelohzk06rXnE7ddJbvrQz7UV1kwMRbvBiz3ot0efLBnEGfBwutK9CkvU
/TUZ8Wn0dLCEs6y7ovf1ewmX+hcauSXHDsYq5wEkMVY3OVATDMOA2K+/vK78JvpPG9m0C2rY3N/P
Jn9s8wjvOprmgXVxpyJMj6NpQOzSY8A7EPgRUBAMNDL1zrt7nKIi+QuqeBhYP3JWvZ+pAQoVWYAP
SwOVROFj/gpcWgYaYgmXzsA8GNdyyNnJ+oM7+1zlJLOrLw10qMT6all4q2Dcs7zeNrXCN9BCVgeE
ELx2aTFkn6Kn5bAr6MA7EzIiaTPDULiXcntywBNFeKKPNITPyS3ImUW7k0481lvuGdTFvHs9W+q0
6dori6lf2Oe631NL0WuYW1U6NqHvoCVxAh3Uo9iUHpGyzcHYMD/nTui5Zhyw9otEr94WdW3uYuLG
2yOp/vDsM486Bj5s7FYo2q62/LtvT5AXhwIjqrZd27MTpHd+1phEeWjan+ZZ7RAOUcxnJRo9VxoX
JQrMcr6ydBu3qytgFv4lHwXk3nn5s6SH80MkmdI2DjJgpTOjCIpCHGCz5xPXIwrjdSTz6PJefop9
iO2JG14tkPwfvF6vwxqV50AyP/dAPTVdofrugzMb9a4MAX5sdlikkEAJx6PwHRRVvXNBj8GI3q5Y
VjWPhJWAJP4IJSEPiA41twnROzQdMI9rPuGhpvgyTV5PdDOVPsy5Urvbd2THK9qU+NnHNb0VY+kP
lImmke2kzxRtN+mE3qCQStl1J1M77KSLHMrnOni7+O/yk7aNuHtuHN4j5iNe8T3R/3/xOkhB+h5j
sxTakRHPOT/+p1mQsUADdPhjgdJ+SVbkLv2s4qMuVxS3iDV05E87KrlvNfQVcgUJJ1mKPdutpJf6
ODyBqeSAKs01QkZtTurA7k25+tQZNolgYU5evoBKPUJJnKsjENYWstn0zKmVFyo3EcdkkaBkS2e6
czGrx5m9rvfO2nWf89jHZ3ib4wzq72MNxLs+huwqkutb2FudKMX8Wtn3LfgDH+A87sE7ky+zqKrI
bd5oXhjmfZILRFfVpwKpVTuqHVXRceTP3MUHz2YIIHPWOPcNaCwYyqCXH8B/3YBVSOnac48sli30
5CLJYWpR22bHQzPP/BWV2jbgHgiClHdLNJadx/ThGeEtTx4OHEha0u5FLX1YFUlG85aWEPuyCHU5
3kogi9oKZNr489OZNyDCCpn+uL4ssjC/y/xeASUTbzoNKz+Cgfmgd6ZLOuEWalsqt2RAwRXjiOEK
pH/VAoNWzcZ4p47SHHO+YLkpO2nHnhWEuy/ZhdqpDLIV0fAWeAf5eHYpXlXUwa+FB9W1tTtxCGNa
KgftWC/8h2OV+A09wehjNvkhPfPEXAdXM1NSyJbb+CAjwdOyAxDoh5V2EqBvb8GxYVhHIjW/iL8o
jQ0fV1Gpqvq+xMiw6gs7lRTleDJFPdWrkSjllp6jWA7AOioZwzLys6/OJb/QX914TMIjkPAZy3qt
4q4LG2UZF8batMqbghw/AJflnFXNgFmCNqK7WGUNFT8oZnIE7CPFr/aJg6kloDVm3zSYGtA7CjCO
2ri9kzSJUGhFuDMZSM8mWbQ78Y907tXZv9oOEfP+NdqsLJmmvQ+TpbbYTycxrqwaL4O+EFMFhLv/
lnmwGOK8seZygnE+SA8D4sqpEwg6qGZNkmtw2lbYRnFfm/KKvAYQFth13W6+y3LDwriwIBX/Q5QW
PxM2kVO1VXr1GKJnhpRHPDiQYO/aEUqpzuWNhX4qa2dYPZkq5daWkE8ZpbYKFIgITJ4MGVrYCOTW
zQmpWUN//h69A4GDf532Gu4Hs6qrOCH2T8NNJNXkNJGgo43kFkXJjS5V82GhCPMTIZI7YJgMtGdk
DLwLbNcooAdXTI+D19QEuJkPRlFkKP8A/kKZ6qB73j08gbGHGwGRLD+ywQdodr1xQ+1Nb42WcbQE
LlwHITDoNRsLnMxXzAxjn10da0LuLOUbOpFmXIvGyig4xQeu7zLdfeb3HOv+hHbq8y2qYE/+7FMB
ji2QypB1COVFTQ53j+e94zgK9Qg8u83+UTOYDBh4SwrRbpD8u24ejLfOXSCgknD/Nal/MXpg4vzW
Pg85bfsfy+Bc8kOFaFXqRlgSOeyZB2pt5A60WQ0hSnhHvxpKBXJV0x+zC+rc9ZMIucPYlPLlCPXN
YKZ7IAsItvvHQdf9kSMPQTm167XsNUsXofHVfwf83ibBDzl6FcQ5IN4Kwj673lC2jg3mbqpK2f03
//PSs9gedMrCc39Qvxa4126uKROpy279TzlPs4WVv8J7aQ9ZmXJz0TAab6w9xiqVn2VKvARHz4yR
SubCdNSdlu9juCcoFGxBb/RY4vik+XYYGSxRoRtSmms6DoXnKStNK0S9SSS/HAYxs1ErYgsIsu6r
p2tn3CQMue8SFq7AFWKP4F3gxOIOUtJ8cccsOe9+c9YSvrpXLtWZ+cQd2HAu6Es3sqOju+uqSgm5
LRe0xi7iffYgH4FS/FW0Nuad7IIAjGSJzkBFEHbadLlBNPxgiVwUcgJDIESmPZolPRq2Lua3m+l/
DYedvUc1/LLiFWeAsajr2cM35chOPqPllP0zoXxTz6e4K/jtLXT6VeGLfSA2OgS0sM5sP9DgcNxp
KrxOTsXRI3YQDBlxMhkNL0FCZRnrHZPLA6He8VXAUnZTtwXzlVCYp/6ygs6l4q6ECZ/YX6fdC0Jl
aEIlXV86t0P3iIa7j9IZLgUbesDScmwxse9Mps1H3PyMNkwegtBAdtjDwV5ka59l6RG8ossykVVC
iVT6J1vfrQkouQtCNcFHLnNp1qbHx0RpnbC1llx/hwzw5LwEmuEQ8gWm5rUeBstlXDKdqmMSPTyI
Jqb2O9SqNiCfXgixDvJZPQGY6nTHwSf5MqPiw3Ov+swokLbylOoUxf8oYqSC2KbSDGU0F03QC3PG
i9KFyLfNhKp7Wf4sDup2ZElXUFs90BcJOlMMs7d7FlyN00OoPalWD8lwNsb2cydgUI55X2BH4/tl
9sc5HduaoMETCgWR9MbAGkjsY1zDsZRRhd7aCDCkdb7tokN8NOk5w+c5VLRm4Aa2g344TewwiobA
a3ijws3FzUYr1JLJGOkLZLrIKVe5kpZ0Ytm9OyHy+LS/gBIaJxcO2HbdH9k4J4vp8DStrMVCHFUy
MBiajyMQcBhiP8Y+zN2O90Iwx+41kp4B6Zxr2VJQamSq4LOaYBO171izCu0pFdg44NxbJS9DxrMl
K+cKbxrxQ6Jux6oBRDsBkR1v+XUltAO1oVjWk+BPRAFtn2WcXKMXz0T+bUqn1OZ9Aytzqe6kqug+
wZ3WQRrTCk8gopK4aWO7V3/BJlZ0qbcrK+c2AV/YJUTGqfILqn6N3G0xbF9EivFF3M2NKAe7CKWL
ed2ACmFxyXx+T1CrZnPqW4/hg8q9rcHm2RQ3ZTEYN2HDtJLPh3irPg1aterfAOx/ljo9HWZ7Nc5t
RfsGC4oAT8UW5Gr+XBsXXgtaqeZOEKplLO7Uh/uGmc3Grptu/j1C4WccXqHSK4RircYIn9YyxNpA
1rKChMHFMK9/Gk4WBu1Gpit3UKQLsNgSKO999Xe7wS52hDpXSh3mQYQNDBCcSZgfQX+K/rnVgn+f
MRxOe6dyqpt32Q/Ol8KIwSk2Ze+tGJVtV24v4BzsmxswLqqD4eGsnOQ8IJHPx5xIa4xhVKc/BJcx
oAV/2VAVx56UEUocPIelrKnD6f21CxiGi6uh9M52BroHwRXxgyO7BAWXfv0wuEaOrG8uDt+H1szG
4PUMA/h+9Jh+jIFnEk1mNsPPaQYrVlGMJuY+8u/XOfXJUjTH+P9d56ecD8F0MeLqwUjjHe98RYkr
hSiwA3jnf7qVm/dPGJDOMzNgG5qcgE60w/8uNFstKvdZTa/LXapHjbt8VSVfA+JBSFB+qosynHuu
qMz0+kwrJFIdTXlwKnjWz/1HW9//JOppXgDIGNsWVMKXS1xU+G82H1ISnAGTVk/XJ/cwbhtzeqny
oAEsiI6fmnwj9NPQjh5SBJHlQuS5lpY/ikdLTOdSyFa/kbkENgIFC+DI0C1V8gTxXWzMmX5ZQBX0
8h1kkqRHfBdgUwJolys0tTtCBqAajM4KOIeJabjv2gBkfDRrZTg8SuTMFG5YQtwbOzH6eqb5h+cx
i4tl/yGIs9QhERJGDFO3IDVvc6gv+ZdpYBm2UmfF11MO9re2EaJ8Td/fPCGg4OgvBE52bRTEGPps
BMYKoUxbsd9viIL9MIvyZxdYIgedpx9/DY30Xa7Aq07NmVA/30qSLYgKx/2OhXuHbiN1SIBzH0Oj
8hnUxBKB2WD112Yj7n4ywYjK2njfU7Oki2sILdHve/T3zXAKQZl+rhNvnOEWgnsEp7ur8GINKFn4
o95xwImnUB9eqLsgG8D63s85F013lDQyvWWgEtHJL8wG0Y0MReZFlAsPAGFbfrcbf5xlnxXsd37f
auX5m8V1gdwxYg5yo/yh+a6MF1X47guRCMaldIzw40ZYFMcCNlw+Mc7f0lKDe+f9hE/urSVaS46g
ppEy63/qeTlaPlWYIQi8TLm9hy1MJ7BQFXndtWcBJ1jWtgkLyg7u1eC2xxnjd1ERCw9zxdM3JEvS
1IhoI2tCk3nqDHRJ8cDDbSYv4Jh9sGXA0cSMJ/a+zAgxSm3VJXV2SsQerN0xqn1HEHSojecPnB4j
FQTiZMydWcZAJ5wUJHrDT7jVQF+BE9h6Y1GRyB9SFfpnDgk4fqDv79Y+1ldjkNP1Va4x1QB0Bks9
dOSjOYftHwR4/sMCEOGLReIPAJdtEM6MwpcGKekLRrJNGWlHtuRxAj5w1a/t/Ri63YUmMH2WjtVi
YiRL47cAyzaI0Wiv8DCOQxHMtCd+bYOgIRi+2k7oHgqberuomNWJ8hESzaGFLNEMRRcG9RJ/Z9Gv
HYWcFFpxEbiZYBaDWnINRePD7dsaMB4UA/lRNxIUazdhDWvIkY4AefgeSQv8QLJFu4ntagSh7GRH
W8TFUoCBH8aINmyfXt1zXWbtU6uTKg9cQ/WnSSJw9wxXGQA4wv8PfZcyKl8IxpHvW+xFrhn+n7y/
bDVMxE9OiwIHP6PJfAts3E+tqKPoilAPU+f3lLNolOvWquxIQKxuvCgmZeb1eP7kxxB05vgWEpty
LWV2hChZM4KrlJpNUSKUivxFvmeJCvcPrM1HGzRsN9goFu9iopwrDyk8Du72RhxTGKZIYh0mBDx+
OvOwmQzzEP7bwRcgobevfsVmCm00sPxlmuWMoJfrVnJ+dNYia25hLPkQHX5laI1wqNEdCHmlqODj
iVkzY0qXwWyg4bjOwrn5pw6IbijxC9BNVGBowN46ysbVHT7E5sID71JPxj+XrNVLKTPP4QtlHp7Q
lmtMwcEiGeUbDbxxYfOF7ogSOYFYk4wmyrGTm7Vxm2IBB3wKWnFBH0TIkIkhMYkNLWZ+hv+XZW+g
CSbjxIBCFWX5oA6G64DvM3YLEGvDroM1mhCyHZ4VlkcBu98PpHNYhyQxHaU8T5Y8PtQAtvrqkHKq
Fy0B6MkbK61jvTsgEZasiq5TBrwyj0yCR4zpih6ebrLW/zRBoS6Bk2NSC0NdSEdm67nwUvuaQq6T
wKNQfhVC7D/esYDMFdbjQEdqOhmoFxNe8EYylDVeZ3Fk/FK++a0Pf3ss3jTn0V8J5xkUqhJnCtHG
taZ4WFRQ8RX/gXrhdYXu+LVefuykidRV3aiaG0kaMieT8yAVNyF53cHzG27qckJkSn2M7WQd0kAd
S4jyT00t+4VmDyL5+dJdfgy8gnj3jER6kyv3fJoWcOMf9Ps/o2f4/R0owZGBieUiZsfxRYyuxN9M
6iJjepEKwPwSSiyml9UKZuN6KxX+ElD8BnH1TVcO6q13WiAwGeWcmjBvAjNXClQRX/owrrOfThph
pekiLJCpVBrLqyXE1+Oso7n6PN5cgHDRPbbBwk+HOR/m6UfrirBt/Nikur4TnaNNu0SFUr6HejaK
K5WZy6QDPVfafz1klxtTDM6RWv4ACCsqNaNe40bMNzVXUVnrtG+3S0r3oyrDMHLvhaclumsJvQhd
IAKdgB67c0WQhw72aEfoVfJ/7iTCOsO3k1AL1FDyGQJwwwmyrpgc4w5em1GU8f0d1/O0fNpSG9qq
IE8gJTCo/GvLrOMHxr1ePKgCPqY8i827S4LFrcFb9Kk8pL+A9uJ8sBnKc5cYbukYIcGU1efm8dGU
AurG1ciLF7flmq9LGNvIaiX7NUX1PgofNTyw4GhSsw2Fc6RQxXoRxHjciygoN8avb9dHcGuDQutB
6PtdkQWBWgAvplQlnOKeQshEmSqNo4uX2A0tNXvGy0Ov7vgIyNxpwevWztnYllpElZ3WhkOBnTP+
Mk3AuZBpwCIwSNkaXqr0MqUkqBrSnXb8RtfRbVsmKB7PK5Xl2iRWJIych0VPfEjXnnmyOV55FZk0
lC4XOiCyv6EUD8FzzwDKUpBnABGV6cCxQEZxIJOaX2fCruRGFCKvRtO7c4C9Vd4aZB0dT4eAbrs4
3jzxgF5zXR+a6Q5j/etWsTd3BKQCZ3iC+NBS6YAURcStos2Nv87gUECVyOZOBwNeoU3fsKFBmqMR
Fi+9wp5VjxIKOub3HFkzC82hiVwOsTRVcBAuu7a/AAnhcpyuDgCwUtI/NHtFM/weJplxsetGRUW/
YL0x3DrnnEm+nHropgR2HnxfKnA82SdWzNi1hSf7jL9ATlpC9mE3ma9nWzU1X9CxBc/+th6xILlk
RzpjO/uHM9U7sTwGQg7dixDH9VR2p5+RNnSpFmTqYsAWhwhbYkCSednYe1rFGcgyMf7KdvEYSNDy
d89WLPbTMemusTwmvw4g7DOgKHRyRy89fl0mv0yoqrvPeDzBl646NW4xNjAbY1pYxJiiLJP6BXWh
bP0JCc7Ia9BB1Ta4GIerj89xeKQow65VJNkZake26mkFOkf4loAPtoO1u7kHw8DKc1Ye/GK0cYaJ
E8jdtdUBVpcA8fnV8khkMStJir+NhGWRwOTwk8wloLUefGUGkKLEfQbE9OI3CjFrmQyE3mSU7HFw
g/a6m9+NCTIjiopQd72itZ2D0dkf/pePdSSXO2h1LQ11gEdpu4koyVpEuX7FzxehwB+RDiB+p4kV
fgkBnel0IJZB/nakNPC2CeNmezj8laKPzEiL7KQ1mLK/SLohu0LpqFHBwC6PerI5xV9ryAj/WJ9Z
2xNMDBvz4jxkaVHFXxC42COGnpHCdHBpZmH1bsQWwUlkAEUovOPQ3hYaYv5aO1Cjj8BFAb6tl4qn
ebBDqW5xENpk8oKQgygg+Ir82EpPPhtHh21pWy5ZS7hVCwU8s/ntDb4nohtiD0K95+aF9okN9pCm
0dDTjeKF2Dh7bhfqAMjuZ3UAA4Kpxlq2YzkeJ4UnPPZLF7LvlRdaNiQitIo+KjZyqZfVRGCmUagA
y73srqk718P9D06RsU3jINwywSSOIcZ0JzfqTLH3Q/q3/Tul6++IhTf/LRhEbAKE9RUESTHIf5xA
hu8kKBS2vwbLe7BPM7iTSKZuJFcOJDTW2O4BQvmQQsS77BNAUtH0tySo/4xwcHi+mHjAUu6oANng
3OgdeFrRLJJsYr3c/4YpNci/em186UmeDxht+VwpGoajbvjFcRnJNktcA/WjrCT6UqAwwcyd5HwY
M2/Im6PIa0hLSxKQ1sHV3SL0+dWRfc1L+nG1mmSGu84vLdSdCAXeS4Eez0982jhAEhylIfNO1lcW
i/oFDaxZizwNDffEeDb2Nnw1IULQqDi4WI8xMGOtuMkdVG3mOWPy3QhhvKJJ+/Njc+mIQJl8mvYL
O4OOhsdgwxkUtfyyEbyQeuny0D7Kq6oURM+zVgYRGZXUN0ZFe8Cpnb8nVn8gnZR8HCYAVV1tqkp7
Xi/3mijkQONSfA/6r+obOcBGjj1kguoUje3RoNRJYvplSz7Lvsv+mahXD16s0rHylbxoHxji9Zhj
xmQ3jtzDDjeX8W+6fmOqmBBY8HwoFWH35ohYDQ4lCQ2JHmlybi7vIrXvMg62ET/ZriCvLYOs15VQ
UkgbQYmWTfo8N7XpcZwlX3rMohKS0w+jUG6tajhUcQCT0JR5zI5ITKO7JKZ4AoSKb00Dv9oZ3gI6
1xpnElNgWwEqAQPAxpeeRwzn80IaxmtDqPuOElQjWfrei9h5E0zaDxHgGvL+dSKkeRIre1uPAljj
BYcCNcr2k0Zyr6lpC5PtlyyqNe+5yeykCAlozN92rB/hI1XUZKMKcFQyjXTM5XhBhRLudCSGboES
IVLeiC4xBEZf5Rp4tGJcW8opGNl/VE1miVrjgQmlr5fc0pN9ISUU7SF7BsOwAixXo5rvMev5uNq3
eNQSccgZq3n5bIMDce/+TwDPbILNWcdB0d57hehqJlieegDwjuoDUM2837BT7xU2i68CZ9YuYJQ5
5mAGOa4nFKQQCsv8W5E9yukTFGL4ffXSE/e9d5i+SiGm8ylCmw6NxEs2W3gXqIXrY5y4+CrWsD/j
n/BAueiAA8ecNsh+gkt+L81ZV2Qdo27Rb2Wh0mb1DBTWIpTT1WMSKltKDLTaRtgbZ7JBYcR8BYhj
1fQ0NYcSVh0MHT7zCkaSUjZkELZK4UaF6gZCDZ//HNv42RcgrKikjtpo1mfOciOl6uY60PzEpSJl
+0YQ2q4RNR1c676uFeFzFt25EBHUv6lq9XzmksTZlWdZSCZTYECAqY/Wxqny/pXpG11UjB9KT4rW
FmRBKGFxbjsfCJcHo8ABd8cY7vmpb0qnF7RJRlFJCs1BY9rlM5QJuggvDzIRhHV2rWqJ7lCto0xT
ldZ4hjwgvIMM3YGxuEiRaJtlYyXjTHzoh7d4/ZKI1Dm2E9vCW1jf5GKaqAdAV9TWN4Fle68rfML7
/zhJEdpxzPPmNGuoKyonA1pkeVOaoFBAqxJCsmGDHIscYLed6pIpwJr63Xod84DX1tMTYZHKKLSQ
rtincvvhtunR7TwvAtsZoAapGmJonnokVStIwWKFhugjC8xZfwBH51chZLumLDyY9gu0FfGBtFu8
UHuFeDR4z7T7FPoo/ZNXl1lUo9UZLd2n1T2H7kbYs0BmwHuxPiWKUmo6J0b7iF7zZwu9CcgyqNJI
G17TkXjTkNVCsnnl7KPkkD21I+4Eb0+2g8QguYqXyTzKz+iODkoTXePx7SrkUSttDTQ3j8Xn6Ccc
ZKP0r6sNe2n0sqfiD33FetBLcHpLluZ6uDnyzp127/f3jF99zagqDxpw/53MDxrBSCeyDYLEu2q6
7HiT2QxlhA30XZ/oLtT3hCNErWEfXS6TvtvBhbzMSO3W7ilcyFc9AqVNwtEQOrZebn79BszYGtJy
+Dh2xdKxY5mbCFG6p+yyBmQUJqggdzYHj2xV7Z/n3vP6kcogNzs9eAwOItrjAHr3rncl+BcPqaFz
BA179Xd/8+ZRrwdMwIH7/WizVjNuppRxjA/FjhsYeJhp1v/zdMP1JQSzVO9Cof0R0ESBttrRwgJy
p9i76X+kvuAFbJ2vHjXN/OTPvfubeqhTD9E2a1NN6/zhOmpswficELhWD8x+Dyq/bvzNrYdneH+O
EKIFpD2s2tJqQutXKS7b86+TGUAtBdboz1vqUkgiPU55PrzPqztbDqp3C+c6LL6cjmw8DI0DfoNm
4XS29Eqvqvc3ALUttcIRDphWbt8IYgZQ3dAtROK3y1Bpd8/NrpTBy88CZMHuPazrjlripowzZUf2
bCMlI6EDLl/XIHdqDHxGEhqaSMHK2dc2tGvfqlrz8yRuA0ivCBqXgPcriobsKNV+66jJJCUSdMpZ
yzDdVzSVU5zjjrYvIALW0jhhNSt15c2yl0pmThxQE2fzDUBhOeknm/xYAQJZZqesREH+nqo716b7
kmlTqraVYCqPKQPIFWL4wkrJUPdYF8M+rc+jvZCdl2lQTAkaXg3+h6tiIlv3O+oaZs2fdtmbWQ+K
M26Ry12ETOeKQlG36t2031sQiVF++o9qHU+a5RC43b6eayivx0YYvABatHq9rfcUAg4ChzmGVAGb
BSh0NWhz8MmyqwORcIs5PA6PSVZx7Pr0Zrr98ibrBgF6U3EE/plJ0+NXQD3PKYnIbNBb3gDRr4kU
b+WZ+MZfdWxzcU3BrltyglB/tPeSum6/2VThncttLCsPGGD0fYR3Ukqd8BcnNOUXXEF3UDFoxKGI
SaKP/VF8/MOtwXBKE/H+T18Sx+WBkzqtiYGCTGt42/flDkyGdae+m5bVf2BSvrNoOBlJa6M8ueGp
bzHIxNymp9P/iCJKh9g39+pp96q7MOjmVozLW0/xurxMNZjk31fxXFoDTnEEhZgaU31BLwQfIsor
PL+uAlUIWlq5mOqX0PUtWVGVdzV931L16uaF7V+PwAm4y6qPWoqk4MenCoL2n+3+yBn3Uy8HVs4B
RANxoOwMR7rwUHQLg/yeOImhlgJFMBXABbEmd4ewqxxGa/XM4U2ApcGX0lWsD1nLY4zjDLWNxS4L
sNH43bkCDuX8zWLiaCzS2JsKGfDPSoShnHHiMnQjckc6qwTITTZRdnP6XXm4FZrj/VeSALcrTG/X
1DwF9XkUKsJqXovggVrNNa+WnmZnpBSKUU7HfRKEmLZ8vFwXnlKJSXCabt5kMmIDdS5ohWrlKpk9
PTsbqqpZE8IAxck5wZF8Hwg/h6Qv/wxCWHEidTq76NQwvb3qMU592iv7sjADqRIvB8/9H+A6tjfk
p9WNgzAu+82KQmOOt/Mrh60kA70el1NH9nFNYpVwcQQDL8MkhhbIaOKGsUywj7luDXVo4oO7q+T2
rgZypE/m7dqUfJgm9kheEgD6UK/ce14y3WpJn7xAA41JfUozIg8QF7iYCCrX7/ftnFwOeAsC5DqZ
LG5nFQGEnpuiTCwxM5l14NZkYegNImOgqKf8wrU0qCALsUalFW9hTShqvKNDGfjC3K6GrP+bZkT1
F7da/vQyDZ/URrfJUT4CiPfUXcvoESPBo2K1f04JCGAwELaGxnT2T8zxoYAgwON/MflAEkb6r7Wg
/2DEkb5diU5zwp27ERqlG1e2WGEfNkGSv+Ea9IUhy6IQeJ3KMjwEyBmIVvJiB93S2uptWfWVRWhU
s3+TFPUBF/zblHCNEeZnwYh8JQnQZX2+kVcLrq9XF7cmF4hvfDmLP5mqf5Go0AC93VF+6LXVUL2E
wlAQlEr0a+Q+SAdMloYtifbUmCs0nalS9VjpOJi01mpB0mhiAeruZPV/fdUN7F/ype0i2umFoQf9
mn1TxJdul7ACaHVcxXEJOKswpNv+HLEdRpbZXsPGiBrnFeukSEGcWMCQflLT1DoBS+pY5VMnSwzu
YVsHarxPaPzecgF3mOOJXyIm3J7Htztd96suPH8HiuXfnVdyFJGjM6/tyu45BmbIoHgCj+B1A5mw
s00T4x1NygvA9p/MLNVJgi5Viqs6Nb2QmDFo5wiCQsSRfuIS5Rc/6MV8YAnLMJq+DHDD4JtwJ0hj
jCgn9zEuQmjQKmxKDsCAT4fvb5GdBL+J7PFMElM/regMrnm43M5zDZ00pFvqrHRl5+tZknQLI9YN
gVaVc5bUyER9PBWGmuLGvaT7uuUOmoBLGHgQRwin0LvMXHvYHk4vN3X+kbOLb+sRNUv6mXlRSCsL
zXcUcM8KA4PUFLEbGR1Roul3QCHZt5X3Wy97FRuFbQXxRVC4UDTqjL0UYNOzoBqn2+ecyctkpMXr
QZ2LaER5I1Y4fAOd/MG5CgtlywcNHgDXnyObJeZS6zmJs04GSNs3MJmipgfxPBsKs9gNus7eUz8C
5w11TB1gUBgGg4Dq+1mEx6xvhkV6F25Zmps/WuXSGaHWDgImkmepRfFTBRHK5aohYcacBexAzyCS
bsIg+zLnj9XkNABmNGhUBqixeA9t8CIzSdyJeiDQuXELDhQPwPPVru+ndieAhwCReUqzQMi/FV3w
NnfCye7oTQ1P+u3zvxLfVk5IY6IGf1u4PXgKlZpRc0lAEOSLrcnmud1d8XH47heUllEeb1IGZ31P
H/WrxZ1atfFguVNpb+XlIEm8Nx3zM5fgrX58XnHiACJ/xuL8Ea1XgPG3zD3g26d8SvjjbBoraw9B
zu/CJKa1sJ68GrAaojXybtd7PxTWtpjmgbfauK1RfL9kCTp3OhWRTgM/4rQPzoLX3zeqI0sdEuUK
LkMYT6snC6MId59Rh3SZAqdLCs33gAJlmn9swBl1Vi4IlZZaRVEc9QvW7eddDDg4A49VPPgXgv5+
V/OpLLOdRWJAv+7kfEWvA5ZnBheQ+N07Kr1caYfGvTahAwDgoVDtGkzvmAME3ryhMvkb0ZELCbVA
I3lSRrjwZkbncWSVUGl0ZXYIxwn95sK6Qewnwe/JWd7+z/7BPrJblNo7/J3QupTLYAZV6Ksr/7x/
AwD3OdeCAgRlhRhLagdYWR6iqN/yubMMGnurajTIi6JUc6DwBCG9AHMSRTD2LmTaw9ThMBclFpQq
DfiH7XD1Z4ZqWzC2qvP1ZUk2xRITVWai7/cV5y30NpSTIbLtNrGWbNAU5jgI7RGlBv7QnfM8Fedk
OpRvUNgQBOEy+irtw1SeBaGye3U9ltuQwGquKTMFlcH7Gj5Cc6SpcWtxY9XGMG1+JYiIcyYTCuED
vaFSqu2SQjvleP/ZfiqjiYrTxY241hfXz2jXJMurojcekZGBTiiGfBRm/HxQPsuKkPA2bTTUNeOF
iK/PYIy4hZxek2aQwLT6AdvjzYsDtnvTBwaaVCOhCx5N6T7hvJlsrRgGguqcmVIcdF1dkSE3zYm2
jOj+OrYAJo3nmVg8+Fvf80Lo84kgZM9L6e0zdK8tZPhH7ohiWxe7UbNoQUrzczvUKP8PW+mAjGyo
n5BKyl+h2+KrgPwRoBJIo6g12sc8zc2wPjoBQ5PbeFk6P33Wf8eeCLCTASW2nAKShs9gRhEu86cs
PoXPvB6XckVyFsIF0do2HDgQIqRgL2lFLdvOWD37LX8cq92xgaXpbb+nZ/n8lgTPY5E0Mt8Sf+/M
ItekP84raPZSnZc0/XL05A6HG1lHLJJ5GjglSNaLC+/5thXSSb2RQifdaPKuXjRkHUoEeqjG49cg
Hxl5kX4PmQtPWmzTg090SWNP3spQHQZG0yGpFfSt3N78ZUQv672S1xPyi6Fxmy+ISSAvi7ArA4+4
PyV8/HWO09AZEcGOMDB8kvXsbG/BPZSaPf/iZlM/DUutr+weNePEbapZVd9cMvVXxasxTG5e5BYa
6FIswK3pyNMAQhj7VuDZS5bVO42HlPn0+3u4/QWnfWHvb1UidcEJ/G23rYv4JNUs4IH88qJM7KWt
J9HRWSKKBKmp87wnyXWy592HS3i6k5uDzM7++Wr+0V/iDRFSQ0JVgbckCQX/MhW4hEPo07pCUTXY
IYlEpK3/6jcvCRC2neQknvLf//m84zy6MZYknwaPT7zBISPtyZE2nwrmh7CGXGDHtuQ4Nf/99T5K
m9THAAnLMqmfjeZlczmy7UOVF1Rs+fZG1S6x8D0Hi4/0KNBJHGgja4jMUASa8b5QVxK0VJBJqbsW
UwwC+dn8WBk7H7L2C2QrIbTMZLz3HNeejEICBfLGMXMtWMPwuIfapji8SFUFe46rHWj0nr/aqz9f
07U7QcI8eOCGJggd27NKZX7Ts7xfW2Uy0YqDRXUPTapVS3BlkeRvZlz5luySRR5G+GDJtj+THCu2
v/nfifPPe/3QU0yXRdSQDcbnnVe/0Hy2a/+hLp05ZTjCGo/mYepaF9TzpN+owZMVkARr+mGttBPQ
wVZqqjdaTgrJLi99PlkV3LdvJkrCe4VWFNBIWfINCTkrDxDKqXCt/eL5Jrg7oyrffAq0C3UKYMe8
OqmEqtcNMBfonCnPZsD1RmJ4bywQbqcrAHBBHJTs5PjSqOFhQGOqWSKPP3IjXdtdE02PQ2gSBF9q
AyHnPSnp0O8J48VfMquoOS+QUKppi38Jz3SXzxgMnPpb4ize5RFwQvuscvXt3AOCIxM9lou0vt5+
WjwKMFBTr2uNwpyq7aiC77d8AxPliYu5yG5WWyj/YMaihie1KPGjKcnNLSJVpeT3UAIH8vHdqDd6
aPjbgHlc2E8Pma0z23eMFST2bTdva51BAQ69tZEvufZo99+zhiGETDw+u7NTSKDIUbjnf84KsghC
q3LwOBe277/zuee354fq+PrvntWCbFzIPvh+Vk1fX9VcaSDQJcbno6KVh1DmC3N4uWb0FLe9UOgH
n8UEwincUO2CNid961KQyOmAmBcM3W7+boH7gv50kA3k1yzcpx22Ny6Q69aRIPIKGhLp1JbLB2q8
7lnt1g8oA06JbAoxFU9h7hUplFvD38QxgpO0FuQy/XeTkGiFVmnRWk8d7SDDQHM7+Wtlvn9UQR/m
a1yAOSld5l28UTcRAdTTgFIClGVBRVH7NxOouSz2gAlYC1hdULoGHZvWFfzu8RnVgURRTNpZ1Okx
suuAuSXtKCZy80ztfoDuYLVnYkotcyJlCEb9p/32dBDNIttRQg/LnULrN20gaxBc5yBQ5CvY0KkO
PKwPqC9NIOK/4YnJOOVQ8SSWKZNcNiwN/wOBh8egF31xsQWiqHZ4L2+SOstYlA054jTQ3FJPz2o+
oaVLFuHPCJARoqfqrcZJ3H8fTjghRTGPfy8BotsReJb6gFf7JrrFpwI0jajQcgw1Z4GI6grgUQKa
4NRnu4WEYj/c0hDzq5kKAJhoGoIB2CAbIZpthLEBZa/8UWyTTEeVDrmV7i/vKvgzvi06ylEZtPx4
mOZEI9Tb2YeH21B8Z0GY1/c6JuGxjr8XbOAZOF7QqvEiSpZJ06lwaLcLAMvosDvNn7C4rNAGf4wY
IaPH7AaDmVF8jUS3U4a1ySFN2Kcd4coiNSEfP2eaxA8YZr0d1VbeFQ2mk1nydlRrSRoTn6kBEYNV
G9Fng0g7YZodfV2VMzy/MeL1zh6c9ZMvXo+4twv2kXrUTFm1wZOtC7EbMZ7CJCQ+rALqG5QeEbKK
PplkQQQiZqS71HDcJ2QoA+9ZGiQZZm/pSbLnqL60gKPUChXOPRRNLNf851QMbEwnwtlz3QXaeGAn
7lvwnaWnpwekAB5ot5JxUqo41T4dRTTetlXQL7epi0MZOwwfIf0reE4Gxjzu2Fs1Hn79SXA29xxb
KeBFlvzPqUo1raV1WVvG9HyJED4LhH43XoO32ebtdKTPoloiQMEw/xxMYdPrBl7DkcNztkBdqZ+h
fPIekk9uSog/7PngiPYx3OkwePkQDa+NBUsq88LB5UsCWPDzg57SuBW7EMV/l0dih6jJA11rOiu/
8WFDeiPo+yhlNIBj04ieZsj9m7ikkHo0vXNf3OD1mHZKhIh9oyM2dpdOySr0sXgnN+30xk5PplFW
D9p7llKBCgsV9P7hpLlp0Chx8TNLGKdjWM9bY222e0gy65klWa5P1ovoOWbKF/iGXaG+y6WwglBL
3re610blISxtVAQ/+xPpaZ8KrJEjzYqwvtHeFdIsU5HVf7CwWcpN9kk7iLqh0pzdx/zFvESUKMCL
r5rTE/uitoa+DKlRihoP7pdDAdMHawTvN9+c2J2x2AliJeHY5uETwK856kKpknEdQXYSzHgHqXn/
uy/p2MuvvYkY5//cmZK/fHMercR9jl6yPR0v22VERrumfFnwjPSfmImFYB08m8M6XzhQBqNBp33E
TUx4zvhcbnB9bw9h4bJZkCG98pQBYPt3HScAu2VVurpSYPHT/XUGk5Quu0yF8g4Ib9mCpGV61MGo
7mRygNL87Oly2Mr3gpD0jobx5cIrc9NVxvWXqEEl16Mx3TCXz1nMtcZz71TRqFY+3UMugIhIWUlZ
gLse7zTqkJXMWEglnu+yawDfIFI5E7ITUIPwe5dUkjygnDk43cu9TT3rRaS2lUzTQLZfWCsEzHeQ
esJs3G+tbvNXMRiOQAUeH+NbbSfwFz5ZMa+I2NwAcVh4GYS6GIlYsWlHzgk2cPJqk4/LYvxEsYgp
x4hDG/arcWwAY+cLoUzo222xUmOmMq+IkdVH4nktAy6RGDW/os+lM7CIpvDjrH1d6uBlGzZ561Yk
jiW+JK6SWJwZ/cwa4c7eRVcn613mH4DP4ngtDjwTE8l3H7/UgoSxOxF4GBrefC0fj+WXtvbL/8Yy
AnqtKP/w5ChdfzV4ErRd7jhx387hwaNAKnRnZqV10Jgb0zSylnK7b4hiGufdS/cb9OGbHTEHknkW
7SdeAPQNysf6TEOOP+//MtElE44twFRcbw4psGpvfsoyytv3hRXOUaCuDF5PnCesooDT6UEYQ4OC
PkYnbLu71cb7Im9mOSpnE7bznZwDeW6bA2QgoyG/IsV9hWh3cw5QYVBWah60+jVRAUlaXcwR55Tx
u249zQmcPZR4dgqI2TvM5OoY/VxlgCck24xtlXdloUn4RpxswHBSM/qrU9L2dBsqjbFTM/guEBJC
PcyneUqe3w70UiT7jr+ueFNEQHzCksgQiLCmVWAIj/oI0bczKYUBpjM0I3urEnHOwRH5OMDxvqgA
bmYRWJuYWjDfpV6eS5IV64PvhwrCgWHvBxlCyXV4Hj/S3Gr4HMdm8XczF5oMDx8ZQjFExkH7KeqF
ON3a/kJ+qOEAoaQJDU1gZP2RpdgiFMacDK3dy163NOhROTBHDriwPL7uxOH5Fm2xA1Bf92kKP22o
KD5z/ZlGLtc7jpWH+AgPJGW1kExdr+KptUrydAHNrgb1fP6G7a/a5i1JzHK1a2SdhO7taI1Rq6jt
7ayYxKTQIAtvivPRMU4vsSBT97DF7r5bhi6aNXLw1ACwL9s4RFSe9uVjqjAZm4EQW/BBRJv2SPPv
rCNI2GdoqzKWmZ+AGoEalY9ku5eMMfPEjeEOODN7GXm2FWND5gfwVmaZMzObEiOk9kV+OEyfx1Vg
1NIMXMhAYPkY9qWew345l6J6YSoY3DqIogvhm8DGYiGiczfb8L37xI8rRJJPzAw2y3YMOoyj55bv
kGbkoVBxIPoaS+HrxXW3HTCy6ZnJLVyItmskGFVZiVEQZTInAtngvtCzNIujS2lamd7O+1aSeic/
fcufzUdsxk6+SuGvHSJzUxR5OXJ9JQ/gzdVMb1OtUhkUaMDSg3JielmM/mdxOURwcjgyjcgGfXdG
9Dz4CEW+nnVzS3I53PTyCvdeJGu9dkkvOShb7r0+CgTMppRfnWwEOkI43b4m5fsvO6GQEfIAzSoY
8WtIV3MDIi6zW1/x7i8eBIs9HlY6FOtPQaSX79k8ItkPmlBmZ4IugEjtzcpZOEHobw0iVso1oxPS
/Em/I8KB4QawVc4yqupBPc6cQ/QA6U6zgBmNnSf2R3q8BgtG8T2c2kp8dfG6gDkxUyikssfwwlnr
mhX9pngn0ykEhpbZXO5yxeQFrhbuDhWRRlHyw4CIRX23JE6/jK/E+7LmMU0yoL4SFFGlwOmCefia
dhznPem+LVFQMwOj0KRCIGZKoHIFNkl+NN21p0g+g5AY245DLZIhKAXJI1VbzwU5jrCRMJsqDXYi
AP4NvQw46ilohBThRChUnMVu0LOZb++IC5PR9g7TFxMl7zx6NRrVHUewCDNNiTLBOG9zQK4cc7bs
mszL0ccnWzNdl7zYzTjOLjy/ARxPgwZurcpYMHGI9Nl919KXeS8QERPoe2joKjpzxBbg0+CmmH13
oYO3XKxztPICkl3fuTAdwfoEVUDF9VyGtLmtPSVPLwl2CLeIjTxV32/rHto2Qph/8pRz0NBh7KPV
I4eOo2Yj+hlt16xIyPHGiBR3Iz6e8hO3oYVk1qXsNk4wlhnhHTFqvoSj1aUbZPf0qK7UEFP6B2li
1UqpL2eG9s2qnHt/Et3fkrRNrPQCaP4/9zh+DhmhcP3vlQnrCV/9B7fzyrcyMAjAcjSQVDcXSUAD
XLZhGYy4zIRTYWMP8oDcDOwVqS1JG7JbwYm0uMh22YSb+yUTfsyeV9C4aSiezLY8u7feKpSl5bqP
4XQv5hbEm+P0Us6/2OAoKkmkNVmcaLxFThKWNkAu0HlE9sA/1PygYKeyr7L8EJYbFzIB0sTfo/Mm
coByI8RG6KXt9Dh1Xp+n4bOUYNS2Jq8sPj/o520yiLgGIe7M4Z8mgDv01nI6zZ9f5LuO0iBxY6wr
SHX964ZxPbrln1fprjw9RbkoUbtpzhIejqO/+Mr5RMlvpgNGbmTWZ1Kva/AXoF33EsRRCNUG+/pr
sZORnGfid0Oyg/tS38VPs84ylZbeSv2KQFMlf1JvTBHorTIyGijiG92Cf20mHO6bd4CFGsUgGXsU
bzAqNL7Xi0P6ieTp/qM3DctfFUoUeSXhAoUsN11ek+Gw+fImnlPQfBsQeLGppUToES2VYOK9me5k
Ig1eSN39fGOkk4PSt5cCV5kjI/KD/4pcNK9poAnWV68dBGJ3ZO1Ac+MCUt40o8yYZg5c7Cnzfe7M
f+YnLLiIbnGY7Bx7+ut7X0kI6MxBuI9OwzLP5w/jufcKqt0ey6a3YSHbf05Swhcs8jnk/5Hf63zh
uuXmL/uoQgtNjN0zAeFSrlrtu6qemFOQPMi1xd34X0K4qAUy8vBs423Qe8qIUleJxC8IklER5mBk
paqJvaTp1QWKQPVu/vB92Guf4VEtsTHaoqGoYbkF8NJi4CGsBE5LVNzNuitEHpitcN0VPZzsaM+1
eX0IiU82FnSej5S5EoD7gFMrxgmm2vA1acghgAWJb0QEoLyATR0a7E3WO+rjZ39484xRaQZtM+8C
IQAS47sg1pU2ONJYNsnMvJBYdtTG9Gkh5M9+3GQG+/szwprTfGE02u/ShuNxAAeSlsf24FQvPie6
S39N9x1nL2BVb+AQOr2OwQOAPkYqZXO1NwEdPL6Lw9bYjntCfRSlTbTGzu2i9x2/ZL3Mar+b/M4T
W9wpZofNnCOXrr6M8VQAJ/GqJK/lmH/kmwrsKYVIEIyR2/Lgc0pXMS9ncDDlQ3lBBYP3WVJbnk0Q
q5PRlg9CU/wH1t8ccEJC5f7imHjmevHYBVepDKbW1b9y5aNJ4j4x4uM0eDlcpUfOqT18SeqUEaEo
RF2dZFNkphza5qH+rtGPbBOZXNsjAuupsylBPpkYzV3qwr2BEtPvEKyyx/UwAd8m5lWYe3GvW0rU
e36kVZGqgwsiHCu4PmfcDgy1GBmiUmaKYPmikOVSC5CJtznnH+yK33SIGef55fYo53b4SGLSfsNT
gdOCwOgi3c9VIuYcj67z+gHXQoAW6PDhVWKnBw9LykYYLJuWjJbNvdYzv4mT+yJ/cObecNe1MO7v
CsGKoxSfpnWTtgOJsNKsaMVrEaCxsLBcalu+4Z0dyQ4dCDbo4iA97dA/LuMbNz2pRbHxmWCe4lUp
7nnJN9W23ruXjyYeWBgmdMuOZBDmGT7y6UcKEOqdPyqyxXHHnPv4ApWUYEGK73Ffc9ds5+vauAID
DXpUpFrLO7jOzV/X/ziGLDMYGst9ioSQ+zI9jhbfIIE5p8xW4DiCigLr0Qfgtc6CM1QJe6jDEmq3
2qcKec9YwCSWjv80AuR0qv9y2B0XsHCSunm0BxgbN1Oi2L2hTiLmvJGz6ya14QUIqTrviPc4b0xq
AT/BtuLb/O8FteV87+3WztTsGLWUKxaPvm+s6lWf2fMq1DAJdTzOQgy9fo0azmysmFLCN9Yik/0k
MpUZ/5E6S8aq3hWezHnsDNPMZpCLqnIEeNivPqCAqJMtQN9INb1Q8Pp7SGedQQnQYL5uHK1JAO21
ftqT5o37RTNz5WM2Lc9cAlPWs41fTK1PTPdwtDH7+VfVVThwoV4pGMbwroEij901Fv7fX237WBkn
vR8rv4IH2+MNzMde9JLMHYD2Wn92VaVbY5kA5KW5UPzWSSOBUeli4eQfWV7waSnTV38R+CcllGp/
Vkkn6qFk+kHK7N7spQU+/T8onEHs8jpVoc91i/dbaKbLrVKs0ueispeWWNECri2NxkdJmSRbtF+s
GnLXbskNXGpDlZLtzVhTgQKPRf3idG9eTo40/cQ6BhJ7nPbbUoDF6oBAaSL3FI0di8HzyOsGhiqh
VnGZGbEXw1wTmps9AtQgVUQlmmpFvl8uDXwkl6TWvwS7Cjp7ikO04tln8cwVYQ2wvsKHr8+Rvzof
c9/I/MhenwSjlc0M0FB7ln/KniAjKEyo0W/i2Oxi4/fshTbhXfhNsSseTyLkJ8jnTWeMheS8NaJD
7glocOLHorKk2IiLc4hqGkAEA17b1aSQkR4RV0J+Jwd4A7DqIKXDiaPLlJ+4f127p23/eEhlNc0G
tHiMBvjRu6+/iaJZor4KAu1XQrRgbBUIg70OzqbFwwozNqZlK4bYbD3iAYCb8S/ylAENqK4m2QAX
5W4FcJ1ExY67I7Sg+48y8teA6M7eQ7xgYGCXy/wL2+1SYlzv8RIzlsjuY7uzXbc4AFVBNpuT7VxX
R7AgmEdGSwLGt6gITfMZO3zc8n2ZjtYy5SDJHLxz03DaDymcIXFZFtCwY5Vz6eIOIcwrkSPIsbkr
B9jrRSBd5jY0H+jCf+QfYcUnrxG2helEFQz0bFuPBcoVzkoo1ZomOx9PARej10GhfK0R2wpvI0RT
Q+oxSm1DgSyp+XXaFD4lUWExiVWHOak/DqGt65nZnpin0BSLCeJTEQI0S/4CLWY0gxxf3X1timI3
GVvq4Vr5wfE4UoWln6M1KsNkdi4094hdD5wSOxpooIDUJDgm5vPpgaQ5jJjVrIG+7LC4y/gsv0VA
0AvlkFYe/++7YBzW3qDjADO5oUMQA3VCL9ov5YjAhM7s3Nk4BmpCAN7V1euondtHv8AzIK/gH/ap
AfnRe7OBkPLIguwEpTdYjIg5DPglyth3579Kcc3TjoHiSh2GZPQKnGrGxS2sjelFx2WYnONvAC3y
xMVfPlS8WX4dBtOMRrenQMc7dcKAGBU/tpD9CHDrI8ugEA3TOl6uzTfhIUUDE+cmd5KWyhZ2oUa+
VLNTYWWs5H4zwy8Xd1Hh4+dU+6hj5Th1S+xlyl/pK7V8/A76Fxvl+MIYP+FflAQp9mjt5ZFhzwso
qj1xHMep1bDYRM2E6+gIxv/uPRLVz0e9OkZoimX5r+5WDD55pfn3Am+8dzbB741qiM6DNAazgbzW
SDNBJlX77RjVy05y78K82E7Wn8W6OTF/KnX/ildvIihxtlBJBTozghWOfcapgcLsZ3i+BLD/5xXd
mafTVEskq+gXv3socQlSNA/UO3vTc7mZaCa8GiwDOkf0tdLHDoeu+3ivBawSLmricR8OM86TCy/Z
YerfvyJ2PQv6RjGJWBxrKUlxKh/tRGlAgoXRI/NHnPZqsns0QbtTzOzeerSQTf0sZwoxv+Q5p3Rw
61S8nDszcrEdSK8+5FqZxq1jzneQVknmCGa0dJs6Oq52YHS4aXsjOdnuc7ikJ5IzVLCYOW0XugHt
ReZm9mEcsfTEvZq+v/b/BjFuLwt1f2PmTSZ0PQM5deNtnHWQHqvTiHgQWQGy+PSwDzCENsON7Zem
cRoF9R/J7liyaan6gsKkqrxwf7jyER8iALG2hega5iiw+4SuUv9vbbbfzj6QvIB0jTmg/GzqA4gc
OI8wYlCtSsD4kzwBi/ox1bX11nBW9XyubvB1QqEfheoMAGY1TbbTbQiAbAnQCsgQzXXmZIQ4UI40
a/fpq+AArtl17kkSEutY9Zwmiarf27jd5d2M0f7Caup5mrvs+4UkDBrrsuYl/fbtEdexx13Fmjzn
g4HW3E15jinzAbFk7+XCV19cHsZI+IipGV0L8rTIy/yDbJyd0uHf/UIrsG5OyhqEdXXgbX/H4vcO
K9/rrE90R1BwhmMuRNcI/Uk+q9+c1LRxTHmN0Wx0JjSkYS0QFm3RSl27MeMZLAPt52q6BvdNX2JG
PZ8iZP+qfVUulTudNFNs+2/A9chN6Tng/bvrKArutDm6t5WlJTyxXSokfBKL97IIPpG1ukAkX+9V
iDeb6kkzSp//e6aR/sssaPHEh64s0u1+NkCdvkI1vaGax55JRIRWC4R81NRULfA7C7IBWWIiIPzy
yWZJcAu3OBVZHg/Vw5znJJDu0C8oTrLiQqValX8SnoL4bGRD7OV+OwS8OSxMMft1briqOY67qCb6
nMOhEFc35FQuJUaJwc00PhI7T+2yRzw7F7P+8VOp8zGscoqqrgejWhQ/1sIIefhhbBaWD5URnh6f
l8yJABH6E2/Wh9CUn16/Znpi17hz3hxc7xIwGJHVP1VgDc5hJdq1cf031iEuMbwkQ8iMKlEnBcC9
eZPDD5kZPxKRMJZBLBaYMccZqFy7zlhvLTCbZH0rDv/dfyRyaj59sIPKINeCbaaf5HumFhINS3xW
oJjvXfvxCkoEAif35/kIUpl1O3W2iWs1cUPvP2z5yfpVQeH30vRTsi+04vdTfqZmrNOaXrC9xF+J
BDubOtt3rSMGLKC0ZBRfLLP8Ucos2ZHcT/XphAKea17Kdn9qSfjPUFXALF28ExFSAPXbe9iDrkcN
tprMWn3conCNpIeFLZPXdKJWQ17e8UuAW9C17q/iWo30h83vlLuOLgijrKcKHeoRJ2ymGH+32cy1
3mHTSbY8HEzuMXdIclBgtnGiX64eoiyyI/XSmMUXGi3QraEk7YydYCP6Lajb4bj5jbQtzjrHUnii
u9Ai5nAH9QdTWWnMQtbO4QzQb9llC/Fn2OXkIBR6E/m5ahM0HxV1XLpmqt/Edmuc+JreapC23vTq
YjUqVugyiYxrKVVW+A/iIfsTccOMGBo+gZoL5SBrSpVyxJwi1EbFAtyh4wokOY65QVv1QN0jlbEg
NWFcsUfG9ZM6dWtgoTVMcMmR1eMRKbIm/UfRW868CgXNop+e+rBJfEi6X+m7cLEm/Ti78mLNxaAB
6sgQ9/RjsJyNZvwo2b3lM87PR0KEDTLmFNXqFjM8LkjKb3gbh5dHsSM/ce9SrvB6uCU7uqPbqbRB
yw0RZWmgzcDqmaUI4/9lwQBZpDfrtPEpmzDo+wm9SBIHuU38Vd3CPI/g6z8szfxe47VRUCd6+/9H
tHBNkVNAYLyykuqjW7Irti1tgHzzV2VvHdkQ01VVf7D7A/JdvKiwYVR+32vr9TmPA7hniG+uQuj0
sSjmthDLAExurMW/FGj/bkZi1D9DYZK7VXxzq0Gb8jV6TASsCyUeKE0R4zpMbd9o8DJVHkfdA/Qj
5PBSVJoan8V3P/HDqBiU6T0ebFohLLyOyoSmc+Wy2v4Nhs61FSSwNnE+0UCktnErO54SC6mFptXZ
4nPVQ7F8egtodSY/Bh7OP6vRjGciQzSOeBPjgm5rHYONmi9/xal1ujT/7DchpUtPov+YlRO0nQFF
vrJUssj64zU6s4OQHmP3ZHFFxnoR/9lIVyvE2DLwj/vtioKfmOxxBts0cmrs06IwI24RYZIic8OZ
fqXL/dCLN9QWlGzs3sZW/OlyOJQZlsKjYM+v3foPhqhkZ5sf4Nv3TRqeoJ359Oy9pvXZeNxy/KO7
vJ1ZlYW/FJmCq98o927DYpd3gml2LqVX7f0bQe/juKDXZXCzvzIRV+DpBIXdU3aYdgv4vRcJubU5
LG4/FvrAD2vibGJ9kxKkoo5YrUsyR/R9HzHd3G7oHDfKBV1kz2SuChJ6yGVM/KEo/EKOXz9v30OC
5eUHqVrNeAcZLc/mxA4UT0lvCo9ZskZD2din4tdv+FHw2+5cocSqLFSfeXtM6XKJD1bo/FviJqC/
pZSLKDkFxRUjwT6FkU8rPklzREbXITmFtROCT3OU2Q6MUg5hP82+Bc1M8yPRmHEY/3bvUJGDxCUe
Jkq1rWqb82vECGxGKUhBZlGskCw5bptf+TcelqtmQMn0MIx5Jde9vKvnUwp3Z/SSwo/NL6wjG9wO
ZfMUr9ZtP9tI+sNeMv175WP1skzaylfEpXpVw/YQ2YQ9+AU5VRlDMYZV4te+enII+8hP19TXlcWh
qPzFyLJPoXGKlfzv+XIKSITHTQRuhnml2R4Rbc6PCjo7ocGuC+U3f9X7Mo38mUwp7qDbe1PHDWx0
q79avjE49VNAkputoXIsvXntu241tDFyWO4AhXj49vXUJbqlGwvsFjEvkdBVAvg5AOvkJODDu7vB
tLImmDK3dgFMg7YFP9XjWD/Xs7GSscsOeUP19wj8tKAaTZvaP05VViYEStGTUTI5nfaf2PSZow/9
+seiXrO34ZEUlY5HUZXnqTaarCmLNOMamupjiWn+zMQuaY7g4zVkcpkInX9jR3DoqjW57BY/Ndna
al81epdnrr9O00lt6BsvdCGhvoWxPSCU/wL2ARxEKAMti/rHBhg0gwdO1n32pZ8NLu9FEvUOH0YF
HcCh1Gq9masLKF0rxZr76BEEzWAM11uu60TpGZ0ES7gLhkMykmuPIlnlMBuBd9zUpoIVS2lV4egm
7MFPpGtSCqPwvVWt29U7Rf1xYatU3qLxp/i6M45GBjMKTJkFj1P09H7yUGnz39TI5rweJ+Hn1uGZ
iJq7U/oWfqTENoGuVabKr1FI81A+FQbzftWXKB+MJzwSN8qfBv3PpgZdRQjzZd2CM3nvo+zN33a8
oMyDTWldzo98eSxjDLX6M7rJGUnoaRzjnyBe51JPwkUGsJag3WoLv+z6l+3kFHu9viwgZ2bwQvaO
Oy2KVTnFbyIIC4ko/iqCzcJifJ9eojJR5lNKuqtn/iPokvBlcl/vtFB30XdLkWq6eSLMV5uIeuLe
xuWOXFlq4I3EfnbS1SnJXcHEnKayudeFNuRvqZi/FNjK/mXUfxKrpDjdIqITHjbqNWEN/Qb1OtK5
NsvMxFM/z/sIOjxEWTOz7O9h8z0p6tobvb24VuL9G0JT/px+OHpRxPGNdmCKccfOjzhHnI1NAat9
8V53uPU7O7ArENjuSEQOLUgdsXXWT6b5V2FrEoxwaG3IMNDB8uEiw92fW0WGIAIxez5xSYCG6x+Q
dWYx6ZF061FVYEW6XNsCEKgpynl7n7a4CLwK84hlRhDtEomcKi8zhoZPWKpH1XPkU+vfsldHDlpB
8Kovq4iMGT7wSnvSlXsMy8yO01fLfgwvi+YA8/CgUNwN+CN5iPOeCSduRNPqaVWBUgcW6yBG8PXp
5PP/oracBcY7f/aj++LRxP7KhcrbLkdGpt4flR4wDY8cXBLDhGGihQ2llK8HoIMsKWvK6D1TGWAw
2pcV9kLIDNRc9LtX7t24Nejoi5Myrp3LG7gwap0x1ImjwfgxWkuw3a0tqoJoRNSQ7lXBsEVxnWhj
kQqYDoHxhrBYSW8ud3OAQbcCQs4EZJIpQTQmzCHDEMdf5tbBAg0ODl9LhkvN2ILnFuN11uapzoew
Qaa4o2dKQELRG968t4upubxDnrZbGtc4zsMWkWoShniMLAQKIP868VPPvF294gFYNlW8MfNiPMpl
H0nIPo8NRpb2KPnRes5r/iMTB9tL1keNY30/OGuPPnF+/OqFfmVKBuD2talk9jO+4zsqtJMNydfr
ZeI/UHauXK2KRbDWms2sdgFBVOtaOvmosfcCbOhzOv7pwZMINCf4rk2WKAPgvi3D0Q1ek85hWFdx
vsG54RT81505WdC9D6CCNrnb2BMc7s7EvZkUhUQigsQ9zLN9woSLGFEa5iig9dwbehRGIUDw9QYO
hL52Rax+2QztG2OQIzMogd9FuRwQxLKz+7B8bjpn5ywNSFCeUolNlYHWQp8/YUK16aX+eh2PpODq
jj7kU2dSJ9okk4TIGUhurdfhe4Xae0rMY5k6wnIsrYkZbSXK9w9oj7w6AYPFFz80zaz3SB19aWsw
BBcABNn/bQKUPEDFFGkoFoh78uU6scOfu0go8maBeHPlVlFfTUvy19Rg/sozOS24BkTSqH4USQG8
UufilEu7t+hxxbTkpGeLAsmqo3iOaNy5VJcRvrX8qzhFCEuK0NKN4v+WkAX0XcpWkKtOaBruoRUm
3jzCuj+LWC4HNrey+QmaSaqd7XBRLXUD0hN/LvU544I8OLGRch3daNMKIff9kx0P43a/3jPXkEEP
lYbgOsC4J+L45Trn4g+peArYUk3aRcsVBgZHPShqdlA5o6tJXfeXDUh0QuxEaoL7KtTVb+1bmJBH
hBqEGM/BN95rswE+e6NuNdx6vRh04fUSCVl+3GG7PLYnqdTDMQWIWGUHwX35OSZiUKdXXSmkyARI
jLiYJ1MRRM60rU6g89jq7LEI6U7RZw1iNbxLLaEsPKzTreBGYMvjxv5W2Oj0ry9kKtHCUbDaZ70e
K+S4SQLt9//S5DxzqIuZZOh0IL6MjjAmLjEIV7kRS3IRwrFPyf0SElgS1jHoPuj+b0/S5Ucp4yza
xMF1kb2HxxuVOovas+tp62NdYcX+03N6VN4XFvecnpmpDaZI6cBvzcEDNmWB1C3ukyVPhADFdSf7
qneL7Z8G/Ur2WsuADf8SR7wRAOObKi8zCeng2EIBIotfdAsw32nuhMdB0x1oDYsYZ8VckDX67UTW
WERDjyElSnIB5Ahx+uQlLuMaizUiVPILSF4rm68tfWo4bhkNOSZa+MgBEdNYSzPSSXFv2Ok/L9Tt
6/WIUGYaJbiC442PKgie6z1qXP7a9RhTpolYzWg0D0zjsOUfBEJATYJCDzc8voAsZ8e3xuMa73AH
8LP4dReBN5VBwGiS1RP68kXsmNTWQdMt0Dcfax2rn36cdYw2AErB9KDidSPt6LXhQT+YS+kFG2c2
R1Wniek19YY6kSbm5X/QuG0zi8y6MXu6RPluoCE7rt8ymD5NQsUPcIlyj7M2qnyKNMzxJdFRhg63
DActZghHWPn/yoXZCKV5dr6da1/KDtEK2dgG/OZwNhhRI/O0Hhie4XHEhWAZFXOVxJRwa4h6IEA3
hliu3s9SotoiOVbkUT7/XD0RyMEOYnQVoTWhte0hQSJjC8cIum6xGUx2rKxDWoUMaJUqVLp4cs/4
gWfuzs5oh9V4od2BJFcBN4pfA4wGBHRWn+MJaLFYY+lBz/ShoFtv2Mf6AguR6cYQlkUzDYt1Lu2g
13/R0SY/PHaAoR5gP7ALx3v9VxkN4j9F3q1VheD7A4E9EsAzK3CSR4SpQp7l3JoAdg2GHvGkxtzd
+7klbfWGMCZBnS/oj+J0Xx6yZ7TzPe8jb+tDGjL0EOePYkUbIK/+1u8QTobkE46nazpk5bjV3xDr
yjUlMFx+HdTuBItyHjy9FZQa7b/rMiYOhlZwI6+MSqMyx5xuxmMWN6b3EhXabzTeqUBcbZUF0IM/
cVHYpZbMQmyV0U7fKpoRnvkkO8Qhb55Yec5aGbNHeWWK8a0QDdzKN3F+1JeogE2U1p6E4qbYi4Yv
DQ8IEx3ogGFg1AN6TS6LLKx6hp2VA+2RN5m+iH+vGQPfW/W4w0+jFZn2ScAR4Op+y74k1x9bFpw8
RfFU36u3Noc0IO8YJ3zU56ttQKCy1bEo2ds8ZxRNX5h6hIybCCkDctztjfqKb7sKGN/Z9NNaC4sM
RmRCbYN8ACJIEmY2X9x6RqoCrSH9Zyzod+INC8FWm2aWc/AMge+32N8q0zJJtfNz6/DeA7JBF5G6
u+b8/TbCRpyOwffE8C6h1kjrH0KUMZtvXmG8mZk0QNCSiZS0O4vbyMZJUMgiSiu9U+XuX72uLxua
Yu6daVxBJkugUYs95ZBDetZog2+aiT6rXZkJ7GuCOGJnR7TYX75xK3C1Eh4VqltUbi3KVr+a51oh
1F/4XdtpEHnG7ChBPt9CaoRO4JHwdWM+dzpb1926hDH7dL2KlqpoF2HtfiT199VD+yi94it7ZorA
YnPM9hxp6M60X/VeWQ6d9XagA/DdRoe4+08LVxLAueG2/JMWszlRB3C0zv6uWS5ML0xG8DYHF1ZP
RycAfpBvVWNy5AHsw4i9QFxFoVNBwkjE9xVp37oxEz0Q82fSJ03HNxzvGuKRTLk6TOiSHJIuFP4M
EijSHnBlcRHmlgzz6hWdraW+Wd+x1htmTDQ26AAQopGEKoE+mcHlbLfyXSbWDP5dRXEY5iPLmXKh
uggLkhnGF9jB+AFs04nom7QhNi0zHL394TbMX2sqnIOgFvHO+jRfQHnzAX4E9T3VzQHxrYBQPDkm
/0HuF7AnY0AiZWVrD1nF/4gV0k67wXN8QKZHm+2hmS8Hl0hr7+YsjhABm/wmhxaLw1zGJq7nXWqN
kF4IEIs5Nlx45rkAC6OYpuKizRQEIIrOyFw4hGexpBSMT1XYJPzCvGR4e/+qGWz5XpScUsS+4CQQ
tZYg0uZ3ZnMLPHB0OdFhxin34z92bkul5vUS+TR/j0Uh827NDNaEg76rZvV5zHMLgsjX7Pt0Efpa
AJLhp5jOAlpI8T9IR9yjJN9xrFmetuxNLGrcB0anzWauoZP38jAbaSSE3G7ZarX2zUfqRVzg+w9S
mGzB9UPvT/89AHx2/bqC+Qu+qri/NIteurvfcM426PtNJ9a2lMzTqx5cX+iM0VzzvkD9ucJi4bIB
V3eF+xwj1ql0c01p9BdegYg+7lEJDrgixh9MCvT3Dr0YaX+eOhGUuu3Lv7hEaNzy4iJj3KgeSCnQ
Mt0ytfBTUmfpeQUotX/QOSr0pyonQRQdCZ020Clp8uSPCEdaingwmH21xwgZbtJfCsrj3Ly7zHhs
JjRW5bdGklXqqmYBQjnoLzhCZOOdHshtFTSvIY1f+/F31KqQMKX2geYn/XNv11V5ka+CtKUNeSBA
xzpiSyB38T3MRfVzEN2FdSXlHTHIPk5lH+wGO40dUpS/R94ydWY6UTgmmH4GWqafl9ZzahuEgbk9
3xibtOXyV0UhgPr51RejELvqjKyttVJj5Cjf5ErkTgzEVvUY/AtqSHrMmL0bm94ubCiXf7swicd/
+41nsZY5RzTg73fXUvzCoW4+NpKV0wE0qr02IUo19XWFXj/3Lr7z9rRZoKDM2ndObHofuB7QKHpB
Jltw8rmXiYcMF3l7/2fSbuzW52wI9OUEkyRrpPQtN3QN4FqvrCLOCSa+E25hS9ppld/Wj/BIKw1e
W4mkb0XfWEkjR3ldBuwRhaMDF9CfNLM3DJNSHFP6UYDFRlbxPrklakB6w8SrEIUQgYRBaeKWTk8k
6iUcAW82q5WYrJtW+naNz3mnnkKfvpqVAvx0LPngcLIdiz4UIRaf4H8xR1rlhhiw+1OLyQxBHn7W
+wSFre2uUkPGg32eJSLXGybRz5LVeK34AxAzx0vPBCapwFKXft3cjGQmSN31QpoTIrxkMkRRHXeB
oK5gTDTFNsKFMdA9O6SXP/wedgI9TVsWmRVq+oRzA8s5LEdKJ4aIBvbMlgKDsN6MUOpcCP7H0S05
e74Dij8lfPTApkfYSCirxaNyLkky+6AmNtn2GWMRpd9ZQbwRAUnHuN2q4fEsB+1vrr2ORq6XJflB
cERdv8UWLH8PMPNteK4LT20MuBbRmqj8psN/YKECwUV4yyt73UakAdUXM/dpmOQml5ELj6cQI3Nk
ftMnxUQIMO+JvZGE2G878sS2Ik5hHi04wh31XsY00KAg5QHqKFoPapNHwC03SFupbvBl0Yy3uLvF
5MZU5W/RTe9gi4x3oh272JnLa/62o7sl1ZkQ3Hg6fPRUI8r7px0GzqbSRZt8FBaW/B5LdJL/oeiT
x0glk31JTsgjx6Rr0/hb8cW4csNl/VzbqIbZDS0hqHtaKHrRYqkP7SC/xitk11OvhL33npF1jK6h
6uoHp0FahlTPqZAy/sPIwoTGFC+9+qOBURGFNMJbcQ5LnWB6XOSSL1Mclig+uj3yJ0TZ56EDTIUt
4a+RTe4/I4jh1iPWmcHFn8CE9NQPgjBXQhpRlcvZ4W0FFOkzKzYsNhhu/ooVD0beKrdAnPwvmWSL
W37H21z1iqSjVfjwzJ6i8oq6uqC70ZDJqCclEY9BuSW7pqh1C3RcPFXXDEYDuXwCaVce/5lSx+AJ
Qh15hkO4kVJnTLYR+chYfwVhB/Pg09yPdJj5XjtugRvRn7Wi1IFlKwI50etgmXKbdtjGJEBID3mC
0CnWEu738ybcrGDs1MC/PyjRP2RNT8VSqHuuoTMaB9RMN0dEwnI+4Br/tMper1+NftWPbUsXZYGh
4Qjf8xXNlrbOcGc+F1K1gl2CDeiuE/4X8cUqAa1r5rBbCjnvwss+Povo6ziFp6gKMQYzKQZQ+vNJ
aTxOxDdV0SYItiXEO3QFJei9hxCgHSs5Z+tjYgcdNVmqhSzL9DuDaZd/4+9Jm1HwY3CoALhMaoiu
oWb99GHYthwbmZ+oBjWaS7Fa1SYKuUi+gSNUbon0eElLMYE4whHhyYFifgoByIWTuep78mZtVsDy
9RGAHXawCh9sbDDWu+cWyiI8TIYabOO6z1aqmMnD3sZT8t4IbaGvd/T0KVh7JFajXTsTKWp9HlAl
FObMkPvSFUo/Zcp5+gHf4kHNmsxHYO6fL1uCGoDLHHJXqwbg7nlAR7xSy0TIk61W8bL0M/SO2eGC
U6j8jZ5ESIsfKstpPE5Uhn79fo25p8h2BVI1+hyTp2ICYRThlB7z1LFOj+dVzd+5Y/GxgAWzhJZM
FmDLOiR3wMICM58RxqywhRy/DuCRYxtuU/5RDb0wrU6AVe0NTLbwz2b5pIed+2Q9bY2USMfxz/gD
LEnACc/l29ggQsQVE9p+dbNa9PJ7Sr7SKwNBBkvMn2KdW7nFNZFXbHOGdg80vJgVbP9zvDjSFrvO
imLxymYlH4f5BEHQa97QzOA1o5TWrfaF5axY/th2U/K86nqR+9w715AP/yFxnf4SLA+M5eGyybim
+S368BRzwmv8JDN1wihOlYhd8D4N1LZb5KGqGVfwie3IyawcreLAKumcK3Yx5Of6z7CWGrlnCuVY
pZ0nVoa1ZeAaN74ULVikG6cSdrc/OdiAC1GXpnvJUEmUx7UNhvhNWpeaB61DCFJuFLK9qPvTrYDq
EmO8WDqZMZgxInDs8xlbfhPYSGj5Ju4sJmS+Gud/MQtiC2aehEakm5D1mg8Nb0+BQ8E5H7ac2TN1
qfSY/Vsd8SNW6vjONPpjUN620YHVZJ/OU9ELA9HRH3mfZdg+ehNzfrNNssTgR8WramxEFs4RlYMA
a/jXGdZSNJkgqGRCPMKk1xstYO2vPfRZGDFfGM31GDBAU2fLa/my2ei1f4LzXg6UhqFz7p6XzqQr
jCtagAf2DxYISYUqoUNauOqWpUpU1wFlxEcFeVexH4Ys55c+x+nsbrGo3q/duFjKiOjMCQijpbKB
/Ls8O2XQHhjaz5nS0h2s4Ow1SK/3bzmmtH9AxAuBF0k4ompG8p1D+If8Gn/XYRbSDiPd7i+MDbdq
8v5Ni5TR/yaiVLwHgKfsW2KqjAW/CjG72c/YE/KTCSLidoEkkfp/YK1NtPnkcykHMjXu52KGJdHE
Hk9Z2h4dVB9PEgYNRH2MGiKnipqJ49HaFpwOarqVw3OdKpJV9zVKlhmgHfvqOW0+gkObJ4kc0PMA
zgw8a9P4gVHJX360kEaVGiczd3S8hKZ78Wu3soed2A8b0SNNam5xqkxMcbG/UtHhZn3fE/h+8oMs
rOa1SF/jrQuYDcW5uYYFaIbhVs12+2WF6Dc+6yLgOIDewViMuaeJzvyEMrQfPqGD5OIZ/3onWiN7
lJcJQNy5G6toe6FGuWW1LmzG//44ZrXoanZEHS2ntXhvjuURgrzvV0iK0tPEtroa4EOAvIoV2jx2
N8wH6+fwkNZdJKy2MlwiZMUcWv/alcoVmn6MPImkk232Pc5h0t5g8RQmberxiyKYd2H+QaeBctqT
24d6Cq07HRuStUboBbACnN6oFjY48G4VIwsCYdJq4m3ra91nviPccO7NqaFpMK257d7QEYUEzQKz
1+5VBGo6W4RpKx7jTx8uNEGw1T2HgOsca8BqSgY/E8oc74pMxkw0q4i3/74aSZp3xsoZF1bB4R+l
sSZGG3uqjMywBPR5HzcBB81x8YUMzHJZjepyW6y/2ZmFE4E3fq9Px5RorTvXPqlE/y19f17tcm6C
oGi7tG7iE4vdzNtRlsWpanRei1tu/Fb/iJBX9lllKKj0mzIY8Oi/kU+Mtcb+5fnFT+x4npk/pQhV
B4C0zM27d7Xfe2T7d9zMHGgwcpFApa+112EZ4mfj3LThKYqR30rBdBBh6VZRW4/S0bdeYagIJ/5b
naDQlByw5pXbG2sUQn/IvmlIBs4I7Wk/K53xfSFaBO9v+6sxlFNvONcTGF8laP8LShozoud1UH/n
GVX872b2A++4nXjKgolXpQlPm0RsQEiA3vKyHU+UCckjXqBWLpH/WtGbNQNoDX0hsXJ2RI74mG5H
RJSgHo1jARrYvzjrkqye+hPUCYnSRADQ0nlBV5JeDhdo4GhBqp4P7TmUXGiCIfPbj3OfcJsN77fH
0fd9j6E+pLplma+03nj0tjAQElp9v00EWV24Q+F5arBsXWuemm6kO4FGqk8J8ZmFgrus8BRudRp2
j3ys8kNZAcodlNcQSLoulj2T1NQJAZgLhTXfmJftjsjJ/4lDvz4SuSLeRjeSqjMJ0ZMTlfiBikX4
ilfVzZ/z+3IdFhV8x95Mz6e4OH5OxRNtRGsvdmraIfvWVakbMErziQbHqk3Wh1KK5OYbS3PyHRhn
BJlJQU9MG41Ln3Lu4VQtT2zAdEAPKX3USSE1pmIAjeUBZIIiBAqWqZtq/2ASe435AJFcXwpFeLZG
bE5l055KNKA7vYFWlVWzuDORJ+NIPYvgmY55xgoSsRDk3x0VKEOaGz4uJZkhzEzpIBZqAcbVHWlm
iBHFZV6FLlIVmns0r01ZvrSihJHeGWWhTibstbeMvAnta0bs5erBtm6J91YpgaeqEDC1jFxL+STV
HK82eNUGa76M+1muIulDWU05/AZPe6Qefg1G/RgczZl5BhxbED7Hr5egaQe/f8Y2h9uDXd2z1eQL
FjTGetuueRrtiAlc3nSeSWkMtmTBW/pt3K/IuoJUoc5qjQTEVl+Uf7zigz/8yvwHqepTR/hGIAqZ
QEw2ihbU3zJSphp9sXDgX0J297jzaONbBDZAOa0Iy+CzttF3pohk+V6lh8m60+I07GaJ6a5uZZmM
Y9xMXAi9jqK1hy6sOjaZiWcxMIY+mhzpmu82xAd8sZQ4srbZ1yHfPRywH6xB8L4wWckbW85TG3BL
eZZh3ex8lie9bDDPNFvJ0jvVVPTfKFIPhwVth+A3DwP+PuYahJHoPsFzon/JLgE2KW2agkbs3UXu
Cm6mPACSEL15UKw9xDXgmJzUIwtsPKjvNmVzOTZLBFv1hJ3eAB0oguy6MKstniUXJ1yIfuM5j8A7
jhV0aLamegEfLEcaS2nB5QKFs8zq+yU5ZImw3hdUHMXX+hZe7YpqQK0XRNPFJSttZ1fj2m483X1y
USPj5vG7zgrje2sjsJNRD1ySjF2l2q/fPfftliAXIVG9cqscLT4sWnap7AJ26c3sNgW4gsCKJrbY
uf0X1E3HUn//2h5pT7qhrj5PtVmUtEedpkRwJVxL7MFicaJDJt3v8PkP3jNNjGhETJ5dOIg1vdG4
6e36ZEkAVyOsw1u1f3w0BYwn5JpsjN9vpQZy6TqJqlrWFiTvX+jGDMIdvbegDKgwEScdKRhWrPJ6
IqOLk0xth0TSisf6Kxky6lahHxmydrliLshuQjmewbAwHVwU/eFhaKOKyQzvdpKvT+M2KsUtbs1e
unPG2KAJ37oP+Y4CgeouuNnFVEotWdMEcNAK49tUAn2TEoybCAanen4MC/wqMO+c6hVEpZjYH/tQ
8+lYm9ncia9oZ9UD2hQ0nPDBMnoMFTUFBEoWVQJ6nPCKuBgw4vGIY2NNGizSgW0krRno5Fgfyh16
qcobnkRLEDwcXPC4mxR4KQgFutT5Z1F+Zt/WBAcdAp9mPciOYyT+CuXn56snZkSQKe3Gs6H7jrha
C7wUiMXX886QnX4VolFQpCYiNbJoRqRCYTl1WRiZ3KWoCSw9ResKUxwBNoEf/w3TWy8oer9SgaTu
nkbfTa80xJt7P2ly8RDDfdPsTVYSKzQxt4wejHuiGeIU4Eia/oWv6MAIdEsVNCBS1FCKNhFs+s2T
hujuC7VzlPsx3IH3h72Dvv4OH28M2Jgz2WhkgTwp4PfRuXlYIKvFxDtf1mtKOSIyd/hfKZngggoH
hbKlg45E4IRICDIKVwoftXWAXgAgdu6TdNYbJoOwCDB2jrjkOOJUhQLw94fTd8OPpJdr8jtoTmuH
9nGCwYHJExdhI2ASs7X5HF1OvP42NcHTHrNBIJWRkxejvDreLRR+mXe2RmwUTCIwFJ3dqgJWWuXH
YOXhJj59MUZ3nKcPujmcSS2vF6wKynv2bDhFQLUD9ngerTQmsz8ITBmkiTE32OHSJryxm7DO0rED
EW/3e/yjCFOmC7zhJ96LmQhuqNgob46LvSkU5s9UGrIG3vTuzJlPbTwKReMyFm2DBmKxAzBgGuxG
VJ8Mj3bfB799pVbM4VM+ObXgmQJyKWZQaFK+EH/g36+2sRft7VXKfXpykFXR9ABlm+3lv/up9BTW
Y2o3mtMM6NDwWci7rVOVHqgfhOC2t5IT2xLMxCsX/pWzO/X/ASOdA5EYKqh3nSNvBfw0rbqk7tT2
wI54uwfwaor1Bytfv2OvA1GD/1WpvwL/x3USBMzbgqkwo2cvT4E5Xb9TvCib+OOPgZvP2v0LPSTs
LmM1utjASxZwnPGelFYVnQ4SAHMCIHXQDuH9qhqp5BgevJEMremTnF27ARhopinVjEZoUcPvcIwP
Xr+Mfl6eVe3WcrcMdfgIt4/5aKmI1NOsQHRIYgOevNan3c3S+flUeCMAM9BXCGhj2YDghVZNdwUW
IeCcpbEOVeUaf8IG9VY6tXUtTArLyECt6c3m9xMOh4tZnBWuqLgFIQGs7BXJ64KXEQZX9A3qkQ7L
Rp3wKGkLTu+NL0p0JraAH72GNfYlUsUrxfm6m4GV2Zad8WiSF9FGmVj8OxOB/6zfq/vm5TG2DaxT
oRYyn0YkrURDO/p6AJSHtO4VdYG5sFFsk7aWwuNNDDXnakipNzPwJR4Bcdv011EYm1qYkzpFswTb
Rorv4qrF+aqXAp8zqkXIz6ASs8ZUG4stkAS+XcKmsyvfcJYYBuTvZpSZ2ucWMcSwaAmI7/HgV+Ue
D4TdxSUwX4tzlEWp/aI30JSgjwIGDyfOXlOBHv8BaQ5tvg1KHQL1SHZIKKS5g7s85d07xo5C6nKy
xlVeU97/36AMwQV5o/kCqD/0GO/9bmH35tWGVvi1IEV54J8tpd+NGOzXt5Sezo0EXO74gjU12o4I
3eEsMP+8XbMmId9yAEIWDwRU7EzfXzjwUyoYRzXD3qUBEg4p7UrHWFbfLe4iamHm6NIG5sVPt61y
QMqezr/5s6239GA1/BI/KzuRDHHS2LO3hjDqMJYqTBZca5hOvJgreWvIWbUi2PbP1Zq74kd/TsgW
vx1xW7tz8l3Giix9NIWxITjmySFelLqeXvIOMIkC3qY78vITtRmj/oa7sujxLGRy1RIpyDQrw6mw
OXk8gOvHmulSvnoPbDWC3OFM29MYQslfe1XeDmufdu+9+3dSeofygUssTq0jtglBPqhkxEiAYobv
kj/I1O0gN/SxTEUmMA7FpfJP6CrR68WiCaaFMQ0Z/Zr1gydFUf67VB4BLEGNCA+SI3czo0lls4KC
gxpYZmEzE4xD3+Y4Dk2ROl3yeqZwyX0Ms1PTyzLzwdXxjCbhZdxO6HTMeANpFnNZtmsvnPn5AJ5k
82M8g81tbpteJU7hOCoVjWrrl8ytF2RlEzwSuHM0JTsxxoE5zrICKreaI8Pdn0a0i8bCbMNxkjPT
j5kgbj2O77I33VJ9YBqmWTrcZ1NmvBcYAQWtsSCHtXhT3K5X00yyT+XGm2JUqS7YscctQLyrBB4c
cHphPHHpL/EgntWU5UchXSyb3z85Ljd4nao5RbcxtFnO/I2AHP2o8kDYDHaPXLxoia1XPSUng/kf
Hkhr6po0Ig8+8LY972QOW4lUNHpoart5r5aNHhPeznwTYjlUQTwffIreA4syWuNj302cuke9Iije
pXYOwSKIJPCAIZZlRxSfJ93lDiqjpOli3yx4VVteCttaFo2mjhDd0QjWcGOlCK2e2F26HfNsrVx3
o6FRCa5J/kUuDNmXYiShdgbuH6attRXG19+FuyAqi818N58JTy9CtngAIRRxcWpFnmZWdO0JsoWO
7ncTBBWyhWuWe/GCojZpv9+yOuXerkVzF1VavxGrKiBNuuSs7zPZGiDsJIrkAq6IOI+/NMYP1Gvo
t4MuFtvcaeIr4s9fGRLYYJ6l/LNlXCGiy+7UJMqY063lcR0Ni/+bzN+nvQJw9t6WIaTdxCGapjdp
DBgSFBo6MBC+Nmu9pD0hYw0kA8C4+0NKKwBvvUd2g92wrv4Xijf8tifNWNeIWgeYPIcK6d9aG9O2
zDPtIetb1gl8Nw3UJQvyu9L8wZOa8HmDqqGtc5XCeHktSMgEEbOxxygJ7Yk2h/2FPquYtiKyDlMx
VJP7HGGnIC4LMxQwHvGUhLjdXwNjV1wHwHDPh2qKf171JgzJJNElTPuC0XqM/dY+VaXTqGLkPLO8
tGqSis3PO7haRoj2bRyf/3tsrrfqXtAekS1l5euYjQi2WO0b0UzVT5DuXWM8RR4aKmO2f26+VtEa
luAfIDFQEMwl9qLCbKSFG4c/NR6K6ADXAV6RBGoo6Rj3XPVgW4dQ9hZ8Ykefn+GA5ERupnLamX5Q
ThuzU3+G8601qJASP/yf4Yn1hJwbAzNrbxjNg6zD607RTrJs8Hnv2sjzYGrzYY85GnI7I3lqKVXU
PUPr3JeL73H/tqFJWYV8ox/L5ICACtAuijNCpm+fJ9IAeLi3G9ICYe3FrHnYqqNpQ8EVUVJPOqDk
fLleLpkBxSqREKeA+P44tHUDO6EcD+As5M7obRYgPJQL8ejmLaRThXyYGdEdihhKuP3ixUQ63Bdt
Tjr+RHbwbng/Z7dNyGPaaCuMsm7uRooXmYd+xof66WmWCHYp5QY3u6oil7+3ofesSeq+EgYi0/P1
RHJ2xhg24Sztsgpy00kQ8H+ztCHNJOcRbeWk+7uSUHNEnbm7oUqDvRK0HRdGZvly/epe6Eae+E7X
7awaM5SNEQUhz4NjCRmYDAbHDa9rkhtfNFt/uqwMaEvqT5I7qWTbcltH1TD5qaGHdiUB9ZLJdCvs
Jer3uOSWzGK/spuV92cGazU7uy4GMvpTA2P2Eqntk+PojGaBjLHnuhXXAD6nUS16Z0HxYHDznvwe
FCPKwIksjcwKcYH3LV1PmYs1C0bYH7tFRAge+XwIDrIQEbu7wpz7+mLxRpNXn62ZqzaZXEDuJhHt
hD4v2LPkgVTgbt0f0EegWH3V9HbAxrpRUsbsFYV3LXlkZxao5H+ob3Dx9GkKLFQAXcP5ugPM676K
/ydHau+byul1q/pbywGN1behbWfB6NF6e26E+QQPjl0EArFU17PLFgRHWMobKrNi33L87Xabwd/m
QmbpacbI8K+0bDiyHFnkuuOghc+JPBtyNeXVTWwBIAug+dzfG4JdcQFkM3pnlserVHaFswd9QDrx
Z2A3YArDLCU7o3FqcNtMuX7dyLLHEQ80yPH5C6ZesKkChqjMpltxkRaWpmUKmpdB9ar66dardF7I
BaS4jgH1FI8QBxmUmZd6C6spav+0F/Gry1Le43AbNhuzbwFIivGwcS5dwM669q79vDTxVjmGBgCv
BLHKQOeiFREgwF9ltiFT00PrNTlDkWgUvSeBiQpuEDofvx9cWAmydlKZvt1EPeIZbTWWGf9us9ac
A58SjA/NpVbcEUNQ/DElPipaAcRRxG2tXKGsPBlR2PtnvWp5QkU8zWfLRxRw9LYEYzMkAnKelfSR
GGvD7l4Vtj+hjWQ3jbN/tQdzrk++nHWri07fg1521jh+0198ooWNBhBnCm8r9erA7P1BGbPwSXAf
IbYrDivofgNvOUxkyAKJGL4q36IdCh0SuzPig3DplmBGdhFFPQapAVLkOsHZ8vvhaBxzyU9uCflA
8auucssAjbBPJ3sQM3JLEwkNeCcP/NL4uV0lwbwr0Kom524ciEiVs8wC7gSh0lOHV3AbnCEv73P+
rNxYuiPDNgigKwtvyqpwtqtlXfNA9n3JwavJgpPRmlYbuyonqFE7xRASwhp3U2Yeb4hiOCRf7Qw3
hzzopd8mwPZGhYnvfkCi3t4pzos3+igSc7JENJrVaJXeGNwk47hy7/sQtDYs85yr4kKf20IDXYO7
+haB0J6W3N/nOtQpJBNanuZ30KOVEg/ou5KLEnuSqbbXota7J2fBETIlZAbIy0JbtzjLaxX5X53u
vxe35UXBufNWsiBrqn3Cd9bLmkgogzHpahs1OFV/0DFyToxcvXssdJTz0JcUF1NNNmBlqZbdBlSq
cDaM8jjHErTGj58it0rzEPfcNIFvpZ84KOqJBBoZAGYFya3b2lsddfb07eiiRRcJScXMH4n1KpVZ
QXDZ1FfNfBZY4B4C1jmUbGVVA41q3/QJqZHmtE6FRJN68YhZbloOKlzEeTSoNHLs+ssrCrVUVUGC
mJ9ljyOZgnPCdWt6S0Rb7zXebzeBzr4oC/oj5aet5ke/wcQev2MaEjYrhBk00D5XqkyhfPhr0uKn
JHY3V4xqhDdwI8apAdMsTZzfGgl96AUIT8uDZgvI1+s5rz1v8+D2bETiu+9HFJzVt+MVLSsHqBXY
KOZQAT86B45r27gGEeJbafVfpMFQ6jZ08AW8O4KFEMCN3+S+21TWrPnoANryTlvVYD2FchKHGb1W
11ARWiY2EQh9ALNbDqES9kAnhqSh5VO/Z4tqzpAUxRF/23ujr3yey6veE69SZKKFFGUbzMa8gzvy
VfJxvaSlQJNP7UKAbvG69YIdYVfnVlI7wOMdYhmz8wpAm6qRdv3Y/YBubPpGYTz/QqJpShAcjfgm
ev10oKEWW4b+SOjNdd0n8fFwuapj38PStX9BTC7tpQNYw52v/ODzU3GNCSywKmxgewsrTFxZCo2K
lSqs4GCj6hfFlQhXuotQ750JOm0xEcrZfTI0+JmQRO/TcmT6shpdH79THWSW/clewIthaafy95ub
tqlIoRkkqt5/yr4iYR/1wU9KIUnX01dP4DU5Aa/okOwqBLuzA5H+2YgPq/31YlEFpelaiGwza3hb
Tj1SuiVemdKn04fkLZY2/Cjbnc08wNxTkPJBQzNFbGosI/UUPk2sads5Yw5hodgJrD7fEKokPsuy
ID8W8JeFyatuTUpsTMR+YysJY7JFhNSTbxNTXzQ/1wgXhnrkqkWcNxMY52VYBbw2Px7HAgqZsFKz
+7HNNZVNqnse6BvELZbuIcTJtqb/hlR9OpmgKKohgp0ywbRQtouY3Efe8u1IZyoEnT0dmyhvhpIf
4lTjpjVsb3TjQ2yEAZshCSwLAYnx6Yk+z7UXV/dJuhqKIjfcjZRmVh4UXOVzB/AHVWDBBu1d0Kyk
eIt6G5xryxFUw0/MBGazkl9aHfQTsolrH5PdHUglx4UcQdSLHk4mgwtZGoXD49RslfxJkT+cINpm
zF1L1epIux+v6rp7S4KzAPciUmXnRU7tx1o+yW8js3IwX64heu/y6SG/iEgqOaCZvkYDQo2dVFsM
ZvRP/K9JWwUvV4MXOknvzb/poK+B5c9SoMw0i/nIC1QZS+z6v9NWKDIFzzq9KEA0B+QTZqn6WukX
qBGjdBqxCbNwRnoLWD0ZVOo6yDX5YIrtbp1BD3dh0pY4NnRC3hINtmbZMcxB42Ydd3nImp08+HO6
/w2w9ZDqOP5viQJ4csJN15EjC4ZgGyMmofsEOt549+d8e4SwuNedvJfZiplei1uqspQKpxmN0gsI
WlAvIIR9LfoIVuwJ/E1sHtPaQtRYyZxnsYLtf8j8EZ8W/ixy+0Rh6DY6zzb7KKlXeEkWAuM3bxu3
NuVrFX2ZyCIJa3y8N5RTB/5iSte2juZC1iwf1s2bLh8LNXIm6PAxjVlT5UOfzpLRVaH8ar1t7QhS
S1jOemYXO/8s+h8SAFypQwRTBsQ2vNEjSB+ZM49+hWQwa7fAqf30ep+tK3qRPCLXMkq6zB/B3LGO
joQjMER4zZVZBfBS5ggU3d59T8lZ+IxkMlnLm28jxlCrOcVVS7dUi8RfNwN1Z2UNuSlGF5PmA6d6
E6Qi7b/uze6HkXMIrCHy2io+a9ddTxsUVCpq7VobuctYh0+C8ieeTppmDgM8aJwpS2JnQkDxlUfw
XNNnBpybJHKHT2uqNeS5HpVgrWbp4jgpwAXvYEp5cliNRI94b881fyb5upqa5DbGPF7jOx2+fnCe
cQWnjPBdae3MGlyGd25//hM8rgMGaVq6YtYm425EndxVViH0TNsVlJDBGcJn/7lzaOgl58zeWYww
SoQzjaDqE2T2MLiQ8BGyO/FqmKWikvi+xtUxQLilqlKmGlB7MpDB8H8jS1gm4eJ/jZctY7aqw/JO
h/PNEcxWu9ybVlpE34DlkbrgQBFlMZl0FprulZdtOaSemcPpEFw88cBidw68AIo4K1S2cuIuyzno
stdHa6CDqVIbSzU7qhXExZdjdxzz682zxc9kABk8jk0b+J2hLox2QMqL1sfiYsHHJe2CWcqQAIC0
vhzfKHRkfKfFgmRHH8ww7phNtQfp5LhmZq/jz07k4q5xqvzVUsKTDUspwYm99SNRGo7hNviNWfUn
LFMquZEZwZkzDiL7VW/HCLhO2s+o7GrAEg453OKaP4eRjpdaRS+ZzV0fB4bJD8dmgwXL3RNldZoG
tGwqYwkNql6z72xjwTJQDNCpvYO3yMg+ymDcGgy2zOuAoIQ35tk+IuEMPZ0rHmjZnMes+RXWWS61
fSR2J0+/bQ1YjeTH6UeYzZwQLZ+IlyKiN7ah9ob4vorkpjcZDdwsw50OBJg1Id88apGLAsiqe0of
aeoVUMdwwuVdXoTv1+oT/hMSiXxch6j1ub2CGPirOK+wiOoA8DGOfawwHseaRLXfFJ/Muie9rTsy
tCap9vgZvQuaUBdHCQyH3o/QA2KOVc8L6VcsqUDlAfK7K4tqjKPzXFqkepSjv/BN9yfKaeWjW//K
Oj1PJ0LxXiiLln+ogVatA7IEEs5rKVCtiyunWWuON4lnDgkOtAi9B4oCnHaBC10+96gI7A0HhkUo
mvxV5V8b5ZX4zfRD9QDl9tUno5ERk5DcgKDIvfIBpK60bVnH2WDVCqOOPxjU86kfepGsRXLf0YHG
XMx0Rfz4IMd8mNyXFMOp8u3CF64k+w58H+zya+pRsAFfa+aFCdYxt75oKlN/P9hwHJ7XtEweH4kK
11ft99Qz7JfVozJ2PiaHHNobhMyi2qW6qxo35JHtLn4wGecvG6SYx2odVY9uzkSrf6Si17JxyB91
bsXsy8HiU7fKRu8NkMWpbgLMHGHi5pNZRTY91oHGRGXiH61Ru6UjljLNh5avVClU40vx27hXra/1
1Aiqn2yUqdcgzuFkQoVE5JQqkNtGuyfDtp/jqQhaG43DwjPHyQpNaK3SCPE+uwTa5WzSiMCCftim
/L30skLUSzt/7FxxNGhGJv6TsbTgTZe7k4/yp0ApSzGzL2s2iP4bVeoZm4byvFwDUbsDpEwtHAA2
RgPzBLXezbnLi72BTKdhq3LdnZMAn9cedMzVisnxw/CKQC/TPllvzVz5q3s7DpPvudu8odR3jmVf
TE6ldYd2q8bRwTt3/wreWRWx6wsGV28qjltJ4VtSRi8W0PULnVz1Jliaj0BDZZjO9TINzN5fnxFU
Mw+6tTqyUxgWDtCb8iJzd3xBg+cccVlrd7HIvxOUsuWzKr/x/8ieBhZehhn3znG5dTceltCy96B3
vi0YVil1b5QshJzxKHqbaMo4eOlnNWBdYk3C+LcWuSnz4fWi4UMRrdL1AbskVOe/GPJEcqCfH3CC
qkxtXMBAqHa3gWqvg5ryP9RgBAr0ivJn4KOT768POqsle4QYJ98H0rh/yMFBFJjMOqwLCERfzIKV
4+hLFkPr/vky2F1/vjT8oDLwV0zyOtCXFQzjZ6kuGrUMAsBIFyzWNo2UKO5s5NWmETZtNF4nDyFu
I9PAs9CXqM4DvKRI9sOdyvpTYyoyvmw3Gsvd9r6XiDZMH1f+hPZl9JK9IpUcJlZ8AzleQocVAiHk
GFJbfpL5ybFpSZdQYWQCrX+23z462ouYo9+vjyWzLdch7cp1Q9V0DOoU7m4yY0lLAV5TefeRvF2j
vqbLlh/1d97rP14NpVGi8RoIJvOOy0sBtNS3KGwkqL+JxNqDsm7p88Yut3zH/5ha7TQ16qulFxdW
6+x0CU6j2kfxFtcNLzF+A9nOPoGvOu9rQRhpo5FRqFAWazBD7I9BMPZnxN262g1UorAf0REqVG8a
/nu+qMoYSSo8zaRmVAHWeIciMKlmE4TGFlmMIIZ6f03GHqpmwSHowvPaQZv7gvguO03jOed7KOn/
FMq1eBR8ZFOCdnrrmPativ2F9+J/zkhhlOlIcQYQlN9OGpGObEu8Bg9Bf8MxTlzjSk+Iq6lnj8J4
0NdnBt5hv+W636WYwK3qm1qAhJonBeQTbErOsKABKZihJcAmbXkuH0NiKshYCwOLymQqnwX3AoA4
kJy/j+cwQ3uUg4BkghUIiNfzAqz9tg2tlm5ntK6OjTj1to2SiFg0yQxHRUYGwi8TySSaYwxnc0S5
Xh3yA93/oHzrkt03Rpq8e8t0kxr47buRBgMyovbqay1l4B2SQn127mTu1la66SPreqCac3psYVf+
l4z8bRS2fLy75ZEwIzlqowHhYPQoyK69AqZnA8MrkfHuIB0PmN2Z6iGr1RyaRuj5XWjBTzZjA5iu
79Cof1f/eqIVR4p5xiA5qQ/SYbweezlLuTg6rLXK1BXHsngdf5VocW3tX/0TxkFqsn9B1w3a8GYe
qllurz/cHHCjm81d33vGVhBqkqJFeD6frJ8jbmRElF70nesUwNPgU0ODJPsg/qAypWTTtH5ovwhb
v1ux3+l/1SFD667ZkuJ9hLDJZKjaPoDCeomB7rytwCf75oSm1gCcJKVXJIomhJjT0M+5dfQmR6X/
/mdvIiItTz5bg0ggJc+MEuyH7mjduzowQrVMWADq8sU7QKkFe/ZAe8iozOdrmcdCQ8gOZZHXAyF9
aG0536uA6K7A2rdvmImttpyc8Dbt7pjX74rIZ8Huo5oOudhtuUUMmEAHC+e1v4esLLIaP94GEicU
tW4SsE6cXOWi4gB6df9cAQ9Toi4PA4ScBI8+YoYxIaEIlJhyl/B7a7qXNPcEVZXMXESmDAyNheBP
cZ4ttsLqafAr03wUjnaHBwWh3+lM+t0niIMElwLqMC/9j6aIXe/ZyyKiENYaCWY0+Lom70LgDWIa
o1v2/tUkf+J+fVUl+NowQw/VpBtVizazMjbzo4lFFY/lH3il+ijaK46Glq10MR0xWqvvXBvXqWka
IAhHCTWFlCWG/RWviuWRWCabPGMehPq0qpAwR3TsFbleO0VGiBFJH2AtUd3MwfF3P44ILg4B8FDi
0xG+/YQPs8+xIsWOljYXOmmzNgVyQY9SUtNNm+cyYJTJOPX+XuyFtNoLPbeRyYuoile1bBzzlMTG
I9LFoLBAAhIBCMAybqrxvyw2AX9yhRcqH+3NHvAdlOCjIEEZ1itMDBKcwDhwDRZaokB9bl1wcEVV
h2dUeEOaSeMnNi+GL0pAP0JxtqYMlJTVicN/ZGjZ0u3h9c1j/VhfZRaG4umtNhtpfRTryw2HKKm6
gDku5pkjIZWBIUziAKdRimZLDjno8P8wE5CZpCUyIPN2jWkxZqY/+K3hsl0rqXx7NMCkmEm7r3VF
XWSxEUWgbb3VSd7LUQY7zOrNDrKlRpry3njbwHKl31KGSI8dJUaE3pjnClE3L+JqPoJXq/z/Z2G/
2plrVRKkLk/2E/yvsY6wqRcdD5NNQtMFHovxes0RuO5+fCUbGjysUdes9tKl1p27UNh2ZpwFfrXb
iwUuZvJb1HfDk3ATTFp3BcJ/U9ch6AwerGuV5doFYXrErNZ0ZS2dpZQVhXwwfhczdbuwpkqERzGC
ZMAbI1L1iXRobmaD1Yaic6MOCPyqiT8m9WRjz8p7qKvbdDsmTog65HgChf5BrQeuXc8HL1KJqGAw
p+JN4YaBM69ZqLwERWTqhS5lzI81UkLfgkiS9yJOUEBZhmgfvfLpnn2DT36CW5P3pPUZEUV9ByD8
yajHXYk0t/mruz1GLjB166cU7MhhlxLE9XQmtap5XFj++i7kx0AHH/rEAOtBt6rnpWTkbHSD3Ulo
DO/o22JwHI6XRgSP0oFsMDlsYMMUXylz0FfOcFWaR1B7fKLMAjj6B6j/n7q3xtTCTFuvrFiPDq7T
ofyhuPVElVdTnoOOh5PbJl3S1fm1P+VtXD0Eq7u6Zcoa68Hul057x2sdsAmCMZFpEBx18Hneu0Mt
U1G1EkYPCJJTnzioUJ0zfhinU6kKt9Q3ZUr3lww6OS9JP/W7+IfCOwKvcOBdq5GvxlBIHdWcxMBd
9zs7KNQO0ZMxdngCzco4EyoLQWq0jhL/n2Z4DskTDPRjtujURGivkwXQZATcc2IMHLu2c9gaoP7U
w+qDChCvMFdYAK6CoCjzrmsCvGQkMwB1mhlNSLBgb35XK0rOti+X+H6KbRYLWMyPqufNdd96NEeo
krhqG2w0CVG155xL8iRKpMmvoGxszDOapvYMsZcXSFO37STHxncyFl0US3+XWkTdmiEM1IBx6uza
wDrsV88C93Nbjtx+D6E47TWqoWPy8cl5zoSUxlnpWG6fA+0QXhgGGr4NyMeODmRYBlBKtG8a+mcZ
jSwAuDYf/GS89Pz3YNAcLj2OSg6qaxmEyZQZRJofPuiPsUdOxe/Yx6mmnDVqivOc9SYOlpXbkURb
9iaewtBjKlRaJx+rNTLi/n6fbAGqd/aY0mvGBfyxJW0U67YZh/7G4bs+Nzo7she/50fL7S6KHpM9
aR2QjC4UwFBUlf2ryXWpH0NtTHUFaxBZ0ZSw61cAo52U+3h6jPto6mTlvIIjJ+SNeUZe6UqTU8k8
bF0YJuSg5yRUx29+q1qEoGyfKeFL73UFHvqVrIWX6AQ47wuYwqCgwOfzrHdq6DbHtgTWCMvS1GPu
A9INpf5JeotpaTB9yugLv3c3o/X01pJ/0/khGumOv8AA7ZmmIvZwhAelgjjW4i/4cysYysqJtYVO
HV0ltjzFHhOdu/tvu3faDvWsb9CQ5aeDVopD8Mcms4i+LGi2EWm0dm1aTgUXKIrwa1Ao+tPdvagw
zAvXMccyh8ZvvQ4LuNLLP7TcpsKzxvrwGK7wQ9lB6vNzMm3TEZOiqz3EcWA4V365sxV33tSMvAJM
blbqJi0Bjngpn5DLQqzmvFHOxOJQvAwMiq7q/Os/XLGM+r7KgQxp41DvWX7PsJO7ONWHP0Ne+yJr
kZd3sqD3XIqT8erWt9c9W2M0cpNcnpVG1INUw7MX8BGSEYdJUm5ZGQd5EFhlV4XQQzI1bdgRs/7m
xtUNma3uxYeZJAj2pyy+NC+iupOnxfBcv2qna37fJirsCD813rFLonDrtQUKLrbRiarQ7aMZQdAK
vxw7JoF09iKjZPskXXXkkO0vZC7w4GZ+ZS+kKtxS0LOarpeZNb2P0cEOSbg1+XrS3lvbNOkPcHvn
czgaMjWKn0BY1dm7cfMQPzw++RYHO2KQHAToE6WRXFdpjZ3Qg7E+LoeaR8vvST3nhK4qR0MaPfS+
4kZ/Xxr68MycavV91OHBiiy01gLIPp+twOcIskrPiyYdMXS9PVI7iC+GVyUS0BEIDbU+B+z1EWLf
lN2NTAi92RNZs8guHsWUArIPn6LGXTeZTc7ubifwXoUrjumERk/CD7yvPOZqwawhxp00fxyZAMln
QHpzVPqGQHVrNXGq39Fu62VHuq9WmR4TsYPtk00c2Sx/54+54emqOSsl8rh1rP4GI6GJW/9aSOHA
IKxriVlYS33O9MCTfjwyShFVf7DfJiTsw4Ie5WYIbtvUjBhxDWLX64+kHqmuCo9TTRf/JXH7ZiYb
4bbdhy3wxXT9J46FBDtiLjju6AMYNbVLJm/WumDWnO5w8Y7u2LVURuCYX2m29ocDyPvhDjWrlAYy
2zlmx/V5R2v7hDknV3TiiYbKchTs5hRHdk9/ZVGb/WUNqWuf+WcG70/BAvqftz6/u2GPvywdjzI4
mGMYusC2xWes6vRwGDVEWb1V2T0QbETVeUeUl6c4l4bkKlkbaP6Mz6z9pOwB6gMGMvWt3v34cN5v
/84+j9p1E/Nxw5q1oh0IjGw4EJkpedDgNr5Dy2uSVGg2ZKW+9Zx+y7ZMoPYu/dnwKQlPhNSSQjRZ
7b0eQTZQvupsoFzXD6dQZeGpizn7oQWKPQyyz3ILknizl1cBz8pCzTsAAVqejfwp5UK7Ma9fx7q+
3+IOG/mxBv9d4VbeU0CDpGFrAu0+GfigTp+BktjZ5yR/xYyXfJPxwjdBs3hwO+u8btovy62IkrZW
e3gtCDpsXS0yynvr/ubEuN3njJnL7AEwRvLJ4vSuJ+hrnalZqN3AnfwAojypfFX/3EC3/OMLBSM5
gljzvCJsUfWbaCPy3wyQULcmWhddS2krVSlYj0ruIhNN9F91u8mXQDk/proA422c4i95aSA8MAKa
/dq9iwPqxCmqS7UtJ0Q65kt10RZWf68FSqS7Do9PE4iIm9zaH4XIZzQWYoTZHSNpYpIkQ8QdjVbV
gvYyORSs1l011B2HJOqRtedeJ+CRg0BclVUC/Bob8akjcaJnx6g043C29GCs4xFRRl75aWLm9QyZ
bVQGygp8f6udg/HysbC+5RrKgz/qCuiqQmfWoSf6te22G9RGCCvsac7HYMV7h/WLyQ+lxSDEnGKC
0kViFuthXnAAsH/NiWozhWN2mhyk81tMUagViHqjNnL5YQRahIXGSFGh2yJWxwNCxVh/jzzvcWuf
FJYgxgk+DSRfHeCTysLs1Dgx3ea3ytJRcsgeiEWWb+uVQYZbQjljMFbphI4eRgkoq0Y27u9i70BV
9bZvbm8gv7r8MzJJnHpPBS4lgbxIbdJC5qqMQw/x6h0oUlzOaFZpbN+mm5tmNoekqnukXcouwc/q
TqnLzLq6p0EfmNpZ+Hrz3lQWzPeGeUAbjlguW+k68CgRS0/97sDLHCpafYaUHHkudAxXICDJnmtU
i0nPh9/X2vCI7I7c9+OZx7+vkvkugIWZxAQwEIJyKusUQSKTdD9Mth9Z8LErAWXDrgnoo2Pkt9oW
6y6lXBCnOAxliANWRw5K4WRPoZvvU/homPtlcS5M0nFWSHCLkEdhbtoFnVm33jjOXVCnVCRBtzaG
QOwyPdi014EQPmecyddTjF23NIYHY0W4stKHVb5OREAiZKsPGHI5pYo205+Ng8foSrDZqO9G3Wrm
sXw1tw273Z/OOMMhkL+FCIWCNy34zmDvrY5wGmaDVb1UJoOfIs0eyCMouN4P3kufwcldMLDj9QPE
ARoXHm10WlLhP1Pqn/xRp2HvnrSwYvjK6f69TVsG6C3BAfVbVl54IIYZO9VWQ8nK0dQtbb0Kk3ID
ksk70CLWfRwqOlfiNby9Lz4LScmE2d5756XofYJHZ7czsuMID68ETUai9pb5IW7GkJmwQfwHTPXa
mcyysTmZjYKAdRCPr4pARSPrPccHvKhUL34mQNUWGa9RCw5G/XYxcvFAG/DtnH2ydcPVvCJ2fp19
tC3d4d+PBOSY5bEP6XDtWH7IbNJMGMcR/BjELBDIgKpb10tU6sBDmFAJu+RZT1eDWnGXsnluij4P
+gKweHivPNYSqXD4X119oymCqG+XaQIeaJzMi0EVdU6pOR3z/g7KtXnBrOXroVaLWHXjGkZcxnu/
YAlCc9xxI8n3l2etyKcnb4ln/OpN4oe7vHFMnoHLBg2BpdZOR03lT253hYXRHrjPC+X9fkgjXL7O
n1patUc6YF1ILqZUokQFQ/UKdJg1zo19c8FcsRPjWZtgJMYvMKqCQrqLLd4H1BV+7Zuz4HgqkCKT
XhcPJ9A6CSvBhNhQtgOTaYkY+Ra/grxLGXe8xrxWhvFTvCCJbte5GROMlPlJQwm5SYVXT6VDeClH
s//jUXLkK8l0hUCZ5P8sqYMXh2uY2AorkeuwCn8oyFMyr87ntJXl7PgR7N+pyrD12pQGCVThFo/l
EMIzUeUJd51PCWSAfOXOHlvf1ZqyZyS5UPSbBJj5XT2kJU8tAVGXRegHru6MD5f83gF97ScBtI2U
Bj32APVsXuEsml08T8Gv2eYxzNPeNZ0eB4YZFa2jfPCf5FuiGUuEp8cYXD0Fl748eGDhmM6FWd9C
/eSKarJGaJY8ZrpT411mBP1h6vBU/FbnKrzaXmeGe2djXXDfcA34XXmAzMIZqLerHiHPXO5he6Ay
E038k9KsJKVB7VF08RR7gwAc0ves+dMTYHwO+uKKRELYncb/gL4LtAeHnUGhJdHr0CKoA81y6ULn
DLNWeaADE5nJPDthGB8uSf+MwzwdKVcsyJe6P34c/fMbQ43QrpxKnecWnNgXH2a/ObaG/bL6Xq/x
IRPuiG8VyoWvxRL/fWA7+rCztdTrAAarp/IwITx1QIfY3mYt9YsFoelVO6A+THELdE+vXlssR4EU
/gLxQgumMGGr2kDNO1C/LVA3PWXkVf/tkP8p3Zv753Vk9zOLJ0TkLrC7YRmx1JA1XkkeEBzkzk5s
8A8jv6vm8Fj1IIXq+Ms9jyJg8K2aByshE0R2NqAzmrTYj81F5iItZynu89q1XFfchcSpxTceybI4
QZiOdHonj4rPjtdm5BSvbVFBKs8jL+o8UVoOpSNHVFgcGwteZek1gCw/4LvwzBVCJCNvnc6dTTTz
8BFfaCYASHnbVRwNHFeb8Ae4bEP9TPnWUc15xcppPwt1f2dWgq+LgP5OJRrY7rBFViaEqTtCLsxU
iXCXW4r2RITI34X2vFCEZbPwTewqz6lVocZHTHUZu26vFHx0aDCW8N/LFPSEvCAmtC1Fz4j37yNN
7Nt5lzX01ZNvgdBCO4NBRwDQge9LsISqTJYsima8yx4Upqs47J14GHnNWd4GpmcCNenkoL0byieZ
vib2fl1WdH8Dmr+hnJA45GTsxM59/y6PgIz1vLTV/ae8fNnWnr6OwQUmwGmZf/ms8wPN+plsJo5k
TvI0BjJh+KMtupX1FBsOc4VpYWZut4WryxqztzZDDVVaQPCwvTEkt1+T3KVtzGfk02Qzdkgnjs19
jscGBIgvuQsace35rFGQbWcIxZrHR8q9J/+7hq0fljh0ugnEwt41nZ+RspWVnTPy/Cm39zvbj29l
DDSusCu4IikvY1TSQ4zHSVFdozwMXCIzdq/NcF1pAY4yuT9AwFyfQdTMLPrUZt61g2Pz/yY+OYub
kj6wenlsJx/lZXeqwOZ2aTD2AZMyRaWzrFoi/YJgRHMbq52kfb3jgjD1FWQO7pn8sgV4dwsTmNHi
jhJcgMunXmp1Oe1ianQjB8iWowZ1A+w7KfZDPO9mXRYJKiV0yj5ttUGPXPcYV/XQnZdwjq6xvrdk
mv1RBAY/GaKvs/b2J+OavCvMYqFsyBQ2ztIMf6cTFuUAuxj0t41mBhXMgRe6GihlKEv0RCC+uWAD
Zo9Ms97w+W/OFq7nUhhF6EdeSzATV3kxJ4l8KhhTj7anGCsoBuSqtjjxOjicHhGogYk1lW3IwmDU
lrmCbgNk9bddN4KTQjLtjyVlCE2nRU+gdFdHqJ3uc89CDb+LfFB1y+FT6Sg0Sw71nb11Q4IWTWcJ
ce1XA8VHr6KQbM0H9yxZAg6cynI/a7AU7iwfsn6Aopy31p7BkpKpAoFCSnUI/QBMLsxWBTknbHLn
AhEvFobzMYMrlgA3Je8u0i7gQn8W3ksq7R2LbtjfheKpoge8MaK6Y5n8U1sMh8Sn93pMI8Ri3d71
UgmphcSGYoY1hdq4Z/KAufLlntPGczQhaiYneDN0BCJYPnNKb+s5LfjZTDeSf/Sujnpy9ht5zuyB
2hI597Flkptv7EdcHYYp3/xY4bVa/IZrQEL01u1Lq8M4CHxeMdSADCSlftItW4nSYg+nicq6Z/P3
i2IgLL7ki4mtWl8ZkB4H6gYyZNaZmrBEJonIn2i9Ut+aPbmiJDmfLiQwjmBQSsF8xGxVU7NNvx2D
Jafng7MtX7deWu8TZ2r9YiONA8z0TIHfc16pXhn/Dm8QPix08xbf8SHIkUKfaHGb9WYPQ04brwtZ
cUDHWzdHtW/wDRaNGWe8rauBDEIRvLXKAfYZUPtOUIDA/T+j9mseRDFwLodW2/4pFrNNnpnlgc6e
O/sVq+/Xb2Cciw9lpZlwFO+HTjQAtUmWqfk2GWKhxZgHVahk6jM8TPaQlWp693zAOlJQIxCNCaqZ
34T4s3102eViCFlqLZNyhSQuyL3rNEIcjweU6+H3QtLN/52toDCdFJmNf/jZxYFjgIHBB+Rp60AC
DhHUASi2JqwFA6GGmwauPi80lTgWHejfsmsViN7WGPxv75hmFo5a3e1EA002AyFvBJAd2JRn9Rni
uFdhaMzLYcRXWmrskmYVn/S2FtgW8QI0wtjWOCGIWBjlZfUY0FCrnpNKBe65F1VfDPdM9mLr9eU1
u5vd0x1yfEeALDULGoiD3ww8/DoZudDSs6qY5RF2zHmAVdiYX/QVDgKf6HgkAFQSeFH5r2CyI2MP
azVPDzePQ+NRJKtzi49mjNy0uS1R6ZbzzQubBg4v0JUZ/lG76jgFQ6sbe1XhRIliXiwZDFXZStMY
9v5erv+07SfH2kcuYcHUXneLYQwlbl1Dxx6dPXPmUjYu5EYyTeyZJIFm7m1Pyehy16jSj58sBdrY
lATS624/wXB28doeshYyy/CBIe+6KukymOWgjlig2foscF0L45U2kHUKqPA153tTdy4vGwpG8Sui
FfRfP6wasq5JkuDOtMcdLk79eFm8FHm5R5bydQ5913GqS7xVrlNRqXSfLcjdMI8l8lhW7383/MlJ
DN9WJQlB94IAZrruJ5qU+Gt/EvzM96/qRuNlH2bwtwwE9dil5EHRk6JD1vhxPcmCI2q9nQafIYEH
VArNt6BvU68m2S5+3Yo0iK22SpJUDNrF73PkaC86sEB/2CfKPJgnRlmBDxmVTE2v4I5cjhnb0ZIk
sK8+lRtkcfMKLCcu7IttIKBQe0/+a4yEC9itMYmwOyRGfW3yPpw8EsRznIywizKHgtxlQk+kgJpP
QHLPpEeEYaths57n/jTvobHpCfh1nTeNxHUKBbBEI9g51AtuCsJ6i32vqTLXqhD0leVh1OX8Nl5V
dJurEy4HgNK8NqQ7I6vkfBDv7nhSlqDZ+Dn7UNlkTYQ+vrVfApyhKKPI2ixTwAYhVsIaqG//blbg
5f2JP27dtHX9GOg447Pgd0qJ1xF7GNqs8BXl8s5N28KdCjRziVKQ5b3xsJNDxkXqymneTExOEYSV
a+aObrinF7WIOBzb2zEKuT9FCsr+yVPmGEzlu9fJ69ti5RXDBtsECzkFro3//hywyMIYGLgQR76G
JoUZR5oF906+Ux1v4qJkGOGGpjqd7Ym3FK+yKIVzj33ZHAxzbMgMO2bfzWa1E3bpjK40RVB5g387
R+86EfHr8ERNzlaUgDlsugQDH7hahI0qaV139z1ErCZ8DzOHcZ70e+BD5nCS9YzKvgmPxgFe0lSO
ipzX0cCksJc/IYAmoYqtB99H/6WyNzBsb+mDjRnb/7xlwfEAPSbgdBhr117FL4j7brs/V3HGuxrF
s5nluwY9Dtu5NG/19LCfMOI+e+2uHd9AaNw271ki3IjjWo6V/lM3DCqPo67ndW6qtSS+5ClNhoj5
JWhwYyQa0ZvS/RiefNd5ZZs/TaAOICfNbODFTTItVj3h1hJgYTLDeM9XAtVBihDi1cJwQ6bY8dFk
nRkakXbTH3qzIM9moolrFRapv4okSgO1/pUpVSlV0/zdn1sEWkAi4RoiKvg4OhzgpimbYfO7yI4S
/lYt3HnC/TJAMiG8ucmVVYb2Fj/3NZx+8krHZUOHkQqiTPjBXlC85UcZmb+AkMsbZ4WTZDrb1tn+
QXk69MG9sm/2dZYSuv5E/eeuDlKCdQhII5RsA0LTf+bpDFolpBMYGvpU1WP2mFu9ua7DGY553scB
7AI7RBhI5NyqzBdY5FNEBpJr1nn5k6waOE7a02Gjee2GjuDp9/ML9w45z+xWNFpJO+8nz4XhjW4J
eTlduUZVjNE6wUf28Vp7nUMFR8cjoJ8hFQXyevKqhShdwNWW8+GNE0Y02+BPN3H8YYuz7vch1f8y
XlBsHfpugfiLbhTOgcskzpR4G5F8/geLg2tZGNAk98sPz5Ka4WR1uAv5mvgcqXVymz9JMivpUt21
PwxPjz3B91Vee3e3em2IGvi8owTLj/EKEBZ+rvjLKJ2NjE1TwCL6k0afrCxftiOOpGyn3zZe//dk
NP7johd1ttDZHq7VZdqFq3ieUYWtzJCCsXZs/+6YRgUMEssiIo3fDN4NjAqOIsm0/j4paa8ak9Ey
VIevetuQgpg67k2XY3bfOdPLmmife/STmff1ltTEn1BGfph/TIYGs0TlVTOClZrMyb89p2M6W7Gr
2RNHKxOUsjxqTtwHyqLxA+6nVRzFtRFw4ygH0Rvr36TQWLNBdddyNUq1aJeDX06fXBN4ZPQxV4jY
l68ycmLmLSHOuEeV5y0fbxHwe9Y86nKE2mVUxrQ/bRP4+7UObn98t6oakF1jjJYA6MQhMlYy3mnF
zFpdqKnta7B+clVu186nb6G6NN+dJVT7kbLdu562sn0anSMslokY06Sg59JhZgPvnaNUEAYP7Gxm
OqfqfhoLMErbvLwgtMtEndL4vFVa9K0AxktYpJrOrIW87CpbQPOvsweUdjDYlfpi5xHCX86PNOzO
5lKb1qxdeG2KMms0MH1TUMUoW/jOexGXO3OdtfLbPjPGycx57Pd5fQ47XYq6CW4zAGOk+uLz4ke2
gbTX9h98B7A+jA5jjF8yooL76v43sxCWZ0hN0fdXU2U/V2AMJc0Qtlkme1Yxj+yUTmfguVRG31Zd
ILIEUXWQtU0cQWmEQcfCXU/ngxozdRaX5FGjz5tdVbIxBFgDAKQ7Eje4UIlT2u0COv02tVlFZdPp
HjFWP5NIEggqEYn9vaDITuq+Pnxd+sJV27zZvcmSeU6jqGYBC2rhJ0LybsgB8d6IheEigf2amvOa
RsuD+cQ12ny+RgAnIcGbd0Q4DH0wL7vv7jP4t8m5KxZMBa8Yqm0dB5GGm6nC1TXG39++pM0B7I8F
UMKUa2RSLSX5z0viKxglKbmWfjAHN1PlyAc2doFhw5FPuJve+wGmgFvrwjhxzixB8RU1N10ks3Az
TSM7wtpf4MYHhhGlHJQh0vXOv4ihsuLrYpngmGyk61e/bcVBBlV5WjUAIQhuVfDdvRlBWd3qvGtl
xR2Vp8p7R60Fwbkuj4SDq2D0kdXawhPI4QYkQVvfKN0i+yEGBOopfFEn16GyzKaXyvHhsOu/7klY
Ih8+S6fNJnIMSL1jyg9I6XJHjPEx3MrS3pa2gwLogpQBJpu0kkEtjCc8ocbESEArKEL7cyQswcYS
q/ormRKAPmP4gIN6/E+SBjVk6lYXc7Na+ZuzWUU7QtDAN2r6ZnhoyLgi64P5MWnHshzl42R7n7cK
xYu9Y726YlmnUGwakrR5sURmLTMAeh/im6wxTXS/+8xg+w+ryxDuvw+ulU2txD0ics45vzex+JrL
i9Rk76WyKrWeNlnSdH14YopT9xMafm9gwzH6IIe4x5ihmzEMOAyc4iAPP4F4mdeL53c65nctqYHv
Rx2mV4/FHP0yasBNwB8QE0YIWMNLzqEckeavmDP+RP1tPiW+LO2IYVPg+gPd4Jg4kclOgVcDSmJZ
iyO8xs8eGaeFQgyy9HDOvvQxdcTTCARCGB3y8m+AKe7VD5dJRTjTfFr4oEArhjT411B6yBwtnIz4
JhXGDm2+ypBo09aFZYWoB5SabhtyU9F5PFiEjtWjRfrwa2j3LSrTJyKDhK4RVrKnZRKRVBT3LY3y
EYW8NaQJB3tejUOyOk5B1rSyh4OUGKMqvF9c5LUJY7GTXPIbHKQeSyGjpVI1Qr2AdI7L0JrgOx13
yQK7d+tEYzNRSHh4CLQsTuEas5KTAQbkSKjFrhmz6T0HlWBktR53GpQ9rQRKACty2Yd4B83QPtKr
5rxAMTD7wSvayt7fpVmTs2JYVQDmYsDjXNYBj/2WDNzr9axKYsc5hxsVxIHvTHE/p1V6JDYDnuDd
13nESmcOjbSQI6JW7e4+HCKOCWf17th9Un9l0t+lNeyb8d6nz6jzLGEVoSPX1Ps59GVxyvliGCIX
bRF0UReTRd5/QQyPkW+3dcycGfY3tmnQJqU8aFzdGS5AFiTcjRJON9jdPcJtLM/X6uDNpwl6yWIM
Ecw1OttlSXExLQSRYRlXiTMC65RNwieD+X0kpwPXbadS0/IZhBJ6mU8UthZG7lJhKXyr/mXohS++
7WE8CgNFjjkdMe44xy3/MWfimjZB3OWqxh7T+myfPAD2Y+Ap0/bwTH673EQVO84L7twRH/j0P07X
RDVEWuSTCHhZEh0tBI26b1vfIKj3zl2Mv9seSUI+T7iIsmPaiSnM7gA+eD7742NDJNX5511z/bof
XTiHRcTJrE9105KGq12XBM/vZpEIBMZKNqGpnhh9/iW3KamsUD1kXOaHN8j7q9x1wmbAC92SdH3J
Sa2PoC1m615EVzhfN4dkoA2DjIdQsoYvBEEse2sZ0avHl5lAL8g/8IQtsQpVUPcA3lnHFsuCFYN7
zVAfl9JxhIbju98hfjlPI0imNKUuPoWkM/5FeCT/MhWVGmxUXW4CT90NAdqEwCjG1Zd7Hr9ga0z3
QIzcSMUTA99TDOkHM1W8VmbyeZKgsCAglKoNCHIxvba00VXyQTxCGtKIqfEJntyNRuDQXmsQ45B/
T7Oc4yk5I5ItjQuEi9+3XMofb/o91Q78NeHJprhkQpxiFmJ7BTXXd//CB+JzWuq3KTqODEahMCXT
YjyvT+qasWo9fzC/qkGix87DssbrFynvj0PGBM5VheTP5MSqTWWFanckaN62Fh5YkznW66W2n92S
6Wj0b5A52lQwYom0KSTddNNDc29eZfTVFK4456/3OR2I92RcIssKtk7tw+ljn5Y28cJDxjwju1SR
MbTQkAF7pYMryC950LH9Bki9FXciu37AcoKG1O+74ZBQmfz+wkJpMjYAPKapbgn/9rB1yMmR538v
wnCkIP8w87+0WcBK49RetEM/vAM9aA4CZMit3et4xYt+xWFR5yxVj1SGvgtcTQ5o5kZmjhAg87YP
D861RM0WCWce8vna+ltxM5aH7BKvDwE7KsqSMj4zG225RJ3ixgUC2sV9RSfW3Ts/71HUZ7iQKUgq
Otc7C/7lU1WMbz5rE1xz9eHWiboA/I3u7a5v6kbZZFba+cKUhaY3hn1RzxVoh8GLUGguqrhs40r5
q/iOkBUOIr7yhtSFq/DqIZw6DmTn3BiFeXS8+OAMN8tBR2rfAzqrCdIkPQiHGtxzfqD3NKvPn4/3
pWzJuZ4MbCcpN2SNzHkI303714QE8//FPHoYJrXnDskH2nrl09sWMgOmnJITB1BOQePRryzfhCAL
l86ww+es/LA6ITW/26jgIvyQw/KezeopwtHgWW4PND+1BK3n8agP0cLwK9sb2rd+ow+szPvkMj8Y
2TuNbe/NR/HiMOKgCfWsB1wg/lvuvhHTmg5Hyn9svllzesUjLeXY8ymUrtczFM9Wc2fr86HJubUE
MQ1nQZCZmIaTBzcNMJwlvy/mb77zwyvGoRf3wDIIABVz8+ZUzoW9MWH8ctvbRvMSZIQr3i51C0BN
y4RFNdEzBGpwbASVGhN+BrlQYPVdIYId0faBCaI6CzshU+KZgwUkHie11v3aiQoMFIc9DHNsdZE6
PH5MrPmj4is5X+8+ztpNR33kqyLKCJE5dIF3DIjBpWqkqlotVnGi0uCyFkbf4YdWDylOf5XsoQ0g
d6yB+ZOS6pPn1yRQQ/6Xzjg2PuQoxbyoQ/rD+lder2wDa5590rm6GXVvZEgRjc0hqwYSlAecbm0p
AHp0RIv2y+jd6GKmCxbejG4T8jgBmISYSJp1DevNXOCztN6snewQh6/b9hP+lDSW1jTNJCdr65Ns
NULLo+h7yWLXQcaSyaYUKhPWARsWP+MnaLO2DXR3DeZdLbT7Q3/n98m0xJzZiDCvTpFwZ0l1wfwP
hVrOmjDDF2QF2/8IiijOMgk/mxNazMa6yg3CFihb6tspT4N0pYUgsIk0nNN9WeBY2nYzFA7Zydx3
KsJCW/ISAViX9MyNTB/aCefyJEagOOwJj1tPTiJ++Pfk3fGRUcrMARxMx8PS/3dNI1YA4RPkiDAf
BPWK0MUPIKjVIPzNSzu3lILxxRXks/yJQX5OKDxI31MWGO3AgA72QyqzoKunpVYUyvDL59B0GarR
gKjpZo/R3DoKn6IWM5nAJ0GtmA0SL0VwpMl5gtPwEV9HjCJfHcKK98kEoc4csBKIh/+nX8NtH/Nj
KVQintwTVES4ZjOiMfKK+whP4ECOf72Ufzuv0VZr/l9NjuP5flDyCoauKqyQcZOzqZDv//HWsqQU
K8peqYMPyfMiZ74tSEFsLfsqsOgPtq2FXonXBEWtdH2U9D7W2dv6TAbnVAc1efKWTg8bJV1rlXf3
7Njs83HWBoK4whPVKkxyTPDMeacu2kCrcAiDGRdcH/OMFn6G8AoFktoEeLnHA5JEMUwqOFuwFeoP
dlnK4suO360Zm8ApL6/wslFcUFS6eVQp/hvMiTjldfKpA5IyzByaf1oEdXFbGvXlt2JmT9rnUu8e
4TD0M4Pd+Hy5aF+8rshXjRT+f9IajDWk/R8rsjkZHEW0FC5G+90PXMfSoqZWrB/daCOraBITa6pi
GlLp+PaoIUs5yp7fiTh920pPpoR64lEVcp/xIkMnv2k4Yx45YFmtEkST9Wp8yT3dm2AvcPs2BBcz
1AAhlpaXVZv4m+LCQJL4I5LTObHIdsk5XX7Uzyz6H7aEhJEXvgPxKJwMrkw7QIehJM3zchNzKUsu
4jGbZ4xFcOH3i+BOhY36h1DXg4dXU12sC0JJfAWigWYqCMf82d1Nt3vQPP/gZwJ4W3NCB3t85V52
++sup8LvBNT+LwNOhnUC+d86xh4pHak3rEojOoPRctoyNxDc+FnAKl3txnM+Utlt571rWY5pTHFu
5dOwA8f1sdaclwM60Fykyqu/dg5MWC5hPINaEf/FcLssyFHrNAa7TDU8/mvWGztxAQxVV/RDVrJ4
xSn7fmKbY2iKSedkLsBTKsZm0N9y2D7hHCyOsmSguhd9xDk5Trg9jTmzWdwJu8cgGeJliTJIwMnS
42LOETNlqdEplMQ6WdjhRiqGYAvnCzPjDUZBztuyN31nU+4R9Y5ta+/GWmy6Pv8EVQwpd34bpvT/
Xlc6rLAOd/Sm6CQgESOD4DPFEnTAm0fSPhquDDEUyrOCpHW6EkeaZtRWSv0AnXHBf6OCmVR4JbL9
FcdxXT4sb1KJ4zFUhwCHdO1CflwXa3TVfoDyybZJmd++aC6WYheigQ9xgydJOgD7/R2/qvh5PcXR
KgChaVZVcxILZhC9QanV6H66Az7rCJJDy87OzsNblkoN8/xSo33u/cs2KcDXHCisyCc7DtTW7Pdh
Z/4LkWmQlT1jaqglUvxFjyF4LJHeDSXrxjqrAhLagq632askFc78rwLrBqtAHz/mOpqUQdTOSjk6
cZEpsukFH6ZwVSdeS7PoFJ3vVr3xfkruRSwnY2EBhhhHq2KPI4NUL3AY1wOpcJtKpmIaifcJrRbT
T639VnCskGmxd+rUe6MFKjt7fuNAwWUu4RGYpJocACHZ6mxd60i/hCPoUNCjt6X2pRyeN80fFv/e
yG2DLjieAqsMAlwj/mjExLVijDZPiqMHDtdnYerS60UGdGNDNoPnczVUsQ50NHd29THI2WcxsIIT
wR56hIe0ejTDsIRe/ikYvgyvdF2rpzn9AOqHOYXUxYjk4G7qC+ikELyfwj16gYELfE2qYOODp9fR
thD2CErfWchHiMUWoVTuit4zEWaLidOme4jrb0xjOJE5vERLnPdPHlxDQncdgBln7Blk/WGBCGP6
DnrvlTR0fWfftHJzFOrYm+omgku9it+rCadamPIeOpe/pah+eW3JKeWGC0t/5yLHAiWsV50S/VR0
y+fN1hmjBUDQh5LoRgMQ47Ojdh+mnySPsOEVI8MFqGXgnWbhugHIsPv5DUhu+g67JUlIZv8HSKgQ
vXadfflAn1BCOa8GXSXoGJrInRXvgrZvjZvc+C36WdnTs9BxBaUJhtyEcYmkT6M0Y34oc4CUV4v/
h/fnOf8N74tZiW+3VrX1TB3cOM9LwJgT+UDxevWsq8+gV1RSpAdMdzcTKLogjd/KLOS/gW/6f97V
QrTb5AYCay01MiRRrcN16HUInO4B2vF1XVcThurswwCpPFcy+5OsK/f8GQFmL8dEQ0P8fSu4Ud65
R6aoYu5lvC8EAmKTRurTUm0cA4L0U7CYbVaAy+9hrnFidmgmwrkhYzYJYI+RNcZ9QCsH+GevqJt1
jlOq3TCGO87Fxx18h6MnTi1Tb5ZOVIdEM0I5p10tgWlmqs8k2HakWsA0cQenS/6rxeM6VJS8shJY
5PGsnB3GiE8zVXnZYW3zWf0H9yiv2ksogs62cjcASDcHVcJkxQZ/MQrycITIOMPzQn7XDF/+CyWA
SizKXLNASKiq+xh38V75DhMU3tQ81SjP1AdBpJIWJy6jSpAA3Y6OxRAac05+L+q2oY4frxmqAYh7
tOjHbyjjablP2ioCibcgRpnVcznPZdkZLzMK7ztT9MzlBkEHQV3sQSLjxrcAGGI6Sv7FXOhDhAL/
/bk/87tZ3YXE1MxB5r2QNe+D9JdtwMRjJe2bFoh91OkLxC22pd/6/dUJ8eHDuTR5h0ZAoAnTgwjV
smIl3jK7qy+H+oilwJEeo47L0FFSvzM14SBiNmxhqT0vkzIbxNx8GKEehPwGUhAdMAQePqzh9h1c
YycpkP/oDH/wNX0DkcUhM3tk7iV7kEf5fbECRpzQSYh2x+iu8RMm5wBVJxoa3EeXJ9DV0rNjGSWF
/SCWQkbG7rgPmKDrHB88bJBFeUgJii65d5gWfhvkr0Yo6Rh75u8CyQlz7eZg4l19bY0bnpaEO8W7
3wMdoAp/zRRBEOgrQqWKJCwCVCG5A/nV4JPweupZHKNCxSkfFHEYurmURAtOTz7h7ADBgDrHQwZT
ZShKvsYhKeFCiUuKXqgIoD6HQ1IeRPMtKVAjXyHN0STK8iREVs3mUvZnBmk3J9yFFn1Fn22cyV21
rTs1QP0UaEKmNM9Oqp99zP4E15u5qztn89cm2ITP0lH4ngCx2QDt27L37qqCUn+7OQYgBq46FHuc
+TMZmD7FsZf0s7LynR0WKDJTdWwA02FFAxYM0bLqnAtpH5OU/URX6jnMf4vO+oNqrHfS9UUzr5oe
l4BCBftV4MHYatrhcWGfSuQAIJWDsyXATQ+cE8jq71Z7i6sB1rHgP5wnFNLfxWEGtl760RJqb2Au
XYDTc3CZBORGd14axdrO4RTF7XUpFQBZB0FZ41XW3Iu30A3mjNzQ8alE/84NdeP2v+GJZsHRfSux
sA3V7or4FBHMitqrf5ujtJxVj1CTfcAWofS5pMTpX33YUY+UfQqcZ8XR0JtNhQk+Lchl49zeFNdv
vcMZmejeBk3TkYhxK+7Qq/GOGGS8VNHs2JengPFoD4D+uWKJEMoj/yrsAnUUORMkYqRxTWP28W8k
vsrbMfvhx7YPULN/s344Dcu6xFt7uahR5EM+L2PW9tQi1mp5eSoTdvCoIcfJkci35dYO3Hha0XnO
FWbV1VY6ZlzKK+aAHZzUgHv7qMy+xezeKhkq8SdmnTfciFdIwflxcyn+KmVI7c9pT2KqN9e1tZbp
If+2D32C960pCsnSuegzOir52DQFxv3UToq+V2ksioeEAGLLpolHx89oMemvOWJxrNkgopmlXnMT
LrQNMMDJTLDYW7b1eAo5/TYwMtLUvmjeXGvm/ZjzOiw00lDpobtR1jHdb2UwwUF1h6ft4JEtunNZ
Etz4H6iRupmLI0/YTf7tvyyrBueOPj1ZRxmDq9Ev9vs5nhWXas/2HBRxzAxDHO9tToOEx2L6TNWO
RZmt1jcYDdcONqdBNfEjuQrEJjUxjKrvdb96BUsT71M/OiSU5wT5aDh3nOE1Y3U3pzWH4ooprymB
8hhcHq8q3tZOvW6Q+W8UxyyuuAQHk/DFv1NauY2/2o84x2L/dYfViJnbkmoCDZ7Wh1pFJLgZLFXD
8KsL3Fu6i+T3fdBtMN4+vdPha3PkJYl3NI6hSo62a8dRUZjw7m1pXtES5H9ahHips/yg+7LDboE7
2Iq2YKCSwdnGdRLR8ppaMYxjAKz5lXyvP8w05mgchSgJmqXblyGCBmMyBG+Z3E5tyj4LzFEf8ZTv
l319kR9/ZBkeXRTu9m2bVCpHqDhNPdmGlK6v0OQSdD3avi/RkUBnQUTjNtIPO1t3lQZOpY8EQCLa
2/q8Nz8CXirOXhCGIVRIaNxgoS/n7BVjHCd5py7KEUnyRYoyjqfxG+WlqNJbfACbx4gMy1JqAczz
86ImL5K+Ff1/uha1ucZfl5Agt52nw/90AlDv7Gt9Npk9Pb2JnPmYGJt9kWftYz44C30FQIPDC+XR
dvUJDZM7sbb8g0AVLZUugPDhCb9R35Q7Kn98oTVthkLVIcch0+wgUZtMjMEGwUwOLnbyR5/wfETp
29pKsU5c5a5FSXWB+MLQ+7Z7ezsDOTBVU8pGYCvYjw1LaSOUbf4LUnASDIOKdIR2mLO7Kcsee4Mo
xJoukMfGEGjy1b523vXzIlLrSaoTErc7lg/o1LWUHVDYQ/ualNlvovg8jP10VUi9naARmPTZAz0c
qBF/tftXtasZRzbRt+XZyBS3iDrl7gHjs7yO8z8SazP/dFb9C1ydM15B4wbaBdTz3qxlRVRledsQ
/yvXqj7GEGsEBH7193sQq+CSd4B+XjUiRLxlLeY2et9XQaosIl2J1Cv0CjcyBAT8Dw+AsMw3Fc1y
iHb7dbxk5Zz2wcDeZBdS2/ZU4Ef7hoPMlmYLgdo38ivbaRM13/Ly9nuFoY9UY1vmMr7pzDvyTfoi
Qbems2t++sh/uRj6wwY2MochB/kwquPgr8HlTgoZwPUvvMgudFGiED8eZwwQUNpKqt1LhUnTLz/f
bGL8AY26/fmhAw0MxAs33ICbE1XkMzydHqp5BOp77n3x9YTHVaq6ou9m7gXImUofayF/DQ5N+HTG
AE7/IHyMMPktNtuBgDwzSnUGUXyglL05HbiyvCbGm7MQ3nK/Gwl6JijZujDBTT4D222or9tWt8He
tI8sBaTiEMlPO8wY+sj0/YFRU27A/4OKy/eYxWz57jWpVn3pEMMSWHBSTuVLj7cvLf/lQ8G69eTD
wH/WiIOS8FcFsSY7x8/RQkCiawGSxr/F+KYA6hEcLr5KmjTPQu6QERFzZKAtLywOx0G96wfFbwLW
ELW5wqlDn8b3P6AMNbCJrdoXtsQgGhZrIRmeD4/VgeycIFC8DHRk6PLDBslYMVra6w/CXQu0tMGS
OPy2KH8LX/pFnIXVGBFYwVucE27g8rO3A/PQPSDSKO233SrD7KlAggs+8aaGjSqd+g5x0eHCoR9U
JTQ0w0Yo/IW42HpaS8o5Qkahg11fXhlQyIMYm7QXCElgIAumQkq4R8TNm8Lxk96AoC+6rFrPkHH1
ck8g+726T6UiLrojr9hSC54+dAt8EGKC26CjduEVwzzSNwgJf2SuJUALjLzCiwrI9r61VLiOHY0x
sMJK8IyVVBK9zBYjyWAZ673LAip05+YjJ+KG6lpkZOhAFfqeOV2O7B0PExuVe9As0KFjwxt3JYFu
qqJjO9ml4HZOgHPiCve5ERT3F3Jarq+edR03jnb1g3H/Fse8NZGN6OQPx86aCCbmsHe1lphgBQGi
6D8CWTlTpKFmCz4pFViFb/wddFZnpRn99/y74SQA2Lzwts5a6atgDQXJ8sYE9iFhn8lcXLhnxrpf
ueZhlt0BxLQE+AFFvt4uCozMr5DhxTAfkXcrKhIm6aZo9Sf8OHpc64jPxtZBsXK6Cr8UbhLfvUOi
V8xoZUS49dnD3WHvLA7erlpRR8SGNqV4+YgUd2gMwma7VTcGwlYLU3oBRdMMwEyiG31d3cctcoOE
mz9vvNqTarra6/ozUq4qho7VWJBBrOQX6qQx/WhuMLSzcqrePGbEDvNDW1l3BMGMuxCBdmUzAk8+
pcGUL7ZzanX2vmbYWLNsf5EG91LkM3+BzUU74HBCgkE/DZobwkNd1PvlPnBRfCS8hG8ZGq/A/U16
2DX6b07wUEBDKbkigdLq8eodSJYYY/O6ZeFtNn7BEy80KAK09KlwBZmtE/625A09P3mqEFxq3+U+
orO2AU0+A33ylicCz9n1iWpfIQieHeTDV0MQ5Rw7R4Ee5TrQTT5mzFW06QLEJgDStbY6tS78BqXw
XUa8rhyXnhdLRxOSUu+v13wGqemMjwsmGWuZjK9KSy6l0PU+gCAk91e0hoECAfEbVcR1WjLzHNqM
tm4fFkM8LbPVFJVP16IfJaGCCC6tgLCAz0mk3iH0obJia1hA/Z1iBfJDG/fMSHG3S8ZJ3snWqgAe
c0mAqAcQRDxl+dta6wSG2yNmiPZnxxuML1+ncI1x1uXyXiSd3Z7Hc+Etv2p5eXDBPnNYXwziI3pw
uMsPmYw3akBTo7Ya6pLme39ADkAC2ZUIkuvL7ym1HUtZbpYv/2kHXkQpq4OJ01vDNPAT70QHUktA
Nr3GtEnglWDmROCzG3VNdYkUwlrofjpFa781HUT9JyIC6qDeM7HoBblWuO+iDU31d4tT72XxjSEV
aY6EKPin3qa2nEK86jTnRjvpR6oAXI1uSjmcbA/NHpsvDVVkp04zoPH+on9wsmflC1TZk0r5vjuY
O0Coy/yjwrWFoVb3jOfCw8qt9R9si0JKgfgbOJUN3ir0Ia7zsHUWf47JavtTFYcNpAExlqbCFrHY
goDaJzTBAR1fvFIinayDXK+YfgiFBe0wOrhFG9fOEo9hv6r0QcbXuXB/TebRfqRcbSVpo2cdRk1P
ChE1onWl610HSqhWnW82tQff3jR/WwrxWa6lEzMDTgHIFcCDQLakSsJDN6JtL1E+wzUiI8aRi+dK
8bdIpio5AQ6K0ItD3kOQTZ125W37PcPG2WS+zN7VWFmLLjoPm5UEqlVj7qgI4nCR3/syYak6O0S2
cJgQLgj1ssb0EUcH6Rd4NO9p50b6bYf/zfT1DUxMzw74CliZHV0z09Ofc/DJ80ShxjR2GTH8VR7X
0dAb4tOz0iAJxTojNenrN4zt2bo53rq/aYJKwoS3AdjtAootJyGlsOr/s6950nVKLORc/EtQ9XMT
AT8hR2w+syUDR582YJDUNcXvtYThUPsnKjqHyITpv2bVZu3RUutkNlDAjBcwRCdBUJcuqnl8tQXu
zDjw9PrxszYLEw3PUQsQ3HVhe8vWMAuKMHOuJ2097IhzlZtSPU61YF74FFNaoy0pApw+zVqVdsNo
Obv8I7q0ROjUEtsoOQcxZ/XLVWglSWaZFKTo49ssbfCvzMr7I5R92e0ILYWXutwNRdO+74rxrEoj
NmepD/flHXI3m5VHX2usW+A0LqGi2yuLcwlynKU9uadPdQyJC66S+6hqpn9xgOogOCjBODapS05J
kqaxgUA7DQGReyJp4lEgzu0KNpmP9MuhYoo+OXtyZ1OPeT8xaCxaJ3dRtxeu9WMJVeMbg1YQ+6e/
AWRAP/KtTG0S8BlmqiP5f00OUufRfUsVOuX2t4W7u3jtlLOSpjiydp3okD4Sj42B4/Xp+XTNdIz/
N51S2o59+S/dIVPuouXPVK3/TSzjzbfc5k2pbZaMtqkoJDvAMgczUqsIqSlCrWbBGMLT90W2HhdM
lUf3VqiKA5GpdSSxMn8sTuIP6pu9gFvnMSTASHJklHl9oL8D+NHHk75wfoeqe7opFQ5Au9SE/NS7
WJb7KiZa8D33ci4hYrJZwlIL5Q2J4Y3tVVlNdQ3I9Epd+8vJoHItf4OalCih2rNOWPeVNfR+5l3H
ArAjAaRUbK4BI+4sbz/46s3n0CxKnPnxaIO7FRuBGi3KF7uPVMDkwKO6NGsy5bv5DqOxS+Gp9JI9
5XDxQSUJ7gMNghLkfLEZ69EdGM77zDjHaOyBIjyNy3BrWbZwLMg5bt9/TPfDlqH1asguSbZFswWB
abzExHjMFbp0nq5YLEpsdT+jziLlI3rkfOGHlMfGPN5s68u2VhRtRSHg35iUZZp3QL93OkntLhj2
tOc4XsWW+jV4lGpi+dA9F31xOukUhTpvMUEhwiIWlZsXhcq72Z3UIalxlUMQSr93BQSkagm81JXm
oNs4ykWg96PspZJj15jj2JbYQ4dYYXfzlCikqq3wXGcWysnvlK1l9Z0IYiZJtco1htuonXre0MYD
XTauHYLTk6F7HCTMufjZF1/VtPCUS33TLx7m6YFb+rGFpYYuRLbjHu3z+x+VI62UUPQ45pT0uHeH
lktN75NkqULnzS7rFqKcIhko2WAyK4s6JKmvmBAPU+oZAb4JDoV8KmFtfiemvdmNvZcGetMLbW9V
esCRJlHpCD6AlQ4tyiwFWJGUiKxqIFLTomlOJhgUx0u7wjP0/H6xy6Ak0clbzQVp+8SzSvyWYy+9
wyfwnHgaIbUZ34QVBL9potIYaqfxbdp9jJJVdS8Y2yJnRQe4klXVahmqJzPqqMxDxkJbmQvkXhjJ
eTwVMzbr3ocErdtMQ4YZWNM+6GQYPxxfGIUtuf5ABmgUnnWClLSJIJre+LxKN26U2VhPS9MMG8ZC
GEBgzCVcZKwF//eMt/jQ5GGXOSsSPx8Kg4jawIp27lgZ3Bl6T/InLnCxLQUIWlg0gEmzy5M19KoL
1TSm94qHSuaRlNQqJVavNon8BQpfkGI+GA7dHRB4m1htwMt28pAAyJNAjas+5Qc1J6Ma8noFPxgr
YRW6UB1lnXOYnnez1qMVA0sOaYG05hkS0jmhyk8phaeVE977kOMqsZYRV6Yi6+Iwa/VkVn8FYI7v
qnkc4iNbcgaz9wTxVPNTbUXYnS1kiZv/hcGibN4io1NDg0FmS5AcKxNWlsAsh7ZPKfB94D+oc/zR
XTWTscxHVOvExkhKi7TBvtT5jSol57jWVvhqO+1kz8kY9qxbu6oso2yk/GbX3y7bO15ydbTn5Xgd
Kihq+gqe3l0rolVShxQEMg9gr7sMO/u6yFGMEG5ctWkK/0NaVdXJsswH+oxw4dsUX2S6fAHKIXlL
wzvnHCdFzVSoI9gcJGWInAkqMcTw9+3RExO7dz+sUPm7XyVCCmc56ENFkFQ33wcRNQMUNhjQ73gB
KKelf7gL4bauodl6nqsKuIxQ+vsujc7ahVLea2W94qi/YxTew9rjIsqrYIjRBcMxjuJ3Tosn7Wv9
84WWEETF1PvvcXQaVuSi3YeK3By/tNlGMBu7VL6DV1DcTLUetLcKqHwlOrt5xsr901K8/gL2/3Oc
Wj0tXqq4vdHfWQkpAR2g3jauBYGBG7cilIeuSWzmAtQK8Kfwnrle70Ymq4UXSWWWTH6smGoB+nzn
kb0N6zeKzwY7ftZadFAAruw6euX1/uKX0U9R+kfD7Ew0CkPNmbQAXl39SclMtFXHnihiwiPW+oK9
n8wCR/A5lK5JqqkXOscJO9hFXni7Z4D6pS/zdxRR03faH091usIiYQ9jGmqMwXQ7XVJbnPicNMTP
xUvZtGVlCYOpyra+M3mEADwyNH/CM0+NCCMpDn6GAMBzfXFOC57eO+zy51lFQtE4/VxnImyxYPpY
SpfZcsT6ONi81qE14NHMYQjrqIJLkgQDx+PYLyNotRzJBdBPjnwUljUvvfT8H9sOgtOKq5/OjhOA
h7PZyj+5W9LfRkEdt3+PijGxUPlDOH2aZmcvE2KUwjn8kim+9FMtfdWM/OQ66YNDOGb8oABs4lyO
mKKDPxKxC9VFrNYSv4zMX5RWR5ShTCc/Q1rwXrMbmIhhj+3Aasp3AFtsceSplTduQtjNmCEHn2tW
Hjtq2Yrn/SC1a8rX2X632N3mxEA4EaCW03PtvdTpYHZBw2p/eCQIhaBqfeBuwv7Xn61ULNKoIbuJ
PskbI5RX0E5YOBZ49XKqXsHcdmshC/zQGAelkYgMoXhUYeL9TCkClu6WXQKWbCiHld1cjQGFq2e9
sgzs2P3Ax+xKXqp9sWphBnzAvkieMNbSu3h6qsNTCTpNovF6zijDlaDiL/awBOkZiE4q93pqEuUC
BUk2/qgNQLyKIGKIaIfGOZujN6TbYVeqhipcmWfrJuwee7y7hWUblysH5qpgqFUuB8DHpWFZWxXu
Hzmd1rvJI7jnEGJGGZnTw5a9ZFdWkiNDcVxFoCGSVPX3zpsxrDEHYLMtFkR10zKT2hRZSpN/sHJE
QzLYVxJZdz2t09/WS+EqwYWcqHiBNxa8bug8ZuXvjS6swTmUZUFO+M5lecoMk+tz3//jNKiCi862
9lESO7vm1Z/8rgfo6QMgClFKfltoTfBJX8Fzx1MpY8PtWefWIQAS9aZkfdKbcZYsx6L2ViNj9LmI
b/A8bmT1+SvTZ1ucgnIYC/3yU6LSc7eoNTnr9H1KJlLDlJnJn/6PphMMhR50YEx1t37NQ1IWA8gW
R/uPrlRqYL7rLUteVFkx5SHpRwp3rMaPW7ZIrBya9poonQ3T1PWPPLSDi8549ApMNpJL0VoARfFP
SVRotDP2pX9YWMpFnUPCCe64JU5KCdYJSygqdp8M4aokvOJXbJoawT2uGCenM8MaSkFJA1T6YBj6
4r/3HHAfFbeFdGcQX/TEbyIr5bOLMvaQzRmZUqi/ZbxrtVfptwg0KMFWCVGyI59okxEZ16wRwSwG
LbYIkXSXg1389FL5RmkP4RPHcyK5IIFJIxaPXY7cIS1hHAABQiyYW3F7PehE0wfC8JBGDEGj+Hiq
ayr/jFpxRn1BIXKzWWT9UvmulY9VT8WN7pVdBGp4lnlNQ5R4Y3dJTbfYOo7KpzgNjntm3Kq3S9rA
PyFnNr5CNdTZ1b07yi6pnIC1aAw3x4XACkiC974uJMbmNSE5dhVQzw3UQ5UHF0ReuDhUp+XhMvGW
XOuqLilhBpN0ftBTcx+JygVgI0Z0InID6278WwvlOCgf8NJoA/tcO+gwKNyD8EEzTSsNZq/I7ucA
NUmWituKoPnwG7Dx+4UxAa408iBmKERpbtxz/1xRu/zhY//Kr2uFKHwFAipTN8xYHX+TMuy2YBM2
OmOnxZjul0oi3vZQbdJHiMTIDMyRBGwjRN+c9Wf0xZnZFE0fgqiBBtg//shcsxVlv6XtFqL9IzBJ
7LIvTna4qLWnwOVbvpzAtm1co/GIcNfPfNQCb1h1bskY/wbLmoyWzHFEniyM0uyETVrnvKew5hoq
WXlUFU7q3zcxJFk9BC3LWdTKYrKoWNpemPCqs/36usKBWFkSjO+yMPJ57/DBCV9Du+IzFcbr7rpr
sCpvtJJtX5xE9Y7jMTDva6bRFXtN47Q2X1IXJHeC8zwelm/koPsl5mBRU60IXiJ5iE42yZvx/02w
f1Z0K30Gn4fbFhNJQvKHLTRo+scLDvBK1ohiiM4AaMwU4GB9F+oQV18NBzkh56CIPByb+rEF/5QF
VAtz1LFBUhbAT4lxkaGLFYBxSXq4UnlNVFcyN3ymIAknPJWOM+YHjvrkUxWnNlgnJ3M2PWheRKzJ
UVHNvFqOIIT1ZbvgiVPu88Y7yOZiOagATbrHea6vlwYC6w/u17LRAX4azOn0AtiDw4B+gPW1VhqD
2OeIExXIf3xDtSyhVz2viNz0NULMBIIeE4Q2r4Qg2mqwXN5Nx4z2RGHj0xTpIQbmHnjEEhQg4UyU
pSNuZ+uVmq8sSCcrpHV727eeMO0jPZ/EaVXRxR0u0cGBIf+KSjMQQUo2z5peKaVuf6fuFIDpPyLL
eSfydtlSnChlnWmTaFwn/LVl/qk92t07CRlIYVrdSXOAfIvz3YpphPiNwoGw7o7QzvcQ6QosSSD/
I2DCtZ9sfKvN9freXi5HlEPdCFrkddOxKpQ5fJ5+ZJ8QruwXwA4GfFvckdlohs2bJt/hpc8VZp/W
UbHscAL732LqKrX/HqPRHqr6PcSHahEM5+w+TODq8Jw/R8rRNOPhIwMvF/uhdw7FcseytxrSSmJ4
e48tGroN3b0udNvh+8Fs8OV/ABrTJ5XGr1R0VM+nGaJS6dMMid3xerOVHEt3B4ZO94fUXKJC2ZGr
dm2tvHgOXIxtgSyNt8i5QJ63KcasBY+DIeWMUKEh1wBZJ+zIE76fKt6/Q65eACJiQUShZKNollIg
LV+LXpoIW1yrtbAG77HmIMxZvwy8iIDTtHqjMaiwGiSJHAjvFSwxcM/owDeWBF7hcJykP1ujUX07
XkUYCvsFsDvVqSjwTUT2s0ucbX0RmPmw7zmk9W0I95A4FmwXmams5attv5lJ7G+lKeJogt9RTCcm
weEE13ruGifqUIy+VlPRqdhrhS9CC+jIWW6oLXx4U1kzWKmZA4oooalDd3dQKwlHveQtq5az2lKa
n64mXP+xgcwTVBJqTSdbj/tB620vWknxSO63+4YdPtdOoXz5GYCN2ECDifen3kzj89JPM+6sJvYD
f9HxmphH6vJPOwzcSYSgYcnxsHt1Y+omCk++Lnwv8h2iDzBOJJ4xOlVqoM+P3UZ1Oqe8z8+Tx630
rCgLXo+sfiz6hDFrGtkqJuGv0bNm+MMPTCHBN3Y7zU6obyUboGElmPMIxTjEF8zMOzkz7pR3NMg1
GzwixkipbnZsbx6YelF/H2qDYCtPotx3EjmwyM+iwxmMCxTPFue9r9CxT7tZLFHqjqYf5gR3Tk87
4fWx8zZxxSqgGD6yhKFhR3EbyLalRCPWuUcx7659uM7ZGcSPpcKhwdQWSqFak6uWElILY2PgSuVR
3ChItTg8kys78bSwuJRSHR8YVw+pvGJv2Eiofjo1a9TiEAtBo7f/2LH6N2CSiQVeF5fBGrDxkNSe
X9xg935xjuQsujiO32AkL6bngDsxAMafssx+YD7WOFl64IjBOeEE/zcezulfkedzfY70m4ncmHtm
xiXsnFnimEEsdInAt7r7WQDkLD3i6ZonjhFf1QNBkKtBQoBo79F4WjCsRcd/fwgxh2AgBzWMVRK2
BRfDHDb9uMTbrTrsHfw0l7fJ3fcYOx7AejWxDfBEzsAOfshrzrCA0hZsPm2fkp5piySNUJBZ/xlU
fcLCY1qGdKDLfWeDMxtzVsuNuARVBRyi794zbgD7peiJqKc0rcLVZdAbtfeVwnZZHnmn/Z/+m6zt
0cOMu28oLqIIqbbXQf93KhtwtXhsDCFUtGZH0Z5xB9dkw+qIQEgBhHFKhgeENbM6obFE/sxGmoI9
TZxoev4j8br2+JegTPl1QXK0p0mizV3CJ8mCsXDZ+O2rA0XFcLcen5uO6OVh3IbaqYm+DKZnavOj
e90JTL3/USEazG9tk9r1XEVxJChTw8IWSG7yzujI4bxfE81E0naZOzXEqQJuUjHiesSbJiTuobgl
gio8zE49QvpB3Iu/JPgohxnHv5zj7GKXaPughUAUiGQvFepr5IcpiRI7Pj2uMYfZIydWpPhrF3aY
EhGV2It0dVGndAAjdCYagrPKKiENU3tz8BKMDVBq3v66LYSo40yOvEt/ohvIoMW/ZQS7s4B6DNzK
22Ad6keIwNi1k9gQlnY2yfgw3wsmOdoNFx4gkQq+349R2qi914oTbcwoj4eaBeSnE+l3BQ3HjMj+
i6UAr1zYo4oZ05kJnfZWAwy4zpEtloFrBPsncwJ18unstJCNvOtiwuP709npu+5qidhlX0Lm6bPK
8a+Ig5EjKwkNbjmfRPFwCLlCyFe7I5mLcd7LSjCpDVmtIvQPF7CeNEl0EYGjgW93UwV20NxFzyCy
yJpzh81X7Zokgw7ej3MT29Dps2uo1ux/h9d41wYFROPjCYmeDbUAMvCTexJvoiLGBpZQ3Fg6Opfv
H9hD/Xnp+mNFQCJtxlq4ZQ98RWXAqWYFrdEVG4aijQL4jrgYLPBr8nUr3JUhEg2W1cFHNu74YXaA
RP9wELNYUl9BQ/5BAIK8rp0EXVd2Fl2VdAuxRGNTSI7UES/rahWHxhadIanidR87MYJ6N8ODzR43
ohEfq3pUNog1FSQelahCnAuyffglwmMQplNb5DymLkBervLg2BvJl/6hEwwkvkSptlLsCvr6/JoU
CO0qAoHW/o96DHJyHM0kVO1eZ9sbSN9c6l1W2DRQ1okb1ICKnqrhHMWCiEWFe6w9CIn8dLC+8gS7
DhAh+PLXHRfLYo6tyHxfhemodNAk/P1K6hoWL/YJdVEAFz8wagIJAqrNPeKAo2N9rqqOD3rq/tzN
3tNFY3s0RaHr++I7Qx16iGQMHSvZDGC4OMkoIoMk/1Sxe4z7ed/2gb2j9Y//ppmcx05cR1L0O3aa
eNkWKrZTF83OQTlZfcmKalahtvFUpbItn0tR/6iOoIoqjlElxk48R0rXUUszKFUxeDRxDFVUkPEL
7Ks31uDwWmJqnlZuHMHLqmCgAJH5/rFpIEXEZqLmZUolaEpTvrOjdQ8u1NHj/Pbtin2beRmGr1z4
dSURfWHpHe4JkC+jgWwDilc3XhgBwOsEwbarG4FHGmE1L/LZ8OBGh5/+2JfN2888KDRmHdw+aQx+
5O7oT1xAqvrUoXHqPJOYgVpPPXymrSL3qkUCSgwEe/7GxC0whyuzJOSXFEPoriw45L78aIaocTkh
hHNQfL3nfRi+XXRhPUPr3vq4vEgqRjDmFHUeI2yE77hER94M8scHAi8zFR3GfOx3/StCJgNwEMke
TEWH/Zaxvh6ZEB3r0gS/EYaaKrLKx3pemBLhZzOwAqKfdLEYpv9ooC2Tk5uYqUPjXS4rGeT249Uz
nBLAeW/vQO21c1lj12HF6AwPTNuqCiiAlZiRJihi7WFB6yLnlRpmOQjdedvYhgPSue4UZnSyY1G3
LoSkv0HURcKj/+4z0j+phuCDb8qNpGmho3h2ygWekVlRQu9U8q5tIUx/C3NKdhgjpryAtZmY4+Ve
boK4i1Kd/E/aYbYpi9OVRSfbq7DAbCuTY+k0c4RoG8NIZZPnZqm4i8oryNdk6/9yVYtNjvbOYASI
8yhLscNCF2BHu3VQxH/mgNnRbU6plM8jyURgchKngSTFUzLO8HsHDDDcxCjBxV6ekixDgjmmcGik
CzzuGV6yaGFu3anYAK3Vhnr478z7NMCePBMzkZzizf6zno2MO7pQDnpgxG5nJ8bQs145JbXO3Pee
DaXtdjuByo9spjt4OLJGBglxalbP6nV3K5u6Kcg6hCoT80gPSVm/HCIVgCF3aZWJai5AjGMFQUUC
rly8URj8vkPgwEqPW04gYPj5IBuT0QzA+fIjaSQWUGeJ/+OCMTp0bsx52xFO6y5w1rGmdd1D4Msa
B+BrjBqrxLnpYHolxDhdp/ONkvBBU8NudYAmXVEjwXyQFnYWZnMHIXttgnWH7w3JZn2iv2sjzA9p
kQFmW9sakj2ur6ocZww79XxS0c+9CPX0bZg6uDltqS8Rw5kbR2aMjtt9hRkzBVwMx//EDSVt0ygx
Fsz/gmxsTSUFOAkiK5tc8QeSafvKNJHRp8raUiC6UzPy/LrgbIrJvxLZHueZmVs33BApOVOBpLqE
dW6WK+q9rpN5gn5ahjrHcC5pvH6hVuogzSHtYZ4ZI8hBDYBrSx3B5ozhu6pco/htpqLX3VHKUf/g
iz1abBVnNelqwsN4i7Kj6oV9GA+hbocyJbkPG8l48afTAuhpbqEHka9z2YG5tB18C78z+mw61o+W
w3pF4BegQUVS+ccaeFJJlKaxcsJZx1UXSEnFSz5k5OEUqP/mjoWwKr4WFKB8q/3jCbQR5w78i53N
A1tFUHugVgf87Eh3bYVSfpeyfexGcaratYXYv/MZImfcZaWs9ZXErzS+Z6KAP7jx/LD59wdRSgq9
ufxWX/HT0PjRp9jomFh2Zpze/9eoWYUCTeFUc37hBfrPeFHwEvixJQvaoCEygUOZ0bVULCIr+Tbr
OeqHYhfZM4iEGRCq/uhfIsBg1jYIUvPp/pBxlH4gbjsbI00jrrhS8Qg/2TsfPO+tKM5pvWnOckLY
1qw8mWNFovwcKWrAHiLTmZhfgQEPj3xZ5WY/WbRbI5nrBlqlcnxjIDKNMfAI7vXDW9vrUKIb9/UB
08VUOyU4DAcaCE2GXflhnnaScRs/sYWBDwj7ps/y1nvIOhr7sMcJMxmUkMH6C7qC8npoJsDvJBfM
LUqMXi2odSzOlwiZJ/1R4DEjt8lrcMp9hykB946Sddw1J4aT9OFbqd0hwbuqbET+lsApBTu1dLj6
dCtWZUpXzHLtqk3D1GnaUJliBz64mJNxjuxN/CW571m+fzfOLvzTzmU0UX9pdQIg+D6GUZpHg/8/
Zgib58ivHYT2RIRSuPq/H+FEyJC4QCjKPoVatjmbPp8bPxSfaKln2JSP0nyV6GpFMl4LCgOExi2H
/aAw1n/Pn9uctAaLIJHHa4LZLnnlqZB8Gg4Ui+ZVA65jK8n2h80779dqVw1AEjiBRTq+YoDqn/dM
g4gjzSqKmUMymbTfd1r5ShbUhR1/J8K8nslCZXFK/rLl2vudw5jgFKTBNuoiImwk4g8aZRdYrD48
n6AFRjSyla8cBE1wXzZpFJoLU80Ys+oh6cd7iF3BvDry7r/q4JnN5WpUZCW6+g8ao8W2SaYnqD1v
jSPG82WwoFzAj3Ot7zM1TVdwd4Ks0KAO+csHX0JuR+Ratz7fJiIzUcTTc1kL+sVUjFqz7gBK6JJD
jyO/U8XqocgYqm1a5eMrLoK2fSTD/FW9+e1FEcoNTNZ5cmXgA4L8S4vgaCu3ey4QZVfYzWdHNH5R
Y2lIesShmEzbOWkHUrk9zqcmGhtCFaSkuOU4+c7TGI4yNUL93YUPHsMAC4kj5XWt3mpsKwjN5Hhj
ZZjyZrDiVs8aR+txKZFu7YStu7zLvmAald1KzjVmscUOrjr5sq7RylCKeOsxhYJaTsBh/MLOO2Vz
tvfs1KZrNe5QwrLrc3DNoKSLurqQScqiEkytLgKqFNZbtvAEM8F6IrdY9ihzBILbLh5U217RTRwq
BK5shJF9jWHIslz+V5AF00G5QvIs+N4mX9yiqsRCuGRTskisqPL6vQk1HK5B0iW+umVxEerjjCIp
jN2ZTOcWh6b5aImi3rLWTrwd2J3JfFKft6r9VcSJbbv9Z6wrbkcTgT/9N9f+myQQJLFsD5DzLpmP
CNQlxoq6y4qgBkYskyKNJ/5VR9+nMwCEMkvapFujd2yQuXXHbXz53nxlgnSx7o0udSKD2S8FTCOv
KKKSZzU/NZzSZIWyEr7/AKjR9/jT73COeFqwDFGkasAojkU/p2NF6QWqrJLcpt6Ms990FbqBsHAG
SPjHFgxZvL5JkiuJeqNjZX74AlGb0vefOr2JLMeQ94wc7aJGsy0NW9/v6XPnNZbNd/VQSurNv4yL
Hmc4kXT1kyCzFPtSsRHUAeHLwYhSoDMSxyTJDe0iCcOAxacUY2dND7kv98EH5JZ41erCIA+aua6K
cJsM8z3LsF5AlnqPFOlmkmPjGFwitV1FofhgDti7t+rxyH53Ytvikuy0yEpCabfr3MZuIQEXpxNG
rlBtn+3hg6gBvd7ophPoPBXm+r1UrYKy1dF7KeFJB8jvYzLv236rdbU/61DUXCM9yVJiyYJOHAls
txBFwXSLp2hIaBP66hkADegZCrAOm+1K4j8MUbiGSbBP1vN8gucKgPdqphl9cLJrZWeJU4iW9ixc
9s0zoQyq96DzbM9FoBBSglsYLTPVy5S/mIiWOJx+832aHVFdny/T+R0LV06aSke5PNZdRa23w94p
5Vb3bCO9/YpnI1sXJ0b2x9Sp9GXpqYHzRHOx2GyB9+H5szidtknp0pLGjUw4wH+Wt3GcMasDzCap
q0mBgPfuochnj8akUe6/NZccTTV4hQ8qw3K/74zDlDE5he6/SE+oTuPmqutvuDJCiAaYKeOPEYAw
AVa8YWnCQomYeJZRX4CgOfGSYqwRKvidPp4mO/gPsmqELr49nUw1kwaYXYp+MVheadaCIrsBI+0K
I8MeokJKWd1y+vpthd0sdPw/I+FS5suE2/Ip9zEZSI+NyeGQjJGR8FRu0X2+k9uroEZv+6Mxx5On
5367voJnvULC8GjteltI6Iudotv422qcB8LfmPeWl96Ajcq0GR8vxdul+MByiyoqZlI+UAOTd8Fv
e6SCJTPSRJdna0yv9FPkCdYMxLsxI+Nm99Hts4xJ6PWnpb5fbrb/fimkk38yQ56weWesriYmeaRq
zc+hIjbXUli/yj61ZFlQuxCaZjaEu1otpVZl+5eRwE2VfrqGqT912FD4osdDPT33KB1oZeR/4xxx
1Vklq0Sjn2Vs762SOgP0rUjuCs1qZPfopAw16ymBGNlOdXE46jCk4l2MpdNuQQwn/w6Fi9W/4jll
MxMTmJSX5oXOgUd5KVpt1od+b804I+hRXxAhJMxkyN4QJeBdtT1HcF1yGXxqqYh3rp2OpfYQROwS
nicbnirgx5vvTtCE7tGrwt1b2FpOmGkBKE4pTOBq8l2bXbhE+RCB/ectEZtPQymnCQAw2iMNG/qi
2Df2VAkAYdYbBZvABAar1a5ZSprIIKomm3zRM6CVXeSElHlpNwUmB09jArbBjVkv6ihRJ3/vDNAA
LM/IXx7OpTMrXp9Y3kOleeDfsYiHBc/RDKkGjY+TNKKwDMqwptb6tb4Xa5Yu60sC1JmI1SFVni14
wNe/dfyfBCQzd/EK8P7yWJnrLxMl9L7dAObrDwbKGa3Q9mtXE5dnfeixpGt4ijZjN3rHKBK3xc6E
enr4oX8pS1VTZnOtzZq8cumyVoRZVLxyu93z2QeNDZ6meE4djFWPUMZpw6RiDs1P3hm2GJ3rUs9m
/dakRmGnFnkihJucHmdxFqKKCdg+Hkp6opwMW9Oq5cjT9CPNH9AKh6OP0mcN3CDvWKeoHmCtSKZR
9j5fuu9VCetRnuS5fHx/TE3caf4XsRScvnoHOem8j0PwMtBZVp9BxnVZQpeT2HDS7wDdsATmVG0J
2SWS/m+lsQVzmURs9j4hpDaTix5tK6Yr08aWbI1a8Rgy71XaH7EUtI4NBDiTp12SB0u3iTpuOAN7
jjjyg5IaRVh1SvlkamY0kaIKLENDSWrarAUqd0krx6RrFEXbmwk7C+uvJBc/nx5TJ42sJeoX/yTe
bzgPoyKqE2xUJm8eHRGuuYokTSmAhR+GEYySqk3ZSc6HjqK8KEDo3JTyGdZZeNImJgNnMZoyTGAM
xrhpbjs1DHo4mc7zYOjOHD49aCVMSf5iSHMP4QGK09XZmvExUJHMTYVbRgIbhtK766EWZMjLRD1V
AIgeFwUcdiYo0UB24XntDwwu+AmqHOwlPmWfFFEcioeHOChJFNNSpWXuIt0omtYi5ij2Ayvz6SMx
ZlbMbJtX2YxtxyPTHLqMG1nTpSihS1onzRkSAnNc0ShbHLcy0g+fw6nOmOM6o7aLruKYrEWZb8t6
/pBW/X5K/GQ8exb0nRX6i8okzgEy1cXRDskwt4gC60LlFWT9tWWLNpgBEFyRIfFkDGaslzc9TcA+
adfBGxRTSIrRxZd3Ex9wQE3g62R7GKhT9LsqQvIg5SsORgFTeJytO7R7FyMpuAQLQhrwlrh8YyNW
+docqJji9i6tLeCx+FoFl6w5F/Iu8Ewm2jAPAKYuXeM29cZGMaGEii2SiAMWp8DL+ibE+mNPGPc7
wVvbf4tSf9OqeSVd6i+udYcCMdhDRunirBDYoCXZ3EpjkjHoI5WzTI7RV6XKcCEoiJAc+gvMjLVH
f5ucl2E3/O7tSyY1g7FeVwetmk70cewO3rH3++VpFcfPpuwqEdQmNvAUNONt0Wxh3vPWV5FrQTYo
Aoe8yZZk8wrEPUL8nrgEXrqJY1N78VybNcTKC3YK7uSed4gRwCxLObgJ7LqCS9ZeFwiZx/m5KB1S
a8EqPbBLeeCeiXlj0EbmmtBoJFFqIoeAxsAF6jge6MzDVTkuVAQ6JPyrHUvkdTmo/hItoK/YMNWn
U9VRc2zLwgVek8dShOFn0s9o4Y/P+QNNVDktlXs6L+oH/9KCiigJCCdbRryT4Tr4exfQK+CxlsXy
o2MrffcoHtDiOFqGAziU3NFkrPAFfwqbXFysjWq9n6e//jysirtP0BF2bBZdz5zvfScQAaNiQjNB
BH+BdIR3oMiqJTNX05c3o9yjoCVKwtNFk9R7kQZCGPwWRQuhTUPaWtW6otBGVpmnvMsFfOD7JVrp
MxA7CwAhwCFO24HJOnkLQIf472dBQG/uTtumGj7o4BzGYEv7FU8KKyZObWzqI/WbtQpXxSwtJT3Z
xgVC42BsQzIG4h/9q67286+2WjGE7SnudGVc2MVRzPQZGSsqR3C7oL9vRSBnLD5yui6GaZ/5YAYm
4q4fOft6dOgn9Hcc0uubZ/yjnvq8G/0j9306+9UERPcfhrtk1DIDAXL4b+bvzYuSB4ct9C8fNAXB
ZzxafOEVnlAJueHl92AH6TQYPQ0lH8UlsK9q9XnWWny1TlHkZ63ieVvj3tRPlLBxiOSjsS5ki1hq
UUmihUwrOGU40/gS7zv2R/0WpOOWOfwE/h2c68HM/yVa0nuYGOttsYQJkUmc0q2U6Fl45WvJtISG
tpTW3m6TbO7ZLGszqNWDhgKFg+IByBExs2/XLl43NRCcvh346TM6wGY0Fop1sBpNXIyI3xPkbJCW
F823GsFcuDXB2rOrHEh6uAVrRrCu7uAt+Rd3BAj3tsNdeLt6ZL8B2vad8j/ujmHMoAp043pmGfff
5sTnZCL0b7cr/kiqiH6zdwC3MHPnEOdCvQA93NIsPGjVzVe1cABYTf0l9TVAZzBhTgHZdFKuI84Y
x8EFD6ft3d8GsMxU5j4a9GxO8fRH3BYoJrPX8CUk4SUZc5wOkR5ajmQ7ey792bTCQWmJkgMYnT1U
hu3aKASt+gtpU/UJgfcbklbgBY2wajIpBxfbvmDUQ7QJDj2hvAjeTOX6vTnBFYM1saJale75FQWg
tkNg1SMfJSuyC6aKR6u0dB9uf6pltLvEdyLPfmYvtPsrtZL+/BmhRSkOVbvOWGJxvKf0zsZMS+5D
jIUyP82cOAvHp6/uSTl2JVohZKzNLC0rLIHCg5NfGwOLw78CfpN+8UDzWJQ8u0hoI9+i4TRJQPSX
Sl56Kxc5kk/oCo+mxKB0JKCy3rhFhk0MCUTxy4SBq0KXnGrP40bOjSRsPjq2OwqLRnAnYVa20yY6
QoJ1SAST6mus5+Qi86zo/21nlCJ95QwNAAvtSrjqZG8aHKhGkgaf30OPUcbCWZ/ZUF9wlpzCgJPP
Zm/Y8/p28ISjlQbPDpVz29wu6DMJrpY/myxCQr65tN9V41Rv70rPI/+b3lzgEKabb+igLaLBlywp
6LM08jEcdCDONpU02c912eYMfPloKdM6zViQPrsV87vOz5Mgu0Cd1uAJG60AzG+qaVe7sY9bdz0G
C0xZWp0sk+1UG60Xcd1pgr9joCFoF/F1dOUZyxxiAjfVVHrE5N8i6Wy9yBW8gdsjKUrZyQlSeRqW
pjEWdoubEs+xExWBdYMoYfiTUy1WmOEfObQnJ3c08aST++wU9zVEtso0MnLJP/audnTl35ekrFOj
zTJF5frWc5OfTCZrOQFqyeBX//ceMIX87FizvgZUjQ0kincf5NyZ37Xx/fyWtq+awDRGwJ1OEIom
XlH7oNlgQSptsBoCZbrIsx7zNpcRT80Ji1s4Ffz4+PSdMIG/0WguH6oHdk5192JfNc6DBLEUsiF7
MfeHQgYp4sw4Th7NVxYwh8o4TSwxyrkMr+O3wjHGSKvpOCkit9a38NSoW55cm4f0lGfIAxZPvc6W
VRbRXYpFEouTrPVUk4ij9aXi/4XBPstTfaJ9TI8bUCkD8O5As1lVXh1/0upiVwEnQJZEim9E2TV6
wahoqbDGpGGYl0lU4fNjki0BMI8kzLcja4lzYa0HWzsOsFPwwz6JQU9JboWvmkxbLnAtEPZ1nbSx
t6Ah7CGXlwFgcbSLp+eNe+06X3Fcu6Ixa4tHwhvEkBLVHMXyDi09hB0KB1YOroolIFMbuZkJd1PT
lRwZOGrthPQpHCcddwhLons1R3IzpNbP89pwUhBEC9/6YDxVJlSdVj7rZUYmQkvIpjq+U8fkROHH
OiQXbsdwufJfx49+vLunepfsxAAdjQKwxKzdnEquFzybWVI2YwMAMSc8ITVof5i3LGq8TduqXfQ/
od5pXOrkUD/cVnhDWXwYrP6+eP0bJf1RNbCc5jzjw2/IHNA4NN1dWMpPY+ZSBuLAwBLmUi5IXpT9
gIgi+F32kb2+UYtlldn0jSKel+kfF3lWmcV0Ckow5qW7l6Xzb+CgUtPl6biOCHe9C7+j+xsk66lt
bXL0wxVHYF3eM+sKO43c9a49lxurcvA3CQ/zNmWGJbbKRVCixnxjzdptlwCMuaicgGAOCRuo1HZ9
EDPIsBmdp3yk1HsXGmvMfP9N+fkd50EsWOH9aQCThGU4+wXYr1uyzuuewn1kHS/x8buWDxvbKPns
kHn9eQWaLRBDMyMY43Cs1wBVsAbK0Q41ckCv3dqMroLieDXsPj7RDDznCXCmLhUICBWrK1AJBSHB
O7pOegc+FpBkcV5LWjTMGye9J2INii5dKf6yOM6WzrKh4WNCiRp701TLWCn8QDbNm9plqaUNdECq
kjziFOcs3nqv8e8snd2gxzkNyZeilu7J6nRLbhmA4exA8kHUKgINW6EvSSr5fo1maw63ZsmP3qcr
NBjPx4opQ627WhdCREaqMKPJWxkBNTrIQs+QCt+nB+wvGlbEoYurK1DG5zBz5FS40hzIV3SH8kkJ
+SoWggKvpxb3Wt3AuH+zXrKUgUWlrAhHSh/dEqyMl1SwgjYQ+u2zjod/80NjHyg7Ll1mqCSmvIO3
fT9Ez1StYMhWoLUO0RgXvzYsSdihaY/cVYSt9YzKKTrBZCATQgqSkmXLlX9HKStt4OUaKRYgLyM2
UFzSyewiDXDQjdPbFKbIwgvhwIRsE1Q7a1Z4xJ6leUo+HpNHwF+TJjxFSXRA0HiuIKVfANTK6EnT
LCC0iKDpZ2s7jR/dcXcxpGxkcW5dFkWP8GIXtEPZQuHuJrSaXl1uAOOrqdoD1f7iR0ON+T/qAI+D
Ce8sstuqp01Kax52tKbwlEcZq00Zu0L8BGyAUDtL0CmXLOUoOv3qk3S6651+8YeDHKNho5dJeIoV
noq3fwCwRMS8K66JiF7HQ6zPV/2Kj6ejWUjTCof7QGGe86HzHzzTvKzP/aY/YBvnFCwkn7pbaoWP
1CyXNLBX2zu1mKSJQ4nurFJGAEihUpQvuo9Ja6FnLY7FzUfyGb1mPWwVdrrUHBxNXjvXB0eMCx/C
IzAukD2q0YJJGGAc3PFVyNWZvZqOQbMK7rbFocLipWMcY7hL8UkTbadpo+RIyAuUH7TQqxG/tVBJ
/2s8l9umeuX3ZK2+KkX1NiJtSAX7Uvqomkv81jS5lrquy8ZtfUquqmn5+8kFUfvYIge7C8VSO5Ir
2Lz/O0X5z+Tsc28oKxe7Fgfde2AjA/OrTo+zH2Fh6L3NUDZU75ImxhS08x4vfqrD4oMUyCKGKmnf
CHTK+78Ls4cENal4xgYXXI6y0nOh+pmMGEwDMntrHCYsN25Nmx/+F8rtdmrUdl7gvqCnEvqNoRTU
bryw0Fgs3Vcla+gI0p89LwPwf8DDlnHoaVFOWPqftGnCWJ6LKrQhP/VLK4mAc77DuRQMaFOPEJBB
A1sOd8YPtwOy50L2KpKCs7dFtuAjGW3TsQ0pMak5raBvPKdxBawpAmGQEG4446Qd7w+KpeNFsCgG
9r9mwf1keMCJpXJb82npaQzZtIkOurl7yyrOHNPE3mW+ZRXlupE9eZ15kds/jkzxWppdcJoPbV/8
Rirj/Mq8lV2ZF0EdwCe1zNXksVxvXe6ZLI2V0PwCjqmzh9oLXpA0VeSpGlDeZpIHRRyjbdly3D9a
kHSIgGBPjrj47Fn6f85F2d64zcHG1Ud7hYP4+ZQoA31jr5zdSPmnj0kkozj2ooCUrsn2Yhn8Nbtt
YD7dljT9kWXd4T051/M9V6rpoUjoaZhkj4TrWfiBi+x2srXxvq9w5rAgWFtGL9fqlTNszUH7PWS7
v8TKCPoOE14YKo6oBjzDVvGwkIfflioJoKfqTe12J5CwoB7L9BG/yMeNmcgDXaj3DFq/NrqIpWG2
dCqUtkOzNc5/VsybdQKx/DAl3erbZ6OO/7IrS0QeI/ANphIPDaNm+bvxBGks43dHc73yCNKZxdHF
V+SOIo9ew6z/pbcl4wtqHkbEbqvt4qB/odY+z72wYYo6s9jYgCmJ5K0FGuQ8Eb4RSAYazsxFf2YL
0WTn9SN8JQu56z5X+8yELzXacE7Td4ltRlM6fEdFoxjjTnIq8T4+hx0EsB6Atp34N84kaxVqHm8c
FaGR9/tsKQzjUN22ssFlYyLteiSlKCZ0tfpFDxzFZa5WPOHgIrLO9/lH1koceEu02bkoSeVWGzAv
N+eYMQHwaIpKECIDTfjSwxEH+91cFrTXFpptvk8P/cdmHep8FC+1L2ABw4vmR7V/Gh3yjUN7MQCw
3Rbnw5h/2U2DCm3r6M022lxzT/yFDCsTFBsUB/1liSl3y+xbta4Ys12HWmrXfksO+oUxqV1/hDyE
pZi+U1kgEujvEkOI748tDzI7oqve1qbcqS2PVhZdB/VRI/rh8EDVqydC02J1Bz+koNzL3JS3vm2/
q0USYtME6eevjAzcA/YZPQY1wnkfYcfiYTf4u2FrrClA639IGoJpb+keFjfNkUOeKzOHKTicgqin
jkej7iPtQvyI+hxrvNec40JUiL+4aojlz0iWDZ6oCSF5E37O9tnvYGKy1xP0E0e8EPPoyqFbqpEb
/LW8ZMz+9l2i2GNoTnzrzZgHgeiv8wMuB1YGNX3iMkGM64OfspWcRiPhII5/0JdcDXrWOpG6/ysX
eO1VSKUoIoN1DwM8lwLnB7oUa8z9X/D/Cm04aPL38cnYtdrJye3Pcyd61Uqzq7r9pxaSJ6mBzXoA
iSTr6pHizcZ4Yc3Q+vF3Npg8+fSBM9p7WFUxiL0PgXSlUkModJE41buMJLixLd0SshUCxha6BxVG
X/MsH0YsXomOwzkyPXwrRe6rVX+8YYRzHpecny7L3pVdoVDP6fY6ticoB09gyJLske2xR3Op/dR4
WKiirWiuELXUOvxFD7sXFnPNPbGj1TAfF8Y2BRDxuE8+0CSEjgxvcNuYmMGaiLcf49H6o6WSsOwB
drXG+enZXgNp2URPcD/FEeTwG2RAD++5gNObGGfACtZUni2UDon5D3dlQh7rOGTZBXGxph4XfGCn
fsL8MvyYVCnPR6cKbsqy/YT9VO0+ZnLD8JHxAq3LPCkAlTv/4nIrpUpnuWw5WxaGxTiJvP4xTWus
Vw/fq9VUh2i9erRtHAT924azh31qBpn1vAMG6IeO2NI7AyDyyHlhe3nFWa9/LtzePFkaoKIRWxei
RiFusHhKuw2pvVgBkNETLOpg2IP5xz/qPpSIm58CYjleD0TGQj2d9yZaV9iTm0lPzDiIUWpDswi3
36qzAPiWKVAi+ADf21E9Gw1b4QK6g+5bVIkGIL93XgRzuDFg3/Zbwj7epSaAc/odm3D1VmdzMh3u
bKS/XEHFHfMBxkLY8KQrxEwqSrDDrmoboniSB1AdoGYDbtS0/9wM0FEjP1J4DyXlIpSv8l3qEeCh
JpWjby66OMgpJuFyuKDZi1R597Wmog9/J8T7vS6M6wxexILqPK2j/mprYR6IgZ45tYLUv7cXSIm6
dzxz8lg8E+jOEBu9ksvk0EydFL/i4q+bV6H8oQt+YjwBdwy5SWa/Y0PXA9QajzOsoqZESrl1Pwaq
vGF8S3qzMkYyPkyHZJh6jLB8Uukt9xghaYfURXyuRiSNIxvqfZ/Bo3/uRYadbdE+Cw9UMYvCBNCF
HzPC9A3VxIdoIloVBHkkwHl/2fPysdkgiJhrfpeWSjhLUOAchenMmXsWxWeZe+5rkWPjxAV/o0OA
gltYxrYUA+nPQoa6xeQxomvP1L1D0ZpG1otEtwpCyeGg/zC8xoo8+UL+9NzxX09Z3dLFB++/Nqhv
gGfUFQS/iMScYRB5QfNl2W2yt7QKb7irL/0GSCi8S5MZ4sBEhaq7NZxOiJJ0bRJqeiDL/n86ymnV
AZo29LgUdTEKoomUTpcBe8Rujp2z+c3GSNy8nsdWWnnIriCR8zGaval4B9SD4t5IPE7yhMf2fSQ1
aZNIGxwPntuvMdHDnH5K1s3b2zcYt9MtBNBBhinEztwgU7cZW3Khc74sqH9rDoFoh0yfzOlqamTT
X321BjCLdIY1Hs7qoztp4IJDflNuecDTZmob4q8UZqvhWeqinAmX2515QsB13wfduo7c47KTgb8j
WvXj8ETq3jr0hFcyyz5iNT+QaKFGLu2+052SMiVmXjNaXfCyJcyWR2AxZsQROgEO/vUw3Tr/eXCy
dMUwdOTYr2r2bJT3ZJYEUcTqWS0ZJCgf0orIqdXro6ivdY/EByrDuXBxbnw6Ws+mBpaXMezDAeRr
cPpYfINSnqxiKQE+cDPLQ4r0V3a6xPlQhzRW1pVzr+eyiXDnRAlIQGquCQI0rVA6yfQ+24QYkkct
PkuZ4gC6XhPtUWjy+WUwTlCh4yqZRBYLqOIpHjDG24FMG4fCc0nqPtZ7TYL4ymA66D3fFNizQDae
wmsMNs4rxGy3zXPJUXiCzRr7yel54tjrld2MZhKRdO5lhKmRr6h9hM1SLFjbpkTbc14KKdfxbP3g
wwQDOwmxPbwbebZpAghHoRktkJvRAffuuP0HQpLpHOxnyaKEN1I0WwNvhx4eSdoMO6gwtV3RHZ3R
4cprUmSOFFMuqzF7CFfLUNoK2UGt/QoFToimuKkOi4C4VCr/orMNg76WbuzgKyqLroeoTXJ20oHi
D7QyxZo1Ebs28gGccF+IVZvJU/T0QgYFRJYGtQ7VgyPermvSNnlQa8TzwrUhvrYWUfcKVApqG/hd
8UDDHWCUpUcSRXLnuoMxbWkt3agrftzOSmrbp2JiZpkFnUYPzGOb48dJmNdB4uN9v32NO9S5ag8W
LXQHCZl8JNl8bL0annxl7fXXHP3HRSuMOZXOYdqvTEwptuNXh8iQrEYSQ+BC3DYTp/noGbi/imq2
bScQm8Q2LdPtNmuFyv5wTtrFBiru8vgfUpNZzcS/5ffbwHbiuH2h5PkhfxhA2Jc1VEmNjdH/FNuQ
6EOPK4T8oCnLBIeU5LH2UyilvHOuam+VKogdOfoNN8is2gmoc0a/gEULg+C5iF8a4o9nxQ90AxCg
zYMMN0nC6O3+6JnbkS8xxQFxDVB9r4Nwl92IkHh1duXOs7NsKXtsNUhcKd6gsWZErDXnGssd0LCP
oh8ptLXY+GrqydWLafYb5QUtWj3dvqr/Uf8I5iVPhQPN+ltXv6tIIcX+2CapVFcUpaaKeMD35hIm
KJScO6jFfwGGsR7CCPYVYrHCJVWCqQr99K0GWNwyKhkDQNYSpYNp404PkUFoGCu4OxojSEvIc5Mk
Z6M9Cbrh2km0xdxoMbhkJuhoPN4WoppUMfSQWPQQckTCr2SnUSGFERswjxDeqM00bPSaghi5ZXS+
d+WUrKxFLfDFWBTJAoCXYxdduHx3ztGg/j2v+ZOGQ0Cz/8+yOxmeVVnWUGMZRYZcRV+qpJ8OL5N5
6hsZLgp0oWB94MN1D6D3ez3TdpIIMuCIcllRQqDPkeiSCb+AJ3pASkjDvDZhW2Oic6bv+sxGDgWU
h6BuCC6OdTFgmRKNTupT40qU47VsYZJIO+7zoy3/5e6tamdswJBILlbWMwaF/r9Rj5G75vxZokOP
7gCHQ6avOfO/e/g+dM7BwbFCKGbZ1BcNxm5Le5zCNcmh43pC6rzWC/Td3nUOKRcK6bcJVOie4hPR
/OWc25V2/6v3BOr1g4KBk9nkbf/NFdejJgccVOANCOYcpsd3cWQuRHmrK38F6jCyjoBsEqIIvK8P
Abc6JRoqvd0lfNeiIlmB0ViXjo+Cr65P00RPivJ3Ybbur8SHYm0lizmLa9eDX5IAbcYUV0ndQY5t
n39bp9kLij9BfZuw23p/z63yYPs8MHtTWfFMsjE5Lbtvi8dbEAt4OEzJSb0ZPzEr75GSsgYh2dxw
oX/5oNChg1nMbZV8Hp5sCdHCITXT3Fi41OcPDv3PpTPDphlVa89Wk69weB4xbzkeDT31nYUYRAF+
tzk5L0QkjjtkvX8ddsrTdCN+dlCwjeGs62mksy3E3aBn5xcAgg7vFwlW5ApehvTuLXeku11vzlH9
JMYdww9SoVJhJ7eKrGfSLgYn5kU9HtHq4qBUNiaA4eUs0mA8gyrA4DsZhPGWgP/YNEvVTBhg8+O2
llS7y35W1FasvwJNDa+VsnyLlHPMOQCcyF35ztSFAfO64M6n4sst1oifyDaS5vMA0kFAWBXyvdey
NTW+OkoW3QqUtbGEZQZgPsMa+KIY+vvUTnn47+M67c5B21OYV6pbDzfZIrw3VU7zh24qFQQ5FPmT
BFK1C0kyoNQFkf0B9ULEuBsUdLhG6sqcXdvGcVdH2y3qWlcyWQPPhaM5XG0MZtA+jwgafyDBpOuS
DVCqJ8UQE1IEgNr1GtZhD9M5IUHyqTeIwdjnRL61FjmCBdxOTqnvqzYgf+X4m2JuGFPOKEfeIcNy
KdR9yOgjmrWkU0Hi/NHdQHFaGP5dCMbeaueoE2RLi8MJwxxszbex8FYYhkr6fZrCX1h0b1wMUnCN
bJvfuOhBSFG2igBn/OxYXdRXd67QHfp56/yeRY4igSFeM3fe5VpQN3WWWRpvkKn4qy7jaODMPoRU
fUhtgPkR3ZYgH34s/NsVLzGR9FdGwR7NuyKl1iDnTzTnSmFEtshAPQldWNXMAVxzI32BLk4wvKkb
NfxZfzpEOAyasjPxbqVfAKfiJMc08Yc3+NBH+itEsAFaN2+ma/b/2kgYusg6IleWU8zjjo1gw6Sg
wMwhH9T16zn2yPni1wZZaOzbOsMRO7L4tkg18y4d2eNgdFw1Ai6lGU2QtYQk/i3EhGLsYF3dSeoH
fyMmdLsSSTts1OGZFqaHlk8kgZ/2ZaKwOhhNM0C4+/PlAgBK0wS+OJSytygww80Fk+piAJlLJU98
Wh3GjPyjdsiLympqjS6yEASjyF42ZUdyyYqBx6gyDKTbJBRTr6pbTJBcdA/+LNN4A3QS6cdQHQsA
Z0zgIPJPMz4uc+8yS5ojWnrFPQnjTgzm12c5tWThfBkRM5iAPwcviCH29hY/ib2P+elJW9GSUBdn
jyuXcfEEIUbnCrC2QY56xY1DEjX7OnUm5g+xCVDVhof0kp9QcUVu3zRWa7WZHSE8bENp2F58iUyI
8WXwCH8KVvHjYqoYHQ4Q0KoNCdf5RcoMuuyJ3QHhSSmOv4aIcgt5XjFb5o05kNz56sALeZ9BLneK
UwBrpgu9UwhUcFt6yfv6YAg4z9O/LvxQNR38gXoSgGwvAgOsQa1AGgx7JcCr92j3RbSrEyh6xqs3
EgBWppVLlO++Wy42jVKexsOGgQgBARdghKeqyZEt25IDBT0mN2yO6zvtN7nLec2+P4rvAk+RBs+M
hNtpdJMp9Un0GGRiem0u3bCh/+Cf/pER1VQpV3k6GJDEr6JR5QEgIHqnv27RqMjru+rEkv6lF1a5
o8WUe7mQTazO2ywYqz3VxNjXdBzTnvi/eVjv9Li60eKqxi4Ia64zpmM/ExZCxrfw4YpHLIjJANzm
lUQ0MSD9E2kdWPxN+NcSNuJWp8z5Ag1BmSGAoAxaLJ+v8IQlDcRYDr4V6X8L5bV7YZKnZAhzDIk0
GcN6W1AheCA2FC2YU4hOmGiGdYUdk9RAvLKhA4g5bq+YEZAbMNJPrpS0djbDXtX92oD/OkQQKcSF
tKsEnBvl0VWxNpn2R3Pij2zD0C6Ch8rxUwv1eQDwZGY06JA8I/JiHAn+ZPPUyPnp4H3+orVGJcQW
1BJiqREKVK7P9CI/P9FRX0jB6ye0u29sh6JZzUMww8u53r+1X4H0BdI0nBwEcbbqN4DDImHjyLTr
+9dlDX2rMD/q0k1zT4p0SY96/Q0TOaEiv/xeZeXcYRqyn3ha+z+jv5gD/d1p36530lEc01YD76SY
kam58dENf7bXLUrstWHWRCzoJSLBEd4bGD917H+kZLWcRraFapcB01qKDseDosuP7vXlFUVrbxhj
P6VQutS97NN4468NGPFO7yRb3v8ESffiWeo8DoDdMdOrO8+Qf2d1nM6SETiq36VvOEGWZJTNyI4R
jSQg1PqyA7HwdRK1VC8DY/+J4UcvAnbZ5nk1H9t2nkJJmLTDHpmNnA9TX/4zqJ5BwYP0M8pOQ8tQ
zH7XitaHYtSvknnSvaGqDLefVCgDESwAUv9yH0HlCBj4QwcII4YhCmsloxqrOm06jl3tIL7puFMW
kPTUxz+7abxfZ/4iwt29vu2e0ZdrEmjlCyTPa5o710B4UQJJu6esErS+W1keq92+PsCVCVfn9lIE
iWYZlwrQqSWUANMz2Fdflcs3EO8pCRxpK2th2QKcb0zrwev5b1+QLStO+VRk6IK+xICUgr9Pgz2D
RIRnTmOn62HpcE6rtuJF42bNQTAzx9cMHYF3ab7nvqkMWtJ0pJnbrgCeYafiaor2DC61F5R0R/uz
Prp/+lQkqbjwz/kICAcUGMQeWLIyXk8hGbTomuVWQi0mdVZP5HE3r7JiAlx4TbnCT+8uVyhssdOL
+q/cvo5SI1UBCdDN2An1q0jExqnV1aQPp2k6OflrahV8CDzeulMm9OI8TBqdDivO5tt6Q8gBw2RS
5CUrZWU4Wojj2SS2vtBSOCvnGWIXS+dMPEitw2LbIVumajzeRFJlz4BzlGD9StrIaK+PORF76ukv
8xPsrRNUwNkaQYCIgtN52GQp+RlUiqVkL+IG2Wso1X7S329IsSpoeneLYf/kQUDf4ZlHy3qGt3XX
tVwYK0QYR6EyuF0Czp6HI2kpD6KUwoiKPvPo9HUcBu5FM1Yl3i/Qi4o/YCZyRCwKHETdnQpvmA08
zqTuTkhQmzBosttBlRsXTO0WFDPVvdu6Gf6TDgYFJ3oR56hZ59nyN3ZUAnXfG1Vo5veuHtX7sNy5
DxWtmg/HFftv8qsfEkSssztcbVsIur+sF9r3tHaQiwETJvOlOiDD+W7s0ruCRforDg5IfQycBakr
gv0iFzoqy2v6a2YvVDVeh+cjDsmUEO6B2vWOAlTPIdMwMGnIhMLFpBuMm43iRwZ6YaR1EulWOJ4k
KB3uERcbsitKngV/FUrEZ5Estg0pqFIY0jfLD1kwvStG9E3fG5Om4uqIT+JZoGuYyd+ttOmVeXul
ZceGlKQgX1TRlC00eV9km6+Lrn8zdXkx7lioka29k5IBSP2Ypkks1/uC57IiDHraSeqUsIE7oT7y
0FKipAG6+HNKmk2wSTskhYQbJT889CcvM2ryw1Ke1v4FjsfA1Haqbz5sSJ5jaDdvmu/zbGZJdGaN
70O5njx3rhY+9rFG9OqKUh5LilkC0Ate4eb+cc/fm7ijbcMOVW74wLXdn/mu7OmFp8HA3/wqiw59
FU28NKXbsM7cs872HerctTKtn0+QRlZIc58d5B1tb1KnqzkDjgxMUrI7I41vSWYeme/fJP3A3cXg
focwPEUGUuF5d5QNjyokfXOqEjtKik1xLFZaRdTsrtgwy7YPoUjsTPvNNdqcZ9nFbd6eZFD9rGwv
DqGcaAtvhg4Oui0DzGFn/k7x4hGJrmCV2qOJiaPwkV7kcleVouvKbsDxn/MAfGHORji69BsS3qmV
dx4/r90vOjqNLYZCO+dZ7YIVq2ncJUl1YNNttuHulDJ1Ie/N8leaFObII6efh2Hec+n6FUqfpvli
2pcVv0IAgemiXLn5sgl4mIIhLiJ0UO7gEh763v5UfOsWtyK1Y1JszNl7GWKPqXK6tIoqZa5lB7UL
0P8pHWyXi6h1PZuLAWu2dOVKPVJ+fzOQrzvjABNxxCV8yuJf6IJKkkfCdWA5GbcZWdpcPg6U8+FB
ZZPYF5lxuwuyC8jE0tmNdVAOmyYWKAP6TEClhki1ilgUyNFJqZPGQkrBoY+22bAnU9wvJlQAnSOY
aKxv6CAYK623Rc3YRmG9+VQb9zimwhHc4ADdkLJapetCoQXoVnNb8m3vZOll5S5aTxQDMzti6+Sx
BMDXYylpTfYzYLjAtsxTC3WxVmhYcpUe+qcpHo/EjS9EC1YMFWbtnUhI6RI4QAmy4XXI8tnHQG9x
NMQLl+6ft/p8/PZiAJlDBTASF02GahngEuYRnLk4+geOhsmte7KBOdAcm87VmWzPZM/FLMV0zQ5n
yJehIeUNFWZy6qN5H1dtn4KeTr8n9R3KVK3iMKADq9/1KihCRKriB3pJgc4EajJa6Yp8paL972RK
1SNXzXS+eDS+Y9ou6IMsTKkmLkdVtKKmRiHWVlTpl9cVxaX0rwiK8Y6DjNimOtZStqzt79TXNIgE
dx1Gf8vr3zZXfzF4WIAVFvh2A61vtyaQyC4VDCwhkzKxUF+0OD3YwrYXuZg/7A2C0VZnjR8vbtJJ
UsF+MgMq9gZt9wVh4o9RV74T+F2RbDKuLNYwlfP6z4Tos2KIMvmjGXBqS95WNLnQi2b5aPCF4L0r
gGJRrx/FZLKMZImggg/hCjItvn4T8sKfpwSfhb6Um+STBWrtLgfF3H/T5zGY1ReU1bX2JED+gm71
s5sj69d2/YUv8TD+KcLJj0IgxoSDWdeSShtKrbsBXEM1CBoscHJZ9we4UlqGh4fEG4+rmUyASP0B
0fTUOS4J6Me1g9L4jfeRO8tqMtn08UdCJNl5lVoiapnEvxCRUv3FeLKropNwVDL+ZeIPM9zQJ3p7
9NTsmDxxW0bis1HYrYd9pwmfbcKMg1N6vkuIKkESm7xp0g8m3CHb/hFxw0wmCdUubs/GPpS62zr4
/S1S2fYJeX/xHMLRmYFLxh6LZ8u3rEDfujSQzeEVGNGnOnndg6h+jqyYAxvOmpA5jFmolwrao5SV
2ktt7k6KvjRMi6BBdDKGJaM9sXRMxXdbEwGMooeQ+2jr58vZXO7kdkRwU5vShRLfeW3xxqjQNsjz
un/2Chdymbis6gsyiRiYGOmwShJtFM1d5YAfNZbQ+Tt+NlLpbjqBegM98b4j9ubQCV53Mo3NZ7lV
MjZTxDyMmyLXoMTRWBGnEsYgPx1xvi2IkSl1ndSJLFfdhEcNX2dI5ClC7VnseQWhMj1etUOIVDbS
7U0dD/MuGXhMyEuq55V8D1LJewJsTRnx+XuIEK/k/06qsTrDEg3Z6anLCh39ViP26yuHVq3egybt
1DehsBlW942OkpWaxAncBq5wK4C9JoZMGCMma8R0eo1bg/v2Z7ztPAEvc+igPY/ApsxUFKPK2/eB
nKO2M+nLpKE10u6iWt8daxxD6S9KGsb69WwCyP5h0Rgb51EXd77ACibNQxh+dYKCs10BlwnUygdM
sKPslVp6fnXTlikTzHFqrEc5jpVoBEJlsgRFc4+iJtCOPAIEPQH7apBzj2bS+CV0Yf1yJ/mr+/4B
4b96g690SvqDiQVMKBw+hzyMgmjRf6wUi99HWr/zrDZKv8Wfb2yhd88Wve3ZoJUsvEtjk13K8joB
DhSCz1EOaHoHmY7HYlPV2pwNqc525Bi2VjrO2zkduY8qgtz0g61ik8r1XV+tuO/XMORqHerBVGD0
AbYPYtuRRtoqVKajXVkwIm7HWi/igxNFtMXae9S/wvqYblX1IWDVZJjjtTzLrGiL38sIhNHgi3Jq
NOUTjuwR2+ys6tDOWrm/bfE/dO34SiFMYI6Hl0hUxTQGv15pak2eWvy5j5UJhhqA1t1GIYI5Tucb
PRa2cgdJoQ15qaO8Q+xIv8FUgduOAWGxVQeHIVdLgKulDyWm+Ot6utBffvWqip1IoUyQ4UUscXN3
FFmvZZRd0TOWIy2kn7rdpf4ea0FsQqPOp6GMlvpbqL7wItYPPzcv9nO6QF9o+YX+tYCJhTuxPvTb
/Xr4omW6m7B1lM2GjHRUO1CaLXx4ehlCAUTHYlf8wYTthaj6pcp+2oEaB+lo02p5ACLHMsBTDCjZ
afhkth1MWfkcG1RmrXPuWAgDi5qI8OiJJ9a4em4QiaFnSMoS9+bWd+ux7z/rVwMfNuDkLcEBzcgE
bGjgWIzpSqfNgm2ynESW5/Ib1/4aA86uYGQ1q6IY6PFcpy5cYMsU8I/SgkzweNiwe/acmXg9MHHA
T+mg5MIgo6X7cjF8FGgu3FWzwHWxsiR05Js2+3pCHMXQcndnvFknSYzAb7lU+hxNSoaLBSN4x4W/
DGW2VuhNsUQ4XJ+mWC476Zup/nSGd7j/RlReTwVr8F6V+omYLxl42I4sJrA+xWpCHUl2EVHs1Ky8
aKumtMxBxYZhbRmv2cSSB5TtUhYo6mqTPGK/6nQ0VAAwNoSMxKIwIZJXzOXFfNUIDKSDKtnHU72e
JNfHw6OzAVBIs1ax/IBYZ9d7Zlx0AXTb8ESFuaCMjNABftkevcpkuqi6UUEvICDnQvpbzAHTnDFR
FimRGI/XZk1kcMzfwqp96FbvXoFE7IV3iy3vTacEtu1Er6l5jcXrYVXDyKRCDLaS3HVJvRw3H2qJ
Us9oTgehTy/p8U3s7z7r07fffpBmz7qyH0oc+AgeunCE4kH3i9d001p7lr3InotNF+33CQYJPFRe
aYBvJgQroUSnjRNPrKf3n8rexIGW/BLbR3HkZiNh3YrcenExGSo6DWqRRAKsEYfeU2g9n6M+SGEs
0H+5hO+W8GwOSNWnNuI7bpU/nXaQEBmdX6GOz0ve7cDUmLDuA92wg14bNCyByPpCMoVS4xpe6V4z
LLs0xQPFhtY+t9Rt03SKTPHGwGD35ayr0D8ak5gI6pIdrj7xMFZeZG1VqE6xDPxJwHVOcjy6lbDG
Bpa37RwkHAS3Ke5XJfmB5F++0UhxkCLfutXrn6hYSJxWsW1i9DBpK1bxH0lDV7HU7XOfLJ+KEYZC
uZ91X0aaCPadSw/zo+o2y46aYUWB1K7W+lYwxyZ+6rbnie/DH7NY6ZJg1/CCJ9uldD5fBhcWHRic
LKDI1V8c2GRqGYO5obkEKEUEl2j6Jp1C0g0rbpOO42aLnC1ENXmbO3+dVlDUkETsF4Bsiu1P7fDe
FQ6mrPGkzQvHGbYA8nGdIb9pYcuMd0qXLiOcWlYPElK/490amSTUu8TXuEsn7kLD4HWCAAYzFuXw
6w8QIdcBz4aBBUJkHdg6kzHlF+tO4pi1qHF8iQgjXeo2SLycPXI6TGZDJCUaisTq7eMLPiP+gu3p
P9vtmiM4Q4PbRDnVCmoh98B63PqG51rv/4SxvKW/s5AkRIiGRRlEDD/0+tgsTK+mZ/a8Qyw8Xdk3
PcLPNPqLpbFL5zuGMF8b7Y+lrrF0C+F3PLTmWG+aVbs/izBDF2xOZdvAFeE4VdL0UNaDTJJNHVu3
B4d//B7qjqNd6psLjcF0Onh/yBsvF5iojq3k5+Dh8jt4/KpcbcrmMKB2pZUqZrv/sP/KF+JuVajj
2jeBR9mDUchvGrZbIwUiSLSAqukvFBMxM+5AcBfZoTiYx3fI5pXIikIzTjz6FRP2SjnWEWEe5rX3
DYCQ09DaIRLc209cXZARIHxPWvsHsk5R9JoQnG22WZ0TVBzID99Xns52WkVg1hl+iEN5K2VtO8KA
qmFPwZa7M1gtegawZ8zcyXqzv2ZP/6JfAWCvjHsR71C8bJ3hmHtD7/aFZjwas0mrZUQ/tpN6LPuN
XUOHj3RnA3WgKOY3pAMTnNq+lXbRvbKoktZetL4UFjNqrdcaOu+pEqYjD9E01Dx1xWPbw5C5ALxO
ADG+UOqgry468X0AD90f7iTSp9Mm+jAMIU9kqNaY5mUkH9p1YWU0+TMPwu7YRY2FPj6gM+mMa24w
khhKSjVncVleTlSf2l0JJgoFfHya+GDNEa4mdbGfyyn8N6Z+Ho1X13b+3m+aX2Z88kGJiTMFVHmL
+vLDxr0OhDPMZlZtK+XyVYTrmPYD864NWqSOAa0iqWOxbMSxsRxHpZsebkbU3DAtX9XHR4ETcu5C
0ftz5D0U0SKGMAuyfm6rN333pGyBHXEftHY1PfBOPY/QEi5ElIo4nxcUnRO2SVWHtsr1ikr4cWpP
d/3wB6sO2LEEFg5O4f+uRYgLv1aV7OyLBgRcs679c3RPYjkm/ll1vvPpkdy0l9pspW+fC1k09V+9
2jGBNE+5bUsP1va+o7HDSC722VewHT2qYLfdaqVbdwnsc8BxPyqRfQQHVpe+Bkt2Nbxm6wn/PL/C
cpyByWn7ZvRaSA1TvSVyO1HXKnVs1l5gcMk2xJ/OEz/EyIGFgnfMS3QMZCaJOZGiXQLBh0KO+PRG
9h8evf+xjDXF/Ek//fihlCqr5+v7wvGYgUIEUGCwMxbzFB+lgrWE42mYe3hqO7aJ3uZOhJMETBt9
nitdHYZ2N0deqL4QoQFzN8KE3WjnnR30voSe/CR4C/RVeffvfDlxpsn+k6Wb/A6bjzfe/8COCSvF
GaLOeqPXDKKyq91s+IF7Kr8wnZH4NMiX9beipup+8SV1utRauPAsglWnaiLX0xEWWq67cUFcUmTY
4L38wYckjXxgrh01Mguf1il9dHomuh37q9DHTQOljvAF5o7fhEaUWC0Yp9rI6EDQ5FhLk1OuQvH4
tNRibKNpNvW9ZGWbpXLvsqmV13U3TUXFwi7FGJIQNMDZ4C8PmFfwetBvGVa1CnZf0D3Fl9p/N/bG
O1xk/tBmgqFAnkzPCCrs0pUNGnXK0gBZ/bz2mwYuonvYU8SO0J2WTA95YuY+15hcnR3T/CcPFN6/
5pXBeFTwz2E1v2xjt4f08ojfhHg0MVAkOpzqgLOw+Fb17FzLPobxk7Qv+W3e4oxfysaYl6fGFl60
VVFtyoHrZ+dQj4p2SwCpLTbelV4GOlslYC0XjRZuzD8XCdjlSQgzUH05uXFMdytS3CUc3hrxqMGw
JEdplE1z4Qy8UlDrnz/UHQwhkKyLz2jT0DuEfZlpzENTd0PQNLOWXf2haNXLbbHgrch1Anyi0P/m
bsHDeiA+HOZ6hxFSsA22mim9SHlwwLaZG2hEirEc8csvcMov7jJPuGxN8RXTqFqSKEvIqZEpnUII
b+HLkGO46T2MYDhH9u6g60+x6U8llu0Oi2bAIlvzLGen9/otFcw9uJIaY2O6mXGfly8FK3pRhVy2
t1HbaHWAtVr057M+AFFQPe0axyie0EttoOwDPJ7W4U+C7WUtk6NoQthmmLbfA/d+WnSr1ToQ/5ij
hKnw181VekS+ZOMbz88FMNGyjN6z/6L0MBXJ8F2uYrdGFq4CwGxJXTRDpoSnfSg/ItzV6xZCd3Xx
JGBn0VI792S74QHL7ErJFgOu7RSpmgHaxzM5qw3+Z13s1+FHxRJUcCMyjHsqA/cSdIXOep9hIt8C
GlyiMn12M3KvUeqlANHmjcMIlqM7uLs+2Xm6vl9dnC6Olwmn/jYu2PPHwFpqrJ2blNgcU7GJN0Wk
ynmaZPUQIfG6fUI6ICKKxpzORGYux8B+f1OBrR+U/LLmckbjCa71RlxyLBZUiHdTqJOThKMWiTct
5suu3PBIhd5/cnAUN51G+2ktdfkvvJJaBP/VsJkgtXS7IVBQHZo7/tWbmp4Pg2CyePQmz+9JjclL
D8nRdyGyCYW+2XZkKMXE63ij6iYvqIzEtUegRbLvIBg/YZtdKkAyf0Uuh6dZv60Cim9q7yRkb2xd
0Ov2MwGDxHg1ol0BSzUy+Q9A1VLlepGuhlhSlzorIVj9ibzxupuYgtd8KMw4gYBHsV0+eVb8aK7Q
zyqgo6sBZ5TN6xad3l0p7LTtXn6tjUy+uI3tQJCGqfappGlXRnEYFDrlLHmsVoHPMNur2s8nwxgi
0Naj5kLSFcoTxGD24JdpRPs8yNncOJcNIK2bz2HMndmeSaluJgll+nir7AwZ/3VI+E0zOQCsTb7s
Uv9Zrvqepj2mBbUQcA/4AL/jrWh8J85H6R7aPGu6myoGsbvFhgRPbApNLlk6ASNTOpe8JzuCeIqW
1t3dD7T2yjlOMkxCgJzXKFtDenqOX7ZaaPUIyCqh0bnXBojv7mOuq+A82nJxipxzG8Rs4vruL6aK
Sc2LiD+iEdTWYUg7NeWBZtnHid8BDx0LtbKVQinXGcKAZBXYAP4QOiwR1Z1LGcKUo+E4Mqi5VUcK
6kwqQ5kxdpsJ4WGu+efTNR+k31qaO7ltlRL+sYrb4oW6236yArj/WLHXMJdPsKEEOW1fMA2qPe7c
/mc66RRWKZyDjQg4J7rrdfIXCwA7z25wSdoSG3tjuP2j8za466MmjktIZ01n2MQNcj4HBnp0RzVo
hkTFkiHDRWe3NVKOz4To8Ez+umZFblCzSCMIjOf0ZBbOLY91WYuXod3Eb+8qEzdcob3e1mlykN3X
O2q6J2lC3PbA2lbYDtm3XqUL5bHILk7hNpNiVBST5Sz9F2aNpWvfdfRQ38ToHnEFS5f9TkRRR3SA
CDZQAvkcopZm7uLPjzRGCBmA+H08uYujtIp99AFnIpob7h/KCspRA7D/kMkPEcakG96dctqNXkny
O3CtCjrhIOZ0e2/tA6UtTl6lQ3a3VljEIaxl5GotmuHjOMJ8AP5s4IIr2cHNJzGZhUgjYvW0AKqE
1aYWtWFcS8nZSCmD78M/fdCFrDWN/pypKzD/w+MO/yQIhe9IaYkGthCGgfCFszHSxUqnBvDUCE7j
9ApBH7eZgWJX1F7usU0OiyBOnc7Yu4UkHoPxb9/TKP0mZ5JPhVvZ138acp4I8iSAosgB3u0c+Z37
267qILfoqS9sJBhJbNnwlLWxQsO908p5kd+tmk0alCgHXuXZrp3p/OYxiva137nP0WJHLbp6ni37
gfVo1gwENQrleeqzhpa+6EBXuBbd9ah57ycHSGxfA6MA3SJN5MnWKN+RAMnZ5n+dKRf0oFKSQBFb
MDBcNgeEw8pV/B5ZOgLaQ5lnAeE9YGClpK2MjS2PaUz88s9SWVydqdlP0N+WI8LWufQRWCyCnwiN
I07LV5Yg4BVnu6XS/3tGCd+9ZNcGA9bQLYKLCHQCbB0N/bKOxS3sRGBnwHPMA4Vg3PfnfyYjfZRP
xh/7ZeSWxpSaBSBbToH8bFU7ZGCwoXADS/3iyojUo4HCkfRJE+JO2CklHPTEa63moOqQM2dZVQWJ
NWY5Yd9s8gbpMIv9L31XNzEI8bgI0xUsMFftx3NQTZfId8R1xyWkUVusE7RunGDcmWK7CfqN2CgF
KIVkUd6bqRp89pwR9EzT8pn6GxqaBqC6v0iDcQfPO+1An0cvKESRgCRoO9LlvOHQiCPdqGiME++c
OFqM50STkuSmJmL1PxQvc0LaLwzEZO1GddR2fImfYQDEVuB0AlC8z/BVoCZk5YUeaGvAVJxtyvwG
Gbs8zS1SNFHUNfXupOxnrqNR8NLqxQ862q6iqnQyZAJx0bjgxJnGb+CeE7XEdi8YeNokReKQghq6
8SAy73/DBoBM8ihwkerXs3zJ6A8uKUJSSxU81Zno+3HvO2ZWe9klKHLQbKo7JmOUmEynuU+NDyDJ
FqOHxo5M30j+7DMG6ENUPvMEHQrgzWbF/BDLe82S0xtWzjjupyxxuTdhAqLUfACyreYxjimc94nP
c9D+iH9GTjD8jfJOeAHS1OkJ94LAxqoRmAbetkgcj4PGiUBTKAMT95rCrsAvJ7wrUlja+jQ2VOtp
4pF4FxUsvyKcfOWHcILxFnQCMDdXwoqFcDroeeFPibp4fGOhoECyw31KEzTDTvecDO1u1m2uHrWA
OuiwDu3nrt3jmghL3uCxHk1thfY31YGiyR8uQIegkpRiY4fm+qqedyyfMqtpFI+3SfbM8ojNumBH
54eyGnm1YbQ1BJt1A22FjCsCizJWaI2mwWJJvffp3/0vUM+7DHb2gwff+Y58OAvVIwWV+oL91cAI
DYGDTlJ1I/FlpkR9OxJnGp8Qxz/hn98W2dqRg5XdH8zMYupXTZaAyovJwfsl65xgRverMJ4YuNR+
vYxE/Mdkq23Os2CaYyAtVfBPfrJlqJDfVkY7DMqNFqX8lDU8eOJDccLbZTdzCY9ijlLei0QrEQUO
U79RFL8ku/aeCuoYFopOeUMiqAcCgQ1ZLw2do/+SaAj+1XNRJyi5A8nuMFVBInbB6vr5DQpaNPt9
yrVgXwjNwWdQokUMd+cbTGQ9K+J483fIhpRHI8JMiTDM4p7pIpCvDWRgGJIfzBy5c3M1T1pXvKlT
jzXEBO/Rsqme0Wyed1qdzLS1L40lDz7nkufCSPI5yefPo85zKCFxEnUOXBTtZNpWXYoVPrdZ6dHp
Oo8cAdWeYHWjnu3ZfhHmHNB9GPHSF1gzX003UvqYidv4GY///RvHCSp4EjexzHQ1kMIlYvl5kVmD
AOB+iDRAcCius8SKdOpxpavSYiOR7EmFa/M8uOnZsg01vrem4zfXmOMp4PCdMikspThmBP4fcg2g
Jr93zyZm013EPC35kMNs7vNfgGxwM0QtcN6jXCLrzk9Sdj1QNdzxeBpSObB8eA9M5U7oLxFQcK70
vFoXxuTPM6PiP12Rc97gcPiftcoqc1R3t1lwN5FGx0QGB4iPatqwqwI4ocK2ZHTmuy086gJy9e2O
Y6rlw3XH5OOjX51F/Ib/k9ywtnEAns3DZxUlInMlf50aNnEjO0jdGI0CMGtf+O4ODuD0lBZKAP5K
vPnS1ER4nmmLsUxMTyHvue13+y/7aY12DtX2EPItalmODuApRy6qFBtdt0jx/rdDYgCrWOPtATHJ
Yf2kNkL2rsxurIsW+3G4oQ4gZ/TTujK6NPYYdwavbf8GnEOYjR9de6ObewvN81IPWXx1cNKP5QIq
nEMtkIS8TJj7eXSpqxADB9tZC4T2x1HCrqkz2lc/leA43KTyJ5nfhbPvlvs8MOTY8i1hNaMLaAfN
8SfGcBqiiwrVeUeAY0vecOHXTNg4tM9Ql/KfEN6x/35LdZn4QXzrmDg8l6y2KGADOAdHxfNrHJ/h
d9B6kgutXqsHB8dRVJiJ2DjttA6JLrws9WpXxqlkSHanY5smm9NTWrtX9uQwyNil+4r8YZXblK4S
AH2E2Hr4f/eEQF+teI/hAbK9vF8MIvzBfpWx5oTeA/oymfNNen5JyKAIENd3mfpUW3jv9u8nGM0m
txlygcgQFaqI7vwA+8+jTQOdkvCUTSq8jYEEtpQ9fjmWRoJvrvMcUb3JSl5O6gpVzk+RiUSWScS2
/bi4u6xJzTF3IuDAjfS6S80UkUaz4YDauJGVezBbgcTVM0+fEDwkISodi7ytGekhf50Ri47nPghY
XYcGixg9W6YBpVMDOMBr7QCHiw6k1U5LyJf4ZLGXJ7dTnpocH6+9WHw0hVO53BZ37TxQyfVL6QmL
vDm2YfD3yScGgBo0Xq52ifBMwQKTiWb88GXt9LfVk2NpHcNfJNf9uBgo4X4KU/DWaI1o/UimIB3j
02rW2KAVK0hHxnETbdllmQm7hl5FzoKFq1nFOZDT/o3iqy9NV9IUnXoBwQwVgIhQVi/1OkR+M5qw
D6ww2liJvvwg4so4HcH6um1cS6v+gHKbOOt6adYLgW08aUDrBRhQGz7Stti0OhYdOZSHr2ZrCI9h
VAMdUdJl7oM+MqzIvoO802WaDhCfX56cTe2BGnTyW3ChoQtlmn6IrKM+h0kmg8ba4qZh2NcKOHEe
s/onh7ckTZZ/QQfJ2gGC5cW9f1KEL23TazyC+v6lUUxsSYfYJu+DXuOKMefweZKg7kYrsEwXc/Mz
3L0XYJx7p93CYc3NFPemPPcNGWSLmWiV/eDmSiIzqa6KbthoUS628LdjPZy6HBLmYqgjIXqKL/lI
kuu7v9cpOL1ccCfAaUwQxmivWO7jjMnfUTQV9EBIxS1txVScUES/MxZd2baJClc8Zt/mx0IQyVwH
WF6mqVyxH7j97bmBBUTdVjkTJGgGKx37iBEHoQ27s2/hz/08TFhXu/iZaO/oiF9dsKRbw/mjzcDg
Z93pAwQR0D3XqsMCh2gI0zj6NAemBDeJzcg38mcKoPN0HdFrFjtMBOl3x8n6CjhCrIRd4G4NSnqa
9O0YCZ4YnQKNRZIQh/niaCA1pt+kg4lmikptRnVHHP5CieFr5cTuyw4pLPvDGwl2f3XG5E8gd+ws
iYuJMvCPDAxoR5wPoEycCck9IyTwBioA0K3l1BfNV7C7WUtZa3Wu+i1jaXNJDDBfZi0oTEAg4KBB
hwmeMvqxR4EFRc3bDAE++JSqEWGf2//W09JatoEFTGmjWvD5nsJKBVZLlJ23l9lTesxGFJPSi7zb
aoD7ngXUDK4NgrNvHFEOSqjrUueFUqDqa+UyKmYt1rHR1etms6arMT6CitI0aRDlgsu0Zx5cqp3J
VzHiiFBb4YsIl0cuNMOzg7Mg+zhbjoAnPRof8u7xvXfkjkg+85XIpb6In6xqdEivCHKHrzaRG6VY
hjLHaNuzzkWhRFhKdXZXPNraSV2pD2hA4hQ7iNFYEQUfb9bD6/3r0UI2xqC5gTF6jM3SNGyQVx05
L1Anlmf1ox70zAqgb1LZdPcmo85Yc/qmAGYQrndkDVC1MkNVHjxOBP7P15NjhgiXJwbq/3OYKT7K
l8KiQLr/CX2+BOwy8X5eSstD6ZyuPEIVhQi378ycyQzl8q0K5qPXzXut5CRcuTaJl5HsGt67KViO
FHbrjZGxsvCY2eWHxP1f4GgaCI1fDUj6o07BajhAkN0EZ0HX7JpvK9nSAZ2fWJqXckfs8pI5UU9m
xi0ddEoak4WPA+Xi/Q7QZyfU1ObjyVHElAD0x/BFSJVJvcbEUA9prsu2RdC71yB6CWynuhkSgX5D
HSbRxe0y3EOgddc5aRxt/1CP5ricM28F6xTF2l8PX69BiSosiZ0D3D60w/jRHnT2W8mYTOIa0g+a
a9YJvROH0RBX9tjhYL1SbzL0/p1TUlwjsAwFmUuHwzhq1r7nuJZlwrzlfzWwzfOvGiGBwI/fUBE2
Vu8q+o5yEu4pe0J57HfqEpo38AuAjJWBUtNIYBnJdY+R6djbtMmc/qpJmF36g2bgGvORcBEVywTl
XLkQtitW4hP3vODb4PhMy11959GVK4jfnJeCYzh0uYe937Zi+Z8Z8hpfrBwafJapLc5Qjad7v3o8
F7I8V1KGyqxaqP9yG7wu6egE+kJedvYwdsgchsi/vP/A2E/cqtxCd91cPOBk3b+5VMQWmNQm4+le
4XHHfhtug7Re1+ydPgUOFBlivvcaK9azmroh+jUH4HIcZRWXPfdceN1i0/EhEjEi4Oxfu8EaMMkJ
+DO143MsEoNCMHoCqEV9sBnVQvnWtHZQLJ8BXUSNY0EVswflKo/vXPIXsKoX/8Hym6xXPV2MR6uD
wwVSddGgHOW7tmzcpZGEylV0oiXAasKOvoNX9JZejC27cBrWhmXQZFsa0u935MD2lOoz5sup8V+X
2cqrT+b9WB+7jkZwJG8R95JO0X8esf8wVzatIiOK8pnYk21r2gucI7SA3A8EFdA2xJscPijPkrm5
fsDWpIe+f+KTZWx//VAPnsZSi2JarQCibiiON2rjsMjTjO2+sWMAy9V14jv1PnEa0L3NYwV9k+Ei
/KZdgfnAnfdgVpSvjls20OTt1cjitsAZ4oIkdO7A+KbOl29vhnV0DGQbEqKW+Nv7BEasV6hG2ziY
NVBhLk4oDKAT88GoqBASXS38Ym+4y9FuE7Qb7h/Dq30+w6HwpUUs0tD7JbDltYz+m7rl2WSzsbTX
tl725aeiYtNS+KuSBSguz6u+d/ciXqIjM1ou/v+XS7gsb1J10p3fPnH4GWg6I+5MnDwvkDiuWz5w
Ow8LKkAVUVtIuicGJEb3TauhdPnM+iYINHX2CmAaqOSj3O/xfpy1//6RmG5CAF4RzpC7hsKJO2UG
HZJhLm/W+T6ufc/udqvVLUkKdPTI6prQT2kiZyTOXjDdcpxzpCOhT5/dywfgEqOP+5NIAnEM7c2L
BxGHoFvhTpe5CKKKe9X8WZgKem+tIYgXrp5eKk4easR4ucw5lHyA9U+en7XkXrUVES++yHnSO3vO
GXB0jax+mKNFs6YgMXoOyqZgbXKqRB40+dln6Vd8MUJGXaSOuw18h4ImSyYEgzqP2XfvtAIzYLeW
VuV+hO35zCFRKyjqMz/ksZ+4nsRTvLB/kDIr0Y8aRKD4KhdajiH3QAY4lAYjb6wo5sp8+Y64eBgV
UaFTQNc5VwR0CMttEYnx0y+FI2eyd5JpgRO0OC7A3NhkAg/e1pKf6rpPYPGlbRBsEmnyjj7XISkH
y5UHiMsFlEFU9HTJhCSnHRlhfCoJylIKCqaEJx6stuyMnenuwhSYFsduGaVa2WSzliIoQ5X9EcrF
wpOUdXp/x9DvLNu1SOqtqBQ+WocI9Swjbz5T6DJ7ySzI1qemjYmODb2k2aQ/hHteYf7A7l4Qm6Wn
YvTFKcAv6wL9drutlywWJw4xbOIL5YuCmX+56msJfQ4GA/GgSFpXMtCN0K5hhGePAdmeHGhASsXb
zbvbvwUgSDNSdbEn3N6264vR+7y0RALgo4otPb/+L/8MINCbT4MllIzse/yjJ3daIXdvBEPqp+Vi
ojv5Rerq15AMkOt/jk+2/r9sZ1TQO84ooqMn9Stc7stNRKWqLJDCh6UZgEsxC0QuXny+LLIZLz/l
57w9RjRBp0YvZ4Lwkem48N6tQSfVt9+7LtbXgsdKHYU1dVuCS0qzhGcCSAQJzKqMnSaJpjkuvjFB
qc2+ypiuW5Cj8+eCGWXV3eRVWjlMKcFb5QUhPLHTSCQcRenahSkarJu3YWDOl6e+dCEDB9JKwCKf
GDzXYJobrT1xj7jKSwPzz/tfyXXKOm5NbhXWRL1eqyOOk3dzH3TYPCa/AAw9CyifauAPctlJODpk
PsSljE6MG6GH0Bp6UMPjdihkKo8/nEi8x2iwjkobXW0ris5l2VPavpraxZfzz1x/xWNGlBW5VzYa
qkrYV+7ejWOm3uvuvE7V/nDUulLZABUi9Ddu4Qf6/pE3vEAzimPl6sX7LdKTh89hv1LQxAoUJhlp
VkNVTWudi4hsHUTD025VkpGlv9Ldt+bcGtjx+sfVFPZGUBP8D8ZRbEmukPRTHZ3pEVC7pHkMqLUA
Tr/ZLNkw+a51seuxT+p6wl+f0z/QsOKrt89VS6g2CxxI6gCiE7mhwXy91/TqigK8uFCTDlY31RTP
iLOqtN3X0Mh92NTjK7jyWBntgh73egR5Bwr1r6JDOZRdddB6nJGX05zId8SSNgqLnANrgNyot1bj
g/Xt76fsIFt6VrOXLQKdFREbbtVa1+0AidYZp94HO2RrzzANaVfwqhGWp1x60Pu83EE+gzsUoyZV
4wU814SI6oNBwwR/IQ4i64FGI5nw7DRFAM3/D0v5V/XpZ3bHjqKKUQBSIucl2uY0H4epXtzaddSy
ozRVCfE9XlubLEst6Z7Ywc5HnDHJUOXTWFbR3/qJFEkE8rX0nkmxm+vYeBdTnHcLYm3EL01iksAV
Q1eES+TvyZ8tp5Cp97FzjD+r8jE9PinmjbgLdkSIImWJS2cSVwHJrKaDuTa4OnHwX+vUIGKzkUxF
L9+ddAqoOTpqVlD1jCb9KZvKbkj9vxJboTw3evM8/A4L9Ur86edhh9putErU1qG7JIq0DA4VIZ6f
Xxow1gzEm8iDscFRFNb/rY9/CaxcgPDGbDbLhInDISVa2hAA9+8Q+crTLRlcvWU/25H5dIut2Or6
eD6v4JaJ/XSXBCat/tih0x+UF4MI2BMIrlnP2kPUfrMQ4jyxF8EhzWCT5SOK2hw9heShDW8NRTlZ
hisYkcDP5dyMTujXK+Up8OQ6Hl2c5PKBMy3QcvZNsscJIgOjFxXvH+XmjaIeGjt6pn2UP7F6YxWI
izmIlJbQNjeVmFpO1R1UnbB+510X1JK54isUNY5TPwVnBrc4wgTWCmteRds9UMWH3pv5DLHoqcxj
HQswM9/2f/TR8kRdobQwtVunm3oJhy+xXf6ynBGbVGpFsVEa4mvOgj+tqTNmKd1bUTcChnkC3JuU
VxsgP/5+HH4Rj0IaDHaFxImYPgvG60w4FZzdrLZj+j14SzbwPFuqMe4oYq3ocbx0Obt6Mg02/ud7
RA+mzePK+PEY0bct1+cQVNU15hqg/qIJK2g+5B2vVriK2a/E2TvBt1C48CLrBRZyQfusVgRMPX5w
SWW0/u3flLe63Dw0ZwyD95qqSucWAAWv1EDeI1ZXp09dIAFj3bojjN7aQj/3on7AzL4aEzHo4q/y
apMOjPEHJik5/dCST8CUfwA6dlDHyEaQAb8IcyeAPJx6zVxSog10ql27HN9SulPGXH/wj00TEhRM
9WXjIHru1CqXpDPpJ4O/J6MCPvWW0mdekz/3M6rYc+wCPahVR6KH9p3qpnWwSRaqF+SkMcmRXGwg
PbEv6qVtVE4RUbg5Dqt33pAp2OavUukFQIMc6mYFJm/CSWxuzU5quo+pPKDJMvWk8jXMH00tQ5m4
op54z6im31ECkfQhdrac4D4thPpVVpoybJGrtQ7LFS0vuoYp167r7ameXv1QxKsNGQzDUZvMBGA3
tJLNFnR2SbJUk5Mrpho4a19MVobq7wiDB6UnefSXJYK3HwVGIzn8RagPG1QnTibmQR3emW73sukd
QxRFPfNN99oGJCm8anpzl0zBEjpLbQ2+IYi52lEjhCmIowUfQLuOEX6fMSxViE5sHBS9fBJ3OcI5
/BynniTakp+40SxpF3KmOFAcck+ilRp8hmSAWiFVDMfO/5BcQmlww1FFN0pnrd9bErnwoEUQAWjt
q18mZV8OMN3KCXzDZN6pxUiRVpZ2aqfYKGVi/8eh4PrpUdTpr1oy07uup5EJfUDKxjtnfUt058/I
W6ZYVOkeY53a1svyUNu/qsns/zVR3J0yHHpMcNqONSChrFkd9Kf0uPdsHCUpXg1inwvgRlOUEQkc
mYKoVhkeAuOHbVSmgSOWPSeaPsox5RlHkXARrBcyilEgFdyl7+X1jXhBBoqFI+s83PgDaw08hnf9
GlsyzrtDEPHQA+cso/37u/l4MSeBwNaRhcwC1nO2QUaVWgEX7398M3076qpa8lBoN61GY4NbhoJM
JCREGSEmwqLZFm++p5MkwgxptECcQuir2/EyWH23kFrR9ikY/+CDS/xbbCIWO5DLw5mACeyva+zq
iZu5kB2hf4IPKqTOAKNOeN9g+6bgCroh6vU/2D8rZevbIAAyIo4s/WG3Exw2r6hvuioUFDliRB+w
SEZpw5Y51rUfpfxByWamTkGxuCKIk8Gy3CTsdISEl0Ej9ztOdN8ROhailXlkK1oDFnfZRKlKa5Rg
nb6fs5iMSXI9/6lm1yShH8ygIGOkGMHqgB7mvratMPC/SwubLj0mnQ5/2GAKDuNxzin0VzS0srfy
nuDoeu7NWHNyVhG3wc/1OdPgVMYhI220GQsHHYafNPp2QqVJ1qu75saOV0g+H4mexQacjq+4gXcv
MEW7NRt0J4czmsXmQvgdfBpicJ08JNsIeOXoe3UWkydfAWUNd2tYNhljm+d7JreqGau0gfFji1M4
CjxvsF9QQXtOkOGEYUP9VCucJSorhRqu3azquF9x/KP84lyefe3+fF68U1xsLm4Y00kaZoAsHxi/
knxyIjt2E6XQkvMqAlLuWLEouwvB/GPRJtqEq2uOk/pB+C/Kj1130KNm80fXvdHSGWG7MAw6Iucy
ESMl09zPYNmwoyvafbnKvNklVc60Y0l6qSsvLtqzFG5A5Q+6d2IPQn5M2Nv1RjNCc5nSaiyn5jV3
OlxrzItfxJDgF1NwFI6RqitKqKlqBG73mslpHD2WUgxXrzyMwiQttGh4kJcdVnKlU3NSeKHBmqvT
8zQ6hQpf3HuLS526aDksxwBy4KdBdUQVWyU3PLyMihzOBPj7WVenk2xfyFMademRB9Vhl41rMN84
22MU9SGUMsV1KQ7hOmST8/5V0L+BIjSe2h9HUR4HnILaQY/3sERf7fpHY5v4KZZj5+ngaJGv/psz
7wD3E5VY/xb+q37/8K0RUavtUfDZ7yyZmvolDOxaORTXdO83hk8wlQ1ceKWXGzETcwPViG9JTm/H
DnzvzJjBmqFg61e9JmI659kZ0Kn4C7yCOAlyFYKZArgLsJwoGNSgJAunesKlQyv8tgTRdsSlpyCf
EwHedUsfzLlwm/EbL3Enz8aEA/+HRlT7WXQR/d1i5Ry8mtXJfGGj3xydmOgNZOdOikAEW/vjJzdc
AViSNtAao5b/kC4O93xxFdDPjF8fHw6dq2u+mqVXKdv2yNcKS6uYZpfghmcDftlGFpTMhFYmuIkW
d+OVDMOfPSJ1dhI1jqDGh2mISkLH7EJzBsYgYL3e/kRBAaacC/UGnKrTc1VidGitKIE1b8HNSbHQ
yZsdP3z0l0eoq0RDpxtcLwDrJWY+3G9WKEdf4G6qX+zEO8YtKoM6NfcTNNx+5orxuA6l9LwtuvqT
58lGybz7Q60CWVq+Kn6B7971IDlBJJ9F5B7fvsvag2QDVFSyAeBMmGmnMp8mAJt+QjGLcZWK+aj1
2AX2Tj7LlVl7e75qz6U53QWD4TW5jUsdgvRC8VYTnBiCrg/RnRKhzW4jXgMW9Gle8CvOPMwJ44VY
CFTeaDv3Cz4LcuelnWVC38gClUBCzbT8JkdA7C+Ct1v1Dc3IGFRnAwLL+4r2WhYRHfnec1qlxOL/
uCHnhnhpdx+qNA1rRHhOaTeA3wp0/nq3zbZbTd5pqPGwer01MSyYvKetBhk4w06EYb3qw0qIWP4F
1kF4UUaBWhJiEvUXRbUd34+wGqBZFOqQ9jPpbWETVL4Md71SAZzGGf/bQRHNBtpUI5E6fatUK2oT
KJNfC6/Jvmx0xpn6WokRUFGevK6VkerUkpg7pcFohwveU5A9gK4HF16NUYpp709ye+tPXs28CnjJ
LKaSUtY1XmaYfDjbb/nchzKr+alAbyawvaKYguHEyMHDwg1dJfLOJ4nsw5GfOi5zDWLp4rnN/Zhj
wGH9WTmh1nAhEG4t4UEsRQXpO6VauDemnmMEhknOPaV21QqUrU6+il+FNZUNewKJdQefzqsLU/CZ
vhVjaK5oW8OkwFpRGgCNf83aSSxm9V0ILVTIWMf+g8T2dUiMRS5Wd+JZo0C4WGDtptecjeP5ey+R
+uchNW5NFoBmeSj/j/Q3qVDWar7hoiK8+ZXDeGojSCCkDPU8ocvGegMfHLZYfKbO+1qPPF3pN0j6
ZtaWkNMQeDwqHyFEXf3WrsWN5wK50LBObJA4JhmbQHjsdsxjZl+nV9g/7sJ5GRscPSeK61T+/Ocs
651EPAUIdZzo3d9U8J+zl+UDcgNsXzSgP8JCqwrFX9Pqctej1uok8hPwUSE729srMf8q7LgAl/Cp
4chv8Fplt9IMi3/YDMk4m8OCFtXISCFr0QTSwoFvsLPZcQ/VtowrZn8/goCTqA4zwE/9PHuqrGA/
gJ89iFYZANoyGGqNb6zbiGImoAoCvMfj7+hxOIr20z1X3MPVfCjlZf4wQxypc5a8rQAMTNqySCSq
tG5Tyt/LphEw93gCeUpCUCcVQWLE5BKtYZmKN3s6W9VcO+6BjYTWpK0fVWAEFfLymtksSqGKbEUF
Vh6S065lYDrfwyinTZnbkWWm5KEAMunM3EoTtCouYZJAKJtVZOdNNc0CW7b5B2Hc5pgpgpT1MljK
PhBsemtT10tqquX3Al1TeVvo0ekL8kfNBvUutGaCjtyLkRYF8I8iquXIO6N/Enw4EJpbPQByQ+Ew
CJLCwdb3ZraI/J4/AIpJ13Ev3LDjoEt4zxf87C7EN0DpcgnZgApXF05Qm3UPpEiP7oj4EMRChl9A
E9SWodmnUBB7aG1II9dZlVBZ/kPz/ixYB7ODNAViHftpFBPAT6NgdUKhpdZp/8HLFgPvMkvrjBzY
HsbvcVqOXhDkeRcggPrb7LuYo9A8vUEpV4cWXjCWelTQWvVIjjwwG6cpvniufcwxZ9RrGz0enqOe
wLeT8Rp4lbegsUVu9L/HfmNrkiK0eSxgTHoCQ0jN0kidWYj1WlSBGjNoBGFY8NWhf8P2czirCUc/
7WPYsZdU3EhwR5U0XlYM2aLwaHC0Qxm8kT00wqfD8vXMogaLFhHi0bmqRBZUEdpy2r8y+NMJZ9Zz
106qKo3D1f29tBOo+8LTXQgJGIsTkjzWaFN91lb9WWkK+GcJz+OHEd9LB9+QRKkfuJp84a/DPqEZ
2uMS77qyCH54itAQivWEtgA6tvjtZCf2IRNmQuqQyXcw0jM7p0K+btgVlv85kynP7rPicdnq6ZRI
iuvJtQWZZss1tIOouFXEW8c4XNDJmbXvbrIMjUsJO7a42Do1zVl0n42sihAqeX9rbWG27u/RgezS
fBYwLMZrapwFeHJqHjGKfgXRSTZ0C0AuvmFCZkBCnVtIV8Ij4kKvy9ZvLb2EHJDhYwAA+MtnMfMV
qc/bRntHjOQ1TrhoTt8JhvWpZp3nPGWvNmHYlLhFLkZFGOpcpTS6Jet9nWlkvqxlded2UCwMITHL
9j/Kc4iKRQq8YKccdI2NfZ1fA2K4bG4z6MScHc4ckDgZJbai4QrScV/o4MQO3xjygk4fwoq7aV9E
+3qN/Vf0wFiclSJuTFPzTIKeUPsbcbiV5RCel8ZUPMj8mmx1pKKdLM2ifq6vAPyUcu7Id+d7OqzI
8HDsPmC6vazLG9waH/vFDLzH3pNwu+fZgXmh0vQaWJ8WBx9cHOs490oFmSmnqXi/UMYna3qwP/Ae
2l4lbuAZH7OdLt37KPM10lwNtYt5o+lJeT3mkhusGhXBdpt1vAYcCiKHHh7i6OfL7xMi4OG4SEZW
rduKdz3/ngpKgUyseE+TU5WNzWCfGz+ZoqSBgFWILL0brs1YsJ1z3MIkMxTSaoPMu2j7tomteH8Y
Lere6G0ErjVbmvteXLV9zS1Noh4IFdqSlMm0xUOWoIuwHRRbV9uQ+imknUxXxJF5ygkaTP2D8kKl
Qi3qFWrkFvtWOGfMTFIime8D2UG072xUYbiqbuetPiKrpVau1fMTeXmD1DxNp26zrHpGdQ50vPoE
Tsgol3F/FnQVXUOGkKNAQRGxzDuo7LJpwtxPFMGPhN9Dnewogngy1W/eZ4djgXC3q3HteDEVMPtg
lJ7r3TuwhdtZQP3jGiPi1aq7UGr/9gIk/bIKkAD97J45MFlk2S4btHh8MN/P1+T7sh4lJHLJHY3c
GjB7UukZJNgxmnQusZceOYsQGNEQjhk6Uc/LzS2biSvqOHWozQMN/TaBEF64AaVmK0zpHE1ufkhq
24MyBf8ebxaWWwSNZ9eIURvhTV5bh+kiFloA4drCmqEUuut4GIDjnmGXDfopkkUOGlNh9c2lD5L4
LI+il2C1Wai1j67Qyf1YzgFZbcuKSGF9u5e4RKphIOy9MlYWK7DZdRBXdFxIj1XgkciqcmZ+HYDl
lyw/dOYG81gHsOWUyn7vzIuiCHdfgvf6RLdVvBSZylL6H4SpqIeDaZVrLOlp8DghBGF7TLhyPnjM
tPTpRMK9AsOkj/XAfIHnqskUr6dxnoxeFUfFozkF4DvB+aMmka9nnSpLCO7D7rnw8KT4dSkq1SOL
Ixj9JeEcT34fdsNinMY2XCJeH+gRHyi7LF6/bY7ZbFcWVKXgF9dehu3nWjRBj/LeTI24tscP5YfT
B9O7fP+MgDX0K/CktHIFv3TJasTA33meKk8EvLK9DYKXL2ev0wCp+NzTYGZJLrkKFa2J0Sp+XJpk
8Z2mQU9vWEyCW403B3Ig3OVPXDhgMaNAoUZTatFeMpKuzKe6DcUpynZw6pBGyw9u1mN+4XhlCVuL
hgv+JBYCfJWGmZ+blh0DK7mb4BnUrBxb2vie7qhLWvXiXoxLhd9INyq046/h+W2BPp8zL4M5xE10
LlF3/CZ+hy7O4197x7MUvIjBlnV044WEu8V2LbkJUoXsZLgdQyN8JsViRxezWSHELMhff5o6YDtU
WQ5LNvxwwrb8dJ+uVloPLP9cgoD1NzsgcA480VwZPUDw4RwT7slbISB8BXor1+lQt+mCmMctXMLf
ptXeadzMA80HTEP3sHOy4SV/k5dgnKmR8QuNrx07BQnV/BTWViNPmOrAKuNneKYWdhvOqOlPhigm
ieIQzi9k0VbQHFv55ekgLvFK+CG4Xf7SncJzXXpt0Ni3891FMV2F2AnmvV8gkU95+evsrk+U16ym
RWN0HCbrRRGbSYJYq1MVOFnGn8lZ2j3wCa2Tkw9OrybKsi1Cizw/rkZt8F4+PSgsayTL1IJiFcWR
gSK87P3OOVc5VVC9A5RfvRHziyMIXFIJRKjkIR5X+rMFu/GtCxPfyclt2cLCbGDs1h7J03DGauGs
XZVegK1ATtJLPsV7uQWPfHtitbAnI41c1E5axHjiLiv3V44ebjGtJ1GnNq/YkHqUpHTRekblclen
QS5IU9eIFlXo/tj+f9d/jAGTbwT3k3Z2MCHdLENxcXKuj+HCHg99xmmwb3T/FL7GE51swcPOOVy1
n6chzyZMPkwX9PqTIl6ztTqVRnZkiyix5lPZtmcIFhxmJgasOVlNMWiQkGeXM2qozICdC+ZomlkO
dKzDc3prMMAMb2N8/QAY/NTq5HSjYk+KjhRiBKia7uGLwMrE9HdYlcF4mTsRjk3DifEZJ1AKq65X
9c6eca1MGT5XkJtgQ4EFyxHX407i6otZp62tmkR0u76KLNWDgKhnjZ7FMGyUEpJnbt4xa2sfqoBE
XDi+ZGM+cpuhqfMzuxf0Na0Opfc3yo1K7OfMzY0g/csOyytZpLfCmv6eXJlB14KoM8UFy5KzKihm
ptOmZlirX782VxplfU8Xfp8SrHSQPCWKtT7VOPBwkWj0MYWSgZ5OAqKbSutiuGsi7RysVL9w6Vi1
gbEdTyt6ct1MtSZ2W7OiFNZUis7TdBGmiZy0TJH+GHolEaOOmU8nP9LE4OENIUdOI1ahfKZ36KZF
a8zL15K1Rv5yizJOTxV5cVWjts54iiHJuj9J9WPIUyCNDKSQKoitB6GTQvxeuN1O0nZ9RDqtlnHy
JdUIjoL71FQkPXp/GKuSN5tkuxS0v6ZjGHS+cFQ7KeD6rVGnzsiUx+cpuY3ObGWX1NTxhuep4mhY
bbR49k3woK5HOZyeyC8BPSQCv+TYSDxDJiGGcGh9xlz4PCqHjrB9g+JmHk9rx436yQUBmwLGapV/
R/bn7y80qdKFnjeezDMam58tkeNQcmg5E1hERPkse5BZqhNi3gyEhcsZWj3JKVlxtkKr8gYiEz4z
S6/8j4DFnj8x0RzbcKRUYvHpFAS1UOtLxd+/9iowkK62NX+ri5EqorW1dh1VFTHY9xMZORiDzQCl
2fqS4Vo6DB9OhaRwo7QsLrS0YK4dEh1iobCmJ8aQLJ1hgBDQpsxLc43YlLk/YocNMnpUT5MmFlRl
bbEV6Pqa4Fuo+lY1pa/kyQUm+We0Fv3h1+ff4udDw7TJXES7DvSBh203e9zCvcw62nMbk9F3PQJ4
Q24TvnPkI1qwUfjBm+zsJZmx+LR4u1KlHsqRCOpXvez4Ewn+9KCMzGPg/CVuAM7IwQUGMnqqrKSX
zBEp0ExTXNaOfE3OVp2nza6+LJtEdjFiSeDcJFdtM3cO60kaPDO8d3cSqkewS1xYEOEaOL/jvfM0
OHrNVIYVuITqnyH8YJ4pgAe79YxSlKyfvX54/yFiZlX5gm5I6hjmG27a+b+/IRjGGVSWuJ5/1s/P
CRu/5p2H/+M/jjN3iV50UWj8fCeB01Tfm0Y42T/PHXAQf0uUANF50glHpEgGBsabtk2BSkQpYJ7j
3c6UEc06CEngt/WBH3PhS3hOGIfDie/1odo6QV1K8zeeAbFo6spnYPLdY42jH8pDVvMh/zA7itsl
SxBEeCWX8VXecQOsYOUgYvJrWvH5ZsqjLQYKORexQEPQLCmt/yP8Q4SAW4KgcFDSIVqzmKu85+3z
Q1Pv1CSLakStPe3b5i2ABQvNZx2QskpdwjrBozD6yESsp++Xn0pUddl5Vs3GIVVif8oA1jfMM3lL
vsOwS29NOKm6KSfCuLDGtpKFqZhK/iL/nn7H+xJuXqyyPrf6cF8Xr2ZwAcbLa+cs4pToCG+hdI/1
K6zyB0B6qPDrzkcL8m3Tb6zOgL3n8t/vmK13Wc6XqgQ6yzjBcA4gJcC7YnagUDHIyFoRQX4TV7Xv
HjnuxWIt9AR0rtkK2oCQFAqcV17DXqN9b2kYKyXz5KIxC5BYAb61S4gOZEyT61+jLioFPjawgWZv
V684pJ3tpNhrv/xnvlPAmCjbtzgpYIr/s48UaW12yl9cSmy9z56yYUAMmfG+pes1ERTR7z+H0m7m
JvmVtWyR2LHMoRRXnwkoQheJQaXQhTRZ1QU2tdQhTjln/CMZDsf5QRujeq46GXrzB8SvjdOXs24T
u+0xivq6QTX7l2uRpZTVOf4EgLgaz2VOyrJj0rDIWlnB6G/vBHfOSIiHBKs1+9I3TXXoUwudiGTw
U3egOOX9mSItNtr3oj263UQis42TiAsJA9ejp/onS61TzqVXPjM3p1UkSAqawIp2oTmOp50EXOJy
WmJhoxya2Vb+gHiUQWn0QoorbXGA1hSoyRDZ5p5nneeXhhMKtzq/H/lqihr7tNijY0YP4pMB9Nj6
cRwPqc2cNxrLDalfhSbL6kI7tAi4r55uDRvTtGy94r7YBE+oSslvNU71ysbVSjtnw8wwEa8ZPbDF
KOKHFgrr6ufszVw/xqrSEJpqjSp/6bRdeuuva22UEfHNC7rwgCXFHNMU5PwOjzvKrWU1N0E7qDQ7
xrqH58RUaN1OQfM882QVSO9FVCeWr3MaxvQ3bEG+LgrTcpszyhc29/jWWti/qT1rxFtJ/FNxvR7B
L7pbcccaWlS4w8cjT5JIt/WVnvYQhwxJrmSiAWtQBlwybuuiaCxidAD3+0cwPJarS9vWSSlNiehA
wFDsWHoYHJEji0WevfMABhDfUAmNGCEkXhq+Qt2daV7ZUs3DWM48LPmsJ0ZxURV+anGDRHCPhHoI
m244d+ciZw/noz4RbWGCUXmSnGIj83RDnzq8T10lXqdpwDKhSkjuVB3/WIYb00f9K5+JDOrPQlwg
JLuyI4wjvcSfZn3lenIcn5glCf3uuQq4weraKe31FkSCawIBJMPaeQ+1e/jtUr3O7Hih35jYiizF
pBXNGvjCbePp02AeIbnHmgtR8R0UKKN04YJukhJiw506HyK5hAuHq3HCkYjgYaWt+V7DAImaOX2H
xftoPUdau0XbMLFijLVqpQF9+WJKDdT+b7geRfMsODW5RNsLry50YJHJLVDlOryjXMjKJL+PHJRD
wqDamuQSxFMyyE3z9MN147zwOx1SvPlsA1+3az/EqXc7MmK5eQT+w6ugwJmTD4SDeJfXrK/I2UqZ
DrKsnG7mVORpJ/0WF+maqR1Qzl0IYE3iadUXpcpcP9nwWXLhkIBWuf6/XyTtJVyb1nC3Fc+Wk2ro
Ga8MF7Lpo6g1kwCTMx51i+LNvGtviqpToZnamJ8iz15SRjYsc2HcakSagKHzzsYzsw+gK44VWwv1
0k2GXQBLP6ZihmQWeEIfo/KmbhrYxqOClcp2Q0mXkKyU34q5x8WX+CpwPmrLp07/uiBANdBWokuK
ILALls5P3xheKq+ez4kP0BXJC0K8ic1w+gLgADYV3KyQjxo2ET8HW/3ZNxmTINsq0kW44WXJ5L3D
wKMWttif6zcUEviNRr40yeJ4r+sz7bXAKSfmR6GELVGpt5tK8cCwaIRGnXIGS54ZNJXDuqRQzZnB
8PWi8Udkoq/xpaaFTH5lkZMd7DcwhI3SPv6Y1gTRK6YuMYQhEwrgaL3YnkVW4uhPmbcIS0kMq9ly
fdd03Xi7diqwquZJT3Bg6x1oQ5lEO0R2tqvoZ4kXfEVFAOEAKU4dUU0SKkxVV9FPMEAZC+1kHUrE
xbDge/REL+H7wEhqEVadME4w1M40a7WbVtoRMkE+sdC6DuaLfIHMM1mAZW7DHqibOiRUo9B1CbBX
6wLxr1WfbmKLchm/OxmPFH7jrAFkAOo4aGUrBlIL360fNo4BvJY1TPtg3aTrMMfaJ3W68jyd7Sbv
OO/J7B3crA1gjMkCX63rSnlv4ns3JH3+ksL1mShNYWjTwi5lHxL4FXtH4eQWyc7rmrSZ5B69Ywpb
orlKPd+MBWnZxhgcXXUx1c2+OUoUa0H0Gp+uGczdvR9xu50qyb8yEPKkGOJwmYWEc7NXMS3KABwK
8lXhmIkv7VSzykIAc/oD9/sdakMNpRUZXnQr1nb7wP7bcuGyBvIxKEIpddv7XMCOoHsvuWmHVW7w
t3b+SsNaq0e8zQy1L07b0rgmPLK2FILpgkZZ9NoND1tRO3xbWda8438INbYfbr0XeaoT9f1rwbCJ
8CyEqREwT2bcMyzKtHL97jBv939Gswo5IwP43wwyNgkV0YZrgF5mVD3cnxuw9msjzVQGScHbDC8F
i4tXUIenVgH7Z0iNZpSXuPm8Ov0iFDyfY6tBgAYu47VsPqKWXVy+Dy+9Yoz1/qkrYj/NfWS5b+Ip
y4MVr2bH8yK507Je70pEtpsQGq1KC1VeN4uR6Vp6XdN5ZiWV2RMKHS/eDXgckYtWZVTJeJRMMlhh
x5cP8L6Ayg5a14plhnw8MRLT6vzNBfR/DxsnGbdOwa78Y5NY20pnSUL3VGYeIyricwT/EMFn60US
hYL1+icsVEZQnNrIx4tPduRi3Hm5dCcfW1t7DXmvwX5EvRfCnmwTmkiefAt+Rvd7ti5r2Hzkbaba
7YcmDjAHFJCm2PfM+KUnEk+fC14Ac3KOatWxQyXp9xsuNsl5BM3avAXosDBnx2YBN8HuHC1VZMVj
+dMY2+vCS6ykf5QEFMHjXYeFt7WvcG/8lQUK+EiW9ANmoN0thd5hWiFgmoXznDsQjHt2MeauxmT+
BfHKkr1kyH6cAy/n6qK59abR4b9s/faUY6o6ePU74zQu2bMz3yD/N7GMS6PoP00XwTryKvhXjekQ
MGUp3Fh1NjIfpAUATZYQvpEGMbufANP4f2jtWjKy2rK0Dhsz3kuaDQo/NoBV1jAKr/oSqz+kH+5c
+GYpH8IMHemzPUjV7XNVHDIHYhS5a2GXcsFpoaJutM2aAobkn6M0v0hR9Wz3fai/vgGiGe5iruXQ
Xu3gkvyRgignDvJujwbjc80TRuGu4J727uUiEi9rSz+a4WKarPK2rPFuKczZCWuLbWCYa2l3daDr
mWwcdFO/Fgnx7ahkjSJXZpSFBLmVsMZ5NN2gC4HcSpG8fCADbHgIKk5eepVUQJwMadxnGLADQv0/
F7Ueup4GI/6SjTvtDQJvmWYX/Jh/9tEf7EAFo3cFJcJ8oBotW/m8qYFfcikpUyN7agXAR7HRpXwK
SWCHuwty69JFn4CTiD5tSdYgYR9SKbnD8dDKoqqRgC5MODntfdXKvnnSyIR++b20MgqsrvLaM23b
RVCvnDryevICG+oWJghrfNnMPKaf74leyLxGQuwyCSK2xm4dhEtZQXVLhn6xa+daE+/tvyCcIDqS
hEAseS3gFrZuboIs0Wss3ufjExCM4RSW7h9rRrC95iIQvkMYuFJ3gjXGa8Xkwp7ReBn/4C9FslRB
hFGwCh08d/WzcxEFH+jc0ddX3QZAFcNbsniotwjbEOjrxHKmqaKncuu1PtlcATVGA4dVTfMNUSiU
K0dxSeuDV40E4TKpg7tSF+2yQnP9sq3ctkKwD1v1v8EmrOCQuYZYERvAvmtixEoxtfv9mhDbSQ15
MyZV8e2DAfn+2ktdwg/QtcWwrYu389Q66eEbMSeexLZNYxgybsz8TUG/vHKr1WK/Q4DhVBJT2+AZ
LwVyb0kiE2cAxbTMXGxNSqoFhLGT+33T8RIZZS+J+f94YsL5Voex+YC2sKNEx509IOn0ndw5+/QS
7MgUIfQQWwE3Ir1e3RreNOKZ242KGWsuBqzM6CbOhPxyVcsSsdo75Rf6qzMclCmzx0r9xpqXDTXX
7XvuZN+Q/S3dTtiH/yGmGRJnZaLviRYcoxdtPwkhw2rhDZ8ZPWfOSDzNdyH2zWPqjAw95qzWk9w0
ZHjM5EyTpkORhq/IXAZaXGRHVjkjEdwNCj1KBcJBahKEYNx0BDvJRT9ozvvNpQ0O0ITs6af1uwBW
MH94j8JgIy1keyMpHcpA/7T6YxTOv0fS8T+5PQ7Ooz/yKkTBftaKiGU5t820Hitz32+RF4NuPq6J
xpUneLHT6DaVafP/OGbjU32gywE84l0e5F50t3wE+fYzWJ6L9Vfkatn+rDNpa/XVy6sMbVMdhehL
C3DYd01uBBCzMuyiwz92Z2wlfg8WQ+HUK0U23k+zKeBLSv1XH9izcAzwVpAgu9+naxZ6L+wVXSIB
eYeJkT2GNY1IzE6pFtVzR+xFcTaoO6FZcA7Kv6H6qFjyyDfRgZz6KEkEPqfk+u/TOl8xA83wfs/z
MH95da6XVvHFaqK6POJti0pPj//4sDK/qSbU9nausGgm29DNzJNlVlY7Oe/XaCCA2fGh9TSOYtn8
OfFNLk6VTgt9WdVqRRSPZGbkEyBEQ+um0N1/XRyJI3HSe6gsiMBfDMWUPRA9F5IuDiy74l8hcmWu
xWFWI/x/UQnxQqL8xrk7Yr4ujydZrHJatFmXMMJ4vElV9ac/75tZ2G15Z52JfdLF6emGLHE2+iJg
VezQGN/k/deF+wAwrJ+zh162OmEFTwBxijsZPHINJ0cD90ooZ8Yz1SZu5+kvfWwJOsmFBMorYoyi
sNn4P3rH3Ck+qOobCSFFNJo2F5ER3Ul0teeLFliDAlqs3e+stSoMTU6yPF0Rw7ZHbwrlAoUCWokp
gGfGV6BLnCSkOQTdf/4ZB5M4CC+XtXL+VyeroVIgMFNjTU9Ssv/l/RTLzD57CTp27QinRkZa0hUa
CHa60LPqreiaekUgtBuZ/LtzOPu+xQkgrJflOkXEJzD4+efE4hhNCAbjl9yZig16DzMSBvLUATJ9
iY+4qaIB/MGHK7GyQAE5Cxf7miuBHKvkahsxC8HVjIMDkbsKHi++Vz6Qnrtr8M1MyFRqgH3tTUMV
VMvIyHi0V1V3bzMIrUfI5kGjK/2S0HeG+vV1TjLOjQd4oyTKikkjgYxpnDAeaCDiVEU1RsP0DXUC
4ZLGzD1PDQsPbqWPwuuxFEP258DEPTIxavjoBwo7D48v/sjgprfzfFGAyXcQkDXH/P1xzsh3IzxO
jvYqYYlGzhS9tQh8EXnPz9H6oNsiakWaFZZOofO8p5xeLua1Qm6scnv/74pEd8Pf7kPDVhTxM0v2
0yzRBoFvk33Xp6OKy9XyJh0oSbi5RKF7Aqo9Ve1Nk1e7Fs/o3Bo+Zkemr5BMWXlMtaH76WB/teOc
lciydOq0BhppNZhV5Kzp0TB1LRnF7lLB+To2DE1vs5DwsLNjgux+EEuZzvSKGnMa6wF54Bnt1q54
XngwWDLKLCSrgE9WrHBBtIHB8V0b8I8rZ00EzW/mI6x4U0pdhkTvXymMOrS91hvbpFnmW6Riivom
cLSKXn0Y/boWX+3Wes/Iawlly0/SVq+Cl5WvbNljCTjj6QvWU620AXj5jXEMpn0DHXrRKfjcJe/N
E0Wojm29Ygg0KHdsiXjdC9/l/95BcwtBanTp2nY/+nT5LgOr2FOK3J9pYYMiIlKVYTNQ+Ttfnbmy
NGL6ORmBX9IutMh9zMvSW70lZUIXI7IqIWHpMms+T3aU0PBSUftOe9A3/mYAzgMKCxGH84CLtRBX
Soi4dNEoWSgiIn5sz8hZR2k1UFGpXNGN2W5OuMB5ev/LIvntYP3VenvdNRru2oa3ntPaxEAMMXXY
ZAIVk8/G+wBAhpM+U/BZ7EKjiSgxpXAlKZejOIBhU1YrAJEv2H7MyHhHsYixp/vQ7aKavGXRWwIa
epyyn6wzaAag/R4J5r+JXwm6pmarJstrXXbESLzxvslTMBPF0yMKRS3FUdo3GXDnax929xBUfRox
dKaiS6469K6sCRoBGLcASRT96wUUFzxq1USrtAmmRsGMhfBTP5emcFIF8ApMUhlu8TCrZ5r2pfzr
Uc9qSJBOFqvzi9ISb3wIAH0NyKFWAeypz07AJJU9EH9HyFF5AdBa30FfH74F4+Zot4qu9aNQqkJM
xffvsfitukh6koejJIq7faV8/Y+Je79bMSdnalcLKG+LRd3klfLOpBvFQm//oLCV5LI+tCq2Tu8x
BOrAe4vYCtFdS6wR/0oXzUoU/qStZBgQ8bSXRoAfqlYSBa7sLr3c6GSFGKSiHHF2N8cZoLOAAi9v
8z4KlJrhDg3JfWAfwz7fq5Tmn5VXMAypJNqL+4W9nlYgxVwAYLi6P4uTQX5wDVnzGrI6aXBwXFCO
TVS3QWF2zJnh0kDyeXLNpgukj/VWVTztPFSdgGO81tm651QDy4Fc8jo1hEDXl/tFwcBM2vJc8yqz
Jt44o1WcYE+HY6eG9XujyUfmzg3I22f8p+cGawz6uiN3B96bVmhKZoxK9eYaC7V+F/LuGmJ+7a/M
ltQjQLmjQWMrmZ/ahBjFbaR+pGr3VPM0ADS0WoxbvluguAFKUee/WToCP+xGSrRnJ1pouW8cIvkC
MQ/mHNdsYkF0ZCIQnd0fRwNQuDOvbPsCaGjfWWieRchGXMyiVIbhgiXs//7jnM0gex1Ee219AL5j
8oZ/6x+apL6r3vOKUan066p068tOIFt5B0ETnD+ElaSbpQigSHn8eVhZwRnxJTlNJozH5w1h1D6H
KgaqL8GFydizf3/pnNeV8r1hMJs9x97ETKwxWiF3F6ltpDh7VkC+A4fn+9ze49hF8eftXR+g6C0H
BeofAQe5M66sSkAgV+bg8s7x4le4p4W7uzEeRPP/5r0jYl2GyRnG0PRHJW31XA5hhKplFrjVe/WQ
PGswfS6Hn1rkqCas65rxVyi2IkSZ6hB8UIgRgoZ29YQJjHNgqE0r2rs52+pYQ1aVV2u67Rv0xqav
mrXYl9VqK0e1Ik27qf4WFwb6tGgEd4kthnzWYWjk6+MeVpkgZSM+ThFjivRmy1qUaad9SXvHcmlV
9XLz1hV7TH6u6Q1bAmXxPLkF/tX2J4Mj6To6xlulFXbIjiiZymUaRM77mGHbIwsaBXaPERoI/U9g
YL7b9UM5jsD6YK9zBZZAfAS/ddW7jUgw4Pz/DqqkEo601TblX08eD9IFDuuGcAin7SH3DsqeoEWe
r0dRCMqWqaX3iWJFkMOnktC7K4bg+pHPqyYFFaGaUMp4q+G+EcyXK5vZJuyUJvuQ0u5phAqwpeYp
oEwQELIyV8Tq/iWVnl8Tq8Ak+OHq3nm98ZjtU4gGJqlMBYJL/c7yvR6HCmiJJXmpqT0HFDdF20/g
uBjGarHTgkg4DG3k9gso5cAtq+M+WUoGjv6cE2f9llm71UFIUv5ryKnKi1O9kLh+gDprk88xNP5b
Hd9oKR5Je7mG+yOqxkMStCHYbgoC+WAl/iQeSH+sGSNjaq80FV38G4bosWuW/gl9IVtvSJpHd8/F
gKCjrR97JVOAe7RPNsCzjiiz6Y3i3erYnjzqLmTYvhb7HE/kWklGQ0DT9IzrL8nTB1EShBpOCOHi
fdNQBwF5IWZSMZd7vcB/a39B08V7X4voQuFV8iXnF28X7+LFboRc/P0TLFs7oC43QAc2sPXazaSf
9M7RgOiwLLC4Vr6o+741d+SlMbhyvOsRUHAI5Z6jXlhjgcQo7CGtXzSJ1Xl5VRux611HMdqVKxiR
cnBIpY0L9FtRYSyzMHD/X7rVT4HS1d9BIc6PvXwTMlwIlOjQXYVrBED8glAEQIgKqJG7ab4H/b+2
dYq6HFqzKoMqE3u3IzQ631WhMLEu9RWtNOMwB91Boo3/JPLpSePMBX7xd5ucthNjW2M9yhHWfq1+
AEa1vukILIQqY/6sibiGXa7gMaJsXop99g15Ao7vK9WK3NhilctL3F53m+LkS4tNR5m/r0XwZ8CT
14I/dAE5e/wsG6UrMsqxxkIGq1h3bs01owlPLP8/EMLPiZIOZlvDYVOPM9rBQX7Rxq51hCPzEA4L
6jzzdyJU77S9SZLl6hP3o9jHWBIJFjyTQ/9FFKm281olx479N2RTi3Gnaaxl223cgz5lMydyZ8Iv
yoZqK3XQwb9x3Etk34Kea4f5iv9OQuW3Yx1ZmF6Btk/FgCmqzDm23v5whWXyCFu2IZ9yg9cfezMi
iudWjO6eFxh18k4NIQHBCbs1Pulh9RHukgmvMOI/YNdzmTza2IiJA6YB6eGW5xU0huK/Gg4tpXZy
zeTG0LW8pDPaHJuYB5r98FWPQz588YcW6+eclim/JREkRbiOzkKI4wGsXw2+T2ItpK4EfSKo2Vi+
dKoiZ9gqreBwV4RDCK6ledPN1S/zbbKsAlXAb9uIEs4qqmWP4h7m+qFIaem5PpsKLb9GFDW4bKH8
v6fBricr+m67EA0GCr74DJvVM2ArKsAN9jnM6fLbpveLOuyXnLMrd42itq1AdWoyaTeL3du4mzJc
gYXTcwKCtTBDT7b9t/w0Uqs/SXqe12HFCj8UuqTPQwhp9v92RL/SMoFeb2XOh4sXTI2NaM9kfnlz
s0BPtmK/NtpBw/ME8VlLcp7w+0pHfAcAJeUrvR44ebgvA/Xa9h4aWsZgDs1yITR1VWDwI2BXkAbN
w7qIbZvFgXgzoF2BPxHnQmqHYGGLGmxFiYAO9ZRKLDNYrYqJvnvPQmNirY08CzNt4fM4FU2FQxQ4
jK2yATCwvMfoyocQPBCcg0uiQqdWF+y27u2twiWKTwnxQ/Og+rc2xCicOeIc55v/08totbiXMC9u
U2JxWvJSqNDMUkejeK9Ck8x+lfG8Pa8o/ITiBwRqfd6yncsPzTkJ57SW+BOUDW84kbO0HWd9WKlW
L1DV6+E80NgfciWZmpdy4/KUzEUSCMBoflc1plY40FEh2MliJf2JDJfUdZRGl+MI1VyDXibw6qbL
LbTbxNBBrbY49VOmsxMrBZf8w/88IoQrDPRmuCEmX3wF4PcgF8v6Vx+J/C6OCl0qHIVMCCK4LLdi
JN8JC18O7VOlx7zEy2upI/zaGNFnYJZNucJuF46vsouJF0MgmXWUc0/JdH2V/he8B44Ln/RVqo3W
l8rgyvTOPYPdLrMB9nWDjtZRDYOBToVnBGw78HGLXxPHIZebw1MDF0xoA8aDqr5FxEQQZ2EGCreq
VvvSIY/Ivk4x0je1tET5R3jYi71rZyFUQwmCtGRP2hvkt6emV2NeBLn9zrl5mmzdXbw8ePXM+XVM
ppw0KlfIWsXSnnfrr0yWG34WSqTw7NlLS390u7hW5wUF/m0IM6/Ka82NWtPL03Kcp2Wlxq+DY6Wa
watZaZWJ6sTXBhEJaX7XB7X7ZpAwVR181SrsoZp+pp1ynfAxUW3LLyzWnb7nPUACwCA5T3bAPkW7
ShbTAJ80AghXAzlQK/6Md3Wi/WwGym9wVcF7Xsbx6kknJeGrFk6O0mOmCPzcgjDz3/T4u8W7qByS
Ob8AzDPq+TgxHEHbA8r8c6cUNyfAWCgeswv1IOnnWyEy2MzIOJGon6CdINwav8qbwllLW7BjIEj3
DTJwcJ2JQ7OJW/f0/0rHHi91Qx5M9gPfRy2MOlsHJHHaFbM4P22CsyGzk9AsbTaXh9f5BcjEZBUp
W6ajU8sW/IY1yO8qvKrykfRs0VzqngfrqJW8JUGFq406zbJs9d4lSC1czqgDgJdUQHQIhf3ZK/Br
Hi6Ecb9neOrplTxXA3fR7SKPla15qsQ4m0Lyp77H6FXLXR+DbjnMg34a2r2z8BIMolAD8oymH73E
T/Qd7iEpFTr7mNnkoBV972UlBNz8k7gHTxhjVOjfUne/b1BQL8/f2AKHMP8VQfiT2Nz1bH4Isb2V
xrIRQE2KzugLddJDXo/mkdwhadu7mjiqOLgWDdNVmwLGQ9Nz+u4PRCFW6kK6F9z5S+DOVq6DJNQz
VZ0slwi01uwwoMDaGNL0VKpT6E4cx1aQN7J3GRoJPtj6ulYZKsnTe8FUB4dBz7PKEM8Zwzr/xjde
ghATENhCDefKVd/uOAKJhWvmtYT/GTaWzDP7U9Y6ji0BkLUSix+jsGtpgoMo9Hbp14CdnXnAqiuy
a1jlqAN+pjPKDKmkHk5XdBvdbz1ble8s+xC6EP8JHE035QLA6c2k+eWk2vSIV34lAn7qM7KFY+T0
xP5J4Q9xAMcx2V45sQlGHw3E1BnTdSi9KeEDysPvE+6hI9zoirXF1kUUSgotVifmh3Lm0wwDpBEp
6aKb8FXPY+qmBkLmMoO76+tno8IGTF0keoNtNBRWP3yn+4ikMoHIjcDKBouQT42+1Bp6hVWuFmlv
w2D0y5xw0thUYZnZpi/iZVuKhJzB65bfTQMLnNN3WBS88uqWJ1uec8xP4LM6lSoTXVAQvp2hgfyE
QfA5ROaaWmuLsT7XhwGrINg9k314/27Sjchj/rgFgnAUHZlgbqumHn6NqE/zTvYlqf1CO8/o8ZJ3
bq8lRmg5V/UGH05Kr9YCrUILVImJcDkezKNUf63dsDAxlNDwFmibhNdxs964cwqLPrvplaqSuEDG
0rktWjuBdMXRtwbu79qk44/kGsI5xXk6CNM6dvxO83BmcC9RPkHed7ohcFSnWR743PVV8RYKm0rG
VcMomhcACSGhXmP8xdkkHhMuWqvXjqYJrRdn/MBUx8BeAKu/H8GKZVdH8o+Z5QlqfkpbTHe9ahBW
heFIlA7wivqTM3fVJSk+Io2bE7MtIbDiqqh1wrabonW+oRLDoTixHHJFFAhgBye0W+r66DSx4VfL
kFsCtgZyDeb1TYvunmLcV4Y9/IyQ439N2mF5sHTeoiRIeRweJMzzQdBes2mdwdPDLiZNv+Xe1r61
OAH7eQ0KnT/SpaFeEDjw0n2bsH8LdoARAhUyc+I4+rSWOXR3Vz75IibeJ5mV3vLeOCHgHVgmvSPy
RjNOwEJoBE9pO7BJhUyHIMyrHKpMGr0QFiaGA98pKKcl0dzkr6RGkgsu4r7xJKJWHtAf6ZIJ9Fgr
nCiEy2xXYSZBpzBnDKjbwyZCmEqE3McbG9mZdqMVf8l5alWtuebfoXa7xMfk5dB54dv956N8zANE
39VQvYl2G9XjbsGVqoOJ8G29GQ+CumdR/3tyFbBtO5l7VbZmaPbtFWTz74diJf85dDpESvX7MzCG
78TE+SX3ZzgVZti6WVtSFpSZDbKOzesncjdV1pIhhK3URgvghdue6363Zh614ZBTosmHshbP84p2
fwfiZ2cleXUOxLXZ8D8t5nPHy4/yqJNNYOnNe8lIyNKOsDaFUdsoRF4gwr5YGJTwy28IR4sfmu76
S1t9oMHxmCeabsXvpIiWvNAZ1LXKlX5GJOh2N3pV+23xwcY3MUlNfN4cRKGc4qDM7ghYatJUoKCs
Dw6IX3k8cDAXIhSCa9WFxscuqWu8D4WkQixG2az+Ipcr+T8wtMvv16MMfaC+FYoSSPHS8t0zD8H+
nVF738Bzkk1PykZ3LxFl3phowGwXIiHheCR1Q3XyXCDydggbtatlfRiN6HGAjBhotae9o7NpyJmk
GLOyu6eg1G9iDIDRW4p0Kg19PNm4A/8BhaqXTqOk/knJQMNPsdL0Ehe1MzaOgCVygclSwHymWqVd
e8oMM4qBM15ZeOVqIp9WdlWLvRbVIaOXb+VUnVwq4M906erbnGiXewVcomR4E+1F/3T90VnWu531
gUHVV9uHTl4vhz0GsdC3oZhqBPYpxrFCxjV3X0l7TZ+bKZlItmhcnQooBCfuD7jMb/iTqVcDO+om
6JqpJj/kkXtwyK/icw+12DJYsH5LxVHFowfHhTahhPiIteqFios80TV0NxaQdrf4X3/JHQpd1rqn
DyjlpH2jlvpaLTASG01Ieza31UFX46lxfQ14HeDP0X3ehBSm9waZOdvSFQb8CSiIN5w1BDZLQ/Am
Qt3NMHRN9fr/78EJftxhPD1fN7up3NExm6EodbmajXEkNDNMfWzeOt9TAxc4c3FY//rNyH+xtFHa
FbWBbUagMWItYbl0rb6t5tPTkKgI4wRUp+wmmOvhJT34RWmVxwh7aixodTEoRybmEity2O+Zor3E
rMg6Nb9p1AsJyLCrcodqe7uNA3x58J9Gs3sVz/P3aUw57BV6Eur9N0/tDiG/ddkGhqi8AAEHqt+y
dFJIuaWEUP56FDApsjJ3PKTBiPdF6/2FGc2sPIfhobKSB3ShBv6ZwnL3bm7RRiLpQK4kAOBQXJ4Y
bAVDqZMT/5NOtEvhWq+ozf0Oai4/X8xVtre8q8qm6voUNjb+AilgNBZptT2vKSbuuyH0MO23s1zP
umLzuMeGBvG408e9YnRgtVcSH1zi8dl9E2ZG12HlJ4U++H80I99UJvZI8aeM7EhtYjBlzUGHZw7d
QFd8d8/np87TXLu/DPvc2g4iNGsUza7wSZ/Gzk53vOUPAQHsiRDy7sFYCajOnpZuV7rC+Ngvg8wB
Zj7iHy5OYPCRlv/098ORMI4DGycToj1xp6PgIf+YWuKPll03JiAE0yN80Mp73MCxvWNru780h2QE
Mo8H4e8sESU49rrji57vi5vCteRzGQLva+KNV4DvbELauTUnzFjlKSEeoGskNqJESJ0XHQ+uOxZQ
z7lWROQF2D5EgFWrSq5xgyeQm81/xNedGJATAtlZGt3pmyxnTqmd24uUQrJIDtZk79/0yAX13HGi
9Kt4s/8DVOidkyXrqhCl8949fq2A+KEaIT6bZR2hB1XG/HqdPjo5yTukTkTxB/WC027+IRUf/WO5
gHiCiKe/vp3uvIwjpwgn61MPGuRYeo2vcMfC6xHD6esfbY8sEeU2KmYkSB6fCCOr9MjUW/rfnsxz
ai1qvQm7ZN/dHhgy27bFl4x3VDDnk0amIOGsw1UYzEYnKYOLjdS62tdYD1UVj0yNs+H9EtpOT7tF
j5rlk7Ic8gTFZRZ+A5ZsRmLM2re0uKFHTIsA/1pz/MPhuRFz90raww+ptiBobO3piBAiBJmPy4sM
Z6QdK5sd/CkIGoxRiZhxVMwYtBzpqb9O87xuSLm1qmBzCi1bAi6cdqMiKgc+OPzeB3+XbjvsK35s
2VrUZdVRPRMY0Gss1C26sHLberDTmbQ6NngzYNtGCgHWio0k3kvG4f9/INFROEbixPtxfh/oPX0Z
EdYbGKIhC5SBcmqwRUiGcMbWxouZb9gi+ZxBXndrjgyHnpVCY26j33QR0UXL2I3LHVriX+jImdBn
fB3wUAiaQq9wQnbZsHhcx5J/uwXQ3bVDIMeJjU0obtoOZQTwDl8RGnDOyTG17qxDxUObf60+LU2m
k7RtyHFqrtCUY1TbpirszojDUJ46XioBEzEQOO9/9eicPZkcNkrGofJpwNtdyeCx26AK1IKJy0Df
QBgcwnR1iCCrsQd/6hMYRJKHmBYZXrGgl3M/abndPZfiQLBUsshTlVuDV5ODmtkIpc+eB8itNhrZ
WoXHY5IeKzLE3mhMQOMhDN5U2koGrrVule24/LoZQYvuVf8xY1b0JfwE6axSQwI3AC/0tmbAENPz
+e4gujnF5xNOlSp5zjlIFWx7i7zmeoNV8e9kEKTS7uzjyN/1gKgWQU4HwXxQX6Kf3Ge4W0E3Kz22
Sq9Px6vfagfWjN/xvaPP4KE7f2snLSt3n+DhixCCJkdAMcM4XG1BHPlpES1A0FHV/y7Yk/3EPt5/
NSpis9s8/DhsEHCfNRn5oXfOuwInrVVFhW4vrayRfuEeMEzLOCpOmqnMi3fNl61L52ujEDL2GF3H
3I+RDK5bPpbUz1waTL0HhlV3D0U0Q5ZuxTEqsg6jJ8+pFKu8FLQRpVSxhlRkOEVjwjYx4UBVJ/1H
89vXvftR4C93/RDaOJtbKWZIr6PDMxWdJ2l/moKXXlNZrxxM8+42fJPP7d/iUa1tk0KhwZHW4pKZ
5qKviF9tLVnXFjQrHQcvQXERdUjdnJltVCeZMVL4b5FNGEX6mYR/AcAGz5T2hlE0Als1vEuZaQgI
muut/JG6F3VtBK8xTszE3MCtKjtZbHRjYsudwYmOzGwbpOKeqBMf739m2l25+68tVF58DMlh6iju
RyqJCDUH3xWdNOcIQquNqaRADHEzY+ql6az2CecNKbnOOr/evZQvyk1oluTgLKWkdbsLOwUdvPeo
8WCxvDDoE8aWMPGx+4vsS+ipZd2dGxOw4+T+kRb+xPBf0lAEV6CdnsuQsQDkKE+8GriXfqKBjjSo
ttUABI8DflZ2ucMO5r05OAMEEUhtDGLz/lta0g9VUwUOEY+ZcGagh2Zxe6b9TQuT5/ZOEiVFByxW
DMXNSSEb2p6hd6VqPjyioJ5xj8cpxiStCJF/D6N9afYPOsXpeOPBzr0Fy9vwXyAKA65hjpZUA10h
jbtY+kZa6NVscKciDrNBmgrzPkG2eseowcKKQbwBz4bxbvp4huekU3Kmv1xAmRzek2fIMkMlkGwF
jKds0KWRKh3MaAoXudpULxsn0i5iDAuYJLvvN7TXs4H84zgv6k1Osr77kURFHY6pZLPcIJj8jfYm
0AlyAreovtmsbdW6tHpkcPikK90BMsMN8r98hPYtPZahzBGd4vokPCJukQwIjkbKksoftTlcFqr3
ZLGPxFW6sqKLibGl8EzQb5zTMF7fbJbLkr3R1WBc/Q1xV7McY2CrsCjfT4BdFFvb3zLUcxptEzNI
E+8AFDtB6VaopBSmJdYk3fGG5d2EbSwiC2IrlBNplLUt+7YnJQ8/3F6MII+cns6Q1g++V3rzxtWi
+m8dyE/RQpuu2a3FxnbGPCB5K2MrGPdXJJR93ch9yWFx1Fbz57QYQt0brkrdC0z8BjL35/J/8AeY
kxF3ZAwDsEgZ6nk7PlVdOdcqgJ970uwd+Y9frbEkt5hmucWrr9TWZjvd7W9/SOVRi2a8JypE2Epz
+0Nd345I93gIn0A2j6h6Tl4HLAbdhhXkOA84wsbmBbWCLfUHviFTlAsCDxeViJ6DEA2Y6OlzDGM2
Jclf52NY4aFaNUuw21vx3FCT77WQ7p0mdjOA3fe+WFR5hcyF0DCydLgchDdm87OCOYsF4QbShMrz
9efdhMiOGqIsPundQJXr2BlwGfNo+ixeqsNYU999tV5iG198brAEBG9ciiRqGLf+0t7INmcj8f2u
9CIU9wW21/DDfb+5oQxtQOMjwfSX9SXOkCcNFBy6cCw44mlPS+ViuUErAUl6dhh260LXFLgP1ISy
0R6ZcuAU2NrT9j1OOQ9cThnIRBPxo+QM6fkTE/PG7TdFbLPK5Hx6ndY3jwh65nG3N0oREjF6kZ/C
pUm8tG2fR2kDCrr0i1OtPBIGoElZqgop6cmWfpUPfcZWrRjN4q/wG5f0BT1WjxUQJw1Hfwk6VtWc
7KIyK9HmnN10AOkX/ZT/MKpfjkXNNsmE8NDRzpfxrhhv6urk2bI9C5cijOHw0z3JUYdFWs4tYy1a
/01BhshkWwCghOC+fZQC8tDA8UTPivh2Dz74isfRfg/FgTs0H4DTEMe14W6Qz3rFqCosiTuUsKVw
P3YV7eDITcJkgea0GkT6kAbr8EMiox1Ar29dOLZIE0SDw+2Vq4Wp0gC9lyMWugkaWP0vp7fDFGTK
W4U0eCkrALR6LWqalRXDA/M82VhhXZVy0A/w4aYegYqAlGa2Bzn7CGtuRkjcA9VkA9T1j1qPEF8m
48PLlLgivRChoSreCuOk2BJx5Azv5e7upyWElENk/gVEx0DZPC4ieSSXK9VhP5A/wDyRqTTLe2d5
AEPGmHhizO5I06BTELphFUo56DI2JNB85wvhqwaPznyqmAVCw28N83kgqQx73mHxYmYJnQE26wiC
RV0K12n2poNHRTiTp+EbQo13qrrufzxlt/G9+AsETnDFeM93BHcEXCDOQCofwEwSUblYd4mU/uP4
1ZwgnyBlEv17J0XLDGdwq/SPZLF8iVuA8Ta8lSwAXSRnXVO7xtCdaC4D2+gqCRL2LQ78FXJNhlAS
A7xL5MVolyCMC4MNZifbffOyv4GwBezjJs7UBrYWuRTHYHtsRo2bTwzzQYYnGXs6vl25BRUObleS
K9A7btLmbjEFmHz5FzNYixSat/HePh1/WBl4IwwT8UK5RflCWy6Rv0qLP/l9Z4fDupoqCwgi8laV
gAG9d/o3ETOY8NOF8ndGwzn4b+i9bwOXMImKUuGX8mmu99k3O8kTuncHmJtdBCpyGO22D6JU3qLM
PAFePj7++xVZoGsYf7R6m1ZwlEjVWn3wQrkOzRMJUNGw5R75alp6Jf6HZSw0HTXcSKSPvnIGdeXn
fpKTOzCBGFDgGAPGodjcXu6QIkVxvbqTgcBaceHfOLvNYySl31nDB3geMDg7xGwzjzni8nrIDXME
yjyTB50YraV+kn7OfMiNrV7M6rdK6IqRH3XxsSxmeRsWzuryaNKnNejyCKwjOOTGEmH4njGRBCVP
yO8DNq4OI0x2Fa87+e9UKnI9unhNmiN5+vAE9JgvSkNL/No/GOKRU6CBMrO3WN6wdMsBtSAiH63v
xCltut81Aezbl1xGOyeBx7MmTMH6VYLJktNpiYXDz/Jva9geEXiEVybKgGGWrNOn9JbS/ur7JNcI
iFlKS0uOuBZ9bypwsfwwItOPlDyrffdWOfRrmwzbWNXur6Y84kNk7V7JvTVHIL8RHF60Ub5W8GoA
xg95iOURkkcX+AuwJDw8LFACJKHEo1ICDUh48imB8Hi9kZS6nc9YDyjanqg9PF9udg6O2hJho6Ty
stPzHBTnEtXGxcRzm2lLjB+HJ3jpUOuLQ01wP5wTCAYuvcdkHWISJMOiyExEfdsXPMTUwhOSSMDW
JUjnG39BYsJ5jyUnXODCj1CRCFX/dbYNUc3fNkLoXEqYyYQQ2v+DeiXEac4zVKk+jUgc2YNb0NhN
fDWvkjbZrqjtLclS15hc3n+ZLfeRJ+GqHKLvLfMHWmG0a8eiSMoNsCtlcI6wpETguDfzwFNQadQN
kt4kut5zzsc1h+vq++SA5EEjJBQ1SJlAX9YeaFX2AR5ld+XMPlpsTDQW/mBRldzASktxIAxS6XC2
8tkPfZDc/w+3B2/EPhTFaKpY15b8Lq3AaOJPLDT60fJE9z5QrcT23iIoiC4nCVcHBZOdXnOChRDG
04JdSIsWe8EmRw4hJx/LEFPkdTVns9Nj4aiC2w300BwC2+ej4oxGEzCcfcfavsStG5GhccLS3/16
xTjoTb1jYX+jSSUm7OGSLVdxvCKmm6J3vNtfk2f6J5sP9jo/Cm48t9uOM0rVMwYrJm/939GvVZXw
pO0FlvHHFmHRre83HQJGtyABOQy7WM0T4dc8Fb03eqfmouo5VQBybGWhfStplZq13O2rNyIPLO6W
C7ru5+SVePl5/85Y06SbBrNym7xzjVviIg+iHS0YbRt59qor58qxZ3WtUvlsxOQoUy2sYfZkibxs
JjvexcqH3BZ2HWV9HW1nWTeStT0qkR6t5n+ks8v/sA/sLfzvXHTdX+yfHiRQeEnsDMe1FH1d2PVf
ccPDcFcKp4UAZl8ivEBuLO4blLpg9LcLCzX2bboU6FRMSlAba+J5+hOLJWAhB9Y1aigehMCCbUam
HBcZpwFPF6iY4gk7PTHw17Ur7FrOB7W8ySnCF5olhZVZ7bb9qHp30QJquy/bTABXvc6fvUzDhDHe
+7SahrQQdlVqQ6ilt9seEKWu0fq4CNMcJoi/53mEr7Bmd4av1Hzu4IdIL5Ub4Yh3LTIF0B3OxNbY
F2qAqMIW+NkksyavRzvXgCw1M92NtKf2c8Hscndt4pKwDwJxhlnKHiGAk40SXW9VKHd//qinpmmp
ZPLktVTnl+jvniFX49RLvagl9tUVNpSNQlOe8sY/AEMiSlQCMAJETHHzYq/RA0ODt9a+Kt02GD7V
yE1wMBYn30tzJ8Vv7r2WQ961uB5CIo0QOQYj79dn72E/Rnw8jbsaJ4QflINkYhFhAJctsvI3YMDA
lptDSeATdTNp8XKQgguWcDPv3/iuDWDbCHBTLkRrkopRvvg0gsk90klPFZfO3wz1G5Ga+BSrYghh
5ws8LNzsCLYtBFFa1/HCcU733f4ax7ZXm90lvcJ0ARXtS+mS34JadrRKp42dYogLlOeWXEkZ5fvZ
4nKLEY4CWVogrlbk2BpS10jCS3ThRjY4iCn76il9Li9YNLH6qClDpmHO3aQIRHh029BQVfwYB3at
rfIjWgk6B5c4RmL5zIGRwQEprCRCfBH80uJvKDJTsTMXU7yyxi30JrJ7zEy39v2OiaQk8hMtPGOg
rp3WOAorWqtA5a75YwQTl5DGkH2tY9aOCrIFvNWJrfzTphso6ANcRG+Q2p36OIp3GEFdN7oODYHS
mtDSi6WdPe+x5ljWzQ9ME71bisfzoaGqeavs3Pi84etTSja3YlJ2Gra0+Vjf2nCYXQYcP9/wSskh
+PROOQZkxTT1cALEcqtLMQ2lFN0HSHlFhjSUltvP9F6z73cmRvtps0N0tGja5p3GSeFfXBrWvw2M
Lt1F6mgY8TQ596+j27EJEJm6PIBaMCsy1ZsrXz6xvf705onbJR/FaWqONY/sOrMtocxzxdiF6PkT
RFauGsdtqBV5cuCUefvDUQvDfyC9fhxWx0MzMVBh3rHOM0C6ehD5FFnfo+891JkfNI1CJOcHxpYf
k86w5LFApeg3A65YKE+DiYyi7Zl07RkNHpP0d1PizofFVXmG3s348k96NcBr8DXCsaNv5hvPs8gU
DcB/LfXqi8hGqM28M5OzuJj7ekcVs7Vr5peXLhpRW4kRMghMkGxHBCCsWpYAw/y2fyicW2AVEhE0
ourL6JTPY3AOcpHgJXvD7JhEZ3UYJgm2o5a0zhkgrSiSJ2dm81DNYWQEECD8cX72TBfnVvP+IC5S
zha/kYOpMUia3Fr7PvxEuRD0aIuRHAVtC37z+zREWjDvPSRoeWsQUuQ+JJW2ggysZHOcNDMKb22Z
EA267uwpmy5+wCX8sGJREg6rm0OUYG1prUJ2+tj/ENweagn2cxpkkllhpislF+I3dpxGrtgAXEiM
pTkXK8Muue7TlrisW6n0U4fp0kgua6mh4JqrgYOckzjG9UcYtduNZPFpw71q6k4xXTx6UScheUtv
6kQntM1Jwe+QjDlinmHtBvOpN2gs/ZoxbPu7yLqjZJvKh8b1ZKaz7S0tkGbI+WwIwy8dW/kVbIe/
/T3zO6k+JqTYo5vcWD6yhBALaDAFH+swQi2P5xGBXCS7XkrgCX0Sz/ClKMwPi2eSKXORNopmgAof
Rw3+BxaoH6JD92CFRwUpF3e7Ac0v9NRgaH7eDglY+vYzEe4+ANDqqytoTXRJHGPFoKUVHnCbiO+S
PTnFdq6Or/mQwIEMCcO6P9OYw2YyEs10MQ4SXeCZeyoXRlLPMoHythWbauDMHppnFTrfhkFP5GJ0
r2K5GT+AnehukQrsx+uLlVU9NHH3TyDLVJIdsYgWUtgOduHCrQ+llyAvYTexF3CsbpboXT+B5LDt
i85UC0g2clzTI6QCCUnLxsFnjKFNUfDKhwzAhqcDK3UYjum0nObpju45SbNuZ82/Bm7FeahRy/Iz
sAG43zH94gGU3kIgvSHX62dGF3dAJqsK3LSY/9QK17d0k+Y4m6MAQVMVK15SP/lqQ3fGo8GbOSMN
4/O6HXkoz7KJUGTwDe6+j+P4VrvSTt7RH3sBb8EiGYOL5QwV7+ev+LSYE35yXENhevTU5JLa3tZK
02QPpzFfJtWumOFG16RUspd7q6+tS9JRYGF/K2vBNPsyXEz9Q5K5EHf+iITpw+S3Zs3g1F+j3i6b
JhP9LXkT9ekr86P8icbDKfLFDx+4vE0ebB0+t/t9+4W9sSBF8TmUGCdnS7J8mTDXFKgb+uKa9VXd
JLdaK0nuCe5XXqsrpKOHBNkUic7//SiImDSKQ3F7rvBpWSWunE0i9GPC7iccNh2diIdQr+5KaYvU
76Yz24UAhSyJbLDvR9jo6LP+4iFKVTVRVuiPPFv4DM6BzcUFNYC7UIoU5+lj5yWW1MujSo/QTb5S
Lkg1S2YVeUIAvfezsbBLs6OcWw+rcD8Xb9miJkwRMj+3EcFUVgwQKT4IbXGpD/shV2ceYVZxzB5X
Gy24yuqE+Kb4ZpL38zULP28vhxMZmPH7GdwDz3T5MagyWvGmSJcys85qbmO+JUTWS1MEPx1pZs/K
QPn2CfLYN/eqt/PVbuBK8x6Qv+GT8Y1oWJUigpGdYzxjp/70NSKToJ8nGXQbQ/p47RVCqocdcVR0
Xc0KcOXkX/ea7s8rWxrKPSyZKBu08LzK9197HDx7naZo9RwEas/crPKSSCPuo8Ql9EazlMs4wMg0
QLmoqlIU/o84smQjHzXrvCMSAu73TrDGtabL9MW6hHmI11iQTnOrFDpvOAbymSmm70Vus3VyWSdT
+MU8ZpwMM04U98/ruHkDIa2PQqqgbZmoQBLhIYKx8n1w1VNaEU+xsGXJzUXsjJXKPyaocmssQGli
j/hxqh86TIOsXmSolIi0Ph067UgHh5lPWLB123hTiTiT8jWQdP+IfqAZQ8OrkQUzfYY6+o1+64CL
boqluwbdL/uGhuFzjgSPwLE968+eM5qF3ym+Ka4GgmsMngge9a0ZS+LUnWuyxnB65BLkUPw1O4b0
kvgqunbEmiJ2sa3Klyhva87r/jRxL+aZ23EGf4z/gYnOK9joVrBoaTj3PwDdggPOEGNTJkntVd8K
vPCTCGlEVM3NQCfnTmQhgSPBjOiRHnEUVBFy8+LlrWIvXhsp66ml1Oc3GT1Ke/6xNqbwS5S/dZ/E
ED8U7/weyKQF7b+3x3DXWQ3wE8cSRQ0qdpEedk0WX4bb9FD5eFvoN6cDnkmT011LQ8CK09470qF8
EVC/nmWcN1VzmShVKpqbZTNfFlHBNq0FHjiM37EOENgmdXD4Jm8lMI1cbhL0OVRjTFkTO2Rtr/Su
dPIkGLVSAT+iFi3MUu8wIe+V2wGqPIEXfFTixVSHw5JKRPoC1CHpvN+9D9anKp7XLnu7iKZ/40Zz
PmemB9WE6W7ymQYt0r+FIG1hC95K0Nel92yC25+eKaFRvzvm5JIrfv3TgSXVhsUqSRzYikSmb4gp
5jJbALiJoS9hWlwq43bugpEY9vknEP4nh0AvmfTUfQ1efzmNWFLcPh6IdXyw8trIyn/PVf3FJhxF
fu/cNa0g45WOP7mzi1FyOnwFOnssMRA8bFlSFgmL6zEvZuPltiLhMDNL7HqnE81TtUzHa58kBNZL
OKZJDovP1HCbEr9uJ/+U+/eDoSH1L7V/islFdQawK2fGIVoVcJkmX6XZL/3TxWcYlEYMX62zjqeI
KByDxPddsDrniAw6Eq/G6ECw2YlSVLgNHBGIcyMg2M1xU0hjbQL6unpLpaJaCBURlXe+gMiw7p0o
fQWi9q8R4fLttVS+95AZ4Wii+/KEQ/ogWyQEr3oG1OaToRrGqeb5MedNue5RZV3g3oHU+n/gc1HD
B2wr6sJwP7+CX3HM3gTKSwQCwHSpyihRfSvtCBJCmXakvpPvgzyobkWHq8TQS/EJWdmOcHzUXJFe
EkuKM7Rc1OILMxQBGMWHgU4jQIB7fYQlhXFlnU1d2MZfOaj9Ecsh/0rTz05cn6YxU+l0FPw2UODu
Fzb8Q5MkIMsH+ccUTW8j7Fgievc72h3Wf+uJXIlXcUCGT2e6YEkkX4Dfe5gG9GAopOIMOyo19KLf
XufrRPw5TKpniyCMsRZVmwes7odzS7NqSM6RLicsmqOCAUtwrHIcvObNNtpKcOBsopJqoZbzAtex
otHQ6Yrli/aNhcQIC/KGgFhr+12bcZkRrfXSg2fNzRnQhI2HkS/hyX3caDsVMc1yS3VNXasXAWXW
chLGM5iwLi0EhOEUEVPDIKdrgiWcvUSfNx90+jDVSMS3+zh99stVcsTNmkU+pkqNRCNZnYm5/KNr
ncDtOA038GSEqHYdi7hyRLqdmXJqfqHyzJJrqzVit6hp0ZIJZOKkhpwWBK4SKs9ZRK8cjrchB8tp
25beoNLyzhsgHW31jQcmKO1WR7DYYyvske/mPxV3nagnuFXzXKX5GwM/7avkkW+ZsPDxWDHkP6EB
BngS5mgmixpRjem4tbETstSU7pdMz/v2y64icibw8+qcYBr8nBDAwr1ASMiEsQTICVPw99Akjet8
uaKxcaSOjhYTRUPwOKs5rNzpTx2n8eivKxyDIDGI5iY3+WBxdiYY636OkQK0w0QFkp1Yj+A4lx1q
1G8ByY2wMW9RHu6ABvua93ebcjPMbAlxS9yOynJf8z0wPDGlFsvHpYLuWFE90RCcG5UC1QFy+fyB
2UANGuEJ0bKKsyUolmOjJ5nE4rQUcKtwTTsrHYx4/WzWAJMR6NV3+Rflxi1a9b4+vovxZ7ZkbJQz
mO5amWIg+DaaKORd7rSD2t5xnMozQsi8eL6JkGJAsRafimhQgAc8/eFE/dHqFTqoOrzXcsfQZ4PE
lbhdC/Wwpx34CwSlGzXimHkeNBJ1tWIyaB9+9prCxGo+T2941fCZ+ADMOEt7IH0IsZmXOTLmSSso
11tppO9NM422N9CpZhOTSrTWlWtayKYWDUha9LXCpBaZWLJ84BusQnEweOkwbKum94wSGEEknhKY
L5OsuBni0JPuIiD4niJm1pfmg0zZTroAYbHDKr+JUwKNnyOy25gtpArHwinFCEw7mrNJi+iTtP4e
juZ5ewJSR5ymCSOfSxy8KPmKOBtf535Dp7BUMcdzFZkVqsvQ2epQfsgy/s6eoN2O2/URxscYP1SP
ZOBnOAZ8Ze/EQWTdOpgikwDQvefc67yXza5Q8xad79R4R7IJmhxdhbGlWlgdjltSgzMKsmr5XElm
jmvy0czTeUL+zOjSGNkqS4bamqPusJ+AXw3sTtEzUxaNPkewDDsSMOUfHwQfAUY570U4fJvfFm1N
iQ1yjmLR0yhEYW/gDNmqUQJcSVaaYc1OHSwHjkjYhzqgmk8vmyRHIsrZ9G7zDwZ/FZd0TnUGLOHV
xTiCf4xskMQKLq83DqiilJCFD2d3FUe4rtwK2epPxSznW8YW+XeSW95UN9nToR94WQyTclo2m4on
wXp3Iy+XmcecfjTXUfxOMwa8RUl+e5ZLOXdtthSPAq3rsfDdadV510w3XeSJI/NNu1e9hCr2bL4d
GJgKbpprdufcpk/Q7pTwtDGjIuPGpAsv3Kxa7f3wRx2utXTBuWF26EGkT7N6YJqE/NsgGgNqAZW/
r3+C+uKiVqjCyXx+Jg5bXt1NQfI3O5uR6n2ehGzBORmk2VX9jCRomoNguEjILAiOkMz8jclEHgWq
KM9rV3gO7/FcTnAHK9zLB7GDsSks7xga6uDqXblupgqsLzhAGkEjVI2Ok2YcXo/CUuL1vQnpQU7m
XFWABzNela3edPK/OYbmFJb1ITISFDrUJGwdcldfpl77f8eUIpdTm0eh6ZImvwkYISN+Aze6KYJn
JE8tJv8bdIfQir5EClVxOL5uBZFMKBp7cosFOoY21Cfrk4Ic+zFhB6EO54PpTCdYSmvX4HvjrS0M
j9fc5IRAHoh11wvTgdc6AGajx3hISapLlxoxVQzpMfTdMSVLN28KgLGmLOz2jeFV0rjUj6KRrwuW
YiW5qxUkg6JBbNHVYtGqrpkiI7wdScPmT4wOnFN/kW9UfGKDtEMxsgUO7hNkXTi5BZ9pet8nDvid
lp234pN2coL07LIR1IJaPqLHHONKGuPNP+M/SPjUF5inj8ks2FYMMAcJdZrVmEUUdQdSZOUUCOF+
Hy9af2VU4g5/P3JW8AezRArSaKmxFvw1+0apcB2Kv7OcGaJHIDrUK48nf3xw7RarmLICXeYPdxaw
QNJSjds4egSIE6HS5+VZHYgPlvB1ixIztFjmU4X7Sdwhh4CKlH7g92JfANWmZlG9dhybwRDvzDYo
bhqeHREvsOySGgzI1RlGUGJea1BAVowgzI8VUpM1/8TWCov8vkDACz9oJ4OeCDvdgo+ZZQlDoT/u
DPFOLK4sR4tjC6qeYPuuldYppT2FIpmd5CIdCozV5sTMRjg2VjJDgNoTnabiLVw0Ixggmfz1jhRq
KDYVhqtXJcSevgmzSCDqiwBm60yznjZtBgZSA+OUOVjIktm2vi0nz0fxqC+FzIZNoChRdWdL/yEr
wQgmHn7E50qvCP7wW7imzznjqAAFH02NfsAte8eWgArhWFWvm+nI8INpBor7eiDqU0JkNSYhohAn
76qhcWaM9+dZfxJBWLpatUH1b3KWto+VrnpZBw5MWyPw3N59/LrYOPgQ2ZH3JGijxpD6Dikag/1s
sRRFZ7R5dGuEiuaxp46nltWcZMCUcYbUSi/F4RDmAEKctF5HTNVg1qnAOhuJ6KuGL0d99RsnD1ko
Vp670Ffo+iMFC83sLf6mECrDfcn8h2vkBq/SEovV6FkD5sy1u1cDD/fhKDYA7dV+Coout8lv9yer
qO5kBxojnH0bo9I6Nx0uCRIoq7H3pn+uF1TVIBCoTg+lU5704VG9A/5ztElPGCKJIUUpnenJI03j
r2P4BT0aejAEv+bzQtrtR5crDmaiNAi+4OO0/8SO8LcBnElvKD8fjwEO/0WjoQ1LZnLaDa9sWSmK
qDPVJMU10Ok68hM47u2BiVIFdtCJobLehvHC+HVAqouP1Mygr76ZEdNbZba7XmcHsNxZlzINhIds
udI9Amn7HqdE0tu4135oJtUCvXLsMtS8CLmbp9r0HDCHVemlrPf/E4P04hLfnKS1qy94KBn9QmWF
AUub1mVuatSsGc+j5HAImNl69JL0ynxnxt3h4pp6nN1dv4m99rVG/Mq7YK6A42/cOK8uknGdTKzc
d4uumAALYxePR0OtBlJbpvqVSEIIYp6Dv3HMLMWenum55PLpRO8mVbSyK94dsQBUF8l9auQwyZaG
p88F8hxv0YlSQCWnprJYuL4bAuHOYrxBNmqF/D093uT/c1M1NkCASSFmulmsiUS1vw3cLr86E9Vq
lWadWpoIaSGj2D6A0RYAMKA3uDndCHJ3Zao0E3rFnEnVxE3PUF6jIS7mJ+ecmXkXdngS5xpJMkUX
LaqfKv1Q0H0Ht52YiPwpwnDc32p4PxlLiOa3CIiW4dD0//mLfuJ72DBBvVmyqHVLQW6+DoFPxIle
i2SDe9gSjfS5SsqgNVNicDfM3pXWk68gnEui+rlyQo/cr6OthqiAQ+j85V8e90XY4JYuarhmzZw5
wZsOrS3fioa9oqMXJoqcHm18BVUTvZH4Lnr86n5Yj3bVqglZDPk+8o6fnFRx6TjZI6FN9bN77JpI
kCGEYZLZ670YsfIbNspKN/cBhEoDbURJmEzcBcM0kqh0iFEzHBUJq1HyaUPxQFND2uiWpGpdoYzc
HyDkhs0gIrzori580xSXfLqdNhc+agz8gi+u8cEm3HaakPbIxFz6z5WetRy7B6Mdu5mRnq5OpQVA
94u7+3dLTVPwwJgMBV4uu7yc/A3uj9WMkKddgPM2na60GwvnD20X7C+rG4jyVSfrWhH/1TMiMPk3
ZAtYNsMuXDTz9lFHkRqbqCZFwz/0bHUNXn4K+6yl1plSFOhmL85wDVpLjaSTYd/tK0Qg9V9ddgU0
RDnOKZzBcfjCMxV4+jZaGYJG29aY/O6I9FUx8wzoUW/GOei7kTwM5EaotwWd0MeIL7X28ESgrVLX
DNFGPrKooYbFxJmdlDxJWutyAET8xCzVlPsdYdophDHTcxxkDo+MTJCaT1borDnq9Ikx7734+KNU
KvfZM14Qg5xajuHu3r1rfLt2RtkCz6kFP7hY7at88XpiXVBgBxNvcmXeHsSDV1/BEWBe2it7FguZ
WxnqLjlCg5Q9ZTTiRCxzsA+pIaxe3VD8Wllw05XQMyhez5HfIKLtIYmTdhzqzfkXxot9aE4I8upN
ppkIX7celfJK9Hspma5OHbgKSZn7qEI/q5EQJfEBAbDoV3YwQl1osclz1xjiWn/cQVi3s8g8ECck
fUSvoi/RtdfiG7rQ8wMBogbMG0CzUFsxfODCiBpKCi299wueX7W+uCqPM7YeVd1MLlssh0m8R5yd
sx0aknaNwF0xuOCBWgKcT/mnHccOPO5epZ6dLq4Y+o1oY0+318r+L+aY++zDVtjb1bKrKv//atU9
068P4Ly4M7aenmpmyrFaxheBemAHgkSEmfe0J3lL8DcBUoPO9dJE+80hx+BEvLll7nPE3aLvHeC4
SvH5jWWJcIqSHVugyjs8u30BjQdppXumHn9YSXQbYpSX+plRNY26XnwNtegTHogJabYaR45B+XQn
fI3a8EjZI6K1O1nXUmVw9JsnsRxOjaQRoW3+XitkUb1EKhL4FznqaeBc/KisbrLx0WnuwdLB1EuX
1Aa5GSE7XWi1hFdSz9TmQ83O3wNIwdlEauFYnLAGdYmLpWKSHPRBVL+33oEYjrXlhBTPfrv29Mh7
zwstZC60yH19LUM86aX19kDSvPqxM+hGorckcfXivZWwmCIIi0k4Cm+p+j+nwVfPAxUTnTmWBRCE
SWD+13EYUwd3AKcEt0zvrmo3EqhTFjvpDBdcUs1Ge16YdkZzL1KhPS53Cxi0NkNV7ufUGUk2XiHY
shFIWfhMM5O2Mehsy7iiD8PgTMf+1F4wL+YLpTRK01t/ls5eCnVf4F0nEpT1mypRqeYXWueJLEDV
6VseW6MfpqKWSLQxRhZG4LN3ZpVQkcKOp1AVR6sYCPZMZoD7Q/TLt5DaImcFhz/KPP+Me3IWcPB3
E6mGGavKzMyZEzP7ZMGS5OlwdJQFiwBOpJjXLNKR1BcCXxSNQDr3ERoJg4Gxsu99YPQJBaaneXmx
fSnuOj63WzGTcgcLZ7SOS90XSWhIkxh7XidTvnXvXGR0FFK1IpYyBAPjSblx89ZeyKr4Rs1yPd87
agrwCD24N1cghKhQsuhTbXZiIqmTJxaoccc+ODZZTk1ZW1nN+bWM9q140Qj97akfdv9MOp4pdSz0
FLuhWAAH65jrggDiqPZx7tPyBOMHTSUaIlCm5nmVf7+8E6v4d3LpLU548nEbLxYRqdGzb0R3idVl
YWDmgt3AeLCyxedWN9UP4XqMfFttA/eT0ujT5pyMplXvNXWBVjfrgeYj0slV526jc9eYtIHwwUhZ
c4ctPzMp03uEh+p1M53NMaLNxmT7UUgcMMMP+QvZWcd5s9ovc4HKsX4Wpg6ZJl/u6fO6b2UB9sM/
zhKQ8pVAlVSw/ui9/Pu8/JSk+nb0g1N4snSDaXl8uqubwpkHoOTeuIL3FFzXuBw+vsKTfI1PrUow
QLyhLv5gMm7hE2jmQHWEph8TRiBz1uJcAQKrI7X1nlCOR+Tn0YTPkdxQDwUkQjXx95oOZ6zfaQcV
PbTTW0VX40ShWNKIDUcTY7DGbVsDYCZ6PG2UR9CI0Py3u7PVa1WsTo8o8vA5XGeY94MmR2XDWqMJ
JRuSZ3VAVggJ8/9DQcMrod63v826Hc0RmQu1zs6VG+AMCjC/nd3ilVU2uqeLQWRNLcoMtRVvcVUn
TyteeB8MwNxSgRECahYYvWiG5BokByVq4cVKdKFMBR2ZRDsxFtI4ENEaH2E5FcoGOIaU3zlXVLkl
zWatvPjG2Zryv5odI2bIV/5zpfLUkaPSdWMB/Nx/a6OExdj9hyrnTDyMhB9w7VWhQaAFRiu2RPki
VTumiweErp2NpwX9+rZG9T1Tg9U4qf41psx7eS6bguGCvvX45WGNqKQo/UgcupzqFYw0C8VU8uxL
dOlpiGrekYz1nbWfwIG+lYQJthGzxKrmam3rDxQT2DqyP3FkbztLb0CiciLIu9Ddbkt7XQZD274D
A+d4x3+y57+Nv3w4nrw41wpy5zILgvRygzdc6UIzDY0F6bRa1MO4yK55p85o6e0+k2r99ZF25yVi
tkzlCuWQCqG97nI0k0lJGL7PjIYt41j4sRV0N6vBibddKHLxE7WuSvc+1JHSkw+7871JqKKtTa3+
P4GFe6wgihjJebgBLpXIsDK9U8erLqktQPccEXXH3E2OXo7/NpiYiF9cHVnNLvEqj35I2uRBjbKA
ZZRTVo+FX/Z6zb4LxOde9pqmvqGD5s6eIXcKBcPFFCVXFMIZRYsXml+N+iifEz1r+dkBgijI2Y3y
zr+6qke2bAsZBZUzw5LnJr8gWzu/iH9U9ZUAcq1s60Xai6e6lQsShjHls30kkcfy5XS0L/EhQBCm
cPHKFTRFreiC5mRT0D857nRModFrNF+JS12emVS9iMcby/1k9OUB9nk8PSEQVq52uYgUk1jkzBIK
PBaNoPzHaNG0YopbuRNisn4olDRD9jkXXVkwTVsU+4Yp8Fy+J+Y+kprmYLN+UaQic3ZwLanHyez9
USWWK2qJ6sXOAFoLZs6JOz3kGb9D2ot6K+EG0urdUDMc2nSAm++m+2HtYCAzO2nHNw5ydlUmmUL1
43MAG3B/lBCWzrNmMpo6LLyNxJj6Xn3ZqkzVNfuZnBvos0NjymqgKlTyqDas6ZXHvFPECmSS1WN1
snx25mCiwCLd5h6FPa5HDyYJI2HkWUyypQ2hy84RPNHkIweUQiENJ+6AZOEkDUbfOI8mZu4PZMEg
cXg4BnBe5Gv+T2ZwF2DvtKGNk0h1uuJpeMsJzLI1xcb2tpCSD7Yd+13rCsnwYDj3AL11DXd8o8yJ
Cfe1ds9KR3L9B9/Iy3i/CJBaftR+GO8pSd+V8VjzLFlOFC/1XITbYNu0NmL8kuIFXHfLJb4qrk8f
QH8rOlIxb/QI4aqUB/SrVR+pBMyJcFszvSMM03zKuztY5ekHl1OjpoO5kddqHgIAOKkSV2AhZEbd
QnfhmpcDDezCXuWwgDPCQKCwZtPEgfeJwdcN4ufr2nQNECgNZ+xtpG3o20qvqfKg9o6XMrmJx1o2
BnAe7kyTlVj+GxHZKvlYWKlBaoEE2QoN0k6Dafi6L7W09fcPZm+CO/DopGOrtAjyV1bh22bPBpEf
iVFoSHM7KlDFxVD7+LHOYvGRhAHivP1+9EGjw/8fXvV7rwZxba5ay0tscs5H5RHFpxU0JolBkYeN
i7bMc7Zc8/EvQIu0H0nQPr1wFXiB9hdpjIL4QGRTBIR+jfD3GR3iddvp1B+x4V0m7uJMAI44dz9A
LPzyfQyr2AGdJq2jMc78uwi2QLD4gL9ePbmLKrWWAC5RCLfe6tDvvKYDbRjt63dNSDS9d3w27Usx
d1LAeyRyIH/6Ej3bOcs+2qNJVLHDS16wb27//aYHOffoRbmXgDQmsL6uCFG7lPX6iFl5/sGup2QZ
zY80QqEouEKNb9Xxds48DGpwm7F6Fdh35nrgv1wUpKABYGTenCYPV/xon/nKUTHuNXO6u3SvNC32
SoDj+B/k6svmR9y7eG18G0ZEekzR6koRr50x4QMR3d2V+6DWjmUZ6rILZ1HbFmdSMpvAUri+TPgl
ABLG51FUlFdjG5M6uBm/gxhvHCFd6kjP0v3xdjYMDFsjynaWnXSkst6ZCmWpsvw5ytFW7b5fVICC
QWByK69A5sNdRlYYpXD4MLocYcS7UlA0aeAFhLugbkMC7uUESXNLaIlUoygZ3/FbzFVJHz0eUIby
vkmkIqYXraJvmEpho/Luy8/3V9+uXOvQMwnGvCYvKZH6XPVbeouci6am4WnXx7cW0GF+mcHe2z+E
SrJd3dAHnMqd7rK35KkjGv3EZiTM9FFdPQMMTJW9lnnBTHusMESY6a0JTACwFjv+Tog+bue0lbx+
NuMSTCFjPB3mAfsfmWwMD3tgkTQ2SC6uF5meIyZK4quMBwVld1tihlz4qBljBpdz3gHn2TYzR9Qq
Lfk1wHFgnFC2K7hnvyq6DYBan42d6npRqGmriZlMCVNHk5XA/1q8SMobu67niRiBMHpbZoerwzqy
+eWd4Pt1+SAsX9NtcpofIwjfXr5+DT58c9YFPbIu6fCRRYxQIvAz76Kf6ubWdyZIgcNhMB/LF/JG
FvMDQ0H1v4Jm0sXAQgeR+pgrdPJubRhIoLWbX7pqeAwuxcZHRRqN+NZ8FiTasZayBZ8Zr5oPfxym
Havd9t+r20PYuorMs0TW9KVZb+lbNvVlgj+y0PFT/ZNpUNIjziDjO/UOCKCZRlsE4PBqZgNV070f
m5Iy2g9u/R1gyg0XmpPey95Z4+BXIzGBvuYc4bN/Rky0/GEXrgClqqFgNfVU4jwEEOjwwt5iXaqD
i7y0j7sRVUPlUSn68k1sqHpoFV+Jz+oAevkq99hm7Ym5LpWKkitoGFf38IY2W0Ecci92MMeODIo2
nUbSpa6FJIzd4Lc5dmvojkVRvNKdoxOHgrDNBxHVvHirxDSbYVA9UiMIL4yWodked2QTbwauWe5g
Q+h7DNQ9VDp72Lf3rBPOPyLOrmWabi+1l/e3zPORIxsmfvel4YX4BxozCnrbP8fgi8IQyxOP7NGC
qoid7QWU5MfAky5EZDnmJFlphPI3hhZ9lTvkHZqIv/BxThluNlo9R2MJRevgQ+ggJZt49aZEcMI4
EmvELhQ7yFh68z8GMSBLizJbL94ESHMWutiB5WRjpw4Vu4zMiI2M/DFJ64EekrxEOrMi9zWfFr1E
9UECL6vSAx2OZLAh+TyPv7EEIwxepegRnJWWXYmAxsD4WvaMIbbvfHOPM/QlNehHz+bUasTQBzTL
LSGg33Rg0OaT90SS+0aDL/fbUXRMT37h3Mwl3AoE1RYBnLfy1EjaMKNmuB9zBvT0h3C8tbWoJVHe
gghcWJqi5qHwZ+d0wy5oB1QoH22/AI20ipkyyHlgGo807KMgo6gN8XqZg/bvbd0HfSC2Y7lMGoQR
FKf1pCW8yIu1gXDE+/Oi6BrZ/40jcKHJ6wfOIEnaMvSfsXA6LY2UZuwVOXWCfHb3yj2AbJyQ5pEQ
okh4yziXtx6WMBAhDKQ1SAgtYq3PJvVETj0oQl6zFHraCC5r+59BRMNCK5yL4RBNzcAmXYB5DOlL
gGDvMyEBrZxZezTydhYlJXR/EQmlmiIKk68z7xCB/2OnM7FrirgNNg1aynpM5Lg3FJFqU1C8fIO1
QStpHMxlTxLvByApuH3fhHbzdR7KBqgD4/0F7pIHmpCp3e9g9atJLiTKfnYq6wcF8l60UvQcDUX6
rMgBW7P5I2x/4QObiaKdVZg88B2rG2EP4peCl5dLXqtROJbm5yWvilB5AIA3jYdBuZI1fOGb+rTY
tAZ/w7+bplA2fuTqHlX1UjdYnclZofdlqFPGN0CMdjyKiFAAD/kYMesFEUpgOwRTozTTVxIk4FCD
J6IrURz0+341A1DBXbDfMJULvXT0CKtw3kq7chjZaED4xmDDsOY+lJWqEIaT58B40mFVt8Y0CQsb
Ns6ZFBz9pozR/CJb4e2hfE5DpImcttowiPOvJe5RFSkxJMuSNzMgzecWmk4zjoDWYPJ1zepmaYgo
ROQ7RbcFnsMNAGqGHoFmxZMQNh+ADkUdz7lJjRrWa0HJEqLNyw89ReHNgcYvxISEeJXurXW3ZuSp
RmZIA1Dem9u0bfPdla9yQta/393VTzGvYMKJ8OT/mIFi2GxCcD2ZtSPsz3Zc+ELoeS4+WDyGmhu9
7I2MJvup9l623KadWboRIvghDSohLGw/PwkEPy3YpxzzlJUKC5b4gS6BiQOrt3eDkmTRNsy2kQ2E
2STYRL45eiLqypfeBkAm2uS/04ivA8MO2DKRTya/G7B0hdHNU2XE903SNCJLS/+SXzhl64cr82Sz
rxUQY5nL2BC98iU1Xo/ug65A/Z3A0hIpq31fm9cVyFt29YWlisCYIZ6ZQSAI7XPOrfBe+o8c1RIW
ZsLrQwCGS4bw2Xnz1dErTsH1VRbpEzBRw4tlYm55Eqr7ybN5OnWNAGx9MvGH7J6keBfcMVb1Fpnl
v6wHre+ym+F8ntaXoFbXWKsqd5aXOTH0d1Fw1brJJflr7RzDi88TqU5QWmAm2b4xz3cueWviaB5C
UoSNhSiRs3YV+NYi3654v5CK4dFmiJ4n4VZUYLe2gFqVqlSsnBJNPV7xdXZNcTv9jdb/UUnCmsCt
B5PrthKfu2QqDjBfxNhKSvWAH6hUe2o0qzPVAO0DMAikuZQuab/VXkmQEVeAjOUc7rG6lGcNy9lN
Zg8WXhndd5bWUFhnEYYysx+hZS7JuL0MRnbfEz/qhF7n+dNgfY1M52pyP53waQhdroym4s2yEQIH
VgeK/MHQ524r2lXCTEoAwuGzO8g7fnMU0s6lSaXXBJE/XMBkVFOhACm9PJL2Sy5McpA8KpGbHCkj
9eKz376cQF/N6k2QF2yztoUXbxdrY35adt+QgtIF8wia8Qcm8U4aBtyBp4uepC2ANLvI4mUQ/fhI
mJqWHLftNIfL5gSbjDX97+5gmjVG4yPIaM7xl5Bj2VEQRbBOOq/3hO8cn0F6RLYL4TAkhGBf2/Km
Mc/yCEpgO5MI47XD9srCasCoTg0IB640N7O0vO5Hn5JPIHWJGqqbocAkZ22HR+7htlfgwup9+ciZ
XX3zn2SI/4ESNak7V+JofTMORR+WaV8UR6u5TcB9RFijjHCbdX+5Z8Rem++ZrnacVSOjFH58qQtb
Cvg+ZTM6Apq5XiX2yv78bgFsWsaTey6lvbX9zEQnOMMTmwc68r/Z2OqIrJ4+wReOnwbCZ5PfWOzV
PsgZpLLgWJ637jI9zX3hTfT6qIeDdzlUEehx+8YhPlpMNZxt9vNB93Wppyd6AeLpKkX7/dAhDOZQ
jRx3rjFy+V5z+gKfHoYgAJDklrssbfug6rtPehzBHFeS9TJWVM+t3Vq/V3SikGPJ9bUciPEjtzfm
SMkV8YQtqmEKba0p6DbK7cKsepQfTaEFz3AG8ils7OS7hIrBCPPZMu3dWCzJ9ruOl9h4FX4PHqAj
ryn+lsYN6U6gkn624oizTzdrK7zmM6IvaxicA3U0NpFL8FBEAOYxDMZX4nd/H1k+K5fAjBaLTY/O
rz1dlOAklcbrjb2ENgOQdm0zHdS9GdhKZMQOYn9P/w3j3DDg4mBZZF/OmHMUU+PALTE7zwuyRxVG
dqlXeI4BWw/AtI/gth8orymAK++3V3dJK4jmPM5Mp9LUyj03sMOY5LZkuV1a2J9pr1fo1ssW94JY
x7rPNdk+7dZRaGe8eXXCs59GAjf5VICLyC3kaLXlfrs8mXE9BhsyUtZ3nQY5X0kry+tbc1doVa2/
3vWTPlx5noTBHlxaK3csPsqLy5UhytxWStwGUwMeCC4w8yZIvesTtwhg4gmM7AuxqqGqbcCXXix/
IA+MBHr7/zX7TSjXOQSH7toGYHPTxFLFDzQ+SP+fhkpyBL48/0eoDjyaMnffcVQVE/BqE2MxMvru
11Zgt8TFo025W2fHhJ1tArolPFI4Xj+RCVQcpRANENrWKJNJ1RLWNf5QgPIbeL2YImffWGqL5Ogk
a2cTMEP7/vchw0l2aML+dlmPgh653uQenXQ0dhJJOtRWeMUhjLo1a3B93wWi7aAshsGjJcm/Djjd
LHQlrMj0EY7YIXE1O8A9+F3pdMMFXZur1+DedUNyr7T8S5Bbrfg+NKG9LguTy1U6izWPdt/JYo6E
BqeWSM6becB1Rldn3ucddAE54j4qfbND1n3FDa7ASprDHgJubz+WEoPoNcn4ZdjotKtAOlDJewVZ
dRuVfZljwaB2iTnVk/q9x88i6d8FotIpOwH4t1fk2jOeNDywR56YOEzEt475glks5AjTvtOJP74B
/x0tSFJ0AcP+WthgoNiVgzGmLO4JslHjnFzuJR2dJWjxyJa3lxLNuZH3y8iC9/fhunFyCWPBYYwv
bjGpTQJZZxEoOwd9JDq4pbI4ZePuxK7wdc2jjthMgNx11oCwTyIMB1Z/FosT+RebuvxxyNy5Eg2S
+zVj7sarxnJdMtUWge7uCFFjuZDJ6jWAmxHtKb84/iDfiQckXooHKa5k/zZusWRCFqHZ06kG12bc
1UOkDDWWGK4JRYMA6iIzBj1Fo0CoEIUymdWr7QUEniBGZ7K8b7udIfXHntw5X8i0fBh0+A9KBFcx
mrMy5joQq69pKATUQlRKga9TM4+sWJ9k2+DjmZSpoNi+oiVZyYas3gQtjSOuSECudB3QeQARBFXB
xSqy+s9lJ0d6myMy6GukMN0Z+Pzm5TpRMGgKICt3a1TtpJlsp9ESXx01vhE8UvbD52tqCXCXK9vU
bvdbifZ+VZZc0mBwEitIyqT8Y6/MITiaRt1YrAgZAz9PdiIij8+w/B2SChsNEpm36sXoLFgVDC4E
w/mpTJy7c1376z5IkbLT6+wXa8GpQWfrE4Xe48Pg+2OBoZEhDfpXHQQLUSCk0oedImtMPLmIz3wx
CWcGIU184ZbGd795wQaoC4+o6qRfJF7p475A3HJ03S+du9qfQsaWyZOmxX8Gn+AENqpmbl0f4zQ/
xFGsvfeMZHe5Bp3u9Bu6C9KqNqYTDo/uqw2FJqz/aWn4zRJI7WJhPuGipjkBDD0BvBwT40Yc2Hoa
l8IlLeNnvZHiVE+uyhJoSeQQ1cNwRkIcleca7Nh4pqPb/LVxnoAvqQpUMXLwRCgJA5OeF3R51Ns3
bQdzI0raWUij9cv7IHK9ZnF1x+Z7dhm69Lf5a/EXMgMEw6b/PWWSaQhRqp8+vrcURTTspsxHo0C1
FL1wEkeqvokfwy9aNsgisBDB/4aUC/6NZccDgu57NtIqyjw2IWX4e3uUKeweOw22NGlxaCsRhgnn
5DeXHVVm/0EB9X1VZAJhAMdJn3jeLXGtK4Qig1T3hqQPeiNypSGbMVbZD6eaS08kWjL7DQsBJTfB
D83jqNBzT2DYm03aGBS6WVT0EPunDJRAiC91id+Fd+JIqB5dbc7H2eGLukEqh0RsDRr9ej9ld8uP
JlekU2fjrlayhGO8AWC+UZmEtqtVr2jpZfy3O7r/31zx1YvrO0aR3EyqeoDskcRUZtiUXScUkvi4
ngZMjEu/+pQb2n1qLfOF7BQAYCLjwvfkdGSxv2VSTfgULn6tozidsujlJkL/0pW3NAkNMY8T3Yfp
qxSDOOUQ5y2ccw2Tfft1EKHmyjo1PdVGMGbApstrp+Dxp/mKcM93o4roDEvqUQOzgoh/6BflwC56
KppGTXA6mARCH+AaGrXq432mFkAUhlEi7+r7JWYEh0tlUAK9bBCOtIqCIgcrnmBMP3WWbJexRob3
HFPUJbnj0BnOLfTVFZfPFyeYC6V6cb83nNpMuWwrFxRbsP38WI9odCcWKKGmNTmpSe3A5gUxZolQ
/q2yhz+e3X3MbXd7i5bvVNUyBVKySxxLzy1OmcK7inL2jrXrgcTAZ8uL1csI2Q97aDZ1HIt2ihjq
zMWVFw581iODHiJhircs5f5cmP1EF61OAOWfPHMQg0ii0ryWLjDWtpg+YHEgU6zNTcDVVSRmAI0q
iA5BRxCTF18i+J4+5z/lGspNopo3SC4grBO5YDD6SdRlpzf4HVxpL8VjtshkGyCTh0o3oWUsMWu9
adg52DlE/ikjbOpWay052iujtAgoTy3/tSOF/oxhfisfd8s3GRia+BMTV2XMwR4J1rS8q4ypCdRk
voJlMZJDZZh2wyjBz7c3tRS9deMgxINXXnl/VvM2bE2NtnyUS8+ijjKBJFyqZMMNzKIPg1PmIqVC
owjbcBz6sY+664XF2C8Z55okY6OUODFzhFBk6yMVAmKI3h0GHVlNvR/IncyZqxXPGov0df3Altoj
SsOPzSMzayJKQ4by36rfG1LKir7kESmBQHGmC4uUlmiEATu6uyCeoQ1nn6V4LHsiJ7PEwpriuK/S
LX1cHfGvEly5YjuqCVe8btItSZKvSF//1o3IOgq8Jn8GNROw8cjAJMoIG8beIl7wViQE4DqIr7Wf
0uOPEUUxvBXGvrggli3aDVq0MTDVT1jJ+Lpx5LjYCkyfmG1c3nOOD45MsV4wOc6vbN8bz2lRQES0
SqXGZANKEiBwZwwuycrYmowrFxyJEFYa2OoRhHZiopbbbu8oJNTjtK+QDPEZzwy0Hzg/5CuCNhMX
i5qyxrUOzNJgL9dbbIkJ1RIt/779PQL6HFx06S6rd3t6WaSojaTNDlmvzWF54pevGtY9tKXHr3Sm
Mez5j+D2NlLLPYYgGJTReIpihvT8kzbXyuTItcJP81hwI1jA+LuElVCV1q8Z39Pc9iJ7CIGQUR+3
2eSp+TeuQzQJG9OYUUDcBNUGiUruDuCErhdRbKKpOGsZQ/E5bCX4EulRVYTDlxeGFekkQVQdKFWh
RLN3fqHK6sdBZOTK13LzaTN3mBbXyiEbPbXPn4EW3gpXY85M7Y+UrVS+K4XZpuKHiwJSJInbrM+S
tJbZJ8Gt1FElUrSzkJsEbrTNjJUMQRwBuWM8RgZ9eY7qkBRB7pYZOus1e5dner3zmDkehL2p8LEP
Pd7+mbuO/6t04FxUmyVzjtCgxy/8YiAylQ+UR8RMwnFdcgpsqpQFrLlVZR5xQnFa7zIJdWZ2i8Uw
qXWVq7b7N71QK6FZNUsChGTRXj4vktS6F9u0LSAC62els1vZ/ZVqK97fetJrfX6+V9xOv7u1lkln
i968cxax4ORlQbfMT1jqabOycyWDYWtqns+9vD+fQlGVIthoSYC/Rz850q5fCCH3hpkddKix0l8Q
87v6mPn3sW7wexvybqthhBlryIdzxiZkGN2gJfouVsIM3TCpCOdny6Qka+i23cFsb9Ffkb1HuyQi
M4Gs3nl2FxE45F/3FUScSiM4cvU7bYGMeDfd+v9i0XZJcAsNQ42WA+svwH9XHb83WxiLN5m9Pb1Y
eqCv5HHtXlPAeGKyJf5ckJri2ztD+utbP2p9Hmsnl8NxQbULWaVO628NXhefdVBgiDAPhFbgbQV6
1A5r1+wSW6zwyac6WISPvbyZONZCbIz38kJa3XEk1fvRHFo6uTeFnEHGTvb+pSTmPmrSwHO0Fj7t
M1J5RZ2yevanJutpuqrQ+T+FeALLcM67RjUqM8ckCcAxSVeQUWjlvUQjTJQgJuIdgDoDP1Uy5Z/2
+IWZbyX2LuKtdN35oLWHKz8t/AAe1bvaePtZjHGcV+uDfJTvaPUkTUyOmvuDVknqr4T5YKt19HV+
Q6ZMG5PfZAwRfmsCPlhsyG541Uz+6+U26way0ZmT3CBnM7sZ5nOdN6qpwGMn0GIaBSGlvQxpeOgW
FBjgBseP/jb+k/NEDR01AbDFUUdoX6eCzbJrdW9rzly97JQSR0jPaH3U8hHsftB/qMCCTHDlt4nW
Dao5E0WtDCVAs3qPFbRxf1PG12Qa2seMUK5zrmFbkh0mwd9lQzFk8dP+vdU0k4BJhsZP90rjRncN
c5FNv8rl5EwW9u0vcSTlOr/bbc8+WCRrbLEChKOyn0XaAGhhZ8TzNKl6XE8saRsSXhbCGUiQ5k4V
MJd5/6bWZohRzdzvLQKs3RE997qbTCIXUhhXxbI05MtqwRpuoc4R1D/J/h1R/wjMchFOqv8kx0Kq
CHHO+RK7bGP8yrpNtztKkFaxyAhX0Ymn7iJOjdkLFmoMlH99711XNLHMgsjHyrhV0XH7VgfurkRq
e4P+ZUwpF3rXRGZ7ABHIl9Oe454BCien0I9FgtN1ESXN/7oqNLVle2UJPfkLGgunc0Sfp3PrpKoc
ThsjqhO2LbQuw9v9cmnDfROOP7cNyQYP1gppG303je6xPmZzlvq1U4j65nVBuLKBVS3KcMY7t1px
W7B/ukRyR9gqZM3yh8Vy3h9FASDHHk4n69m7vJqBbirIaIuUejlwLgYfH2DV5FeEHup0FHMq2YJY
xvJy/s2yIexP7rzyOxA3Ikm5NFySfGhrKKqxpg4uUMw/NRshdTzWcwV5+7AxroTHVajmHUHHMNM8
DYZT5GDNwYx+RCyt6c56ETZkUA8rODmMjyHJy8hb3qRLRDjRP8LVHVsJp53rz91E4OZUaD/9NSkH
ESoo36NkjOmCBAsr1FDOAsjhhL+/tV22mp6NaGKyhQM761lvnNz0nfzsIgB+PyJWH1GPEG3bI74n
M1+JHiPVeTetvDoa6YFRHmJNlGBGSYoZ5dX8SGjaQ1NUxC1SzZqmd/0cxaBF/NdFWw1LZ6PjTJfK
Q0fTS4uqC5hXVYcqlgKQoJ7fJzX5hgJgl4EfQwfAStw6MazGYNBJCcXbxSPpvbljCSoSybWpTb74
nhucmg843UEaZftQZfOQYM3wed89nsw6qiGHubtQxfPQfdvZkGWVdzyCXaAOr3blhz+KqtoP+MFt
aHBvIttszvHCLADOY91h/NUam08qYpI6UOFMbd9nsfb+A3CnFZoq7hrWvJnhjJgcD9MKVgdIKW+8
AYGTn54CFhw4howSWk0Y2tAmnBGlkmYDDrlApkrxEpzDaBpwt4voq5pbx8LxSylol0oh5GzPemNf
s+GmknOQRts68oyJ5hN7CaFDLDkLy0jKqCg9YnWF0Al/L6NW4PSqm+6kD3zKdS1BTffCnVAIoKvj
9aOUDwvSRlKmFjRJMkHxksjz280D4MTsRkjjwokSjG6C8jeZibFXNgv+ag4c61RQEue/wbUjipKn
yfsFyHjDdB/hj1PVgYuyjt7BsnzX4Z51yQcHaUuhmW6ewtZm2SC0IRFs0tUr/aD35YBDaabaqzuT
E+NwFPxG+Rcoyde1HCA0SCBKOoDpRiROMpeLKoASC+2iUJ/ZnsibK2/bm2LcGWn87nzpLqiG1Xkv
Md+hZFHS0WLx7Px8EDX9ZpIJjx6Pzey7U5Xm8sy6oDe4Wiiw14U6mV/cMjsKHUO0x884V6bZIA2H
KVYR675txUxFRHn5o4SfInTBJrIk3xWHngHDxT/xSOaXYuwjTjDk/VDyeGY/07CjI1Dm3TAHdOsk
AJQH8fM0MDFyg8pHXLe1LLN8Puv7kMwMyoyfgbtJ3kElk/fAIq0+UdX82it34ew8hlilwCDON3M6
M/P6yfM5JYK20BpWTrOmiCABfTm0mPZZAlZFl3gDXcz3ONMsFURZRlaSh4RJB2R6vogQgtDpe/mm
hx0fOGEZmKy5MueOZrKLQ+F9SYTFjVPxjxOo4Xcnc/Q1PfwiSPWvbdbY2/MLuOPQW33cVU0+gQzJ
AyV9vIdaVDVpPqeBqCec+xlsYKMuSk170PjLTwocY7O4fjL+I5NCach/sdOaNkxJRByYeAowK+p7
hgf/M7StLz06lpR/tN4FTzaxy54a0+ah/RLufsilJII916b+cqCqLmg30ZLI+VbRMah5CuX5MtK8
ProgL3PJ/02Fh6QLXmueL71o3/goBNkFWYN5gjuhbsKwI+8nKIUzB3MYx4aKFF16eGgfaY3CjZ0A
Kla7IiNk7NKekw9qns9hxA8N5D8atkD9Hzyhi/WXqu4NC7txb0fOLocuKviuyb1RbYGyTiO5qRJO
2YTX8QcOfBK+MtPBcCvqUzBHLgT4pgE+AbfU+Fz9Va8ogzjcIBarviSlCH8Gqg77uTzE+Q8qO33K
2BcgBvGVdHr8664QZ3dj3O/MmDx1JBx9aw8o2AX2/3wlgtMZmc0zP2A/wBjUJxFK+rIsuSb8neTH
h8/8+zosYuMqG4OyEspLnV9/8akJ9j6tbNPcXTzBXKg8O9y7CJ3+sVTEN8kOkaKHUk+Fy491DFAD
xFQMWteqOcziwqUrNGUm6HZn18rckhrvP0llpvjxbqNhQgmx2rbxCTNBZNUURinur7nKbaiOd3dp
N2ccEtkVL/61ybxM/fF3rDwSV5lpwdcrxG2JzHWxCkgyigx23VDQeoAZffmyyzA0lF2+0TIsKypw
zT+NFwb2NAgopS5wWSYTRphkjn4RpuUUhkVWBgccavtyZrsX9X7GU/69VOUZh/UhFFtrnI2jAbN2
NtG6ZiatZ1Hs9mOqXbxlu0h90bB+0idsdAF2Odabm4OVRCAsFpXWmwzL/HrWL2ZZkM2ZV9EipDqt
m/KU+g8En4LjSN5YTMgmFBrPJkV4Qv2M44xqoyFsEkeSrzKJZerBjCtYwzclfbE74+nPtnJWp/b9
2Q+Fm9NLrmPNagkkXCHYiu1jXIvrhaj5XayVGVqSJUGP5Q9YShKpTSxftqdSbtxW1fvnmB6m8MY6
FXVj2ELCb31LOzEyQ345W/fD+Gqol4ppdARP9AXIbRaCpvKkpRMOJUoF4t0s3msVuIz3lQHahDF8
pxhGZVzXtQ35nLQO0DK707Ut4B1UDobIQkpSV71mAq9MMEwKU+CuZrYx9gMfYrbyJBcNFh1PYgkQ
SvBin4ewQnKLRTgEHFvJKiRGQC9XL8Bs7Dhcuhffr1CDERtQ7Y4UlaSVWYNXCbSstQhUSASF5oFV
t8Wscf8guTVIcvRJBFrl+4D/iXeizElXUvDph+DO3PNLXloRWfFE36b+PeQCpx543bcNq1bt5SZF
yf4bp75SqU5eqMUH3RFAcFOefcAzTV5OdmJi6dSVAvOSeNqBRGlKBiVau7KIODKmaT33PT+jJehM
MzsOtv+7rBKsL0L5W09RpNl/q9j33re2EE5UAT31PbnoqLopFlCkk5OOb/ecKIxcZtXd0VEhZmVu
YzS2+uQnvVGMH5Hbc7NWImTeL2ZmnyqFMp2YhNskU2Ed0L5ljvMlPs2+BxIS4VTIO+IKi/Zt8Qp0
/gwFRIl8H+aqwVL3tf8KeMMl4WJZDmlWcycjAGRf1x17WHxx6t2XOesNrSm/yp0K6dxfxo5iRSrm
v1FsYurHtIPjkwHSKmqxOs31YJ5lidmRXqgGAyHfa+z5PdyX19aAZRxrLVqgy1HrSnEixPXKBOLj
5d0MYFk6A3bS3ZoMnIhvI1ua3E14h+ch2yQjV5IKxVZ40+li53lOckAKL2hhlYHGIhfq3jA25G/P
RPzaRMHWBKcFG/vsH/8BUo0wUOowT9aHLzrvwM8d83lYn+iXf4uAOhLHTF/Wwv79DaMN/Lacuw3u
BXtNWwrjSURpz+l+BFV6sKdqJE3FyQ3ZqGvYS9GhoLJq5dR4aHEdW/p3PrqBNokuO4V5xKepclpQ
pPaEthkhwu1S2tmTa7zTFk/jkuRZ1NzoGdAKj8zVzg+dWNboVa3mujtuVU1w/QUGW5aiGtLrVDe9
vEiDdTUQgBTiPzy1iwmc0GBjvbFU4zPW0JL652QivY90rrSq5vJFF7lyRkRCuajwm5V0WC4bVnii
JI9e67FrxKhB1m/gtEPBcUtE/oXC3OMHkvUqVpd6RsbeZ4kBvKcdZ51GyZ6uxQZuHG0DQND+3Bta
fBvkfnyUjPJn5tB/moXioNQXwe0CYNIeDlINZPblpJw82Q/ApjguddYDZWTH7JdAs0H+78pxO9Z9
cH6e+w4qFUIsuiHyrhzojbMBM0bZhNOWCOpqQE19hrePsmNDoRb7/WJ12WM/T6NaB4cWsWxVPSd6
uft7Nl2DAM0Zm2leR5BqmHoeV2vBDONUIx56yo7zOGGuAUikScUHEb9eK8OcU/UFpQmw9sh4CpNQ
Hrixp2jCtvMvGrrdHxAf7oDxXoZHXUUn5Ol6QIyqlc/muqR4Qa8UHOU+AwEtfnHd2P8sKmWOaX/f
7t4JJYGPdV7BAz955pPze9wOoUFAez5mFtVvUeGGNnCfZkBGFSxyD8z7ImbCp64B8iBMwMmhdkXH
4+wgJrOMuNUsl2m0B48DnexAWGd8S4O0pHmGpiC1lH2yxE9PhrMFg1y4Ae2pPB03Q9+8Y+zn2rvv
DNmATFXWY0tP/8rPeyK8AT11j0B6FYM9OnNZfyDNWejJ00iURFfy3wms9GjchRe/D19YN22D1e5S
5o1B5exs413RTgTib9YCrA50yGHGJxDHKk3YTwrkr0RlHOUQv4bQicgOyWIwPVgaUIWFTacfqJe6
2/3FT5c5jSxlWh0ezYsQuFjz9t2yHIQOgIv5QTsaCCPAV/dMnGXwLM12F2Ilr6xP/pA3Kd9vK3e9
R62a8vdWlg4ITA1FzGZXnp6c81f2StDcRBaq++37h385h5lbUQmzGZmMP8wNC4HKCQSHUzXcv2qb
+sqmlKPL8SdYaQcf2AGk4Fd78K7JNGV7nAMnSFXtpMcgIHrxw2DvN5jxzufyc6xzIOTjz5ygn6m3
2J3nDLxUuEvjl4Gs1BmmjZcnAyu8GHPUm/PeUI7KFOq2YgMbx72b4YlbD+RbotAXMBX4rXGP/VcL
60OpydOGUl0w3G08/J2RvuJqm2Wmnb/1P6SBd88EnZA2MrJvNWvBLTN4bQJLsJ23tf8bvx1vVDtr
cQ/xCgvRHqb4xyM2w5nOL+ET85ULk0jO6+jEH5WbEa4vydNR/TfPzyRMf7RNvv31GvKAbeOkddRo
oLA7hQJZpk4kZPvRI86SMrmouPr6I8YMaE3zN0T6ElzBspxsTKozV6AP3PgV/Opi6THLyjm5cjKL
TjY05HZYHObORU/bf9wVoevD18Tc7Rgi23MMKQTTremFP4HwYMCsCLTnipzh+RnY5t1+0IMUpn3Z
8KtqjCEaIlt/mjI42V+VGdLbieCVWOoCDWpo4OF1D/YSCbtZ4gzC533kkT2rl7EANIv7up27zCKr
RZW8+m1chX1ikFIK5SlkRb94Sg67rbz7v3OgOAMf1utcJQA1gBXTZZ45W/HXw0PV8BUpAFCoRN1c
B61B3uvnxjMsEf/B6uc0ycwcAcVXAmvpDVXzsXFb0lzfHX1XJfLAUE+2UyyTuV/oqP3crKPHE2KY
YzR7YPUWvCZGY0osrteoMONnRB6vw5qNzptfZ5G3QHOPahW7BwWqVDFixqydj1b1v6li80nwiHOM
QxlYkqw80bE/5xj14F+uojJPMxEAYZhnfuM38KPU3SnLEM0TtgGTGrgfY1q9BZ781JIPkcjpd78a
t79cmeZ3LyW1WfFvaIibn32LL3wpXxQ1TMUY4Nkfy43lQXVE4CKlymQQD7fjKpABfLDd/0d+SF2f
tvrCG+3lj6Ko4VgmKB89pv5DUY4uMcXaHXetrXE0hiJUXOhgrvUi18R/ncC6XGSXYZdOJO6VCymh
y3u+1zmXm+/g6mdL/+/1BZ6fB9MG27TxqyXaGJH9kWP5tbBFPAlP6E9ri5XMar1igw8YmZVMAFkA
K7fGVEKuyrYDsuE521q6jw19hAvZaKonQAso3NmXgdZKWAlmDEuPxpYg3jXL1+w/2O+CjaV4xfn+
jfttA5zYhxypIKsN53HOqDogxr4qCzdGVW08BfbQRrvfu+HPLWiYvTz1wH7620dsPuqPegBwRXrn
KjoK618usxGazeWz9sW93ibJ3o9ha36HNB/nbDkWYj/2zGw3c0kBghZb8qzWzdsit/UI3JwyGonz
Z5Av0Qipeu6HMpM4MkJFQsBlrHPME5ISxenYUm9r2JjAeK+RhczTIKY47b7yzE3gQzD4AdryyGy2
4R6qJMV31Z1amE+Xhw9ZU1zlMe8yM6D0g5CEwC0Szb8UE0YSV/ecjHdavRJPeSNxUMO0s4lc1nDu
7wuhhMpeiJPzyhH1BdeisfETRqaSTjWY7a5VqL1sF6t1pupLOFWD6vSa7+jOlcq6LqvUmN1NmsOG
F0o6dRq0kr5dTWP6sjHTTquDAgNRTikWLkzSvM1rN51qM5u2MLcxNT/vdJMHoumYuYnOVU+hjwCo
cy9Tf3D0g79Tkv7nLrJjPS38D8p2SCkqYnE1dmq86sKclFjthSn1Kjqsjf4E9m8yG8BCZ0peG9w2
Of7cUdWEXqny0vZzYlDfV/XubzZiErWCP0yn9fxLFPxKqDMILiRyiQC8h9O64i2g6u96KXF+uB5V
klp05GOfg8W/Ihvlay2YbyD5WO+eo6q6zc3FCm4jta6Rry2a59T+YFeREUa2ZPHH1JQegbhlpvuU
RoxtMcuoYJBK70KDHpKhX+Q3yQ3VH5sxTUA9xssjojeTWItPI32PQwjTV+z7CbWUj02aXTo8pIPL
jJMS6OcJ490LXSDMTqrqyVSIrsuRV1ZY/0+AHdIn71J4LowG7nNPt7rq3kuYPlN5oLaanPY6BodQ
kpzRG7kax+NrrHG6zZ3aQ125/2E/14MsAmCTVZ57J9vWp6zrPsnyPalLHn5VNx0qxzPY3uekd05Y
PBkAhEPf6PE3BX6YfBEufJWcx88iYgRqBCklnxgtM/+DHW1D0HmbWKQlYYsSFS5Nm8PZrs7mWFyn
U1JDN751+j2d3pcbY2RVqANInMSULB8qixsO43W++ilvb3/xqEo5xigLAyjRGWykkDcbteS0LhXV
S4Us5hasb9blQqyW5EVM1eg1h3lfTONJ78OSZHUpp4IAjf+sbHZwTzFwjvvgaSm5BLLcZCDOaiqu
OnmwaDOhZztB0yQcK5S+EDRxfXBP/nMr3mV+kQzayNTSFziVXyoNHjD1vE6vp0lznYRXJRJP0TIm
phHalPGGtOEJ4xFKQPLzV9QHo9ZGIBHZu3etw9fE5CDu1YXna0qxLQrkcBZxFAxB8Mh8gi8dsm4D
0BpcB/YSpzbqMEGaQZU4T4UI76Fu42CXig8IUK0pwZzaAZGOxWkv9z1TMVDyWDCpQ94oCBTpTgA4
vIjnvjK45kUKbEgWhruGl6mBab+kiIbIrMfIc1uR3ojaTmXdeR9bIFenlO/lhJj+ctHt/HhbOG1l
/HGfcVyy03D2DefoJIyuIQxgOhuWyDHelBx1L24Lcg/5/ZxYj+gQOO6kMeUNCcE+DicDOn4assta
uaw5NBKm5r8mqjQZkSCOnQ08Kf6+H8RQXVbUabKlj0jdqVA79GhYXlIlutMVodc/4Jiu1YUxhdc/
fLvCQUX2t2ywcD9FFdYJFfUtbjhjRMsjv4BcIPGJifVkEjAC0rsasMvzndHBYKOdyKxjk6WjPU62
aXmpJaLYSyiU/Pu/XqPYxJVCBbXKduB/qQnoX3wvM3muqTMhaQhXfnePWLpGTujuCyCzDDJ4ZRzR
m/6JogLlJaH6o1k1CUpBwqTkbRSI37meb8kOmHuZM6WC8bdB/SALO2XLIk2s4yTlUhVLYHyf710f
xvtWAcLjMpZI8jZv8viSnZc7jhqz12BCXCvBM74Dr+IcDSV0V4FqGHSMW7He0WyrHW8c1FAsxAkO
MU9X0jLmbZHpZzpNe9GFVP4YpNQn+GwarTpCzrQBCWbQn9L8xei6N9fvQq1qCuR+eQ9PrExqcZTy
rJN4Dk+EpgLxh/EP7+ti6HRo2e/3hIbsbEV72GrCwiY2TBCe4hoHcglK4vVrDt//YlDakKi14JjK
QwpwoWTE/vh2jvB6oTqlJaitgvUPQOVCv8UZvl3ciCp2H+TZmy6iFffircYg9J8rgjS9rV65rVwb
mJGqN/x4yy5e+V8y0MBvNcqRqtj9VtcbnlglxBQ5k9Bq5HhNytCNlxd4leXtlEuFpjsYhT+0MFwl
w4QFyFPigagCAiaaeiHmRYwM2gs5GIKEHVcSA5ClgY+gGpy6KLYr336ogn2jpSjaBiYKzHJOARNK
c7542XtHT+i9AZ+EvBlC02/jSow7etTvUM7trw17V1W3ft47G0le2qdPGOR47Detih1h2iGNmq50
g4qA/W7yFDunxzDOnJSJooH/MjxDKkbwx1udN5XveS79rMu8ECQX//xGezDawgMCOShppLbIjxB3
MdADGEAMMx0Iao7V5AjvAs2tIYUrcIbyHZ4T+PDnp6hA5odPzs1lS3uyo/vYvnWEVcpqiz2w/rKm
VFo/kYPIlkemHnTYq16Di47bs/FgDR9gOngL8Vk+KamxQFgPhC7qjQQ963hX77yg6X7BvdB0zolf
6v3GyjIbQwG3FAdx8fiyZp1xRBaL2DmPRaRnYCYNVyZfN13tR8LLaxPo+7zU3AU6SKJ7qW6gJI/F
jk7QdN2bMAAJCb2qdJCxdJA1Ob2Z+t40WV7j7NPM3ZSUYN7FlXHFUObM5AyggyZuYr/Z026vZrqq
U6URGBomKz76QaNvhB7bOYQjTvqX/DWhVFL10CdtOzxfMU9OqlOuWYkQzCNTyavZArVEzxjgPQ/9
O0n0WCf/iPhykn5+5G3hnoG93liXy0mN+Ng5q3HryamX6r2YlPq0GTpPTjYwZPvRnGWAPjDxau+O
m1K4Z+Vvd+Vbv/EuH4bUsZis8i3jsgFdSXOXKj6xwV0/zZVg4lqUPQhGhjLBLJrvQysHb7rvPCQV
CsnQMqU1i2XZI1bc6CVeBoZGVV1dU0+5kbqHPUz2xpPyVQvjQ3mRd2zYVEQihLviyDK46H1Fxqij
Zucz4ZBS5ZVoyUNn1J5rl4QiwnnNoY9QqobBi175rHi/MlS6exkEzuL8lL75jG8wIQingLrs9CjD
sXJgWotph0qYQUnXJaYTJAEpFjxgf1tCZokrjdWPw07r1IK/8Is1XGOk4dPoEGl4j6/5tD19nM0S
ZoacDdOzcQCbkmrmj2J9zV6txyjCuO/uooHcc+Us3HjMmTRUuctncJmb2ZBRsR/QL57hlt+6vHYg
EwMfgD0FaHlM5utjCXRY1/veULAc9XNQUfmnatxD0I2+tQIXamV3GpHM/67jOEE0/DCPML8bd70w
uR3mDfOia5GC+49XFVcEdN88Pf4CKovyr3bt6JDbbIyXQnzu+4ysOq/NnwnAPh3Fzoinmru5dnA/
EwbBBs1s2Iq9+dTPczXDX3y2L+RSOBo3Q6WwrJ9mj349KVmbaIgx1F28uAONNXFN672Fl5m3uSrv
W7ObumttegER7ID0wC7OZZCqPtSSvBhm8nvRTXar/gBELijSwWwSNN8jodl1lzsM+qwp2DNNfmZF
11pKbdkJGXgG1ETKLEhCiTtz3pNV4+idij7lL3hpKqtxd+BGPhCyv/bXCtUtGMrf+Gs4F0aZ1HRB
QpV9gIiqCh274hAKKsxN7hC9bhq/anNtcPQraWH11Frx79CnFz0RF0I1rog1YFtrRlIsBC+0Kxsm
MYMA67g5hBzLLgK10gZjkv8q0T6ZDZAu/2XlE3Bu7G6BPoc7NxlezxmNxC/I3f/mtpInw0XlNCK7
zemX2fe0UDE6j09B4EEGT3ADmNYjiOHbAfh++7E3b6M5rjxZYXSXlzAF2jjEOPDuLk85ECciZJIO
yvjbHX7R5En5Epov6XEnWqrrNo2yubhiPb4ySW+txWm06EtY7V+VIT4pqCx7rcUZpMxB7dOaqeZl
jOdKZAeReUOIq9Gl2A+guFIiBFQQ5qc9Uql9q5PLs0FrUjWf1fnofEabnRG2IprLQDKLb1GEn1bs
k0Dg06PMoCweLVm1tOcXmziNo9UQjD7/KLG1tNvu/iHolDLFs7KmSH4iUQQxIp7C7egREVynT5dj
HnP4HH6aR7V2b8qS6XXlXp5gChRf4QvJIa+kumzkP5+l6semzchPK/kKpfdbX4nhwP16zALXS5nA
klVRYioTxDHGWN1z8+io0ovegiDbdDHCZgB0Gl7oQSnTRIGAohNdhm2xtimh9jnV27RF/lbbtam2
xjehIiBlK7muFrfdhCOCqlQWQqWFVrKV2Dzv6KvB3hxSrSxcNtGUebLMU6bPkl6iFqgn5CmDevxX
ScRMXjB6BKyo89s2K77Qr3eIhpvnqXvyrc08G4UP8nx+gGlHXlzbUI7n9rn+At6/UgQkmvZW7QjQ
r/ST8iTH+SvmRgHcKHjpLakxX96gcdX+Rgtgk1NoVjqkho8TPjsh5vvbpMuzuBHl/VKNwz/EAfgx
8bvsVdJ+Cv+h7cphKCn4l2+nU6vOmHfb+fSygsGQ7XXy2cy9SPYDbgrSsmLg3AUWQzzRdSUX/Qn2
VwUFn2vTpSOTbvpVLc+5sRJ6ViXFxGe9FeeorqzEjUxoOkf02vO6RmX54jd4AoeattDkdBfaL5az
PRjLga1RBnft54EBQO5KK55SzOwDgZ6F/SUVEEA00EVY7OLe7xYJN6R6R0mioUJPbGY1C2GdMFxO
csG9g5l8n9Q1ITFKnSUDI6PGppZJF3im8jQ2s8Z0CjM+GCJWlpsHL2pX4OjXhlNws71waA+WYwbo
/gHvzROk0u6GoGRW3TwRTxijF+jH4Kh1ooRlrOMX31V+o0UFDCWhuKbzTSeGpnF4G4z0W3+RuSMJ
D50IsFFKY7wByJBWpnfuf40GCdOnF1X/vEo/kGWYG89tCyWIknWCtcvkb03cyK+FAPU3ucIWd1ef
oWo5l6TRXJGifdsbGrK0/HsaJxp0VXVX/EE9/SHIr5T1VM4AUSokw3njYu6o5B19UZ6V9RJorIkF
aio2YjtXtP/38xh6paNQhIWucKDpRTKFt/k46LgnLU+ZHm8nSheJthhBpyUh5h8tmeN2Yi3qhuPZ
IJYtDRHQ5ryoEQnp0y7ux3CRLPELhIF0XqH8nJ2SA25Xrg0Njm8vaaWnwCOihzqQak23AOJUZvfL
i9gDD06q3h2xIfwE2M8eGtpeDUZZaIVYViGk9CvSfaTt1vWRUn0eLrCvBdXi+6xnKmIIqR79Ht3b
q9sJch8S+UvfDMS39nucJCorrNs5k+KiN5sBFMIANXDS0P5bf1KztfXl8d90lNvf+qsjqp2RoJNs
EIA6AeeTHrMlXPe3pkKOorKl0Kj7V5Hwqqr4G92zI27+md/rHDd+1kN8/DEjz4Soz/XAhwMicTpF
oqaL+eW/oJkvYmi3x4KU2lGQ+Dz8RQ2ulf9AZSrJk82TRyfvthg0Xq/l7lhLcTYC8+6N4niMBDF8
r9bykXWG+COFfyH46FF0pGCc0H8vCSZjYW4gqsMxop/WTF46KtXCfwqRJsUdkLN1le5UlxUleIqn
xX8pZmguOat51H2evBTeTKcbj/Dy4InM41LFPYemnHzA+QkgBcjnL4NRU3Xc9a1PiKE+sqh89voC
W/9U1RryQ40fvi4iogqPBiW/wZGyisu0f81U+4JKQwwzxdw0v9sCubSOU7NlAJGfEXIFolWGBp/c
z2LsbSB6G3WwmC+SLra7Z3znXEPkJxgEIY8MKSzYbXB9hYeW8KVpBqqi277Oq/e2RC9eN1Ws7pJr
89wDEk+5OpdAn/6QF0m+cD0byIRKszY5LrvaPRw34SJX8fzus7K9ouoluZPITD5KPoSjPAnrQ9LA
nAh0g+Ik8EmkAPJgtdSunXVL/XjjrxfsCiUQdsfRUjYbBxz1tqKGZGkmzqb8Nr8UgHSchwdZvCnx
sNfmLPGlZkXBbwojScx06+KcADwPw95BSzFac69F68fyZOZSWlJjrqEzetIYH9JSFsTUM2cgWj0x
Sjj9aPhHXhg+HNw4SEnBxbeKFmvgn3xVlAGF2VYqEExcRnxIF122YLs3ijFuI5ljdEJTQTknibSw
AJS5pU7j4EbQmJiwvC5gu4ATkKwiom65ak1nB1xApLir6tGcwF860PwqpUQF19MLZYCGovfOIdxX
eGYiVX+hJn6I3+kgFoqpJrbPp0QyL0BEvdSIf7iVQ/EZGSdJAZKdH5rMcfiSvQ1D4P+NDNgH/TOr
SnVWsEZdkPjSGdM8x1xDRi8CiOTm/EKXf/Jm39PI77gtkQ6c5klco0eVphQCNgu7WpZluXfu2WHx
+psuIOY+0DqHlSEdLXUOEWROyFFVCv/ogkuKFjP2JhdYtIbS9lkamF58qoAEq3mKrjrxp0aYsHuu
moOl6nCNl6Rb1IdoJGjmJz1TFzW2M8vq7BLyOSpSrS/femlena2oRFSGvVfSE2JHHao/8GsaJ8dS
XvFckuwu62PZNB78M4hVsjQ6dsZHAgDZMGQC/kSUahtMEgRGI45X17XeHUkklGo7lptnAXsffSRi
lF1XGn2nOrW995ykId2hP6zobOPqJS5Rn6cq9OCUQUK5xcUxZEA/6bYSzUeCLaxHxOsVZ7i0QvkM
8yof1burUJ1iiYnlpnRkevMKUnE6VTxyHWuf/E2RTUxDh8yhpLTsos80xgJgsr0/wt6pNg/G26mm
jxzUabgxx5bQAIAXvQmR8IFBRrQtMimt2BfmDm9JcokSycxSzYJMJ8ytWDCjgRO4SYACz61145mW
8PYq37wAzKJq02+mepV2UxHlgFT9KyAK9wLqvz5fJ4+Sy8lQHLNpXik4oVG4NT8Sh0lzbQs9VqDz
C4YmbYJ907EnK088ksKSGXDHWEPb/e1oqc+WCfZl2DLQCXwLvZiOtm0G3mtP3nzitw5B+Pd6+3ZP
3s8ZXKyZLaxiy0Jh+jT+fphvo/fou84MqKNMcfWCvuFEutuI/ugTqfEU+RU585gZlql2F6lw4QUg
HGpAvRbxayCnWR5CY6xKYLGFj8l9KYFGO2ulScIKiSv7Bq7fzTgdq4wvjb07BOBLWSN9Gx7MGCqy
ssJ6poG+uuc7xXZJFZBhVDtD/lo9nwO3+oMOj2+1QqTvbMBg4mgHNzRCDjK1IRAvIdEm1GErcgZT
PZUBQnllpvguORvf1aKCJ7/Hhz5Pbl66qw0ZNbqddnymppKQxBRcIo3QueUsqAsZ+1DYajPX7r+j
pgSnw8nNUbYzep7A77XSuVls1ccigimlx+j5A9IM6v6EMho/JmlzQJ4tcPEsGsIcy/XWsRhQYo42
F7Jcn3psCcY1XZicYI6oz+TmwKaUM1NlQABWShNWyOzOvgo02O1/l32JaZgfd9ZF7atjYlUpqYM5
cq5tKdXlusnTHEqa6/2r5bM1q/afE1slxmCJdffo2dTSA0XnyeKvH1rLRTN3DL2xcwcbEvKYD+yK
9rQphS2fE123B+u0CBfAZe4X+I/t749Bok9x1KFEySrifPoyLSS4gKIBajIA0KcaGgczgQJU68XV
p/Kv5NnIUVA1/x5b6H1xa58jUsjdXdNAT0Zwf7WW36id6TpJOW0TFqffLliGe7SKjpaBpJJjekwX
XUCpqNumMv7jcBdUn9xeTVO/KffklFOGG/48C3VLjJvJfHgFKyGRKmu5vbroQaxQhDtmZUlOM84q
D2xdl5/p7yXXlPXjgadkVqevz9Pzf0Z/LRYbQpd93di1LZInu9fX32pv7jvJb+OzdH3yE0sdq6qv
xYC2p7cnOvIPzzfwYpEw7n6mdwc9x/tcB/46hSSZiYE7reH5/uqRZ8L0RKJcgT5a39kyh/s2DJnj
9C0TUgqh8heAhwSGW+mt72RNlE8Nf3Np01oYbavRLhqHlb8ygVPJR/h262m/MuWfDH8Re8K7vpmp
wnMbLhUmCJ9+sCni7ZOwplTqrAaUqduGnn05plbYnIvTSUYLp/AOZSStwb2nIWPnKJH9z36UtELM
TxiqukSxjMe3whVK0p+mCSN8UlY+76vLQc6Hu/1Wk5EHeHtqEKPdIxZomoJ5WAJy1N7n6d4eWzpn
9X8PJARVBSkxsH2mcWz+OQJEfx06Wmpou1uLZdHwzm+IlT8oSXCPeEsY4/jDcivPWkfsCj5WineG
pBTm7yCF0HoMvXWMPmwkdJKpb6v5/zUYBvknJXQfz/uiaSmDzqeC4O3XHxORBjSk8dDi73vl58Xa
OVNHMktUHLZcnIrer0aVfoJm/a4PLT0Sa+i+zzbDHpeUUYyFAOqLGZB+2n8GOJFJQez1SerxY4hc
1cLI0C3/SQVu9KZrJOFstG33tEHVxvfMxKzwqKNKJBMb9yaurhwlTygYfXqBSVn4t574FkhPw8z2
st5XRwbWsfbj5ikP1cwTCQW2kFzAY+JkDVzbHLWNGXIrPIm2Q+f+BkS3/bYlKqUXEvavqzT9e/UF
S5Jnu5vjkf72/6AF9o7ywJ5jqLPLTUvwtCex/pFEGG4s0ZWRuDyUIXhmJK0D5Fv86yqdzMxBaJaw
Erum88OOS3yUtbKeAtMGPNWNUzodxy+NyV1o2kmC9/L4iW9W9smdWgGn5iRb+AtqBSDLGcw0YtEX
pJ3pzXxv1OHKVi7AzB2JOKF+jxKPYVHTcILAL48AlDRUElQvq1Pg9IkxqrYMYd9Gu7+Kwin+IaOG
jYNCd4KH3kLIFFQxSnjj5whlL1Iku5GaHZ1Sx62YjK2RZSCX5kMOffOa/xqk+uzfuAIvNEXpQE1I
A8nsWorogokoeGWeAVvMLef/Wr1GItddigusCUGX7brp5eYbR3tfVZL1RQrcurpVydkISk0qT899
N25ntOhBypT6a2T1e3OHPWZqwWK2Z0Er9t+z+ARKBt/5EzxcMBQTPN+OTwNr4/HSJ90c0iUlTxFc
rbIHsBfvPWhbV4Sqy2WNtbNe9ourMqzdzGxF78gbOIffrLYP+NLolCIzqGWW847s/NAhDq3og94i
T5pFDyYRz43inwBgLA7n7JFWExcK/BmfVIEzkDj7LlMtc7d/EMR5Apv5tx5tm+gS5zHSi8SM1TJv
3YLZYlcnwwxjBlkl5lzPpgk2XnSd5YyS6e6Vm1ZL+PI3ofe44XLZU/6GJMvhUM30uohT0m2kokIv
3iBtGHUl3E5IPEwgScibnNBT6YLS78tDLxieEXEUMmB0vG+yFNt52tzZtgF4wKepA9pWOgINQovL
WiELpOoc8fDaafXzSOh/2L/BPPiEiHRWeHNTCGunY80pSYP2ix/chGZWASEdDdSSG0atVMmqqoQE
jNTN3sDPv0wgHXcedGnX19X4hbT4WD4Z+EDt+NRGNtvw0NR0v7hzdSQinKuUkv6Sb65iRAdIWKXJ
+Dh4pTUuuHUMfozMsowfJwdCkymTXRkpM63cugzv75VyMrt1xEIL7cNqu6AhZR0LgyHd9VitlbEK
fcOWMoE24yHH3lnTmx5891bDy28MiqFymIYzP01R8GdKBD2pLTQZAC6LFI+x3PF6kEt+9g7ih994
DVm0jgtDRS0UJ6LPLk9vKjkCGZCGtNID58eJdgpb4I60Uj+3b5+enkLyB+4T7CtdJJMlYabp/0+7
oAEhHrcL7hee66/K45RD4IUnbx1VdNwvLS9/6xwJEGC1cxwmqGrqaK1SdlmD+T5zWFNXRt/gKn21
F3jp0Xs4lea0Z5WS1Xo9vIdsm5ZqRx+jHcHgSJbKQ9D2nvjKP+Ju6V4NJKskbKPkUbWZ+YXMCV7M
QM2P6nVUbqiFaOALKyMQ8gIUyo/Jh+gxhKVwXjw4cRbTRX/IJJbb9gBze2XVibjGg17zc5iwkPmp
jvgxw21Xloab2cGI4omAa/OGnVmk7xfX5L6z8ZbjV043+rxKlBfIhLs2Q/G7gRq27Zom/v0sSmTv
MSg8VcfjT+1WDnnwTDHTFJe6/D8nHavbwcA3FH+e17qHWtXbWrU4X3mzQIm+SzZAajgsnvLb4MD0
d/On/gZ//H2cByN7csj4PdTMQP3bubxa5nk3u7StQFydiT58r+5nnqGE4zA8min1J211UOldnjXb
yHSxNLgJ8xl8TVoF/PTaIrBoZAUaLlapNCJp+HJGxJacTGUVPl0TY+OEWrLnhoTkEEtffouWgexZ
FS8j/ifOnxPds2q8upJuuwK8PttYvbSdJyEn2VQ0S6dZ50pPKqndeIAwhcZXvib4HV26486OuVfa
uLMLbD0cqaH4wb6m54z6oAJ+Nz/6wE+ozfeigX2YkL8VUAZnJRA3pHt6hfkks6D1Qi7vaecTjVmC
bmI/s1DmtBTchYQBUUUXIMW5jJ8qHFRPSAsTGaW4HDGBSY2La1IlMSUOkeC5EbqZtrycbW6uWU5D
7hXnN1LefmwcuySjsGUfPkMHM4eSjUFpwkc7hx0SI/137UZ/PYjsaARChaFfCn0VdYU+CFhsu6JJ
Pps1s5eVblGCZoLke2E0o8mfvnRjxZMY3C8m6DqDejUxGCmkjYhR5xyNDE0rpNuP4DRXLX9UB5CS
QLIzPadbnDU6FyYXQ+3bV0ap43U94QMFQvw7OgeVCPmw1Wc9f30L7uWoMnZ1J36138UlUhSk1CwN
prnnp48pios11HuFeSmflRKE88lVeulvuG5w2Ctj281mIJ3rHw+IXmb79Qe8+tGp9kfhhSCb8yP5
cs+EoomNMZoZNKIXQYKByox/68XpxlKOOmye5cwlo281n+8J6rJcYMZ33vHZ71UES4HdmJO6E9ex
UrQlvVrNYEwCFV1XdVVwPBV+eflU5O/VUPPxGkIthAWR9DdhXWNoWkIRXqCU0ahHEnn7iivhnAkT
ox9zpjEqoCCQycZfOmXXCve5ed2MMqZOoS8sFZPRaih2ce6H/ZFNFHnUpnxwgpyRiwpgOf3pJSwM
iLFFv7OS9z80/vu4K6I1qs+Ithbo26TZoh+MkFTD+cygp9fk4mCGVRBXhlVlrt63mZGMaf0bjfgU
nBU70NuGwEOxKCe5vhKjBZwvYf6uJelyKQB4WRdZ0OgVoTvEJ45NouBrg/dYLPmUHyHkkX8Bdbw0
gskSTTpYvcYX6tpJqPuRpBltiOCt0ftw1NID5AW0pNvsged8cMs5R7feZYPaFgdnP073GcTL9+vx
P3d/mcU7R0oLdXA1EyFG3kK16k3jy64cqZdrhWKldIDR9jXgHug/bfPQLWjdQFjbP0BHIaRNV34G
XR/K5jOUepUxkxyXiVtkAGKZCc2C7HfQyteGM7Vl14fspv+w9/zj0glOPO1T68DsmAgTv7KdlGCe
2RFY6MtsHwIZqNTWphEjGIDzBcRp30f58oW78OU9Z/3VzV0G3q9Hjl8t2evH0rIOoQjzQpIQwkAC
hUrUQVnDAGusXQmy4uJNF3laQJrb3rSwhw3TRzfycTfjRqIghfJiLjXB2uKNTR6R0TKcDgWVSugo
DYJA4tbOLGiqW4F4/xa9pql+s3I3x4Is7wKqHDt4BeJVLclXyanM9TNY3Rgy2/+10bw2Xtw7qtT1
jjK/p6vjS0H4E0L89PMzsA6MZlAui5SY0CCM08WxpXnluXZ77FUahLoc9jPsSe7v1YMKnpZlVSFj
fwUS6DTv7GrSjWXqhUmZVs6s2CvmE34d6DbIJYevNA2hkj6Od7HgQozlVG2TqALWY/N8KfX/6Yr7
iB5BX2H/aStqXyXqw4LA8AXG1ZzgEB63P4a2kA2EaM2Ync2SLhHHV1XtsHx8e+7cV1mFAwasEGOT
/560Jc/gZAOGRdM3Pf/iVaUgV/zjH/AVhJ01YaMtiV8cfpmTT2tJGuIdMKc2AEM1PNPuO5LcI6tR
5NffZDM6TQpbsHh4Y2k6uUhvWaA1s/KBQNJQFLvmxb8gO945YBwQEL0QvWl7QlSsU4EN05qMEYBE
peUJabhZHSbCGSzMyzfpNua36vi/vFzgLZbcoj4/laMpYMymD7/V5UZ2y2/xy8DbfsWF4MKTpvOF
q6Jbgam/KRDo3VT6y2kLEaXfvXwdfwUlz3+TLMRc/VDQew3J1LNLlzenIcYtPQTtRGoueiskc6E7
C7tCfMyERF+/CYZintjJEe/8/0roeF211kdJ8Nj9kGsWwY5Yr9e9hT4JQQUQqY4vQGH3EmC0o0EF
JivVDo7AXd6p5bKkErI8NHcEktqb792yIw8liLtQ2mtJl8/eNbdsuNKS5hxEs9y/9MvgLELpu+Hd
3Zk6TAE2xN65Lw1LuccQgsaS++q346kGN1YHQMLMJ8fmY/hIg8CO7xvzSMNlcskOeU9YBO4lTR7R
h6oHyojQcK/Lb8c7ujvRzjh6Yg+nlZ99wBO7TMzMJd2vZ1uhFVHjLEciKSVdwuH4RiC3/zN7JTt0
RKYlnNKaQqVMBkIBPDlY3iQWk+TZ9AO4OpzfX3UqREqrLDZI+lZLRM6dYED1zlUZDTOGKKg5tZ3K
RE2qn1oEwAY1QPFDhPoTeM7Xsf5JPTi0ciLqE9quzS45egEWrQRhkchZhqvQOBmgiaIBRPzXMcth
K1qFzgPRpAWYrHWFeUDhy+xUuYlDC4m/QJ2EIzuCcScz54XDR8IDgHMNFZHglm/oRMlPGyWLG1ml
DYIliNq7T+blxGo8am8nplueqP9XWi/NXlNG6ax9qVa6lGtTr3YEnRpz72RdWQTM20N8tKGNgMHW
C76X39wm+40d7cLA5zph33UBW/KhFND2jdYrpZO8JzrIrdLW+giQcp9DhlgysHsoIatmtvMJAftB
lRhc+yBWCVnqUtCGyOdNSKj7zeOkDbXmpzxr4oW+h72yfx3UODi3pdaxbW+6ISxb6mIFxAcAgwTz
le6MaQjglRloprmJzdVl7qKeSdN/OmvqQ94CiBtgRUsyYPKgV+/ZCSsuZB1Ka32kC0ZxIiXgV7DR
WEIWfJqPQYRO1GjTCIV24dFWcgMVsDqAkEkSVKtNfgcFmuGfVPmT3v9Fg6mPlFSEHF82h9bmNx2I
T/bGw8YQGnvdYzrEVgXoY2/LEbGwkknMd/6Esy5/adHKjW3ILydvZ6COz94yrZ+j19CsSoVqcQ48
U5Qn/EWrU2VRqRcUYsAGg3GGBc3WXV12NMzRyGIEh9vje61c62Pw173CQUNNJecrhVvxnNbgcYWL
ozWb5WnyEoE7MhrKJD5BzfIJ3gJlKdSgVBG7FCkL7RXGav4DWYgOdsAZkSalk3s7Z0eO65HfQ3cL
Xhvf9piFuD8yZ3k4Q+TJvphm4EzvRbxfbcpeRCi7F+iEz282vLVSmz/5k/HQoCt6V6A4KJ00Y5yh
TvU1xX+IEgl8mOn/RHu/oMPkBH3x3M6pBNXUDb4rxwYA/fbcm+txD8Q/Lrh/A7VWL7Bj1WHTZj8k
jb0GFI00Ukn7HvYoLQFmXp26T/5PDAgdB8lWzIUnV7aT5z1yz4OHGE2mQ9R+OG4abVQ7iNgGzUuG
AJ4Gi9YqiPq1lrnOcH4gOivBZSk15fB1UnIPebJTxzIkN51z9+HctfvBWvqNMzsP3Oc70jZboQhv
kPTzqeQCBXbsXpZjvptCSJKKLS7afYu4cLJanhjaEpsHNI6Ji5O2CdQYZF9g69DHrfzOOhr/8i3b
eEjl/GVvggGZDGa3/t/kHv/tKHSYk44Wq2FQnIr923PGc4PaSLubDqohi/u7G7aot+EtCGp8bC5p
gJI+OKGOTTj1ICsn/mIxV4MSfLUV2zYBHzdEpZIWMlzVHM7u8/4mDvwwR3EWxBDApTRVim6haPPO
z4ek4/W22J8oDqyy4ad36IL12frHj7VhFXBaWBe8HtswsbygJcz3pqGEXV2kLQxbrudMsW9/S1Mh
wyQFMgcRU6OyRoOHc4WowUv3m0aADUi/0wrOJw8G5gwt3XgT0Ym9eFENIxSIxFNQgC78pi+uRSka
3xJougivVn1Isu8WaaA79KTg9IxKfUMstgqXLtIlArm4DvChLrHifotNgMd2oS/ozT3DE0ymcCeV
vgrDxsjs6VTgMw0TyvZoo9RmtHoUFierOVxO45AYIrixN1WY+02Y/gZTqvEWwyGs4AKKQ4PemEpA
dRbpc+ddsVwfD0j7JC9zS1NXF9TCdaLZtOdj3+z9yeMh+Z9seRLfVNRfDjCN3hxnJKgBBGzoBlDv
jYAsSYjPl+whOrcJtfhc8CNMKg0MahpU5LGW+lmWPluux7+RbHhhs32yXrtwrbtlfM8mSY5T3KmL
GD08T1uTvQU/VkBhUWhnhv2jOiAsqk15x/Kp6T8tpm/g+ukWu0v3a1QJCxsadEIAl6m+Va36V1lq
FhBRvwzwG8ijf8YkidgqKl1bZ8dMB9LSOtDId73x2jnTVWh0cJnBdybXljO+M3LpJ8Bdcjw6sbGG
hlblwo/Rfw+5AoaenCy2vmOmvie8fVAswU8ckhRME1UTgp8zJI7OXBwxsvTdiQnInHccgolCBjrH
EjWTiNsOkPrxletE/CVbaA5KjfYISyiyEPs5TbiyLB4Rlb5o5gi/A4D/+mNcfFDMpnm6YelMmxTd
bOVibCrD98is6i7j1pqB/KJANTY8HdzRcrmyihGLkRT3RJR4hK3uKWBxU8cLNl1+MZxGFMgiWN5I
VwnvPK2W9KqrSOqL3fLU2N5OkzQrb5XTWXs2UFYthy300IHYY/RjH4uHjCwhWGqdRFh6ZUywl5pB
QmIT8jfFfKW9knDRdxLGafAdKybiCh6cdW9+WkHMUb+Xuk3leEwP0VyYvUT0wTH7B1MyF6X2QKBJ
y8UpjgqJtzK3E3eDEQ7kzVMHmgKyn2nj++DYs3sIdjl9N2ZB75SKHfZeKsamI9dnlsv4lvodvBqe
gV2qPWy0L8k2pAkrjlxG6+O0UC5jEDauUNATF5oDaObdg/zdXFRqMJBeFnPlW0Q+wjsPJfKyAdzv
QwMqve1zBZD+JGkySahGkWBDkvNZ1UqG4zblxuyUpV1SC5CEnigF+VH4ZmmceUJjEYVxgNmYywq9
C3J5XJ3zIocSUri6e5OuDsLpK/iROFBjc7nCmN1PPLKruXktZuVH8BRv2tYnvEgCwTmFqR7ZyWJZ
1soyUUJYchigZOnVSBsxtxXUkwMBctbCZSceFY+LRLN/mvEuTpKco/HyhxriiFDU7fPtF4AH4VSw
5xpVQuLEI93p9yeGMym9pA7Yx8N4MlhK4vBpuPowSHSKsN7eApeXzr5Cgj4fP3yStV7VdmbYF2OI
T7RP6XW2J8TFheQAbW/Rvxb9L5iCKFN5ZxDFEkc96GE2VVMtCrAXImEgE5p2zjud3hayEwhaFhub
Ed1La1Uuq9RRxx2q/RwqnlAtzhN8ClC4hz/Y9tvvcPeJRJYJwS5Q0M20UmiIt9DhInhjTifXgQZq
nZbUP6/ljcr0bSMyRVP/3dnRlFz3T14D9CMf68R1puCBPpejdonzB9kdDybM5Tu4fVCZ5/TQbRbT
UIgcgDKxXq8lb0zRFgwzF+1XQBSPHdH5CH+ozhs8MF2h3+wZMC7zl5p+lu86vWSUREaGVNphwgSU
5QFKG8r4wVy/EE3W/VI/orcjNrnz/ep/Z69S5hYfEQYKd8rGmCvEX9COac8kgJT6YiLItr3lxOoN
OGyDpq4WhPBxI8weGLGev6V9EPkkGxHJLkpmC2mA+7Llz0BakoVgFv3ny8D2w/aI8ADuMsF6F2gb
UvvVbru9tP3OnONG5unGO/QKmbhXb9nYgpS7CWDBzH+yxzGY+wkA7wGyPJhOCeAyxit4LWjwaF5O
NnfVHo1UliXkkzLKX5su7bDRt+4S50v9Kg2k+utmA1dfxEoCFm3/6Fe+PnWv+sWkM3ygHzTcQGZQ
6ibbXgi/bsAA+OeGec9Ev/rFgFEqy9OsDM68AQ+PvnJm8XE4giOEAOFejx8wVZxoX55utX/h21b6
32yhgGbrj8b18AnfECcDnlJOqrcZO3J+Bn2QX5+Y+a0sRrmkCnOge4xwgvU+tO3Y3SrDJGrsSQCI
ihXycpjpzNLG6zbPOoq7MzwpB7v4LhTomI+0mjNIN+csr5KUUL1+Wap2rFcRk3Qh9DJpx75al/DT
/TWiQgsRQZeGCKa+DTBerH3vtGjSOhkxzLGUIJ5gbC1fnx9Oy1QLnQuDczEmm1B61ZP6MxcLba5s
4sBIdRjS5er/mZro9fcrtqZOC7r6rc99YPgOVBDw4OReJ2vRG8lqRYQMDThaOIBaeISGA6iw3Pkv
u9JoBQPDyQmCjdNj6FRZJ0ysZ4OBVwpjGuIv1IBGsL1ad+N9UAAVXuF5sqKK3Sqt1lSUkiGpCITV
XvXEJlEqa0LPw69ETiX1iDv6u7aLTuKDLUDmsy0VMI1vKWDrChTM7a0GEjMAu6UeqMP1STOREyXx
4t5q2w9aGTOGAUSiNWCgmkL7jyUMY2b/v/lhf8Sk0j3cq8rt1PF4wQ2G051aTFwF06UyvBKYLOJe
jIbDLcO2SIEcPPqeq3GfqAdGPx9iBSByfuIGt9uRrPMX1M1EXmURYYVuskkQZuXTad1S7tiFUCJz
Do4JQDHUM7o9mgImpysTc8LIMYZuvrMbvRPeDElufgJ0tOZyGjjHqD6Mobt2QvzFykcEgSDj+MNw
3+5+omGIKxYYv7loXwUhvgxYawDGq9kWqz0Lr9MKexU4EL4XKSYyrOZsYnY4MlbobH2j/Gyse+rx
6SqOk5APFZ5DICxS4LLU7mhD7WMkDBeXid8SAFIIwInPmF7iQn5t0xUw7+o6gLGAD4comfKCSi+G
KjRajmMjc0Hg8fyaoKft08K7NEI5nMK08gX9swx7rgUSde7jQdq/ZwM0u1TPuxDFV0+wZ6neSAm0
HJaZDIeaK4hXHQ0YfKD7j8h45lH1qDFIqT+XW3HxtLvskocSp99e7kufLtIegrjI/mGpJuNTKS6J
9ltLa4QtlduEBPMrGkWkD1Pbv4mk6yAcLmT0IxsSnvfuq3r4kWtkhvMeDAw68sQSn8liSbDrSJ6A
udIfZ4pxDOiM8wu3K8Yee1NrE4UB0a9e8CreDCVmc65NmsDrB0hcwoQfgQ+nb09shb5XO/QV8I2R
StE+17zAzWv64sM/4DolyI2bT1v3R7r6a9WEsOpf6TNcr/KaeqVIJdV43Ycr5f+FI8C9UFIYVcwC
GYqmHELifXO11JvuEqMgBQ1S6Zy6sBetubLKaUAxHMofsgesY/WgXlYm6XNLwvilQ2aIKCAUmfXO
r0dsPSJWIq2tXZCI0JmFyVkny79x9Med/DGCoI8MPJiGtuehbbkp0cNdmjMPgC5AaXDuF7aQW9US
86HNPCskh1OfmLpfRxaqJQTYTSAwLmDfmCX2Mbc0eY8GFf+FhYTAzPnd/XBfvSLi/vsIfYoyyF+4
v7cYo5P4Mn9m+8nisVSLwSRQ5DoxGToHrEB1JqYDrZsLxAPCLO921LFLnuFa/r80g3oHglG7F6XH
z7QqLS/rCb7w88veDVNvN03aIQwvSHEsbkt5Zo93zpLtf/Nf28M9C4KKOkGjF2yU6dvDQtYwLJhy
8rem0FDtE+N1HKNgQ3uW0bExaSogiX2pVpr9sTWuas6ls7uMW72y5sx2ZaopOYzVrKtdL/K/3qo9
YDbFO2WuLH/FQMYMAC3hSNoqX/KgcQZtMmSucQV7pukA1wYwEFVqoUypxjMarJK/BEtd8I2PaZh0
yjmjKB8qNFj/hP6TLfc2XXKg9tXS5KYk8nGRwt3UwzNUqoyONWceP5LhssTc96E40HrtnZwASYgy
R1+FOeaNeVdZbfgnDK880LiMU6iwxKsa/Qh6IkAgWmb3BPLN6/UBT70Zu7s/fa+beBqri1TNNIYq
0U/Fgu2mY2ES3LkWcQ/VXwwo+QKPL7yKj0heBaXrMypECQe7w8yNzztfMarTi8MFIyDoZtfNwE7K
eJ01tunU5uqiTs6T8/HTqsOY868r4DUrTD2astu88/w4Kagcu9Q+LlmRBHLV1Xt5OGLkIeVz6lS5
xCjUSPNyGZhyv/dvJDocltJhwsl8lY6W5I2WEBEsmDMfkjZHJlNnkzjBaTivwE5VlPN8LKeINh5/
W3ModAQ3DjcQxkU2dDq6ahgKtalw5DwojOYVaEGPV7pBcxnfy0r0pEi79WQFZ3hT6/Wm7B0k9OVR
rTgtoNA+fhVDpKA1gXaIp2S9TxO62qbNiv+X/CraF0fP0XwBRVJko/q0+mzECryrq4imDXOT71zV
9VCZig1IfCKqgJrqBI4lpz1iiIkRv/jI11sJogldfTKb5IQ3r2MunxpwFrmhV1X2WYJV5sefvLYY
h0n97qujuZgARls7gWFT8gCyD03vcmUieIce/e7qzAjtDiqfeS5+j3Tb4DwO2TGe4r+XZX7/y2Db
zQ1D0YvBC/IthbqFJ4pfMgFLNMRqCGd9DBVJ9ut/siau2e5rXH/nf3ERJz0uQhkyZvjCrRO+toLP
aGWObedV4+UjAD4y0QFSiG7Ql92ANsV9xA4x71WLsDmEuphljBecEP8aIXovXCHvkLX4sba0DA4S
CutkkhhQjl5MdvhpCENfvm5LdzaLh+GpVVPtgLRBYgvzRgShhGi2xLZ9xPK7yvlMAb51l3B/lfYo
2U72ltaEv0RvEvdE1dGlS52s1VNFjotYqIhmW/NalGiPi5DogNcAUPmQsw7aS9nP8zAlnjV32abW
yESp0amf12cGwVVHvUG48slyRhE0w/BUhW77RMsPEJ/U6grcQDRCym9xXO3eWWndGGWrga9upW20
I4aqFw88n6DHVLdIYfBgF9HRxLxnsmvrb9h8mZzFqpfeB9P1eoVkrpezRCOdMXJLZ/hs+M9J+Kt5
epocfbWWQ38E0NqQMqzGYzGPDd95JMzry6gyp6IpsmPk4M5aHtUDuVSGP3yRmKVshxDbstRgbeQB
61EyFPaiGJjXN52ZB+pQd1Sbdj7WC2BlQeBjV5A6I/jgF8XeD6a9DSpQwM0ZTFwss37OYeu16PPD
6hv+8E8RW7FcrZGcEgJkeicuC7DZl9o2C34fFfdROf0aQDdmkPKTrwp2P/V6hBliYcw9Nz8J3p34
Fxxtit2gIY+WUEnXzU8Lm1slhVxtO5I7WpDcYQhxv9+LLU0CnatKt2eilBb9n0D874SENZVzS+fr
qqQ2n79B/BzZObMkQeLQfEFXMn0zClubU3gn0sWC1c3WqV9E2Ri7+7WQWXcJyid5OepcxBAlf+1L
pYuAy0C4LfupoybHw8hJgSmUr00aLCEQqubo1Zfoh7xdg18kEZWVyjIj6jbsECrmXkzFTh5Vujm1
MXbLUmJMtmzegfzYr0o3LBkgFA+SfYRwAjlWS5FMUfLHpQInErT7UwUbToPZxPZox0AoGxq6yjXE
wvlsUp1Ks7XnMY1jjxBHtIv6QCq68ZUtY7c38p7yKQfLLfEGcyiPdqV9iIEGoWyFGsHgCkQ7TzPM
2SrcPT+F+44wV2LFHWQ+OSj6a7whzua2hHecXY/tlnVuroPrPsSYt3YSk3qoIywUoU11BO43aFjf
BjwpGNLv2rRjONeWctQdBho5AVT7/rCuBOlUU6snzAenOnzqkjoUz13e/8n5R8ffw5gdWGpioWzG
+pOgUYcgnfnbrFrGyVvw0SkUQGNDnfqe83/lGaJfmsMH160BJGgsf5aIoqNyvb3ommw9ubBL00B1
ZE0XphJeSOyzK1wAzI0SZ9t4mpOGVbUtjEIgi1kQYC9Zu/27GiE2tOmt94bHWedPBbhboCdy1KT3
SqRDEPwx5mgJWUBT4QOLmdhIUxNAEcyjCKr11msy6W6b3nyTHieQKo9jiED/KlyxBDQvgTzc3a8+
KHkK2+gvRNdd8qIPI1+A+eVW3XwECgsR4yxKz+WN27hhjz4MgjMZxEbdcOznv4nZBzu0XEK/2ha3
xG/f+L7mMiYLu+3nO6kG3p8xmw0V3oupb+Kh8thX+rw5Xb6dpUE2i6g1jS686mSr6dgftSEyR12f
Jxl5hQHNjXhVTiSpMm3FVMb0beFpOLna73QHvqtN6PdUvIiFIzK7mq6q3Pxe2cFZMpjMghZ8Fq4m
IGsJh0d8KsnDUD2KF/4zLzImPYo9LZTVji9xYqt2on3gAkPj8sPnpLWOP+pd5BchBXgyxIxh9PV2
vqCMJob1Ik4sbVf5ASjbh7o/HiaPAndgbq/G9VPRdXIYFBqAtF9Q2KdQYp6Z80mGWR09iNr/SWLE
0ky1Xc431XTrDnk9tmoxGj6trCBlM5MetMfkr45c43huOKZ6OrsUwg/30+QpLXiOP/1uXsVn1hBb
qGVJswY5+gMHc2dzzq1cegUb362UsZ8epdqfT5yF72BjpLnifA+vhPWVgoFfBowyWB5X9u0hK2MO
tIMvDGc4nWZG9kNNUm8jh0HOmUlWoV6gaOOUG2PtSk9XQvZc4gBTwcETNJz0TEmhR/iLC5q52jI+
Rr0H9vFJRkcMvKKR/aIeDX1yFvG1NI8x6NC8l8lQMxm/ycFIdW8LSuZ5ZOkH2+T6Z3kpoq8yumTO
LFJ8/BODyK0ENKB0BIh4mJ8Rz2VRKyYslQrD5B8YESTMPv9GgUFzH/xJyJDMAO4My5gm6ki3YqPE
zRWCnJtx7ZXXykKGHTk747Q7gHjFJHDIHStAx/6baoGZJeCK/Ob7KYeiIE38Zqv97/li5LtdESE3
jLwMHItCTM1YdLnpJwOTbt2Fi4rs22DH2EG3mNxrEjerKuSBiJxTiwfJQZgZb5JI6JfJUP0GCMez
5w+pjmjvOrgdjFwH/d5e9LvGE00YuiNVa7gOkhpj8TJYDazvByUfaf06mJwUFM8lrn/2QsrCeGHA
kbtVdqEAq7+aDs5nQfsTWWlPkee2Lmup/vxPGf2CONT0ERHFZe+ovS5hzGerm5wu5owGctSBnxcx
LfOgx4jH/0LzPwTHokZXK59fxL2wm/x1bOL0Urbzx4I8yBfY+BeGht6PleQID+lwYGBvDwQsWc5E
GxvORgizjR6B9Td9+LnKVInxazDpuNmrR9qaLANuFxL+PTVKznwkrBp4C5fqQLjyaLz+TO66gfja
6AlQ/waJsxz4CY6Vxp9U3X+rstpVBxYL9yzdOaICkCZO5Qjczcz3NT88lwKlCQwAjekd/dKxTliC
T4wuLZwuwjtLIHPla9OahOPgowbxi6Q3E+bxDAgBxNcO6XDynIYMIEi0/rxGbV/EelRhtdqADwSV
ARnzfF39HlkDVG1YVWO1vqOG+OXHqbw/bSt4XNqyn64qZ2TjjJjvqxWvjCWNlivPRPDBzvBDLjc4
h+60YOH3viOJm1RwVyWnLyg1u2ct/2onl2B9Q6gsp8eruIyKHsD6+BoBpYgLW5N9k22+k84IWxcU
HFmItP/cuvZHqs/28/dwyCOYBj1gdNM+mNvvGFjdOzR3z3razP5n9Kxl6ST9s+DptSDN+/pYbdOV
uJCwnnvthMLrY0HYcm5P76xg3FKsluVaMPv8LGUW6djVCUVt+xVD8ae7o5V0DXg9KwED9JI5hRaV
77wKmnKFQn9c1a/ODYWQ9VWWHYk5f3e+D3Ogkdw/TxBsm36XtD5VlhMM2zk6gRF41gGAlVIYlNZq
Q7+m5luGRKRAnGJZUeokhBULgFMNqT5qJEG9zjNpU0iwP64Wewb3Ef9kiibYSQDdDGrZ0n04jLtL
+AN85o5ADgMonMZR7wy3WMOC+NFyXcmq0aOEGELuTD8JrIsnBkOqJqUw26uOmdOj9ab11XpcDN+8
FbWgrHe/NRVvg5LVFBQC6S1uX+sYt2kPM9hITaEBxUwmX66neK2YWpaa+fCtIVr6A92rRK1W/Z3w
k6b/CKSIjHMLGulenLNGkKXXMGLIPEO9RQ3Wx+llzWOHjMtLQUzErOLMJmwvwsOlC/7KGxHprJkl
9RhBa9brnu86N2q4PMCvXQtkOJvEQD01+Tm9EjHw5gdnOp8hWLejnAhRJIibfIoo7hXrzh7vsWXK
xrwfZ1zgCKHXH4bATqzR5itutqA2rLO5mCRd3psgk5PZ+TaUoaa4lhrJ0SovpSNJrtEYKfuSgMck
6me8iPozbnV2jVeit2B4P0mE/cUCw6B5cYBV5/mbGdXXYwydlxdVBbKcCWcfYT4jkGnvPuqijKGN
Slxj64Y0t0mnMrCnKLCJ4i9sbWM4Q4PrHkFjw4O9j6ox1GAgD2y24/6EljTLVmO060gWvXXzinDt
P3mWV905UdAmGJ6vI+ucXSAFQim06n1JqXyM2xoW44fARSfFg02JT0F83QJ8gXBPXJGS0aw8r7HM
zoiAfOm1RCsJ1aFPNmTRFLnjxXMMD5Qlt+nkw/Uk8LHxK/pWXutkql5tpz/5l4Hm0Q/Cnx9/H3NI
POeFKPqwtJ1OEelCEd67GhkQ4BxFC3WlEZ+uE8lJ2NkjtxA4g0Mmo/peFrsFZnwC//ut2uLZ+50g
Vh0pIKiSFWi/1j/hNUxyaUsOPSn6frPFvj63j347KMafrekKBf37Opu06klf/vouxSFqHssDj9KQ
lZ9Ucz9oZXrzvtaWnhv+41Xbtf6n+cSMHlKwl5eQXqbvpdpfDA8XAli19hyV79SU7I0evgTMzZEy
tfWsJCpIK7V9AxAx8YX7PG6Dvt/+AvdmnuXWHk48EHjQQHdoJuekOUeB7y0U0bSPjk6NzRWN53Wx
zDI55l6/TGT/uVEiDAcVa/fdW3I7IKHv55w13H5h/tc4cgFZbk1u63OdqGOLLBDy2B3igljEGQPw
uz5qp9v/bKIHaDcqETsY3TRn1b5fi9yAJUfR/BO7HJtVp0hrJ8W2sXEB09ZwQrg2jUr7inif8BG7
ENhnx0kDsnjA3uwfO0ZdFeEYPRbe7IH59pfVB31d95ruILNfH75b0gYEToNRTawaCiKBEa4kQb2J
yz/jFiLbKMt9dK0g5PS+wIx2AIj664uRI/E0zBnJ6opxjRAeCjnmA/F6rcWFdV1KtIEOjlj8/exE
JU76aEL87+6CB23g+yFWa1RhXXoldyqxeIf1QQiq5yoWa5HYsdHoJwrQImwLg/lcZiVCG2i9ZvRU
Axk3fS9pDthNHe1rUi4lyL6NfvjVW2a4E9LFkVa8bBWNAq9Vz5iubajp/yA/CTxRi71ZqV/BB/lJ
RDFPLfWJHD0DF/JI0EAg1PnUrjN3sjgTR9iYEKEXV7a5Me+u/nsb4Kxryz/XD8BX+G3t7/WWfrJF
c4UvnaJoy5M39RMElcAkXIUeAcoKxFbpkVOaLE7KPXd9GUrA6zspzvEwLjIAp6yY/4wYe6rNtYT+
BfxGdoVaJ7C6QC+hwclFHnYDc6vqlw6e39AQsSMLW2c/fJ6/Y3lzinHw1cyzCGe2+V7lY5lEhyWh
y2JoU6gVc5XwSroJUUvYBRCEdLCDwYZjwKE7S8VRS6N9oyftgR8Li33tB/2+fkPinysaEU/eoiGA
q/kn05ShaA9WRRPBXV+TlwbRlYaBhVYIeeM5fsoTjj3WiKqtPDgb9GzFuAmwRlF+v5oIPu7orf8c
fBEuz+d1g9pGfunfU7oQs3c5ts9CB/w2+vv09OSWYxm4keJsxlkXt+SaljC3hupx4h389MXEVRcl
Odt/jWEWA4oDmk7sM64+UsRLF4p0rSX8KUAVq+fEZbXcN39z4MHpHxUQOJF13mlg3M5KaC9oyCrw
0xvr6rk1+Z0NJeLuLpOPt2m0NaOJiIqtsUinuQOsl3KPVnWTnjQjO9F3unmWqhl3BhZTEMGgMBCt
ffKyGLcwoTaQgOB7QTfjjQFywOJjE245B/jbiiK8YyTWN1ipnBcseiMyotTeGtgk2J3jDYzzXfUt
rDOkSYqN5qrfJgyfJshxdVW3xKhEq2HC7sdpK1kKRbOXsvU1fW7/ZCWSrfrVeY9gMOO0aInpCXvr
HT2wJq9gyQGZVUojP6vNaGgM77KY0ujjIg/Al6aiTPXWmiSh3d7sz/kYhT1/RVTV2e7QLWx0xk9u
UV+gEepVj02I0dpSY73UpZ9nmNi9fUHlYvMPkWDUbGDEzjGLHrcpd3i3kx5lTIUOTV6J1PYYzDPy
EjGxCat735V5uIsYhA64HPEB78Vxmkg02Qr4E2IqrvGZIMo30124t4nlAXI8ISU/OcNY+skdraT2
gx585th7sXNOW00X6Dt4Obhqddv18SYVY6X20tOV8/g/nzPgLo9qjyo+8GgJuKCix65Ldo0qscTo
wRQTkKpalRQrjk7cUML84grdOt+qbxS3RsYD2whevKK8Bj5p6Rdguhs09je1iM7y13qtP3JJ8rq1
LiUL113Qi5rVY4o75EVkJK3sKVb6pObXB9++FfKGAFZl1kAXmpB9s8Fipmp9F62hd8MdyOBLvx7o
W7x9POTj3wzsmzay7TxN9ikAvxkmkWOq/LAKyINPMtBqESnH5prRIc2vkeUmYOoSO1artLxXg+4L
RHEthm0fc5YDAa0SJSjjOY0mqWmPrOHUIyxfrSFLEyMTGcgNtyny+Zjzf99wtqwa2McWV4L5wdSd
u7YwIwbOk9frdAmFsVYBxoAgYGY2ebEm4YeqiO2sgHu6+HkrEb+oMUB2NUXxua/cNC2CYzff9k32
MDiPSDO8evPaVdkcHw1jPQ6BYWwkUTo9ht8TzRvXJh9MLENmYgqKvu8EivdL/LrE2ZOpSet79lvT
Gc/gnw8OIDsLVmNHdnMpQi4Jm0HHu11YztDAYzOs+MetVcPAGDz5y9YU9XxRP5yrFZ++UnuWL+OQ
bNdTZ9owRXIqaJybfKQ62uxaR25KTqcvQgyyqLw3BYz73vdU1D5rrFyqbZ0i46Nj2RxxtuAS8aMb
MOODMrAQVE2Z7NcrS268B9snVidTJL5uuo+Ce50RIBZIXKW+grxG6n18Mpa0sl8Lnv4Rrh8BS2PF
LY/p9VWLYUTGDzvmf72F+z45fItw46LF5IERBjDQkP4MgYhMJiLBV4HkTU+E+aj3IjholsyJKQF1
dV3oahl60okSdkQGlmR9rpFT7ENHLsLMpN/D/g0XJUWFNPwRCJm2HK2eKtjYj5RpjP0UJkDGJAiQ
WKffupukoxSFmYXVeIDbJ0tThho8s15nlDmiwjHt3KIykrbbS5+CjMKDcbhbbJoHhEmI7s3i7K0Y
RzcXMfIEAUvX056/L0VHqqk8dVpZfq6ljUhGLV43+uZqx1R9HRDrOeeiLjwSNpH8aBSjXkJQJ40l
9LDm0EIaZJJZ56PXRHBxcIMwCEEg7ny5LHjOScdbmnwa3YMyuEBZ04mHnDe7B0yB54zl6D03ceQ5
8mwG0dxPfbvFcgunDIjSfx0APeFp64uGa+mzoWaapqNFoAu+l6nggh2cIA4vc72vjXhf15/nyd+L
0+Ytg++Qur0Smhuk1LgwueQSYAgvTWsRIDLOVs4zxsjNDUE9SkU1eBDtgRn6WsBHxXkhc0dvNe3l
aWcGaCwzq3ShGvsNHIiOAhpn9bjihNsbKytArELzS2RDrnV+zXNI9+0JN40WNvsqBaxcx5nIlcIp
AXO74DvkejU3S/bwG3Wmjx5PSwwelB2h8I8sfxu9QxMhglyauBLP7mfSpHc9tBJona2Y+8XMNHtf
2eYs4l+cXWwuay5CHm3YkwEtwOy3f520MKJFYvv7UrFLG5Mrc2WpxeeMxzFdDgLXfTQKDJMiKKtX
gz2vOK4tH/KmhXY9nh7Psr532+BDjI16Q/WDnMMtoBuB8L0CMx7Gr60mvvSDH0wbx2EMNS4Pf+fw
6ufMlg54v3IsF9VRtnpgUCEb0o8sFOn9rJBnp9lrpfJuBJkzsfUv5x/Cs1qJ18F3XUPqchwEL78q
qIN+PmJxO5YWXgyAz0TNEuC2mE+wCvxInF8uF5ckYjeSVZ/a1tI6wGNPSXwzzUc8Ck+1bn9sJnc3
UNvA7t+game1ZtPgbI913T/NNxG68cZKg1qTYJSw1DtQ0oOmidjK7eWH6MBVu80TitSpiIWHzFSC
0ovIzS80UWrFPlAkt6HUeJdCFCBUj/ySNGdxvxXFjG3OYt1fdF9EKAwNUtRq/poit+SMyzaX2ysS
ryFnP0YDF933UnYoR5ssJsikZ/KJtcTU1/GTxgbi5z72XB+pEnHVT4ndiPHrGTVM+M5Dd62n6q1f
0b3nLOYy8OV83RN6BIBMtU7/2tCrTPNItCHZS8ln6bxM0VIT3oGqjQdgSGqHd1rYGe0m25gqns8X
ACaMIgHmT4C+LCEon72WtyCZtNw9sdjYR/iMbOqYFpB4ozNi4F7uMHSJtuMopT2YY3BYhiPSDT0g
Tc+go6+Zgl2D7goJmUYi569Cr6p7Lyk8pAV+tbLQq23JZDBxNzbe0DXA0HXm7xiF3VVrnblUoQ5B
fGFTOaf258siq6XPWEYe8lav+68iegpwTn1noeq1Q9hQ82R2Lwi+cQkP8D3zwE/YZWNj3NHswmIz
aDSQfMf3jwUzHyUwwR4z7gTPrI7PvwGEfULcBWQ5vnXWO0RrAx2FnjC7koLabbsegBWGt1e7sqGj
czh4XRdh2L5LADVKHzCDs5Supr//s+AFkXlkuwM0uX/gcQXu13e4SGE00/xP1vi+Vaf1S5Di3ekp
lNJA5WArbUZpHExMDrXNO9fG5aeM9t0bpcD3ld103RVtVh5axgrsx4avUbqVTMTPjDHAuo6lsPmd
BzBZdXTPGLjiUF5hUctFPCqRCiq0N7vJ+TPvWSxAwVXJwnwjkVUhXVLLruaxjMeDmVkL0UjtC0kd
jOmNXJDjKKkRhd4YcV2jvQxy2vbMolOAgcWNepOt8mMmtnG42nlJTfCBLTB+f0ni3WdSDwn7yQKF
T8VWMhl7I7z1jpVHD396Qf0Xup4IhKLd0jScSIl6KWc8IUZ7HCA2y1ha6n/6kbMsjhHnvr/C+IEi
W15JMbKQvSMKJ1FWcp7iyv46HUJHtp0ka08Q3jxJefDHXhDWF4JM1c30sBh4DMWK/a0Dd2nrI/LT
5fBz5d21WLguYBBj95e8Wgyipd84qUcG6jmzsrDkjkyXvVZftVmDZ1ouwILotxbMvV6YsvI84Fus
/0UASqo7SLM4wlyNucaF+PmI/PY8pELL0nhJCA6v6zlHsct6tlaTXxKbCJflcMlp67WuyIQbFaxy
IR+9mamY0rgIh2KDvdzNU6xjizxdMpgSOR2adLsnH0LK8RvngAIZ+IhPGV6/QZCdfspiX0j2vVZA
nfEezUznzZsJUyvDM33fGSKjREuPeps6PGJE/xR4/LzyIeC+Kh75vhzBbO1Qs/bpsQhelaf+km6Z
xrjl7Cb2A9uv/cEItVQlWOuHETqccb7eX1AWtyp+4fcxAVEtyVa3Omgt6SU23WWorPFS1d+jcb8d
0BY/EZUou+23peR1fvhqHnl8T3l81sMwXVS2q8mdbCwdq2jgGSQQcJEP9osh8Po98GGV1yz3SWUM
7JOAR++wYSbDXBjcn3BQYpYCz+63bfoYuudfRkBwOvE2V08uXoC7T6Ro00FN8eZ/aExA6N3wxAYZ
yD0cwbmKGD1InUvt4Sf3X/Sj6jIVaJG+SpEDmS+J+5e2xK2qvctrvqGE5nsJLKa/H810tIVhTHkO
rmqxERVhs4XvgJmJ6xgcYBGiakDqOfB1/G09R3VdMgwAVds6kCpnSnPgHKl/pa33RUrpPjK/ZeV1
gdewPuF4WKsEOoVANDCigM7Al5HRbIcgaUETdrMfd7xFPKdYf2DwTnsR/fDl2QbZQNp4HtnrA6G+
5UcEmZ53wKUDohSGEDDy1k7BlCkG+ilo9PV1dlcHBIEj9i2RhV+snxwcxz/9rBKfuxQFZdb1SbU1
G5nbABAanXdjFY/FPlvhYoVkUqqvnx5Bbj4YgXWeW4RWR8oLRNThorY4viF7SFqAzviW1DQpRLuR
Dqb9aJvLJHHEf039cxNLKO2AnEyidHpsp1sI6+ZtZx4iyU+n2YpHBpEFrcVRBXT5xz2mIJDTR7s/
PYq4ax5TotCP4PK4YZ/9fsa82TH7fpsaS0Wga++WvEkqc7JnGOk56T90Fj1LYrPSu4W25tgWjzxj
caenfWFBMIQ4y4qa7ViG8JkIp4qH2B5lIPxX9xGVudTlN3ZTJ+prqmghOrFLx6tjGS9eY6odDTyK
3nTh+UDRxJ6cVn2RCScctOkL6GOKPnADaDiFZq2iIWs2ulx3ICFxOWhPXUES2qdY8apNeFJYQX+G
iaxwflWKFhXQQZMYlwu2ZElLc/h4IR5n+UrC/c5uyS3qmSmF4I0zojQgV+/V+/8yJdf2RnA4wz97
n9q8i6eiDYYsH8aexSxUqwifK+hJ5qg8uWZ4RkoSzkjofp9i4RIRvZ4qMYWuFbXmvxzIEhI+wpBs
MldVqNObiluFBBZsoAvZhcQS86wlyMkwzlAA6Src2Io+iR9sAGC2qhFTdYTDTF49zp1aIFL/TGQx
zrlawDY/UrjI2sVQceQGTU+1SHs7UftyywsQLRN319BbF4sHjPXLZ8SG8rXHVGRnVUbHmxaO2R9z
Gw2zbGfCvspcV5s8Tt2tZyRrelv+nTFpteY9+y5fQGGpla4rdWWVMn7mWq7vbqRM8Wx3nP3h3QJE
V+ltlKFuzmJ1DhtHhStAGTTvfFCIrUXn2jde3t9oQCzTYOdy+AQrFvqHvpNB/4qwgGd/jQLD9pnn
RoNUXvAgd2UAQZ1zn5KgYXYtPKJr17gmhbdP3k0sGna7HzrtHJWnt7sIVBbRzq5ow5tvOEcBuxAp
MRjsH5fF6wI929ZxjNmV7u5zz036jpvwA1ysYvMJSCfG2CXMBN8WtocOIfqF18OzD12avAko0DXK
w5EnvwyYji/XJRLHW8d1l/PbvSYb1/lONRK6Nm6JQ+K63HlN45/cc/OhTnMHqXXh+UmUY2IYGWi9
u2ym+ga3goTb/hX0fzpZkRJbUJNa+0RDXoI5FIwexVJaRLJT/FxI8jFEnK7RE3ngRJOlXLtIxGPz
L56quG5aNF7ON3Em03p5AaT5s2DM1UfB33vy1MXtltu43Ej93fsveSPpI/7QhGRFoTCFL1Y2Y/1J
bMCBKy8gQKlO0UkgFjPi0Q178rlasRmXgSvbQOyzcBXSEZcQTdPgFv5UeWTcmfQV/Qw+BfdDpecL
qiA6TSfKZcy3oZp8XwqK/Jvtk500FsN5xap1GTBw54BlzNoXxykP38dFsm/7iI40JsazvRofTiEB
UY5p8rEDzAX4eHVU7z1aTBFWF6UDrOf9yoXF5YeXLwLkcEbMLoa3D5mK1f7R+qc3iv5Wr3keX4Qw
dXnktZDFvDMy5tXqg4d00XxknZ+ETHmi1Hz1TGRBWPMSRoQZxuo3WoXtj89ycfh++CZd/SogQubH
hH/q+vM2ywwmGkk6x+/0C72Iga0ZsTeS1umhR0nyJJeqfN4G0a6KyB3pTag0QGB42J67vUdcuzRw
CuoOB43Y8T2lgqIlBNPywXMogvZmHYBln7wp/trvbnxK4w3PcegKxVKYHZA7C3m3+xyIqIqYs5n7
p9Cyo08xuGy0T9/zNzJ40qHVCb52IYh7w1K88YI2NLWAYF0FMDxFM70e6p5T1XBRAEl3pBehf9LF
FZY36zUmVAWNZmgbNvD/X5Uu/QWWBHflrwHp6DImga8+BIvVNcVlnRpl5XY7FIorRWOEJ1eQGQDn
me31ymyTgDpFZwzh9gAnj6Q9s8O2yTrayZ6ilJII1gTtENG6M2ueQMcAVLBKJU6Eub/6cOETTPAW
2DLwX/BFS2Iwqrm/joQoJPXKMsg+5aNmOlK2HCfBVJUHJepfuoP5VeoxwblAZSA3A09BjQ+OPh3T
vOig6rN4kiVQpVpl6DqFmiqLrzhPwXUBLn+6dTKKBPEOXz6iM0WK0UiiRdeqve8VSpeFx/9fiRth
N453I2c2TO8DV1LMl+e8zWZnSeCUqcvIWSJpdf8sYNvs9k9qTFDUAPSG/IpJXxj4Q3a6lgLuR6Rz
AV58tC1r2yA5b+YKXlj6DlOkSz4julBoezq0fmKT3klgqGyppL+E93SRyqvlrTq0/6H9syEqpZqB
a86wilyrw7KeNCuuNRfnXqkGfpXu4ojezWH27dRg5fELbWn64wBfsY5weATeUxEO4nlfxbMbB0os
cyH1siKC/5O/3deJHvG7nVdY7sClSgwIbsTRH6glo7TKMW+4SgcxWKdn0nOaDtq5aYQq0RuBlhp4
aR0yVG7ADA/x9nYIj3tMJXLrTEVlckgGShWAk+oESbdkxkDkMFQKgv6P5oqa90GMnH6SRMipe1Y/
sNwWlfqG/wDX0RjilQuXnVoTsc0MrsUUOa9LfWE4BsCKW2hKFi3C6vO2RivSp9N1WCFyxFdjZzk8
6QOWCB2GntHH0Rjpi8r+fh4I/mDl8HdAiWhR7jHZPmCEIX7/VbBPTNFcNeuntXjyWt82TaWmSYgj
4HbBkWEgqYdIWkYQwpkmNsDtfSA7dXG+EkKs04N7QM+Nu+pP0wFUSovaw2ZOIR2z1mY8Hh3ccjGx
1ScYysUC8qQLTlSuKUwS04JlXOIjGGKYSRxn/JYo6FdfK5n6m69Z3MyIq4NWx2O6J92qJ0EbN284
1f6ZjShBcyIciOO7XbQesD8s9pQKL+NV3mwKotfUvcnxb2EojdhO5VCAY34yo53i827FpDwwitu0
+dK/FMd1MULLoHVPmaLMGzszYixUYt24s+jOECVPL6nwSW0d9TVbor2gmcSsxFa+u6rxHM9H7rdb
hX3spj4kpppPGArn6UDuwMy303HbFps3YaXZgjwtMO5sKoE6FnByeEimPbp7DNSqaN130CgULLqw
hMDQONopeTnSycchEXgkHiRb6w5QDZ6Oe5dkRYWYwIcDkDzaUo1iSPJcbN8/t/UczejZ64tLRw58
0Jw1g7m3DYwdrAMD0IjOmHQF8bxCxvyLWTipMXGx5ULcK/ycmQYVkD7xUHnBQj8j5zMqNhLcFNAm
pzEMML9f1S/0nfsWA6gCxp29MeAktJBcvti7SxFF0v8jTlD3502Lnk71VtbV22mt0oMJTXXqGAnj
dbkrrvypBWP+E0JNoBp29tYKuQH7rHtq/Vtkk9ZQh7RfsvvoRVVInopqD+xPQo9eUFYyyiW+4aUQ
7M0W3zHlLv5hGlgJdGLs6aKty1YfvNJ6zD5i3r83Xlj9RQc9bfsqmhhq3b5Vc/kLxP+Xi1eQBMAO
W3UZ7/M//+ABVrcbdPLNLyDqGHdpISS/+QMCW00w5xESRK/oXuE1lyyCxNPfY1R0dqJQ00Rz2tvl
bRWchQ5Kmv00D0T84taUG/JDF3s9vgekEbT+LAY7PQozG5sFGmhYuh7iXlTmNKMUlA0pELeUpmC+
36LMEYz8xmxD50k88fjMFfD68BkBs4rd5yq5OHecUq2Prc0UrL15PUNNkYEQ5H3NziktQWPjNtTU
hMW+ikDtcvLHn936/jyQsKOqwQZpRJoaswLvOuhmaAH4NoHncoSXItEKoHJtDHKezQkHNcxBfb1J
XL3Wf/K2XldUB3lB7SceRWyTlj66HxONecbrWPazvv68p9evNqbY0kxVnm2mA9b+wIdK2bFAIw0y
B+8jcGQ4xBUYfiK7jwLCj+q7WVcAhbgtUeMR95y7Pz+1uvFUKXtujnDeLZQhOBlCXUL8z5cjUTgY
1912ME/nOvH+1wBFxt6DpyxVLn9jZW/QIXxvcO2+pa7h7D/C4SUMAUaS7ILy6JyqLGzy9cxNCOeC
zPdyOU2lorqPD0EwAz4eCt+w1BZi51eyaKxSEX93L97/d+kxcrlfCvFQc9ZvYG+i/yTjqqkjfYTh
MLuGQ7yn0SEhz4qwjLRCOZBhmZ/WOe51r3WlggXtrpNtsyluhaSViUa492J4BZywnu99pCXKuUup
HVLK8eg3kuA0a9hW8nc9Qf9aoYhous1bNF1iUFbqwax5HCEYdqgktWbi4oybai5UQmHXPD3XFee4
u/651V3oVNNRmrmvGkVCgxDVpBtcCtPWQlhfp1TU9oQ3CkySwcig66FAaJXLMF+X2go24mfJD+ZX
NkgTwM+sJRQ9WyalnMMjNeW7nErKKaI8edLuNkG8MyqUY8knKHzz7qgE6XoELJJwZ6n3zTge9L68
ofH18gHgKrf2G4yvgRMEjCiOAgs5kJttnrxj0LNzlKnGmH/SAJYtDGfAgIyYjXVFYYZUN57/DR6m
h8hJD6DJ8c/xHdUlgyjyImtMxEQ683UlTMM/C0Yz5JaJ3Bxsaq5O40cWhNK+hA0VtV0kUvaDhyuk
/cyCXLMKLzdpY7fCuxqD/C3Z/d502iMD2JC5WKcsTZdjRFpFfe+jrBN7qJ4OaBKVzJDli+6jqLxM
G0wa2Ztnr9yUmZvki1nFxsDYfQYTA1bUO8jo79T17TTSqtVuEb15JvMZ9qOcSRownhdskNKkYDeg
K6WlQarMTDI42v6ciuz7Y9yW41cV2KDO4tQ0hYrLmjtdYNAfBTD1yIrkBuTURhwUQCFLyCFAR7lY
pKrmyr92wn+w3QR+0GHQRvpgN7hKtgmWde9hubcD/mT9pg8S9rX9QbCEiapMkO5UvQWxvZPdlwWo
723KQvDKO3HXzV7OpNY2IuiM2kovFCrXwaluzM3shvRhrx+hHDqIOE7vMqZyikZEfnvRt7dSoG/R
BQNbiHXr8ja7zyEQuscLe5xZfvJcNlDXkBZNDq7ZKkhM3IkfA5pUNh8wsC92gZ0lcROifdFiHaYp
7t8Wie1Ho9wEd2bEaTjHEVWtCb+3yASCJLjj4Gce9lw2JBCABSfp9eN4NbndY5Nw9CBnsVDqVUZv
VW5uVtuL8rsxEnAXaWQ8zL5LoWnYvEXSiD5ab7pedxd5KuJhOLQqSdg3OE80Dgt7xM8I2EDjNbYz
k0mKtC3wPOag8wXs3qOv8GvCBFDfk+J0hvVF3cavZOo3cYujvmLiCeiugnsJlUyny5TySsdzrUFx
Ucnw8GZAe7SBFn76I+XI13nT36NdSOJ0LdItmmVAevCoFgCZovBf5ICbbkjVcGTjbEWLpFQCJRdn
pKEofZZpymr240FRX7HMrmnKFu/fg3xAikEQBLT4gQJTSQiv1HYxep7yXaplPZYGuU0K8gpp1JUs
iA5KDeIdh0KThFbkQQwPO5rWV98jbeph10g4Gdap+mIUQm8qQY6OVy9j9mjfAdrz95z+m5Uxdc4c
O5VDXi1Xv6Idegq6YHiocjtsZdMuEQYv2icfX3SuCNwq7YwI7Mk/asqqqJB33L20Vyh/S0Ss34iR
vWk0h+NDbJpeG4v5ZvJaUA7vLnGV9brI4PnIiGefe0yUYsI9Cf1niEBzQXPobcWBsbRa62NBFzXj
8RRygRxN3a40MM8fJYWrg6STpS+jHzZqRcoqRwCpkc82WszBpEVcffTOqmtepx8UIpZjP5XXr0qy
8PPdcLhw7p7G3tnXOWp/CgekCjv59w96fzrhWjRJya3PgQb7BeujmXh88WhSth/apbtZ6dAvnQgt
voFJURFaQbuwveWOwmWo8j0IaC0jE4iS6XVXuFeysv059XxH02oU0yKmGbmbeEX/8VrJmky2fOvE
IU4dnWnNuhbOvmxlJftFedEjw6Nq9C8R6hq43cyPmUZmih+S7xgkdTcqiN6mJYthsHCxA+2K3Z/1
YRsrvOEI8AFfNo2dX9ZdF00YSAH9bj3L2YAq8znbIx/ga/ZlQN24lkEqr0nYjE2eMucx89qs/Suj
hcRcnwVfhZzwMvuIu9UEvl07eSdgpoZ5s/bw9XdEbz7u03oddRvbGJd1N+Byqj3iHtmmvg+HgGWe
ggDJaw1Ok0IWLknMRCCxVTm5H5kFg70/yQl4/4653WliLLdcdebv9Te5Pk8FtiGla7v0tihASBPd
vi6i39rPR7IhxNaIlf/7+Esx7lfSJLPaqcignuVo1Ygp3JuglyLru26dWM3FelcnxwvhBwWbzkNH
i39FaWisDAXZGm5bmmizLZWw4V+sp0XyY8v2QW4B1BBAwDHTRg8r2QWmJUMy4JXupa5NlP99i1Lc
K8Ai9ZJTRo2e0hm0AsXHZcnG3GyRFegD0l13XH2Nloc3/TwBdtjqOFULY8A01mLKSt5a4bi/9brY
vrr+pgxiI1mlMj3D3dYMVKdbhVNpj0GR1K7+8qi2JrzwAdVhqfA62EwhOTyOexyxhTVEFHvhI3LU
Czn91f+kMgF2dHQUcm/LzgEPWHPSylF3Ks8dij4xwGlsjvbpJtHiQq6nbB3XggOYG+Lk4UiA/r5/
/3WAfCbgEVHFRb7Uw3wN+vw0ADzltXcuka2rKzlEcKVR5VDc7qUht96+F2Z9pXrouq45Im5VI+P8
kGvZ7EejhYeBmXAxNAeKYTKn0c6tRSxA/nXBOV3gGvKdQVeRyRtDomgDdQAr2A86CyeKl3Olr9NY
U223p5PVNNOMSu2FwHyhe8W1JGGJm0ll1uKYSwZzniyJ/oebyG2KYagjZzPsYarYXclNK5/prz7f
lBPSZPu7hCAFyRTY7BiKbnR10kYes7P1fSDf3snh2zG34m08U8xzQ6KX/au30JdWG7DH0tlsro/i
fDeBR39BiYPbqhZZggg5HrjKhHVyWjVluREjUNXX0zdAWb84abYb9hTiwXJV/KCENSAc4v78PDAy
USO4mCFwkecuHZJOf8teArbJIZkPrCVX/Dawt3hBhZ/sdIppS6XhxNqgOwi4ERAFASaWxNqZGaTv
1BunPTX5B3Abi0+eI3cT7hXs9qhdisXnsrxDVAVkZfO2RIo282KebxOQXqitcAWlCSDC+VImpvHp
vpIRQtztxuAIvYu9LHpnBIIwgv8V6ISi95Ug3bVbJr7qkaF+dUWEdv7MjSLw4AtUQMk6T3ZbXWLC
0SpZgm49iSDoC1/vbmAtYfoZT4BnFB3W7C719vx0Zoo5C+kGNLfSF9HB7M6Q4Sfu01RZ5C0kimXd
iWGikFr2jlfD1NgjjJ1QKGErCJSpU5DxsnWYrLIeI6PPkX6DirgU5Wko3j5VQOoNim+3SqCDzYwh
vrOWqAK9ve2RSqdZu756eQebR34B0XVcDDnlbW48VDrUFoJ4dvrOvLWdh1WbaRnBCq3vlQmzFp6/
tS6FM++WhnX24/jDZMeYjblQhFOKc7ce+St8zo14BRyJh94CJ7D9eQPHYbb3iMc7Q+gjZaU/lMgv
j5/uBdW1BDC2BO5kf0HTfy7FS855eV83rDGcvnVhZnTy9XfL4G8dP214nypYYKWomlvkpkXv1zoy
d8pT1cv1Upz7bWu98E4mhrTY+qObQanyDgrPGiaV0AY98hDZaC1yypTBbf1CXJwalNuDq6w02iA5
Nmfr/uxSN9bZhM0UB3vxhnJwdZzQfSCkBDSSyUfFYdubyRreZiSsAvVfuyKmCi7SEKIjbFXo8wTw
GruUCROZn7JGh38Z1rquQw3waGPx5SZJANOqhB4Nu4V3K7GDmXLXbt8gRUfFD8fn8oN1Y4tXukMy
70iFOdIo1cszsJn2kyNQv5o+ygeuSXz6poKNJPcPFYuzCa/tfXsu9DdzZ5XTKYgxaN54dBhMdo7k
GzlouA06eknoAVhGjtc0pEOEVrE0NLLTC+ckgclNxLNBeJ2gymS/b3o8tkgOi7h2cjuwuTkX6qsd
HbbJU5WIarNeZJfaiDV2dQTI3qCQIjxqaiXhJDak/qQAvcKcUXbkLC5CzEZkRSQPudH/CN9gsQ5Q
pp0HKV2kfdDAaOY97ozuxtk6ehmyzn/ThbQP/6WvFZwNj75ldt5rwyaVuHwwL205D8mijG1VKPn2
0oSJx2N5WdHAzY/y2cw5srFlOWawMQI/mtTF7aJyb4OFBFTNF2tTdtU+kNCSF2QKXvcxaGP59nAc
EvBk6xrDHeQgmTsysxipoHkoAMQdwYv0J5EQ3Vl3kKeK1rLCKWH6XUf0Yudk9Om5gOs46zK0pwFE
X5e6BE3cnG3RXNFqeggItGdLWcj9kHSw2aPxC4a1ro0loOYAaiOi5hwuOzWZb0Rkdq62Q3witdx1
SRF8ZDJL3Wuz5ASjfC3STx7faYuYrYqDRF+aJPVA4TzZEoYALhkct4xEnaurfRiFom9eEwEvYdzJ
B7DU9g5m+4Pr6PQqcGxZ1a5w6DcgO+GTmjOP+VZZyzJqFiMfyPiDtQJMF81z1Vpglv+9lKYvV87b
K1YwMvW8R+OrnkIX0iV2+pB0d96rHAN2y1wR5z2F+WhG+d4ESQm7VIgLZaxKPitaWqKOM1yW5l+O
etdTb+jj7+laDrp8+VLJHvQ/mpn3P5Nn+uI78CCV2XS3jQ5uryxBsA8UwGeE6xV2C/Blx8YAlpZf
Yx9DO83gJrrO52+mb0hwQAbwa4zXNLUobIFR81iEFI0nEioHICmOIy4U6qELSP9Ur7VOFElAVV+A
oueM1wKUpmthv9ZBULlnzAm2yMxgRhZu0wdOMyJsGELkw8Kb7NfDEFhifC4UKvU+Vtu9dPayXdnb
Uj1M2xgLUYiRqNFjPqmrXANPi/yeBw2X93v6GG82Y7pDssJQUKTs3Pg5nyN3fzYuORWaXiOhU/IV
UyecRlgUcWYweVwPqDKa8oagi0HuzfOKldKs8oFl8gT0Tj4nTy/rqXMwa3z/ZsM8jDPfV6Qzfo5t
Y1bkj9MVsT7d96uKnKkFIk5R66yiTJBCCuEm4aPbSjqIwObw3NxsLMHZAuTZqVq1Ms0/VmF9s/m4
62ogyWMl9fxy7UGwhxvNco2RkdFg1UbJim3UlhvfY8Qh+/CBfVBFve3KCTr+CgMwn3s2n/xKkxpt
ikSLum7pXwnVb9gN6fZ//0Vs4u7WyhuMqc7JYGMwSaLGrFObL5+oPUK44/OTEMiAw0Xouv9bybpB
AchecPPZqnPegzTQmYYHhlORP2KusiuHXmriuCi27gp3aM7cysFm2DmHXPBZBjGGIAwA6gYYJYYR
fvgtenimv2nqVXXf4DDWY8TkOQtoc1ItKRSKlYDbIcZWaR7u7yBIOSq7JJOCOkL3usk77GIqAcRk
3YkQ4RMJxSaPY3KflW0JCI56AVxgUVwIxC0DzijRhSls2vdbfkxQAq4jkDE0P3HMTsOH7PRpFRrU
E1KMXcRfLptPAsbUmVcYzmgiktjLds1Ya7Y7Ys7nHCwGBbzAX3E2TKbk4sJZW55lFQ8fLG6psFSx
gp6atn3CsEHs+ZziOvb4BXcFLcqT5r+DjiVTMeRr4Q392nhnaph0k4z8LsocElUBfA1XMGUubwU6
c8TLqA9wVo2YMya+RJK5wW9k+xcAWMnxmj+v12xJYyqvIzGTqRDvZ1ed59NKn45qNf2ZCZ88AMMp
TGbHYEC1QgoFoIiNHOmXoO9kmTLO5erHmBlL5xQ37snSTzOcr3oE550RVl+hUSbsLyJ1wW+H+GZA
Yb6oENPH3snQmFTLDpULZUERg88LyCKiAzMqq2EPA6Vrjwi0m82RwoupLeQHuNP0gKOCk7ZvvY2p
uxqMxeqtgaDqjQblx1AXF8o0C1D7OIpLccpFpwd4ajjpbbs5RHPblHoaNtpt4+edHY/OmGwfKXAU
RomJHH4KheEHRQTslABTw8MOWIk3uNUhv0NWwiwqV+yiu+FjMkSi2NZZDjLD1Axn6HQy6tWDRCYj
husbCF78IF3YveU+nwrUzWaHmNFwwWLAyigEr6HLF3ol1MU7m0kmwjSdL1Pqc7Rdv660/qBYGx4n
xyp/6IJMhxUpvo5Et5BMKOfm/DqDV2xA4rE0aypeZl3xuqfKa8mtT8EWBFZTw9MqPgCyAJ3y5Ule
tSr72aTqK8UhAcCZDLkj2n5W5WTwAoHADtD6jnjIy2DxnhVwjCQ3b6hOu/LErILLWJ4ooxtgh2N1
zowTc35Zmn5e+xJQ4EKF7GPWptoqLxMtOddV8fxQYqTwRd/XRTWgGlKivyEIfDpkMy6oGyg80O9Y
W9TzzgaHePh1ONBtjCYLlHzxG8skNcSX2EW1o+tKxO2AxU3aONZwDSu6ph2Rgfaa6/H9l5JmWfOl
cJeMYZF+RTi6CB8yPoizQfb+Wo0hM/O8lFUYPOLi8zq7ruYsr/Kg9LA6L+ToXQqbgVOW7WleAE3v
lIxkRfq+tWDL9MyAp782eWtZyi0XxsABCC0cSr6Gj7NDwJvPwPPOlrsdaQ6FzgGnqV/8U3TH6Koq
dR/mFmBKLoNGM7+XQrYjVFndDgyoe5ya/KZdMwHJj/R96M4wJ89qQnBqkrM/iLIAF2R7/eqfLLuO
H5MLNBdQouSZvcDE5e1783iozFy18DSoDBYU5vGoG1ppQKXzaYm6N3LtLpm9/TG/ztCP3pOnVUsU
sabegTslf3WqczAlZ/c42x1tlNuMVHTR6uuWu9mXtub4w53NjHXitVeRY/Jo8kECziMMZkk/gsPJ
TrJyIpak8d0ysO4AhYolM64B3c7uJwt3DYvk80wV9C3i08BBbmAyb03JVJ8zWpgO6RlywSGsreap
9sW9SLkbltoDK5DxSblTQljUIKKWlqYgQvDRVBSpprcTlh7TWtStvbb+nG0az0ZJJqJzZMGb9Vx+
jbSPOgvqdhczIbNsI0wDxT2S8UChWLiJxP7eq3bpUJCz3+0+Vhw+tc+OHqFPQBboHGIL3pwR1GVW
3G018AhFJ8fBypeJ0gXB4k0hAyCMPt2HHPDV/T0O22q+yi2qXDmOTE6a9AJWjPCmlcJ/CvX7DdeS
S+nPhtKiHW8fVEZxXo+rZ9Br+ZxEpcxzvUyDqy0D57pA3/mS+KlN3a5G8LaVd0tdnY9YGDeJZ0sx
5u7AJgUKWl/bfkm+t9Zi8uEaH5WjDVaUtV6pOFPNCSeN0n34PWem03zDlWINepH39Ld+sqll6gYX
2FdSZNsg1pvJOC/gof65tIBq0FrcP9KaWJ5Ccyf3pZOhtjqNEcXg6fG49g5om6iaqpRVaT+AtGRQ
4rVGqP5MzUiDbB+Fzv+R/Ff+za7lXLWMUTEuvIm4Zu0HAdoz2BZtgizO45zq4K7ie7vWcIMbuLqS
IUnG4k2mrNXYmwHHJG4RIXnmjh8T/1E0QiMKZPoXGFK5/h1xaWTPDcymKl6UksvJ7I105mZGfhqC
YNk2LAA5wUQHb2YURvhmOziK/d62wQkL42IR6gtbCU+ZXvciBM48sU1wK6yLPjcDK6HayPBZdbDk
sattEaBm9MrWu/EQwUOEg+Vnq2rrUfSaeO9sExYt/Ka7JoUNi3Pua2SWYFadzFyHJWM/Nfmwbd9y
XyKRthaIyGhMlPFlTvLli1wAXaWAOqb58QOo8Q2A5DDKA1SLXo1+Vn6comlPQOsKN4Kd3g8YdPuU
6q/W76R7cTjUi++aW1IBt1qgnHLVFo1K5YycU0R4jLA1e38+DIk95dJxkqYkZ6xMeQlrG6rSbBtR
jzp8U7d3VapCeDFthixpu1Dvpiz8ZZG4SL0LP0YDZSgumvmTCdVw5DBItuAMaCZIm1r355NJ/Tck
T6DO6TntwV92S6lcZ1l6LF4fKGsR9hG6AAXiWZVfjWuUthSIv1oytk39bfZ30OcNLaqEoFPcAB3j
tVoKdxtGtWH/K+4c4cv6eKmyQCKkkv5BqaVttScna4YgvbhRCZN1CP8P7YuvXFv5/g993gTMTR2c
cj8oFCj5x79I09IMobA0DRHpTV54vZobVwGVUOn2zDshop3JE5jngUqXNJNpedoD7TBO/1/WDo2W
vEKTdTV/znY9vxHINUujdxJ/oz+yYgJGlOQNWbFeSKFvP3I2IfIJblqTBSiLqrSMtjoK6GL5YNCH
ModGrRf8t+MAXtgpzIvmICXievdUG79RytbQ8DgYna1nQf1uEL5KiRWAQRyJB1OhlNjgbOsbAorM
MsLIYvwYwludxzSnaVH++A/fFoaYSJI2qPu8wL5nBgPedQRuTp9f8Bv7bK9951jHdR5MdL17mGSE
2QdfyR6Svdrx6T3UTVtkJQ1y640rdX0Z6/QnFZqWyLUkyj47OneiaH3mBVQL6AIT1vZ53yim22Gp
vqdqVifOc1A1NRlLkaidibiWpI+iJVBHagMKRR0bBCgI0oLypxy+wZkYaQO+g+YnbjpHRjnsSTNm
6RS5uwsv5iyukDoiPkbFZ6JjZHni4bWaJnrE6SLZTkkDIfHCuqiJFmLA6iB8qsuwfC0TNWA7V3as
oLQLdVSQI3ObC9CFzrw1jQIcqoMmVKGN9TZuYNypI337d8QuFWWneKJhKTayWwwXbPx4it9d78g1
FQODvIj4f2pruguIpxgx6uiG1Ireb6WIXF6bKxiXLBDtBX/Qq0cuTSRJDO6J/v45fXeqwuQ65WdX
hu3LRVv2Oh3YoO31t//50hX3wLFzH68CNDZDB0zb05UD5goRxSET/10BJpxPU3uF2T8JaDFsjYQv
uf6r27GaSrFqQBzCHEvTG+jkEKPUkbU0q+WU7TkR+EZEOXu56TCkDSI28A0QL6nYNNi5OvEhkJXq
gV7pUxpkZUbVEBilKOZUj4OrfrlPtq2r+A5eQ3ZHJGSbBxRIRnVedyuedeSw2lNsqgw1eX4nqtLV
UxH4aFuitkrcpwd6siRpLOZSSthmHPw/iGCXMRFSe2uL5PiJLOXywFb0efg2gF14G1FBVnDkReZw
fe45ZhFPfi6TWwHcjate+YNRFkc+BVMDCbjlJZ63l1sYpi+iBOyAtyipG0vf001ahZm+Vukn5QsX
jd594mRYXvINBaIQNNttuJaK4MVt6L+I7CAxOMJ0L4alHkzSHlrf6oTD9pKDuS10oAHqv7+9tvsh
nvu5eKXF1FLx9wf+/YQG4BnR2WMb8/aFcup8da5oFvFwgHtxjVFeJTODTidbnCaHcuBZwV//Zd9E
0PIERaFKbDH2Xkj7wpU1zznesVoVYaufRX6bClLiQgV+OkQOfmXR++zDA8tjdhuVYlyzV8R6oroj
IHILt39JUwFMpaJ2q3wclYcVag36cnEyKVtZ4izl1uvqEN7KUda/CEV8iImnOd6eFFgb5V6YMZ6C
2ScZnGCGJufVcwZAd42OuQrPV/80h8U3NLO2rad/HpnbX9u6Mxx48JUOBw6wMMaeh/0F+N8NCf8H
DT+Ifl4/FHyDn+JoCl2+mu98Kqtc5WAU/MCo8youz4RvTOx1qqI8wZa2TeuiuESd11NBi04wE9d7
lKBcv/7SznIhiD1J4IVvdfK811CxDOApchXnypZpd3CC5lVYcw3pjwqG0+aKz5vii+mejFxbCoQ3
KGbaly3sDWjYQsd/jvnJ1EBEedRuUdudlbW7qoUv77uGrVzm1m6h4jefKu9ta+/rt8elHpxkXIrn
O7+kadUlOZy9MemmD64/arMqIbjZp/I7q/MYjdAr2syX5BonGQN7r5mnaVbNwXmGF8IRVsZeB+42
WyzkmeRPYv5DUA42claI+gFBHkMJ7ym4TqJ/Qk9vO3IHOFGHLVlQoBQYKS+Jor6KJkRf9TH/ZP3l
8+qTD5JV4hlvBHiM9k0JNwQh80x6pEwdd1/pT01MFGlndbcDu5T1yI7ISLFYo8UVArqdqLaKZqr3
8r9hXD+ufN/ZrBJjqU1E0uaz8ZPYrc2GWwfpS+wn7pGfYviTmhuzr1lATnbEkZkYhJPnEzHGGT1E
32FXZqfqsR8Kddp6IRqLqANfa7ifkK7hh8VQKA1op5sbGxE5/vYnJfDzwuBOjIIg1ayGCdl2GKd6
U1VuiIXR7IzytazzZ2O8JtDasEgWrknf/h/w8QyTGsVXB+N5vUHILzfNYQYqtgzOIDNyIEBg7ReO
kOSWW1MbzLwMohRPCy/Q4j4Xvo0NjS6Yqo5zNOuLdVrzx208ZdYpjoZ4RHBeO1xn8Ek0UJMqS6A5
gYx/m9X98nRof1zNxLvSJZb2GbiJjRWbuwFP5PySLZfe3J3PpKx1R7YkkpTCQ6D+SVJ0HBNT6hHC
rmiD6wkA+gL9GFgvtS42OON4CIhxogy0GLStB9XvvUXh65qy2wO/rzShw6TXL3TVAI+xaB6czEg3
GbsejN5/w1EjNOM/r+JDVvSjDXGsrkZGlprsnwzGiP3jgqkuwvE1/oRJU4bFWfLza38ROIvGkuWK
RGbk3TtRL2Np+7YYqAVwEhJKbPVNchk87C/6G8CDwzD59/nzfGFA7majdDQwTlhe+gmefyg1jCPY
Ke6Ek7Ht9OCs7oZdl2Ie+7cv+XD+bLUmGSKHNnxCEu7bPWResubfsUK+BKGf+ORidVz3mBt7XDei
KckQToD4wRcVJjX21+cdWlx2XDt0RoHFe5G4rmcTJADU7PjbBSuwzTVqCLeeIRqosnpPINnEeSI8
E0hqAsqJQA8/jM95a4d762j9lLp/wrfOJhk7ta0zAy4mAW9W0vfqLLuS7QF6+V+9W0d7UgojzyyB
2a03qilapKy3cmLLH5A5F5/RaPgevaALVUWL7hRK12dq4k2EjlbxSQaWahKP3YFaByI5/eeHdZBV
JR15FCR6fkT0fJJDP4y+oHDitxPvvyXnuT+nsOc1zUuUgiLaO1zHhHBMMv+L9RqbKVLBFf1HBPgC
asgw2/kWUNqOY1ifMGz3w7bnJNCMtmmtFM/zQ6dsRNJAPnbV7jgscNq2/9J+EzAGwrSYnkzjcxk2
qtNvV7JR9OcMB3ck4QhAFaHsjJ69JEs7lQrZwLc19rqVOP0unjyMiVRGE4P4P3J//YWBFP+Tqil0
Cty3H/XK1kl3cp+gKznkzVSdMZPbHs1fOrN5CutlMz3D6Hqj553DYdEOsffOp5EgSJ8E64wpD9wI
wO6CMKL0mYrnGnfyyJwFVjp2yKrBHveIvxZDwzLZuaRRMlD32BDvRAIDkbfMTpQBdA8M2Kuk1Nrk
jYruwKCE7qtNp9p2U2onzrAmbxEiI57MHRP2a0XSwyrvWCcA5Y5xK2fbL5SoO33/e8H7GJzN2592
jOicIaFLhBOJQXSmNPtcPV3KZF23SAGDTyqBpMSrYSOgiCQPEsYPjceW32AZnhxvUeho4UZt/dBF
+yTSAedTXCO3cxLBYPnReQLwJU9Cm2CNiRAw+ChR1xpPFwn/TS6zSz1Ho5pA0vmgmSffQpFtxFLm
kqazoWBAemSHQV15oHWlTZoH+6O3Vvik+Fmtsu8Pk4AvGrNxgIdF7dMUwZexoyqGyYD1EE8iWV1s
FEoe9iUXgNF5QPgtZDfyqH3RHV0KWulMtUrn95ft8j38euZ3iWkjuGqBJfQHZZri+5O4YO0vDxbz
IpaezMirv+yvOfpSfUQ3570VrQMHuzE2GK2ylpfoXtrCMbqOqjRyVBjY6aGpO7E28ymQmx0pyO/V
fVZ6QaF1uYQUrd1PyGpFIDHbNLTi3DXztB99jnRNYSkLT4gfTy3NerNrot0KOevF9YfzUAEbiwj4
6pG+LcMcEI33e+oeJiJinUrMmUZTJa88V0Lh8kaqVfUtoNAgFjIR5DwB9WIoFUsd3gGw8mkgHD/p
ktHlkg/Qrz2Fn9jAh0tttb0bLmAiaQ9EBPqgyutkeIn/kEiXbd6ypJmtRfaUhEklbjVuqmGjs4By
uKkmVz0FXriq/jK2qHMhMNAnO5x3qvzJ/m8yV0+gV/8IMkBFpgzKhNYccNIBTGM/i8pzyXmaz2eI
IyrwZf+uiqjSCsamlwwzMU6GQ1ukRu+sjksj7/5qlRRFz1orVoNnZsoRjXOoA9vIMd+kJXEsO4rx
9siaq9xWaJa5PN7dcn2+PveIs6Qk+06o5w1t00R4BVHgGNSjYEgGaXCi5CrMFSjyautjmK5acQ2n
ncURAqXUlpbPEB96xyrc9FQYu1HnEu8rxtn3qt6IZHlpwmimYikQAjtf58H4L/oIwtGW8hf9lcOM
gq/agdTtBdyVO+t2Uc7y5N2VY6z7qC0jgZHG+4wCABdJ/ywrA/nmnGQAfE5ypuXiLxpyMZCrScbT
YgOIbm/oFYO5GJ0tBVAwPSWwBom0/DA+M4j3EV5xNs0x87fITXNxcGdtc2GGN4Iu5rGm0MA5lEBG
SwLZulClxdtu0rm2IBgzmrzLEc2jV9WMht/nUIwpOrr5IErlR/pBuTmzQtP/1D62Nvr0PS1/1W5q
KUDGapDQTG3FlA8FNRiO6ZMOIHisHnWcQuTVBUFm6GzGzshB458jd+1govB9CftUIf4HgI6GK7h+
0fqHJpkf9EEFYJu1POqPrXSCq0K70GvkJl7S0LK3wraGRSFUglN3P9bEpT2llYaIb0dTwoGX5DdE
6xOD8yWbsNjx9ctzr9mw2eudD5c6BmMZpZXo7EWuueBhMr3VhWTQCoMROF5YVDMRQDexqMm1EvIy
4/nN8LwYqhVP5ToL6Cf+i7rL/SonIleE7bioukABE3a9Nd/FtXvlZfRdBvZZAuxSJVcSO/7AJoz+
kP6o0gbT73JdNIthDAv6ObCi0PK1CZZVlQ+A6CXGeOAM41tirol5V7p2lrvrBSZcpgfqdfFPDGJr
Hp8kvVIZqSd0ivddvNGEnlX557yGNdTkV8RC0dMvFa7rx/jm5ZhThp+agJyWEZCMShjm0RsgEnqy
AGgQDfnKsFObtjs4+I8qW2CRtOanOH04fePBJkqViqRumPfjFcMGdbXIysL3xKv8J9MnkXj+jj+G
m4kbm3NoQJUcMHMxfhxkn6b7oG5ucUyqF0W/yH7m/Wa4nUYUVCZ5FXRTo3dSAWlC95WHVU+pyJH8
8UZ6ElQzOFniRJcVgO7xsPVey0PhBcq77mdUa3YSxRWAgQgRygh7xFd5uMjERjJMSgn7yvIlAToG
+hCOJ3dGZK9FsPnbFHzfHASsoRVLCkHG5OZb9Ht3z8xB3++gHP1KGiIdHIYNOLaCHhw2ryrwd+B1
Ct6+Qgj4+AbHyVesb4xuIqlAYzQbp6rrJpXWdq4sH0r99IlUFa8LEXA3p82MV0XB8Hzjk2RO9I/D
nvKEHO8E0JDawuTxONBO+H/PSq7RRkrPHN6+3dpfCyi0pufobOFk8n6gPp93SoX2L3CIak4C/ws1
qhKxF1oPipDEUHHeTxmMWDAJX6G31YxTZXjf79OEM3JtKbEXkXaOMTY9vEe3ULYlrDVhGxPxCj8+
zx0FsHknoCJhjkA8oMMCi1KLUFapMy3m1c8CSD/XNjs6J4i0lSJvSZ6WJY5sWIdq8MD66osIfpaF
b1fEmxXEkGfdDcERR0CP38KctWOJShYse4yuo91m/T3xDNZ+YMGsIGGNO4tAP1qNKvUTGsVbFmyl
DkzmPsytkRnb02RZg87grodn1cxbI6W+z5L0LiQO6ZY4jHDkjR0/CrvCotSZOopU/8fu2/OBCtUY
0kNW5Enw77BQPjoxecrv9m7ewXqcOMD/UOWQJutlHmcSvYHqVeMjm2z0iDAjOpehglgbGThUdBfT
zc7M6W+RjBRtFvwSL4l1VqM37bceDBLf3xyY1MbC3S3bIHD3mfO3rwKgdDpXty1IFm38fP5Egtcm
IYEZdcWQl2XB8YOK/htvA1HjCYgGY4GpqGLs/3D2dZjTt6KUl+bs0SHobE+IMYHyq6aSmKXI4x7w
M81FM/XrZ3iENdaiAcyyJU3m0uTWyPdbsxnl6V4BpZPhvYjquZ3+2Ps2RC52RMf/stPVFNi/2CrA
aP5AIBaYvAhfWDaLv/rVktvJoRyZg6us1FLEvhVNpj7K3DmNktdVnNGml6Ji39fsILRBB5q0zCRS
IAM8UdJQVsUjP7eSTg8DIEkbROaoDmTS1DlwGb4NfpWigMlKObXeaJAz6wXmyyoPMoGW+7DPf57s
aEL2dzsSPVxYuxfQPSfretC4bEblveMXseOOwVVKv9jqi522p35RBCDfonMedjlqSbhW9HiNlcXK
Vcnn675v+qco/kFiwDsiEps/j9cMeH7n2G6x1KEJSClf6JUBOLFd8aKGpneUQyF7jSMWxYaGy0tV
s9I9BuggYQdE8/+uOBkS0IRr16iUlEXPtZ4OpYjR6gRAPRxyHR/nzgsVaDanvRJDPNUhICX/5L2W
vsekwj+bqy4Y6nfvY3dEdO4MXq7elWNPaccpW9XXuihw7POfDDgxjCiGScFCyq2JsrsJJGL+Fa0+
1ErzrMqu3vHiaGy3QcxCXBUVI69O+Bf91isznZpw3A/KWS80HACEglpqVG1ZXfrOy33WHrGuOALP
Duz9ljU3Fb2HbQcUPBbqf/aIDBLe9qHnNEY9VEqzRzJns19NMo7dr4zmUPGdNsEDkZpnc+Cp2Lum
Lrl6mxFEbQ4mW8vHKIVrHKJQUhe23Inacpzbpc+5HY3d3U8bYhY9Yu2RbtNpCTPAAIZXYlIvM0ck
PGq/6vyLzM7pa6X9AmMY1eE9Zq3BRedIq/rokRdiheWZJ1vXX8OUoqh3KcAYwQTUed3Ly5T6QeXV
f9kag7i6MUJ8EFl4tEQ24H6O2SlhGreI2ansZypIXC2N1DdntehPatmeglPdiXAop2eJeLmENeDS
SSWNmH9n5j72mR4/qCYA7f+zxDTWno2CBwUaFIsX+bx0PFqccyNZnGCgZWbCvjrSC27XeEMD1Szv
jaETHMSUclrvwx3ml96UaWwzOITbhyY+iQfKK+5H63cyaY5+boo/7ddI3x60rjnzlddDCVZb5mmv
J1s5LeU8C3VoanCK+oEfhcHbzPiCt7BgMAwq4WqJuclvELLsPZ6Sn72dTVkVrk6hrIeabPMKs5mr
v8HsVLDLup6NaoZrdY754j/k8D8a7uSAeenEZgFbJZAQHkuoF8OSAH7wtJqrMIsmMwHjxl6Y1R6v
el9DCs+IPIEKfxe4uZDbN8jdZLQCRHSjGgtq7eoQQPPI5jWoGySYQBgOPStrTGlNsBz1t6tZg+Nz
1GsWEvFA6q3CBrhfrA31a3fTeMrhudpaX6nGDf/wEmTevtsaMD2TwvVq59tGPB0vs3Rv5Ll9jski
Hbjch0puHZ5tZoUDxMi11j6b/wC1Pj7ThTWuZ6/Hda/iyex94YB3oOWOydUXcCpkktNWPx4A3Tzk
ma0JMvG2R3vFSNMQpj4uJM0Xuejfxn/DWjeXTtgHW9GC64sGqK+1pXSWiHnth6cEc5m93yd9L9mB
kDAdID+SvUog92lTdDRFdHecfIFzM06CBZzVqnf9iRTJjPvkdVMxyCRllQSzt0fLLiHW8JJ4SjaQ
BvDNYdgpm0+6aLc3xnRTQE2ssZrFQHYDegJxpNptjSEZNaUD26BgZCcLrFmEglQ8Yu8d3Tcu7usi
YsyqWEgjVsRPdGbmLjB2FCD6ggU5X2qRNIaVGZdr+Kr4rhu6kgvbWLvwIUWC/N/cg8VluxK951Yb
WVfriXDjOpcOzC+AOBFCDVo9g6nKUlXmJMj1AKcmzHdsEuwh89UCo3yD/hANQY6gHxZBw8IglKGi
bVeICmtnG9e7OxBwSLI5dW2IU+xqHziFFTbhVaXxzdJvw0VFkL+gH4PLJrOY6VHwJpyhAKGOrvuf
pEurobjJXDWaM3ceDGscDn0m5vwrKudvW7LQRPY4rxuKcTUc5AQ2eOnKPFbnie0pCj16mph42InB
Ur4dOSK2GmD7zVtwCvq08EYH5Lx9nO56Tw4+irZlvh/lXjBb0iKhZD3c//ZnmmePxQ2MVzKaXtPS
Gqs1qJEvypVpchPIXeHj1XT64ScIgaV8DI9595j27s+dfOv52qUW4efuSXlZXMM1j0JxRRzma0SB
qnaoaGcmEUmMM5GD1ClQI41MRk2CoDKo6xTiTdqr5/UekC27NEEv5ZqsOhnlza1qG+lR1SBxF4Qm
qq35215La74Mgrw+8Hw8B8CPXM5sT9DlfmoA64cjuucgE57XIe/4sqJDDNcXw2duXotkudNvBqOD
1MFhAaRa1i9sCr1f73q830aYIP439tN/6YYEO8iMvEzS+XFYbnGnMvvauUKDLIh41FpIVPnHuwEv
d/JUZpGy1WEPMaTk+ChuMIQiDUBv3HQu39HxJEKwubKQeuUPzTHWeUDgw7d/oXIw9sCxCnxAB6rE
Ov8bEHnqqltk9rsgwYqYkqqLUUZB6ORIacf0E+y6Ipm73F0oGCutBgeDU5SFD5146hX4I1LmONV6
BaDKW+QGP6j139cuEaeDw7+dP9eY/EQOv49b/uvqGK3PYfOwm9o6NU47pJP+KdXiw6HcH2GkpTCU
VkbQkDG5v7+UgeljXB9tERyuWVQSbzFLqf9hd6G6FyOBuP4OKoMwbfC3XiF8mEG85FUS63DHecqZ
SrNC11wV6AYuUZGyHsavQcIEAMnLPNfHyQ5x95UeF3lxpxhPioLAUXs/YPb2RhfIgy0XAuA5IQEV
NelAXYDfuQPH9RcHe00UuvQ+6JFVRKyJ8Junjbg8BP0K+q15X5MPPSQL0b+00bGQbhXeoZkNIzb5
t/1+ytkNIgSLF23Jo2umKHtP1b54+wZIXHTlo7PSHWSaVkazfk1vKfpmReAB4AggWH6PI7QIV/L0
US/5fLitsrDmjWrc4RleKUTHXUJwZodWQZ0YEcKv8XpajQ4a70l0LT3WPxs5fLBVlvfWXNisqwkA
LQRfxkN5XvLnVeK/svlZOYr91r8vWeM4Z6iUQ7e3wnDAyDlYAPMHuD6TC2WP+BtGkNlNKYA7dqji
33vSgjjy7bBfDRgN4Ot+DLtY3pc0isbHiSk3AUjugHvesGLmML6mSpAG8qbtX9wipOv0tqoew811
9/1KLcEL+kXatc5gQXkhX5bLrW11KgLuwTcT/qKNEmaGjUBsZKeFvyK2Pp57p0kflv4ZsKUH7HY3
6KglQ4z9LXwP0v5EuOCLqenqMW3g1Z+fpF60AYLNm/pkCmn+rh119pDn6djhVxs4/0URpSb/Ie12
xJV+y4oyJcdfmYTosS2aL6RycLzbTbYIpln3ALfXgUKekfvJb4V8j0/nyI/aWkLvtybl+71szXm9
t+KdEZBblVJvjpZcESNfE8BzMV7XjX0srp4GQFTwgF2+KAhLyRfi2iCeP1vZ9NvfOFTn1+xl/edk
XrmF3gZcIIWyYn/bZXcBhGF7gZqpwRdXPgWYTFMrjD+axtVyPj2jDcyxvm4e8+G95Lzzl4DR924a
16ldCZWwSeoPgKjjUyXvQN+aHME/MaPTWyaUJ+XEyrFR2+tEN3rZYLUymWr/2d471U00rVpLyzl5
HxELruX51uYZQLx2DDP4vK54UGkhE+G9rHcXyzA+GQu5dl8uQVw6h+03rX35kE6SpMeZ9/rWqpnu
uoXfXCvzJ6q//hB6TmrQco6yv/R5vO8Qke5MMxqGikggP2Ua49Nf3N7ICeGB769foEp/lqS1GLxr
/7oy/faED5fz9a3aleyHMz4uY+E7K40v9sahds4Z3js1mc0cSgpDR4Q98EoCWcnlb24uEbaSK0RI
/hF6/3aF6+zZoAZXuXLDgRhLrJF9Ar2GY1NJ/F18qXidD8MQXatYBqi8ZX17c+uMiCFzQx3a+OLM
RevEefKoLfL51eH3g201Aql+GI59/pA1i5MzjboVM9ozatAOERz/I2cB52NCXEcn3Lw66dQxUhfr
edFMrctmr2Qb5DH51ie+QhPoa2jfg/KKW6gH9PZu193dXooP6s6goLc27YjbRHzUN4WLoWOGGuMN
SGpSLxa7Bzyf7IwuJAx+1VuD54NtczxBKUWo4SXkxRTCFrybGyqkgj5iEJ4KSiranMCpuRjv7mwO
7pcMmlQqGMNLyuTg1aorIknyDVYhji5q9d0MXFnSN6AGzzU72Z9tTGwXx9v0vIwg0FXJMN6VLGac
tUOuW3NpAvqOQjtWVINYWVjZLczRTvfBvEITRkUtyTLhU7ITZ5d74zAaX23C6VEAT9T5e3+WvPYn
Pel0+5qH2/HuEA3CPlLjC5Ox/H2QRZ8vQiQ081E1WQhGyxMDg+zW/Qa2AqzYjps+4gbMtPtSE7cd
IPiivQALCwVwUo0edDBCAZKSaNmu5YlFRZ3pkogyWYI5QS6mZwSEVTo3CnlnjT01QXb9dClCLFos
nBGjRjnamU9RSmSFaDsCwYKkjS9F4lJq0NCfZmguKIlwUJlQ/Ysr997g8BnCwiKXhP8EuWgD/cw+
DIvfBXGsVvSTzJ4aAFtAM3Gu91YELpIHIG5xSTn1Q+6GtRbtDHyJKrWx5272/jjJ01uF+JKpUdN0
CJkIuo0L0105pHACDHx2+QX+qGXZp3quzRzChUZ39OdLVltWqw9HYCj5hwCbKtMwDGPqBPZuhhEr
vyW2A6Zv2dpIPnCsU2V5/o2bI/+4NR4J4fDki7eqo+/YLqHKYLeVHfk5+pSNRyMGh6DoQlJ0MDX2
hLzf5b80iaWZxB3k4mer0HsGx70KEOPvNfu07x1RMyvK2+HNwZ1C3olWLDYmAyaKEb5SJfTxXOwU
8TXuUwzUuTSh5IhFp130hCvD08ni9qj8Evy8hS0o4vjpo0ShbcTgbM4M9C/8z/sVwsBuy4Am05f2
pAXJRx+FqU9+QgGElMMxLHDeE1Kn4zhU7YxyNZJod/vE26ZkjiIBw7ZE+ujkk7yck1UkbO5EJ0Jd
xFckXUZk2/Y2dRbiz+xIOWM7zyE0UgvBkw1A4Mel5yRV52WB/av8wrHcvWy0fm3/kpkKXrAuaTZY
rQb5+IybROEGOWeaQELiPIjV+5+H/EUQkjz3eUmCuvHjs7FeMzywxJWQcEsdlpjbrfSifyGSDmVk
Ln3coESBpf1CQsFHCcBQ7yfv6IL4RT2E24knsY3U3IBkVAwx9G/L/RNwXWNy2mxaMy01mj/5wX7+
zDFIws3WylY/NNPMPvBnoWyeYkOYKLlycODMYUunUf2dkBO4iASLuv6ziNDjk3qW3oeHMYO9S0KM
bghxnS8LsXZYUV27AwoBMpMYKKJHqR0j8Cy6dUoR+9JHqmEAVX26kqVk1GUBiTf3RoNgCCmmZkHH
cF9Kmpn9G+MhjktMgxfcRgzTe3ywmPebPNt9UC0wSOsRL2FOpMhBE7ekO545GUueGYbR/X+dbC3D
aTYzldWyUfZoyWn3GUxdb9QdlMCbKvw5vBEW9fZlWU3jZdbYCHZ9HjjGdM/fAUAPaOHUMVOi5Rq7
lwcPPBAab+2PHO6WzlD4ken0/PUDTDL/AnmZ19W8ngB7VnB6fNDjyMyXmBhxAZZ3NmrxVyIKw19M
mXZ94Lxo7ooLHWzISNzd/SW0dK+fVxJl24LcKGY45CBO8Askla9sPvZy8mWdToWHFPL+mVLnK6bY
+i9mtcvEgk8xiPu2DdZtOfwxq0E1leBbs32ssufbkVTVnBxkQL5/S1at3/lVmCd7Q8C95S5+Hefe
N1llyDsw5vFOiILtrxlfAHtebOTV3NO0tnzwy5WX0XK+mWRgrrOo6BEFmrcyziXJvZtbg/GFKFHM
yfFiSGo50Te0jloOmyUwrdSPjuggucEDg3klMIUz5sHITgTWhYi5rVQkhfKhE7DUsgu1sZinTqey
1QZoFbErqW3zp44R9gw354wyCkNGgPyy6hpd46+tLLpiAK8WQKvxmMLpNoaJOcZrx0DIfR7a1/KZ
Sy8SCgv+w1ReCX9/bim02n+S0bAp1d5N8SSTbtM84CDm4KiG8Jh5iPqPE3Y0fR7wj6ffCSAyKl8A
+03LgVygqEZQh+59ITDb03AbW0yaLdOHpcxPM4sdIu7RPgVmCVQkV8AdajWSNlT4kq5PbBQ5JXxF
XqZy62aYClL4riouZuT6fvF352MW1s+fxXZtS5BHzYXYIrGimv9ZtRQKQqXI5gbQxv/BUzf1jxvl
w9GgaJX1fyz8mkQ+MXXGoqtvQb/VUYxINqaJIJKOg3RwCW7J5JflaAfFAfFTsbvzFVDIcAqFy4pJ
Qb62L6SGjTYRU5qaeW7N56AXrwvC5kGxZqEZyBCFDFAxRB0uoYh4IfCntikiugKaQ8maWrSaYk5E
raI98MmjjuZ6R4Oee4pTfqUM8/MQqAmaL4tAWkHjnnaT5W80z+XrOvjoP77BOD1P33W3CsaQp4d9
2GWIdDhlVgIGJ1c5Mm9+SdzN8XJatzYBaRex6lTSPIn3pVnotHEDPGbJZFG8KAgdgWTh7yc43UcM
23QnLI8Kx2OFEjECXPPiGpYcTi9d7O7Yn/DGufRPyA0FnjzdDjy1s+OW17hpD1RxuMtmu7YeKCmO
+uZnuuolTz7Ud4MKtIuIXASEhefzySPdANhI/0DnMLE3uzWSCP+1SCzBMmCVb6zUZS40FGzvToZD
01o6hktrQGEwry1m/dPjeLU2fg1Boe9v9CdSSAlDzDTFQTz+AGWXaDYMCTQbZcpWmnkCk5nOq+MG
67I84EvOs9lzaQ2OJSnP3DSo5QHvuLwsjWBB+OjFErOr58FlRyBhAG7PB4dI1jKdc0sBobsvpQuR
ftUTSsVmTD1G73ugH/70ExFr8SLbc+0QLcAviFg177vBR0rhK+iCgwY3plo4eupNl56d1+qNq2/l
GtiWnRB2XoHAKWcFgYmN/XZ6ezpH8bovxBkaKh6wb5DLV3nKR/Hxm4Pg31wywmdXFJulW0ATyLhP
sMRwVxssMqnFQuMvZG5fXllOnTWgtPYrpM0GQHHBrbLnV2DgMzXGK1r9W2sljazPDwuww+Fz8Hb8
NTbbUvH+qvQp1pkiUuV/qdAxF1IxFm8935XXHuRCuRNOOVPuwoRkzk6SsnJaycSquI3Tdy7RR7hm
RC+/8g6+GZ/HChdis8vdxecd4Kq4m+sC44uCpIZkcRlsLqpwvdpkZMpemHNhHUdOVdLKXbu0o623
u2Wa/2WatqHo6v5hP02u4a71hKOFDVVjllstLfibwJBssssxyqXnW/M5gpDw6SRSoFSW7neIkM9J
Vflgb8y/GDuu1vg48XrFujdexWqGrUvaxuEL0Uq6OCgutHDuvQ4f7rh4iJacyphRAzGyVvuDi1+G
aQ4l9f7ootvsOUt72B6xGeUWUtkp0pNUaSQTGu1oRTjvARky2eLaU0Wl+i2NbfWueOG/CNJTo35i
SNGPnJabkvxl3zQPetNRs5Uy4niwu3WDz0fo9544WCuNLMkOSIVlCJxwiKcKeQtDfEzJmWg1DqXP
2I9thyDVnnO6c+bkyGD6u7WTIvhBzat4ZSaDEScPd7NT7g6p6ZQlRhbD9DuUAAOktn4hvT2EN/Fm
sXaDgpTyCkffzdVzSLhl8ocIxHQqaZSEW2ORMTgs3SClF2o8P3iKCVDHQ9j/fS4nZZpClapz6hhT
u8ERT6zDshwhOm0jfExx37qIQEL9haB4g9m/943ila6ixP/nHdAVv1zrvl0gnMHLGGLN7Zn8o+Sc
ElGjY574HdVkDY/6be7qWKD+QVt7BKAkJtqabkU6OS8Q5ZbU3+ZWc8VQJQEHAZUTNma/Nfw/nIxd
Xkkcvkvbt7QI9t5TqCJQZ0nRzHKveAr3qrPsdfE4GQqDsQTitvAmYbVxaYuHhx6Am8pHDFxlvLgm
agc9QeBqbWWo/YJidZjRn5oseBrposF00uqPFU505r7gkUJzZ/OxGR9vhPElh/XXPDFxNk7wEuW/
l7blnwSCeIEVlQy/z84nx9eYDm9Y4XU7r5qU1VyrDAgqyWTHaWJNan5O9dGNEsbrihhPPdKc9sR6
Inp/e11B3Bsqqwil5qVHMs+01nd2/YqEg9gGTdKWbWTODHpxhLpApv9FyZzt1XCi9WucEkObDeAk
kubx0JJyMClKHIJXZE6VHaPqHCBU45b9Rc2cMyXT3rvXW5QcXmuljv+4TLZE3tr2sF8ypEKl17ZM
36fMZ7/ihygsGOnsYQR3se84vy4Q65i1Z8oLuVdHZzy6WsW7UOQ/DQBO5zt+BORjPiUDdSbMPg02
+rQGTriLAsi5iRgar+8ZTd0r0baUQPJYdznRyO3QZ3DFIkmE00vnqD5ID+R9TKoHgmkS8jqf4Ev2
fBOYpjz3kbrtS52VbJfbM6zzteerqofE1/5NhtbAQ5FkBtmF4jue6SU1r5WI5kVAFwniItnT4yRp
fMozSSqcM4ufF/LVUhewW2MQlTdzsOgPJUVH/mPrcgtaith64K3fSPm1WotyeyqS7sWMq4erllB5
FHmyv7BHEEj3EISATcoIKSRcVtKHoPFlxIN95Pvd+sL7pyneW0RE+0gCaZVramzcm3NarExyow3F
pCDV2sW7K1t7qAhJYmdo/BYygeqJuaZFmujOgUVPLwVd1RN4Lk4RgqToLluZ4JjuZtwEwe+IqNz6
R14K+O+SN2KBBytaY6exvvASrbQ4sciNEKT72NBFMplVxWqpFQLSFZ2FDliF6Ith9kilXyz6U88M
3VTJZ4wIgOEKgVa0vm3VLXWcovttaWqCjeuTh6u8vRXYMAvQQRBnYW14iRIua+BZ1GWYN7Gs2Zht
hvesVvrrVrE+3LC53vm1VGLkXgPs2WG4Yv7Gnd01RNJCf80ZXFJb7wzZisbSihijUUpx6m7IeW0Y
Ph+2OeXb6ysLjsuLgUgpijzWiPdM1rXEOkE/ia3nxAKqGUESC0ptrWLC0kmA2/x1tFPd3BXhsey8
nkxvm2HWpIr5T+hgSHirAqqG6kSEoTjv02/eCV3pl3suxH1emvVWuJycdI/gsgKws/epUc9Zp6EF
xPoUq4eAAOtF5Y1GXXFEE8S8Ul5hi5uGd3sLt2ZtvmzVUd7YflvrPDNMBQERapr2aisvnFwbEHOO
xmwuM8k9TAg8AgFF4s5u2dTpyI5VVqACnnRj8AAxkrE4nRvzOw4BP0gEcsY3v2xef6YtTa4pjWgu
bzFEHORJl5AO4SFQQ/LJMIEH6FbfEvNytz8RYPAuK92NQ16zPkaUP8ZvFLDodO8XmCxSRNJCHlNZ
icIR62CHi9jsAv8umVrh9h6/r+txPjzvmT3/Ny+aUw0nIaNGFzAtBKkhQlWkndHNQVruK3cH5Y0F
B9Qpm6s9FhSuQN/HiTJpc+8zCWG6m0pKp6zOhYc9EwW46PzFw27Locto2CiXO0nkaOqmF5naQYX/
42cdMshWJ1l12NQPgoxyfCPOzEYpBTYaC2o6vSBVvPFgDM2WyTshOONwEnzMMFvPBColy/E34pfw
W449vWOXlqgMz+DBgxtzAZWPd+h7vxujREclv2N7Uq3VrG40np0gTltvVQJbhPLsoKaE2BJAqM0A
tuKGIw2a+OQcqyeCGnaxCYKbgWkCkH81DucsUO+qEiYOo3ZbfZ0gdvHxt2pz6Ux2FcokI+58la6x
nWfKP+n1hYbpr6JJtfxnLS+d1cXv+HnsPlw1n3thxEOjZqGTi9fW60uJXZPMC2HzcqD5pG7CF79o
NVKVY/JRKA77leQHZKVpHDyM7/q+VVX2GibzYtyi61P/ggrws+e9UWJUE9P0ey7qKuXPDgRDGSsv
dThOHqluTZuQ7lBjAq4xBdhGc7exNtHWDqaVrO2KXsQXK0jHgjU5KmNSw+LySqQuVgh/SKqGmCth
xtZuEPAqxHxFNjmi6ti0p3H/uzPbpHoZPpp5ZRByOCigbtjHip1m0Eo1YgABFG7Z21588UAKoQ5m
MdI7514mBP9KEVb5AMFYdXcc84Q7xLxXqJY1rhOPEHsLe31h09w/2giJOAwu0KzDP+5utGlhjLz4
7Pteiseo04rBAQSaBH7sp71DSgGnYWtdOC43QwnbXDWOS/9mqPBK8YWFVi70KLaGsrJ7xCGcbrnC
/fyDNLFfqgt2r2LJZu0oE0qnJtUsgp81IyPwyYdsZHV4ymkUfTyF5nGOQc+y6KEkNc6VLpwFoYJK
rOhTzaZnOMfnm8NX9Hgg5O8/PUWrQ7TOVom7BdTg7vJeCFgqSIjqs9EXF3NYkA/u1/qKvmUbQm74
bGK6pzjYQP+GPEBz3JB1PjlA2cNIzMCRkB4Cr9o+EeZHPMsa4aoof2US6FYTR8h4+KHxtYYZe0YI
AawFY/X+u+EUfakvNJw5qgVRZQtr75IoUyNVZ+C1E5sBHJZQR70nHaecA+Jt49QAc/paMVERZt3y
00NmJKTd2DNYttD1n/TeAF0iVDdVBGixqv1co/eebYmHdD/Il8YllDlD0rQGtLxDpzFHQbUxtEJ2
gnrSwBSxRnoffzPNdjiNAgjf4lzFVgEy3lGAA0fWS/4p6rABoTahmcHmaGTGwtj3FcD0RbSretnJ
bQF+yGt2Y/iVagQ6WgGfPvdv/XMvEeJ8VpSHyjN+LnfIfkUhgqmu50AEhR4rEI6GpT5eMK+oFc2C
l4XPaZZANTe492peh/S2Yim5/kFWXjp8jKYzk6HZTLrD6ikP71UbhmUf+ORid2MOZQ8JS6yKqLYF
rC8Evi9ICv4URn/kG5GElyCGftkuD3yZF3iSLh2ocCskXTwBovVNuq3zh77GnWYJDil+AjvrytTw
RAMKzR+7cYtkJ58gm2miLzmFWtumlzcCRLno4jeCw98baTf84E7vsVCdcZlR+Uts1uUZFY5pX2m+
R1SeaaFdhjTIP3p3n43sMobATfp4a6vv9XR8wde8bPPBumZoDsy81yIMkInvUGSxjVrOGR5pTKCS
pDpjSwRXtWeNuMkSPU46PTmnpACpSEgAB4Irq+DhAdem2iWfPG8q9VSWKiPjdIgKBUV1LDxS33kf
GsIxPXmjCqNAY8GByR1k25ncjh5D4ui7lkjI99HGazlMZWJzM5fkdcuxF6kigeC2SQrARP1jLREr
MyRCX5flR96Mezrt4heJh5c5K1f6/2MpJEFRddA9MpkcJm+2B7Jugk3C3l9KDA3bFffB1q1m1Mrz
yINGECpIA83uWS/VNaXLwpP7ORrsgNOLmx5KqYhhCSeF95zB9jWje3zP5sAeMkJpQOPVwymIsf5n
h5ZtN8wOj4IRIkz3obMPWiR2ADvkMf8kqsNF/fLb0evAH8w/cyQjuNVuVYZ7RnVYdZdvn62qaJiR
FyBKllHTuyCk5Gff+wW4N/9lrwGTW04ot2H7J3llMgosdMmHbkrZ+wVZAFfEceHYqUAGWqqzOJ1j
T+hqnuKexIFfEw5APuD0sirA3g9nj2ZfqFCrGNhzXrfW/2UVJopTbN6rp4rmFpfTkJJFfuDmsLeU
FcDBp2fpIZhQtiosMgSzlnJwD8B1kY3n5eiNKVHI+fIa7M5QoyfTBKrBm3MFqwKHlnLuNbxXNGcu
JrVGR0f/olh9iDSntY1ktUIu9yPC80jzH30fYxU4FXgSF0EVJ3YHohpiOZRl6vw23UmIHjHMge7S
JnXJgUPI7b0J+l7HEdNv5ByFPRcwiKE1XYszxGvcQ3DFv3YqleCFLnqmHPVON3Vr+8Pbw8EU4IWq
W52XBhCr3KKawWdeK80e32tPrEz1Luriwv3cWNIHtwwLBUrek7kjqvArDbMRG1tZ/CW7Ej49Kot9
s8zD0X63EYL5yC2N3mWOd7q1Md71kBV77C0NgQZnhCyMMqJuMVTpY2uqAl/uyA3mqQMuKRkjPpDx
CSWr36KZfUpr8+uF77fK/LrjDv1GWb2IHvHhusk6uFJlavzgcuRpa1jspMcWNi7t/OqqnDCmH2v9
iVelonEDNO7Ue0tRTVS7Ps30DXVgoJ5Yq8da7O4IckdnHlT7r2t3XjKKM4Hd6Fc5PDqscSWOoSW/
QYPEjfODt/hWqEVujfQio5Bt2RvNkeEDec5rUGsfb8Ap/O8sZzLpyy5KctO24mCm1+KBsKoC7ZY2
awJvJ2Fs3l+EFd3wFAt0K0GK9YKSAYr8GMzEdaUGHp2TkCkjpNR9IsJUZkxa07XkRNnwVFikgv41
+oF0x9DdhsON/kXiamo0inBE/WMxbxWV5jSxo5RX5bgRFfqJ43fQ52iz/I40YItHudrk2ofPJg1c
Cj2i+0DrhGEyzY1kLEh+NMHRysfKgG0DFV6DPdbMqOCwXqu745C+lfhEtoxkGwtG2j9/Px6CxYeW
kZaJkDG8u5Z8snruE/d07sh3SuOY0ikJwmxKtBgnEgzM2zMeEC7oO2TSi+gjne/f4C0HxYwJrvgA
/8UZwsK12y7moAgh8MJbomeUhkqWBdfgjP+MwD+AigU0TCYv4/As7jq73nM8MxC8B+Mr02dmUwK6
zeuTjL+s07SIZOls/Dov6FsEA40U0iLAjhDFWOzYinBy/YHT9RAl+6wvdVT8rNqKeNCYWchtqFyC
MaDvR3WrfbHIdrFHOUf7WGvlb1pNkc4fAHz9ng9XVs+YqWa+WJMJysaO7eZoJwsFnlNxml9wM+yY
YEFC7kYmViy/QfcOVVxf+hSA0ZPyuXXtxc0933zSxBEH7Qvz5AHhfnSx42gd/PYSHEAbiYQkpyFB
JYGhrLgvrplP4CvwarBNfjvXQkhiSvg/63ficqh3uxEI1vL3xtkKGYMgQGKyqTaJkkGi3JxlYWC+
kyQ4I0rjmnuUQMOcZPtPU0Oi2C5mjUQbon8waZL4T2H+lEftZh5l69SAfn7gdK9gfm+XjtGQiUOd
J2RMRTD2acBZvLXFHskQHkFjTYoQBeqrkU+RnIDxOYOG4bn03/AhmsAgZvEtT0iKk8HhbBypB1Yo
EhkZBEoFlSZwN74fQOyUYs6BCOgsT683MoilXmzmNpDhLpZCcfSSVgOPQXBYzYPxG9zxl3sV4v+0
aieu+4OB3XmFEwDvPg1KVBXo+uht4j3w9i99zwbJlqrahaTXQBGR+3VPRW4ZzgkmptI9dfZLoxRd
BtxYObbTb04/2y+bzyaW58vlmYrvL4uEO2hGNyvaJAtMoOKCuTLvbbrQKW57nA6RA+Xl4bGZE1iR
+kbo3hpoxTg2+EBaGdi/X27EPiFk62ElIE0MDsiMOeMpsVeA/LAgYBaUVPnu0059hxyC8Uu/xDzb
t4AkWmnThTu5VL1yNYPbCjNNN9+iv9iIUr3nBgPDnse/BvqvGf6/SK1/qfXtq+xOJKyNmqAplrGW
JwSeZ6emJ8fIA1pIWIsMltO9xFaRZkEBXKFcSAkRORMYIvUIxc/OFgffab7Alk1WQhXhmxiw90li
4woLbcvsT+O42B2jEE5Bg4Hpuoh+GZOC8rgC8zn/fwfnH4B0KRTyyo/V6QaaVbw5pJB5SNh5pOWN
daFhO5Q7OsgFa0eYxb98zw+t9TLoOpue9qtOcyOuPhYTZpqiyg8tAzb4hSF8yLEwDHiJQUDFHmlg
4m5hvQNgRkyoKFvLA9Yc7919FSCh1yI6ys7/HcN76uSpAr3kzx7O17n8baOIvrpKtaOFXQ+y8Euo
k1taNWwGujee9ghXOUPaov/zfFQ7WY4wr0chG2J00a52RnU2tl9bUuItensRVft7hRsxwAm4CJKK
7F7n6YAWMUXYezXJBsNH2eF3EDzIvr162Qfn8LbQJq9uBs0/yGf682kNB7bU6gtZ+RyJPGZq16yT
onFFixN+8N7IuOpxg4y9iU6JAV0hlxgbZWohTroGAmOXM2uTms9kGHK8Hjh13Bw9Yxu8SA1IV5Ew
sUSC7DO7Q08Kh30z0j0YobUTNh6Qm6Pn217Dzdu+dizzGkKtn82Wd8Ms7N1f626ZV9sdTJCPBjVa
6mFHGcWqPK+k829IvZyOK1uSUlnpZbSvj7nffNVBm/jNO3MEFzuXmcPLYVMgwwV+g7d3BZj/CjdK
rF5t8cH3XMCoVjljIliW/WqVFHS2YDAslEmcdPCdztoBS6YuXcb/7jcfYSZJ4HwJVpKUeZFVEIFV
y5TdVMY0CUwGkaKNDgkqxV0LfxXeAR2qujM6vJ7ztBNc24NLpS12d64NHReMCxgCws8gpJUhc+Wa
gOJ/vZtPq2RuZ7PPxISSRTAt7iGCtLZgiNXcxNWM4CtR+edEqsQLD+56xTM+CvbrVX9r1LXfLRcz
zSxIQvlPQGCgv3bg20NeKmO0ExmeRKa6ui/TOeQ/8xzsEYudQiWHY7Q6xoTZ0Ud3JwUYEBSiqCHX
bjY1Rw6Ns3GUKXtf4GX3vFrz7MajVUSN5ulk1iqB3LIArVAqOKDFe0AfUVRctxPDfBwS7LB6XV4G
spGBJNv1TYQX9jCifTbmKY5syQUuc9kYfbv3byYAwgH684HdgYKbRV/KSGWHWPNbdj5EEZ+NPfyA
p6BZJd8JCQa2hILB6j9F0z/LaRTr983LydUWIH0ps83c7sWOhTjsJrRlrS9NnSBRoo2rNJKEyNWV
PuuZRfxvTAF9JUQQbgHDILW0xW/H3c8jGx7TUxT+xpGVl8iXlF0MtI9H+70Wdn7QoE2xCO4qQyEX
Ut+oP86AdrAX4cOV7zmiqXs5gcy5QjzCPbN9JOzo0BeGXiTOfaiwKRtPfwCb0XvH53O0jskpboOO
+4L6Hk8lJ+R9CyVP50lkBjaDritV52+/1P6ZhcCjoHvLXVH4j1+11z5mZ+PaLDzOkvFemb1pfMit
ilypMr7p6JNiU7P6Cy1UuBUiG4reoIHPWqlT/8tU9iefz33eK8ZIXhc+vtFL851VBiKkKmVakKTP
F+C6zbEF1N1amUwPQUrd0XjeYUj8IkbczalpVq4T0Bz/6en1N/B0ihDX+2znHIz5wBkR9nZ/Se6X
FKmnPIHFFDf9sV1yEO5eYIxts8w5wKBL3pPavZwjPtQ6HG8XejnVgGMfSaUZL4gibFB5XR8+h7oT
EH1YiQCyEq8zgmP6ymKkQiOHoDZUBPhjAZdSSZJzyxUgzODJrD4REAvCMHn1V/a6Df2ui3hTbmGr
SCkrzyLlaEAYHDSD7R9EJuyQ2hGS6JjqsK9VjXIvp9ahr+lp/t6Xvf/x9KLhd/8+XpoU3o0JdTVQ
wcV8cKneHdJL2km3Fs0nrz/J+q1qPtog70EsIANaTsJIQEqOTnc2n4A31dblLjgG4+CqevNpCnjd
bZl65RHGMfkJf5fZ4QHS/VbB2TPPP4tiN9olruwULTv79JgrrLpRD8d2bUI3eNunkoyfIY8tMfyP
2Y6ruA9hn9Wkk3vx+YscV0Al4Mb7TFZ5IDdAMzWyQLoJpg9GYV5ZF84OFy0BcWMA6GDHpY8bEgQW
jes+W7/lSPQf0KaSo/s1PXnDypVkoHNSS7ulM06jdIMBIcNMiOJ6ePofD/Blmv8VRp/vqGYq0Wbl
YgD7np3tfqCSTQAQ7rN3AMK5EAkC2BTIkObymokE0+MBIR1vp+hIBzhFcXPTpCZecbr0ighmORM8
+pBT2Yhxuz0iK+duDlmpuwOo9D0vdeRCXPLuWeOMZpnMwy9FBN9hjB0QzI+6nrD4sq6VG+tSKLDN
zqn/XGtf+uuoBUNbxC8cTO3zdu3npMZB3F7u2bQtCztEDUXlhgCB1xpjHEKNOzJOtrlOk3uXIYtw
HCk9kmOF6oT9kHyBK51tW3iGH0MQ24j/1P3r1YJaRiq6Hf+yjCwg+u8VohL6MAT0rQPj7MK9fkkK
6jjJPUlLfiTj3L01AZAld/Rdu6EddimxCe6ZhngUDXF0ES7HrZWdl/GkBDmBCd6BVpmlscd9lbpy
TuP+oZdFMafUoC+Q1ccX0Vjtka8P2LjCKB8CmfBMdc6YdRvZH7aRLNjmCcFJfb8frM68NoDO/9v6
VxQpuqPO9WpKR5TE/5BaSck86elGrZ7K4yC8SWH+4AU7XTNKJdvg8dzhCHrd3gkKP0Q2Hf8IELu6
YIkG1lLdHwb6kzP+qvhJbKGSjkg0Vw0u/IOoCmJI1djL00Lf64NZqDhvyYFotkHkg3SM5AE+bVvd
CFJBI2iKZDj8jGo1f/U9r20zLy2gFfeGeDCs/Ft2xyb+QISg0t9MWrGuDwTvzQq+TEUcbhh1CdCv
gJPJg5zzdsoMdf1f/UZIBDAF+AxA20OskE+H9RncJMgZoxvaH5SX4kr/e029Xryu2WmmrCuWWi4N
HsBlKjHKsucjZqel4H6oXicocj2TgKwHQaedKkQdM5P1NonmLXburzrte7MUGXJSy7Tx1olK5wOh
S0rC/aYtqHwtt6XJOcCNj2FC1sl4YJwOarOzi7/sCZ5q/XStcmmufiCCHPGia4Gsl1p0eAHMfzu1
LanWSYV+z6uVzD+SkR1ZCq033pjNpDKYFdXxvXuIbbKPU/0umohbcgdCtpklQcBalqgh1+4grSrN
+4YR1Uj4K6io5a3I+UbL6NCUcOJWFid3vEBYVEEIs5+07RKAQXBo54qBkxonqING4lz1TuWq0TuY
aFx6gN7PslEbhE88xrTGlVW0ctK47WrbSpq/Vn23UchMZQWSl+1AbCFj4khuZCCRj5+Gc4sreBZx
tG81FEXelGJvFWcspiFJ6Y2kI/dgO3SLdMh/37G8J5hI+Bs5XTcCiOPl8Ywab/AO/GkCIepKvVwg
V/05H6YQelY+8tWB3lO43PUmGkgkZBimrMNVa5RCZK/wt1facCqiDpprHNg1QBXVh2GUZ6KFsfdS
0y2Z8npWg/3vCoV/qXhKOq+n4XU3w9K1yM6e7/NlqHt5T7Qo0+NbNJJ4d8D1i7LKo8Ntxlgo5rek
kNpIYrXk91AGelZK1uTUvRW36IanCpWfkmJNVYkOu2VILyT1ZyOfNm7pMdYG+UCKjOdpNisYyVT3
FFlzqj9J0G2C7bA6Y1p8u1zDlEcFLW/MbpflTIU5ZVmNJjvlK8/tOwaqM7Wo4la8Vkl8db9NiJ7w
NqnlXzdBwFvT81zkc3jFzn2DimbNTji2U8lwtaPSwpoXwEeAOIbTTfNdHAq8iMf8f8384LvbRjE3
Z0r9IfLbL6kriB5QGL1UzeIovZTPNsE5j+KiYnQPuXrdjBYG4oYUsaKRtDLExNykBpAClp4CY23b
U89jfeTltcN/LWJzOxpaI4SQrFW9Pliz3rbnfixmf8jC0TbGqhQCFcUPCqSiaO1r/lFI3wRbpLU6
c6mKCnUwjkQeApthl9TOn7JTuczHe9fWMl1tl17XYswDmAqBq0EgDSOFlbN4PfkG31SIYLZl7Yya
wWWcg7xg0+ImcMWmcQqD4ajAZK7xJNx7hIWATDvne2PbCRLIfC1NpiGW73rUJ2dCJ0nB0P9smmI1
UVPmenLyub/Y26ho14qBdOeCLagIKO3tImFbBSNsIxGqBm1dApoSUVv9Ol8XKMM6JSq/PjTgbuEt
iJB8rf0hD3nkP6DVdm+pR5yoFguVx7dywv2biIfqmmNFhqhQ1cnOmdkmZ/y4XI84YW4VWMIX6An+
hvBcXdGss5ueRFj3b2mpt/46IaSyJs/Fn8T7H7OQLJgqIsz8RsATiCGpRGUhJ8JlYD/EtK2u/9yU
GerNFYcjRB0QGdo/wsEaqc0Yo5CVBkBeDf1HAcrL+BbDytCjzkrgixjVAdSBmp57Kca4yir287JZ
xHfoxEfbA66rir4u/TNDzQ0Yx6NJnoUKv1EkfZpI+hMmf+ZBCctYxQ451UEEpw2gzxPIKwfFvfZJ
BxhaERR7whmSrFLTM9SKMlRVsAJdn0OBk+Uzw751PB0biT+BskbUyl73HAxbiZLGxm1pLqc2vfCd
DjkXc/r3oPv6UsPtSS0I+QSuShpG9sqpiI+WhUo6/jELuNz1lxoJ2UFPVQ/ooJlTpg/P1Dvl+YZv
5rUX8ODYGDnDvBYS7ubilpJSKbsHnClC3uoeYy1NVJHpafYuqybxhirUh5CBp7MnrPpxhqTsELhs
613tyFg/y+Mmb/AQpL9yO6NWVne4uur8J3PY/XQaW0X2I7M4Y30YopfyWaZf3FVElbxUFDHCnGbY
4+9Bo3JFzPUpFzJW66E04yemTqeWwXqFtsU5JMErYaHE8vfdxm4OD0czuMjhHgsKJZc/8VU4kl8t
PAKbAHuPNRL51W8lKfQn3z9LSYCXhjKDkBqKijqoizuUsqxpEAjhjEbTHmnJHBPDtZlEZp1j3oHR
kTJKTZag8VPJpKbCjbTra02LFbckUQiY+DpETz5sAsTLNlTCrxn6yc0zFAqLRokLF3vdr0zgTQdd
dKZHG9NEKaWOcvSFlJIdjRQvKAinmTWBV26YeowMbq8JkgEabTmWdSPFe59R0lZAGJe+vIpy5/yq
g+n5eRXkD19XZsStE3aLqoQ1yGCDwNW4OHP03nmXFEp8YuszIU76B+vg0wJQXBjV8ntrK9gOoqzR
zV72/IxYfKDXmd8JgdyopSXflMHwz64Zk1L9pU5blkYWyb2ufwuN66jL6urODE/luBSVMRbTfnhV
5GzTtBpJwmcSrZJzsSDUexzOJ0Yo4My5V2TxHOoLuA11ZjSn0dQCLBdrJdc5FQEd1zPdbpVs3Csl
84aI2Cu+0RaaCEYuPe5fB/HFtSBx7wsCwjoVAzxd9/kLK4YJP65ZwCb/DiNTy0ygzwz6aOjyMPfz
inAFVoc5P/B8y3Y8spUANZkHhxbdumU1ncJC6mOY6CCFKL3u20LnuocyMwgHX+YQ3L/Kh2QCeWal
qqPLiUQ4hucjmJkzQOlSqkyVg+I4i4/xDT2pBH7zuTuCgbDq3rMteEFsDozCgr3JkdRgo8ROfRoz
db31+E/QH87mSwbHhl74QRZI5q90KHyU62qswrRvkMEE+8ZtKeKGs2tKGCCDd/vIWH2YnEVbTfbs
IpIwenMqh6NZYwVAsqFQkZq1/SYY8uhstC8tWwgek9bFQrtZuE4XwZ8rXGhk3387EHmUWHFltMCO
KFnpyY30GzHnjcC+0I3d6+Y1sGuLSTCD6wJqi/TYSVj5vnq+iT7n8yhNf51LIobJLcVjWhUPumGm
zvFD1nT8Fpqjm8NL45MWk+R5Hn13fNEcEVN+8Mxp2SV0OcWyGGymPTiSLOFEfg4i86hUfkdP7/9I
BInit2sofpqp1LxaBWDhS/1nYcY72C+XiUFp0D4dqt2YFbc1Aif5/zicaSIjONWS/L26mxgOgjTs
EWMZpIKuhgQ5Cwg+NSy5CJ2e8fEedQ+TX/m9VXvFqRgDIjBI2vPToUqSir4X6ratOwaLcopcJHDm
p35vb08Wrg12OwHczWwYqWvUzppLMfys++l7NIn9SRIGSQ3txc728oZ1H6NnTdBWX71HLcVVbjEq
OxS9spUYxE2KILAGXGZaKF75iEUQl1KVi07kAMt5F3By6wN2xRrIvFytPtDstV8Lo/B9ZFMIEZw6
mTy6AMuNxR3rQCxFkjK438gqsA6El8eKSiAcp+18I4JLsx2K0kzYoE1pRTcTEh1u4zxKYjEm7k3d
iHJZ5NLE/h63pQKRGPu870qmxj1d9gk9j/PT9aRwbchX7sRksqzW/R3eVQbwggOeeKSjGrkz67iL
+KuzgZ2VetGTftAXUdCyX4vl0fOq5CEIREm2Gi1/2Ka/PCkZRlFlDgP+dit2VaJ/E2GGSYiC0zo+
meFM0wvB1B1UCNKqQvq/Mjhg/DepEYuGZlIkzI1jtMvUnYOJx1VUHH2GKnxpnF88rIKLrLvLtLZr
9eEoD+SiGImTDEs4QXeuV4sXXVjyOySdbBK4zz9L/UWQqB1ODd/PIIfr7S2bfns0RMLSuuyX44PP
zGHxiCQ58ekMKv8Nu8VoSGj02XfhnhQstaI4T44JSpLvgZBZ4+ag1meNWPaE6xsnh9LkUTcNU+vb
w8S1Ra4pQgjYe6o34EgY70C9wNu2UhamiAc3MSsyrDzQaJCjx3Zh8M/evu8b4txjj1vkEGTR8NYb
hHxgB28gA6myhy4pasDmO6U/kfIeuYvKfmevDdT1nWo+agkvbiQS0h51PCMMgVSE6dv8YT1oVKDf
yK9iNJDrrnkQpZsMGClJNoSTEkMtJhHAkyQ8XheMATrWUYqcgflKLT1U9X9s1mp3DVU00RtEVC7R
ulldBwk7O6YVgxXCFdE7i26rRYoAI5Qs/fxs4O2J8fys542i4pUgvNcQSGvHdvV6g+tQcWJEyglr
zyjx2BDsN3qTv7KVP2hvzflmu2zLLQfdUuTJXlw8g4YDNQkgwXosXJPTIpJ+R7vv6xd1LGn5PcS8
Ww5ljm1ROCyQxzWV82E8kn2PSH+y/ZaWKMSZL5Eor+fklzn/223Ua9P1b9LmoflNF5EsOYj4yPDa
LTwK4jD6GckNBskQ/6TxXpwKBFUKIOhXWxvxf9yny37BwLKIId8qN9sxoE8n44F+dCO10ET6mXcf
6bpCuHsDeHKVw0fxDUs7O1r484JpIB6x0k+STtBnWqioq9RUwhv+I/7MtEJUqJq/sUYGjshSS1kF
IuFkOVHp4Bo6Cb8s6v7EqN3DL6EdD/cCDTsj+v66l3IGxEwLRu4GXEOG1CCa0ETPD2kwl0gIFfom
DZ3Atwf2xqFJ25+HNd0cUus8x2vfdVi1ctbckwUUOoU/vlc+KfwEyUbYL+oRpKDTcN9uZ15IF+mj
Hvi440hcHYs97ibvjH8LruRXehFq2nF7zoNBZP6nLlWONz+d0VxdU5SlIE/D6UHOXgEwJGfHPudj
e5dEdsTHvWjDzON/Zkc1fLcs0NpoQB/VaK1E1rOYorRpr5FsXN0xyzUj5Y464ARqVXwollYnfT1h
J5afFD6NgQ5Bi5TZeAMq4ccFwbHOB4tDbBtREH6bFRb/k1Wc7Bbri8ofLWg3NPzayHZdvNc9NBz3
6ar2f/4qVxo38U+9hl/tB9PsXOLR2CxntnJQ/wU0fhslsCDFBIIMAcHF2mDXqLaXTHKO1RLJgxY7
qRMUtSa9M8Gl1+sm3ESYoB4KsdCSUdhLi7wqfjVYqjK/va79bWupdJHW18s1kRNKP6teH6QI91Fi
cKqOJXdU3Uvknw5ZKZY8rIwl/0Hbo1n/L8CeTI9bQdAzN+cE4iQFbFfMJrUd0bnj1MH7dYHJhDnf
Eu/DDOrEINppYA7v8HaFxOqrAkRC/USn99kneP4sYKxAEWy7e527OGIKuPFnWjOuR3xtXNiacgIy
2qefMRcojjHbRzqX3Uj/u4oHLfZGWGeO3LynM3320SzSl8WyPXmBdkHRt+DF2ql0sghuf79HTD2W
X4Q6gsXaaNXIaiN5Ueyg5GarwI+PAj/O29aFnaTeDQcj39tPafpIfhuZ3eXbrqpO4NXzeDEjYMk5
g4RSoosA1NKDx5MBgW3ETwOfK5Vh3G77WaVgbiVOAkGJMlVonwkIXQoPgx0ljGTz901pOiiS7VO1
dkxl+26zJ0mvwZ1Mx9w+JOLFXU4xWw1EXy3hwFAOSLTqUz82qBdTIm2CUrqFf2GeKzlqWS2mEKNj
xJjXxj1n4cPH3yGQgLiIH2xvgonrevrESUkib9FOPa0m5yq37opESYWUelwnejP9gjCajVOEf30H
wSXR3hX6cPQP7fO2amWbWNUSLLNgRqrQOAsADHE+KDxZp0XSY5y+aU0ciJIN8z5G7sJub1QuCAcO
ZrGmRolYn9geZR+ymwXy9ZKyucYukUKbAUJ82kuWdkWF6zdSUC6dW6kYkCqeru+DBJDa/0kISGGS
ojn1/0oLXPUTQPVM59iEQnQLFcnUdKy5dcovM1fzQ+PLJ5IAuYFEz1JOkDs5gTr370AykVOPJdt0
UT4EM27OdEavapmy4c/uOUA752ccMSaJbf06RxEqru0N0wVK0eRfeImOpLgiRqVpdQlUv5Tc6IKo
pyrSKcgfvP8T73CM4TvIDP7WTQZAgaH6GAZXfPXkt4z+lK3xg3cgfGNOpiYADxLSuB9HeP/809HT
BnMCIrgH8gCaKAE51pgJR6WFgLd7zTervJEd7XVBSypPI6Dud2SSFBzCwZj7DOieLeMk3S4iiate
RjG08qDnWK/gw9qERsP8oaSglqezX3rvCbRkUsuZrg0opjvhBJNie9FarTqueWRM4ujoGMGB70PM
l6mmzmqPadzEn2TgtJSk1FqBhDzcfW4cv5/t2qBJheIEas3N36BgEG7n2dBurD2UqRiKaziRMCYM
vJxkYG5dr9HYJeLTbjR/Q+QoPgUk6dqBN364OvYvCUp5RnK8SMUszrRHCEegW/0OUZ1jr0WEwTvq
e3WqHjTK9GH9Oc0NECu6E4EgWZv7ksAytTfXdAckSyANeDYk8uzw/ebZTdc/r6fE5c34q3V7LRee
8SOJEIcg56gZJQ/4T0Ylvh32t4zFBWn1Tfv/OdC68AQ2ssWOG5Wp6iVoaDdGO5NLshWNSemQft41
9JjhdgXJ/lvMoL3jhyEUuCZxxubWqc3FGsJQZEoDYxNPMArd0c8WfiJ2gvX+0T3NDmwpIW4EXT2S
Urh/ypbVmfVUqOdtD7ySb5SWZm7Dao2+RNaJM9m0LNMGJTb/ei3mBXyxrOEWwoQPA4pFX9t9MX82
jiseHC+JEMrCnDCvX25c+IZ0l0fBxlYSudoXf7dT6W/rmcWayTL52wHVGsEqC5C12WdcxTc8JU36
7+vRIKUeq/qbd3dpLEqVhZ1TpXcuGOyqKEmGd9a1sJozY/RZIZ7+vesLXlfjYW4Cx1HUn/Yr3N4s
G1MuCJEqLXJIoEXYeuM5zhIR/ONurWbwZcvd+qD0ciRKA/Ntox4rkd7zkLE7wGfB7XhXqpyyKAhi
MHJj8j8pV6puLXjpWgN0z31t7aMCjUFWuLkXoidPnnaqmB2PfWnSsfCIRwZBgdabY9qbdEkZRQYV
8Ntdy9IkYWZT2rVA/Al+UHLNTP9mZRMWKduqGxewccKoqEMYgGxxL0Qw5xi85bbV9xdpiJVtOeS3
lfYKAnaxPWFVqOGWl3KIiaFwqQZR9EVHAULRy8jGC8JrWMt0c5JgBL4kIC/Fq/dtCItMn2UceKgT
uVdm8buWoanOIl9jB1NZXNoQOaNnzb65VxYI04SKkzvHH15JmZKw0kf1ViPjah5pCwNM4T//dbyh
tgH06bxuxGfXNQ2eULOOvI5orqp0FuqYjmc70mzXeVqv9d2Rt5BEUuUqJYfHm56U2C+G7iiV2bH3
tFpI44rglRq0INU+pDz9Y9p+eTsqqepNIxxa786zOLLSPzYxDf/feA3AK+TbTuwovZWWI9JkNOug
3TjrgadxKWVWDXwNrz26Lxend9gTOnL63SjaCe5c3Vi4MCYnWrVFrdpY7LzWLrc9n2n3zeSXTLGp
crjanwHGzO2uIylcSO55WPG73nSGEHQV0F/qUslGdfovpoGQKtu29s/70GOILTLgFAZbDsAHeAEw
GiGqtL+1Y9VOsIlIp+0AaC1qxQtwS4cOexCYVDAqa8GCNNaWGsog6sxZJqpPLOWwE/3/6f6q3ZxT
o+w5DVXCNKmXRP8eqTV1GojsQ2AS+Ptq6t82gXPxTVbs+VYVNejvVtZ5vv+K315ZpQI09AS4ek/r
1UfeKpvXNcDGGQMpAbSKQ/sOkUjjyVvZm1JsU/gyuRJqRRi8ATt3BZjnxlK4In4oqzUL0NgCrTJL
3F8JidIN2b3CJ8ZTR6V5GC+kkXUjeYPB0Kja8te32KtBGbwlrpgihcxdcp9dvL9j1vMPawujbV+U
Yvc/LnZScTWx6pNwvDcofH/T/QxVhHE/P5qMoOYHTpVOom4B5I23PpxuzO+SK7TwltVvQFz+S9kt
myY1NvpJ9A/4gTQ5UnYHR964GRTkZCm6gziPuRLX4Sv5En6jiifVqJ7rNhWpOGOdhLx7m9o1nGYM
Hk+SrEUO4ZBbrMJsvQzLQJpFIlYMVl0V5wUDtnG09BOGhstxLQCueR2qML2fBF7i9TnlJwrksa/J
BFVV8YycTAjMDhnthf4GnSoJxm7RSvyq78Q2AaWbecBxSurPtJNhFo394agVbDngbFiw2fmDt7rD
knC2Rkv9XndugRNnRjcY+y+J+CZ603ecqG6T9AsxzaHHAqVCh8pzhfEtfnfJKNZ5JQ5a2GRaMDp/
Dqa991lN0fjVcS/UV91FJF49os8p/MdeOiGW508TMhC/r3e7eRQfD6GCPVHObrfIeFWIagUCIbTn
RWpUGTyrTLIAQyi8IiTabW04tGMl7vKkDPYGiIDZ0so3jGtenQRHn+a6LJv412JGRNuW4Y62k9c7
eIbKIuEpt8tSBuDStF04Xc3vDDiYSIj5AdG0ZNnUNsK3TOwEaIh1EjtCZoRMuYoqlQ9Kbr4MxeDi
hMIK7O4Tyx8P3rJuwhlEc1qxg6yRafBkJzTmlbzisrzS371EnMQNJt+uUJRY2uKRssi2JFtEM5Rm
REmzO8taRazB7MMOaM23vUYNihaTZIsYZ5GWxLlx+YbCBgcpm4YzNjTFtqcC3H/B6Mnq5JquWWI2
PxZMtm5odTgy8hRkuzbudMnvovEtoZmlNO5HQQtgp51DCsPgt1o542ZCeP9N1uaQDuwDdFqsoZXn
+/Cn3I4yy9Y6VvXeUKuAYgT02rLbNGISYZWbMk7KHu6Dw270nYO6eNcvzqkv2AqRcD9I6M0/kZts
vRJHdKmemfjz9pa7Nn0pTy/yrbVKvg0xl3/gjU0P+NYHemXuvPjRApbbD1i6+sEGuQJOKaBTUKqf
8syEKaNhoEC7eOu7aZbPE9EXPyYT1xUvFk2eEsNsp3aGim0xVL8glrzfaojnXW94U9jjm8MaCxWb
F/M+QGEPpyMlab/2ZZb/Z4AymFyQ9yC435ECOqUF5bdrozrjErWL/5yZWatESTvTxDphWY/iPPBi
JNMI3WIfFhtHCrLzrvpkYeHk4IecPhL2Iu3O3MQnOeTra/tilebnWkBwVPpI+FFtZRdiSmqQN67U
CCBXFrJK+y/1g7c/oWzUQAQ29KRQmbFPTYbcik9/wD5OHcIKXvwkssfU68iPEnHPjku1KJmZdPCL
uHn+N2+jPU4pnb6Jz5XSrVPZKV8TMP34t7ZYHvGQssFANGn6foGUujp8HX8STbtpBAesXmG+Y5r7
zVPYdqNUFSR2JsK/MuzUdoP9beln9iicPH3u6FqzcJr5TGVHK8F8Xk4v2+SXrgoGMupT4kFYNbrk
puYRTqlHfiV0S/6qGD3Ag9t5ff7fZzyVmNL5ow0theQERPyn3eyhGqOc4ZR8vxDi4aoU3bewWGLs
o2AU6fdj7ALH2i34GTVifpZX9iC0m17QQFUlDC+kkRD18+7w4EfwFh47zwZBc8A0qK+JEAyJ74cJ
zVrOu9QrsfUWHp6AMcX7Kj9Qu/U9ip6bOcJAanskO3v093lct9pUA2R+LJHqsF0o+S92ujiV+Wzu
tTl5o3RFiqwqNp/mmemp6BAJbL+llkaE4hmGFknwl1FA5rNneoezeuUyZ/Ua0sSuXnext8ODaYgB
ce5+rTPTXTI5gFhcT95LLh1MYG96tGv+JyUNPJ83PG3VCZqGiKWafFDufa/eK2Sh7rrIDoinWbrW
RlNIgiBGaseebb6QvYjS1bIM6pQDQYsZtEtNmOp/ll+BiLy5p0H9Dxp9ZJZDrvhcJho/vFjfaKi5
31udVU+TwFlSprBaQQzuKngvCF1ILw+xyo15Ic7aXxo+kb86EWgDf3rthBbYXmBZTasB0i+jG6Le
yp3bmfCi+/gTmAuckcEUCBZ7BwZpS7+MD3riY3uNrHJP4Ka8MLYjDnPVjIBxS1gyy2uL7Txu9DrN
C1MUe+0x9zyZmMwlyqbBoIZk0sTFMaV8LAw5TRpT9UvdhDllH83Q2k5BlcbzKC+L8OqBW4jf/Ynv
y7ciFDQYYk2FRUPxlIQNeGJi3OPVOahMJWBAUVhbSGXe4CZYS+Fp/xmZRjbtA2jSZu7uqlQ3az2Q
++a8PmmWwC7+L3ygPi8VGYuIbl0MipUdAz2g8vZuAhy7bOKcWrfiFmB5SQXyoAaTPhdSWXZdWF7p
Zv6HJkcgk/egN8veMGB0y/L+x5OOGxTgsoz2OlBT718DV6s5MjFjVItB7AlrbTDRi5Y5lp+WT30y
Cgdr7zY5WXSuB6tN46V01AGFYPxZzQt8o/HhU0/XrIn9M9MiCSjl9DjOVcrViameVl9VMFkvWY18
az2rCmvqSwIny53Y+3/l8IctrTt9cmgQkX14JKbalcAnTMNRiekXAFUdvPbtQXk99EbL4FBZt1X2
t0IRe98fJcgefiOKC/Tlr1JT7Z/4lMiIBVTZq0FdTJEP0hiBVttHFB/bZSwQjziNhtdgoO6teQ7/
rbpTTe2UtGPq/nxiHTmKOZJRr1cBrxP9Z/AX4j9Qedp9CJxp5MCicsrA2eDCs3ZCXVRCR8ii2AV2
j4cnJ+9d6iARq+jnv+REB/mpsdD8mfuVdFt3zO5GN5ows00t1qSjlOCdnXkrWOUAkNSNbwdFdCub
eAtIamlDmDY0Ffx5NdFVJLDRmrPolbVftxAcrYE/1YOECdL1AW7epc5WVYkLeE16DX0vj/AWrl4F
4J3dq2h8LaloyNSNk5KutHFbketB6pNnv2iXHNBYOSlAHqYei7zG5ZfbK/7I213kcyZVJX5R6coc
1AB6leeWaYvNcchKQ6EsJ2lDS/dx/RADXwgq3T8tngsgCKSEKOCyc5nbORugOyJxz81h5r4gdPrb
HTQkCIMMMQTeE7Z0lp0XscmikMgqDobdL1JhoIcMt1KIfYa6aFycfe5KrZmhuYVjQ7rMnAdGl9o/
FWdkEgTJkNyQkF7W1K/G2I6XHPIGDxxsnGhmmTKxPR2q5VB/K4471JqYxXfojG3qNq7EJ9iqO5RE
NowkDUmEaT9ypkFBfFQ+btTgNnTQH+iKFKjFnnCKXnKwrPiin2j5CuDIefqILfRlmGcYDJZfen6A
UGuSIil2AAPRucSHzakaVoHVt1C8BKnduw/vtu1SSy+MHFafrsK5boaLgjyAYJiInn4KREMh64Kd
0EU2fywtCeTwZ6eRBUkBfzY4y5HF4bZQ1/BD2QWN6jcEyh6wlA4LhIhSm3+sjLjEBzHjkOpTfO8p
GI1GDYpp783j2cxFvW431T2FhOSswSz7pLKRC+WxYNzXBCxfNeytkY0y8xO3yIFeUyQgHRDxml0R
Hr1HCN+y+UPmSNYrVRO2nFaxmVOmecM+arca+N26q1pcWreyqE6p+IrUL3sVBbWv3mwQTVhEFFxe
/EWMInyS3kNfhZ05QzCPAjwEoCBLSTW7NGZ1dMYF5sR6/TY7kKbCAMsF047OizXxJYHR3tfM+3WX
hxBAeqZW3BgxQ7MwD8leGXBYH0khTspiDjHzCpCAipAirO8/vcEEqBfK9e3lJbuSQnePYMn0mb5i
F6SxfKmD/FFQTHnK/0l8uJOEC5yAH+K6mX/9rGcSAD7h/KvSuSPUfScIo5tyWFXF1ItEVxXVthnl
x3CFVDHaaRKhB8YkXit3pfBAa/TXVoS6jyxO+qf5bongFMy3vWL0af51a2+CxxfilgUeHAXJFEQC
QbxUx3SBBmPvxjxRTF/+RPQ/RMR9Wy5ldW8X8ETrpp3rIl8QvxISO7hUajYDN6ZsteeREM7EWVjz
wTyz4buS4I9gVlTT8v7yY7fH9W8exn9bsa1OYw8I5EYUhezg/PfDkRaF8c5iHSLo/3L8wMdBdSFw
yp7C0Ni53P+qUO4xS2KzqAsW7nirn1axLOOPESqxYyucIfHjnTtNdh3a3kafJF+rEyAExpcOAzI/
wLHxjXPVw8aP4eJeDq0oY/dz3glRtLtrqE5egJIhPNrthGuPxNgsYiiCenqz5b6S6o1Q9HTqU5l2
URhTsKu6IHPqoD62vkFFTXnzkHj/vIIn/gEgfk5+dWtQxK+pv2BtSjxQTXh3YvgqCqQRJSHWqaUX
YQMBE2qjSQSoUnJX8NCMGXd/NchhWdOGTqlZlAyVGYAkyqQG7Jauow3v8rmmEQ80iB0DXixzCZhr
RGk7Q3T/XKBTEZOgac8qqxYo13ShFlPQTMifgYocmiJ8fnEXJz/X8N9XxmBAqkekCch2r3xxecK5
ggH2wYUJxqt+3x9xgIJtIOxWF107FHeKrNKNE+Vq5+mP4lT8PywuUGiIjWt2O+h9S1IMXz5W6wwT
pf3r4tBvhODiu5fnYhEVpl5kuVqAHCF2KNN3m/rosmDqMrFzicI4gjsl1QUvrre7zeaN1ZLkoIbH
KQTlLEwajvMyjJWHhmwshKeGPMZrPWQ3YoXSvEhUZgu6VXzKruvHj2QToj4hs7w4BL1s4CICztO/
3IqbG49qkX6kT/lTL8T6B5AUoxG5l+6UtvFLxaH2XYyIgc64MYr8ZoY3Ojqz89bef2YjJjFfN/VW
eeIQEzsH/Pk5COshXPDd4u9l8ar5xN0oXQC/zP5EpfHhAhKrcc/ToP/9sH39l2ZMd8ys8uQJkQkK
CLJJ8H2fT1raq/+qjoe/DVDuf8LIvBQeUp1Doz5xKHbT3fNx6Y+f8zW9EmlFy/Phawj4F+8na0x/
7D6yHUZWSERZFjq7qsfa2FYxAyVWMmaM+qvG6ABsngkh+kGFA1Dft2slEOS8yGuAuHiBekXahJlg
+gO7Vj5omWOABUrIBwiaP75a8qwNtgYo+pT+H4iP1PnyDUCBdhATRtzD6EaBdckVg5/UbbDf/ksG
wT27x9CHXCNxblTcG3pryQClIZJZFdSCvD1oUGgWVw27dW3+6qoGCqEc/Am9PiZT/BTmRGNudxrh
DAI43WaN4VyE62BJQyQRMqVUlApij1DKDfJESH5Ww/SzUrsFRwHXmf+ksuTvRgkdyeAxNUIifmMd
JmVZ3M8ztBeTEeS8YbtzbZT3g7Tqws204rN1Uzgg97JEVsD3kdC044W/LOCFg934sHtMcctiqMKT
0fCpkBngOboHwEzO2ni+PPGzbdTk5qGpm0aWl10TVZSKbeQQyqX63RvVX77d8BCHB2YPjlNGysph
yTpKwc4jwW2FLslhbvO1PuuNFHlNbr83DxljKP5M8GcZRV6cAlXOOj7w1sCLiMxkl9j0TQPAhOBf
znqZ5plXb0q8QQesQpIuxtW4c4XM8ZBHBVhZINWC/PQ6pAXudmYgJr5tjaXF2uJFl/qsz50+WOos
ep2uXhDu2l8ObrhrhuKHnIKQ/vynUOp/Caj7TP/svIC5nC59pYHuXHqtsWcTcsehk0D9OAs/pE8D
B7YLf+vs+qhwtV8Qn4tVCCu/n71VGLiT7B80LajSp033j35p+F78/gmz6DVn1X045p6Rc+aAeLzT
zs4caGH8/llQHnFB3TGkEQ8OfjJjmw/7kLnL6XJB0KMJzh+M03lT3NQcox9wjfsZdnkMYk8eprEV
H3kgniqU8ipMFCNVX1AoM07qtwa2Pu8B/Rgw7uzmoV0p4QQlQ4uFK7pw1DQxbNdZDH6J8L4eRBuk
gaabAqKZZwWu/R4qKM9GNKoV6kQzhwuQFTKmZJNSCnSNy93xHXem2dDGlvzUNuV09WJP3GOY7aD5
qy09MLZgSbEN5V/RU9eR1hbbaji2XKwCFNdZJSBHWQrv5H9AJ7AItRlmBFmcUdgMAbkwOWGN61Om
jZNQErBzgo1uOQawb7v3uzhJewa5uP1nVC8ST9+rEBLYWb2SbMYXy9yCFiq+sdg0RUEmwZi1ffdx
PAJK+vbGmIvae6K2XnsGN55zYVs9deQyRyKm1EJP+j5lEikzHmMyqZ6jaTjT4HyjXgLLPReKkwLy
l2/mv4FqEeMfaP1IW/eKXdvgjc5XmyI6MunBBL0ZsbDkIZkOLWKF2thSOf35hNiCJPBNeCIlkPX4
r/nsouWXZ+VVPF73OFsmA7xgF6SxiNx+UgZpC9aeNfP84rzQVBq4+I00Qha8AKXgA5ZFr8NP34LB
xlNyLG2VBLsavq9DOjwVb1ww1/yR81k3XXPUfN3KT/sEfXmq8YxOxFFHij/LL/u7pp2iRz5nIfOt
Zt15yZnCDqkdKuJK4mlTnEploJRvHkqOPU1u/7fT1YdujjBvReorvMETlmOKUCkxagVYD7vCl+bI
ym8MJ/tYztYH0mbzKjXfmeQwthYrJzJPnYPZEGu3WMUncW3ByYMPjmeoHf0dIzPWjdpoEZ1mp3LT
UqClk/F7YhghkRGK6m6QNlRgkufd8qempERXRXFfPDlxRZNQy1BZGRn+ABaM4lPRxt+DPQ8wXKYB
6xQtPLHj+4oQIT2e8wvlgAh0WGISRAv3V+hSjW+Y6qkC3w6xhf5x7vWjiklcljCYp7P1SWf5LlVb
Z1ZOUYH6rJV90bvTuNpsllnpD8Wk378bBeCnbEJO4Wq7DvHPCv0no75aIAdrzlvn0AYZ5DAb9qkC
ICCns2M2wQ5MzFgejRvA9t/HrMOZCxBsagJJaRqMU+Dkp811aPHxCT2SniYlC/xLPR0GWmtrkNRD
PVK6uXVxZWy3T+yfKktgSVYQaA7ZmjGUL3uAnHqSbZ9NiunzXsNrr0XCuKwc2/bredVrQvlm19FU
5lq5ui/Gp6D/3u9/sCdpscxm75BzL+1bhdzHGG5/+z8Hi7+ju2YCH3BeT5dr25Mjhf5ZoUsiHp/i
OXCy/lc65HD8AL9tBx5dhrTWRoN/swvxRE9q/h6/lKCVb1u5MqUU4K+BehpH899TeEIKUFR1M5am
EjVLR1/ZjoklM93RksbzOVvs1lwh6QJa1/3ScW69HKtgDrayLNEcaYSALNA7OUGQmVliYSpRONnW
Pr9itQIpqgHTB0DnyCI0hb/oKTU0byWMonTnAjZKIpqsBBalM5VPJdxi0TPtHLeQBjHo3TV1gKq5
+B4Q4qJPSfUDdN2Y9ZEJgKw5xUgXN4k0JWPJBNiyQKcM7MIH10KnkWb3yzsPvaR/zVmQvwB91pCL
F9sSDVyOG8OOSlbYwSa56UfE/ru2VX2LAoVPZoQtUuv3XbzW0B2qV7AJ6vpz/XWbCFzsD/LixnzX
2ykhR1TT5T5DsFobKFsImPfUbhzPX4Qf33/E+8q43bh9QqWuYPFKV7ufNuOWkxkDKLcCkrGuTiYo
ZcH6PGYB9E28F9AgVwsFBWZy6eByhLPC31CyBpLAQGB2R8bOhD+IDMW4UavyAhIDXalCvpwDU5Cc
Plt0zc3Z6TgIIkQ1G9C7sN9rLERz0OOb790TI0O8DqEUm9AWP6kdfpic38fDZR7IQkp1dGS4ERLX
Rg2Q+3fX6mLI0QneRyoSmze33SwujBNKCT1moJbqbc+2j94DFI73TbFuZnSIdpzdRkPZLp39eqbs
8rzbO/mgGW9RkLkDgRGlA3cqRI+NuNND6PIeXqRBRngMvOGYqYzWuTYDjUKhcVXbcZ4UFfPtVj+4
EBdP/GYoyI38S9a7piF37nmAcsrUp+pYEVUbd6TymN2xw4pa8HGvK+LoFAIqODdkketDoQzVq6ko
TBkcS1WDQdvIIULGpBvmqQdvtB82EPwRQGjNyCw9QBTboB3rzzhZBR/2+zRO8W/BgXakLtENVoNQ
4wiu/SMgK+Yj2SujhU27sFAolgkenOL/CpqIwUUJStvrPTXv9x+zNPjlc7OHkuJlOXYvpd4ICWge
rHgabMbKEgHCZz0R2NpdqiLPO7EB81twMpI72huUpi/RivvweJqB5TxwDVpJcscp3pgLPyByJbMH
T1EGSJy54myYnwmaxQKcOWRPLswDKXOxuHxUAAbvOZ2V5YPTI0GLa+NEds5ageLuH/f8eXLUb8Gk
mUqlrPnNJi0yfHW6pnQNbMkxXeerJVpsgAaBHMRNlp0+8ro0KlzXkKwA/AHyo2jctLIuPrPQPWQS
QsksM7oaoXi3MAhCBZ6z42l6z7b7VrMpdhZ75USVwB1snIY3WcoltcfF746Hh1bm/BNDnzKJTKzn
TJcAMtSP6ed8dWR6akZKrofvwXgeDsC0HTrg4HRxiv6olfRpPwuyr7X8y7qZA/v09ttHoDlf/ft9
jih7vlAv01QX2UsF+0OfB4xamJm9+P6dOT5/ANYe5n9clgSd3zB0/43bgtnbFH1teDKJ7xWl8pqf
ah3/KsCd1f73R+BoukklsNtYv/cKgnBXfMWXWzxTSnJQtMGFrYbcuC5cwyizt5GUu/6YhIZTOk0T
BaZx7TitMO9DW0cS1ACNQB+48/P8mQ21zi84+A+zBB8871eUI9F6+ACEJZQHlyLMKAGMil92FL//
UtAbhLIR5Zgb4fRwb97BI2O+x6+d9gwRveiWiegg70qHyQzXvxzJ9eWCADIemaazyHKtXgjYJ0mz
8fHFgaPGu9m5H1t5tG4+sGkxj9O9jT8GMDPi1BJfer/r0Lyej2EhukgaNtFYetXKFczd/BHOoF/Q
EuTuxCVoGPFP+iW+0ZlBqyiXInEMolJMMaN7lXMlHdrldQVXW1FJdlu6AvCu9nWzhMxs6hpsKMhn
vVzCd5SRIqRrpRZezDgQZulslT1AWhUeM+fsMCk6MAlqxUxHInTMOMpKre3cb89cACcU/0OPsKuL
BdsTm2KmT5Iugxueo6wkC1CsIQv0RJu3XxaU/uohrYi3TTXYJPoFocRaMiCk6FHWWqBRMAedGoYj
6ebFMFFPSJNW1Ra8Z1K9197nIuN5ymZj3q7UqkjcnfFtHEJ6FazF/WxKVlBLiQJ9Q0ZjT2q8K7/Y
PGg/o4ElQhDMO35Z0N8800geRcPTL6R16ifcVSKvmRu3hcyXPoTmmfZyJUcrRWpNGYODv4GRIqqA
p2+0F+tK3Zoc+qHpLNNX7FDJMLwBQRHu9u/pkC/DTXRT6UamuZzcSQCpY2TF21Sy8hs+KmnIXJLC
/8Nt4OJcCMC+jfx60JsFDdc7NiseFRrHV4GwG5aCO2i+HEj3QeSqwuGOkP6fVe0LAl2HGvW8Zmb6
xkBAcYOyWFpUNt1S0iYz3uD2kHtFkc/qjELPWnjm7RQVCfKwTzvboyYHJZTjeSBRJswgoBrVxY8i
KlBGRetoyUoSGxbp3o2zmOFrrrK1I6KZsGzeOcmTqk4p0Fy/O0QiGeA1EEOL8jpQAE8Rwld50EHo
iyD2YVT/1Op6DpOrTLexqaDsmKmg3LwCy5NtXPwlN4ynkWkKSrLTDyzIEFqiMqYBeq2AcwOkZc2I
AgJffNLQslzVEY3EqKqN+mgXew/YzhJOEHAIE3aT3T0S7Y28wzT2h8CLygP0pg2QaT6h/DNY6ull
SyxRuLUmTJM/uUisD957+2NAJfBBiK5zpGUMDoZ4tOj3KXMdwVjKlWwP84GApSA3jqn1zOrWTYnv
oM8Dz/Avj3fTECJ02Eb6rmMsoxKapIcEACqt8AlAolktCkcAfoor3SPA8w4jjS7Ql4B93Dn1iNHa
5c5zpjfKMgQepDMHah96EgBHJ5L/Njnz/NXMsLUBjEj1PaMUKuDvlqkODsqFUGuNsyK0YE41fBP4
sFhzQGY4XmkSAA3yQqvUTuweAxD6G6tpvgBnlmFiAgK3RppNlMYO+w053/+Ht7GDymJJ1Nwn+gUf
Q3d8l2WkFbi/sga6Qu5jeZG35naQwLCGAkNrRYzZ0m2EJA1xzhCkXRBklA+1VRZJcp8rT6wcT23V
yzELDSDZGfBWkixbqxLDKBAcYWKBj3sSrMqlQI2YCKfFLaIoGj5Cdv24eDS/T81JHw15nZC2a2Lp
i0CLkohfWWEdrB91I5qYkerwTqJZ4+U4H/RkrSJaxigVE8Mo7LZJkoI8fWGm7hvHvWAXCHlLRwUy
qVwBQG0xX1saRBJ/pRgS1aMsvAJzEdQQDJWsPm9hvHGU4G0lmLjfUbDooRJW6fwkW+tNOqr86Lwf
gz1eRMBYK2Rp8wTgMldS+4BOBVggi7HJrnbzVtpM7Eds00FoLrgphxNwkrxxHhjveXo+1Oq9ZVTI
cWMbhQeAXepdpy62SywuSFPsOGP83IHjQNV5SAiDtZ01MwgiljVs/AmZPckcJ767R0DbbVeFe52K
q5TosUziXNk4XbmipMq+kHpnTkCNjO2MN1L/MBYZyvhqpNXTuLA/ozVimuEDKieitVfoT9Ion1kW
1C0d2NLI20yjck0XWRsj74Ck6D/2J0ED0gn830Bo/b9Qp0sa8Z+PizsPdxw9CWFQDFKIsfYLPypH
8jCh5VOHHisuT7fRxbQUWROPCI2G5w178xeu5Wo+B2jbek1RVv485ujSujMIhGZ/xfCR35piC39w
1H6UmKAbvOQLVESyoaJrWCn/TKaM5Km8gGl4faiU3QkH+jMAxhEhcRJdGYL7mpKsDbRraml1xX81
sh2CZ3BarsoGNq6QXjN9kA1jpbw/z8NcNoUsHbmxKhgkqLWbdR1J2Z5IEULInJQwnYLiKg3ySL9J
S0Ld4qWiGxbsfq4mW311Ev7TnTtPEtYj0nS3DG3c//LR7VziyWphjL3/di5WllqioqT88PgL2dCe
Bg14gyLyNjv46ugWKmtr6Hc+wIwMWhMCCoPkBcbeAnPyvO8ekA/rA0hVgY3Lfu7R4FaxSpQY1+i4
zeYJOGcKXCpjjuBRK4OO/xmCK0KGef3FE494kz98mWirG1tNOcW5PfQS7HP8HwvgqNbtkjfwx4mL
BLfNBWXVokUresmaDQkg4ZKrUY/u3HTPLArGuJH36MpR5KB2qglhosI4wMkAXAZQj0n4kEc9K68n
cvh5gNIYbohgOIEyrjjmNK0RMGji2hOA95XzDpmXwzAE2tShsS9FcJX5YBS9FvJV5z39FKSmbD5N
vsrCx/mCAEuMKCCVyTSXFLlA//uBlYuc5/rr3qPj/GtGblWMnofM16DoLpHjWIpP0AqjmtgLxwvb
qgX1MKnD0xG7VWNWm78n6xLg6vuUMy/iIlU3w2FPujpCTGFd301j+hoFvw4JzTAGPqWhkq1OD19+
VSHIG457ZuWivENNltn+fF8Rh5hQAWT2gzmp8ngrUgAqsY4940siema/17r6PoZyY+bZzrUcPW9n
DCAQ5S9iqRojgVHhjvQBgPLKrA0AxL18/Cm3B7lRyDIaWJv+akGwS3rqjwBiU6d+Ohp772mXtkBw
+exENJ0u1KTHPZ97OwtNsnDOtLVFdkALv17ZRgsgdjAWkksCCNHQdqPnIwvD8zH6+5OekKljwOPb
wwXETK/7q8FNAjBLSTzMUFBpxWc9tPvxGWklcQcgf+tCBPc3wsyOIHnvhrBuKGUBHAPyJsz8oZrZ
8vzcLthJGd8uFKGHAxPUWklR7JI4hYgjRWKgRUuXb8O+vDjAF4BEkxmw65S1+JkOK29qC1ifF3Tk
ZbmSdPEFK83dFESYWu4IE0ccRJwPIsGzeVsRWja1L69d5O+G3iwGTweFGfi5W8unxoaZXhVp9M9U
LS/rJcOk32SN55baHFCAPMN557dew/lX3tqPvNURQizxgm9T0gbeDeBx9ByKkIEpi7kNo4F7CteD
QuwIDH86O017jPN/pbA4kFecKaywT/fhrNDQyDy8tO5dJHpNFWIzvSJEgP32bAVR3j/kugVYLmT/
xLvwYfrSyznvKEjMRBIA3v1jIkEv9TWWYjkqLVWvW9zOlTPQVMk3xxr8a9Q6bAW4ygK2QnNwQZOM
K4MqMiLKcJWuAJ9LUCrq9WRK9z+NVZTo9Aw6ryabTc+dtTjxdyAw5AYSuok5ZV2wfpqKoUTHGnbn
kT14Yq1RocI2Ms9gnyKqEs7TPOiqNbEZTAWhNa0EFQCcwjjEw7P1Cb873p3rUQGC+isq1GXPxGCg
hgN1Y4hfLr1u7rreaB8rzJi7A+wnB9mPWT1nryGyqq0nzrFjfi0FCfd2mOCpTlTFLEtdZRdNFPZS
xq/YtRJDb0ysmEJENyenl7QKTX0pQiRbpBZ5lt4vFyQpe7kzjn21jw7eaZQbwnsMr08IvOMzPHlz
lsyPq3N5NcmwMR0qe1dkPbKNXgvVArdGrmGEp7Apg3OyNkg5SvzVB9z+m36bTqRxEzuHs2Un7ILB
kWLw+hr2uAcwl9JQO2eg+tyji7Jfo6jSkqBCNwajaD/0Fbta+X1wpV4eTv6eo1dQMkvCfk84yqnr
5McwPYBX6747Sc4ZEbUwe6hCCfpyUPs1Kuus5TWzYN65L2E3AdaHVnSzfQZCcga6cCeEaL9kHMFm
tmV1X6Z0mGJcpR+tKIkAZ+bLPGQ3WMuz/PUzawNLo5ZjBcBCevxbWrGT4YQSd4XvRK8mJY5cCui6
c9tnbwURIydS2V7kJZoREAVNKyoV3H9LIapbiC9sn9CF144yy+2x/jzxLRbV070Kq/tKTJFWgA4c
B7981LkCR+yd0+Oamho76K7nlMuc2adkwoTNGFoGsyjvvsElMGOiN5Sf63e011czfxtaJreC8zIa
FfXRAa398xnim7wWK3fIvncfEfjXMNzcw+o8xgU4T8Zf+stuOVh9Tsxr6jovjqg3PYrXVTSGDfE0
+Hrphfm/TDBDz0z4VGW/DQ6tZfySX542CanxiR1MSdgmJna4WXhaBIh981Uu4d+xll4yZzpCi3+F
thQGMm/H1uLojhKB5AGqbYj5ITWENHfbnNHQBq4CSjDMn5HFWq3T5NCVzWcFFuiBwsRJWBY3yGKG
Ig8A2Ysdy+2xkZCEc273Tp1mmlIu8yRoZ9VID++yaPvUQL0/p141y69vHuxXMYk0UKlSNYbuUWml
BmW7K+cVOzAm5tZL4OEiPVL+rvRNmy+x+/D4NW+cca5HDfyXS+oddxvW+mxFskczr4zw5iOo0YX7
cDqnNwPkQpbxaqbZJkneAdlIUNsUSXYQ0qNb/5j2e6928FJlgQfaVTfaQOSbGwCPEqaQ/5QDiC3F
GZWDcCj0gkaCzudHCyBlf/SLmdnBbZ+B4I1e5gcL3YUf/OGhtZ+gpjfJ7Mjcv9sT+Xo/SkKhao84
7ardJZARvr7ABz6B2+RdjG3aUDvx7QhCy/QuuZAP04fjiy+61v1WaLfkQs9vVRWc5AXJ7yLWFQKc
0a1wl952A0KWKzc3D+okRbosZ70UGXZD32sS9rOKJvsGKX/+pZFcQe+kubLNrfJj03cRECBNGiJy
N6ofpYjGUYe3CPqBqZBzk+KH6C4rhcDF5W29poSQpRUL+WD5e+g27NPvBdJg4JIBKDAH78a2RCKY
cqlerG7tsWKQTWDeeBOa1L0sZFOogSaDCK/jzQuPm6owwI9fNnaYK0x5BY0Qk+F6NJvAyJPnRhJ7
8+bdizIQJtHR82PnqRyhNcrVQJma5EAIqliBbz19jgAbeRZQ4OEcSvJTCYWZuYZimnGwnHJlD1O8
EC+xYX2jt1VWUwGi3m/R4TU54OGG1LFpcR2bpdlAXQ+/fphpmoxNbbCb3Bgrfv/gmjb0F8Hi5uov
/8R3bZVohCn9E9jfaGC/UJmwVOU9FeoxrwapYEVth7lyGkp0HmFZhaJYQ/cwI8ZnyC34PlrWCoF3
RQjbGiGhRsP5A5kYjM2k3S3kvZRraDKoWdWgU2bSPT6LXSSurQHo0qabmAGh+wRZKSkqqqvXSR1/
trgH+mkhd2Hv/N5Q14s5WhIlRbN2GYf4znq47zatVzDLGOVvz3Ul2RKMUMf4kNV4JL3C/EQ2Xo5s
t2gW21Id3626HQHBwI+2dgkzr+gznkEi/HlcoDeK3pDiNXFUVjhb3IlbGlsS7w206oGZMOAfgPYE
aL35h1hHibzW433DpGTQP0SIHfF4BumQF8nrzu5IiHJVaYMmZow9nKRRHU//rLQrNfj5WZkfgy6f
Oo9fgwxEuvosFBIasuhYnls2hqP0mQNdltz/Nu7Fn4OptdtxcBrKdXd4+tld6FO69kKSVAJN2buz
haKFN+hwN7CK5xQVeySw4xbPRDAzR1QmkxCCrtg5iErgVDSmZDHTtrCuiG6NgI0ektNt2Iu7eSzn
Ps7Q8zUoB9z9ZcxuE5rvhOV12KLss0KLMhZ41WRdn/fk79ynW4g5PQDT3NZeYg7ClSwS03nLVhTP
/cxKf96+a9SSwD13PEi8dMF+GYZecDyVQ8Npiqz6gfSQrXGSE4VqEkcHR1O3vSBiINHCA/Pqyj+a
tFg4l1xCgN+aHMGO/dg9SD7WfWrb/NdhXCYDurH0nyeSAnuE+Qp1iVMLwVzzd94D2smoZdWSyXRz
5z2IvZOku/SAsLwI9kJloRLkkivbXk0IHvkCSMA8GNO48OJ/k3FgYmNGybRCfIeLiYGaLKgI3vYJ
7Z8NfiQwBsEetFX+AILutvy8gCFau91fUOqiXE3FZ0l1xAS+3PoYbqegnSLcQg3lnQqH8AXqOF43
aGOIrzqqq5zqcjnNCraA5QnomlodqyP4NZsxsJPTbHPF8jZ0gi699UHiyuUp5xtrON4xKjl0SAxV
emvmJuEN5p+Hkl+PKtNVrYypo+JLXiVsNdvnr0f2uZIyNJnN9jwU3mTrS/8Ek9GkhNIU4igC+d17
wjpDwidf5RJ0ImbrbwxBVuinUT7H83NNAk9QGeuNMXgInQYo4pxu68ozsEDGy94CJEeY7AD9t1pV
LI9ISVAW5mHDfKWEL+Ccq01dcgOsJb3ThELOCXzx9oWHKyBngQyUDMakYZx1qKNOWcDkl0eNCPTL
ygmyz0k7FKZ5eZ96ij7SPOlN+f979/9IGhjg2raZVijAvinlmifCs70mrby5Lt2EF11qT4O6xd0c
Bo8QklEToC7HOAAhjpCSgPy6/D4j3vMnH35e5YvMiirMUPSAWUmUab42xItsZf8cuY8eJytFt7xT
S1Cdht742HDb/ricQWw4RJ2hOXtwv6kZnXrFC3t2QBAfukPrfVt9CpP3xEiQit80KqSUbMWgi7XC
Pw44fUC6GmGkbQc1pXxuA+RuIEKpqID8WOOILrdmJbV1PZ+XxmJerJqOXrJ/+Yf803W/wDaAfXWD
KBMMLG9cpehYoddTUU6BFO3DARt40LSlFRzVnodwpxjSPe72SAn6dVlvXCyxXL1fqu2aw8Il2Ryx
VMAdzxCYge4PECMk30NRqrtOkmtSl6+xb9fC0HBrXdb5CMVJD10eD6vg9ymNZYyXlss71Of+SEs0
RUTSBtTodBLNGj6Q7KB4rxVDUSQ0zjs5xrxcxw7Q8lvzbXxyJMNQK3vEMjEQT7vgaESQG3HkNVBV
OFacfkquBeedwx3e74JlVIgYX8HXD+sckbu2EkRVAK7dLg5oGzrhDSqPoWleAdFTwHv8jXYczI6Z
L028HdbbRuhdl+hyJVeedB675f4OPyR9+K9Gkaw5mQLc/8Q6/362WmwCqXuDrsPGlNI45fiQlJqS
WT4mEba7cXlHX43PxtiAHE7kZ1M5LHUDNHHNAjAdjDnZZ+pYnsbX2ObxAg0uKDMr5TV7GUsUGkyU
nW0UNsc6MIG1vZigNp10hDSS63hiGsguN7D83KzNWwLR8nTJMGjNeE41JCPvaWFEytI/XFP/fWlq
NSYPwDzkabBXIqTls8z9JM9fQ/iUDoOiwuOXTQCqvXoeSVtT0boP/f8LOoY9ZiGPIK6IMCNvCbOg
STKsysJZ06U+GMcxGmAyAH1y/XKOsqmmsLL/p6m4xLl9cr1LSwWnrv1d+Ttt6dQYvPpj3+KXfJMx
+TG++2T2AYgY44TTX5CHvMXuXoJsv7bsqPKMQsp9Mzp9IK8GGnzhfkQj4Ti1LsAkVEMcRWatU9pB
WEDGBXzpmTJeFE8C+xbmjMgkqKGTYnbQd1W2T92P4rzsqJE/LvqsaGpia1znJO1vH1rfqC3UQcIG
S44jbEMMfAK1PS/iJWtsgZNkzlfd6sOtoNf0KWoP6L8N+GhmR0QBsFCy/cvtjvf1LRQ2y/iHsXP9
I9zU6+N62sK3tAZUVfY0u8Q9tZNH5gpLwUx7dnB5cDMgx1wagNr5OIqU2YNRWRtoDD4YZL0gaNLj
U9aXpNwiw4AgAyUxbVwyM37Nyzb7dufUX9z9zgpLpe9Jrz7zOMWs+AqXvlqUah1sIUVvZ76Syypp
lbZgSWpjskvp6CwLb7aloVUrygYODHj1vAhxkzzPPogUieEmNaCG81TQt043b4r56MtRXlUzp6GH
B9mtmykwoKYqXN776Pyfpg3Lnd+cM6hp64mdSG6irEDx2igYuPub3/orIIWUekeL2tDvdsK610sF
ZZcnZDbjhI4RjQOqWH87AJVTedEAIy06NSl+YbHNBLOdnAceA0pbS0b3+k6GgQOVrO+d5YGuA/3n
acCEkIvpMQDX5WJJ11Q62CYLHW93KCPvCOzydOXNFvLMfC73aIRkNoOKbpEnJmXvEsr2ufhWpaPV
DyEBRnR32U6IuYfT8Zg143/ORIgeVDh2QaeOQ2SWMLQwZ1ZeGRX0kFoDO6h8awfPH8tW5Km/TuJX
uY77ut0FpmF0E1iPRDXTo0m+P6SrdZRw7N6e+XcP/XgC29tZcTX8MgyeJdyAqBpXIwPPoBBss3Na
ynbkY3lsv/AwYnT26nlO7pEX5WGM3/S+g8aWzM3bbsqfs6WFWzWlpRJhvml6o0nrSkzs9CpAVfMY
UuRVCjeDGD8rblKEQG1bflrzFRPBY5dJH8frw+7WamRjtWSVcf6f1StwUumWiIAAidSzWwOiYwIJ
YiSrgrTlKoZMeP6HN91ySp85jWejnNu51mp2iXSnHrZ510OvjO50cCDq8iYTsaje1kRh8UeagUlf
hXQFfBpQnR1pN/0+KSAjGLwvsfhsnVMCREPuZjCp2u2yDuUp6IdekWqnBhtRtcD9wr4br0kxGPfl
28e8sq4IujV1lbea6h5M4Ng1Yyq+rjBunn3ZZvLJAW4a/7Bt0lP3S6ul6AYTNNFF3prHbeISbuUQ
087kVcBypDdRtoEGOiZBFI1t2zvUmL3ypKGn6rFMQBM45ShS0w4BExDn0TmICbMXq3ltVAds/yQe
G/JBH3T6Lfj747KdDyr1sIw5z0kD3Hb2OoPrnnRGQ/3ywJGkQb783B8iMiHfAnQ9s8POu8wfnATP
dbnzyraDhLr6YFyZ1dZa7kE7+1nXqc6GaqixrGKLuqCheoP4K5PfuQCHJqFbKtaQblLSEbQqRAa/
mT5qbuRzCUC1iuJZ1JatRu+uxte16jANrwSaPRhQdL2V3HpZDMn6lIjwWnq6R/vEyGQivYKQwxkY
GhI4P7bVURcipbJtn7YRtx1YIaEaY+kXR/F2jKDorIKa6I3Me3J7qZLnd+tbCSHnKGqa0kfv76F1
XgIhMHA4xES77k9PePshsoQqOlZHTEDYRhuJyLPFthN7NcQX/BBVjhq95MgqYW5f2covmwzUvt3c
suca8pnmk3k+eZOn5Pf5I0MBhW1ptUfVefxoCwurt6k/Zz7MBFysMPwTUNaKOMUF2Xay0OK9EPE6
wENqEJrUw3SnaQzSd9u/lFCyzaGmrrSvUkHK3VxxeVsZ76xycNv9/9chJ+DDFTA3wJyPydiGXadZ
hYGqHAaOmfJBs+CrR7TigmHkzHl92lwlN2eR6grL/tc/SGse60HWFgMfChrUvpMmb9jnqOmcfe43
U0lAkPrxlZAQ8k6Fee3UzvbAenhtZvfVedKq48dthXRaXgC7DSAuK1YpY3AXxOQtpWZBiTKNOb+s
LsbsAO/Zg+F2gW22wsbcLke6buIGZLKbAeDxBzZ8uN5Qt6q3vJNpqMHQdX6fdKaj9gmGkMhTTBVV
/384gsXiAzKZKLQAUkz80Fm/R5q8jBAYF+Csp3UWGG3twxsnhhroY1gHBscgrfwaXMX4Lc90M9oS
QL4oxEBSC5aM38mqfwdjB4GRutRyC6O4EaB8PlZabVqW59x/hB781efj0qrxUhQiugtxz3lxV8xV
WzlLijU8FAZKtWB2GanyU5oIMfh3LnYsg7oYpWCd6PVoBlcb7jHA1ueQ6BPgiuY7CnHHuWw5SBlc
QPTyWw1zab3C6faXwBC2KCAEr3EPQnW0qwY3HxTagF/jzJcktb8mBLIqH7jIakfYHBdp6jEo3J0X
T7m1qsUaZKC3NndaRXdzkjVXvjUIVIO2CclOo7KDbNKgEjZVjw7AwbRn/+1ZDisKlZJZDDWhZ22k
XpOz1LXb8gNMlegaknm1vzPrX7j+7HwSnC4dBKMBIyGssY853Ay2qRSW4iAt1y1WwnrHkehxWWJY
XofkoIWqdN/8t6APYfDluXZ0XBazNEp7DOdzikQ6uqxK6cTY258ss6IPYrVNPoTuZCjE1yJC8OKb
ZRTIJ09FnG/PR1CIbs4P+f0o0kYp6Y+2k6j1dHB8RgCpygJRiDSd0z1fgOPmj00Zq/cfHk3zyFpp
NDZ0Ue3N/0H0iKwh/wpNYHdAhkBrU1TcAREvrasMWD7gUpLPeMVELaMGuZsG57PcZ4J6LvU9c/Ec
tEANKPPRHkaS3GewXGmjFNVNUzUrKt0q1d1Zhcg0EsBVdZW4TYovBG10dabRIZfczfqaEh+1YTVz
NkRRWVB/rx4eUwJszwwIkEt5KaA6aLY6IXCckqvw2AvUrmmH+XNMFNBXiBKImjBD1+1hqJHFXPEP
k4TuaPRHrsSSsHL1XFaM7Ko/fBCxSJbKr5PDZylqWaq+Ws9rW7LMQJneLInon+tmNafkH7+B40+Z
5X2QgavqrTN75rLPmFTCcsrH0COypyXrn16RNTDtAs1tywHcScP52u0NU0RRZyezOQ9Ijmd9Ui8M
zn3V8Jbtdk3A/y4cYKl1C4GxekBuu/0Vvut6ltERs9jVOeJQ6k8CRFGPWDA8SWASv2tPVtUac0KT
HzkaWimI4TSBz2TRVnpbPkFy1IQIQU7bjh/Rs7xKugE3jJVY5iR8SkEFx6x+3ZNtVAEDY841YDUj
koAlqNDWK5yIQuqKSCBBkWr5OiyBCeCNGnnIUCYyT2uncCaptWubQyr3atRNzj8nbzXxd6XDSQ8e
1CQFtx+VzL1HSWCXMmT+TvT8PlfSW2wPe8Wzo9IRiGEQdLN+vD5XeV+/Y3qRGchTGHmqgMjnE2d2
k/b8gAB/v8N12OSa9gix6a1HV9XYs3gl3ki2+b6oOaFsucjuo2VgEQjA4QEYCzoBtB3X1YVSvxZp
2+uihty7CJvuRIeK3rHtvyTwjhDUl9+pDBC5JZlWwbEOlLOCVWowA6UBSgB+IJWBI+eQqPC9HV/7
If/9Nk2bJogElTm7T0lhs6MI/XKl6v4aFC9Mu25rnZc6QvIZC6moi+XTSADi4E8/YfZE0gwLRWcO
jk20r4oBbCGyr5TXJcY7g7/8eNXg72DqfiQFnlI2dxqTb2+yCytY8lK/9yAJf2jfPTnMyzYnrvwU
vglsXdQyVyTJx46EVNeLd+aCBBWKRBS1MAZPSw0oLIdyjl3sRGhfv+sfRH5nNmoLWPlpccwosZ+V
gKblmETVpixwunUmcnL1UW4grI+AV/GIvKVZo2SA3Yj21HYVfzMoZyVy9x0mwZnehm56NmcnI3bv
VG+RihJIVI8dBLp3OZCBUV5YjedBLukF70/dePWyCuT8KQCNDuJ5avVZdqcEydAnqN2nYwbT4ixK
Q4TRl9pp81L+kT2prmKVMOvLyKpziP0qEB2xZbVZesnS2AEydJWwzZU3BGoNA9gxyuK9m7mtxziM
VfAycMBbYnyv6jlHWbR9786d8/HPpUgwVsmLaVQXJMZGePSFccpJ31Ce7RrVEB6hAAUfjKmoC/Aj
Vj78eCZ64aBd3rjR4M+hMAIknj2sJCwuL7/ePx056E9bpzwq+1wMY/+ULWFlpbh83HQt1zSC6M0n
x7szMxDB6U94lSUZEfGToJPw7yqHStcac8t3IQfrs3fIHy+c05mJOhe2/EICmbX8vCcDHiNKkL6V
TlFeptpPLBFX8WouoryoAZZ2OMtI/7HFEFds2OY5YSAjhTNGqWnXL31xb64ihqmQw0+nlzmm+Wn4
g2Cccnr415/pD3qk49TILv+zYBaM4tkurvEytRdOtNGoMZRpegCJF/tAxyi+znWpSJfJ0E/RypHz
Bvg+hQUmo+llEcGDQO4ls5aMSFyYEZlsMu84xuFnyYiD3aztfYcYGn9Gmy2hlyAfFVbkVL14D1PS
5KmdtE3h8x0YF7Cr5B1XQtlmNzIjnQNWrEcNZ/7atR+A3QbQC9yl9VXEh9ScmT6R89GU7u6JlEWL
NP9CkA96R9+xO0T+7LFJHdVZSfKj0nJ0OPV7rLIhpvOdAjb2xYVtxmXdArGWBAstX1sy1FSdbtcA
crXIL02kiRFM8opFdh4baF4mfmmFY3SWG42GKWZs24RRdfJWxCVY42y/uA3a1hjVYEDsQvPu7Q4O
5azlNdAB3xP9/Y+541XQPanWWsZiEnaExQIRYw2ayxTIvYLKNOY6Zp5wt81iK1tYHQvk0ERaDyUB
wRAIjYdAX4Ur7jc1EXL/EX4htTR5J9sXb5U1WL5ZUBiAbCb7s0O/DypjoII/630taGpNp5e7aGjw
sIDLeW3Zr+TCMGyQBf3i0mj0PSsN9jKIPvV0t9T403RNyLnNRZZYYGAcnQgzV8lRvFpHM/YACs8B
KZbsU+95ZSdKNW5gBwHtHA4qDlCFwxjSYeGQQkHFCMarvroSUL53xL6/09mDOyj+PE1glC0bB0kO
qRjP+ZvFvye61aoLXwPMjn3AOMT+daE+qk2h988ljdgF2IxWMRWjiCgbDVvtDoEXNAudAne81+Gi
FinrqqMKaV/6SC5gSTkiPVpSzACPTmQn02rN40tSvGliO+s5+DMIjoIa5CN+RamxAmgQtSVkNznt
A2TL+niRIat37lS4xz3gEr1q+a8Ros8/T/ZvA8tdB3ctKZwt1u3Frso1QqvuiRBd98oJw95Bxm//
6RixkUey6jIcCq/pbtZiQ7XzjhHaQ4ciSu9qAuiM2XPkbM46pg85y0ybVJu17UolDVXZ+qT7fLuz
SIeF0iUmP96H/yYkf3Rh00vMZxbP/bThNwz8P1SwzhJ86D5XvrqyGBSRIjYNB2fwRXtpyppya66u
hskq2w7/wkYA0hxjBVKOZ4RLrN7+CtxHvaORDfkeyBKjPhZiOFjVhAxDWUT28Mfz8O3x7F+OtVui
y5VT9xVLdorvohgiIWzEg+YFgAYLysKAssbUc20IKfURb/BAAfJKTxbYnsutzwCsRTPjNtLYo/qF
0Ja51K1hXAykJeg+CCbXj967z+nyQPvNk8o72HEGisqmmVFZQUIbAn7IfScU/a0ndnbKpPgjfEKn
UckTHPJj7M0yGNeAfrKHk0gsJ6okrloJiAw5tGUBTYsQhiEvH7tIyh0TKEHk2KZ2bmV7OvfDeqGo
Z6qJPXo7EbhG4kY9fVbYhQSMb8jIYn8am139HEsrdYzTKkkCFywINiKHBclAi6AxnrNWcDEPwJD2
pigqom3Q2jtO25aYb7k/Jeg5bjk5viB287Q+KyBJYzu2xbi4BG9qBsKDs4SuzfjuPntoGy79uOCQ
juxsba4+eNrW3oNaOliJKz+gHYCyVjiBkjCcW5LzSbvcAigmwcRTfa5qExD3/Ep2FUG+Zwa/+lss
tcJV9eEoU+pmiePL1uBpJerhp8FYkFUhnDLF14I74BOMi+9FVp0IeqPu/i6QijYF5lEhuiZbI+TH
gFUDegNDlBcxg0jBwICcORGCYVCxbTmezshjQg17eyPGWnFsGA0/o50WYYrX4LHYUGc3THshqvjy
pw4V0Rifqs46ydTchXct9Abr+Oo/q4VpIfX9fJa80h/p5gTtBnBPwcJl114UUWvDkZMjKyagyRFF
5yDictEVj7kitP2X68x4YDlb2iMKo3oXOj4Nca3Hx3rssY96jk3eQ9phjZej3nreqwD80P35IH+b
a+K1RR8QZE5RXYO9ITzkwYGNcdFJ1FidVFQF+G+2UsfAjDw/AtnNBFFOsxH9ZXvh8IZNQPV93kB3
OESR0MxDTGaujI/Pia5+cNgt/4QucRNKx+wo51ZcM/EVq6XG6LHQAoBF8+foco3vXypCgXMMljOf
i1Zxr2ccZsVnJ0TroYYBtALYwj+Nu0cN95bFuQodwbtLItrrMRFVhaOK+26YkxdmunEjw9xojMpL
MzYmbeahPOAdeIvs+aCNClWkrVjreSeZ33sxxuCZAixImYW9szhDaYCeeJepyfTwBNUa0LYEjEBl
vfuugMwUNECVCJq6cslub5wFwV2JyJir2YxtEAn32aNM4mcO9BzfMBe7ap05mmCB9ovEFF0+TSKB
WvHT7G0eI69KumkxET+9nEtFnlVD3lMLMusd6ePk12ovvsNmcseHlWii/8+ucLhGKj69S7GOtrsy
bajXt6rlYTMsel1lcSpf0X34ylwj2cIPZyhTCNC9JMp1zScJVLhNQUp3Z+dRXnsT8TBTxTDKhIBT
PVqfnkgOwFHcrxGu0v7r2CfShPqdPipopiefsMCKzuSA02vA4tutP3AAnjIUqRjQfF6RNFNCZcud
hPhY73oS6jJmzRRXfXiu+l1yVdziVTYHrTjbrcQBLVBHH7miHx5m/KOjARuXRcl7UQOyMQUjzx1+
2UNsqEbXbLYCjatGb8IL1S0EHETAuDRuCpfd2HoBWAjo55NM4DMOqhdtzP23ArG9SEBEvqJJNcY/
euYynzidssixLS2SoE9mYnFmzt0A6liU60Thdwc7ON0aIhNaLejgM+cqNaxLAt9tBq/gtNoifvGh
dykItPjAqbRbAYowWETsgWyk8rqHBK1JgJP/X8LWKWwz/4Crzumzgtz5NvnKtwUyOFW1oco2q0ji
uYTckGwdjC3Xs8+06q0J9wLLBkHe9QBeAa5rFqpnhtHy+D22mhIFNmzo2omrXFV0hUyAXLbWBPej
Lz2Kvy6ZkoO9tbUxQoIgPz8vPt0n0NNqcZtXSEsuHm3kPtwhTLPjArJZVMOyxd+W99Gb9RUolaqJ
vBjAA6GOKR/feQk4gXsXi7XHXJ0g+v0CRupQrSs3zgXkczKZpuQ2DzUOKwkYgFsaGHv1cTkC7V/O
cTZ0KSrtaYoXoLF66I2oNEYW8mv7r9A+g4IOclc6XxmL+B8pN4P5/lp6Ng76hu27/OCrmKvI7Q0I
+ZapHDiglVx8sNsugziFoj570zXwIJ4TihPnRlNJiAKJBiJ06p/oSYKC0Q5H8w+89wrep+BU2v8L
2WQxTAozEuL0o97Yc4DxgSPMdOpvJ7r8uiS/ulRs1ZYcWsOEdSVzt9UVnrikeFlvUgG5BEJyK59o
o5o/HlJU6GWPcCgbN5dRgMlUv4V/O3VdvJ9OqRmPf5MpaTG2dtIW5DpWG4hHs/6jtuC/KrePqrkx
e1/zraJo7j8nBU6ZHYchjHAZ6dqS8Wgsi0s4Uq916EAWTtOdct3OySSruXBUkBZcR+StA6CfMWro
9IMHvGbKDXZKnphagDV0xA6oJFa8RPnYvq8BSAEmU5+whzH5F1JO1WaYHfR1DfPV95Quyyv/00pU
WNoUfHSeID+JOHSQUyrElP4d7R1O/g0cRlTi99f4qDhxvLLrXdK0lnwDMu0aKzx1j31/GHr9wXpR
eqqOgLpNOPcpWj/szt+2l3c9Xo/dJedQFGpKRcrrkLksf/8lw/JJgjFDm2CS7hebcaPgrNMQFErl
+1KiDEil2tJfVk4PTMiW12iNoHs8BfRdWyJITw5iCEdhbUmOD99WaiKD8oiHbXnsXdmOWBTf8kzo
G7IexN3IxXzUdYl4PagQzQRdgToV2xVc+pu34/EO82Bx4LHgFV59LpUCrytRXYMlYFXw+jDg+Jnh
Ai7BWSDGpjkUS5Z4Sj/zaII1SqJ+MfYeuCLgRteHi2lDXHbqPH1dVFuyeX1hwdTmKugMe8FrsFzc
7yOCaN3jD+7eGgrn+UYG0BjGZbsMDu3L3M6s3Q/pR6nhnPR20vuU6mzrBVefp9GYQ0ziabCAtxlF
2/OW916eK0r7VdQEInudkbBldTfbEe2EHr2eNOiZJEWGWUiUTghS/cVStJKGu4znm7fTlXe8XXmz
J9XHU9tuJ7AQiMoQAD1qnADpFkqN9AH+g39ZTqicl3l23iT4tC35KXADAi7egZkNwmNl/6X5Fumy
imLQZsd8/zSbituJ+/8Z6o0bGx6au/M3QxfK2S2ErrXMv13vkg2GPaID+T4lwM7JiYr3EUp8h2Dk
Yek+51qmpXgIjGadyq65TcBg2WQZj6kVowNB9pi21gnzyxC3c4bPTws//pQTDqLHDLf9N8yvn9X0
ZWM8ZMwsW6WSBJHqn5R5ghPscRRVGlpqDVj9AUHot/Pe9vUhTsnE0D8CPB5IxdFIko+35gUAHQ+P
JJ198f/BtyjCmD7tlg6/nPeAQ/2ChaGhFQORiB21zikFjnuoxcSxNCJsNREJiF0R0G/Nl6tmCvBY
6gAe5UQyap7f1UZUjt2/m5+eECzEYLz30zoBgYytjnrgTIDLs9+X8Y+EqQzppnaQQPAARJj6up5O
OuFl7nQlMgaR72RHgc1oy2QJ0rN3TPBK78iFE+72JombR2HYoEMjUmPaKsK5MonFd+CR9y20KdR4
z3XRouV+J/O78h/jGu9LUiomwtqXjVyMwM1+Mycj2fcrAiRbsqBUtVv2zMTGwFoguYKVIcP0JFHc
txNig1kXc7NtnY1pijQdXDZNgE54/UFvSORRQIyU7DxtOVsV+9S/AF1vr2u1h5F1YNLZvNsMoezI
OjKW/cZMDeIGoIt5b8vbZd1c0jjEioTDogSGxOzhaTskRBrr4ce1MvccrsI0RZZF9xk//w4v0El2
lcFPMTj/caA8pFrgOVE0ditpBnF/tpw5U5BK0K6YaHB+2hHBDq858oH3z6/yRgGflIyl2NCU1PoB
mWZXF8bYP8Jg3HE1BIatZjfy1qZ+gGkyIm//yUwRYxjDiaqIBhoUHdCiR4+gAUhzeK8IuXkAWOsZ
wk1qIv3i0otfCjND+D3jcRZSEj7NM5q6pMMw9KICTu1VnNusTA6175/sxsEugEn2ELxgDDHiGowD
YrybdYGl2LxuUxTcDywCTSdPBjG2X4nhQVVUGCVvXNV0xQL2AIpvSqG/zYp1/JXYNgY25EzH02Bw
BAELiJommXOEuVQdAKIyV7SU1oYSQdCUgM2n2pDcOjEkaQBfeJIbh5/tJT8Vhuj6190PBO12KmRD
FnTOObBWK1pTsCwmX9CFsplblWWLASug/U6ZKcNWrZAPIe3BPsBa7INny8ixQ8UehqzaRJvBtg3u
ySw4I25diGNVGvWDRnGlS/he2UGFSCUNC3aMp0SALV3F/0IN6VFN8BfNPiEvlQTEOcBXThMfBEOg
teUhKhEYJyriIwi3c3EEjIn6NuUX0V4QX9RgKtLqnTmnjMX5HyP47dT5QpDALFdMvCWzJ4nhKUX5
quaP2GSzY3NBC6mRqvb9k3l2Gsn2N9Ur8xia/Qk6qQuD+jtIyYootzk2f+Ngac5ofoNAfO+7Zr23
yjOojdd/p30OzuQWiZPkdaJNjGbqvPSjLENS2E5HbbLbRjSMAQZRmG9vkr0ABoSb6Rj8WUQkA7IX
qzp46/HgFvHXx+OVdHbszBh6Om2nhVKECHGvKBG39VOrfFOz/pFKSQT7AyQl0AIpqRl8opFJvoCk
W+l8trFTFvyjxj6Ytab5KRdpvpw1YgzhT2hKfzRghTmP0i/Xwdf/zmMfjl+8FXtD6cRkOpjw5rIr
vuj3CeEtryZjqbhmYa8cmCZ8Hi3S9BRuUF8kJpdruVi00AGQy/wzoyDyTeD04R56LlIQJoJhVUrP
DGDco7IwOxbCFDpFEpoGMwDfwalAcv3GvaLoWoWR2NJNbpCwM/gmojqhjqXZxbAzKVDu56NutTD0
qcnRszLABLvx+neEKUZGiZZypDfU6d75lFGTBsOtx/8iPNxqD0brhkaY0e2eM6JNXyl7Aqyy3AOX
Yh86nxS462AvNO++G7ApH825aOQB3nxqW/XH4bMAs2PYGge2DGB3sAEGwB9Zas7O/EqtRgjDABVp
3h54/VoCAcHDmDuFhOAZLbd2ZO0VRiDMV7TiQQ5lKLzLKAFtNt2+jhPvHuAnjw4wbeR1TaJDfnLp
6Ipg4af+QVyBLQkJpv9RC3GryQRqbJ8Y5gB9NmwkJPLKm9xmGzhuSSJX3i4sOPHlOkNFCtEZ/+eC
mmY+jYI22NTK4CNGxFCjwhh4U4hsfDMaMblAZxGxPvd03VO2ZLZ1K2MTouFTxPB3lF/9TcyPKp9O
PGCm/HmFu7BLw7Ls1Kv1BMGjvVe+P63aeKRziczcmklS9OMtc72FtmJ9wRfWqMaMLNqykcqIP+Xj
oSo1YvB/sCnniqw8dIxb8qzAaKNlFhLMN1RSgQGU+aQxavW+Wxp07lQtz9eodF80w4qsUNsMKvTX
X/3c4voSQv/h9wgOyG3zi2kOMVCb098/vTEQyP0nkgsZxohgvudqgAX/db4UVxeL577iYPPT5DgV
xIW+JimsNeNbn0tlVxdpGSI2bkRBnw7lo6biI2X8z+BWkDZllg0Mil0kO8DkAFq5wpt/pm3DyT2t
C66p3T13kAR235D1PCH/JFAPZEb/s6IwYGhIVzrzybrdL6WOABuJFOLWSFJ45n6l3zRXqhZt3t5k
mu40kqf4Xs3o4QFhC3XMNNYFg5vAJMcaPnfCG23+6ZbVG5b0chHENTEahTla4QEiBtIxrRlA3xTU
/SU3Vp/MuAz6Uo6EujRK2wcz3z8BtlMnqq/S4Sa6l6QOuxIJ3OKAv5qFauzgIbSV/TTTAZ0R5S7m
g/OK4jC0KX2K5bTWmyDEYbyZJGxkgFuaSSxs58s/so9slIFXjJGExEXMytzxZid9zPeU05PhUKld
8l7l0GUaRoevEIREsRzwLiGudxSB22EKsRcaE06+gDF/tSsIg+X7GO8SXldt1yj5FNytHh8ec/Ki
8g1uL9MGNpiz2SFZNtXVBtUH4Uj1ItlUVBfVqVmL7qZ/JqOB6XHLWWYIK/h8rQX/KbWA7XZDNbzP
RD+5naewhWrWgnujtbr+nrUHW1c/9NIQD+OsfCpWhKG2xJ+nuhImveAElX6MXKaKQXRc1VjXmIWk
ZSutYnrYdRo8ieMSY/y30PUGUirqYQHVE4bR5bpZWIhagq9KpEEIuMUkasLhjK56BIX/Bnw6A10S
gzTft7CeMN4vANrb35CTLT0N/ZPBX8CxutSrcNpa9CTHIoQBCE//R/k0SURAii87i+Pu6sCOq+op
j616DmTAzpjlDrQ8V5vzdBlSfYIe5kx8sn1dWEWK/HAPdXwigSXEdeNM1fjD4npSHBXW+LsYTEwQ
6fNcpwx9MjqhC4c/YBqjRHQRWc0tJkAc3DcX7dwfFsXSZF5QVFsBhqddLSi90l9JU8qcGtPrH0TR
lhOlzcW9F3qRrgfRHSYQtBMWNvNRYh51kloQeoh2iApw1zHSAEIG7Ua6XRMJz497wS34oNGDIcFh
dFUpRoRWjM+OYAfpUh2NDRBil3RTe45sTCh3vCsdfcDTT+Lshq2zuDJ95q1gvTpon/cyQTMZK2T+
/0ttPT7QVTOG+bpJEsN4KKULLA3G2tHUrQWbFb0b+llBW4O+kN1m08oqacRsKa13hOSiiFrv4ncr
oeDkDYmg6koappCTLz6wQ/yIexT3N0IAc8iP0KN4LBHcYpOnQeYDatYJdH6qKjhWJNnaI0zk4BzB
kt7LGeH5LS31+Y3C/CCzxEOA9LC/hPe/bHpiCQdP08ar3W/3hCFvPBZFNnSMDISdu1/uFJghpz4A
O1c27G/hXziEAnf06uzeBsuhyw8eUj1sZ/AIoFQGCEzyhO1gy85k8rg5Zx5VLMGkFW3rFGEX4K4c
Pp/RcgT+xPRWgowJJtW588Vp4XRcGXb2pQuk1rd9K+dvvustlPaexrvJDitZG23VCPwwbte0PCgt
gpRrDbQbMQE09PKQ5CPBqQB6iDG0or6jgyU8xBDC071OHOns7h/5e8Uv83HWroLdl+nKBFwka9L/
Fdcxe+0SfJ7Xuis6WNMepFIYzsJVBd/PNTHm/40+5p6K2IN/072LWw/Xz2HLiWq3Q2CzTQw4s/0+
LIfLdNTNLpPQ/HqsRIi8PIcHs3KvULrC9Qpgn+4gfmuWhaWVs7yAohvfnb/nVYQiBPSAQpe2rEpX
25fcWezKz7pcVgp1NkFoma/a8zG/nU+/HhYbiTDgVTfcritEBykf+MQjXLl4LsTftbaVetAwBM6p
siQIin+e3ST4xasFwL1v+QLYFr6lYlhvKwPCYW1XWKt0qKNjHK0pRt0F/ZQHbXRR6I3IeXXNRLbI
EFRaiDQ7Wn9+P1u+EFSF5AgAARfI5wg0wFBo6m9eAfb21i8nrHMJ8c4YTf74VnoQa1APNJSta+pj
xARWgOqxTCKHkDCnIqV7vavZLaNt7d2mYVu5mBwWuW/9gKU4Ov+tvQSKb8JSmW2aIiL1fLIOZCty
Y/BTFolbG7odchN5V0xeI0hNs0e6+hfBbVvi3YZ1go5xd/EujzTsOmNJhNvkrKsaKZAD6lQ1zfk5
3bok9u+0UAB6fwvro4aSzJuvnBeVQV6Dw/vHPh9CgbG5bf//M9MZd6eHmGxw8gU8Gy+wdX+kIila
jBn0Qk2vD7tU8ROC35RFOqEZ7AYLNH5iCQIFF4W9630lGNCy0wroErGlQJNK0SHJBzOSlj3HByIR
45E7DyMhh7ewB0yEJ+BOq4lrtmaUuCNFvfvs1T20B2A9kvTmjBRFUfF96GShH5gMrMoNdLHM3fln
aZc0iDgstJ4JWihkmW6PB1jujvFcq8BIW7QTzP2qOF+B0VDwyONxEzPz/a7xlxUZ+p/sqUdvHIhm
a0HXbwME1w7Mhnjvx4ajakk4ayTQLFMyuQDURIvsMNdEY8cIkbCzNvIXVLg1v57ciu9ZLQ9lkprO
8EmtLisnzWD43lDRGDyYyEs+3J1GpzvXzkH+VGlZ4xBL+AHdUFmNT2MoIHellMSsJ67ojlxNs00T
IEGClpM+TCSzkpOIyY5VbipCSOhORzsSyiSGqnM0Fvs0AZar+RKfa5fAhicwLulzJTtGtxIWQ8Tp
CUTz85bGXPfGlx1VeFASj0T6ebFx+JZvircjB2g+8jHsWW7GfRMUs11GeaqtdIJIahcJtAbVMir2
fuKk/LgRe3pZSRNLQViZpB3Aay51oSepPmu0T5uuZz4AwZHwRQamAKyZQ3C9OiL+aKHDF0OGZGqN
Lb14fB7A5DNbYPWcIxyUULzBFFkP3t9o5p5Y9fxhqoutGXetN+lR4oYBkiRyYOn2cLRllAtL/BFm
CPcn/f30ksh3vsUvy0nDBZQfJVqx2HC0GmEfDdrIFDICAwa/IHTgYqHrwXvrmsxnpSwHDJOPMMD6
Mga1MakT6cUHS4EXwgcdm5o4pqGxiaLLwGxEjXGSjjR1cQStVM/yqDRbyOae/84bOnNR3NTBnZFC
Sha7QZTv8KCmpvfur68V9s1PluVegMYM2PQ8dvuOKrlXX1DE8K2qQSstuHTPpnEynNYIKzrC5DcB
6uWyXXXNDW6AV8/s5tRgSeb10ipAPi2eukX+LsE0w2wC1hj8pSUBDgR+NgUd9AmrCAPVec/qS7OO
E9pEZoU5fV4DtXG7uC9XrtsxJQCytgnIPlU7WvwHRpuMjPUXiwZi6V7P5lQmTEgn80NsPz3Z955U
twla1GgWKTSi8+jhsXElsoR+6Imav2BWesWGahCZ+8WEo43lAmz836LjliF7449GEnwAyAf3GMP3
CBzukMqTj/+Kfd4UJC2qR5XOX4RvHi+b5lzBAWXbQVK0/uvZ9Jn8LdZZyIPHVuB7Y+7BsA+r0Bvs
9aDjPJXJOz8XnNw15DQZCwIy5KOK5lB0QASCLtP43BQCkZ/eWgKoOpsYzsqRJgSWKu0kuWE43Iua
cEXJ9lk24eRJOYW39QMs3MlaPkLgcc5fgqUYtLYYYlesJfhy7QUIa5j6U62iwemRHONbqU9s6x2e
ALc9NBkdwgFJQTUIh4vAqq+Ki7v7zd9Hg776UrokI43MTGCbmDwCmMMfDESWd0+oSowAJlMMUba2
hrO6INtaYC+X1+XpNC3LR2l19GjlHOyujjeT0GYWftcHxkhfYa5b/GllBVz2vS1Ai6ZFu8GeunEF
LQcrL7S11oLEvIAPvceH4bzKuxOFsZX1x3dP7ar7XDjuwIzyg92yiwQlL3UO5Cc2RnKqKSxBHHp0
3ZxgJ9UD41SAXV0EL26jLbEb/8UzKZPZw5GDR8n16q39LKBYqshI2v3Zia5eZYLIB5mUgJUhWhqL
GyPBXcLcqntyXp0qvjtTFILamrPtryklAbjCfeC+oglZGCJvsYN36vxexjGmgbAZ47wcrTrZiGiW
wi6eti7ROTx8hh3qaRRzvuGcaPpupyWQhoVCvzMnmCx1fEjOJiJ6uA0CL3unmk5EqLFNYk3dLAE+
0SSv4RgSAseWzOBE9joCGfHGZKqEuZCsaUA8dkdmX3Uz7LH96/O3/hoezVmJK2ADwa68AFXO3HmW
OnV8hL6K3so/8K1O+heCw1T2O+pqNGiKHeg0Xe572erXwTL7soB7PuAqHChE2/9KG9m/K9N7TJY0
Bw6q+yr7w5AvT8F7d7iyxDVbVntbyZdTdDy4rSnZbZdkw79IpZ41O9VRoxKXQHYJOzItkgfihvl4
FtLn2El1AoWepPmY7vFw/3MYO+KO12GQZk03Z/naTfAeUwpxENeg0rxjjnfvYEbxJugv4koXlJf2
WV6YPoBSa/HGEmiXXDLo06GiRQlVR/KaqUHDEM60oOFeZZRz8vr1X1IccdIznG8AnzSPSMTuS1gw
jEPj6DyuW4iUAQCAQb2qqBUD0Qz3mFF3A7hKOggkwh8Jq8qHBDteTmPrRtJxrEP0tbHj4CnzyDwG
/eR18kJURsBUCgiPs2yLiUKF288Wr3/Pr7gPcQwDV+XYddo2hYSDNwpOCDdvM/JQcOFh7/rU6fgX
KrwYAWtLgqx4Us0ILeIKn+IJ+lPT4XOFkc3Dq7YxL4B3kNau9v2+R/5BzwEq+7+L5mnW37fwRBjf
URWvQLJWp8qJVxAYRNUbk9dLcdM00qK2DOAXuN4WXZM4s6/LaWikaQegrSTTiRpFPVBy67jM6E2i
iz5YnydQXUyS0SqWq9G3xPo04L9Vg5NgO/jvERcEF491rzapo8KqzdSINF4QLbOkAFR6OaE4juRU
Ufa9xhZyLUxrV6GgYh+V1JKVKCFZFTIcYzgRNfLRzhC3jEr3j6RMcZcx3HV04hRL1zrFBCcns3HI
t8hBJ4mcXRTSvtC9Dz2+eSlMOm02mCIicNL8p3nv8NHk7gAZ0EOBJRayynz5UEbzPz/je3THnSNL
C6oKUPF5fZQaFCVwpuzZRbRyMnuYS8ovpJhRxjzP8owTrj7IaKxmML3YNnTIZGYakt2aMrFXYBBe
emEFL1DlwzF62kNnV/PCx/oNcxyCF9d4VLsJ58aPkdQvYzdxcGaGpw4Z0TY4BG6T7MmCWWLLIz1u
GNqIkf2aYCkP7M582xPsbbXIR4WgZelFJv3ZJQ0l98MF986bhv0TgaMjs8nLIKBKB9EBV1q0RdHR
Dkbb8DZOlaPgy/ywiip7GNjSumEd8nbzO0E8LCwPSeYgsZgumZjHCDjTk6qeIk4xdyBAWIPaX5Gj
PR9v1mqBkrLcA1LSNqiMQvrjNmeDiPq8dnI55ufllS5U+l0fjDpkNpH7w19PxQPfd4tqioQFiyg3
/IB0eWpXWe7k7tfWOlkwa93/pTTs5vkQMmHTzlwYAFaQ8oHJphvakEchg+RO0LrVtfqjSevm2PJ7
XazwfOFoul45Bi5gLywneWnH0t5UivHSmxqCe8JBAwnn8k3Id4F1Q6VhqdmnUB1OXd1Hzogn7Van
MkiTo1e/6s533bzwsjsbVBxZAqOxxyQR2s+EevV89w6cA9AH7iMHoporrJVxbuI2AYl4M3RZnCen
q0e76fLMZ2QnJ5S0tAOKUg7wq9MagisxheILNsqEALywGmAcRdoOyY6VOC9ARkKAynpXKApTPgAC
TxsQD3dRoNq/JdTHTHFQCIcYOBZq4G4Aj+kpEDxeYOoeF1SKRffU4UNcN7oJEn3cXpqkLrs4tcxs
6xmKDASEhiSEU+HAleTpNzHgpvzmhkW0jckFZ47oZihk9OO5clQ/QZjSpYM8C9yggaLzsrIwXBhU
1SAPODIxN/jZWZjwtd2HmnReieDYBDxK9JmS6X6XRqwZmQrrs4z8l6NNva3h7Z0Bh7tZhKAewTBR
svPL+4YoufBpxoxRbJy9yw2O0KjTU2r98vtw1RXLiaZYwX1YI34Xdsm3UFWF9qxj3DaEJCcKTN0G
FbYH4sZG+RWt9kcxbrb4co5W35k/JuR2vo6P57/WgPvEIn3JvHzNsNKcxH4VMCuZmP4Q5t0nnwQ/
EdkTfyBhr9hlia56GIDvj6ZhbB6KayA4mrV1lLdHMgweYAUMIJUerXBqYDP2Q12NvKzIKBuXgfpG
i598ziL2zxRPJil1ddP5yP2Yp2XDBUQ9HNcS6zjGqF1ejufrFBoe/xqgQgDpzrqMyPk1sIeNOr7u
hCavahgwLjEzUFrRr338tI86rKZNS9SuDAAxp0BxsqUgdDBXOmckJu6eUDy5QJYkc3sI86rWOLIH
ch/hK378m0iT7VfE4th5sSLLRECg+Cem0QdUoXHSbZQjhE4V8FllooGua2Xw+k4UzLJPYJOrsVZ9
iWJC7DI1Fehb2cBvMHxs+Wb23WQ9YVHelMtgcPUhhM15VC+UF6MbEhBHULnxOAcASpYDf930oFrt
m+IPEUo9BQS7OSkAkm+3R/yTgVHSfaeu4c6Dx1S/NZUEYJ53lToBM8Y0QbeggraEv3pSypxKA/Ir
kMD/kqAHxa9hiaIcPwihhIYwm/SPZJDN9TyWoPqXgxoGppCb7Xp70A0xY1InCb9aM8nYjQ/GbBYJ
0W39Go/uR+HBofn18YZbXntalpqMvDbeB/EvAthemm48AD01UtF7q3UO4EkYYwtryk8A99uWMlFH
zB2ycAuLH9Qw4dXzPiRjwzjpteQpx7fAlJElDfmH2PfjMfRAIsLLAPKymgCLkMBZ45Q+DTHjG8bB
X2JPfLF2G49HDocEFFQyTjj47Id+G59IRkLmh8U/ax7sgBtMRavz2BnLy8501MMSBEDpfQjh1Mpk
VcaZQ4WAirxT6ojhTItEnCrta8Lg7APQzlBjhjjhrwaE7x7Z0JhWEu+z3YmMr/uazXNCVeL2+QHZ
KOC0UUddLIDKS7KzTIG7wweoxjYlpBTt/r/RvnadCwEGam7330sRMkHz4vy/v4a9qSqjIAxaukKU
iluz77jLXMQV3Y9o1SCZeEiZKRCGCugn6sbE6ySJapKL+9p9L/ySpR0YR4gW2vfCS72lta99BWj5
VY9+wAFhflKnAdvvubUsQV7CopHbNVJUplasjCtB5VfgSZEzJD5HRFe7zETIFxqhLXzMWYcLN+Ub
xScoGpeiw3WqwBvYbAutV7ShYXG5v57tqUYz6wORv2sATEKi1gMAZ4j9Q2ah/GjpoFr9MVqctM1B
FH9vvJ5fCY1NBnsn++JBkpYOaUDljAEIfbK5gxpgZFouHjuupc5jrGVUHhloER8CniQWuUtC2ku/
rtQ9H5g/bip/AXbZlkIjw+h0w8Jj4QdZqytpNiwir9wQGTDg10C0H1hsyMs7Oi1uAnmGKQBOS9Ca
QxkB6K0wMZKIzhAvMe/kJD1vZY4rQp6veD4zo73Qo/qeSL0+77KpoBLscX0oELXZS/y5GR5w1aB6
+PxDY0jokn/7ZH6uZzDQNveYAu3u4qc7BacOMkvqbyxJj9PMMClrdn8PKg0t1OTDVeks3uMOp9u7
YyVN6+AUyXBhC1PPv2ubpsWhhiY1z3URTZQzSY+jfbRysPCKSC97YF5Xa4dyQPaYNHJbxCD5zwjD
BeoemAorjwKh7g2aYl9RbFTWir2zINja38HQGGyQZaQ13f0QkhRypHlP+5F9vco7Jub3ZtufEe25
KlxzfNuqnETQHZ+sGNukJcc0CPpAsRH25LE5H/ZmfkarFREIcOedCHZY7pcIQNfc/f3WIpR/hffE
Va8arIRpw1nhohCcQ2daovb9d4oESl4wEozYDHilMcTxU7sAxuJEXzIlkD5RHcAH6UPk1bmt35x1
XOch5n0b9GrdgR7Ps037sqr18lwdAdqMRAkw/pr1RW9U6tQVo6IvYNsgfUfhgmozl2SDT1/ecf3d
coHbrNnkCIUYbOihovDeE+fUZU8u4fYHL0tmazoodNYDWeGPI5YjYs+xpDZw98C6tsMLjxJ7zR6m
xqqCxKD21jiD8baZ77DRtdxrlWGz3DxQUVnVlfrN6HVPPAVviSt2AWkCtaZ25j/hDttUoskTz5m8
NR8DXUzExAkp2tsE8LDIHYLFj9EbbiFFHdOnCPbhdX+fADTuKHnCeK9qwgL6fPO+iN3CYFK0PW3P
mEkFj9UoSJbsL8kODNH726rF06kTzs+qgGcVO4Zgo7K1/AzGJxQyJFQGnnCi8iIuh3eLv/ZuWu3W
KQlvCxh4ZNQKdKchMSxPRIrC0epFCQ1PFL3dK0Rvyd244IGtWfgF4HDG+NMMBIPaoFYwSvPFtW8R
bXlAZpxvqTbWM/NnZLktHuHO7ezQvwlZFJZeLiBzo3cZraSrqWYOG4PR++EAIebM2NbhSOxpa6vv
7lsmseqq+QU0IyaP05ib4TYMXJoyNeMspo/+TFzlnHXBWn3s9KtP6iGXlivJ1Ji17L4ORMzHNswo
vCCnaNWS5aJnvsCFXOkUhQ4T/+5gGsNhizPUEFSZiSXooZMilm+p8SmUANJKJwtb1usE32L1hNMv
QRKW5TkpkXqZ0k66WmaIOvyc+thY3mvXzgX8aoCDcWsBFy1o+KlBsplAVqRv36JOghmZ8s0PpL9O
OAt5Tm6P3jumNNEn+hxleCvPXn6B8ohZzX9432WcY3jr9hYuVJd6EsngYnjRGm8skfXUGAa2yp1P
1ZYKugbp37kaFcQEu9nYLPwJjwvaZo5wNnrdXAs5gbDLEbm0JmcB6/7wYCO5uS8E5q9ICn3Hd6+0
mi9NRSCT2EmfGVu2nAdzjb31t3c1XM9xpkSq9FW1+vhYa5P6QFRsKN4ZRbcntiGB/bMQF0tkKBs7
qKnyULPrNHnqxXFrka+P39pKMoq6Z3s015im9jZgs8MyAzAd3aMbGdKwRxSdFnsgj6JkUKS/PxVl
LcU9p/qoWL1ZK/IBPcB+6SA0wbGAvxDR22rz1SqQ5eyW1T/zFJ2TWwmi1I3Gi0e6I3JvzAIqwPrL
Iy++S/RL3ypF/MmJ/yn9Bx8KGi+550TUrp2RYZ45JZCxS7ETQfFeF+CXUJf0u/A3NRuGTR5wOTQR
PfdWyGukwUp9054Ts+I1pJq7WL2N7cltd27jFQFOhlG1Gfd51aLuRNNwWcstqNcpyLFZFQh/Df0p
gAXOjfo4PX16lIiJoUWnZAMLC5PWh6qhR5QVw26TRhUJF8DgHcrpGoBntZT15kKKCaslaEYPmPVB
fMPWzDZwRQdEY48nWnXJRFcngO/rpnj64mX1McW0wfaqApkael+5RtXO4NSJKTB3wtnFOC7kk5dK
VrAkqgGOuvOpUJEDXCYUHhAqByQive+C2ex0y+LAI6lUG8nMQRk/My4bq4bRxWnIzEhKhJs1LHYR
LGrZr2EWUFqt05eOx7o0t5ggqNhHNB8sK9DfQBnOALwwAQP5Ok7G5K7edLLBAgWgBbONyiF53fLc
nv0a9CEOOj1c63mm4811Db/cnWN1HVd8M1tkbkkjG4dilePm027lABmXYYhQ6qakgEwS/n0DDzia
kOq4P5HtsqCTIQA9gTXg22VkhYCof1sCcLzNrWPXQZb1Y3XOdbTf3ieEPVJdBdXJpFfz2iT49t00
Aruvt1CHTvPB4NE+SP/jPzy2dlV3GTmLUDk/W/XRF0C1ranZ9cWGgYaXyN9T8DdJerFZolKdtvLV
56aqI768K37aCLzE6MjzUdU7mxrDlHaFNEHIb7A56SPZqgHWgPw6Tti/tUn+ZIikcH2dhUa/FOHn
OCW43JHm1R8yqua5U5FSNKpI2TxNtBy0gc95MqmUb1mBHs2OITI9LO5a8OFUq6GZALrbdQ7+0B7p
rni5PUtBzDr3PlrB27Jy+CT6aus+HOzJVZ2w72lEQXt8rmV3R4BR8aDf8t9aeRS+19sEw1oKWy2x
ZXsQHZXwinbGv+p9rAoBlTkIulQws/xQKjLuzFv5c6Bo/frvLIUdsEEKFMP7jtfpGbJw9Y3AzcXD
81SZZoU2ngoTTDTsfi0NUINCDEcCjJkrZ9XV5JQZrzsTLIt9hR1MheaS+pyxC4uzUmSqYmxZGStt
rFsIhaOeZmrUknu9ePUJeGm8DdjwgUCobdEJGTNX3YuqKgCYfHswJLDe7nu3OfH/xLHTFF8mKVXk
NIpwRH1COyr+aY68V/yH4mRiM947JIy8ko3Dru268rJNsg347OTv4JjdSUA9TLUhT4w9ZRSPHUVg
0+FT+wTnJUReQI7ou2acHyreKSzuB+cadLH9R7esVjc38p0kkwNmFjoZ77ri6HHh9xag2VSiKbsW
Tx5E6LtTk4BsPkiFQLZQStA1JCRE6EsUxUfVezBzKUEBzfIBMLkVsystlEuI6bvV1IM3NGDfTliu
OxXA9EYsQ0Q5omytDtpoQri1Z/MRFubYwZXalD798OaCKI1DuQUEHwfGsEs4pR/xGPiBfHmNgR46
zNQ6aMtMbN50rOfmmFGd+cbYm50vORNvGw2ITrVxaFiz/erQwxa3v/RRSZ1m846vLFTVrwCFsXfD
tNYg50JOfE95jc4jh2rTzwc6e/8nMLTyoL/0D3IEcDxU3sUeTazGQ/WVeDHO6CFwmOSP1yXyLqwD
s5a3ebuwBSUyQcphpKDkjyeDpuu/Od6K6IbrI3KZs0q7vrvSJUs/V7LvxEto+mcTrjcOAOlOzaOB
kvbnTSzMBirwuD27rD2lQPNOnPa4w79zavk+CB5ti8S/WnIpUP4Cuyl87bKRTq3ZuyC6bKja+5Au
ICu5hngZWCaTxKlARJx2aWVfsRMG8tDY7AW2MjW8E5Jc5UiWMSeLZwx7N0H5Egh8kAYl/MLMCCtG
uSbdB0L2Nj+HihMvbWuL/AHryPfhSG2NGtxwf7CFgcZZ+OqzXSEhmKelxwlt6A+k8loXrsnZaY4R
soebnvdslOFAnspk9scaiJB4cwLoTHBtQ3fXzpbROVvT6WShwyNOMDqLHp+t9gGMshWJj9XyxHeb
ih4DxxqSWhjdo/eB0OoysdgeBKYhhRowlr1FIm6g8cFGfc5jmgW/lXVGxXUq0jL7iROgn9015xL+
L3AIkHT9x+ALo1av+IMJM3JrgrZVzKH8LnnwSjk2Aw72j35nN5aIxbwqtpBu0rtU5jlvezLvcYtY
QWALiUsLTnTOi834rUZ6NZJ89LYMU7I4xaqh5z9K1lYa07TGyqIRhyUzAvJauybPeduZdixREkTd
Y7wgKUhApEpZ1nUYZkyUF7tAUgvHVKlGdNTjkFEqOiuNSRNa0hUuYWlpEtLJFUVh+4DF2FcMuODL
UvkQNsg5KyY3fE0QxAxaZFQuFDcxDCbr1Iek1XIsXeoi1iZGFUqKKqwricDbc6VLsRLrpuqyhWEh
+AzuUTAIMw5h5K868M2M3VJ9sQ01BsrSydWQ2QDCkOB/GctIkMjNMnKhOxe8tPn0uSEnoYtF1SVj
nahf7WvjDft6xt1ZGb5XgwdGvw8+t87r0J8/vFETwQR0z/vxF5AZWL/QAMRzpeyStgbiKXwm0xsr
oEnXYf+tf+/jT7itWq8CnXpscAjWTqseeFjWfB0qGJt2uH8SM0fWVu4q/ILf7oqKGKvEd/2xC4R2
fdST8Wi56hDUQ5mvzEItmpI/xtc3hCiNpkKObmSKeFDt46lQPNr3cgEZZN8W7eWcgfZ1yhnbDPnP
03QIbPhqPV0P8f2GLVOhxgvjUh8wnunrZpIP8Dq/TCyw7WF4gVUx5sWJIeHB8W3GbQ44JqEK3Pe0
3JzaC3sOe7mxYa3N9ug4KJk4W0QAKoxqCmkG/CE++XmnddLhs+m0Lvt/3vqPvGF1hr93hGAg7Wct
2olcuFb22J4VYBChaKA/TPhTrMFyNcXH0cFArUFGTJSCn9UYNa6+JwNj0GQU0YjfUsnZzVubExrI
VpDl7Icq7Ty/1o967Z63i5mKpbKOGfBPwMSNSAgmDVtD0FUpm9IcPK3WDKp3JuiadTsBKchRL19y
SKP9ajyXyT3ujhFSQ0aFo6HCE9fWggX/IU4GoUcBlmxDIYbhTl6XXx0c/MU8A0vlE9F/KykrjarR
tJ6k4CkxxGBT75h5CICSjy1R5C6V4USLEM8BtGMN4amZHjS/KZQf1dyH5qqwMv+8jERncPpgeEYG
F7MV/FE/bCSb0Jn4UQ3LKYrbXhT2JWBiF/5GznlN3npf+lKmwy2U9Vy6LyrF/R72TseTs3o/Z40Z
PXA77zAedlIzRJAkMeIUB1Xh8Q6jINp2nvB13Y+mSk6ByJbDEhR0TNJwOZlG95r0njJuCdoQt+4B
r1sRoqou6vLVUdZSGxyLUzlsoQSaC72tSOWMewvq0a1eUZ8YEn3EKUmG8H3nGNORg3yUfBru1elF
ycl7WZPebKhss/8TgMFEdasiQF/6sEovia/Nmm9Dno+GghQGWjjN0XU+YZFn/haPTmWCb6jWO5pI
+xMQURBOhEPV1rspk0E1Hw5S+S0+y4dTABAeZl0e+wdxRsIpZZG3WXUEc27H0h4dt1cr2eK9vWbJ
usgEd2nQALVK+4+4f9pECVPMoyJggEt95bVp/c8KKtz5z6chpkX73OIs7OoSVOwwLBH5pvDWZVAC
TM+Q9dsZXcIDEyKAMWGLaR6T+Nvl/ebWyQcxjbFanK5g6HU0EVL8PUGFoORs65W89t94GJQw/wmX
vIgrrnZoJHz+vE0E9GSyyVY81nSPHo2y8G7iYyMu9dvv2ZI2o2EAlbzaTh0CwnRmcFCXPuvJJOQF
VU1de6RkoUzBOFJl+7qzveihuLFCOh5FEhPJLq0NXr+wJKz17Hu8sCBblbygs+7SPLVhlLtTP2kF
y+JjHq2A2eJp9py6h4hU/bgHr0wcNMCW+RoEycXDGy8Z7+Fzy3WN0zKhC0BuvSPK3smEHIxchFsr
cRQuH1C+284RgoVMGMR/3OTUCezeIPrKf0oCyHlR5bJe/thhxKlRw5R/jD1rqb9KB5xazPONFtbG
0UaO1dH65z/49FRtxZqY5UnfcVxp8XewKtJU4MemBFYQPy+mL6WD3exWh0lLdPcPH0WmF56jB/Xg
cu3oXXkmYiB3KZGq+tXcgtLxwVIs1UOonCicrTjyNHnFHkw8fC/EQ506lqDAaM3N9gk55dz4u+FJ
s1hEao/cM2dvmVq4q7WO3spP8PC9C0bkTqe5v5bcyt1ttaBnUmZs/AEIx1z3OgTaZdN+a/3hGBf/
u7vychrOJ+tedoOML+cEKpCslMQ0Iv7S3EJAxyH5RiZtU/5JkbY2w7SI6ly7FAA/SrOhCXYN2lqt
Ta+e1YfintQAMfHh+36GQl/PDwUzQXfe9dy3oCsK7nkjlvHLjxQxxgPuQ0UM58oqJwhfJbi2hUir
wEdWfmNYrLfdvLPNZQDSw8WMZYHXyVurpFQ2z9V/nl6t9IuHLLDMDkT1cOQmntXe2/OzOOHxGeeU
wQUaxzheRXe64B7HXAJ34xcSAs8yxYCTN1EGlm44OW+w7HAwVYAb17YHFn3xFnWL/DSOstawSQn5
RxnQrtzS+kujyrxcgTR3ci1LQwrLHsCBUyzdKltMPbhrVe7qm68tvrPNXX/EmKWJtxGMC2yhwamE
ctHVEYLDvwjCdxsaGRfFbQ/X+3m/z4g6VbMPnm/9EIR7MGhz2yIfYeuDbu/MOafp+onotTuzysZ1
wLufPmGJ7Sd+OgsGkrgFVr9GTrhFCmjMrDaU6nO6n9mUD9OW9oMYqnNxkqmekVfA2ryCF9oqiFuM
vleicdfwaOcYlvGIYb32eDkV3ZW74arCGopGXUApk5Oy5h4ueNtnMIv4PodvvCV1LMgXrOEA2N2O
jEZIx/0tjVs6llP+iFiRAaCB7hSB1ayKzagCwHkewMBTPTmJGYvXlA0j6tbeZdb1jC1qukWRLrtJ
mkE3iI//cAT5+vTFJrqrIP1FUigZUDRWNkT1CzJpgtlcgTW8Xzf3Aet8msFBFysSuTyWWAq/TzYe
kz9eeoy0HFurAWHGXVbEkPr57ip9AkG6UTMhhpEQQmW/c+DSHLJVT81KIQpdDVtxl/XbOFix0cmw
6HvvD9jNnQWQfZM2NBfeK3h7Oq8AR5oEF4fFvS/9lTpHeYB0uoC1hd34y6EIgkH8aX+VMjumiOPR
Yv+LZgk1ZGnbBUOTokwDvv5Gas8YxhmazAGx2ROx69XdUji310tiEpZKQMT9jP7JKtPQnA5fTgqu
E8L0FUkKaLCjLWekFBzA6Bl9NNP08LgrKXUvf9wRV/TCNBBvJZJ3AxRl03b8pfIF05sNvlsCi3Ls
omDaqJvxnnlHUWBwuQBQZ0apMFaeamRsGksEQHEHso/O1m4FQ9z9eW5cSzlUjXUxH1iWAWlhRuAY
OKYTXTFThRhKx/z0bEdne8Sahj2lAPE73b+C4vLG2e9EYfyH2HF4RjbNeE9fB6jc0wIyGIFBGvTA
DY2UkyXi2ZnNzdDOdI12LaN+baLuSrl0WOqBlkJ3PYiujHYxzHOxtwosMav2sqI26h1StkwSbDsU
/N04wfhlz1hPtMbQbdoB1L5/9IoO4rETpXGfdYqP00nSI/fuGToCPUYyNHoXTTh5d9FL12/wdc9Z
8tNgMUvbsxdisi9jjusYiUYEQlwh2MTMIDvvlYcC3Pzx28zg9P4lhqfP0c8klPENa9NizbCjThE7
fwQc+wz2gMA7O6qRKXqgqmQvXuYCFbdE2V4N0ug8YyYtRZcx95snhOsfqltwJQhat3RfV2DPxumm
kSdYhGhitQoSsdjHZIBZeFIpuQgtzbnIyN+VFxj+02Lsf84wOhZxzqdjy+1BIoyzh/1JpY7epmkX
ygxjqfq/xP1W5RHOI+jUGQuAlOWczZzua1mdRZ5/akgrQh7/VZLThR4Sh0k92iNcVs+bXnxugTKq
KPGQK9VbXp1z+PYpLLglsaeAmLYRslNv5bEkQTG7yCfXAV/0EC0A7Y95UKnjHoze5ee5LXA5FzLN
B5HXMDl4fXI/aE5hvUZoQGfjdaAX/Y2lRLFf56vEz2mpxRohavsfSmahydz49F0wVjQAgEek9nzb
/v9AG5U5EgJ/AgJKZkBix6yr++EL9mSoOhW6IP6zCShY4T+IgrqQc0Vqrw249fWi+Y1OIggxvr+6
f20hWVaFPdBlGMJbpiKkvc0SVZD9UZ+yBoYEo3t5UZ6+ZJIU29N6BvMTZ7k+jRjAWIcvbrVl/XMi
NUmSzmKOSLpo3CTkHNTpXBAOsFNMyT9nOfO3pwNS63nMHLNFmtGqbETKmkOMIw8ci7Th3QCckYhr
6nitFNigBXPyDhDQy13DzWWDvnHH3+be34uzhfuuTtUYGetA150pPMawH29xGPLih7j8EDl6wYlE
JcFfHFQY6A0HIhNB5pWdQA0kt7pv9FhvtWa7eYFZfseQumM4lA62x6kQFzELFYETkEDFr4/D7SOp
HS0freTyRxO5weHEq31S7ZExUqrl8HxjqNiKVMtq54kLIjdL7Z5cdvcmROutjM7qX0PiWs75ZbCr
NsUfYCHypBOvrPuGGZZ2dI+3CnJ/GKDF5QPfiPIHpdDWtjYKZiAdswfP6b1uyIXLQJKHMjpQcoOt
GeutdyR0vRMX9OI9R5kaZ+qXW5Ib4RRqo3TZqCotNEFHnErg7mYCHlFvT6tfrubIyOGoOtD4oeDH
CJzJZ285+tbPGTfN+Us0Ov4KjJtu3HGqNA0s8bDTOND1V8ZZZKnDcywdAUyNIhUdVCZoIq0QYjQu
bbcVKGtG5nUk4mvtKUguxHrz/yd7WdY0svT93KMrd0H6bhazy0XDmbvUFTEil+xrykn20bWaSa7U
ALzG1xMvT7TFy6KTz4jCMCVRTrgtjQyNLspIIBkXKc03t/GCl7a+HcGOweHBlkQEPLPy1K1tfL+G
UCO6zxSSRF6EaxYfQDvPrcjNgJcoodHY5cU7jNzJj8rj2x7QIW7CNjpwxbTN7y7vIHUrB54o+lZ7
MIQOIYIOLeuQgAqFMksjW2Un4iS4rZKv6m2E/Gs1X0SFvEjU18dj27xey5m2PKOuyf4D6OQIGVLE
Kp9T0xwIlMXOznBibTpzUVD8x8f7C1+9fAH8Z7QsQuWCBOZnMSHiKnIakPdUNeRhE4fs0+IJN3Qe
9K0cY+hD6Wqt93TLID/eEbyEWZRq1TRyJnjrZn9JrsvGE+zucq2+vqgRLwor7k6iml5P9F/3EMhT
WVG9HPxveVg7SFxqT2m85ajso2a7QCk9aXxTfVYTYNW140CKLiIsQFsMFSslD+8PfsdM7Iq7VzTP
rLVrFDQIS4qM28YnN2K9lqYpz9Uh2MRtwXnx71ymJOXgeynmJJCngtwf779sjN+Cu+L1qhoHK6nd
/7OXFLPG8am5kEr33Uyxd99UtpJgiE8ohjM8JIQjd8+SmAC0SqTH8b0ydygEiLzokSVwWlCJKOp5
50d3Aw0IP1TKKk7C+divsycpU64rniNXqLrWSkP/ZgUJoqCAJezmx19xqp/gmxOrBd2eaN2eQpem
wM77tDr+YVJ/wxlweixPnuOnAIajACDHVS800p3hGEdQeNmmvTUOdTCGBrFLFPrSk2XV5XVMR2Qb
YkO03qjNapIGciCm5TC+HiPr8qfcB6NkjK2jlq37pzLm7yamSfG/Gh3Vkd1hKY6eJ09cH6WK3za7
ecmDChGPRXY5Ci0rMg2GiHmbaoz+ZwQgw3shy2hXh9F8cKEDfHJJ5Zfa3CvNpke2DmZ6RX30LI6+
AG1HBdbOyn329mCqYDn4v0oxAUwVupqFYNDTqrMr0UaBWNVLcXb/Jg4ZdSN00rtjVwJ89AKH9tFo
JKyh0fIWVMlqz5lgONRHFTMHQw6pGqB0bxZPcUVGpWTTpgMaU3LoNR/bceRkLr/RPJsnx5In0kUV
TkukDAaYh2cEMihugn46q64fhq+JJKZBccpmoafLvPOV9I3lrdUnX9c3kRyK7gkDUefozrn81XKN
0Nk5NXivka1DZGXln26pijuQkTvY4r5VvSzhlBLaWzyZCu7GKv5g+cK2L95m3bBTneC4j92xMX2H
A7VOrVwCvMPKCJ+d7h5HESSHygUhyBWkIgUcT72f75pGoR3nHSms8v4HItvYwmVUQOT1kANIymNv
+K4rd6sNe5eE4Q91EeEmu4lPFqUvXyWm8qUxt39pZTrgKxmGEWF1Qd19JaJ0Cd9gMVoHNM6qli+Z
qgSKmUaXoLv3QyjOlO7hJvCHCe2Z1Q2o3zjYFK/tmAnxET8UIDSilFvsD36kKeTKUPKI6SLfsqSs
ixKxCQXeoq/GFzu5S0CzspcXFwdjD2FErokKKlb+NEdzmokbIbSGp8cd+3pYXs+7il8u5SFZeBYt
aI8zE7rwBXj0jyowDfEq6oRqkdTmc1h4c/vYldi2QzIcJ269E+unFVBqtLPSX5+nExOUYZehq5CI
R8qrAf+J291uZvqpPNOVVnpt9i2RoqgY0cnqaubna24pH6Hmm+lcnj7PYN59rT5CdYVWms3czYoc
GbsYbJVRUUUOu7ESmFuYQ+9iErhQW/GTXmI9RQESOVbNoHxHEL+BI6A5t6IGcU9+1FVBX368KvXp
oqSJfgtYan361MZjlTE7kIAZlIpP2jI/wya7bCZpcATswAMcLZreiG+FwmSMR/7qDSIqF21vfCau
jBpWpklRZZWTTpCAtFDeU0fhVOdhaDnUL3LaAANVa3xmT0vSY+LPBI7/XMc+UGZ35rLUm6SwJ9kq
c9dRLTzjVlGqwpSfrQk48/ci2cFaf872APdFfEVn52UOF0QxxOEXR2xHzmDsFmec6cf23Kw95VMY
myxMMyNCr6nAKBoDfbfzc+u9Wo17Ihae/YkQYt/5ZUleaK8j9qXSGJetDwGsib+nCqw1d327/Nc9
zjoxf/FShz1f0wiu/SRvvPQ92FV6NpgDKm45D9pB6OWNR3q5T7j9trrzmCCEaswQPiAUExbNIlYv
ixu7qQHpssGB4JKZduDQsxYTnvQ5wAoRUqq9WAsUqm74orADOnytVqYTwoupwTgevoVIbtpIK0za
UEaP8tonySFoKrzJHfivIj7buJgx/MnoXhvdpB0qeFbdhUf3BwZMZ4691P/3y74aSSXFicihpMXv
1B/tvmPrVe0Dc+xSU1xgswTXd+HfutjpElJPwuzzDaPOVDtd2SwpsmbWQKE51BXigfUwQSEYbZhs
SYLiXP90UxpQKPDLyuX5vC8nTjxf/ZSoFIIB7SKXKBcqJnYm4ABqV45f62GPVm1Q2B9kfx2GnuMC
LJctfq9BepcswNIQQclelg8/1ESSJHVr65XyQuD3SXDOQg9pmnlpcxp7kiT6NvgvOhiLncLdPZT1
ORSwORkpAdDe4aOqu3WHFVvJm2uohvutly2yJgMT5Rm972oVrqK2+vHiE1UcOdyyf8K+ZzOaLdE/
WpIf1nDgPAyQKp3SQS8hlx1Bx72Nj+cyjxiC4qwBPTAeq7UCw9VOpZFTwpoIYCYet7qnqZkaRTzT
j1e51dt3D1hsrksmxmr+F1Re7VS3NX3j7fAZG79+RoI/v/s91FsVvB7Pjd83ej+gz3R69qTtQmQM
WzqzczSW7MspjAvG1z3yYS5DPgUS1IMsjLBFm5zZ8vu8JBaUjUpH8nRd+8mLep+XbenWKNaEBFFW
lNFHdmH3otjcoxwsk4J6/XsOcF/vAdAQVE6AknbZt6aNOPyBxNxHWSxf9KNC0K7UYbH22uydEv8v
yzIz2R9NQZuRFioGfuuXkub2esG4MySADq92XS6EnXXIgId7osR+yGQwZqlGpmAMzbAQQ+7HW5wO
E6AoiT1M1B6sGeTBAny5P6A+jziR8AnNCL9j0L0KSssNws1C/bpOitqKV04YMfgnArTMalBP/V/I
gM2XbgU/fZMbbAlYah7+Mw5WtVeF9aCRSI5a8sWqIe4/fmh+yKv5fMtPrkIbfyMJH+My06LeFhDg
ivk9tqFz63wCjn+PbHi/renpg9MnjIHEDlZiY/jwN41OG53O1trUOh7aog9kvp5goxercIcEAwQZ
BrzZISAXEFW4JFiseDyO6vaGekL990ptWY1GvBQIEg04gLSb+YgBQijU/LWs7HH5XjgqbPg+YnDH
mK8KB5vfv1e97ONA8Adk+jzXgIr2CY+vBnC4IZ7wg+z9qXT7UNXSruC+y8j3dJG2vP22lRPTqr2z
eUFCA3UdqawyozncW/7lzxrIDucv2kl3frHLhNaJPwou62JzlfIQ/9pzx+FmhrokVahamS07cOTk
azUptiXk33uMOOPJK8/B2m7cxYMErUS2YHF8RgXTOLQ/0pO2mNUcp+jFd6Q+Pfobv9sIbKjMssnk
QNo2AE/daZwHd1ClqUiwgQ/NznW0aZYBNAXa0981Jyc8D5IaNKSgnPydcHMMWxTwfTvU4qO0nl3/
A4nuvgWuT96+efho1saNTqdI+EjbWvuHvvj/rP8dDhuPEKiiokFifSus8jEt2HQ8xpt27ntbP4PA
g5Da1hZyj5h+Hgx8ORECEkpMgmSQEcWIg8IrH7K633C/Z95tzVu7/Xv3lGpZbsVa1Kna9SliXQ9B
oUz2dgUwJOcnAOrNwYSZBxeAvOj+RCuXTSm5BYrDzplYxJLRmo8lo3mBCn4vpVICboNDzcCoHBMA
GtE5C7hT8uc305g2jFfF6nNLwb0A6ZpU9wjUA4gm8nHkYG0nlj4CTcXBjk7l8dvga0LM7tNaeogw
INnCLQw5wTefm1eymQw1SXKcGQt8QRMNTR2i7NxrTgpXwJQAeKNd9bcwdRnz38OENTQ6Gsuh0I2U
gCKpwX7+T04RSHRNFboof1sA8GyeCbaYDY6aGtqTSLs5FXAotYyz9t2XRlGF4LYNqeOKDBjPAWLD
E1ZUcGGSS3WeMe5QW1ZV+1VKD6WdeVrmDSTa3wUU8jp7hefAdZ3ZntsaSuZReZkd3SmD598zy8hu
PgjF1FkqfwLe2F09ObI3B1tvOY7jUjs0M1VwRQ2VeDyYGTWXX+aMbUsCOQfXS9xBdz+5ADDhGAug
r+IPFLOeFAnV7yRM++6/TX5gv8yzDdIBc7PUNPshmmPfXmsi9AIqIFPI37Xs3DkDm2vQEB+hKr9u
rsxEri6qd7m4gSh9p4VaXTia0Q8RqKRZ3NRTmylcLlCg737hj7uRxkgsibkT5MGoHKn/PG3fyria
Gh/Lblc2XQ6azd3cTz0z3L5SZG3PwGS9U4YQ+2M3l1isY8jzJ8ra4JCZ/WS3FAGx+IXv+MMmHaug
EmxRR55JldBnGTYpc+SqR/NKbjHlBxCjbUKU2GVd4CTylAK8fwAwvmdI4z66L2jrpau/0+7goK+8
1izqEc55Jy4TsrokrX7V5mXb/c78pfTzd1EmC29g1BVRcc1B9cyFMidP5UHW5NPge/pSIVZ5rOyf
fxBJMzWtr938gQAK8ElfaGeuXXWP3Mconkcx9Bifunywsoca+ZL+yLPuWRr2E03zsrpF1oqjLLzX
Y81GCkAxAGstMO+CWL0CgiSHa8SYyndqd1hA+vuXQ/OJ29hBfhVCDs8JHp1dOrWFMOLTZkkaI533
b77KN75za8J6hLm1+7fzUYvPavpf9GqRlT3jhhGPFBVKCltj8ZwL3+jf/byo74emFcG1ZOcJyXpB
MJyUeOJvBWDCa/K921Yox9h8lUcOrn/QaSeO7MByP0zgbi/Nly4xfLqtSZ4An4XqNWt9DWN7sGXh
O+vQqKILYRrvpdSbjaokXFCgsaBfUGEgqKtZpQl0sAida0wc1Si/6u8p6CmbWgOrdR9ZGS1ZzfDG
9PGQ+v8OwEsY8furstNC+gz3xZfa2SNzrc5vBSgLdJHkcHDALdutCxOc2oEX3hcRQZIUNNsMlXRE
zprBBFr2Pz2qaNav1PYrWgpFG0VHLLKH5nIo1OHBfxa0b75oVSDxu0VFaozbi1//7Vbsr0JlTfqr
/EuNTKeRmGEJ1s/+lB80AlJKdkeDOFcA0FIfNnm3rsEjLHxkOc/I8DTo7PYnGDNvUEEGaP8y0Iln
1ucKXw7+g3beYxpd2Bsn8uJ2+VJzKBo1pTCdRtmYvISP39hmMh25ZHtuh8521nnVvDh/0LGOUcXn
r34Jseld9U0C7HhJT+eU5AT9Cr9RrogsccmKIOpqhAOAH0S5ObxxBwhHKwpno+Fb4oTXWTgVjQDN
JCdEImVqTjVmGJMXqLXbKSaTEUaFEBSDXQHEjXHOcl4oSasgGhs96YTuAglXnF84HCgXEnMZmqGw
EG/TrLP4zjx7hGjAdm6gxR/VU07ZIYK9bDrw5KJmPQf7d4okCwZcPrC3IQP6FWUijkl4zP2X2c7x
8i81CuHmQPJ/ha3VUNFqFxF+rhacO4zLMmdlIcfUBGhNK1lMb4FslKeESEujPGrb/HjA+q2xRPUz
BYvVyAxEFy0gW0h/3xiiRXpaPb0DUg/Jdvg2LRtC3NC87Habf0knKGn7kad9kdVXtX0qMm2QIh4G
ZsKCK+bbRkMNH2V8C7E9wbtbl/xDXnLGK5qR0XqSTyvmScdM2P/9RF+sO99GIO2qD0NQP3RvMDTD
KPHW8YxaWHJde+WVRG0rxs7gFThbkEECgiMddaKIGu6Do8PwhQVoYQGQd29qbEJ7vYd4No8Br6gU
dzhbwz6DIRx+fOKNfKRnMpi6fNEhDuYvg8x6kq/YSXVtPmqlwi5vmekm5I4sfVZVWJu1NPL+CGFT
vutYK6QVe7ElcSK6WWNJh5yjQ3NHEjueK9x8ZGpoyavIB86/shNBw+ebBLhy8fH1viXfhF6TXEy9
Hk0kLmVnUNHOzCeN6eRQ1pgw/V7RV576kIkwLLu4q9ZQQc4yW62u7zP1wY+X7KszWmOwnTDdLE6I
odfZ3CHqtkAvODJQ+zjeOGxcMUDYnA3LdStN6Fg/DCOMUJJSQViaQE0ysw6JJ3k6sc2V/CKDa+EE
Ef2FL9MqPSv/4aMmCNPUOmAUNka9pC5OOhl+OK1acA+nNnWEETIGxYAcRs1wMvV/OC4rQNC4kA5A
Bn5PUAeQz9xxt2wZnZayob0CjO3JhtOHdoXRqq/xvZmMNlky2IcsvIwUYnVSGJmyigFfwlU1Nb6C
KB0r9GAPg3CuPd02m3E73zppBdawcJJs1th3IladHoK6z95NKY98B54TfhXlVZIYmCLFlKbstWsB
ABDoJc52vWZcO3CW9Dkm2RJ0hGt2gMlj9B31/AbvX+Ixw1Nxd4fDtbtXrbwmofynqBjUQ5bxEb/u
CRXZ0N9ETOyZPg1k5LrOpRsD8l0PCfJDcMgykstgr/QsXXs9Z4/ApjiUn9GQBwFOAHPJyIRvv/3S
zlTFrBKq4YaoijJST6X9qXlo+D/Hgdh6jkgvMr8Nyd0A4VHRE/HhOcilPhJEA5KFJriDwoQAaYN6
Tb1smf+Dr8/Q3cOA1MPdEpSFvG0ls78wtbBb/ZmS8soM07vbvMr4XTxabpFya13gUYfXZjW2zVhW
7fhU3Wm8bX2CRtZalzrePGhQx87hOU4n8t6XqLVzYILxmYhjecO6xKvHNBbPZ566S9qgZxHy3Ks/
K6NyTxJgNHrRRClsyABYqnpAa1XIOGx7UoBfZ+N9lgvloknTA1es0e1KBMrM/Vp1JdFEGlN+3xUB
wfgm04PvLgaUvNstA6LmTCo3+kl3MRpypwy2Ewe8xRGWs3S2yNcx+OlO9eHhTaxKCTDx+/3ftOPc
Ooh70gAmLmLsxEtCHnQo2Gyq1jyNnJeGTI1ihPwZmGm8j/8n0r7qC7+Ne9TDy7AAijPwSwbWD9Jx
KXHtQQ18Keof1B6mvhiRq03Z6fn7IHnD4kD8lenOnRfTHZfzT1vjx4yzIX1Z7UXRnZiBoQLWkNbV
9cjuISLedL3XmAZHsIUdQjBx+KDTJZKD47/WdjhC/cJlX1d3ldG9bv/jYxfSVz8geNIcUhi/KRtT
1pVzl9gyHHwmmAQFDcxJP0C2uWaEeIoLuPXJQA/k8Iaf/6aN5FbmtpUXNuXXxeVcka9l/uf9zSNQ
dTPATGLaWPLbAbri+VJwMg2GyBFDbDYBsPVF7ORRNY/bPXwrMpBqYgEIchYaJTpdFNT1alKtDs/l
7Vckxt0WzfRcL+vwrdaVjYOTHRA3dErZL3JDx6AKj5yle2wSYKcEd2FOURAPJ1mURmNi7w5XARnS
4I8THpWYtRsEgvnyQv7avwh8Qhallp95MNWB5kYAqYLsPSoSPzEbyoy7U2GmXQ5dJImPDtRrFtY8
MwhlYujRDXkMDoSK48XaU7aPrVQ7kKUpOxV53ZhCPVsKIfElY+uQujFmt6JjSiGv2OzgZXy8hLpS
W9ZeOealv4a9WTiZRxCZmbal9VikEDmRmly2pCLDQjrNecwbh5L7vtJftcRovP0WQ3e0GnuDj/qO
utp/FgU4Xn/D+gxacdAWEXFJNTCmmRKGsPFonpzVDt25YosIN8oVO22n8M8q9V/p5Te//7ZW80JU
ckXhpyHj1GUNJ/1d0UNg3yyTOIBhOBk38anE2qo1CHLl55hR5iKFYWYma4O3MQxoTC4klxV2QHNC
0i0Ind0xmET0bQwD7ZuBw0nQ3IFq5st6J+KVEkLrj/IbxdhgXrEfvpqYufvYL8SMdmTNubsHAnzK
ZIeeW99lBmSuOLtLXYwnwQpQV7QX4/OhOZhOCO9M2R20vRiSsgZmeCCFp36FYM3Aq2Odya9j6eE1
Z/eFUgHU4nly6fwrYTjWdDls2YxJk/Q3C6MG7Z1YJTK3j1kEaaHqgk0CpS79EUik6KRzUcLifGIr
o9M9uAIbDuALbt/Cqln+NaAGdDJepGs+eirLQXsypbMW56HKHTUSMh+64nKV1wRRO0OlT4vDw8Xx
fo32Q6qgmC6wZGNDMNDis13vOcvr+qKoY1lwhnUeOVzSuyilM5rjA70Ev/bMhS34rjY7Xq1K0bNr
95rRj14aJNeRXkPBVnzYJIJZtetSgDvEh1KpZ954VoIwhxsbAfGSbfwK6LCwgeU/OlXtLasGUsqT
FJDvaWUpShBJvSJLW3o4dcYUzon8cMp9wr3KtzczNEBz6Iiaen9iehT0pt+JT9ucqB42ZR+jDYvI
lmss589X8ENAdMzZITXSAmeZ2Yl/cZS/i5EVHWIRtEQl0bSNEK11+9lL76d1/W7L6OInR3oCNeLa
qUb72CMsn4PW8Kxu6hrGcH6VmC4y5GyOIBWpOIsvmKXHqXhD9UgppKvTeZYuGoBtRJcPuNiwdvpJ
baKzrR/+0T3lTgiVM/prCKMl/GaLh2bmt/4msXLsFpoWSmT2JMYoypQbx1s3v0SmP7CFyZKeT93o
2pr1lLYDE+asOPICaXjVxazgrESfKm2kVnrHWCc7Rj4tz60Dkc18b5kTYmp3C2UiVpRanuq0A2hD
rr5PPsS68WjreVoYnWzVA2Pfcp3UeUMyW/oI6LxsOZmbAj78TicvNlGC9M0ycqo2cOkuE9lk1Bj5
koqCe0k47HL64Go0DGCLbUDuIgTHhVrmU8m1qsdyR1zZjxQrUgyamM7nuLGU25cXPKY6TVbzbtcc
69jEV4T7M3ZTAyiuDKRnNAR/TTwj+YPSQ2kEGRXchtEghMXwFGA8mWLsv+jPzazjYk6LImILuLaD
Lkng4aXY3Jlu/4FkLX2W3cm8gMKqzHt+1gkcxMIzJM2QMQBIF12816Ur7ZAf/A8nz0ymi29ohEDQ
xYzBp77cYgGwHBPFsqtumPmHsPGuPK7URjXMCcpNHt+ijtGI1B81lDhjGYamoAIp8KU1gEUCpBNg
Qb77HusQ9i023ilZOiPllUe4MSemeDV3IN3TjIogs69UlXoS71SIP00trLWoPZIC4E9QwpdVc5J9
LAbgee9YW+dDYc5aSBX70hldF4J7RftKQ3cgltZHascbKzF+C7xysQWAYvPwJ5J00mRNdtUZnhZ/
XTou11V6OT8TBuTFvVZrFOwZHgwF/sTR+0tTFintvHXwfV9jSBORtsfyb2I34MuX96jxYOXDoZrP
QqwIqJ4Ijov0quBQIHSAhuIJDRqOHHWP6o6n/UcCdpsX9An6GGClT170yV3ftwN9fgBpV5FBkoTk
158HHMNdYvJYJhIG7o7HLxmNxG9bbSL36TkyG/XW0pVfl8PsKs6wor1y5E+YeyGGrm7icvTp3ZTD
OrjNqFGJ4zUh+J+QdIBHTVtUFNY096ASEOqcqwdITRnCK7YhMWZk4m6129akguiez1cS7O7K32IJ
uxpB86aQXE9LiRqBFnlMG/wHYRFG4Z4gwlj7gk9oH9L4UViW39Z/iPOeC7DqOo0U04yaNBmGdf0+
0WswrW0nxTl/K+71DzxcYKDFu8LW3Dj/xDBdesaRJxix/Di2MNEJc3GAjZ6szTsP1xY8UTaGkREf
m94jyAgg0YR5G/GuudsYf33scapzfJ5WuiFQmU2f7mQ0YMB2gTTaUdF7RFOgJLuygvpI3RxAImh5
iuTUT4KACaeOmucN+nvsd0DG6Xhguo3BesrcUkJrqO7m+afhg6E/rVfWwBlgMhhHgh+BSJOJhrAE
lvxdywyUbgbKlHfsRVDRORc3W1wXi0fKE+tiNiCEAUEFHf88ndJUx4RasYtmSWomj7nfJVllBipb
3hd6GLaSyW2Rmkcw+RnoZsiZlMPhQhu5N3jPetElpPcn2cC+re0LDZxt6qlan28WGzFkMpSRT2NL
Ek19gqUtBULdYxAJ0YWHpAxpMGBKIPpbc4ipwC0ZP2Y9xy/KWhY8ZiCYgV04vnQMJq2QB+olBvfY
UpYcTWj62hBb6LiayIUBOHhpm/45ZkHjlc0zE1Pvcp6IFA0oZyKjOsbz7kqolvIkZk068Hsp3SYE
ZS9L4iHCWYHgr5kom3CZ1BGVPslRy1gck2FcevFC/OUyBl3XyYGuzAZL9/16tKM9bpVaAZWbwtP4
CSToU/gMDFHjNaj9xza1mdFqswd3dTS2d1KmgBZCVT517/sXCVoACDOkQeSDitCMv4WtUBwrvkTI
+8G/+IbgR4iPPd6F/1zrB0S4cX45bNAmg5oG0NvIuq/5fAh1+w6QCV0pw6Pk5Ib7dgksIOegN5xB
0Br2nfpfwZrHJmkVH6Omc78Lm4z1ffzJQTdHKcg9Ngxh7KbFnYKLsLnZRLDuUvYztpVqyHJd7pY+
awgcIjJ0vjjxR2/VryjDH3/8VlPDlsUCjPchvYrAXDxnmCHRcOfUmYGF2Jt8h4tdWq9CFYrnoIQC
PWZpHsT2s0doBD9FD7VHqUP3ys+IdghJDuRFx15kuq9De87s/XzhapV5UKmTPXlwaNe/YJMM5cSD
MDTZUY1r3vbqIVrEAw7OS+GDRm2FcLD3PeY59Q8MXommw9YNWbGPoY3wIlxO0hc3wWfvzhiXaGOo
0dpy319yQgdDiQIa0ZXLjBQHnlHJO2lJe68BMRh+iVdIZbBuW3uLqsiYDkyakSGesVsfnop+ORPJ
19BIvVTfDIH2FBlykKpXpwR2v/JD18noESlgZ7iVP266OXS+0VLqW4g/nFajZbYhE06+d4OWOTjw
6kRlrUQ45hGMThm9jRzPZ+l7BhAtZefQiYKFssLgT85wVwMlG6alZoplFjZY3uGdyn6uRCIfbs1h
Cy+d37E+ORdiNSlKLXaUla6eJTgoQFdoEKSJhINRITarfujDmFSXAXQpfvAXkwupxTfPk43D6gv7
oWVDbCzAvt97K+t0c/GbXF96y1Tia3rwwY48CpkA+45RdgApQ2AVQFvVyx9vkpsROCT/pOMYsVkC
JB7f3ipXgf9xtvLkvS/aJvi+0OFFicORRDJtk4Ag/HOI5c4H9UfOp4S3NjhHk5ugFYbae5VcKC5U
rqPzZT2XMmvta376vSdf2RnZq0q2yGAPN8FzBtxGsCWnW/VFk2YzEOHRJit5vH3jp0fsJu1nTg1B
l31RvqoHzWObr7dM95Krj3C5qOutg3vcaQV8zX56+gmQayL6ikK409MKWO0pv4BOzt4tbQ6Zzosm
ZjASzaJacBGPXufHa+rkm2JRP/Qjnz9bmHFg6F7d0obdYVtc827qmT4My8YIfIXsX9apZnmNf1vQ
9DXx0iONTNNVuvq2oJOUQ8zBOdD+RyRwKu03nUnflWupBgnHxYAgKNfsH3ZHuSBMyCogOOVSPu+q
PjfgPYbsDakVGOIz2BG4yJEYhEW16+J1Cqgfqh3caZLWePESa6o6Q98xFE91KYI0YDTOTh3rj7eE
9zrGW4rogeK7ulTxNy2WrDQHbI/FHrBIUWj/z1CifQwwMpEs9oZbvvKg+80s4YSDUceptiN1mmLU
V91zWb0ELh9uK9whu3CJwMiROrtG4SKqr5rAIp572Cv9hEiWXnM6HheOqadfmAALhcahdB5Z6kOR
OdCGsnPd0UzWifsRTAVGvyq98hrjERhEJwf5VeS4sRdA4MNUKkCR39PXH7GnnJQsJwG5Zjff5NsF
+ZKzSQFtwt5ZrVVGFFdoa295JnyZ+Nm6v3Uce7nHs6E8n2aYAXzRCRW+cT7/RmkTJFdGDrs6V0s/
vHDOPxKb2cEKzAVXoIoIhF4lVGBEMgkWtd1ETsVxBgs3zuH1qe+aj38EaJS+tVaQI3n1t/BSx27J
eYRc84n3DWCjmK3D6mHpobhkRA6C2PmhtaL2EZCINVlPEdNiFGFpf5jPaDVDzClsU2G6X4Bt2ngc
lB19QLaqSytBg1d87WobOhflOEVkvki1bDz8mXabD+Yfr7PgHzB7/GR3oYf/KIgjeg1HYExjORUG
oIjs6ppGcj1niHKfs8Fhd0XFJIBzaWl4sLN1GhcOkq6PikI8vfURL8d2Qr+JSA+l7ApiOYTHwc4X
L5yDvHr+Wi/TwVga2GtvYUsn9Y7P3n+HDgiOr2aF9Zd9UgV8FZCYu6igK+LwL9/DTRgulFIFcL/2
ydtc1NTpzvFHEcqTMZ5vnnhIQr+Fw6zBtNTk4qFf79P+Q43BSnJG41xEhUM/Thwkbw4b6eViwei0
6U/JoX5Dxch1DXiz3icRfNYhgKK6ooah9aeqBPEq9l1kQLJ+KCG8f/mLYqONCZcst8PHdT/WaiUd
exLjp54I/AnvYUIBBUb60/CrBuehbZnIySrRmReqV6ty4CIYOvi89D6ZM21qXSZg1mbZrZm+/w1h
nI8jEoWymeistg5mZhQpTGHNZPvB7yAYYQZHeLpIZnxPd2HTQswUzYOIw/nQJPwNjKQ9u2iUMyCZ
pkLIcRyq5nEX5C6J+ONnPxAyoCaxhROc6iGsDnznRgooD+eDRltURQUyVN/M2PWLPTqIqn+co4Os
TQkOp51ow4IUxBJAuTO9XocXE6/4IwnPl1rN9g4fBdFPywnMsB49Bj6w3wtqA1+jfcYQuTv+/2RA
D1h9yVAW6+lblVCvd+7UPvmvFc84dwAp3cmQ4BEBaSfAytQHuzekiKar6TjzLpOlWeKMYWWBI4A9
jp4vPq4ZgZEOXecq8S/iWCgARLq4U9lnFAPqEiLN9+4o5gi7LrcfXxLItxypXrakTporLpcXkPJ8
zW+u2pPnj4RC0cS5VcteTWTRveAI3awe1Dd5IwPQmDbWZNP1HILlRD/7GfUvGs28nBXcorQglrCu
6jsHmgL6cqNIlPZFUmaJ68TwKuFjTbG4kBkoMH1xdsmxr9+7lItWPEXp98nr/sWkKWXzbTFBgVpt
gYMBxmV7zdckDswHliUo6A+8wl3wYgjFhZJIpdxlKiZ6ZeUu/jFIn+r2jbzP56umuYtDOkf2zvRA
tdtAM4KxoIBbhy1EHkdURxzJtqNUXl1F1oKM4gXQDEG2ZSvQ3IZCDji/UTAq0YtwIbSDZprjy9FK
mehbaAASvcEl7iaNJloqZ4CCSF/v6B0ZmW9dMZIfNUKIWUdufcx6KSwbHbBUTJ8vVScKA/7A9oa6
sPdrgPH32RohV4VS8USvx1GW0/wXC4o6KO3j9U5fipPFcvExGRrCnPDT+M1gbCrmp2Id2fYkbvsD
beRh9vEU7UCqaQHBp+/2xwJf9P0vUG2gcWVzN/xVtev1KNCHAJLsiQXvRPIF2ZUR5cVjj11nqQtE
HW7mH9iEFht74dZR2vg3mEnafpquwwz3ZiuGLGHDbktI1Sgcx0MY+c8Gb1lxzW7HIr/Mc4L1vdBD
eq5GNngkT/MDm/r3rmkgX3NDJndZKOpHnPjX1OIZHvQ2zE/dseAHRr8iwUPZHu2an9wFs4Pv+InG
JLchqdZddCsK0zsA9wWZ75vggU3lVQFB/LXWhYnyEVVwA4VSCHp17u21lm/gQAhQl3XCGywsxxP8
FCPL6bdkEObz/oB4sUYmSEvAwGguj1PAL8laU/IoADZBecjr3xfRjrMjGTiDVQT5Xs3EZ0/UO4sE
cEkoJcIDl1LI4AzHauvHdTvibpi2gBPcLQ4sW+tEY5SHR9zPgoGxgU41euYwZ5vht96RTlqRUt7L
3GZdTzuntMouIORHp174H+7q/CnCOWTzQFP/La6sWqf4HDYI7ehXd02msKW1/O9kh9I607ATCTe5
5+zROH1yd4qmBmkCJoKepEzWFaxSfHURwB9Ym6aqyh7qU/zCppwkjbN1BkyJbpmKP5Uj9wy/aQFI
aH6jyxNSFVvUIXLKKat05/vnvScxGcziN1b2vghrJPvo8aMzNw9KpamL6PLPsNFnkufBIe/nNlt/
GI6aDN1ODNFjCzBllUt4FZxopCEjNu+dW3idO9Mz755uuSLlPBPko8oRde9frAIXvB70sMt85xf5
n5w6eKmfmkpvSMUvUf8q7Ozj7m67/LFHoVPlpSy6oIR7nKhh57fTc8oaOT3OOsjBgYiQQcRImWNK
UCyq+bt0/JEizdkIMBreWS0sXf8CBBu7pvr6635lnUt+foMxpMEroDZbQpeFB1R2KbHYplXUj5NA
ENHaEl9kxLi4aQjIwoexleHcrwzCwr2qLGUFe0nppDntnNZ6JbFdOr6icLwz8FpNlDXWNIW3/tRG
Bk3DwYpd6oVflsEBM8KLi9NyThDgUUFWCFsdgET4/VEU7+MqjyZ0Kf+R03bdRCodeQEmFb4cGURO
sNT70U6dEUjwfvdftMvsNIq/rN9EKwzyv2ljDlhk5xJrlaqAlbDwxd8egR08syJKvM7Jb5UCnbBe
qXWmP4QDp1dg6voaQJSIbNdKB5WN34vHqp6nqKZPwM380tThnRUHY0OMe8HRonc397ULFgjMKNWf
lzix6J+f4CLrhPAQjH55qjLed5KxzWR4ZLSZXCi8Nq83bc45ht2H7qSkorQ5J0OfGhOofhrjFJwp
lwSX0QVhINA8uQirjDe1ss4I7An2/cQMyHGYcFCa9jLx3vjJzclOF4rrXLGw4GQgpNepOkbgExmw
cFj2CTvYjgZK9R6NCvilzATaYpwtRYIakMFNxT8wgAF1zR5aIjvo59a8DpTpjJNqq8rvGxQyX97D
5O4SssdNTqpATh58/fqblTAVtmLi00jYSPZOur/n6/38Fjo/VbNfOzKHJjN9J4Jrkf8uIOLXAzMh
vvTKeL4IoS3ICL7xG0G2ZpAKDY3NFJHY2dZElW9Fw5VJ0TbqAijwU37/91oC8qhQ+Ifc9FEHv4oa
gI20OQ2Op7m9QW1Ih2hA/ygRB9tcxqoEewaFYq2o9vy7CIw1jfXdVXIGTi+lmFOOtpkDDue8GIcR
njeq/KA6+abWHLLnajRp2uKYdb2c3ewL77ToD0iCvcxNcePQazckvBRsdap2shrOOFWKTz+loAss
QGiWs4burt5fmfjkvFBvBTwyJj6DygPkl4ADVoCOEXz17F851zVEkMNWGJEe8Y8+xgmGGBN3dYFJ
x6yJ13UHA3mYgGxOiIr/fZ+rj1dMtQ7KfQDHOmjdLNMKfcCfhEzeb3iqnQgW1onh+5OweaM+3in5
ANFHHnzAmajtg8PsW1tekZb4k3K/Mw0wxc4AuTyuw27d1nfpMUdbHUQ/SglHM5Tv7wds8+BFsCVq
ulQ33kBLqNgFVjLVZb98iOghfjwCzKs6JAorKazppWOzXOtBI7DIqFshuFD83Bkt88xMqBu3l5s4
Y8WUYgP+i6h/a/z8ORVcx2C2rdD6+u98VkUlhBxuz5T7igUfbtJdcHgf0w0AWH5BUHSFrZX++0h5
IyLtb8ed5ai5JSLC8FslLEXmKp6b3FJr81Y/ohJK7MFIS7eJd+iCQzz9WMmG15L22uVJI7KMhBxl
ynG5VcSsyQUtKpzfKioigISKAJzz09nHG2Zcy84NHrn3vhAti8CL8XamI2wpMNlwQNBTO4irk9SU
PqPWQZAh+7ExfrIv2crvY3SaOZb1ZdZ5hehoHFeXz4jUDTAmDlhs0m9kzOdfUpvjUlj/sL8Mgatb
biVoExtk9b47ZwdNtvTX0Sb0HrfLgP7X9b/kJj9bIb4FpFnIEtI3DK95YaqmdH0CBA8/025eHy4K
9Wo98HkIrxqmJyI1WQB9ra/1OsGLGKpV4lHhp0Bg3iwDD6+6gULyfq85UTNSNLhgcxafJMc8IRxW
abc+NXag2i24hVQmLlAN5wCRc5vrRuZukPhNuMqqZyGFv0b8DerhyPpE95wRu7xA/1it7buHSGJJ
AlMhXTU8LpPmqpxIqao+dzGxlAYnb/IYh79MQ1k2k+/pwxs2QdZ6oh/0f8lmQc3HPAlyoRu3ln2c
95URjgz0iCXdicDs71d5A2hYayiq9nKzd0Z66Yka+kNEVBk++moDJAplb54faM2u26e7+IF4TNw0
1whXce3pMNVmi+jkV61gvPQ0Rh4ehpBG61ySA042ywkq+SLFDBOuudcGrQ1az/WCRw0AY//N6d2+
HmYDevnDmfpb0jyRLpi3WULO8La+zZC6nrbuTntqJTnt9TC5DIzC+uSZz1AWd8W4Eu4Jr4PfhpFG
NxUGeAn3SwlaH2Xy4vFLjd7i67TvJGx13tkDdNVTCZu2Zs/pe/leem4cTFwm3Wkq63wdy3ufSRfz
wqqfAVYJfXG/fyKXAV8kST5lJbJpKaKI9YG/WJtCq9EgxU4vaJ5q4cR/ird1o3+DwlbDAyssxjQz
2ORSZqCqDUZHBQ6YCVyvsEPo8fgkbQGsaNcrdcMCX405sxSOHGBFZfzwzQuWfOruRw9P6NSvqS0p
1ccQH60ZW0Od0PfC3ZVPvUL7th9S8KXzqpDnya8m72noJ+WLeHuppLFScnexDh7T3D+n0llQdqfU
Rv5CSs8obKoWo/0YBpI9pj86EkInG+9Ou9zjhlOfZIT0vNI6ZF4Pbur/vkr0eGFmRB91Iu00893Y
VQdH52Q4HG4huDnGkCo7bZJqJLqlrHmsq4SMIpt4x5w/xmnhjknCZQy2u9g+zwUi6TL+naKH6caM
gRIHuKcDNjtHEHdKJcs+QXpq1TDu6gon19an39Tqd7UzR3fNNCR1sMLsGzNZi755+xfSEpirUxVv
3n91TLF5XxfdWsEUt9NksKbpzMtO5rdtSrRsjZg5i3rIcKOXyxNF6N1u4bgbrw3hZxQNeiFANcHc
RSIXy/wVH4xbjIMUlaA3OAs1D1cR6mC/A0vtyRrzD/T3TF2WZy2IoAry6aIWA8I1cp/X0meS/GWC
O+zw0iSH+V/I4KpYmqRB2+t8WwA/gaNTLm4JvntTKtlM7HYaMgviObXxWP7utk5+SaZ7Xgh17MsS
7B8S4djiNCuHhj75NIoyuZyGzAcoTwtTK3Ry4BV0gYy1BVXQFvMU3pHP0FNwGtw4DcYi5qZMXJ8L
Jdt1rKqr7rTNejUxVVJgmksilZwyNGrnFMWc5X3nVHIOsAWz/ZBpCQmY057QHEycEfdCM/O0brZA
oSDNfA9nRFpQDk1us0MMhypwEzSeoL7CfnVhQHKW/ENRESRN4D3h0AwxuY5kPDVYnM+eVnobEMiJ
SK6PcQe4rzte7yukDrLWbwDizxXELzzyYqqjYcQ+aGi+aaLbY9+/65QAZdJF0zKJGBQwBe5AT9uA
lm3lILjhwqJv2yAqxSdbnMhTpnor3LPzNZlgLWE7UeDfEMBVgkpIn78g/REHu+hoD8KBDxSKywyy
QjI8d98/HxcF7cWepl8EA++HJ7twNoDdgw/bEItDti8LlLAnN9n9dU6AbifnCI8Y3rww+UnTSoOq
c0j8UI+9rvpwrbH4fPcHUcK20cbDBo2Eslb0Kt9BbMB94gGRxpMwuzOmRnrg8XfqMNpQgunZmlvu
HB8k2ZAZGR7Z1ABfkjy6b6v1rEwDEFHxBilJxHpjYBWtIg3tMTZ7ZaXhaZzpqR93/UYvBupYyOfY
aiydu7AdKHBULTxYZV9IBX6GZCo0Z1PB8l8IqTtNosEdpTbZk/sVtp+2l8oY7MRrM+4bJ1ONZ5oo
Faw/pYH3daOXsm4Cu9niJdzsjKQEGnMC39K7RwHgbVJneA6+27fVb2gWuld8nk/J5pmryMdN+/KW
OIwQgzva612sUmCHNdjRHpf8cLwfmrURaevl91MdA9F0KFiEq8odMrCQvfhmi5s/8PsrZZKjFn6I
pqXwlb3H860ST4Dw7q5sWEMGesBzuKL1Ge3YZusmnppZ6YhMoYW9jD/SoAQCtJ2rSa8asJv8WH4B
CZEf/xNAL2BE7a9TZO7Icy4qmRHJ8K0sz45mt4JATnQMgHids7N9nEEO/bzPwj+tOLI8A5xFrOQK
1+AwsDnTBkBEHWRq7a6Sj9wHZvVmBKuIkPznlG99lVeE4zu5ShlVjwS3ixmPs4Mdcf2E4nhUCPim
tIyd3w7azAzC4VDzNhruU6QYUfK5eU391ibB/fSYQj3b5OS9wLNiLThhKvAs4zZ2iaelZeSD27Co
YjZIPpozRx/UY2RGe3RNkKAg0Nxhw2RMIEVeP6C1uJRpQ9Ot52ZFfY/obAUBxMGBFxvIlLQIxlYG
Fc1cV9PDnNE2jvKEAF0miOVm05TgWQUBz6LsNLWnomB4Q9cTJeLYYjC5fTONL026Ik0G1UaiO55G
bmw95DWQ60VXLpyVMVMsPNNnykRykHEWqfP0ierEzsjIaHE8lUYF1HmvlOYFQuBSCHWKQ+qmqIFE
0RTw0J+SJa+59qmtkA4ENI6xKprmyRpbN80H56ioPkbPrLQEXv43lZ0fq8bFFGzSpcJdd/X74NHq
nhjxmLKdsxMURtBO+lyYGwbJVd6xYWVWhLQ/KtjTIAvD8MMOuIQEu6drrckWsyogrDt/QFI+Ucry
yInJuPcV6k1LFyoMncUWXe7iVKopT6OEPSnPhTiYfDIWVfqze7hrrh8YKtU2r4KxSvwSKWOoEd3D
LO2Y3ms/LZcsY5v4LRXDQpb5kKZC8cut2gRUTDRnIfnyzakuuqM+8s1kgNG6C1Ot1S7IuEHssbf1
aig2j3EmrDR6cGMJXSraVjPMgByfPh9eFTx9hyIiC8a8xPUIbgfjwiDaS1k/nYV7C6U7EHkh0Rlj
PO56pc3EZJCuJMTXHVUQ70QeqdFDCrFw8uJUY1Bb1Y6D68BAGd5sAyVNhoHPBao/SCMO9e3YPBZb
extgKDtVuAOy3548B8gmF73tRVsqiQkZbGrp7D5MPahA0ZwOrmhmqsTjZg55fxDOs6Eo3Bo/BlTU
VeSdf7iEOmF6grqsT9is3Hrj/gl56gRO6pHdZP9BTB+110pOrjtPLLrF4GVZ2+NXO2CB8RW4Dpd1
E/6pejp3qg1/WSOny+7DmRfwAsiDKE9JGtRuHHFFotpn+USiSnPKCmzd9Hc779dtBiN8OG0VR+0Q
mTvBLlYbwxFSWMKNjqHCC7xtHMVsBmaZ7Dbv1RA5rFVhqbboicUPpPQasJHo+kQTpHueOkOXxFmh
Mb6fZqU45UQ35cS/kztJh3loe1BUYZcJqIc+QxyqdO8SRquyHgphh+np4TyscNxSnyNy6yIPO9RT
t74JnHMEUiqI1kAb91edEGd7xYoE9PGpMLZigmowAnNQngXrEZkfBxt1Q5pHdeZ5dvH5h2NFG2kP
Gpakvv/ij2mGDit+fvPHoskkGedbCpLXXsYK0jPr2z0mLhswPccGEQTYrS6ph82eR31l2fA8A5eZ
vWw2JQkyQZacS3SAqujP/5EClqmovP6re1cwEIXazLzXw+2o75IIuMBDGQuD6g1laehRqyJi54Vh
xfW4Vi7HNwNtXFEKGKduWZH9YiqiLm6rjZP4n+dZdVMLhKYrOd09OMbmszqhWw9oKM7+eZwLSnSD
UuIUfMphd083v4vZ0V2+hG+IIUII8BiT11ZiZ7ntOcPS/zi/kvAs7NyXu5KAcvdrd7R6cLUlq9wD
7bbqDjrbmmdcEhmpLLHrdWT1eFpaF4Bgp/3WqrQEzLaDq1v9N0MDYHiWejpFbnO2AFi4uQOSBKnC
N4Njlv4Ux2RjOSug7CfO+cy0XrK9UpwLqe0+qj0SVvuj8AvGcJDI5Zl/HDX0Ew3hBpIriPLy63BH
wBDMJQU/byywYgSLD4Jwu0+cPRtK5DE8R7U0RBHhLrGCJ4COuDoGfKXOGJz2ifgoGZ4FqszE2RH3
/gXwlw+wO1O6aj/eh5nHO/q/vI07j7VooKCmje2gaxOOy1lfxocnxCA55vDDmTeflaujuCC3oem8
2QTQJpIpWGww4vDtVmtaV4hPJh0JtXRrTqEexk3loLB+sWp61UU4g1KnGLuSQZYjpCG9vSktbXC3
tLYqNEsdqRZbefHry/OpR1BG0sf/oPiK2ZIoEOipfqz/U3o16cxX4U9AlxGdCHD57FoA8V/TJx+n
V7NNnFiVVuEk7IASkSx6ic9e178kBP4uuZRtw6fUkZe8KhpJkPXKVjl8I2jQMPzS96PBVS5F73tJ
2dEuef+egeWnoOIJyD9n2iOkPGQSIWSAAdL1UaFjxtSnugYqVEOd2OM7Lt+jzhZaSGmIovfrTvBZ
5AAN5sL0WTlwbvzPR3oKETyz8MLK4H95CnT3lrD7HenJp9BevTJnoq/GPOHKIXQODdrDNVzgQgS+
XgtcfhbVKRlyHaTsCSgebqORhRzn3fcuUr4V23S0TNV4ezOrJT1t/pKR5blHqOiwFoTCdkRSt+jZ
AuLcXIZp8z0Rkjzn2xcYllWcRzJVJbfQ+oLPOk24/p2BY85r4VOldmX/G/4olF+rmENxy7xaLwsI
tUxkt8LeWbxQe4cFbEATH4C+iM0+b/y1tsXaGXXpwFs0ChpzSBBLEEAd/Zy+4m3wbWJGxcEB1dVw
oqedNcNKfR5Mjx1uYUciFT6r4aAMX5yjmR+Q+AprqWUJOlfaBqrP+WLcPn/vzVfnPae41m9N4S2p
hbX7mACd3mqCjmecxA9LLcWgHvZRUY0t6oKu43GAbQkRVbww8JBIMdtk/PO+sr8rfitspXr8XXDs
GQm38N24+afl/mYYMdMRpjacOK4//PcrRLwRQzbkK6mJqvJ/aFRCsaGViv+iPAIAVEkcQNEgNHQj
vjGknBQGxiUHPyne/ni8fjtA5k/vSS5sogGaaxGEu20eoxQreayIrGNhZX5wQkZH6w5mzL2168tO
4I1+FPyEWJkTNRVF2rwwA3NO17vHF9VPL6Lb/gk7JKDpu7iZNGXnYckCOTooR1ic5zjZiHapqicm
e0Abhnr7/1u2iyCmH5J96SeLt4JS1vsK9jeJWyXrrvsE/cIR2gnbmKErDBMvwilfzkgmo5xMXL69
74Q2Jk2S08kxKP++Q/EInE2m/ZWvLapK4m0gVYE/IiuRGOBFTkg1NxgF590popWwUGdFVSYRdgDX
TziVxqZ9Xjm4h+GVRrLTu93OeOml/5Qq7mBa5rfLKOMdyh4T7yGIRkzDnoxgKsgvhB9F5gt7gA6b
ZWYnVaaqB3xrl4+lCXIHpHWYEo0hEfJY17G97JM3S8w4jzXUhsBMMUlbGpOC3SwSrHjZXSm/mvKo
m+nhrgELzeESzxmt3f0aBjkNOsluGnYswhrLnuEk2M0l7AsSAQRAorN/Lg303u/Xl4mt4qKw1HOi
1u6osxraWM03U8FfuKd03PGHMgQfU3ADxzydlxDvCuU6qN0bmWU4tzVEQVZHo2INCO4UTp8cX0bo
yvOCgGbhlDzfB6tO54GaU94bc40aoJXsIbAWmNjcUiJs2l+ocB20/HBfC1EzmjwCgIpQ8WuNr24W
HJGlt/tpx65mFrtln7sPk9C13cAZhQRbXuuJlNa6YkDoOagqZDQAXT9lfWvDc6zqsSI0JZsvRxIu
LHErdFLIcMN4uQclYD/njlWdwN5ZD2VzX1n+dTbd5U8UjaJunuH+av7Qg8F1PUGS3cSGGZyNes63
E9H9pOpklG4dst5oh6ATIIq4Jo0iwNZQgq4+pTicTNphlChr1T9ZhqqdmBXX/IGJVd2HZAr5GmLI
0nTLFXswxDflpJy1wC4OV/RFOqwL+MyoX7+3ZV/MxUTJp3QqUp+iI7z94oiiOov85PRAxHsKof/Y
82kXmy48si6qjx0HsaQi6A9WcDR07xEX3hii9Fj9/egiEALeuHgUT6yNXKz9YZVAGLZXlksC8d+q
BGSyteCyj4AiETcK8MeHu/hdVXNRXuXGQwUtfoDwzfiXh7NHX2WKWwG9V993m5n+zo6zI+OJwtGm
yEjnQOyBWcaCzSTHmSpUs13tEY2Caips3Y3iJaAMrv0x2QK0lzb7/BaJnljdWjEQ/30qP1FXGzIe
xoefxEuluH3dHi0J2X61OnzOpBsbEg2cXc8B/oA8LGdxJmD8vWlRzMUKk39QT8yhNnZ18UQL32uP
02gCAwLf6l3uKesqa3R2aWHvRy5J9xdWRHUab4rpe1xwUXHWD3rydgmNfR3+9/KfNAYxsNFM89xP
39srQHXJQJ9aus37Vpahq+ViUiAnxfWMKxPfQqk5INyqwLYHzlE02eYm9Pwp8AkVQ0nfRpUPa/SF
5m7Ud8MLgOxhPXYz3G0e+Th9H/u2OlO+LB3cX6eqSyksufsfxoi6VsaIBvbXV47pZ9TuyWzplLer
gbI+6emkFQ4/E4UQiy3eVTbMDC0z6iaYM1ZMjyXlgaWeyPdnPBwEM1pGv2ReL7HZgMVfjGyOYfNH
sUbPgE6gk229IhiixOkJxP5tjTHUI2AfPsd3sFOyVWy6b3EQRVD4wJ2n+bYF2XWb/TX7ZRLKCZOl
aGfP6kKqecfrtqn5DtxJ8F05XNbQy7e7hFimsO+iYxDlh1+D4ikUdw5Gkb//8553kJse8KzXhMSd
dI7IltHnX19/B0TMGeXCcgM5o3xWwPH90rRlGbe5ajvrDy9oJz3ky6P07lTEodPKGACyaHIFHXYQ
h9vKZez9FdHIQkrSZ60pbBr/rwo+yjT4F27cpqbZYinuX3CmI/07n46NJni+V1A9xKXyN/WpWF75
fFGbqi9YPLnO3c1fBodi9Vz+c5PT20UdRqVoz5pO+hKs1rR6JiB8wEdHg5nG16jw9RmaGPevdddK
LcGdsjtysrlaXEfC0UzDR4PUnSGQ1chRYgmeae46Qvq5YhsvtCbmX5AK/+IIs3pTHj7pHtdlHG7Q
Gh9360AZGl5LlCdO4Ve6P58Y+ZREtfmUHSiOiu27zn6w+u2pF7s7sCvNOM6pTzEP7PrUeybjQUod
G0eu9OujwCy88P+l8X0W5MkVmxoNYzwF5bsp5JwacP14PuAOkyeh1VqQUifcxwaR7VEOIE03IA1V
NimhfaCnyRCcreCtJKKlq4X5yim/XsOBXZ4oTDLQzBbcd3VDjblhMi0+Jq2WDW7f7K3GuoHsNPwp
asUKsTGO+pg/ujtw+GuiJ2C8DaRk1zi5govvR9RBm/C42QLK/3kypC3vPtZawpWD+SfDUU617IoW
qLXP8KvRk+NPMTFcMWWN22AljW3mjQ2LNIcHP1pyzPn4ZLzAgEl7JiUuEOLwqrkG9l7PfSXelFZ0
HB2gj0rGUtgKJ432+PdVwuY6XKl6yvfBIBMmoz97zRZsOWY1xvbhA0tRwP4lFUh229V77ytN04fF
lEdCS0c15PrxLfwJQK9GzFbMxTTn1FaymKcoYhuaRmh0+mgQ3laOiWRpZyzQ7GewauJ0ivRL/zxV
GKjosPJ41dmVbT1daTbjgwjY3l3cnRCKaTq9zc27kmdFB4wKsVdBL1XHd79N6hDGRZ32IoGZdSl2
m2fxBSOewPZA5g1Q7+nusdyJfy2U7e6DSIHqOlU83HsdMnSygNK4gkmaL2gfBtLOs5RjrNRoqXUT
XIVRr4KVIb22bd7Huucp9oHIL7R/OC5gcRGkhEL6ssrMoPzCCvygxGTbM+YtPMGC0iU0szed4bVc
lljpmH/xSQ3vqU7X+H5LNjiNQEJ5Z1+oH9t542lIodX/fu/5Ybu4e7T70qu7FGl+lGEfRcYB/09X
EtquL4mOzolIVvohBYWD5p4tie6bYEo5EzYJO+la3lNYdl2WZ3xvnExnVq/DpCF1QfdIr23fIlJI
TPh2GOrRlyGzcjJZQWaxfSiasUL3R6Dw6C2fdUxcD+2hBYCj/LkPH7JqiB+UIDUqCg04k0/QFU06
dVSxZccYnFBtzqCz+sDEwGxmqXbau5giQcXtCMno/yQVvki8Rypem04+GbhNevOFix7CMfjIlqpk
hXyOMw8u3beaWbaUisKZiAlVXuOEyUv/pPAR0ODnRqzu4fmDHHWNN4tbOU7ablN2NCufFrbU7rnT
HW/yrnOsVPl9ThUcC9HTzLjNb5w4DdQuqEPJAWFJDPfOYLt3D1we2VIHvQmSlNRWhLrj/0Gu+77N
wLwVlyEPMy8KERYwhagisu61R2YP5sbFB2gMH0blvamYdL73Q1DNr/yUHbkJ6buvvFfUF5xcCS4M
HW4qPKuUXP0ekvQ61Kqc1FJdMSMTNBq1hRK0Fxldu2YA6AwixJgtYkMquUXnfaiBnCMaFMnRQhC1
tHdYGqBha/Tq1e5rtfT8DLF7x2zmLQRtU+mrgovIOiM54KbErkLXzJpPsCSwlIJHNApJ8ZVy3Ed4
10DNXcrZciQjIDSE6IKGQURxGTYQe+FEb0VwVWOLCy27mMG3CRn0LoMpc9bsuH9uX39wSgGYyaRc
RL4NCPvcI7c2n2GWaaXkebUfEcv0VjMtlHVw18H+xFCIERpiTZdP3NGs/czQ68xrbDIcQIgdrE/2
P8gfg++4YD0fF4RubBHuYykj38AJ2rWyCaB9MEI9zj/gI9KLK+O9mc5jU+t9XACseZ0bMNfc3dbs
4IiAWU3s9PIOGjL4bpfGqPkc3QqvxmbS/I/4n/DulaLbBwB2XTY86/h/zdyDJk6eaktbphB0KtT5
h6TdrWxh7Dx4oP3i06rLP8UAvOIje1em/74PUtKhjYLQIb52BQPtjpqSLMF1FHCHKzjekq0jw089
2w2miw+kNmii9Xoiyiv/eO0RoMByf+aWrI/ZbHiyk17oGEdz9WjCCEg2DSpKp9OFgte7ajGkauP+
N1ClLsD2IhW9bRgjsVQekSBFlF+anBtmv38a7h9Uzu6dLPQSW8rYbggGVdEBh/mAyOQGePuDghrw
Oh6jv2A/ZAR1voYhYNXQzALLRHk7HDihrc1Ts51M18W3Sod8NGLELkw2PKabhgKo7zmZ3CdDoXMZ
Ck7IEclqgc32/WV+9wYb4tw/HnrcFfhQ23t4rOruCJpqvrWml0IULKsm3GYPMZ2+o3mtg30KbLQt
gs1qBaMwNdSsn0H8lTJHP9zvh2INXXltrJw+jwSuyLB1wsEHc0SFrDL4/JAlJqlNG7qRamPnEZTd
yWNKSbPuB8Ww/TO0h30cTFuAHPHL6fent6bryhgQCry1kyEd2km7Fu+ilg0v5Y8QZMGnZQneM2tN
Dou/2XckTgZmr5ixIoJWOAzcVdiPUE+xcSBpO5CJgzY6zE2O9JqGOvYW8ET4RE2YuGlCstsfaEwv
2iXsbkoGuh7fLqPO8GDXuOy5/cdOTzmuiJPbZwyyBt2XNIPELHCMHxfLhpLBuUxvp43u/qHUcE8T
LQ93e+kQuZrjjnibrh9ivqHGFW+Au0VjMANv4KRHjSCocczfD3V1sIhKCIGOlf4NQyX4sGv88/iB
RO8g+kJNgSZxV7nxpSl1A9GVHC6ryqSnI9YmyLneqpbbS89DViSGZj63pr7BwNyG9tKp8+WYS82y
DpdvNR3Vn4t5YdYT5Mtsu6B+ajdA3ukyruJgQR+0L9krIXPR8X2bbHQJk8kWPLjLpLlVMfzEkMBY
NkVkzl4PyfNZ/raNoMAudb3NKspHZ+2qxA6EDDkF5tSsCcpEx4VaKwexYhmvP3KhMRpz68mT4thZ
wR6DhvkC0egc2Viz0KiDIdNtmXMkKVE9VeIDBAZ6reP39JW6DR6YSj5r1NUClOOyZw2VlKkE9uHf
i13J3mOV7g4dxBljkEOWUE11xhn7s3Ntbc72uoPYnRPvnp40GV87tKaCGd9K4m56HvDIYZYjqXSb
YWExL5v26vLiQ9hBcO8eoARrj171gzpnZMuN1ajgYZVZKzt7+LIpRL8jXSaqLiwP3ZiPExK57g4S
DQdZa9oI/mreS7+SvXJbSiihRaqF8rVOG+tfYE4bRx3aJBbm/ySrMf1O1j868Qz+fQeRyuJH1Oox
Z69or937SiBYl1MaaHpLxE/dWZPAUH5arMra4rPqrWEozPFNthAlRjj+hkehz3pQTK6zM+ur12Sv
5fYepkvq6Bn/sbIOt/hNmDryX6GsF04f1w1/P4PsJ+ZyrTCrXj13Flqn7hZZ6mX/7pJvsjD71B7r
OBj2B757WqVH7NZAnHRcfIl8reSkiMW0nZaV6gvVvq5ZZwHdUwf9hHGfC6pjEwRFMMV1Fb1Nh0z9
EI1BQlYM00nG0F565slEqH8escQY5LA/P3vkr7WjsCKVlVQ8PkihG+cMS2qlxLt5oPJfpstAUglv
nJFMmyEC9Xfn5kK22YY8vK+Mi89hZO6BRplnM8LVj6TmMKqStW5sV7xZV69wGvfzQVTq3mTMfouP
tz6xYfhvwrv2Tu/x8hVPZlUnB/WRbR2N0PqB9f6yxcJ6PabK2omXH9+OFt4I4niqHgonV6RObspE
wOcnwS+eFK/Qks0kpth4qcUD9YUTI0RLF4SwdSbYlqinLzk4mX5TKTPs/JbGIqHT2HtZoPwliF4T
JDBGZg2Az/QefaiHCn4Xj2Kyosv+WxAxXLPywEVhdIJFjGJhAJ3UQzExmVuihk6dLd13xsn6fvte
4njyeLR06ZhSds6w5cSd5WLO3zwjTr3/2STQs51EpV6fwk55ocC+eznXMQtlPqEZpF4eObItgoYN
FqXcQgwm3gKG+Y4nIaMxnfUyg89tuuJ+1+dbQOQz7QvgU03QSGDusH0Nr53nOt6AY0e6/fmoehk3
2WFnpmkcXPvfKxNHJsh/de9/igaEQfwq3codhYIaF+xcL2FSUv9mLz1QZiU5sPncFhxTbChoUiVx
9thgKMfKkR0vR0pxrkVDiDoXOtkWdIpgPsS7RaxQn9HshTgA3YZtLkMlNqMLlub3xIZZOUCqJu0N
gSqUDf0oTYroGKYiXJfjPlCJ97V0IV8+WQfohRj+8UNvNJ0V/CROgsk0AeGtVRVW9WO6TZ/P2HzE
g3lVOxpvjnxuw3NsYHIj4iyD/UAWzv0r3DuLQS6/jBxmnF5Rjtw1IvSdqHc7ZmlZnNaNhHBsbym7
3LQW7SBwB0lC4TOfy1DbqP5hjC4GdHvZhQUu+Xs3qAwJYkv+PO0S8FQuzAB0FjeH1CezcTgxrBBJ
gARiOlPTlBfm7tx56bob6Qr1OKmNT4bMmKcV1MhKPTZUnKKIxurNJRnX/41RlIoBADjVpKdndqKT
tv3cOT68OhBhG1PWrIYPCSMYNfMToDfBVGulS1i0C7QNhJp19RaQMrsG8U1SfumPJp1pgG9uHPR1
KIX7gke5Ic5amNfNPNQDVbkkMqC8haxxhxl3oOWbwfTevVrve1SmceWq5xb3Lld1vQXKchdHhcKZ
4nTDabP80HFGq1hhNH0O2DmmmPnv6/xIZ4xmJkvBOFKk7yzDyUA4u9HB/MGQRIeKonP8K2jzpLc7
VRAlvd0tvBaAs4K3pd9Jq3DI0K/MG4GrT/BdDJ7nUhq1wYuOxBd1AHpVbu6UsPzV7Du9HRZamRes
6Ga4fjWR/rfAdFjwrgJSZv+t8uiXkXrQNudwELdx9tHnTZshMKX7NZhFX2Y8bYLJy9T54qyQWiYW
MRr7ipz7M5A79prwwTUKgucCOVVKcLO5RSl4h4accQkisIxVeqnu5uftMN2u4qDA2b/zhmbvIS1x
nE9x6k1PqeW6wSNCj9pyC//PLBvLPGURbP9slwY6bcSG0kNjGDgc4Pc+Qw6OCF61PT/w/u0yngby
rZ4onRJ4/5wye3L+Vg8mU3JkFXLgkIUuVhqbuYy1l3g0RmDWsq2O7dGHOGrtLdVgwqkPtBj1icKq
selZaVtnsU64NkZKD2BTzzZquzkweRJyBzQzB+uUEM11XOTaC6WYBIFy5ECfNbWUP9IjKyxEq2qW
02Q/EJEat6TU4rbShW4YpRMhAlk8cgqNDTb922rwDftgBdSVwjmDIVChCfPm2kCwK20BWB82Wnvt
PzPplf4e5dYYEJc7f88YnPTxSwVopjHL68m+/L52QxR0UhuVuVTjMdIjRAKYwKpQLUcl+jij4XBt
FNg6kYRfz0mNkyuBGsS4wm3z6UVDsR1w7hJ3v+WCc3TeyyUN9kT3+CE09bmC+j3g8B/jqD3P+cuD
pdDN2+ex6RpymVukv9oYwrYEyaLbtSX9M6SiBmJzOLeWLvFucnuvQODaAVZt1Zcf6U9la+AxnUs1
7I1rfvGdHwgo6oOD8JNFqsGwDkoHYPXO7TIaiQ8sLdizVjp2yEgaCpYlfYJVVps+QJWQhTYuo1Dt
Lc53j26Cwqp6/eb/7+lU68xr9GMZ1WBgwSODBZNx1o57Y7MAexJKF0WGlm7Ro0Z54yNqFazNPiXS
kMCYbGybiAcA7T0FFUNOyd/0EaGeqjHLrsBxmH4V6H+Owbkqi5eSShEDwqvlVwAYSyWhWVD8MW4n
JjSXRhTlkzQWlBmq/AxDhyzEVfZjyorvCFGqGzTxhsFel/uLrWPSssBPTgJOMord0mm1C5oUDqvV
6VBqEraROWP2hLXq52gq5+9nnRC2D4Twp1p6d0IVl2tZdIteHNXkeQCzJrkNLCLaDX2LiOMV9rac
pFTaFT6jqIlpyQk/SFScmvJ4W7G75iDj4+gKSZ6P5zLHBKt+0f8i9/Gy6UCVIRB7+MkwYGKMB/3f
c2pOoq6O+GiTmMBS3UEPFG4zextudQ6litthiq0caWT4RamMM1LtGaAWTckZ5/ittlgKp6wf6nF7
LAuRkY3F5fBJbDZ/MjWImVA4rYOHlc2EVT5YaaQEugt6GvjhrvC/LVCF3ejSTWMPDCrEDVon/yr6
qIpLZV/IY+VN0wwAJKZan2e+RVjC2ZA5d07DMyoW+ldvAS6mDLD7ick9RwvxZ9ov1LqjpZopxilI
xIfHGqgWCgtvPa6h6BZvmJnqJ+5VV7o/xgDjZQ97tZDwh2vk+a0IatV7x57qQrOdW3JJeK8W4uGh
fF6wneY1BZU93U3RQbXbzK6JlOMTwIGKZxgIRIsO0ku9H66AaozqgrACxo09BGfL4nbILOT3WCSb
gSwJMbl9olDG38ZkmOt6bK1vlfVplFmFCbR00NEDcgn+JqV0YvxAs7pKb4WapO1TEXhMMtrtYDge
ydU6IFnuW0Q6VH+VOBveyZXf+DakgPdc1FDtfp16MUNMEv/6VsRyIqi1XfTmwKsQf6vXhVEMb7CC
NG0ROexXeDWu3esGaQ6iikx+bRHX/4NXz3Q4WtbbKEp1IokRSj4tcfY/F12k60lFe9YR6T3z6QbH
5d6tdIOox081eEIYA2LHmCxJMKgyl3V3depcsCCwBqUe7CePpqlPxcWheieEay1OZBgn8x3rrfzT
N8S1FXQ905+Gwd9eF0MSYD4wm+qmr/kQYaVM49IhTxeCG5gxDR9RI56xbVMHfPWqjJqd/ssyvpxn
C+15JwidBAwIO6qFMDCqZ9Fvibo3xwyfIdbEM8MqyqPoE6+dloY6BMi9CE7kKSHLBNbbvXktIoX+
7S4v+iZv6eHYPovoZQ03MBqo2gOUuufh8roJbL3s2ajJo+XmmHaZkZcfX1BfI93AezzvKTfEm3dU
H+HIhRzZjMfqB5xrzD3q7QmGmRpSNvafll5ReesHPKUNcTQObhx8ctwQZQu0x+JUpVnfNvmmIdbl
mRZY8E68YRqRdbiBUAMFo9ATGnnzwEbgxOKlxkNKpbPuk5ymhF1xscEfzRUDKKkrrUw0fpkrocCn
+pEjuPlMfFHPt/K1csIYYbuR9G+q2UmCKm2Ax/XmjsP0jpkQhoKDFPZCAc1lHVv/dWJzstoTEZGo
RFmqZ1vqjM45T9aJKRKyFT0RMY7P7y6M3PikzLPHP9BVR95jXajUcDQf+pShBRuH1PiddF4oMpfc
rBwXU3EWKd5pCGHqdzlEQdHFpv4kwnIJmkOfYIhdvjumXByvHor8pGAuEnMJDtDCb4LaePxFzHLS
G0zOG+V9pAgiyiBy3hKRdYSnvLdCe5eDsWiS9V18C9K/NigtodVGBC8Pfds0DveSsS72qrZiZ3FW
vfwigIs7WaesdEQLmLT8UReK0X/N2rQLYDHRZfULBA2I6RIE7QRtNtn+VdEBgkh4K+z8J/vF+asZ
1xtAwkpw2jOCFDZUOTzM/dwPwxphlI53VI+mbX0hAuMmzBK4RMEdBje51qoMAvNxCiJy3og5JY4f
s3k1KN97oVBLh0C2AddDb6HjC06mWDI0kqWmnRQLXB6P4LSkk2JjMdbGNins7kMLkxC4A3J8rFSx
8wXY2YE1GTT2dG4u7vM6Qk6eK55y78UgQYFTI2gxt3WNi791X6VuXX+QN6xrEM//6UIVsu4TGxsF
SzFPWArGHPRCBbZmA/c5RNDxTB6Om5416bwXqBOut5lgAkXtBXC4+p5tEQg4P1aLHMfa9kXZ3ZkL
1rO5p6/xgU8MfeaZVtYDKxdSlJXsrDBB21BqcQKKd17uAZHdTbNC+b+wHmAD/EbGD0B0kwXSaDQG
+kM3CPma0y5l2TctdTUzUMIovXNVvLhggslGaShOXxqeVRgsHEOm6DKxodcxqgIIqrZsHmUMMQ+4
8XsqAVkSEIpGslUvLJS8mhzK5hfwMF5cOAoModxC0wdxKV9bv3VZcqsqF3z4fbb0CPEFZRSUHBjT
SKpCnSWIyN4c4zY8SbqaONTovXL252Txaks3eSck/gMKg8h3i9r0ZrPdlv4ic4z0rIXmyr3jlai8
v1iP0jUesDLI2fFetpOrdUmIAMhA9s+zHAbuv/nPcukRAYdfzawBDnQzlsgH+l9PwtcNH2eajRAS
Pkm5oTyWMrbj1Z6sFELJXXYFJ5NZQ83SYwvbOr9REeBe4lHqTH9qxaHB3W0CBkZtNK/Z1CEMKv1+
w4yRtb0nwywl72dwjlG9vufxRhYy6kntk/5y1PdrOtzan8jM0lQufnxOvQCvrVKW8ZK8wefTsFUv
8jj4vFitgx1sv3IhWABWRQ98r2DChQSfNOp1unLK/75yBKUySvKRqXWrFDkuedMJ4o95ZY7kiP3R
Mx7GOAfo0XNo9ljQ32xk/uGztDroSboJp0OUCpEaathmuRYzM/SwgmUdOXztKebGP6NppLPyULM0
6ElecsTc21AMT18RGMcAhbO/wffeEQhc6L26JyK/s0LP8hw/xSbOwJYF5MqGRQzwXQBziCrfw8A/
lU/K/lvi9xrJ8anjrwo4QJp0ASK6COg7Bk9nLJnMfw85IXIwJ2ZiWCkpQIExWS48Uxse3jmvQQFS
PBUHcJGHo2qI74XIQAChTe86XyY43r44x7dhrNXWqzmdGI0btKKnoOMKp/3gVY1pA6amhAM5jAfY
IXTLTrQpgBmvHT6qPAN1rhrNwiLYc9IebgbtsQppvknlyJXmT1pqUzC1PAW+r0ka2zfeh/IIykp6
WhbMcpyXNDA9wALETss4ozN7IexTvcxoR06TVI/dTQzHrICJ9azE/lerAIDQ9IXpMvUCXh8jdgvv
tMr3viA7PoqiNvTkqm1YII7Jkw1t03dgOwpRUdtwpkMdmgmikeHa06WUGmVDJnei35OfUh3UQ3z+
FY3hm9/V/ml23ou4eNDSJ6KiE/xpaoM3SRChn1EOekBl4XJ0MJMIK5Smci5ouMAWJwJlCFQ7wG8p
ZkCvUc9Md2H9PdTau0AfISPnMKMWJfY0YdS4VTHCuqo9Oy9GFbpnPC48lxZM2LPsmOT+6Z9Uh7hS
HcRHYo/l0d/M0QbmNnZ9/d9cU4bCFvjzCX0dRaodh/9LhsRj7AipwbwiYrQU0WfrNfpDMUmCiWp3
pQAyYOwOL/mgsacd4uO+tpOZYr+PiGe+47psMD9c73hsAv0FHWCckBhm+YCB9uUtf7AvwgVugWBL
JPlYtp3ahjhZTwrYYLpKttg6k3q0frXTt/+EJFKjzH2QdAFKfltH64I2Kpijy7MyMHrZKI3EKQ6W
x/sNnqdbRbCDKTxNPDMvwBtFeiSrrblvy5sgrKMWx4y/YVLaVb/YPFk/sJNXpvL+i99JjlGnvfDM
d2syjGriUE1VtA9nv4x3BClqAxEYiXnVQJB49QMWqg/hqCxQwwi44uTbObfIgrfPIn3+YAC1+49Y
2w+fGBtoYKVNd3bS2x2rbMQPMM5KW9pRP+UMgPAYzv78XnMqIFAt6tkrBup6duGO0GuxVGbynVyt
dH9BxrOVNZVUxQNlUhicbl/Z8GbBYCRzd+sX2e1zTvOVdeqLo1dFpIgRLzpTwQO3/pN40P4R6NPO
ndWze0T+JIR0VK5CrJAz8QH/xL11ahIkaiJaH13x8C5avOTpZVVV/ke7wvVZ7QLPaepHrmKCoDD9
34DyoTKg33emmf18WURYSapZ1XQgL0/Ie7cCY5jPLr/5C0jJr7bmweJxPbu1Ysq8nng4Aqu6Dctw
OdiHDaO/AJJySF01v1KEjVxKtui1xvDsUsh39Bukd3JOC6IGZN7GLtW5LlCK1MGnN8awFoQv85IE
YfTBeSkQxO/dmZakZ7KkekuSwMfoUS5LvTPQImv5Kq1oox2y5ziDioEWVxobnsSB629xKH0xAiN6
cpqzOQG4fbuu2eUiJFWPf1ail+qyfUffK7ixxTpgUBkGWZc4mtA/l++YaWdL0G6/1hvqfTEdIqQ+
S9sx6paduWYj6GdWdZygEXnMGVlFjks5+M+TjpSGhyy+sStjrN1Gu0vJt5DY6QaMza2iGOjfTz+h
9/q+nuok56b4j9ewkdr96w679lCN/1ETVcV7RdnoGS7xK1zzEdh1em7JnNdQBCACT83Plvcmcfyt
gbg55ECq9mbuzsXJNxlEIISP2ZwPeOWvgRzfav5eNu8i+ryUM/cfW45rBe6jiFdpKuNhy+8ViLDh
Ib5r5jr3z7r0Y8puZ+0ib9GViAoqKAg3u1xcJY0e/J0K+94Uy1Mx/HP4fcRlRHRNP1Ozt1ChnDxO
u3h6rd1cbWf7cGdShVINxBEtNLn+/dmvidtCYyyQ43nSgUj5hShJeBAnJDn2bLxuXaha1Aemtesy
FAHI1f3gtsiBhQIgbQdXCPylDh9evnLkE5peWJ+NQbDDQF4QtgTaN/Kyxo9tMFXUYSPBzfJrD7lX
4sJhVS0AekqDbXJ4FzIlNIQj6k5dHdJ9J7hYT+Dsonsds2N3t0qHbNZvjW6pMYqD4txuJVYSwcQB
5NF2pR7BRgFLEoTTk/ueEU3GFLgZUirhDL7O1zungGxtbrxGfh4rFhYia1rcZLeelW8ejrYGXMFm
lqJ5VfBppLulMm8KzLN+ahmnnpV5OI/MaNeFhQ7PdktAdXlcLOXPJB5JIzHxOdXYwsP3KzKdHyLB
fDNJrU98CAJ+lvS9r0CpRZkCxCzUNY0GdhmNCC0WT/xYzHj4kxowQAcZOm905WHydCsaZzcyqlV7
kh0vY00ygrMeWUV7W9cxI3+VKvxQ/aVFZWzN9ponHIogNIqt64YEG79oo1aET7YafqUQIGE6IMYt
ZlfhECEALfc8wgJbFSOqLLwlj+LyPxxF67Lt1TmJbI/WRk0AYreZRiegj1viHLbOVEEqxNmQAwhp
1YpaiZyDJceZxSNUyk2Tb/42G7soAYEgmpiT498/uEZ8Bn6ycQpUojTmQSuQnCXcCxDvrv6p/MGx
rYnLpm+18iQQCTMcieYGoJx4Tq4ezDzcfKFkiCszh3Kyr6aX8x7g5BZzL5XVcD6F2eTbJDIutbaf
1HgQm/LFzzy3xkiUvGw0JjfuUq6PLQ61g0qqEH+QH6fcRQpm5eebCWBAgkqsSs7ybS7WHAMa0ZB9
fWBAITXtpO/JpaB5AVKpAz5IgIXZ1cgSUfYziBKW4s1TTS11iG258ao5SP/jQgmXReyfrJe4vVDz
A+azL7X30AjCrhPZt7ix240a+xmC7cGg1UkrxjBmJIESJ+lOkKAzG6i/u6vkc+7v7QAe1WR1XrYl
13CkbeOsezlxUbWSZ7K+c6GfqllwIp54IJyw6yoW7upJr9qJza7HuaEJm+Wp3B0bgr6EpFaDQKu9
BRWKt0Fb1rgwKQ8NBooZj0Nkk0RYd9QlAw5SJK9Mvf6w6nOWR+6yHRfNjrbAj351JB7OaKPkHr7s
j/MsZhfQU4T+pbEZvr7ClW5umeJgcVq4ZYGWW5Qr9hiB6yRhSn79BULBcN/yddDu6/524QvpOO0h
+LVhejPyOZS/pCHeZupa5jeps9XXejAfoEoAZJC87aiXpBpBUk41imwGh8qCz+ipGOqYONpRZC3a
35/BwS23YYpfaPwadDR1M43golGR9rqbJvj4QmkR6kGdN3wWktxT3JsEdtq2DNEA+P7T4gyoWgy7
vImLQpvescLqBVWfvPr1FQs5FtdvREYdjwO/owNEra3cIO0cfR+npkTPV/nMmFpw8GqU5+a/UTKj
IkUxFsUkfuhzKSMkbi0+eDftNnq473ySRxul8JeWJsSg5m2Jqj2UV6kMJNSzzNvkyKJ7r/XzlxQ7
94VhBFfrHAzhclkz1WJmx8EYx+QwBqXsqLd9GBFJdLKN2/LxoYHG5WjHuBDAJMJTgbJZRSW0XzWG
za+J4/ezSG2V638pJTmQp3dH+1bkbaB6fJK3QCgdMiwp3a203Pqj/nNZwALECpsiy2mEx2cx9DBN
6CDP9RzpTSkQxxXVq6kuWHwq356lItu4RWI4BMw/uaL6yHsuozjdsKXyDbMp3njFQezfzCNAxz3a
wA1H4p7DaL1+Yq98hfYqFnbMqTZbJO7tr3WNMdJCMmxzN6xVANWqSLpHyIHYKVPFvOtfY2OLtaRQ
0ktlvZ4RL9so2PuFWM6SgWfIPFxPZBj0kp3e8B/AALXgVBxC7hT8Q93wy2sZsoqr8Lhwy3iuH5iW
tey3xxE2iiznkczW5pUe6CA1mDq4rFcgotAtzpiwV7CTwk+f9p+G9xOCvKu2XmNWJbz7ZEjX+KYd
GB5Jcdu/FWko4WIwM9eCNHB6Dp2n4XAPTD3Av6IrFOur+DElO4NCe8f9zWzMBTCddmtQKSYfHN5f
0/hGhpJlX1lz2UHQlXITorMwedGff3jeswCp1aMeULgiynLdb26xi6l8I0QrO5YDMPvFklBEZdgF
Ec2lIzGscaMYkfBssp7Y5LtnQpABBCn+Vxq3DUymjmov6XBub8t0H0iH1jnATsbZZ0orJ3nIegsR
lV8UZ09RZGSz1mnV0Y7esuMBA+mqNvl+Y9nqCNOwXTg4NICCs7LEO3HPE03nHOKi3wCRn5vWQrPe
v8tMiWPOquuaSnO2A8GNG7dvqQj3nEwvJsU/bBDG04cvESxw/RC3wmVLBtNjVvojvFN9ID2v8VQH
6IegO6dl7TrOJd4trbCM77KZhR5QyD5Nlak/v5dMUfuWBPYLPhObnM97XahECm9LnGQtWEu/2w81
H9PpgeasOPVrupkmFcv4WOSQeipjsuXgEyOlus3Z3XvgJCauqKFkq5faTcups2zdtrfS5kLXhANa
WORwqF/wO/+hrjGJCzwnuajzknqtWQFkKIy4bIoDQUMBXXJITBaiKb/Weg5BGCYg8phlbl4Pc4Jw
jVj3TIubXAhC1VCKZ4ovdnE/Kdyd+oNVq8sgfPvkwa6frh+QqSIqldNUt1GjdHImJQrDjfjoeauq
8cctyIqEc23JrR4pwuTmBUq4kNzph9u51xf1uK22soKR5TmOyfNbQLWVOIKfEemePVTOr5PZr811
YagTj8EhHuwzgB3FAQfW8sxE6r8XGwoSFARqAb1BmtioYtaaxfYGtB8ScJyOFhEOb1CzHhu3oFLH
miTxy+9HOghiRGxnQ4/FN3OBqO7B+3GcRms1yKjIZtJzEFLyicz8ZfKXE25qyxA9WiRegOfFSJ08
EE5kWW8EddOI6PA+YKCzzLVj2yB0L5euoovqvvyzEFz77OM8sm1/Q0WKkkrXmt/CtCDQksZKJKPI
5pPvLnfPd5nEe+Hy6KnaEb+6ql7HLc0+n+kvHYuSS+oiQ6tRj/Mq/3HyCfMBDpoPpGuF2MWvxjnp
cp4Zuh2VFBGPP5i90s1wAIEMRAV5yJWcRguO7uDoRq/serfxvVY4IqbCHL7QsvbXPEEUwzKEkxDq
G+iQFSgGXUHNqSR1A4XLUqetDDsXgkL72r7mKzU1njflWp4tkh7zQoHzvAepbvy2g5WStZxDlR6+
IGiU2UV1oaho74TCGrz8zbtr810cGyAyLzG6s/jQAZzwXCMN1a3qy4Ir2ZSDzbcuR9ZPlvKwgrcw
fLVIREVRDSb5wQpvBmGX0fmtZ65U4oQ6nagn9O9XbDLAyPixBLqh6xQH/ytCpyE5BNZw+Pp1/rf+
dHS4jwW2qjdYDwRpwBiaINgWRX+Hl4ZNXgxeprkhp9KOiP9BIbu2Mfw+XJXy9gIG3xyBRNHqKv30
C7PUJfoZyqqDu6+lOjQN1aqYEZrUEP9i0GlM0xnqFNWWpj1RP4Tj/N7iJhMT75N+lSEfblWeX/FB
J0WW6ZSJoZTSQ7Lf/5cKGS+9Vj59hwK/ukdYJ97SD+vkBgDDXuiKEGwHRyvinKTcAoX2E+/OBjg0
slwzbjsRHAJ3AJRZINDWdUq4wS+kIXHBpefcQqBR9HL5aHAqFVoVTgeyOQgn3PCuyfsGT4IOehy9
KeG9KHtMF4syFF+Hh+3rw/u1BqQtHyxVQD3G8QCFhS2JDn5uOgF4irHZiZ/qWR/WnJxlY9j/qjX8
mUha+bm9Aglv2CPEq8XVq/9/2zA9yK3IsRo63+IAf3/C3uM1lZsyzQgiJoz+hWFjHH7B/5u3DyAk
Py7jdK+EfzR7tMfPzMWiMjTOmqrQzupxy25MNNj6HLS1TsOQWpb1+ZryjJqnbDaFSkU1lb4FNP3k
WaSUjUr0JsP1vdG4K4R4IW3U0/Ys9YIIoXKxZDosKAZLsMd75mVIY33EPVb9hoOO5PrnMHiSklM3
ADlbEcw0EqEqxAvt8we08wW/9ak+cOmu3TXwhxSfRiSHBTGPzHFT5o7xIDXi3CSxrrJYL4qrwkRF
yNogqfnC159B0lrM1SbVctWAgnIxxGSaF8fKDQNJF4yOuT5i5l6WfGngZUSWRfwqL2VhtztZxZtg
6EosX/mT1KoXb73rePUmYfmZBvMVxfFgCId4Ge6neCw4G6kyPQ4a5pcFiEGKm5ea4F8LE8M6zCzv
I3I4fwsuNUuoFgHoHli1ym6FLoRE02+hOxqjqHb567BDuYc1NSoRfkx8T0oweR2D0Z43qhbP8N22
PIAE98tr4rJDMwSCUsYV7V6APTy3nu/nZ59ZyL49uMlBaMnYpXU6QymC+b8SbEawVTiZVMQWMH9q
F1gT+8lNWZSJfTIh3CEudaC2gl16oSc22sxohWemImUAYO4r1tHwGWlBU2tbRecij2Lh3Rpv8900
f4ehdN3SRejPlxpEqC5ojw4ZACHW1zvIRzV+UDDAi3y3Yg8lAIGTeqMABiJOxf0w40Y4MM6DqTuh
B0cvhltgiVa44ZBfGrnkEDoiLlaWAYcJLDjXMhsfFn8wh+VVQBFKveE9rYQzgPmZAjod2v2gN2Ax
tG1AMl24qnnk8If2rJdzk8pK7hfX+RYkLQFer1XfSIoXAJOT3JAolrkGcbGK3sePbggYhCOLr5Gi
SEuW9jMs9CMIVd+hOznWI9PmQFUrpNPXIyDYSXLx/4fDpNJ/cc8IjYOr0oH5O4Ii3ti5XsqfwNGH
nDSBKOqie4M5b2BDBpqZBlI8kSkcT3StV8CS5+l6XP2U2epEnPrYGq56y78KqYuG+BA8//7Msj/l
2lGr8Bp1pt3W3wME7LQzsIT/f5BVGZG1ybG4/m2up1jnPLDHqZtz9PRioUFCvUTqc2tkYKUt5AM5
mC29kGt4UygGGfYle5al5FDhlTx4e8Pe8tE0HkRUHBfQvJZNKtfSvkucg8zlTmKPOZrpGfZt/JjB
qszXg3Muqouh9liI7wjlf8ke6CCsghOdlPNolNnl97vsNf4wpPDVbjAIxBkEAoDg/tpKJXrRHjRa
mLCPVMeopCkC470cwcQYcDKgV3Lgx7Lh87aHjpz45TQ6SwbgC+LbVSR/jRCpLxQGY+XU0Zu4p+h5
W4701EaDRysdf303vuVfTwJg8Tx+nKAkqUjyQdO4D7/FTvXQzJYKSZZIVd4ZPPkkm/UvYzRNdQW/
LQ7BKVxD/tUsKr463TolfIb2POZpD19URLDjNvWWX08D2ngeAUTkp7w3erIILYChKZcSpd4mN+sd
CyC62hCVs8x6a+VdNg3KW1Cs6nnFPyACeWswwhCkT7E3NpHx20JDVy8Vdw5udNy8LsZGWXw+mwif
MhqXvAzClJa/DWlWspGQUu4IWte6SDGPObt+EvdTUuvjZehFnSVQR58uNLUT8Y6AXHw0NlwUtaLO
Z7LczWHsky/Fk1Xp8dAHr4Bo7CTSTWQWfAU1EUnJ1GffpphMoPjEmKBFoV4++hjJgE754WjoMzKP
d1r8IZX8Y9J/25Y58JRsKs2QvVV4kaapU1AvQK5/oAKAFrP34L+3EC6J/wl06d9/7BhbKZft34Vi
67D8cPdNZSDu+J8L5tWAia2eA0wkXDFBO8TpiNATYZnW6+UP+/ivt/FQFX5oFGNQW5aykepl/bWo
uijvkOe/LpIn35y5vZ45jhU1AYcNKkMiW5u1GZcW2d1NAnmIEmgACOmOkYpxA1eQ3PxJzQrKr81w
qDCd8ruiiHCE+FKmuFq2bhAsTsphR38QB4kFqKKGC0q8+rylMhjqxwNv8K/WxMlSrTm60jrIGsDY
g+QaCCYBuQxW/sZrHRFE6zHodzj91QEFY6aXpNj+58vbzuVGO781+LI9R8ajA51YrGEo3BZz/LxT
0SHB4jUlQRtBvrdwcWL6bHh0vFUo5LQ4tcBbyHpqwpE72ZVeh6N2gwM63Eapa0R5oqxQ/n23lLjF
j0ubqHHz4goZHA8YgEgcwhHXybisIyldnWFhsodkNKLCOEplxqI148kQKfRgqxsAbDVyNrABrw/z
hUE3ElA3ddx1OI7BVc8idlrx1LeKHDRet9ZoApoWfypyXsjvtuoWZZVVF6TOKl0CJc2UFhBK91pD
iQ87oaHo68M0KerK9f0SQUHO8m9uQMi9pCQ+RrW3PYxTJonWc9fFWdnrs85i7mXkS9IehUJYZ9DZ
0wf2PtUA0bGEHjgkStNRLm66q3UR+USGXBsR+T2T16lOs7u1Bz1Hod1VFfJ0fsCGCKVvihWKS6bN
P8SBImII58QwXLRTQBi0AX/g90/cR8K4pipDHbjQL4D92IeKSNnsAFqlQTuu+Z4ywD+r4wVh5MQq
rzJpFzjZ1EIUyrJXEF0bBlvUxqiQdxAJDKbw20hpGuGvVYDqQMZFyp8zqMIYr5R3s2vSRuIURw96
Iq4c0554fqS1OoxmScInY+gELomG8TL0Jdn7IGRrPaL+04NhY45a+Bjj5hw44lpDiF7kC14NxHHU
E9FlC8yTnpTLSjaXn/qLsGEfobYwWhctoF542wjcfuT5zSKzVExODw3ybqPUec/UaxL8YXzI8g/x
Se6ygPQzcyBVwq6QGGMn+AfveRyVLMeHVtB2P7HOt57un7v6geyN1A1YCp/ufe4AigX4++vjlqmX
Gpjvrt138pVWUnqP7b3TdFxfpq+HXwmkKiBVEtEITEhT8dZ/XVDMRI3nI5+CrqTv8CgIX4JBh/8t
riL5Ex0+OpCXbVrSFJ+FndiAvGYl/DLFiTb6tdPxdo45KScQMIcWGYq/AAgKPnuuzYmBJDJxjo4b
wb/6Z25JRmCbycqvF85Df55FT5vaj0bb7Lfoww6yrjKIfoOcguvr3rOvD65ZD97sJKfR7FOEnScc
ySPfM/2l7HexU/7n79JIBJZq6Bn2Qm5TXcX/Bdw8p2m6aijGK2JySv9MvqgWnh0UeC3bB4ZRMPvC
xjl45PJWrYACEyw9J55U0mZ5eaZ3ZvmzErYiEMITA17QJyh80boU7/V6sPbwDzSHQNHLEKCjJKfI
14UARdFfgGqEOtNWKg6Hi9D0APKdC2osDvXH8QKeua/PkVwPqSGHWp6YsOVwxkFFTuQc8nd32Tqb
1SVq/BAIkMlYcB10RuFU+ARO9e1/BajTDO1bgLhL029Ye9eEUuAXIeY5zTVHRiWrIblAwXjeB5Qp
NzzgteATb+1e8SozqN+2fsRoobCj2eKmAuYWsTj07aEifNAy8WAxxfsTBk/WMCe1GvAj+fcegWGQ
6oDPwEV70u09863Juv2GAPp/ETNntPwiRkDUAlgC5YNCMAY2Ge7qiaX02hj0fw/Xf2+x4ZfLGcAL
DtRuyUlABOVSYeIJfh82zPlDSUBzwVvNhZ/mhIf4FEM8hixL0yGDwryOHcuH73zLanL38WVif6uT
+ZlDd+mMslQeGXT9jLrAjDfBpTuwEpRCSeqO0mFUBR6dZGB+6qaiOpZA3iVe3DWqvxqW+qmTTSJg
7HdFwW5e8ksLC4XH9/xk8JRa7AJpgssULK2R9OFgfN9ZrycOGczwbynM+qg//W+QxiQhiG84JRLu
p8ezsIxvXQoPUSh7r3dVndkeu2DvBFyIR1i/dzTurtFrR+EAaLEHqTsgzq9BjtoresoHRoas3G2v
xVuBBrCVrrTyqQnxj6Xb+QW4m6hcsl9KmOcGkerGxikZcg405/Wf7HLbH+uWKOVaVqiNo1K+oF7G
R9TmyphEoW0gY3y3UXoqDNIg26AynGxvD/yGO35A/daylcEG9NrS4df6qOTVCmPF4O0+egKuyO2+
/dANPQdYuA4ydwU2N3EZ8xE3gMQqTDPMhDrllXIjHiuHVqJoPbeNypP/H0yfZxqyL3CvQNawAVdm
MKqcWjrskGdWSg5vK/Udajo87G+WNnLoZOvCC6nUKdPUf0srPA2pbTV5THtwmSgespULEA8w6pIC
icyiqhNxZ91o930sEWZBWBkhvL+yAWUPoh2QC78mABkZlY23+D9vjHKv5llKhcEF1LXCOXJHfA6h
iFmbH7j9amRb1KyB1n+R1heEqymEEuK/lT9tbrvCmrFpkYEYV4EW3AmLG6Zbv/UfO7vdOxZh9Llh
/Y4fnhoUiiP/ZY4t/D7OyU1Bxf5uPv8xs44gq5WrBQw0g1TBU0xFRaZLYzLlnoIfW7W5ky6SSo3b
8P0yu1dLabsnnLYNX+WNhCM2nZaHpqSLxiSiIrlfYo3X5SMNSvgoM5Mm2l+i/sjh/vLj5FegueXC
akt/YtwReNQfl7Tp4TCnLo/Mt1m0OQ/PHqFu+X8H2TtE7/Qq5zCyaq2BxpaZWqsT2yCES3QjpHbG
2pIS76lda9HLIraY1UICHdSi9Zvt5EYLt+4BWZYxWX1+WNfzVfkEzLK/WTPlabY7UqV5PDUS9lR/
lfgdaEvtmc4r+d5W2OlusB8UtWEmgrwJoL7/IjjxI3wzjFhtlXDnIY7kvEUjViWaDDRPcCUBVHRg
APuUZDjKuCzsLHFBIW7hcM2CUNbdf6iDEkvo43Ry1SVNg5v9zOUttj+1+MIgF2gN6Cs+8saB0iBt
t1sga4JqyUXCsM1qz6ueDPQcW8NWLhe2imEuCBwyZJtCUCw92xdZ9JAEC3BiqEAdNE16Bo7agLrW
wTf1icn1zyDOzyjNUaAu8yFgg4BS0rNS17aoeLTyIAqxagH5Xv9qun+aB1+Jr1BW3LTIxiWWcTK3
JOVKY6BemjFnMs96AJYHvQw28MNDCsS2QZdE7zeK0At1EJ2oUFCU23cQGc+9CClUTERs/d1JaImj
MyLkcRemolQDRi/z9uuTA1aPjSBhGctVMeG5+GHWYWIswn3C9gUZUV0Th3XErS3LA1AeR4LLgVOG
/1DDNAomEcDNKDUgD/7HY7S0jnH/VcG7SesIP/eb0An2+mpTohS0drPJn+sSpkRN6BFQI7uU3f5C
N3TMT9m2rCMRzqoqonZfQgoOwRZfkaoG+wFUxYPRq5Wx3WhV96FLpaE6zi4cnKnZqqEO0RtwUe3T
14q4uFoVFdDjuTFqVmAbjn/okpWvrwWa4t4gq4yijxpOH59iqF/k5XoHlaGRaBmrgx8eQSKC0NaJ
sUyGl5s/yl0gQUgJqy29CzDlgGKlm5vuupqn2/RF9/5O2UCktLUTS8eJW+0nJtP2hGrNMFVE46ow
JvVEJifEG8/pX6ZNbcnX2gkUvolNfPWwWeyhVNMR2+DAzNmPfg/1YG/qhjIZ0rSesYOjBejtSZuu
z3mJlP2+IKw9xU2AVmC/iLuH/9MEB2dVvaMdxL7sWP27IsEd1ZF3cCDfHf8VxNFGSKAy5VemxM0j
dkJQR7R9NvD6I68TY0c5nza/IvExj/dNJ6gfyYiSlDBaNueiYCHFK9Np3O6LNJ2BTN4AElrmZKK0
5iF1daJsclTjmpNuAFLaJG9jvfrO+Dmn9vGND9zqCfld+J12DwO94MAaDC9kPtf4M+NxVjx76TZm
bGwN83RiAIXFWDdDyYFoAqT3682LFHYE4eGFDpy1ctLiviU234tPH0UI6NNwr+2DQq1G3pFdupnT
LV+5cZwjFvIsplA8OuIR51sDNVb2z1F7ocPymRrFWYPb0wEOdFAsBrSmBgqYg9SqD2vDxqlYTEML
x52BedsLbAo81dNzRddIMyA/OW46+qAnxwt8cKL4G7VMW0vyVbGhQKXpUzbp7bt2/OlXvv65W1Qq
nyn4ajc4ppr55lMl0db5wkyqk08+SwioLQXYltaQBWA1x4+oUIhwbB2Gjelg2fb4bxX+ulfsKuFz
oL5+SacTbqDq3Q3EXXLb51URiwyGVxL8w2p4IqNgPULKxfIfMZqjzFIMIfSEi3TfON3JN2WSrCfc
ZPKE2QJ2ZYVyIarkcaQywxmwvh3wJpZEJSY+VzsiO4aEzsMdocukiN1O8FCFljNgfVuPx1ZINLxV
ONPv8POokxkYguPz+VdpQIfKOcukS9xnCquaXniTJ98wKVXLLTvJsogPpjEjta2jB4SgGx7aUn2C
BUSdFn5KiJGIbgF31S+QLL91JkFmc7IsKhei0rsaykwf01v2Hn1Y6AVV+os6AZKQHFjlPCz3uDAZ
W1/sp3AqYttD1O5D+L7cmLvUPtRXzwaUyx+KUQkEWirSJGags7f9L8arhL99Ay5k2aH3NwejosA8
JZvzUzo28C15uTe7c7eZXS6zzsGFHTcXav9aUfyhs9YY8P1xQbLfAv3ykU2Thn+yNuYaXqebjdqU
xMtuOml+S3T2hwl+E9Ys2Wmb1m7HzdaTnG/QW14yqgSINDga68dWVpIC4/VUcRVtiXjO1cx81L8g
Km8Z84fP6yAc2jH3pg6sEcwuCjnY7RbAshfayl7FcAXwaYpKQp5XD2nbnBipwNHVqn1NxGy53lNV
ZDzc8Jt3knDv4OzlzzZlShaGwHGKye6y1AkzTQJ1ndT2nGeTdqb9TLBQSEQiL5882Q7AQSXd5Pn3
0Ojoic+4pRNR20/KCdJFVy35rg80HPfDdYjKNCgr5so8YQQjBIu5fc/KJQj1kw+eV/aQAqMIYg82
jjf1vADSWUIRy7/6IaNKDVwfnTEZhDNu7bAO8cBXypBluWRWwaidgwkn+JKL11PqWW3L1mDIoaOz
Tfd2kaHyoRhw9XDhbF/EmAL70LJIYu1KABGjywQQs1b7NIIoFTw/5ALy5fkQeiE+C1ziOUB7v4Em
juS9cvDKdkexi4F/xt2At04OJDiRh8XzfvIXYA5SS/KhqbhuV+SOHGdrRCeYqgL6e7VwWsyodsJ7
S+IO9NjQgtDXi0KmY9BSV5SzrhrGr0FptgT3C5vQ2PmgWe1A75nxMqjKBnsb5wyPsCki7N8v3ZnX
NiNPaR/OZ9SvOZPk8c73F/QiIWdz8eLHmZmxHJDnDgGtGbxzIu4sNZMylNreZpk74ObBv6WZNAlg
p8lSeLew6lcZ4jqIEj9s9+mLmpcKrgmZ08RM1nghQYkOQxXO5mmaiTa6VY1SFTRFAgPqk06Bg4bN
OhuScygeMsuj8+ZPoQo6nRl1paxJoB2lg2iBmHs5zaQzAPLeJ7Y/k9ipHxUxwcHH6MPFOAUXnreW
HPbaCg9YOTlCf7CpD/IJZ9kIXi02hr8O1Oi59j6hp+9RvCCZVLGVmlSRrzSEtWVKOCMjHedUWM31
Zb5cufC/dEJjRPGc23N5ytB9P7O7PJPUmVTf0zKsyMv05WzrFVF/eDW3l2BqLICBAUxbqqa/Bjwk
QzaEZGN4jUS48s2C/mp0f91RVswF9+QSjbWrGRUSj9cT+EXa2JLkkrbgbVnr8UzRg7GXOvBeZddo
z7KBWxnJQLoLixxwm3u1FrUdVDZ9v4P9jOt0CumaUAUubjwxHhmX91pYoczkROk34gpOcZXmlQRU
b6PZS7WMZFKJ3y7rxkYVA37ze6gUW4uzbLNRQz9N6nhWo2k0TvzMhXMxD4ljCWxgE3TAZ04uhOA5
59D1OMB8Q1CGxdx19XnYrZCyfw7RDrrRpXKufd/N5XUjRr+UjKocoCLh0ZqDCmMgTEl0t0u0OrEB
wetPWq2g01EG4kzA3CBG4waMWEXTx6OKRsDz4W9DL36FCKDMyi9ms5vf3X6XiazOKtFZrQczQqIZ
SCv6NxFPuYzMXu5zIFsOVTQF91GkT0LqJxTZIzxSBMLtQV2HWKcR9bsaonpip8k8bB6OsE5kE7R/
LC0TuJnxEzhkx63P+b12s2LKqTBBv+9CeO0Y3TksWiw1+t6rPmH2ITTVKScptne50M3yK3nodGtq
qUK1PC54QklOpYzXALf7l7SjIolM2l9oNR7tf03JYngaFapRm2XoFEQTk8VyzUJJ30UelFIcmK+v
eoHCuqHLqVpRLOc+YyKj5GwCo+TXb2eWdrVTD4DeayyK27KGslfX6zLBkct4gh/zDol+np/n76Ko
YJnuULeAlYx+zRXZ2bWi8XaCPVC70UmUVSWuaqezo6m62MY+hiLakXxFy55c7et+y2Rj8QR/yGX0
HGCZufZhGIyr5K0aDKukoi5sNuxcFCahJ0l+GwLJM9Q4XP4KiwHORfaszoYaTKCV9uyxcPEFhjfY
b2H1PJ84+49RMz6dBMKnXLtjIfUdTThwK8qWz0AskbI5REjTZwjJnmGImzZWQNhWrApsdc4R5d9Y
Gxprxbw+y/jVSkftwArB7BEKszutBvujl3CW1dOEcM63OpYvPK4d2oGPOTjcxNrr+OeY91Z9hvpG
Y5iCh35Ot62E3kEu7AOI3eWx2trWJUcaioLDYFL993Cahk+8kSTCDRu90BdchTroABBAfSy7IvZO
rD8AZYkpeShwWX9IzEjEbGRpBnskZr6FbyAPSYmaaENVYUiOb7YKSrYA0jwTq6HCb1efoWegNW6D
0wgvBBBhfmajTAdunjEwk+KIp/vet0OeIfpn89SwAMJVhtxdSMSb29QgeVtmehPbFyc9Q8zhC0NW
D8/lvhPVygfW3SAr/hfFo0usUOtOWHXDgoBrUV4SQ+OBNxbjHriW5RtV69psuRT7IzBbxzIqVHJy
7+trpm/VkBj/xAsQHWyfKQ25+u1424s5xRq3wCjLeis4vYieqeOqvXFQ0weElS9E5L1Xmc2A4DyH
xgSbvs5q09ZTEX6Gibsbao9emWgdF3ncSDOIoGrw8Q2W2I1WetYie/TTxKaB08g4WMHF2g58+wGO
3d+jUfdNRSRldd+irh087eFgsKHcW/B+SHd9k0Ta0584WZDU+ZmTuJyJCfHE9eudbboHI9d2Q64E
HtCYvyPxkgOyv+r1B0g00rZXgzfqbVxynKkB8Ye7PFLNsxkwUN54VskZ11sHz3cL+wEo1L7mP2Gg
wrxbZWpQbu9RR5hHkwdOLEYIDk/etyjIiIbLK4OCmZskp/hXQbpWk1jP1d/xDuzOGEwCP86kQG+u
2BEdgLO7Iver2Dn3jWp0uAbpsDEEH9kQ2e47w01klj6hk7M++LYH9KqwXlHo6H25BVQizGtvj7qd
Mr/LtNlvC1OtG7mqEOeiBeWgq5QZP/deI7xQXf9Il8IMh8uamPz47ogFPxYXpk/MusKk38PxLdVS
xX5EWl4xJ0zAGw+sdqoJxWYzR4t8qMB2EDIcSUZNU+3eN1TZZ/6wEA7wcWClW9eMCgM0MWEUWSip
vefzMC/XDExbm2RLDmgjJ881CWfZ6cQC6rVyxK2J4ODDgjzXz4gi1HfeWgkDvGdnoo6fYb5s1bq5
KxJsebNGcXW3Dt0ofwR6KfMTWmvoBHObmgQA7n4DLNF0qf3KhYio2FWKsavLNJDaUrZvZgRWApOZ
1NJurlMecijpoqSQY5WNPOcpYHIKRvc05C63cyLPxJKoDGKXh64nd8WYz+uWtMXFtoB2uvb28RvR
aU4chWzt//0Xvxwj5PeAvY6zE2s9AvVvF6FDuXPNjgC9iQfF0T01EuZ1Uj4KWAfBChh1L1suvaeH
OAUTvW9zf2tT+gfsTIm4U5S1rNj9FfClYcBx7r8ibeOsT3VADcIc8vf7JMU5IYWin08REzX2nBvJ
qdCzp3NrL3fnc3re3JGVVjxdmlEwH65dlDR2ZmkyP8phBTt8WqEqVwl+hrrQUoX1tNbGENRVp+8L
3twF99WUEYsi5DjS9ena/KIna/fqjC9f4hU9s/CucLf88jeoMOf1C6+AbaAzMwWwcsBbsqlHOidL
uY8Hw9cshFyj9Xr0ih0Djrl2dLcSfnXzhfRXyJUToSeVigzTfXeXtH8nVw/2+VsHrzCN4bx85AaY
ayAw2P6wU8w+lecqcjwWCWEPN3tulvdk0JyAp8F4Gd+ZFHNdzpmDctm1nb7y9yDrCwCRrjuexnxf
aHbHkFnQ9XgnuxSML4HPVMc/s6KAI5B54BhURs9Tvi2hnXZoGv688l/vRU9oXq6HTGmvmGmbz/na
8Sa8Gndp4lm94m/B3qMHZFxxaMR9vYxTt/ZonPy/1Ym/M9ii3r/wdnysHJbYd0EVAUyHBaBF3+2T
Zkamd5WzJjfrdJMb2JT0VElsQJFEElapDPBhDTK5CfV31idnrNnkvMaT9J89EfWGur2tq8YrQyss
d472Hn+BT2AZBGp6UBpLkH8wlFUNfIAPdfu7TbRDagrt0iOJHOmp7Ig92+Uwz778Vr0mzBEkfYAa
eqBnu9jaCh24cNOBL8XqykLJf7y4wJK9PhLs9WdyT82LLVd2HipCX1qK7SGcCMzWaTMPtc/Ll3Wp
oOBhZQA+p1LqHHzK20Dsgu56WdOdalsQn64AKeYdl1w94w4VUGJUT4RGVSFEo16HcQtr7djVEnYp
wFUMDkXpZMLbbI2L27b5cPUJy9o7uH33thKCOBQu9wf8JP2383bSxYJqO+Kg50fZEgSkmpZJgxYd
M0Kj9YulnOfmmkhhbpfNGlfUeDqHpjPKdkQvsFal7GjtJfk/zC4q23/lr/zqchMZ/GiQmczZIlQf
ukFxBEwFTWUfIJmujE86DkAxoFx1Q3w0EWW1Cy9ayM/G5ZEmDKKve/zvvRyzZiHqRRmD4MqPbO8T
BuDLmxYQYSDNJkRqFgsghWOT5ZkyoveqS+oiv/cyPhgRqhUMByHzLrLwWLUx3DHjvnpa6ArVdrNS
N/TO/fsg3n9Y1yT5NjQcKF2GPS+zNLeuHAobMk1Wc8jBKHuFdXWglbj/wGtD7hh6MslIgNNNI8Zk
kIFe5+TYJmypwI3p/iMDDSWkJj9VA5WsncH9uezje5uhK7WeRKdzQ3tKeACWAcxRS96ddTuMS10P
ToBMmyjTJc1PGNmzqy0kT+fftx+5/G3RV48RjQ0rttLLnVuua9OL6SADYYvlpq6h2Et3dComTRwR
r6JU0FANe2/NsUMJcfKUrvoXwdwJnXn7ABhxglbzDRwsgaEtee/5+Oqgd+gfPDNVLTAyqXgOKxOi
Oazc9gMdtJwBh8RVgbcSXlMslHP37K7qrBwrbiZrIQpLFHUDreB+cZSHAZiHJLOsWXSRHJ/vAJlg
Lt8UKumal+A48Oum/vGqGbec7ZutSqm+AvuF1sA6o5ndK8/tNN1i3nLMyUpGISxN3ksT9JoBNxPc
d2yvAeAKg6uK257V4zA/k6aQqmR4WtNVuvXPVhc3U2TOg9MnCm8bzNFkTQGDv+Nt7utl0OrFUc/P
22cb8J3ODOnSUsaAdIKd5IpfdFQQKOxi1q0pZp4Nd3atAF/BTQchtZVjuzsJ2XCnHEba85lP+9CL
rut6z0WCGvUlSGlrTXCTXI1sIFcSbA/SqimCIYR+idZVsMOvGIKVvJ84gLd2CNtbWPx3yomWx5WH
XsUsMACtcieftqaTviW6sYiHaMFoGA68jy6nH2ir9vWFr+tHqJD273snXsuSh2+qZwyCw/QJAfcU
idmF3tgIjJcjmFigrBbFSrOWYwY8cKCELsIikKqzpEdCFjfJg/J4hL0bKp0j0cMzrQVaNwS4yst1
j/U//h9aRBSs8yCl30X6Vi+R2ZX39P34P5pcZ2j5C5uCh+tzT8IgKJpk0hkOBwV2CW8fFed0OIYz
8vJbevRKroJiLlxZDNqsswGdmLg4DFzw3yWMf6PbdIdpEcVQ4DHMJsgTslFPNMCrTpgfDyGHcKOY
FwwRE8x1isVM1SpBp5M66eVYnelQnK65Db1jW16q/cuN2O4HQYtTBM3O954Td5rikEDBVTzevXbu
XGEw2D7nwvOZSe1lqYsmGpgr6+YW9mYTK4TD58ABk9OD4z/ERkvwv54E2jLMQku12oBdzx6NNaIA
3pL82ed+vPy0hQzqyWUWsGlAMMI6GRJBWkNrefYdeCS876N4HKtCw5IZli4wTQlZ7IMiZG9EoFIL
7d+brAb24eL3GwGRRWk2hWEXF6Mr8dLOq8FADWk8KWvT5MniRhBcG2+NbAsmZIpLqcowYxwKBqNK
lRyDY3Z5kcLv9J2l4nP6yX76+ynTWpMkF0tmHrFvSsxJKbtw49mRep4SCuy7k6qdAbYToVjDdsuE
tteJdbCS9Te8g1U0N6X+u9EIMMQS7IS+c60Bkc4JRlZMllShLYHHfNijUKulC+UfkOzfECi2u0M/
SA18zDq81e0cQKC+0E2cMSVCJaGRE279lgEEJJ53bfIrWhW4+PfaOFJIw73QumZkgr3wykYCr6SM
V8pA2kzjj05mZXG6D8oWGkjBHcI/p+28fRd/B6GHGQbtqOMTAJyg7/pO2eCXsmzXxZx9IE30q/rr
PJj6IRjciqBirSDU80jx3Ytp+UK0R+/scMhNQvrB0Ffu9wD/UkjjiUPrGDPYoZoD2MnaTWFPgOr0
I+AKsvyonLLGAD0RXjdyoOaUdL4JEA6GpfpIwvtNRdrBgf7OKBo42rl1JUtM0DNE7CLgOUTIVEFu
/RV1zvBvH6QZOUgw+P3Y2ixoknplPfSlxrT+ac4wJ+8KO25ovzrq7n6fHXoR4P06ylvodx3bAoJn
CYRWqtEr2JSWTP4m6d5fnJRFu2PhBTwpeVSPu4xV8C7OLhzvf7IYJGd/Ao/T18cVx+tef/x8zq9l
pDAHvK3pOCIQL2Gnahx9iBI4UzSkgpDqhJ84JaGb46VisDkejzCB6eB/LSF8GH9yEw9sgJeO877R
OmyUfhzShH8ugDf7egsTK5i6vfEqKIIX3hYBgUbAB6ZIz36uQ4vcxyEWdXH1zmMhDEOZQsGainll
8yCw+IBhW0PwuzpiFYGjgybyvPn+L0UY0bJ95C5S9CFG3Rv2w1ISgwhIiSr2tF8fgeTTgGzQ5pzv
w8/TrckTVG5eMQ1fnachTJbpUXXFtS61CV8qpKpoVSuzzqt2gHtVDJibreWs4s8s1uYSzduqT4Mg
Yu3RQpgyvKIKgACBTq/39ja/uFJurvjOa0YiIHGNWtngyY0Fol6ja8NK0OteID08fGJYMjFN28at
c2P1DHRJow25gVvymAVgkYkI+xmDstO1WV1SylCJTuP6YHZr3BBgHZYzUY4ruzK4thnjXcuGCCL8
zubBFitnGmGmKrsAucAHzk+citEqaXZ2PhIy2aB22FnBtcTjyoexfA0MEZha1BnalB3YD+0LbQmr
jKCkm2EJZ5WX4IjzCcm2lQO6YrNPX6nTSAjgKBdwxsppVfkKTyU3xBCZRKtATfuFxjP9tRZO6O58
3J/Z4OBebJkj0RCaW1tj6xBp3SKc2+9cStxGvhlx+SOl77XiF0Aa1ihOR83dN94XqO3+uNYw0UPH
nmqe05MToLrXuwJljXTx7KqMdZTMpMwiIzx7NHUcnGNkR5hN0qrP1kpaLpvXzv6hp/cm5Ciw+tvd
e+BdGh12eMFEi6IkJCK5QLo88AdeG1H6FTSpbW3KCMMZL22+v4+FkNLnvRXEEtClwqyIcTQeVdKX
e4kLrh650qzL703d9HhS25H5T+Td+h3O8zMTEdoT6rHMX9x7mQav/WZSVv77lqA6TtSzUQnQJcNn
fSvKq+73MSu3xyjwnhHgvnzo2nznUvlZJckDuKq1DQb7Zxf9R5WO+oDInZoVqyFxsHMGbSNXO5Al
MCPhNiF38LD1kRxiTb0TUODNoJZdqk8VB9uw9P/U81sSMrSpZ9pvcZ/uHNq8AOjkP19FT+LVai7Q
BHig375bYp0wDJ9sUB5IBWXmvd2mLMeL12zLTHjSFL377BDOFubCsHQM4zS4hdP7fqVsTP4lx7dP
bDpDdINGiCkcAR6x7W2FGJwtkZa+T2kaj/UOMEoCYkSgthc7FLx43pwyk8dkbpkGw/V2OmD6KRMy
yoWiPMDu6NrCdG4MBNXiDvn0h5yRtnYn34KbKhTrG5AnIACycnSQKau1Dmas7fcsc3B7iBTDOiMU
a2PqWdOCcW6SIxc1YViNpTTkNkKJg4RlOmXDze8n7O3KMo/sNtvOXH+ZilfCDK3DbLit6186H3q0
6WPlrCO2i94VavYDAzphf98fb/p+/XRoEjJKriJrKWuyhL+R/vZiBy7yfNFxQd2SQAVwumuf+RiQ
afC/iwkSSP+vkMrwTFbSBADEPaCdNagCRM1QIRCcCKdoae1Q2o4CXLmKQm4Z2l1bSjcxvDLir/qm
FtpvyqmBd8bKJqjD51C3tP7PiTxI0p9cuaOEeo9txw8Qg50kC8ZvZ+aUhKuSQn1TvS3UOON3XQQI
CDLYIyvn9ujLkNvKtkZCi5EFGGJvGrb5jAIC50KvVQhWeOcFkag1wpQRXlW9a5WppjhWqv87ljM/
m2JCQRgRLbmPxZR/s+qRfN628xs25kvRneNudZB1su49nDfleWFPIONrg/aI7yguOwZLYNcNN48o
T7tyYetgOKniZN6wKojHueoYbUBSCRqQ4yUKTmYhlHcUln4di+YpAxuUnw1J8RGiNxxMAmQt62gu
wi0VGm533LpnsPxA6P1vWuAMKpTAeuWW4bZUVZjCXYnBTVrH8UEYNBpJey+mZcZLDxjnzfDWV3/5
SoEwBJ+Hzas9fj+8All+Jcu5GpfG2e/EH1xHVLFhTNrlWJ5wT8do0SYlz/PXFsiAk6aAQa4jBH7p
Y7uITpAgse4bY1KSrWLznYa/xmqaxA6eOYP0r+c2Spnf8+UHMh+WUzbe8AQfzdGVDMVjmLZoI/SG
FaHoi49RlhGh4jfvZcn+K/1tzOOeVHkXEd3m/ZfipmpIjfggXB9JniAqRWDqyO7qASdRlalMdjJu
TTn9j018JmJP5/TCJGiGn3qg7w/OtrV+5miUENT2YDn2Jv0n0cR7VDZrWPYjM8AG0TK0f76d/4aL
9oUJTjfxETIWWTEPt6etzpesrFbvg1Cr1PpFTg+03Ii5D1hEC4d1y9SvgbHiOHzIGY90kp3XDHQp
DvlQZP6+a3Z3T3pA3B6zCyf5EHMXU7v/UTNxH4P9nb4zulLLcrwgDB1pftlBftFRi6nw3zo4BHJG
Xce5H1mSuzirg75K2/YD5R20VMHvMxwcurvPt2731NG0hQljbPTQ3qWg/HaF8jSSUIqrXC26CzXQ
364IqkMdXCzdMsLa+4HLn4cAwwgi/wYOKATfUXNsS7eBEeiCr0U8DunRFRXa4mU/QQU8ZCNzDsYd
ET6xAsrVeYxYsi7GBrhwsddffXMEAiyZvL7ZoW93qZ01tCHqheI3d5ytdlz0EIqy6+PP2QZHlpEc
1amPZBHo8ocqPAlRQJFE2cYvxVZNAY+dElTBZj1SBgf2gcf7vdDL2je1KxcW34SbpTkT5YYYYMPa
GClrhy7d1N0YcUSzdu+ZaEcQ1GeQPaEaCNIsAMP15LYvfDJ3KId2ndqi3AEMGBNaUCNqoHMsdf+r
O6RdsaOWBqsNSBN+6KfRCSciodTYsbzYKM0Ggq9t5q0Z0MTXOoX4wm3kRUYXNjOd47rqAYN1RwvO
BuFcPzUBSuEBKvoN80YGwTr7dBtq1mLA6Owlx8KYpqlPYocktUTSLbPt2aLYI/3XBd1cED+XekZX
yyLoQgxOiwzZ0NTw11OgmcI+w1r/0Kyr3fB6B0HHcYPmtZvTzhJi/Ki9KfRNm4QmLQQX7ijysyVh
MWRQQH6CdmQdnXBNZls7+eRZgNWkXkxVPRtR+F07f+RGiSZVNQbPuCKAFHoohjbz9SV4p6agWYFI
9vlFicVyhVurTybsD5n/hLCxBpxoRoRmGsO37o5TrjAoa7jBCtKxr2jY+uhkGU3e5w4qnYpmwy0p
DThIzoA3PItji1ngNtJSttedtkMqAVS1IdfQIKTfpbr4AdtFMrRiAo1n3MIkviGJwrNZHk/lyj7z
O2pJITuuXdqX7Zlvx9zHia9Ry6HaRocQr9qP29SH5kAmW+zvO4Yfr9+ql0Ys3D2jzBdNceZYmeh+
qlLgIojC2YZdn/U2yptLRCT3tPcuL8qOB02HMVpXFhOvaBhy2vWkWlTTh5QGDh0mKAmn3SOYie43
KoRJys6kxP0T4EYOk0rYcI4fLyU4TQqUwMrklqQRXG7r33D05BaBhORLs8l/cBY+TbXn/t/ziiRl
aKN52LTW8R5fMy5u92V/ZMlrdQ0ZssYQobK7qVUoHV5NdGem4R2xt9wr3xdnCZ0nioLKrebWXV/8
FGQUwBk7pP/R7xi0ULRB7qQ06aHExO3aETQmmIxKaOGbIodn/8/cmKQkvUq74o9tctJKIEp1sb06
fWwLkkjB/C1GZAroomx+otj6O1t38p3DJ/ySHn62FHIf8RVposYQDTHVlsnVdDI3F++brzfzgYtk
U/GTzFdoO5U99LPc1uL0KhvYI25f3Rnbem8BhLOH8pHW5uMcL4HKmw+cp4ZbaspBZO6hyC1wy1Wx
D+rHvYmus0upe3aOca5AAhNXJQIbKaVMk4WjXd3Tke1+XZTM2xL2jEcU/g5xlx/06qSFPfOiB0OZ
ZczDcky1qFpmpBqeC8UyvkJ3//IHt1xaS58Ot0iOHlaMdyPJnRLem64i7SQETERu6Y7wVYf/dFEX
GreZYQFR85wato0MB/tZJ59/h2RpoCjpe+QkIaG6g1u01S6ecAIR/IQbx6lq0t56hxAdyHTewD9K
NsrG+rKwZaVFRielvXplMcOdwFEFYDmHyn7Gb/X7tVV9hIz6gHe/vAxAR8nE1vB3s5ClBKowqW3e
8pxrzK5t4IBk6AP7NoQReBVqsw6Rn2LYRlureuNywwoIIaDvPGRbSqZQCo1ziODfOOW385tKu/op
eGv8shP6+YyFyvivQNgo6Fb8Gc9M3VTpwFOGCF8P5pdHVu4OX60CN7+bxblSCRmcSvAH8uc55dNM
G1cFt/Mm6+hx/UguCv5M7xaHKCw7iwSovHqKV/wTflMdkeE4aW/6+JWS1RvsHWtotDqYu9mkQwYu
PdKEqdACgXU508nbrOvfyCyrxBSLigaS4OZnLxtQEXoKsPFInuOYnUUau3FSzu+qcsK1GL8KIeen
hoOzbgvXtLef9/WEPo+tkawWI7GzYQ+Tttl7p5+PJ1vdMI6xsr1p4iOu+74+zNe9AbAxX/NW0T/7
KndJG/uQjrzKZFHqP60e/1q9SiV0KJbER5KIt74RO4GO/9eAHGH0bnT2wI6c21jrTV+U7JxWRUqE
P3G5Zz4cIOIIY/xGeWYuA6YIdBfEM/GJeMv8PV0p7/eS6vfi+kZ6cXaqCfyqSxp4v5jAv6U33cTZ
DRj44Zk198bADZh6HKt2QCul59BsDXn9AoyYXFuayvbbXG+B8k2+V1jV3tt/SoB6qVTM1pys6H/x
36dxwPNw20jDCz3DYee4mXyzCxwae3AApXfDirFfHrRB5k27SG1MVmg62nRFnJ1FQpn63ZrLQJD8
ijt1dFf3alKXi+Nw9ob/oe8I47uErVrBehVn5JvQvkR3YPOkWd7jmXTgoHtrghlg6A2cwAq+7xqr
UnKMSETOyCAILvJ+7ZtpYehe8bGDO0pBCKv425WXVyaHS/GOWMAmn9bA0MQeT3y6W+xlcpXGWvxh
v8jcoSbbG0X1ZolIvOE4kjjHBNyAX9+8i8r7Alcw9STEK5mgXrppHHUOP37UE73AwzYZexhcElcV
BSWiRFviHCM07H+zxKcyVoUnF860ovUJC0M2pMb+rQCerDHNKvcUgfbs9h52YPpOyD2mNDdXttkU
OoEv0fgI3JecuigMxFy79i0Ucz4sYvc1iIrykNcWs1/J0aDcypNPjJR9WB9aA0fBkdYJRrTnmgsq
XHoWMIJ3MmLhwHPOSJX/vJU+UCeQ0CL91iNy4zyg/K++iZqjN5LBuFlHWlARmAAi9bRSoGsN7zD0
mfNsDRMmUYQXPH/i+tbRhuHxTazTZulshdRIbYuAxyrhz3TTSum2ylbmXQyk8su9uwOlFLRGSFwi
Fgeql8YIRKJBX1Gv9U7VqHCJJv+Jb9ONlE7nssAUVl3prYviTG5alsrpSmKUgK9I98qwT2Kuei/z
Y91IG27tZRn6nDSrO1JBpZMZck5ZLpNzzAGb1GrzaldhjOK157hTcWFwQAZmKu/n9AhLoIb6LPiG
JRezSrKbBx7XbTm7jPCI7rZMl8A7CGhVAyTL3A05T4aO0exj/JqPZ5mDOwI2gKklbtGfriwpZGLn
lIr/VEr/oV9Cis1YQg46odBeG/pYXxV9eWEN6nIMDP/+9E62dqwTCgMegE2a+Cgd+LnRN2Kp4a/p
EJcX+WawYzsgHLRzBTA9OooEAwIKZkJdETpsOqXO7AWEei24hEBX7cRWtRQ0YLoEfb5E+gubsdnM
ekXCEZXfCu6aNYPvgspfupTqRaqwmbF22eTj7POiYUX1DIXTGswPAKJLJfw6h1IZNY2kyiau2TMR
/sOdx6A1xy6z7UWWJa4ntTuFQLXoOFYW2BKSINcpIEf2OWqdlvEpQoH/hUjzhvklE09edySdEwX1
4jzOIYuQG7RAUpHGXfQukozkObQxaQZuRKq4WAUWYZFuTqYuFt4NZiPpqSgd8+87y1nyrbxslvOE
UGFHCZMdNP7kX+JkczyO3+ZvEMdhod2/54G6APY/VxAesQAzTvL2tYqmoeiw9nXa0tICcKtTDsAj
py+1AoLfAJg5a3EevOYBQDuVCOYuhm/nzVJ9/kxwVdh3RoHAtVkZ6BG7u+UDc1tBpl+8xKF/epfq
lPbkuUxLOZOdiHo+3xR+7ri15HpyOMlIfUlebFyVpa2MsfVEDhMWHfT7oFqivw1mc3p7Q+Gdwrji
6Ak2nW0oa4zvXks4Wq90nTGkyUsQllggWPDtS9KSz9CZxVSCmOsf00/0g+Cc288VwDdvDcauyz2z
nE1PnDhWe2Ym5BoAY+mkjoE8rujym5b1wInsJzcfnPBvXdazrcb6FhKziqTpzX9fUeQZoTVjyBIz
tX2uWj2+dYhs0Fv0Xh7dTyurlnMLHPmYuuRp+0mGU1JZhQStkMkAsQ4uaBSP7OrIk193Ew9kpFUG
ZX5Cn3IoyJ7BSP9U0cwHUXfURdIGuyl0u4e67w4aBUSUD7n4lk+Zz93pyLXmq5GEza0HiiejXT53
9JeZUlNWTEJfah28e5A1D6FcMDbANORkHygShrYRAZPtgU29a6VjAt2cS5S8hhx0hKlmniWNu/lG
1yzzcw/q13zD5rN4GzJIUQPZxGhAbIyX9T51jtDPip2ljyFCeNKVHP2Y59ORUuLhA870Uv/i0i+Y
hyI2Ds3rkBvk0qvtMp18cVvqGxp44Q0AG/r516hgR3Yc72xGjOZd6QFuUa5j9udoQDBjxFPS3zSV
dKhTfpjFqY/8ApJrUTstbhpQS5VlUt18pc+B6WHwG8RR/NOQkamY+aqP0JfWU5o8a8naVViOxnmo
cMwYp1J+szypeGU7HAlcmK3MdPbJyxwv2RJu3RYRxL+X3z5lEs/KgEyUlRqifpz7w5IZo3dZHkhK
WqijO2btbaHMFDYfh7Sh7lCfW3fGSD73DRfE5comQqae2TWLY9veWuiAFCf0UK5ViH0AuoenLzvO
9q2pLJ0UB3u8cNxByYfwbCicX7i9w77Zs0ocbommvcgeJvvd+E8ZVJmPYn7ebicd9dF3h787fKdO
lds/HTrziQryX8pburLECOLEHMsLkK++6TJtzK9WDvLy+Ob9k4P1VsXGEeSYwKx5llV0AAWLVDfh
UCcbtBbf9leg7jPGolC/oYTfemZVvNw6rm5ifb94lYwK5GRk5ug4ncpZa7ZRmOfeqB0hUKPZWLez
OkTGoyxhnSiTcuQorcWejt51Q88Fo835lnNqudclPhOK8U8HIHf7+Sb0Ii3CZRT0xPuGx9vPghhY
5oQFyrX9C5P7izDAaRDHh/qtG3387drEUsfKBnNU4z4seDpzx9HWdpWvjGOIM7oFxXMF5FeV7xQz
gEB+Ml864++GMjav3TOPcpHUol99aKrzqPVBK4d9ykShFbNjCqU0/uhXNDyJAM224H6+4TITVCPe
AIUR7VxB6XWB9Scd0DFKJNjnLHSq2ACAqkXw/BpJRFGehSAeELQoPibc53eBkRILtgRMvR++1+i1
Q1YNkAVg7nqxS/rVS0QMhxxqnDrATzD2q3r9ugmBemqkTOpBIgBbsin1Ck0mGap5oDG4sxPYae3i
pkFP9bkh9YeohB19VC1zMZ6dOweYCcn4Q2ayYUkjpCMYAzr6VfCSxBvvGWt7IgZjCuRX7N8PfWTU
s2wcZ96ATTgoJysTDMX51ouCofrM/SfwE0+UFcJ3UY7k+88ZPKczClW7pU1q5gayB6nEcYJYe/kK
zPYOkOTSKIx3I0fgrrYYbK+1ynWpzh5JIBw3KYuk8GqAx/NOXAv+UGWQAVbErsQqMGtRubWZmVKR
o5irdIRd+P239nPS3nPJ9WjkOzSUfBVmL2pwWhivyd/4ZLI/3KgEIPKFoc61SrhWRiexWcW1y35t
cE0xg0jrZbC+k1TeEffVi/lQ4OoKQl4OmZFJ+AviOiFZN0yTb1+i8oSva2RgoKFinV4tf6ZAwlt5
trRf2A+OmJKVU3kLbqlW2ZmuzG//5JhQ/TjN3KVSZX2/SsTNnfZbi8G5VfrAaYfE/qe78mtehR4x
FDCpVW3FFjiRnJ22MTnrvH8t2bFQsI4lVQL+l+AGEgg74Ludmbzt5im/lcr89ZinDEAVa/u0139T
ZwIH0iq7sv2hJv4GWtKY/VDZEKehj8oJHJ22wmKYLiRRF5jl9SwNZ++ewZtwZYvPkSOZyvCDQzuo
pSDlbP/BXNgDswcSYkMt0CdmDzUlkHTkMMfGl1IdJVTbcc3iFf5oOnYJaB90OwNTk/IcD6kayWR/
GerAmaf529/AjW5FnswQJ0pk7/dacJBGV8u3lsN1hkzAEoL/lYYgLCchhrjxGnMD5x5w4gJjz2uf
53sdLJuQxU/o3ZJOhUrlL/K8tQCRhNxgSL7oXplW9tcyHifGGYrzHRToUulbTMDTPUruaj1wskZa
hWn1Sbwt+yjsOMgI88j4uLfd2ZYbDvv0zFVWKnRw7Zl5rqZenV3f5uR/pF3Ri0IM885b+xMrlwpR
IU5CXFg2IkM4imqJBec0fJ9Ii11v033YwB5zwr8irrI+jwC2BwPQuVGDCnl4tOis2FgHig/m8eC4
L/S3/TTBEMzw3UFyeCVoPU2j4ztvQ32XKlxIJbGLYROvg4mCuXdP73Z3RolOqC9GTgzyyHkULnit
VjIuZenH1KFv8zWKM4NyneI4ACpFQ64RUVscnqXWokI/q5jGWNLv55ca4JbBmRbphlt3nWlakuHc
HPyBtpsk6geMnnVMrT4IlegpLWGHUSNL3glraMnIMoX5xkge3mPqZAkEyN+dWiVBKEKDBfogkiB5
loaLnbnhx1G8HVXgTEoW5roCQr58XJBxCEY23GtaNTblPuWRLxoyQdjCORDYtE185il3hqdnv6Qv
A5uY8MRAl7MnJujms3s4J+PPPQcYmuT47rtDRibqEoLOhV0fPZq8UQf1+xOSkTO9Ky8LbBoAvTbO
dejpsHeIMlWqBab43qHX351zy8TZsq/Rr1ZDkC/MLaBxu6XWiPKebUnIu3R43DNpBSG2yB28qPcZ
uJMfgQxQqT7T0RM0de5wvrJ8tLVGJFft/nGG3yYptF3+HNmXrM/Gxp16fwx1lZFxFTGWwwrH0dS/
zAttlds5M9TjdQkq7wuThRnYnlSEP95sOkWAKcuLAIS1PRIciy7OHPXH1JSxV9wkCxZPk6MyhPwQ
bh+tFJen6uqGvw+jfYob7nFFO1unwWqHaikFl+Yi4AN0VOY3umKCvwo2AaMYM2iLwHNN52or0mUT
LlfcnJI/5UqDk0dWTXQjNYtoXhes6StTuRJkSillV4Wc8jO0SnVZ5wZJ9EZ9bowV+iOqb0dBIV3l
JmM16tZ3sUvNGCmAEMlBgindkSkDlyaTLjXlLmMrhPf/aFt39EDKmLJboZ2HMTwr1L+cfepPeeHv
dhQi6wSumzAheUWg6mGorIbgd2MeWwtMBw+oIMRJBIX1mbNb3mAU13c/OsaXgATdF586lKDgu5LG
fg68C3wKymp0Y06mmUTFifLptLqk9kG8J/oP4BUwVCGTTbJ5Q3UGhoablpDVtR9gIIQR6trE0uOO
NVDDVpT69o+K8n2VS08Qtz869VBIfKRwG+BkaxUndY171Ii+6bAw2enBylb2sNlIKw70dvP28ANm
GlicrVjmyV35+HekVHcMnQpMBjpo80bctbauKMiJkGB/Hka3qETQ5ey0W4P/fvCXeHKOcWMDPPxl
Ikw0Edkmgm3jILrF0jdHWQnuLqeme3Vm8D08fM0pcY+deqKzTMZnn16HvfCgjITslBV58c5zLWPt
1xqgjYuhzVExM+WildDNihLlIroMBf0Dc8UdBUvdxh/awl2OCG/XRO4BwJZvPGfW/b84KErPIwy+
ADynl+C9wwiI5to89Axcez31S9bDM+M28aTJ5WEZ6R9qp4b+6P+JQBYjO3ciq+ZE9RhaTp5JOj7J
ZLseKiwK9VplKlMeeKni5WiuXs1YDccFhMg97zuWBaL5wai6nZvCo2VrpJ5ao+nitPGTpEG9zJtn
hcAFVIdqRQAyaQKUbjAnTRDXGIN7DtP4bMWMozXqZHJa/rNp7P+KGoi7zMLFH9f0Z33HwAXK9Pu0
hQ+xKlQUWGI4Ot055auwBExn9jIm/gZRYEBk1ENwngFr+FVBE7IlmX6stA7zqXTIIkEGoA5alQXP
JCcUOAp9tpqi0CfqdgmDRVo5i9U/7RpZbrmoBYgUTM54dmsTgRdtHK3ZrRtgiTwOvEIt6I+AN3C1
W3tv5uTKnQZ0SHeuzx8Wwn7KB+0+aNz12hYq15xicZf7kkSXAwFQYQjEWUshXiEu2e/VzaBYRglU
U0UAH6HVerrn8M+iBbTu2nD54ZXmJYaHCZmOoMLg8EJfDGWVbv34xA+crUgf22uNiRdbSbAOXkNI
WvWFwo2J0u7kDtgS4q3ovsLS7D16aP1UsFSID5EIeVeoFPGQpNdtAs/N5AmpOZBi3IQa4ec9jAYJ
r7OFda0dYst5EJT9YUlIdWABUW7fAnymajXVT3XkcYp097KeZ8UjrYSVCz68sxItdQ+t0wH7eU7k
oCkNitGsw0Ty7aGIHfOJ1FTKt/oHcG5GIiQNBGP+lByrwnAzdCTtNTek40r/lmTcdz2WUwrJRX/3
AGxtquzjlosw+H/qKL86X3GQLLz7q2xIL64ipRLfs9jpmQyEaNIeCv7dHP3AGFX/yS5iPAekHjBX
IzVOgKqU0h9L0KuaxhclWjITE3m+Ia+tVNrZ7OhfZLP7EI9+HtBVufW9YBxfc1HAlywnC15xEk78
Xpa8TjpVzdFyZF4VxEgh0IPS+7U/V8bIU1iHSOau67sptPCW3K8YTZZFnJ1vfg9KIRDcwPGiGo/m
AlOY6EMqXj601Tvfjq8M0yW5cUCd8LDc3PUX1nT9JkoWS721esGyDeZU4EqtrD32ydXyVSDaFI04
9TGqqjtXOlUI6uQgIW38TwwdA/A1i4LGmybdtXFg5Em6Su8keHcWTdSaQzCmYR1DJTS8TUgjMddG
s3NKD8vhS2XZn7l7K00hZbJylSK9T4A4or4V2Hog4Mv60TyGy9BtGyRhDA3NVas9xxGYdMiUcpBa
KVB3FtQuFaDJoAMVw4iE293gyjGvmjiDx0AXpUTX6/IrNh+5UbbQgm3Of7CeTe9zDd7qMamXgyuA
PJDUPgW6I91Bp6Eat6ahT92fWfXfIUAKpwH475Vm77Ewl5qX3OZRlM3izFCb7mlRjyteibULtNWe
kLlbkDE1tF6f/tF8Xx/4bT1O3c7Wcd5VZrJK4l1KDWYQuFi/EMg7b3fVg2kTvBLNPDh78N6ZvjNN
eRCmBPutbaP34qqqWIkgk/Lqhwk6V/FJQvooFSlA1hHQtAtcXFH9OQYOxWY7CbSNBrS9Q89YWNNd
M2KIXclj6VxohjgcxBPKr1UQiT8ghJuoM6PnUm6q7GQ/76ROPXO3seZbHtP2xh/9v4ksgU0iWrAf
+4VyH2yltFrLCVjLkL71T3koIhrycPv2f1UgQi5oqPieEcc7CABZa7LPi0gYh8apzNnkiBareVwR
gWpd5sYqXfU6+jciVD58eNMHzJjQuJgFeo3Xn2s4QJ1UO50LaGu73UlpkXrVVHrvqqENynI4z6Qb
4asawM/m0zluzeMS/58MysrqORFd9Pys84KUd+g2ZN7ImksrglgfloamCEVtVIlfoZAeaj/A+pon
Q6HKsWCigJT/dY9D2zBKn3xiB/5aYBKeVPMxpVBp5sAcVzqveFUdGtQRAMBrrLvSZxLESiq0z2A/
84YccYFKtoHzodEujegMQX40CqzaCy79oG2kSL9n9jdfiyxaTDiQux9c5KSwCVjjO6vBnWMMioFU
DSslSJBFh+8XgbnDi2DK1eQt0SPheO7iV3z6BMQYImEqKWLBHVrQSHmcuVDLm2/t7azJYlljJNuz
MHwqf/HqkinMTGP8sN9alg3nfKmZhR3xCynX8biDpA+odeHhkOijy/K3j9jqOjSmC1VPL0z5JVGK
v7x0CojRy4qE6swhCtRLMi6wD/ptEpUaeQODDFppZGNo5XGn/BPcdbkRgGRLJl0LiJvE2XWwvrIT
U2vKim/nyCmsd5ZENtmHEZ7KmxA7GiSEX7OoRmlSWs5x+3LxDfS+eJYyQ9wQoYhte7RZgjvbitR1
7/nD0Oeyxevgl7UnK7rOPYm+BwAOk+fLohUsSWAsTl2GZFBPsTVnv/I8D42GgYiFM7wA2+KpHUZI
nXQRps6QFWVsJmnn/ncQ/yapGV9m+m+YzoE/bynxyg9bM4Qx/VzgcbRyoyZ8Y6ecDbysQp2YBSLv
L+y0FwQ7eKmkFEa3QoU39hQGcYmyK4XuKowLvx4+3vvs976qRJkSHww1uCcQGbqN8OlmYVB13wjD
mlzaQXnpQsl3zYhfooOF8Kj/+M4hqLU6lcjnSOW2DyYRsOaOoYBYIIYPEJcF9m0tWmHPOSnQkUkT
hSiCNS6HGh+Tkr9ip+itdUcIoWs7D0fThydP7nakStA/bMlNntFgsGiD/1q8Uc+io67OfJM0k3go
lf2z3H5/Ni7DVMlWtN/kiOB4ic6w+efvKKVMsV6pRVa7FwLa+WKG7KIkb5qtdsutPTruJBbleS8g
NYdESj2cuBfazq1oi3jGUpkr9c/wi53vMvMj+1PXI5tPoh6Wb287X7+cfGeZ2aNtppXPd0u9JmoQ
dNq/LNaNQnnrkQjPrhav3x+b1IshzhILKgvEQHnQE6qr9Q+XIP2O29Gs1YdmkSpp99K0H9oxCGK/
d1GD3kSJlkYVpxOba+bNCihN8rSTsmT+1tv6YodDWAVFR1I2gKL/1wOTejzzsW4FVrt/o/Y7UCEJ
8N5kqV3LmC21MhUiGAtEzvFJnFs0r2Owko29WZ9vt26iiKiqqBhyvAyWtdn3de92tHe2mJFe8rle
ckV1mX9JAKbPDgHxZYNvrafr+s3rw4XlW7OYhlS0Ds5REunaEyYVsfBCg4sURc8NEg5a0i1oOEAR
VFTD7uK/6dmI2Pz/cPGd9CAZnyq83bMwr7jTJvFzLH/870kGgtUON4M6FtQb+xHrT2PmpQys1d3O
7qsUJytsMiTwPWnBSCcP3G7KZ//Ngym5J604o+umyA1LaD9fj7TQEIBv5oCbV0/8nCv8/rYIrgJJ
yq4JnGzuug6uuustqMUNfnH21updDRjJXBe36765CmlD/cjn6PTvNvkoe/KHJZh7geaaDDZYOCjG
AYZTeh4+pDH/WNModHE0wOQKyvmMvwYnWwbJvEjDJBOXMiUbu5vptBviIx91IMn57anikOJUdngI
THx8KeSSqBVu3hjsaRopBeamHHK1fk+3o1/INcqg2yv+5uoqgEJRo97ij/9Unx8nkEG1x1xg/4DJ
EoGZ69hsD9RTh4Qd6Uzf3TsoF55K8/rf+b/EN3F7XyAg88rx+CKUUaukQHD2wrNlLVtluhpcr09F
1QTsiotU1cehhQM2JlulewrKMEjdwZmKXAa1M/FolLycmKCrQXAzMnPaz9sOMzwJ0lH2C+5CTEfN
jKv+VJA6snQ6d513/NZgaxO/hA05EH1r6bR6HH7L5NKJ5N9JZ3OswBYdkZsu6y+fo4soGOV9Zz5X
C7wI4TdayVCYU40YtiNQdR5aZZDB7eg2dKwQpoPf62nHXOL/ZhkAqo6bBCOhAIOh8j1DEOBOSSIe
jqzl/M+qf6dQUyXddG2TDAbA1cLob6s1wplQzKnFW8KLbKmN28L3TROKJUzDq2yyNNsqpEx+x/3M
HtITMynXgfsDMFrTcZ7SWxzYKsqSIug2eMSmZfye8TasfHrv6zH5/4kCcBJl2LrjnI1te0zzAzGn
ftl1cq3aI66q03ChicElkRdywbZxAHDTvBXfdHFYPTHSQQLHMR1HjI9nUKIh+Pcrcu2wCTmLwoKr
pd2IawUlcE0nOo5JIsobqqo55onLSbUUciEdwX+kM+tZuc/bn47xMzJlKvOUesKN8ZiwBblZLVqa
WCmGzcqY8HW1aeWos5TRzyKVpA3Z6wsa15XUz8rDoW/SRF6iCxEPB+42sAL41uuQlAAUbhrWxBEw
1xjZmReeTF8EXd/eNR1RqPIyK4dBA0c4CwL96c+HSkrCO2UE1jW+Nb0CMIGEjscy0ec6qHI7uz/M
DVIgdjbrf+NtvqoB0d2rCqKydLGrK0ZwtXn0iKsbyC/HJMsjZFKFomPrJ/IRcin9+liXvN10XwC5
h5Tet3HIrgnzq2XZGSg+RMWQxznyTSXb2RRS8RGjK72JpQRG9KFXqL9Tr6jeSqvZLIRpmd9d+ES7
n4PVYzQa/aVNa0osWLibV+4vO0V924uNvuz/k4oAQcEIdSGk1jZLkAB7jwNgdfnjoKrB/Tco2Z8b
RyL344TUGKDhKGp+5IvK3k9+0tx2f+GMeQ/BIoyBZfYMWWaqnIpCpTmPD+b3OncMhW8j3nLhmfHo
aDfKZ2dz2igFqFxGGUAQJwnDpJdZ4QXrlipN8LdvGE2RrCQfyPMVacYo//Zwdoml4x/L3dUjf4Pv
x+V5QqGMzBFYHRHdvi+pj8eUZDgnHEG2tiqqBEd2W8VSl/VLUQuGOfPTlaJzNbyvkPHsje+yrVKi
ENnZ+Kr99ouNL7xH92CKzTZv6B5B8frRyM0+dTzZk34TeooVKro+wR2+R8uQvoNOq1+PgEYOwvB6
PnEVZJbEXr/9efhDBzSNCA35AkGiUBu9VtIHaqY0rbixVwN0BB6puL72Ux/88aX68vvUxkvFwbFP
O9AIGNp/SdhR44CiflGsIxzkK1RIIwtyzgi4dB3Fl9MAUkW18Hl/dA8BhJPqRG+tVMbb4CNwKCZH
ubVXsfRyZ8oCDTdQ54EoKS+7jGkidIAfkWSErpZKtnw199f2HPv+5veVIUXaLP2Nu14BhqnPhTBb
Vw0FIS0QEKb+Gv7yrYXWRKRqdN2iyUF3HGB1Z/CgieR7uRaACuOGR0qourLLjy45gkDTT9S2qiDj
OcTjNK1t2b66Y9lomvL1KkDBSOwcZVtlRwJNSX2uChqUGfUK+YiUk5zcaA2OYTa2IuNCH9AoJkCF
0X/DH5zR8faWTXK5W5EZ5a8KHhMkXFrRMPDi+7pBdKy6UqQ43gmMORl+8i+6kVfPYDo4BInU/rmT
yHxoJ75Eyl6Os6mTzVVVyIUolAK/+6lv3L2zA/3TUXMUyqTcMFGaGyMtnaSwpGn9UxIglnafvwty
4/VDRRXfCs2fkOcQVtjE5ehpI+//xHgPhOhh9D9KFlW4rLfgnuqRU9ybgAOScBESXRYSLFV5nxRh
bV+ZTNZwhmAOAZv4w8NY9vuupRGWSPTPXmHsk1VIunaUpkqxzuoVskPQQ8VM4NrZmmnVoRiJNQut
1IUyNmQ3xdBgIfuXf1Bi8N8uENWIQK5RMEi0ayqSSjn/gaN9cxmncLLrQ/opjvJK3drvbIY27D2H
0KjFLGS9SyQwyMqqnCjJmydQjB519UjEIntaVfb7RtHrH+feVoEE/TBzxAcQ88Cq4EkpjI1dJ8d+
Yib0L5TeFlNBnzCS5/COJtu+5HnEh0htnVSQL2rc/+VL/5Wj7+iN18yUmYokGatoQsxD7XT5ETvp
W5ce6CLeHTgNHeXMB0mShJBNZ9J7+rkMjxpC727xRqf8DjvxDIx3uP05zdNVOVL+YBdn2vwgJhNS
tMDkAU40AYQveAAXtK/1fOjPZoCde+2kfrk5lB1ILkTjUexJkVhyvu+tKVH/8bj6AHRHZVkato5m
V97wChJeAtWZPzyvmDcMRW8mGxCW0JttlNqseXVlBpiVxdyjil7QzNhu7N88YfOEw4ZuDRTDmjUM
Q7pT4PpGJ5zfhbUkQqsrdTCDYRA6Q79ksnRFFNHcchpRLiXIwjmCcclIdAHFGd1OQow7b/zyw094
FmFGetli6xIOuc4tCfqkETz4PXv3zRGnkdybUTNGAkoSZoHpLAGuIVP6WzxXLapMgOWiytrv28jj
oxFha5zhb/zNpwzvoNb7bnU1dOu9p5c54J4iIGhbM2IA3i06Uwbxq63XpRmyA1SvW8NVUz134Yoa
NK2BkIWyRkPUWCBqIa5X2QVEL3948SxLwf3Yyo0Inebc6DsQ5tmk/27MXmyUJ1xtKyTkioKDxmHv
cM166ShWhkHmtKs6Z18hP6I52Pxg1dloJvLHFgJb9lzpqxbmrZ0/CixHNMTGx9onaTHVv6fm2qLn
LeCa+FJ79mrJJPPwhqXScs34fnOjjxJ8Km9U/cG21t/7ylHw+fSPefjwdnAQv6WqMYNe+beuQLdD
BX1F0371jHSFTOHHeYi2oZnGYxs1kkhjC/l1fVjxjrjgbxsZxxmyBAD805ejQYX2EXZ+4rFBjZso
x8p7dBO6hpIajss/zRb2hYCzzf+mIGHCW4VQ0c7Nf1e132Q5Ml5k9pfk3VV1zcx4XN2VOvAdzs14
JUyNazyDevnUIRdt0VsG2Q+TKicIRz7PB2/ASts8UTD9qHc55GLzVnK/yeEce3Vj7jzU3U26O+SA
Dv+idc0MObypDpiO9FCcaNHKxSkHzVfOdn96QNqj+j2M3GtuyCnH1y3bjiwt8qfjf9518PyNa/kB
dk92oJwkrJdkhX1weetAJQv1fvAp6azGcIzqvzcvR2XGrH+tIvx9j5QD361OcnZxzLQHaP57Bs4p
N6FNDilF21EPp9IeCYB3zeTMOMyeWXzwfq3q1XH21cdZU21ag0WPDaT3nAlFgxpZwAQeDjLxIgjS
5d0NFSiS/lm22wflIo858DmcuGGI/7trHEvRDv8Hc/ncLbWm4vvQNzWfPVhJ2+fX8iAiREd7h0f4
8RsqyzvIbAba2LMWjF2Er+/ihXOrO9e0M80rKvlPa3Tgsg/Q64MiVElzIX55AXDfJ06xFJ7hujWo
IVZHSakEpUo8xI99go18M5cjtH0YB3P4TFkU+6VrYX16lM772ixCOmtHKKl3JiVI8HGGQ9mUgpPd
B0WVIYOIqdWZ9QhJuogweWqf0tZsq9WskrKDAemhODZEdFPe5WRTNIcBiuCqnBQcBH+B3ItmtpqA
EDTR7/8m1PyXbJFA0sLy6aPMDZpkZGIGvHvUgsEczx3hVuIqjB/Wpd/NrAqVUpwzeZru9ORrYoHc
JvC2WVGwLDjlTiqxs/55CDm0Unll3kZs6cfm+g9OgfcgGIE0k1syLm6wW7+crnxDAay795UJU3ql
B2AS3d6xvPfAphnFJOBHxbT543ZB+b7Pps9W2BsRoWhdNxH/iLlN8wfNp5SizU8E62zSBzqwagmA
h6Xc4JCUjX07lwKU6T9P1SVt5frg4qjauYh/qXjB/6hp5nrHbPmjZW14i3wpPHEU2kwbltJEAL8p
2SFxVSMWcmOx41AA9fB+wiKjQyO5hOef3vHVudeGnOoQEDl4p+iaNSCp2HjfRc5KdU5qEm2GzOH6
eUyfU1xXBQqXfg1vyHhNQbSCNvgvCNGibCNxx0tF0U0a9X6fig3nStIe5rw2VzlulLT1HbDKEd98
s9ZUZagXi13t6pVMe0qmNJHRVuhCf5eaePvk0qTK6oYnFoQq3lvfOJuF5DilzIWRe5qYc6PrLR9g
4HRQNTxB5eu5u9ItmcSBDY2pSoLd2sIb8DvL/imXlRs4BdmO1c05qJaxgGqzThCv9nL1aKwxEB9E
uFBqRX+7iFqOrMgELSQtEOdV9csralJ++vCc9ct2hn3++WXJ427bmTui45JZUBPEWO8sZtGz15qD
DmSOuTVxFnPFUMWIJaZZdeXCqwzabcRKSFo+Styqu9Xwqoa1LTCRyE8BmyNF+WW8kx+1rQM3TkIc
0LY7G6ZMNbhUzyHXK47iSwncw0Q9pjJlVDWUQrzwQeY5BZvzDktwEbx87HFwuRN3uoy9USReFdpC
KEqqijxz/g01YjJNcVlpICTDAMlO4qOLmHLJP5t3MYLenCVfDfNJThHpj30v/pf9Lfqo00lYvVwS
CMCqjxKpZs3s4sT+TUS8FWIRQ/Sb3TQpkn8/X5jMp8/bkMwwITqNVi4vfqG9WEzcx7yXKYmITUMo
rGFOrUCdra8WUIQLUsOTjtDMUR5i+hKeXjUDO0ToYdX6pNHk1dY3BxJySQ3iS7wl2yDOR0t3Uw7Y
r29Mb6z+GZEtegD3t5Bz/GhRM8L6hT97ih0p/9bviUvY3lX/WLf1Deyxp7pzZ/kNI6V/BGqgdXCx
8GtSPiZcACBRFs+S9t/tw3jHTDUo8aHUEzaP0mt29IKHfO1rgRy4FogrHJyiEsYCHKM8n7LGT8k+
ExqVrOalSFYN6YQXdWPhMVJ/Yt9d8BBRxaMID84WJDGRBHqYjkRnhexpj8zXj520SgcR4LHzlVKz
tqpF18Kns0GNXN1Z1Uf/5nTVo+rjg8pREQVqxGQ5QwXmK2HRLMAcDLDXdp58Nzhy608NXTCTQQMH
DIb2HnQk+mYl7MF4BO4KxMl31fEPVIbH2OMO+c0XJDDJqkZwP60X8iXkhNFgug3lETRTECCYUCPp
ZbhGIxovwWXtNAytoxlrm+fbsOdGG4zUpLz9rKFDTdl9E37pmzZvlKUg5uuqOWt1MmytPAqfrMID
0YiSWxdkdVuoW6tYniCWWli8sxIDwAqkP1uiwz+FaAuj9d8bof+aaqTddS7nIOrWzc0ZgSdir8zo
iL13NdVtNAzHEf23DBeVZw8l+kvJH29xJ3BxoI1h5iuXk5OLYJItSnlF22prohApYxOi8bubFIBZ
uS5cZ5Kcm1sjwnz+aTd34YU59igrs6WuXTNAYjPNdwTmvHw6b1scsDobsPnsuI1PIx9dRCCDwWD4
OIEb1+nv75CYfk8GysGCblqs/KxSQQxTEuPQPLVoCiL9iF9rdFmXFXVwnZ2Yp49j5/4+2OU8PJkW
Up8767nKbc6273cLnzYRomradcGjPxjWOERAqbTDB90lqxZjycHRIotl5IpDquk+LdapQbXWhJJ+
6NWr7BMaDO/TA5gxiAf+N5XKG4NTlO31vYFEOBFeqQSDV2aqDq7Xa7Y1c5KuFAMDHQR8ngXFVX/s
M5+xpJxODumwUFLIYilI3fwcePMXwA6TPqeH6h/ahGj712fSH5hFpzm8UZtpbVlYI8vT2oZVDQiQ
zJ65hzPDmKfGyxONoQMW/EZ6dUgaKZA9LwWbj7+O4i8ylFWWiCi6qIxpLHQ++tSUUNWNpvMmSkSA
SEBRyMsmFjWoNZAbZlEvSkGX1tBsxpkIjA0vO72g+syLso4ZLtWknNcHdCjgp8yDQZh1cJrDc2pB
CLIbb4GcsKqVH1Htc1vPkYyQRBqHFjx8AmjRJwZR90StjNlIzHIKGHfcGqkSOfoMjurBRJknq0oN
S7ScW8ne7AjC9yatzwZkpU7QFATlNt5ppj4uXelaCUF4/b73+PxPM45aA2u6eA6jAHylN6TN65X0
M2SS8izXCRBbO9S2G4GtohZs26oGbCNy0Sj1YseWWei3UJkySlxgr36bbxUIZ0p0ss0GHXzll/af
0WyPzoT+FHBCXh/1qdq6Inxil+KKp063PPtEPQf1vBeFyYZSICfr2CbJ5J9g71YG3v/Iwj1cgpop
NtfT7KPoQUcJzTbnO0I0zDT/cQ3rmDAflkH2tH9mIcqgEfwMxpe9ReypIoID62YumlJIeQcT/ahq
BwIpM1/6cCp++WNP4rOblK1bhyNny3cuiDXpk2ualQZfErA4JicA1DoxvaV4G5mD//VsMX8+8qx5
QdEkxbn8HGYvyzaepxK467xX9zd6Sx33SQdqcL7eXBAyNaeAbfhSKE1yHJ+JfeV1Bu6fh+tc1ViS
FkdoUAP8mrgG0h+AFy7qjdDVoxy3aQ1zuNI1w6UcWZQOq3SP88wWZfs9pJa0BByjHhXOGlrLrMKQ
qr0WXNXoCjZzi4JV/YGGne94c/AbhGNvHV+VM6n5ViMf+szMc8JeSEj8HnBi2/rNug210NlHzYCs
5KbN/v3Oew52it7r1DawTPaTtqIbsMcyTr3p2QGiUNiqAKnEiKfwMbDVJXTv3jZjxZWinBhaBwKU
kuZ2qnBL2mAq8mbFmDp+jpY6mvbZcTanUOEQEqtPn5BPhMHLksLZ0nGCdhU/VD5j/HTPQ8BCmz/U
LMXl0sX2rgMlSF1ysBUsauOxEZyxzNMmHehDzYKDuZ4bwWoYuT9RRUbLrhSE7PmH3NttiUuUTaQR
SISDsNNg0RIF6NFNNqo/8A8zruhLlpkLEcqpor4QhpExNn9pRzwT+mD3YAEF5+2XphtwXwNLQssS
sv7hDl5xQS1e7qBVFyQGcFBxc2NQR1Mm6yEoNXHCuoqSVgfdVzktIaPIZ+3NziShQ1jezumGYGyj
KXVW5SbDXLTTxFprKvuub6Z1iQz35wITUoiRE12y/plODl8Vv+9II3kvqR3Rb4eZ+4bvNBdJpwQI
RFjLmTyZE61q7r6Z2YimLrh/xEMC354I/6Fg6RWvpaB6pTXpseq1iejR96OjDguA7XkVXqwF9Hqr
E4RUv1HMZq6aogdrdujVDYP/xCbgmfMc129YLfnp6jE2Yq+ihOP6VYkz59kpiDuvBfp/zyu5cdy4
JyYz9qdalEJjRUt2kzylZZw0JqErxnvbVfAVKKo8k51IFWgmcdM4xBcLD+6BesEYmTHXUru1S/WF
5ZoXG0+o00VhEJVGg1kO1X+T7Vcr7XhMjuag1J5a923k+UXBNIlkyG8DKUuDoIM3j8z7cwDnwrU0
FhQ1ua86R747R35FfVRCI11pv9Doo24rUFopT3HIWtjEr6TFtnmSC0SWg4TVxT5l3TAhZlCkKBCY
SDE1CCngcciH1qaNLpm2snOneilHyy7VUwhJnnL/EKeRnprYRrOKans5FyC8z+ZNF7fIHykVzXk3
Q3yWTDASVEDRODyHuLEmQJ0mwKdD+qOZYiPGxa8nCN1gyXZ2z0vLSKMtQkde2a5lYVP76zNMLbUr
TKCWW7UgF7yE4Oq/XBVQb3NXf39nxuUmQ2+zIxd+M508mwKrmXSoq8BZEj52sPXKGSQP28gNiOUI
FOaoZ9YvPFSsuv4+ngkYvURxcB7AR75dv4DvYV+pnjqIe/ygziIvr3S2BjdaWR+OUG3SjJIrnh4x
tYc1dQk/QYPspTDcCSWpj/DO8y65U2q38m1Z2hnuFOCn6XmkD2A1uJz8EL/Hnsn9jKSk62ci8+h4
UEiTORAMBpMnw8vt5zvcvp1hb/JhFCzMDNMDhSpdjA6cDwqWF0nj4s9cxaL6a3TCPAq6UxVZ0gvG
wGjqN+mob0j5gveiwaL6IIixyRln+NZenCPDBMWSEscaoCyEZ0vWe/jG5pazvY/zUfRVpSEIrbvB
NYlDZf8Y5L56trJfVHA775NCRit2T/kCcJrkPXUkK8SOSDNOzzJypuL0QZeaGn5nRaO4w1ZCougp
kxR408ysGUGx/m1QCUqJlECEMhus6FQ8x9XFXjLBYcliwOBKM5gV+DHTyh0c4QrklhfnujyeV0i2
556UC/ryNX1RC0WhuZUzYDKkChcd6nsUTrQ06569FpU/HZxzSUFD64tmIRUJVrbPMJ2wIzTTfu9O
OOhKmcX3r5yZMtngQwh/NIIxXU+C7FG72MslptKvmTjHelcSxrRdjuLN8cRZqdXYNv1TD2f06xzX
zYq4uIvoEMBCqM/i7VZY6SeNryOiFWWU3mMeaKVBwDO+9/6xHfUaR2q0qEr6jkru03kaaoHHZpP/
y3578K9HQHWTNQZUCF6gy1r88lyU2k39/lE33zPnEX6bUWfkL3U1lsh7bnHxPZOKZuaiX/8Pe8Rl
EsPugz30AgsNK+XkMVE/kpEu1dUN8ZnKu0wStfqFlH3tHoY/60DWaNF6PlM+5TYpTHuqNN0LhEzE
mKhAf8agDtN/dPMnIC2hXtvD/I2EL1I18W5kSoYZNnJ9N1olimWmQzoxFP/xkljCWiJvA+QKYE+i
yxm76tuHhmb3T6cmCoynMfrSnCeTuUwFRaGPn+So5Kavmfz4bbywCXOOe3gWM9xWIn3i26O2YYJO
ZdASTybfwrjrw1cTmkXyeXNA/FokDq3Lsd1I8xG6C0zJAFDmuCE9naJoJBhXkuhI9erDmRsZXDET
LPFgyPWI3WPIpmOjVbDDraD8N2PZ6rIHetEd8onIzwLCwusb/ho40bbf82plXMq8pFR6HvBGdf8/
cYl9YZbmozaOdARuOod4Eaz8xHgAPbJaddTTVuutJYjhTD+lCooz2aDuE26afr6UQQhcMXZFuRaA
K8Vn+U/YU+nt7b828OuZNYt9XVreFtX/ieNe6xsdXkX/F6AURnZ8cAU/ZNgiTUuF+DQ7PjoIoCta
Gks62fUeML7/1BSWIPJvbUErusGX5nzPbbprIvICyosHYkmmYNVz/c+h+OSiDfSsZwC9+oh/MlOF
xDO/sy1lTDpSKaHi5QzQa1MNP1b3HYV6g+G0ScMjxKzUYAi+Ig/9rEA9cbsxg8uc28BGEo54RFCI
dUnqi6Nv/KdGjTCnofqnwmNd4oq2ABoNv8DyYHXs6F4J8nAFwTusgcsNCU3IlhjFW0SMMqpPGzFR
0eSW9NI4srcU2X/5I6N/dptBD7fg6EX2JOGEQFU7L80onf08iV9hTUT6rBwyvjAuOWJjfVn0nOKQ
jSDj5FO313Sw035Jb0r5teMOP8GtDW2NZPyr9KTJHnUhwoqHgHqwuF4aW0uc76Kak2WdD1aeqxYh
2IpHTfQw7GCf9zLgrZv/BQl7v1j9rSw7zZSDFHB0Dh88wzgHVLQ89N+cIs85Oh4lEiytt0YXiS46
2egfSSGqFgMCclomSh+iURHSu94gpKY6RqaHBorn310P7ULhhaNRVX6OF5djxP+OhcybbhNzVRIS
/Am8OagvFLn+NimhKEUKdR4cLuev1xfgPU+XhidZlPRpUKWjY1qDV+xczLy3hGGpUDWDfdBTgha4
i60m3VhL+tiqNYILyVwW8x28HvcgLoV4XLsrqWxjiMkKJy8xyhNPK5s+kfk0Gttm+/p7aTuYnZ85
CzhLNmAvIu7PGBfWpawqoYY+TWMMKhvudALWItY1ZMkjLtsy5czpx5sIhJky3YYa1ax+kflYYpDu
W6YpBtx/I/wpi4ynK7Pq1ldhIotibpOwLAmSbS8dHdeL4UUg72lUM2lg4Q7sHmyyDzLcbdYV4+8K
+abzqIFVDP7fUI5XOZEU+WOyPVt5jZr/xmf1devYZ9uf4IwER41gaXfiabiej8YpiuGq7IvGYx/Q
GsfC7viHOHBVZ2AtwVs0QtilB6iHkLVOw9CsbYIv5SY4/BGeaCZXkiFVGABWU7/a2Lprito4tcsD
bhwIQAC9P+Ao9Bwdjie1K9QThQe55j9rUCwSxjGynInjYa//ZxYh0uWY0HlXlxnrDeek4RMMK9C8
80yS65OXnb6W13t4ZOpRttV27qWjgRx5igETdwnH8okiaMZ5f1KpdL96vDSdSNLJjqKW5I3Bh2bw
0Z3x1/2poMDYdNDPNxLsXkTIiiHfP+DD4A5QFroGWlCAMVYk1JIjeEoNICleeEJl4+qBNRf8orWZ
xUpR+QbJCw1Ro0Bq0d/s+piRfVHHQ7OuQRggYgnZAk5lahLN3HX4gQTOXDv8JLTEX+4AMY9IAt8l
1WLwkKpQKwt/+do92+ItpxFwb/QiZ2DMlY2okbvywzwK21DzSBNFr10iotzySTb6zxnEpGZ9oDhb
/tnCs/2C339v6XgSc/RDLBcoJu/GOsZ7fOteVp1+hEsru3MJ0rTORcCAx5Icnw2B+28AiMLEnc+D
u/Y7PPRd0qj8r28XjgSbdzav2k5rQZKpVz93UnzmQt8QLXX5CWXHYb8VGVq6nJZQaNj0HX8OzbJr
phqQ8+sZD5ZPJGYB4zsWihIJGJjdzyoENg2zJ22L2PYBu4mWDdUMNi869yBP8ErmtIrdLLBI+TgG
XkN2iRmCe3mWb1EoYoTkeaek7gNA47lzO/c1qX6ktFf/R/zVv3ReTlyq9BsGxb0MzzZaGQCx8hzO
b1OJTGIfwdWcuRRKxLjBxRxJnguox9duOlYokBSPtaVhZ8aihnba7KxhaF5l5umC1C/equYu3wn5
6bRE9+FjnDMIRVT82OiGCUjwGcTB3hk+XD3SQrNkMzVv2rCUFgDU0wS2G3CS0FF80dJDVLRmbdAP
rA7A2StG9fmfRF2Ng0K/eZKUxOTU8Uw4EC3VmyKOzQhKApM6mHZOxy+qY02CYs5sNjx9fKkwoS5L
xZZXO36AhCydK1yOYpVTTcpokgt7J+QAHcBW4eCwtIDq4sTbrbdhB2kns3Ws22DOFl4dbJvvNQPq
xCSrxZyS7cK4YkM8V72J84TNXG35XnJfcIXZN/WW8ONu+VAnyCLXyj53EtPDPLdQxz7QPayvH21B
C9a7ppiZAZi6vJZVDsobY4oEsdHRaIJl8rHwbWHVxEpUQYUi/6MOF5rQDKZPk92cIfO129PWQTpy
a/9bZ9GqNNl8DnrQXVe0NPzRLdNpl9IG2FolncOqHVePg2svTI8ZyraVvtT7cs/5R86o8Y5x4b+X
f+H/YNtY/DJo7d+uunqRN3XAXg/LQwYnK4IsYNTc1ioXWM6bt0afjxQcqSsAS+7wKAcnPYdDk8I4
xhXotnKeguCBJ+H2iqQVDEQl0Li5gn1QsOKI4u8OYcn0O1nXxoH66QDu6C0zMf8fTCpLAH0IdTP1
5vFq1HHuE8Dz9v3bqL7cuvsfHC91gKkusNb1UELFLvAwRsC+TaPrbgR7/pfEKCBqCmTuZmZfgoYn
0gPocM558tvZP57Ijs21Q0YQ5Q0FIVzQiJAu0j/3ezNj0cT458ZpLimyDw8J3Pcyo/WF8IHEwOpN
JorifSYxkDkPN/NkN6UcbbKW3Gbv3rI/jbE5IOwUMC0ZLVFwt8BbhC20O+RNoYP5NI8gEcvaYmxJ
DXl5TPGJeed5wJOIrAzgthaGOtO0lHAmo8dzsyu94mAqGyo2A5P4XOea+qiYjiFf6/ccosOH9exs
4hWdS+tarMqSS2SXKboiPtPL2N9VT/SPEAHRfjrKnEaGQGg2Plm2VFusITBWhgwDJNNZZtpq7pMw
0omjuqkuKMrsxiZRE/fzFxAGUBWeLUDxA7CBeccyVnDfdXYv2iKjsdxJVXhnZmhN6FIn1b/EMuDP
EAwGezi3ztw7v7df6hJ8hSMX9hBLHb8DjHoVS+BLl/oAHujeZ7+4nH6xtDid44J3ZdD4VXfAA3wq
KcsFMzVzfM16Xmltmq0wKaxwpo7RMLfjNr/ati5XJBkB2QnobACm4nG83d7/3jCIBqo0mr7Qjz7V
SHRUxqXV7Ghsm3CxsUfKKcNHIZhTre+pICIMgU2qAbLycv/6+rZWNmVaQOqJw5bZPga/EDWj67fB
GYKy9UIR62WqFu+m9pQUYkJHCP8npsi3yynrBEpUA3PcBj1W5yQ1EcN8yJur7I/KtZOrSKKRuuSm
P1mJupJIPs0p543ixTAczuHM1I+bwJIa2D0QIGk/wZtW5zq3M0RZEAkN43At9KXUEHsNpxdh+DDR
Nz7JO5NYMofoaLq/dsrCPA3m0OoiyEV/YyW4aIMMGP5FuusTc/4A0Ec6HrGWcN7o8zfKT9/8pele
OVd4qcTxdlYjSiXN/9QfJpRlfbHIHvnyACuvUrqR7GZnVEX71ylVNwYW8SOks5VeODvMkQKthMEB
UMsMFdsMIWQT3t4swqKrcUcVom4ZK0Npmz+lnrBop/yjRQbsA09kWScOT2f7IW3kvb+eROi9OFob
OrAXYigMBji3v4EczV2r8nehBcn/vkS/Q/k++P5yhrjVBz5CtouMr4rOIvQO+86JHr7CwXzRmHvS
C/nzuONUnQzqxnfcaKWKCvduw4T7Wp6TMVfTqle9ZtMnkzIfrlFPE4Epv3qSXiABovORo9348JFB
nDWvJKqtyRyatPpYChesvK6FmWGdAdd3Kbpp0yYRFYUa0Nrcu95GzleCQ86KNUux85HATkNZKEFn
1fj4B075NJesTE6MmuC7Fr57lboc8BZBJMmf4YFQTc6fEd5BY6Spp8Ra7R32W6xeCSJCRzBhrb2n
7f+Ao7vMfb7eQ/ns/ecVKzA2x0mxe1ISUnjRq7M50bY3r6k1gVl8kAqRdQbPjZqky9irWO3ZW6mj
veTC5nZHx7Y6ndmsnYf4oiOrXt/eMKojPugDiW3M6fzlswA5CpTSlFD6VRRrjjjn/rp6pGi/ro/T
CnjgGyKjyjNzNXp0wl6ml5Te0FNnm4+SVXgU61/a27nfzVf+0WwNldxzu8hGLAlXijoIuTN0FqLD
M5Gyid/c4z1rVaS6g5ZkJ+pGHEGMk/GBhRDN9ciluTaeUdjxMUGnFcq15Q9Qdf0jg06CvIEh1OSd
abolc+btN3DsO7awqoTUx2waIkI8WyZgzSWPRp9mAI1XztnzwwI05tI0eaL9OdHVBgMwkQdFmDt5
OKH6ppWRTccBTO92Bla6nRGHXXe7NwZfzimm0Sr1Dkz+T9lxQl9gZW2vj8Q37fe94PNfpW7ocH09
05lnVTI0NG0jMn/5tL308nnBxmXPKMQCQdjbwHKrYlHnGrXmOODhaV+d2bB/sC4bR1yi6bn5S7FF
dBSWxZ8CtdB4n98vJd3S/u2jBAZtcab+dPb+tsc68nZmgP7F3caenDGO8VskzO7dWUSaYoy+2MOJ
WcH/AaMG3+RAfQCiHGH78Oq251Rn9/NoKsB8nZ1KpWIxzcBzhafTl0fmhcYam+lfYtRVu0DSmINO
2qYgugOuqmbOSMYEq1bbgNQFmUD0NN47Vw3qGl4MLbp0pnb4KN9/ZjGXj+GjeHaMAjp9vEgegUNG
yvoQD9JZyIDakay2LNdC2Hr1wMsgMGO8LLCCtkRDkVV3YAsYTM827TgbrH/ezLunCz4ndbk3FFsh
l/6SOb5VnIyQRrAXhzIXgPxcPETAGvppdI5iZ/TwB1g2q6NGyHzIFNnjXRkiBKs/b4hxsIsw81lP
jGbE1bagJYq+HXvDypI3RKcoUq4/sHy2zjwq9v4Xkelyxp3ot5EBgh2ysNuOCVDcRWlkrP0ibzNz
wQxhTd3qDrAvVgf0y/xGlHJTwK8oXQhtdKz02LaWGch2ew4qm6gRDGfaEugMpBwY+T1Hs5Rhzqke
PTjlmwIfiZ+ZBF08cmAQBKC2A97BZUri2Iac5KKsOfyYFGS+UqWfX2KPKF+jyO6IwjLrkNv6jJei
DG6Ym+wIEg7SANOlLLSBjMIVfmDb+8OF1GsURoRLSGBwlBe7C17BQPrJULpBhJu0DDFz4m+SebOf
9ETEiXA9sZOcPadbNfLanwAQzyXEms+7KJ4b7aH5I5uBk+Lea3bJZCvEbfc3wtGpk7rWGn0uoz5n
8QICPhedUbu+nyiE5wsKdVpFTKFMSizgYzphLFmumjYWtXyazetZPoE4jooOvIeWHJSzybxJIaBz
dc46WwkruO/v0HW9dJiNKGvfUn8fk5eah+RrIVn6sQ7uReXFCWXs7i5fNOdpquRWhsVBgxOlE6WP
7kXjEDilg5ryyrBWXHQU/NdWhIpYR4H4R2XBTL5eBFHQ6h+n9JmGATcj9VlZpVi+Rf+6JsvgiNzQ
C1d71Z4MRtSqJbVf/0RmlA8k2MBIKh14r/PdgUglrNboB4mch0mbb8AOL8aWLoLO7ZrBifUnFvf3
1IY+QhSCWLXgVL3M+oTN4YFYq7XAKEyxLrbozPMH5JBXHRKa5MEcfemYazhXcnEXJlHZ3a7p/3nJ
xRjRaAYUll8n3vPbXfQXac6dgKZrJtxXB+ra1ZZF7kS5pWWSVqHv7pfEisVlXTrpvFC/1WN5A3iv
7Xi35ScRgVVCvbPRoucAY/wbYM4UmamEgdY+6V4ak/InHORrvi/PfLs2Ne7bXzipT6mmY2w0GZck
zl025mrKo2dw5i0Y4v21XsS2pZjRFH/em3CurJdUuGgvc1fhW13SasLF1PZvDyXtVU63X6S9wnR7
fmfOzz9vU1l8yay9rqUtUxXK6dFFSI9ZlZ+/CPWOFtwuucSyr33OIOSmNxrHb0HMCH7JwlklluyW
J1eWfUGWfeQaptuQBQTnN+CIdPG97aFK//L7xVOHV6ZQpYDVcoaEdwD+mqB6ur/XATVEyF6xlVMZ
BJTIVc9Ja6ztW+LrAwsgiVdzXaa6M8644MWckGPfuHQi2mqecMB0hp0qbaCs2/qRpcpvyaCzwt6k
WdvL5wX2G6ngRZ7hnNMEkBV6/73eCrrN5OOoccUh6awDRRAp3bsRFex5Rp2nz3kv9/aoLcyPnO5n
HXqHMWbKymDfYcvK/yAXDNjryfEY+EC22DqwloV6QzoiEKloqmy+mpO9dSQSNBqKcDmlohrHHM25
ATAQQaFHG8JHqcj10mH4974C6ggAojyfn6mqSa87jPx646fEt2V9nQipa/6SrT3EBECIPPsn4Ef7
RUq+pjRmaVhVtakist0Hm3M3K8oZSmVIH4LT3wM1thCNXn0Fs/twpUkKu/BY8PGELp9tD3qV4gqo
y5u21JXC9vO0JzlfM44uVgqkJ92NIWDN4CcZN4dX1ZoxnRQ8y9z/+N2NStJVFHDFg+n5lbYvtO2o
UZH4gcIk6f/bR/mg3nJfs2nZAhCkLPmUVye+kJ/VdqPlaWp5ULiqojD8b428qmfYPMNdodMBbIUo
gjVr6qj9pNs4IOnEGOy/+g4byXXZMKp69CewDlFNKEI/b5StLqT8G32mHSFGcxOZS7W9G05AgHCP
htebJ95syuh9K5TMde7oRzmi1pP2HICzIDwm2t0U37p03qGhjAkiTGTjxD2FUAHPm/0iGvuwJ1fe
AmDNN1BAKVIuJkPERgGEe4EIYgqp3aTLNVrC2eDsQsGt/7YODhtSgRHqGAfXrh4Ejx4iOYkZeZ2G
XVF/M4A2EbAbVvdw71lTGDzXvBXiRHTMf16JRzbpCCKGBJPtIhpAO9qqsnhcUcP55S8H/ijXyTFz
2fPtNuZ3Ek8tqfXEaVnCV5SM+DVf25icqwWHDEgqDb2vwTQ30Ch3199KchCtNWdlt5kTI6IGrZfW
8dkGydeYH+ivACtpx1c+ce9BQgKJGqQDsOkH1qK/FnfEOlVID4X/P1rsIOihq0k1322bPfbCXQBw
yBCNM68nJ02egAoB299BUMi0PEbikFXVt8fImih3qxDysDhv5KzowLS4w89nM4n85d6sITOqcnpF
TU0ujLF/I6094KJ3JjZ4EpoitWKyg7XzHzbf8tYO/H2a6qC6g2cYjN6FJyfwlv6AA+XiuH7K1S77
AgQcdbyg+/8Apf1VHasqPMrIVuh+MnipuRKM+YiMvQA0ZFF9AFUbeJBTZIuUOLfT9pLdILYtYEBC
xsM4/sV/PHJf/JtbxK5bSwPEQXObly7avVwErXZr4uJ0qJJ7+ixxV2hiwQhOJppYYhRsT542kCkn
7V8jg5nYvf9nitevhoAYUkO27QTBeZe++AXjEBoR/m6CsgGJ+FSlZ9ElqnoTUvf1bEWwbukxXjlk
/AyMqwaDJwwnGbaaJCChPed1h7tDWf+YrwSY744B4DtfieBChhxQz2wqxWkq9kBp1LJ3a/Y2CGJP
BC9qV0Zmnf+0iz1Og55bBOqoEhp1aBGA4oVLEGSvFSQw2ZhrOCr7a7BWIfhQaOJ4YsgHufB1O6Os
fMc+ZZIXt5psdhUUaeAxCswWTJ9xiID1bSVydJYt2+/h9eAes4DLiNlIAQrbB8kc6xGosndVk3e2
GYw0q1Iu5jlCMrnh2qZZREsYLJWr6txicpgR4dv3lbfrwLpnUjl5Zyi7MuPureLWptxcHAulJSq9
eYpS5kgwS9U8H9SrSZpqmzVvFWXc1UPGS/EBHN9DABX+jw0wOZHW4BXxSUTfsyKFLNbYDDC7y7iX
e74UgwZBvt2r1343DERkeQ5HpWFbvNwjtZHTmpx1OnS+x3fwTA95b1HSZR9K+7acefD6jQR7JXox
Im66dyzZLbJkSQ+2P2xwS/MByzz1BOe3IZVFDN7fClQ0/JsM7zgyJ0cnHNbCejMertPXJLR2eV+m
O1enTphgCSqHBITdL4nlyyfed9NCbB8pMBikDMHgack+iKz/VMhWZ9vjPBSLNr7Dak/h5qt6kBRP
EFV+q0UOurEznF4QHuEl0ciXrkHSGY5IJ2DzT9VsQKZHAqA5sPciSiMPhkVHQfeH8d7vhJfMg7kj
1WSX6CtZLVf8JJrlrshYyF8t/oAyG/baPWPFi7BJGCPW81MHk8QXfyzSJGuYkwFqF6En3GzkRSII
Y71Mh/DykAmwEAlnDvo3d1dREholivQnEKE2rvzBX51iUk+lHhIaMcOe2aOYhrtSaKHwfOpbKhI+
lVzWkBmGh9B9QDe0n65W6QW9qxRmQhSJfPF3WlYjQgMkHNbi/UEKcJa38dQG5mW4RU4n3yHnVheu
UcPiH4MARemVOsVAdoo+uBs1UMOrebYMbbYnEDNGUVO3yUZQYPKDVXxBASsaf5ZUCmzoNi3cfjrj
2RhqzyXAT89ryCN6OBaEL3zp8UC0XYtDmkpOm8sUODcSuB4UfDoVRf0Bbvj5VtVSp+F/7xk+479t
Ucsp/+SQoiP7sbQs3IWsmfVerRc0ZsPvcQlOSEyvigd3zQOmflCdxUPdGhVvQgqjDIwTO33PxUP3
9q97g3g5KuiDhZY4ginEIT7se+nFaZzX+llYFok7E3IPzUtT+CBhbYmBRypcbyVDAKYjuiaOl8wJ
c7oLfunqMZbCjCLKSsFDDiTU6gsKgBMvMK2YOxdqqzwEN4k8fIUu3e46UYVuhPNI2jFUSrEgJRpa
nd9dPVsabn0W+tgHyhbxX60a3S4TUpHjy+8s/x9np9QKg/atDJwBlfH1Zrzca6JgRRg7sudo3v6N
Cu2VOzziSk6AZ1CsGfEYp4ZNcxZobJl5Ky0yKpq6r904qfDjkcW2r1QibdB+a8q1ufivXpp8iqDj
I9TQok7L57jGvalXIuyPFvfQUxZycPKIGYZzwk/cccrGOqkUVtIRO4isJOGbPwEdEDKNoYiNz1S3
yqSKozOShkd4jA5FY1S0TfqcT58zXiAbD3GUaPZW8tp5io9T+DSvBjJnun/3IAYJMXV6+nXGPcFr
dqlNy96OU4oHV02Nlfilpq8tZJKDewsoimen9P5LByP0bcXXOwEFWq99Cjh2pAR321AqrPvqljGV
Lm9uxMzn+pQMi1CKckYXihP0PXiSe5Z/eaYIRmNqETlki4cpDJQP4LnsOsTMhU2HUPPrgMtQMCti
UupqB6Y1b+6w9/rLn3UlszgVQSCYr7pZH01OBqPehXDeH2LNfQdDO5fFHqtxLTmq7qcJNvLSU3pW
t5cTSRT5I99j3hPpt7qqNL9F68UEp1+n9O7cLTtJhdK4FF6ym6duX+OBUK4XsnCBSp/vMlIOEiFh
pPNU64NvVa5lULVtFlbaJaIwekGxl6E72di1jMQylVENP1S6g4oJR5H0b8xODAZ9S9jjkTbN78Xe
BjdRb8cMO0LQ818gNmerXSWD5wjBV0KAkvxiBmeRPjAhuUW4M7WRuc5xmint5u8D66nOmJFcmmL/
u9W6TbjVkIiKPrBkbYKdLxtejzz+US9tM94vFXnRIi9gEKlZQXEQHwDAtCxgCOywhkYYVnKQ4rOm
ivU9uZVa6ZCmzYMjiMgKtlrbX4vbNWzZ5URh29qoVMYqfZAz4v0U0gt4uGVDrbwsJV++9Lk05NMH
7lKtGXfKa5MokrlbnW99dk6wpu2m/aqUdF3ttEUlGFUyJEusZcv/Si4F+59mMyPtbN4GMTPqH061
tLgse5CE6Ja4FZz+07H3B+HjtPNv04KtweF+EAWc1Et1v9wYLudRPkfy5Gf8jt96pTCClEb1oSf4
j12UMHHQ9vI2cezrd5p8/EZPn5M1QG6ZiN4K4AW+V2UTEqErdbXovMAMIF2b1E15CQ3HlgQ9VS17
ElSn0MlUkdBsNxC7ZFq4sFQAqy67NkY323SklbdNW90Ft3kjvoI74YZ7DVrxPQfeGQFqGqJK1UV/
KRNQH8YwJPvi5VSJZFuRZ37vIwqfTqpt0Ep1Ww4vaRxrFxhILTLqPva5GPqDyzFs1Rets7pFeqx4
Mqo8xq6RjRYMx11QdMPilOtpDCTydoWtM02VRmxHwSRZpRxpgXM/rXbYxxvr1wuF6e+jFC/n54ru
KUAm8FSN//6hNkb1zlBhG/2g8+oXweH2vEiaPfdAc6NJl4KcJa1EinZ0S0CsEOk6D9S4WE54ECRT
WncYTOtXH8XSLN8Tlft2w9WZDBNz6on/29C0sEw+R3zyB902GrO+qxQq5hXlmXKBH/KNvOoyGGBZ
um2/oz67NFiRBAQi3GwBiZjJkqbsE7BjYrCzUCL5MZ6BmEdeUXsAS9yvT1wy7dw5DDZT/VXJguS1
CHRh4fO++kw6u2q8teSj/pz/981NbjtsZdcaLIJrhb6icnpyixyZNwrlfA2q/qJF4DEmtC4bwB53
kp7f20JSBZ4rBMyjKzTHm63KRClSvE4kZW/tth/7Ziyc0hxSLuH8/SXDlo6cbFWJ8YmOh/J6YAge
8a8TCuwAxd2h8XBZf9jDv3/95zcl0c11Fb84Z4eg3BT8gimAXqe4XngaK+EoGGTP6ypWquPmnZMe
brMFlrCpnvU8Vas2Ixfulz3of9PDApSM1iG+k/9Mmy0FwZjkXplakYOXC6/zXPKXtTpYAhYathLL
b1HhuTUOsajNutWEhl43XjrjMYDdoOl3w1hvAz6TXsg5rT4xmOivk5ow9sX2HrMwVgU5Tn2JdXso
UXmw8ocmVxHXIHwIZI8iy9llszfa7GfXCpOfa5mI1fgBkjc+7Y/8ZYiI3lQbFLpN/PuDrTyCpoJ4
BOn3VRsP56bpBzpI2McFW1XeQrpUVeHdnb4bckYVhCD6L0x+CDW64ZoGIeZ+D8yPpxFCNmHWARWi
b0OJ9I0L0skhEuldoKOuZmxJeVNw1fo3O23wFw+ykSCvzea8yAx4kZUy671eEusW+8d4tKfBgIC2
JV4Pg22Kiu2qTo9Yt4ck6XEptvpAuGw1x1KNQzW9Kr+aNdN13H8U20O/KLm6NZVgcz7UVrbsBdFw
RujhFp9H7heuUsknjeYd2FOPkouiyWSS1taEpd3cARZofel3QBXercxN4MM2HBoh0d7Hq555+eCu
2tH0rFIKVVVvCjFNaBS5Lk0aILLhhqqCaT/fZ7hXhtft6tADEYWMWtvWJ//IwJNtLW8CnJj+ws/M
4fbCAdPgcThZR/YVAlqFF9WbaUv5gj6T9MEsDJsTKA0UJcPDY904fg0zvQUD5q5UeFejEW9iC6nw
yRZSN2L57rGlkCq3OCOlVrFtwX8ub2SeNNoZyHqDzHD6Em66Q8fT1+SkKoFJlKwYHVp56fY4L2gL
H4OXTMeOe3rnR0WsLdrnkghCPRy2Ha/DTi50PxS/GgKHp+sHKVpdcYRfqpNu+JqSs4yY1bhPvOYS
n4nJjgDqQJMpoS0oD+PSnvZIP6AV0VUsIMr9hNXU/tgEQUI+UdZExwZcsOSTQRGew9YULpRzrm3I
QdKL2g2Zxa00YP69BOQ79FSv7EwmTi9uOpA/v9+aTqLDCCBBWVWeJ2vWpq/HHH3+mZzEIJZ11whl
hZRRiyGs8ExITqYomp5JiFKvfxiptxuSdGEbTVDddNgg7l/c+aNEHXg8fZtvli7JMuNSAkWAcHJv
gbFKo3b/Nea+cXfgAcVtj59zcL5xuhCBFa3oaq2Y+u5mT6HkI8OCwxYDRKMH8OUzTdvvTw66lMqt
1gv1gFqFKqcqFzF5o6Py2Qy9k7kNoh52kIXYA0cM1tavY3WL8jI9DgGvtjYOLtu7//HeDzdn3GIk
B5X7QsaJCCVGnmiY0mPFu7eyYu0/jr1yGiEMlO0vGg4ubTJjzC/QzdIsAbQZIfWXhyqxpbLw9Ptt
e1Zosu1yNnPXyF/dTa5JZqnNeCNBs8rVhAjBMu2G8yWnt5X8FQqznfNmUN/QmPPUDaNJE1Nzxr+L
+KHIfr523DJZfV0jxJYfVteNPbMasxKiuNSsXPKoSZbtEyWT9y2xVImLT2vwoRKvFX1N6OoOL9Kw
gSGta7eoyTbUORD1FwEZXfyzMTt/xiSN9axsKcw0lrhhYESrK3sn8WnuLm7EN1QhhmSIOEt71f/u
TIOuNVUQuq7+CIuzL4GgX+9RfywWvcycF15WmZbdI0VFfiZhc6uXMWLhTVJQZDoM8/aCCAua30WC
F2ycou6k7jFjj+K6CmRVl8Axcz77TV/TCfO/yFu+awh1q2t/+PYJtD2HsLDb3TBH4BTMDfzfJ/nJ
mxPiABWhzeiy0xyWbUD6Oe7dqq8I6rqbW0HqD9B0yBg/oO+bbbIb4XntOEc72AtAnJlpWqlm7Rd4
gjqFFg5hvWrQGOuvBli3HBTiP3QmFgS6cyzrppat2YkYoUvSjSFJOkybAokGcHIiBSNFPJ/VCc+7
ktYNCxh7gs2U83sMReatQjjUJyveJSd8XLRJcBhF8miPTo+SSF3VPYA1fe7XTUX1ZoJ0QEcvosEQ
FIae2MrMPsX1gpHUSZ/cab2aIS5CgmiDgjIM6tuxtxdszEaE2bKfgnWUr0L4IBKOLcGU6Ukh/1/p
VYzn3GCx+Qu2/JGmwGWysIOgpsKxER0sey1Xj8X+HoqX5yYBZgq2C6ZzquKW4Eh7yiHg43NVWc5Q
rxn7j19mTmjArA0g2PakejhQINpQLcHq2Gj7gliN9j3NO9k0Yosz+AQiXc/9Hc8xELwDMIijA6IG
4XoQXRuzNrRoYsilO6SnQ+H7J4Z344uJXoBWrbnMnjSkoSn6oVhKVyB++pCToG9tQ2hnuyXTAdAe
AvcxsfBI0sv29yb58r3+k3PmvT9R6s6mtUS+/A/ppRtmoNc5Qmmqom7pPqDSq5p/YiVkrx7hbM/A
5rW8ZFzbeXRl/AooU77CDShVTM99fXfvzAsEVxCAKR1io8VRv27k7wl69qeWEKwTyypQYAa+qffJ
Vy2wfXWqd3XIP+jkbwTEKS2IPrU/8VLKKswFhWwUA0N/7lGWxdgtheaEBId70nurN3KSUM+5D0Zk
1zJ2ZWU15F0s5vexc69wLSlIqQlWUKo25ZBDjTjVYOHv3AlCpELBuz4MeuM5xz2hINZKKWzFqfQX
dtgPa6btbd1ILbx88KLhLFiLyKKlyBlCqKOrlLbfRqzGY4OLBBNDXqkIco1HU9qfd9H/PAVECo0c
G32mbeFHzCmModD5KR9WRc4MuTf/bmrrctt1b9qzQUhsG6W8Tv/J7VFt/GolGDsGjk/CY4pxnP/k
r/AsjggBcHLr3SMg2QLQpfhjSz2QoVYDIOCjPoOWeAmC/tkPmIVoXlOuzmgaCj8BfMBUOmmomYfF
82rD9Du5sXOwZJ+rwNG+bgc1lbB6CAT5yZO/HBu2RTI8/mI3GNp8P4f6MTJrQ1G21nbx9RG0n1J+
VilhBojXzDe1WYFok8lM/XH/j89IInQmUsL3barXxTDE3hkBDDRpp4pToHT+FysSXTHrnhZUUPFs
ISVvd2QxNeL0aBe03ayjieWd/Y8PJ3+y5lWN3z3mag9moHkoPkWoeJWEr0i5YH7NWQn5lwuASpvX
5dJs9apWAO7wmdexDPifGMdH5DEDUY5TjtrOgMHDs0cg0zP9UmnzbNHFxZ8AWuLDov0TPk29PKo8
lilCJEhVfaDBOAO5ToRWiDYe+DU64KsKiPbL0AbTFZieEjg71QEAx37haLdhZKXCKcIBWvS27m+k
YhGl34EwNSy49FvcTqbKjWovKtTjxdi4a+eOq5jvx9tFZmhcGDQP25k+gDVAtLSt7VCF8fRCn1Zs
wfM7QZltE/Zeg7FyO8pj3N1Q5YxXlZMyJsxteb3vr2OsNIngVfMIQEuxPU4ie67U5wJKUBscl0Em
D9sD2Y6uTh3wBADGfKxv4k/y49n0pVeCSCI+xkT18A5PCTcY1IvgxPbxpiVGMsqiGOBWwOR2gmSW
oPtHv3huJgHvGfprZvTd3Id7lfvY94ZzDl0r+YKkrH43YjAl8vfIu1Z/0T6cVm17THPTe7qorStv
HcBkBB9fjlkm/FHfbhgFIMeMiSmAo6V9Bs95xU6RI+PZRZuIpYwr/U1i231nV/zcHFgI0puzDr/u
s/4iDRTv0S5JiM2OlzwGrSQCeasz29VvRzDWruna5X5wMPDsY78OmdbqhjixiVggfhWzuHs/VOAN
25r24EE5i9/dz8jF3dskRtRUsoRKzj8uf9tS/qYimFDnRe9c5mz8PFAI4xG3NZy+bpej2dhGjIPz
swRHC/7oBuZWTPZP4D7F5HnA3MR2+UOGiSxw8k3Szr1UEgfbdYCAYIY2dVQ1pAuivszenDczubho
MWqOTXTsHw8tGe26kcNNsvbKI77CZjsslKFDke327iXWB0E8J5LXfJwrFme/yWKOtgggidEHC1//
vFfOXgwsCaermMRMCJ20Vt0yn18uhvxVd+5OstwDT6+S/BiF3FqgiRjA1BKZguwoDozWq+fMfLQz
wDajIVLFMLf3TrPUop4jG5g0s3/aBwQJUC19PM0sSGHfFNUVqGGIZoCz3ffuGnjO7lyLqekDRvBI
y0HnaPAwALpFkMYvUgWNnhgdWT/7Ts6ejxx5wUoDKv8FSfcj96rh0jSHsvpPeqsgDuokFoIr05n4
Yv2VyZX/S8TSz0vkosOAinV9McYxJdbhD0Subt8mva9HDh0bBWoxrLvZlf8fqbd8pj0x1DRXg2K7
Z93bzfR+qcJQ5F/cztBnVW66+35C3BJ2OXVWuMoMF7TVPaVmAmVuPqT6+dj6Cw/14Fm242zP0RGj
qXMrMAPQHPHrCmVL/oBUAvADcWBuY7HODEFA2ecJ2M6DLJmXO0Axgmi5kPuck8LVqA4Xa5dMEt1K
deXSdwQ8MJrsC4pm/8nycz61X+FqOVP6JZ6/jcV6NWhwCRbT83cPa3aY5ySnE81YazK7pF9DAiu6
X8xIb92/sls/myqS5ZMmPA87/I0jebyGV31Pa2mv+6IDlygFoU/+n+MzoFQQUYxKZLYqBW158HH2
kR1Gs+0t60NdUsXuUp3x33UOx8k7CrInOhhD0J/Q2SuHctv375E6nVBe8UoeCtgmM+Dmv1kH/y3s
NRz0hVMdCJ4UQ3z4S3aUanLmB+nrkK9vXSTDndWCX9UVlmrNlSEFWo4L+9tanHPPAeU8qUwDAgwl
nD9S5Z3otkSAvtS/nGu9/2NfEW2B3AowXvI04DAq+n6tpVv2B/FpSRHdI+paV1Z5dc7dg7knEkV2
JprqFP7ITngBYPf96WBKqpfpIlt2I1wie5P8sFLMINBYPRjH6RAXb5Ix4cYTkhkRwJQEDoFlMJb7
fz6VaceNnnaCVzBbgW/olmdtEe2dPCdwcS6mog2a0ytzqsXbsp3Ojn56ZNdLdeMrIkmeneodVLkK
G4AO3ou6yodYIJPVcWr7t/AtQE85Y+eSyubas35rjmFiTN423vXd5QNzh9Cav90/6JYGDGBGZFSq
WMFFojC94yVt3g3kx85yFyg4q7owl43kNzUqMf2C388FRngrQcO4Qpzi1JD2dncIXHIHqRJIm600
tYv5NJjhICVHvWOwVOXkYMngDtF6Xxvbu6WiH0a6RfhgDDa5eLCCochORUYkWwm9+klXsgKzdj4y
A6l+Sqz7fHZhReutqqCq2VdoWdvqVctoF9w5djp1W3gfYEuyQ9cUZvKNemNiSYYGXIkSvocHg5qm
7rSKoT4d3Z2cmLucM4zI0/p+hrELSO/0Nzqe5bqqAkPVcuTyByr+/cfFtq9tuh3QUO8nVsWoftmw
NbSr75Yx3ThH7SVDEZS+0DJOnhhpPJW9U1kTU2EQXtYRtTOeR5PqN3l1AoRm0Nj6XRZbTIZL/GQP
Cp9vs7cypFyg45MNgsCaASTs8vWBhihfc46WeWxcyFiJn7t2H8Kv9SvOU1A7QxIPDoRB1eOc96kn
v3f2AMFaEGYE9svC8+fx7SEBA2FUcP5VFWwMQuoVtv7Rgfslc1dJuhj0oypjC9g1qo1JUSLJbmfn
NRbikYAygoGzO1AeL3JFsMgGg46yL0bAltcQovOJBtcEA1o6apXsj0ccpoUbn9PR9+B4eWKY976v
z7Kyn5sru0q1GvVTXnCnATA5PqdIkYjrfWanM1bhyWmoySwhUuTCq9rReW2sMcYmPdG57FWwdHIN
2+ostwmsSfbuYSpFd6SG9dYrRsR1UQL9ajaCbh25JY5nKA3V3bAXxhja4WJe9AG27ftEHtF6u+Y2
wskxwam/F/v9YMW/40NpzwtGRN/yUkqngwX6rGiWMggvp9OsFZJJ1hsWDUrbu4Is+6LJsWo/1w+Y
jaqnXXQ6EwzjPfZ22N9LkKFrHvUaibc9yDtTyHAsmOBf7yYPDRlUz+Bhrr9P7u0EzX4fNBnsn2ew
QWKIrhLsYFJcBUauvBoHB4liW+KfAWnr1zFXmnR5bw2AKdvsHIGcqPThYysOzPq7hMKSRMCgDFcp
R8Mi+5gDZlIwm98DnojJ5DUg5Wyk9yE2CtvCPj4Jrl0f5NVbMXjYENyFsXPqVdGMAkIImFmqsjzA
ksQCqXbZD37Kc3VdQX0vcH3Rr0nw7bpp0nDEO4XhsCGZZZw9p1cCCUhcDaYDl8KClKjg15vQgebh
Zke2NkqFPEGaP/F2rBMKYsGQ3I9VRvYwsW3DddP+Ww2f82fymgG4fIRXVr8E2C3SBjpJe01sT5GW
Ag12bsaIF1qX0XaTsLTnEJEtjvfI0yzo/Ac08UPfwrq+nf+cSDtSoHqS7AQfSQokfP2X2HdiB/+J
BBIxv7TPYfAY1fDXj1sxBPgZn1NkgVLfWywchorw7M7YI5ivRVCAE2xkd6xmB5K1bq9zubfldgiY
RiHgSq6Wo5th/BOiKuWaCNPs9gZxWnOKkwz2pXBo2oZ8aFsRWwp3Y5tvIh0YbE2TVTWfmviE/N6B
MaLsx8iwO0Kddu+A6fxqclAA+AR8oie63s0xvYjqytY/0YDu2FitHjAaI+A8DX5wfSxGEx9fwAvO
lNl2W6XsHEx2w3zUbP2XzI63QNcM3XimE6mFq9cqmFR9QfG48XZol1TiTRz9VoEwAFZEJbxmtDV/
HESvt6WRfgDfEG5oUs/fPvxF/nLZyh79hC2BdnIq57iebKCL/T/UiTGc8GkeebG5h+QQpJZ9FNDH
wmi1snj+x3eFKq2Ejz27zdX+mYnW1q9NSrmr1PzSVCrXPvQbBRDCgq7qdB7BHp1DBrNhR8eRbd0Y
iSS4rLXruacsWJJMB2L+2dKP09/Tc+O7foioaKp8vu5DGCuBONUYa42OHeFjqr5s2wSyT6nlIWfI
lJr9x51cObYNLjAdDYHUM0f4+XRLiQsJfi8zG5RLNHAU2x4Kdc99n/zvobYD4518LvJNTh7Z6ulR
IW1ViWtdCw/DANdazKp4aPj/WM+GlMicq0jFVoK4FZJxo17de/8oTF4kpC7zd5Q6PrhPEal0AzuN
BuH19dNu30JZfdu9ywMw2x07Qpi75Kx2RAWsuIGdeyaGh5QvOU++nViwmPvuDMZaK4T5OR+pTpPc
dZyGAX+Z1tGUa2HL7HgenOeRRK09pMkyRPmw9IUfm28lVRH3zPwv3Y3QrKlIlA5xPTQ4sCtSBQYw
CGyEGwZXGD4yYV6PhfVUdxpbGBgAS1tdGcjEoRmAmC2QVhcVmG/S1r/kbTqtAY+Ux733OtimhIDH
qjduF//xzkNhF9c0By2+ZvAqxsBv35PN/odgD6TuVK8cQgYkYJFjXV1xwabaxwfcP78zMFcOGeZD
NfuFgcYTJ/I8bUqqo3cTYzxsrJJTOM7qDIC8ujxQJeqx+ibd7BLqt3jebiFYfkPlWN868xAj+jTt
ebvFKVJ2nlfXhw5Uku/NcaBIei0fhnz9sir5Esjj4UYGY3J97Fo15w0ByVkPpmmPahZR7vOYC2KM
iYcagTyYiJu/l/pYdDQr2KxBFBrM0ewDNZVzcS7qlCkOX7zrXHJgEyOoUGBedpTY3iKSVLUvxR+m
c+GyjcH7viLjkDfN550VQWNy2dc2sLc/+dBJf//nwPNibLBM6Y6FPYYxrJPWszwC5/tGRWOswGDa
0XHHZY230qWivxphYyug+bAHLKXuG2+GOq7rSusn8J432VCIH+90fg7raanshH0HBG+sOjAFOQqi
8jJPNHCF/TH+ZKGr69Q2k9IiIb94XsscDi7ufnn1YEee6Nt5Niwgrh0KU5WQAEm81HOWgI6q9sbT
e5lJJQq5Z9gCS4EzKefgoQVkcvD0cx5KOXJeQ6osYHR191rojhWb0gu/+CbOw/hXMajiPNtj2kxy
pELvSicEYxd5TlsXTyP4hGq7N1/bwASMMTTOpMo3AvJX4AHnDhFFyBOT06TSodumYneitDq1MmQb
Ep00Q4pcnM84N00f/qpVxCOn2gWac5Rak/IaiQ4wELzeHZQTYunnaT4v7O1LvAtRpjigbXH892Zs
OHq3XWdKqOFqMx2SCAYCFPYdpbRYqOJgGk9DNJgQUbEDJKQxl9CtWnzsatkapUyBWLzewft4B9xe
xSYKbMuUNKOnciOSo5iHCSO9o3chZHmt+UC04NZvWlKfGhlTKT/R+R1OdTn3QeZ6PkQa7VtqdW1b
GKy3MfmmrMQI7tbPKFs7NxhDIhJYg7g52TueSTrOyJO15rJEubn76H1gjFm73Ix05veARyPX0xl5
y4W0+VS6UOQNdZbNqUARGezscSh/gaILxv9h779P4oyBfBZI+F8Kiaa5jnYz3gUItQdxi6XMIFCO
4+G3+pM6DQaQoBk8EnOpRwx2IxFtTsts7rDutReaYX0UAS0nbLbeIcMw+wIAsJ5PskJT0Pbiln6L
1qimySFoj3d+AwdQ38auWrtqhg3C/w4CGPZ0bIoMwIHQ+m52vH+ikz18Mh+CzRuBTzTW4AjctQCI
fi3DKFJJmTd59kk0WFpD5OaSEZuj1vJaGPa8yMa2x2HVtgjHsIYO8CK+MU7XfJS8JDqCHd4GBPr1
QeguQAkFckgFUn6oVEjnbPYOs3LFUQhwKCpWieRqqw+youVzRAqm1wWTj2Ht2r2BXqQYhD12LtUa
n3maXbhW4964u4eRHsPvu8rHbtv4ZgXpQqoSnYpNCqnCD8Smih/cvHGzl01AR+0xs3VYrjUz8csd
sDDI06aVaAYLGvJPu0E469620RJvn+zuq32Qt+FBkMsvXylTIm9lnJkgqSkOHPecPNwvIoeiO0HQ
jyY/m4c7hbI/Bjqe86xlA0QqERvgb3dEyU3ofO89zA4DCllU/bSKEfIkZT7vtwAk5VJBRldLT2Ql
5x/mpzFCQDOTjO0Au7SFfbz7iaLEF677yZVr3WksZ3xTUHGDGhch+LhT7ynjRTCN2+eoNMYmaiUE
f3rYxRtfEsE2BhtPRu4aU7AZTRDtrVI9zCRgQRR4BA/VldQCwWTFZzeJcBZymSq0toUmwtvkBQA/
f3YZVb/JEERCMNQYN3FQIGKLFW5kV+zQgaBKzLBQMgObXaANjI4HWw/NMcvXMpjNrdQQwQ6SH4Ya
3lSSzGk1WxwYNcJHmGbAUdlwuhJCFOPwjT4QzniV6Ay3q817YpI6baIZSubePGpfxE6W6GpdTaIq
XzHd86mqFwChUNIP1a+DwR4bB5sleEfQp8lf+1kxrSMbrHQSZSnhkzhMTiHm3OTyLlb+sWPY97J8
QqarujI1Gndlb335RE43uLLFbXUj6JHx0hXwrtgifx3V6qaXdTqhufUFIDtVDQ8NApXIDF5WZj6y
g3rGNqtR1HKnpqYHY0s3lhjzz/HGmkSv/PY2OPzOx06exGuRiLZp5K4Yaobf4XGjIl3qeUcfyH9Z
5eDoUxsXy8jTf3fUQIMyX00p1F2+epwULAWmLVQI8SidLSOIBjc5MRa06q6oaqRvMelG0GhG5JAz
4865vzMjzW/3QoCnJv6LGnPL016xm5iBoAnXnTWqZfTKTny8JwN+T0ZUxqddvOoqSrzcFfr9j34x
ADr1/v03FPJ8FjqFv98X5CWFqB260x8/lmevi/oqum0vMGSxJ0GnHISmzFp+nRDddOv/v6Dp8h2v
OOD8e0h7gKHAWw16b/EsAVY7RoU13P185Darvs4+qOvVVXoV/dtbUyQaepdIKKRXip7wh5zEvCOo
h+MpcwjKnzoSaXgTItRnE/Pz4w90X8kb+EnFamALDM9HE0SXZOzu87RdiX/1leZxeHmdRk5/uL3i
Zhf+OMRUEOho+iKHTZxrejrY6KJ7aNzzooSKADMstmWxwA/F0m8/fr8bvAjMRAAXZf3cW1CJrsin
/cuOgOtHzv4PwelQl6XyAUszn7AgXcsUoFyAM734kBo0KFRI/VngxWYb0p7bT22cbGmFS/OoLDIP
TjTgEtQoAMlFl74xf6JefFsEnodoshatUpHygmvVURFy9S7o2eNhwHE+M4GxsfE+yNIBQphzbCa6
v2YzzpSZNwO/ctpupfiFxDWSUEgh8Il3TVnxMawWIgn8QfuRYwFHy/zU76xf6Umw62CMGBrVJRWd
xBfppeDyhXiBYj1dO5MPcqJnVkiXTtWCmuvGecgT/kwiHhwgyxBrx4LTWDVC4JgEv+Wucek6pH1h
MZyKU/54o1b1cPfV2TlfQwSxmsNpqaCEIClt3IeBgic87S4nqLVVvSCvbVTx2m/Mj9+crp5Epscj
KJBGBp820Mo2YSIHB1XRfDMEyGE6xKEWvsPV7QrS+AVtXzOZZKsLH6h9b/lbRDOEpAS0EsxqXqLl
iz1clfRlzUZ0xi0p0Ofgrtr5Luqq6F05TClaImWizloRbfzGmpAy+BeN7lZWECQbDbNZMSePRqGS
fGmmKoA2CxuFpPlrKFev4aow0krBK7E2aClfcLFyy59Rz1fhoaREv9Ru5gHBMwr3zRVFAY7to7R0
RQJabLGiZzJno7AwWnRhaAf41gBMLSsGS39Xcs8HCNyhEFQ3kId2jTFy2KOmu/4w1KlL6shPCunC
5PE9nLlg8BUkbNPAi8nffATAdb1b3asmZBXEBuB3HNB4fPVg4vEQomkE3YlmleCCIPLiAhB6bGQp
TYYISjb5jc62W3V8c7t+tGabrpJlo6mVtgvsbxReqxf3cWRq2g73OKmB50QbBQSC9QTthZIzGkbh
HAen/87Ece/ILvFmO8WNk+/OmpfBiJARJKTxSvgUr7rNt+VRgDTS+2PB/SvSnNKqRaosbm53UG5n
lsmUP0+8CQcgjEcunBK2Qvz6cEn7AHeFxPqDPO3U1mYDlBBO4EmEyzLmj+/pIrYJJoZkE7H7YHag
MbZfgZ2lRpGNEEv/A79vjyyGsfxepTsHnNyQUlNH29TAXfuiLbkCnvRaIEmvZm7VNlIUNeas4u6o
4VYdULlqit90JdHEWJ2YRgZAIo3i1F9rr+4xAl+H+iEskR/PhKTPXM/fNhKrifeQelfbeSowXVaZ
jWK9StHb2jAgWaCIG9invDe5l7yEUiIPBYFPD7o5jn3NbjxZsso+JVv02XQin6RImXl3YjQJ5s3W
q9YYMB7pZU3Oew3Bl24veZprIFS+5eILV302et9lxBCP6S6B3OelqmfvRyxcX+s496X/jJSeZKHO
bfHU6vs7zey0p0mSERfjonJkI29d98b/nWu5CE9eN0Pamee940loQOKFWukb+REhEC0RDrAhVFTC
MWeD2J1caEUPCYyIhvFdG7SqOgRkdJRPyo9fYghnMfokVFooeba5aweDO5M1Vyxh07qjH6o1UVfY
MxzfT+jcO0uZlIuha2AhPZErBrhGra5mwAUHF9am7Z4Eu2fd6TWjNLmQqdba21wb4rOiIkY83qBM
22WSAXS5+o+vHRUVGKFFAjTcjbnPooiGF6CBZKFrF/T1kaOe7nMnAeyijOmScriosTemQb8lrUcD
RAPJ4E4Vz0oUQq+zk/XrdFfDwZfG8bQNpogmE1JcV9YF/m5FiAr+hZLXVlSr1IMNbWwZve91lzhl
GC2hnbgG5KTap5y6fWhXMbV5XEjRuaD3LAhF7SJIuIrPC2cokAbYQxhkUct8HZvGAXGMi9OTrGmt
TDVCnVPARmNYqgqN4ALhy5uKnHIwvHbXXW/zwWzZfY8SK1XLl69T4Ykcl2NAwRlTzUOKGojMW+ho
jZy5SbKEuQIbmUU5bzRH8D2GHIvyt1lYaNXqXrSZeYawjWXkyUfQ3KIrLlC+cF2jRrH1f27PH+gm
wVgj1KX/XBfmXQ9SNQg/+5urKVPx7NW6nbgga/TiQm28Lk8hTmubLLdDvZS11tPb3F9ydpRcJm+F
eJT89BPzIOnAtXziM5qAdR/w/aM35rESnMHq2+cHoWP/zGEyVPyLLDrK55Gz5tym3eTxa0PRSrOK
dBBPgVfaz9F2Y6ng0kyhUHSqS3fXc7wLEYDiEPBIv947hq+c9u3sZArwb8LYF6dAU6uUKUj4RIXp
/usjJuE11/zc2MNncVIlMziY9pEuHc8JGPxLlzqAew7PsBuX17Oq4NPQgjQZmEs0Y9SBMKljdOJ1
DGeU6CEBG+3YF42TtAd1tZio3DuJgBCbvnJlg+7qOQLzuatgJVtCF91xLI23W6OkZntcer+Hyc8l
b79x6nMxvYQ9m9aP/y2rJIZ8aMJlAU4sv4hMdrlPfNycO/S0zCTWyVbgCWnDE7ASb0TRz0thd7yP
GkxcRdSfvH8ZtzJ/laDfYQ9rQhatvEG1FOqW9fa/h8rr95h/1x689jqoPHcPrH5Y+EsJthny9kT9
6F+MO5hOmTEuQhMHInAFbOmNrTvfwT8LqAWwA5s3G1NbL9Y3j3rB5qsPXs7KsIH2t+Ym98ZCJylz
YAWr4+kMarh9I7hzGhgophTMUUfcpwS2fCpu0YTiEP6FfxS9hDNKRdXOhcKpli6flh8i5AEx7kq+
FVhZKdVcpnopHGtCqOhju3lzMJtwqZDHBKhu/lX/sOsW2DoM2L/lAcCtqmi/iOj+mteq2cI0M7mQ
btybSjFq/pder7g8o8z3t0im+/X4t9lvHfUq4+cqbkmlFRdCtvjFjFHXPgEmZJJJHtHpCEJpL8LW
WGRuOqFN8pgQzau31VVGl0MZWumvIz8VaBBP1EVcW6MiEKDW7y0YFkUcPdPwN4CLJNNxWP0mEGeE
T6pERdk+ypj2KPwO+g+mpgkPttBxD93wNt3yDm2Efep+8xhfWFbH+SJKyjpBxC0EVBZd8KZZal1a
ucKBbFHCVlAITfmiZrj9oKVal+H4NqBr+8LYYB1WBzNDuzfiWeTeRlk1Uc+5pU4WY1eQrlqyMOHs
+oqVl25lVTfp1DQYsbU91D2pMLTHWqG79XFmz6YOsXRXgxy48oJvjeF7EGj0gpNKByNh4XZDXZy6
Q+SgoKtFi7nsbZJB51sAy67AJfFz0u7dNMM4J/HTx8AEtFqQdDE4I1o+sfNGmkRzO+qwDvfSEcvM
Fij16at/tMPOcn8aomHWJcbLA1PuOrTFEiYZ6kpeQqgrVAvDxdMbBbq1uidDNyuMBMn4wYa/Vya1
lCISCMfMhPrXEKCxDQuXbW2kb/MtBKO/vk9NPAd5nz2JtBRM1WVE0yODSwkgk1fIuGHN/gMuaAU6
kuh0vcrKmhk+xzBWtRklTwbhNKYFHA/RGMSAEZxIdBunODfAABUbRnYxOVaf2RmvwzF6S307+7S1
nVMAG4150Kg2tCUi/lCO5a8vi5ZR3TuXyZHyckDZbFpDmu7kFkJfXhM9rgPpJsaSQZbaupWaoSZS
D6nF93YqgPkU/gQeDYi0EKzjgjU0J/XFTKeY+mdOZYYBLGDP+0WPCwfm2NXkpcDgcIjj+WjbGC4R
6EafsV/nqemHEq0T8qWRqBOV8Mt4IqwDfDDRAZsqSFhz9C1PzCopYLl0ljvmn0cyAafTWHMZYAOV
NPDk8xpDFp+FKenWqFsxe9ri6EBPjZskgS3TEhXDuDBmtf0kORLd8OHTndJ1I3yyThVjN7YV1avI
ipYOXA84KoDX3DPtJuksj8klz4drbvxWjpaS1zIPOEmX9Pq9gUt2cI6MvDVE2EgUHw4ZEvp/Q0+D
lFCd6FpRnIUgJKcVAXTB/wS2kP1t1godRc630oiDjJnNzzUZpqyDYkRKiKfI8lppmzidqpN7B6fF
nDdFkPZudZOop7A1AIG1Me+OlN4ONvW/Ci/piltBqVCCVPpMD0FQ9QSSFBhE/jGJDKBfpAKTsiGi
fEHYJHHuTIrQw4PoME2j26TdlBurT2qPLF8t5dVnXGO201Pz6ape4mBLamJwlULl5RRK9eYLK6Zz
3eBWd5ONDMXMEHShafQR+TomNzGNFwnyJFN7A2MpgELIvrytvSq0dmZgS3UzxSZOOpT0aCqqY0zN
pAl7R6Su0lhF2tfShHiqQDiM3sEX6VZvMa0+pyW+kjujIynC5lQMG1LVp8I8RFg3uPOqT+Ku8ieR
VtUH/1bUCQKagaEZ9UR8yRiVVxQQq85vMrt+STODPDzvec0bGLEdN0urE3H5cRS/Xpgw+8+wHSHf
OwBUOe1B8r5OfttTbsVe/XLI3Rfx1/dw1SPLOaoQfNn9wJ+wXlK9OlJUS6VKhX+neF9DyFOS4hIw
Z6/BxfSeiCsNWvu3GxQVkxsT2QVdypYyX8Z/0hiU/SRNmL/j9xZkUBCK2ua1l30kV1usY7Ucvjcs
ruvOhh/tTS9h2rfZoPkLPD9lWaCWifVFF+/5LQcMAbZyvTk9AYeIqCLckFje/2cczUPOgTvvKScu
JjgWMsZEQa8wI4UuECoS2JVMO9YETBvvWKgWTvh2KFnPF8mnTpyijqR7c4xw3EGKm5t71dXAOF1L
6KWprMF5ewP5j2cDAD8osCfC+kOdQm5EhWpaQy/ZRmgruP7Ls5rC/nQBFyxUCgn6NBKOfUurJ79C
EGhqRdZREoXLWx46iQ0MIvTT358ihQCCIO+hjGLplSW9CtkiAlmAUXjek1jmpa/ex5y1ksExDrNr
p6lRUJW8FeNko/uCX/3sFGyNFfp8ePhQoAJu+aN+HerW9J0TVq5YQ+3Nq0Bxg5C60jmr7TLQfsZF
Q+Cbyyk+XbBJj48Qu1fG+npda5NtzwfTbj82qtD0hCghAuasrVy/Tia9YhY7hyO6OMQHen+xsrcg
L26aZXV8CdWzsMP8+fln1wM00nIsetRC13hQyVGZa1U3+0n5fFAkVqMSt1mNc1171ijANlbXzIdi
hKSeh/62vrTPowceNBt7D+ag6eM0hl2gw9kDFsQsYO9gNdp93fB/CojSSh4QBPZ208Hdf4GwpDzo
PZ7EWx7dit4Q14IKQsIHx6mLpxrsRNhL7/RVfpqySLvtelVZoTjZ7J8NpgCg8/98xDCt37CRbXQ4
WLhpHcM/bwJRwz/RudZG+vvuZaw7BtmiLbGNYNVz7vydiJecsMFXmexcc7GHQF9k0DOmjdN7T2wN
axT/vGn64+IcA9ghqRv/Ep3XT7kpYzJnOaZFzIVrmgRsNpPOiD0B4DwV9ciu+sVypyHhTuo48tGp
bCEMKzZR+1Qj3q6DNzf0lDVrLp25HEQ4mR1rKriInP/KGHrijhYEYM3VvxMlDiVYJ+qzgr0AESBb
7EeYv1h53Q4nDv4OGeL+BlxzPGr0I7RsCXJDslfMsXvANBTk6LZysFS9ou15OuN1EJh/SR4dxlrb
OcvkNIawaZZxgLnTCiKhKYAs1u9B64WDtvIoyplIwx7gPr56FxgxDie5jERusAMZ7rcEmm+Rvbnd
vwvWj4LcxubxMSTHaUsqL+qL9pNzafizqbH2lujhqMB4vwIV5ZhJblooCovQ0FBtWYNHVowc2ytC
A1yAhtKq0uGVUoynU+EvYvoFocWDu2GXUPwkBLCk/+FaqFXBmolV0Yb/5vXbWMb2/3AjN5QeFZ5X
nWWEuWi5S74ZMCp8nmst4VnKnlqCRwvc3mrulNHD0dXaC1KX2ljscrWuCTyxJM+FY3UBaIGokCwU
D24JSEZ0DUdFHDjd3oSDBjmOHTBNlPJu8R8cBDIk0XteIoBAISVbue/dcrnazIezemg6VDFUtNYs
rVd16aE0e+QDSeySFbjSkuX4P7xv5SVMVnqg3dEsZBGBkjDLyhRFwvhLjrs6TqehXLQAPQHLWmk9
TFGbNpyFLuF13Po1lKTm8NVNjPjs0+aiNUVjrrBeQyHjgOTrNxXmjlwMOHwN4j/aI88zJ7hY060O
6rQNWf0Yo2gld/w4XCrPSKwSwi5xGIstGSBecNzzmCUC7yxnYqsd9RmXJqEfaxqJtxuEaqe50Ph0
v01QjyFb5hWuqrc2jbDfF8EN7C79unfmYjDGg9nzlNOCADDBOC4MiQBbn9WJf02Byhk68DUuf1Jn
W18rE3y8bSVM/9fHKlyyK+x7x8P/LyLcCsTiEV/4Cy0w04GBt2dBfY8CpXscCcFe9XYzm/YRz0JX
hQNMEx28TW+Burlr8GYdndttui6J7qxvZnBvyaRdO6dA3G0frMlwW0jViY/wf/OtUS4AzDL1sB6J
+BlzjnYjwEOGvhF5VzvtyC3LYH38IlXh0LfcTZa6y9B6162IkosZam6noDncEo0g92VmUGdLosjV
cKDovzbC6yKht5QOS3plV7bKxV0bMu3OlLe71Uawh4SBSpX5zpENk6U2qwCH+8nfKh38L9WOWgXa
Nb0JgjAon/9RxkOGdS1HO6CkC9kk3WViWQiLcNDrYbrtzeGwK3MsrDqxjP0d3ha9v4ZalzNWYSl9
sravwNQyt03+t5w6TskG3jVX6VvL0nQOY5wE3zaEtae/JeUVT4/Bd9E4ztXaXbZ6x79tNfaKZItu
cuidPrKys2fzo6Z8bsH2EF383CuwbtnlLVpUhL0im1d5fqtmDRBc6p/3VeamG4+4m9DGrSpFgGLP
aryfHz5ZMeJlq1KY3xKB9SyMAL8tnM2IY4aXrkIoePSf31L2cUf3kULqZjMomcWIc67AfFaRA4WW
hJtac0U9b/qslIGkq7UCb2T3gX/LNe6Pm2Wzl+wsfQiA/HSRPFlbh6uDXKZ6Zjaj+ynEnh3Y8WOh
eCd9eoLw1uZ9wU9LhtEsDdRV1wf9psUim2z4V232BTJgdnmomQmv1OCCjNgSjYCAs23kWmlf/aLa
4KyASH7L2iNpSgQHsLlohBtrm7C99VElbfSHEf1uODSXNJVlpa0GOv/rtdGdtfnmDuspFKaSw5Qd
wwwoKK2KPhRcO8X1UbQKytXvjhWLSbrYaTt/v6YJ+lO9cDctpZKkuopf+c0WzzLoMPA726P9Zr2u
nggIp+rXomuAVMc2EUyRnJUCBcD5wKtj2naVfCI6bqdFtyW7BITM7VbJU3zjg0+VfZVDQNeSEpEW
PY3p5HdEOFWQiI6dN9fvY3vPNZOE02L5gooBhLJ8YjRE35i8qBB5t458gSAhn235nZOUQakd+hWK
csd1vF4PjNH5WmMj8iLAjC4civlJb5GaLQvov1hxCpbH1/5dXtORHzleonyrO8C0JBvOHhQP9HHx
mhMD3rLb9yNxrz+8GpKku82z1aQuP7/wduhQ9pgLi/MsgwO7ocXNKparpuBk1fcJLj4YYOE7FFiP
NJiS7JwPbwYceV3+B3/D81oh1mm/bEPmMr8sjt90GAkVLlap+8frn0P2cogH6pISCf11WaA/fUey
WkoYQJ1z/5/yOaAsnQrhwxYDIuq/I9WJUs8/SSAzVyKKSQn+34ufqm6AfYp16Y2D/+6GY0xmKKcM
tdLmzZs/O9NRWysEvlRyLnoWt/VQWiSbXMU2B23KGACz0Qbo5lBaxIxGf7Dnzqby60ZGF9A1XQjC
ECbj0YfpQLB6nNJ11BnxcQLv56pywhkG5FD8wEGCVmvHAOSWNIY1npnbtzaEJO3DC6ayqUTO8Odu
bR4OZ0szmdPNZiu30TiGiqC30T8Em8tpJkil/t0JzqvJ6jEnqQRDulQmorC1GHSCT30DlSkVPtrJ
Wh6yE6bP1+IzmiWLMAg5ZGykuK6cpQ/HfABzb6BgjeIrAbQjHoDGxKyAklx286FQLK7xmVWQFwJG
Fy5dbE14/vQp3QtpjZ3tmpu9mJowcL0SAUt0Rqoo2S+8fSBsnf/9HbKrsMyLo8hCvCqT4DX4CAd1
XBG8zjlDrb9ils5O4DfvC59Q83lRkD38wKYQBCP+XbOleZbg75MP9pERbtHy77eJeoiPnIu7+lqi
HfTdSVioD//F1HlKSb5cODcoqraxD7CHr2KvBg9sE9vELfkXQh0NjIAfpfLIrHqmCDtEkapsb56m
fhwPJHRXVXAY0yEuzH7XIvbDAe65YpM9u1IFRI8l/SH58XI8NfHxK0R+rGmQIXhGygzXRdkYUa8A
qw7TrWl20w+0Jm9BnOPGc/AJHFGpdWcSXKSir4TkY4bjuAoQfgg5aowqay2J4UqQJ+gMIR7sr0Sl
gfUzWRJ/g+L6jhh8VxmbW8oTOA6eP2+VilLllpsmD+S9sR8ggWEfQe34+HcongEU/w+UiNJGaD/N
00tRhnefmbyJ7dxo+YHGBjAI3VubSbUmJm+oeJ5lXhaOq65DoMn6Izdd5EewQE7IYbN9HJaLMpxQ
/39HMwYwM7DAyQqOv+n6xc3+RX9yhRBn+RnVBZMaVcPOoSFhEW/PH2dOrQ6Ma75BgNjG4FJ0iM8q
BL7c/DZhf0rgR8aYaGmJKX9UXk316A4wqo/rHaAAjBVpc/gJ9lHaq6SyqWMxiOY+E1S8b27xx/39
hK4QODIVZq9/QInQvPn3na0YzlbcjsMyVvwg/Fv9HWaMAKl/6aSRfwVHKFfY1AK8H+PHREM5Hf8v
lVqhw7tAJr+NxoGbJE7ogUpyxvTY+bd1bdwt8xQnBvBiM1DytdKYEU/akUXvFb4WwwL49Z/rc0ck
iZmGMsyK8hqm/vpJAMPY75gGpMmeK7UpOz22fpa066uvbNgKq2SOZxSUEl8RAZzFlAotSlKrY7j/
EWm9RT29gUyhalzTwNn327VbrXJbqBVLaNduJF0KxYrw6djZYrZBYb2P+yvZ+Rno2t/XFu7F6pVl
rSRa10u1UwsQS+iVtA9+DqeY/4N1QdSKjPFfH/+/md6vUNMqgUqkj9uYYT4QGPvbkaVQ+Wodc1zm
HsoL4nxeDdK9deWFF6LkDWlW5DjEr3Iwpm4reLqrvba1w9AhAiGOiTwO94GqRHUP6J1JH+b1op3L
XHQ/pkvrGSJmsCHIqum9a1fteNWMLOFPMl7PIpmrP8vFu58yejrwAhphUfDzwCBRO3kvZrcg3OqF
cIM61iS+aOvY7buhglvbKquGxPq4o8FKLiaZ+8WcbRx3T1dKmxjZ2Zr+py0pbJaRpZ4W3esfZrdI
An+VGSUU5gd3rP079nnyLPT4wwphBvoRKjoiv7eYxtDUxEgH7cIq7t8TAZTrXVMnHCmqs4eiV1hO
WL18c51PILmttOa37Y/1M76TGTYknPClomohyBxWZCHXjQULv//QGyb2PdyTA1prXjUISiybwmOm
OZr3Ux8slF9LxxCZdeSqWIISZ/QmczfQweIbdZRBuQov9+t6B/f0s45tnGS++91leOz2/LQ+NrbT
BTEwWf/Pgf2aFuTrsdWzuWhmM2mVufRjArDeNT0YijsTlFM6+n0G4PZjc75qCpdNmvNzmHbwy6ZI
mVPsFYyOqs6DdR60K0a1HmAItN3XOALTcJuS9TKmcnywpJZOn8lSTZ2REjOfv/NXc3e3emCc3yON
eqly65CkFXtKCpcxypMid3PlkexJh0WlqfllfPxO79deNJxk0kDkwHEwdHDDNkaaTlFiHE3+egJC
JXiDWI9WlvEFdy9DtNgeUc4baBhwcYmvV/SoqE7xxAeXPHzO8yco2krR/ySKCOcBdpEet4NkIwEe
a0oU1JWLHNNmdPTR81EnHGAMmcs1i4NWENA1mCOcrkpTKkQA7vDRZnLA5XIV/MRF9xwW+dsDgsqj
+WT3+RXhNWEgPMIPaN8uRwwajAHXeCUgyb6FzjE72H40jxRihTDsS9kRrYKeDNO4h7reG2JHD7aL
83nDzRG1aP3UFmQX5yVYdfgNx2sq908gZWWLSRWyokg4STwqCOVaTgLDWBaDZimPRMhzuZ7zqFGL
URovWhO7m4CyHmgyqUwREEUx3Q4XFW3nawo37DlfBOTcOE/LeWYszhVGHLj4aOWlZo/iXwR2G2+7
eTs4vQ+XM3/w9gX+UxOIMHps7wInnKs5LbRsoyPvYHrfMRAVWsfgFQj0kZWvQ0Kn0sScyK1R8Jcl
4VeFOg+ai8lmM6cyQ6xZB40NWixQLf26SNreQvd6/Bg5YNtKLV6W2TZyXcUxtYzNs1zBBVsbkFs/
uwBmE003KELDgEz1lRJuSLkVPQWcWjR/tmkUGfLeYiA9HGOlJ1vNZ3TxxZ6u3EeDISPCmLBHg7lf
sQAz1849S9RxicZKTe6qCVHgKZmw2JsN+GS8P0onBf1GnvumXx9mhxa9GtGhrbqDHF4jR1BWhRBB
rETTo+jUyfB94JYocwm0JXrSVsTVrEEVNg7yntszftZNxck+4iTbzrhjPk8gyfWVQGgYmE9Yl/V/
VrsF8B9Ri+xqnmx/ibhF37HhlHEJBxK1C2Jn4yX2oTvPt+ubaw7WywXv4ApCyelef4DwEakoO2YX
vSfpaZHYmOPiyZyC9OdbOB/TR0IkQJvGXihvgs+z+1AXNX0QMuy8VgDF8Cj6B2ouqmZMxDtIGdpD
WBlZ6EyIxD/L+HFyvgtcm/8SlkHfAjiMYNhV2j5KSTvqpN/DtNXq5upWTJlTSQVnp93wl6tl36p8
YX4tTq5MrHSVr7T+YsqaIIVz915D3llsW0xvtdcddb3kokEp4uEbGz13DbHahBiDNNMCpO6ICPz2
dtb7IZucIyn4HDyMcMwxY8mZUA43qlVl9tWSejdC0psmvjbhe9zrOb7UmlIwLG+i0eO17t9eAvbg
+yI1CyXRt601xB1pFtAA1GDZrPCPlNMu3YHQ1AcHxtEhdIzn7RCufp60R9z1VObHOGXSP/UxaC8p
Heekw8Qfqy/sQn4mo/i9s9b99AGNEo+E3Yo4qidtEYou8cbiGQigQssTXydkRx9s2Xl9StcVMITe
UcEqOF/aURGXgfqWMRwk9yH5YsvVugY4BIrErcVL1g8YUR12mgdmM09G1qnPtiiHlLIuAGJanGAh
GYAtqZgYIiJAdX0ucIxFn+NFJyEdFBcuiRpwMwxIkmhPLcTBa5Juzh+b8wLz8HTtXa4UJSklX+2P
U1NJ6p+Nb92OfFR9wqWa5Jqes6jc/FC/cY0lijmfOcdTJOJsOLDxcN1MLs+gdNlkkPQoRWr5r+2n
Fc/i+uxdwEAl8ONr9ag5N0ouYHKtvehNnGGaJlRVPSMZX8waweywghP01MUhTzIdqzOyunSDAeAk
/zGAv8WJqGVdrx2kktI/GkaPGutSn9rfCCswpBoq+O1Lx0jmLzYFlF2B1psOm1+Vt5IeI10rr+//
7oht/6YkXWTwgJsFL0ktyAEQsy/t/aHrXFzrKH7o+2pY8J7mDQ+feet8tujDQrRgKRez03zOT2Wy
VF+vfqWBeKV49uJHDAmHPg1W8FfBh/91ExkApwMxY8e9ha9dEO2o78QB6/DzO6J/q++RljeYFqkK
KzVgoG30uR0EqWxFlmJ7I7nzvE3NyaA4KeKyIc8BNUNYAAujo7yCSNKtDJeeY2JBj/g5m4aK+oYs
PrijLLZf4vgLEXBV+Dcnh/50A8gM1/yfOYoKbC4sNq6MJT7DrYU0254qKrTDpX7E2z/vSJOdxuN5
VNLNQwHOmpOGy4jXNJESlYYeBYqgqJZlJtIHK/jMkBZTv0MEmw4cKy0uvJ5+ia18DwymEXfg5OwX
jKMhf3DFuefNNk7TYr+vKiDunmHoX5Kksp044iWvxcSNHym500OkTm9dvPKNWhfbzAoGYiip4eUE
ocspJFViRQa1gKEY/kDV95nKpuR+/2Qhr5CCVqiWKKjtD6+vy3fjehF8KdGkne+oSTNuONpBMwrB
bM81vqWxXfS1pIGeFu15fUgUcdDyTQMzTMhwMh/dOaRHDPtBNb4552LlDuVyVpM99C4S4vPmb4Fe
ORke47Os3O6GPDSz3t7VrY+u5GTjwWXZKLOYW4djQ8sxDjt5tOpTyAG0CralghXoWdC243O+vzQ6
yTiRML2/duvFOYbpl55mpiXi2NuDzmddlYAIx9SoTEbruA3P1LlIOhAZcALzg18Mz4OqV1hj3VK0
zKprAutoxZgFcojNpuEUuloyChXfjXWEjoWYY6Kg2EPzfZg/eogp5/EBrMGRzmHCU/bQX8017YjM
5FMZmRcWqG2XYxOpM55KRtSvtEaL8sjGnK+jGQgWs113xteJr5Lbc5G9TVGhLILr9Db7eB7Pb6Sv
wbDAuxGHe7SSjyUK80liALZs4IOo0Sl09DXNs5sZUrtUzNH7IuyV1ySETO/LjsVOvOFo72Pbr71K
V6PtJIPAnVz2J3Jp0HMAug6xGwDlr/ldBHdkvfvR22Ue57G2agjeNRie6KbIBUCLlehXicHktiGA
km65/TEdd2ME3gtaY5VbdY02iv5XIabwLVq2p/jKyRadPKofwH0AKvvn34fOasKE+DCLzzhKBrzW
Yp9UhkonKy7b38eLmCHx+n9kMcOAkPM9iixB/npQ1ZAyojcZm6dDpTcxM+1oCc4kJoaQvxVv7iif
XGPKGytMsw8ktLmjgC3osXM1icleuTKPlfIlEsExAcSNyKOCnytFtcwcjEfW+AAqLHV8DdpGbcat
x8f8p9n0vNhUIwD38uYqYQ63NlfuxH5SITkXpgh/j5o/Uz3MW3qo44uQQZYYR9MFJ5jxDX8qV4eM
5q9E5VAZAeLLh5LWN94YbMHI13YxGcPg9d/c6gLBGzNJmnAVRcgfQ0co9plwq+DAPT+jafmSTZEk
7iAi6R4SB95fbXV0wu9YkDFgTo46oHT1+FyKlJRX/wWXkZG36OP0waF+FiK3Sg7JAUq6gyG9SUDS
qMTtDSX2Orm4N8OSQoExJqQTRym8ODDwiLnvzzhQ6zrd2borK+6VUSoRkLLizB16e/nKvYBtKN/c
SH9510fIBMLGmTopGXGpEvug5YORR5cofilgFKuuvInqGcRF0daOpEmsoEfBWNofIJigp1K55SR3
DwufqiaxXEbeZsbGDzgXOIhQ/AYZDnmk8+HeJoIafycPqYZwWY1KmRP1oQk+PmpWnhTrJ/HtPbZq
eNzM04gsotoT61b7WSdR8IhptnVzWkCb8F88mTppp89iW+fV+j73tkZRIPU7fu8ErUgu6So2AFQZ
5iNbAkiZhLTh24SKkNukN5vsu+79/f6elKXSmUQgpeWamMqP7MD48M1CXf6UAL1cF1G9wwpwtHbo
c+ZfvHKA3Aee64O0KWs00jxfKc05UENmZauK0TMs4EyzD4fnb85FhJHVFAhF/Y5PouakY6Yz89E/
vEqYEP9BJg5RItmymDCNwzp2u5axNGaz3CeAEYhc5HwUE6g9p8mME27G3DcvGoTbjzSsRbKdh6Fx
ijRyh+UvETnR9/3R9r/q+Pz9UazY7DJm5Qa628Ahtbm5AJGZ8B1vTvGCgpLHBhiXKkx9UIfYhbQo
yp6fb2R1iGsisN6lsd9R+gQwojn+HMF/9N52HbW5W4BR2imbsmaWh2+dOvaNOz7ZLj+LWycwYOxm
yxUC02eNtdHHf/tuuhukaRC4adHJ10pA4tlg7GAifBMUbXITXUCJ7nXe7emBQQu54RCM76qdldog
t0i/QoA422rWI3xUNV3Hu3nMkCTZabc7GBfYbmdVK5co4RSP6D93Xa+3mYh+c64Wj5o2z3ce7ypA
d9i0JVSWQfg/9P2ospyyGYAc/PDvX6dl+bseDRqsBnH8RJZbYGZNUkSNTltI498e2Djq4QLAj/Fd
JliHp9msz0fYPa4DnPvKnQADwUrr3ln9KuOq3lrhKCD3D0XxEWLJ8m69nwxSmQ7HA57/hi9k84M5
8pNI4zU75/CudjAhIiwlGYQEDtddl0lhCkEchVDXCAIRjcq5pfonvivDQaYNwqpWIinKodEozWmk
DGuuj2An0nERNUdMotoaW/UDhaIGTpJLCxg2L0c2fgaR/ejSiLhS0VOCWjnTFwiC29nl/TLTNQNy
+T+T5/m/Gj/AAlAQY1EKHCaMNKdj65YqzrSqP9Tqlx8M6Qd1wNKxhl5iclTaIKqX8aNeSJcKtebL
C05q3SZvBPSYwfLAbdzXZ8U096pVny3zvJ61OVWgViwewWI1k+OmR/6MYmlOmDqAFze937cfBFnx
+5pxJoEM2uYkvxisy7+CnpUJSh0j9M4fAYx7OnYRb1r9XgmWZ4eRqe8D6EVQtiNkWTMSFwHwXfM2
PSjS9VEnfhDNKk4a8KSakS6k1FXvTeLwOZ47nFCJFZyoH0paLI4NeCjs3FwWxyKi8HXHpUDIKg+C
rXr4Ly7qZbBXgaq44j3gp0t1JRJXagr+IouNRB84sg6p57wNaYEQEV2Yy5q8Randw7koENrloMX8
GaVrOaz3HgMOOTQYHo4uyEDE5p6Jov4IGyCTYB4L9zAomIx+rPvrYD4jReu6Km3JGN3qXLL+WImN
CS+FfhMQncZw51/jCjk1Znrz3D7iSQtkNLIueqAoQk7D8TTR7TiaeFafgDdegNahJvpZii4qN/Gs
hVBkNcYX62BCKM7AZWTZGKF4QqF0o+ombEBbQ1d58ZLw2CyxGO0KajQSmX+l1xJ4rmAdAw2BaGay
S1bwW5E8y6gIQyM5mz9J7M8IvGfkSxexn/ZDYt3MUt5t1r4dPBNQ1z2uEn8X1VfKsj7kG1c4bn5I
hzuId9RzfSyn2CyIgaqoImB+6I9m6fHwZz4i7X61FoHa85nXdKAX0f5xLHqtFRZwophopm8sriBp
RWaknlE4YuCSr1EwtoHg4H25GhAe1/k1m8C+k9xhLE8uTKGC8JwZ1KVOA58ALCyfzutLxj1vuhpa
cbAherFiuURXfKZu4coSHmUQTvm/lKtwpt6N2QgnY/AcBx1JFHezOlHJWNoNeVgAdwWa84HKpKhb
YxGtdSIzrj7amhpqCAw8EkAaxf2Wloey7jlwQtcWdqOhigzGQQRQ4FnpLLB0qxUdUA4x9cVUwJZA
dZ7+D5o/SFwpg7sWJ7uULJ2f0jwuLGTholuvfFC8awc8Vgxoui7vKvHVFQsSpSfhW6+VeO6SoBEz
9Hmh9Q+1Kr8HTg35KpBOwFfyHxDAj29BDXpAs4eF8xPeOppoN+ie57HZktp0illPR5GPTo6DFxrx
wEm+SlWo8QmYFJFE5mchh2f07MI3SpnbrJO4a2BrUvdQrqWgqxppAgg1JI1yRFZddBwxJtPV0j79
hJUcfZzMlzXjdfVIy3ulI1FwAb49bU6mOBS2c3gI8EEX7+BPujHgi6ByRr3Msmv+V9SL4VKFBcdu
FWATOpZ66cZb8wZtbwjALKUcD36HfnRJk1HUmiUi0qGtXmbYVatGGDKJiBAnrAbsqIEzXZEGwMom
eaBeTpUepuBLx3LrtOBmKPw3tfoJJl4Y6O9hY8HpBy2uNMqGV07dJ3pXSCqh+GM6XvoMFUfw8fg7
UMee2CsC7NJ9wrpiYQmJirRN/lrnFflUeSMPpcrEeD/Si4/OGIC6UvGCTMHecGKrCB1yzeh1GVAs
CswZK4zfp5//eUzUuSxoMaVAGERsL7FNOn910yXpuBoPtetBh4P9/Gn8HwQLTC80/44VJCOPNM8a
XaAUmbJQIKP7Y92lfdcPmu13+7m+VBmvsZaj/RymiP9d7sNibWsQtR4TSo6ZmXPXIn+VOLjRo4hO
oQ2QQ/bra6Tm8H68Ti5Ka3t20VXcJcDRyZAJjy+IXj5IJHNoE2BesDaVmGrtCQFAO2WOmJbJm1k6
EgJ7pArTLWhoeke/M73BauHRiE8uGX0B/fUgSwXj4L8J2eCgif49SCS4eVv/bVV6/VOmt8ZDsvdA
RgeECGQISNob2ylkMpTy26UCwDASCY0yConDKONQJ7BLv4RfKXML8wBChdHAlrOHbXAoFFYPHj37
6WKDFuClEN4vHgGh4HsYh+wWabgiokBeS7Qds9KzcQLv8IAM859AVf0eW+4pduGP2rg16WyrVc8e
8i67xpMNJ87qTZf/9a9mo4POSIIa4heg0ZcKssIPNCsOOQxU4UBx66dSvbuUmLpFKTww+MNpNJvX
NJoC8LiqqTPVfowQzSm0wjCWQ9ry8gnzx221HzIzEnhZ0ugW5eb+1NjKzGsEheHyYd2z/G+Btgfi
E/1MhAGdbrtuVglSkmAq8IFWuRstzPA5g4utT86is9nNCAvUib/crzQeRZmlxGpQgM8/78RzYv5X
za6t51zWqlyzpKcXoaVmc6BPZZ1Izk2Kg3iOs47gqCACbHpNT15LKZS6F51k4mSH03VC0ux1WcnT
+5V0sQAWk9PNL1LaTrNt+FfpeTwmvrQ+bM6BjyqFpyz7Z/B4o3T3mOUCPmNY5oWitJVB48xaD0cn
3h/VqCeRN/yONkekH88riQvWXqyRxatmRFIo7Hs7W9Ao1Ev+LQp7RXJKOM3HEThQfr8edcB2RSnQ
tMyVOA6zmeio7PpopcIZ9wquYYl/xpcn8qkCi4OlsNAhyu6QulJiREoW7DY8habuIy6BuYW9cI2i
R0uWmfE5623f41oPjkuNgtDk3WU9TZsjm+2SoEnM0mUFiTTMmH3I+iwy7ikuk47g59I3fi7oi4I0
JhA4nS/EESIBXE0YbeBWrc4dFWVjMJ4v4qjYeuGKvnfvRqMzF2waE3XXkpwIM0ChWCOajBewCtNH
EdV2KNnWXxwm1Haco+BLr0B1bzyatIVxVK4Un69cT2Nta4pTtrXZI/QYucY9J73kSxXb3K4GBBQS
enNHreJSl6urKD/CgRzHkUS6quQf7sd9bVeDCfNFjJw5A7m2dZFqEnosMfWHBhZ/i4A5+4YERyKI
dbE3aEoRCf4vnefHXbxGBJiwlN1BZlotFCDI5L0rPr3X3e+EGfj58rj59qJmtjkC/ikKdsBKAsFU
8kl/hSk8TCCyePO6KXuGkFyCsPt4wcj0AOKjzNVTD6o5xQXy3F8Xxu4HOeRVrIJon+10ZPMZ8KaS
tjcuqXjA2i3AE6pq/2YDWimOQB/mYrVyoJQyx23Mad2hnw3sVllDQP60JUvu0eeb1Vm3/jywrYDk
oM4gKCad5Rj9iZNA+3YPc+5BHnEBSFc85r/lkCdk5xaHg/s1cDbLRZpg0DqLYq7kHbynNkfFPujp
UuATaM4AoNLOS6skyKnCz8W2jifK8UnHnkAcIO87WizGBo4JdAez6J21eAO/SHf2ASiKeCXyVIFk
4G/fGZ2OHAoxos+9CeGz29FEG0kxfBMCyYBgTf/aT4ZhMFJyQHUGnqnSDQ4tCx8pcmMtq2tk2BEm
94Ny/h7e7w34pHYgP0/iCGBNnjssOswGPHjP8D+95OKuA0+Zt4aZznLIDeBCofawvkkwXldyYRcQ
NfyANjyG/E5CwjaXF7mRyX+WIpguwqUkqkyNMiB7WVilxpRVsJB/XFEMJB9HwUP6QwrnLdHFub1q
0wmazbKyzBdXPbUHohcyn15A3NX32ePlc6pNZlgTpePjfDNBH7+aPcqMMGxd8Ad69dHSZejh5+pb
O7J1q/JUdxvM29bX/b+m3aFdAKKvv0WfwyOGkYnhJFzYG5dN08cKuuhGEc2qbDBYMG1+0AG50vf/
tzEwhQEjQSoMjHj9EeB9COhqIfOt+qjlOM1W6lqVJYddPWr331Jauwpvsv6VrEveUWHHS6aVaAGA
NYeGrlQN1lXmD2icKOh6p/bfwXVqcgGI7IU0EWjuLgrrgXp1Wrr3XYb4T9utjqvRO+/g7u9j6Xek
lT/debJe7O5GRJZPl4j40ej6UXWzT3HxSLK2HJtyR4zJjsyw9fFbH2nemRN7xwHEt/X56vkBn25P
/8AkqAWzNL6hRUh+aHGYTqczi5buXNfX4Tmyh3n4+nWIQip62296zDdvkG8e8iFnDlK+zH+0duZX
zO+weZ2XgnRogaAGvxOIOLqoMuUR+5T73wmb5MPHSJSsm4DpvwYcG5WmMcD/zZr4ZmJ6zbQNvA/v
MaRLQwaJ2ijBNcWGbTL1YEslq1oHoDwvOxpYGSJAcLNZLR1nZ00/nTDHPLn/XrQsVYMILerwOHdz
/GMpTfJGdnYZHPGFtLNpFFlr0w+M6daBqOgM9+tHP4W003sDo7OprjkxIoOjTk1Yk+8a/i/t9sf+
2IjEgas5wJCdaXYgP6VqK1QGAicMRk8pDWt+JM4l4JisfMC5RAvYajIJ6DaXbIE77txTPr9u0Ae6
jJ7pKbrF0+EI75QL4n642BGTMbCRsATh2uEEa7jG55uVRL/L+sRfXdlNkPZ7L1iGCAeGp9VoUhXG
cCv8+Iu+n9QZNIlAaZdt31/NcUrLXjRrl12+ZBHYehy79s09OIBlKnIXXBIIulyufpYlQpNqQFzb
JWaXu5Wu26d7dgxz0x6IwjPuDuy469kHPKxfvUZhBqVlf+CHKRPTeu4b+kckdZm0PtAr3DpRMRxn
C3C0OmpTmzYgkNPgbk1i3jQErDL7ZEHXsIcF+JkiUGR0w54bzI1T3LxPTwbWGMjR9LpFzy29O9TS
wfkY31aH4RMqITK95x5B4y0HpGbXpG6a0yTVdkRhUuToIhCDMeHig6UQO4aAymjYkPEJaOLsvtaW
XJbfo9CAoDe/V/lteq4XTm2bwWQzWtHml2ZBigARSzTHq3NR+U29Z79Ii/J5oUhXJVtWtWgFSiGj
hcJpMFcPoW3L/xnPdvkXtD6mRg5sIRW7zVgDQZ6/K6XInE/h7W9KXwg2Ua4/6UTQ7fftTrEcC0vT
JmfwMqTbosRa5wYTAfJ6kQjDS4/WEMbfBe8ssmIuSAgNjIqsIPEwQV0Rg2A4fjOLGS2+dVI7zLSR
gSIkzqrB8p4v0ZILq20yW3vp8sAk+kYuODxt5XIqgfhZeTv9HNdq0ggsxPLLmBhgO2DogzwdqfEV
Jp5qQOZg8T69DZtbGfD6NPxKIOOTCElT0Ey9LAcVDJodx9qdB+dAKUwvNvTSkd75L+W/Q+rFpHXx
I+SHlv/rzYJD0Xu4+TiamF+JV81XXnF5m9pBt9rixM/IqaP9zfCEsfM5MEd58PyGxU/dfl5VQ6UR
gaq7yCpL8PWWtIRjF90LpNWYzruZLvHNgmARwpmg/VYvHIkr6qSrjOH+nnK39TlgfLwfCl9oXn/M
v8JZaxupbwgoQP55zIO+It9B3/OTNLqTBYs1avfC3U8WCFvInFob6E+l7KvyBEcqhagsMdZIr3iz
Un2MKTj4jmknTzZljLplaAkDC7NgjzKdP1oBaau4h3dTzSsTM0szbpgHuH1aFxFw1JOAfQT/4nHB
sR/cJUw+vlirrtx7lKZOX8vGJXPfLctvj0LdsXMB5X8t4Onviv8Tj271CB5B+x38w2DdJCWFOYZM
qs+7ji9ppugm2EZbx8eOpdFEqPWixrEa/aC4IsG5mdl0FKeREcbGi/QKfiNEH9lg0VtnM/iqL/L2
HxoYiDyRvMTRg6fLEnqNXdgCMu2LvcNITNmgqY+7q/LBqfXxh7j+YgcTnSWtrKQTWyjhxtu3XmqL
Akr3QSimF1POR/JJ0Ge4PL5zgfqrZbsWUdMK9UBYBrLdHP5cXhsiUfXvr9soSfv5jX1/9b7TVCgX
TZw0OJTTsClNP2ZyVTu7juItMoJwgtgLZegacCJAf51eaTpH7aXS6U9BCg7pbyopP5tH7YsDkt/J
2xIrq0uuZa9Ug4xejDLdT72urLkoBP0MvhB+DB0PVGEthxrRjxZBcxXB2/WWQajTwynxp7gG+g4f
+TTKrqSBozaSEVUkwAwC6ozPq94f2LQxa7y6+RLT4Y5M4zJ2IIdeIKE/NMLjLzVUF2+CNfSZg+mb
mzcCGavuw+czBixVDVeUcwsT+tbpm//s/8uuPp9am1OgmRgNq/L6pqbJ8DCGWnGUx95sQaBmELEG
jhtHuB9Ak0V3CWNjyZESQzFV/JHvr3HW6HkK0L3WDWH0zxjBzhaytcRa5eMplETupadzO/vWwaFE
SacZgnnB4Yizu5UiGjdRY6BRq2gdYR5XTTNrThp6HTwpuQwAwhK2/yhcbhKLgzQ24DCR7shGYImi
XFnC7Cbd8GGrSfF2LHtaPvvTD908fgvIALOU97h3KU1uNfkIsTmFabIRaN1PpNTRNp57n2N10wWe
Ymy46QlRxUJvQ9AmDxFbzo7r8RDE8mbnIGu7+MH8ioyjwb047GIR7eBI8USTUl8p9gSD7splQGbf
BngRVmXNjsqUVqruo3eSMq4pi6ChnhAzCw6cc9WD3pQkLez4aGUNiUyAWL74zIS4QbSUPjxy5zgk
mniW6vMFX+XoEFIxsLR3NK2C3hnSwPjzHCEHvJJxXw6gf7U6t8ohcQgqjVaKAQy6WRSE+Dn+Prl9
exppYCOl3c6sennmLxssYKZxCmLIMJqWkQkFlB3pTxSud99J9EPy21j4xM/1fL4OQS9NQlH7dDOf
0Xgf/zFEtrmJVeJ4ZeEi3RuhKiBalQx1h7XNH0v1wgrgY6GwdCbP8hkiSPkVEAt/1DT1BhZutyec
DbX1ZBaO0ue66ntdfgoZJFzo1eM9xXWFpLOb0VHGRgvgotXVGUYSnG320cZ3EZYWdA8WhXLqTJ0y
v6GaXBUqSuWW2U3HlV9CrhpZOz5JCzPwOTdLltYovhEWPl+hpzhvRJPQz0ilHcGs1ZyftaMdm9Jo
zvDdZ3VZlm3cWj6Tj2WQK5ktCbhTnKYT4HfYbB7k3+li4ZKuLfMILo0zu5dM8B466sevB2C+aFKI
FEn6bKqJjBvBJuv/66z/AvSct9koGomoI/FsekBCixAMjNNuhIusdhcgfYBTzzeheDFQoORuKF5q
PNg1KS8pZ/CsEnHKl4wiEPdX0pLyUelLWjnctHae0VHQ748UVUgIIUHPb5uVy0jPoQkx8I1uFPQL
EOX6Whw44echD9Z5H+dpAYFVE4nbRYjTfa+CaoUjEAoPjNpBHKmTwQiKdVCwQ1UhsLoR9OR1cjR3
b6YsU2pAvbZ4pw4Xzfla+mCUnefbR2nyItO5M5LZDlm5B4UW7GkE2PWtJDC71XeHLpIN1FoM+KHY
UmH499pbwlqp+eu/H7db+xMkg9rYmYMWvI2BpPndHxZd65JfQBz3eSFB/v55Iy3pQutQgOUQkjbb
HC4DYmu7/uyq/JkFNP6cfbN+5sNBILj1k9pel5TU6Cn1hR320nk33njgcJT2zmii2GG67DMuD2Cl
NATZ4JQ2nQtQN2AIP/fsSbNKvDGTQ/4n3iHNXUx97ny9WYRib4am908u5rtOCExnvPNxGAjQkfE3
CV68eOJa6Yxuw/G2j0vzL7rGPuPAIU8kWvef0tellOcAN7tzx++vS1bnZyO8t9XEM/wngY73otuN
8702fhICuW6+PW4Nhn0/D8NVwFR/9uwpd3j9DXcwqjdqg+OmbE842sFueKbE7esswuSRHwRWLIIs
nNvb4G/fwMzV4a2LM2P9weua7p+F1sV6Z3/uNo59IkNbErSe3gOiKuNV4yfwbQyUBKKquGrM+E4E
h9mtaCAuz+wug5j2Yxdmjddz4OGeU8pmSyag6C9AMeznJHwcaxMaRa9iBuMjRsO8kl/pZGksxBJg
ZndaUEc+dTkaNzVTCff8rKrIXP7ONN/feXoFUVXwwYUZMqwE4IjCSa7MDD15qFE6YHNbXyqWwBec
q1EEL+f6exzRh0iU4Z5pStdG9uswqgf9GwUdu2vVfHb2NCl8/lbDlqs1dRfSVgMnrT7umtsoUf2U
fn3z4UsXWCeiPZSbHcj9aDNobbmxhW/ECLicFBaUiTuBTMd+9DFJR0pZs0O/BpwZkwwL3RJFDqDv
uVgs3PuZwmMugap9+Y67oBhOJvHgWJZx0JasX9FnlI8F9W7yeSBwAFbAnTuh4nloHZk0z2CEikMi
/AsXFjQev/lxIToLvSkGyP035aF3flqZUVDuZBuWNTV/53FGXKShRlutQqZgIhb0X6LyeIBJtty+
bs+JyMLi53sh6k+WKKKc2dmHhIiMyYhprPA6o9OQpX7Mxasnak3atR5BzlM4M4NM60d2LMQ93rwu
huZi6dnIP9qhW6OvKTDhpj+fu+TFC77e3c22MwUeEA/MgYqqhPnPhXRvgVK210aG65Hx1ZbrjCNr
OhNQoVSfWQXvarX/tkwxdlTQav35AalNtBhP6Q8FKL4VEEJhhf+40NQMEuHf2wC9IaYFu0nlINAA
FjwyDZ4jPlMDoaaVHVAh2IaGDoGXoossvfl412ok1lwIWHHZuubgOjRmEcuYe06WJF8O4p+VvOmZ
eYAgM+zuaVzWiJF2Pr3+e1ySwSLkMu2s1Q9l1DUrvXO6ziE+ycPuiGZfy5bRDTqKUhK8Gu4k9YCB
IwEKwXiwE07KrEMlNvkdaBFa7+M+B0w2MOhdkOD+xdJOuCUGwBP6KJ7DK58y+tohOqF0f3mlbVef
IabXZcEC6+/hgb+iFC9x0xQEYNU/kbqf/6kP2QVzLFI4VggjbOHfiTce5kmbhY5aSrM8jA2aDWwl
WYZHsoadfdDHuRux6+1gbylvQPxGKAi2OkprOMuZrbnVDlWh1OFPIQ2296BKuZ3tnPC0KXLg/AaW
sk9Ol9BBbw4ORQpjbvxHP5rJPdmOIPiLO6+Q9j1wr9+/ss3SStCeXWnCJTqQLmKD/LCEbhI/gShr
cYCqhzV1j8tvuBXWJP55TtrN69yp3nZ27UXGwjwwKVIZyj5x4ascatp6HLDrfZESzrkL00pZx5Cn
1Puz/eYpb3OExBU4cbkrZcdMLoDvW8GMpLUz738vDEVB60XjIC7gixDYizMQQzs46EzjHTpgLXtv
SczoZY3DbGKhFpjlgGgqdbFoGOJ2u80fd3DGdG9ujkODKvhYRFirWnGiLcJXaRvlHZymdyRcpXPX
rAbmEjNQaaW78eXq/r4EAG4HRttyjyhhcugp9vlNkD8YI4iiaasiQswglsHrk32xUW0aaBGYaZ9h
jnUtZbtwNvCKGDd1SnsPHz/MNidyLKvPHdJlLKYoHTKiQhzeFf20aV7qenrXDkI4JNgFGJCVTwI0
HYGH8QV+XKTKDEzQp1B9fqfmScay118Lk/IUZArfo4FQ5oqkMJ9q6DAY1LvmdZpqANrWFm+0dN1e
lcEdmWQFS2t2g/JVhekP6mCzw0XzILJwkjYMjIqHJ5WPVxgznGdG0gKFCeUun/I+o+qWlFYRY9GF
JOo4XFK8VXY9ZyE0pmc0ZJ8GVuGLhh64HMObsw+YK4qLEXf2X+f1cZp3rAU33tzQAzI4mr0BnZ3N
hSmpMvRJ11DKmXYjV59iP26B03yTS0Z9AVuFYLFq6yEwoN7jMbavaUqTWAimaXfN+wKEyRSKdcU5
zP/eAadN9w12DwNZYmllfwDxQYPKoO5LapH6n4b6lu+CoJdGPtpLn3bu3s24dHZy1jSVYprifwH/
EORrkU0d1uJSVBKaym2XNp1VDEmF0xs6s2dB5M0UOzkZoVpeE24esFJnRFZ62HKWY1Pt+9r0WHsG
eSj01ExkhyFQE1+W/1+1/bfudfpYXoZokkkf+bd2e2hHffcY0oiPzmCg2RAE4jKI2Jmc6vlExZJf
5wtWIl/XLWEZVZk8oPd8le2Wan9pZqIF+Y614vUXz0JQz+5E+kJazhDRthL+mStr6DarSPNQrJhc
EmhRpDmMy+PjgysC0boKqNRZ30H5Ik4GbG6rFpeeL7d9nSmL7rfdHh6zZbIEN07zIhdKcwkhqXXy
mgFLqiG6oR/tT/Xd2Z8fgJnx8EZfqSiEvf02+Ba8aHYIaTM3BOdqN9AbBzYKPL6XaMcOa+AQhxdh
c0P5pFZGzNTmqDC8rAilYsAD9h2aonLnGQSS3LCm7uNQJj+qTw2IPHPBAdSnaLoAqLEpfZ7xxRfl
nPvOZAI0ZDd2gsxFEGLJzfmc2E4aK/uR8LPkQJokALlTAJBWrdkNCB9OxcTsvHibFQdGeVrXStGv
FeOHFzIzeLjfUOvpVElqE8ufH6K7DRAnhcx4gOSbNKt7Z2A+azRs7fkQ8ecsjs9803I67mQXFxpj
DfG/A2++M3zFQznL5SpQqjZmRLFjPLPnIwfdgZLa6caJ/AuSlEMLs6CNHn6zfUjf669Ts9+kwZDP
HcJ6kKVwb3iC4ocYhLYd3h+Btueq9KU1x3HJM/X2TY0BFJd+AxndmARcJmRq/m2I2NF/ZBa0QgX1
VYMfiAW1O87SL0vAsZ/8cc7UEfx73G26ZWOVYUHZe4sxVc9BcXFnDMQ4sB5GqfB7C7HnClryvGIV
PDVEWOWAi6Jq/yfGs2JkJxiCRmx7cKF6lLMQNJOAZ4NGOETen+MpzdUUOoy/0luPfsaLEvbz0gMl
/s7E/TtFSoVkZ0hge4xQo3ZmboOErPJBNyphDyl+wvuqLV8ErwZ0sk42Uojc5rsQ72hEMvCrCbj/
aUUV8ghnlWeCU8s7OGVJJXqrcdOPOC2vcbPylnxmPFfjb0WvmkeJSVKEkdIaYnSNrVD15GvpmLdT
g4KCfM4b6lblL5gDfG3CiyCQi1LxMofXlw3L9v/01cS93wxSsrCIdj7X3R7VaOLG72if1LRlPq02
+ttUA2Y/vzz3N0HVKXLsgwhvhfUgNHCws9lpviKkZw1zUAAIQK7548VknMkxgBljO/iHmBgfWCd0
fqbVox+K74BkBb6V9WSfJdBt3VuNVp6OAF/KliNcOtoKsevcBbOLwXtRpeIrg5UScueTD7jGkLgK
4SQSfDFbs34AIQrLziKxJwS/laRXWS4dJ+2Zs2l8wguH9pmhccUQinrDcNmfs5eDyJjrMHqdRHDP
/RVQ6gfRxIG4DIDN53C6rxhpredLBwC01xPubcaYFwhqBUbxgh3KZ4xBX+E97EWKlwO0v0z2cIhg
hxzACIn+UiENm4+3g82fS+fqUJvwWe6X8KLKEvUJ4kLlOBMa26nT1cWUKjXi4s3JnIpPhih+st4S
Tt9JZbbwx3bCo8pY5pLCxcCXK93SY1pe7Z+YhtwQsJtm2sqBjillnPl4/wTMFc0BM/zK02QJjPaw
vHhA1yJHed2yQVBPeAj0hL0zmzpp1BQ0Oz/8ZfvOGNmsJtaX8C0VoN5phDXWBq8EhmOWeSfZ7Mp8
IWyCQ0ZHHpa1jLI1ncoqOqu5e+pjBnbxLEMdvK8v5dxR17qoEyeepQDZ52wrJxFkpcK1r6iYE8Z5
REga7VpwoW5t4O/DEf3pg/llq/pZROry/+SkeSFRiTneypQL52fjhFToiY/yPp0gSFQ57qJgsjEw
gzDNxAk9CfZt60s0qhb1QjymW/wnjSHE3Au7tIMrIMrCEfwWPFR+WMnvzMrAsFHazlTN+28IH8dj
WXujYxD7iOjqQRqvatTMvQdxtSMHTPTaUETo+iJ4gIc2qp9dFIwunqfATMBDmgEccD7SzVlMdq3d
u15YHiYGzDr9OX5nBopwJnBl/YsJ9eYt+k5/n8gge7TJm3DKak+Hmz7qperAxmbuM29YQ3vigFtl
oFFuOQcFVWbSBHdMmgGqlcDqQSa3WnAUpfjvluVKJHEMacTTL7T5cvJdErbqBt5X214DCPI1vW3Q
J9bKGxNt42K9roQI0B6efmNWY+GnnCKaAXDjnYCa6A0TxQjlju8+tqA2AcY7do64eTFDS8yKqeHD
D9wnBTRzWimINfGeowcselDFC3fV8BhyCYIADsSYu7cYPhQrJXYnsQRnFMrFkwqj0HzBPxC0VjjL
tGKyAQpivlY2gNzLhVRYWrlp/ubUgy47klmASQ8PkRsVfk1jB+/+fS/hvguXFzoxkZKwlWjrFajd
PAiZtLevjdhpozBN/hgXYjUB87YYjbZL3cpjeirqiVpJRBQ1584m3xvW2CBHrYAAdP9Gwc4bzHqP
/YpA9vRn4DXF21mAp6QnH8TGoOA1JFWtx0TMTvY36ufARMRWgxkjH6vQ7OX5CoWpQhbmtzehzsLq
yv9+GXxhQSJt49pC+1OiKZH2ZW1XCs5ideSWPh6KRw38a+a2rXbpdUqh+juR5cZoXVGe7BYFiTPn
Rmuo4z7zpPWBqBC9VVlvxcVJztt++Og4xT49sXo0TFKzzDCXOnJL2fEfo2uxH1+GTZC3fy3QydxD
VMkdTowKOqR9iGu9tz8msJT8jlHcs8c4ZZKhkcsl0RZPJ8t1r3MIUDMzagS+RG7TaVvuczgfionZ
UBkXzYU49RwvZjkIkSPO7rqg7cmpd0Tc7ZPFWbF5btQwyuvrfC7leAUUOdijrDXr9H0NJG4PsKiy
uK6SkidN969lHy4/3LlCvwe26ab413/5+s9zTECouXksATCosNpPYb8285YW+C3Mju5J2swZGl8C
hPelPl9w194UnCYE1iRij4F7dTWBdOO2rnj82HuF+SOfWUViSnQCc9rdpPZNdu7IirE8TjdcI3wt
Q850EIEnRGC8CzAQSMEIm0Kc8SsM0XaiLeMBeye8gnAZPFnzuQYDdRHi/7FwzgDapjlWBqjSlVx9
WodASwsegW/YYSJjqZ82qGDyxSDjND/d0ykorg3n+gmGroRVkNmqOqsbXfqdQAkMtpoHIvsmMfa2
/aDcrzV3AlPv29d/LfzPlW9auSuxvG4p+42ERTwwSM4yfztt/Zfd1wGiNa4EE0LALQ+emqX+cbM4
llUuV3tDs6fVWlHxRiXGl4JT8HM+QQUiQ923kV4AjNgDyB0C9I7VmdWUjXx/R0Aiw7BA2hbadaXB
wolHnITl4OFaPOScVHlD95ctug6mmUcIcdDrt3ECUOD6d0yVQF96ZZLF3R2cKeHLtX0jx324LqV9
+vrZGdDaYToBOPpCq4e4jFGiBwHOOgLTqo7ekTeAbbTsYqZxF+ccAqjrfDf5U0rAJ+Ta/GDHF3PT
dXrC+cCfm30+FyMHBM6wivZqhNM+v80sbGSgxVx4K/7Whgf3mh6+KQTJJbDh6dpcBCmC4V2VPqhb
OlXXdF7zQQ6VvbqRLAJ6c1olP9VBLlN2gE5m6m53TG7tOLoekqw6YIVdij8/34AQ0FYSPcmePNOP
EwqVdRh/QidIfU9EaYwhqh4b/0ntglHquA4igeAqiFM6JU1n8aZ/5JFEui0g2s67iCmaE58Azg2/
BoccvaqJwTBDLXqqiKUOSYvos56IKX4fI7OlgeWpcyltEjoAPaBVijuF0eVLWV9XrBsNNfFF76Pf
bTgdFuyf3osIvzZ6z4b3AtRLu8HI/8sNtpjD8f1QhbCUMBgChayemKTDuXbQkr0fZ5ZcJ+fKvz32
WDjfnliR7U8ly0IodLt3mbD2hJTtzT9/wg0kO+AiEHYndmsbBUhhvZ3JrjQ+9KQcENfHoXhADKFt
yKA7OAskHYjZWrKHJILx+n8m60u8Ma8nBvQFky67yp54cIPIvkJxxsmZd4H2EPZ71HsYZzRUrNVA
B9qkydmI9abkaEqHBPNfi64c+loXWpxO0vhNeu/G7NuU+5H2zodGnx1Kn8oBUv4lWXFVK6O9nQTp
62KdkwWFeDfxnXe13YKZxCmeQmhqxDmZzNverHqCr5egu9KhWqqPwtacvzxTx258UODLMwyAj7CT
hsiWjraNguMTru4fU4/k2msqk52bUYRzqJnvf9+D8CurAQGjVf8pIRsTdSBF4zSDHMe6NP37VJAc
DPNRrZaoOjHi6k0h+jWJLMRAgN1zLIfS66nElArpnOfODtOOhbDpC4bqHKlzHjgGGTMT78oNK+9U
o1viPwcxcFtoInQVZyMJFi1w/B1uoEFQaRjTqEeVwCjIiVLTr859GyHD7DOajK89SQ/HKK8aEnbx
PBRoBn19/z5Omx+Hst2pmhGeoM89RfnQ/mG/9IxJA8VmvoaAPmbhUDlRJFxjkew7EGqDhIbtr9oW
ffZT3LFyC3ZAvEDYNQiWOLUshLaNZPd/ME/Gge+LDn+7rDhqeHAesnX7o8NRMHtpGjzlgBo6ACtf
aVxZbFOYc2YYXemOVHUw2O7TRD1IajY8DBONjlwfl5MpWhR8Ir5LMyQ0WDF5SHoEzkZPokvMrzhC
JaTCBrHnQWGQ8xlGOgOoTcQFbG0XWkChgCGS6nHwtazeOUMZ3D1CBG6OsXQnoeV1bB8Jtla3/YWg
e61SJ8RBBg5l/OnVqifb/I0pNGAGL2x1hzt0UEB4sgS918YB4CBpHNJI9xaf11oCz3soJ41WXgkX
LUtg/whs4ZxmSHhyw67pJoOf3teSsgicCkWjKohQKfWLfo9VoUGTzFrIMJwvgaYiBQ4zJvYH8E81
T0xDfhGB5gHSLT1b/u/yRq8H2YSzqF4Du4XOUDNz4GRzVXQbMEiHTqHyrl/DOadkwt3LitNaLzlV
y4N+xx99VtRmbUQQFgQ4qQjTXN1RLeAk+oV0A241S4ypTvc7OfANoq9GucG932sXNkcuJLxqUcmR
Qeo7mvTzHznxf6U26fPGMPaVPuqjy5BDwg7miJ7IYhBFl4j2fFFxTlCP8B8Rnv90x7Yrvq0sr6ZX
gROEy1dBB6PSdimWv6QkLJ6OyC7+Qvssz7uyxUa2BGxEtVeaI8oqbsQgMVr+bkAx8V06TJdVrHUX
0/jeMXP34KhdT506JvYMEImi8J4a7mOXnmaAOhgshkM+XobYPFbfZHLhR8XTO8XZAFEOggEylyQ6
po71H9YjyU9+3F3ogedkqr4tWIpv8bcZusIoNchme73jZIuFK7QLNWqXBJ7M8DQpHTcW4aUKxzXY
04Cg0GPJyQ9yiY9DdhZuV9iRqK3y4Goe6nyVtcrrT0Uesi7Ql86Wmnyd4xQ31zGZGVbkalquOpjj
gnmLVq0aAkoKNonk27y+84oL8fxgzKxS0boOZXuF7XcrwSQiJLkS4Hc+WZFm8bZeTW3IlKn2oXCI
cEhLO1L2bhr8MPQy+8o/sAy801D+IZIS3fiC8NYTlOne0LYQulDZ+f19IwHuir0IMxtRwm/EDwHM
26GyztlBzLHZkoELpQGz3f0wb7l3xziEBXhE4j6cj8SwybbqBV2qFGMd07A2ugg11vFpNEVJMjvX
cqWR5gqbBLvDd2dMl/W5zQ9TsHaZyH9bMqwJLNdKGAtmVsz51EwJw6GCwnd6WeMYQBrP30A8dgmw
hEsssu9t3HznS+rpbqSg4D3ND5O2lyqAHUcM6XTTXOHZl5KtQ4sNogWsh9dYmBevjITyL46JvEiH
Ea1Xms8AVT3sh1k+k1g1AAnL3K2Lkw4CL/H9axhPWjQgrGsXNUgzSfHvzY8cDRU5fwt8/oH1/KTS
sNao7NvfIz9/U7MMw0RW04PmuDUGEDPFAgTITjYFcwCwNy2CgG+ZqJZPfJUGV0AF5bn4Cq7gymu/
fj/nQcPaGI9igxIVv2Zwmod0oKuN69Yr5fyBt0XzeHo8Q44DMblQIABqSfCWIjlQFbrC/9xL2SGS
KceejxoI+xFfaLo16UMZNmb3kMH7z935Ui1u2NfcM2x9SCo4WbK1yrtF4VamK2kbghTVP3pjUB7j
lnxxgWcRbUydqCXwcT+yY+CYBTZKz3j2vngSXlzIiSpR7wQC2Q3xg7wEMXqH9RzgkZB6YxPrVLKd
cvv6F2XamQ1AeJF1BFiVeNEXttX5roJponscz6YI9iIWQUgWGuLcASRS7aocdt4sZpTKZ5IqwoQz
7qm0tv4LeAjst+/JgkR2nmKx2Ok5OlM8cVY0aAHd+tcpPr6upurmbgdu0CtYi9O7gUP4vn2OhSjx
Suj9Wje52Awv9fFIuQsSwAnlv+dEFlihMftWABsh6SBGV0185StvDmgO7TfZ0XmQ2y0OYS1JIAzH
OpFUi3XQbl+LZTyzxzVj6wFkDcmHvWEBxWIn3OniF41j5MbB1VdorJltRlY/3qouoQ13qL+mF1P2
IM+8ozoAB/T4Gn5k0gj3K6UuqmscM11zZuzEtYd/ZYSLvgf6Kukvx7XPtad0VbdgU0SnJBzNEXZv
MF2M8utCaNFxDz/eRs96ErN0NYoXy+K1KNyNgJiFbEe3n7x2Kwyaq/OW1aELZ+8YVFMXKJnCNjek
ynQoj/Jag8pUu6IRpqygU42G2Wv/Yl4acAhoA2oLevtLCIGdaKnH4VrCDC3ZqHxu27/2G2ETFIxh
+gtQwgKHnfAf1kIKgj6ULdW54DOL449ggys4ZKCVZszf3ArM1qgdV2E/UccvQB1EW2xPYZYi60hP
qHSAEa5yGt43bEAQD1NBhoL9W2AIbEZ2L0+xzQ2JRddv4h5IuvQ4yF27GUL2198t6tFt+5Qv1DLz
YfWeCgEH72GHAjmFggl6rmq5G9H8X+NLG9I+kDC0i3YYL79kExxZTim1E/czxV4lxpXONU/3FJg2
Jzz9TOh1h6awga3fv3LAS3R88zYkIgjun4v+SdtRzOiRrMGlpnioLmCZc64IucrEdFoTdGSUdwIg
n5WfacouvHVxzKZyPpvl+DxYSKfnXR5R7tgLX9KFInxola1NONqajXKEFH2bEg4B20zx/oQRlsXu
6APskt0GlL6nLNe1KY1Q4xrM+GAZdQEMsv5C2y82i7UjDi7iThm67EYQQDqqQpSroB5jfNaAov1v
EMoAwxgSW2I2P82Tt/Z2gJY0axynmRrwbtIeEl9boSMaRlwDsuTqAnlaPyMfFC26OnkRX05yBjKn
iV+5gubEphSxU5mhvTPYEmiIbahlYbUl01dVu+kGEbg8BzAi/DJedRATHivSEL7CtrSKZg4ALEIC
VoJ0f//7JqsnFZGqO+4K2ngGhG2xfL0dSW6xPMTmUHGpZs++q4wYtWq77hz2dmJIJt3qyvgMQu4f
iwD60SGW4mrZcaF5zE7tyIa0OgKn/5i9Z5ZtzGFrMWmsjFcRoM20TjzwxulexVrXPjXfjAEr6Ct3
H+7cADh7EZbljnFi/AyAdSeNDU2M1bQC8WOWfixaPJqqSivUzbRDPK7epbTdZpVN2fd1ap27nQgY
O8CKLx5mLSuekroADPAozjJPUwlKtXDK3v53jOKbEkErFLZ63w0POhawcklkvwqEOsgx4X7W0KNW
v2Xa+tem0ITkabnQ8wPo5pvGNYPQevCXnPMIvHxIADMtiDhitk+SJWWzrKwiHpaJ+RnkIFDSngQ2
3WwTrqZGMbUqui7HY8bq6r16f/cLZFe+LQbx9NHyb7X0b9lUkWzSSgvaI+jiosaDlIM8Z+qnOU5l
iXZyKqZhdKZ+1Ic9LDnPKGVxI69mzLwf1Z7nlcnb3nQ04Qgsqu1eXlOys6KAabzerC6v0e4ktuTr
Zy6Iz7Mtg8dF8WRv0LTas7qlCktKdG4K7QYHhv9apQ3O4RiCNyN4e4qaWx7Bq8m0qnlmtoC3+iKv
dwfdwzBz3tmc3bg8KK8jK9YSqUNPtOXKXaUQ4oLsU1WhrwpfQ+mXwqpQX9iTGpjgkbDg0tdhQbxG
UmH7c6KNOFXOsPrJV4/VLJMH20BLtmRM/1iOWiOP94C9zGOfDfwmsFKxi2HgmLa5ZfdvXGB+4QUv
l5gbADOYIemOA6j4YDUFXHMaeOQ+1kOsXWGkSPltJsOwfBSRClXQHrpz2fNxuflGvqY/bFIIxGCH
In/mfbakDyP33RAXnSfrvj2UvFcood2afrOaXqBHwKcgCKZmC/j7G75DlsJjUkrWrLqxwPPLBtw3
HeJgZ6WknEGosXIVAIoA30IdDmSBnvU5w76zFvPD34Fb++BuZpljBCljjksg/+GtxlhGpRJFpfwK
FSh86BFTy5hjVoLb2WH8MputXnkdH3A1T7dbzfcCiSF8yjTe7VnDKyKuvvlQ/JBoXD2jaAgCZS9g
/hqSiZ827ZzjPbcPa9k7UIrx9QbTyliun0CBJhD6mPt7KEoH7/eopPTRc/BlM519peTWnOEfzPU4
g972NBfV7NM7IYTIUbC5PXEpbxtnUhOHp/HKOOEMmI/WGSvF+q14cJrQl1L6fzk1396qXrbprf5B
W0CnHdFM6Q3fpNXOePc3VmO0QNanfQmdNR8TYGw2riuNMUNp6cpF9snDy3oUDgBhL7yWopUfn9XO
h4xcif5XeE0sGzlVys8cs6qBZzsj1EJ0HhhL6bV/GfLXJW2xiqDhkCPWcgBiFgA9yUmtvg/HglzR
NfmPl1U5w4xHAyi3/dZLFJ5Li8szM3+nX84XLrV37A+G9UrI6gM5lT2FxQa2lLB3qRGpSDqdEUYv
do8KG6YRlFMn7Qv6qV3Fxm40OlSAe1vOEBHJXooMLCw1VyTyUReLU2APFgyFGyNY432P3FUQHChu
i/gZPeJKCn1CMz8XiOe8s7iinYTg9d49GTaqJF/lN1IWKOketiGVH2aWg00FbK6l/p260Xi97iN7
Yij3BBU5ND0OlJ7+8/xEUFfuTWO/PLjBaaO8AQtY8oPjdH4UhvtGJRwJilPy/410YoBianSjTE19
uaPGQfU/2EV/87BBCnwWDK6Rf5z/K67VNbvOidttK3XMYbQOVFZCnluAEXtHSEBlwJYFFOgzyhBa
BmdWnyX2l4tjPTrI4I14/KGxClPL2j9HpRJ3H1a4E3WF821faOLwY3xMld6BARb49awen08c8Grn
OHoFV4OaEdPV35g7R0mxNT3pKdW88vszyJsbN3HGDjQASfOqpBEZs+QtB/Xsg0nxodTFLD4qQDuk
1jGBnv6/8UEjYs6Pm/XKWlYLbuiXMClPky12TsDRSRobWW8cIJ72YetuaQLxAt6R1vKsZQSYuXVe
FP+aXo2OlwOktG4y+FRa9ArFqgbl1kFlGl1biJZGxWl9KdP2aiD+FSLQ907FlT9DByFvU1gVqQjt
S8WmhZttGH6D0A1F/2kCkO+/im4xitn+SrEqGh09nUEZ4iLNk67HqR2TWbOyzWsGYHR2i/QrXTSw
4vqhGpeQ7Zkmbw2P2lRw3Og6+JvTZGwcgxoPT2O6cW6XRfS8Su6OIXS5cPLOFTbS3Edk0svcLfdY
phghcaBF8n8yILPU5gSE4htMDawtYrupDiulDfrnWYcWcIQlTDnw93NFA7X9kujRXHJ8Ts4hltyV
kvqcEStBNBDbE7GV5pOuasjEXFlpIQgCK7W1grlVKBeDpZHv21UJ26EJ4W2NeDXxUfnGV3HkUc3L
4UdCQ4Ih/Rqv0izmsGWrDcqBnNTW5bpEx1HXkgXmUDkmeOvNrD2bpmwL7YpA5p2cjK/TSZoY6f2X
uqzyUx+IBpPeOxQVfsWPs1ITRPENZIIHFeMvpKPptv/TRT7WksNj5gJkN7QTbFJrkvYlKS97AoWl
2XKnzLdmbUQ+Xyu07DL9mPSov7FnqH19ci4np2ztKfDL/WQ69ICMI8X2mS1twaJs6SL/lXXCG+1f
+HhupRy+9pWf4jGjfxSzZj+VRKE1B+bMLWQ9vRIheBd8G1uJsCsyirOCi18EoqgvYo/91FW0Y2bE
rihAcr+fiZ8Bv1c3VeTCvEImZH5SipoZY6WGYLx7Tpjn/598nxEUKDwbqaHRr2IqigcI1TYmoD6Y
AoJeBDcKOgvI1YlgYqLks38mfsWcBr2xs6KdRZrX/+30hC8WtGoj+0D8CHdVc7igbSh5pzfx/l49
dU5QyEj5S13Cc9aWSoT3H+HKvgPcOaW6/FbwkS8f27nMnIDO7xCQsl4neRGWCn6U52Q0TPZwfzaD
RCLQeXrtbYD1Pius+h+Q/GGSYadUMKzHLiVuFpqKN7uYQs0y0s4r6c3geo+cyeuPzVH8ULedW3G0
D6H/xXmuZ0s8YEQBTumCmF7IYvgN4L7rdMYH+aq+LmREWYOLq3Oerfc4dbvXagOiV/NK6gjVhFUW
kBAeTtWyKrTV651moAMrY8crDdOhzgcCp92DGjOMSsoZwZtuRDkKLdUJ/WXGI6AHxPAWyJQTi0Cq
hl2xu6S9bmFXdN3S8frAsPIphdpewe4mxGpxe4MXg1x3SDvff1gE7vTzJghHGjKkqDYXx+IkipHH
Zx3fUEapMgL5oPBe/ugwm+jX9gTzGUaBHcaTKzTHYtZuc8Ryqel7kclyX6ji4t0S4aYXisSAI1IQ
EAuL1qpuYQYagUxMRZCB3k6igMvP3pK1RcUI74JEEJQRi/Az+ZpOMsjlodN8SiRNDaXs4E/9fjuc
Kr+rPxreLWHz3q+xMdsac4KD2biXRKPykMcwerB4P8Q/yfXqmgihlOB+z2KlEOJEIjsfW8roDuDv
49VYIVGQHZEQvlsUeUOoHuKr+5xF6RlqEFpXyirmaXSz0KT6Vf2tfledVZ71gFI/qwNxSCALGG2J
X5wkQWCmqz089pdHxF0g8cDJJYU9LiQKY/0AxZyeEa+n3x1MAx+oGbDfckcHsX6UMv0XReEiyFn+
jONtbFznLjaF9UscaL6PvQOfdASkfo38+PTvAM6zKaK+GJI0kz3GsWG3alwNGu1PWlt6/QjtSw/g
LVwCHp7XLDRouSkHWDJbxwVszzw57IBLTgwY4Nz8GY/6eX8g49UdYXSIX/3HYDsLw3NVp8WCcCjR
XExDwyIiVEfXn2Xgpzt45UJkvf2IW29EzquTqnbFNpNwNU7plPb8gjCcEjdijaIdNJSAhZNEXKKS
/slfm8wMfKRQW8nyi6aQbETEl0veLmLnamVt/B9NUs7c7J6d8SSRZBlgJ93VZ8WJoZkRNNegfmBs
fN/gQofviLoFPX91mPrJkzgs9qqnicloU1Gj4w6oc5v/W1qZAfK6GIjGa8QRm38mm0Du2wK5iVPp
o4odaj/JibEcpAWNRHdfSeruQv68wXzOhoat2HTRmTsLZktkSO5vV3oOBzNJ2zR47TCXSCtxH4r+
94cHFUQND53FOJG89uY1ZahVg4GppRCjeBVkuCOC20zix+4uiXM5SshbHz+FlGpmz1EWPJe+Xzai
wEQclSIN/CaWRyHnrhVJY061LZVFJhG7S8QPdYLYDC90Wwcc/nkZwn23l7ENpa383Zgr652BxM04
8rx+aJvlcwqSWRJXlQgo5JE6aLZxizymNhUPoFQ1Br4tntQbezYzXzqkEJqocUa8IbrcUVzonUA4
0QAfvRkpnlOxQCb4avQjaEr7k17EDaqkn6/MlxPVL+4tFlHByFKeMrFIzB0eY3OzQ29GVFR/w52o
S31QeXTeXUfvgRNfKIlQ9P6BTdqXEomdduOsFWIheNkMarDMZDfsMMTuZkkbEKvpmb/oh5aDS6yC
FccoloVKCMGSQKuTorJ+d+wqKvpha/ms4+evEK0z33bH2woTBlZ8PnazjEvS6gyxTVsHRRBotznl
CHLt7q8G4WlAdNnNZS1CssAdbw11+e7kvRJZ7YvsPMce45JCbT+9NJrj0PWRa0SIRAly/nb4IVD1
duO4X0B7WaOtm2FnoWVbj5Ieb8sK3Mr27pNWN/D8bekknBT79TQRcESxc+DAdzTjWDdzdyI378lY
NLf6VgTGC7Jkt5xSoW0jpKxfknAL0YTqMWzND8nwlHl8KLNyoQ5jW7UMCb/0D0RVKveASG6xuT2Z
nefo1YTlGcohFD19tUtSHg6RWLsoAclWEtV5J6noEuGK6BJ1nkkgUJ7npYZMHcmyEioFB9tYxwP2
wHedH6AoHMv0dAPuOjaAFu4MrtnCe990+tvz8D+pxii5uh/PI8hlczhfAl3UgnoPIaoobvgta+/V
uN32FjHR2lBSqA5GZabIY2qEzBgbeA7h9D3sEeRcMsIl8K6FGsJqADFb4ghfEnyJV3h9ew5PwzxY
w0eyhd73YRyYVCZo0KMQ0S9d2M5Zp94XUtJXrxpBJkEDSEZ/qZ/d46V/uzKPeKI2WflHlvX0qgMZ
csuecgqjCOHW4pBhwK/rMWyjvN6WnU7Ftf35abtQ8KYFZDaAm5TO8rsC8Ve2q40RX0Ztv1HN4PoW
hLojxerXsGk95Lnw6RJwtCk1osYPbKHS4ODjunnDBGwbwsza3ozKeAL5Y4OkO2CEdOIG8jcV180/
aRnF5WWZd4qno5S9uFbM0H/F0ZL2HBk+2AiDcmkAaOhrJeNc9AWfYJEZa/FXJfC4jSkhU8CEAep0
RYt+4xk5C36kL39sieeHCUneVsJl++wrssIcyUwe9Nuk8qQhgFP8+YQV9XeHAlZPBeozFTQQPkG/
yqc+6dtmtmdz1K+UNB2cF71VVr+Lm/6Z6P1qocwrNFDnqpEtZX27n8Jnks20r3ypF7Fp74TmON/p
/ifg027nnjcWV6FFK+5wDjdTemA1pZPXJCDxquKKFhmnRcWTVNQQydhWyhjQHJ7L3W/elUseDsJ9
MCc9A9jTrB51Mfuz+2oLKBPf3x/LE/+4AQaLBNBk1dQ1/srpav7IJQqKaFONBnb0WdF/WADKeOL6
/RsnT3UEIoK2ofuSirnrKuKa3uQuaUZbA8u/oXI+EfDekOSZs7BvBSiWrj2zRwCBGucsS972Nj9X
flKWIhp4P7QsjcPDrBfozk2W1pETjTzj4Mibh1zfdTq8BWfwvdppg18nLEbzHM4Z5wui19LnqA/k
lhGulVnLT979Ucuc+9HeWeVRFXXODjoXiyUxjO9i/ng2gf5BpRETdc33Y8a5+R8/7FBiFe+My3KS
i/ENFcF5+YmzccWv+QhfDvbnzG1WQxkfUN1F6QQonz+kvJ4KP9ZHI/fKPmteyZodcEykFWNvqEjj
gcWkIKe8WwLMruBFkWEPguZ9eRmPAQgwopKMlb3AOWZSQhC8ZPWRiyPDrs7x3vGStyu+pcqrVvbW
3oIsr7ve9/3yy/MLlqK8DN13yARMW0/vzf0ZH6CaGlNObRiUlVCOYu7GzC+Dt9sItgQtVdOY/V+5
48mcJKzaxQOpMGJr3r0cIPRlhe2ORCakZjSgUjL+U11HAILLjWvfOAk/Fla7h/ua3JKSUadKZWF5
BpW8/Ekns0PH4mrWKig0/Yvv8sQkfaX9TqoJuwefk6//0kUhIzQLrrhR5DKyDRHntPAcXzGgmJfW
2l5NwjgGmhg5HJTQd0pweuTKk8XravzuITiQJK9RnU1uO3V5vpPLy1lvsW2/hGEj3e0CEjUfIY1I
qu3qBWODcyi41gomINYyVnVNkjt5RZmsr6oPi2q9UJ6hpw5USXk2hbfp+wafe2pTglvIPEcIv7Gb
q671GScEwCY1pSo/cgOnnKU4GnYY7QnCzwjUQcd0uYr62tvBXI0hAfEcZWmesvqJJ19SLDIHAoCB
nJF0ddWgNKkJWOtkkQJwB9dZfAROnqKPZHr8NmvEHdIrJVYoCLZAJAemPcsVfLMjmtFG8qwz27bo
gw89tdFbS9FMGUpZTJlO9ZQOSGQqi6ms4SFgbhBkb4lhrjwdrf1fWIKwsWyFdmhLS7enEOfhZYOx
RIlEPZJCTGUA64LWAR9JWWitPt6jcupT23q9HjXptpZla4XOx4555NyoF2gGrk9a8kF5grYDBZU5
CqYpS6UbEUc+eAiFFzDM42dWbp/QvoXeyqNR19f45tPqByREmIDMC0HBGhMh1Micum8HBVLMPK7Y
frr62Txe5BWc0EqNfgxPT4s4JyJ1YqnCDwz+m4vqGaDAQhbQHpbaHs8eVrKky/1ZdTQxpk+PFLMR
aDsnHGlucp4aI8271/ARVIJbq56bYOp7x33UC0IJSbUJLwLsEukPOjviMoIfv9VFpHv1oapCvQtn
MYi6thBBUgpcGRDLdrPGyjGmYqBvbK8lak78D2cEkVso7EhlSrmOp7lSNJNwP969O41PFm1lnTGL
MiWaefndIKz0/KAbr/NWa5JeNu+lap+wl8bFlRM8vmZInxs8kEh/goKMbmVUiv/PoBc2BGFxES2y
f04H+7P4PGXXAiPFHlb5KHlT9fgMNM3znZoQvM0H3LibSfzt6qAx+XlW+A5lE84MFzs6OCIuYG1a
V2Qp/M1vcqXqbZ9BMgk8PKWKy7xmBfVhuuiCvJJuntPOpQ9NBwiDIVYbWW44QjmCfqV++1lopFps
w7z1MrYa+qzloxBaS6j14XRP7zgvhXemYKi4phSdUkv2Zd1spIjENKo/VgN0DdbRHVaLHC14tf4N
pwxk8jviqu5uGYFO1of4lc3VUSPbtOZxDkhCcQmHnOcOz0E2fMofgdsJnAQGs6sctcU+cmNdPvNy
B83CGbU1l9wRH6a/hHdERwzfYcKJEBykBdWszbDFWyyRhj9L7hH8D+rzayhM9IIbasZXY/Y6nFYz
V7sTSMOchKWGSDB9ksH8NGqKOec0KVKEtY7FV+x48An+v9IZSWG9quyemkQoWq7sOIfAF9G2EfhG
PX4d63pzVvrtASUaGbr2kAsoJoHurfpOIaAqRcKPrm9MPnFJECH8tWMR1l3W5W3hay/arABLIpYi
HZxzfNqds5wT8tnDKqNwO+ZwoDNRWWfdUR/QUlfKBD4GLBnN12TWoHHEUzyyRRkrRH/LVgN1WJAT
VK5bFwIlP1FjW77V4mRrigk8se/MX1wlnrC5FNJe19Y9IguNMnh7WqJ/Qaurs31JEe2eIfoFf/oV
kamArQgFFlwNWKDDDX+riJggpDOyUGOUBEYMSbK1SHrhu9O1Wok5KIkUNCtpMWKrhJ6KmwSFADOk
s5akhxGHV4/Z8eKV4EPD6J2V0Doj/a5hLYkry2UjkvOp+RF6zBZECSXouBcRi3Dqlf3rQfdh3K/y
P16kyClqcclpK6Em2/qimTxhxbwffdB6SJnmCc8wIfDQrA4rqSiRAbX6nl5vZNl7YcO/6h8lkimn
NrqrK+0s+EnnPGive/84JSlmSmN5fgmDnBfNmhxmjKfKlE0XSICx1g0Dpqj4ljv1kubfY+3Yi8tt
i40m7GxXagjQvpP8ZSfxBB0gzcnClK46R6UE9DgH9wBDy6eikORDvROHhMKW+VB3q2VyE8UFbw0D
LC3PimZCMMmTgxmhfQyiG18sJiaGIGDP3eUVZVZcyc1gZ1M4r3sRx3k+nUAyG4205z8hRN/ruqHn
iPxmnw4CmLP6EZIvFTE8Aauxr/H0yjQNwx9cx+gJsspvU1TOGphkiD1F5PTQk8Z7oRqEAJ/wVJK7
tk++RX/4igGuno4WgVLIi8Q97IMqlxg/NyRsWaAH+iTCnN5Q7DjEZwe3KnFM4hQqrjHAAstxsjSe
TWUODvylQyBs7QtFjxkzcrOkZIBnjuuzsAD8H7tggjy/cuccc04t3Auxzi/F2sM+TWbGqKrvOPxl
IW8Sge2Q/NnC08uwDroHxdwWVUJZcsNpL3O9fyljN1z9LF93ISEWzub1lPLrHghEJiMkRTjOxtnn
ooSAT0s/RWxUJTjnDC7Euov9pWzhcvW2wWxqUBORPFtSZiTQCfhJW/HFfyD/tvqWo273xr8b0pbu
vNc9Bhj0wHojNw+L2kQ8GKgViZgTNEjUV+/QhPVK8Q5wKvg5R+acxx9At1CTIvRfsM97CB8Pz2Yr
EZGQVIO+iX9ixOU1IkTBeQ1mnsytTYaWBDVdTgkc6KTmLAH39cloGLRiKXbWpMvlvc7SMnYCb/GG
vozWVbd9bTMdw8hoPjnYMqz1Lxe/rsn3DumQNB2EM9BeOO2+v+3syrZZT+rZvMjeCJayS4EMJSVw
SRNuTwfiVskwBu771OusgTwxyStif2k79DcBDKJdgtVEZJesZn+ykaFquACskmXuGCIzPzLlEyC7
n4HRByhndInbte8SZioSPh/o5MHmKBOIu4f6bzETQeunAHA0k4h9rP2enoNi+Auic+bacqFQdIKp
PZ3w/0qGqFZ3JV/i+9aqu/Ai7x+U5D7/Jo0H3grFy9iXG4jZJMTg6xXcG+yHBJyMhTFDTcibY7Ea
jfvpWr7oCGWvieTtuUaAIS8J3SL0rVTrEp+raLKbcXB2iPCn8yJgi015PgWpuEM5K6zcq1FNSP21
TRGfHjJvXrQkNN7NAacKi08X0dSuh0YfTXT9pzN5aO1w1+Vv7ZCISMUDswpXHQh9sGpWHvOuQ56i
kYxGXhx9nNCmCMmpkAG1ggIAx/53+ewBrVcl2bRfQ0z1/Q65I76lVMkfCTrD4iOxWPJG8JmCRpy+
P9yWH/pnj5LCHJiMPm7+cZ6f6pAdPjxKWPfarXSS51wD+bm1yUZy6pxC2hDgx+rCEXGBqvqnK0Ax
nxYIMq8UExUcF0sBhTau1NST1JQjQRhmgSCcbiRK3SylMmq0wTovhtzBgrGg00vaJpQPo5IbaZmh
Ky+ErxJxnt3P7jqIo/GfZdCpVJrokPW4BoZtGzr5DS7my0Qp3xn5WeXmdDpXbTXPWNEeeQLN+WOB
IPjQjHANKuKBDrMYHpQUw3Jmnrz8otKW16kSZd/lO7auOwVWeYoaqWu82sPk5RVJuKb21M8JV+2U
yPnKWjfNtV/WmVos/Mca7CiZqnkVTJx2STWuHQbm4Q4QHa2ll7cXAdWK6a9G5saflzRNRIJ2GT8C
u4S5oOpd1E325ajHRDUwTI6Ses5XWCymSmUwpVwJcjjQFYPYnc/YJPiXH9eTweKQVK4bVcxWRIlS
f6qUomfXPIjINEqbWuYCvq8YZyOaOONOd3rIscZv/JrU9VISWZfPvzmFgWIIVRiRgHPOGHQwurXc
SrmWJOtrCAFeSxEVHikqHYcDtdljwZgFDlTflCzopkr4d9BZTC+ExUNzC+a9xSNVsr+CMJYDLrfh
zf/MsVHpe9sAPqDSU57ZcXM29NIdehIhfFhMoU7aNwHMA2AVFo2COyIYE62LAwBmC/BhfAUd0zrf
Q6tAfB7tAAvkkGgP7j9lf7iWwfi/Hfpz4SCB2TLyLtgTJM855r2qVfxg/JWJHFhzg6O/TxmPKgXb
malDC/ySt3NPyY4hl60Z8ZswU0QIEMA5rb976clnH8FNyMXSurOXttbzpfi5R49tvqnkJClZht8/
kp88Oj8H+tUiSx5aWi5Hg26cgyaruvhA9Azu5A7plOvy5Rga2vFzTERXHYa4xsHJ1jJn1A8lE2O1
66YyhVkpLD4Lri0o+5XmmQS9nx3AtyzbkB1x9H8YN9zDuToKfyg9pOJlWAhYPoKxmVjB65ohxOgS
9yNLigJ/DI+DSOAPwsWVAapdcsi388kx57W8Wvvn6VX8qwFGknQk4f9G9WsYeZPIdPsxZW1ybc0p
cZVdzpQWL5iLt+qIMD2CaxT7U9zmUX7SMIpFXB91ewz8iQcQTBLLX9xWSs1Zc8BKwTkKwpxsyRwN
SwmS+rDdxnON3snXtb5OU2T11sBf6Kufb2RcQjFMlB0YJtHv6l/zlunTVhuSthnfH+QW5ZK065eq
pfJU0HgSpVAgf3GimdpGup/xgoQjv8325E//HsZw821QbfceczEPrNdE4emQV3QJZWMQea2kkl0y
4bVbB612sa58vTgW8HOxnhbQnw4k8wkjOJINQDVq8BgKte8MB9u/uyI+hJfeNuN6SCbiZ2uUhKoH
g7Vyit3U9jYRlAIk5XjGY8797FNantBwHCmV5xJwO5nRbtCS8aSYsmdFw859MBqSODDOdWOxAYf1
/mxDpyj39FvceIyccCDy4vG2sROxzlJM8brGbl6l9ARUHY9d5gQq/pOdkjw2Q5L4Z31ZAnSD+T9E
Cz8MYzUOoDciXjwDWv+NNFocjrBOPqd8paITDMgnEbm00JgS2+RkU3XjNYWmnkXYUvfQrMnfkxFu
z1fn6ewAkb1dn80qLXaIzn+Bmkc9voBLWSjw9IVx6pZd5ZQBtdHJXsDWLDFzs6wuDcT/nM+sGtLd
WRl+3qIBO/4oXIlx+qh74YOhPxZXMSarMeWKtwyvnGLxo9PPjEHp8Zaxtfsnopmxdqu8JEuBX3De
ZRtf6Ja/FnlTBdrQ4wA03bfEAHZSwmkNCz5dehPtPmSFzUOu0ZEXUBirmD81IWhxpowRksK2f4zh
+EYxmAhQU3Cm0rSHE7SAuPXjS4LdPW2iDLbQa8Fb4c7D7Zn1xwy6VWglw0yoQ+cCCEzYfNaYwZZz
sZwQa+6PMT4QSp3aX5HYTZ0rSK6onpJ6VVf725nU1dMQpunC1sRbmf6FqjIrinlvqByJbjEAWV63
8tSRlzOeBPGzy6E3arar5z/EnqdD07QlnP8VmRzfaJ7+elQTcOJUQSc0JP1xzpBLDXi+yHRZpqfa
Zp4bKOOzJewb2h8ZI8TjEwd4mQpO/eyA8ZA+8h1xQnrwsoOt7A1U13FCLBW2eFVhID+hrZmCW87n
LTd5Hg7lftIrmzY6gOwEgNb7Y0biSZwv6lvxvPnPSZu4526dFCM9wdwKHTdffzk6lXoDczXpI1+K
KvuJryxnhpGOdiAR80h3vMAasVJVbeRrYYFsvOhXcYWDeW8zGdIn+uQCIHQ57rqXqZKqcCDNX8P9
krodS9gEPoXJ0wilBXSK1E8Dk13fzAvSxX0JrLgpUCn7Qtetze2jrgn68eliZIgV465AFFBWKdc3
DLMViQycRpA/knnykvQWAQZD+O9UhB4gWquRFqf7wMzlf12aXDDZ6JuBIfwrnfmIsJl2BoQ9SoGH
Q7B/g/yX8EKIIMhe1Nld6igkJusm0MjuZgUdGAIHgZ17FUBnft4sgXfzEKOeNNGyzJxC3gwAUJvK
/oYLmTd6hCtXc72j0m9Afv3ARQAyfXEP23U7+uenzmOzG3lGV0EdYinG342ldw5SF71GB9mbisag
aZxKVXm7MHH49d8RTCO9eexWMCxjSSx9O+lcV+mgU6SUd8odg1bWsnVjXwjoGUzAEgAEKW+L6jgn
ZskkZ0DYQkAuseiYPUe8C70ZE9F1tz9kID+FrJW5MAd3tB/PEHKrwHdataWernYjC5JGEleZtIU2
8lBQLR/gbuPnufAQWXklmrfcredh4eL6xkbTltKbs17hGCj/91Kyl52yzQ/qjA3CNkoUOoFEXjtu
SY4sLppNwAOzefDtsAt4cRmofGR1jbwuE7F3wtu338QxaJPqNy1hgDehRafsTg5EyJNsoHrkpV9j
ZhtoC/yK8nC/z4oEGz74XZD2vJ1I92NKJVwjfLlZCtFYaErfl57jl+1YPmqcnYNld9jFb2T9sNbj
HEvor8E0WPBd1YRhujZtgCHtt1nfb4GOwBog1KOMCLO4OZ3cXs2y8SrFLwjDIZTJWeQapmfh1djx
JFV/lV4uoq1+5goNcxUlJ8krBJWQAXwMnh6TWVzBHdNGR10/FD/tQ4Kv2MhF9q6JaK5EQb0+nwy5
7xfrGnZ0pVT0X/DmEVx+hXPUz0u91rSFCOW8CfZ62vBm6Ql3gm1o9U69TEov7X2bSd2sUpFCqJgp
OkJEpgi0nmyym0LfKP2DamK2+GLVrL9vmvSb2joJg2nOvCHWRqiAZkJL7aayFeNcKkhImtRjVKcs
UjBHtEMdokifJQ0HIYrc/lb+d7Ic8WGqYb3dIoVYVgAczThrqTo2Xq5HeWfbJZi8NF7vvQkm+24l
0xzfMmG4wq5eNQn98tZfpv73crH4XRglxWOCOkim8t1wMIv+latPTbeSxErrW+Z+LRFQl/HeK3bC
/DLiMGGYRdit6h9qL4f1seD3Zj2k9HYqHWY/KtIjgGEK590bHs1+ks8fsbMpZAh3tXfE/HjdwLax
FX8O3VsbzVIP9ECPxezsfe24Mj4fu4qeeZ189enmezUrYEuJ7U3GlJo9juHLXbBRoeWNdaNPhSD3
9XfgRq150yPYBEoyTNA2BtIQ/diZDZPpyTNc/mvAiX6c19xbKO+mcGSGUSRxE7oOOLTILqrvxk3f
77sRnZ/8aM8aT5rKillnuHVhdHrn3KEwdddlSdcwH0h720HKG8k6/TQmv9iqCGXTWjDSVZjbIdqc
06CNkqJ5tH8Gbo2q/brK/XJ3qWULxxgsbp/KZlae996BSdabAnm9m06eulFz0IWSz5KYfYQXkIwy
pMKHg0SrtOr6sr/az307Kpt7hvKtX1CcOavVb2cYLqz0C+OkT+xAzyHE6B90WohO+OIZWSEHHxlX
1cLXp3ymKHOX7USaY0i9JI0HShbpgjkitdE1cWjUokGx405pg6sjWndNGdJ7tb6nB5TDR79IAIsx
9DnKblMOPCyioKYImB0OovNewMkfbazasjKvLHkS5zgujnOtNKC46n03kidAAgWfvtu+TPhBuHtu
fJIMhCjEypHud7r9pQ5cO6zUljFQGdQ4ilzuw9F/X+Qd+o8J5KJFq1DvEhCL/QaETiIg1Eh1xBYK
n7DlL2qHtAJzcGP2cWq/iS8JE4tYqidhQDs9DvyQdXBBRYTZPJjtz3bsDqxix3BmjPrJtW6smDxG
UgoggDHcJyCVSxnXAbp9SxLktO6/iwamje2wJDV9GTFFUM9TAgwJ3PEnsM3FeWO5J0FVHVRiZvhy
xSaeLkT8diU4b4jlBkxtdnMEbocSJ0W+PruwuZwHsvkZdL7715+1guO2sjWhronPoaIPH4sJkhct
yIUUhS/Ko0jbYY6ctMM+KmDPl8AHZvaX0NrDHR3RWT1WWFI9GYNTAZtbQHkEnzzaFzdERQCHy+g7
4en53+G3zRTJXBovNVabJekWqw2Hhnj4jI7X2pJAdB5NFUb/zj6T84xpQyGbiAqJAkCCTcLDZC1L
MiMn2xyo7pwFeFmKK6DQowigFPhcxzNGL62YNLGm3npIrVp1KxeRzrGiLR6hf89fEYMd8DWSP+Lg
aZbYFVQmWnK5Xm3caPpSIBVSr6bxuDcb8ZBd2vx9CJ0sqFyJovA+yxG/YhKSDl5j15e5uxF4TyRM
5idBazDjnVqd8SM6JSIjsNa5tic9DGOKPxbTmXcVabV734onKUz/dnAZ4J2DR62qiLRaxxOTjJsb
HLuuJYH47ULKkhwU8CwHooVsqu90vioViALWoYUNouHLhoC8gOP62o/u9XLgexcv9LkK7QTeGW95
wWGnnAFxr++53DEsLqL0CjxFDuQrpNbubElMWtUNMZmISEV7k3hims+etUNJAn8dr5JLv6S0O0zP
8+5VToF/Opof7CuJ4Q/1PPMinsMOVKnrMdxmyGbxknZJTibPCAA3NLCy9cj+ScRpbB+ttGjfSE0X
ucGn68HYRVgDBOGKxaopfvXhYqU3r1fvXBQleKean1blIFJ1ROFjCU1UvTCtlzaXJO9IrDZolc9/
mtEgpLVjRjprZWjSRGrUNCC0DlbIQ+hRa1GVIOZQh5AZfYy4GDBUob+bf3N5W+C/3zL6ytsuKJCt
PGSzUzJuxj+POH1tGvyvrOz/aoe3kdlQZM3vkQjGvDq/pGKsKYrx0Ux47GE6vFxIvZGkEGDEjrsA
JZ9jnvTrFirJJsWlId0XC1t77iPzI8ElPthKVFgM5tGYLuspIxibhve9zqM6aMe48hJ8mU17FK6S
QFy90u+x4uAGz1M5QcfTsLaD/NDA4EjxiHJTYxo3hW9HnHPWv6U+4aroazCCFO0gnmyEvSfGdVDa
xyIhmFhG19VycaYiYVvlLk4/anL6hDxpksQLfmQQ9xj3sqeRoSducedOewugNZx0O/o6ruIS13Gb
uNG05YOm+CC878WjFkQTMYNBli8upFPBC9KVwjSNejQA04nacRTPYJLUm/NeMjJwVonxaP9hXjgl
XbdY4c3UACAqvUNI0/l/C9GfWZp45n3UjHq33LBtB9sJxaxIrkDeS9Mn0jsuUjxN0KFncvTbTO5I
Rk7ZsO2q/HgSFDD0oWuZld89emLKd3JHED7QD2zCHlQe2+2FLuEuUo46NP19IwzbkvlwNrwGuOgY
5r396QYenfHCHKSoH6YjTchRknLf4vwGNX0AzhDaDx77WBaoI4RUg9BExGl2+UQum396k/9jXZ0u
0NqACuihlbUbMLFRGYCyHt3OiK4y489SNXbhCBf/2lhFx+immZAE3RNpIbo9eEwZU8LWchGfViKs
0ZfB0BOxQ9RQHcGfy50+DalOTACYQJ/15IMf3N0wO8vsAifwQ9A0H/Gym4aYxkMhSXN7WJrd5w15
wGB4mDNl+y3WdJVxUVwZbLMWgQGu8UsUG2JQaxaj3QRJ8cISnJWJhH3Sb0kZvE5+c7Fhfo7P3dld
gWqtDW/SDd/E8LbqiYHOrCTahghlepUwDOnJ5E6+XOi+KjL8jN2TjWXbV6kaR5xjlhRlSp7iDodi
70i4kIA1xClzvW35KpfIkOmteiKIh+VzUnvKwwR7UIScHlZbP4DTXYUD/J/BcJ7SZP7o/HZZXixW
GcnwtMKne3VhfDBdHmivKSLDY50T71jeMDKuBulchaHFrahyjumyOMoVeYrXYwjbrhNFC4ynuTeI
rPEgfy10gwYjaXb8LrHHCoeUc1sBK4/TOpV87KyWcqOYQYWUvnV4NYaFt4Tqbjypt8J18BmQYCuO
/jDvgeo/6JVnO8xwB65aGbqGFaERXB8qmRK/7KODKoAKYcimx2k21JN92CMiaG4YVMgDasmPDU8N
oGPUs14JY98Vh8qnN3LWcclmhDZvCr3Wlb1wo9Vd+pzNV7XH2DsWXJAq6MCUwb7nZ2waFRo3swrV
gMfzrAvkq+WZcuqWXC6wo8dMRnWglo53aIP8TS/LZDUJRHHOQooCTxVEwhKmLvYR1nW44rJ7a0kq
+R47YBPCr0VFuzM+1+NGGyoKDjKtD8szjpaz9S0ReAQBgLAeVV8nmMTlom2KcDr5Ko/sgbwIn3SK
urTbBQTfm6l3nh21BWIN8Lky1W84xXa64cQyMCOlyuPJMKtDYkfm7IahVhAQIt22L0U7pkEmWmRw
X1NU26Y2SQjUAzpo4MQmxCeBJzmbJqy7y6iSqWszy/865jgPHP6F9uGNhOQbX1ximZ23X17b4Xe5
UMPOCez8a7w0bmOj1SK8P8FrLp4H4GMUuIv9RrCttTJPX5ERZ5T4FkhsG+iBORuqTujFkcphOAlh
JqpV7A4aoyBjelyL8Kf6CFDEr91yNLIE5BI4WNEN0mFXS9DPxjUmj2sM/RE6xkCgC7PaXE68KNYi
35TOzf9Zj9rmaSX9Z98i2z25VA8sCxMm698dBq6kiYd5YqrLnZ6xm+qFVf0y0anmIsmTK5OIiHNv
bMjxjdUPRCrf0X+rxDsYRHQA5awU0ds3Ajm87e5RjUDzFp0/KsL4dZvFjVvyN63g6Pa4dW+Nkw6d
f4TPiCEUGEgX7tNbXcoVWdq1fAwdGv6aBpzD09RqtSKgQglEV6IuMdjEH7Br3H96FewZCph3RUTX
HaCWAkNIy2ZMpJKzu0ePfhIX6NveGTSCM50baoIIW5tsAhCsmO2geOL+Tx69ZV8EUvU+O2SCsalN
vkH7BvyTefqWkUWFfj/UKlODvXGsZQ15qhEZRwvve+qgB7Z1UeJMc1Mr3JpP9ZQKj5HHE7Aeb0BL
cd2jZFZFUQ6AfoDuyKl252pM9CIJiQAhccT7zWBbSY5lBSI4yeh0vU7379LSAom3RXhekx9Zlq6L
B42XXHsZExSj+JOcTSCSUhn7bKigZSTg6/aeeN1yORX5kl2Rw8S7HDSEF4GOKDYCGgaoIS+Z+S/4
tyUOpvIzcfUSyS0IXpefd9M0J1wdcbZ/Fajkap72dag0ZlQCQHeyYtmel28wuJ42OnoSP/e8KESD
KrUDeV8J6mtSMGQN9X9392DYs3vMWxVztBDT7FkdTBBLUXjTnopZ1cL9xWy47OQixoOlvFVakk5n
NLfNjntqxn2WTW1eb+fmcXE8vsyFasB4nIRN1DkrrSM8btbVGc4EfFoQWKm0YnvG9Jbin6sVYr0Q
GKgCsMihR3zzrbUzDRLv3w7isF0DsKowwuLvwLNEnHuiWTUz0sR39CGFt0LG7c7tyyT8ulqOWVZk
+FwexOADFVbFWspKNEYA65erCifaONjFzTKRGzoiDGVaCTKjLueN2VC7dDSqr1FgUPoH+64xkp7H
qpl3H4PJ8uxzofbmNWKfsCoxk3qWDlJTyuA7zaakQoVNhrAMhpoBYULEB3ZZvnUBfKXm7n7kva7D
SLEzkHAOfsPhjxKp8mcXGpIoTaVL4zLw1I8l1Lg21nvqDq/ovD8FXcU2B0gT9aad9hOiF5nF8yiV
uXoSJQkszCrse6fAAurcBAroGVA/qz6nsRjrhXijQxgen0/lXbk3l4R54goyWqw4mhTf/Ll3tD6K
wKkfjPgJ5ruIDj8fqGr1+lFrLVUSg2LOJkPXAeMx+HH50jH0jgtby4ao+yz8zLvUYiVnJAv7qTRS
kFCqBOSdVsujI/IIviB2WJvJnVC13zQU5dvHNh8oD0z9aFbkfnM63hy+hBkV3V8SGdZ+vnt+SxIy
lnZ3p4cfwxVn9Rr0jVogxnl0bMHws9CzRS3wGMZeBIeMxWiIHt+YY/2SIThpkLKIkneMiZonua8R
T3XpxfurG/SCC8JHeOTa5c4HU84DBtKCjpwYjQUfZNDeGdTE+5tXFgCkgoGVVkdbBHf5oO2l6+SN
5++4whk8h5shmpEQyjCV4FND1/PTDv+DmZhMJKuLbHx3ynBiYFpy+IspYTZcDSFGxPfKlWCEh2Qd
L3PKpJDuj77dXpn7m3VldP3hSloNMrQaqgexCNCX8xtBGr3slCctYoYx199gMKF8UPjqezUAdSCr
ufp3IKpyqMV0RgBqDqlhuo84XIAvwEH9lo2hoju5dxgihc36cHLRlgJS3q8iUfGWDZdPmsPm4rmG
HtqlLzKqAL/tF7yvpd2lvF7AtI85E+rwsPssdOAgI9PVMaEkh4EmszBfp0OlIXoHBM5N0B93tyuF
Fgrn/Ycr6P13n9Y5kwDR9E3c2ZNX2HzQMUKT0fOo37KbapSslHKTUhsFTopu269yfmNFJHHeKQ7X
mM0VZIoSFB0F1qqnVO+c26tsUV+bQtuEWlRDdBYe1ND6BtiLZ6BE7nGk3hbTYIDG7nGguazvBGrd
aJLTYD3hKmzT7J2gb/0ukxYYNjZix7Z53C5XQV5uap9rJEAsHbT/2l3ZUD+evMPn7GtyuBTHkNeZ
QR1eDee7JxK9DuYNHFa64U8d6zknRiF4CK/vIa9kUbgS+22Fgx0v+qDPg170J5ASa4y2zlJHMvZD
dtHvA6Tz6EnxTTcdc9AJ3zXummzRKRMlCy+OHA2c/vdernq0YJdevKTP5zi4KX1z6uwJjXmhRhwX
lnc6pxV0H1qfT0HI44xh9gB06PCY9AmG8kthVV66ojAYYLiXbjYKMjC6/3WNWJOC5/87DrLt2bQn
tSseoUfJXXZA2FYsqyDz9DlkaWi9qWNdo+EOixTPkkq5HFJnyrjbZNJLirceYnscj4sm08gotAui
wYLhNPNdKLVQQxoZwajOGNgXlQToYr4/pDTaCHLFPtzs2ZQ5ztpmGUbYoQ30xp3+peN9nLX0+bu9
GqmwAz2PQ7tcY2hzz0zXoc9sI5WGeX9lCGWvIsgZ2eq8MuWFNwgkxJ8L4ZPf0GD0qLkNBnRYehPO
R7ihBS3FYhsQCWqWTnLEEGZvDoxn21D3Grih7zid/pXjEilYzYNCSuCHxQxuZvsVBNqj1Qus+Diq
SJivLQQdmCEITk3wQqLdKpkFgMYtKPTXpfs2/0wYM8pCRKqUYhza+bnzwBJQqkk655wE0HdqGV7w
d9JStmLSK7+BseClvmaI/n4xgHunVzeTvL2JUzZoVEl4DmGNnLuL5pYIpmj6oxERqBeffkwM0jnE
4ngQqhhmZ6E2pEq0JRkBEDQ9p0IGAPwR6b93ACV2Qp6ASCHD89fG2PLNZvCaeGzx3m6V/oUh70V2
fxA6bN7GK90yGfy4O4glgykgK+ymfrRp358q6bJ6HTpn0pAmHD9SAYEPq8q5EMhaRS1kWN1MS85k
tH11F0qfyfrfpviDvru32hmmnj5vX/t0Pzq0RTjgTVY9CuxWd2zyYvebHr8hmJyZoYwF4/mSvR1n
mea/9qQm4n0+e38aldePiuYWhXcanhnC/Ni3Qale6o4TE1p4OzEhGzMv0i1Mq43xnpTfaLUAstq3
ZauKjwme697tep+SNEpwTzTVNHo7ulBEOSS0KiDYLc6ypJuImSmbwG1nkl3xPQ4xupCFSLYD4PUK
57j+fVx2BtRqpIXQQrIEISaOCoxq4Eji8kmoJVMc/pJ7cOcXW9HkmsvBYYkn9uOXdvFwFU1mamxA
aZVWI0VaLa9LBzr6b5S6i2YKxin+Beb6POopv+knnMYRrxkg5Jo1MQftFzAdBJ4nC5cGSVvWvRGh
OTslTm19VK9JZrt5O0RcX09gxTC59c/6jeihbBysMeu+qZ2NCpKCY0Jt2y2vLCsfa1yEaqY+1KXC
8JT2L1Y6aY5/wgLzOfvWw36DQIOqhlr+U4Dk7yTN6vBLM/4aNKwY6MxC3iYKLnUDuOkDKtrpR4vS
SZdC8Of/m4GTTLkaoXEArXjIlyuYYuTweFuri4T3q/PwiGiCnRCZz00CUDGm4DjtpyNaVL+FRP6I
P6yqXvOJ7vCgdK0QPe0dhbBSCnOdgj5LerkV7820zguzHJh2GqTNZMFRVjgpk2yu48LyPUqODjTc
XGgl5/1IaHKWtIh9bqe5cFPCNFSQMYCKGc3Cz6y/KvDWYmei7ONnOAfJeX3Y1I47JiMrK6J3mmLZ
OYCU2CkAMD/OT6wV6SgLLWu6AOimvBiPQG1Y/Pj75qEucUj7jweGKFI7O49vwsNizOauyGdieipB
Tn8+AZ1GHrL2XppcrlmI6kI0e6BU7ix45cfSk/aIakmHpMF57MGdUi6ZsQFO1+xY8T3hUASpJ2Om
9dLYqtkowZk3kt/paZKsqFjN0uZAS2uNiU1I7u/Gc/e70QYsBmyoMDX6q1ykA3/K8ARrQL5F0sJb
gViIvFZ1xioqUXJM+tbya+OLZ0Jp12v6JoNMDXYe0XsgzWUsult2fsxuAV0wMHKp0sDgAxUVY5l3
quKkc7oSMAlzrjUK/GB9nVBQde5eLdZzT3Ax5lrkEw4Dps6SqqnMC7KgDuU8+Hniqym7Dy0x3KFN
ziA2KwVIZlYP6CJbFKvu9uAjHgUjMUo66pDXvJyiaHnCt0XCf9qT4aV/QELVhPByaLOVyz+mgkfP
wK1J17meo43WIG1nozZS7wiPuLrQOlcuGnd+QRBtKZcbZ1uqJObGqJf9ZnMyl2cQxZ0y833xP+DA
vY18DgrgwRhacaCJVq/6Pe//4B+H0o/RGA8UXEE9vixPUDzhXyXCa0EBDDd3kAv0VVQXWagSgIjH
tjrDjFFzV7CtMqSf7kBlJDRKoL4MMxE+mTaTs+i6ltHc3JnAfsuydht1IkqWtr7ZTtWsaJF6jq8v
fiu7Cj3ciLXVZbrA46L6cygrlL5qYXpjqy6TLQMLigvpvFcbfbq7emhcITOxEP1e0u1GQyXuuOos
jn0PyfJIwgZDkryTyuuKqo+23cODSfGIecg+RYorgKOVWuK8Rz6p6YBUyOUvDJJxeFz5IASLZ6+C
hTCcv08F9YGePeLJddDi9CqrJDgbzwp4xFNv6IZLONIaOAx7+/BrhJboBnNaaT60SXAu2/rbmrWM
fYA21eQ8h8T1u4iqbG/9KS3wIIfKeNudbFhACXWZxyMt69eQ/qjxQS+F1WopyBGgy/0IUMuH6Jt2
RoUm5jdUk6Y/KXJakcgIEB86Bul4NlgitIdBbdO0fInbC4tZsLRDp/oOTmwK7+D4hKQLTdhB73w1
dNiECYCrIagfMN0Wq6kH9fFfkWemFj39YrCZv64s4rQXn4J38zYv6crMPvU+32Bghu0NNqf45IF/
3nyxJGdH+OIKF+ib+YiaCdHWHzRALocOHm9IkGj/BsIDqvXa6hyyTQyij6T9gom6fLJwK+NHfjPM
oiElLFN7kpW4t5RUG8QCCuSqyrqZBYPDU3j20H7b3p/yZ3TTOBg6bYB+kgMKMT5UmJ5XQyDxX7eU
govf7z2ZMZl0dVOUBDAk6c76pUAHoumSr9PxGFoYnpplHE8ZwUUuIw8EtKld45xZAa+MMsuibdqz
VcS75R3Sc7CGvd93T8MRTF4p4O2xVnQrog4Yh3+5vWLX7LGuX1GKYyyuJ73XjFvPNiCTkyeHps3t
xxakQRpDmkYti3mEbAGWbbjgRAtHzxjb6nqhizwOjvdpuUYOFpEHOtE1U97pQaqyLH2v126mTvYa
97d+skwkQ1eR02DzR9dvaU21J5dnP4VoYBIa/Dx4G3wyQgjDbWzUEirHxRIfUIDusryFnBjmzyFO
Ca1d1OjdWdyDQz0KcUdp2x+cIptaRx56JzQggJpzvE8XrNh2L3dLwLtrYcPmr4j2kZCEB/nzlbcy
JTN8zXwaL3u3MGaO13i8D71DxCMMs+/KSXroXI4GIFTOZv8lucBnbupPEq/k3TXZIxcAJiVcotHV
6D+tWGwhZFxiWopHgowX9uH0BL66PcgoEpGt1dBftHYDtHtop2Gh64hKfwxZdIagdqgPowkCUdDj
27LcUb5JgAeca0Ju9P7CYGKJ0qGyhYO+6qzELOVFHsvLvuOzrcq84b0zXbmKYgN4tGNTvwbIu9l0
64DWANtQf5qA8XXS97PlViL4ctpZO1eZVYASb1/UR56KG/XEJ+YXXnMxEHDphud/N9tVp1WMGCdc
t5tZeVBPIhlWDs6kW5u/qTMr+0oQE+0mt9lPLDQx3Gmtze0rzmNaF7hk+XkZxJhH4bwpLOB4cV+v
6AlQHuzk6X5r0zVi9BZPGCScNgZHtSfMfRnSgDl+5AvLFun+mnNHdWcsJ0WSl+bR9ARj9PFtMZKQ
FCA9p3xdXaNYJ3/+LjHGqddKCcovL2VK+NpYfDYfEqyXOMpD8vxeId1mgtwrMfHQH3vk/Pp271H9
a0Ea9RQw6+qCnAK2MxzZ+hY13O/KCJ1iWi/MuHd+o/anhUk1CYx+9GtoTf9QIkPj3OAyMU7/ochM
XNG1WcqDC9RQUlHHG2BKZ8Luq7aIkL7nIMwnuUoEZUo0AEmR4bGnRXZ9cNBkUJCeRwdYTgSqES/u
0iP5ypBwUa/bk2TwVF3uPew+YyPxaEnBsY/PtX2IwOenwLLYPv2FIw0x/a7qhVb9Sx6JsO7VEDma
3YU6Pur6h5gW+SbwH0DiQvKHD9WWhHr4gc/Mj7dd9pYxrtUjz57I/EXe+ofhaK5pcTAzTkH27lK8
4NogoDBd1iZMGWDDJjEZ1Euk9LOYZY9PZHd7imjBjgx/oIum5shGYbF26fDEjlHyYRtEvQm/5wF5
NgcBchA2h/5E90kSRrnwVCTlbDKIG0TAx0jJJWaXa6GEKwVdOmdzSCuEL9iutLQj1gx/svae81zx
V2CI/KrMOwQ55JF4m7PksAahIX+rZMW+sA3ikXJLrXzDlLEqGrVmIerbB3XRAUmsMbpmnZAAV3El
dz/1kjLRnOoNNj49l2RBz21bBklpXLFfHsy846y1xZaWIWHtS2xATI7imK0mIKwiAI35PliLWKL6
UH3L+nHrYyBlHgS2bNT89clUAww721hArrBW4mSmxxNdMhW32UGUsV3ytDA3mE7u/NqYZPAakv8O
hcamJVGEMBMOQfrf/YJkh1u/fsnxpIxWvfyVIO22XaRYQrLGuFOVEG/sMxK89k9LB0bHS8z45m+R
QlwlJdqJISCkh4A+ZC3anIfuqL0XRAwY+VsRnyDW1u0ezc0VBOsV0OQ3XTwzAfjDZVqy6mVQoDrg
4hDlgJE/Y1vlKbk7q1ZQ4DvI6fqVBWKy4ED6RNiIRZHcweMpYBikB3Du3CfwSGUG7HIRN4GvWhC1
Ezo9Xba5sKwArMBmisQszqFc59A6l0rRVcsap5L8e0/WfxMJnEL/+YTRyR5uOZ/40AXh/7m3/7+F
Y0LYmmyWStRq6DpT8edBLjSxpb6xdIfv845kgKmZI5GVbBhbBEI2yEw29gE2Mva5By5vgSrG+C2p
ZuvPHjdmCYdy5Nuh4qf3uv8j4WVDFYp6hi6bIXwGf/vzgc7K1SdWM0zgx67zRgru8elhIPcKw2dG
yqzuL7ESu75H+X+v9dcW2h1o1RRoS1mBH1n2wiDw87lL++A0gqAaqN8dOF5jeLlZ4nsrnEKnIF0U
SrOfHIjsMrjTL+fEN3cGT4YAh9TgTPQMdTQPPhLzuUNBlXFtsWr0q/9hrSbJNhGs+VaJqeYJ7Ow+
7NRR4mAGJqtd27DZwTOYnOnXJTOjBVco5nq5Ma4H2cpH9eMLg1d9fjNnpEW2mKSqqSOktf2+J0Ab
RnR2hbnzAJ4g42Ka7s4gCp8yGFf4Uzk0xxW2oa+Mbx0rqh1baiy3MWR+X5+DXxP00mUgqo5NENUg
dExOTXqrMTECcfAzky4av18ZXHm7UZCEYY7LnxVI6DrKAmEKv+TSVH94m3kQaO/pucUzHyT0tE3G
uf8HQ4o6I5l9pzpgQUiuVpxxvYVuwpv2kAC5om/hBtK6Pi1AkqWv85CP7txB1E5e2RS9tNdh08i9
ONN7bjAjAO95iT/czc9yjxa+LWf6yX1iLSg9pHY7q8KPghaejE0Bh4qbHsjBIK/6DD0a4miiMbLB
gs+wdmkRyT5mj1GwgDHa3HczSufy8gotC0Naati+aeyvPQHBTpIsbpB5TdRAoLAn1mm3JCaNjTLt
uWprNCdpMTnwa+lYmmqYib2JgwNa7ks5wiA4RT7WVhoMeOqEls6EK4n3TQMHVeKwxQUWsCEjuyHd
91K+eOpQZHbUMK+5JmXDD5gdawopm9R7QJpHss5iKd3KZxRvGSlhF+8TQQdVJ5aMxLHT6NAIctXF
dwJ6tjZp2NLXvrspiiRVEACcSfgmK8i6mWSuRaqe4Cx8+v3/hJT5ByqNvaIj1cORanP2su/i/ZP3
aHZXJD1nLc555Y3XUnB31h1rK6ezrzgjEIESAqhek7wzY4BCBchk4JVMI3MqK/oiVoJz89y3L4Ek
uVl0sQXxmEQ2gpix/ewpCKhO+E+BejUN7cplGD3obJqFbXn4PhEbTmIuzsTgGPCv/cxjqXPkI8fZ
evFBj1kkCsKpT6KmMYr+vXgWW5UoEtJBmYoGCwLMH0eL3unJiE/6zUoUVGPjkWUveX0SIVRCOldu
0Mnke0i2igXDCQ7RlRd9pxvkd4p1VMDDRrHN+tDiNKOvfCetHGRaYz9Pn3kWDmCgtlJ7tgdP05b+
ULpT1VK94d6sCO5dVEfbsTbbbtXyvUqghu3Z/EANZG3DUy5dsc2Vr3lktm/p3cIuo9Mb4UV46wU/
6f7ciTNzd0+8DnjwMW8jQWibxvOmi8ddQhHJ00VhdmYNF2p7kLDwBsP/ncshQmdIDmcMHwHLpWS1
cnmR5Bn2eiwm0IIAx8Mt5zkjO1hDGz3A38T8ijRVGhMzu1y7TWuJR1ViJpgMOEudgNQRQvlmLQRi
jMIb0vRKtG5NlambFtrwXP2MIZTHiouteOkZA+blN79YLp+GsiwwR0ihj7XX0YUQCucT1z4H/IXl
aQl3TQN3EMxgUeOlWHYnRptzoOiY8wsr3Vq7kH/K4c9+xgiH2W5V29UxhI3LZ/xZ7Obnd3dWj+7C
OXSNlM3BHfNgNnvC5+X+jNZA3GygiqKbaTFpw0cJK1/pfZrbu5Fs8HlG1DYxBO+9IBpB/EfYztr0
+xwPJqubKwP5aIuaZENSYqYONCCwlPmn8r+Rx0ekxEYQfLIWlEnDQOSP9MwN515M+oXv/ByjyiWE
aWONpppzhjSmXA0/T3rvEBWnLE+R01NEzlelx1xcKv/pMQHmjZ5MIHsRS6LrQ6H3pkwF8/jksCoP
/ZiGCFX4GKybtRlkCW+4WFoJiLXDMXwdxFugPsHHAaOrzg7zeeLcWdLYUZdVAE1KbFmiTTLqa8ZU
4OOf+sAaAO9Ga7UuLYQ79SWsbWCppwWh7r3BK1AJVwQSfHKs8xLrp88+ju6qsUFVMuDPNkULRiiC
d/I1H8den9wZen+LjWVZnVCwSlcD72ok4Eu/5ztxLDkb+/HOYKxa4Qskabpkt/Wn4ZE/DEQ9JnPf
kOfX3cvlvva/ZQyTvSHdJ4l/z8iy0w0HBGL1CC6T2CP+kTQF7OjggfpdMmUFqOXfTLsCJSl07jHt
kvw32sx8TapbPS5e2DtdY8e+T4hyAO+6RTW7yqesdiivWo2ViEUQRYcJPLWPFnwzyEBHvkHi3c7+
lZBwN3WW4xI3YM59jh7PNOvSw+vM19+sMwl82iYodv78P6boSTJR3zHeFDDjjfDc//l2QBrKPGMj
/qaMQZIaIBZkch2aUu84bNuZkAAoUvDDWgcTz0oViwwK6Wt5Qd78UG3YnoHVUX5oi+vH/JxI/GhC
shFs9mm4UH+iZ37DZ6Dlz6i+OHkPV9RTv2RldXj9mEVCj+f6GwbaWpQEMD2/Tk5hUDQYZS6agfUf
hO99W3Wh/DRvwcZQlfC5aQRYQAkPdVyXdtTTZSDwvbgTloRv1NhgQSHsCBCOA9wXnn8Shiu37E7X
8pwqT+zP6DQQxWTXkCqESuN3UmBAi5iC1TLJT/SSgzHxaJ3pTm49fnpaO6b49Z5hXPiBF9N8vRxH
ShptPj5ELqa+2EPdKmPQYYsPbUqgLBKaY/pxtC6WPRcTwAtVhVinCkeTMyNt82/vOcjRPiwJUPEv
lkfkuPo68py6tkf+ib4M986g03eiJcBfvXACc1cWypRu/+OJST6DF+ZcOJtlEBU1YsLWMPw0opVh
VvK9soty8J/uXDWcnl8HC2Cm6ASZboLXAzS/v32XftYG4xJrRLtmG/dqt5zcqR18i70/7OqMhtlv
4QkIouKiRWSx/BiWS0R1OvUvH20rx7DfS461Dr+qeT/buquqesy60b9Sg9TP+/rKzP0wrn087Bus
T9EWy8SJoxrwpByVdkkUI+5VDtlHxZXxj4p9hXkWSsomPYimbfWrAbznI1uvlg2bgbrDXDXaz2QR
dQSGgk0QkI4kolZ0ca8YVcEO7GTAmscmOoNcCh225rSQRbt4nyeK5GSpuvciFf20Jm+m7CxCug/g
2tir1HvNGG/rwINkWl2QoiKLZ+vzBKVLKFmcU9hQ8eSRZZ4ORsNTMmrtzVtwSo4WXAlcsWApycUV
SKPHaOTPuUfrG9lr0mphcWgqLVtqyq+UTXi8rRP7LSzVU6x5UoAHRZvYWtRuzhlVuPIm0oNykQLF
cI6rHrxpkpMyY7vz3g332YnkI3UuXVJH+ljTUG86aNUMFZxkTpsJAhhgzk8i5NM/Fj92z+sdb2VX
rBmyPtHAePH6OCfCGhhVATKSrmbxPS8kgVwas3TPZSzExB8lD+dl9+U/+DGPHbRPz9Tb+WPKUbbn
CynwqezMeFdQgPelLwArKlDLdHl2bay6MwwijrwVvqgwl1Wm1Y409zm/ABhpDTu3q4V9+mIvQqMs
vZ7sK3Z+3h1Ew7V5SA0bujEYQB0aZsIJItNe3Fag6F/sD4ZOj28iTFXUvzHM2vh2N72pZcjrWTXR
ox+WcBsFkuDWMIEGMIV0TLYf8NG1kT+0ZovKzccp9LaP2V6mAwVipwbsQSV6X8b/Wm5cHvOrLEO9
fvdMe27BpbdsEBSQGPRrGSWblzGObHOOMA4TJCeHlEH8AXNPDdm18LiqVUGLtVHWCZFJLkJq5fBQ
1tCkdaiKyyV6ZPb03n5t9uEhEWkpf4Mu1+wiusxs3Ru0KsdOse7B29VPAoxMuYvZz+mu/up+LLSN
g4icTU35/sNLbQdtyY9V0KsC9RHH8XIPDpUE2eFAzSgE+YPUZ4wtFADZE/egBWrzOgJZYGHHyRMN
b0MPA5FRYyjwoQyc23f1noYIGMXxEJ+0PUpquUiDrMcK/Wt+W+p61zbw3eTnudoEX43iNNu3+5Bs
TsL0EJe5dS+i6LlDGui2uznvfuCApIbk2pwd6w0fT5K+Cgo3uE5Scsf/YB3ycjLQDmIzq0HQWOTv
53fORnBwiRr4GaGgKJJcFkS4EsfHzPNpWxXPWHRzsy3m50Kyy1OZeRt9w8Ut3DGfw6Q+r2KlnZ4o
Ph9d9wKfw0jXEfmW6oL2v/g19cFp78CCfI9aEiALShmNrmxC5k3ihTMgFX0xraCITp8e5qx69Hzo
nKdiNwYD6xn+Vv+Es6Mod2OgwtKz9zsB4VDp9dm8BR+qWcCaFOgAdFITDPC1wyA90Zw99wd2j6K7
NHUC+TNsEUF66QOqV5y+9Ysrw9HY2MIoO+CcFmXHqtMiViX1lKOHl+hPJwv5VjevDaV2npt4IFLO
r89cPtCNoovwdkC4P8iGrsDJAPB+dQXwqPDFNx7lz57EJK2u/sYPVG1gEFQuUmrG9VdQM+s1WK7w
y9QnYtjJ5vM/dj9BXhIwYUYVFuljrM8NqgY410g7Rrkzye3vGVnSAgigDuJP+Mwiu9Qn362rcQuo
/pgkpknzwYH29jQh7D0tfP3oLmTI25NJKa6obBa1pFVmIVA0tLsJgfJFaHlIyw6lgEpSAds7mYhV
mXLz0JutrOysEBar+V0pXC6xkGzHx7MA6fg7LjQlPyIlBCYzTgbdncwUoWb5eDFCd+k2SF1KOpQt
KnRNp7a7vNQwwuhogvn2iOm8LTVU5/iy3kS1lkDEOEkekdE0LM6itzvQug16WaqnZ1CQnKzgK6Ow
M9JehGrRJ3dVl1geLoGBivmB/b5AigxYOJT+ICp3zrjDlGOGSosDultaNMmWPn2eneNcjOomVaa6
LPUBtD0w4XvsCphXuHUHqh4On74tITRqCcUVIHgN2xVX/t5Mixvc+enbcg5MKiAQTATIxQWtwWu1
uOfaUjO2v19t7/Zunqvpfd4NfdQVB0qEXU6He5M44cEtfPg7HG8n8oT6X2AikzxRm1V9Vr6ZTvDg
Fz297FXHid3khiyc1kl0TIMJAUsJcligGg9OYPS8wqcaeabOYNzt0UK+PJakVqA9/56jVrxAZkQT
O8L+zjag8nBiCo4M6bv2EBA8El3oXSXviMxppHrqaQent2N0LpWvwaWFqmEwG0IZNHdwWqb+yBBJ
nOKhU20rJz5IKI5UUXSxOT8yexYoN5wiExkguBBeSML9AAX+GquFqXkk6xZWm0xmygqPpMl6B+eD
/olHUSWg3Y8LBEFFUsFRLc7NZzcVRkWGlESJly/6Q+/Uats600hoGSY6hT9VbJu4/iPcNjk9j7k+
mmF4iLDQ4pRO9gQc9EKANMNYTHcwjUKDtyBN/Thw3UUVz7rlQYSU7In0MfWJVuzaUDwa60mRBfkN
NTKQgx+8gbzXFGz4jUjjCI4rmG0nbpeMfQOAM39TyRAd8I8lB5s6PWf+/47BFWWIrrtEewJmlfaD
g/fT/WEJcWs0Fgbk/35ovb0jFKFn2nHPMR/YRMM4rKZEnwWUSa04q97YTiS5N8v7bnqxEGgpFZb+
wH94GkXgVHpmog22TbCFF8D+a+nnctwIdjCWIZw/v+Z3gYDzpcCpgWsRkKvXXuEtNtgbZ+SFOVPW
33duHawLKmQPsmZ4WLZkNpNFpdVxY9b8KAI45KVAUrzAWXZg9m7evI2dGMDYHHDkDo2j3UQ+SdgU
gPIKXoN7DzbjVQRYmaG5z6fLPAZdwDbw2X/Yyun4VIF65PhpGKtTMeXJ5QFYHqZ6ZfB/5DOVihWb
gK+0YcQF59JpZXQofxPre5opMyZs7EYmiYQdTtozaHvh1DWqAsaSMIWPAxJnaQ55kId7fA0y7xjS
TfJUjhGUTQkVj7AAl2LhhhRAMLumNbud/Z09Gf8iOzdgMfF3IIZnclN3IXTSqt3i6a5Au/FPYBcz
mdINh8rKh1rO235cRsBJeUCfmvHUFmzNRPxyovc0+g6AiDJSrgPVUWdcgSfzZRiON+X8bqOkXKab
xPUZhoOXdrpsKTZkjcB0zzHvr67O3tTWRhHeNhEIIixk7o1IOzboens8oO4bvVHQn6h1cgv+JJGE
2IPlgMbOARu1HlvQWna2ApJF316hMU2mt69ULTV1E6JtK4Lz9Nuys6pUAShHstS/zoVyMea28ld/
nV9AbecftkBlv/HCACNE2zvv/O+/zg08qppupTtGBqgfUq9XjqYt3mj6VfUxDIL+wE+kmRkXoGgU
B8MTT8uNrM6FpH/bhOccqTK+gWOMMdGcxOn/7lXgjo1GETnfhq56118/UhOpWgPnS+jkVobH68Jz
wiCHJ3YvaN5ET6BfSZ9kNGTUsznZhGsHP3IYaMmezhiza653dtyf0eRt9YENHx/s8MQx8Qnqzi2c
z3Pj1Z99hk5y5EQeE6G9VY7heFfzw5D8urzhH/d9H/Tab59dWsNLsLWv3CBswzxj8w8xjNLfR3UY
C/pPpKjDLGTpMAwApfKbFa/rwp6y2rJ0q6SSoMXnwUx1EWg6KeGv+lpPxlC4d76OnJm9Oq1k14eQ
e4QsrB29in7nR+K1bo5X0edV3BW0q/h/UCfnfcA0yD7ts1C2Cv18q20tQzHz0t1189sOGho9TeCp
oRZFPS51/5w3B6JHXwZcj1QwvNHWYQwz5GE8Jci81Fg5aATPwwzxuVatWDJG9dyVX9NbjCbqFQjx
RowkP2JCq7VONAShyC9Dj66Lq+g8qv+GRfW0SUc8ATZ7P5rsrAxnObcr1KbiG1rjWAlF0lWUzeZO
2FGO8dKZvJCWMhTRMsBsYjHRxIN1AvDjz/E+GqFnVQBndQT2Gu8nsgSiB7nXTd52ZoQ1R3M/eIRD
x1645++NYHBGq8cwVg4dH4eRLuZ4UEUUcFsZoZ8LxwS4UrEKJqEnfE4ojBRzdPm5e3RZk1LiPyeF
SWx9xPOo4nmUbGUfEmcoTWO+2xdGmslwc1meuxoFGoQH1dM4F8xVbFcTxcu1kG1GPNNhHnBRH3Mu
/aYRn1M4hr4YJLjB5itL2JwtZYZObuxqWa8gZGk4FXxmv2LqGQCii1t4TGm3sNRAdJ0IlDGzKukv
8dXI8K9QrlKmGMSHtq0a54WD/B6ZF/xszMRsRdvR/F3SxxI5prxaA4hsStAAgODd2NtUo0MbyGuG
+D671UVLnCManFXaM9Gm3ShLQX3dBI7iAmU01MnuKj6mXNh8YdZjAY85IgyGp/1eCkK3+ZEZeiGu
GOQ0kzoJBKsMFvkj5T+QgLAlkMANCWeRiNjl1x2nzWxGScOmmyoj+8pzn+Vzw60yYsRLC9lgLzEp
JQRDCtV6GJLfcYgej3NxCgoCI3MbFkEirgYWIhSq0oIBDqd8nb9+wCr9vqICd5vuW8ca6fCXSEwo
J0Zyc/2vmzybfHjP+Dd0mUSQV3ycYY6X7OQ4B9aJFQhgnEWP56hO4Bgp5BnBYpsMwiLudLMns/Mg
zKrheFGVvap5olX4eMh3RYN2G3nDQfSXYDeleQEI2KaqbbliC1iPQoWQ/P3cLLFkNNff+6sfr1rk
KnmoviD0/9EaKN/hNNXMqiXBChevlLmOaO/0i3WmFP5HiE3e1ds4pGAR4yHYB7zIloyR/aNO6fB5
nkAnzpbjJlCbpsA2T9Cf1FjCUauRMDlG9H05zFNFQkVmMKZklD7PCKFYa6I1cKVDlLhnol5iRU/+
VFv72rwHv8ciL9onnwDmL8cqC5vZFUwbS0EY9v2afnCr/TkwVXtQQS4mVYyTaa9RFMdo/2K3cL5L
Wa4tuXDXa4d2JG6oOs7oLGrV1KsMek8pz2p8WS+j2uxnIi8hOJy0ROsn7hVkL4RjNAJDsU0jmyfK
DP/QbE/ltLNX6kJQ9vxreWN5KrwI6ZK0QTXTS2nG0MESNLMOs+bCdMAJPMscXPW9sVodj106gzE8
2fWlf+gU2QYpDsG9RFW71RAhenxmnKJUzV/w+Swz1yseusfnyc6FhzdQqpi3xnlaVl9tJaAne90H
DTje7W7Dj2Ia4yjRyluTtkXYC3Ugx9b+fyIWfx3kAzBkC8nvUPKRmaKquPCbNrz+Dsueu7inyngu
0CUlXOzVYnSMyzNVs1ZCQXFzFpKOweBZ5CKHYYDeZqnZhDJijlsbMgIVJAq/8ll0y0USPoL8PKPp
o6md82D29bfdJOrjkxbOn6ZZrJOjTBMlzcnpsUk15oShiRGp7lWzOg6WGtKLX817zkKsGtFnMJen
HuAZJQTE9IWzJKH2oGGQQvB7iTczDf7wxM27A0ntl6vNDwn5cqn1IqXh42P9z6VgBgNnpQYLhDKa
Rabho7EDFq0pzGPAMxXKiNDvWq3OKAezeJnMS+FCdWlvTKvtfs5CwApk/lh0XFvPIOZtO1wf5F6w
kgTUBB6pNniafcbl09C9xqHlMvvib4f0BxFh1HZOg1GhFRtRHeiyS+ply8SepAjb1PAn5J5JYSiv
UoCW0GP/x5rQXLuvlOJ8dsqPlrAmvJIyTxiMDkm5Qmjxd8oK0Hhv8GGaN8l7lwbJY5KZoASoKTrd
b3LtL/eN7v77uE56YIej+Hkkg3Op86yY/ZE32CQ/1JCfTFrsvn/vHr6glZOIKJHR8k4jAzz3RbOP
cqZztlrS5YAG/ZhsrmFqv5PbxvGmbhQZKsB8QAIc8u7Y/QVwGFMPUXVE6Mz/lEc1OoxlqbGA/UuO
WPJQ0L1j+FUoFAGTvpQxf9vwrWNl/srptuzXtbS7PUna1qVID7EqODPVq5MeTK2t2wPIjH+FJ/xO
8FJ9BMo6NL4rsBTvpGAF+Ufx6dH4V+53fdjKt5Dc3S1zE7I+M2qoBMrpYZgEDLM1PISQOSJABinz
BQKW1yW6VF0rXqv0YunnaopKXzNU466o0Wd5ntmNoOJ07s3DPRUYJZwK71PqkW14wshcYDXmud/t
DYAkMxIhctfrDstWOhvHLWiRbyG5nl9ji42G9UN+nlUzOOC6Lh80mfstH7lPbTTSK8chmEmgEcK8
Etp1IM1Jd3TDchKE+kMdGYbk9l9PbZXcbnTpr1+mOwrzew5CAqUVBSb7FEGIvudF1iXr+IFzHy8Q
cp7tjpBmnH+Iyix6plcYcptfgz2ofsbKZAaMKiqdbgmlKWaDet/f3DNZbwX4BrYcGc0xg0GABwN0
mKPtoRNqEtX/geeZoLQ0iU9YfpcRb1umC6yOKp0KnSVtWMomdMl+vFGeYIcR/SFrsunNeQQP5uN9
49QneJgno0K44ObNIPJu4IAmaULHUKXZsuds7QhpwxY/eOsKb5bCih2sUIHOzKdXntwBfVgcn6zt
SzRVVtG+4b8crVb3e8ds8scag19o6cr8J6WYhuW2bt+6hyemh3PA2pc7+fkmxpyd8PMEAUXg1A4h
legjg/mM0ThPF3mY/0BBdNHyBHgYhDu6MVVLwwZScn8WbO9j91PR6Idy0abg+OxmaepEOWTKss2n
TG4vLgXnZhzw3TDWKj6V6NM0Lo5VJhPw1RQYmmRdZhj01KupuSpc1K9EJGeia2Sf33JDQPSpHQZz
BQWVxnKYgJpzX4tIwZxVa0hDPLbw1dqduelDyzxU6qj8mFsSWraYbcLbCZ9JXAvFfhgw4Ar6nvj9
UcNoKXrUvDm3Z8ig+MhEKduMiqvGd9IPFfKJTlKpjZAtBLc12nAdeiTzX3Br4hph+OOkbprdOE5O
mS6IfHdOm1h2ny9SdRXMTC8neMH2V4kQzC1KLUns975xwhozhNJ8HCx0h091j5nDAmBqvZtLKbNX
hiOSkPgqVwi81lyR4M5Na4LjsNPMB005eYKsq6Ezxfa8n+8SXHfgrR5w0fdEqxsU1NZxKvOSS7nr
WbFvFpNXpq5ssqU1sJ+1dNHAeZ1dBXFjHYHZfIV8XITsE2s2WxT7C6RzyjqNtqVyC081WdxOLBXm
JwwFZ3cFndRSp4fDIlDOB6QZtvTQzz+lKsMCwilMh4Mzp2uKMqHsoxNYJrfm92Cjef7dDg8cl5ks
1DDDDxzuT7t7FXu/3N2v58GFBX7ortkACuRPoNnAdrrjH0VltYFauvnYgOnI0rq6NrJaCC/xgdVU
wXvjHFFQzTlAHocHK8iQSBba4G+OpDbvdHFgmhS69N6M1BOhNPDVs4nvzSsZzlZlGw70bboKb9ID
HniVnJKznxkASct7rqVTwxLCYECw/q1AroFhoGYwg5uv56v5lvwligtoGfbGOWC3Vf5jHFIHs2vu
dOoe3w1WCHzrh1Frs9ECh+GGNzCGCSFyXaAHeuiuR0icUjHK5DscGSd9byt4YsE/qpegzYeohy2s
mIspvDGQ3BydYgrRWa2CdOvhbKHv82gBNVJHAlSQOFiHhQ0nfqqulId8N7zXpxRoMVpd/D1G4lD4
iiy3x43mMA4Uthqtnhia/a+/5h5tauvt32km568COMIWGgB2qI4yvY8/IzO6lum3aqjBrZotbIC8
KUhpzUTz7pSVGaPebFAzRKPeYHRjKa8FxHK02fghwByQg7iQd0U8VNyY/eDmJZDO+dGWSEwmKds9
m5dQzpQ4zYs+AEiUyiqDbdC7eoIzwlLe4Xgp2xznTtKDhQDg2KKv5JYumVAf3mVGPndYLO/0/J7b
aHV1OJ5LbpiO1MDNVUbc8uFZ61WNms/o1MpsOS5MTeVNwRZ8+5wptGXcQta3CDzL15xup2q9m0+R
GxXGfOHBt7ZjDIIHr4ZoRN9fysMh56FCUuO9oya2xyxdMTb3nDRE9csvHTw4uchKFlSwR//p+nfY
f4J5Rqesr4fx9itjTxtE58dLWeod+Jebn7mRr7hU4R66zeDGQ8kV9ghOMWWFwtncOTF67Y/tMG1t
DShuZakU9K8RrRgYpd3VJ3ep/Cnse3h+5YMpMhwWqTYv2qVBsGdNjIVQITc45l8JAfKOcscgomUp
C0DygSxQbyzAkXKkm1XD6OfDftywZfFyjsdjTud3z7hiAxBe5IyAhH0JA8YsrO+Gs4nVDSuxtH1c
H0onHObDVsk2c3ud1ukg1abNgZ7q9jmMn02D+EB4aceKotnxIOlgM08/zbJDBXzfCBF0Ik4cKGR4
UHnkp/j105fuO8rg6V1BENZ9O6l52ZhkJY4wGrJqP6Pe/gAaMLa8u9jWDqa2QRemRN7R4wd20Y5W
MJpPl9wIglvWqNKJLkWGHNl2NRVeC3+u2Q6Ce915HUXG3Am+z0v04rR9F5pUl55eQSs8lL1pTIFA
0rW0W96c6P1K+Ppf0bZmjeYWFnYCGbr5QXbNq1ygW0xHMKpOqQUpZx445ISEasql7DbroCAaRYHl
ZwkZFkJrnsUE19LprPG2ExctgY78e8HAiErssQaAEqaBd9Pl+9VJNtUtqicGwlD7c/srkpfXKPL0
6szSlHOBqU+d0qzPC9lVsQ8OnPdGbITzKxP3Pg8jBfBoTTWdXEyt+IRLprPFL8MkHE9IIieMhbxe
7ucwGY1ybliduRoZFtHetZ8jO/JvbpzGv18WLPFbrcQEPTL8qA7Cga6DQ3SE6b0PBdZuFa70kkut
u9xTtUFYYJWw8zlQSDTsVNe46wUlYtAdUY8OWpt/Yw3JAwUeV5xApT3tz7V/AoOkEAVV1fDDlz3e
K3xWwqX3nLV24ToR33T3lQtvqmIvAPrl71lmNReIABBjphqjsrwCScpRHFee5hpr38ZRrcPWGYtz
v19QMeuUJkjJcc3kO4gzBeQGLkLLeRvgiQs6X6/X8hQDIu7NGdLwI/fMtVpcHxFACoZfrHvrPZuj
jQWzbomfFzExG9wWmdM8kHQAdmikah6d+MURZV5QTWbaJIbB7XSp95zjlcU0QGya2kjESUEAaEJw
DxZ3cCc08gRkqqaFdUDNHf2DWKp792PbNTdn48XyoYstzAILvEnOGMwC4uOD+AvhfRaNCDmiFZp3
0Eg8eGvz2YoOTAjsiHG16RLy09GOfhCbyCYaCn4qxbya4S+CzZY9pMPaprvRjHIrbwBrfsUzr4KC
VtO3Srexe4ZqQYy0i1E7pQjqgrHaOpLX7wXL+H0WuEz1a8Lh7C4ACITOycA3X0MDGUNVyYaLNa9z
jbQDVVx04ro7cWAPez+OqO5JZk15WNOQOkGDkY60ii8XJP9lQ3BKYjPwYf7M/HzWsdCv+g84tfqS
9ANgOna5zllpUEaA43ENQq0pFyAavHyNI0dAVphDv/fryAdDzDRIm5uQYzqqp3O5cocBOf8IsdSn
Nqm+0HPD0XLFB/YWByI9s33AsZ6m3keFT5hLH1u5WXPLx72LeZXX3wQDoYfqpF0dP+rkkUJRO15y
3rNnNrlQIqtmrpuJaOgkwmErZanpqNnmcDtLiLr2DxI8SjlL34TDnBynnQ44QJqt9uKUvA6PJnWq
D2mo9kB9ZGMW5fOMnqv21pkJ535Fobh6mNnnFDhKCpydstqNXAql1Kg9vICVm81DuthuT+b/9LIb
hM+LEXucRs59M1OXuzlXGd32CvcL9Ny+cOBr+GZ5f0sHBHFwE8wmn68553hEZttd9tLt5tziYiy/
hPKsZBPrTXBQSbFxSN7PUwuIkUzd2KTJWWl1d0gAOBcVKjRrGf8I+Ui3xjYgY7lmIUSthH7QXh0U
Q8My8cckuvMbLkUe7nzvu5nwKSzfNgXjhrpVpWhxKv6XqrUWQ2VvkZwu0ZuCDNQhinFUUpGtwL/Q
1rultsGUZhL2nZ5ekQaBLFRUiSbT/i3+aV7L92Ez9TDgXOSq4U7MqwdHtu0cF1B6nKHZiFqekBCA
5zdah2eDFFT5bcMRozdqv8N7avoj7SsG8dm6IoS9rgoiyMHu/elBWAUMN19yBtH/5VJNJ8id1rqZ
GhOdC3GngUEIokknuI1eNvvQ1Ez/ptorYvzeFrTQ3h54fXlMXSqrKt7rhAMK8gtOiNXNL8WoS08k
F05btd4Sdg2bqCmOtoqcFV2MoD8/N+Srb/49pNvsjKhfs0mGX9BdKjTnU9GO+i9YMiGUHi0VY1xC
ajlWDuz1jMIT8/akSYuSpgydnVy+ReppBiusVGkO2eUTDEl6q281vMlkxQGOlumLf/1m+dQAZUkD
tmyAh+1hMm+PJ053yFGCNrFcNFUGCsBSB7BhOWPB7kdmHJxkTkB5pxVGILB2OdqKBpCS9rb9a6Vu
tvfciIxRTmDD21ynJp9xZI+uLqLRZFvzBvqJMtSNcWRiLTyr1tl8YB6/pUqCKC01f64b5O66lmTk
4DEvqEg4uGNp+fhUXSos4kXCTlUIrFag+9uOixcVKV34ICTboo0Bgjl/w/5ZmwwiG4KBE5Vt1btd
oyO/cPKXNcG+E5rbmx8FZRgSqa/FfcfTrPNnoBBeXbXXEpkGNrE1LvJACSpq92qIdsMbBGCUHbOF
P6gRw6PdXsGlTsqrp7VMhTWCLYt01efzNI8/BCa+1jryEMW7gwidr4U1fBxQVRmZu5MgoYrqc7Na
UnMxVQNdEQWMi7rZ8rMTNuORscMFFq9jJpAchLaa0SUbIivqD6gwXebJihNJr4QTYouDR+HGRudl
NiYjRIDrJKbaXwyBJDurHJBepAx72ZEe943IVNsCeVK+CZvB/ua/cbcnnzLQRj6TS1AtVocih+lT
S6TOuXfM9TYpUO+RZJRXkiufW9u5Y0HO/4mdY2210iqpZ+0morTWxzkDG7HcOYfow7Xh1nwqZ9SO
tele0cljogljH//1LKbSm+IU1XKFD9nT+p4Rqafgymx62ivicmtmR+mbKXQ3JerDeWI7QwHfMkax
uDnXAEkHxLXrcHQJ14tf0BN/v9VOqMYw3KgwP4JH79dIakBo1f19sS8BTDoY8xf+kodSpt8rxSz3
c2hVRZuMrH5pKC3BjFeAJTO0SdXVxmVP1jUeDwLIckB7y67gGJi4u6Hi88SS5ytEhXeX2ZHW1hoA
VDW43np69Gw9rf5k6VmtO5pgGSFf5WggIR+azCVF9naxjq7OFtQo6V2Ej0tfbMeKUXpSfwYbdOCo
unWxkyDwkPc3VITckl6yuuC4/mXwE0SbHv4JbYBzfmdodE/LQNSOp9joQWBH+poTkwDuCezoXr0Y
NISaodfPvCU1aTF9b5zh47v4ntZjvLfhQvX5PNgVDjPwiwIy6FErhmnBZ6sViWr3IotIihzTm3v4
F+AOhXL9n+34zcBL6sJsNFF+tZm1U12opjUCT4cRMsNlHnRVmV+JMEKMIbaXq9F4VcpNi1V72ges
W71CtmFr9DYLdjZ9iPS5akxi+pO+iVEDjYMNS/IDFxl40zfatKvR79aes4VBsm5uOkzHHQMVZU8A
lj6q+S3KMZAGhhFCU5xMf3cfg3wmF7M/ooi/ie33zHVDaxZTq7Dv9z3x2pmbbg0RwjiOy3DO7KXA
KGJgHhm2ia579nemeKUieXCRcGSX1P8liDjftiqk+sofliYaWXKgXlUv2eFGF8kRbkRwMwjOXh70
DgR70p/sMD+xx+OwJA3oq8pZpImbvDpt069W3yZHwMfz7UVZ1e9q9Sc5qlyI1+hGapM5C5yGlxUv
akfIdKoXVTih1S0KiBArhhWeeShUKLekmeIMpzedC1waoHBNrb8mldIj2EeeijMuThUEV7YpOqPk
reTF0zTREjc2DwviVNAAQnebM5gpOFCfyQ9yVPPo9eDIkFJrlG9hrhdcTvhpLG5aZuGQo32nAr+T
ucOGUfQ9jAmHnIoPZ5yB5hNripnki07TorRMgDl9XInB56yvHzFUMuZ0sIyeS8gg7ri+r+Cfx1mn
P94OO5g7gBVWrNTFy7WL8JKwch+HBlopNUQfN+LuPG0vyiQt2jORo4+pYOmjG3tqvZ4uIDi/sLjC
W0I/FdLFM6jGS0fiBNnNS1Kb9LQX0bAHikNM0+13q8z0trNnwYju6/uYwd11dIR2HrSgAlyA+puc
8O0yz8UHX8L1zTa6dXaY5o/DXx65AvHpYdnqyXBw5+M3aSJOjFXVOtLAPpv+dOO3HRylKExmq+4y
qiGgLTcIclwmYCVXD8qIirI0nXw6PmT5HnNLj3MfsZocQZMgpsrkBauyPNOXNOp02HKHPJR5dLqd
Ij9uxh5twd3l1MXS88VEYT0EpMVYzqWmZcdfcM3uo6N2nPv78yvKp6zd3I3XQfLfcmtwRwwkFR21
B6sQcBA/3YX6sDa2iN3DiuEssKA+VTT9wJpVn/1MY1mDaq/8F+41KU6+nBXD6OpDeCEbsPyXxo70
qV/ELFjM9rec2x0gjynlEZfxW2e6gzXf9xF+kqyMZZ7C7hjPpYYegZC7/Jx+iVQxEB1O31lNcDb+
N/dTN5ClxjLbuEb3pZ4SkSroCmHAmfCPxw/Hw0HsISn+tWP8MchUoYh90f6mrKsfgh/oxVVPX2w3
zZJab2Xf47JUAECY6+3Yq8LIFrRZmyjM5f7pi5jHk/IILqi/JWZMG0xMOusQqGOlNveT11Ut4v/F
d3tt/iXrpeb97KPISTPua6yCCgi6QMo7mOKl14VbIMgGoY89xWQrPRwTH/6q4Gy78kjoK5xz67mw
0K8575AbNT3Hdo9sQZ8DoNQfKmu7D13FhErBBbu/6nmoOXHaCG4VC2iUzxbCsdjkCEH5r6A8+vKs
WkI2AyFvJXwb47sqKg4LcmUX9MgpcmA62bQYGwRHWSpSJXRv/BCqlsGJNJ7jQsauUC0aUcDuAa67
NKoKQjCi5fd2owzYC83e5XlTL6hvrjoC9iKEDKnNQYTf+8ZlyUOL+HTI8RipLuQGKlJD3b52JiAA
wVSONFOigtBiSa/by/F5+mVuXUf3ODQ0RoIG1X1G44noyYXmxP2eMpkzjyLBQpnlpkNv18/8oxYy
AqREsV53Qn2qIBWui553mUwMX4wsyX1xqYU56NWmeSKI8UGYZ25wcGpVaHkYfjKy17y/GF5JWb5p
mnpU33M0VKgOiTk27blyF81blVP91dhdNVuRE8ZOwlV0ZjPNC/3U61Uq+0/fOYFrFwfPaDm708qR
RgjzZLnPzROhVfSDYy/9480kkqXOs7g9Gc0Zd8+V1piwWP3ckExgXhlVOVALh0dw5vVHx8dq7Olq
FXuuze81ZgA3/VItkjIZifmphvxftp7y+E187Avph58NUYpWRtTojDZ4vrarL9qL2gsljwKNI/O6
v5Jr7oRlL0JyPj7DCp6Y1tU5Jp04L0+cgtJi8D+/+y3+MQyI/zcGAK4REcm7fPOTxuewtjFjUDJN
qKGyAI+kxXIES1PcT7e2P8SleREWofWOxXMJNvb0bs/h5shN04gucwDxyyYPC6lYqi9xfivtrfJB
KmJ9HlEbYEM5kkcBlQA7sdvwj5/PyC10qu7qfntR0xRo29eolN01r7+Cq3oTaP+MgDuBhey2W1XY
c4R53zGXqEhVDMmrV2fu6k0fI2mUiB7Qdhg1FdTDqelZixq3LoftdxjLOF6QmFHPhJSdELSq1lT3
4OwX4NTlc1MRPBxkaMFp1Y/ZMPe8AYsCE5OYxC1ZWrRZ7+hOGYRQtmr8F8Gn2PI8KYTuV6yOYKwL
aEH+6AjYw2R5gk3DNOYQmQ4XGAHRYGVoakX69U6R3kMPTocM1eW7urdJl3DZnE1eDm5j2HQKYkTr
CH6Q/p/41XiRwaWR2C1XF0qCsOxqRhDdcQ0RSC9hNB+lSIU8GHr1HEP8n696BCUK4ubQFg+hH2gr
Yd5EAS87HjiNpCbSRN7ZNZW8qww+hHAI1NFdrq8Vmyn8ajTUbCyPUPo6QkbWedfDduphYYX5/p3i
vpLOQcjb7t9UQeh80RayvkNlUS3TRvQq5T1kNd5STXAMxt2no+4VWRUsQEQINnsH8YzWnBu0LTKE
gKUUaI6Z6fCFQkw/PF79tHL8BEwFQ0VFxG+RmBDp9+xmb0FQoQwuaA6O8J9HtlxkNvi1nGo0/o4j
uGU7oEb6ojLF6zZVy5OB0DFkOkYDr40UXbuYM6OvzWXhlTocDa+GSH3UmEML20uIuvCAzhziF+46
0/i4qVSy0Qw2l/6VkxWwHa4xgWcoEbZFJAmNGKd1DqOfatCGUJkvzcpxmEmR6OpqgTLdLoyOU4O0
LooWl0CdI67OjryOHJypUFHtVEwgKYgc4qp1OVsy5RlhcqLXYKvetzOyGv4IHSns6SeY4OXFd7lF
DPHHt21HlP7lcjiEh2kfQZVZpvZ6RWsNK7lFeb4fIcyPaF11RywUi8PBS5lHhMoe4bYMGDgVP+zm
9FHqazmoDgYxpeq+Ccpet0B2YXPxXt/+kxKdqtYrQ9l+nDsP1UC0Vcr06mzd7+hgn6NXuOtaUpMs
rYilx9Y5NxRo0X/CRI6IThPeMKpLSg+vWacZxbFNvYeRrug2FZDyMbblq27i842b7Q9KwG6DyAoj
uCoyIoKSm3WGRiOl3LgCepCBVftlAvIumDGnWYO3UsPHQWp7eimykZOH59Ct6GUEYhhpobQL/yMn
tLSrV6XWMAR1b+06wIlawWPrRXJoLCl0/io5WPky16dZghpQEvNYy54cJQDf033jvugXu8ArgSU7
dBeBejG+Lz1WxvmX13tt2g9Pu+kd8PteMFd1A8f0UlPpmheyCpC+w9YkJKz31ni3yeEeb1SlIHUO
b5hSjAmzw/Z55I2DZtNK5QlFCygWcv00eJvvCwQt2mlxQ1qCjNc8cGz7wzK37cfos/5kW/DWTquN
h0/48oMQH+PGYV54LCl1oOMwcZrTp4fIVpJG9EpaKcKJdN+FCykHgxZ4cnfVWlt5WNECmaoSk3Ju
4rckm0H6LBXVx+gBoqikgzoO4Iov3SSLZhiFyn2e97rATo7BC3CmQThRmDqG0fmY4dk30I5Cxu0O
wa0zZ1RU+Z7OYq1f/FRT7dzkPBzXeydx0SKdUpMYdJQgI9IuOMLEaQtYsQB/GTvVBGeKytme7E7i
EbRsb15cKF8yRcLM2bKh2T6uOmvw3VwwvN+aiJOVb+0BHgc+QrR+uFGsCG3QDOnJWQjy0PMGZoIS
Uu9Nn6RfsUH7QKa+Q7Wo3Bs8P7BV6gGyOxpho5zz/zNtjsl7zQOK6Ohn9E/lrSPBBNOA/EYWb2iN
U5lyxINwMmjdu+a1ms22a6fzlnulAkgpTGA4ECx5utEhyGbvcnoGQbRPPzuSsDiqY0tgXkGDygQv
2qONstty19aHYXEb9OOQhMaNm8PQRpQwodEWuq86kATlqJAsE+tvchc+Nc0ymYHVFzfHGdrX2IWm
JixgqhEk1w8cwgrkOhKAYUUMYpdaHUho3rVDRYZAf80T7dODY36u0NQM/2HyLewb7jxvxBM2rDD9
UR3xkuDWpGkIK1oP5sulAD88vR51yg/kprugKJOH7tHDlZDkU1pWF1ytEDSX5Zuujj+NEeeEG8gf
wEUU41w/daV9fu9JYCJEV3grpRR0j+tuIZBiNNfA1QLrE2HYePMu/gI0JMp+DAinSVKYNKxGXuE6
8p4wzliOpCE4l4YcziLWZHiIKwaLdcqN8emKyeM0r6hBJC2HskipzVxQ3mPoQ+5/cb6NC5MGPuzE
mWOKzMBXgSpWFEhxhCMgpP3j8aDLYsXfdVWbi1UUq6Sds3+M6odw7SaQ1VSR3OedlbViIQPQQiCQ
Q7qrRkc1IQXo6rnzvthfcBeoORdd2UYS+XtpdW7fWTWtDupDCcQs7kjMyf+lYO55us0JKiEj3OZm
3iVajrws1BNQwZaH96S/EmJZiciCpRtEyBPmgiM9fhHmQgc75Dm8LfF2f5F+IFmCZB/ugQr6quHl
H+6kX/B/pXC0oCjWOKsXirpzw4tPM1tsGj94uKjgjCIFrwBWIFoSTs3U6+ym8r4i+ebx7oHKDjfn
xOQd/tqtSw3LPZ3S/Iv6BvOV8slOqaiNwc81P3l3RVCrh2pAOxcan8WtX3eOt6yF4LsHq7aRFNkl
JqSEeCMSJgEb0oTE+70naKCySKsGJbwmyGSo6a4DZVoe8yDL0oUHgoAbHWzVZxEroghJdJ7jofpT
toYf03YTcgFLMxpbR3sSoknegOCWBnUmaN9HyTtZifJTQs826FlpKRTHSM/V5DmWI9zkI28TW3nL
snPCBpTzks1d0s9dntt3TDI9WTPYwNxSo2PVNPwEyuKGp64kjn3DaucKlYYsiG6ES/fSagycMblt
vz/87r05zjqi0PrLq2MsgBrugBdt3hfXaIkFx9VDOxexyPF3prZc9PXgAE7kHmNGXkMAlcshu/jz
I49DaumFuzRTKGIDB5HZMgDwvWpPMZjKBaUStZa29WlQx3vgtLHYyKssUAtdM/0sKSMIs7mw8Yz/
ozGla6N+47omLn8w7IYl8GK57Ee8o27ciq2MiN6c0HYq0XtzhkKjk5K1pDMhf9vxCLNX6E9QaofG
FydqjYopsmAbsJJGU4Y8tteO1YMjvoe9vsBBb2ZW4YoiYYneIp5rWdp7GmcYt3wmQE9ujZt6BUSL
yCh8xUk3BDJDVr7vm1IZKHtBtetmVdKy7xbfZ+LnCD8QiVU0lZqpU+UZj76h54SxDz3ZaOfvegxm
CPpmipesmPYaMtn3ri/Pdb3FoxHF4RWPqXhjlX42rZdOX/2vl+WpvYkQV+5PSs2Lsg6iGX/AWN+f
mY4jMbQ9vP2oMDDKau2sBmLz93LjhGiK3ThNOv9ownX24a5yzHt3oeiByDdcfuV+FQeH76sq+M/K
R9Sz89aHyisw4DEM+rVA6uxy6172FqlVF7sEFoRs9cqukjo9GMQegkT02g49KBtzyZDVETtJaqsE
XRL+Zcmzlg6I7GtewaHOf02kyLAoJSZdvCOHn1Un6IdKn5wUQDYqayyHe19vgRtNa0/InLwe0zCI
n7bEcQYgrLoslcC7oxf6H6BladwYMp/gfgVa2CBc3PQds4/wNXBoSTMjveNExFuNeFoQCs7gL13G
lPePywHZBqrIFgItuhEhCw6X/pplo0BybXwMx/2mWCT6vjwghSTu9Qmp8HzgnzhOhC9Btx2hqP6r
NuiRsYAE/4So5bOz1IdRC5VEo5Bn9t1HAi2CQ0s0YzsYCACsaFD6EsoBXuAa5aOZKOs8TkB491ss
ty2bqWM6GX1ZJkDbxaiuPjZycRIsvu6MeRcsQuU33QRN7dfbWjr/Qxny8AUE4BciJ5ulOzg1EEiB
6oJiTqbOpebDRjOT81VsIdzf7dmRO83RVBgZn+SoB6gF9IJjXkgBI5tYilI9rjzN3ew3+0bpMiM9
D8Q3i7OvWaM2rjifFcd8kIxnNApDnZatp86DiiP2/0nMZAqoWhRYYsujAgzrYkmK+trx6SwCkPkj
pFaqFXXLJgk9I0v8mes6BHTYU+SDRmFCYwjSJ3/wZbl7yKk7JoDz4gy5y+aVt2RyxKNXHUkD+DjW
TtBchSuNWN7kCUfhziynK0M7hQ2Fj8W27Kz+HBBRSb4GzaIRG391N/kfU3pD9TPz+XcPoXkpZy82
omCdSjuYaA2WWUckbzU3uOezbuIhNV+eqSjwvP0YIpw+9k5sn47NHFx1znV8RcccVms4O4c5nk8G
Httq9ReQn9b3kcFZ3ykWTcesVccI6vQa/xdF/9gjn3YvAOFn0ZmqBo/3IXay9P9toaqju/2Muwj1
kRtgafS34cEw/3hweThWTMhe9EnYSVcw2+T59ZgHRzhrZHROTQgx43vg7xO1AWRulFD6tvFdeeem
Mtzdb02oBmHWbkdbDg6Nz/bK/cgQNeLAm5dATenFoQrwsdiXnDDxsEehvJnsM769DTcadyXIQpUw
MLtSff8PHdcPCalIYQe7s0wva3JPCHriy53FficgS8JlbN4he+F2iy6DuB2I0FAo5y5RRjZeOpDr
WQkgXVLAAb25KMH56m6Qvu8RGYSmg/iIoIk6oQEC0PgFVJD3J03uPB+IaZc8O+v81obLxamvd+fJ
Pmk62oRXgU/Pg0rxfC7DeiNDbYBrk7UbScmYvpPWW5Wy5w9zX9HRxSEc3JtMF/c4c4WFypXV/Z8o
D8WTyIDNCMJA+VY2SSY02T/DO5FpKjKnwgrK4g1wZVVt3N37zqEz2LwfotWxWqMUpNtVdsNK3caE
/EoOIH32JgezJTEAz1t4YRaYEQ06n2RyF3/vPNS4WdVY91gNj3NOVzfe5F8W2e5U3ML+i6Rq3cqW
lyNzSa/Dd5qUt7Va9ZZ2FsSc1Cg97rva0rjHgOIOundpv640WL0CgSbSYZiYYsB6F7iTzaUKR+Y2
MUPaemXTrQaQRvJ9Jau4lz7rdjUAhDKM8UqfuPItSaeObiDh8XE5iQFVdd/UyglEti7VqN5yPWWO
aay4cYlKOQF1pspfG9ghdCItSPKhFk+ZBkATwKNG8C8fOkybIwHqikK6gzduq7ipGk3ujXWfFMYI
Gtbel+CDcBYkOdnlGBX8IF4dsV3eraD18ulQewqM7+ENYFtvuMCEUUzHTkB9I68hHPU/722oAOfF
fYbTKkKYPLPPekxlhgvbmwLHNT6GvhqlYdHHSrQkbvUtCcdkm3YhTFt8FxZWhKtZgbPNjLn/yECc
Ps8n2MXY8Cfx0kUqh7O/Ew1dSbCxHlAkHjzzTiZ2ZMBSP2xTm+QpRvygHHIVnHMBnqza2SRQesm9
ZHr7DNSN7zSgiTyy//CIgTFxAuDoeAxKVq4PvGj3xxuCRaIPRuqGwFp/5V/S0LXrTcuiowhKmb01
o8NgCZcxyxjdN0QnHruw/LBuo9JjKkLtIiMq+ii5fayOmXZKnXDoWM02AgPhr5KqOFacFNYX60qW
WWPBR3uMcMrwDk840tvYS5cg9Ki6NHSl4oDjhv3JUvcaHDCPawl8Zbxge7fFPL4TGHmxu3OcSCQh
wFz9dvcMNsXKRyi9vu8tjUGUNW8CY8AixckK03pmdime+h/6YZByBmgg9++BpDeni/55V5Ekw8mN
GfZzVbBj2PGOQ5hpIJjfLsea5w1Po1U098qxvOPsEd9akmNBk3v7ULNzskWN36tzXTq0IOZPt1yT
ukxE5XO/kJCmlLKKIJmJdZFe86Lq2HviMMglcQqD74bFMIinMhS8znQUPKQiRC3m4dsaQMdnaER1
nqJbUmsunvjaeybRVDJ9oK5YwbJWRZIcsbLTY5IKcY/gfdyv7TZ2bw4OAr296mCJiYun32ffszmA
spXsJogAs6qUZrbl+kjHZPmFvtsauhFT4lgS6G28vbewBwYcVT4rIGE5p0h7OTvclWK8knYH7I6G
VEVKSlgBiTOjzTWz0RiCjIzGR921P9GVGAUnTvfBm0mSip7vQNUZtvB9CClD5Z0wg2pokHAY44DW
LAs5JwGqqcDGza9wWY6x2MJECZoUX5AQ3VkRLNNxDjk3OnsDjoAlHLC/xGqE88y/Fc1021Vwtsnl
ZZjYr/T1yx7J7Lz9nDN+nGFQYv2tJTeo2c8l3wheole1ZQcYQ2NesGmd8TH8m6RDo4vgbxfdM2NC
pkAK939svc9QpAqJdYeJmR41kE8Q3SkdKhtNXQajhU8Gf1lwMULe8v4+gh5KVAKh/jVI3Ytjcx1M
shS8o5bA9fxB4lOVasdTDkR6KdVKtn9GfuxT/mzDYiH3wV2CU2u4L9fQ/zQPfGhOXpoiHynyZExg
GlFksyb6GwMnZuhznTereH3l3IqTfSMPOHxkpny3zlEhoonOyX9ho6d9dPtTQgTgZu5bt+sx2Iu6
LDkWQSfS5eWk2aUvKjvqyDpyiMXSVOfzsy4c0gfwXR63S+3MOU9lhwyoYoQCaymunZjxO6OjzwX+
AAeVORGVSVc3Mtjvy5CTMYxbB+6aoyKyB3rj6y08kbg02jS+HBKvP+vRp4THJODwtDkosiLp3Zz/
5GQ8CENeGQ6CI/522E2ow1bAgu54Najh55Z5skq7L3f738oCFKylrLHTZqwOu+JiBGEh2weDi3Az
N5ITQd38MvqfKKlQBBE1TPUhLA8Dou03xcoXr2fuf4c2RcXCDyt1pUg2y+Sjj5XLXMHtRY3p6oB5
d7bdWg85AwJoym5G1NOZTtVfe6j5H61TpeFEjH0GcBHoIp+G8IW0C43HABFkABST1N3lCP/PRdvh
XcYsqQ/3u3czvB3gBo8VaWz/hBzKp6pSuoedmiS1wD1KIgsZa7BKZ34qA6m0LKLe31TZWinUgMpm
JouIT/4tYDBCRl0mz/GjL0cg9y3iei67q/jYNE4dQ1/WK8dY7yyMb6HLrQXdql6ZnIyozJKiEZ6S
VxqAcchhJ6NVKfzJK/bWVKI08hKonWEO0agtUf4RH5fvLIgQGEIzo28a8qjPqBgh83wMLeT6pvqL
tkzoDQ3jpdSQVxVe/pVfZTfz5QmM0pyQQ0ZCSRW/HMVC8koLWbIB8c8yhicz499xDhvQUMFlHYcm
/D2TQdxsnKVinOmCT4UWFsfuwZAKVGiT5RouDJiWtz6gonphuVaBk6AvI9bjbqLdIseQXJxHvII0
3CyqmzgAX9hAB16vBWDu0/n/R8mv/QFQ6ueLDPnTk7OzdN/HNmySwJIa7Y0lyfehyG25clliV5bO
wOeiqxasALa9HVygGTgCqKgQ892ZuB4HN9O4myl3t6mAlt97WDNNPgaxEmGvovjiie8vuzaFwYwY
XRuZ0bJ+HhRM6eilPvxPHOl/OwJ0xqywGTujqm+I3KlW+cuYVfyo8vtFXghp90jYG8qR61rX47iO
zLdEt47ZR0oqzaYcOvmeq+bM4ua6VLKXy8VpvuEOAd+yUn0XP7F4oUPg35ppCDF1Jt628Cjuolc5
rI6HlXKHHavrCdCaP7gCTAizluKI4b6cKXVbMSTi4RLu9ZSvytgg8FQB8WKIyiJWwEBVAAEV8iNk
uJFaAKu/LGmZX1tYP8Jj6vN4DiTMb+vadNHGY6xHuxFwMQpEOH3G92/7+mUS6hM9AKOFQFlcXfjN
KvdV0EsxfH7HYyOedos+HqOVcmig9vIYlNqhovIrmlhuePLHJDG+RDwlNV2Fq78TfJQyZwRhfGGi
hAhkRkO2Pnx4Czz0TU8R+Vr+TCTc/eBPacbJyssaAOBP1gWK9z4bzDvWGVt1wrBUfRTvx0ulf5vu
6aSZHK5hx3rRVMlpkYJPU+yQ9N1BPWNDS3PC/3+Zyc8mY7tHFicT484AqygGb6egmpWcR7PwzLhS
o4XekM1W6ToIC+KWhg6x2lqGAPkg3UieTVwc1prhjP3xQH7u9g4DqUsytOmM7I8krqz++WjMkc7a
+qXsr3HxGsJCzqzJ49rZlH+fQ8WVFZPJJuywwc8Ue5ivOGfi0kdx/Xqs7uweB49V9mvO2w/c9c42
8OHc+HUU08jUTndPnmF7DZqnvPx9tj5KpbcCcJH9rd4/MlCbjiOoxbKx9H/FNEHAXPwW1MwWAT6I
sROBbBWHKY0eOTkxo8BQ5nIvXp1h90H40XZNBtlID8Kc5245uN3Ntcix0ILCdRnDMBEkHy7vCMKn
EHk58BRHWUOr621SEY7lXcwGi+yH55TBFBf8r3/fVYuzdWiXy54R/MJPX85KKiURUNXf215rorqk
aYIGSknRcUuYl9RihMZmOsM0a4HrLAsCrnyLXH5b/xpyRr9y6rq4tbj3AYCKFPWCdqGzO2LfQhcB
S1uBP+4D7hUNb28V5QAa1R3LjZmq9rZ6XVbAxgqDKcX+Taz0GkihqFiJu2DjjQ/JDr6AjclbhWsj
ONTslaQMbHoJ4o23Q6S9JVlA9Qfl8rfulW1JsqIXbezu/89vadFtxK5OLW0nWMhUAwilqe3ixi9y
t0PFNjoNjP+oSsy+wn9iZHu1SSWcNaPXU9hcI/M1EJoYSfgk2NBkUwrYizSaXrW02+hQCJh/pQeJ
wVH6li5KxeY4/yhRHOAEYP7Crnvjr/OfRboCtfamiSuS+29XJxj45pxoI5zAymRr9C2MXkvxzSZc
xigfnuwzxv3ZaGra8BYnHLi7keNDuCEz61mqvPDyjbPG1j5H8KNQWbZvCvG8Iodzyde7Zd61ogpw
7vT0tsyRc7WUewMk3a7V2Cx1lxdTnjVCYj4WzsmJ5zsTvXBfO9w8p4nkS0xFgC+/FJzFIyiKQVrk
tuWy037Ee3PCA4RZR7c9Wl4Vpli7kZ87Kyl5N8pKJFFpWRoJwjZRsxqSabCv3jFugIgzND26sLRF
BVzkyTWFXSzoghT29sPUxe90gQ4i19UVwFC2n/3XYuMO4lmvPWG1RJde2b54aBWLToc0okpX0VZc
HuL35ihXNwsAr4gp8vGgGt4CrZuu421u85sH5J2NDSfHW5XiDYBZz3xFK7t9tk8O/i+FvV2sIpu+
vPSh2Gjh++rLDsQrN8Q8DeYgwl71YD80iy6DPxAMpv85Sxsu3PY/7C/c+VNjVtSAmU2ZEVzBaTPE
6EZ4O2ifbBDd0+xnVXFypuYLIFy7tKBAKqt6+qiQH+RXcDWLT44ZNk5WmSAOjHQD4218Kn/Jh6LB
vYq/cf2SQFHvfD3zXyuxalX3lDfXPYp0i5ClxW9Zeu9I+cepxJjzNlZ/n1bR5dBrbJY637CmDe3u
n3mqwpugattriIiywXEy1MyyWMp26Fk0MYzwO4CaiFTCKEbSbnVwLCH+3BGO7PyDGB7Nz9iBlDQj
/1B7C6X9dgifJtxesnwyJMkbUoANx7IJXkPvwY5qSUQYk5zGyj+iOxecY0T+s2UkAWJNz7ikVtBg
Qk8ehNwwilssa4mZZVNkqeknQiFO1FRBTcKLazuvXpclr4y/0Ults6u+6nd8akjC4GpgyjKkhopi
KuGrESoDJqlcV003LteAS5sUYElUmyLD+3hkRBkZKpwSOrdRdwZTMR9A3W/sL6pHukjZHXKp7i3f
At4Dd6DJJslUH2mH6os3WUsnmvaUR0qycQva74UfzBfd0am5Ru0XCc38rOAelXUX0X4o38oAJvQa
Y5H2ZNOqpzqEm9UR/uJzoJVRzX77xbY0u9ueKXQXKwQoStbBiH5rnWPF6OBVatVKSqYgmgkWKk1n
HoOmir+k7IL9jQYE87ZarxkM1lRp81IKy0tfshj/USpgdMhVesly/oZO9zODRtZsoAOGANNtuzQo
4l3Tazjb8u4wOuNYe8TnweWmrnFDNwkAEuDmNYSkM/OMwQ+6UZRbbC2+uKQ5PENwzFnZGvU1rLzy
9iMulkfiAgSAO9WFIcvErTRJI5/oC1L3rNdWFvpE5kCEBZeQuouJpImTlp3KwS9aEDB9k3qAa+Hl
lIPkgcPgoXTKPDPkka2upQ/N/VX6LzJjWvApqplUKOAktn72GXEmqQzG3kLqgVwGPfYu7X9cVYav
AWriCNEBjULBt+X1io6QvmFCagB2z091fbXJtokIdbmKZPOoBMmJH8XEulwdq1nSTv61ggGJLC5S
Ie9WyHmV90Z9R2MI3vfSM09CQLLj15ifzTlLmDcVfAQkI/lZsRB9lqPSqbPSnfQo1fX8XWIIXGEH
c7u0fryUndSyxkC1gM96GULqXgCmETQYQ5qMenvwB/JoivHzfhVIBydQJ1L5eXTbHry6VmFf+eAr
9jdOowug18yVJ5iKKmQpLvQ91No2YJucL66yAtQLGlQVH2gSDWDyNPCJLrMLBNrElik+tz1mF8dg
TH3KvWAi0dXHUO9Fd9NJqsw87PuEtnhoQmGQejBaHa5MnYv1Bgq4r7xTUM5xr8Yo97LFFReiTvWG
iZ/NMJk/RvAAinO6hClapQ5M8zltnH/waEUG7q3LKYvTAolAbS5QiDhUcEBTVmvMAxXUrs5rY5kz
k8O2JuUJ635r5bxhJLJA97C6I9Wn3b7fwe/4ZwIzAFv5As9wIYYgtrF4/a3v67jRNs7J7pDLLFMU
KAv2L6lacXEZrfgmMK7Jxnv2QxtM+EidEDgkNKOo1eVRTBWrPDdPVIfrIIBoEteISZen+mop8Y7O
MAleAknnSWM4RRvlwul0bWzpMDv+203kafIHDoQv8UM5zyIXEcNjcPZqiTN7nihtEBrHV7RUYW7o
TVU+2GVIK/Ezmal9Uq0jGVmBOGTuJbI8ULsXS8vkElsFKSjUGe4vv3aDTI8HR7pmVDVpKCYqzNY+
mmmwNdmviWr8SQZuo5rdlUbwWRgObn/i5Syj68Xc/0HLqRA4At6kr93Nru/t+rxuTcQcG6WCyQwV
lgRL7Y4/rf8TZOcb+6rMTCf0dcPsUVCuExjruoU5vjs3n8SJNxbTX668fgnZ1iegegpd6mxbD3pV
razgotIOvu9LzvhS0Sg+oVDdqhvbjVm8I7q+gnZeajxo9l7dNR3wP2Sgq1sMhOAdQkEU31j/hd3H
eyRVKy8V/77Vdg9oYO1qTHxfO8SriqjbZTMaR/fB6hF9i5FS4Uc3YSvp/1jYgGpSquUjXbQkJpWH
mlsuWhB1eP0tICyq3BkRYfoMtjO87kjLFqZ4MjPfDbVHaEpC8nyC5Jiw1Y9X6kGw3DHGL+IJ33BP
EAblid/oYLHGMTQC/6INbcVVKBqoOAz/skskD3/vjoHIRgRetrezfw9kY0du899Q7CuE76qW1/og
/x1Yecx0iKn1w6lN7/zYyePZgK956ALDykFEzzcliMkL6A6zCdQCS5EHCcnNf1yodtwHrEYhHBu1
lx3ki7Qsx9OOfdmBAoc9vNf3uz9fIYDttP1z8YM/N/M+xSQhDN1P3MwoFyX1C3g9rdWFtIK9I+6g
+kIrvBMWd8VOsOM8saTQcaHjl1W4EIgwyWrj2IJ8Bi5mhxYBD0iU6iUapbQxSaPYRVT7RGL4umT/
hhYS2PAufor5y+OL/i/BaXm4evBplbI9PkNAhjs6a4LX8H2UT2VuJ+Llbo1XU/f6jMY9I40OWtIu
gN1l/z4eLWi0kvBJ85mLLzbp4fYo/YONOgJZbmtT5FPky+iDpnoskS9/0FZ7y0/KLd8Ru5HUcuYy
y5hCk+HXpvrqUmnCarcWezOCiFEeTNq3SOsRaJNAfojpYrdpbMwvBZTi0iWzzieSydkG6kY0wlJC
xGE//UbVhicStTKo8oPZpVMaD96EX4vO/2ZFKSmkJXkC5YYxHaGoBDbPjVMC4ghfGMc/S5GA29lw
5Y4Z4Gv24O6hs1RRaybl+mCmGmdYgUOiFPucBlnYomNd54A1XVR+R89OxQec24rXdVlhJLSTlxqf
1efA2Ps64+jYIhN1sBDr9OKv2Sd/OoPnmfOFZRba+1RfkNR3kXSX9FEl3QR2OKtCN/eIPVZEiI9J
OmzTdIKAkZEBv+GD875LrjKAQSbs+4arL6SS462o/pTUInrESlke25FTsphsLtdMBoVUVh0NcSpk
ezUTi2ntflKY2/K9dwn+kP+18JAOU4noOc8eXGqiiYIK29dyF6M6cPCt7O5syAI0/7cCx4y6QupD
KSHq033pIYYEiMsyZU5MwJAmueKiudiwpwRXfj52Yok9reGmtM7DoYAmT1A+EEJ0YffKKnNI4GsL
0WAgfPpRHq2N42JTHnFrHlWIZ/Oi5CTvG0KGIPp9Io7uPIZu/FBihkwymacsiF3/ROZFEZPOTy2P
YCypm6G/Bqud6vF8ooy/0vE5xGJLoYrItU+Ku6VGatLmT9l8g5zjvd6D3BwcV1LXlO63XO/SqhnI
mHL7INXaXtyGqV2f8j9cubY0P1cwOPcbuqd/OA8u+0S0W36l5li5itLgINw3V6ASnr+HAb9koQWs
1yaVrtyeGFEj/B8SFx02Pd3NYm30hVylPArDQ3+iYu3ddXrntR/8dDoAhgDk+JvrpjHI9fDcsr0i
r9+yjw69SJ5VbgHeaqe4JrNuhmC5H4sy8gLsN3mcPZCngidOYjWLDBPLyy505oDd4eOv/z1c9iMf
8zTh3uPtLVR2FjbfM+s1uGnN1RZMYE0pEYra7jvIdSLqAjCNjI90oDJ6fN6sXt53RDAOXN2bE/wC
jkwICbroD2KtN4G7KdlzJWtj36nzS1uf1HTpRXnb8FtPdPHaF83PJV+t5LpUudHqaHiEeNtjZENs
DCRtEJVYEEzRtFg84jIxCbeZu5T6qfFRtkygxOKXVuUTGEI8v4sa7LafvoVwDmYDQJ7hhVuMoklY
SJ9LcYyH8Tre8dK34IHzZlYWpXIsPuQDwaZ+QOU+9DzVPmUfQy1ULrkQrunqKbCMJJrNVmt2gVBB
vj8Jhi/nFAAH3J8hZiPO1silz4rreFpUTdYbwipMbzi0tnCREA7DirTzfTN54wggFA0QFHqZZX8r
JAnBOV0HlEKWQJh/CKwbi+MQ+qG8pkNUQIec88uEUXBeVUXOoOd6dCc3mHHp9O6byu12Et5bIhxO
XDEUIzIdKnyZZ8xY1ftsWJNStdQo+vRrgWZ3odiuV4vN/QJvFIyWKZIJwJdz96nCbKwtZt8shO4a
E0+2zhYmJtqZpmAq35nJl5tnNX5gYD9/TGVk8oXHfHjPfCIiqSZNblzdONf+ujX5LhqF23gNSCaT
0tc6Uunw2GZS1DuTr9py4BQHvFsD3YjHz0eeJwE9HR/gdhtzC2+vbXVKEaYw1esXPnvoup+ZI5wa
XeOlwSL/+DsUD/nmfc7ZGmixfVDw48Ex1dygbwttPAqjziCxzis6D9njUW1UNEJfUyB7w/5H91CS
DxG58w5TSMFnN19HALMzyo2YLHdmb7PfUih2HWos8ypqEq+u8dXytM66NtYJdD6JasjOOgxVXNze
iA3mPF7+TE/pQ5/Qf+W0Uv9U0cJp81Qb4poGQrjMS7fIR90s/YuEfb0Y5YlWlfaj7vqZNeothYgp
sYN1pDs//AVVVW45qG+sMpvpUyACgVbFhYiJ6lmHkM9WqvbP4duGPg/cwXie9+48RZXX71y1tSCE
EYeY7Qfo1mqAEfRaMJDJSUHTPfbNTAxyd2FoGRdZ0e98CYcDJAEzBSFKDmxbCUmUq8pS5T7o99U+
7JCX8UJpEPqs3mYKXxXxIkanf9LwOlpfewGRzJb/TJo7FWaa/yYP4uOpNnFaLF+EFgkLPysCD4Tz
BzdeeSDL5wBRUM/YutAxxRmoPq3JhrpBeLkleIzbcI6J9qveveDSYFAx4TxpSK4bm8IEGQkwnbgM
+NmE6IMh9JxoydM2ji/iIW2fgz+mnd9FARxU/fmxOm5OHS5GBXhzxAOh6mu4UphPPkhMxUZrARf5
BtJcfsUbJxf3mFv0Myin2ovYrsFXW9aWuE8VHEz3elZcYxqItgC2H68oSRlfeFnswSAP17m/h0yC
Dw+z49y/pk5UB3vo4TBRRHqqx8c107bRChGnWE2E0n7SbShreHDIpaSSR+ASrZeDLIq3ScitE48M
Fua6CqO6hlA7P4Hp02blar1lRZm/2veHUeaKXSIuDRwF8GYh6KZE+N73Lrd19I8SeeGhW3G6H8Nt
pb39wHBUg1YH9oeAfNdHQOOFUELCNRsGhdSpPQcE1FDl8ygL11EeFIGechydVBokvs+TXdLThG55
mfxQ4Gss5waedw7gQHPzSF1+Q9r+0BrXEhOOKFGLpB8yS0hE+iaVXwriyXxNINh/isDMJS+bH+FY
rQsb5i9z81br5VPTQLkp/IMYmRnkdEkqjh0b/1lIQ18XPwXJq0ai88HF074jaNvXiXcrKgAx9jfP
T7t56LfnNQ+O38iJv7ORp+v298dWzzb033m26q3tuIOTcK4jFY9plLUT6BFZRtiTyh5Gu42Flx+r
nqwzqgTYT492yxUU1/xohqSXdEfDdp6a4dO1qBqa23gf3SGUryb06/SO+cQwilDCF1/TgFExWxHB
GEzLWyxK0lD3G+fHcisrbtvkOTJNiZ6t6oxnonk84NMtAoWkyrZ9/6BVS88LTyFGIjmI/0+ei13B
jUuwJpvrNWqjNrAJNDYwLOIxXwa9+6oaFmP+gwva/XFA10+GtUtfMaXTq+ic4HIWkLsEeJYaRj1e
vaYgPwlATpgDjQRS0R5H+maNBtod+csMQ3UPKJVCyHaZMMG0YLQSFKEGET7B74NjwYqWWakrZjNv
I1F7iMc4J7iJSmKlOhRbsJ/sI/AOSZwpZa9Kisq/usJR1beIKxi4gaDy6wAa2CWV92AMm8wOWs7X
CJshBVPIcvMR6kx5n4vbw6yQ6f/9sFkp0pljPXmOkpGFO4r4xuXaJNzzVlGuj76bq3cIBugIt8ay
0YKSBJndKUEzApzoTYHNs4gX2Hcmki5wEIyOfNmLZSatV610Jk9/PRC0GfeF1jyU50oCMYohlUdj
GkjHavWIOdsxh2Sw7pwAMRH0KVDZOePxPdBiOJC5k9JfVfhzBbfhbFGdYJDolts4sAxX4lKl9qYo
gPiUIk0ED4CFioAZTJyQMbF1TKs96nqcceMQL3dxFtQUDI0Jw8kUlnCE91PqBeYUae0KSn+ZTPZa
ybT73eQZzxSXv9uu/WtFimKXIw2A6IrtaTK00NiXiqUOkLb4Dy/m7atXbLmh2KHjCKltv2rzGaDM
zTI+/l+hOjS8o2JjzkdJ+fFrBC7cGF5fY2BeO3iJQWQezMiMWX+kKA8U4DmbeyMSbS5PVwIZJTV7
z9uAGsPcVUbYH8H4+TQbWaOW/xlbvlWIm5hVaHVEdKnXQgEfvVsrgFMBWZQtdk5x313StQDSKLw8
VmtyQ8fZKnjkSt8VJuHfZUNXOWgEtpl4M8bTjkQ6GUUnVXK6Lb2FI3EcWlIVhtBm8rtGB9W7kEsj
PM0Y+KOgBL6ZwtMcz8nIdDAoICSTbNG8W7vr6q+hb+K9lmI5DLVEBdRo1Z2qNW83UAw5gj/fD01f
eVmBtX8yYnhF+veDpRYdziGMrOngAOg2z/8iQPuH6+Z6AinOm4hFvmKE/XcH0Dqr4RAm7Mz8lcf9
QdCD2NYFeePh8tzeK3u2GaeMeo0PsGkmpU/z2nEl99ZPzrBD2lnpj50C4l92iFmgHE0inQbBElqI
ukFRljQXthprk9kuVkp28KXdjHu3/GKC4N9dlpnY4Hc3/u/uQAkinoP7xhFEmk826Nj5vR80kBTi
WHV78++ZiB9vJlh+0aJV/t5/S7OOJwqwHqXq3h5PcyIYUsKS7r73xQxJdxmiRptbG3WEyi8D5MO5
iV6nfhJW6mm1awcWRLjbLGuDcmLk4Npj0fR1Mkd6tG/9WtC+gsdLIo5S6NJYwqLnznMEpMFsIcRk
ZqI4M16XHYsBQZiPqICs0YYs7oWQ6M7DQfeD+vYooFaWouyWCQWOAVRzjMbJoD5KAA0UoNECD+hZ
1lTjiAG+oe4kotWW1F+mwyz38mDX0MW/V4rRBxFAe6fDcvYARvZ00SEXkXwiExDeD9Kt3uIJ4niW
Nhrk+Z9go6dYOxlk63UVpy5tgRawTb5kYngJsP/9mWwOoVKr9e530ZLZOM9PbJIaCFRIELHqw3uh
sMiES6B6zMcNQRlIL0sdhwwwmabWzNc95l8WHmtCrAHP7budkZAUTHzRdRc6H2+2/g2iROvCmZUf
hD3BFkAeRqUwdGRIW9a+YMg3gvIS4xz6MpxZ/m8OYJghU2i67lr52yXKfkLpt+xiBptePg4vZnks
ZyfVYrNyvN6aqADDufqbnYq1umbAUMVBkh8L/YkPKIbaeRm6bQC2/qvvYUT5EBgs/s1jX/ra5hiJ
Z8rkNsRbv1Syy+QbKm0NAlz7ssvWSBzUnKP+3FRa6YADsijpFdESdxbjg+beOO/bs4EeYARKwNyX
JEwnyl7N256XfARRrFpNmaiYkU5P/kuj/iKvEeuXMoYC0ZWD1QBBxHq939mFJK3scBynNl2IproH
Dv5BjNDTpZIhGyehSDd7V2ivzoCDMaeM8ooINYbfR7U2HKydj13qIhGYaBPa35EAF+iJDOkoeq58
zG+8VG1Mm/ZsdNgWpLfFqd+0HOVsNWiAam+DuWRyPeU3fq5/Lf9qFQHnUbNZEO17XyPXSMr2BseM
6ClKcYD/qezWiw4w0uBrm5fSav2agtsm8E+Fuax98gyE7HU5DXZassqZITWPkt4ZXYdFx7Wrn8K/
TICuLQQpRHyw/8Nn2okimYI2olnpGknnMRAoe4q+KUP76mcEPKMBEhSm7EmSb6rgJ8BXASj4Q3bv
qzXukWtD5rzmJWdo/to3rfMiX677BbGFrwZdJt+0+1lBKcFguAQ7EX4+3aRwrwfcrze9aoG4FrG8
6inJAtKETOW3NkZKUyuUf/Afm6KrXtljG7lqj6TuKTtFnmSFCj1U1g+mQAepMjxQXGitNrAbZ9mz
NkQnJkSC3rgvjxxcszoqrHnC5isby3X00TERjY8GgBfVIVbR251wEC4oRPB+giwhVUyyt1vjb6Da
PlTvyEPYRwzHdnGBVSkJMoqoWVD+IIYP4QOOHOxtSS+l52LE9HlYwKpcVko9oy/EonIgmtWri3BW
hls+Mt0f1N5ma5Y+u1JE4yDuglGp+yVmo8X8oqruBOuika4Ecayr2tE72w0NOSMrj7VvRboSt6MB
VT0FggaRaSwxSDtE3YfFMA1v6faUGeesw0l4BFLHXYpUgZOXIxmycNe1bQA3Ii2UV5YIIpKWD6IK
vnC7+khb5DIZaGyjeDl7Z2JPO86ex5b2Ytep72bxS0eR4//tvtXSEp/E68kQQmhLxsU+aSaQwUj5
D8Lgqgw1pEcQt4s1EYcUtNhqDJ36qp+GgGcQX28S0h+cgi94tvLR6lZDaogs4ynMgR++mze9Zc57
nFIjvaCZ+Yqk9jlO3dgPjTUUrlkThc1NzkdVKtCGzMZr+NGOm4X4A2Z1nHRnT+XYfe4IgpDy/d4J
NwcVlxIChkBO4aOkd0nOhUWOQv0U381ImsoSrbO21FRpXftXLmgv27hOcnnsfqQBKYe1m8MdbaRq
p6ZZy4kgLjxSWsGhVGYDC9dQ3GeWRGSwhGKxZ+KuJQRx9GYZiPTy7ITP7zZh0Ux8w4dryEqeD7oL
6V1MlmC2A9Btp6UIfrnSY8SYsF+I6ExOHAL27z1fpz7E8jQdvQrYZIYz9j4wQdeV6C2TEWLyFDo/
/x5KX7YqEKw4GLICIi2+/HMmj1VFJhqQTxzXfCnysdL0Q4514SQGaeuHxE3QaRMuYfnpTh/rrhTM
DAcQ2P0UXUdDfQ6wAliuOWC9rySCCZfSEdb2yLR6UyKeMFek04dqcMZyjSv6iccYQ2cgPY3NjPsJ
EPmupcuD+q8f8Mry8dFEvnkyhj33+NW5J88sACNHbSoxa8E+mt0IpavDbTah+iryBjA+4/CXHsYR
LQteEahyRhpilvry4XD2e4qIN16UIxtP9tdZc9YIFl4pLQwkRiZaP5PwRs5hkZ+JNZNaRzCCYLsg
M5A52Saqzp/kVVq/1Z5oFWWwgcAoRf/mCA5+LlseTiHlNWIm+OjNKcGv2e6eWcNjVE25ZAo/SVM3
nPwad5MpD4WxC2DzTPLiWLK2LwAvvHu62A5tQNe8jSzHM8p70mE6ySK0oQ2Zc0VhU8YlbZ8hlqW5
r0Vd7dCpd5P2hGvhvrOBDsa8HUdJBUU7NIRgkIdWpiv6Ni/x6J/E5ETFY8iFjEAeVLI1DrH6Bxkk
tw9EhCD9VKiKqbsgpsB+HbsNxAepZUf+U0op+bcaUKXbIbgrzfo6Y1hmnyFuSfAKI1ONPNxR/1x6
/QbOcbh1Gr04RFThcqKsxrveBNrcvCCTzNiBaX1/NkRTLI+k5Hmj4HKjVflengzqX1Qm65LcbRzo
PwT7SOfj8flvLwbN1hwM9fwXujyuY/DEXBEeMQh8VFPdCC+lIdRtmwapVpc3ccmWnrF6TFI2cyNQ
+mfInyd5ylrWjoJAUpTm/9sNmHgDur9GojjZoboRcMfaa5jDdQTDq8kVvNo4pXGf4OrglbI43rvi
kwgjcQm2y/ezS7fdVuBBu+gezpAdEgIOl/5w1aadLs1tm+TeFg3A6ZXXGkWXCEDGtCmwLK+6OT2Q
AItwtKLwb+dxmiWCcOv9H4ehdA8aI6viRtgFProMZiD7ZQxEPpGuy+OoZEP/bCEgLEZ+u1OYhvgg
g9in8piZLsyV4oUCumBpjsqqu3tMDBnTI45CR8+Z/nOsI05tsd1rkHU+/Bwq1wv0aap35Vd+5C3w
H56mlZwh0KlqKaE0PoDG6soqtkWEmCvW34DzGIlHWty3uJbO3JHz7zwF8SFGy2H7J18sYk/OzegT
PY4uGs0+VRCoj/ciLasLygryrbcTLj9p1Ir6EHq8TjSjYs34iaEBFdhubSh6rFBr192+6zAgdCor
dihtWvyyIdzTjMg2fvJsks0IkWLF/6ARy2kP4ttf7a/hZJNj7229ROkIxCiHZRGfWz+dn2Nf0rwJ
SzUhc42jvA52c4jWaAzhA80RmGg7xYws1dvWKBP9m+H+8bTRcQhFFDTqSER76vfzk4C0fvxFR6bS
nuCxafA9qRNDRJHn2TbcOG3S+thlZRa8xzZXVCXZLiyadtdb9qd2L0GXnfaXL562z9lYAKASS7Ph
w5ypcBh3BjFlCrBATvw6nX0umQ4El9dc79zIYKzg73jqxM/urMg79P+2cSByQw7HiRgZJy4thkGz
taOD8yTr0bloNw3Xf3J0ZoZ+XqBENxWUPC857XqXkZJGuA/YPdCypJLxuUf2eSpmiJzoqwMj2KSy
xe3MRCstgurpYd4hrC4CpX0FQpB7h5FjxG4DClo8XYC4Jx8pzltOSjrXMc32Mlfb6MUEUo5l+Fwq
1Y0fG1Y1XZGQRbLjFeiQN6F6OlIhh01VICUdfOZu/XekMIjnOr2GMtPMVTsWvh4ZkqiNwScWsKs0
hGB9isT5dGF7rfE6m00x0fEisssWE7+aQcAVNujPx1954TIBA7DmKhqiIimmrvM1lKtYqSiBEYiX
E8RIzXLvu/uiW9+bNmh1HyGUT1RVbCimFUnS7r5e4UBIh5NfqjQ0EOntw5f3T77pQ/pcQLwkiuAl
pzTKGXK4UrUYdcGm/5bgwhkFf75CDEo2GXOFtOImDF2YDudD9J+tAVnXU6RPZ8D5lRDjTaR8sIqv
GEBTOS+tDIYFixj/RHoXXy6QiOoCF+IRFPWUJqyTbm2KpN8U6bbGxtqwch3eH0+bIz5e6tWaoX4C
V0eZQmg3tPFiWzuFQUCimVb5wlqcrB5kWTRjHK2o4fsGrM/9aPhr9nvOtjXji2v62RQ04h7lHKj7
EoNj6G2fk4A3eait4dtFk7/sdi+ha4+JCqbaoAgpu28QjajjaoI2+1otYrNIxjvDR2HZejfkC7NL
vnVKBIOdV9yKIopB0JxABciGkz07WtJiMIo9+ibYVVOzaDyaxSmsEBNlraLlsbyhKOKsCz7ZnT2T
WTVF+2R2EuVSg8/HPv/gi2H3uS2G6d9+mhcSDuMF81BPKKpjcq9gVsBy4tzFCQ2tl63GKb1XQYoa
5FyIRP08Jz7LT9uhttqSKhf1iIdwc6TRTHrexfiEeldGvFtOJAg/6r4Q5STo3PPGadMyLSdKIkzD
erjYsMou9mfGWxN2YksLznOh/i+u8Yem+6BmZSdXCqxVq/dbfw0AHft6XX59i4EJRWyavqLerlXg
e6F/sIdcEkjD+GY1NdrvraDG0WDlu0UdPiyxaFcbGSb65rrHErMh4Qd2SKxxAXNX5dnAlnWLAgre
MqweCNMuWgHPaHMhv7aC4tGmX3YZ0T/TEJaKZWNaTTsAqsIhmAMZLB+bmRKV7ZGlNWMTAEK7sAMt
v0RiOSWOvyqjAB0HZTblBMwTC58D4XddiGKKboUyN3drh9pYyHWlADOPxZ8wMGzcAt75sKTDfMWg
jxMnStLXVv7plgPE3JYbxoIUk5j4BltqYrC8yWnxW3UOxiaGWNwMXlTyS7GHZssBrGVU8DZ+FKcs
0/jHdHeXGsyfsczywSw1X5FWkVcMOkCQRqLv7wQ6afqar+2Bh1eDOYfsPl+sDnDAxzSrTk1xbjUM
NEFnX96IcrMmtkVQXxWwCCaZ5Y9Zng8wwnAQieDcW/Os526lglUhFC3Rk3cOP9Dm0vAH6/e054+5
yoYhEevHerafOLHEpynG2IXVxb28nN8jix60uzGrr8SSfzMtjWmWevzY39Gh6isMDWDBtTHaar4g
RrmDg7CdLrAVJXWQIy10rfs9++xYxG1FCBQ0ZNBDigTvFGMPXTz9U+kspr6e6SIQS+evOyK81ltX
QmbEGw4AzXyomTpjfuo+gS+xa42azAOjxPKwwUdRauYrkfZAVoNJfB4kG7JV7UVWGIQ6yK9yzyDt
LmAWn7ug7PXeeMV29PS1JDN1j3Y0xs2sqKdMrxxmrTSkjWi1qUvoCcGd75sZDcdJL54jqMjSpIho
d8sS2YWN06y4p4sLWRczSyDK5yfDPNVJzcmUNp6ogrzwGQJleNjfgdm+Bo/r3Blm89x8AUtjC6wt
/V+3XYymmfgsvklmmxeBGS1ve6cHcDEdXpFNqXZaKS42TzhRyxUEDrF4MZr+ic9oEZk9PEFa3p8f
HK0D3QcPrQrr82FJvpl5X5/F+xo0AexQY9GdDkbUKA2ojs0PXygbBAWJl8hEZrJLx5BE51Ew5uTz
Nd6Yj1VW++xcTw65fcC63FqzAqOyG0inyW2p080D2gMmFoZ2gEnnZYrD57Prbg1I2LURmikUOJpO
6EHsszgm/5SUoJzw51ngMgkdXuk3tIGftG8/HkNJf+Z/nocbCeDz2ymZVhLy2MrRT5mUhPGtKwbt
Y8LSWr54eu86kz0lYj//Cx3R9DRPAHE7c7YwSVzM9jsJwftrsmAu+HE/5MMwMaY3A5OuVOozgix3
XI6SXX2BuPrwT//B37fB7LCSivSQLzXjdY+wXN6jBCVDcxIvwk2zIjJztGZB5DWo72vtx4ncTJQx
kmugM5xZqTZ01wtqsg/NBPb9FsQgDZrYlCLC4Ud1eJHg4LykH0wHHkIMrzan0+0X5wDrfNCauF1O
V3127AGkZviUvi/byNtykUCrs5i+SXjJmWVhw35YHgrgZdCQ/o5n5dG46xW6UmTkx9COw4OFQIPs
pCMbdBf84TxR1V3Q0e+12YJJ66KRaqrHy+3BUSgT1sHpBZk7bpAIIa+d9NfU1VMdvkGR+iUvra2d
hWkhvpDieO/3rq8WqKAAWGIX9e+WytG65wzIBGZcXvpaCGxqXMyl9/d45vd9a0Kzlfp1Mc7VqGYP
a7PegfrShscBiGIliu2ewWjGdL/ibzLl95Oc7OdYbaWPp2vdVe5yo/Xi2DRToa6W7HnokiLMEfEy
7szmYjHjkTSy6YNFroLL1mlZEb6EYXX1D8Dqjp/P4CHDM0CtFq41ExFxncTLkI2xT91Gx59bQsgw
nE24hZAtp6s3ZPg4iwfQFYmWnGEQXzh93Nn3Grdl3zCdcWFPpn/XGh1nebDlKEO3dX9QAVsRp6Os
2+IxeJnoy67dtLpGudF15Xpli7nyei4MDtkTTyfuTOdhjtbSkg/6wVefaeTR2oVmR7ob9JLc5NCe
44lHgkUabXo1H8F9L+kOLpgr5I7bF6LMKiollMxEEXHg+h7F3W1IzTfzHx1GltgVRSRvYykFDG/D
EFKuPFFFQrLnX9rBzZ53RUhRJ0usxevfGZopnyJLzh0laMXkAYaLTqDNoymwo9GeitXlNXovp9Jz
YZjZysjxQpRHL7kWB5jwe/S/gkfj8aQoLxErwNXUqLkFUQ3Sz7BlEQRbpFJOqMppi0nS4+U6hssQ
g4neG3x+DFmJj5/F/a2cHPAAyEIYYscGzKbAKumiDBfO2OYCVbrLigkocGTuJghkPg19Ni+xGFEN
QBTPIhjP04gqsgXJ/wRuP4jhot+Wn90wdubAcbSyWb6uYbDIAwsboErW+qWcoSw1CO0Iks5WXvMP
2PVKDTW/GgDzxE8tGy9fW3TRrWclxXWOHQqbVK2ZnQAz+K6ut93R+FX6qMOLITsaTmSL39qqTNod
Tl/uwX0JdA635F0gzyPo+yc/LhxS4ky83HX2X4UrLSFeWPHD64Mek9YW45/zGY0e3mSiw/OQqJeh
ENoUhemNEkDOrVsxYzXgetXE6roEWhAwJwsk0adDLYQPZIeFuNaYzpumTsQTPHuZw78XcpqBjUGZ
kFbt6qNDoZ/fvpLkYcKvj5/0s86YVMRP0aZxhoj6Je1OpYblRj6jSngF31H0lVe82DjY8aMoCcCT
Vd92hphMIoqMGVkFstl2zhTLotXLCusJmDpKGwri7b530h95FbOBXuv7ODoAbL/OOeI4KDlNMN4D
HxKFouQH9xM3njTropJUSY+XylhlMsfMN8gUL3FGMci2DWX4xiOPqRM404+be+N6/gjNFy8XoRxI
41Ai3D23v8RGpODcMXNOMardUixbcmhOq6H618QC+CuX8nrpfqVAMGLSE6otwAo4dy1V0mmHISu9
s2cxzT08oq76ARHLzL1QBz9e93EArjThbtaopEit1oWRtJFuC3eZyN1Fn8F53I5AMSASEQkFe7xU
MGaOoDJHWVFUd9OBPfWXXi3rsaB7B1oQttuHmQ5lBpSD0lpMI3hQBHOB+6Qcq/NYgV7pwpys4s5u
8zaKxCGsZ7EnWP1FlaLjvQFn4zQ6Hvb6CEp2WfqlUet5638gP4ctnkddgMxMrHLVrWhFBMzvMR8O
E+qkXAvRpxKaA2d4DcM348y61tI3RirdznoErdP+UKl/J1HaGujs652IxdamGwL6r7OZE9WV+lDi
dkqj/y7XPpBAOnUE63xDLZyiALBdu0DqcqUTI3jybn94LK2Tdg3qr2w7b7IK6cTM7yi/UhGpVSj5
UGn5Si2HQ3ut4Ec3aJLNKXMEe10H84PbrO3Pem+WCMit+Ftf9IkFKJRM7E8k+wAwz9x47PeKgAQI
6Ddk/Xlh3jTH+5kJe7rV1ZGtDrcgdIfTON/to3InHGPLGFBzQ/n4GOY+ID3EtSc9v7QMTcE/OhnJ
Ad5dUggoF+74PTh4Sigi4EBw5ljj06ReBM7rQuXb0d5J3cldXFC8nliPeY14h7afsTixQhIObi6G
xOsp/ES6vC7+9dxPehXwCI4+LVcRxqvGfxtKoEIP3+LZwJ/huNNQ+y1ZA5HEm7DA2LNiXaqEmrQZ
csnd3vJ8X4I4JbpJHyE583Ap08IsJKGOotExMM9mJgyG4dtqPQcH8b6ig5Xs4qsO2AurCSa5Ei+j
Ecf9DjzD16HNqB/AxXix/NOzAqEd2ycQHY91ZqFud10Ln8ZFinSgwQtcPLiMiyGjgZDFmHLFrmEc
/O3Wgud1ohKLhjB0FdLnKVm6p0XD19b5XcB+QVKlniD2Dy5ziXjmlYJRfJS2gh26ILnnYlwK5sLT
V+mwfvE/CJiDsiMQP4kR0Q9FXSaXNa5qXlw+S30g/qFbyCWwLxkIYrXQzXb7I2qQ72jYKAaVM3AH
0YTUvt/H/C9pyI2Lz+kC01mQOuQYPkY2sUXzETaayRZbhfxuXsa3P2z7eNSSPvHG351Pbi/3nxlT
wuPT6hU1Jb7mPJoLzZI2mhQJPszwLimSUX7BtZUbM1rkBOZGU2gxUJjoISSCqdSiXreiGM5yJa7W
OrgR5lCydI0lCWNtXLEZbIK7Qym4oaMozXuTfXBu9Fe//vMWrXM8D23bhNFqeN3160+wXjo2QW8t
p58+I+A9B0qM+qc7eLkpgXYQBUTvSr73UFGk92tFIl40nrl5vivl5Kg+92WJbxhZrSXurtfmyFoh
3B8ArgsthZyuYZJMYglBvcMjPz4HmngKOC1SkvCyEcpZKy9H/AgA+F1dCh7Hzxs1cL7U++FZjB5k
OBlXpNbVToSUoPKx9zcRF4do9OG0hfrbiU1jLozmnjKBrTto/p+BQBg2oW9j5jlG6JZ0EmS17lKQ
XPq+GhjxaqScJaEznr2Bm9PAxrURUs6le3AqGFenzGyH3TmYNI4vjxu4mjqgbtglb9sQ10GQU/2x
SvQ77LGh6GIpkRrXtlHR2mGLLy/TSwB7YLt92f+QYTozyWatCdgZPWXskSQXiAXPIgckkKgmXxzd
pVVFz8Jy8WvDzOGGkkCTPovA29MPO1QH/+VVT5Frv/2EEa1enmGD2qOrV32xMfVmuuF40RwRaAIp
C/AJQXpPzIC2fJ5gE/R7sBSCunCDFLkLk2S8Zye9gJ6kGSMUL7y5dPioHdfi+KTFId+f+Pd985Pu
OmvonWni90jp4Y04l9Z8s8CINd/rFeBXFb1UMMZhQRNcOLeogQ2v/A5lItK5FnMcu5aVZYDbqUbr
6y7Ldn2ogI3/1qXtXte8BzR+BIeN/hM6zwPOsvzW5X0bfLlxIMhL4U6+49yHsKABvihoilIumGRC
lK8S6+j3xbX7bAcHEzbzgcMusLqmghoLtv1gNm+EeqLC7L4PdG3tuhE3NLb7hBJARCqjVFh/S8ix
RLI91njCFC41DqEPKHoR6rWw8afKG/R227SQBYoS5cMAwC7qa82DsL80JJUS55Q5NbZv4isOHd1P
p3AKNXAvoM7o/z9Q7dDfe4bQw8egf1XWoT2stdRwJnYKPafoL3uE5chIrnK5P5j6OpVBIijzSbB4
zvYZKQHwXgx2qnO1gQsq+o36Jh+w5LZ+mL422qK2yq3MBdwLEG++yo7fKy56d4ov4MwadNzLIdoK
Wylb5UXAoFA65qZsPr/C/ktSjLX/JDBugi1w1h+RUEb2CqGwe7R73SJSzIG8iI5+bmfQns9CIBJK
StEEVc7JneKtrmncQsSm7zMSoTDYy/gM3C6saZUCCsjXsrc/INxXhy2Kmm1LY2021leOEf5K6smM
90hE5a1X4/e0fvCtPkBRr7kOTPdbvfl5S0Zbt+8NcadivEDQnDoYmbo4Wjvkbiuo6ZF9bmqGeFI1
0NPt/jqk/4AllamtPBcNc/1x7lpyrWk7l3wez4uzJ1WOWvviZ2IO5u5/8lOCf5jkTQH6eVKiBkkS
39XO5hhwUKTREGDx5I7QKuCZn9i7suGnwOng5JWrsHF6b0u53aDjVG+wiiY2+VwJnyDMZLZvrWwq
nTWd7m8Q8ZxPoUilXYXd/qVm8UWcV4c0TYaHxkeayFQA3crQnYb8/6V8PPwGk0js/y7YOmZzvk/s
VTQJlQaNwJRDiZD/TrXWCbJ/pyp64c6YMZrs0UJkq65vmQ0s4A8i1EXZgaELM+O5jy3sBwZ/F/n7
aMuMayZvIfXd4Dl2xZxCn06frP/glLWySEtMhvYfspiVugU2J/zlYwcSCyR01dRQjpn8Q3jaHVyi
c0fbtGikFYnGe+NBANCJqqEh7BxV4FiGRAXqcrW+BahICf31PoZ3buLF9sUgE74AxTMiMSs3Z6R5
+g+Ss9fh1fg1a6y/DnJNwfE22fy4+dPeJTBJ5SGPQRSFUqY/9ZuUNEGyDCvYCH2SfRFJFIlQLrbg
GzzIMZMHqUXtmwp+ZzhZ/lqzmgS4lufR192LS/dda4VEeLKRFwLfp/yT0hVj2Htzc1nEvHE05hLp
j/I+6Ihs+m6l5NndpyvPJitbB0j3yBHHHGqT9Ev2Aq2qqdbtuOQ6xhO1jcnx4JZj+EyXbJsrYwfk
MwlPq3f2W2s/aL2TMLm9OQAM84wlhJSxA5kMzGJHI4w5jsDgkuPKho1W1vrwqdC+a31qiekAyk4X
ZvQ0GpkJy4X46Cp5C3a1qEKXYVyXDGPI40Fa6QDqqmPUMtkm6333URBDvP50lCrYkUmccSPV/ppC
Rx0OWMPeNOzQyvOanfQKeeLFIeURRjgTBuRyq97KkU7SZ4e39I/cd0xNruly+0jKtRCWSXwG+1hE
bnT0VlYAVkaKmWXn2f0OOxWtqxXOtsJORF9PdTX2YExYfR6TIAXG92a77KkurOKOtkzmvZE+4HvV
DKfIwgabTGPsRq30vpCsVYL52gzvaimsR/L9mS+AAr1+uIaHVu/16RxDYefUjRFFt/rttfn76b+s
SCEQqv0+CxSgc4gTlaAI68KKj83lW+/x2t+AS1XRDmFXfAUpOM4C5GuCsfXnCXlFnzr7IEkhPTPm
IDbdpocAi4GQw4h7/bP7PkGVgXUAk2TtKLfdy9uhBNwrnyGeMNvG6OVToKHyjqpA91yLEuE90Mqv
EWAU3DpKWUS1Y5qVg0crSrvv+qzQoGixA8EMuvCiqnN8oJsIyjh72ewBd5c1I4pSEu0Ywg5slZZs
Cv50QLnCJ8RFn7kHymIuSDVQYeG3dTyxNF0HbcimuGMAo07jjnZUASVKRUMbAdLh7RPFneoRG4Cj
grpP/3SY8L9k23o8FkA9EmpuzCOZV0SlaqTacTpL6aDJjyeSVGTGIx5X61A9l+CGSy1du0Ipiaie
5SWiOUpzMz2ZbUuG9T6l1E2J08ZPEWrwqP1YYLGZJ6eNnI40qhWjryIw/7Hpxmg4R72+TgItEk2d
IAhhfMbZphnp4Lgo5z5au2XP2cu8FbNsxVeY5NBGsEui237VAP0AW1qZcq3QBC+NKwV+czqhmdGl
l8Wuaiq8//LmWRA6T//SBxI/oP22aLGVGAFjWaxpXoNXVZV8q0EpksRBnA/0C4wr9w94H1mqccUL
Pdwx5eAf+1GzRujFgW1zbTsYEZpoNAbudiSIh09y4V6LuMsJndl1yK2m/LtgGT9k8VM0CcvaVtBA
ELaoIh3Qu2wUiZAqGrG1YcmtvI/Ag1DW1v2sQ/vPpYcjMVpg8BKurOlR30DPCuqXU7M1zHWlIbpu
Pi7VzkUlc8UKrxaqdMHOIphQ6YzrXViRRW5X0t96HAPHk4XgY/RkHH/bkcOMwl+jp9EShprDEF5Z
bCSM6HM1by1/8AuTsSYbpfmSKy+WFi3y7kLOocECTMOMHdwXRdL3mu7ggKhil6ij11kHZ/bJvHWW
HV/KPqbUwkm63rPzWqZSIEtApqSTHFXKRgtlKrV2Ruuxr66cLYwl5v5rV5A5djnvvYNw9rtXsIW7
DI1ajkmEO1eQDRnwmXV+ujV2pQ2+yYkDqg1mbYHo92FcV0xP7jYr1zGNREmKS9WKSQN0+URNVZDU
CnpjrYS///ETaUj2pkXiEbUT0aLt6jGGMIJTiSL0dC1MyBSWCFYNlHBib4nB8meyHIR/7KB1h5PM
/u4fSAUCGMsm6tiCN+lwgMjSeXfaNtdB+xKukSxJdZq9z6Hwo7qMsgQYXLJQ3w/27YukBqnSfT7M
2eRRSYSAABn3vAASSVYMN8a5/DXfQUypD8A3D3ZiXGLKPSHW/0jw1E1cqESWa/hjdAuz8T/zfY7x
rYfmZhbMncSGyihkUdDNA7MEH/AzzUAB/PQqy9hXsCXok1BLgOs/uKmJnci37SwgOk49Z9OHGISV
s0OqggTvxEV26qOVEb+f9PXHQ/DnUM6HeaRkddTQ9CuLaMZE/m6fnHHCPr8qbqIpS3+vZFBodZlb
pdZyadtUPQyQlfKdNztC2XmrRX3yrZirYCQduWmaq9bNf44BSYVcxN9xQdxVpljrOlb9hNp/vCpC
z10hq21sY1A5orUYp2XnvENwK6kGZRf1seZwarMTMUImdnbv7hB0jHnFTgBL1pTHXxRWKSNA6z7t
yzHuiSJsyySmFxBkRKgPuX8q6ywUoLpq7p2ibQSMzm1Jds0yfb6Lby7Po7B0n4pqQSdaOaS6Cbf0
iDVo56pElIH44pQrM+PYRNbVsTKm59p+AdSVvEWpyPWC8V/iJYyIW9Wk/5IAyeuqCDjmdkh66xKb
W672VKTnvmgdypmNa7AkKzrc+j2epf2D3EwgiMExxBeVLPNIVURc0UM4Syh9LF/S1gEwd8mulHf7
g4P9FZQJki4asjd6+YYz+LdW4PIrSBvgDHW50HAOvUGu3z4ZpGFPl/tdTTAe1Y8SVp6juA4fsD2Q
jABntLmD2NB7+M/FzPtFXKpL99irAltSUHGPaMbqjTz3XyttNJ32FXqinQBcR4Luo07cmAeri0Ta
ulHSNRKT98aIPx4HZKw3VaWVaw9Z+waazgawGDFE6huqVNei4brsHGq6rlwmQXIawOrJIkYu04Dv
8iL7ne8izm+LuJuFH/GbTc1Lk6l2/E1RrqJUeRoz7Xbq/VPSSlUTYU4gveiJ0Un5OlGxjceb28jt
MCawx+l/pLJX1hTpUdOeSiAlKN/XeJ5JWvzzvqfVIN2nmyI6roj5AlghbH8MTTxD/MHCD163PePJ
Fgwf9z1vCTRQqMJdyS+ElOlM2cLG8/Tqd6ZTh31mfT0/9UMnlsg2Js+pJD1fdqQzyQy5wqv0Pq86
zf0675CfFg5fPGbZTZvP5MLWbyPjBgKM0w7KWj0wcinxNpc/+nYOw+re/aunVHp6I1J/2BVNr1Tj
DnWvPQmHy6oxNFcrUkGt4UW72LkKmTKiD3HwBWzxox3kbk5HPEzDSjKFAUuEFm/jZHMQYl8NkcHn
kEwqTpluaMdO/4cdLfnZsYSwXGAi6EwlFLAb/AqQg5ZB9cSQrq63DdLD2l7LR4oY2m5f43KrxIr4
8pc31tFTQeTTIN2D1yKJVOrSNb9RE97SgZVrDHWcm3Xx1tvxfefd6SiTY5DEZ8jlF6RgfCd+AwKN
SgZQIJj1gkxtDLtfX4RoGIOwN4DidsSJkKDkRSfXTsHB30WB1pvYFoT4Tq7Qfg4jVIkHDqVA6fKC
wTi0wiAngFBbLbQUHArvK0wVpFqnRg0n/GqbjYIojZJQr2yo2KTIhfM0rHlR2Wb77fxGX6wkPyp4
qB8EhuEhUXXNzdbA7onKKI/6xqWGFVQavVOCIx6WYOZ7cvCYkeeTsvaxtj4gworhTUvHiRXUZoyg
pLgZywv1vlxVvmT7cdk/3PjnUKebPG60aEWs9vSA/vU6ZLu4V3MAsnbCS8TD/PX7GzVYD5urqV1c
eH9pJZNr6dqH38iK21cnL5X3kcjaUFtLhN0VpQ4KPOk4MrxJCVIN+DLiwmgEkSbt79x4wUd73CSN
5yXPUkGX0T+MW3GyUCudakdMyAzpMX6ETbeDmsAd9WEMZkCfTlRyA+CE3DlXb+KV7hMjWmCc6bvq
+kSKExnPAIcZEC9R9c3BcnE/hGyLLDUjPS18o+nprjrsctABv8Y8PjECO79Z8fnsCdt2lVi2Vhn1
FvO2vrs8f4uCZkpHG6uvz04HUcrMnIceQGx8rzkuKZ4Loa/0vl6uFlunrTO0HdkRMgKgnyywdEkK
6/u30PeWh4zoV9CwwURxomcKIxhYtUcnz+VXgwbFhn9ATwyuf98YLtpzLgl/3FryqPUjthyLdFE1
hywzUqzdnIjj6zDnbU700Xhl/2rkYKzbT6crDgrgMJ/l6Fl4mHF0IeR/0vdsRXTG7PU2zol1Wwz1
Z8UCQvTf2Qrteu/CZj0eIuwRcQHhUJxviJihm9EOK3ukVYHm1nfVyrn4FUMWAqCiqJKBIV6xZD1t
wJ1hTnfX5LaD5ftfe4K3PFpMxnKC6iWx3LubvxnrKKSesAeFQp4iUZNh7GWSI3lbL0oNUNxzjg6i
4MmGIdQf42F/nGgcMRdJ4r01RxSb0qT4Yv8rUXPwHM0GWe8Ght8iWrCRjMYPWlRhBzybjCbbz0VX
5PT5WFUELE88uxeDa1DadpLSKZ0HcZshTZuBTElhCaAHc927PoVyTwL1H3o0hKYhaQy3UNEQQOwS
mfuNoqoaUcWhMdNxlfY0PJ2N6WWZmi3B0a5AlYngizASEwjDctqGlG3oyvGSSEF+ANgsUmgcaC2g
uOb1AZ3Ldxo9wPFP60ACWareUlruT7VPJR23UGzkGqxelfQtolOMVhOssLwocGrE1XRJ+DMGIxK2
kujwT0je7oOMRfXADjJaGn9I0tMoJ49dSVbDBkkkG/dV4sv26qtvEl1OHFv5SEWeaE/PUTuK9a/z
G10EI/WYx5zc5Cne/CRRrGnVFijHNmjKnWxeMpXwYnGCnrT17TgN8rir+aJrxVQAX/CKyxMSeFyn
oiN+X1ZdkK71LKmjdWlpChwgmoXLtD4QO6JKIMlRBbIF2D7otM/O9/pe9x0xuDMZpw9/Xgk/vP/F
CTxIJPwzJhl1P5/tdgQcT2BSdskKoZuh6eyfrQKP/9mjFDHh92lswPWrBG+56bzAOTg+xu5AVFHZ
UkJA5W7SHjyifP283wjdLajgC23t1P1gjdMtx48uOHujm5gcDAWnR8epbaJTTG4YfCZQmj14eji3
rR+nqRuERKytDkSUP2rfW4IUMH8eHeBWWX7cXq7XcIU+Fgm4RPcl6hueZQkHWfLvcL1zhrt2xjTp
cJQDp4TulDxtVM3wnrTM+Uka73OnZ0Lw3MqnL6WHc+/uHYm/NuR7bL0yEqzIfIJrs5maZkFDYkU7
CQi0WCNauAI3ukxzVQZA9+wBM+5fWwRQaX1hF7TJbIZJBgzz9P6bHy3GsjwvyrgVvM7OlFt59WFU
LUEf2rHzdf+kDLtzleRECZs/9UDp2j2x4SDUQO7HTRNU+JdpjWw4te5ZP6024aDe+h2IS7gviEOZ
J1GNCZYSmH8++q6gM8WC+8krhjlXUCrRhTMs7q4EiBxk6NAP0NLlQOyDGhlhDqZM0iQLBOhpvqOm
yUrL9lXPb9EZSPhhSBa7zGCGFjXk824MPvEa99mgeR2wM9hIWSw4WeTErpp+GIew5+F4jQCEBbWg
DpsKS3iiT4KWSRNW0ERSl3mPsVFGafsduT2FEJ3Yb6k3ZO9bFjQ4AnhpiJhjCrQZcNLh9ufTeXgd
xuOecrW/fTfOv0elvLX0PJDtxBnHX2HJ7Keswn6j/w/USJGExzP1sJVSNd8HIiSX+rcyK2MQD3L3
2rQSkkh3OrIUXyNWMfZByfzKrHIPM13rDJPypIBECYPQT8V86yM2mocog18Y5jFG12uFT2RQuRfw
zKDfarkKV+P/g6Wcrix8sxQfeaD9J5UkNPuf6nSlqmOaY0DtRDUO2u8B62EqcSoMY321LQP6qRJo
lpJK4DCIjjPUPX8th3B4MGnC8qGXrqRQTQZy1T18CHLOhKg3JtcB/AdvmN1sEzSYoF5mjzpL1vlQ
wLQZ7FCXDiENjIqO2tKleTRnVg7YOhC02DAJtEh/aeiXnNuMusrNcn7Lp1SDAqrwHa8ZS2aiWaDP
MJoyyRvMysrcUED+aCqpQoYDa09qTuOODst24pxBybAueRCqDjbn0IfdTfAX8hCLIRrB8wj7eHKp
Cr9znknd5o6CK17CyDdxcedHb+VxJAxzx5SMRqKv4eFXf/OdHRuApF/DNGDfwfSxjP4G8fnqUUAZ
DhqHGaHTe+ojDGwuH4qweEmDcsJHt48p7+LpDq+fBZrNKJuAQ3fYeC/9Y0yRjeoDg7i0amkSOdFA
8FFagdL6I7YqJyEmUc66nZ2KFHaE8Dqw2zlKZzrYxlkYFnRgTpCGNQFTz5W6Ab4hbZM6nxaga/V+
KjTDzYGHvtTs+KhAWBDeSBapjMrRa/zMgh0RwZ64itJ9SmQGabkpGdHzpa9s42Ql8rYMseRkona8
AHByup87j3IcwoT5cwKY48DGa+WoFDHzh9hWlEo0KtD9Q5+EVmdFOFN3QE9YxO+QP+Hb/gbg6Ynw
2IGgJ9Yg6PXIcgWcAOo6vv9pGnHRJCzEIuyznfAIjdzefYZHj0vdq2kYxx08y3O+rV7WeE/LjyOI
0IhtqrkForjdHAPErlJfV1RW6FdfYCZpYidQXXcINvEHELKSnq2vNBNuDTOE+vzbGRJ+/pK7wWWT
Wpp+ZHngufA/YlcdzBeNYoZCaVRzqllQGGf8XONjv80opub2/3XHjE98QkUMSmAWe4mvbs+PJObR
E/+8yaR7VGIBv7JUxYkde8f9WE24SuNzXQ1dDZFP0y2ufB7MXWMZ7w52pzEfYv6RyoQdrCK3VNHr
UIj651ODtIPiHmKSMQ26gjEhuAulfqW/uFgJ13/cBn2/jtom44EC9tYPSPFgHhq88+Ylg6tS9IwP
GMTqV318el3FA3tvp3k74G8Q9tzKZdNVKfcq7EVoPO1gfjqzhgXXoDcjaOmvwh4FIMa6okXaurai
+hkCFWaAVYhMLTVxQwFRekzg+35+vQBIFwFEvVM5vd9liBE9yagb8Xop5/p8KmrqaeCAjtsPD+Bx
8kulscXhTj+O4YrdvLSYweFsJDH+xk8e3ebzPMCNwdXMAkisThUEdGxv69M0fTd6AzCAY0zkUd1S
pQzVnuZH4UYxkMNj9VimyqB5MtHWsPaKI71b6ZdyZeasWBtZsOD7Rs/Q4vhqEe4Ab7rhH419dncg
z0EkACrIkqgF4D03bkxtou+EWsfBNazlW9C7ekcR3+BpgkFvd9nJLU+rqquoOYLrFsJ2CH8ipwQK
Jl7fYoSmeR7uYlb0z14GjRbWAVGAN0KP7NlmLGjCIEAeiSuEzASmSmw2AqePUX5cpMIkJ4iqHCnI
cutB4NX27blkZIvdkp1A9x1Pb7D3vU0iU0o7k49rIYPi0WisdsU7TiXtpBPb9rXTsmoLE+6MR0pF
uTIMh5AJdxsSQhW6bY1To+qwoNTmVJq87pGPitqmZa15wX8WMsteRzQfocJCd3t0y9UWNjwDQw28
Z3T767LFyWzNVdrrRMIb4Vjc3IkJTBfQVBVh1UUkDBOWdghmEjnksGciGrU7IkK/wYmvoLEEPiRw
rzxJIfa/PsuaUlHS4u7AlJkDA5cZuDyjErziIn3n/yMTpUHUg8x5Bz/Rys9GZ+wX5cZaJJFACJqZ
OthuFf+X7wikFcn5H1mpzlP3Q9jzsN+qh4nPGOSQlwvLpdVtneyMOGLWqmiFUbdrBZpv8MLmgieA
0JGp3z3Ffg7cDWK2Pa8l9N/rEXQ3ykkae6LgO6J8WDv5ynT8fXj7nDCn4t3+JOtZsLn1YXPYBKN7
Vl1DzXaB4jgWsdKcJ7pPjyyd6RyfL77npsHlM7ddCS0EmlLToXX2zyhwp+vNU0Oik95E2PzOoe62
OFgsZYvmEWp9CgKWJ9lZwehTuNPAshpFelUBj1H2L0dyf9qXVpooodTwy89nzOuyJL9W0gCOSU77
Rq0os73h1qEhtCMEp1wcLoRcBdTr87b6k0PRk3RR4m82jj/0ma7Z3v1xd23JCUxAmokfP7xt/03q
mMPN9YgyFZ/8n+QyBHJCvGsKboutwseEqvm7zz5zEXxz4FZhGqB5atUvP/4J8FbQTTUZel4zLMki
gcVi9RXbqcmujJ7bAy5GEfFQzQTWaO9iqQRacxIeV00tNAGdsiew5Th+ps4EO8ZT7NBoayBq2p82
JQQu6hz2YSUMvX9PvDTS8qzE/VIbEk2ZgYYXupQXGdTDVdHuiHy0gUpFaFFsrbn2pGUHWXNmcE1o
kd9GcJfWS05pDyU+9hMAD7YucnIL/FkgYZLSQwVfEpOp1oNi6TMtVWSapscStx+nrt7l/yfnov6Q
iHrkMwUqTyttIlrv3NI46MwddHqS+2vVF5ZYq/Gt47bjiUci7L5odk9UAQKa06S4y28/BGNWKMTe
BatY4U7ZqjAkm3yC5M9FB8D5p7YOwgf2O89IqxJEt6NLozlYjConDz3kfXLdMR462gAh15b0Drfg
pSVULRN40QUbmi5em3ilNF25402RAYXyVn8RjuJYE08L0+Fxewe+OaccLnb2KB5JIE1aQ4ag5kkG
6LaxyJ+ieH2w8DMMYMrJhH/xInPOPX8E6T9rKI5NLL93E65QTxH4sj5k/4c4XdysMsDy4aDBwCAW
43OkfRJsnXJH0Wpc7U5p2aTCPkjtWLuRTlnie8dkg/ygW3fgNABc8/s5R1C/Q0KXib0F56N7HzuU
JhCQi6QTbnYK8PKX0BIxzCEepu2/af41aGuWBx6jHNo/Y8odsvCzpJH3oYt4bkOCMxAqU8iogR2l
ZyRf/qSmIFC5sM7HNT/vQ7MUhfipEFrcENGeT0YWuJmZqroM9qlEdtAnhGFgJA0pMql2JB+habuc
4q5DRATKEnO0a9aE7FixV1nB8czAlubdcP8VyaSSMSGGwCFe9VnV7zhsSujqnJ9R26rh6yf/rbQA
49KbwMtWBVoZcc559mEscbGRZq1+Q020xswBGlwKWlSs9uf97O8g8GmhtPiSIseVtOcb83yommaH
Qygj+EONnW3fOCnlS26q6nEMp0Ibyp0zvLJPblyBCy8MPKkmPIkzSFfZz0V0lll0uEZQHnAHGc9Z
lCFWRmkospY9q4/Fs5KqAdVIOoIAjCGocRvcsYbMnDRtwyucwp4B5hGyc7S5pK3bmD78fdY5rh0D
+6M/DEr17W26Zi/QfGUUlnfjq9Oz71dEBp/OUl3WYSy4RvAZkyd5VTCUuzJu6T6sIJH5uFBlzjrg
leumtQQCq1W1oSBNDFYEOlJ980D+RLmFdMuKSaGk6m2gfwdcqmKtnrGfA/YhI5TKiFwZCI0bxScT
XlmnAfJIdRLwKrbmYaVm0zm2Lqx791MO0AxV5rnSBh7ZlSEb4OLkqjQKP6LA3sKoTG59QmGz9X7j
vClq/o00eyF+PqldXmRSxNQuNTGAQKCar9eUr0hV2xVIfG/IWpu0osSsyS4fmE71rm+4zrs2MyaJ
KT+g1WHbuK7gMwwTG8zHU7S2UBB1VIW70+IGIm47GbjBWLeFyAeWntYGyY5MGk2G8fnXKvjiVgoe
PjTG/PUZAeKlrH2MkfP3Xr0/wLTtJk3leA9PKxnK/A7HTyMIDaJgTzaureYKynlayo6+jrKnTa5f
hOlaGyS5cLFhMz4Qc2aV2w1I4ksp210GMv5WKV3jnj35pAaCjj4uLnyj8RoUgBa+lf4YMWxJam5P
mWu0ctEK6nRFoidaqD6lggUWKZCdMB5wAUp7BbCd0UtUPtkXba3KSkKufbkOjfi9wf7TbDaEXcS/
tpDVq/0f+r6AtFqKfa2S1owu0hSDu1Ir13uCPeo0FHqfZ+SyfDgzgIsXCkelscttI7gujPwmoQQ/
o4fah0SbYtapQW1vAkCfBeTuKYvt4GveQOe8XIAGFdmrtbHILzrXS5rPbwAexL/w214ME25hlX8M
1FjxWkWPrO9GSAA8Wh+gzpZ1qhafCzqYl2p2OSKqvpnrlr/kXnkveT0AiWgMOgtB156yuXvNXZ85
Sdb6aTMnQpeTG92rdfMWwpwLN2W6z3Apo2kxo0MM8t9E1ZeFrzptabHTTYeSLW9agCEmnFjmrgZQ
Z7h8zticBeU0gq9DZkpJ+jksOEhgcyL+vK1tLsfpUQfKQ1nYU/mtLUR7FjTFbnVyatoEvVgz0FYT
w+fQVt03TQTugtqXjKUhXbH8b9YIzBB7KO3i8J6604yC/LkMzrARomOgaf/rD4YDsvCwowVrbLzc
+/6rKcA7ZRsUMfSAh9YzEms4oFkFRmyz+oQzDjlDkDpx1O4ECnFNebqRCwLFmRRTpHcbdGrdrNLq
fEhaL6+g8RSCVl3jQ4T7jjW6+s6qXAlsCT3xKn0Rv9fJQa83JFEQ8HTuVwF+cf7cjYT48L7E1ikD
402htwo/aRH0KSXr5/NuZdyN+HLl2J9MqTG4RzzU5P+mL+rGCvDZgwGnVmZk4iQUEZwlmD+qEq8U
lsUjkIIKjn/NwmNBDWQ4irqZkZhYAQgkqb4Lu20rtSH3oqvKijR0gnsMJ0k+CMdKI6mcg3ATcqiG
wYolt9fgmffLTyHDgQWmFH0sZpiCdZTQYvCRyP7V43LSJ282cAawUcxJTntdYWwBW48tzz3JVV1L
pWNJJLHw7Uq11gP6pQUVDkSTHyz9rYMn8AI0SZmvC+umEuVWQDLeLjW3YNVdn7p//XFmsrPHLG4w
cO9BaAwoxZHa5VkBR5jkbOZMbmCvIMp66jZ8gnvusiOnM1U0Xm0rK4hjRSj9B4Q53HvHuz6JwG6v
HCScIHIJGchCwmg0iALtXjMf2ZMdVo/rF5CWaHNkGndir16ZWYGsmi/lNYIR7UIP7LHxU2rRVhFH
8r4pUmfWNXlCBtP8jcqtc3GELeDNxoM7n1jIn1fNbiysGLsF7V2mf+YcwRCTeUfuR4f8guyNlBIE
rVf2aXcs0xs1NPvfXFxcVGgX54P6+dIYUT3cYfEL2J/wLETV1kbQ1yc9qBHvt3/LUSS9ayborJLF
mcmb1sQ9x7vIQlQtLfmo/IR5mIY+/v8/3RGGLyhGjKFG2l2wN1GbY9VjC/m6Q4ahIpVWtKVR7iqj
aPtaV2OouzZZWA5D0heNuf4D9LS7Y1q31T7Lo1chqo3dFTQ/kf6PHhx9Tr4R03npuitWWlqgrC3w
draTdT4Q46S8gtP0dzEWrbuvf+7Clx1ksPS56F3lZherR+K+/C84YVC3dCJA8iSeTFQPK+JpHim1
KTzMECRJcd9xbPkasDpM8wEesXFdoMxMJn2NZEAHKV9kQH7wG1irA9Q+xMgc1z9RVc1EQjeFyZAZ
lpLC31wVHnwlId7BC58G2G2PS0XMxkOUpqMOthj43mR6ciwlR62fQyTKn0uK/IuV1jViQML0BO4e
MXzmC10QUbOj1LHT3m1G00/U0mtu8F93hhfAxc4e0dHTgnJYeVB7Uhoq4nwv2EvKhEZ32WMWKHKG
d/mh18bJt/MfIbEaugwxTOWCJttXkvWGhxEihPDn6B9AB13/Hn0ov26VwURxlyZbzWvbTLwZ02oR
7dG+78Rx4Wi22wEEKZLA6n9cT/1D9eNsUg6edlxCeg1lu8Wsw4LOHKh6aMvJ7swR3EUkvUpyiz7i
r9JDHiqHRBXexJ1bVqXumlrf/SkDd1RhCE+MLK+i+fdc4gCZ7ow0+tALFsixIML4uIqely2sM51p
5ILAZ0m0Md+wPS8U5inRtoj23EchVWg8+Iy6knPuJdfh2saMfIsrwh+Cw0XbfKA51De88g/wgbB2
+7R3UbdPfiJk9DfORNGXjrZEI8cpoEfPWNsO5VjEG0d1yHULV6tkQiixdN7TnC6te9cycxB4LsXc
YmXO9RU9ZNzT/3XFwZ7fTkcktxeHWHLyQWXmNqSrDxvRzg4VEIiL4Gwezu12E6+5B7AWM3mrMi5b
Fl1h3LKIoEMYBsZiqyoB6ac7SYOPO6xrAfsQqVN6zrPRVP4MQu/ptbFwEk1u6DWeX94XkFgy835+
uvrV9WnIiVYMwYO+4xT/zVmUoFfY1YN+bYT+Q5tydSqCm4aidyZDl2D4FYbp7BLPefPbP8BLj0On
5DrEOk9fIpkbn3gw/TFjuhv9uJ4vHYbyw9MlgS1BX8fUBoWAkqhHhpuT+kjoFfRRnGRAZIuSKGbB
AcIPAPQPkkIr6tm6HMo8taGR4YNb/iVgygqbK3XxTEI84UtoXjNX6udqWv0iNX7Cmllchs/f+V8t
k1mMpgpDHsF/nEJRhFXlIXm8vDkiCWpp0UwyIR+flaolmZM4zmolTciE1rVAHbO+iO0QAc4Prk0m
UynEg1OknnvPnADaTbFi93NrnIHg9GCbrBDfbH+qsvmvi1f5I2IYDhWtfOw8iD5ynZA4P0zjNMSo
LjjFvXKxohdq9TK7rw4oeNJSzFegm8TzOaKi5Aqq05oJ/VLKfBw5mMPqkig/4C8Gaa1/MWFqExg/
YR+/P4baYU71OHQFnGZ5pJKpZQiYRtoA5c4wh3VYquOQKQKCX7Yk+YBIcDeto3usW0/ZgotbRTpO
9ae+sGcy10iTMGylh8sEvPKWPVjbaylwC5rIu3rEyANz5DpUwcbQjeVclK40yK2hoVuKBh6sv6bC
CT+WyYuIkskxC5fa5hSO2Q6oapcxYMH/olFckXivfmGgQP7aVCzHWSChI0AzA/7KmXf0kKagQwcs
GZs2E7ynlTdEH0FSlDaL90bEgYE3eMA6NuA0X2ea4uU6Nhe5JScZr3mY1gGQ8siMaLCohqtEBy24
P7ZDQrCSAMHUXnUkegjForli77S5VHov4EVzq98qjxBCznq8h6Jtbwulq4ip0zL6XSdO66dM3sgJ
tWu0ACUhQWlBy1UAO+jHh5Y1g0+e30Gz57jeYw77WOhg4bpLlVKQJ/+Jq6ddi+A/FDtbWbdBemkv
hML0jopjsA43cFr3Z8w1xdeWuOrcNCRia5UihdHuTFWgZcDGuNp9YFdu0u1lRK3bAMebfPv0dXGg
/UUTpdhrt4ZnHbAkMZwFJIX77qnToSiCTlanVfdvEG1i2aWwcd/DbgvuChu61tH4TSEVERiOlpmh
FhMm4kfADpbdAYTnOgH40w1fg558q0vPjDFPlhD8iyqdRxV4TgNdX0QpW3ljauQianMZZdH38vi2
zVaNEjWwm8kL/6kx8tZ8mIXKGhiE9CRUm67PEBT9kYg+FeP2Vc1YzniZAEydfOlqbqOl6kXy8u3h
EqI0u3GIE+rHl/nIX5IjuwWyxKy+OqbRdouI6mL1Mz/Ek792NFIA53C+5Pv9AP8rVXV8z2Nw5R0x
0493y/MpoUDYVc9nbE2a1bfzwzIUL9nClWzhMMGWPaOiSUgxRk9c3wdEwlg7Qx1C8lS9I5LHe1ZR
wxybljVIMyM+uaHVbJp09lhlMT+sdVeAL/rFI3PszgvcC29fwpzudencJhomH4RjaPD64/9G8bWQ
VVkkyLcJWzpguWY6zKz1/2m4P3fF51EliPMwq6swh30UL0QaVaWpZDS4xmb09kZQA2Xa0e9RSglH
A13Q23mG4ftjd/deXHkWzARwOJZJjknRLh6wAb8xJoBdMkqTPk1Y7nkuDgaYSADrTcOO1/OpiJFK
mDYObekhYJzPJRS7e2ZrAJ07XL9oNgLJjFjJU5PQlSPm2E9L7U2gCwRlIe1aMOKXVpOl7L/J8E4C
BCCi1WEvC9DdT1O2T351jOdasxrOM7Z9P+H2k5UygJUFuBQekPn8JarTnRbOMUUHUbgVt2onL17s
/qwGgMbeJmqawJ/fZUkH40scrgOU0V1o2ev1js2QR2E0GBPcb14OBABJ15A+U6wHViX0pEGBd/LS
szg2hfKP8cJtY29Cw8Hhiv8W4VJ2eVlBh98ZHk5NSOg/kHTCfv223d3pQl2Q0inkivFxgug3XP98
zE/9zV5mDXJrZp7isgIGVHxLVkLr5WXgDQrfz9DSBIp+LWhyPISKgdftFB7teIsTgCnrtLWwypte
g8TM8xsENQOiKHz0QJBfL+XG1UIEHjAYX80LYckssiQ4no2+4uSeOyXoxmyv2PPa3PDMwXNirMOc
W8PWVyjT4BnniuIMhPcJVKBmOVeqohSUVTR7DTid5w0BQMsTB13145HDQLzUYREqcvzLjlS9H3F9
BilGdJvE+me8rGfL0zv9UGYacfDt+IMeF1wRKUs+QfkaY7NlkKeqARUUMNS7fbG5LB1WYy629S8v
C1jJc61yeyWf4+f/gmRSw1JG/hQHxBHIoDTHWwfNjSWYCPOXH02MNGiLJqAAEyQl4mIRsC7sUgIw
GJ70/66A6kX6Gc/6y6Zb7Uiknn14WOAQIuALQ7vJPbxRMecr7TAzlTMcsjygB0T4L4D0WytqkDQZ
wpI/xSjcu7xkTToU3zjttYWK/gWJKMVmRJaEtvcipyKeODIFrxeIFTXX5B6wYQk9JUePHTICb+bf
M+COI6VfHW10EHmQYjBFyZvUcCGzaxEGbMqG/uUy1tTm6iKdVVR7tzyJDtovKFPCj2Ge2LeLM6bv
qrhe40eB0iBOSdskR9SN2BZOnfgnJ52sq74zjPm9el8/N5V3arg2vIY+rgZ7FLnncW1/uJuKt8dj
lFfSQLbl0HT0nElkBnh84AYNYk2gLcALaDIlAgONPhEEzU9nzj86gMogunrK66sOI+DppwqVBM0t
BSalztJSI4JDkU7pAkL9++bnyXcL2xuBiibvscLS61utqKFqzPfUw5HaR6Ogzj+xBQbp5QVM3uPI
QZhubDSt+ulLh+uWVn/Tv+zxrXZUbsKL2GMC/0zWx+Ht0l5wMh3qgfTgXruxyEdN1U32J25lBYOv
qbJBBZizW0PUZ6+dkCVwPFttIWt0CfdyNuh1oGnDzJZyn9hsOUXJP0WdfmvxEu2zd4rUOjLgCFDg
lilDgjBYqQ6UWSTJ5raBQZQiv9pl6hNDZsqAzRe4M3g2nVw7Z/unK8wjBfdXfzduvI8Do2dicSxy
8R0jeOTHeUQ/lsc2dP7yn2sO87eZF2IEdl17sOKIMSSBfTfM7qWU5THKjtx/o/xuCX38nbX7Bps3
R/QwBqmXW4blInKCNseSwTEedNhTGGmFOKi9lR3AMAB92BlH5DltSFrrM472aiaqTqSYAewb/yPw
DKCEvUNF2ZgchZ33rMxgHJnwiLW4cVHJ7lVgq7z9sfkPtlNQvM/F52rEsErdDGDDoWX0SMacAxfI
wL55HjOb1MNsmtwVeQ4xGadVH3+5QGtNAVs78DSS3lsDe2EOsmMjQY81Gmf/Az/8Q0AdRzC8nAcc
AnKLlBfOtR4RtYk2+V5x0bmZTjEVTjkeQxr9EqTaNUCV18UMZbIHJLdkX+fi4TIrOp0Ytn0JdE9J
J3sR3h97bz9HEj/54EG8yK3Gm8jdlPIKnSskSmkWRmhviR4LsDIiCDZFrOV8HS1oCVxJF1NpQaRZ
bwfaW2iK0MuisAqD/BMPGsJThCVZGER7LSxBbQ6n7KlH5arxXyiKLCf4MrwUr0FrVy/e07Q1cWZU
DXPcYjH+kZd8cmk1NZcO/C6HyHelFPXHO7MkpxeZxGn4T000HM2llLDWmNSadaM2J1sHUO4bD80T
7QjQTo6BQG1UNyuyyDRqFCrFNpEcvHH+Jsr5FtYz6sU/VXVIjFirW5zmsQKKsTlJ8jkeZcGXaiKw
/Tpk9QsudKJs79BnWBpgCqi0Tkn4aTzLGIrpSTwfXzhC3c1cdkjqPlmUsya3vFiqBbXi/OCkcced
xnboZ8DyxokU8ieU5i0QCvZLf+eIyhUaP1OSvHIb2Zubaz5zeP97L4293/AjkGHlhXO5P2+QVeXX
ygFupYKWGe2sZLOS8tqHBmIh8BKbfJZkwXmM3gvGEvORiqF3X8vs+TtzFGzh59f3GWoUH0xZKBpg
/DhJCNAaHgJmVrrluvnXtRs/mPQ2eEYjpiBjUxZlxPaeWkreX6YsL1Eka3OIKVrOdnSYzhDWId8V
DO+ehNlTHWNMOKfVztQTH9MgFBoSo/GPM90PxKz8fsnJNHZ33zTPn+sIcTizIIwNYCBXuU+QqeYM
15v8HqkjmK7BPODTWmvI8MVkaOGkVzQyJ5kfYwSnlGPMvUjWJl98USX/7XOITRnY8AwzfLV4GO7I
xrHNNiW1feV6byslWqW0sI2/EFP44Nii9+AdpQUftyuY/pw8wHVEYNjdMRnWDAk6uVtk7rSNZxqw
tlfZcigRul7cr3tPA6uB7OBF2KX/7a9ZYFu/OTvWN7Wnd/ZYdYQEWr9u1dibyanM0StPmuuTu1ge
k37sfoxoVfbSOPTLWTFJHmOEZxhTklKoxQK7t/kAGSKIMdYFA9xZZ+JP6sBLAWtHrkby7XYsadTL
wWy0rbNHP1DmnRab/wBmVTeVeM8xDgTBocNHB1e45f1DrrNqxWM7hAvhnpVaeMxUCJEfIwkw2TYR
5WBI0MWquRud6UnR/G7qiJ6bywvA+PvOEPS9FLkq+sRtJ/H8sVbuiVii0R+Sze7y6cDaiOqipz1e
4Fm6o1zchbkVnxihdHl/pnG4tFsE51i27DUr1/EwBMmyObNMGterdj/+w6JaNqqDUTWIuZ5hUfaY
seGLK18AGcj8mbEs2ZUGb6SQtt/vZyCJbNY/jBvyuAZmodc9jFVkm7dehj8PqWu2cMs86uT+x5ke
VISXA61AXytHv8ZjcMJMsSAHxAtP/qIrUfAp/ze7jOjTW1pQIBglT2jj55pWQRRbyObJ95t3M2B9
nMR5E/PH/IR5bHMIK4f0251ghC7QD3kevlCHxOBRiIv+Fbp+YjGyTAPLE1WXvIv04IujyJU3hmCS
2MV2a0lA56k/Pd1O/tKDuId3nThUbaLtloaCKr5WqMyEuG6KUScLe28KZ/bds0wyLk4vL83SRgP9
dkdCvIr22IP3ZCg+YUIPa6Rr7GmFX33Q4b3fFT7q/h0w06ejJE5LEwE6X6p8Y/Rzo/LEtGn4ZKHu
WXGwLeVeZNOioBVxtlXkR9fX+h/CG0HY8HVI2lv1STDQEGNv5zCrplYAYPQNK1zqahiLzm11EUGj
TLg0JQk/qCtBQnXdNv5H82MEIMkgzNw9nJbHrnERVYvXC+gDu1AJY+nJHtvu/648uqERaQZn44E0
7/Wyu+uTVUVoxWmFBeiHfT9TrY9mrllJfEv1Jq0lGrlZdvQY2UyNvB5DRUUYquydKo/xhGIj2nM/
U3O8i0KpauadrUmlh33Wxk25gcVLT/O+mYJN7vmVO86gKr0pha/fWjfG7B3QS9Lnd1l8Sp2zwQto
3k4e+xEs2usZiQ5e4mO7Ha6GjxUV9+wkVh2tgQKFf7pXMFBM2g8hcIKgOXELw6+AE9D8KmV2ufdN
f/AdD+LsJM99INF3ZTl0a1KW9DmXhQYkqp2scTkZyJcPTHgA+bUKEqe61k9hYKSD4XevHuYv/cn3
/hKTNCHQee+q3XpXikHT3kRYt7WWQhdRpKBpWMCaY81iAzIQYwcQNADu1mh0hRo0wOCkyLobemTs
A3AZz5KJu9pMr3l7v7qDj7V5qcGrN4P4BpuxTMi+0bc7+6zuGl8dJcZq+/tMZTdXZDhF+9JDj09s
sGB6yehclyKo8UCrgA+DoHZzDhwpq3I/iyLzZ+VLolNErXDV+yPv5XN4AHEuQEQHzASYQPGrk+Vd
mum2fjqoir/rtgPJQ4lU/dfwqrqq+4uvg1anzb4BgVDVwDr+Zlw/BpAyGMxcU3Etc+Cy+kyHxjfz
rhmviCMANXtKQdgp/bzn03blRfOXx8nFUTdVsR+BOn1jYjdcdrhgEDBok4dn1mYWwqfqJ54jU2TQ
7IOoHVprybgs3pAr5UMDPv7LoRnf+6DCTtvXB5vjenDeFS7EKbXUgwKP6ajnubCsbINK4doEnCmv
bvoZgumtMr2U7JMdfCWxJ7kDZBJiTzsenqH9hd06QYVgZuHmC5rUzFtK9dF3paJHtMLjZXvGxi+R
bOr0GIXTrw6VE6IjK/J6Lq743siYpXd65I1BZudj0cHt1J50OWfqJ9ddQ7AjC4ZQcWx3Asnr/lSK
gAjpUTUMBP7lPrQC1+LBpb3X3dE4OIS/J0zYV4PEcZMm7BxsN6Y4r2pTrpqr7ZKp5Q4/Bp07UD7g
si7vzaOrRHb7vpoS3Rm1wA8XtbsvHjDVtj4eUKAmdY9sGeTkVO9b08cecMzvfKEEUo+7YDaGmKg6
mmE1NILncizbbDVPpUbZu3iILUJjtDJ+0udL2FVCEGg6ayqwCrgkAumU0wni9zidLjYDVVrS0XGt
iWInYWwfWIkv/aSPpmC0M++XguPnQBkmU7dE/pmhQUrY7uLpZwloxLnhC4YAb1dlClO5BXKJp6st
3lHooV4IMIe4n9/D1MLB6lHOtRt6S6U9JKxV71Ll5Ro3K3yFsRzQSzhLlOCyVh18i8EpRWQDe/KB
W8X/axiKrFJacRTWoeAkAChMn6RMAvWmx7yyMGeErhDx9L41SW37MJJtnubSqRJFCBGZuZ76ZfhC
3roCVw836ZLL+hBfQV8iNlZ6nDmRcl2Kk2aDMJvyzawHW0I+iqO2VJZbTwSCLjc+4vi5Bkq8JGa1
VQA0tRXuuH2qbUqLTHPCyeQ/D4VHz7zX88SJitHKr1n5vHcUz/kg6G+fE7Y9myhpXxqqHb1RyMJ0
CQN32AlOhig8svA+sr/YIsBks+//zK1L2Ytbooi377sqadRAWXtcSjJvYqCDrPBd/6YRMg59lK71
uByBJZX8epO50+shAdddRjSce5KRiXUJMblE6tI5M25PRxh5q/dRc6WjzCUvhmlAcDKMmkPHRhdE
7Fo25kSEZgOuzINEbswAMByrPDV+1VRNglMopsD7RWd26BzzPiAbu9RdCnvuX6Hz42I13fFAUyz0
PivDD7ul7+o8N6N3BWmC3CrHahKpvfJtDTU8mv1E2VMF9FpdRBNpWMfWk3da+7PbuyQ5gI+omjk4
amHuovLxA5e33gWwFvprf+Ei4KcPNIrr432ID88ZVNpdo5WlJ5rt/8V/mmD5Tc+gO+EmC13mfjQL
/GsvGNfDH2GpqZr5Btck3XD7tOq0yUbc7+LHw68zUACuIFBDOZZycc0fLbwEg3e43dbc8PG4Urq6
ibj4pkfRXsDov3a/1qbz+GyTmJ3LQD9201J/msg7wrqKT1/lQkVyr5LIZxtW8Owj4XZ1nOWG7CnP
Zw7BH1fV3YJgqe5LAEDzgYAEeoEmkCyVPPB5pZ9xKr7oKt5NvQtT4XNCShmD5Dx0NfHJjEr70/dQ
rG4k//oqkl+6F0UggMmtj8v/BN+JlpsynCB2pw1mGVgC6HFumMYiZfgHyLe6l1DhPt7antSKJGSQ
nAaaGTLCw0EPWH5XdArcicjM0QwuAsoXiGYBjdAQWeYoS7qpYduCwUPbVVNYrKDHwK6fpfIof8qH
U79hDntfT9UrIDMdSWfWsHxoyfs499YTy1wv+xYfhpSne/ko/GjY4+10G34nqjZAbC1gHhFsTEs9
3auntdJ+HbZal3dLSFNjBTs5WBFsNA8DLDi5usL+nPyWIQqjzcusm8TN/AhTYVSvgisovgiO7XL3
cxTVo5t0Z0iz3st333sDM51co5x+XSK/41S3aMGEXHfqBx4ehw5LH+LA5O47MbqzG/Hm3YHh8FGQ
7J4d0Fvt48vGEH73eZQAzj3TJ7+ymC+hAmzf1OBNKwWcrYpcqaqHRzZIax2grYndAPo4F1Jf8+ex
UCjErrKIdNDe1wXXK99OfSUiPAYKQ1zwE+BRClS2Wjs4rjkNObQ0+0xLhMScoHAfiOSvoiDb18RO
YNaICvRQtgLdTsoEu8g5iJ0T0nTfQRcxu7UxzXtUpEaUI75GZQ9N4kFKyReF2YoaUgVPscqVqYNA
u4jSrVHzcR9lYNhGN8mDe4o4KhYWFdl2snSn5spiT7ygzFX/qhXKwKdIhOtOcn3VnTaA3zQ89pZR
cJ/Wfj3wAWtNLvAH5CXdyrajJ9oQ1vn2HEyUQeUzbGz3bOnZoTQfkOyuWdqegQS+3HeJUzvmcaM7
ZMQlHhkMCHSMrwkx2ibJ8EgkTC7tlynKR19mEJqC7zMjC7dqkr3I9BqzkZb2Kx3JceRlx5yYoAso
qkB+R3lG6488ORNHx07xeDzFeKf6CjAnxqp6EM9eYrnrEzANsAYp6ot0hjdITF0cNf3kp4UyvAvK
P+k8UwcQKfKg/STSsLHWIcE0/ppjyi0z3EUnFK1jZWha6dDM9lXSmneSUYEcI931ylrtBFcANWG7
HbDug1YntwScstg6ze8RSariAGAQ6XbLHO2x714eMRhT/HE2dGzNtma0sPZl6nZ5Ndqki6ptMfxC
fMqBFee0UPl5F1I7sLszUYp3GeAFbIy1wSppJgOYr/YUZjgJg6Sg1j/ruKFyNIv02vabgxty7HyV
P8nR33V4GcAdtniL1TgbWvUheU3HNrDXfrlLP6cw6JcyGod0LG6mWSn/gCWQH2sNmACkcmRHkgzg
uNXUQ1WOoqvE5hNgVRuQynuyzqsbYxq+Yc5I7ETBFh6HsfwzK3nGU6Li7E9dTxPLlryaDoCI6P29
PIPxDwHUG8OMRekDklymC0323sDmqoTwBuVEURSyjYZaXMTr4xSqCfytOTfktNJCjXXF7MJv7X0m
2Ma5xEgdePS9cwMpJKiItb7WeHL3dyIzL47y/jFLv8zGDwCUPRQGd+OFU8bgKx0LoecrWQl20e5N
Ny2N8hbjg2bCeX15aRy8g4hgJbAek+OeAqdIvTCeT798RxP4yeWIwjDfe6ZG67p/YSmf9Kf74/qG
7gIAHNolTCh8HNHu9zOxcWQx7NQ8qFHTWuNf2FIxrHkNOFToZ+yrvyhkWGncIJH7XlpGqng7bJTn
YU85EX1gJCszp6qy9Fe0YBTdo9cVlm7lApcJD2u0B9glZ5QhErF0EzUDfluTHJ6hxhxLtPoIpgWJ
ov7QJkWGhGgO0D1x+G+FissghWCVa1VtGqCzSSUDjIoO37qsT5+2fgony64E5IZOvXUB2fTc3vhc
uwlkwRTZ1oZePYm8O5oSxYqR6UWF+s/qGZRsxQlcxHOoVScxbgdCxc3Dundll+2NPYaC/W2ppRa0
qKyk2vFOjyROHLED7lvT1kcFFoR7QTkXoS8LmNSmRj1bVdi9EMShXvssd5aBEWU+bDgVXOTtvKxR
DjoSduD5ZNvLUinPd0DzSzog0BsQFNPb7GIBMhtHFwnLgBzXROViglgGGex4NDsGmpqXtbcJhpe1
QBGvl2N0GWeQcD5R3Efq51GBj5WharJ7UL1uZks8CgxnWMkJROYKaV6KcQMYqK0EFgOMkzfCg4d7
qp3jfeN/uESn9NVY7W2xDPNWDAD925uZEzZRfVATs5EJ+ypAEEnXVjtYhP64Y3mWUFEyGp/E3Nod
ax2vjWzvcTwjapCZR8HHCPiBh39Ufx+rJV+wjKiDxRwdAAybWnzKsAGTSDmORyjXX0Q90eWEZe9q
i2+q5+ovI3e6tK6VRWDM1ci4l8cByrv+ME/8AmaGLFpQiL8FvytDIlJPNJ2cApqnB7Duevsskyuh
poIwHbHY2sbGiXumP0AKPLebJjTF4ZzEnDD0BughWWGgymn7krRX2rwLfL5Djs+urY08G4unCdoN
9VqmYtWO0RfLMoPHyasHc1Mf/99cfOIBjxj3DwB7CuXmgW46TNDc1WfTepsPdESKtjo98xh354T9
m8n9NqE7O5ahgaRzzJTVswde+AGvg8wrFQwUfjJ/Y47IatNgLyg1MjKfTDxjbM/Nscyu96+XELht
8ERVG9OEsXL3Zkv7KVagomAiDXB8Jw+bWX7kYmMOxgcOcDNSyt1ZzS/dTsn20g5OTGF9upr4yAYK
X0HP/99iilMBJLWTPpvT4jOowrc71nyTs6ukqTsRdiXhvDleOm5qaW+Zk+VgtOD8VjVKeDwgdEfJ
yhEja2o3DPoujis8VpfkAW73wPMguIBYbTBkhR/rDbkKUY+RgAnOXGAlfI2xNk4KrpaNYthwk6Lk
VnMQOdGMae+vThTCqIAOgA5KxAoM09HdimmLktypaUedgL1hfnJEwq3Tl1mf7yN/rmjb7AmBHzwh
/Tq12C9wjyXkEwRHLIeUa7Xp2ikJ+IVt6iYs8N7cjOOU2aR4BsHgPt1ayGLxkaLcd7DDRpzNxcnZ
mTSSOoiRmtIDUDCkzC4thoAbtPwIG92FrHP9DZ8bWQKpqMLjWqpvhFlh37wewsMS4K9X/hcz1qx6
A85dpXZqjEHSVmEC20hzDdqRoDEeF8RT4BYRao25Qf4zilOfV1hzuQzLr7HpoqAAyEaJjNToqBuP
eVfbgaOsj0anuskX519Qgz4l65HaDw2FUn/oo+/0Rd8oA9flhq7siP5fM7Xeam43yp2xp5cjP5+j
uLpq5n92zccWgv4rO4tddeCUMxO366de6ckjCuGcHxbZTtLKtSD2uu3Q+R7/XljpUGSVLCTMtLSi
L9ifXTjK7kN0MRTFpRniSuYjuFt/M0/nQTNPkCk9UdLK2loUIvmrx+z0Rd72930624+ixE0X9z22
9b73KNESKYXqUHB341dhhj6B1HED6x8bE4jt8sYk1DCZTMH5Yylju/JzwbC04vHqQRgwZj+jg7ur
kcuYdvhHbVnL/pNCJk/0w02tZHRo83EFShEM7tbW6syWWHRPen34MKRX5pC8hnUUsY5MfpbShsDF
YHn0jj8fdlcFdCBNZkh42au3Q/X51nAaseU7Z46/FmZCEQfolsyPwtpevLYFsVnCTV3zgg2SS7Gh
0nYUNUVmhUdSa1bj5s8ERTWQ0ER0KwrGuQptEf/T1wFF2FImtVaA5IBvGAiECDb8VYuQbyaJDg1x
ZYuiXiGTUg+DkwZdaziTFwzFzMGI6Kzf0VYFt9+mb6cq7QpjmGHCdXMIumZGAuCDKZzBv5m4PxRl
uMbm9Ntp6x/bII/YLJPofBYzPv5pKks470h1rrQfR0FvudL9cFIOCrnTxcczOYVGKNRW9Wssd6HM
6YtuxYB+y3yinAU/NwPO6LeoHGmvoKxekN8uJQ4rPYpxrRgjVuXODju25bA+jRo86HCMz4hntvRc
TbZi3ltogltJE2T3kliLpEfsePbishjXEHyZ/dCt/9670kW0xEoUIkSxssgYeQvvFRD3PBaFQgQ4
Aq1ZWQmyPN6HPrMwIkTzRltLw+bjnQNwuAslFUCxM8PzcexZjWdpUglP8KxgtSZ/+xNIynA4h17G
aGbjfLSbCxgzKUeYVwFkRgx5lx4shF58PgJ0KqIZp+4Cpq7OJWTvqeW0OTEN1TlwBUDOr6/JyCAj
VfZ4b+v719Mg5VO2jcVt/GrmcD7sXVTxYDc/iBZD3/qBZyMUDUEBAnFwrr3i6Z0MWa11WglicSmW
LpnniTWVlII5tGMdGxOhEt0fHK8w3ow8krl3a8jV6ncOcDEN6SKshY3mJMtKJ6cv/uCFMxhJpqkr
6kDGornQN+MTdlSpl5gil4mJw5C9JsdBGlgvvnS4e0Af132iPwI5UXPyikyCZgWBsg6VfuLSF6Vq
tiBECTslxumkkZ8XVluCStvAzI/+x8Hncaymvokbi27Sb9oftzeq1pp+mYfjhPZ//I4QR5GPvyud
1YkmUwV206CS18OZw2ixQQwI9tv5dOQHiJgUHFlO2JQrPircq4xm4fgId9FQHYf+GQ18344mqXPN
j47/gBc9IG3FZsbjjJTk8E9ssHcSSZuu3wYMIWKZ9Q8goApjce4vx0HaumTSck4E8s2fI1Ib9nsz
MnHsb/ICDALrJscXA88pkXlGtpdGtVyNgOhefd47WOVMcBiLQNGAcYSseDmopCgEShlkENhgAcUA
mGR9mCQ81Wh+ERHBtdjt/qS1sfzD62M/FcofG6+8O2lk4+ZGu+ZauGJeKP+xgxiBGCPefd5gKBxP
8LwvAMvdwJQ0Zc4OKWfJ3NtYzDu43lXZJIybHOUDG2rtZRD0qafm8Pi1F/sP5YzBQykBGpPr9OXI
l5d4AyhBgpZQSGXlnglzsWBLXj+KKs/mdyuPbeFPWpxZ9y1IDzYlKSQDok3Tw0h24WRpqHdQlSYc
RnlmvE/JcFasIsuhrwv5aFxQ99ZD4NKJvKCmLlAOJ+Bgrq2g9rDqKEReSjYUIr8LKmo1E55EpQWp
RXGWQjUDoxVOKnvgn2FIw6+UPgGaBpBmE6CF+WBHFC8PB8FFeP2xkCcMEhe9eWfm0ZxHCZH1+LQ2
PLZDJ3lXK/0WgNOtT6eIX+jjc+okYRi7I1TsvO2IYKqqTktuqy6AD29GC4fXG4juhokm5In0XE5f
a+XXOISsOUeWh5y1xELJGl4/ln3Q8pIApfYdhAAKgcR+yDwvq6vkMvD4ZnOfxByjp+murefm54He
OhayaXQcDc3ArzJngyzryo+/oz1D3vOjWEoIwNPuETocUDmvzyjGPiRBtZKLiJZIVV3jaTmdse1K
eyf2ck2S3E6Huqbmq4Itln8HhyIL5z3Clg5yOkyJZuUYFtt28pYmZ97TyisXVshnGtAjcy4NGdq0
vjEmCs/iya/mDXDX1rhMZ0qp9iYfESNEQm+w0NXIAre4fTj2DWWycSEtKeuWl0x+0Jy0XwY9JE+q
v5Sk3l2TjYihHo7FVicUgG9loqj6X6oeTr/bzDvRLe8fgte5iZGO5YayQdehl47yCeifg4ML7Vat
J7SnDj3l9N/MPa1m91/d2KvU4BMUs6APvGoKQGIaDw1r55VxSKjlbnhB4bM/jLupvVRLKFTU5Eze
egeght57P/PvVJ28AzCVYmchE5mg5UrgH9WAPeqFiUZEjO3e6qzuPpzQeoQPyRkbKSzeOrfjTtpG
kS4JJjSLKhRBTy1vuSSCRIwMZ4+80BI6SIYEGS9YCitIlNg6RpmBWUW7yK3FjPyWwVsNvIVj5h08
5dX+GpHcWzuzpR2QjAelIaOTsTzgVzLPYh0c7OTOC6Z8p5qwGj6GGefyAlLKHxNb0Oa+4wBp81Hd
iUKu+8+qVRuFPaO7fT4wDYdMUmrJT74YoMWkcKoddPue9s6Eqd5N2hhoXSNAbB0ZTnsNKO/2q240
MPELmg23neWGaAvJcUea7+zlpDfHMkJmRIvIsg0lQDWAGbiExRJRxz8oIfUumsmOhQ15C6MSzQIp
YpnyMNIBGjOPI+lQi++0ELQfYQQm5oTB22LyChX5Xd2m51adaE8Gr7PAhU8vBBfcjRfoCMpuHTey
bHtPgDVgoy1NZkjJcVvn/2dkLHBzlC6eUBv1tnokfEFtHIwCoO6B+23n2NDlcEIRbkGqRjEW7ZZa
r5I6wuq1YtEz3eHESBTieatvL9M9QrboYh5JZp7uJuY2cF992Z/vE4dOF5qiY76C2tdhbT05TUhT
R2Fk7luBgAE1r0AmS/ttysGJ3gCYB3xFHGQx0Y/e5J8MFEGRogt8WkOCeDuQx15XnXGt/ZMXFsjv
FayqBq3fkCjJddYikt4FZhVCyYetfrjUX4eildMOzzaiCknHXQquMBtvYpsSlD6nSmu/rMD7ieIl
/MQFpYbgY/XA05AesND2r3DjNsoETpbMwxF4NRb+5aeo2mD7VZg891h/Z17wNZL1ySse42V+1LBw
9+HsDagD8eqVzQZ2a84sbeqTCzaLxrPWfjyUy9zIBEzoS9sWcK9GvBcnJZH9u1Yk1nMThDowFZ30
po1R8D/QEdLsIm7BpfzRPRZArMA+vC8R52RdhRcV9ZqdgAm3aJQqYblbAE1bl684zs4wnMH+yE6Z
HiGJMQfqnsZlo42XY+tSpEqqmZTQxFcMoaLHqMJEvjlxrPMttPgEKrAtANb9Bjzw6VrEsMlnr1SZ
Rdn3DzhMnieH9FBY4kje4S1IBqE+a/bW+Ei75jpvb3hAiVtdoJldDxhbmO0N+MBfomPn7gde7I21
zPP/NxkowgG6ePCBn9jZwWWv13RHoOe1Buvvho8tZDqzBLiRMdHiPMJv3BtGYQQikUEJysQJuEbL
RCdydd8LP40phqYLtunbKXS2ZnaITGZuJfBTDFEXK8xeN/SIbWh+vzFlUYbcdxPI1IQjw1TLmYhI
JxrcqT34sgR8i5VxnZDe0/wmZkREcFge/My97+Nh2nfqMG7cDC8IKhYNR0cYcobT888qVkkXurwt
HmPcd3p0ww14G/W3GJ+SbB3RyZmTRrIN3+Q81P+grsT4tvJdwVEuck8LxEgGtNgQGqadCWtgHjAY
MkxK5zTePb960kJZAQGUcFn1/If7GgMaw7py9LdS6ObN1RFhx9vCcaS4C0BfloNfAsRSNFi51mOw
swe1J87mCmC5A6s71lcYkZYBV/ZCcINXAO/0TAf5/BOjIGN7BxiUAw0jDVKp8nQ+3wNtO8/LD9ZC
MGOo57cbTkHMi+V7cQ661aEOYSbl67zwKgRSvNLFi/GWfPMDYnbYUV+zfseR3CaAZqLr079MOWPr
tOf7p7yXqsbSA9lskP2JfticnOXhUbL9MLUtzEnlmVdcSWA0Q7s3ww/OudfiIjNHd6NfpguYRxxb
z+Hk9Pxf/WMP+j9Ys3wLnkq6affRfzzQ5xOp9UIYnqKUpp9L4MbS+rDaCRIZN5jODBnw0rCu7VEF
dX1OMDTETsf0mXd6gAub+UkDU5JKJPjpzOkzg8vlBPFplrbmQDq8e64cOm/cD0bMwkrziJx0nhZG
lPJtnmm8dWAajmZuTJizyOxnjpA79VPS1gHccHHd5Bl9d9zi30bD5V97s2f8A78IXq42PV1ZRtSL
UQ0sx0is2uASRdu/r2VpPP8zvhI+WVaCOjLVM5vtLeKmikhrcp4r2m/wVYekgpMe9z+12ms3orOW
64Y6LeeZA+bazddjf9Zlt7wz7Dr0yFXTqq/8+QLJuCce51oTmCe5f8GteFNe9XOSvjWh5NUp3vA+
kiSZs21juef1v43ULV9/zSUo6WjffgKBFCRKi9Yl27Vu0Dkto/sRhFtyvThKfLKscZymVCAvrKMj
STnOjnqAWW1re9ClL7XnF2UEnP8S4RXVkFZc6hOXFy83v2sm0sJrd1SFeyLqEeAnMUybmDDNCN7K
93RbPp2yOKKj4xs9gtGhOjst/Mi1I94xBmqa/iBrldH01kxBiQN3vAIFzLhdZ47/5jdT607jsini
l6qu66dFOx6lSSOcaPBwO02PHpHGpCuh7TSeQURNkDKwZH77ssgr3ZqnxGHFxWgto/f+O8biasu/
caGM9UG/Mb1bJMj+k/P4dQ7KzOdQUjY4Wm50y1o5YbNdskVq9v+2ukX9gFR6VmFe/tqYurPM9OSu
mohDT/TqNxFwjAcb7DHUeVd4nxALg1vWn5YWFYNPTT/yhSpmbme9f8Rbp3Ui9hi+Qssl5v5o6XSO
kLyl0ewJC1FLoui2+Wc8WjI9AIbMiY5lQEiam0jz/fqynXY5sVpdFfeWhstZjServMJPdEg3RGFW
9WXIJ5w2zTp3mG0oQ0q4WhpNi0tnR/omBfCXUlmbAJu06j/Y8RASkvxb/au1sxovfPmeLk1yUW2k
Yi2Ezbn5QIBvW1k+4w3YbJQypb1YRNd/PHR+d6CdP4DIvcP42hi1Xr4O6hwN0uN/noodpWiKUyGn
L2ziAmyVGNMyyiZxEsIBbohDppH3TaiNxLRlRkry+x8E6imXgEpa+AL2WNL5onBrLQC63uVGO/t0
qpXlXzP/Us03hXUKmO296/EaUtNDcm7q+dVo0ps52aVEJSuEQCoGySWUTeFJJScFR8H8/avtafDB
aL6i7jMxnDyp9kqPM99uZyqkjw6HhaO2Pkun7gAq/XQyFU69zonPU0XgGVimvRCgFkBDMHSNIUSU
ByG2Yutyxbgq2KzszLEpG9cjkjuvvMn6dtHkKxXUHabp45BzPsA7B363DreDKY8X51DdlFt+YiOJ
puu4U7bYpvjiTdfNAAzw8QoddXZTJGGMQpRktEbrakfw8Z4IXj+hGxgLVfJtAeap6oNeXbEx48jc
1cT4aUJ1lPtoche0mFKlxUwIgmuTbSa6sFeyXt0PZyUIN6rnMPiqke8JIypn9nv5a0XWwwdPmVtA
Mhz00m+9Fhdfn7UgghzIdbtNWDfB/H0iKbfP0Io5adL5CF0QtY++UPBT4+Lotn8P9Cora/ZhgE8l
4EoYhQTuEsC1FY2RJYwflLhv3N8ek/AW5KlVpvnDzOGGj9iDkPSSUtciG+ES16Dyc47QSSKl01rf
+knOfYGkvSTcoirMVLDENL5KiPHk4b4LyjxM098Mq5MkTGl96AAwhqze5bVuPtbOLwjeYTABJgHa
A/VHS4HKVR68SOKDDd4PcWkqDUoEoM5sYxU/CifXm7yNrOLets9WD+TXYiMmYGeaOH+pUEIceBC9
8kDWbTpzDlwK2DLnjThS2GAqwrApVTgL35FCihjLjB1jApIM1CRhImuFqLJaWVWmN3qZCecIlGan
1R4a5PqPs3SqjsiX/mKoPhE6Z1pOqMF5/2n8ho45YXr5pmIe8fLXoD/T6yY609h9SZSQgj1dQrdz
g2c2lu277SMFN0jiYptpsX6gv109FpnacTcKX3gGefCUvnxLKAThST4LiluF61Bq09Pbpl9RLmIr
PRM/vHBv2AtPUhxxTdzoIoZ/NKRQRMprDIHh1atVmeWgB+emiHtWsC4mvVxw3nVwjz9I/QR5foox
/OzUoXXQSkcQ5C1KFruxYabEthXOp7kJPyE55tYfwunf5nsPFXiwtdjpudYZh7Wo+m+gaBHvUusg
vUv1+0c/U831dfAY4AOU+NsJH0JS6hKGLqgFe0WqVruvOBVjtI7TcKz+zKrECQbwNJuEAoMxvpNy
iZmOA63fGpXKq7rXhIak6wOVP8mcJwghxV/Qxg9aGYxkm2gBU4KKNN1CZfxzuzJ0NgzDfDnro8RG
cPCGN+Rkdg4ABc8kjnx23jC/S2CB+/JpPhNFm17iwOeOHY+oSVm7MRei8y200XmC646a9jkDIZpQ
novsPUjKqugjL9y6gnSX9/f8lvQ0i9hTYr/o/WbnPHnh8lP5s8yrTALKD9iJUBzhb5shCXIWGKcs
b4cqdbQTKCEEHZ5Qi2p7MEhWMZAvnLVcIwCiUGAmaHBOnFYTo/kV5yP77qE2d/uUiG4NL/TyBInd
/0f1trvE0s5EVwIxe5xCShJVt5Vggwd8lurX5OQSXc4blEvqV3qUIkAdqPNPIWk3sDDvIaKQ98yT
ayh9eH42ZGYOPzIDK52FWFI5cQBhQvGL6601qJCu23UXovq0bYJfKjauwOCuVkWCXv/JQjKb05eU
z7oueLxMzXiA5DqPkZIRDCq9FILTsGY0olQOIFVNS1qHpzg8xSVy9km1sL8xXn05LHwwwn231RQt
2PjQm+12UUNRwVRZb/Xg1htq/MJJi0B7uos/fXZBPEbG7obg6Cg47LdFTwxBBdFqz8xQatS1Mon9
HV7CdX24BEfK1dHH5O6B7wABosy6U/n7XDhotljGkYsVoA/MHV0SxT5bCfhIb2JEjKJ6wHmGlsac
IuX7i3uT6TWl8+2lFlj8UMlzYVfISUB5meTG5kQOD62Nx5gch6GLFcFQ0eEMikPHT2pp3BTIHWkF
3X4wMyTQf3Mz5HiVml7adr1ubP2zyspWiCs9zofmA6s15VHoDCxVUdsAGw5gsIZ9za3qwtZnHyj0
j4DVtjdsHboN02rVTwxD+lRO06XiPUQmbLvxhUL5J9xVPWcrQCUZBp9u5VEkt0KpstPgWJos9n2W
DGQNzsKBeAN451eBjHeuQGKUACi3lsIjtoaAkOqclRJk7+VgH4FswGEGhuKb7plZ6+oqy63SwKC6
iJoWquKXrfRJzX+9lHrPs5nbBYCL+3qCainqz7gtqgdOzb2/tYJExVoMui48szU3O1SyyuMSLP4T
tKeH0OUs0hGkkw89zo4MSL8X+nttvrlNKmpg+YHBaVAXQ8lXePRrtFvRKW+xnMUyx/N+J/GbeYkR
NHN/ieEmJV/tyghBZMuNHPLYnpUSM6/UwIXMd1ypfIwlwsKixxFRXZhbGi6QDVNX8SOOeabJ7Kzq
FyNk0kenKHFsi8+ZK1kj9u6GbezgCywxJKdq8tssdtwNRMzt3WkSOLeEAjsMpjfjsWXpcNPHLpOY
6/5JEvX7/5LuLPn93ihzPY9izGUPCiepfR+J8SwKFLVUHnbW6rTNKbeW4vQx9i/AcbGosgUu3mBk
n9n5HcYH42YTdwTl0NphoZMrFMa3o2gWjHzhKAWb2RYbKXM6c3S9p9/aUsN7XTU7KaMinI688KOJ
7TZ4CkVSE9VjiKO4h6Xda6RuI9SlsCvX2Abg6BqaBTbHIqwNpj/rMop02vAIm3KGtVr6QjOqzyls
015ThbI62nI9hKSXldAkVFljVV00EnRQ2+P8xITBRVraJ+d9dKz6ed2ggVtWL/kyRiWVWlOV9Xse
IiXhdGb8fDO3Pb/1nmqCr24tdNZjdFe41L+vaj8Ti4pNT5kbSx+hE50eRsdMGE68bk/yYZXM2CDF
KL1SB7jnarcjzv5SwaHYjQvtKBlMlHQy1wBKTFogkNJvp1i8fiJCtqDZDQX+d4WQOnX7XYhHK0KW
AaNN5tVX5nbzGCh63t9fMhoGbQsnlkSbm0ApGG5cvFrwj3L+5WwQ/yvOpi5CG1tsbrttfzxuOBgo
GWcIExRQ4hznDs1r4+J8bjMR+92GTYqX/zuKfSWqu88JsNvR6ywp7w1z1SAsvxywaIeteGhQeoq3
5QrwGLW4uZEil/EMAO/GXjicYhGSz//CXMkTYN0AThn7oH91eSIZppwvKPWK8JCZ9NXFzIefPeQO
bSA2+xZgPAfPIaFK2qV/CHEO+fhqN/0dxl+i5G7m5SlRUQZJYEdC4prhagjdn4syN4zCMYaaAFp8
KUHJ221WvEDG/5e138lT3aPF+/O3D/APjFu6pSGRKH0gz3jX2eQXSS8aksIuXTUaKaDacdt0MHPX
MQWfbZK2dvR04k/7CRJiaJfND+RnNMf6TRIemEFWHKPimpMYOUy4NlZWyad5gKeIuNVXFv1rLzWS
N5bxN9mu35rsiPJPaULepO5W6bqOIk/LrHMYPv9GZ/vwoosh8ETkHRhfduj9/3+1MLr6Jdxo8blX
yCrUvWtk5ZdLcOsEco7Z8YhsJVqFKu5HMY2stCEVBhi5HBxWNwXTQAa/K0PIugzLCnSQtnpdvXVE
qtQSkQFyJsOo0iZjrE1nTX/g+uflw0gLb0fr0jvraTEZHaVWUA4vKvUZrQ3UBjn6mNAX69H+cAg4
RG9h3LMwhsaGl8/7zA+yQy96W9F2FDRUW8tGsV3zTdZoFazzKc6vHXaZ1mkepUUvPdNJgN3FGblU
efakYQjOXSeEJyTWkS7Pt2aNbmF4w0QnxXNWgCL+9vtb+HWcwX1DkIYSRXw+REEJbfIC1ApxosvD
Fi7B5W/9/y6XQUaAALUmHaOzJxlfrOqQGkHVBbJKWR7QiK32td8AGfFzEZMljsvvuERfibutpOZz
BIzj3S7HGaQHNXUFtx3u546vUtM/Lln+/oairdScAJjaBdD1kCVeGOASEuHrigLwuP/CwHQWZNs4
JER0FA6aCfUEvxHHSeife3CwYslA/yI0yYtzYidnVfKbFpgVgxyO5UJTqwDqRK/DLGRoXidhaKhF
O6HdoDIk/hjteZ4Am3dIM/0HZMlcn3JToLinp10qPFAUTfwW/3PJY4KbVq4oOk08oLSXW0XpX5Vc
rfoIPM6/GNJp66YnO0w3iLvz+1sAWONzivy6/5bcwrB1RN9bgGQuX90zs9mdnbmlnE3AtEKc5bQa
Gx1RZ4gOJMBBTx5xDRUBpeMvr/iEcLXGXuM0zEJ9VLl9r7Ikbuxrq8CXCOckC5qxQHHpp7ZpxruS
Zk9PKxJRZpzSzIxS/4SZRxf20eTXxzY/zxODV52Lp9IIrd2d30oPbbiOtGVZvsF3tlUA2DoJcnvB
/gw//d5tvYDzcKqcsqTtZfHTk8nqAc/eeZsgqczeZdpzcI+KA25fpajGjXolpYTZuFc5E9jq8shN
WGb0C5cy7Y16X2HYjO5LrXa1Ytghv+vHDGdP2T4yCuE/5NfaEC8FtXI/m8kZp/5+JqeynJNXqKPn
gRxKUHhj4mgos0D+/Q7FVS+XsW97dbM4fAYfeLfXSemC8TQVbWd7J0pMMvOe86x9wWi4cxhoy8cG
AJm+HYXD8+elmcirEuG7KMjBOJskZjxyYX7kq/B4NdC3jznHR7Qn/oNnS28Degdke10/c6+4R8ku
kRUYfNs65sUf08iwRIeoKCVTfFpuGpCWKz1j9HJE0wcM4ouldIHPVDNmUW0z9n1u1XCsk8A1PxTI
nga2yRLGvGhPu566jACnCL8nOb8R7307+3OTYxRd/UIvtH2Mh9R0FdmYM5UA9B0oyvwvxu7EskKW
4Ole8+FizGNCtNpuD1l1eFaAME0OLY7/z9uoUPArlmI0oMIICzXu7A2dfYz5XjMMNfvthScVUJRB
8SxrAXXKVEDfaMWq5uwYxLcp7wkQCo42voKaqVTpSqHJGqI19spNgAxim6ZA69REGKYqoOvwQCFC
34GIH3RVGF7TciubUegmQXzz5+25Meh+pPjTo6fv2rytz8ELJHHC2mtNAEbUx8w9HCTi/Nes5S1B
NVqX62p1QHzqwHhShAuq5N//rAZPsOFeiWdce3svvaqhN393Gi7fFMYDF60h0xI3Vy2J6KyA40Ym
Ez1XuLYJpaJ9Lx86rFGdn/Rl2E88JBLFAUTNomJoGXn+d/C/7TFhhtpKhJcQwLey69gr8koX8jfm
mh7bY+D18qfg15DqLrdBRxLEGks16F8ZDa2t1xYeI7FgYkLfX5HGS0LHhyIYlnzaL8bIkdZ3GEaC
XvNhkPGBgUx1a1AYrTLmfMllRERJ9VX4UJSfCAbfaV+pw78SJetT9ZjpliAtVXRFalaK+0Gzyqm1
FJOQJiB5w1ufzIaxdVevIk4DzIcoSmHrx9ZBgmtXTjkKUmlSEd0+01iKSYwMfZJ6P30WrzOP6fOP
YESyp5ZTmj8DBCgSyf8G9GAfkY8BQyy+K4jRZwVKJKjMky7gpv/NpfCUUTZeUrCn+7nXvkKZNV4v
nNTd/sJFFFmOOll7z47erbCMVNdcxhIVj3RLVQX4Z/GoUGPJi6OQcWu1Zn1rn+qfEgv9bnI1xrx8
0rcQw5kGPGfCsvaAOyF3q7DNTT3A92uC7igzZ3oj5uLViBgLjLD/CxAgOXoMfaXSTaX57PpGbNap
9nh+qmURkH+bx0mOB7/XReeHnGV78ALQsp1MW2yQBzT3g78zOeymCjAVuSzI1sZHjtnBxP2ZJMW9
OOhxkW2HrhFuOB212fY55RBEqLNqjWRJHiYZolSrg49rl4Y6HyjOdIACuk41IWa1AJbGkVwjT4yJ
U7J1TYp850bbo/5VzdsAYFPdP83rmWMUBd5NSKe0DyGwJjes5S7AvYkBiy276JSsLxrg/Nn0evxe
bEOJhQlFMHTDUHKUHSVGryiiihPT30Uz1sdlqylLvyGYA++qU3jB3AQd8zsjZiM+XIocTVfcSMRG
D7xqEfmOCCe/Ztipmr+bmE9Tu+HgR8NLZ48tkdeKmDH+PzLkc12N5cVV7zCZCpghTOdUYJb29qI9
ePt3lF3z0G37LMJX5UitFOdvXvsiqZsIWnAkkyx4fWEvXufElhNimzT7ihVEHe8Qz3olcRYg3SHI
n4XswFCYv4tSO0tx0mfj6uZfJ4dUPKCGsJlnpsIwMPktldhqoQpDc3pC5c7HMbBeDL9ssnpDMOFO
DH+SPaCSfmBrYeCNe4vQAzoPVkrGthuFKmcfqzpInJi/aQ2Lpg7EoVG9rVOSRa2mE6HFFT5RkeWz
BN21py18nNNmfWhsLHNK5RPe3lZeabhiJmSU9pluBWKdRbww9cWiCzjjBvBUqf3eibwnxfOjmucO
gjcUJ7CChoqfowv1LGazHHnrus4NGvWiqTUTucSeb3gYhdMKTZ0cAuXYjmnhwOkVX28aGIjXLzXV
GqD9GQl8O7MbnAEHp3thfvrIGApjqsmtXt/PGWsv5jO8I/KH+CpOfmRAuPrwAuoP3p628T/K905n
EEAMvkn4AE3JIGIVHgKJtgyh0pHJgVDK5LNf39ArVwQnDMQxKMdXSs4DdYln+GDk6oGwJiPq6PXl
MOZUBs46grhMbtgGjUX9pQVVrND3IBbjEahBKmBnVCrbloHLM34uN9OktZLdtxfTfhwe9T+z4ZTY
R+Kh9a4FRCef/jZAYUwfbG9FU3IRL5rIwwHHhfyeUHXCfMrNeZfWWqxY06qVhtKLv6SFLALgZQo7
JnL74Gmvq8Fx+LfTlGsoh/XXMA9MVmsNMnRNzwOZkDJFpHVfDH+hc4pbGgwqgruF3BizrGqhJF5f
djMu7bT7ep11/L62u8m26SdQ/rsNBYTFVeEVKkhP5VyRbfQuvASGX8KgcSL2aecr3pytKoSNi2c1
e8PxZ0wsSMhkF84tLlDlz6SUiMxng3m9GjVO3CbTW4m7Ek9AIolFmKm1YcFSDHdGzpC1ppNwvBNg
uDqbicII46yZfYFJTCbKGm6DP0xI00C18+UUSJyS5ME7lyynLrvJFqJ0J0x587U3us3V8MRYKCsq
W5PktyAEishOGm/btOMOxrACl+WKZkpkaPpqG8tqCKq/kiY71JKo5eNhOLtysTBqMTa+FfPUMxNA
8ZlM2yCq6ToDKuFEmFQi+GuK1VQBJApgw/TlDtxJZftUUyHvkycThV8JTC/o40RgkgC1uvaBMyKv
CPn+VEouYHYfN9kOZCeMMgHUORYd5WzcJnFuVKVy8iQ4nVCzF0hGr/Z+ieQXm+5kd6Ys0TUlZwPj
x4vOtwuAGxIDYIcsg7Xr3x7j4eDtVVdlpE0VgWuTMTDMEJF+rEK3Q86l8PpetfwbUiwHBPHBe4g1
4CM1p2fvL+g30bL71Lu6XKtO//Zk8dXFhZr65Hw+jfbJo1yfn3kSHE3LKVhnmUZFhBaQ9IEiH6iJ
UlFzxLvOp3GwwAZShk45TKO5b0rEdtTqWywgg0qxC9lDPRYmcTsJgde6lJAo32d6HcOzkCGUb+Uu
OmyBxdXKMQTkRX+34u+CWXlcEmdJmRX4RIB8oE8skPoVMkRv5VanWhU8tO3RO/cxe17ljtMB3DZb
BkKQg1NS9z9vmMV8qYr9/zZXwFp2Rb2kOLPGR6l7X0icVYQwdL6CZQ0nDmwf9gEt2f9UgSF6p17w
KrOkFMg2NuAa5nmRLy7DXh5meoHHtIX6hgcjllTL3UeYNPgOaNwZYxQyhIFStvwy++FRilGo/41c
2WQKYbPmQA2zSMppGecX1D+JsIwEv44Q96x6XfLpqSkcMgsBhw0bhcgJYDuJKuhOsZwC1CJZvBJT
M+QWbTVqNFqpoLNi3MFf4NRpjc7sr/TjmX/QW2mkVMYkDOACVPLOmaAjO81jRCiR9kzKvhV/8Hbp
fSybc1xLwGrEg4//4h8PlIPmFpaXVH0y6EIlyCUl2NK7nmzwdwSX3541t2KlZn26V1JsXuPKeA4K
qx8lSBhepx5bGBGIeStCDe5VJD9rZYOMb63rS7ttiQBGKzv4HEemzb7OBL4KOOvc1nJRpnPkCeW8
sYpRGO3M7uaiCc6e/GKOQw8XyAe0chvP5/5ZdXR9213U8/qdriyT3B281BU5JIz8R9XMEfMaoQQM
jQ1FieOYRxPqCjUFHN3oYoVLRKZGALgwGUwRHVSDYJY7yH7RnRvfI8yz9QTj9bhbRhNDCVpUlC7Z
H82rjwZgyJnjEo/pjMzpt8atrZDJIR5y1NZGofR8quL9gHHjCRjT3X4k1y8v1v3TRuL01zFVDLN5
2bSc0dyZzoGVg3xlxA6JOXGcknRwcDeqoiU9RLpl+KG9BIg+TFFg5oH1YmEea5h+mAf7rcVLzwi3
WAFYxJzwxthuueAF4u6UhkT9vtOHunfyT7ozC12fLholvrrOTNkArl5jf6U6jKClat/EapPRpdN6
Ama0HOLdun2LB9whMvqNjVBIKgzi+RNrw7hRowNum0xRJnbMvFPtZpSlJZ5/kAyp9BBwGI1bZlaK
aPU4jApa/KGzUnOnMIofsVMZ+DxPufAZ+whZ3f3A9FY5Nb8i1DHMEyYMJBO7et9MFdhgUZLV05Wo
1TVXlxlp+uub6oTjtlfm/usjgGq6U0LCJn7OoBNtcrxLPdIxjQcwxesVdk7ZiBBz4GUNuHJ4Xrcx
2qH1qUpwmvVFPVb6W6FWiQNQd1xy3MMwCQfhtlX5HFD3HDdmtV0z9nHBMvHXP9KJFX7ABZ8Mt9SK
ExAyXY62Euaxj4RGQCuBRPCZwFBWeNO+cfzQW6p/hegQBS3j9G8wBuYHvOWffH0acRb01guIfvqI
XpO6dAOmhvBHRgBMUCYXrVe4fMCrO/Eyb324yDyDG13wPXXqKzO/YUqFeBZ3/iQQyqBK/VO7uiNp
gGfckUH+SMGujsFP71T89Zc7DZLIrM4YbgnJ4ACzkLr0yaMRAHA4t+QssURRwYf4+ccv9d0dJEom
T8GEh1nb5q2NO2LxzbBz8lsHhSxK9wkF/jWiYEkeH8ntqZgT4IKfryvfqZZ+kld7fFSyD3YKqn0k
PlE0bv8ChOl8JqHvA/gR5BsE4aUlfjNTejumZA6nSLqSk8hbD/myvA+QCuAzY44USttsnZTwE2CO
Bus59sWxOjQCBQ4iG7dm9qT0EtY5UnuuKAqUZpLprLy6FDwip5jqP1U1m7GiepEikghJ69ADeu8s
s7aiBEa/0Hklk6oAMsGjNUc+NRR4jtU6nzlPIyfisIaZhsNK8KoEw7/B/1iDZvRYth+3wpvT/V2e
gmUSrI+bAVIe+mIlHrzzvg7Zrt99ohuo7c07GKKXxx++fn7hzfGS4vV4gwNDWrnmiJ3qoQphDOly
LwJVr2BPOvopQqO3WEr0IaaLGlQKQBimwf2aNQ9kvQQoaN/rVtz4JHAA9jmcgcX0c6hRAWVxPNQC
vl0XoZ5yWO+feOFCwuWrMmbxnuJThpw2zWlLe/FCEIatAcnOh006NsWxzbOZvRjh9RUPVHl6S2aC
m0O2Ybue3dKkOi6A5iAs9llo0Zaesp4Yuq10sJZWC+Af6BGFQgFQFtz6jYYNhBuwZEzsYK1OTWqQ
D1CGjncUjxC7OhaZuGRggJP0BMgUn7aqOCxOzL6yjDHVqFD+fk1YAwwIsklCojXNhmnmCD7MHPwX
W5RrhNxpWQUvkDCDwizJwWEc4sKVdYH/Sy8gDoRtGtHUL0uxa5jiH6NrFMpY0GiLwVmQV66ubBF4
Dezb5HG5wZ8rl5flLasX8SUZaRlTSV4gu9Ot1K789het6NgVfMZ2Wv3XMyOX1CU62fs9pLRzgAFg
yP5XARtsO9+iEd9Diyx2T+ZuvDI8mpziLNwhMiW7HEo2mq2+tJaqEg3MH1aCLcNg056ojY4X8PeC
dEA8xNoD7BiYDc/WmlVoddo0RW3QdsFJm9OtERErTYth4JxlEs+Jdpr4TcaWeBYdH16u/WAYXO2S
wyX/4TYoO6HTWI+iksJFj9cmg/Vk0kEGwz+OxRRzTCKNMyKKqIDsP9NR2FWiaFZPqlYIRwp34Ptb
3DzZXzrmHzYVqf4xZ51a+I1gDrBByJe3Ch8+QhvakvOcVmVMvR9X8je4j4NWuvF6KBD6jw1xjfZU
G4GbyemAAqXCxFG01xy7+ngTcp2QqqX6X6sD4UAgj1rSGJDmgAM+nZeoF5iKDIkXuw0wPVHsoxtu
RQwdXYu9GTukz4JQTTDQG8LAuG7tKuQdQB+zfRoVX7+4+Kpg6xo5dokIc8xnMwldZwONVbjgZGFL
JFSbjSB6UnLsdYbv2EV9oaL2ERbrv7XqdwNR0hpXeQuf1IFPojSs/TiltPX2ipt4+7hoXVxcxAkI
UcRgtd+e14RSE6U8helh+tuteM8YeGJltR+DSB+1++rL4WtaUUPvpQrt1G2O6CjEvPYVm7FP6KDl
5Jd3wgAhZpsV2BNlydzgid5kwkcOqAWTzypQufqaCJb/bvBUM3P6v7L4XnbXxaIEy0iz/lNYa9vO
Vq6c9P7sb9dWDxH8BQxbvqo0o207hUXkGzVNt682sorpfTMNFhutUW9BqQs7Q8AnabFNpSPf8RRI
ioDXMbGd+Z4YTbt0BMRZvSTukyP3WaRU4nRDYOSxvwPEtijWcMBoiV2J2qADSrJpiQf62kmDyHnP
BhVhjlgXLp2wzUS5L0ivAAcWga4l8fySw9+viwerB+obPHbbKtzFYFHJnyqLQoC1h3b9mEO7ubcc
M6OzAcsvREr2hWM/ydCMsc1Gc/5UfADh8xYkHo+VFvphAD9GR2pW6y/mJ+46X5LndeR7A0c4RXSv
pMOS039Cmg19e1g7x2SXfm0gIAydgpZRh9XbynsfIHLLH5Sq5g0DtD0yCj8jW0ZYAPCEFOf0bTbe
vixZF3Gb6vkOILim/rmUcp3VdM9n3nnYErg9WAoZBV/VrX1zV0D7yXLjMjiFXcosOdmljpq7vF0q
Ce1/yLlclLdVgIZOVBhOL2jPr75a10eKOZ7jf+Q7inI0LMcXPMMnphzkxs3wc2fW8nA6UDulS3Ot
TFw7lZY3L54yaEoyI5c6B+mz9iU10Ta5FR0H+MzMopBFPdkKkIgUD/lNwh742XV0qmKndbp1QQoD
YUoQDzSF/z1zYnCSMI6BkWlO6xj8DxcavHviuFyGzrX8I4k9Kp70JGdMCL7KMbNtoTRBPlAAvuBG
pGp06OAbNfP/p7TZXu8bfznsu6kh3pg7ylxOakJKU53AczPGdiWxd06wCCYgHeuq13K7Od3VXPrI
zvvZh6kg66+GKmJkvSww6hHn5qlgTaInUcCjysm+8yjI9oZ3IMH/7WJBgsVa02B52WlMinI/+JHA
0hkXXjARhIcDuftShlihUUr43KiSH+rCMMznZRFU//EK1lcQA/KxxL/rAOaK3CWS9qQ6E01EeAWJ
hX5I5LZXvDzjyXTKp4Pck3Bm7OCwQkoOzC3CC0vMhpnqzzMmIm/dyxRAUHIX4ovYqphuEMzEos4U
UI8vkMPKwolBljGrK3JyDN+8t9yCul3wv87F57n4k922bSqgZaijh33vh9zL3CmIBdIdTddmBLnP
e8wO5yS72LPKPPg3ztfveRrJZHp63d2RCsNbcmtIrDvUkrOhbogcUQeqqrcQPFzr1+vO9FQfcZ52
aBN584ghXp9oZu1DUqLP3BisIP+Vg5FkTwN7XV4lMV+KPDWgygH0Oe/RQuKe8LmpvdYu/iCj0g93
iaDXMzXYNAFfE41z+NHzvTjB11b8zNPxBmyRCdASDW6OAy4FAqItxPD8nO3QA1mcNfuO3VgGW3q/
BEmuI252PC6v+AQSxgSPGUDbbz4E2fetkayxp9zg/Dd0dIdwqcu1J+sw7mvIArFyjr5o1Pu09e8C
0OazPm1e9tFnAgDPmgSrps3lt6zSUgEMvIPXrqvlNFHf42ER+bhKwOMCuqJgoyQrqRZJO2HNnoea
fg+ii36lSRIH8X5dJGlNyaxsVXqim8od3Yl/jQJJfocXFeF2U4rifh+WMlunlpYcRsBCojoGeyTm
0GmgiTS53laSuw2UHtc1pV6KlJ2KBB9vizpUmX+ILKKdvE1fjykmX48bwGqAXZ/hrLk63i9qbTxJ
bjBNjgPsJ4wit46dFGiT5Den6sMW3e0jSacvZHrx27+FnvgJDKfCxmeKxWPbdzMtQ3EAL8F4KDzw
GuwT2rn9MGb6wEwa9GaEo2QpOUl/vyNNhtJDFLGTv8xNC8sM/ulNl99F7MdmZ108lrUNyoq1Vokw
hrfd3clQW9wesPx8Uy5Y4NZsSvYnuWxKoAKOGsZcfQechkaILslAAW2xU0vO3rKKirb4c/RBfdeC
c3M/QpdF5n0HuXLw1luGWJ5kXVUBK/T4vwQnTGFUBijrcV+Q+l/a709pFA2ljdT0hputp3tThE5H
8HxrSXh9g/KrdUZvj2awkgirwV9O80Oumuez9h7re3NP26FOr1fx2E9cfsXu8QeWVxG6JNs07nje
9jvbQaMcotyT1KTq9dH/KlnZFwMRnQ6rErluQyZ/QMG0HamTGm/zBNYMAQxGhLGGB/69STLBJXfX
KfCLLQ+nCLgYwHSuz/14NtLT4I2swQsg+tuj8y53jHWV/P0rrNvguR6hjIhlZMzolhqkOlf+VMMu
mcArbHh8H2Tn2q/dtHG5anm15dTagRHTzY2nzTzUn2a3Yqw+KDcFFwGiGZ1TrBUMP6AMf+N4Vpap
6EqeDi+wSZsI+dPG6b5QHiAwkuPnFXNu2V4bEyf07vOtgEsZ1XBxS/07IwZ4ll9OvAUKI2yX+ANt
HjCtK9ou9HhiXfwThZ5XZy3mc0V6aKmxJmJ8zDIe3ge+Jz5VK8Do9s9isXImIR8wxItTHxvSybGW
VHfJToPOSnsqxEcKW6m2pLxCNQ+lb0cQfVCb7GtZqXaxLNDJD5iMp98FvnTwVSnUOoq2BxE8FFw2
aNa/ZOj1zYEt1joThZMWgMnO55SEl7/xb8rO8PfL50wo6X9uZFLiyiXUWnZBpf63qHCZWZArfrs2
lYiJHpxQ5cKTnbs42mQjOeFy3SNaR3cm/5J1MAg/DBepSklls+jFVz5qpS5GmFG9QOcCvGLyIoeA
GZ5KGwbg1ha6Yx0iBbDYYUfmU7qzh1cXBbSOZva+1ofNmw2NXwO30k6wyinxibW8/0AVfsqKbjfL
GBBR8U/ZHbsR5TBO9ZuBWlbWvOwcgiixbNcawcZNlhF9DoifB9REewElBmV29JvgmKP5u1I/zV0m
opUlEGn/DWaO/0eYC7wacpBy/hHbcG34n2SheLGuL9XP+7brXO2JagCRKAtc1lsZB7/DhNWNbNje
rbBWqOqC59SmA9C/yU3p+vldGYDpPS6i6ZOnGZhNIuoEqjulDkJ3dE3LoBjOuxrtqY4W28EdIz8P
c6s6ZS62ylisjXVqAxv7cMlbkscv41vu4g6dncnE+ZhUW8jtkMg89qYdWIbLg1i8ps6q91Bx+DIH
nWmccR+X6dn7TBnGd5w599qPRCDM8wMJ5J6twDlv0okyQiqHaPAGdGVbhClekcDuzV9eLyZCCygV
Iio/k5aZPfxQRwXCc2qqt0/iYTvVtOMuqLRjkkFNoqmWkWOfGLigpw9sH9v8gb5Mu2cz8Us72nu9
HVg7Y0FsapfOpCA9a/jmZXDhhYp6SgByexB80P2/t7QWDIz2/EWLtPr5oQ1zAD5nI0EpZI4AHUGg
zGdlkAGuEaqV4idRMAnivSZGMUaOi67qt9P38E4BmhmBCFqPx/9IcQdCi3k+4MgZsnryyEyH7h1Q
GjQSwu0p10c34oHOm050+iYOAyafEKxfj7Un3TWZ4PsxN29UcOoUtdwQWT3pBV53Fhh1YWAPcHYh
IuXp7JTNV8hXX88b8sn7Li4BhzoUgPvMZgb433JJveLZp/QqvoT6Ldr7x5DuUbBmtj0LDZoxxRpF
XsMSJIa/JRxQwg8SIOYnIqA1Gg8pNCDZTLlgs6O6ob3ZlTgP8EGTBdIVZrE+6pybb2D8U/iQpq8I
iZbwwSbQ1aeMe7hLLdzwi/pjC6fAd9B1Oxh6pfZF3phfn6pAtEpow8MVKrqf90CgjYAbAFrEHMEa
hSc05BajjMxpXemzToEA9j461GzVsFLzMxODBzmiqotmx7mAqcHrhFv/tLucHvsPkzIj/PHIxM6r
Aq5SW7Sfgsxd087LqhrtTAKfCYfIJw4FmvKmmsDmTNU7QOu6TMDZf3fGK2CvoMHX2Bk8CREy2ObW
ip3fUS/83qDI/KVcCfZMf2S3VJepJhsPGJfu2tk8XU2M2kXllvDa09EDJ/R/I8XB6dIf1kk+7qeo
igpdykt27ttcXpjGj2dpk7X1zFWdSMn1WGNS+tte54qC7eWbg5LyAjwn6bLIo4VAU3d5Ctdqtmcv
2LYiSGdiBxaWFH3xjRgqhGXCGRHvB0+GbhJqzUQcgAzwUWVLpjFs/0nd+jawnldRd2XuyE+lweE+
nQeIZ0kcYyW9bbZnHJ3ES3etFKDHYbhq914VAfKx/DDjC3WwdvMalgu9Gp7PKdNZBNALcLMKe06n
lvour5BX+D46oHo+GhD7B87KHi1Nj98XXGLT4yzPz1Fg3PQnLBf9VnQ5PS2k6EVzjsddynobopCl
oTLgGoKGoWpYTStd75I6i8+Gu+T6ZuFDvNKhEQu1Fh/oovqHv8dNLSzH+FraZblxQI2vXTA924O+
bzyRlMtE3BIa/H2bgKkQGbalJ3niASxmdXOdgeUMl3OJHmqlbx/nMF5hXN+BWNkCXlVuAE3+QVMg
/dROnaJenzkDhJlakgVbuXBm6vWEXQe8SFfTH0U92RljZLty93Cudr9DUQhmYbhihi1W7N+5ZkFS
uFyMazCw3t7F8ALl9ON3fmQ8Hq4cztnpp08m9w4kE9go/KKUugwnCPiDacQJMh3QB/aH8vGaWBeC
FkApJ1zh7dn96RRk3uL+QrIAY5uNYHWy9hkKneeaGSWmHxw+6tu+kLZznJpmOZsoKpp9mIZd5wd1
Ah/YBqg0aTolXBDolme28dEY7ikr7nIYTJESGZEgYKcVyRHsJw4R7Xon522VbgM40r6Xx4QoS9oO
SemqIZHDaY4V7mnm/G5UdO3+yFPAHqN1fx95Aq9fQWxSPixSN0ss1fFhwcX17F+3goapjayMx8Cw
iUEhJ6Q4ri9BUe+IRGYaHzQA0ym5T3WhZJrbXBtPBuw+t4V1EbNkzJb2/+iqa+pOOC79s8oLgJCz
7TDpB0jpB0N9nK3GhaaJYGVCkeI/0mN17zMA3QuyIibhpHcZZNEjX3/2VjuLIZz89rtWXeHRRVzy
FaF0ZuZfSEyyMZ4kMBZMyiC7jgenmSbbcds4vzrGs7ZuXy6b8AeMFzAp/hZYpyXlOqkvHBCcvOZg
pOZ0khEg1GM7G6651/LuU2TYDUvmEerxM6hU1PvdjXfr3LmBzTYheb3qtY+kDqN/zO2HcOak15fb
nbrJJtcG0VuEBiIRCYh0baGiSgR7Xw4DE8IFOrnXKlbzrUWOgt/kyDOFBwoO6/tpvl7aH0pecZrd
cP83r8vZAoNfpimZfNqgPk6MJ0KwIqFMLwSFEd7aZSGQfaMV+PyxAwOsNorO01FoIMopv0teg6NY
2FEUi09BrNfGtaClPtz7lLy882AFupXvxrRutq8Kf/T5AhN1eSsBF14e2ygBuMWT75os06g+8vzd
AZwGrT4W1q6Sy4jbDR85OCXLYcH1XzoJsao6LGnSXgvFJd0OUlbZfGsgMpdn3xG1xiCT0q8gVh4a
s0fZdwpyHf/uwQ4BVWH0/7xll/dc//bfIjpop6Skf/gGINmgzbFykORH+6SApdQVHDomQ0KFfeC1
TFoG8N09GAZifq01+RxVyOlP0SgvHoNmQ9vrDoGukjvi9xRa27YLnnv/joP2akFcH3BE4pegOJ6X
QapDrbBTkM9vSWVidbCNlb0muiZlTqEzYHMxkz9FqLoqruQVgRUy5mppC0so83V4ml3NAUz7ydFK
lYliu/jD2VcyowMH1dpIfpYzS4bEwjYKOhPeP9rseFQbRGOutqfSiWF56XP+Y5h+KY8QjwVN/vuu
iemdVEc2CMshwdNxemjKxfAqfTyfNoDEkPTw9dFIyGrdKU6vIMPRqnQk4Wm+5s9HvK+jl5ITPJpL
Ax50QzQTLxchl/EFMv3tq24v0iEM116l86vch4R6tOCuIIXOyQuujycb7PLNWReqasUzKI9TVzz3
s89qxwenFwXsz26HztfqmCLSbcaHTIop5ZZgiqdk614MCcW19+mABmBX3cG0ck6B6S9+WdGVlX5V
zcj+6EOGlJqOZqG8tsdAarM6E4bbA3393UJLzRiYSFjQfzNBndy/dATAikN+SjpBblZ2Y0na+ls5
2Xs3YQBfnNPwvDsE/niB1+GCCXD/Q0jM1aqYCyrMIK0CJP2ydB+vr+fqiGShEgBlfza8vpQ1Ceeo
Mj9qi0YJUIHWPetleBh7Uiv9HHOaJRBtPEw0v5lOVw2d7S2y5gtQbUFf/bK23SevuaChkNgY11wV
t0URzPTjzxqAv+SRyo2pQpp+nPWop+tmjk7H4asQXma3ARMAlR28M2avHwDm1OznBSpRYIUhb5Dc
O4yv2y/mivkem2xdnAyhha/fsF0UigY9coB3KG/60tkwzXaABNCdsGHq+JKxytL0fd8Te/bfA8pv
XYQjUGrmFoSXPghkm2WcYVSsUZwDdN5wTS920vcgVs9PcFfHo1+AeI5520iMIWUwiQA9m+c0U+OM
uvNpJWAO4v060vVtqfAsc2HEuYyRK4SvkaFTHY4PAmtfuyc5hggDuKet+M1DOOJhV94gqwIM3gWL
EG4jFCKd8thKV2MmtVjkCAk3Y/ln9tH69JyB6cmEErHeqlD2jsWez2OniI749F94L8xpsPUc6RDm
QXA/mtSR2lL6CcoLEJgmMZ2812POG2LFGHXVIjO5DJeWuq6aNDXecxQ+Q5f0EHFPk4alx461VTcm
3wtDz57k4S/ms5gaGjeLG9/aPuz6YEKK1+fyy0UM5seuIoRAhJDol7KL1wHFWXhsfTLBDMu2C5ye
PmwMO7bq9dzIW8iilhzsIomRitMkDv8ZtMB4OWcqTCweijY85nu3B8/UX0OHKRTigNYqK1t9oImY
Vdkx6sPF+WrGxvfb5SwkXHcOdc/OAD3rcz3PYIY23uNhX/q2DDwFZha5aytf4pX65Rk/v6tqXkE5
4y5L1uA/A1y03j8nwxmipEdNG3ZYJ1PUaQmnJkNxpf6Mky1wVDYstr8qTXpyFTM//NopruCKvEh/
AIC6wjGYdc9zS8r0Gaw++l5oU+HWASIk869wA7UuF/K5ATvFbQwlbQ7Dahe8v3yUBRh2G4fa6g7o
7gHd7Yta9zJVr1mi8Vss0f9LnbABnGkVfx/PxJUdn1D2FqS9JXrK5wm9ySJtzbJ6g/Mk1G94Gcgq
geMLv0wGF0QsZX5XjCm+o3J6wPuDqw5o8I0HDGR2Bzd5sAxQYoJV3kG1tW+QpCnkaeHVZ3AhhiNQ
HlzzdD4QFCAASfqAk8lg3V9kFfWOWs2++87pbbDIoiDdDN0z4gC4v76YnOGn9wy9YaF0DB3hv3G9
AIaQFIWyDRyIPB+oWZI0CiPsEqQs7s02NmPzZW20XblDTV57oIdSWQ4NKaplvoSEcDmvLTwLfvao
jQXBVvYBeK7TT7U9OLQHhQ5Vr42SFaiZRKTwA1MX9clOf+o9wZ6J3h9/Nu4CvSVHfA9XYA1J1q2N
9XmUC0VJhETrYLYojE9Tp/E0LnGPLWNXH3+TRKKSoi+q/WRJdTCl6azxVtd+yfZS+VMxtRR7UV/2
Q/seuIZ61xmGcFwVg99INkxtdhNBt9iTcxxLyAvhLlztDzIbSflHMWdijSYZeQZo+q9NpgWZI9sW
9nghEx6kC8zVi8n2NI9zHYvIpHL5aSLj7zF7aMQxuX/jilxXmQ3jEKe5+iqsuvGZF6hpIuEHtQQt
0Ddws5LS5lQqPs8+m/sOwa6Jub6SgUS6SKlRSP3hNKZPaoZKBDiA2Xc4X9rCh6pw8tRsK++Yj87u
JKlad0gcyWbESr5aAYWm6t4RkTr4/ef8/vX8f7D8ZgvgwT+35TkhxdMp/2my9xqrJ1C8+DDCL+9Z
Um2QT4JcyHvwRCXd/CS5RmFYtH5M6JBDx1BOBKzpoZrgS4631U2QStN6sHHJQukYijTDJ5f1nO8/
zUtm951Vt9TaTMLvostXx1g01/C9f5R5n90FgXTqnvr9R5oraUkUixO9cB9Ujr/onDSFHucs24VF
rAcQnqZGvE5ohpqxnmiXOe1/g286L9adKLV12SLwZt2cnMd55OifKGmWGHNsBMfmXmRh0HjQphQ2
M90lwdlEeD3HmYXZhOgnNHGI0CeNc1yGSni/F+PZvdjQ7COkTPApskNRDlra6n0+vmh+xYmwJfbY
MiruT4JI/S0Xnne1/mWNRWoIG5O07cAjLAdI5GExRlHY6nts7jCSMEL3YwowYMcwMMQmcUGkPCIf
JlOP4RYtjSBvkbbrsRUbKI3/pzHPj+A7ihutWAWbIOX1o/u02LdQaWp3qsI+O7caSZYENFn8jsVu
1tMywSn7DDnJVF9AX5Lb7ROzUAGfaLKO9z/oxVFh2TEYJYCnmyGyuaDTvsq0CW7tXjo0gObuAdsb
LLR3c9mqS/oJFwtkoCRQ5i9T7QotE4ejzkHCDde58XWlYwBYaEd9mcMyYVFhbwyswH+LrdxjtJkA
sUudCQosGgFYarP+PwdikQCn9h+0I7JK8ivRPqLTyT9WHDxGUkPjlS2UOn9emrJLal+mu++00ZRj
E/axWeAZf/1BXAL7PIII1SI6c2wvN+WgcWe9NPgfxqRwxCsH2rd8UXT9b5zdjCpkyzE/sBcz4SK7
2ySr5QuDfVp1pz6yMYONzwrSsbF6kpvijIoonAFGGA8DuipvkXKnef/Jaga5kn55nDrXJv7JZrMM
IetiivxXBF8MVX5UCmq31aqI9EKO0HBGhaEaHgDQqHdF5mYR+dJTaU5DEWPRS+Vok+nAx1da3XIw
4E34HXn2FG342Cafy9yMYZ2xTP/zeCXjfiLx8+FH0fu/oMsSFdqCI5bS6TPg4HRDWN7UxniofbMq
vmHDDGIWHYoXLHf/SGl6lHIJ92q9qzcBPGO3W/m/YSCeSOdiCaUnyh5QLUH/bz4cUSfAWyK/ojPJ
BPpg64RMzOQs+wpQMc9E8dvfukWwTC3IeanVHTVO0z3vEzCfLlr4fK0cZPJPoiGngcZouy0bmeLP
ZNEEwDMLmWp8fUjd3tJGxV1FdZQ5FhCdubhW9FByNVjlV1NGCAYd43ZGZlIdwlhaB53/3zcc0/gw
5lY6zmJvkC4purvzUzEEfUabu3TcPrrBOMRdMmpLPB/FpxN0L/Q83kSI/Y0u9OYGYcd99UGxEI8n
IMY9eIysAeqhWyBrBVnxOW2m0r60o50bjIBZD2/X7r4y2Qhg7S9Ts7nzb4Y6ZIShtuNgHuaMDcyh
J0YssED2+AqfcmBCzB5OlagXZyY5s5gMEwmv51oVzdU9n3AXRJxG8isNm6s2cLvVP1+2sPwNht6c
BqyE2Aq2NKEwlSpiFw7ReNckVIUzqcMXN6LA5gRt4TX9/tVDhTP+Kc2I7ru6X4DpVasMdV0PM3rx
SbpALwr6M/WMA7/hkOgV0K/9W4jgOXkd4XFz7hLi5CAyAoQMMv4nq30cV2hHDbzbRIcwy7lvh75H
BiD5klHvsw4aVZ84UD/qwHFV6dbwbKt8rpnLaZZkNe9BOMdQvIQd4awi10oZvGtc6WS7Su9NimvO
Qf8CsfsH3hRjSGZCRd+EpsT3fCtR81JwndMfMwdG5NCVYcHlQ78rfan/Vf4sh120vq+lW2g3Lp+E
ZmZKcqFf65lcHzQAi02T6jRMxjmUdojAQHTzzpkIwiE+Z7igtF80p8lzBxZ53zmWC0o9RADETI9h
GJE6wFPH0n9sHpyCCM9Wab2uJyYJhMYTirjAb+YN1jnBIoAryp0FOmGQWzYxdU0M/0ORT/QXXES0
uTfubpBgaILK6ySGugOzvm57kP+Q+kzlqc3Nw4AuF0hhH/Mm1AmkTUvyoiTbt+cQqbUvSz7SIluk
fhX5aeyHEqERObcjfhDyGaHzGme4b8v0iRt5rA76NppgYLaM/UPv9/e1pTgDZZUyKq6Rpc0JRXAB
OIo4YkrXGxGFMuyaW9o8hwgju3+ltA3wVl1jYXLj5Miub4Oy9kQwLh5WSs1jNYY3cz0sYdqEuyaL
Zaz2zHqT1Z09q41uIpgXI6B3KHmJHOwjSf3vSMvi7b6S2Bc+Lg4SQBbomcBv5LgsleOi5cnVu0Qd
mU2hJb9nypILN3hId8PvcXXcE9MDRr2Dgxc6dkMYqa24ZRQltiew+Z2WPbOOa8VL5FS0zpgY0Jt7
r3AJCEv+yGvkHGgDo3nt0XFPRWAyHbl2sMnt7V302ReDs9AeZW01v/1OZr/KCMq2Y1YHfai2YiOe
MjLzIblkhz/FXukMEK0b2oWLn6EQ7OCXjIWe1fvcdhoDtgvgB/7jDXdUlrF5gxLjwip/7yg8Uqx/
l8i7LZWXq0WHtG7jwupod3uwfZyHaaoyHRSQAcAbnV/xTnF/rxG46vASvzxC7fXiczi1iGwGD5nv
Z8b/8m9+WYq0rAH5hgGtx7sFdhlq6HI2tyM7Lx1f34ZOXfc//0MQt2n4NtdJXna1tB11JrXTCkOl
k2UK7W4b6GSZDnjeSyiQdA3qRRYwOb8qC7jXwi99KqIOvFPEdigrwcYJaGSgnVmLTZp59WrOOj3l
kRm/S2EeV2752veuHso1Lw+tfR0DneQWoV8YcarM25bbVW49hZIkjAhgTkzNnBAF8HZ+9tV6OBBn
YgRGv5TTHae2bwQUKi8R00y70Svc68asz+l8wirsGU39ihIF3tFBOaHLRCAl8Y/moVuNc5pWGU/5
hXv+K7HN+j0fFd0L5MyhmZFOHn7S6C5P+Eb9GciJwTyJ35B6B+12DvYT3WE0COHIDpT4vHC38Usw
U5S1LSRJo1bqsakJ5s1WRvKzMoCuDtkUKW6keH8i/u1rj7uIYx+HIcZPpxe9XeTxvfnpE69Z88qc
7PkP+zsIy3TUbX1qt5SUc6Al+t3fA75FSOT+NwadNfA15xL/FTQTBE1UGrV0dr1sZhBQYfAlw3a1
XsqWDR2/Ozs5eUrKITUaV06IHqLWwKdh4F5QwVlljabA5KDGT7hAe+F9xVYlqivN+XS78xxfB4XF
EUptazFgOowfN7eKu8C3oYeIIcppI6pHGr4QujrECg0fKFH+sdVMERuh9a96AT71F/4L0VTq12n7
I1zHfBeKHlxkpYHwxJaNNZmNZcvrNbB3msGnHgTx0YXyvOsQ55BbsE9TlkEgvH/a/673cZCvAk6J
Vb1AErgc+jUlBBuKJ2cLglnvYmEqhlzT6Dq/D2tAgif5ifPsGEy4ASaRDvNytqJNstSRkBmK7qTo
5b87khj3fSH0DUlbVboHGJZjC3Yo2HmnPQ4oZ/6NPYd/vrZsTUZWOC7r5glpfqi7MSeW1I2JJuID
DLwpAWvmHMJUrB7FkXoDXiNBras+GsXESR21YztTNV4oQYFjtYpYFLgTIP9e+SK9mSgTK2FlpL06
4XuvrPKbSFwpQFhLzHoOMhsFx+0Lp5VZskY0JMwxk+Ln83vLOPHjglQozXb+VyL2LuEXHiItZi8q
L3CdfECz+Lkj/vPyzjceFUV51OzvMsZcglmzhAQ3jOATDSL/4b9fSyftTg11BGqpNYbRcVXQRoW4
M7CcJoXVJE+/F49zRROo/fLmycFjnRITDYZ8dPhM4F9N4+SdNPAUaQi++rULXbJjyNMtWOSvPEMn
bJmnRVFzMXUgCG8yeyZ+dTqhYI5wYuUsvMO1Ed0aWptzUnYMe01rjD8V25LI55cN9IhSS0eJkftV
uoGWZd5HcN/yaeC3JicSQFlqKNxD1p777eup4sKm5dvKpo6HvGxwRjZHvr31oTeiF2aUKhrNKGon
bHVVX5tnkJMCEF/G0Yqa1gdUYpNbBpmO/6lnshVZyzUnQUans4VjnOEcwiKiSJXbW5mRu13G93j1
eaViVGBUZDaVnyLxpsx2AvZF79avPCc8D8lWvnb05LWZflxtuHJnfhZJ9TS0aDR1SgnZxvibXxLY
oaY/7J7Xo82/W0rexjPBdM4jvr5H75n1kMSjEVU8brjZpgiAQiH3Q6b6AfHbbiwjJuTcg/3D2cD/
ac7y4GwVwlcUMwfBWI9BMn7oDJyVVazEc/LoO9L5lIO1TY6hcD2+ybAF3Ac9JiDqSkHdV2TZOH1L
6yR+gHoC+qQX3ij8Ukqnj2phRslg97+jtmTQvlOOuIqS0FLPxoa8V3bQmEQnJ3YguK/DPrDLxgvZ
brtxB1fdxn76LSSkplGEj/Re/QgMRYAtM8ASBvaK+NsUwyp9NoZnuuVzrUG6eF0pdtOsRVm9WgXL
M8SQ06vbJlnwCiZpuBwz6kW7SzF9IuZrkKIb667fAWdWWpB2wCtN2WoIut4DxNmsP5EsD3g+yBPe
0vKscza6bzU4LH50pn4a9YBkszMXFQH/I32XPzLtfhpBr1V0eQQoNxhV/Sk2oDmAdG5rhy2KZ8le
UrjMJHXAay9YshP0VBu3Pe6FpEeQqzHC4v1JU9sWOa3b5B7yJtEyb11kOZhxGmzSIPLLai1+fXE6
HlLkxw4T6QoFthtb5e3ceMBfWrJIGCTBlGbZhk0mb4pLoDTgRhYNryWFKbdtAVugtUK9SJzPw78V
STk/1/iC+P/dt5lm84fH/m5brpMwoN1FenFmBCrDodBu6fAhmqXDL6YMPzt0bV11iMleqfUi1JM6
67B7sIBNdoOmGtiKjhyXP5NeqSCvGa+qFjBSuDhq0pVb6wsnPhcDXZVA5LxQJj8Bq8sdiG4Y82vj
zH/ATeBbJZSb/kCuUaSK4MWSqQw6s/QmtGTwaWbrZ/+FL5BuvgvDPKKlURlfwQYQ7wF2cHXyKnNU
r3lShwy6xpzFu1inLNBGFBapBYYAUIGTHEjro82t0D2cM5LFD80Kc95iTulJuPXMkeyTTVBnk6wu
iBw+y+leCVZvnQQf18fdakW96WUE8oKUA6J6xjTKBJ730P3VDCnPVWaOkihX2LxK35LGa3CfSPdZ
ruCqC7NaVz0ed6k1H3u42oLhXdQTMkgaTarq+iUNFJ0pQmCtrZ2p3qLfY706u+3HZpSTuUCa1m7e
4q+4wcqmzwssJSeWNBrV36cinPCq38X/15co173gph+SltGBMPgGNdinjY/KPrEeUW8dydK1T5LE
wdaxd5QETNzoMXqyiac/wur5+02ueCniRq3keGu8OfTAlhxsMHCpamlyqtohhm3nLYZFsGjGl3FB
JwDqWiEAUo8R11PDkxqPHnh986gfPK7xBGNESpzE/HlCWekQAm/JkrOMwkQ0xkFmAPXF9fBZNUyO
MeQSvAoRpBUyDkErGj9WNEJX+bfS5Uu8lAiptx34zwyxwFmAKU2GK6Dyeaf15UXzpRFpZ8s4MadV
ZdKWa/Kud2XnLUai2vc2apPQX9hkqkNhI7YSlcncHhyKXweXGZaVBIRrbIcxyAy8o1qedDO6sAyB
g5BayNGrRwKB4oNibkDD3SdixJZGyc8eB+Ky1hQL6mg4vXsyK4KU3MT9LLTkZXeZ3yNxsR0zurAK
nGOJK+cUj0YTFZGx1qo8qb4ctRDBu7yB+28d5w6S8h7xjl5vHtU9bCF56QTW7lTbI1NB/17z87u3
2JLNXMYiaNug2HiJPF6hUQMw69hYo7xZ9Vm1o3sSwcxVcoMZ8N7h9NGTW9qGtWJfAtddW1O0LQ8r
gKMMPWkukeVSsOMEMUsKRiiTae+GvypL03AXAHWrGDyoHaC4/0h96ZhOUTR/oqJd/L38Nm5TH2Vz
8JAuF5ihvxkPaql767Jf1KAYYxogd0OxJsEbIs7D9N18hfw4wrWj9NZmeOjPnW+KDxpXJSikKwCm
YvdJSHivNl+ddNDf/hz5lMUnl6pCz4rQTWMg477Sn18YtpbaibfyxqRD7Ohookj+SFVsAODSiYQk
mJ5DJyFJyogDMKWUeWBgNep1Xe440e6DPp0Ds1tMMzl5JP6kRzg/e86eKK8iMvybZHvrwIOHm/Vz
zT+8quE97ALVzreHDkaWHPU/jYVD5jCqYq89RE+VjRBdjlNM6HBAVfHhOZCxsVaCRS7WhzDGuEPV
ghELQJ5TIgWPphmIz+dtFoTvnJbgaPITHko1ul8B/FWLoIvyC1tA8i5kZqkU3z6hkuwF/Hcfsl0K
BZJt39rBNFIzhdxdhPUgdqAAb2S3YY2+wxjBoLGTJ0cXCD0w/uMWHPEQPuKe/J15qyTcAP3XYMwx
nnPp1m9yQc0kghSjH+4pRiq+vouDanxloUe/iyCAoZCnI/Vekq2ZjDxFkQZjyOwPQHUTprkOEEHO
+COeH/js7r32QajUx7kxd81SQfU/v1uZjl/qjADU+0u6e6CsIvrLsW3T7UAjXoWtEpUzX+HENUeO
Er5XzWVWj4U84vFqyPDt4rMsAbWVjrNfdZMQzISvsaW/WdOcAOhqs0+ESw/JNvOLmYJvedo8Gakt
182jxU21YGTHV96Zx0eGXDgQA4BeAktIS9Y2aG6HJ4iQeRNDhiRyS7tTFI9GldPmwRoenWan4jqH
qT2LlfCjgGFb55RsTJ17KRensURgH30c+j8xoIzAeK0GTYRABigm64iEBFjHgv85PpX/O328sjye
ypeFui88QhiA1VCAtQ4K+ez1UAb8lRcuET9UcP9V2zxDHKYU7igS8TvknaFUqO21hiymQYt3R1qT
VBbunji1KCNMpKM1qdbnduEfDQvfoMVE9BLyJrFB3aS8O3i8vIQfR0fbCUQ7rmYgcYAF3ECwTbyI
ZgqHDaU6cbK3qOL4LFFYQ+De6ZdD9I0QFEO3hdMIUGZTfOnr4jmuL8EJue8L96t74WDvtwjsuzlZ
7U5sw2Pl3LY9/zVWqzJIZ7Ij7CEQrpmZ3oyiOnj9CatpO5FmhYnXWoUkkDsBzBwnOKosKXu76UJh
/TBJEM+dSJ71bZqqfbCvZIuQ8uCQgdJ0ajNRRuszWlYbsvwfxU19mzXol4olIBpwZzua54F99fzJ
L0SLQ5w2mmMXCbpbPATS2pWQR6Kj2xHshJ6gtXAhLCywXReMxs0L/pDyfolxyC3a3fkuhy2/6Msj
gQnyCadfpKLDiyfw7qsml+LMvhXl9+MjX3ejLY4ngl6JDyewWDJ5XuN9NoIk0qRuOsexLjfneL0u
qHeAJZLp0W7NhbNDnpmAi7n41ErxUdu6AXCs1/7qwLFPCxhj5skaBLnebnSpRluyk4HZOk1dBzh0
5fNUNjPA6/p5bnvLLWJUpY3U8iS1HcyZ8awqmX+/jU8FOhqPN+jsje7hopzV4J29gvBcz+lnMm4A
/igaZftPbKnbO2NL3I/5A9q4BljXCee4YZhq6FVf9Gx1fP40ZZGku/JhjRamhXs3SRbETJP3Pgzr
m+O7SLitjePP1K/nzH/AXUL5Baf7Beo1Ov5rhlmfHq33gUKYwMHBDltJKvEfCjlWjHJ7etZmeJkz
PzSto6Hewhcz39YDuk/61Lfo9xIWTur2ocqjkOZ6fra9ZjHdzElywoe8CbpupHmCbxCic3+tRHz5
cdEQIAqydOtM0ncf6AhBFcy1sxNaL7SkA7cSPUY21ota9EmW0P6k9JAmtqsI85cHB0exkZYW3YRB
0xZCl2DNwP5Lnt627rFrVERgr4D5pE43X/MKc/H1deX76PSWXaZhCRK9etHDK/4/Z1Q+anOTplq3
EZHNET5mtgQu14uy4ZaAOn3hyKujhWPhRf+4vAzEbWXmDFpPyf46jG9mrBXCduc/cxEWT08V0x84
Mt1zpl3fosonz5ynfK0g+pUGDOo07gwt6KW9W2OsNuqvqoHvYEZc1Xa0EDa/GVzzwgS+J4ElQNrx
OfQyPeoy15oEa7myxHP43MrdPVy/I5Kamb/ZPzGUCa+tbSWVPBKC374g9BR61xoAF6WyVeNjjVlz
RV1rs/sWN4wWDtz0ejm/k2XYU1t/jb4nKJxh/3Ym5pXraobkINPUjdbS43dMLV6LD2cqi2nE+Qq5
H2QiUDoa+6/GrH8di0VuQW5e2eFay4X7HwCrUzoQx4KNr5PEvlgdgNOiu00+Zi9Qf4UxAfdr+nyv
YiUEv2h0Hxlb1KDNNZzBhKrA6RpPBug1PfO6y5sH23Srn16aVbRIyWyJF5Jnka39mxkFbdCYix3d
PbQi0OzHkkR1i9qxwtt1TpMEAmljA64akG2NMfTM+IAQmH4dp05nEjHgElGfrhy9gTiY4tads86R
9bWke2m+jUckJAZv2YwbK7M1PXUf1plBSz4B0f+PRIM22LEvf4v8M5J5kdjQ85vVpz7QWH1WHA9Y
ByOIbft85YOyq1zSGnuVRvgVXwmnc4+BtAkxvng3A76swUww8LLcR9sLQO+1BCsBGZ6X561DhSFg
uPSwZbTJJmLikT/bgOzO+cjTtqMkX79FsFPkGGSkJ53Vo9QzMpb0Q40fJ5EB3bIOg8WbnNrJFs3m
jm6JOnGuPqEPsNaaGZknE5vs8hYoKhlICRwOGp+avxwyAY9gHsjR2/iMsIGAWbqL9bn7z2UiY9qR
7kG86ZfrwOnyO/FvtXeqy1M6wjng7fbzjXyfjA1hm5pIpTxy25nxnRV1LeCzIT3C613wZJCSp+Rd
MOuArGCHthD4uT++D1QmkS9YTGdBXJjXG3bgTfN1b1StXnCcSbgHitK3qC12KMDU+kPlSpXb+V0D
0MsLrVKIpflGqOH4+gib9rYenrchDsM8M1lqsNzoqpcI9iODLkGa0sHVdRGdJT0+s3zpxWY4BBjZ
aVLwKXwbyPLilmqeoheaw2FkFfiRgfOQxcUUiZF0kQmRD+eeRuy//fdPp2MSXvzO9ujWzyZP3K9E
ELY3EVGRMsrDGhSLY6vzTHUK8extfHz7d2G5ERBYroGRYokkhNrDmD5RAMFPV2V/FNos71dt1wHH
K1WMEeSfz9tzIbbvz6o1Pg+I7O+bhi1232qu391oi2ApRuTQlxI6uvwESjDvSSzdq5CCSwSmy1gq
v/iM4ug8gTxTiMVzY53sNXif8nps+Lq04yCo4NgDxAGg0+UAjvfOBrgOsRPc6L4StyFp3YVHSsOX
oc7wBVkWyZsCUA+2EpMgXroKCLtE82aQljo6uNYF2XLavTq/39Kmfw5+5bgfpbiQf683ZnkfoSJ4
naFfBn7nf/ZKWgiTHAwcuI8HQvz9ILgRRKO+mSzRZux40xQsAEyA3XjINhIGN45e0sAqMzb1XdJ9
vRcyNOoZNR4to7V20fxCaxnv3VnC8RgO09LIlPTpRyCSXnWGwds8LTTRLtirLVHN4YMLlr09N9Cj
NgErX71dZnya2OPlCaq1JOpbxSKgxd2uyM8mFmM/xEwXPLF2AWvxPnU40Yi0kZYO/4SqPuJiFH2s
6kgYClsE6o0cEHpJXvfiOXTVNl6GyyVIZ+3rVPhhrkwKK5qBhz/25TJpjF9eHkYwO0GdYJCecBrc
UV6OgBXSkx0MSPgKYtRQKM9jiS9eeb2Bb5frCh93TptbVZV59Ak+P2wXKu3mK6XfjGRQ0EqcB/JM
PdgpZOLayyuH/5Qs1QnuKBun59In+hpYcnDv3VuRdzcumIBGXyros6lSY2mcWTGi33omXL2EX4Sy
lZ7BPHcD6+4I3P9FdVBoYIiRFyx+DesOgNE8EEc6z4FSzaLKhoeLAJLgvxL8JHR6fsMHuRU1nWob
xVg3CsaP3aECSk70uWF/XQXctPRQTk74r32AirP4mEfcpx2Pzdy/hqLwDhL4iq4mH7XCdqT5ugZ+
T3hBYCGSrxvAjS49zGOp6b8RLSszIBG9N+oPLNL/Ny5FmVT5ocfML3s2VdzOFT26H/umP7WRyo7V
WdJvGT34yeHfEgdjSxsrhzj4GWR3SySYgFB1kLzM5muJ+voSr8MNAFvlyqEq8JgsAAHkUU/kswUU
tHtkNrMoKzIuvlHQAdqUxOPlzUfS4/MSX9bxO0XtAUhRA/wi639BeiuJ4L7JPldTvNf/3yyXRtnA
qiX0LxC4zlLHv+wz0qdJdDdYjnLrZq3JHir3siROtWcGF4wr69IF+ybpmCRreJaJUQt6qkc3UD9V
62qY8oRsyVnFjygNW0Hkq0hzT4oosNY+O9EmsMlxLeUYB3U/4oYtoRC2456c81stJ1HRn+b7ys2F
3HsvPd5vfv2/mKQ6FD1LQVHWCxmWb72HHCbtxwKLghzBLHn5dMQ6Tx2UVtDVuSyXGVTUmdjhasFq
bbO5k9hxF9WXgNYd7ELhNdXlLz1suMFju8ZoAQJd/z4Qr2ijh9o0xeFtui8vs9+nueh2IhP0b/2o
nB8uBVn8XIJ0pnZekDTReWz9UM1Ms44RXX+cKruZXNHC0DkK3NL9Qxl5Km/Y2ERQ747Oj6S5yJrk
IPIBxtrM66teKxxsQ0dqBlMVxjhhKYMeYL9ySQBNCcwByEDnsiizVzZb64KLXK5YyjsHvx0dMpLN
mmuHCiOsiB0v0Jj56xncZjqr5kAsLvwCoOFZy9G2Dv1fy2z59zWo7n1OpzkFTsX99KBXAWjO759k
2H6XFBql+UnXn2HEffbbEJR7VE6EDqw7qEcvwyefejRlmbWg2cBGExefI5NL5884wQXnXNevTTdZ
NfjH59d/m9775IuGC4B6zFaJ0WiFuvJCjo0KBqX10q9ZqshjTqLZOG8KJTYhZpTdf3uYNdHg81Yg
mSbOADnNNPkI0J9MAeaf5z3yhQhRQNW6h2BoWAXVyu0XgliVlC6c0vt8nhMcyCBKBclTgmzIZwqg
ECpuIRdyeoJhClksMiRq31WgGvnt/HjVqy5w5kL+lej8IPSxfFsX1hl+zs8NzhKL9gH/RttA2ISF
U1yJzz3mrr4+kYTpMqTF4k7wNfY81lflH3TCosf8gwczUUkiM+5NtlYrvua3/hgg3BpAh3y4efF5
Ph+UnQlCGbS7MjuXDJcvFFI+cXM4zUOaUv4PS21WTJTseEJgbIuEGrw+H1DKl2qp9XbLqkrMMh2m
XNdIvcXTgolUhQNEIC9ghAZFprqQvaP1BwvlCfpyLsvesOExSta3tywlywlma4Acvi0mvffk57+r
ANKkapjUsIV1LD/PmyJpZljhvv45p8c8zFDmPV6JcBuDqWjoOzesVB1VRqHVLrDcuJLMhmRaGyQd
+kHwclsYqkvbEK50hZX1mt4zBscDnJa1dOOBHRpyRmBNtaD/P/5UkKg+zjx/BwSJh2gBZS4fOMed
7r1u3zD9MySZl7+ZEGc1mJ0yTNmYTwtvpinF6otsJYo1aDv24TUyG5+mgfjj7cp6Fweua+n/+Amp
UaC5LPM1+kVLtA4ehYW7FE2OnUl4irlbgSm21aiPZEa8WsUqjwB1QgbpNeRlJJmBlz5uWWWRjZrS
O7Gs9L1hLhOVia62bNOMT7le1OGBYvlIzX8euIz7J1uo7HSDN5Uji48Gsf2jOvulseLiWAPXvUPH
qVK6psm8cI6Kns49x4qCX1GpVTfKG0vIRqobYDO0uztJr42LCrHPGFrjRwz2WhSXCn0aRo09s2Ab
CELyZVGe3YiB+vR4ygZcj241BxcIdFpGSnrYgAMybLF06lOv8CtfYpO3+oB8WhlYK5Y/qkapHCSV
acYf5wIHaQycPKVFkfguMNQKeaH8ywx0OqwiZH9Kt7k0Qmdnhg889xlkvujUiJh/XdeqU6JcU/tM
gM1G+Wybw1jb67RjK2LP2mQ2cPjnnDlZoAegDNg6HVCtGa8wsMHiRMFc6mkIiB4AjgbygUH59O12
1cVbmnVoIhb+E/uD7BnVkP/uF4K0DdlQ7WpychjTijL+7bGON7t9/PuAm1Yw/cmTqSn06zS4ndRu
IRWVGBAacj5nOIWpscZMCQqeXSwiRQPrPcYC+faz/NiAEuHJciBkH08miryzhRCIZhbkz3E6rf7E
M67gp6ijqmvzgtUSjTYP4dRAj5F9kjC4+qJYb02gEeN3hQvLf4qCY61m3yyhM5tg42ATRg8eDKTu
X+pPoL7/8zR+4tbCEVJ0U4zJIqIY4gWcSOIE818xOfQSrBhAhaxDtYnKmru9c7N8FFRg2fiGQLJU
UyhjYwHNKPFRNLIO4wAy6+zeI46yOCvUSgKVgLJVeNDyJCOXtH6gK5RiOdo/3Jv2Qx2/uzEWBQ2/
BSR1JtxbPUu5WyaKdgBM5CWX8C3eS3D1HFiuLgzfmQEepcqv5p/4TZhA0H9gaxh3j+zpXQnhRqLq
4tIQJ6Tg0VA5opt/8G7XAngde51dX5my+Dw08qMcUrIY8yrD3vI1UX0CXy6XUJo32tFGLw+8cy4R
J79zShk6APoefiyYpVq97hqttAGzKLLIONHNRDTnfL7JYy75B3aWSoVmRRQ8iHvCAq4vOph1IG3f
I1W1myL8B03h9cDT9sUMmdgF47qIozyMUI8T8reR+YZGanZD5PdSl+OiK2le7LRWZVgweNNzMoI6
h7sxvS4F8uIKPOzb+IaaITPU85sgg7D929RDCv6+izqFZbeqSnbaiHGmybdWR8IQPbiqQxkSkdkG
BL2ZHz2/z0P9AYui/C0aCUsxr+p/tMc1QYkUkpbsWgmCi2uKx4Luz6IRxsuHJWr4G3hQG9vwz0/8
1NoQnJnEQlkDkuy4G0g8gLi+ClIfAVcxus1NfRe4CfccfP7NOzUn2H6yIrlG+sKxVHwR4AiTRUhR
U4mOdeJ7umu3onz7FZuWWxRF5mgFOj3UIgOYoCVUPx5hZtpzfxSaNTs7+YDK+EqaCmxykO6ioz5C
BcMkPIZnvVsh+20IFTnKDn/RZpacCuizHodbsShK6tkRyd2SZwtw4k0gLXajgrWMkiYmy3WAUxCH
JZsQMggDQ0keit5Y6he6bojjbpkcPR9h+e5by6RYejKDQPRJbER7XwMoJ40mCNuJrzw01z4zWinK
jq91pT3RewPMLb9WgFSnd7U9rBLuFJOltM/FQW9lTaD4osrovKwXfafJ2hnTh3o9LwD7s3Dec4XV
t52n4VTJOBGSl82sCc1Jun+LYftAflawPSoYeFUpdzdiNXM7VPJSZn3UA9UMBYFUiZO3LZHqJpsh
uJH1+Stup5MaUmlnbu+AcpxOEXCnhUYE7LtuhQTI0LDEnXZ9CqpLxI7uokxvwi3+7k+5UVk1KDlO
CL9CTUnUgyszOhcx/J8YO1s4TBvrHFlPJHt1NTJtahZxhotIL/QaROWY7EGfQEeN1KcZEUQaNi+f
W7bVXlMuE9kA1yyayfK+CiSl+kydJrvx1Vhh/q3aY/ODoad0BB1asMoy4ZDJKm1Xw2g2dgUkkQt1
/rOxHO/sTI/Tx5iUckJZ4CxrSWEcYVAx03HPfK6Vj34N9IM3f781VA5CPca3aq5RPj2pGJn5/WnY
nGnvD8yadG9arw8DaI/JHZIs5wn0MF1A/7zEoCSqwD3mbOH4eWTDkssZiriCZi89pefbEfe3nNoV
EhwpXPKgh2R0L7wlKA/1i65cADsZnbBb1jzqeaFyEIm4DR5fuUw+UquEmPcMmh9UT0gxuPGYI4u+
gbYGcFsrGOD6fRBGqzsWGywDSojmNzB4s0Jk26dyWV1huXPIIZhediypS0L+cUSZgtlMKPYQ9ikM
ypJj3QsRSzCV38YiNtIk8k4l+tcpN8bSPv0XM411jqBEJptTubwQyhNSwnG1/rNthTRaJjk/hOIK
xyfWdakhr5gs2bYWpCOy4s4unC2dWh8rmYjT5g5DwCivwwNs1LqMH3nZHLN90xsQc2Nb/wdIWJWI
wcxvJDlP02cyjKgJhf6qhz6YLLewLMCioS1820iCGM6YhGmCzyMTmsz0iTo8jxYcxehCSD21vGs1
mr34nyNH0wQHB6nLKJR0hxWlZOvz/Io756niDjWBZNCeWfpUfmj7xmL9z3tnUQnV5rLgxcdtSlU8
XZXqPKiUoy86JUiOhP9h3vVopRJPtNTJcby4fP3MuvMc39yUQTcbEYFrR77WKLUS0zlvwhaJQVjk
OunOi48c6O5A2N2J4SJJAbpEVenfwgzStv3EIMzWE5HiawWl1abFzlArZL1txfN7QjGGjYcT87U9
x88bw6LHoUGFhaEE9yTsmo0xFDcX1Lwc7X69LAmkjvMMoa998oT6LAVHQymR0Mx44EipzhAisIk+
j8K/lRIwvGAYoLZN8LrI1A7PgOF+WvTJnuBm0LhWCM2qx+cInygeBYqa5F+EQFaRjYjHZ/311Fqu
T2DU1H6GRqTejqxgIuO8Ywbfe63m5feFuGX2kXQinNKAggT7GuK6ZWBZNs8shdVsOR6ZrgW/JtjJ
gua1cW1imSJPwdzenSrX8SqAd6Zu3/e/Ao8yDEeu4SRVB6ns27cYp/sKWdZXbV0cmLmE+NkkmqKd
VZgyk7rHEQWzLY1Yemg/A+NEdP8KMk3BS1fek5AmgmJHzEY3zBbFldDZlgZY1GcEylkn6WXhBSG+
4rIrJUZTxr90C/xuDSGVQSr4++O69BaAuxHPADsO5k1mxwFffhFjX9iB9hY0+L8gJSNYo0Dkj8w9
iJ+snlRzW+RVrMOowPwaaOdREtpiyNj9aSdv22qGGXlNxKshtA0BL7WabdIW5tPnjQk0uYv9jNS4
KQ058X3avTqEEB780p2d2FbRhwAtrzWGheAoygxhwl9YOM5feDFyCaNCtpKbniCBmVK1YTFyvWaH
zeGq5zlIzUqPTPN1iXG43H3YvVgRBTkuyq5ZQI1EzYwlNnW8GOvOCcpeKOILF6ebEyYy+iVi2Mc/
pVQfiLyQlJl0pw3w/wlR3OZtkaWSQfsed9tbuHWTetqmMxbj6L/sPPoKqUiUJb1BQ8se08lsGMnX
MzkXz5ld14PgTpfTzOs9/4TUwPH1WHbndlAq50JZ3/myglNNCDzUoLQAXTe+m42+0/Xfd8j7jT2Q
wqJU2lvf/ZNSXee61sEOzajnJEhRuc7W/YHRlJsqWM1biBmP49rKx8LarI5HClvPrKGGof5TwAiL
daj2kZJptF9mS+6hlbz8lDydBjMDFfzMagl0lnajXrgWoKajEHFqau4UuL90MXiHJHshcdwbZKZT
GAMZurBHXokeMgONGSMlBMQz+F7zQBGkEh8bSWqdSCSjL5t++2bx4Xs3fqTF1ESXTzjjKdaIcY78
oNw3mXi/5S/S5eM1x0WGF06wzzf4hr6Q0Fg3qPU/hlKq195Pj91T0y9yyDBQv08Lu4d5D8YU/Bm0
+/CjGWalFMumz9b7pw7Z8+NvXMWJHsvzFsjk9VvGzfu7nwM2LXzDvHhmK2FNk9IYFxp4B6vrLgaz
q3YS51OEHteY8lJxwEgulkCfKuT503xVz2kUzC3n6dFcZWEKNPmlNukLSCiF7UsakzjcOtfo3T1L
b7p4xJGak3lyAHBgViUbmVi2ZaZ6Mpwce2UDsYyNeeMzcpmETBub9W0VI4ZTU0Hk+EBpmSC06NVp
4h1hoRg87gzB7HEI3BIoLMFD/ZM8bUYkiC8o59GMUbSwV/x8uG6thk9xOZjkmor4BE/fMLWcATC6
A3njJcDVL8nU9enbkkUyoWkPjlvKdLNfT+ixCj5g5C8akOZaaYlBfo+slEJqISj0mGDh1ONqrLEA
OdqbUsW2JbqiqSseYSxSga8yDjMfga7M/5gloCg3JmMmlQwRPCT6i9aDDj6/f37g+E0lDo0a8M1s
di6uKYBVNd8meIK6SMU6ECqdaXYHdDxiYORdt7nfJsD+UzMp8eR2ieasu3PyXLd21H2FV0A6KgRJ
OId0gHe57Bezw9Cjtpgv+YX60fpF364hXPy/gqA3BxJ5uC7XClBXutpsdlAcOQZc+e4IDSfX1XTr
o5pinV+68NPA9gm3NX06X+dHDvLKKjRt27HGG6RLOFmYeR/T63REVDaAkMe/zlq/Davw4N1KIC7i
iuSLaMyTqlwvlTtYwFoNdIVkAXQemOpTEGqC/ZPJ2GJSKbnHDqjlGzuNjBcpEquj5okuZgPmTH4s
Xrd+S465FgZYldRHADqG/6HEW096ew+2IKZMN+X+wZ9ubdsqC9TVLH4962HC8VexP+0x1I7fbw/+
G70FZWKrWWvFZ6XAF6U33CNr3xrAK+5UYscf/E00erRjCrlFYKDSx4uvYi5oNw5a+YJ8268uigG4
hZJmjUQP7cV+VrTRUlG73h014F2SIZBDrHq+7JDR/wTyS8wTBU1qOZfahE5ypfPMcwr+X0q4ckud
RpyHoqLW/XX5faFFROTsXO0axr1y7q1bDufC2jie8mfl73+4sPVVHEdHlinlQv6qjcqzYQcs3/2b
eUMPDwMqUK+9RIlc9D16SqKwZyF/m6acHOm0bDvc7/p1o15ANmUYZFTpdHIhEqnyi5qFq+6/jOLt
BGsDfM2E7h+nV6xbHoRcraJ2slTcu/hXn57UKi6ky1xrbM4J4Pzi+BywmBW0OL4JuyvZGMk0qgZI
0Ky8uOFTcJxYgNO6Afb14JxmPYAazHJhSR1huTcN4jFCbZSlGm6gSpPup6LpDKAhG5Ey8pAg3rYp
AayKEsaXHsutHwycwQSUZtWBvIKsKVW/qMWpp3Z+syQumk4WUQGRt9H5hfOh3E0c640oF1AO/o5B
eiuVYZeWU3Ng3JY661o5komMlzTOeyDvxXOYRyifMPnIzxF4CmgiWPh7+DCqZ+qX6r3T85mhuqZi
rV4/BPjSj5lZyJQVIxPx3y94r8fWV4WbEH7NFqmgj9hhFzg3Lknm93HOQgveBNnCOAkbHkj5msEx
1oI30iVzOoAx+yv8JQN2JKV54CK8qDbQuYqE3D+Eb8XjYlAZH9dMMNyCp8Yg+O/mKPirbM2AePo+
jKoaQ1cPoyNjzjKt5O04Z7LRXl1+9gPV+b02T97IUJ2F0JUXYS/ql0I/55W0VEWxReOdANqWLtTw
1Y+thoi6P5vnKvw5Tdn0oPVevd4QLHV/YJs63yI29/vcP1BwmThj668g1e4sH7+sfyqDYsMEOV94
q0wuCnk2PFZQ4kxzjeQQqyDvpe323GIboY2QWBpWXDwoHN03jexyhF/AIfrImAcNHWeSfuTf3CIz
mh6Rl/XUdNHquSGClgPM7vrsukLeGKPNhvZrd+98nWZ4XLFRjPLuNxrHaRZFsfMU1HBZFz0/JJu7
kqgSKZ+T0WX38tuWIUDsCaCGd7iuVu3nVUxKY7YimtYemwIkMYEMcTGk/W47EJlbxrtsWlpW1ka/
Gtsvbtpnq0KK49iuA++YrFy7QytrDcTv/Vmla4us16GGvptRX550nDeeBx8rF7Zoo8LWiTpepUfB
HCZnx4bq6nVc7xJIlDCzfcwPypZ3U21ug272RO/48MzmMloG2wM0p96fex0/s8wknpiNQQ/4m6lX
UONWedMwFlIlklvPCz4opLwiZdzRInsrvfw1F1FWXqsfj10aJU6dw3fFrpQvLWfqMcJ4abQs8GzL
/u1KyLAa9X9/03MeDYBHt8/NtT5brBVOqld1p0Ys9Q0c0s/KfVmlm0X+MVVT2qsBpV94t1DhvLfn
pI4muquiM4DmvyEGexwiEnJIEZc3pXRHfQlpS65wq+HVSeV3pOmgRL7aq3/ZZYUM2Qub/XQSvz5b
W0EmQvvj2cs58OVLQLgZxSmzjl5U8CTt8AH5EEk4mj5uNgPP5mC95n3mkAktwEOFUcSYYLknZUG/
E0ZgzNIFWJraORNCuXkCMro+ELKRyn5EZ5UvQlI++1/MlAqbmw9fXVNg9sgZwtyBc+zQ9UKOxjxI
Ky8tbtMoxtps4I7X+PBlt5K0NfoaJne9E96lyqT3OrBDC3ZR23A4X5DRDQPv9lKixIwTjUbUpSKT
L8AylpTgZd/0tUY0L5WhD52HsMnU/KwGuKKIOiSUsiPyVQXySXLcezg0+E+DaXg/6eAWUK+gmBwk
X5tFANeHAq8c+eFAsATkIxa6qhNYflJoW2arplHVutyPRkJbrcCEr2LN9WZzWX3ZwGhXKQIO/zk+
ae8vtZkUdlQeNGh8+gh2Br/ausMu+vYbYCNqC/BmL3uYNnOnr9VxsLRBQS+ZmDROMZDx865XBGy2
olmBsZOPP7XRv1FR/VjKpKfCCUHdoiG87IlkT11dU9LlssAAZsAPhw41Sbkkyc+5HhHleRTZgZnP
XESrL9QiDxQmQR8WKoehVEjWINnSMUV5OIIh95sXXD3WQFKi9t2Ahbb0vTKyw39K/slvdufQwTnX
La46c64o7paatimSZqMrFLePg10iQ9msQ92L7Z8wxSe+KzbTMai51ar4xlv5L99+jjvT3flNLijS
TDHVPLTRY1fWXpHUaBTLe7d5RumIJKNRjyKYC1px+UdRusmqGq4wkn9d5uiNlS6dWr6Vk7OEUmjc
ozJ0kCbFwFe2eiEsQKZBlIXOmTUyEnS9oSLZAw0y+tYsftp/8X1zACCfskilZY6YznbdrvD9vxIS
DdpKZvGbEqE0t/N/Fx/A+UtjYcOWGPJXqOUzJ9O+n6obd0z0SrLJDsjjKS5zJ4Bh9oeK44u7++2B
iLrPUerOKzKI9pVwPNaTOy8Yco7vklbbAReNKSMBEIEmPj/WBI1+66Ouf8dMXs3ALEtGPl0vQFN6
HZUuRmKL3L90Ty+bilyyQWzkoivELA3okSytvrbKhJUb13ri5S9Uj6CAeDrt8VSmoC8TcjbMa5q7
40ZcDufv5NJ9KguNnv+x+k639odjBfnHtWyMLFCgDa0ZDY/hdK1YiINR+kJJ0gAhV7vCAIzlp3mS
dWlSNenk63hqund7fd58SOlS9dHZci5B8ccLMkUUaOrNkD71TsmRgLKocK5hQdReZWInbJQHrIFo
9kpktNSvVOSz79FkVLh+LPUTxC6OqMmtvwwerhkxvvDD9VUvAMELw3WNvvFZAfuK33v8pPdlT2Gt
rpSpBl+cTpaLOTN7LMDMhX6iskBKR4CAZ65/OxHjHY1dtcwA7omgyDryvaw5+NpWZBUtSeFEiGzi
niKDyex7cepdFUDe+0w3UjCuitKxuHYqgd1R3+77VSwjZbHghovSpx67c0PZ9pTnn7Rytv7Ie9su
NYHaKf6NJ+9GoE1oG52mKTUEf4c8F3u6c3VWasOsyhOjPAs03/WqJEay1bhmhjARGyWHjXc4HVY9
d+1a46coRYZ6le7KTOH4fF5iLi26Du2zhjZixGSrQwONIK/sKKda8BGUO6Pcr4zDPa2WGsWWPYZO
hMF98PbC9304CAquQQqKEZD9edizbaLAxBeYsMFjsKd1HrwADJopGUj+tplmLB7nrlf5KjJ9MvKG
dcbrom0oNHNe7f/7vZBFOegj7iRTOHRFl6FcUmkelbzZjMdR8wjRNBgGyfXbhTvvKQZTGVq43pr1
gIokGa6mEtiaUzRcozclbS3/qtixmoZk9Vuc48JhIs+XlZGoN4VvqgRzg+P7LRtwSWXQFHGKyKGg
E0pUVSNvCVprne38ic3MeIzAM0JTCg07mt8wrAJ6UiXc4b3IferLxYe1J/lLWE5qZ01FLtdAgDqN
CMugy+v4HdOjzBq0i4XQBkcOCdV9KuegMviYqWB51ukhU78I7l0hMlHrWek5AA8ZkBNxHI7pHwbm
N1JBEj2mCqaqjD6flI6CUduQti535Fyc8M3DQulC/nAIbux5jATlQnwPnTco4f8oaxDnfK4nnJ9L
GfQLmtve5yRIC0cp5deyHnPe5I00QyJhSy4rRZHiCip8dxDhGkIJhk4MTnYtW1z3qjdXdgvUF35c
0Pg7Bb4SnNYWDtamRswLHXNrqVHqFwC/KcvXj/hVL/h8CAmTPGaETWK8ebyAApDMPkaiJTJzFU+D
0SUf/jb8Vl5oDFsCsmf6vEG0x49BzT8WVQofJ1aGxUiqr5L1VewLd+2UTUnonZXJTK1+YkzfTCPu
lCBd03e1mRX2pGI8p9hSHGypaNE5NbLuNvd/rZKkAsXPx0ZEJSEm49+do92HgQz1Ezy2zt4U6/3Z
m2Sl65sz8qd5WhAEn/kfZjHCuaeDo0s+minA4HUkCvgil8Gz70wnikNpcCl8MtGNc2i7NkjQ98G1
jwHhBfAx8JoXcAA2z+IFq0iMXDe3eEO5kacp2Odmu7DkXkhHNXPdwBwTyNmdg2D+u09YscQmp8ZK
sJqGgIYTFlopRzn3U3HgdO4u8uv3NtNrjSW3bRKhOqMsSo0XKaOHPSzpp+SqD2I5aMlZsMckyiv5
XjHFH4K15lcigC0M7FXnaslLGBn2tlWiOW8q3kBOcK5dwJQF56raWIxe+biNyoNWRBet+uTEzLmr
VVG8C7ObPqBOIBaWfLxKprOXJZIP7CTw+Kf8p3Zp8P3I7mb4oiaWrfT8RsNSfTeIWLYq4Yfyr9tx
DHuwuaVd48dAnsk2mnYLZnaJ1gS4gxw/97mWpkcZje2OIYrnzrwXx1SGK7tFn49wXkWgy11OUoLm
MnAYgK7wGhVNpSHXX9Bu9yAEbVyzfJUBPt5ga8kTtC9eo2HtfCeD4y7XmkvCAkLWlvOWAr5aLKXX
s2VxP9RUlZZlPjjTfi5Lf6ZHpyEVZTkzgwfWksDjsrTL6lMIZxA4GpRtokXojSwV2aAAkJhFycOo
JPF2vUAPjNsXZSjt+PFsXr+BF3YCx0Rc5D0zsOmHZPB+JD4DucezdzWcu8fBa/C02ad1IX+k2a1C
+XticKgkM1USSrTL8LcSO7//PyFVJytUO6jWg4pMwrUCdlyC2ox+ic3ddLxVgzU00/yaBmTFiqy7
i7nWyLIma4/Zzi/tMnJqCdK9DH0lbRg/VaO//LaXXdz1nhh06FLIK6T1PMKRPfu7cCXa76H6PFAy
dx6tfIMuT6s0r7rCdTODBZgYBIe9KHtmcRQE2J0sK6kFdE0xaakN6Hxj7xzjhBijVyNilvzrgNOr
YIqMimNgn7ntKUf1BQBDFdWfd6n45+0GPqGfmtXyRUt7MPDfuFSbqzlseeRln0kei4sNNaUFmpPQ
fq5QBrfh0lp7AJH/XPfDdmUoG+3uKp+Zpv7pvTBNk3wRBJmCMRcopuKDgIyOtV9Y0DoN/stNovIR
S7PyIl3iDEHZEM+B2CHZX//BY6mCP6TQd/v8DO4wyT3XDtD+ztBhXapiSrZsmX+A2R74zVLIsuP4
GH0mTDMpXhZhfYfuFcXIRB6k9Ur2APedzwBudkegtydLnt7AqOTRvIn7oGftwEVdzWkIQdYMM68N
bnUgBlLKVnBB7ItsDFhuii4qGdGXhLM+5IJdQDbG3tv9+gPigkDlnqXcS2ywMotWTZhhnqIqDybn
CbajBxCfikbRqCPYKvJWnn5ZghviQR49Y/7q1SAuM417T1Suun1fUFUfOZ3OQ9Svg5PSlgaupxc9
k0DxGccwelRDV/h6kb9NTtR6qbvXE8mkMSt9Bl+aVjYa7L9vlylTec90ZQ4zkqTLK3sGP+NRsVWG
gAexgbpfx3eKeSs7XsdC5ecmQ2jXTf2vRgwXs7Aw6t4UK6owIfIeNhKjp5LkUwEqnZ/F51OwslpY
F2CHE0WHtxUb+wXdA2LJWAGhjWWjrOfzMKAZBjeDQy4HA6wRq1ZbizXcecKAtVoS8v6b1Ce+e7Bs
yLG4qHL2yxbg2Qskka0cxTiRi/f5ua4VrLP6BprMVHE1ipk0zpIdve32op7ijBDo8seSI7I4pSNq
EwU7oPNCD9n540oJmKQelVxCfCQz72+hT2rEobAIBdgfXC2pXcai8N6gz4HU+R1cOT7U+zS7T6gp
DU1XayWPUx8QFtSPwcprHuZwZqPbuwZ2xOI9Hg+BTOR5Xes5k5rOnqZ/LPu0ke7+fg0GC97No7Hz
rSkyRjyDCnzJGwQuf8Xmheo344PUKjuGifgSXg7iKDLDjn7Pj5+rjJaOyGwHmzi2UbcxbZUjolXb
gFaeXAqM7g1FGoDa0h0UTvKKt+KtvvXWSiMWJYWJu82usDVurN6EcjVWpcC5v8e6Xt7vQNGc3Iek
dGFOc+MWAXTPlAmUTS9JC5vZl5DI4BXx6bswF9gy2cAp0zwX6JO8VPiYzSrTSh541UgoRddb6Cql
t/OI2Frm86ElH56WjMgHoM6vcpuNfUnd+87iUy2G20q9E5+z8/T2rgkSr8hZlm/ZYLtWFlUfOMHx
oAca0iZdqjyzLMLuStxsyIItklsjc18JwGeDtJfVTGvJRi/Q9+rG9PNg7OQ0HsBcGpwqNNyWGRBa
NNvXNr+qbV0kr9e8Ucz6e/YCWL8FD8/8nYv8QP0NFdB9O4+HyOFI92tPc0aho/4ZP4i/X6cF5UVU
CITku060u4H2+h3LKvqf2CkQ1Br51TLssAD9HVFYyIjc95OD87Rfb0hPgSiJovAqmaI3eDg8QCah
8uMlTgoj4j+JYPGYpjhy2bjQI4eEiVZf+njXQQNMClWc/uMlLY5PKQ/mdY88I4imi2k+F3NswfSg
It+rStQhHzmfOKODYgkYWhhFSgDcjCECenVhklfjs+e1YXNbcvIpRTZOVkInPKe0wiwmNf7Wp1Ij
/kjux3vQJYYw4l4B5PNCR3yBgdcrvzoGuNAtFY7MC+Urp6MAzDW2ivAvSV7aPrGpB1noba7ZsUxw
Ezq6C7bGCO/xsKCNZ2XZEEWbiM4NwJdJ4iKXJ/C2PwE2cCbn1sPnzUtkCtmgHZwCKirAlsY81pq7
9F9b1ZHyHrBnxxPCO9XHmqJ741EjIoAV9U84e393pchaa2M47uJreTmf7WjHvOXVXYMC63scAJeg
2d97P/IKULXMD4clgqe+Lq2QsMwq4RXZnduMfXbVXIt298KJxG0fG7RRkiAtjhk+I1iNBayAPwEV
mKTVOLujwX9I/AgTsGjTHsYcI98WHkMbG5s5UCT6YILlRm6BCzvcWsr1SuyDBHuf5s6fwzuRi8L+
uEt9SNWLTaUcIHVCJ5x4wwLbQp1XSxY/CAYkBtAjg9VKo7Kknx98JoPWOZGm6Dyc5d+lDHSn7Gya
OwbpJMd7wV2LlCyReRgjRiLWyU6QeTTXWEltQzgqCzvgr2UH9I6Q/w05Dsv5H3lodXiYSmgDR+UQ
uySGKO8QXkuSir47zXMcVU5NLYB1OuyWUNB9RdnSnLmoQxo/dDwEzZkUgq3Aa3DYMN/qGYvErO5X
fRgDw3IPFiI+P3I2j98ROamSem1rMrX7t4o8beWFM03C0hVudqGEY4xDzfJ4PEAekkjGHnWBATOa
A8EAAsPbDoGIB84MT6ivipv62N/rLVhopb3Nw8WW+iTw3KPh/mGSaB7DiYbbfge99hwOYM7PlPt2
lVCjaxHJsKXyVVeFQsPST99lChBHe6xwQjr5ZJfJC2wTfvxgjpNjjb/fNxlMgJAtBnsP//UkOd6Z
fhj18pab1MRRkI5YnelQDJqj8nGtNv3YvwC4ewZaWF+VMAKaZgjOTP6A05rofY3iq33PpzEC8eV5
eWyXoROYeXY8r2bsXtMerAIoVVROUnhvRzkwSr1+JRvw9/bLfRlnIOE/GMmtrGLCQ66cDh3aJeZe
SXiVTsuG8Oq4tGNhMlRG6JBeuLMGiGshgKjXlgiOdomEs0WTGEOz8iu+JlccvPWLguX39QTFIMkI
5X9YMsfv7eUzkXsXW/juUFJd2iOCfbTwKqkRi3X3yA1drV0looeuPgJk1BSAa1ea03OwfhAsoNH1
GLeEMxIO5jIRN2rmq/lwyT8wH9p7BaSs3+ZDlgxVnVv08P4mgfyCiU63SD0tMvIXcagD8EdmnBqC
SpjCoQnATr4WPCngJ/kEeLo31hwPeXE/GlaOXSrR5iSVYC0J7mpjk4fXSnbPxCQMpaCdY9oMswIb
ZNhzqng3mcN/hpmlyf9P8Ay3vXaUhe9CwW9UlRud3Z1cN1EAxKlTDzGD2uEVsXzThrT9HaWCX00q
eAErICIY26KLfu5P/2GGTfb8TjCYwYvhqV/d6KbEEdIsmcbUdi7eedRCzv0RZcAPthfOjQ+YD/ri
0vTv8tNqOlJFchJzV3XT+TSvGApKx3OMrZbN0iY59O8CHgmzWUMyYzTEJhBmjmJzuq0cRxWJG/Cf
vRN5Y15/4J1XEZLK80ZP3gdGb27+piwOrSspmUHk2ewRoalVIaEXfH7CwTd0SfUVJ6sLDTMfdp6F
b+xr3SM6T49+hyIMD/gB1T1WD0PKz1hL66l7ZD9+N9psX/soE6gomq/CK4SO0bz2A/lDsv5L+Vij
/ypWJIX9Mqz2ppBQUWBrcAczB2WFYuQb6TKZ9+H7CYfMCePQQf4GE8AxkCasXIINdfoJR7Ko+RFU
XkYYUztfp9aOwu8V4USHT+jbwvqn2a2c3NbXWsCAuO6XdoCLv1uroqx8MlgP8Hd3Yx12X7VLX5l5
AYg4zETsxtOQb3xqoNYhgfprPNsKNBUwhHOPZrz+zdwHgDe2SI/whMHellDp2KyOfmitfH0h8gvi
VNJSEf68WVmp0UUSpILn7Sy+QUzCI7ta5jpnizR7pRfo3YhbFWPAqjoIL08pTBtg6kUoiRRlgZlU
EOvQBinqG5Oio3hC4pxc4JsJor+oyu8V4Es/PDYj8qKszw6ojcVrBMfqc/4JZcMXf2lVs/kIQsYy
VyQdeZtKFeHiexFryz9FNJm6kFvH7G5DLYu6QsBzows8j/HuaitJyLwP+F9OO1beIWQ3uy5F+5ys
m1Bhie1nfsmCBGCgOOBjfspSvlHhKHowp5IDrNy+TSwVEddMW6pSjZNyEInfEDOarnJnVkP9Q8Yc
oFkJhtlW2MQZ4FZH//PAwvIoRWkyuIW/5trNvKouRbzqLdfkvk2Lsw2mhB/Xmv/oK1TLsC3kCBsS
hsIWZ9kbRaGLfRopqRmEhivYfLFd+pQA2JCewflcxDDZn1dXQruNXigGSiCSO7zJPcyqMiavPWSN
GyczHhUcOnlAXHza0QSJKWJJbMjQGiVRlaQfZ0TNToqRvI9v8bTP662AH7iztawuO94fX0dHeQiV
OB+b0DjsltgMv9ABxtU2G5O3zc3v0U6VRkbEHmaV+ycpYEinKxTqE+mtG5U0pTphg+kRRIK+Wk3Y
b6cDkYrysFAUorF31OsLMQxR4Ify/14JDYVH7ptyfqWardAfm1ZSgvmqtqNq7SnTqOLA7kK2hijE
zeUWMv0Y6jpF/uyno2id8/25WbZi0paZrOjZfpgCil2UHUBqkyYG1bMplgHBIjk1oroiCAfl+n+p
UsgEBWq9nnvM6iqswv4FBcFswU66+JE1O4/+mizCldCSzZtW+FzAFWkRQ/c+TGAJOU8zgGR2dEVv
rEW8B26tRbSnlJbQVIhyBtBWV4yz1skfap6N9E0suVHqboY9qpFiDCHpYWk4rllBqXNgHZ267fIu
6eF7VyMkfQzGouE3GZGaC0RUiKRLX8JVUwUb5cwdLd7KzUeSp+/d9C8j4p5vNiNuPY2KPf9rre7t
fQdvjUzTaUEorGJy6W0BLqc0cD1BCOMmy/GpTSm0yGf2UIIORwpFtzVEj2lJwOsu6UQ00vh6u6B1
72J8zG5PzyuruPOQgnhhG+1DMZi56MEhZSr+frYqUx5ZX3BllsoDma9A8u/U8EecmTCdpAUpncqS
EJynv7d58oXCqcdLG2p82O9gYCPzH+iSINe+RrNk99dCrubgIwJAJ5k5o1HMBGVbklm+7IOPDZSP
spX2m0kPV2uVf2juapd2WCFuQ/lpUa01+kfzoO9iQ2azi3GvvhE/oTVXxcQNJpv6UKimGYOeZTcS
oqlI+JXSZFi95aAkWvY/lE5nnhdQAo7/dEJPvn0spGFxV7vP5cHkKuVpHYxJJVPPvKB6R2cHBHRR
bEmEboh1pzXYtqrozjcaXJtworvywg8RtUw6j8E3KTpnKimiDU2UnZqJr57adHjhGsv4Xmsyp0m9
rtMgisgHxFRKiYGGaCujtJnOLwTHsCvzsUt11hQqbKqZLAkxn50RReQFgrAnq3oOhvL+IrPVzLJc
tu2J0TzKO5bbC8Ct2DTj5Oi/NF53HTspS3ULoSzrB4MGSR37faYT95TRmNsyzISULL8/PbG0pWDB
ohsvXIvT1N7jGDmNRJafs/Jm/geMzYPfVffEZ7sP6BDaQBzFB/XuVUz4Lp7AODKGlG4nLbLVVO3h
OtTyoHH+Ai0gRUUtjZWixqwaiGbNbls00HD789m568vy2iTyRKNqBL3ss3X49oCoEECIO7DXe5Yx
4PGAutghQaEPYxAQYV3uR1niqWPxbAa2RhtASNgJF22hT0zpmy0yMUKdEDUKZo6W9pX02ze/MdHW
sDk1N5cTlNIZOavlMnBFB8plhof11SkuT8GkNxgJg7QzKmMxC8VWXFbzobMM/VjHGXtLK4jFTqXe
S9pbRoD4eL7CEKCwZSEXAVOAtC03fR1pUQxHUNUUzFPVKmTfUKrKOuZtAF0e254mxCfM9KwipYG2
5OxgXfWprlLoPSRgH7FpGXuecrFSlqFXsqUiTOQuADJPY32bJ6jvP0d/SmDakP9t8kSwFi2zjhk3
FEI0wSzsG9RlOM5AZBNrdDp9wDQt3ZFJtz5Var1L4haNSOqDowYO9ApOwdk9a2/HqIigejnk9XSd
pp+7UzSuSK/cxFtZ+AHZVn7iqwEdC0VOriA5rFbxxVNvcqqvhC0aC6fpccCKsfDk2j7BGzjUt7Bf
qRzAVib/t9FtZdxQj38e7jBfIJ6G6ZLnqjz1cuirYv6upROzkt0822AF46fwZvrLaiqvzQcFKNhf
+zHcv4abceuOYolK8UEcxKJ0ETZ3bi+Cs9+o/yZbTIv+aoebgFlFktfgDMPA8iPdQGCl1eKRPWUB
33aakpbT7o/1d+S/6jUwCvxef3eaiEmkpG6TsIMQ+LeEqAGw1RpKSrPGkhenyWk+xVr5DqgxgiIF
n5ruL2ZQTG3HCkarnqFwF6nBJWle56b5r6duKAdrSNcTBT5UnSVBLMhtHijPmL7Tm45qJJNuSz34
Sgoyz7euezcCpxbZyO4AGHufTv6vDlJrzI4ueM5zVu3YL/vPGdtELEpBiCmt8o8IIGMo2YiULa9u
3lXnhjryweSLDC5WSeBSuk4ea5BgwO4SODeUQ/Fn/rujODOVlwBpCLCrbdliWDegZWJH7oKJWECZ
kFOMBPS6BiJMfgvZM6H3Za+PG1c/zq/HOQZZrQnwg9FBoGqyhdwkUQfzMM9QnZuYZ04K+8NW5yo0
q/GF+w0puH4QJ9Mc77bdcaqhrQcp+XWw39qs8ClqI/EhrqQ/jV8bjrOQCFV3E//sSwwF4jrGCd91
USkCGXDwe1SqZm8IPhxcEqSHOH0V7b3IzmrAauIUHE3fY3OM9jwSuWv35zDkO9B+BsawblnJzkyd
sE4mqnpPPEMRDcvXWoFIojmHWlt6IuiSn3O14PGafqnSERixSPcpG4jj+ke8m4VCudxrRvW/Mh7O
TZIwXaexe2ii+KwgxYHZrlrrnuYrvJEx7UM9kfnsjSH86IaUg0uWtrU3O5LXokW0Cw1s+dbh+mh/
eUW29z1SeRW1KQA2pkPk56x60JfFMbkjjsYQ8AdUyCAr4WCaoNajs0ixdPwTTf9L1cO1qds8eFVt
h+wWJYg1vUGbkpTYzbRzhpDrnagY9ubT1qZFFvPfw6FHtVcdveaXB0Udj4ybKn6Gj2oOQ84QDdo+
YUCycpa6EV0+usdkN8je4LgDXiIFCelpDksnhsVT1+Wqwu8LAxEuFrszNXg/qVgg11vbU31bnTQp
OsF6ae0V0onmy35RtHbDQ0EANnHx3aa8Tv/5jELU9fHabFW7GenRmRzE2W0QMWzW/aookJB8JBUG
OP2ohFoBpC10vCXuNBrcytgb1Fn7hKSJH5Ii/vsXyug8inu9UGSX+OqOR9+m2+lfpI/Cf7Vq9Z+S
N5Tci2F4VEMbvfzmrMV9zN97BwjSnf68pqDrArIumgiiOBluA+cXdpK7zI+SoBpHt6w6nu7P0dvC
IbMbDD6ri+F6j81jdmkkRmDqX8F5rVexwdWYetI1CUlb9hS9it5VAgWUIpt6j+L/2RgwriZsg+Gw
k815IBaxyvSwgiiWgQd2wguRIyuurdWzBjadk+35wf7+UUJQ24+jwOFCtseQdOnpOT+t3Y/Hf/VT
IKG6q1rFpxZGYZ4CIKcb5xJZvKu/5ExPwRued9P51sDnLIFTl2DKdfITimD0xeiT3JRzd4xUTIo4
VJNwlc7PmdfHdqgBZhK3C9Tm03zrz6jbDLS07A8tzY1VS/cIdLWiy/UINJQr8yHOcPrK1nrTRp7i
QSmcrgNPvM2c5swZMEHcFUZFOLOluXnpqR/6q7LpC7VyrBVXjSmVEPhw843Op5RtS/USxvgL541y
v+BE4LBhvpVSjAf+6o0uk2S8thOiEfGMFlw6mfiwhZW9ERD3++da57xVwnxg+V1n3hIDLq2F7YyU
AFLZpOBFnfCgWzC414hpgxLiW4abIgsX4+uqrFNXipt64geEveAL0bEmQSvy6oL65tLQLx2LYU6t
OYW+2H+QOjHAkA/rnqLOoNMlxwTM1Ae9rDcXjXZDi+V6QwnXuf6qEkHflZU2nwv2vb5yxty5NSwP
RtsxdWQf1SC/TbPuKOo0B64jxjPDR/k5n5h7fUh39QJFaUUCoyBEJ8aD7+tqj3NcLD0PRmWa7fM/
v/fd2WYLGgHxBpxD/CHa3LiTH4X39aHbi69lIMeaeT1RN9dpWI+sjCZYkg6d3pvYc7rKzoAVYB2p
Ey7C1sEy1CZmclqD9H2ntUOJ6X+uN3Z1Wl5Lz2hy/FnEY8FVdTPbozLCrm12WwbnGCNmseGmlZ9r
XX9bCFnv59rRpr1aTNIYKIMzqG7e4hIap6C7hUABBMsIViEzvG4zCoBVIyC3OqLWaaMblDvztEmE
nXm5ItC24otHi2k5jhR0gvSVYsDnjb1XETUMI32sFY7rR9j55jSzuM2os/4N9u0mhEVpcWi7XchC
8k1s4favqbq05FZkLam15/Hd993WQH/zDw0AwfdQD72RCUPPozMo3zNpJ/0ES4XK3B/0/Chj76sE
vTMFI4LW8ken5CW5/gRWlq1rTe6Tqe9TVPNoRtKEk6b1p7/lSA/kPBj5OkynceHErwrGctZc2BRw
+0Mpx2rb93GOvIfTq5fbskl3gNVS1QHWw21QT6DapJStvCy1xRgDOJACldElj0dsrykh+D7kX4NO
iA2GlftSEs1jQbdGUgRW/9YNjkQ75sf/OpfFUwFdWTY2FfjniQ2w/c01TnHrIHYfM/ZuIYN3/sgN
fX1LwQvLqYp0qOAJ7uWd/jeTm5MekkFvGviv54heincY8Xb1548Es35XBggNOLpEvN98fLz2rZjq
vSCHWfqN7asQzUiMK/QQFYxWNsXpPc+TIYFKVRusRZfgedL0jiXG6RpkzRAjE7EaAwMJYrpCWvC+
ssZ2XZiVPAKnM0q4StGKSPrmk/9qQV8GaL1/4qyfMmgInDs2ZJU8Wu1m9efF4tQ7qGr6MuPbvPbo
MHBsLmzJed8U8oUTUk5fFrEZz8PMh0/oGwAuq+qO0hgJI16hMSUklTYLiMg5LgYtngPI1r4/4aI6
F0SpsEXdufHseDXJAPWf1068E7GD5NAPf9cAIDl7EapzvzL4srKf9lmER7a2hdeCwszX87Npyhw7
YodczrFcPljjuSIWj1a+wo9lZAPpteeuyzzofe/4H1i0hNrwqCuMWYfcu7Xb/98u+hktsCW1ctuE
EnFseNa42B/as36bMWgIhU1nuQsezWrV9aUogfAsqZuUUxBl3zc1fB75cZt5RBz3Wp2gl/8F80Km
cZxWh2GYcBqskNKXqQ5IILmFEl46tiTkKjlksI2jwYOERQkvP+BPLocKcmYWiobwsZ7a1YCgiiSb
uV0J4EJnBd3ynVehZw1TfdSpCCiwommCkk8apC06oZgAkSGpNHFQ3/ziNW7aPFGUAoP4Bf3JetZh
+ZZYqf9KRNrU0x3iWGPkB3lDiOD+ZjeCP3DXV7hbD6cbsuncX/XR1O3MIPscRqS7TRXidHyXVG1B
SyKFu9NjhI4BuHbEmpgW5pJPPBXlupHB2hAS2+bP+vNmdPAHKA2vWRj1QKefYyfM76Ah8ddD8jA9
e67r1D1fgcmLS6itPA3zJ1VWTpMaCUEseAftinB5x4f7dG3b0GO2RN9k9O4c4EUwPmZef3IF2i/X
/Ro1Z0CDwzCpa0JL0uR+Od+xpFPcNYKhNAUH56fk+Gm3x2JjG20wkz6RW3Ol5R8LHfHCFDMSj9VK
sxWBOmmusA9ybvbWXLxY9HILN8np2Jm/4c7QajHyjfM+1nXtG7UUijaWc3ij7utyP6jVAOdfKEcv
AJYI67stQNOejDB6H+YgmbksQKN4q1720Bt7z1qUT+rGjRuk1sG5qejurvu2sFC2Ytrfac51N5kN
X4oJhpcR1kqAiKUhMkC0mFsTZlyf8TeFtJ4uJ7JNFq++YgZSRajGWO/KVVW7JwcPff6HDridN4px
2c6zWTbMlsqpqJ++emohn7t3hyV6jWznvS0WmCa0x5woL6SQ8sx0nnweU+sq2nyylNswAJCcJ8y3
JETgW19x0Q/srr062zOEduMUgeDRmWl75uyvVbR9Dj2WSwn9sspCJaCgjRioTeNSJU6/bu8nYvkA
7PZ+vman8At/HVUnGRFkGko5qLWwAaGApvIGm5x1WfB5qA0UC3LDbI6V86JvCjFmykiQPMAxh12b
nKBHIhcrJkpuA8UxuXLu1tl1GyqINluRR0VsamNxJd5Y3ZYfgBcuxhH0UTEJ/LF+tK1xYZQP9Uh2
SxVtA9sm49QA8hpLHolcNrNXEowpfeXh01ZvSBYDlZbQnasCw9eDAVJvtqVqxUgXOfscu5bOXrr/
IuO6rkv4yTM8UyShCVXeJZxL483G1Ik9HVjJ4Mrg8de+CdN/OfEPPqwB6VGQtdKaqU/XPAL02ahJ
Prf15ffkde0grnYOjt49MsLEgOfIp53sbkMLSR8CpRToZi6ABYZeusN6aGapp51f7SGR0SpQi+0g
t2wKZTQq+4D5fHoWkuB5xoNmNJTukWCw4BCvQcN2BDkci31WLlr9bjV/5yg4UU81aNuwqcvX06VH
H5P9+nimGN3tAkWCxFpOR/x50HSwoEvV9Qd1uGau3+oEYzNkpppmN2DkjOcX9hcMWFOQmN1Pp5SH
eMfo2OpQihyT4ZnVskj2H//7cb1X6og+h6CBmUx/yCkwA0WvQIcjUofIIG/j6BMuwmoZeu0HsDiw
zOS1crdrCdzQ3Wmmo0RwfHKKKxpMx9k8a9DPLll629MLRwm3Zg/NvVA2krqNjKqSz9xur/Fv9HnD
DW+Qbimj/0+jpEnlXVy55QtMfPYKWP6lKqMfgva9Cj13x9rEGw0xgZ6lLsFunlw7PsV5xb+ttodL
M5vxonvTE6aeymxmobyy0nk7Rs4f4X+NrT5lPnsTzyDGhhmU75jPdvz0VFt58J7+JpqY2YMKM2z2
TDYZThki7mom48J3+jQQ46WeJ5eZz6Yo0LAPS91gQ5h7DPxVGyc3nTD6pho4B27naITsyRY/SFdE
HdMtQ+2WOe4VOjeL301RAJfh8+/iXPSS8cqA25I6HqbVezshUnaMFWFSo8kJcirjR5KK4iKcHF0d
AS4ojfiIz84M86iWLZd/vXU9KWtt8Hg9GV+Yi22EdZinyBYFADIeTpQl0MgKrdBjLr/b/RYRM0iA
V7fwo5iwN3geG4AF2v05jZb6CX8F3v9vUhvvc0pXvqRZi4K3mBZqqvlPF1JSW+LakDBk19gdLEP+
RFQdZZ0p0FI7TJxVe3p8bKTZoS/Z9WnFsdKATV0C2CuZJVMS6TQh3KaIkHWuNmCe4S1RXOw38av7
0NpvjQWKjC8Alja+6zuX/7+45CwA8evburTnrIEQXrnob1BWEKhHyx2Uu0zSP3rIdECNLARpxmXf
lmHT385DNi1Jfvbj05FPqNQ8lnB77IRgoy3mo/YZYr/jdAgbZcntTVO5iOqXjhpCp3eXP0x+0HGo
grMtVdQPyNBxbvZFD64VRM3nlY7XkY+vI5/LspSngQW7grb+Cb2Ix8EQpzpQg89Scy0kBnSrAl9n
pgk1TVJ4JmE+0N/d7B8JiwbmZjTHJEbdHcVEf6Shj2bcWvtmWnPyT2prJOdHtMjov84GrtT4qlQF
YNELjKkAzYZo941TUuBb7PktYHaBQCgyHSRx7BxG+zxfh5j94nKQzR0Cq3t0FysjoMEdPOZKAigh
i/cIH3Yv4Jd8qWt2K3UbGsYBoUurg39k8SURR6kltRhvy1TOY0vC4MsYUGyqYW4W+bPri1A/dzG9
Ru22tI0Rtg66nZbEnbWxgFBKIGmAq7qT/79fp+skVm/k1QQO/43a6Ap2hzQtIj838Fu7j6qkXzEQ
96EkXuxeoabR+FbOWTEzo2IESmdH6T6i6NWc/3ECm1PfuXnmA9bUHsjFNUpFFNqcJpaODCIwjiBb
idz4S9JBm3oIBZpIr0YPkMqP0i4wBHkhgtvuONQ3my4oeIeCEcBKztVh7LSvUId2rNcgIoDfHn/+
FRiAJUkFa5GB0J4kmW7dfDYRbegRH75s7SJB1I9YImfz85elwqnx/gB6jySrNMxIJsZzjn4La/Ym
N0VYvZz//vfLO0K92My1ec6kivVtourldcb8/kxOqg0yc+zC00I61DLmSkhhq0vkIub2H7aiH/61
L+Y/Ey0lEQuvYJ5SO/FVp75+jLgXkq9V3gmZwVty8/7mNZvQ9e4e5/Gk+QIVb3Z4Fn+/l3kjVDdW
ZtUUDFLeq1fpfczCx1OeLAuJRsSIkU8V8PEpEdw4d1kLXFK1JLkRmuV0+pajfW+OMsAVcG6suAb2
pWv29beCGnfIdKRyVwXibQEoJxa/t8PJzx/oRciSsaFrNXeMKvdvpoVBey1GA8064JFFPkMDGqZm
R9Rgsf44IhDucCMNNKbgkWxGBhyFaSaTqpkiBOYCzsxzGvjnQ+uu2Wh2Uj1v/OhyTy5BmiKwtlv8
KInIsXlzUk0lpkhYJ7kc9Iu6RIFNFAmU5zbljTTN5Sp7JGb1wInqEe/lnGnsuf1IwsojyLU70wjC
ru7TVyvLN9N5FeIrbSPU1KX0T39DNjGkMpPP4WWJrFg59xj04Yhd8B/MT3gysCFOIh83SO5BuW3T
prTSGrPXqT8AhSSsFsYn3btEE10PfhHWzv85kwBg+CuYPFHwsQTRgoBPu7Y2t4VebU4yGRFiP3Zd
YjsHcIOeeUko2uAljvVcJubBbZBp2uIzB/lWBpNn/zxUWos5VIidIKwaI7lgCKA8D2HzmlYfQcXw
gHOV9SlBlGVLVu7UeAfSV+gCMf+NhyrP4U/NLCpqdim79fw7nfW7SoQWKUjEQ/5ZvIkjR/SCFJad
8eD3TtslwQgwA39sSI7q4jEWPV59c/HIOs5y1sEux1EG+j5PaGiJ78ZnQSK10p90IcMj9obvD73X
LOnvTativ9/CyfUjAg+eLR4yBkgDztBcutkB5Fup7r5bGOQnQjd16kzW+Ev7NI11JNmenSClMDjc
oGuraAUa6Oqye9oQIC+QXpwAxRWKFwnMVVEfBjSKkahXu+mt5uL7XxkbVnAXzrMVlhDQ6BLRynjg
CexJMnPChBZrYwojSjB+mrAzxMV91tGWr9N2IFRPVxAhRtPrG6znyHG4KbWeEsHV/Cqs7TbBJrJo
RSbTzl7crmK9agukL3eHvxe1/DoppxsiyuM77afOQso2NtQso3QcTbjYcYBW+ZRsWDt3x61G6oGt
vkZ6QITtV4pBE2jIHmpscZ0MeV06t21IKraWEDSqWjj7HubSwGakXnM8jvzJVJdQTXVk8NREAK0q
rLVDn6ha+91xe3ylORBMHqsgtOU2solSo6zlmPqD/6omVXdhlXsgRDqusgy8+h1NVnWtiEYOOgwL
ZvsUibBBq3IS1wJWYHxPGjBseMO3D0a7fMtru21BBZ5zhwv78d5gex9dryd3UrUTzh9e73gqSWe2
WFxMGRaRdS0jtYNzzYbDrN5UXA2VbdLlh/LAo1asyuXizRwZHXAYEwBKr5bpgY7PrD8p2OJK+tDL
gPjclpRkQN5nSF1O6twii7JrVXjXP5ggoAZvPV6jaZZ1y6AxzVVrhtu0kXAjKCy3dmmnZ31BUNHT
/9NHG7Vc8UQ8bZkcKLKbVxY2NWjtIwXjF98HU0Lx1SHwrNV7z+Nq5IrhQcnEZ+vjr5wQALNQnrhn
nFUXAYD1xp6iBBKw4Onno9JPIoF0X+fGAtDrpWhjyL2lw7CjCagvBF/xLf4AJKSiKdnHsuCF+qJP
wnT8qPSWizLJ1gDdplgvQUwUA2RTf43RMZXkupvF/xLH/FXaBYLZ4M8GSPh62C11VgplNwUWgN8s
ROZlMnajeuojBm35zhkRDvzrYtBUNU6XcidJ7L2wIG0+PVHvjf4WfaeSq5JhjotKYtSFqGP4jpQ8
DjfscTSc+RrJ9bCVvu6DnAYpBjtHVVEhicie1MB+9GzHM2XHXtZ8oLHCT6QEn3Q3XigpFBh0CcRa
7+CQFm6vpZGXWcDri3OOdtdvqHu8JD4Gn3TYVgX7tRyoEcI1sYqo/4+3WkNQizw7agbS3CBhI/BO
HXCsWzMuBzgX+X0+jCM9gowDxCP4Ueqe+x3bnjkVyGWFvxpJEidRcEWJN0XPOi0c4jpwHXDtTED8
VZmzASobwb33THj8gJ4eXYDIvJ7DBtcXBKGV90Kk2UdD0s065lUpE7dV+a1SHLOoBG6aLqeIbIJL
KzOm9xPEue5aXSzAuYAlEqRhnBTUeGn4+NFINFtOujYijJ/aJERTG+spcX0nRX7d0Qb5p/FEy0Ay
nVoNVwIuuEEBhtiSLXrqMRxQIxIJfTlKDY2HMZkxmuih352Ra4JWUVqlwae/ENa9S18GbiOBHhzF
x5GuhDDJu5+srY96oTU0cdzTa07GkGAsM3XbhWqz4F4mGRtK6KQSRzHcYEenixo/Yhv/dUG7FwpR
ol9H02020YmWMCq/x0P0haEu82vjwIvqkDc/Gn/nxIxv1HAGwo1TE0a7VcjBwly0C3xPcwUUB3Q1
LgKcqX38MbsS0QvJVj0k3NQGIULZple/5kWDxIpr23wvZPeX7FOS1rNtlDIEO5ubsvcUciQiaEXC
fTRJaFETkjUSofdoo+lyZruKwixHRZ2TVbKB3bFq+JVCnMXHYudJ7wc8olEnsDDPm5Zim+FS/dWB
+SCpdvc22qsp+cbSm4RFBWRI+Fqg0MjJt/Dl78CBgGFL6SYr7ZIXKaFR6v81NXMzfrPWC4/crSLq
qnSGgugVUAny5II8Vf3mvbc4mN6z/9K4K/sxpYt50KGdVWtubYf4MSQ9DK6WPny0BL+fWbOkY4Qk
m5/cu6ugQ/Gp8PYA7q7U9LpIfD3AZSY4fJB1iTHH6NEXodyIC3CcZI9gWLNxXfPc4/t3lnYhmUmO
X6fW89foTj0KnobClnUG6ExzpDsg7qiEo7Awu3knvv+WTe6l9baB1ny6XIQx3mrs7abOcqb/j0ez
aIkSFf0FsRIcUrCkwR2BMz4V1wvHhOEGFhiGhgtkQfNRWfXgnaCAqUoP2D0409zZV5iKW62szBFT
xpDSx6V25xHu7oyxPPcZr6DYnVpBoeSiFpbsLCDSIEWdb2jb+11vEEw62kfk+3wqcppbUcl2YNKI
AGkcFpA7YZgYyikoqG0jAA+GpW4c+llN6sB6xniRV43dFZ0wOX5LYzVxGNm/2viEdWC7Frj7P4As
/ZDzFWhqU5EqhtHW05iXGEh1To4on+c621bKpB3Xp6N0vYMzrIn/a2ypmrPI25HwE+wvbDdOLQ90
ZBw0fe5WfaFoNf18S53pcTGFmNDtNBkhcrYO8JH27jwtXop7D5/Wor55gwW3bBdIw1rKtwDN+Srf
RzZglvJ8YtWmljuYaLgNIgubmB/7HEJKycIEYa+ad/wlsdbcZ9WsegpkEr98ztEPpqMxy7XYdStC
fSbdqoFMhkMFtNPnvvSuwB5mWVNl9YndgDQBclM4QiD8Vb77aHyylswSxCWXGExZ/mfgJuiMq99k
UHuFYF9SzyWTapX5J22MUp2BW7p+1ZBEomiSU5sOfFes4pgY3PECTpwvKxt0okrkGEBxPB75JJbJ
FxfSH3MofW4wrvWr9KkNgoDVZXYj6oci5Ai8dBeLtw12Nksl3TqdaDBN/mUXVPkdBJTgu0rNPQVB
Kzz87OxVGderS1e12c6xOhsWBuMa0+Buss7Mx7nZccaK7WpnlbvO7VheKH+ORTd9BPjItn5xSM0W
S45nxsX3knsvRrnNNW2y7z5SgarKT+ZdGt4aIxI6K+WQBuTuE1oJgLsnTzDPqV7xOPHruc1/52ET
2x0L3DZ0qm2wn5k3USt84wjzV6OzSoP/Hk3sCrNh+cRMObgq0nHfeNXomDWQXluOrJheAVMJh5oN
gm+uDdpFbxXuL1p2SoDHylC4csBUaBuEidpHpxXrJbRoD2jf+1kxg9eu+Z1k+xQ/TMNdblELX9dI
od6g6+jXF3tPfa/egeWorxy63jtO/k1zh9PvztcqDWphwfMgnC6V9ZzcPKpHpLrJMHdFTi3pyvTK
xqBGQSYEnhYGWkMKQ0elPnpt5CMVQNY5RRAXvFAxHGah+u50RG+Tx3Gubyv97p7TiBtI3CQJIE5g
cHd0z9+ZzEwCvD1gZHKLKn2UlBiQn4GRywe3xl9QeFGqxWW9OcsB942bcriafV//SOEDpY0Na7sh
pwSIcrA8zhgkT5ksD0ZaDazKRpEDPA06tLh6+Y422H/FZ4gqoalwB6b41UQN3WolHDHUXONCJSlx
jHc9suW8yl5QXD6R2vEJrtsUQAhVas++JzKPFTu6HQ70seWC0kaT1n7PMMQchnY4EkaIOu7B6Eu6
M97Xpg7O1zrbipoPsvX3kf5Qy+dC+naI8gHW//Z2vWBbMx5W56saP4SwLfX6119MxJetZlggJCwi
AnNiEsI0L/cTJlabyOBL/1dK+ZQBGm5nWPOz/Jpb5aznZvSyNNY6izduQ2TmkY/3dR8HbtXkQcwY
8WMUCVO/atjR3gyKM9gmjiWhFYnZI16Vhc9PDY4xPOy5M3OAjbU5stVQO8X9PwpCg1Rz+PRp/c4o
DYGu8iibK7999UFylA9w2IVdQ4DOvkcUvePcm2T5DHfHxyhpCTyHlKhegiY70L3PBh4YvR5rNzf6
vDN15VhfIuae3bLOZem7ITWMWzhzmkWy1ElP59I96vMaSOHfSG+XKnuxPrvlgfLZQOrjmVGNQw49
xP+JgOMs+TNvLCtBq6scT/HSL/HEiEN8vVHixNNxqMIh9QPdORcx2WhIO1eaY3QZ9NWuehsi3+NG
owFm/37fSfsguMu9cWJJzc/pNIDtjDuj1n1zjO47waEHtXgofmspRskxfVDPJwjsTi7MwV7O3Vlw
Z1k5Im3Siio6lDE1ZueqauHQvaryuWhj2nRQL2LfpJ1mwrdu/5d2fywv9JVZkkN4Hr0hCCb1x/qv
dFiWT4xPwGo9EPkYPRfTYMGzeb6hxb6lNq/I4eHPnqf0YnX43mYplG5qYAvd6xcxZM9vDzR4HjO6
UUPdqdT/zh+js0Q1Hl+7pg2En0Xko+p7G1Akb49CvIBNGA3yv+DWRpu8ZEBLJwL+pLxWfr84bznZ
hsVr5phcZZe80TvL63IOEhVwO0GwitxhgX0vpnirsbV6Vqxq1I7Mltto2xu6675YzlebBElIQH6f
LF1mbv5aAr/4aw2EJNRqc+pBOBkXl+KawBYuJ+GKjV873/dDRzjHvXPpQ7z1Ep16F7Feg9qWNe5w
Y65gd5ANBP8ai1t+mzs5o1zKxq8bnc7YvksuBU3Yk2hhR3hEPrwY92R9MCXgizzf6RZrarYIMrq9
tQvyCj+2IMuLErL55Pqsju2ORJBQcCqw2Txh5X0MsGg+m4afJkak/M6VuQ2Xst+co7n4pVZYgJbN
tZyMh3nkytf90OdSchMdgQcz4L/mX+GFNyKZ9jF4rrCI527Ip3iy/75DEhI1OXHTobcHPkH7gfPd
BT4IR32jzb3lEXA/Q+gdW8uMeXn123Nja7Q6dpIvr9q9irj6hQUtUjXlQG9oecw3EH/Pgi2AdF8f
pXvSFiI5NbvvQUqaZ6RafrdpePIuP34AvL9UbuhlxkZulf3tEwrhmxEEtGHhIXUm1epSKInAtBhU
mcZ9jNXFSLXyvSq7S+kMPXYb3cjyO9gUA0fgsrpg89TbSxhvYHFCmsU+eom8h3aniHA8ut5SbwHv
zLLx8C1Sz9atJ7EkiPlDiB0w3VmTf5S5FUrIV0SHLbcZMcvonIbk0GncNA1BLnTfBmVKqexH0Is6
AZWHdrUelmeXHPPJxfjlLnDoldRcAPWDCuY/q+GC37zB5CSodc7xkmQsRcv4NmxGZy2mQyev751p
oZ5PUtS2UkPwMepgo8UqEJ84s4tVCiy6nJKWuVq29P0zF11TNqh3HjwvVYvaHzwsNhwchylZho6D
2tPCI2AdXii7+20RRXiXjCUay3cmDknhIU131Xcd5vGLuOxVC8b7dlEAOm1TmK7Rlu0vNhnSj9wE
ih/bclyRGT1e5Tklx5i7k5ZRrd5pQa8YIx/XcIivd+LwcudDlWJK4kvS9kOzr7pXJ49sbWczasah
y6fMk0S1tzPDu9GM7aQyyJo8kPLubJqV5CCkw7Gah407qWj6mNRONWoZFKjGx6cfi8g2C90Tpe7R
bq7X8j8D7+n7ttVIz+sHF1dKuhodMp/bLgcWd/gKErt13lU2uR6hqsWPGZM0pLhqhTJac6T0Jpry
zJsPWGjFeeu0xzTQa2AZlPBGMGH76j++QFYXxBhIccVuXe5JKG+cVhGges6XhhCQGtPTSSfPHAIx
QOpu6gVJIz9qdL60VvCgPHdLXWsMP8py7GeY9dSXvPkeCLceEoL2wczz/gqtNmuVgS2nOEHRWYZe
tV1E9J2TQq+Sh8McrdrVPdBr04/D/T1MkIjdCmLzkHFxmuZ+qhWB/xMFzH1jauLwoT9aLEdX2Vwm
+sTtmp7hee82XstBeJF+NDoGgZ3+M2K2pOrVKt+l2BHg7a2ExrkFJBds40UzlZzUKskSpcebU7g/
oOj/1chpUiHW4KZJJgSTYorVhCi4Ncke9t9Ti4sK1FEup5Yv5McaVyUdvw3oS+1Tcm6NfyRpJrMm
8PezmjrFmiTvBddqMBHM91+ABczAR84D+x1nY86K7ccSVipGa7Gt/y/qiiRuWPezOGTgaMl0ODjZ
5DkwS86lqnwGnopd9c6HYjvAQ7pbT0zExMuNWABQQmLq7TcRwxlQPMXZ/7ip+SIgwnJ7gC4do4bJ
qpDBBLjvc92fWZ4Rw7CF9Y9wvWbGADHHdQ5QPRuoWmTN9Jc/vAxRrCs++ZQ48sTXCzTZsP38+/2w
JYoeXdg3ukA1w7fhxqybKJLmcnrynSMnS1rYCskAVOcDStQazT7N1VqDoN51cAtbsXppnmwu0pU1
f0UGh4zIos+FANsIGM2oTG46wo0+pzYehFdjzy1zSErzeLrf2ORVTvtgPMf0i+iZiQDNNMnnLHmr
IYP2Yj1bAYMl9Uch6QX6xyNe0rZLO6KyRpqo+EVkoTv86nQB7uhpEOA9L/PzLT7Q63j8uwZLfWx5
HBrhHVOz/+GFSR2I93hiXVJrg4VIqEjJRAY0H14tf8qTMn5Gj0VL2P7+hfu6bPiEdH+RmLU9bEKd
dJXY1Z1m7db2nasHbBV5hPipQDGOknk802WCEsSSrAeJFsBIHUA+aAh5zXRVFBG6qisN3mthfGx9
gLQqQg7MTV1EipDojEOMLGRG/g95Ivrs/qUEAHIi1XW5f4BdiWoOJW/TqSrgUPVf9q37EWRlKhI3
ZYY8j2QxbCt8VjkY5rXzJugCwB55kYNgTNOPvrxUjdNTmmPqM5DpQ0QsnWYd7Izo3c+QLMl9u12j
OPdgw7s4+YDes6j47wo4Odq4l0xOfDVBARF6gnoC2XqORX1GRj6MUG9HeOuq9qyY+4obhMYqhbek
7xT6sgbo0eD9vMOmh5AGKxdVzBNwU6JUKl1R5+bOCVlwlNf45tfBu0vtc1J12FPHdgh8sIhuIKte
hJx716ALzzfxm+TkELWfBL66MXNXv5NoFXlBcBoO4U0eHzo5AQpF1bQ+gXaQC4Jzo9/+no0ShTXZ
LQQrHeqTNKzx5dh9SVeQdcdUF3IDtOcpH5hs/SX/hos05ctH6G246qVoy2t1Rv5IA8+ms+A+TOSl
sqKSaS5h5dWlQ3EwudaOcQMdhA2iSnDaQeb93xd8/nq+GELn0RVcM+gaoE/9JmK+ACCufPU33WSQ
ktB4Lgmd+2eCm6D7cslnmQoeRqBHFEf//B5zFxh4VdPcSChcqEBx5bGZOMHt4Dq+6jH5Mq9KwujA
fCWmz8/y1tNUroSpoUhpD+jqcpTixJ6oCp5K+QcEbBiBozHX5ZZtJ89lBa9zNqI2DqRHxdFOh+gW
8TyYW+jQn8IPm0fD8DDP2dOe5bHRZSLgAr0n0j7IEnMH2L80G59NGk6sF60Mb3oTmV9M2KFBTQqH
rF2R8bycJMSYVeNplZEBxKvkon2NLtOHZ4xKfW/FNCJI1Hnar+jkzBw+R9WCXjFs/92hbEPRbi0t
LYcFcntwVH01EZx1fp+x9EI3OK3gI36uRTLVSZTUJrUk1TjStHl3BjPMaDEuklmhKTv2kcepz3pS
FxAXaVIvvxtdnAXA9VAbQOmJc19V5Y9drX1OAkkmJhdveB9hxNuQmXzSggiBt1g8mOi7eYZaqsCe
5oCvQx6nGAQjdzx9WXum91xmadYd28LhKTuU1DupMBoaZBYYQVm6pRmgwHtv/5myFya4T1ua+9A6
04SAmNXc/lwF1tsQVnjZjGT/G3Gi2KnvNIBSC91rh7n109fEkftooolczrBFkXkPazvNi8CKXH1o
BB1jk24hRPZjspojEXuURqscavtXeYEBqwqR9Ryz2cLxnUPZ52A/OXxh5bXtFpmJ5c9p/Y3N0drQ
QaVCsT6POpev0DmdpENKPOmfaBJ8bezul8YgvB20S5b7qQTw70tHYk8qaTWKNLP4cSxEumw5VTG9
mOKVBAYRmUxmJAT2CY3rbYMAGVIQZzB23VuiJ5Ykrsk03Po9le/7F0FArAh5klH1QMANzdwh7i1E
L7LJyLPKyyUujF0IvTXIRcpOYYZJXefe0ek4QGCZvtpoDR+q93sNio1Sq1wwB8R9XwNpFRVo3lPZ
EG2P0Ikv4r+eRlnGPfBGgJUYyHi428AGtNLdHPG90owLWz8Z09HLGeMj1Co31/D//DwvRsmEU9N8
9LHOG4/C+qZdw7xsixKEi4BLfrz8HUzoof2weZlJPAPXTH+Jy7yrrminTVTDx/fTSEOKL+uiBcMP
qEW151BdqmNiMmT5jBEw5Sc4RHY68XiKPUWOV6U8OnoqpBd4eHOLqsUiIpgcn7ZFutKq8b1G4Jaw
mNvUwwlmjVO2qpdbfA9AV/BIfcjfA+mbYcRI4OPydhbKwmEtpBiaXvadE4bhnmmoTgYJpeA2F1vf
g6fpgu42wzmcP2nNpmwSLvConFr/T9I1rSUxQkr434lNuKrw9brTcUSCecVl9V0D6Ba2+W+2c7Aj
Msjzl+LZ00HY9isP5EwlKc0YYffGcRkHJcuhfUstotKWTSbDM+C7Tr7XLU45C8bjgEHZTlYHFxvD
GWiGp8/2rIyHBQkfwXPt9GJTxXWyCuxUNgB22pHbSewTgKuyiRsV8LMTCch9FxImFrIXt8fjGTqc
3rc+RYUfP6S551EGxyYS0sLTBHllKXeD8w3uf5cdnF7j4A+1s9kR05TdHxxdtBPd32O3pxmz948t
PFTwxuuZQMLa9KbpFrI4Zzv85jXkgYC+EdjLLnqIrpCnZF9cTHGWQr7rqQxr6emXWKFKFfvs8/0D
nBlCNiZVFk543w3R/aAliPC1pwbVhjDO+SkE9C/6Vy+2WermdrNfox8B7msEj+aG2js1daMFrvdB
YYt+cT+hwl0iICDl4sngdvd/wkbGMTyhhMBHR3R/twFv2UrFfbRU5zkXOfTZhcvefsc5y+wcMYd7
pyQjcvw+GLY7cYKY+xK7ybCXooi08OrRpL3p5lmQmrx3HVomVm5NyF689qbEgdZDb4Ey5DWN8OjG
BrEhl8kaxKxo9VF9quEyhjLufOWYEEse9QdN9mGSjS7uCdntuHZ9/gZMV8UGh4Z5Ej8lzCzRkrAd
xxogxIJh7N+6792Flz1DhdGux3fa4KL6pP1apCqxfm7V0pV85FcDxAXt5t9wv+BqCXlQqVCqOtW3
C/e6gwIlAhxMq0s8qHFjWMH3Z58JoHRp12cxxVc39i37IIKJ0ApWsonFxleojuqI4p9cpG6vZG+V
uIwiBuA5fswECKrRpgQ5+paeOjnD6sl++Og8JDdzkwGZy6DHa+qKd1JvTsQqbqHLy30CKEDqHbKf
juzidqcqNsPDXNFXaHLG7Qh0CD3UHkbzWlysP6nPBXUz5UaLQOUg9a5ETXN69rvYOnfCzQSUxeAX
vQlj+FFz7imFdqD+UJQr3rBSm9C8IdwOFg2ulnfTHrvAaQ3lIfURNMgcL86XDFtbdLfoCozciXyh
ZarfDN7KBGdP8J6rvSVSYuLf0XVDbPIzZL/Me4mf2kO1cbvCNwq4YDekAP2g3NrhwMqk/k+ThP4W
35VPGYypZQBbjRiDSrNs2OEI622yBK/+d6pCdNaCANKU4pEh/Ht9lsU8Lp1iW8it19gbvIA3qyzq
6cSEi8X8sVdb8sBllmdntItlv+wofW0LTxpV4jeKrRYl+nkr9gWBvdTJJaiZjZk0WRlrN5TAqIPv
lrI/DGmvNL/3d90tnI/7KK3jLoBYME2F/9OKeoZiBWAYip/ErMOuqAbHS/TMRfEnnsulV98rziI+
zitYz/T7IEYVjikEo8w9HKwnljZHt8wOflmkoNBDT9DsYQGynV2XIalKJlgfQD6YpjVfr9HklG3z
A4vQM4ZTxRIKjWq0aGT13r8pvtXYhu4WiyknkoH1VpK4VAFT5+fQPYdiQU3W528DdTiroEuA24U0
leQIYPa4aEeE2Veg6nyymS9OgGWCDXnGAMTg+KEpp4gRoccJRsmXYpxvZnFclj0ZEbIE752aPwMD
RJmCIKT2kV6xNRrWHMcVEV4p08jr626V5P4o8DbX70XQ8goRgFRQ98KnVv1Rza3tnji79M5cFe2Q
4MAG/GiQHP3RJh6QFsMbYyvO/k5gYLOMEcT9lBZjXH8Lj5i5cjckYzVDjJy4MlqDrYrwBbEE2/P7
++EF2Je3+m1xKsKLs0wkx5cmH10eEYj15pFJWgmWmqP8sRb+6ko2cd3cOC9K7SO3uCKaCal0cDkN
KxKWnXTATMmzA1N6bFPewpLDiM7GVMoXGhPOFv6HGUcrVamAXDUnU8mO3PMM0dF/51lhIVEeGhJI
HH5UEermslbYyu/qPUEccEyIcLVKf50j9U1zk1WdhGsD+9f0VaoIRxUtU7buqhUWcjYsBiiWhuMb
uaXxmTxkLKZtFrT45iFzM1CzbPz+uZLGE0JlHnewbO60d9m9dxJ2KLr6Ut1h8Vbgo35ZqU3UVY7y
2Ik2RU6ef/d+iiyTEXiYHVaEdKVTzAJDOSWSa5DtiLLthDYuAxMXVwrD7CWa7Db6Om7pMZt2uI13
8NOxTBTENnsTy7hM+IG5/PVXlNNVVJquBI6WkPUq7xxSTOnVvPSL/d74awhZagtQQW3oltoUOYMh
VLexajZqKP61m7dqWspmmw5XD8j2i9//LT4mtuNCMguNjimgZ9C/kHIkN1imhul+uUTqY9wxppHX
+vqbT74ywQZSp+9tPfrx+az766PMWA919jvlzdlIRekcHCTqCEuHfnD6zzD0bxAXvfzPKn1Vel5J
T+U+733+9XKorGDaVXOVPZsyX+t/qG6nMpsLzsIvHkpRhVX8oSZ0OecKGE/BB+FNT98kwcnHcPiQ
k6SP1ZpkBPp4AVyQ1mdm2oEc2Oo21XsOUth3xG7Pe0VPl6JYnOQ0g/WULm+qwDovgskxVVvcVuEE
jD3gYddXZUW2x3MEeKUUeJ7LBtBXRH0WbzFOwRXekGl8EU06W/3n7EWxKrHT73y1RBhi/mN93EHZ
uXEU3VpBd8yfDJIZwML/HpuUKN4HYMeQWQXFAcWxhXNe+pTyw+Y69kJdXH+amBFRYEbso8btVPaf
nBJ+kNh7kqG+s0QB92wVqqP1P2ZSovb3ZlzBtjLZU/9H4+iT14hLxfq5GJJhOnE8PBZaidV73FMx
nKr8l64Kr4cL4stuMdvY+/aYm8O8Aal92/Jl23g8uiCzSD0owyDmjOoa17xOm0/FAWT1rK8OggnM
7XLr1Q+lRFG7e6XXAkyBbHiaFPPN+jGfndl8h0UKlgoXqqcQHgCD0aFQecAIDpWxNk6G2ujJdYrb
cKMoSE7hAbJ9hxRNxHt+rGu1njhJSgRK2M81ZVZVSHPCYmR3oRCwa73To/PPhYzjOH+Gyavrmxdb
SWwGGhikrEPfDeXjkZ1OF6oY8m7UHTW6/Qqnx2ood4pNeY9u8lsAuOJFxmKuXEhQ8YUODrFVyybk
7Ky6KwSTswznMUirZqRiKHqM6M3ffZIvhyhy/kNYyaSvU6W4JPOfy4El0wrMPpwE1VaW57eL9XCx
+UCuzZ+XYrjsIntQfoozD/mpSUkRQyMTc1hQyFltptbKKlZcbukQpERb4NRSMd9rEt6yhW+GZs9p
A337qHIS5rySxdX9cvGWn5YjGdKnf2W3RQNrak2hpfeRP92kX9yBE0ENWBZod94VoJ0VX+4pSX1U
znr6XL91mM1id/LG14mgjjcR/f/rfmhr1wIWkocWs2fihpjRGvuWLnMHgwpPEjtf7HxBym8jqIZt
7FY0MMy6SYp9SwbNt4w94iUjvH5GHzwQ2aIkI1SmBr71OLTAECDe/egBNs3KeFGn3lWZnkOUcudF
VIkfTmeNO7GmFTOdb1eJ9HSqhyl5qq+g1xKRCblLwZumr5Vb8YYi0q/uqzZn7r/Vbrp1o7nFeXJ5
zreiFpb+WhqMaToopFQE+IvqF2gmLVPP71RW/8BHCBp8sZMbNwHONA+Pq7tNEYrNDGl+syPqSCt9
qq/wZuePjN1uRI6SfV2ueFPjMLW0c5cak5DdOM3mHjjwTyVQ13XVhiI8H5XtwAaoi3oyd+iWynyx
kEB09sY8Nz2i4Ineb33wwLDvWZXVDEAEZ6XS3q/23JbfPJudp0SV0b4wpr8UCVmpjibtCwC8HlHv
XNCkTipV2CdbhBW+EggJuraKdcW/g6cjZNHMVxBGTCTTA8vq87ZX7+LF8PkwlEbGx31oFKuDsilp
5kFNMdGrVNPw8hL32plp6xg+jt7h1w6SZNiSKFB1CMG0Uw+CqEaqWouXTpCQs8QaNBWlxCfg/KIj
99400csFYbN9D993Y7DxJOj+oSuAbWSmv4Xyqo+E97yUd5d3vtWbT82zZWnmAtZDPV3o1+3Dsnxm
HmmFj3tnMkgHtbShZ9QHOYsmfuXokPAKJtOlmi1SILOzvaYN34HcNU/tN2T5WAzlj6MkSqJN8cz/
J4QMeBgS4/B8cMoWd++lnl86lcb4d70KuVfQBp/hCdjP49kGk6ijQGj8Oas3f3QMO9I9K0YA+CJa
OeOCmKqmLlKc+1kxoYcz6VB20yBjQbWaIkiAWrYLl3RGAd2xQCR4He3vJtkeN62N+2HVZL/FxR1s
jo7fEwRSkEKxpiYXcmDunWZo+qMVesGywKVtZx4+fuvsFmk99b4tfqUbD6ZyDz1WEcQjmaKgqKOs
EqyDSBhvnj2iw+2q7ld0rTx2otx30YrhuI3x1w9tFyHznWZW+Hi7JfORXzd03nog90wUBWHelypT
bJE6bq2yeI/1A8lbZoLvOfkjef1Pvk3waTxSIb5ktj3wrPUM1dMrclBVA/RHz83FJuw4HyGaCv2d
MSPIDSXNn5jzk9KSWCd7GWxD9E8pfANb89364fT+aMlhkIOBZ84BgDto1NAB6xKiU126mvUHc++r
i4xjy2FLyWJ1zBNYJXtRoPU0XvA9OUnhIm/Nq3Tvk0VKIvuW06V0WqoA0ZmH67weuDIs/MQQKKms
jS3dKQBq1m/7Asa/SV1ZeSQvkm0xMSZOFguBUS+nm32GaIoUhdSKtF/occ52o+N3409lFVTNOHSS
Zu/KWLv2eI5Ge8ZLnI7LLXUEQqw3kGUdypaSeTuWXzYdrXoTRkpkMHZaG512zPpN6BEj3CJOVyCx
wkxhN21Ur95ARIsNAnbrehGHapmDl/DTnqQ5giy3HTFvfk9D1RLD3W502eJr2YFKiszIEb2CtoUy
BoVI8cvt0CMwSkR6l5KOfHimAY7tEM21QpYZ58ECHJKv9YgieJLZBDo9B1/rdWYTEM56rIPpcsRn
Aqo3LFIYN7x/Rbwl7rr5zgZEEea1KJIRqKyMbdLyucebB0F3lwAraNQXcEuLc1A0bQS9svX/NaZ6
VLs84Gno4gwh7JiYGhXDeL+MEiyDxWfGQ8IC5qEC8Yz8xK/eo5cH27NBySmf1OUNveh9/3j1PL/q
8zIcc5dkk9c8nC5PMaZPIjfs2ZG0PgL5V6AK4YK9mLPixAFt7oSrOMoSGv/MzJTyMWlXkZAVYdEl
Mqk01pR/WAciOMW/17iiAoeV2WZCpoUkMSKCeGvSUzYH3Pkqygw3P4rDkwq/IQDaShFJbi6mxy85
YcOIjcYs3tV+YxqcnUN2j7Nyr7rmPXnpROKRMuGIS2GozYHhc+T6U1l/VJeOY1ccWUPpogTU2gPV
Jze9jYurUNdZgv/biI8ZgaZ9BVJ8CTumSAlWji94/9VOzIxGJNLcKls7wtjIHpcGdEksr4Dq5toa
lVu76wFYE863wNOQ9J95E67/ODcol4t/DjfopLsj34B34Mv6IbQX9iy0vDXoNIStmbdL5MNyqKbQ
QAE8+L4qil5+ecerYUXq9XaJXe6vz6LzmWChmHNmfUwzBEcppbO1FYDtfiZL8sUpCz4ogJTrCgpC
Le4wsOf22lNhUBNl+vdORwwmVwUqTIB0J9EWxFkOR2MmVw1SYGENIS0vmOoCaFcwvAOXRXcw8B/v
6U2ryWfsCnDhnys8/cfqBaDS05PVcgsZ+3O9lZzaWaNOhPAp3oGOLCphP73ZLbVEPVs01iqeVPb7
HVjO59V+8D91t9rqZi1DHB0JX+wgsWXl5A29m6ihlaWPrveGNFTNiXmu4A8MtvP0YH+odkBwYdEI
nhq1dmM3NqY5m/AmxAieBw56Wp9v88FAmPxltta0a2fJ2P9xO7PmHzDUOTiGlFTL7C/la27/DILi
xSRb1qAhzwS6JXoQp6M0emlM0P2YP081rv75HZeKhem1Y1+OVDW1f9XRJm6CgcncIm/1a3vAb3Kx
t4+mlCbr3g0daL/oJDnuqhYZHvV3CdeVvF4hBNzuiuZhX/efR6mSxNkRNi4q8tHvkCdNogzjQ31J
JpJuIENpBMXDv8qIzYuGFult544LuJGRGHOtZHCLJq7wMBjniYXAPsGH8XXWPU9Cm6ixoH0gVVff
Q+/ICSZztsaQs1gpphYD4ldHe+l0WL6P84lwEzCTXYGikWTvru/Oi3uJgpqBf3tGvsyDOqdndztd
i3dzh2194COqGVl39VBxBQhb7PQskyxKsDEP3c0onguKcfFGHGHuAdiMC8WHZVvrzZ7+W1g9UPXL
9Zt3e96+HI27D/WU4an2VYPWI7XTpc/SN5GS7BEy4Cvk4XibaAYydgrkYbo+tPNFxNo4v4vD3ccN
3bV6kmtG0+RxzXnfaXt+AQGlyLI4TPv9L+9FGDckoRlylOdOu6lZvCOq6mYAwfvtnGRcWHcJPIBo
QpGcBZFSkuJ0eX5WYliWPZgrqT30HpJku89HKe8PRJDczrnMzj/z1Eni+LKi7esXtR+K2Ws79UKZ
T3rF/QiMk7dV6Y20/307omcxlgdXw7ZX7gVSyhXV5eq4nubsBjrdjECjv6zgLiJcI0rG7P6SzVK2
lNITi7+DzJl9laXddB0meIfPMhEGUqJpc7sYqyQcozy0kbA5WxzLLgfonOG0A1eZe7iZsqkbcB6v
bhlHdIEPcs6ziA84Evb8nVa1u2fB9lHcQI0pp3aAPtNlSW9msGh7vMYGHggi5MKeYdT1cOexgVgC
K4zFiKt5oOVdCQ8JeyLxzeVNNhiRzmw/UgOCllAuKQsQRR+wO44/OraI5nVM8oQrkNT1nN4Vzamh
tBy2+d7cN+GHWJek8PKeKaYUyo+7LDYCDFyRC1nUsPDFjCnunRHnAzWEh7XARvI5Ub1BGJbBajJV
rdjGwBD/0mqxq2mTdfiwc2b5qyKDZXG+s00Vw2HWQaV2FgbUPGyqnqt8BgF25JrNrSq2qHG2QnGp
H2osn4+VTf3/HOU7AUbA04UMhLHg0DGAimuxcP+tX+RIB5D5mn3atshFm1pldqz+bgpRm3KpsJMc
OHxQ711GpEioQT+b3odjEPE4nEcKg1G8fIW7hwLfXAJJOyIiYoqOm4ivglwVpXjTjmj3y5xyuzws
WQOJv6Txdvx9Qakn0eFyPJby5AP2Xxbo94alSP/fbdDFnP96ItdH/eAbq/LDtjEWp7iusrReNR2K
LZ/Wo/QthD+k18neFCkqySVaH1898ms88huFOQyXxklnSi7v3mQ4gMPz3DB5j2RE0ImB2Vv9cRvB
zfhZd8BcChUye1iR8Yx6/D2L8nWlJGxjG9/q+E44MekKX7zjBk4SJlq6dSibeXjDdemSbFkWhZG6
5Z+h2VgPuEvmb+u4gjJuibBV0QM6FG9ZHC9NsTWpY01EtKZHveceTAV4jPXBJ7ddM1fkXbM1RuWI
AppVIZFOMC0LfxghBIXNa8aAoGnQwamLWvn4i2QM9gZOtDNy8XL3Y6YMtTDNIXuKuarhwCHIokIH
Ug3lmcAYqHv/lJZvvS+XyOXEDC8obHmsXWDJJ/Dl2hUk3OyGgTsKsuMhvSjryQWnoBzb2GjnpIEY
ae5UWyTh4nbS9TdT1JD9lD+0elykX7NSpteMZpWeqm4qpYKSD3BYfo0HVNytv6bXPU8CHwdjeYzO
SJI6/HwKmjQflYG7H+LkgoFr40JyeaRpEzx0g3QVpHzm+vytIaI5u6XxnPi2p0yRTFYDWOjenZlf
pzwTUzWRwx1w5avxLVMuH5nMnEe5uOrfIgf6q3gpnqL3AlbYWkY3mOVXNMz7bSsjX5eVgxUpTJZ5
PeEPsPp/OKHUigTr0iQaiTNkJzVv535mugmCd0c5BorkJ3kDRmUuakAX2jjv0wD+Z/58YqiyqA31
5UAfcSQP7uIJAH1rSk3vYtiTl+qqldL7bOyOuAF581PFKuw6bfMn5oPCi9SCG2krPQgcX+fOmNx5
i4/q3A2cdIkHiLViqVP4yPb6K1oBcEsSvzvpFEGXQfpxYinzFmEDO/nbTky5/hoP0HFpt+z0V3Qi
GhAjmcyYaQKFgmaoAaSDg1p6aApOvdRZwBHXzqJ36varVOAuyhztp9rYHGRehLUtGrKayU9ZaGuj
Fov6BiEu6FPmvCA+sxhTtSe9ladMbZUWMyYoWCmAGw5bNcuAoifGkoIMi1Skq4MH9qSt3viazM1x
0QH3FmSHh46v+WTGXN9hiYeXdvgLAz7/Z/nmYMw8lBGFTFeitfX2l478/5zWGG5sswMMCpZZjA74
N0PJ8t+dKoTayBGRnSNE77LNMtXEvUu79eXy96jXSMzzoDUUHonf9CTQ0Utn52kWZGaMgzMTZGlp
ZRSAP+jTdqQBFpaVl0+fngLf7SmpRvzwukDcIZ772+lFMC2DAXSbqGCNpcRF2ySW3QP7DYcoFoW2
NV9da29+LeNRBhQnpBy+KhI7JelatzqdodCw2IwDtS3vu62xn+aNClarJtYX/+rapvzYuC50p6KG
SdC3FeLPdjsZArgikEaqq5i0TZNb8RcqZyiD9M1ooUmemwNZyfG4IPKsIhbuLnBSWrPKphM2q/xP
pLcn7mLnXN15eb7CRoX4n5BzfoI5RGg0PHca8x59JITLSrITxGgjOcFlvFfjwH2ELGwAqBp3N3rs
4rS2WrkBcqwnGMGur2OGNiOsCSWhYMduNCY8MkwIVo4mLoJHuvdgfQqCwJC5SOAXLzYX9V8D1MRR
/Ydqeb++mVxKgPHFZ+ZDJyR+vL96uv6WvCAUqvyi5V7rKk0kHQtzA+ElUAtm4TE86NJ4AS/Q4H3J
eLpXQDxW5x+RwlluEMAwtKwvO3lSsY/MLQv9WBh7PlGWqZWU5LezvxCz5QCgMVbJUSgZ9+2N/GEs
xgGUdXU+CUIhB9m15GzFRxv7NgEcop+CjpANrChf372NwFTZJoqnnM0uQWcvnlJcRFk3EMaIhqVy
JKLlgga8SLL42T4wvarNxSXpW0OORSmzzgjI8//FQYZdVt/1fRt7RrJpq15+oBWi6TrjDNCv5zCT
insXopg9JXS9lTfcN5HrJHOwM3eQNhapWwVpKZUrGDSz2eD9IwRFRWIY3i/vcRUBLnPbtWX6LEUF
B2xElUKGRuK7VgsPvEdof+wrG3yl45iv59g6B2zWx5Tvke/kVYKQkAU+rC5a8lRqF7ABuG3vUbNB
2vbJ3dYhFa7cWUmvGmIqhOB7TZHf9XfU0NYvMbPqW6XZHOROfkRDu0X/3fufyKzCFeS492QoY6bs
Fb6ASY2xUSslzBmkWwh36xduLmLRNUiNP6rTdcE6PsD3C14io5dBevMQVaFDzECzAS1b8fAuh6ME
0m2RjgiVqKsJFvrL+u7TJfjaG0b9vUZJn2nr34o5yp9ZzawypBJPMlBqKO83ndPD8mKxlIxF/ZOG
b5Jo2k+uyjRGNZYIoWM1McGTr19mNperfXypwF6UihQTm8D7k/5qRRjwehtnp4Os7rAM9Gywpc75
Kt7ncOYt3WFtEclCWy+4JJEzphH9q3I3wRkJG7pvMpUtFER6J8k4TkxiTiWyVFMsi4wFfT6R/6LQ
o3ya4x/Hv10cujnZEOFY0XzBUhWtIavCNLTeHc3JGQrn1jK0WTVMgjXZDVRcHrdX0MEv84EPUmrN
IU0Jj8YrJwqvOamnnPC9D6FHZybcokzdgyeGeTNvbBm7pjMZxZ7ybYp0DoYYNOHEq0ZXfmTup0Pn
pgzYguI6H70gB3Av5dk3Z+FS5jF8YYNtWMUt9Fx0XnoBatKk8TIPVT7bvE6Omxo8bkp6dHJGQX0e
Fmou57NEbKEaH+J0zXgnFAUYd/bpjRmapmkiDlCv3ecx+Z81mXqeWgPgy7kCqUfc0S6l+diBvXN+
UqHPOUv8xZWS8RCrbUK4HkiNIfAK+nQdwyALLs6THZAHcd/dcvPMU+fIqjBPJNzh1FZjUTyOA2Mq
MRAzF0WZyMv2zQMeFE9RqiM1dPVaA7q3IkyFI8lb98vO5Eu5IOVokQS/k5lT/2f9nSLvV6k8+5n2
8OGZI2aOZ+QANUbe8cM4lniakJlcMtiz9LvuK0Yhv4B1IVSmLY2tEEczHwkw9CEfgfYnAfPuOk9r
Tr5K7zEYsiNnBVXp422oP37X8szA5k+u8P3bsZTpZbGtb51zod0ao4hJ38FMmdIUhdfN8xqTkCqT
UtM/JB6OpW8NyYVVmh8jrETpWwOdoIp6MU1ONAwD5kluMSdtDLmLvavQPMZraiuiBmrD4z+k87LQ
EYPURtssmUxKz9awMtckCT4k5vMLB0T1ncRdWWRfaknkX0NuPcwQdoZz4kSigrA1lI1ThU8c6tUC
zXsqpYAfMFlnQCPZ9zV2KEqUHvthfKygxzrd7I0Br8OGvFkN3nRhbLaVxrhPOq90SRm3+gTx9mqn
HL+DjXIGoorEZVrRURCm44rNfpEB5LerJ/Q8yGlnOSEk1r994fzefqCMNhPOG6RNrPmgEW2YXaSK
EHzkW+P5s4+rbGmWHxkcovY3sEKDv1sAKx1WwiyPzw5wa6UBZhgjDOJDobR734hgGwQkvcZ1Hgyu
vdmi8/XmGz4s/osxqU0bCWrHco180ibe3PThrwPWWfRc0Jr97DrQ1Iwm4m7AVqvK7bySDarRBMvo
48LPS99p3kQBghGcbNE949EgUFvD26q+I33OSlqIaduR+fg4pdrJsPBERV3ES+yB3zJhTBSCvCck
L9F7CSobdfMQkEJjOxkgUmet9w8VVKO9DxRKmRSXdGLzfiwbPNr95fyHWDrONE+YBl+ei75om8m2
EEar7TwrQZij87ygpssQ27y1YYH17U/Nbgx9vpPEO0qXHfGSRfhSpHLhokjipJflk7uuJETusy6W
kKR6eh1OlG8E0+lVFQ5fxE/4gNDYbCyYvXhG4hcjej0I3NT1DsL5sfGgdvaC3P8uCIqHJnHSXCI/
y2zZ8k0BVe/oG4izBmRffzBC6QQJL76Mne9LAfN+zy8WdDqwLb/xz1rI1R4DV8XPvxi8R/5ETOQy
R1aMpI0P8/CQmZOtdrk7bhecPqPMsr999kX9dpW7X8s+5X2yfo7o1cA6MMxxgt1yePAQ9TzPxtsa
f1V62ncgaoN1QTMCxfcW59TeK+gUB1g/K2EtDdo3+sYhmmFPblMis9VaO10K6NP2TtY/8J/oZepK
kEhW5wLtslljN+4U3cumz+4fodGvYf63lx8stLcvmEYHw51m+rdHI0qr4By+oevl24fdV7tfZKKZ
Rr1OIua8kch8cmgVuiscF4K3+J/Ikd8mxdfEAqqjtcsaGbNgMoWwhZp2DQlLE0+UTrvt/2fsnoBR
k5DsHTY9chSOVdoSnsildb75I3hUtvFdhlTGgLLfDFYcBYVeyVvzsxyUdl0/wvGAfs4pgPjdwTAG
SnULsFXCsNgO3HGawTEwsqMUL6zxGDR3lu0C/TOmGPIWzRsSOqXcgpY25XGfjYpm+Y/4jf6d39HR
HWA9uDCHESfKSwwqDrus7xTyPheGtDgoYf0tyCNaoSX3d2CBgz3AUjE4Ri7WXAESjfNtJg6B13S0
oOb0A+LVFsj0w0bOz1YmhGYUU6Tr5G0/sfQEqwLwkomJQ9B+L06U6wThbH+au3CB47yOsrbTDDOQ
g/oXuVKJxVpZeyymQ2q8O1VQAFxo5Ksg7Qv9DVI4i4Zz8b733vI8sKoaGKOvuhlGm8AqB6CvG/AP
FnAkWNxJyaRL3scyaSJdcVfyfwc7SGUXbGOEvuYo6qCxRpsbsHFubtJbTpHZ7gx/oc0kOl0awTuB
EIOrSa0SAfIUGj2Kbjpl5sqhNTJYY831n9kQhO5iVlBhrmKpqraMF1ulNlOldY86wRbNsv25K7Gm
eg/zgTDqJmdPRLDnU8Ra6YTdgjoVftDXsQ4Mj7FVmIkeK721ESs7jhYjO5nudK1c8wdks9c/Q+Gz
PaK8raK5rBDEMj2lBmDlWNB6lEaR/XzQiMjisV3kknod+G3tlPFXFbu2OaSrKC0DtSVIx1ULkKHz
plj+oY878l1MfOhj8bYbWoI4zj2slkw5NnpujxIo4cPAnSHBKGvLyVqK9job7UEdMpeSrXfITDVZ
V+AKf3uzD9/PGnwlVLO3Byqhviq2eslSj3BzR04nfAl2tYejBRjDf4WamlAlwoEMfUJAwn4unQl5
TokzjnZhc+t47O/nmdIDGlvbs+8MJjiQOlRmwbu/JNGR6UAOccc8GraswwhF6Ys6Ja2L0v5M5V7C
mIoms+K50g40iPhuGaF+rnwqjVhG68Slf8gdXMzaMW1/SeOp2gjRTmyqq7+CN69C1j8mSKgCU0l2
DVHt2ijKMkBwpcyX2SGavLYDO14pUQMADJlt/qoyZyzA3BSxdvIufrjxBcXWElah3sFORFmTEIhG
ImNKg15UWt9sW6qnTyvws2yPDnZQ34cbPQmdlKo/Qfua11ztF45341furqUnXCut6qCeHjSHP8A3
Iv6MpA+f3/HCnvUG8ta3Ha04zx661FGQYz3xAZT5B17QoBcadl9JAUdaZdtwLFZENQrafNVYvJ3S
D9GtPljy6a3AJOPTM0g0qzQwgL3X+YOObzmz/q7y8yvfr9cNgLly3zfZE7hKUL9aUghwOoa53QNf
RQ9iTUybcv+Kx5sBCvHXXRFgSSuKHl4zdIzIHAwBTdBaX80MxO+4AYKtcNb8ZJ6GR7ej+UTV0iCm
P7kyv4SkScALleG+YF0mz+5Apxa6u9cwHtYoYPhLv+Q0tTd1jCpurKAPbP4N+gl81yn8ky8GT3O8
G6hKd6Xyw5Ql2P6pu+jO0HYELbCOXpNHhCdINdNjXxHbdu5JwTEdYGAJG4/4imaoNqlpGzlaZzwy
jdzw7FhJ7tQidII2eX24wyxUTZ6BKkWTnfIiS7c5f3Y23cPg+wU7lv1oDeWXT6tG9nNsGgNUmT3A
fln27K2k1z52cwV2JHp6DyCy/94HeUEKyJvZcIMA7drNuSkqnu9nC3q2vsGzmY3X0+a/IVPSpP3M
Y5CqbWWnL3ylfFsBrML4Hmyw6i8y93MqCne1LCaEm7Psp+Pb1hw+fPcVQpqG+ushy/7fhIO46P6B
8EnQIMPWI7QW3oXxJu8AMxIEja/BNNNUv/dyJcPd5SMG/5T06sY0bLh8A7XUe2UO6hSqqrTo317M
nB/G9Ejv3IxRYWvfFd3LTYOVVIVXgX8NORcbHJgZ8Louv80/jHwxbnFpCQAnI+3fTFvj77FFgoOf
Bbe94UAhbnWRuJfzsVHlHwmwva6dIFNdvvhAjbH3JHpmbNU+BJoAP1T8G2XIjlII9bpLk/p+F61z
urWv86KY9Nkk0ghyCeysjMOpQYcbJR5rfDpFx8zGSQQ9I+Z8zMLG8s2OJLBHKKiF/UfwRvWTzkp8
Us1q8DN3jQEUPetlxcO7hS2la6Eqkb24bPpxnK8Zbcd3+45He0oajABYJ1w+9URhZZvNJrOGmw9a
QhrGHX3jMZ4TwGHSmFoV02VUU+cJCUPXPr6STqWWL2APZOVq9TJKgSXU/SntpxP2HYl7LTmDW0+V
5X254Q21zYlo1mEvNyNybWxN9kzu2wk4SFTiRlSByUOpYOH5YpUGDgAcFhZmgp1pH7u3uyCjcImi
QCbbc0qO7AonjfwRHvu59cmB8E0w4OuSTLCVYBh0EerJr8J2UAAkFICQ/6RCIxWddNgXNZXe1dGn
v90hn4WdK4e5ZCVT8giaz/+tlaBBtj/ZcCxcdqqcvnBRtycMSDTdAV0GJDfkUw+HNoSmqW+oRPCw
PRmUP/1OABnean2XSAio/fN8PUj3p3PxFemAhf8+omBfKhY3QBYyQhZS94tTp6RpcBN8LqggrDix
nFMWV7KnJbd2XNH7OHnQCazdGWizNhRhft5nvFPJ/l5y9Y8kEe1OkwFCNfexv3LR0JlGmHwEIbqC
Mc7p508gCSDo+dbT8RX6ukb6NaPT5jDy3blJklVeveefZF1u4OtvFd90pna0P9WApeKqJxy4J9nL
tTKy4F9Nk30OhG7FqpDy591jXSzCzk+yy89sOsx1eU/NmG10ILRr/Mx6OZGxYKr+U6Jq0c4e9z2t
9HdMzJVYCMIQ+rPoyDxjT5VlndwMNY4YB1l6KqOJpcEhDTQLZqZ4ACg5j9nE/xqNasuvaFGyhaJ+
CE7XhMYK9cj+31PIu6MOy4hzTqIJwfI2Z6qEMzcJRQ2R04PfONzvlHcgKASOptzBjm53rVLKnHyb
/V87kDgxuC0da0e1zEBgsfkzwEX/1SWh7b6IM1KDqHafCbNdt6b8LYfNOj+0Wgz1IWec82TuRxEY
Grqq4NHxRhrLUuqhh9oOBTM8VLvpGUOSzhFW1hqXYsB86j48Ni2DmQFHSNGjVJjjSvC13GgUitwU
m/yePxOsFHP3rCRCijYQJr8J4WHrYd+tLWqQmnEMUY2I6rVaW6UcYN6MWqEWzl1/IAjguRqh1SsK
901uapCM/EskgULXEB2DfA7UDyE2iso5rIUKwx8l7HwssjOi0NbUr/XBBdww8O5V1LO02mZAQ2rO
QdPsNSth4CIB0VM799iaD6VafPky0GiOymO8Z7nu8jrR+YGZMoLqjxVginI7+O/8Kn1jTVv+0TGD
jY3+slJEt4aJQzfLWkGstWWWLuaSOEc1uyYuVy12QOsRsmkkmpzOpNbbkU53NeQkXVTMXZeBRGFU
1Xlwi3VlyPZNePGNYe3Z8AlaQ8f0UsIIeMl1RkIc15h/vWo9yHkXM5uEFVhux/7fyvISzfZuve+x
7buhdQ163paG4heUqe9LYnPX/gperLu3xNDLAJbLOFXUwlmiLG5giMUpz3qEhdPif7jA0htwMqC6
TzknLX6u/v6WIe4HlObm78x1PmnuoBhV9mkt7LEpi77x/SPFOw46WSiH5Qlp4rZXnm8en973nvth
/eUDOkHadhuZbe9J7YIPes2IxvMRtQux6kzTTBh01rz66yTCYI1P/yoX57XrXwnb5MnJFEq5lVaD
mGZPIphikWLxo0gWcqeuHTUgD55iw0z8R99Jep1+nJ/osERvIaHanyBluVZfEXVIeWX0O/p99wP5
v7hzRrhgYqhx0CU8r0POACclMl45goUuP9sh+lmu1vH2eYqmSMhOEpST2v4wofTFfdS4gszSlutu
yzgtMJPY5uKmMfSS6NVxYaVbKhFRK0BiDQF1BTblGtqH6WfoOYIKgieotvccrWMmEVR2GtoiKcGU
Ej/e7bzrnABTylZwCgFUOKMs3WK4zZK2O7m3iieFLJildgXhpPnYJtJealy6+lkP5lbVpTpWs/GU
lpYZmW5AJxVKzyp/Z6IN38px6v0PpP5pFy7LflALcMJbkH1grl+tqSA2cOwubYRD1giNS1bgaRpF
2bwTluRIxb2F2Rmm/HjnsAzn6zB+gqInltWufyL+DBy3EHy62AUyIRT5mPZbg4APu7iyI4AaqVr5
Q2xwgKoBOOtMCZkW23wDRyLxubaAiiQCMAMgXHxBIVdabByAgmVqrBdPzbxHk4nF6oz0akM+ZeWq
mcRG24Fo/J+5TBT+Ta9KEKRJO0S0K0OIW0IohyylVpg4VcNymse2Z9+xxNYZ9hBi6pzH58GdZ1oH
P9SKhkNMpIT/U3P9WTdueKvO0BcibsuszGdjPIwj8hs0EUIWKAE8ndGq2+nuLwEnggSs00Ubr2km
NEHQk6MRlfIvJF31IpqsBMFhFm4RDqS308wU0Z71C86tediBulYfuLtzwdijkOTuI+VeX4Nyiq2h
7LxACGK5cArr7vnDzSJ0xusJKcw+b1QOVGgFmHmjH5H3piVgJvPeHTjoXQZtoQxw1J/32IaIz4mB
TGf46bNgk0cIgBVEK05hYmQNxjc37flKchLRgNFYbMsM8B5kFghx58NngMsVxN1ddXLTovmbtpXR
Dt1ZmKDhhgmHJzkdiBuFtQICgKP84j10WKnhTMlFheuAuSRbjVTVPmj2TqaeX2QLsgL36n3QwKVQ
+hQ0zHGR4yonkKtexbgxLa5ktE7yQk3kRbHSbBfFTajN+pWcTQe27aYiM/81Ctcsf9ZHmzuJxqqS
HC8CZHtfsukJaKRWBCylBYpNgOd6DDot1vxcGC6HM89/ogRhlEKAdC+UW1irIH984hx+VAFpklRR
5T8Ul/jDnEJoFyuIpQ0745jsxSO/H2w2JmWr4Q9yZD7vQBAuJCes0ECMX1VaztEcu32NZjqzgnmC
yQvh78wND12xzL0gHnuQSH32+/ECzUmeuxVN5Xqpr4zNPbbrRaQAr2iCeAC2Uzaxm4Qfbw+Ut2A5
ppPHGnugabZeMT3eP/MMit71gdOfzYWLCF0n2dHLysbA/LK6zhnmZPYTqGqcWFqh4NBSYuzcgiE5
Vfjv5wHB2ufWYwUhhuBRd8UjXtkArG8ZEzvddTGQJlmEqmDemtT9gWYEfQq1E/Eh97sd7GlmDHww
mqe1Y2LMiPt0cQZA6SXa1AqnHOpMIjN5+kOU6pQuAkwAZRQc9bSfvB+nNjxf8iiHtDceJPZhlKsP
X4f81gACOPiu1QeACc1tT1d738jlnfRrtMl+cfYn4Or3KYfX4hfJgUolGtJeWxIikh0b5x1TmkaK
6HecOzKNfBc2xeCF/NtU28aCVIkdXNXl5fyeNEfPTGWfahuRGKg5ML7MuL3cNWOlkUCtbSY1UOoD
tOOnLDRQHcEgRUZ1hmOfI4XI/e+mrE0m01pG8pKfrFEh8a1fR/goPhU5ocjHIp6E/zCx6eZ9pm2d
RKJg/wCBsD16gKWAVZBgWLjKYGpfqSFGj1XKKh9PpfN+EaQfG/EmNNjybfK2OGniUGkBMGuGAwji
W2WliB6zRp3NDL1FEHN/Q7AWxiwDlomNz+JowcE8PTB4TZWIb+TBOZvlvQ8Mxg2z2UZfdnqKXV51
1m9sri790G56U+Ai2IMk/vw8OwC2vstwIHJbn23H9kTu/cW6+btKc//fLQ4RuDAk7mmlVfzZ+our
h7d89f/UaX24KQzQraaVEKUoKfil5k/dCEQ/REaRJNPpoOAoccE7w66pVRDg4puaE07LnlnqTgOl
YDE+03fleyNmYHrvy95LSM9cnLttLOI7HklarEtDzZ5ZIiFH18eDsoKpcvFxHF/nVEBiR97i0Me6
EIzZFhn1Vky0rJUL8hvhuNnzycF3kT0E1J+1O+Q4VTcdSFNIA7CVknbKdmGstDczNmHO4W8nHSIa
gwr2zpiYf9Y2DxQr9KvDuCSvZLsMYA0//6F3N0To0TrvUycq3wb+e4FctUTaZmOdgwoN+r/4Hh4S
99JXNKRcgn8P0Apyp7lKQKCEieICq+1OGV6YEEFz8fhUE5phelkE/V1Rxd7s4Bd/ESXcGFy1pu2k
21ZRWkHmy6Iqj+pRUOIVU/aHlYx1X9LwmW5Om1LWdne4aEeg4k/rdUfy30EBLa/qi8/pjECRQIXS
lByGmwHri9qfefpYZVcT7w3kn9CIJ+gtK36BNy/TKwO1OsDOU6PGDnfgjs6A2xZslJv4FRtI1qQD
ukYE5tbMtDZPcSdL01NEWv5TUOx2g+qsZQd/LeQ73RJJTXQjHbSVU4yrfBXQ3eoQnC49omQIKahi
L5jqtdw0++Kq+RILohNFfQ0BZAyJ5CEpUcf/xWirQyvx7/kdy2MivYHBViPpsU7O/Hy2hNEq9olY
N9U7AUQLKfHEGaAz7eqZ31Xhh6wR9LD0/7oT5nqnmPhaIrfJ786XnE6v+5qCjM1VwQan4byl2YGL
xfDwS8fwGoIqfrkyvBhStP9pYPJaXDNSpqYx4H+9gIkMSTMskbivI8qjC5U0QeOxj2utIu7dtK8S
V6aPJKDMTBhmhC8T+FCoKoh5uNJbJKmFyIdp2KEjprxYFJ9hXsxihRp0iSpqxP0+YDNPoXelULzS
m8Kx06uzqxm1WnyH62D+SDEg58LxFOLRRUX/XgXJ0W2zWrLytVGdrvNiCWdSw1JgXfCphxHd11cc
iZ6PjKEwQNPtota/wx9N4DPpiIpYR5k+Q850jKn1SvyTgYlvVQr7IOAECQI2+EMnbH2ur8pWHSF/
+djE77YwgrQyQQGzLip3a4vazb3ORP/Uvy3gfjn5gyGFwYCftetUfM3Km7wQQLC+2JL1+R/dbK25
/r+icjjEvduQYvyC/neesjelojCokBgWGsYJGym9wZeD06x9XmouV5QNS4quTtywLD+E7dm3C7E3
HKpz4DBRAPzAcitXkMZEmnDQX2mzSvDa98XOojrV08/iPvdbQv2HcYMSb0fpfFKOwnUZJp6GZe7j
Y10D6jZzMTD3rNYyaFAAcSGP85r2YhNrl8PhPA7fAWyBHXs3eDGkuwOHVigyrZmIPW2ZwoStIZQe
JpMfKsuztH7fa4128zLhTldx5tHnf2umIyHrYgw3DjNylP4ZhbAapypOOmttX8CeVPK2YKsY5Va5
tZFPSYOP+ANqFDdSHFAuG3fQeiCOongpCocKILlREz3McrGQs1STsPOchL7Ue3A3PWotYfmsvUCW
x4Lwkcz6+ev/6SudoddPFNNKsh1eoOIczJwxoymI0WBHBbrPEm3/tiRyMYfnJK4E+IXbcx5wqfRD
yA0BzPIYtBGnjK+VYb9i2RtNNuoD5CgE9d4KWX28K96+CVK9aSB3G1uJrXosIX+JrlpLRaJBBt2G
HpA43Z1wRu6VZQ+ivf3g5gOMyBrK6woMK+BHSOVywkjaFWUeux7SuzBoqGHhtG+8dk2LbeWkasWi
bobK+ohSCATcu9iWElrJ9JVydd6TP3H7UqgU/Im7SbA/p9iYz6yggwWzA7Ck5w7nna+rwpMhhgcE
ORNfF253BlQzS2Anqk4ibS7iyKst/g5eK96APqaGvtsQ5Uzf03Ekx3zHCCd4Ia5wxZLGXpU7MeHa
j/KiEQAkT7K3i6FFSNjsytRKUKji5cVuRH7wbkNXv/hbj8ZCN+35tImbWASvx28QZ72YlRJryL/R
yi9TK57k35gxxfV355EIuuiaM7rzQLXYRckUZOz56gd+LtxWJB4P32Am+q/utPtxO2AOGh42RGA5
uJ32IRgP+xMJNYk1z+KCV/uMmw9y17UYPi3KzpV7LQb7/uqjZ0IqIKUR0sVFzGEpOla7C15YcAkK
OcPQnvsLsYeJ0mcEy3fuh8P66AVROp7t3B2oN8Xcu8ArthG4GzNpY8YbluvdLG3ycFhqtzzQMssM
NrUQ7QCzidI9mpHieUGNo8pnw6Omlm/1GjWiLnyA/A7jBrYOxCgseqtjZuIbZYfzCFSRzNl4Or3o
V645U4gjbcJfgP90ncA6IKe0DotRQUFOAGhmxLex1isWK4j6fWRb69xYhr9Un3wCkoebm3CTOeuZ
nzCKsZBRMbzp50FAo7GeI6fcDd6xNt/5jv1RhzVlUaaB82Zz2x1WxPD9YOBenj8IpR3iZsY4OV7h
uLKsLnsRDUrliXS4dsc14NcPA4nwsRzFP0bdXu5zjHKGI8SSY3dv/3+47Ny1aRYYl3NN2dwTl5kI
H9UBCNRBpV05W2LT2zbq630TQDdEdwr+TE8Yjj/V9HFXXBna9Vcx92tDVV1XYXiG2H94jOg8/ZSA
4ciuwBP/Eboe1S1G2a1/s1xM+rtB0b161kV038cx6jcDw3gfv44hwrdoNfMAaMNJ6+2flKdETvin
uA//otMipQvEh8P/+Wc5dUfFNpE2uWvnN0SS5LcOZB4pfLdts1q3bpA5fydx7b+JxgPbrzYznSXT
gttEnDv0cY9ET+TiNJ1ys7bQ0V9Ove2WvKyU4ze/WL7EOYGL76tFJCO92DjChlql9kNrg8sgiuas
b23wz/c1QikTbQiEYyP7XgcnX6ZQef1VQ6MYHo7x1F2dnd3LfNZ3KaJswOSMchQcXlGFYFFsO/74
tFujK0xiO4+SskFxNwUoNoc3JrTJ4SGLunKP4SAsmklGl/aeIgFasfv9ydbgj5/I9/iQuctCkVxe
7nZB/QbWFnuDG64MVTfY5Vso3q2yOyzl6x+rpde2bG95rjFeG6oOg0us/KsHs7eQV0anCXQf4sS4
7NzrKOxrVg32RT9rnwPlQNyHuUEmo084HjpJJYr8S/gJ5sNmt/beeuuLPHM1K+BE7dsDM/8xuxYQ
sFwzgZzRsw8uYi3pRuJV774pFfQdYIwdDMEnUyeacRJqgietSHSULT+2zJNjEWBlPIpLw/RbO5nB
zB5c1vYW6NB/mANaiXPAPSsH1888WBWwK9BEZ+VNIuU+7yWyP4iqBiCUfJ45/Sm5xbLkEIdRTcPm
8JZxyD94OdwZGu7eInbHHPBkhQ0rIPxtbcy1tUTsdUR/n91Ya1whJj8Xzel+ghFBB12rEc8SdG32
yBrZjFhuPAt4XCMykk0h56xmxFgyrTTg6Z5XQWjZZAMfu9P8KvmZv9QnbQZZgTNMeK0Xbw5snq4F
ALBSqdyGbsb4oOlDL9xInh6fQVEowgZHq/CmEl2Sq0+jyPx82xWKMtVw/i1WdQYiP/NzA8EPnQzw
9fjEj1+Ne6SiMSb2wUScjbdQ6rMYeDCs8YvTfa1FLKdQ87VCskjBcQ0TIF0DeNlCduEwjlUPjFMt
ZMgjy0vE9Q/adDdaaB9vfPxjY69WOIHQ8YiUNgAdDp3M21DkJdzFKRKx7KaC0j8E8Oo+4Pi7OWwo
WbKSNrE1hMUqjEt2FzwqiBL/i7VG+TKa8/weBA+SxqkgbcqV4S4Ak7/DOtcU5qz8z878YsD2wN5K
M32L54NtNpIQYgNdzAGmmHoAOtg+8ug1SWCaRI9wKIC27odxaqtDkfDNLuZE1Q/hirHg03IkdYKn
R0b9SD1V7Jwvaj4+iKSzz1H0Hrqxj6waz0nB9OoMMDYEivUJaB3jInUsfsRT7+Qgnkh+Vwjvf7Sn
jRX5xmqk4kyv9uWglnBAgE7yOr69IeQ1SzRuQRlL7alYjWbJUVIKTdriCO7QadcYT/S4yuMOHmTh
EkoLw6JpSSF1DZnrJRx3/29eV7znCuUhCI9hQdxL2cx4uMH8ND9F7EDMzLhgMZF73r/E5gY4+n0X
WA6/0hQsmQ7fkmgGU1JaSWmSgWL4nxqH+8myfDH+lGFDT9Hqcx3DfJk/Yy9SD0Eocm5cBRiP8J/Q
wkmUqh1J+95CB3saCfIE94GE9GSy6nGdIwaCHj61zxZUu4mkipvuTf1wcTAamEYa4owroOjzbIDC
trV68Gj4FPSO92qXaBD5wRVGo1+PklvI2eLirRkiDRg0lPS0qamZNlL/n64NY/rIgzGaR66Q/eWn
1rHDt4/j7NlRR0sdtlku4PTYQr2+In4dbagjW5bOupYXsuVvoAG819l5ZO6zZWKFhxlCulzYpROy
w2W95s7fVt0llneKRts8wBouMbUzjp6HSG7n5v/7EO2gyzmLvJib0btLxOgGxklq30cf2mPVzkdZ
mKzDbYNDC8yOz/TuDvcY8lk/YlgbmJX5nNCUUc2zsh6OwzqD+BFXAZavJFjybhC9OtY34MAqnsgH
9o2hL0uvP+LP2ZAzg91AMp7w8irTO+Chh+vcCVD2IT2C5q9c+FNxPNuaQfV532R2XcyEYvXjkuAh
5DF+sdbUB5Q6DM0FrN1c4ldIerqILihAIt5CVym6TSTtGsycOZNoCjsd9ehAfbW+AA/HL1h78QX6
7Q+/iuVnIuf9T2VnvXF9hYMyh988eb7UxFWQtBTbamLJl/KwzSFAKsJCkrfaF9m3P/EhiZLVPox7
UN+HNkqL3etQQYwDCLOqqRN0x4aXCwTx1FWxMd9Ma/IrMuXsWLt786aVx5q1/XLj7uHRcpuCEyDE
un7reS2GiUxXeGnnpzxscsEeYi1chKLupgER4lm9jPYP8A3RwEhlttg1FejDYBDbHR1DSecWURs/
GdIo+LsI+TkE7nDQS0cV3pA2rNc+qKzmCeVJGZ7eXDNTpkIHbzCDQagm8IAmFEyf01YXgfE3uMLD
SGuDGYbMZUD7gDfcNPGJYM+sKS1g3zLjWEGvE9SW9IzQa8RAzUqT9bReiA/wabenz6vWawGGekt6
oqFy0XX2sm0GHYKn7iEPeDE4NlPFGC7m7EcTX1w8okrXKuXKEPcKzULJfl4rU3IdaMpfERv4/ike
9kEZAWbw6QCxOcmaXczFVxIG0oTnyp73xsvp9aO2py8IerpTS9NUlqtMYXZZld5v1gJ0D8dJzvDn
l6kbqFs6t+ZbFipgeNAKV5G969X04SQC+Rsz5dzFlM6VtjhhXcPUlmKOyX8UUQZxaSCj7UALQUXH
86Tc6StkyLE6rbEFYomrnx/dRdnAeaLtOK2+RXRLiOVQsD3+5eavyba//u8UYio89lX8DFcc8/Tt
OPM7DlzvSO7kb65Fu4bwZYzdm7+eMeXCBNGFordNxXB9ev/++FGcyyU5gnjBExlvgfJAAQKL0bNd
ricM3gC52EgpDytNaFMDIXmYmKFhS80Oaf4ho4bTC5pR+5jtvQylRWiM5nmYqIxo9gM31VKcMQmO
EfznTexYY0ObZuXTn3IehSeJ2pxIyPj1c2ppBdWpGBuR4idf+b7OFip0D4x6EfMtj1QpcpCkaQvX
OpLXOScYS3RD6NzfE0ZrXHA2vvz5RHhWG3YgQfRSUnpgSWpf9Ieu1xL1I6VjYyd1GG2phqxf0VVu
jO4D9qHd61KJyaBr+lxy4pEphw8PjcNmznKC0phqVcJBwXa9XJ5/Yw/wsAk8G/9BtH1Fw/PfhmDQ
3vfCFSzzH1O4xeYqbxDAdoQL4vKK5Fvqdoy1HtsnUygWB9WAjIkK5DeonG9CsIkgNklKpFylNcm/
XYQHcBZugrCI/H28qcdFJNat5+aRhfcozvqR8xBuq9sIMgxoDje9Ns1cEXBkPYbs/lonQsfOkzCd
iUaiH/qhNupTos8QFZdQGNRo/ggM/0IVZMlLTJzHm5yow4dm0q+PO7A1BBvvBUeKJJ3kxiJDAALa
3SLLrnrxmF17Hjb8KzpcGFf3aaY4c9E3gOAHtQ/fkDLsxucCGxyMDp+Pxxt1GIGm+jlQzWMdVHec
aITajtxkkMyaIWlP3AftZr6tk2ZB4NbwsyJqQiMfwR83qiSUzZmze1OfyARnLENYT2jxgrwHToS6
WN8OZFDtEDv4j4anxGLIqmM29qgwvVixbfVO38fvsGUsMJ2NFHeAtEZ5zA6gcCSgeHUGrJuVohB6
sp3kPmtVPmzAGjajZ/cjaOjIacanzOqF6iBaOFfGIGfGM5JEpiwHrJUog/2ED+SrlUkcQC4BVH/y
nVZK5N1fwW3nGIr0pR1/umjWQy+7z+rvlf6fBgY8AIMcgb+jaCkLttErjtGyTfNFtnStHgAJHXtE
K06xg03VRVGhZJbPOPmxePbeLsd4hA8p+byPKSgtheqIATYlIFb/BVpIR4tHSvGNWc+MHx2Q3Yvz
OpNZZkiNkgSWHRKoH6O7mqiTo3T5Kxa7ahB6pjdfQ7pxunswIh/M8DMohyb9wmjTJHyoCdNRGKzi
hcVQX6kvFKNWAq3SH1yacjn9CbbDbeG3/Ue28qTNF2sFtxCCLp+2LHsEwGzNvkfLIJ43JWDXJX4M
GyTwYj/YtJw5kkNtOCqN/xh4vny4ZNApN4LUKWMYATX5JCt+sXQvoZrZbSLedTuHPBj9Q67wx99I
rIGqSXuFhfLljrUgMxDV7GXXZmrCbiAGNsbXiTCtl9L7WT2VN9uRZsxL+plmCXceb6Y1tNA7VPCI
YjF352Yjn/Wk4pEaQ4iGx2QXU/394IuOlpia6VTFCVDw3064OV8NYkPUsSAg3UqXKWuFdfw/dbSd
U6wgaEtwTammdukOlqZ4+plgo6mkVVqv3IoPW1M+qkn73oQZy2K4qGsCKPcslZXesGz8Io4HXzNp
k2toUJejPangQP7uO5W3vtjty7jwv5klp/w8u4eqSQyDTVT25Lt+bv/W/u/YLJrQpawgJh+XsCyc
+7M6tr5iVOfi2OCilq+g5p6zGbCwrusfH6yc9C5F24+Kq3IaQ6WS/zUcEOrmWXgCf2JviOb6U8i5
VJ2yOq5Mmt8yevqJl0k6z6dxt8LoCnszcC6UE7uCbafLrxb8+S2r7aFAetI0L8mVBFYa8dfM/3rB
bOcBVY6nmwpXWk7856DkfnjCPezAO85mKDrjdjTmyYjW8eWuCnS30ZtCoeuZQLg2oxw1/h+Cv47D
AvL/ezQKZ88s+vwdgmJT9fj3rb9CI78RDJR629wD1GjGQ3I4M+zE2lkY58sZScgUDo3BZX11Yyo0
3vx78CjoV5jO14S4ZRSjOwBhi+nWorO3bve/KVqFBAXjRJVGnqeWlc8oeLPhTTNAravVy01J/ZG9
eWePFwZOx21CK3ObTXgLqYIWLV1t8yBXaqywOwFhUet7nBhmVLT6tSyVqSBvSjMLI0jwmM5FF1HC
yWUqWxVtLZjRWFN7jLo63NkyJR1Kz2kCe7njp88evdefkZReIp9qCgPbykEBNvEJOBbRMc2iatag
aG9OWwqnBJn6fXi7PKYoUT8m3KA23HsEjWTtS1LDUa+QL7p9Fpk6KzQTxdw1EUT8+Hh0Vme6PO5K
G9yfZzekxxK+m4wQDbzMiqVlQs+k9tRDJWq1eJmhOaXlXYGFdo9aF3wde9fheHf9SzfXoWpZNNlc
epPNcCfG9kTtCY7+INv0sY2oVdIYfMiz/GogOiqYud+6z2vyfkiNcvlYtXZBFoGZ5Kj9YtjZj937
Vx13XwNbIa8f7kTfCVkLOiYh9vWwYKtYsm1JruDC2q7GIfAXEpSY7f4m0T9jccx9UgDvoM0Vg4Ks
H6oeijl/omqZ5ZjXiejqgW4giMyTQoSdIAGIWw/K/FLC7Gmii98sPZtUAOoYx/OYpC5Yn/ef0anR
2Zc1bXgob7sQr4T2PkjPN4v4p66wwPGd9UTS3b9P+TUAvdg2tW0MZ0iIECy2dYXU1YnBj2CkzWnl
ZC8+lmOPG2a3qbL6hTxn0aVVqqBJCerYaUCnAWjPGob9VhbsuCIq8qLi7wQHfR2WYAWPijVhKeS/
NGOe6cScgFzgu9FuDOhZCqeMuQaguxj0LXfwsCILQ1Yldk5yBZZKjadKxYyJ0/1aEgul4UtRZT2b
p8xVKrW6+C2HYpgg7q1pdJeIi0S6D1dWdHHYT1tDrue1HqB9R2rtwv3ZPOtIGdB1CdIJdznki1gB
VgnjEUKgAH77xhpziV+L5IwyjRtlAtqnEJIVSRucl4dpLMctiYXrh8A0FXZadKA1uPHqP6C+zlKO
j6WGMO3yI//tQGSem6Kz1S2lYhfoivsXpbCgTo/qOQppbijvLYsr/y/Lo0r6jLs6G7pV6cWvc1Wo
X4A+VgpsWYAiMai3sKXfN0c1kUSd+glJ0wLZUlIPHC2BQ4j43qsBHtvRVe7WLtHyG2x50a6j8mAq
5iq3djf96tnyDTuGhLyu3vXH5iwhbV86o6RmQYzR8BpSTLmOQHqji5E3BE6cObJ8U9WuWT79lBfn
Hxdf/HJwZqte9tE/YbWEyAk+qUktMewMV7gxzMqUW6FbReO1GXK9iQ4Z5w/8EP1H97MthxxAgy4K
m7zqRZw42xfMjfSdAHRPaem4XgdW68gMNi7b04zUKMEUgRpGuwOtL4h4rmeLagVzZYXcHRm42GT5
8qHQ0A5AfOLUJBg3rIrv4BhdyV5lp4yp0o8ylT9yePohx0dHQNLlj0hL/t0Y8x0Mmovh0csE1Z1z
zWkyYIrykMZ3iiQzxyzaI2MusUkzTJz52n8A5QrZMLWCFFzRYLOecB/96omfVVdpdiwsLnn66Ios
1XmuwyAZyPn89FBRBNCV4ugFmyTOm3YCwPZUp5ZnmEC0eSNEVJYWZJvXtdC6W+/s6OlE+BCqfhCX
Ea8W3NOYhGb0Z0vBwVVC5gBwRZ46oCUa3/HSOiq0Yy9717P11my/daMnIaH8slhgRMqe8boUXYvS
TBuLwr7gFqHMmSmGc7sf6B+AUBn08EasIri1wF5wGeH+CduUwNrcBrgDmwI8Ta/4wm8GhN19KW3P
208jCaPgVoKL5sLHrq7XIXebr/PCxerGyT1p4WMcUcShrjDqNBsHdyHELta5hJZ+sA8Fvou7m46k
ySOopg36t5MKt/AWd7lAFXS+LaIHxkaoCelz18saRfSOlR4+M2z/mP1QKq9ssB7DjS7bGCaioIRs
/eDj+LA+DZfPIB2+u8S3Qqx/ALWNF3Ob35dvxQQPEwQVpxmiazK2TH05vdY6OwwI4aEYBjsgCYbt
xUvKTMky5YDMiRCIzcwiqZQD5xyafDPyuEhtw4RqDyc3Ar2wQGuHlEEGoRBdiJqFVF8oh6VOa56E
WGBU67jwzu4SfwbU+OQTdDdXk/XM3ACeQy1TUiAqv6+0EtX7e11x+fGCsgCtj2oCvMecCBadFiWN
HkxAebugrLZVkSex16Fo4/PwyEeUx5QAqgsBV/XMVdgpLtxA8mtx/+p+Hp/momjNJSk2HCVZnW9O
4Zq0VSLFPWj5QQEVxtNbVdTHB47GQzemSPLPfEt0OxYwCqSKdTTuORouJNNyPAmJNalexfpdlIG8
ULGzHyjTSr0cAuKqkoi12f9ECwaYddz9ErgAsEBE7faLy5C1aTtbqQaiNeDQxREAosQOt6RdTizq
wyX3bSLqQIDHUC7uvXp415WIoqVJW5bxgJTC07dzdc6Bc+dAJXzW7yH+p3gEOe/EHk19gwMxc+fj
1sB17F6ecDY7l1cMCNIktZfqO3+czOrRFU2SYYEmsQZAXM9lk9g6zvQdd74EkCKlC46G1nYZh2cZ
DjIdvdcFwfz/z8iSoo0I/vF1u/9nTJ95oi7BC7PQ6pV/rtu6jcpK8WXQNNmTaPiUhpxeYP2Q4mT5
F/seM3N+I8rAoUcPsvtFLaMdGN+/G3gBU9t4TmxxWUvYsZzj+Rp43WhbXpjIxHrQ9+KA2uAOa9vF
+ySQuxcostWbeCLTTo5bFxF018F7Q1RYNtmErcEhzohH5In2I2S3vq6H0aVZny4m/yMFMYf4WVVG
sQ0JB1QpqvTxojaOD+TRTicPfmaREKfD/N1z47/qzMVNouM3YtI+AsROyYTK36JSOVohCI+zU/8s
LPvp+A39tRDytvGhCwDtTGc/FKNnl7kFqx71Lj094AEWmKnqlVv4u7Cw511JvLDtjCgQ8fUijMdV
TDxZMvHEm3itlRAexQX4cuCgjf/StH233oIPKUIBP468C+WAMp3Z3PMh91pH5+Qq5dyLAZd4rb03
npkSu8UtGD2Bz2h1+K1g/YFgY4eo258t9MhZxoro5KAy5NOuc7x1bpeSPo5NzH4TixqpEH5ETr7J
fH9larmwTIXkOFog9qfZZfHu8jjv3RDeLoxIkUtZVk54hhh6mw37yc18dcKkiaBljcag/OFypvHy
ktTFbCRsfaWBEXHqLDb2ne+OriIjMddhvakbg1CjU8QcSvl89LipA8qkp/rtkgbV6C6VjXcxnrlC
p+8YU5WUNUE3GiTkRZIUE4i92OMKOsVo+UpMLMH3SZ/dvgWlQ70F3fEgDbnBeRumzoQEiwf3lcOp
6FNz8n/QfpRt6HvYbng2ZrfA1s309ORQ71rywO7oxP58eKangrWPtJPztGv/899ORRhuyIP42IXb
F4e+904AJnBrtYTVNu/iWg/uy4+1POUGfNbN3/bye6l/sP9KVMUlkq+JUwxffqwJRg4wTULi4OWj
Px8+UN0mSIqovBbPKl0Yastls66Xe7EBqx7HDBiF0Yzh3Xs6aki++UoNcLfQqH2BCUlGO8V6xc7R
HxusB/xSiaP+NiZWNGMAgkqZFpVWGzh54OOIcWbffeYe/CJ2FGI3HQ0cwV1uh3uhVo7f2mkm1qeh
nrn0lWwSwdSqQi6nfuj4ovvd0+5nB5jZ1nMgYWKAudcwIlpFIj+N+34WxfecjTPy88WrOs3d2e51
BChqZOysHROZd+mP3SP8c34aCwZxhAnutE/rF+mrpjoTt0AljduMo5mzhvCGfmiyljNaeIQfLrhA
Ye20ehMK5H4DrWRhqYfgXskvgQzA84p4quVRK9Z/SMGzX4RSTUmCUxZVw8TO8ZmdTUlvoNvgX/5F
GWyE1GJRjiaPfv9r7Vq0GJ4hVOvieKTkMDlFT0r+QvrmC7p9w5U9zVvi4xypiPuYIGnFTS7ZGTYs
tGJigYV7lam3ET6t+RhgCoJHucqRMwYcoJP12Cfu1XV/gqgkJ+Cc5PI89BtPYniZVsNQQn0NAsPD
IBafDzNUFoNRt95Ifit5nR2fjsoS2VF8+YiP90F7jPifLZInPFODNChe/lvKqRdHsyDp+Mlti44i
ANDiKsjNI/Qydm4hO3rKb4Md9LnkyBrkJ4YsJIgINpSdql4gceQs5OgQ2cOkNBXvbP/s5WL2UX4h
ZtCZTRwadJfYEPxSd+oklWmaocv4edwK8TwjUNecLh0So5MqjFrTDIKnSE1CRh1o6vZNbrTs16Ls
nVEpN4ILq8k5dhr8K1Mmf2ZGrPcZ/uDeHbK9XVGVgEKIeJsu7NW2lRsDGXqm8mvFDichvEd9G0sw
FzXIGCvGTAN31LifHK8RWpRNxJvnp4IibiFYVCbVADOPPzZzOq/ga9le6ZET/7xQzKG6HDCNn1KI
+cBeDvoEqDkfiwfrW4Gb/vgEDCdTF+yExRhZaK1XInW3nlTr8sDXes6xVW0zWl+xI8eoOi0C+pkL
wYaLJvV+mRvQpznoAn1AngguxJPocJm3EyQGR5mY/IUit0QDaK/q26sCggmjny2jWnUcGZVp2syL
OR0oPWkoQFjqB7U8s7ghNZTlIK1l5X7bwMQHopbkCuAhSomOZh0e4FfYvwfg5hx5HxolSqBocsQb
zMDTxVo+VRecnN2MsUd6Ju+MZRfz3LKFVg+t2eF3vrshT8R5pqjjqL/xcZsNBlczAqOwTgopOHk2
2F0W06ahvxq46txpQMm29oqnHoBBUuUdYXblHByoy055VpGpx/4bml/0UGKO2Y8Ccx8p5EeigJhI
hOh7sQv8VFeuKqDR/Cwats+gC7eEo/y51gdNzbZrarJo4C/JCl19WL3lVaIgy07B8TZqHhkcV8wm
8XNiveziacSGlzpbuRRjkyVi66oopZHg5zLIOUQHtfWzawzqzCAVvwIYYDvRdr7RhTHQnsIr2tZt
/DmvBkML4ic1k152lLAOn1fczcRWddD62c3X8fE5wC+ParzyfnYCcnTCJeXi5CM2oLewNsYUB1xH
hsvs8VQDEgVlmoMi/bWPvOtphEz3e37K9QOC84SQ3ZSrIuzAxClPzmJb32Iqu8iINSVgjOwyX1VH
32HU4T0U5rwjyF1rv5DxJekOQMAoPkIaU7n0HbA3uZVSk5KyG8z8/gFGoNjD6RlraEUVv6b/FGfY
TOwM1TUPIenCYgEWr9imKUjGtN0UF4Hhigd4F0Q0XBaO2r/HTLPr0MP/C1/jVeop1hVe4dU4udBh
XSVwaXx6LCVEQ/cLKwTnNnHQZiG8al9vxM89OSNXpcHEohAaG1XuDlr+aGXeF+3AYjs2QlMPDLrK
ZoPsLX8BiNQvzU3Z/KLGuxV+nw7UGZwrnrDXc5cjwYL7QZKDnEP8zOXzddu39fW0qJosDgrpSjqb
4ACm8LX/dC5Mtn82X6HE4oUApEIQ0Caz+/oLb0j9knXRoX5+1bwZxuxws3RaLIfED9sY+SwqjCb5
emQER7ftOH7/ZZxIKxwo41GX3Vh2TcVDccdz8Ywu9u5nRZ3H5Q3+nFSj5GoU6T1Dx+rOWTIfUmhI
5HPzQ/rK/XoKfOKRWaYZL+5f9zSkpP2kNmQeeETXFUirb/NYe1Oh+R8koiFaZJGea3lDrRPKaG6e
OMU2+uzrKu1VWmUjFk9gvF000I+9DxMjxt0+jfEbNhRvx39oZZ3XZixsgDJMMesA2ZUhonmfzInA
AA64bF6IKgdY3pK5snubYrlVe+wjemNlKOQTMNq42VP9eESV1H7bSbV2OpHaa2D+rtgzje+ql0kx
qQ2jWbQCRVQlbh+Fv2UkxI9BayBWYSVsl+bBaoygooRZigfiuMsiZr/KmEvwTCN9poqRdmtONWI0
sxdgVGoWAvRuebpY0H72n40UX2tfQbjCZoUWnW8k4Wbwg7T74Z9UriShAyzFnjNfr791vVywxYdo
8zegFH1J4qQsSK2ogGMXsCEaygY9aTDEE/ZXYDD1H83QHQoqSU9XEfGHFpXn//5pOv82TmCc0KoN
q6jrjZZk6WHgElHNtm44CB4Ca4B/EdxcCKvf8aCg4oo0UwrpMpbBAF+x1nl9pglftUE1IO4mlPMO
t4+m1xVsBZUIc+aZvsPbyakqsoDCu+ZV+dI/zTEEehGP5LRJ8pAEhb/xBprEZ5moiecWpIC9tXCX
JsqtIokW7gExoqay96qnSlqTgEhDOgODm/LeTBjlC4BENNqeUY+vyJcRQBxw4/bopNYQCJljirKn
ancVaV6vPcHpU5TzSeXwhzVkoDdv2+WAH0pA4hOKq8EPTL+5QI7wfcXuM0WCc2uR3qgWh+IzOF7Z
6n0ldEYFwLc3QPvzQIew17QRnNVJbpbznumkiLRZkgNE8C7eE6HEffWo6mO1OyjLiPuJ4mGJOXrw
6Xuh5g9Y4yr0I12eG9cBmasiZ8T2MEYP62xNJrWyuG9VAMzWYj5luJKWazjasoPv212Gd4+PecFq
QtiWnfwtVNC9+aSPBoZyLeaRsc4luFUVxO10J5BcZ5Fmu/BhKpt3u9YDZaN4UbWksUTPHEhiMIFV
c+WZiVW1Zz4kUTXIqcHAZUFnIVRzfc8y9NGpcMfFsSJgyjjbjODZGky8Luu3rUcT3eSkQFSWrzBB
jUsbVKXiH3CmmcnsCbQyCd1QL2eA7ni3JLJPcgNpRvqQ/A1KqehsDxndN0LKwiQc7xYyZRxAPXIL
kcZg2lTOpn3+4c7ehfvU6FrJ4ZkcXbj6F/DR9nRTx32kd488oknWu6SYRQx+DvLF8LCME/Lu4xeW
a5aASBKcuU7QOa6BSKJ8oM0dAbrQFCAVTL8AjS8CC78Dvqdb94mUMPQYOjWKSeTajVcLs1GMud/n
VNNccm3QIkToUnNvM5rMctKeUZIHbXjbIeOCl2+n+E0QgoMqER8FOJQhP5sagc/6Co0XMqGbltMS
zaHjf9zBcOSs57k79JlTc2cOiCbHVvep/L0yvMsLqChql6jESPBJVmKwHLS65vFY6GIgoZV9zwrM
K4wtxmEfiyY/OM4EgZ4AnXA1rpvmNvUo/fyidEx90C4y3W1olg6teq8BKec+d6/kBmHfx7rgrYrX
gxRiWFxNSSS7Sjy8BDLQ7JF+bzG3hLiul80eaN1j+W72cmiPPRsXNrrH7szchTmXz+7VJgjT8AFV
A+QG3j2KfbzKMTpyE7/O4WGrVE3glAqOn7mlJoqaGnxZGKFOYx1XWnST5Zz7jZVMjJXRooxUQ1Lb
8SWonfJ/H1NVUP5nXSpvV2q7gykdRO9Vl1nAafkkk6kdhuLssp4jCaPkMWdXYrnud09jNJ4SwzOp
ZQyCP4grGq04Rs0INC+ORMYSSjOZ0H6TE7THZrHclRaCwyf6UIxoJ0AIp+WmSl8obIRUgl09rqdk
EiM0a3V9gEcuBkVT4bV25a5YjR+nP2fefJ2J9gOo9S7MdfUn3+xjH3uQfo017rX6jLtq0bbT55MA
vwdw9UD/USWoLevP5LrqQc8cZPKQQcp/4Gb/tvnrIovHNzZA9Pyz5yk9PZV1zXUHXK2bjLlLBQ57
nGfuYutWY8sJd1ATE6pOh1rGmV8sg3QFqBMffuZ2vj5FSTe5DYfVhTQxrIhUvnya4oiclAdR1JeS
Y0hpake6Fpex3poPAdIaFHzDkQgK643xVEKxXbxk26Ay/h/qOqBk38s922xHcujIItb6HyAT+IYZ
kGEGCzPd+ty+hArGiHzmtM2bJbqBQlUSP9i4zm7/tMkzrN2g18lky2fdSmfCAXs9EeAWkdYNm+es
+0381EjItGJgAlcQoXUJNpsypu/lzUzVfrV4flK0aGq1Qc59727xQn2kLCpuWph3yyEBiLyLoXYM
bg/3Liwp7ZvVg3GiEygXF2BA5DBZpyfqdRp00fIgxUqSAU2swno6wAxzGFUrocOhMi2EOUNCE5WQ
s0HagxtAw7UYe1OF8YTimuwwkO04adnWhVvcJ1ameuHxzU8kIpTCBzH+DEjanjrtEUDxqHSsvP22
fr8zn+V/+Baqh4vsfbjMIPOu43fvM5ZLXa5CjImugXSLIpj+znqjeEmketpOmSgV5vaO6NzUlfeM
4zaESM2w9cLfUvEGOUBX7IKDOZe4TokgNl/UJ4bZlFG+G55xnkTAZ3Y1AXzuLWLOsn1pe/U6rw12
IRkV8/sFLhJVtpFiBvYv+Y4sx5SDjZH1feSsb9lRz/3wXxA4nS+R3X3/rnO0PV0QF/Yfg10TqnP0
fSbpEkpwZJyQYmjTwNr3o1dc1inbuI6FvHS6FBimr9oR9ihKrfxS/yvzKw4dYlCmSjPkUukUrg5X
JrKEwRpUZYCeO5WBJ0OJUaEXZIKWnbvC1djdxabRcKMY5jgz88+HCTulXY+jh9iA0cfRh/Wt2X8Z
5jIbOP1WvgiZPL7HBEt+2HApFmTbWNoPAilXUf4NZcn+7gcWK/AznSS5trtt79aN7zs8Juj2qIx4
QtUfD6YRIyF36ecWssI5O+Z4j5c0xsbQth4UwZm+gOdTc2t0p9qsFhNsjh1AI2BRag3K2ujOxc1C
YYQuViGWq+aPpcxxinb8TMUqwPxHh43sBWrPaDnjoTutwNE815wdE61x0gLwnGuVuGULcWXg4RqE
1tnnRSLyFdds/RKh/XKC5GpoP/AqD9zqR0t7aS8FPff3qoNjmm3eYP+QxcWpMfy4a72IJHKY1ygW
+zo/ZgAvqJvfc/DnH5lZ784YjpXfRO55BKl3irvaws4SGKkgUYTxMZGiUIuftycWwfPF11UxKzPL
hUPSy7ZCiZbxICx/5S092DVrnTNeNMrbi+TbzJ1Jl5kN1Q/aWQOGmq+7RgPQHAySGdVB/QLCd6QU
W8akZ75zuyLFMIxHAl9MsJkDLeXlNjhCOBB+vAZhpfd6o3y0GvzxI4W/lYGwbagTNrPLvZ4pibc8
R88SLIuqKXTXRs9W4SHgpgF/RpXOObEx4SPH6ZG9aLIIoha02KR6XlgTxeeZCLH0e3ZTnFwe/dpK
/+H04X2ULu0gasmvczLajCAthhmeF0+fzG9Yyx6KHMV7j1HV+O/mQ4CPy0kItjujl+PgKbGsZ3Z9
tmW9e2vukxYGNBmv6tc/9JHttftZ8yhT3JcJZtnEQJY567frqVK+ZHPRV2qhJDy/o9qfNLiOksxt
FqOt3i7DvwPkRvTnfk3ltTzQTbU6VgG5wcuL3pvaHAFExedBNLtKZL5aG1MEoa1psj4LPwNigFTC
biLnEsCtkZ+FKy3KkFz1U14Cc+f1/4+5FIy/TYzHnL7Y/CExVQ/ovwF1kTOWYnf+omTGXzq/G247
qHUQm2MoeUQlXNCmCEqRq7Y3uQwMURlr1balYMUT0ccy6slulNmBhvX5T13wNvhZsi76L4CEPhfk
pAwMipciiSVoNfiOrP9vUBrvk0jR7sut6dXuRPdzBNaLFiQCqSVymd1E2Vu4SYRU8LKFkPCqJ+GU
z68x6mF23BuLlUZFCRkFtvwHTapgMZo4O2MIzMayp8IU8GsSDquU2XHnJK8gaa0l72pFayOrOboa
D1xFYtnmpEJDEP+TsYekrUkGFlzP3SS5FZdC6LFS39iH/qxPIGuioWxxGaZaJOGURe6FqmxV3AaA
TUTl1mJyJEguuLOrZ+jzqs502EEvwMpCc/szoYpiTi6qptBeEvjChSYAGBbdHR807vuESceQzEsW
TNNnFiQob0WxkktsXt9Qj5mg3+XnvHaidyR0djYJpUPS06FeON/jhk7+hTUCQsjFLgdw2XUBcFPB
/+YwnPzOpYaZ15VIa+pH5tApnodGXVG9dAAoPNPGnGuR2ZrNBBvCw93+O66FKz9+6rNjeVY1ilMF
B0HkxxkzYC8NRxvTxERd+SqzfHX8n1wv6eKygMMet7dzxJXN3TQn9SykncFbCr4cT2etY/sbUppj
FVKlAS+Omuj5OYgPFkV/FlPQAE/jP+cE6do8BSorgWIGKPsEYXjcpjLcjRrnBQNFq2FH0e3yqHYL
+rgZCEvu058zMQ6IssNBt/t9/PK0wdtLgx1dzEPhDYVBxmiYhI1BnV1e4hhAN8RM/rfKMxCZBKW/
0Mfzyv3a11WZmwkQZK8UYUBhsY149r516mxpl0beEXPCkjwWntLmN/xfQrClAwyhRpxwoXoa7l1Q
hNsdPbc8kl3dCh4ZsjTr4vAxEFX1sp29Bm7AZOZh5hMPem6xtTQD7ZccgXLvZtPS2XdiAo+COarP
+DJhhePeSKgi9vurYtqB7S9f5H7Sq3dY7rx+G/R89M8rulaJh26pZST5OrkcKFtDmdLWcaJi9SSc
RlRv2EW5zO5k9ewXFj57aoWg92sWARwZ9xM3XGgK5GVHa4OAn+kBHmiWbwSTEzbq2d76GXbcTIbQ
XeyeOQ4HfWuYpj+DSWKSdlh2iqrjaGSyPbH96MlSx1GtRgfOyHawMhKrF2MBff7yCM4LfOmi68XJ
3hrs8jBS8BZIH68+decJa7b3Bh2B7a3ajaze8O0aHbDhImNZGcBloEUs5io5Ql57X7ILP5nm+DCD
VlAfYqaW5N6OofiypPBuJzhoFS4gF8OKk9nL7h8qgOiljWOyscnDIxAhkBNpf5mNbcWl98w37KKo
XWm1ML0EKlDxDPrhRzhdHdpoVO+h0+6xuqSsSbVaaQAFJ+f7cXULqxCgPJ9wN7e6TrV97D1alsdP
6u2Xi1lG2Ns/WTBKc2T5iHRJnWYhzTGEYEj93qTHENIFZ1gLGNhsTvCEhY2Kavfb9X/E5LON9xAM
tDsBUrHCrDZIUAqof50sNIatJ9kjGjvcaqNvNmzm1DmKS11aRTgFdGhWmynJGU3t6ENfEQnIpQ9I
CXmecuP/LRlpXO2TDYdQ/Ag6uIQqDGl1mrgL59+jw97x5k7l5jRQd6RQjsA2/KPXtiQrLm7jA7dm
tzTya1X/JMeErsrm6sE9MG3lCaXKnxF8JwYEVOmP3vULlqTCwV16Qif/1+gpvN+fHWs94ZDnr0vr
da35KZP5QiqpAR8B87VX/mP73WhPMxx9qZxibVVgWJSY6AtInzHcoeyKx9Cf05YLOsfirJ9fdvxO
chW0lENtEu6DpNvEYZ2Q4dZnTusZqqypY3Oy87rRM67ytr0WBogSseH345IRcagvV5iZMnD7M8qV
uPOCwxvUduBp8mGFNdTxC6+y6/WMcQMGRc5BGWRYp5QBcLra2KFZ6Hs9RRqrS5FVu0Hh5JJwjBMs
z7Eg50t3/RLJmJ1DxPfGDZizHuISakBQbEFOO0IkmrFlHc6P1IfeCNZiRN1skPtLjMa1qRrJVUe9
/0YfZzOfgLydWRiX/z0HC8k7A+dt3mGMWVLLx/FzFDJQjdAleFw8pMLU5wUDaxOUsrBBxyC/abug
CLGcafXWKvdYkPlkMW6CZwiUXWIwfYGJoypNcuuYdrJ8THLo4ic/ey48uRhVwbeCCL16wL5GiZF4
Q/BSeqQ5hzQ1k4eYEr/Ir7VVwxN8RDjH5RRsxsylCp0kfKy6NfHKvO2G1wSFduB51GgRMygdk4yc
UoC5aic6ikFS1yczBeT0VYylencnRKkVWM8WqGmn511OUM4qLz+N5ZA1pDgVEXeig22yHphCfwka
mfoCIoA88d2jMBbGG3RFv4Du29WSURJaFt4x6wFg6rahTEU3IzAQKZpD98FfVR2EN0x1//pBmnmt
RTykf2sFclBuQ2dQZ532vYj/e2vTm0gUVAQmx960ORnibs9ruIF86hEo2RAj9Q0x/sAtmP/TmGHT
4lykTcc7OHpYFR2ZPDpXedBsn2HgBIebpwKJi1dDGNxrJ8vdrsrVGFLsfHZIHTD6un/tdVWxLDxZ
hmm5ZZ2i+KEP58hmZbt/HmLFT0oqnUBf6zE9sYAGUFf7nEWPKS047TOuCQjMKS396p6ikziRvaAH
1w7hylLQF3RUkRLe3zAwss7fIgEbqbiP7Yz38s7jUcpZDxc0w2xlcS5sBX8BVIi0hxp4oS9QOZv4
lnIypGGq0NBt2V0tQ+FP4GgTCYld+gcfmu0FSuqa1vF7+bnyonJPxarZFKYJT+X7HF8m9sJmqhMJ
M2qE2j/khKeldSBhnuxqZF2ulVPWkkrTuFwPAhPVUiYnypcQgu2m53/DhjMzmdPhC/FoRrWKy5kb
dK4/24b3AN22apcevZiaek3u5lySFZrepy/W5ciN1ZqneresYoc2ux7geRixLVA1iJwoSA17LuWl
cvxiPjfJge7iPg7OwNB8X/uLXTxUbiwWOJjZkIY6NlRxvK4GNl116BxQpNbF3SyV1OuK+mKwrZg+
nnTIlVlcLLbe+Cz1IpNo47YBNeKP/rRgw/CBlt7Y194x78Qrqto0zWand+8OSG0zJPbwV5WOw4RK
YGp0ceRvfdH0CgWAriYtdce4FoDv7ha7NDUVsiEoRTgqaM1hov/UD8iVuhD2WQAC/pj2pS91KmqN
1xt+0ZMjrdB+It5vD3iVaab3C1aEePMwvILrfyfBC278bDei+Xyx69HjFFDJD7alinYkA4ne+Fk8
wwpPibU60mQN1acfePyAm6AnhJMICmwaOrovzBckfjHCV6joi6/9rHrJDL1VwLj3yOXv8NUAWbOW
7Oh0+rcpcAz5424xUF1lEqv2+5pnN/1iA5sC6LV4j53jldcyAhq53OWFPJzHLmCwbYinX+vs7OAH
hehkleQdIqQqncQRDgY3KuxwbvLkcRL/kM88ta5AhtpolMMm4RrnE/HP0epHYKeLzGpiwg1ZRyfE
4fHB1DCWpMptxb6RChI08ANrhXTojPqnX3PO/2u98tLjnxUeCkqs9lbWjxIJR+21vILCjz2oSl9P
2RsB18fDnsRGVQs36wlvlPzUsbww285CBdF+HVFbhFRQlI0XE0VaE3XxsOSORVxe2zlNwIdYLN8P
TaxhgcCg2JsyVUNUXEewq0oUran5hkmqkP5sbNUtZEo1/G9WQKZ6C1d8284/L17fkeYEoaTOLoEv
BB+vl7EfaBNLutQJ0nt6IECHJ1giinSm//4WiPkznz/9qZGDcCWZgdoqwZR0OlsZgGPezE7k1b7b
zlDWZtpamMN6vbK61zZfXOTXeoYZCMvQ1Z2rrpDQUnkykVgwsO6LyCvcDy15BLMKqZsuB6DjUEs1
D2JYTTzEXpKoDiJ3gqaodZNTRNVOzSsj4f2xK0yU62+mXBJCkHBzvq0dxeXFitx/LS3QKmVZYRWe
G+fXOMaZUHsWt4eFAcuLAyEF5pGjzvIlW3u64oTl2P119ompx4XJWnQ+lgXe54K1Pq0TmF8LeWdF
JW8LmBsnDfeuxJHp7KNZxIOOkD/b5UlXzC27esMz2xYcxdE1NQsaElGTFcjZgnaaOAb5EIGL/9h5
tluyNVnbqYxwnZCjeJ1DyjzNkm07CUcyRqznV04C4b8isd4QXskky2kX13CJqVDUTxFSO7CGxHG8
2KxH/4/xnqBER2NWa6cYFZ/H2dYNKrQJh1e3SNHI6H2PmH2QbOMvcyChTP5CTlv3M5HzwjWUUWAx
XH4qc7W8l+Aru8EuSi1xd46SkW/cLS+3IjzcrMCuWooaU5T9aj/kY15SQOM7nZAcq8ZkqsUm3HVi
JCzCICU6hqZryIMFUEJLe4ymvPx+12Drg0CGo6N/tfjGQvSuqD3CIC7k2PD5LZ0UcPOsyu4xI/Xx
reZ4+8npr37ALTgqxvKMB0mbTfrHRIlDPMGVRGW1zPIMPgmhmZVHft+US5p+JTmNnte9tKc/Ven/
WF054Xwb5ySssp2PhAKKcMw+vqqC2ww5dLxSdFo7dqHOQd6rCBunFKETZPzhIsYSdu+WRGi1/cVV
rVInvJlKh3PhQ9eAKu4f16WuepLXw6i6dLtY9uybIOE5Bxzb6zY24Z8t0saOmVYz/cfSn1+kJQ9H
f35DakcvcBfGZIzY0nNyA3NqZORDmqhHG0soAhaayC2hD+c9GyDePL43ljoJO0pWnJXNfO4GFUzt
kLcSwW96anyG9pnAI/KToZkkCMrnCVJKCPKx6+JXj2qhARbSCjssgWkl874JZCJ6knNVAuw1Q9gj
EX8vMqFKBSmQVeko8GrTy2D7GXPLlGrG+yk6hbPbaDsPYWn9Tr4RYhsd70PpkdEMthngkthJpxIC
N4DTvAVSAFYofw9d4BKm/QnwZqIUrSGSBP9CPVPKIuMw5qgtZ7NZESoqvuhEl5M8ogV4J+3ljFYd
sv6L21KrYvg5zne/rvGRgZBjrsv+pm52/5kqasDP5beeLB6LaMlzacH/ZebWD7pDb0SmZpXmsGpd
mZJ++k4obiRDeUA/bWVNtCtqPJT1+4ugfjm+SzoY2wl0zfULS0gJKkGvlgt2s0kOYmBgkN9TlJqA
2JAJ9q4dVmCkwVAfAgIufJVbOUeEh5dxHu/AWmR1hgZneRJwI2vhiEd1HySdaLhL2mn9Ral4c+YG
Qqw8H2PMiEr1JZQkkPpsaaYap2Ihg5M6EDKIC+ZWZfCWTBpCPu4YWE1Y7A+CoR/ljiwdGzuRriFv
fbCALfPjQDK4hCHkfRKVo0hpFSxIoZ4Ko1d7JDEByk5QL3jIplbl1i2nVw3X1uR1tewVySt9iPKT
IPuR1Rz6hRfIg6DC6oQAItBYK8j7tuLjIZ32c30WhGgDXloJTyQDClVNNTgMxNj/iZgnBU93/BFT
VYXaYXxAeKxrhR3Bbvp6mAImjMKO0eTrEDYasoo4SU3vTZ8dSFWUQ9EFm8gXHcSM7uKeaX1FK4fm
d6lKTWA6yrPANOqwl/y5VZmnppVnCZyUMwLCX5sLAKosJViFMLvXFTrMQq30/UCBohZZRUQBjbe1
d7gAQByxCDXFEQY8nD0iVOG7bPpUkAzZSsomtTJB8wQarZ5bxgZSJIyOMJ+A3Xxn4zKCwnlWBxl0
2iBp4oL60BhNh0aGp3/R+1tHVQpehvnQ7O5FlMxPzHafIUMTDJ8cC78dBA55K9Ihw3A+zQh4gaYS
xmoy674eAgsR/fLkGFHqv9L8dYDk3pBpNiy35inrw7fs9LnZi6zsggB40FPpvoDck1IZiCXhhQWT
d2xDyVk7my5g8LJue5y1hg3HN/kMkQ2To1Mh/8BJJVxOYqZAT452Q+wWVy/17fhN7gvTc+HoMF+i
2+/FVw2G0IBciESd4ksiOp5xRBjICLkHUytDWyFVfN0pUDx6iMD51dZOqfqEt84VihD1jRA8QWB8
7oCUqgW21qGJNTln5UQln+pIL53ErISy53Na0Eb1B11PsYxluTSzFXIc//wylrAjCZA4kaDRf6oL
p6QNsJVnDhntgBD7GFjayuqCKdihJt5I8VHJo+SfGoy1PsYBlngMjqqi7utEprk0GL4ZT2+EPF2l
3NTPy2p2NTHzdQAuVXGVnw25a1XDRTwjTvn0EBw5B7LWyC63v9Gsgqakc5ynaCTwEUimKLytvN+E
MZkIx9kzvT0HwVNO+IUf7NdvVg+n4R9mrb2/cQCRmzO9aNswLZH/Bl5TmFjM12d7oVU59rST86se
818Y+gDMmEF4xsXVlafD4yb0lKfS3d9psIsoLOQZO289c1jqlW1eKHkBprxSPqoVkZ8mI9d7kNse
hEyec9e+QQ9Vc4hybv4m3Cs1UoPgDky7kC1kCV3FOCYYhqV6gmdpi9/HKrSGxz5qMbS7/c5a0hQ1
LYgTEAQPzAc9o+0CG147uMutHPuXBN3b9tenwbRFjT7FxhTXSVWKXtzFIxbFHgZQZ0tiSbljRTz5
zTiierWuQOmmWxUUFAw5sDviV7pTqfbestxn8zv+33XaROi4ZJJPyT1ufqg523A4ueTjmmu1c7Gy
sZBCTx2ZqzJiU+i31Nwb4i0O4ntOHG6lmmQxb+yFqYecxOacgJDpy0i9NFrCn0DBHXLcxQ+kIAhz
LCMH1qUKuoMPIaOt66EFF4b7mKl8ZoxUvaEafCiiu2NQJ6wVnk1w3flAT2SKHprxzvXL+5F6H+p6
7bkXAQjtL3T3gpWPTtmjyIcvXrJ+BodHJw9c7x5z8HNBspnUL+h8uH4r1ApZXfZnNVtAu6UGuLND
0wrUGOH4WoqUb2BRE2W6JvtIU43W70njqxY1ARoKoSLVh2UNtnM/JIM6sTvUKVgzwifqo4QdHmPQ
aYgtoUxDsTgKxUUEcj6JMuUmBzfDVj5zOz48b+tRCJdWo/HcVM3nYNMSA/A4N34drfq25ubMvY2W
ac1Yqz3Ivib2My3/FRJ2RQfZAVLn32rL0JD1HvVIST60S4d71w2WCzBQ5bERuzr4TZaDZ1EzyUFb
iInNpE6/BXWwvOg1X2mOvHjQw86vAn9wxqpdKXu6xflpWEywMpl76QWZ6ftuI27sOO+FCOoi4rjP
SvjS9vNraUHWwHFXkeVMO2mHunHOZ5E1elCwy1o+U4DD1kU/bYHsBUsArhnG9XCWFSTsL8gRn46+
GG64+hXHzDRECaU4WCqK4panS2RiJhYzljshz22Gzu4Lc+Ojfd74pjoPL7xd9S4DHTGJCu/GgzwN
2jfULB4XS6RGXnc5aFncUxjWplpzge/wiJO9W4xTOlBXmtFjIPoSQMiePiTg07rwVdFHbOLGyCUM
w6MoWjwvBSuAzqj/lyLrZtMJ2SdXhaENAMXI8JGiEIBu53/yzQWGIhh/OZFo1se7dN3p6lLtKPaA
7NgG3XkgcdiQY/XE3RG4gGwVcaqYna8TZUmhZ5nDKH31feBeOv1sJx1I5+X9zWFmAmDks582HLFV
w98RRD5sCM1Z1/dqWoXGsO0yvFcuL/ST2+tZtVQygXgq+5r+aiMzIJ+3Hki4MTy5yMcHSrQX66mO
91W7FX2NzpT91z+lZ+RBihpoVByp/GHvY8wAxewPb4tCBJxlUI4VWV1DI56+wW2Lh2kaCILN0+rO
jHYuJuvwTCe6Ide80TjfMQGSwlkizXbTfM8SS/L97fs+fRlm/ryyktncl8lx6NP1exsvPLVYhkpZ
XNg9ehyA/QIREAa90kj5osavKluAZocR5gUe5zYrag1VkA8tClyF7sxmbUjofM5K2a7QrV6JZodv
8m9vJIuPA8gu2WVEOzSik2Nnl1ttCyIMuOH1ML7pE4pgmkJRy/wWIgGQQ2wK5YmloYVP+zmEQTT9
d7QKuzOu6IyWT4EnvS8tqYVv5M2On32TN7Etak6G7jvRdt7j+kETDyjZZf07FrgOTClJZeZ2BKJz
9VDQgGGgwtlAYkv2IEhrkmoPiC1UAoJFa0oy+vliiM0BvtIhJZiOJ+kpyVg2pzLAscN2VTPSXa3N
+b+48drnRMQLjnu100z5rchostG3602BWWPX3lqjX9ifJi/eznxFcrlOUgUwTns06XT9WA1Fc1Qa
7Fhm+8zEddhASS4h2QumpxB2/fpGDqSsg67K6nAC2s5FH6WEWBwwDhqvQzSO5GjFG/+Cddstqkio
3KsHp2tHHaJ9KNRObilsc2/W7svXndbPEZbL45YfBxiC64F1OPuDSrYtpVKcsX7g8loU7bTm5B0K
cfxJsEdSs0fZdMykQZHE38mjywvibYQbEGKgrS0iv/XFirN9nUk7NLmCQdjQLeFh4lRyJQWSdpqO
IgiV92uplnS/rG4/ewzZK6BVfzYZKTIHXoJmb66FIqs2JJHOWNXPrPd48z3di+8+EgmR1jS4b6uw
C/uJdK2xN4loW/rlNbuUp7xAOrNubbeJESsM8HtNQAwbwYyETDLFaH0Ho1V9jUSTA/VyvlPhbmRx
G9SR20nfMsX7iyFfXCw5IgE/SfMgVxQuLJBzgmrcLpH48NtZxmm00G0I7uriKHCOnXdqj6n0/ufv
rfeol9I7DxIcrhhvkndN5N/dbFcpTEeeXF5JHyox8kFW0QIjdTmkpN3PUdjqEkwScKVT8RZPNyWK
dpcnT69pG79M+zfxdt2xxRtuur4GIoVA5jm5jOiihsLsaLxzEdFyASAexi/L95W73mxS+IBrQ7wJ
aZx8ckc64fAl7cauTzgCdqmhvPrqELco3mh1ADyCsmwezrMYD07Sb7vSKPb1mjV28Kj0r2NOMMam
aeO8ntq+7MS3JGSuxWwwWqKukkSamrbvTR/7ECBRFfm685htohmSnMb/xEK+G0iJWOvrRUeAm8UA
502Q1Ix56a9iysjRadVclseDenIcHrLgzGFYQOyNyKcA5aYrDgkwcrQteA5RKXclBPUegangigEc
UwVWdMzptf2+xlsQUz5A62jCz6g90rLP5YeBtfUQQn4SMFz/JJX6PO8XkgF3JZHg2X7p7tProPL3
CKfsDds158DV1muB5pEJtCJEIqi6dFcSkkWS3sae/Mo4aHZ+65BHL5SlxtniqRTii0py88LIG3Ul
L2dfir1PvxNEJQwWtrR4sH+QsNisTxZBkN/i4jG9ls/hEhqoVyuYZIPqlniiuvfhYW6sWq2a0aJm
hzDMrq6XssgeHt2O/VqpHFOzJOShHlB+5n3eC+xm8TagUT0uh1yxpCdy+mzoKWFDbrw10VVP+se0
33Ldh/kCWFIYJIrTj2SfE+vOaJV1LyiiL8tpqCM11KcemQmavHca+lR9/4YaeWwiPgSxAdqIpAEh
22UsWxgopr19Xcc77XB2aEa/l7zljuyjTrVSXzsY9dulBGx9AelIRJ99kyvfCRKxg++VHpEtvMHI
CfcG86Y8XVWi8VV4Ja9GQI8PA857Byufs9TTUwbvl9FqqFbr0qJ7qcCwlA3iGsFkLgMMd7LXtE7h
eEhWlQd94p+45dorDGQJuMBs7W1pyo11lZJbBMiaONSff6uQu36LbK3CPh5WlYJd0+8eWGoeO4Dq
tcwckTHXKK9eHh0COD48GLcGeXX2ZCh5+UmkYZGuXbB6Fbkgzgjtq9CCc10Y6Z/N3YR3V9Fq9G2Q
bvDgofrbuAkF0W+2o7am9AMS+X2yKaTiOMlemQiavhH4vrjcsdhpBrqXxiWKmSXBkNcqXO8oep60
/DW7hhu8DiIsaMIzh2+qDnZOXTtCMpXSPDCTqo7YtiSykX8LqXo4xoQUoMDU9NQczTqrvOE1+wB4
WRr5yxjlvCKAPZoHtAl5E7twHsfV/Y+mJGKXc4XnuKvmvV2pLO/PLFFwjY4BG1n4auGXZzc2QGBH
ifazF0Pz0LNpjTO3qreMT1g6u+KimZp/iGLfr0txvABxTQWTJbCjn3wX7r1XVDMGsBRCq+osUOxh
S0jNDHBKIhWYP/LFDZXr7viWoe9OscjaQulTmqk1IYIsW1HJX2sWOuzVS1COXMsSWj+ZTnXXzCm3
AVtzkIBDkxOHvZYHuAytCiDStO31xgoLG0E+LunDvEs4gFt3oQ55RdaI1Aw9XS1MtucSL5H8mfbT
fESVOfit65H8J9WZdJHzvnXVq0NU1eNvJrgrIczWpJQxJWaLQSEyDPk7qef3XD4005efVU4ib56J
SYtGghCniXQCN3iig1Lszt7k0g6aaza0RA+3rnn4MPUUxUMy3WYlhsP59pZu+lEcbu3287C8vdU7
xbcGaUKH71Ngmve6KoXhKP/BkSFsUcBcEzw7nyjbsLhH7RecH6atoJg3HuyffiPBhATL9vU1MLhW
2ITcpQNYbw7DDuTgFAMneiETT+OhQPZlRDocfyI3aegF42dPLztS5tdRafw/4nfn2i0KXmUFt82u
gZV9orYJCDCCAcSWKEG4QpL5SXXVNLP1/37li+5DGeQZ6LYhyJUal/+tHXOq5iA9H3mLGh0DMrf2
sd5trfisdiqNzrEoW2OkOI0ZxywrfVfXL8W5Ls49UDbcvEk4SjZTIZt7aSes1a0EpLWDzCKBXktK
CQwq7wmQbY17NN5ghM1qDVuyWjgb4spMYQQO4hTDCdpfaHfK9IX/82nwfnEXigW0czyXa/KVi+Uu
szWj6zfKMOuYApVyuI5Tu+7/S8ZJAm0g84N9qaRjJu46ZIL/28iRi9SKsHreY/ri9rIpopqOccbO
4x/VGOGfvvy2CpDlQqOaBcYLNE7tPCdG0sjyoroomlfQOo+XzVTKU9kDSvWKwSbf64u1tROjy2UV
9Bf5iDQbF4knk6rsgkHlL5fc+dZEiRyIAi6QKyjOPcl/U+S2KSca+ly0JDuDb7fPAoN+nlXK00+m
Bzgv3DUMsTyIkfn1QsqsznB++87re3j9r8xjvBahXNoWZFAAsl5vKm0F80hl+iaWP0Vkenz/u09G
mH0d5ksAUM3tXo5kvgpJeP4PW1f420HrexKkRSIwpVpL+QfsSEplhBCuObEevrljTxa+pGxhEdqX
oMtbVxj1hPGHyUSFksWpZns+D2xxV2COzhCIXvn5aZgYqBa9904g93jyimw7OKzI8hr2CoTiXgcH
Toxu/IyJmEM2VEeW09jeIxSG1JjsujDz7lP3jMUTLkbRIM5PtthI1+4EG5KflAfy/Zq+NGw6swtY
HtiwrKuKgL6I1YDg48kaHqkAaJ40R+sf7XVm4sGKB27hbX+uGEYAY9eDdZF8Mctfwe+fPwIcg04n
0o4MVLIblsDXlaI0hsnNlpTxbXXwiu0TBdeE2EXBkxBv4j4efzYtbZZCQaVaswilspCD3ZT5G0jc
ZI4kSlZEvnk2TB++AoHFVPYLucmMbADeRjqGyuOiS2kr0XrMTjmch37OQx9/yP88ccg5Opfnn9YY
6BHtDWtKrOVStXPFm12pyZxW5TLpdtQb4oeBTsXCbJLBA1Gwtec4tVpWipwrBJplwoNuH/Wd6Urf
S/w+/U7FF8f/KahAsdge8TC9tHp46TaBhXsqLYIDtNq1JkKYeLi1OSXiscPgL5eTEs2hrnUBqnyM
ywtT44nh4C8bPL2dfdmmyBIKty5xQ51QxsIX+FfjKvhPyEPb3EckoXT5AQT25Si5qbahfky3Elk3
g4vogQYq9GlOYcduyYwatCmGuPViRG+dKu87xsrYVqk8I6YqfaDOPkKrlSITDb+fBXmbCuC+REAf
tRWnFKtppucY1p6g/Xh+eVUORFDUJH1AejiRs7enhq4qz6RrfZEWZRYrf590I9Rji+nNF7FGX1Jz
n4iW8MwJaMGWsGJxrf7X4DF7MWMEfdj8xGvtyVaDYP4F8ftNDhkWRT/z2ybcWAWLNl4y17vbqYHE
8QsZvqaGsUxW95TiBdzlY97G1CEip6zWnLve8BkoSJCdG7JX274FpQKAOz0UG2M6nsEkWh7hKjTu
FYJGr3AYTgIcyzBdczk/00RvMa7k0eaEVm6af1zKTegzChb77dVCofoQ2GHyHV5JivraeCijbwIb
TOplYtGwyfWght/eDWajVgNel+qR568V/3ArdLkZWndHlRj+N7tflljwcH6FIj6OnW0EkEQq0qS6
9MP0h8PcdughBlx+D7zJ2s0s/ngJLu8vXvNnd5zBS+Fg+hn/KTa6bVUXym2zycRkXF/PKU5D55fB
8PI6CRp84AY89y2CCgLJm6nQUrxuJjeq2urW7pMr7cenWvMojDfbODehbcDNC0rBB/K/QHxl2hzK
CNrPLUGlA84zU+yYh0oHyo2XMhSBPa9z1y/eKGMmnTER/7Cd/Iw+IEs3uEJrpMAkbwtz5L5jH9mG
D4YY07zakrZK6rL792EK22tK+/JhQR1w1jMZlmzFg9x5L9uK327E4KAgSi4SpK1yhYspCxqA7HXr
FO8cUxm3aOr5/Q3xncrGsbai5jYn+muRa9FafIgoeOS6WsEKD79JL5HYqk5inMVcVwkmb8+rEWTA
Mm9KoEbpmqPBZLMXkC3INDlIu0levPVDag8umY846AC8ZJdSjkPbSwwZdXj+eumT7NxeqLSdXmLb
td3tJBuf6SBkrpJBarjfNVAv0+7Cbp5S2PIv8LGfHAVikw4B+is36KFvFqDqII5gSLtUOxRRkkKa
C/kQ5RH7Q41Z5cA1ySiFm2txhs1sACoa/vN8xeqqjCCI25w8VY8YAFO5gih33j3tvnaWV8TxxcWp
At120ARcU+3pYklCQ2hW9lBVQACLqKEAz3DiXd+vBWVGv2+Rs/ihwYkj9JZoMu2NkxMedJVAjYZH
AEXwpWDaEhXuFaXINNe/3vuxgEgwy0o/f9LoMkgRu5fUMD3RitRoKyqC6ZbdlnHyJruRaGv7HGD7
eS1mAidmVi2hidhtkPsMuOi2vDmb8A70hFTJm8inBJacrcKW0wE95ISv9dEX0Cd3xoUWnBdtPtUa
q6XlhCf3WbZ63xyAU9tHhSQwg0R+7ieI98aKj3z6mSqWGc48dhn+6DCN+lpgYAEq26rRNqaBFSCb
etu6Rcs8Qrog/1yymisB7KKhd8NyhYVG/GvJXvMk6/fgXqJFhk3WtJtvDq8S1H+5i2cNxQUUMTJJ
wSPbpIHZOBtAoQxvMOV8Js5Ak+PF6naEDRZhkjO3FuRwJkqocxLW8CYgbT6LIDuLc4vaTG27rNKz
csNrlsv2wACzTzrkr2vONwggVzDYXQnHkx+fpwfwQw0tDBR8+dugYL0Cha3YWZwaNQ0la3hpisBJ
zGhwFhcJurZwxb09/Bs5eK2ywoxW68nmyMua/osgmzRxZJVBJf9hOb4Ic7PV5VPiICiKcYeuFz3G
Un25VaNXeXo1UMY34koRFYWLeNL48fDRXJ1GyRPNlW0gAhXIpw3wA1GmDp1pBQZGDkEtMwyG7pnE
HwbX75l6Biyx2eSp32k9Xt1tt18AOIDnFBw7ld2SI5FcIHcb0HMZzX58xK4XTWhHnX4o1Hmx/5nM
c/Y3xY3mKL/yuvlbNDHPUFEcj+K7b8kzsM/zj068Cm3k037q+/fXtCr+BhX9Gd6lgZl+D4KH/4dc
+XR/moyJv3dMX8aIsV8TFUkHR6bALYjuqFKuube0ljANp0CvvZ+UhkaNnIWIrQi39myTJb8uF/Ck
wxHla9PpsrfT1tt2eQN0pYHWWCYUYV30ncOVLXzBTO9fIQtGoJf7jei6H8rZNJ19WBFdYyML9PFI
id+MEZuQz4y6mblcpNqqYTiys6YcLTt/IWs7jzkwxX+jMK9rSUeqsPWgqKJcQ1rigGeKbZkBWTIC
B2+WVFgCCd6FNgTgPqI6FDQt1gim9Il1OhiBYlLXHKFTWdUQsZmnm+zSv01oovzPl/q8rX7eu0hD
QM4ss5zv97OBiWFWpT3SGH95xf2TqkPw5Zx9WhMp/MZoS+dl46yXzV5dhajNiy94Fm7iL1L55D0I
MJGeTK2Zpj2qDkt0UPcDTBDrZDYdOmgNuz+ghT2O//qEp9+n1/svIi+xN3SAgmZfYGc8Pqiv4XIo
4ZKdckQG0SvokFVv4aAohXUFzO1fxW+1xexlXCkiNHiUOpgYdca94t6GeTjVSK7yNblfUu29ySy4
NEp1CHDIPuaNwfrUS2Zv7BOTVUyu+I/zSXnjZyAWRuUeLsReZaTHw6pSLOHKxG96FzcFamfvx9jD
7FgxHbM8PVWQWaLOS50crEWYfEswoLOjlXnqmySR/sbYamZ5w51msm8qTaXnr51WWsUQpJNi1vbz
rNRLytMEW7AfcRySn1Cd27EeZlIg5ULmxxnKZl/dc9XjdGtnhW1TaKS2t4Th8rUUv/TdTO+fp5Pm
rUG1XOSFiDE3N8j3Zbi0Q7eIYAyoJjiNbcWPerneKSD4g3YfG1pRSA7LkFgc0ta0+umkMekRoX7o
pTUs3u7Bq/VR9q2INn1tfAFS4nB6CZfUB5H9HlitIWC+uZsrfCYT32NTeoMRwH/dZunB72LDQQJ0
L0bPUU3e4ND/Ox4YRG6dAP1HalxHxbQ1jqvEVpxoH+w2JqMjqCQAeN11lWst9s/248PP/kPKuqID
k/cxziJT9UwaIGIVUKC9OqV8jgc3mq2X5lHSZAb/d3UJjL+haWn0mmzQQ+GI/QsMrWkFNjHl/q2g
xE6XSmPvZe5tONMzQFupr6ae1hxOaSFIIh9B1ztmFGAHkIz7Csg9hR3RV5jsy0/bNek340dIASts
mtXj6W4CGdSjqp9Dy/OLLeYsLzE04kAfA7hEoO67cw77SxAPSrEUkU2UL7gXySRPtme3heEAcBxE
wzTBEiu9mnGdxDazkNMpgYtQLkBPwWFWNFNlpII6OXLoU8Oc2eUJ2sHqjiBzEz6wfLpScE5y6I/4
yintLsVfhQKIPey4HswzGf2rvPkIFQdG+v+9CJE0O0xesNKxRtX7v2UxWjV46j3AI3Sfib1kOQp6
rrh6LRqlvnm46j/2i67xY0kByMY7Lpe22ySw39kdpXV+fFizfydrpHhV21aBh63IwDnVphc/9qrC
0FFj39YnWXHA/H+hLI/nKVWqtljpuueJSXecrHVEbaLWN6nSoCvpo8+ILjtDiNvZvZ1I7kzM7JPq
C7neFLqKp3XIhbNczpWwbNDflwK27QK0BGIpgH2+xYS+moko4i1Dez1shcjuZRY6ZAIuTwckqt/z
nDzXBYYyB4/mgUz/BKhfrGH+8MICxb4w6tkX1cN8eXaEvsu9VEh+jtk5E3VAV2OgrVn4NviEVmYS
FDq0z2zVGMgmh9OHuSVt9cvp+DtGCd4MvvWEmlXCNa4CqZZNsZWdjF0uuqnx+RMXXVF4KC9osiN/
CAq5Ct0GP6hN5AvFmho5LaCvO7ws4K18hcOPNO2xI+xugXWT7XQP0KpPIgUp10ZDCQLhyfN5qgS1
svOaAPzBgQI1HQcixSZYUPr7eQ0B2O83CBRsEKE5Jya9ftIjka87HtCo1nCOVXUNKNWmqUNLeqPf
oSY5GvBbmMTmNW/oDt6zw6/uMh3fyLsfczVKXhRrV1+t3AOu9Uzuf6/d2di48vX9ZKPnNL3Ne3Jl
0fBYH6UPXTQygtUE516S0NZvfUrB8AceBv3glld30J94kGEPmXXBWTLU84iTkACR4o3M3e60Q/AI
3O4onSgUx409RJUvxNCTUdnAZHdkBH7K5K22RfWIu+oLQspnUWkOWY2foYWsdbNuL4uySB+Hm4UN
urbvTCSq8CiaFJsanoliQnpJny9Ipa/a79qwmYtOYE9IH0RtRXtIm1jcZOe+1cJ+o0t2VLzjEGq9
1lG05Syk6c85sg/yG3do9H3mn+NJ+XvMqH7exB3vCiZ4dOXFpjm80ihp9PnpjB9mxJOk9hhhPnNI
qy1NiU2XR/IhDCh8ZTpKBd4iSZuvW6YbmRTNkr+K+woU/KuJ8f/7u/NFjh09R5SYcHIObTCje3Qg
9GnzGPZpnB1EbFHdQzIeqjtxjZHiXfD4TMHSB2yqIPjxi7vI5vET8+aY725QCqEIVvPWpzL4gkui
ga7m5yLkmLqO8KbMK8q/wUH8cOuQu/cjSqtKBx7G8UR5XOvBl69qPP6Iuc64oxSiIHT5mrHhQOMF
ZUa0Faojf2CMp1fr4z5GIzq9ecpN5YCFeBigcCBePgp/muufcVaHHBekGh+jitqvcxHaAS1Pkwvx
Qro0TWTQBp4/xknyRQoZ0D5oGSvIUWzGuZra7eNvxOtDkDo8w3em1lz8vGuQFlwEnWLqgOg98TEn
1eOkIUOeDpUQabeiwOnX3t8UbeaDCDrzbS4D2FAkuqcTgLb2DNyR1mKcVTwby5h1zqveCbhJ4epc
f8KV66qEdcxwgDgWdzjQY1DlGtMnv93EDpR1YHJKUr/jHdBiRIWAS9Dv4zg37x5Aa4B7JBmJPFXD
qt2WgSrzrVMntbgYNVrtF/hZa2kkPaSLm3UW0ag/YnsnyonbOQPv1o5ie92Jv0OtpOb8QIt47JiR
/lHDdDKCxixQZgJ9lN7W/XdNAifFyDkKoCcRCNPlz3IDRWfHaVKrlKstT6bFNaAzsmH5VAKCZL99
aPwPw0np4gWsAXQk6MWiSWBTrwPCU+2RtHpyCAM2BMSB6CkT7i9AG1rVeDvQhiu92vTAqjsSvL7Q
sb6n3ZDzUaoA50EHLhwxAncQ3N4KCz6TuxwzPAzz/2219f5yrKoBGnJ8TGF3e71UUjGVKa7rOaqk
WiZtgeaaKq8YPQFUYDGzo5vNkn50G4naHaZ2CfvZREfm5tTkCpZOQK9VIO7QfmZePJbKiFQiBCVv
VZmfs+8HSh9nR2odXERN3kjF2CzNbA016K/xQyarUCtTsBvbkPD2QW790C5tbYlW0mvpoqmSzAiP
vyYnwjmprTNxbf7qbIgnSMLnhaDGHZWFGE9VZs3uULcRy/PU4HJ/bJlvGgXBEH+tx/rz7K8dvBsZ
gPtpVbxEdUR4f8uS/KpYjTjdqRmqzUQTcqyNtiQc8oLiqfPgkMeBzckRby8apd22uZx6b81aEeOe
TZ3XjSTX3kPKsXoOBY3QIoL5MwYn0iiD6SCF5raEkOeOJoE88SYjV7VjxVGTyfG4kbkuYZLgGGNl
VbuZvIyj8Ap5P9GCViJuLBryujChUUAU6OlZ1WOwMuyUppbpQ4kKRZmv5koYOQWbZYE5/aQv45kV
iWzvIJ47TbloBiLKhOtXUv6fj64vVTnUukPdOM2sODXzHmLD3ShmZT/EH6Kh7Hc0Kmup7he8Zn9F
sDaRDdMtaJf135OokhPtMsSpe6u+ujAruQojlnrnvZgmbSO1LO5MwSVhV8dft1YlzoLUE7aMFxTW
ttIyR70rb7hQBgLu5kQSv8DT6h+TOytPAYK1227K3rCRfdJqsLkRKZaeFxnBAsW3YevBBytNUSTi
nvS6Ys9tcOIuDfgkuQQrySuNC45+OaVxwsNeHkOzpttrJFAkHtEJuNFiGqIvqWiOtXE0wBDxzf7P
oaYjvAhfMvgfkNamgQfz+l3PiHxLI4hCLti+pZ8fA5oFmxc7he5uAn0xmaxUa6/75zAoqyZ+ehob
Q1yZObUpIrRY8jnGaQTNsBkLuZrEj5W9kluPed0Mzjz8it66qgZYAKJ9DrHEMX1dsfV5YLYTacMn
w1wQeYeqteGPqzKKYXu7SBDCbv0UXvalQgJNbwMt7K+VBNwQyF7y3hHmv+hETiX1D9c5H0fjpq4c
UT19ho4JgejNLC3B27iy4d3cA3aFzMH9H9ZjhjMV8+g7nmI/5BHQdjbuTsyw35I2y6frOtD6oX1P
HYvyneuHzkpcMvgocCsSHBFo07eD+uNw/eCJjk2nmCk8K5PmUdRmWZJCEgbh3FyCbVd3I6Vzpkas
xqSuU1Ki6/SR1svABRCbaz1yk0zfc1LkomlW8AisO1bPm/V69cjhFjeJlAshz7c+HykulI5doXNS
I6OdMaw2Vi6sTJ1DisXPpOQffq7HBuIzrnpjUJQ4j1mz1V7BGRVp4s288SCzv46gmsLJj02xxO9U
1igvHxE4gokfbilq2YJ+m/k27KO06ZooGcdJT5yDC4EjIHmGRx4OTt8YEVbTxhy/wiqrR4u6myY5
USUZhJtkw8hua0cReinl5E4jcP3diM9y3wfbhTenNmPKZCT98WKkqcoI4zJ2YSXJqHX8jDenMGLT
PU+SI7Ran8jMoK/VPT0u36PnQO0XdXdM6CkCMEskSHokitBhw+oLk9drZbURlxXJfYZWERVoo5yz
tz52GERKNzov6IhBvDUvw+XgPQA3FwZdPV3sIWytiKG/y0stAUp/zha5g5sQq6a+Onrqds+CFyAG
l8nJSmt0rA0GCMe8cUrlK995IgaxZZUaCHVtIxNoZRvV2EhzDQW+LytpB0pMKJTkH0W51VnuUH2G
UxULTDm0ktJnWwujoWVfnahlborj/guvMddpaKGGQzGgSOhXR0Io7nRPUIDuFNfyP9B19oJQ+us+
2hP8vqx3JvdcO1VE4lvHS4ihJBSbVbYkb0OpbflKteldwNoJ3aa5CHcY5f+oegdrZ6iki+RyGRFD
AvT4waPFGR8IMIiymShRXy1OFk3Om6naRcb4HNqBMx2MKFNY0EIXRYrKwaNc9blHvXLAGa5u68kF
ldQ3qwXc9YSAYv0QyH+ixtbEaLsikCizbO6OI1MweuoOBIAPa6DDoKCQ5unPM9yqZdW2I0AkJu94
qtKahB7HXUmNJw5mT0WH1QQF7MxSdEQzJB5usAFvrWPawJX/23P4uLFmtIlPyhp9oPBT+eYxjLcv
zHekSH6ldTyboqlr5/84K7kuZmjmbKz5m3CVjBkyvI0Lg1wKog6R7TN5rtyw8vw735UNwc1zM0gk
WX+Y8WwpvJrUC5dm7LAgDc1lzsqZ8Pg/T1Xro8/XLGe36j0PKGqJB9D5u7rKHqzQFIAH05OYhEuq
JeLeNysoNqvIsfIsZdJz/gUURxr/kDCQUSqyTkyrHYM9/MwO6WfSQrKBhkeP0saeuRfzuCWYxFPR
cZ3HACL1LEPDD87eCwRxt3JnGqrz3GaHtw/YhHPYdcOBjQRwhG+GmJ6L6rF8dcyyBKcab5R8zXCo
qD0bNifDtu070lSKgdgVSBBRg2Uw81G94kUD/wrz3o2s3DoOYeHo7tGT9S4OWxfvXGJpIN55Tx1g
0vpMU6LEdOe2ffkgjYlWz2n3j6DrAGtkkUlz5Y5v2uTGGTyzvuDmbiFGmnVjh09kmQxyUau8uBqG
RRVYSwyAYTq2hsy6jhXqvgLeFufKqU+9G4NdZwFqKYHoDTsjnxMZQ9ukXB9NoKN1RRMqOcWva+tA
HdZj8BHgHAm6d4LEQdodZBBEnefPaLkJsEm8MiZ65RlfwmBj1vyYQg/sE4ho1NfNdfz5ewME3n54
nSizIhT2EC+rvUWvWBHZjHrTfZG6SNv13XGT1+FFEfXUxwWJRzFozjgSs8yoIkm1FMbCm4LovtIS
OU7fpU27yNgQ7oeukDhmwrtzHvVpsJufmFtsclUV2Je3liVLAfR5+M476hAcI5ebHPhFLta1suEq
2L2qithec7yP3Gx5yC3lRHL0BiZGBnvXsUvEmRsIUl8xCKksgpgwuQmmK4paA3C2o3IQcb46xdKv
rhEm51ee2kwTEJtyNMuU5ZKjl3/qC/8jFyxuPlAsn131vnTJM8bA83NNvAhdwlPcJH4YNYWVYkIW
ZX1BWfIZp9odr5ZzqAt8fFKYMI10rOHLQq1iJF/2mJxU8lTIr6LonxGr3PF9x7m4l3B4Pzexlepf
0GAz40MZe7DOjIE8Bw3wmgjG4rnbiLtq83NOIzv1oaFxcrjpabYy+zl2N4YBqjkappT0wIHf6ly4
XwKhhm/12jvI+9Ywunee6nTC7EVDuK9EuC3PD/9aiAuWNynqIW34MehdvqQsQR+PklVj0qOCYJ48
MqPdxrHDfdqRnZxnokzENQ5dQUkeh1aUiCDl+wwnpKX5ZX1PgGVMLuCUinjlmmpj7AgiCBavv7kO
FBaMbtkjQxB3jogcIKy0RqRYLwxyGklZ9xV5m9P/ihPHysFtp2hEhwdcjuGL06svtchcEK5nLMM2
UyVxZyhYcwG4+ClmqRasEPBoBRHHd1+ZcMOPv4BMenvCNH9l6sAh4V1CCzxyamuAQEcupmUXj5YZ
R/eJ+ofpTY9e4kC5wIY/n957glbmIQyUN2yJIklC/VrVIom9k0NGp3L77vKmLYrCPwh9RcUUUv6A
+BLLdJXvrDRhTzHCi2xMeTnei46skb7hSBlmk3k4Tbmz8RB736RqWdJDRNkaIc7ALNt2CkP3LazI
8/jtgWZUGiV6Fj3aK2pfejH0sRvJE9rAxD0Z7i71Al2WFooA9v50VMznZntZJlO5y+TNz0cBiMQE
dpqqBYcz8aLAOkSvtjJ62Gdo3pgI0j9LpdaN36jEc5qzlvI9ZD1hMpyWH+UZrRYj7tjZpg8HN/YM
y6TCjUaCm8XdRU9kjiDiLfVJaxcQapDwFREhl/AnvIKFhC0DTuCmpM4wsLZS2HUmJn/MnHQA5FG+
TRSJowaYgSryvpAoSvKVI/2KV/UjlvbbSF6aI7L1GeqAkYxTgCdb+3QOOfg0ij67aC3iENw5zW54
UL8aEghGUdNVs2oczQPgUo7JlyMM0mBbHiJXGOMzRQFt6/KQpv1Z5KjPetK1NQlbTZMgJLavp6bc
DTw7tM3fHxu45bzsNAmaACeGP8u+/nKRg17vkVI2v5Itnq4Y83ztgMYHz9dJ1gfHW1RgxyenAWok
1wOl/6VTD7Vgs1hP4ct73LHDLvehFegKnC/osWuAGX9tWGNdy6AFQIdhM711yVqdnAISTGE6v1D7
Expb00Ng2v1J/+hSBltA6nwn0RiqJXXglCo88LocMZyM0dqm7bqt2cZON77uRYeMQN9S8ZyMsbOd
4RENVh43UElDzHt+46oZe09xUp2lqyK2zcjUmFcFxoHACDdaUdcXnPhhZf8FIkJ29x1tmtPtyGAY
mLx80OmQYC2U6hHlj3ksBxQieqzqw5m30UFxo0UuuJbWhmHWNDccrN7WCHE8R9HLA/kKEWCpOneO
BXEQ8/xg2Z2gsleBP02B+FF9ONCBo2/pLZuAS1lcIv30bK/ducsfneueX54aekSLyj3JhiQPQYx2
cBTEl6HhChBCLBFuq8QVlsin59qoRvgQRdL7XQ7slEtb3v9HrqKR2ydnXfgOCJQy+4JTFwBmDCtB
Y1M+yAo04EtZiDT9BWUF1gp8xc9ZU/MB6NT3D/nnkl7HMA6QcGJQjhAtfoZdoltZlkpd0g/LXhdh
fFw/HgvIps69dFEyBPoalzQYiMvBd7UtUBKmn9lKFAPnUrvigAXQbqDYh4wEF7FQ4SsqGTzGtH0x
s22PyOfY89zpjAD6Xjmr8jHl36+MKcj9xBAql7jueuv/0Rrs51I0h4TdfwDaY8rdg7rRT4tpFH25
Lb0WerAoQxzim32yhlWCDNkwTzvFkNTux8duRZcyVx7IkN3psGmh/pxVpdx7cpy2X/XTDBNeXAYZ
7LeI9Ankj0g9WzBcfjpNenzZ4x3xjdYflx9IkH0RaZBdX8YY5Opt0+tuxCZ16ok2Cg7xfFEHErAP
q9kH5bqloSfAF1L7eZpDUmcq5YtR4+C2ElyHZKwsI2rFl3LjKbBGkVRiB2Z9GroE9kWlsYdt2qoG
jYh4XJiM5TMEmBo8xEouIzD5nv3aaaf8zskklnLLg6NgYDwZIVArd1ZTrqCQoyao1EhMF7QMjISC
p6JIl0jEB375NPWmoRLPuEyDPNWnVj2Rv3t/nA4ZfHxbK630hIfpv3zA8SXTv/Nu4gBy83EoTweg
IgximWngw7WTz/lj/meW3xkWTZqRs+kPM11XWHbzTlU4i+aTqZAFK/eycgeo8NOgH9W6GFOE1Erq
yT8cvRlUzbczKHDupTfNOr77aiU961o7Z3rf1W0wVInVDvEpf0bTJPUMU2VvYes8dhfmPVD1e+4y
pxtHWE8EM03JPv7CBe9M0h04Y0nGe2h3CvgYoyB6mQiiSihEhzRd60VdXZ/dxFA5D9hXCubofX0b
hoUexIsMVI8C7W/rsc0YYSZvtZ2EaI6ibidt+yzthAU/NdaTrKabJqu2y5b5b9ufqBifid/17ZkK
yTstg+pIboH/tdzqTxf2kevNGuTmPa4oaOePRZDMacN+nhZA4X6XMdmDJjjvDJWHct4xFefxl0Od
lCLbrqWHs4rmgGa9b8hiadcfO7NkflTUBpGqpJicGepWD0aAKmkru2TFojeh0mPksiBT1TrDxRLg
1Msp4v49bB5OwCWL+c2OVMPbtsjrzX99Y/kEC7fHBGnROeifua5xfhdNpbtNTvozkw/nDT7orgfF
O/rPo67OdG1PleOf642s0YUahZpcdBPPHGWMo4i6k91NRb+/icmAFYcRK9DqA2IxhEwF0q+echW7
j9v5dT8CCJ3znJNpFiGx8mM6sN5cjTwx5EtgAMF9BEjhsUmSlP/I/YfMrPsfF19XksqUXX44Cn+Z
Z4fVrgfF0qSDHX/9iT5+J08Gbw0K3N7qxLWKWG8FGrKxunn0DMtjyNJy01MjevXHfN7XOgiyHPQd
Ka0/YwGbEoyfRdigi9RgrZ60+M/oyy2qmxI3Otr9xwzgFFsNU/k+ljzbd65j3Al5wKHhRUAb7qFX
eDa6OcIkJfNr32wSpATOaREx1C+pSN5ohaOFfDLf0JDzGsFHYAPbAKkOmICXqb2IimFZwOmXgN6R
2zp6ue4NGbQ2JHMC4MvTNpd850nRb45EENgtSo8TPu8tI/aoHpoTLiLyjynzpIG4PTJYC+v7c/OD
+r+3irUHx3NeyW4atn3AwT3nnGiZ7GfqLpnqKR9NK6243lPlXH7zHwIQXxAhzNowQ/qLNsBZYiSp
PxI4/h+pU2UMtmj4H/MS5gZp+DJWXhIOHWmZb5HybxxJf3VyhBos8gUYNdPKM3IaIfutTerjx9TV
5Pm6IeCxJZA5TQTHfFNICasLKanIfxmi4o2in5XjIvgIDDKrvqZNuoNN19dGQxgAymMqrribFP2o
Y/Fnm193P1AX5mA0AKhp1bbDMBufnk9xx7s6NPV/gO/hpIjd6BibPJBI19nZaw3gjr62/fGm6ZfW
8IhzkTR2SZqLSQb4UHyoSqTKnQ0mihJ+XBGEcLzOt70DvHBIwPlxhBWSahTn3EYV7JysYJAmMVon
zqW+cPOOT54WKE+/E6z5o5dMcS6zOuwu7GQMvaxVPt1DL7i3cvPCyYcW/AAr+7Hpr6k9uBDoX2s+
AT1TJVzWPR2VIu4KYNA4hdQpd2mC3IcM1bnv1Ylfk7ypLIEDwczR55jKeL1Blr8ps4rlQtX8OZiL
4ET3y7JrL5kZc6iqa+5FNtfHTakLQB2rf+gU+s5vq6a5+19cGhF3N32/kUPTJ8dwKdjZSftJt8xS
Z7B+XFYNjrG5jG+CfVSKNJY5gGi9CPw+mjiF6kpeTPv63Er38h+VOLCyXbBAus62UPYrmRIOnSIJ
S6xGn8YTGYVJRgMPqjYrXaQ07rbScsTcHZuX9L5hTpaJAMVy6SV1zljs1SebS2JT4J9SmSvR/DSC
LIz5huskxShauyVcErkx10RM2DFv9W6K1PmCYNdctVXizsQb3ZSU+uG/MkzqRpUxYlW4F7rNZ8yc
GLrA3yDO2CSd7/RyScgW2SPPTlv46vQrx1RSt/S80ouBQkvaZ8c9ACp2aT00noE5TOHiOmH+N7ge
OUsK2VW3PxCB9dgNBi6UDrnpBlaBfhPat4aJsCsVx9ImXtgC92Rei1wOnvvj5E1EfUHJlmY1RZ5k
uMThR8XJjLhofXy0vO8nuI6C2h2mDe/buCmtulaKQSssO/jMatj23vrrnznSEuJGiKwP7UGCPfcx
/35arZQG4PSGTwT51xYilSbBScxLmDzGzdHqV5XmKsYpi26oPQQCEIDG5qzb4eWx3R5NJogRbBVy
2fpGZTuYS70vdKFXo6/vwtgo2RqoXeQM0Gx6w+FFmXCOntbBFRElgVp1SHT99QRc/1LdcMeYvQuc
nhTlvTTvROUyv6PvG1vB1onoEZRSB9KISmjSUpwS19jiOF39VQw5TOj6NtegdF/1xwfKuJmvpR2O
RTRAG0EAJxafKecuOjrhFjQ1pZetkb969Dm9kHUrwSS3oRRAeWhRKZ7Unl2X+99pr1hWCDwyt4he
425MbioEo3/i9TmnMGTJtDSOYxqhbr9kllPPbSWGgz79Mdl2xmj2Dfw5a0Q9+sRwhnb0GW8diYTb
sHf7gFpPpP68DQMYJHY3hpwp6AHNVu4sSxVG9aIPglEbEd8CP/sjmHtyuZneTx8ntC22R6NH+ELC
TFmwUf9m5E2kPf456k1TSFGBEiBXgcn5P65oHHX1OLJpJttCkQmr47fC/s3wBfiPNmq5Ov8tjfuE
Vv2rjJX2MRLbBf+AB5mXB5/WiJeWC0djp3tZXKruNItpjVZ7WWB01Vr+tHEyR7VkiWXRaxP8e8Fw
AD5Z03YrQbd6F3Ez/vLTZ5y3Sxfztc2UQlenDJ38delk3Z4H2pklcX7zHt8jvb1qXjqlc7xWzBPq
aBSYmQgBzoxMB46Y1ytGV+agvsaT9emhiUvUtMy3n2j1hmGSzuqh7EBrVu3QYaIhgP/+2udY54QJ
ztLRYdrY+4TWA88kI5cSZNp2/Pdv8MXwoSi11n01c23KkiBO1gnh+yym8GERL/3uT4yYQzPyddjK
AblTICmdsfm1f0yV8RIWy4wTQy3zjFUbCPUOUd+Xh7hLZ1e3KxY2/KdzCP5IfyTXwli66BEGAnzz
CeGzLdR8i8vY6x6QTUeRn8ZKhgkJ5n0gEOtsxODQnYfKmdBRURjjProKWZWeOng2cfJC6WIzrwIh
W3FaDNffQSuJBJhvo2SO9vno7gVi0I2I8wHGyzFd+HJEHH8bNV83hWASlQV2YxzFv6s1xxeJv3Fv
/7jM2XeoAxSuyhoP4wuUsTVabZbmAMSItir9wHPttRYgadOZgJFmVyRL60ILO1JybO+SRybRIYca
eMix+wPk6Vlxho76M8wgjrENm7XfJ5dJ6egPrWVr5szryo9d1wSSIZBl84WcdKhA+Pp59MeKdIrv
fzWITdR71oqIvE19E/PAzNyJxypFHDuCtn07vKnoGMjMVBUsLZeb+uf+fr/VZTsnINSzBJgBvupp
IqjTEM/nmBKUQey2PUxGWTelw4o9msmlmh0ZvnrFJjxE/Nuh15IlUjWsk640y8jH2kxXvQoltKP6
XCNU5I+chJqlClo2vubgyA2HJc/g/vYDO5pofJlhFaJXuFBrNJbMQwoJoqaDdSq14JfQpTE3Bs1I
Hw5pNmu+7ZXnYffjVk38mD1r32/uwrdBnQodLqQ48FAJRaMgRqKE/KQkq5GFAoMUqgxVnc+l49P5
uwb5H5Ic1Yl2+jm0B8wViR77EKUZVVbYKWeSDo8pBEXL/POeNgohzSMkWLAYzEIA7HLPKV2h37fj
J6PzUMRpsHi2zFnuQtFSwEzZEN+VqLz4ql5HtSYgPvhejYEABpna5/+xhdC9ObN+nQZzesEKy2QL
krWjgSrm9lTOUFhvGuxmwoWAPcFQjkIDl7PijmXCjWIPir4pAOYxpdhqFmu3Bj0bGSDmTCl5hPbQ
zEQpgW3Ssc+bAj2xC1Cyy0vgiDUzViyBk/d23fnJQl41fvb8R7+RL+xT+/dkqUD9imnoLjq2qJq2
/KBVMsKaekZcwIwutAMQW+WSBgQfkm0Gh91/3v4XRJcLSSv8DdkGMEeIIBUq+JTCmf6NL57JlMcj
ozlW/9Yct5l4qobNyvpu4UGEhG0v8lMqJLdMb7kaHh/aRLYwz7u+HwB5T23CBsz4PeyM+2MYL4DP
ZFZ3Qe7O0lzfJC5F/40a7pevnBjbmH/3W1i9EyGPfwrtqVDiar6qzNyehtqiuUlmNR8ndi884ylX
T4fG8uuN7+Iny+FdJLLWqDcvNLDtgUVPkyZXgSEqc38S4SaHYAULn7FhSPMs0zqDSyMOvJhCOlcP
RCJRkf+lMvGPMK2g6BnpTxhUSYanmKZnH4vxY+ejLF+efGhzfnnChD7qJLhvIYjYtTbpg/6HjTIM
ry/w9A76M+ggTBUgj1GYesqgAOBr1DuWQqnPRhTsGxrDML/C9m/iGeeTJy0jSsAwkqhNpbR0o7bA
ROolY5XmlDqGyk6/2Gt6E9wDteBNZTDxiir99JLOK06MrPlqS2stygkIGnmklOD74KLEnnJEZE35
OprMO2Bqqnyn5s+Bj4CvMOol7XxiSy9npfhfAZVvCvgwHD2lwQYksx0Cne29XPblWbBCJRlHfmW3
0Gz+FFXsPHYcbgouo1Wq6FBHuvpiVdgw9A9nzeQYyadixbBa1y00wANaaKQBmRRTDNZaqiFIf06n
H9+40JWBTxDkQ+O8KGDSAesxxpibiiQ7r9RAJy5KNrV0rq7yEMeY/C/U9JmmXEUcBB9oSwnlTIyN
M//0TOeybx0OtwEG3KL5qSexcOEAOIlJ5gE3ejv8YWsiLro7Or9s2gddoXLEmcm0tHwFAD3slF+g
GTra4X4VZwJxh6Cuzyv426ARpT4tCOj2fJMH21pT30iMqNPu2JKWQkxeJIODOYfAgdIfJdymE9oc
9n2nme5MQAlInuK53QAOJe+HPMRrcWh/qyTKMSAwfGk7OF+J7LaL2cw8UPsS8S81825oCH9VpcYT
a+bTLoJ1gqPcCqOIusrc6pjbeWwFRjzDClKUNtRe1uq+dmjs4Nro8y0AT1r5uKM51XAVZfchnf0x
JGxipKTOekZcYrAyJTrUt2GKH8mo/7uoS1cT9Gil6GNpJU4PJtssLHsEyubbnn1d8Yzx42Behdmr
sDSjrYxOrpZghq2SqKX/g/JB+yNeSzomPYonBTrr5f0HFdxeQ6p+kZCW6tdH3TLQ5LXH0dMdMbXg
yMXdI6S9Zzh98FCI9WaGOc9zP5JK+DgSLJbiH+hDvfF93rDQPo72YuLw35Em/Rv2TRVeheV+cCG9
GY75tTRleQDQKhKG6h2FEWXyo79HvzXRQYhuAGtcOZmyi0oCj1koZ7CEqnpVqNDRaZ60oEHdGKXy
TM8o1Fsz0gETTAToOpYbsRx5b4XH6aFXF2FbNoI7S0vCFHtIGpVlE9xEAYbMNIXz+dqg6FmIuZr9
myFMp0eexj19FTqde7iu8R2r4Qu/2peLnzAlo/vGwvEoIts+r8my2T2HNRJSGQ2cuArFFocBaY5Y
EqXnHgIbbvDNV3ROS14NafAqy6K02wrbAQqZb+W1dueLakE8d+QKGuUt0O3XGlYRKx/PIWremA8u
srWQ5SRLxh/uhPEkt1vd9vVjuPpiIoHxjSVi2NSKqigLcTAClqJ9YvAfS+D4wDqZoEWqcRYf+Q56
ogG7zZQSI11rQ2FSpJh0BxnIBDGje8yc0NQdbXdWjbYwBQz/zwrB9ZNCv7so/djaoantkOOa5R0W
vp4xhuayG+NK3b0dJPPYKNOv8HfYcczGfdb+FvDGD/8SHqn26whbU17sge03dxZSnEhfmAIII8V9
5deRvasssTCFl3LOo2xYOs2i2fviSdee/1CBHUuaQ99QC3MVomXWjyeJUsGj/WU9IsP7bA/QHlrV
5t/SMCJ+ZRTcWp1GXcVJqGtSzcHggZnasFYKxRc+1Lgh1R5nCWpq5/ufDuTajuIPYeymLLfbzW91
DGkN/1yYUc3ya5RZgD7FJjQW7HXHwXLURsNxZY7Dtu6P8pONXGfHpebw1bhZW1yq4diRdMggnO1v
FQ1zSwI374I2s4k0vsHQKLUwAjdJEQOVGN1dkc3zaw+ow+ZUURnRSe1k8tTWXJ3csG3O1gpL7Od1
BvIxOp9U5ZO2h9zpG305JKXsFHdMcqBaUPZMkmILkiuYLrnix1InjAxUziQdwXR7rYPImK66UaHN
2uJqth2ksjbsQNXPX9RWAqR9ZtkcUK3LHtJhofzJsFJacOXzPL9ZuLM/YIEZDWeRb/hnHMO7R9aP
4qGVgg4fI1TgpRDLjY83UzBVGCJGQ4rfuvDtQpcNYs+88NlzmcI84wQEuapbkPydF5ARlbK53gXM
AIcaf+yaAojH7rAZ8MPVR8raAf01rfXoCpUjvUW9A/8qMzZjrRKWJr0Ge/8Jv6hb3UTvbmky1U3A
O/qupSGpa7kQEJUDJbylyhxIdNuXXYZb/615okqzVJLZamYrzhNwuoAFm4dq/3syI05Q1RVYcFXW
sAwjsY1s9aO4dtYhJgbDy6okS14Fv3ro1x6nzRMeIpW0FDCzF+ueB4buAA8GdyhcFOvFMC24lXll
vfuWsARWHHwij7k41FBJi2TIa0fdsAToC4HwhcTsXLvuV4AN7I8wu+cYljrtlwt9ThJAUc6Gftuo
Y56SZegG0TKj5b4uaWpyVj77Atb8xsoC9fjL2U/7XnF7p0A0KGklETfV2laa8zhRUK3rV7fYbDYl
r8U6VI0gjiEcr53wJ8JJRwwIZI5/NrHFN2Ip6tQUr62B08HgHDlTQPRP49giKxuyYEjXKdsjX3Du
AWXu00ygwyPPOGEcpHa0d0bqlTouO4UMr9ShX92y7CQpUBKO0hMbu/x7lRCElZ5pxUVVT2njfpxj
YWw6RtHyu3qsbJT8HXShxl90Yyyop6ZilODaIdhUFjRbRoVtBnUviMnspM0Q7ISewOfdjiJ5pkGG
k8MUx/v56NU7sbfnaUcUvrt75RdqSw8Y39bQj+ZwuACdJZSUjPdEDawK5deJnFkz10Nn2YUKfrNh
QxWaLzO490woJwKjtz808jfVjHMPAf5vthqyc2I8sc4iZ4TvT0ZBiCFFAs2ZUPqqKI3rNDt4IG1C
wraLUcJFWqAAFQqySFFL3YghSap8+8eFesBvM/VQNRML6Ih8APLCPc37oD4XH/L9Yv7wmRSWunOi
IzrkQdmAIcJSkSqBzp4Ih81R5R3guR9X/sZOkRIoZaQbG1XGYpRTnuedbx620ZEh87hkg2DafrKO
auMRLOHk+3DsCOVW7+qllLPke9yYb42RNhlVS8ayzRXXbOB3JVW+/TR1xpfB/0PoYbmL765c5Dea
Acl197gcDArAE5FqWIMcy+rtXF9L7xcyNLhf9UMzT4GLRwOaaIRlpSACoaayu2KiZbv5QPrrWHTx
saAwQkJgv+e3VVfEUJameebD/S1DVtxy7n03qWmpEa7onQRf1gnGkkueC/9YSbCsZyFRw9K+bBsJ
O5uM9UWmwxb+6Au7Rj34JXPyJXPrwBJJaKh3JtKxfxHGF34hmAyiWMmHZq/P2JmO/b299ng+kEbM
Kwf6/RmlRMgZjq/NTYLFtrMOKp3dwlim8o7ZhAChio5Xf0O5DHafiU8jpA8F6xYNtLohzEpCQBGt
TupqKPPY1mLb9RvzEyDlHoPFivnQqCwbA6b9CXxatXgt5D06NBxKFHcBqbuW7qHFvcnfFMUy8WDu
1zPRiSuebehMrDT7TH+D5OzPazuh9iis1UgyVD+T2EcTci+goEtDbtviiwC1RWSfcEQMO6a7kAs9
76C2ZTsT9u5BTmzKSh7WvzB3cqPJCoSh2W0zyPUifLUNBheD0Ay6M307coZbbkoHZPKA9Vi3KxLs
DCH6ByODzxhNZCnFZlpE8kmon4UddNowAnsmSypSHO5SiMH8tzs34hxugA5z1hq2130mEg4WAC8n
VKnEVsn+QhClBBV/63kCL4ZJPnMJBAz0JZ2+sSoDnRyqKUbSPagWrZish1k259T76RFd8U56/PmJ
UhP7M1tHCcmVHorqSPvfNDDOzCmIXOM9wvnhN5c+AOvaBR2CgPnzSCR62BeOUfLb+ac/I+Fc0Axi
oXf/HrOAioex4BiuG0XNmwrDR8QOJrXGgcW8yuUZ/kKFpH9bNVmzZMUhmZgPe3DgMQ0GRlsLdFJz
UGVsUq1R+wGebQnJjIbvY9Lnvo84fkUsvxidL1EGcyW8+wxtJ2n3//taKuzXOr3eWg8yVE3awkOX
q5EFk2CP+ufiQcfbc1jKtBDz7fXqUSj8BRIH1ZXcamj9NEkMsq9IVrDylvgXxjX8C8z9bwUDz0Oc
+m0SETdhwYyIP4sKCRvwjmAvbyg7xF65mJHHhu8Uk/tX12RFgC02elLk1vxHfYVjQLkei1mel/fZ
2DDUWUaKBilcOnlPtyj6o+lvq2w1cuE7hI2Ud0dy371GYQFREwdwnX2JvA+2NLSPhkkaH6WVh9tS
vqYi1Um63XCccAAK4yn4z7kpk2EHzFACUVAVJYOcQB/Edyo0EyPnqOmD2kjUdc0yTxgysjLMvyvp
Y+0MS6F4YYMu4CJ3QXE4saa2qcBJ9EkF9y1LE6JDFhlaZODVv8nSlXN/4F7ui6P7aflqOMHLQLKg
OATl4DEebXTEKfsEhqoYrLMI48BGecF2XmgRcNl/m5EPLtfv7gk2pQqtQCjkI6l/ZUwHKKZ3alY1
wwStTQuxZLEQpXcoHjP4qqWymgjqJgnM3bfJrQhngGnYFMNSJ+yY6+HLcVbhgBRZg50hZuDMHkNb
jg2nxeH+hSFlKPKqdsU6snqsjdfEugD+GZ9KCk+/ycYdycDNuzGUjTHekQkUoTqpn3oGoUsrZIb0
nISHUpzCU1puoYzKo3QIkuVhUsv+8ddTutViBhyZDKO8iU6/OqkvRYqBvIEK0Msv7ckQxNiusNFO
a9nj1fDwSkeNEkhTC1bsjCrm4yhW2oiRDGab+3GxFMoQuuWR4w7V0yswGJCDlyv8plcsX0hbEHnA
y2HnEtNJ1sdrGTI/WZ/3qZLBJWj56KKMZZJZ5umqKRTMwDx0N9n6EQ+V0gTxLDwW6b6nNQkybcLQ
hGiiz55PaKOqKAq5it1kmZVTz2cIYVcWh7nu/5lk0o3bbUa2PIqEaE7bnyyJmGIXZ8V7ryWfPqLw
WSt+yjlJ0NfeHW7Ntsd1zrqncf1CDzu/2mKAdEqsDYauoLNhatsXCT39bNUE7aG4727/e0/q+jaS
K6WrHJiwExBmhyYhOHbmWUxf+pRwdPiE/5y4ByjsFJzYY4yPhxcH0zvOURly0d53/hkwcQbLPi7O
cNaKvHkFyRMdIowLs5eX4V7KZqsxAszNYLn8y4nP7eNzp4riLGFjA09TFe30Ztty4LImvT9+j/7z
H+6svTuMVt2PewcsWjSpDyl7Tf3zTZQKq+FkfBCJvU/rIJJa/15evmeyUIQ/M3TZUjSw0OBae9LV
KyHcyJ2sNIcIxtTknvwJuqbfbVJyKe3RXouOiEISBNMyEAL1RQxWQH2CwSs/3fOWkYeidsH9IKd2
Baq4dooGEOwaZ//H4An9wN6tfZ8DYttVWaZGFdd7MDYgWR1vQldg+tn2bTkKaiK5bE6Ofypmzu2F
lxw9jBVmNU5C5XT8zDW1rPPl9sZwqNXh4z+EYQDo50PF4JYYLnqtMUVwYzPgZVC0j+Objgn3T/O0
LhpjQ4Mw8cdOwAhX4MHzaJ+Re4uaFRcCgLjHnyeNqC5NBKJ4L6GC3f7DmsmWKFUYzOKoObAG3y/g
7lgxBeZUqX+W+AOz4Q0df+0NWQVN4FG/N3khDAXNLY+4Y8BwjVaM5khnhWuRn0eXIsygsg5QLAoM
0BWSNQu44BUibUfl0fNYZsVXwUxWd2jlPGOX7R/9bGPB7ER6SYoUkX6s+qBfZXH0Rqto09Nr3Xuw
J87u/K+eJrIMYLwMjmeDycTbUMVGWdWmiVCHOFOGRlfVIaRDG982PWQZVN4D+sSAHzxcC4kRpqWp
S+xL0lHGEaRGt1A1LQBuXXimSqaBGqR06+7zTRLOynsTA2qjfy3RkNX205DDJtU5w5g6kKuZh6qD
ZlN4Ey7/DXg+uXDzmSgNrWP3+wRUZa52MGbBnIQM84E6t1veF6HTSuPi0mt8MuRmbA0rpAiT2CLU
q3qmeI40VEtTIK9dMzQ8OIXe9kuHJcX+jnCValtEcKZYJNd7CsfIG6yPU5vHOR0ZtYC0Pd06sPya
LBFxCoyLdCvSCI/9S6bQmUNnP3xmAOoyzvw1J5jZTXk/dfmhRFcan//ovr0G39VIohNmHQcDkNfY
6U28GTb0ClZcvUrdQr2iWER+X8x0faWGQrVb4SiRIvf4+CSzTccmkfbnqvm1QRjxgseuFnUGkNF9
41H/d0NNA8ZwDV6HKzLDJ+26HUPcWSGa2EawKtl2oqaIKSciK027NHAMRUkaA1OHfJiwZV2hS7Xs
HjwSsTLN5cBQ8ac45/zGz4dQyrwWZvvKCpbkMK+UUwHvMeegQQMS3vocFUI/pWzSzZOy54/4RZQ9
C1YeYtPkqz2wmdF0DHIuQSL0niB2h8UsDjw/iml+WC8hrEKobw0Khv/WoKZPPcVP54Y6b00L9CI+
+8z68HRT8/qQkiCbPMyPZhDjXy6Mj0vtMEjAxb6+9lc5UbFY+nBDtSCZrClZc1lqED3KeErfZWPR
uz06N2ump5EZhvt3qu92+lz8YRpvKVeVwVPRplyCdA0EWGWLJ2AOvSlrUFK6zu2OMXHngc6hnjT3
tY71YbiUfMtlykPErQlgnvJnks6fncI0zmDKaXRtfrFFI38YVqOUVIfyaBxA9yoqV2tUTGAiEI/f
EiogyHVsB1nA4lI0Jsqto22LVUD1fu+R419r94rYdSZtuoMQkAdR565uUR2M4pD64NdFzPTCQU6T
Z0hSmbE6uqlWNLwTDRJRs/K+ecB9YT+XJ/jAU21/ZdoM3OWykphzcyrx3/T41GJp2JepT91aCI7m
FbytNtINFzYYDU/fbPcs+0FfzL01SdRLtc0jYxCBBWGYziAWBvhZkrkaxbQnBz9dQ+9mVX1OhO96
8KlfkNckLobvprNhaQkWafcV3UvistUy6IpKI4IXbqy5ZBrL6WyWEI/6jAI8ijWwjLJPbtM7Iq20
znvPZijuQDuafWmUttumL1SI4Xe7gF25IllsVCEFCXwkgWFn79iLd6gUlPgCdEbNTVstYmmtJTkR
fuvVryZLJF/10TPm+pZ656PIdnKKKepPxfzf0ZM60wMDTH79SU2zGIwvODCDP7kEFx2uX6UASyU5
9vVJRETYFWByx7Cpgf0nsEzknJpHOEN6IHjIZrdJyR6UP9Q/7/K67KZF1KhxWfR/XCPod5k9b8eE
TW/bG/wUNWRcnqlNq1HCjLPNs2Iyg/cVC0+rg3eTQIWvWCCd8sjJLiS6D47PBR7SwOBQAZtunej+
6ipsubImY+7wS8RMQY0K/xTlRhG/N3uKu3LIMpLAQPG7ywqgb3bDa/Y99/I+zgUQsSUjjvuSGNX9
2V9eLglCXirRbJGhn8GqUCh4+p+h++Mjy4HqhHIJp8jTtyUWQK05UFOrzRWZOq1v1bj0NHih5HKr
AMQMSR7g63/KyGH5c8ruJuJuZUIWQ25Dq9/ZUwjV9cZGt8gc7M5AYQhvQxWgFlA6mmXX9bQLsUlY
h1vQcBGa92CI1T4tXdJAt4c9t2nz4H3b9125v1gHsM8oXsMbPJ8f5YwMtwS/wxdvDYjbrEJMfTOa
dkeSaOd9PeozLUZEEqcVjVOznLXvKYvL0tHvbMz0wESaYtcNgDVeJ0M5v0kIf3NQnFkTeMasFWTI
iO4/ozZff3b+v/9mmq2QSQ5UdxdYjVY0uW028tv04f93GEHH4656WvU+/ELNoEoQOM03U/sCoolO
IgXuem/i+UwXF0cL6GR7IznkR6t7hRM3Bomzlonn+mAhswoND5IwXPXux00cqgSlBqYMrnq5Acq5
OnJIXOQED1KPXFZ0PT0RNDIHRn4PLab5b3h81MsBUWIyZERnL3CQKRG8wO/No5ZHaTkOXGXFGx0Y
yme84sKa2uKRb0Cp9Inlsk35ehnVKNImO7xEgsFj5AFQuKRln+C9anG6DdD1m8nZctD+uHmSD2UP
feOweLXEc8ppy9hPwjIGUVMTzTzRAsawozdm6pzw6EWxRT/4a3H8wtyZ8omi9AMRgOKyero6pZ91
RXOkP6GRC9yk6IXmbA9TEIR/kDOOEYOAsRQ6WHYHJ29tsxQLAvkS4U+7CoRSOzrGOMt92sZMiSW5
elNhii03VqR3kinWpnwHfV7P7MoK21hHu5mkml5HkUawSinib1akxUgEy7aFrsjg4JgbZSR3R6AY
wtkTtI3WwXZguHXQ8r5HgzU4XUfip2ysrUYXjgl+t2aPTYySNr76pXjsaEI1dHsQINGqsiXBx8e7
gbmXJkFfxfkGtCiIG5+94bqBRQ9Q8mtZFePYmVb/+34ac1lhifRnI725xDeZFYCy+tmCHYN0+bVZ
fGvMshp5pk+PPdINa9G/tHJiZXQxNWmuZsiBcmlo6xncXGqoZTWu3HXpwCzwnDrbKmks4DODsPfM
5Bed1O2/LmhtWZt8AuMj8AI+9rpLuzu2emH0eWTVpL6wcJVIxLLXC+nKzkrQwsIvfU9YVogin5rq
rWN9qIdYfemlEM5EmJwdr8ao75ciA89ytcnMCdQMmnEJJidlAiQXdR3DfwEgfmUhmuVcQ8Z17G6Y
6/mpiiIn6oubSRY3C0+esekeWkeWPhM/xdasaxOYMRLYueJwgnWqfTHUm6igsetnKg+fZ15Y9Rh6
kDvnDjOBAhaq0sVAzNAWstgbb6Tut3zTjAJnMTAjPGMI0gi1FkxmQgxlEkj6kCZQUBkg4GvEzblB
VuDwwTOb1wzJbnfzAmoqashtEX1C5gveUNIYDiWl3TCI6QstYflKCQY826PRucjXdpLOoKOWXwSt
C0Ov0IdLD4fpI8ODFc5KWOJo7cWB/u17KUMCIZgWoGJzz3/0VQuEmsQPpfVsqgKzwuofQMeSLKve
BLJthhfIVuMsP0mAxurwe8sj++Iu4WlEMGTvCVOI/2kyr6EEGDnfvWp5Y9lkQQ/hyslajSHlgD5z
mP/If3csIPSgO5UardMjMAdwcrl5h/jggnItrk8Sne0HvNGmepNDrXQvO7S5KbtGtdxj1iS3whCF
/RIMcJv8lf/7MHfGmDqECwRTZ8EkGdRj2icAJzjKU0yKXI2s/f2Dnm0K99awl0mwzwqukNeKcp+d
h0EJmJ845fKBc8kJVIeICdpq+tVuJQr49U50Cwsq3av55AsPd5EBfi/DEFCzaSXy2vJmuJGFZ6OO
ewilenAZMZbz+gosfqMIiq/s5gRehI1YRs7MN54VFW1QaLn7dmm8mBEIy+/DuTZInSmCKyLXW2wD
CTmltX0jYtBIXXKitmlVOEN5FhQlSW72nUEQ0p+lsx7dXaeZekl0U0YfnF90zLU+9yp/26PvVcwU
OwTu99BaRSqwM7HNHaa0+mY/TcEivNAVn2LdrBvuvzQThWxpr5LzR10yERbfLa70R+Rg9CnMDJd9
KhlNI4IzLq66Y2VNgomfEBLZKdBiNJKWf75tiHT7gtkdTt2E02LYdHYrNjUm7KThiSjGvBn+xcNC
dxpsG18w3IJUJHRDqJIR02KJL9MhtMXoCPnYuIWDzD/s1DD5dIB64IOzzrDayodeTQe3t6wp/tJi
4itMLmY1xkA+lMCVH83Wek1jBP4i5cpUC3/Tq5hFlps1cVRXAbYyodG+g5gWGTp0CI8VrgGzT2Zs
NOPyIODSWpocH+3PAVDrmjQ+JM1KAziz+GMHsesBp2oJi/MBi0rWIFtXBF2CBm4uy+jn4srt2voO
g/zSq9z6OeCFOZD1DjR0CcLqUJmq7l8RvlSxD1s50xgf8F3ebPHBNev8vex+0TCYnj1I/jgSL3wQ
E/8Vb+CwoRd/fSN/xoAhUaCoo5izGcOymJGeiJwGhzBTZITsYbXalq3wc8MsRVfUxDklYhr3U+E3
bpcKNmnG4LOHv4yqqWDW1/Mf4TWqPmjlNsFv5flA7x75RjWZBeSusgdqxtZMwgiKxCG+1bpL6lRP
tuliNxdfxCoMrBVBLchO6CB6CUNOIFRHHjosJeiVUOZv7YAMO9gfG4K9wX0zJRmi1lnEN0rtqEvt
Yw8umH4zVqD/xbJdy1aQzeh6WJfg5/Mw2i2IZQBBHQaf2liBVBmT8KLHj6tvJ+aMKEbWp/pXy+fR
bRNTfE+eD7LLEUoAgGs+RipcpFOBzOzSsz3FOH3vwSqrgF4GUs6XfQ+ZwP3qxkXb+hWgj3DDo9di
NMxF5nyVx5nZ9rXsyafPC3ryNruIpRb1fcTxGxS0oJTrJtolSlaNMfs/aRbvtXKRA9f1B6+gK3ya
H+U7mp+Et4TVV8vKPNwFAqHx07VgRaGnPbCLMGRQ0H349iwE3EqvSmSjJjOiiwvraKuYHMdsBL/j
KUk5qaP0zVxdyZwogJKsgM5RNVDnuaWWkFfhO4yYAMvCZ+CX7WpNLS2+yBLXyjuGiwLNqIP15Kzo
S+Yu1HGAw52CdwNVAWZOXeY3XMFj78hBfY+/SiNZAqE35GsZdTwPdKEMMbGT0pwA0Z5vOEDDttaS
Kqu0gnJx4As0A0XGJrEeSi67OuHl5KrZeIu6oW1qoDsRlcVlJqF1WfI8QkxbWN4WSTR/3x9Z4Fai
AScfl50fnBF5r5CTbDIwrddiHzWiOJ6URO9mm617hSNFD8lEj13ZNkN7J2cob2vUtw6MysIHDfh3
Pf56Tx6F/CmovSv2DChbQNWUJ/TnvhsCXaKFReh/zsVD5KKHTKo798fXfyxi53Mt3hl5CKVoc8Ll
/ou6u7jJiqruIusXP7+DrEi2fAZWKnB7OwfVxdskFIV/s8xFgSGLZ6X9oFBsUN+CQlnNqIabvQtV
3V1PE0xgZHZfS4o2O2Ogn47VNmXzScK1Jb/qxRD5QYbMNxYYmE3ZvOkSCaBaF6LR6c2e59cMCYHc
OJHp/pDDlTTCoIVHeHCuPrbIwt1PDblEAr9yVVjUYwmO5ZayYDKsAXpGA79I6aO/sro5mPKJdEUm
YsBrEsJCLLXVYduGiFOvKalVahH3cXyk3T7criF0FReOUczCND7ohQE8fdO6DLAjfy/QQ7GPOdFr
adk6JZI6MwlRAQXUFpIeWh5lyGNzmbxIzIPUua6r76MBvwBiEc4OPhDGmaNOyVpW2aiZYZDcTFo9
R3WZ5rdxK+tXuOB7VOiWryZ9rXQDTJBSO6p1bTge1agz9zR51DkXMYVyKsdOg1hTDeyRtIRdpmwj
WJ77krr3VZbsWi2ypCgIWZlFWWYgAr0cBgig07iPlgJ7Hd7hgDyVMgGYizCk0D8GfmCc2LPA83vg
yyupfyjlTmIajQENxVYj4od1qDd7qdQaXf0/YIJPRYAGTnA4eHBn8aHuR5rrl065q3ZVhNGBtbvY
9pRVFgp1cG10ZqPLWANYQPxohicQ+QelfCakk20fFfHqdvhs05Lgv/evbXQFoWYGezXFmBjHj69S
04lvtWtBhj0ypTyHwYfBSxR+EABgdU4o6v50M/QeMlYuJxUVnqCIBzuLj7a4OO364PAywQiufagF
VQ7TpQo4sfx4GXIYhFALv1v7Gl3LKlGOR+MU9HOZQi/T+hUmY4XaK2BGnxHoWf46n9WOgd2KVQi6
wTZUFitGmeHTQ0DUGdNe8hY2qycPR8LPch9N2m7RWl0BZiAjTU44b5A63vPrkQoy4NJbfRfSxEq2
5QuADy7CMRD09dWG0NCt4x7kPi5G5xe+NZvcl1nvFWz6M3l+2KmP4D25Hxg7Us96xtGvtxngjJT1
tLctygEHcLFYEBSPMJOX0RL9U7e2EUHEu8CKsDCBpJFUTpFfN5ryzlsOxwG9uJ3/Wqnr/ljLTFCF
P0G8Rnla40aPt08IzQF1muebi/81KqSnG7YYS7HXfNPeVujMS9v/tWw0EeVYtltmJ6x/5CJ1o8oS
eUeoxXdR4VD0JIRTnDQMAJB0Fiz/O8wwYNZ2BONJwulObYT2Rajzs4z1oh1YnyaH8xuoJ+8Q7b00
TnakQBt4VmYz8hbmZktdhnn3yN9/247OkxBmm+f35u9IZYREtRb8t/+MBjQFmBvydKxdsCQXMXjW
gKU5I5DpjzMwNFDS0rXQLdnLaMZNTZp6ZlQHJmMWGykr7XeUhaA8ov8o8cN4DdVvZw++ntBWE3dO
TT4OSUXQKUigkis6k4Z9dM8Mb/QiR3L2Nc+/+MCkaxjBAAqMEJIbcZfBFQ+Q3QvmA8sligLhcqCW
UspI4n+fH5IsEa9Y4gFU5FWEZD3rM3md8IA1BAOuZQC8LvBv5FmHcNk1Aw+oXpRKRDIzCZaFf9Xl
di8DDzvbdZArx7XzSDOR1SaQRSAekcu+j3bMN6ClrtNRnXoPf7vMK809Wpmz/m8mKfcE0lmjVT+E
t87ronUmsghWwavE/5I2/nUkw5JHd9XMNdqYMjWJwt43CCl/4cR97ljXt+nhtzi5Rb/2k64BCnTK
Xb+SbphGH8jOmQlVojCZzAJjngP0hqobOIkVZNg9DD5aztjJTDupnMn+1uw4l/XwAg1UIDp9QvZq
9H8+uwS/c5CAC7d+r+HjbWzP3jZKK+nEQqEHQO2vm7TBscxxL1jo6uCfsqi64ZTkstQOBOt134O6
KwQzaoczXjlci9iB+KIER9rng119Lpxn5ffy0v3MkoBGe089k+mV5uTQqrOKiYV9/e4Ve9CaPfMP
+OAwFlch3SeXoRrfMsghuf+zQvuyZspxsOPqk+2d212ZktP3Ewx05G4FQkzYvdmEjIGJ8THvc4eI
ybL3z5dpLkcLwkrC9WvrEJpHgRA8HKUDhwKUuvEGi0r+uSRydr/BSbE3A5/xL5SX7YmhAr7YT+MK
kAACQioynzdaz4vJg07ta4erA+9mctzfwjE4Pe7G6vdtVxaCNs1gCz6RXWzwG7r0FN9aSFAbW5Ed
xHbPSFzCaYZaOESdyXkxe2q7ZglumHLbVqJeCctlFLcnAdHQbyET2ylxMAYiwR1sqZFWZNNGozfg
tRyjxfNl1ojtb+6h7wChn6f2xtTWEGZ/iEIScBOgHTu8ufsCHL3i0H54k6jabciNPKdNwFMVDOW/
240HaAJVhF9fmkrnUYpftzBUJvWcUO4SLF45HbGYMc4ImApbFDCKxaqW11AwqMvBI0lrncDQA8D+
otDdj6wr6cU/lcgpmfbmqL2QiUTLpr7vtuc4Lms++k20ITjMdGIEqUTTQNNu0YMwzkRIBw88ojjx
0tLXFlU8VbjHTEVPZDqCBbFSwh9eXHlWLSxgWoWCNTSlPCzm437Wvg3vzzB9ZMfh5zS4CcTFgL1i
Aj+h4omppFhtDzby6InCLA5WioWuuI7M2++vM1oMC7Q74GcGy8k1TCqV07oabxVNJvkTxn2C/8ac
T/iK3PT2iMNPYK06HaJPpjv/0Jj0+M6Wu4tp9Or3MvVC87aI0Czjx9dOgGv1sdvbXqdIh3T1n4/o
S4oaRmBBYMSGMtwmHU47xPb0wzn4RK7ZT4XNdd0XZ+fg7mKQ5dvnUl2ld2xQx3LbawrKgU/6ytKW
mv1A+1YEBGcnzMnqn5ZH+FN2KIqWfziTUS2x0OR/MgRFyraeiDxmx0Yw68NZHGXeyyRAI3m90Lsi
KY7K0VkqRzCv2qD3pHjHuTTKQi/NpMDE/3468xj4fkqSBpkQnFSv93k2CLimwE80+RJqVjr8eHPP
AW9zFcfWlhiTMDukog8nRtQQ5S1xzV/ocRbkCSmUPds1ggiybMRkyz12iZPfXCQ2JWuIlIXCRYxi
GwprYKc8G+YRV8OGHouhpSS2Ea1YWlNzCQQp+IECwRP5Gatlbvuom69zKJnlQ6E/TrypaaZNqqKd
AJFYJHgdSh471sPwkN/uPWMiHIv1FP3A9+MOVBoEZRr3G+xAdJdtYN+/gHSngKPF5wETeWBW9VMH
SAFcY2DT0p9jyZ6AGppNHXbWpbUZFxgZzq4Rav/60GoEwB7T1ZuIMHXL6UB4AGPNm1uGvLSeUomq
9D5JR0Y30Dcnr9GNoPdP2mOytlgACpWVFpSkPwz6x8RaI79ROTZXsB6A3laBkxNbLbHN2it0c1Tl
OqF/FLpq1Vz7zwAIR40Px8SHxP3o33Ogd1G3H5YrykK5je8dVsFt7asJy8C08OArXBls86WJCfB+
NzmvYWCK6nnRzgtFHjTNCUJcP+lblST/C1/LaLhhwby/ic44BHX52PlwrMMAWILA+nmsEIX9F5TJ
knfFsRhSq1Lbu1L/96emKt0mNvqm6y32BfBhOj6FoMTYGYTOzza7DF06vHF1J0mjGomF+1e7dUwD
zfw85tiP+VKe4AtcVjbHDVmIYaMCO5GllaCMzS7fUA+8V58M3X8nlS6kXp9DshUVvfBCwumid9PC
p+LKbdgKwFdJOt+ulILgTeJDR5nguEFHpDO8djgNfkBlUaTsgaC9ZXZQoLexPKAP027MWG0peaF7
V19gf+Wbp5vRKgQwD8/5GoiXXdOijBvhGmn6rrKPSGcM82Xd0LtiDdUJsmkxXVs5t24u7Zrz0abF
AZXqIYXXelkIiNE6pze44RiY/PBfR/YP+dX1iM9wR8THALsVdQqUIv5wRCxIYnS+8QmQJ71FYVQu
G8g2xHTthXvlf3ajqLZ+bXnCDTiQaxdcAlC3e9z63H5oUYmUfeVcSYDS3Xc9FWr9zOFAcdIfEi2o
+y3HmtVsw8o+9o2j3Txa3P1G1rVtP6zBDsxG3iaQNKGxw39MKLEZQ7G5j5zvPVPrzL34Y5OIfQPI
kOVL2oTlg7Rw4ksC4odte7KOHqE4eZWt6SfO8ygQ9ZZVp9CcwDQv3TqEXeITKkZjBZFgEl2B19/5
W+erAaypDGrmNvcKtiPIhQ58LZoX+iUDgn7pd5TYgdaw1v5RElEqQjeOVnnHbKnfml/T/tvldcQ/
PEzG4bB56jdagaUXsurJG5ZR1CD4rh34qlMQZepxzcnZmLu9LP7eTyANnLp8w0CEgZ66SQvYjK4a
2VVpwojVoCv2ZCbYKh3D1xc9Qop49J+m5UvKvhRkCeswNgMwU/Tjvre8B8ZfEeFkWBIDfvdvcmZR
iPfscJpYS9Ar/EblAfmhSzFnNT2BaAYZG0IC0uotkEQJRw/0/p8Qe0FeJza95t4lT9OAcBrNEevm
/gD7PmCH33qZJnfE9v8lFgBx1AAlewcL1oZJG/vWy4G2AZ+TkatNiDkeXw81h/SPxTGhswt/ZKJk
x4BEt367JgBRNurVOLSz7ABRnZorb2jvQhfAyam++e20KPU7dbNlEwvbc5cEt0WPr/B1Sxm3rjRj
SG5aFYKL7wfiZnPS9KUPswDb07JC4T1AmEoLHoE+9oZ/dgo2NJuYTRwFHJYYyaOncNTyrF5mGSQI
5Axe0cg2nPBmK5THls0vPs8/KQmlwfU9KHd3dlbeZWiwOK8j97crWWvC8BT9u1eUvuPxrBbQyINB
AV2DHfT7/jcBZK4R8m6Li0r6Sji10QfYEd0xy9dHN2SMb6PNPihAV7pYRTZU2PL5dyxDsatxdO8R
DhS8OrTpZIXljSMN3PUhbTjyIAFjpXUZwATlH8d0egPfaF8QkiXAQm1U2MphagatbO8MGvfzs8fk
FLvp3EmyB9orhoi907HqsWHtgAXNgdpMd0oKpPTVSVaY7xDC2st87fnL3DKGlwNlPcZkqhrZcK2h
VaidZ6wNM2Mq/3VwSEB7k34LABfC5+OcVcLFb4KhPXyhxwKhNa26NnepVte0VUI+zxqcD6YembW9
r703taxlcVC4P/+7Pp9RcqRQa/3r8V+N0pLAn2rgqBlGOHFgfgOQLwU1KolbbgguWHHY0IoAhdR7
4IdsmFTPAzJnbkfhBDoJtBz7HAYkpiAvonMtHCYBPYkTOZByRsXGNJ3FvzpVIeSrzxtHVFETevdj
qut2HkuOgfRBNwc//ztul9UJChLhVZXAZO2pASBxjj7is/ices+E8uwi54QQ9cUIRSXgZedVs71K
xc3vrdrowh+AOkkpLQKNX2GLlAgNJGR4mB+NYKOTlXBmlhF7y8LXylquh0cAdf2lsjiB7raNebTb
mzkpa4XkvpsziHYD0ZEIAw1jHv/8OrvpbFeTsum8mTMkriYPvzKpL+qsZGKAXOmBKpEJUDf9lC/y
tFy2StnD9DCvc0T5ha6n4w58UEHApPPUk0CvJWJxLlqCuqzt1gvwNScsNaPepkl9cnVgjEZBJT7F
nr2JAnRwwGn4lC2I9dhbEH3Ww6+qP2F8UHslLr8fFVUO/Xw8o28YfELSRmCKP++fuD65NvpjtkIZ
NNkmU8pR24gnK3Y2+DqBCgd2LfURFAl+q9sSxgI674ZGJCcSexJNv4KqcONX93fq3Y1czV4AOyjj
kWRehy2q/9sK+emYN9h/UBx4bPUWUMmvP6K7Y3yxQ98wmoX7ql4I7fzIXuPHCcJoqE5GKliowWEG
Z+Ga7BCETq1xTVPV4hZTSNj7vbKtltszfzJoHeQ+iJAEbYLGGG8FHHXZg9r3A+hjp1nxJ2rQ/f0Y
COELAROoShmKLNbLQxjymLRGm61YjSNmQnEGJVqAKGnPrVKIWkvL1qHCWielMsGQeH7NDEni4qAZ
6m5kGvBzAeOZpkVdVbSRifmo8BYB3h8VB5ex2faaVZfB65pPs9N3fWSUwLUu96rdwvUO0ly3nJkN
nqZmf+zawtyMemiG5c2VP7xxLsJAAJFtli65+Jd6y0lNlqWrnxYEJzZqMebfHMMSWajKj4tURxl+
G5lerP0F/DTDlxqbrJJjfk/OEmSG3V5aDDFTcFrzvSZ0YwAcTM80zWzYZ6dGu+uF+uR+cJcto1UA
bO7qjx0wPfdAFGOMoQLdupQnOQhr/bazaNkXaszQGddiDPbYy+yiaYCtCDazCBmKZgpGBjU6uQjm
sT7DG4j1lubTLfJRz69w3tpAbqnVNyCPw4IC5064jFuVTZ/vkAKG5WnY665ZuRWjz8vDO8CmPXI5
o04ojCrNGuQzMa4IeFhzGm38IZ+E+22pFDhNwi74pXnsBoG/jHiM933PjKcmomZei30DnETzGJ35
imw2eDzV5dIwQlTDfXsTHd1JbEIzdfBzHPjZD+qMIHJnKNmL7HjTblZ67Ft1UkF8VFUUXbHTIKq7
6b7gy6rLwvCkRmvZFi3AgnPlTSMgCBdi5YmeucBYF9U8H0Qs+3uTUU0ihPe4lUDEeR9ASTYAjJpI
eXrFB2SJySUNKPZuixtcsJ4iWmH1n8nHwHNwAKd3+HlEEYIbGQC1xVwNWoXe0UlnsKf2j8PWP9od
9W5wGkJztp4KQnfy6uxu/xhVBrZZSJeu6d/0VO7ocehBuKRtGqBGqGvUeCekLSgyFHpWVwAu4RfP
btMAkTQ9A4kXANuOdySvOi8FpmKcJ3PtLPxzcNepVUNZSkvycmsqp/pj68JcCgGMlMPjFAe/uIHc
JB/h+SBjTzS5s5JRCTWX2+3ap9Y5vtA4vnU91NcBxUG0wCmIOVGFOjZA3vgkojP+pqg/Wd9u3rb/
iQQYxSRAvztXwUEbAAORnhFEbr6qZarUmFZeGPbaTiELedNUy13mDpnOgNOZv7FsKR3vfLBxyQpv
jdnSDsUA638fz1vh/EfdmBTjaRuYeazC+qYVWDNrScR0Lqqb2T8bAhyb3Gb85QgZwjkX5G7nRQta
fE6X8RWMnDd+YeJgLES7e0PcoDxyAJug+Tq9zQ/ZxbO1KCkSGD1NQP5KQNv0MofFQISYrOUAnO7j
NFdi4/OEeUKQdmq98fpUR8wfacCf/pv+Ozxb3KJU7cZGaAbS0VHoBItxGydWqa3XuJeSLYDqdWft
vIHLuI5GK8xIBATAc1rOcntDx+lATnwIvuajWZ8bjIrcXlE0zxi3FviLVHgcHREUjAdrmCwZEmnL
xfoYrOYMIEXIEDA8npfUfdTPYt2jf9WF1YwcrmurLYUCDORdwCnQNl7ek1d+c3YFipQgLzF7vUIY
uJRP0+1beBWRXYAD8ewqE2hE/XXY0vOiBOZxpgd3ttDwtewxaV5uvDv2Uk/o8BMKMRf7iE3lyIFC
hL7C3TVDaOWuclfmUzsmovWIW6ZXFnLnkSaIfXaJbcsDQAR6tP3QFCaEnwSR+sqrALIGU0IT4aHW
/Wo1+1EcJl2UxzEToJCRSxLK5hkjsyOuPKhdpKxSEqz5bs4HxX9tvl9SdXfrqbP85kb+h7XaIpiQ
2kxemQbVXqiHYnFpDIhO+kd8IqO2UcAxUEETc94t56CVHtm5a09HCXysB3yUmrRW03aA+uWxkDA8
1Hengo9bvwKdKSR19USVKaaTAX99YqnAjGCaTItrDC7gn4yCdPKP5wyYcvqISw5gnKE4cW8y9ZpB
aGvQiKOlu+iw776/oxs1XF2tlQQRtns2YD3j32tk1aDNwh64xST5kM+RsRsGGPAX92TGNpG1bgoh
psDlY+rKoJlcSeF/Ajut/aXRO/iyAIrFKbgYLm6rklGKhVm4nvlZ+adj5HW9M2ZNfp782hG/T2U8
jDQSzQzWjiMKN1JzCypesuYOB7m+anhEYGibrkKb+DTb+wKRtjAR5B6rd4In5LtlP7PtvrifTAQ3
ei4WeikEuJK0ei5jdr2lZRmYVyEoeCAtA6OIMMrDmfQQU16eEQxGRyv3HIiJA1hNtNGzEKJHYw+u
XFGXPDs7Wt7jlkDAczv54xW35MUJwWs6VAUD0dn5rg0Ag/tp8faZIeV5++6tDuqIODx81tvOtCIv
r/VKGcBt0x+51W3XgEyK5+Uz4unDwU1PhhAioyXnlWv1r78aVMn2Fe7M7zIjiUlQLU0+D2VkEaIQ
NWk7lxbwPQ8zj8Bqgg4yM5SovHRiNIqRvF2nWLRLcajsEmHFAi7fx4mk+IdaSl5nPDvJj4jsHn8A
cSL+hFHQhP7rx4FgcqGFWWU4zgC+xSyyX10qZxy57JjwJkSLpBnLfd7u1sHi74kkIzPAepBkXtKp
fZTxu1M4vSRqObNQ7285Z7VrsEJzUQhF+yC28/DDiGS3P1jaYrwLWnRGrX5Zq314SlO4AIqa+yh5
2QsMNMM88PCAi3jVD/9h/o/oLxwMhGLx81jbXGdJLclEAyMz2Bod50EmeTA5BMIvvMaoJw6nJYAg
OVB804NwahB2rydukGhf9TlVxxDjD3VzBZ4cHcNbj7GP9fLRi28HFR3ZicN7qg0zYsrjXM8jGznj
zZRNqhUZSpdRuqn6ijrco80fjYFav16/L5ZYaf/dNO3sZQrXIVvlI8dBE+FhIF6s7eHGIYIY5MX8
dXMZlss9utVo//N3a+YkYakRKnDUfvooF/sONmVr7Msv8WmMkiDxLorCDsFcv0haZhJ/flwc1JVO
chCbmIAIT5E15bjuPiW0toPoePI5FCbhUasxVygDgtJ5Pp/8Ax45a2ndS5k7nrwx6Pk+bmH4lQPj
lgWbZFjeUL96kzFzdnJ47xgYJQ0ufOI2QTsbgNPa3Gn86AVWqkoPbNXJh+njvp4zoYN7tWqAfEIo
wXUCIMwfgzPMDvEJk9ISWdwNuRiKTyGb2sSRmbJ38sUUqMWpf7v+F5ndHyuWpwFovVNPCUmGM8qw
Vy3J+BnVIVUYu5bCIpwuZHq3iUbvLAP+3ndPfE1Vro9qM+WaU0KeNu3SIvr0yFjKIdV9kRt0mBaN
Bsxy38Tq2NAcGTUE589ZLB/3VAq87YK6xV2LIzQq4f0W0enA/feaUJXTn1MgLd/+tfMG72AHHQcw
INilZNcDWrsURoF81OXHu0RokhXV8p4NdsG+201Gvpq/t5R0KWLhseeXKRfPpsz1K8C6VjTcNH5u
z/l643gY1hpFCeJmSJ/YzzGaniryqwXCzaMA6eqbFCsNDQ0WCf1K7YUb0HTMqhD7B39TqOvEtiN7
BE+P6LIqHsz21pOYerlYjuNEzd99h+msT8QEK1GWB0tuN7tKElc7qdR2t/w4/AK52CpNgjMgIFPm
Hibl9qJOZB52BLFBUZS973imEKCXfkjQrC3knT3X8KQivMYWwlZ1pPBEouJLD5yhBfWsidH9Tsyg
faVp+4mNEx3b7T8nYaiPaLi8Ujgu615QN244PYfNzzh4Ae9jSkSL7NFbKdnzQOqchxxl7TN8KCLQ
qV/3cBra9TGK9xsbaBOBJhuXrWOQjYfSNRxF9b/a/dq3UmVFEv5jZNSU2/+Arnq1UHmtuoNaQEcl
aR11fqC/lBR0V8T1dhick9W6/mGJia9e6irLLoNNjb2IlFU0BG7RuEfEwdopC7XPpBNpxbRrfrrq
uouh3/q2hs0lGb4qz9rwP8TbB1I4Y9Im5+WC5t2S73qjOG4qVyY/P1x1iFgiscLuesdNCio8cyUV
Ya8sfvnhIsvDWagky5PpVcaRgNngbuJvbDrEHDdsn2WneXsLaGgfnZWyC0fOjAd/cowHEEmm4n67
L7HeqWdvJYboYIezCZBRpkVzVQptSGJ/+IbcXTd+9lh1jBaipbof1Y6pBuIlTFfyMZ93Jkq8kN3r
P8uwbz98xwaytrtvlJXjxbhOI0BfrlcFEcmW6+ApNu+fn1ncEV5UCFc5DOh53Z6KUKqM9PvOmyi7
EWSAUQTT/7dAS11hx5MDa13dC4ocZ8FkONWs05DxenkekAm51/5KItT4EgdDf962muEH0ARFZU0w
HRKPPB+ZQzpICzMTz7W+ERvLXYM0R6m3wneHEdwxQlbxeLJ5bpkAwrrV+Ip7r7rs6cSiqmA90/Bp
+3sln5RaJOJE5AwAZj/1yRaFPQGISGeq8ERbrvlOll3XDJXadapTWRMjSo9ZEk9RJAAYzLb7GgLM
XDUzX0aHpAykwUEEhAPnCgq/53/XeZoI7hfch4C4CdGTcwZNqftarwXNOyzqKfXxvQVRd0u9m6iG
zCqze7w/JeWJw2wL5JRkRzkSU8WewFegBTpU1DMT6yOSi9CsiNh8kGryTPz8VmBebuKfYK3SYNdx
C776jnS9QkXKYCJwbAn3gaTZKXLQB8I+ondKjm3bLiItfo34/TJ348eKpomxqTxjLRVu287nPLv8
AQdd/G7CaT/3S4IqSxvwKuMXJgOMBYcOzLMbgHEU/65d3CQqP6xgfP54irtE0L9Nk1jKI8hE+qtS
iWkj/3BkMbErPeGwQ/yFe3Y6bbrh4uVGau2viU9keC4fHuGrRi5/plj2e3FCH8hWpN2sMcjIUQKX
KADutHcjDDg7o/nY7wAl1WTnzbvLAHPzDFgUUwKEdD4oOEr1kyAKdH9Iu/eX6ibf15TvBVx43B1B
sRZD1aBy+CgV7Jm8DGOb8LOjW2Aqedi37fiN7Uyjgq6jBlCWvnKRbODGqrjOU0AegWVPoeiCFu96
y9biZO5mT3lH9OqUuxC1Mn66hIr1qSmQtrMSUYhultgN5mCs++nSWqyhw1xkXKudGt9mbzHWcKQ8
C5kRe9L/G8a8Y42y1q3lCPi/dkSaaYYTaHkoNHt5Cp6GH0/JjioMYG4PXySXoEdZolTByfeJj4n8
m2gkGCrC0C9iOV54fSdcqQvjLoM007p0xZ7NLxjGxXXnXBgsZPQDcSu08veiYVJEOF0mNiiUu80U
J7A5IXQEBcvflqZ7t4Zu18RPj3xmrBb8o9rRBzmZlLb9wz7Nyc0CbP8PfQNW9K+u3vezrza2mELh
fnQ7huiJDcC4xQGSdZrVU42o3l4Lv8qXMrHLTngk9q/pCnrVmUZkcVNi+dvVts6igOlSuL7pm9Jg
BdXOrLSdmGjP8wM0nHijBokdQexJW1AcYyTRVoqRQq5p06fLZqGbEIm32a9yGNDu5aYZnJdhNMk9
mFvaB2cC2I0/YXAfDYv0u7AF66mVrOaQJ6TQVUD413c1ZnjKx/ejMrRRtfUqPz/7jzx3LqtLHN88
6RyovC2oQFuXrWMZdCRRRvsc6OypqiFUZUiBBd6L0f5PMm9VWYT8D7MWTxfJC+giL2/rx0HdeEin
KpbIsNe3ZYkwT+ySmQ41FYD+RWaiTu4UuhWLmcQ2MoJB786wW+hIKnrGQLUE0jkDzkCF5dYPESAK
IIVsZLxUQZ2b/dgJS0mYEc6FdUCO4jHaUZApJEBa02PHDxeFNy57EyMmaSo4CDJ8C7p+hk1puRrS
nHdR1xDAmCliQRZBxBaMZ6nFwvIL7LCWXUSuOgjCmFSFCVgrSeXu6dlKUJtdjsEgejJKS8LXergz
X3NE7g5FPE+2L6fPcp/Y4TW+EZgxQvdpEbbrFBmTyvgdfY3lTtKx80x7bcxqjPL0ZCJFb61Nc6GT
urbFyqdXe5uFjaSxXYL3N/o+Z2fkEob6D7rOyK69hnKP7daoLVYtJMe8TzRSMgZ+wRSlgkfcOgoM
6WYMUjR0dIvgkc7751GyKyv4Z+40GGT0FXYvjbU1MZua7XnHIZAMLar/aV71hd9MU9ZHVwQEO0wk
Mq7MH2NILdeve1mYLuxKYbINvmh99b3sWl8TTBk1h1eemuKus7uXiJK3alyekfV0SZpiP6YgV63V
Psp8fbl7C8RZVmizpfkRNH/nDPuqovqCTkfX7qTm/PHx/Dz8e0Luot7hQILo/coUCL/H5LBNf+wz
/Yc+RHWGMkDALHcecnefidqeoqiCiZ3AAuNwAFGH910f/8HVeQesfCUkksyetN8H/N8y9mbInjVk
oFA1Eoau2zXGrWOpx7B9BFAwb/uP0N1ylfYqCRZ2nCLwrLLsq6R7PhZZW3vKmcKAJecSCDzQLMne
U+KHiRa+LgEJIYQnHlCpRiR2J5H0DHbMna4BoBDMIPOPua6dAA4ei/voqjqUpJ6WpUcQfluNUTuY
4fnNGU/i+vra5cn9fOabDoJmZoRZjbCP204OabWZnxd5zyK4N0Tsk5g5E/FqUvTdCPYrNRNqGlQJ
qPx4RLFEsJeaMnEbeGQYGXR09i4OTyYrzJ3mq0fbR1Y0/bw91bJOlg1uF7yTb+FB10LmYJNWTRm4
dHP9GdftvBJiOTUz0sEU2U7LcfEzuUkTYK91qtUwlMTvzm2CQcJq706ZlUVEOmZ8nZ5hbqfxQaz7
4/MSEBUE6L7ybDayVSeINHr9Ud0IJhOl7ocwivI1hjMiMUuJvL48fHTkTvYiwooLU1d/Q+DMlAg1
YloJ5FLCkwFR+TWT95Ln5E2LB9wQjDHsbu8sYVXm0jBJusAX01+1yruejuMvWQ/zBrrVQhM76vQO
M4AnDigZ0F/4VW6ElHZ/XQ0n5i/1Z3MKoUCB/OAY6dvROODVuR8TIq6JDQ1Gy0eIdjYem3TeZnZ+
I2VW2mezzhmu5u2A+KTSh9sgrPfGg/7C7YMlbo1yqQUD+dStqfre1gFlxRS0aJgGRk4hi4roqRQ/
zSQjViA1SL+gCrZ2o8EmY/eXirPFzc7kQxMAVhm3Qe6CW+9RJS0jNz0GbndsPS8goxnKwTQ5WTac
DgTzRIQUa+dAOrBtUffKXnO+Zb1CDmoS2/lNatQhawgdTKyhvi6788LbbuFHs+gE3bqVxUmv+Dsd
bl8PqekE19MdTwF2iY39RGkYX/QLgNR2lzs9X2OUWoy1/tg2n9c1l4Dc5vi7RT26kdiIDsPeYnWc
SXyx8cp5O0FFsk9mkn3CPJ21/9ZPXPrdzmhnU2NmpdkKz4AI8GI7/DNiCceEi55SOSVZAuhmskAe
MK9G7ii3WrWgrXWQtRd3TwwfJcW2yNW7ByNkhAE1bTXRla5gS6WL9txU9vKy+vTKy8w1Tk9rDSsL
BL+/G5Zygksv/DBKafK7LM6TBmMhVVQPfqH9eDfY0m2pyx8EKpokmXeWiDzUri7J4236ULX07QAP
midyfOA7Q3wVfGxf7eawFkkfUOVkUV50LAjnKFVeigfqDC5k/li6YSl1WmHYJ2S7v7kXI9JnVR1D
0M3Ipw0DbwFd3BxAL777+pRoqyaLPpBtRxAu/Y8o2gs1YtO2GPryW/RGDDJiCW3Mi4jVuCw/B79G
Kh/3+yiwLSC6397//4AG8MXPBxOrnvuybjWVbRU2lEZNnvLz3jFGjWh2DjjK53dVS7BAMnAjXjOy
9MqawpRK3VzrNBTDQbxc+byaoAnjaJMwYw2CJEJbroC3fmV5/m1Ci5P2XqlEFMGndlGS9XNoejr6
XtuWrlk/JHzxkOLf+Pyxicmu5B8lc7Y5olMjknqVqOPpRkKly2JMAxMgskk9NRUF8q1PqF9PYlBu
BJhX9r/6DtrgY8PXAyjlbH+HvZpaXjGEy7yO9cw/oRhG7E9TiRX755X3UKTng+HpM6VSE9AnwoMs
fGRJlzBjgvcgEYN/xQ4nh5XCsD/2IY6qGNpfQ+5Ucw9fnhaO/53H4Ut0hK0LDWQ0sCTfrdEI8fbd
bf3XNmMPb3BnPqnXMyVZ0+63ZbeLhc08T+XzIXdin8fWe6WJjSEO0n9oBY8AW6xW/j9pYftKpOVh
ikwimGF1ZVDwIhP7ZDU+MhS4wFxlaQ+JB97B75oQse7c9X8+UqqFDrYc4Yd0rMIVfHogkQf1cC5F
J5CTm2vdfzxvax4LCNl3BOl0i01xHnUQHkaY0xJfs1oprrf+Uao82QgpySOHR02SUKDSYg+L1hsa
qrGzIPB4mH3BunskrjsjrKp7YDiIvoofqu5K0qXUy08cXAQ/lTPGxjjEr9CAz1X4fp+mDXNSBqVI
Wn3rFmKZK60HO+tYEAbqiK4okRxAuS5LiGsdE4OGTd0XvZw0Ngwf5zZuadNtziob2UD9NCAtIMVE
bcwZz3KM82NzX3ciLPyrZW8kjxM9LuNXC/i0bpYPVaAfPlmO033/VyIGmJTLilRcV6yeyA4UtY5R
wjNblKFcSM/yP2A/WdCSiIk++kNWlb0AUzfRVhmNREqMEupclF67NQJ0oQw65IhIGjjJ1Rn/PA9k
H4nxUEnp0+sfFnxGlwbJWyHqKOCYqy8ELzrDK8kErgQ1QYIEpZQGbMxEuSAAnf8qa4lUe6OMs1Eg
uBi7tgq4tY2FgVabQSbyXftsFyyMXcLeIYH06d1MIL0e6tFZDKXtXTUtCNYYFp3S6JwkiabPsuZw
kA2pzA6+52tVgVh4n0mHoPGDabl5lB5iJehtMIMzj9l9+L3xghG9JF20/wOjzExPtKCeCzInkDMW
D7wBcrUmosgHgu7Q5N3LHEnAaR8q05nIY2b4iLUE2Ercj/jVSzsz6o3kR9RZeJG9h248eXjw3X3Z
vPjvo6OeeSAtr571+K3l3XN5T5Crw9NBNRyNC+X3cj4EXnd+wfxn+HgFbMNik3crAPRwjkbTWRFb
c/qbJ7AQ+VHt8fK4+0NNs0KroOOkWw5cxay82DG9ftKUMV8VOm6jiIJbPW3qGzTzsXxRpIXSpBTH
ZhwV7OWheL7b+d9W1ddAtARgDS2ZVthEDnSUmQqkH5HgON9Ac9DH6boOpH3DxXp2MUcDP6J3/Szw
13tdin0yqbZiMPLzPsAnGHFqB/w0WqBvnJV3595KUjqhURQOZr9gnHBVIkEJBe3EgQzWnSSU36fE
n/i35m17Niu7+xnBd5vXmMxfugs9aZScOTq34iLfNV7Ix6em1zjol8nHbcPHKR3/wPtf3XWyDC3w
jlNFUwwWv1VD8tpD27YCZpb/Lah6xL2nj8fOIHFnZRuJNduZ3+PpVVWBSds1ZfNGKpkR7if2skpb
KlKdUUzjxDm99mgzpHh2G/LtWQErA8v89nC6wIyQ+P/3Qp+TsTIVLmGwy/6TFZxX32bOlbNHlIje
pBu6MJHJYfCfNoEv0mQXnsP77kv7qZwZi8V8PLp9ewb8lUMNwwRwVCxZkH9nI6PTF9z5BJGdJvQo
jztpWCZoQqJ3WEQv/HMDgPY8c3h82IVIYG/6lCm4CGrwd1ngn02OTXvVoZfGnbTQNwye9AJu9MJc
JG5nvUZh1p66EKY1kmgoL/gQFDAVLjiLcAbokcJoYzWIvnlrGVfBtDtMEZSGLjs4ZLRdOtRr8aLP
47q3S841BAZFdhInVPewTvdqAB+2zWaN8/Q2lbjNS69185eELUFXwtn/6HHlI5xkSQAcwM84bPIk
Bzs6sh92hXzeqHvVpSEU4rMuHyWBvNh4jrulqcSFbXvJU7lLNaVb9X5irpnxMtO0lO2Ce3I6iCWE
IQEvj1LxLRSTDh0PL0djznQMaHMUNfr9QxZP+twVHg5RxGncHj/+jEueCJd2hJ7uu/a6XMPlQbAI
b0nd9mTYWhB2Z0jI8jddYjO/G7ozpIgiUndmPUGplMT8VrS5sveNkMXWLu6ntSvDB/HDXGhQPJDt
mFZpHUF+PfX6Z8dnriQ2IkjqNHaZDzJlEOoxLXYZoUZ3wIHKq5CvhKIJL5DdTYoLHedbdagB9E03
Npkcv247574XhPQUw4saru0B+D0sGcicLoMI3TVQV/oIYhj7WPcW81PKIrvFa1rTAntjZdJtu6uE
ki5JbXZDlE7DIszLOAGyRBYKbCSRcb9FVoc/kuAiyI7fVQb8UjqUX+E1YGuDecyeqNJKx9IdJ1yF
i4ijcXNBcxOJbci0hk6TDIjzyn+IalBgmfCLifGPtvbAbXnvuLexU4XJkqSHAxPZf6htAaT++c84
bcz1SK/MVhEWVy0flCz4n1GQaLXy+Rv24tMr6AQZg4J1jlCp+TXH+/CcTn2kOjx5vZx0OGGLwhdt
zwDT8w4F89qYcnGKYwYl6JYTETAsHp1fsFNAoS1eu5wyHH+qP75iLCzLnQTFR9ikVpfRKVIYukoy
xfe8c6XlzbhAG6AuTV3aNN4TltoInbi1z3c1EPgZClgYipXoU8yH2MZOjMuxyMg9LShnDEw/uOqR
UkQj7Ii/3Cs/HhhXO4L1hMMTjN6tkaPHCX88GT7UF88S9jlzfYDbxrMz1XrWMQrF2fecZTWO08RQ
Rmj2bPzo7xhIZ+KghOb9WIxJgPacGseEvRbeYiLaxK1Wz/l+iROSUglD7pUILJiH62lMKTiFq6N8
5Mz18juiR996MwqhKErXdpPzr/96OJ3boujv8vxPx6pKNEPKo1uy6jP2F0c/DGPO24HHRIPRtoGm
4w5erHVmIv9A3yP9ZfCIA3mSOJHQ53Xr3k0fohmCVHQr70d+fy7biI3QklWAcG/4RQ+kEGt9jdRk
UJqrz+7UU6PoGCpMOgjqGQIedcVt3zw+1Bi8h94WQ5pEKCkk1frOo6SmSMV2IQrmlKrw5QF96RIr
bMsX6ienRCStVXS8O15Pg4L6N2sopsMTWiVIgXTQJms+D4c4L0lpLgSsleOLhr3IQYll4sPpwoMV
nnHvIluH87NqHFMLYwK7ltBOXumqzgHqXpdhxnOezAK7KdNfIgn65Thx2FHNFaLvQsNtRfyCqYJS
+1Zl4AngF162QdaxjW0LjQ54lYhNvncMTEm1dV++ahQjpyVPNG8Jpm7/1Z63y0kqEQzPmTP9xuiS
nc8+BSJ1xO/0ZrldQ4BbKbQOOlx5/8+6V9DZTAfDi6uX3NGenhVYsbkWkrOY8NusJS0qPMacI0+4
WyY/PlALffO39lUwuc7o/R+py2v2Y8BcsORrEkO3wqsIqkZ7fDcieFPCfneU69NnZ3jQS3jZp+YT
SnRwfxLPG2QLohXceJphRXFPrgqQUtD+8bedAI+fKRu5gndP5EY2C75D4h+nORfSbuuLkbPatjRs
Bk/c7ogzBc1OgFBczvtYN13WrEMAv5GoIAC2YsnZOjihjxyOns14pnVqNJOWsHtehLP3vZnrAhO3
EOtKWPzCzu/PBNN4MVZhyU65Vp0itdBCjiZQzm9CBNws2VGw1kFr/ughugxNODV/jUoGDuwctDcn
4cUEiPTost1RpodpLAcDnQyhBq6m7LLfhNtgoi4jWHgDmRCCAIBsbdonxNAg8IWcW51W4epuAkCA
un+i+yhwulq/vka8sLZ2pYt12nMqepXsV2LSS0S2e+gwpTq/Z+ADqzCruOl9pUmumkjMLq7DfAfu
mbbABY2Q+VHMM3c9J+Gzbuu0WVV7DfEep1w8YyZHtTrLHyrhKIK46CYx1xhDupoY2laoVgCKp7fG
CdsCFEZNl+tNNvjqwQuQZ+lCEVuF7b8IkvakhrSH/lsoyWF0cqNR1u3inEIUoIpVRayHW8MGIohJ
vJgkL0rcOBhC2U/6kt8mIvnwe8rhfDRLQO0hwVbAPFEjAnBB5yNJb1QnFlXY0wSOWTdqGOoKh31T
xeCh7+67pdsRKZYOSkBvcSUP3xQFd4YLnpi14vgk79UoxBWlR6+EuGHRdC8C/HLh8PizQFerV4hp
A1aRkRmNWhI0t/0Q0uZ2qN8Pkvx/a5Yksgqd6F4LpeqDUljZQxKtePHmembunmCXoWcH+r1O+faV
sBLlTkY2IhvMh5jEWpdqMuEmGKnQUc6WpQYhVlv3PkHR/AV83C9aM7kyQRUHYul2CNvk+jNQoOWO
IYGnf5lrEa9dCuCRHL/IjQYlO1OavyHBBL23b01Axg6w0a4VQEJ8jhghHGtIVaDbxVKi48Ud1IXd
Oi+OAl6p0NFocqFTV+lOoq+TxFM+scDHqFCNbJjsSN10I1oYb+yna3Y748M5fQ1J1zAizIkyzeoz
PnS/5sy1JwJ/lxx3kSw7VasGRqrU0kGC2V2nNMNi1V1OMpkaHvXjp7gfcg19QDuuh3Fr2LgsB+yu
/tl7i4GuxtE114QapA/bgoSd0jcRwhl6zTTps7BROyFqBzKSXdFuRoMDlqyf6onnLZFArAglgX38
2Okaqgdys0SWO29hKYNkuXpiJH94ASUz734V/zGjSufDr3oOWlAHy+ARuvedQCaA+OW9H9564e2z
LIz/YeMbsgXb4bunKD9L6j9LWVTCcCvHRF9yZGhF2T8Nr2aEclRGowqCwE3ZrW5yLgYBNXM6Oyi9
zwJlnubUrLOlUe8XHAW9c2fKUDpteR5VHEVpRfaBMFcc1BSVwTltbghc6465vp5xETW7UsWR/CJ5
b+k1N2vOMxMEXRavwSrjXDXtIkaHFuhMJez7KVBoS+vU7n1IZ68lq/AOgWYvPoCTkTUV/YvwaZi2
CqPkwdqNXFW4s9YEjD6QKXYLnqLRufFE1O7hSzN47Znsaw5qlAGjvmX4MjRFuRfe5rhYkAmp9ImH
3gD/ZQR0kJUuBJkGV0OA4bPZZUi82FErQP8ClOoBJErCtyRH1JzO0X4+9u5mUUmEJLogWgPlcl6z
YLe5LaJnKNj/aV0dGDBPqt5pXmq7IcSivq4UOaWxijmroNf+02aDnZyw5NAxFoGRNQQPSDpwcmKn
5Tc4z4UiGOLckJZD643LRndeAJTnDZ7VSgYD+lNxUXjdxm7jBTxnndVNbkjrWDCqKWa97+QWZOZg
JxQlDyGGQOUhDJKS17iNC5NKzw6xzdfYH99D+oaacqHRP+odxyIq/OfoIHsbT+6QuAV2A2oQ3d4m
YyuBti/3rSoV1mdNxul36S4Vje9NPh78rygcYik7p3s2B3iRhcD5lkfORwArEZtcgat931DU13wB
EfcFac569UFufQ6OjuVz5XaVvx7c5fM1yVa0jLrA8NI6YbBCop+Fzdfoh0Dm0S1av/si33P/9zvx
Pgh8SXrHy9E3pEu4OdzPam0acqF3PVSd+EwXNPeuU/KQR7M4TGQ48o8sIc42UzusRx0P/QuEho9w
l+t9k4zzQZf19+Op2Ke8auMFOJl2qFcoLKdSwBJ6ZEOKwOUrwMOZJYBmTinQ/7IQ6HC9ha8LoqeO
Jer4TvUX5ds4aPCgDC56L5bOO0VABIVNTpmSb0kvnLCzwctlMJNY4xUGvQu+ESr3EKCU/25+rCCH
h8j50Xr1VLcMUH3zhvRihxB77z67x6Ugn3Ol9GL3QGNRTI2xfbsJVzIQ+qItYZ7uRORQQLzzBe1Z
ytTBCONl/0lKM4y7nq5yzKaNg8zvaQ5HVenWPURAE/arNGeZ3B7zQRh2bCIdGQjW44q/EAp/499V
a+6wLniYwRfVfXRdp4fRZMW0C9ITQlhc6lNjTmtHmnb3eYapZqqXDRi7qdqfRt1gVCqkwOQgXKpu
czBxYuAARikEuEWikquhbzTzqBSIsycPi+SllhDnAcXLGR1pwk5mQHPbPq665fL15xSR5I0nxn5+
APg23WBDS1H97X4YCfLdzF5VLgwR7/E+NJc/UMavNq1Ks5EPZugb/mtXWAoPxQcAVZgKPH0Orpj8
nXw6zGxCavtn8kh45rpzMv7PuzmOpWWY1l4OEhD400DBA1FFRJ1LPE6XA0t2+OA6h5WJuBt0rwTp
5BNmVmPk3bOId4vbDvXRKBBNs7f2uF1H9a5HWlCdo+l8b+UPd88A6hcnu+PMxhNJt+p4ABAer2h+
5BlP0zXyjTO5YE+dw+6DCX3vZAFCkwpQX7a/yAe+gHtcXmEXP0ZhMxKQfTbp7Yibfbd1us8BCk41
gtU1LY/4ConH+YPMUaWaEADKFGcg3bqXwpspnz7w4YnAywRqlSNhxdGPZPEeDD0wsg/IiFLwdwYt
fT/zO68V6ARyC3B+xdfPAU/jqa0w0Cp7hgoW5btGiq5lCyx/qgL2XjK177gi2xUhhvXsU2sdQni8
Bwf/N0Eg3dll6Jw+VemhdIFVTS5LP9a92CLenhvgG7xp8W9P/dHs0W4DUClqo5x03Y420mPozLJN
sm4u2wwqc27VXKlygwzdh4sxN/I0VtYGoAAVRrTo2lpSx+cWT1xbim0OO9g9igcbKAKSqciRfgDq
62tTzExJm8Ctk3tvjt1jD1fv33IEbZvjUpOb4gm5NWt4dA5d8lnuN+WWYWV8W3gEZXKvhqnbcvVK
m8n/98F0R7bBf6lW7uRbs38gvxQ21fO/jpWHfGTEtT5TUxHbaZKo62RxJl+MZsVDeRiLdLd5k3+c
hRpiOcQq7OfLkW94t4KhT5FQ07nQf6xxxkz4+MYgBM+VuHhSK02wvuKDhCq0m2QQh7BGpPkWKinT
LmYv5iQvO8BYGgJgvU7c34EPVSp4ToRJ9RGHG4dA/1fV8xMXEaLudkGHqb9n3Iu1OZUtF8bpR4lB
2yDnuMxaRkv6QsjFoAiCkadjpvfqbYI+F8dJ2nqB7cqc9HMCkcKmEm50KcA0oHwVOur0srbo0Y/g
W1KA3RmDgi5IXWlK+tBl2QPZ3rhFY2w/PPKf5LERFSPqMu9ATeDWabuNtQxwn1pAOK9fTln67Eya
XO7xBBD5JRHAjyM1LJ5TqWrVg9Wy7Js0i6e44dwxN6DSVR5hHUGrtdmpb/DT7G989EsZ634TPDvu
kgaa5nDesVosS0YaqsrD39vm/d8gLzciL9KL0EgpSLYJ5It6f7LPJw7CCdlQ2TWCqeUt7+a/6SJx
Kmif7ssfUlKjCSTWxJLOn1AUgTlTKd0F2RK/kT5mM09yG29xrU1ZU4Hh4QwtNoQeQS4AldyaUfAk
eooTnx8aapSQb6BM/t91uZabW8t5he7jXRnN1b61Yr+laIRgo/1OKDCXhx23Jaj9N6QhpoKHnRA4
C9ilKoNCddiL0G+y4jpC3ga1Im+avWWiTQVO6lAFJVcDRUzElOwBbBSCXRVpTkI1Exo0OCUv9yta
uDgr4yKYb0f0EQhYSFwuZENM1D50F1hKh2XI92cSBMK8pIxONtswClWmcUJ5/4rS5vwavt7Z+H8b
oFO5BLYdX6ZxYrc65PA10HW/sr/KmhDUPIbJ/g8WwEm05gIZE4eMDtEvYd3muTfpgzzSGhBu1836
au4KnrljY3f/cx7peV5R79/wGDOqsBY6yoOUCg23R0SabdYqy5XxyDydJMFNQ22O4L3srupSK2ir
mod447ejcTTiH5ugDX68U9LuNkdp4VqSXvmsWZIfSYJTl695cgsaFXch7WX2bYis/nCE1nnUT41n
pEtbrD5FGlt140Q3KkzIIKDYToekN3zweTTEGVAGyTHsVDPnY46tOrdMWr6/WR7vSBuKQgsjwOEV
T3kO4EgR6hxpYT2LONtj/d80ccFNeIag8cj1gP+nKzE873XJwAmbNAe3nYBaHqN4rb9ql7un/2jD
VTzVYT78BD+/kUDGBQBdTlRV5TfoNZ754WLt5qyONSUKCgYbDDR3sETT7X546Tte1OK1MoYlisIy
ZaV/yko2JxaRXIyw7r0QwtH7cvLVX+w99giyKRVm6+znMR0UbmosxGxRRZlJgirbK6fKcsS4y05T
/760U2jW6UJIcPOp/opt5MhzgFOL5IL9QcOQPUrFKGpS33yiohkrqb8soc76MSFH5W4gjGZxIZYD
5lVWcbsFNcqzAGaoHRiDHFao+t5yF1K8tn0FVjKvrATir7yhyXrdVs5EkuFG+6MFUhbcBjT7zrDz
yQww7Tt4HJ7teXGTAtoiegMOkf15uljglMHvV8ZmYtmTPGzRV0M0HEcz6OdrIOrUz0It+pJ3Rh82
9yUxlXF5wFzxyL2oshx6cCY22b5uXaKANqyrOFTIHIlK5gJTzn5Iq9deicnl2Fb+xG+qPKHTLJ9n
zkVYMFbdY2zqByQR548zjB+XUT0feLbvVERias65ywV/Ov3ulHI06AmMPQnFC2PAw/7uHWvW+0X8
UXqVLBBSKWQAsOHZSZYlSrIBHE5UhG/hei4qAGFSbBDKIQcn+ItwT9JPYL3bZUYLcqOb1XEcycl+
jTjfYn6dfPj1mgGY8AEUhBbXQYTv1uyMD2chTU7TnbiZZbWj1GvNEfm3PaPRMnXowLorpyBPE4EQ
MzJjr2QF0+oel2K63qmk8xhJO3Lr8ky57NOBLLheeeP9sJyi2SlW/wR75apBPcaR4jpId/jTqWZR
o+uUvSWXkGpS0hNYy0T349mYL+qqfKOL+wtf90EUsl8zzaoA1wu6XntcgwxeUZjhCN48Nmyhy9aD
SlBf83F/8+V0qYuqLY/IeNhiUBoP4W62kFQcKx51tGcU8rTjhtWV3sS4y6BsEQjG9OwWCWIQIC2W
YXcSKeWL7epxQc3BuLS13fiEnPHthsKQDjQ4hj4YfM3mcib1k3Mt8whDGJMIZhrvyqGvqAeStHNI
ul9ZmEnI6DfHQPzQKudS7Ot3UmNacDJ7C/OoVYq9K7xmqRJtV21c7q7EkRkZxMDzyWGjmOxN6Zaw
ICBYo7oSdLTrfmvLZCOkZdWBjBQu/6FDzQVq97NnK6euz8ArJF6wKsnRg/X87+J3cZkOzLmwfRso
z4ZnBPTn7B6hcTVK1AALbesc9NBrUmtsXo/FOR1fw4ugn8ifaZjHJB4cZxHPt9nxkJ/buEpQ6h46
wi+//ZfdDE7MC49Zy4eRsmHX8irXa5MwsOvrg+aoFSDwtLaoxC34Rq8BE4zVwqIouGWh/36j+hUR
8VWfgTbGbskIe41I18ozCk5YwlW36cv57fpKmrUkEJLKqsRlpqgXZivQhgCiyXxJ0wGYmtWH+/uj
rpEAdIxrE+E3w3ogwbvbTiAaByBM3/fQ8qrcqJJyRGmu1eqAOeuMtRuatCHGKwlO6YfRQ/z0Q1kB
pM364Vdra5/rlxli1LJT8betg8iSIMN8fEx4UPq9JaLIVeBeWed7Wjrrl/lbZfKGvY4t6C8cT1Eh
ovaEg9WXeQ0ZZAdYJSRFqpfTPstJrU6YerwFzwEtm/QfWWkdIeel5acHYg2/BrjFFM0HJriCoogM
LMhWrc4UzZns41MWn3+coNIb5Ln1SOQWAYvOzmlLdzocVVPsXv9D11imn4uTa95aHzwvm/NoF+ND
w7bNxsxqcnE3U3tUqvkSyKNkgyj1/3YcDlLTp9Uvr77XsEIp5FNZAtm33JjAADboTpzFOGO+gTtb
N79NiuAclWs462RLstjXrUJ9aqqq0tCF3GLHhZhgmpH8mrHXxv+MVMBYJchQXLn7jyg3+IPc2+PM
OQRLysxBSwBHWekvp8J9jIbBTIo87m67XqTCAdDCToZZ9or2x/vG5nDHYW2Xat901OCvVVdHaveO
FJjN/+bRlpQTyWlIkA3BQh2hbowW9H4/yvy01DcMMTtsVPgzBUwlLGpOzZNZ5gTAbH/I1BHegcGc
Kn41RshPVxiPcfAL18/MM1FRKnRShCyBibtws8fAxBcIPHIAoT3rL3b0iVUtBPIEqKHBshjKf417
isF5VbmRANh5EYn4FtzVdwTTb7ine1/pQcTyXznCMebmx8xeeZGpMv+pBS5MYAdicDUM1zyvxoD0
7i3o9ygKv3UO/scJ2nua3NWDtH9UFsXSX9cq+H2DH3TAXFJKTdG+XDFCrkz+Odx553iKDSEYRcG9
qzhWVPpuK3iIBDdDUO9tXd9oSzEUCu+qQjeGrJyMww7V18fO+Wd6/aUBpRL1yMPrH8sGgNmcuA6x
c/Et1dpWAYfPiRfcEpN8rcXHMuUTNM68BWWMtKCgSpfYyE8eK8i0kQRzb98JHKcxA+/PnJb6Yt2A
zYcWRjhYr9Tqs755jYznd1w2OdGsVlr3bnOCIgj0uKkYmH0JAoBttaenEWTt+sYpdxuqeJC4uEfm
SibPAkSu8MBpJ6BxrzPzek4MODmg59jYl65s+gz9dqdpTvb3NK99P7zXM1vkFeuIVXVsxFqHk6A8
lPHJNV2HVBjKAQelO0v7NoXPttCs32l2UBTVrHWOSEBS8ul7JrS6jODkc8rV80Oa85Nb/15vRKYe
lYX0oaGdxChkuEcBYM3f8IxhC1bNhMx2l2YMfQRymVYahqMQE9fRMv4VBgU+00Eb4BYDsXL+Qeu1
Jv8sXb8mKLmrjSyzOcL6dKapjpooXZsjMFH2adGaKTvgUl1eDX5ojigVMTMEwCEcVUi0GZ7idhVS
GxWYvkpgfF6BIJLLGfLayNQYk/wr/fIAyG3RXpuHlsmRkZlEMeXaitgx1gInG26LYw354ABARe8H
03dYY3vQS8qGmPG2y+3lR6JmzAmZF+5YLHt1O6qfgw82TAQFCmR478Q328R4HgYgTDX1XBCAdNGi
YugsRYE+8fshvFKDLROy4hrklRvCdS4/jqSfgcRrcFUK0o2KIuLGQ6bqgyoW444HIrX21AEmuxL2
wfAdTTlGXPDak3kWwa+PhkVGVRuZEwzVzSSweAwCbyKjiwHLv0+0k2os6HuA96OsspPJ2iQKqIjO
DYg08WFHAzYbXB9lk2a9wREUtDUfiafF2RB5OcAXAJ3JW/oIEE3tQc9b9Z/L1idbC//kfVjXZNse
gqLd+r+O+UB1HxjDnjdOP+WWKg76WSvkPCyqmuiwIh/PliaT2RdE9w2O5mY3FxG2jgWXU9bILEO+
O2U9GSkHQS3S77oVybgeW77f/oAa3umcxCRjA/8bUaNm+L1Ua1c4wftTJgdORgekujAVutKfRVCr
fZOWv17AbITecViDOZtUYj4a+EC/7J4KzmHtqy5/U32794RjoJMJu4/r5NveugtokvDH4Jgq0kmB
oRo36BrCPR0Tbow1SGZKjwKHogoLg5duliIR1I8tqbrgAgNQJsa0qk/FFqoGgtpimtx3HoPPNNjI
LuGUdmGByJFIcH123xcoh0BBl8z1jZ6n7DnE6f8GmJW/FsYJCMWffjMKi0DXRKYbDb9xSRbX1Bxh
9YG71cOr/zvQLTSpclIugccYAJSLVIU/y2hEBj9HIwslc5nEdAeFhwWvbJSzr4dX9SkCEk9bxStz
e7YEs3MIWmHrg69UDRJJnF1GSRhyLW7wk4NR2T/6D1Vu3IJn62slORwkFj79bCMw3JzH0n0wXgf5
03xVQ/besHR8DB0ndBnVXFuMKdpc6uU9enL6cenYSuSb/A57dblscHuNo7gexUbQcVLrqmkj+YoW
Up7RIF5tDPOiN4GEqpUZbFtFNcbukDjMvZSC6cBFb1ZCYBg8SCSNu+FhR9uovW9aCcFEPNnauEs0
Bwh+wnuGCuC0kkrcXsc94SO5Shc3Yz7yZJxuLOpKcxS6cGQ6QQYZ5Uc5moTry476u6cSUJzj3bkU
7TuuzIiQ4oLx5FG205hp5vSRTaDrvapeMYksu3cQ+ctS+Q1V1c2PF5az42A2hTzSA7tIKT0xxBH/
/n96qm4ta6Aaj0gFlSN5v2LY4NL3KOVBD6u1nVZzk6l8fm4jLYi5FmQDMuDuDlDDZ6Pltkm3Snyw
1negNfRCF+IYortWOqprtTnIDyBokP6n4T3+xitIFqXWtDjlUyX3Zp6S2A+h4Mv9R4rieBy2qZlS
HAYnLABZerB7/27tbfUMtxs+7rXpe04i/64Lt+6Bj0ZGhE7UaVBabJCTYZtAkgH5XTSoZTjjToIO
z9A/evwrxysuZVTKSjty+cdAyt3RBJmKz36O6xICwcy1Xw78HZxnl0IDR/yAwIIyL0r3UEYU5RtM
Hk8sAczlM3/kaOgPGbVMIW03/pKupM8Ma51l/kvOLjWLeI37l2HuxhoU5Jk/guRacVMKaUKaNXxp
kLnT6FhGspSN+C5k4bFSd+LuLcsv5PmK2huxEHcPU74gCrv8wsC59NIcRDkS3EEDyi+wKDJlXxYJ
GFbuGbGODbxXO7Ufq3UZATCEkr1HpuvhO+Hpg82gfUm/hxBz2SXO7mG5dkx/T34As6kf0LXdhW4+
1NeyY3nZ7s5ggbJvEcvd7G4wLvE+MT9feWIZy4uQTYMeaCnWcz0opBrxkj+eFw9r0q/B/zIuJTo2
QF2brQyeskRO2q1mYLAttD6yYgpnk8Fd/n4QF6XstyOMh2dFZHbgiNtLbRKDocAiH0m52cKLl/Co
acXJuO/qJiq8CO6j2R3urYCOEvIFik12vvm2RD+hVca78ESQYNxNhdiIMPMGzrmJ9Sdorvt0nyrX
STtW/m3xzuvq3cMzlD110FZFhZiKCI68f/dLNdA8FRJkIRnudjFFrvLyDTDC5lqlC5v9weL3JJLD
ewRPtcD7wwVU9MigTzShhwkqJwFByw13I7YHjtJG9/A/pt925ZpCpZgOZDc4JyLvTWIZILNesAj9
Pczuidkal1qrgW0U7BzjN5YVcUKFx7fHRI+Y1xmix3uNfu3jNHXTevwHVjImuMlExw4dagu+hQL+
XX0YebmZ7Az25vzwAVSZwBzK024pppgyNBoUSrwx3aPXhjfzavRgsXgjmXVcN1LHYbbIaS/j46kT
Cg1xwzpH19ak94DSfjT1CWDJYB9f76SxURUOqGgkJd/NYW2Ve5gDfoOv1BZgjXUS5TdWC5l0g9YL
SwaHBWsYr+YiP0RrmReBXsiYKHZLkAS40Tw7cIIHw1MCzFnolWsSBZ7519zpx7G6VWjcMqAVxm+b
WYYwX474ElryV/fYDx5TZSgkU/IomROh2vNzt6t5J/oj9918643L/Nmh/3ysaXp16Pxy7aeJWAur
Cq1F9LMfhvN5lwyz1ewrnZ8NiEe+UXlR8odHLgHHeRRxV38iSAaZxBPNrouy3X50e0pvHMCnZP2G
T4cDMYirF1TeMNZARz0jNUrcQPZy7+z9ffx+E2ypMDMVBOnXvvQRdGDGOoGKXP16NTNmDT8BzwsD
AZ9jJO6tR5kZvYAdrOn2aBL7sLcD1xVoWDM57UUHE71qkZFA45UES1POczSpLZH127LMaqIHNzAo
f2vk4ie8f0v/K5XAsW0AqqZw//q9VFXiQrZVHs7pQjc7bXf93DahBKpKLW+tLMbjbUvYnoGcc9Wl
ktRqNdzCIclF5w4ymAeYygJ1DGRkvO/GTSZZoGbHO4NkTqg9Bxm2g3SO2AF49TGsiqkvBQrz14JN
/N1itWzLMhC0fNtmVs14H/FvVmuqz1iTnodlELBPKP1is5k6Gm7NNLMb/4DHe938Nhe1NfP0g1Q6
XjHQ6Kg49uLZu/SzAEZMcgoDC8Ds/EC27UAzoDg9uPyfuIaG69hGOv8wrafXKAXxYLSXRn4JKtlE
uw5hlgjznypPkpSEOZ0Q7M1slAJuqmRKB7EuVbM4afmjiWc7C3AByUrie5zXS8uhiObf27BrZaWQ
CFfrh1gvILp+yQzdClnK0KKItUbUNWApMhHqhnsO8EVPfyxr/DDMyDBedrSER83mRtAT8iymyc68
mXMWtQ8s0V98stmQp9XXxth3pD1ME8BvI8FBuWsv2zv7vcSi2Zcn5ICM/LCUQ5OLOOvtcKjEoCyY
llwSY49gMCXPRmZ1cR1CNwEkdKWMNSTQMz5sW5NSirXXIAf0GZPFmNG2IZSaKWVQQ/w328jCJTql
iJtbnnAx0/IUc5p/XwytwvbpjLmrqD7D9bKZxfd/YrfbhqhxL5MHdnW4X5QG+d5LdkWSA45Ybfgv
TyvSQJHoo6dQJ1MSaxnb3R1AoAjybt4Kf9GzvNWUAPZK/UTKA0nZTfeJu7lChLIGietzNH8BGoLm
vQNrq5hhStfL+zQQaB+WmOZMEYCGCjjlwAsLPIG2//QIuwvBUliOKmbrviYgsCZdzO+3o/ImdJB1
k0L07SOsPr/783egzWiYWW7WzVwpk9bg5laUZMUcav1uowh5VebjTwFtbJ0HuJVM5VlfXb4OiIgT
nRQ/47s47G+FOM3y1BsaQice/xeynYdyeUvWrAJqFtBt5usqnf0dkpHB7rwctOqPI8i00f6N3rHn
MuwNawLDU5Vg1Jcj/zaW+kFZuAWC86Eo6iQhR+OSDiuHZY4moTNPoaQagdZFlkHUsYxKyW4u1iRV
XSl9VdIXdoyjyFhzDBl3jTxgE/gGKpGyC+0oI6P/nEfpFHZwDUs3fwoqIUkwSDkuMDqRRiMwjpau
ywqLzDY21kdVibqEybWbemH9jo4G6IZu6U6HxXqjjQdzY45JOHC8veApH4X5VWPtccChXxO6OMLS
3S9z6hJNhz9O6bI6D5wP2ErC9wSlw0Fv8IBBxHuQw1f34rcK5ufSo8UH9oYhPb8jYaqUIMpXORv0
ijmFBfngW4nzIPFZec2fz5N4VovcAxvB6TmFAg9G9T0/kKgk3SiZcMIzGTsA7CTEBhC1y9sBe9v0
fJuYw6FgsXoBtQ+vI41T5lg3hoM/R9KlTqZysJ3jQu1ckRAuetRoz4k2wzXUTb+lmvp4UVwR+1yF
HEjanLKJzvzD4qw/66ZgX/FtDpiGRKQa7nZWuKq/lpIN+3Q1vYNV7H2oLABOyHOsVr1E9V/dmshG
rM/+ootA1s0ZW1oZ1r3pb7zDsWz87xqBFuIk0qVfamLuKjrWN1ioyERQi7L+w+iw20bXuaV1dw8z
fHlZrs3+Oao+GYX6tusnjWxYkSHRslsyNZKngG9NamHugOcZVHdZDl13k/br52jVH6riCQEiCmqt
4n1g1gjsRyKVMg1mIaBM58Z1XWL4G7VEZTpUZKHXWOqVuHQ6l1QK4SmS1iWBexd8TcY6ei2U7rsS
+7fUHP9GC+StjrT0x7ufeeEg4H122OPIpDI9qhcvMOq7ef5z/dxoHCzhFoW/En7mef+ykkwiPC2/
3RdPYiCCEBD7cEgUCo48mO0Lcl6Rf2yCi9wXPRNfkJ945ht5kp7pq/7GZTYtDpp3FblsDVYZURmw
kx9ZmoPJOcBN1JZUq1kaPt3OFgFo0eg2XnmaZh46tVTRHfb+46v4lqpki9yVYo8SwsXTVS1cOvpi
YrsswMIso8D87JeL8QjXQlDndlvG7svg0G/bh3xKpnEI6dXkuD9yX35vobNTpiY+9QBUpDRGFcQ8
t1cOll/hTXTvqK78kVFwGZX0GfQ20VGSq4PReie1eVI5DPUol9Rm0duE9fjRuOMkPa6jx1HWC8Io
zF4cxwK+vOrq+J6BpTmJvvSjfooLw7+Qw02PiHHRfsYqIVXhClaQIYm779y8C3ea3MIQda2VSWcf
/7xuIkMETKyljwZBaL+mSafhXRxArDq34u/K/4c0sp1NULPAkGoRi7X7lyYwx07DghdtgfaUoyAv
fQ6L+ogwCDhAJyN+y6la2xl++3RAXg3IIp7Vhppa2iSgmB0SVqf6wBz/n2boUQn/P13pxsLi/0u4
qq5kFxjMMHWVJGV9LitWB7hY3BuwJbnhsoggNm2LLo7XJSMKBzgIDJuIxgJLTLxHWSGfMeq65KwV
QgF+7shF1LctFHwHsA/TnprLZGbDbsJYWSYcDWCdInyR4ttzZ2h/6stgr26KpkVScGJj/YzfgYBq
xiUAgcodEsGIiYMV5OH6niTMNx/WBC0cNPciSKyvVCwZ/9q+HOS/6lTrdUac/HrM7nQMhP4mMZzy
peWdymN4e8O2uu6KDqI037wPrZ5HYs6CrR3wUrZ0Jcljlrxe30fDIvochi6kIxvEKTDaPYcsD/uT
tWfVtePIXDivr94F/DnkJz3/ofN0e/PQ5H2zyeRc36HEeBGgczj6VxKp3HIP7VrpYAIWGvKsiHGx
d+jSYuqTAKbbA7Skm8Wgq/KxHHm+rBB+KBHjXbVBtGTEPf7Wso9M3Y1JNYn1ft2OXDGkfUvVIl1W
3fzBQEQhXkLWFc00oQ3pDHWbDZaUGfAYkyGx7r+mdaJ6n/UQU+uP5/sQuj8mUmfrWYtOoxKoo2y1
oghBuqYcoZJrJmBYA5IRI9A5J/ZFAWAycTgtcKodjF4maaHyvakfT8NeCTeewJAdxR48nS+8Ld+d
Onwbte1ebt6o0fNkTA1HjR6OrCI7MkI6ub9y7Fo3X6vKYRLxKbAgc5aeSjwq6RV7LDpsymj/0NZ8
HfyfqGEjwhcXGISkb/Sjq8/Untg9Gx7y3af4AP2eCmCQdwq9zfmaf2F4RMeeMH70J4Z+nK4QFauo
GEcvtks1UQ/gqIwndRswcPG8VadjFl1XwnmeiMfMiJhaG4JVkNfayTjtqIBimTDQtOJobfuBBsis
VxmwvjwApLRsgj59T7Fm5/r7HKUyaRcb69FzTflRvpIH88Jnkh9cYifxXI+O/GHcpSNut637vU/T
WDltOs6iFQs7zifZ+hd3TvjUIREFu/Gu7lYOQHkOTCWhG713C41CRFjSEZAWMlvUHACWRG8oVMg/
TnhmF1Hvn0TFiFEkcylAhk4/52hTovmUJJKKbRXop3QThrnd+RF/UBLlScoKDIJ95R3uNurKkyRj
0uMRUPyiWnNk6FO9Z2n7CT5XchbGzlAinSyqW4TxufW8A6/Q1xMD4ke8M2xCWLMyF80KSNVJEh7e
zGO9H8ccucHsbxQ+5OU9LfAtMGT7lOe46rSJ5oTrAb0QaT68s+G1Y0AkXjxnWe6lxZgngGVnwD0B
kH6nMUg4MmuE/0zT8IvdIQyC7fm+4qqdOHV/tH9Y+CMq+3le2p0YZgV27IuJO18RCHI3yGRTJaDf
Jp25RbtuhXCHehYEcTvspyTEAvhKrWblTqf9tXnJwwlKBSBVhcWS/AVMprzwjFzg8JwZ04+PfiiR
3v+NjZ4cUgHfCFRZ7FJKFyH//ed1fNKCfwa6pS63CALEc5dnahRLn4F8/8Z/O6FxRKz/djgsBpjl
KjG71CjQhqfbzEvK9cOdETijbf0g1lw03rn1V/N0xu7vJL5zUyl5ZqQ1Q8pKvSJ8sV8wUlNhGmDf
4BH2XeQ3GL7nrrShxAKuskiT7DFMw0dDf0IPSZ5gOsvtdmKKbgvy6bALkvlJgqfsizuhaw8d2GXn
9vkvPV7NZ2qFbsje/Jiz1J50Z+TDoZB6ODiR9zQrt4xh0QknnsoD4loR0nXu4K15o7I0PR+vjZYJ
0nUZkeqD+cJOGLQWdKJduivCADYs8QcK0w7a8cL/fEC4t3rAdxahBioKtf+UHZqShLRdLiZRSjpg
gLikDY9bJ1hVQCg0libs7w4Ul7Hp4+jtsaunP/VN1v8jvgjIsnVxsfyxqJxNDq+fo3ksCsZFEsVE
Fybk9V3oYXkS1KuG57zFRIQ8gCUXqJ7LR7uwSxfGT1d0g12S2nYWR5gTsMYURs9GNx4rDZEzyI2h
PYecxEX5muXzORozGnGyrWjrputEnXbxBIZPsyOlKY+/sj+yPakgsc858NUbe0wsG6FiZebCT2np
UbGWLssxVkcpD9w0ZxA7y+HiJe0JHrmC+6zUMFmqH+RKrW6VRwk/kj4Xw6fdH0DurgKq9tAdRUFv
+8wlnESHGrbTbkKpWOy0fxF0F8tFY8DAyoNL2mc51U683RfTbjY7PwBtG/2NdxNC5kKN6E+hvB29
6Pc17dJOYiGRaXDhM0jnJeJwy3JxnC4sVRRbl0H9TLvCHoStP23XDQ+h4AgxkK5ugzuJZjKTOBX9
fM05w6KoxW5yiOBEN6wOOYk76QPTHaWD7iyHZdGf4UetNnN8S6lEo2vIaZ1V986W/SqoPpTH2zoc
8ajNa0Ye9LWVygPJ1Nd/dthjRMVx75OpV0/uMficoTPPXAopQDIJuqKmCp5eC1m9EPy4MBUpkCLf
nbE/Gbm1wOyxjRaGZ+Y0Eop0E+UBVWeNgXvZMp/rQZL9alkyGUcOPMjMT5TRjOO1Gy7g/YMrMy+7
vCDZVxbM7h+tR5TgNq+Kp/XLX9HlC8ObPpRf8I1mOwiLKTyDPzRx/5ONnBQ2oET4BrBCMju3mjWX
+bmsY89rWjxzi4lZj6BBaVwjHYohyRhn9aCT4HNJg2eVnNlzJ9ngCGaG9nVEiTjqVqJ2zRHJ/hcT
/2xtrPEK38PaiEUvWGdbfqTrXM8WhlT1FqSOYUuJxQp7DaX+mRkuKrofn9hVNwLx47OhlXDDNwz7
Kf4oata7Na1l2wSsrRVBHgCP0mga+Jjg36PUxmUrmAn9R2qJnizkNUJKHB2FMtrX/Zi2imegp5Xo
6B0rCbdLOl5zOSms/lM3grPYFr49CIMzhIBN0qLh9mxT/hCTXMUPbGSPu1D59z/F7bOPDG2iL1B0
edeFhaLnb8sk9ctyGvI5Xli6hxvs2qZPdrZgt7hdquPUM+B8bSw5YdcMqaBevutI9cLtafsUUr8O
tNQ76vCAxBHgLH0C1nlAPAGqYm+oW7z8dfPOlKwNqrL4OnCbjzgc6WnC5w/hj3/5KdPQ6oJAETwA
HpU+YNPO9IwE9alZink4MjpU3r9tzPPlJk/D0AGeuFhe0BaHWGPfBr6EpNDeAbiyYkR8u9TX/D/C
otoiX7s3fG4VBDRuOTeus4xl63WYFmq5wZ0MX1WINohVnUYLZ7eBT67N06C8pOOD8uWQAMv36ldC
aHXN7JNpfgbgwdPQOvn+DdBHM7RpkK4tBVa1coV0htDYzLuAqw6kFNPhCVesDvl5ep2gU4SGlvmF
2gv8G+Qe3x+Wj9VbXJ6JrbuXi0QQLio58Zd1YTaZLh1J2jfGj5rGrmxjXfyj65fbZAFFJn442YTG
9LyyUu1xbBYhXEU+dmTP74NMvI6hwwxPgMiYFglqdwfM3SzIKwa8V/aovwgDnzG2Ch4BxxFwd80S
Ng6Td+eC8aoA3qdLgpWFp401pWbxqctqdMlw6EaryvcJFx0v+V2mIjY9Be7XbrVmxzwLa2WHxKPO
OrKB9YZGZe3sw+8F5aQlGtCruvcMTLurCuvUgCgeiTuSGdd3IsNM21LHHzXjD+FAS1LD2fPE8PQ2
1GoVKQxAhXFkR0if0tbljUmkG2bkuexpmVZ0vZ74yRSwWPUlRt1Adn0dPHI20Bx/NrfHxNQVgw6s
dTEeplphYHyA91S6T1GznXHY3RhAMUZVCpUrb0vjKwZF5uv2PzldPAZvZI0CLzuCKTu1CzoPs31G
yt5m0QCeXDQUpMFFNMfFu9RxxGifj8wlLPuNJPAoDR6rjouPdUjVsVw2vKL/CpCLWbyMYymZVkT1
IakDEKbxKHCBQ3RqdRamy8KBbQGPJDwj2U+PByCMh6aa5jdnpR5tBKzruNbqadBWZN1fKFlvT4fv
Du5Iy+H5bewUgxPLmbSZFdpnssnfMTIRJOPDgVMRLE/f6RqRXdDVAbh+MTkWF4P/3nMNLXkf2OEP
TFqFZY9slg95sTYXkqw/r5vUxkn72+RD3XohZOp9jENhDCsAubHrKi8ygjt3eakzBQ2UdsvEQd5Y
HoW7cuBR6x+o7i+y0NKjcLo1kF2ZrkffxtylNOTha8IiYBPH1g/qVxxPmZMQG1UUs/aFDgSJ1LTi
1b1PtWzkjnxDN1Lz3cf5OahzbvErGT7eBbZdrA/FzWRw/cunDchZR0oEDfNBd1uCQjwK+csrUybI
ErGzlZnGlHT6D9QJyx/SIv+4W0ED0FtPDFTHY4D1MyktpQk3yzI72TsBPfICY9y0k0G7jNZo67im
WyGnomhUeWQ4qFaDqlJyZxb5scXaIjJZ1Imxy9f5gb+6hTDTFQ39pPJzJsLrWj5qF4E4QGpnTnCB
tH6jhyOvKw6gUYEHoyYsTyaFx7lcipKPuxN6AwkHdL8MyaW8as+Y1L/mElsG+qdcXmM7qAf1yJWs
3zhBSh2XyUkRro7L7qWDSdTRmJhJQaMWRCpmSQ8Wzl3nhivEkCR71hsnJLX1X6BPeVSn8nxH8UiN
V2PetXxVnWm2rlo9Wgja+78h06GijLT6lgEruZY2O2p8cmznMjfzf2Y0OSlE4bBA+3fqBzYPcb/a
R76HsS9s1EMjeF3SRB0s8uL3vIMl5Y8HNq73CoGdCkoL5Q5v0+CytjHs6PXJ1qbLvRXVAZNd0JZh
IXnFcdRJnEnyJ8cyG0m3ru5FzH4u2AIpBSqEKgxE6m3WuWnLZ59dEtnmhJDh8EUH7d9tSCZKjP6Q
tm2C73S2wnHom7sr0WtF1eHkSyP5eRtkd9y8ymUYmxcC8wtia6G73Od+V//ML5s6E/rOdExkqsa/
3P9FlJUiev622AZSL9SZJyRE4BzDGuSQV3J2ZiFjAjgT9+hIYh2XC4Z0Segn608+9m9bQwzjH9V1
MowlE0iY9PoUqETsfhsIYmP8XJvSmjs+OdcIMOY8c04UxE7tn0skjo7b/7FZtE5NPIc4eO4EyDI8
vLvZojsJkx9WJU8JhOC+yPdz+npZVGYdr9Moz/M6Qehj5qNCzIjA2t9lmZH7I7gm/X8rR9urlFpy
q+g0Jc0+1BwpZssJvJj1c9dfVwgDgNhgK5DeXbFYgFu7T6rlZoaB0xGXmfcT8tDSzmQfaivlyn7j
XQypFLGVW2LzqyyyeFVCCGNwjqLqRnygxZAUOAexBiyObLoIhBntw2obt+n5AgLJzu+PFJRUygJl
Sxxz4LYnBUD5Xnm9gP9o86CLU3AXN9+RH3yxMS+YYddzQ10XQ8dVrbpaAIrDcYAk8MJIWV8DFPdS
/988oKtMLXADrBfOsG1M3cQ5LHoI6wKyf+5F5bWaIwRQqZcF3YhFucq7tJn5SxCVkOLlooOPRN54
Pa7lTOWLcYP7K0gTOnrwGqJa2w7PxL2TyXAy9vucBHnGCPYKEZnr63wEeYtd/WBQTJ6H8HsvsYGC
/5g9Xi9wA1scHDb+t6/1wlaUD21EcEptb97mP5vFgpcxKf4DZPuw+yHyd6tcxO9vumImRttaJuaC
DkGj+Kn5hEFLwe6BX4so5QuvXwwPzU9IZeSRodHxLfg06Wbciq4+lDwgfgOBIu3YBbwZblzSvIFW
Y80hXvVWiFYxmXciY2UHC+anFrfgxyjVmT0m6tbJNWayPfzbojyRonRiFuKlK69epc0z43/huYCu
Jks7G2JksQBN8OUA6S5XtCa/M2qeA4rBEws3SN7k3Fob2BZ1LdCwBupfpePWkhic0WkmYj5dfCLZ
bChusjYwVTq+Tu0DZYSa/QjbAWadwnSsmYCTc3/P17nqLIlpnip2OOmZg8NLHzxBvjH8So2Qx6YT
7/xwO8OQq+Pgo/4XmXmee7tXYo0dSmOqkWcnA2D7eOeTPn9nIOn/xj1c1W3ENwNuB6+WbpxVrKga
RrcoGllNvg0ngSNyI0UsDGLnhkKrjIV64xpvDFqmkgjNS0kAZFl0ykOLv+65jVXhBltDvQBTa5lz
Zn75wxsAcZE5E2FgpHNyGNkRxDhe274b9HB3TncBtWMtRVV0U0IywbJ3t0IkueSQpHcgLg5wlkS6
hm4BElncP3QmW9+VuO8oEFiUtx2cfLhkTR1BimbEDa6t4lKk0J8L+EXYfFRLtxfd1Q5g50gRUsnP
fNTwGudqCQWPhkXWcP5oG+8UX1wCDNpWAgIbxzZ/BaizGGbXy3VzSMGavEQOng3V9fDmZGYKspSG
fkhCOcTLQwDWfm+dT28O4KDwAYQ0DEzIta5EC2kLp0F5sVbQ6T76kD4hVT9fORptScZZfRap3rdI
hv7ui2Lkqd2fi84OzQbGhxDb9E+Y2qaEz8Gfhta+5KsZZG3UfviyIxqgGS0urEpeo1etlovPkfc+
kCoJXuKvJtauG7/WVYFP6yYeQBYU41Gj/GmlbVaOS7wUb+jpNDLje0GCJU49oBn9lJkOIzf8aebB
aHfK1rbwCcTFux3aE+hE5ReZFhXAQSq7qwhUWwQZ9x7BvcRPYzxLZ+sZcInt8taCHENHurLxDFSR
S1qokEdbWXW8occJ2+lEH3B4UJ21kmLaoKRvsT8MKf9bYxLhPJx2zQXRVbbkHh+xQve5Sv+kKIoW
yeVxVyM3A19ZeEIx7jpdFgqxioGIV0J8XpQs+dk/4t4R+icbKqaWnayEITeA9gHayBnd2LHbjo+1
aRgM8Tnv++jE+0x4rF+Ci+WHvKnUo1Gvw5TX8yulc/0YiWqxOYCKdlFJFmootsiHPG3sCjzrotUY
9mfyT+MRintVm8sEqrRYBfgRJQuSb5AUFuLYoZN6WJEsHfT8vI+mDH7t9HXSSeQlJQzW+ne3b555
ow3f79MJXxqqRpwVcsiCLwcfLdPWuGvbry+qw47nKcJUK/7Tnx+fR66IoCsSoqxs58gspxbNShEA
pRBGY8hplic1lFjFseMwn+94T36vG6V4HDWNYa/qiRSR0ownljXzLXK7ge40s7AOlEfNu8vThDqW
UjA3kZNxC/yt7g3L6nXcc+hu++oq5OCh9RzYnIa+wJ0Y+T+oYQvIX5NWUC6L9lLDZ28jF1oWA5K3
FyiCD0BL4AYUEWKd4L0GG4uuUaw6W5keaZnbAZhCouJeV50kNsRxNiyJeZva2ZmfihHxaEdqbaZQ
AyxJJenW9YqUz4fd9FHgMd3rn/FmVnd696UapOGdUUkl6FFTp0qUAofyJ+q/4vBLsLOPf7pMo+WS
vEH/BNAeX+Jm6hJ8P4TgA1pxe8posHlae4yX9wvA5gXQNVxKrP1ibk1ugvfErJKbKuMOdrbu5SMA
1kpB1mHYubOXWiw2cmZC1Y7nZi+QJ5RlNmD/yIAno9RR1JzyXQFEuBmwVV3IGK9B3LBpn97utgXE
o1m9dty+ukyrcsbXcnRw3voBXftYPQzqcBzT0fv+kCSSTDoNDCIkqkWrZeV/nkQx2O1mYpE5W8Y9
SGXjZT1SS+U5nQ7OmKXHOxVxaxiH7BuIG/RO5xkjDygT72OzOw48xmdDIsQQYAzpexKIUyqveTVx
8FYKuSUoKG+zfQD9bP6fIdfXMu/+ojeYXuEVBs9mwFJt9tZ48hzta8WSf4m2EIrwjSFdK+/6vrZv
bnw27gf9by2wl1tyE6Zb0MYE/Do7vFWKdpoKsTDC8A+GkVBXQmje/EE2bmqjgRD3z5+N1/RlEGZX
voJwNqbI1FKodUVmP9kyO3CpC1eXR463YwH93fIAHgoQHEUSWlf2xcb1FULQCb6GMDvy5Ww0bwPn
pPxUFRYsg4/drrGPLeIYdbWYRx5J2HUqBZpoYvZ9zh9c9B/z6yW9/WmWipCmFw1Nh20EDA11Ckum
Ti04pE1qIO1zLwKV9KYoWVshglhYO8L8qpUbRHoCrSffpMouZy23xmJVKi5yk0YDamisl38x9/5a
sVd05s5RZjzIgV/laUMU5GND8Vz8ByJVH8vZCeI3CWJ9COjwQoQNWMXD0gUzIOz/i+8cPaDduuI1
FMkf047OnpSOInCzVInnKWxPGlWCJA1s/LLhCP+NTSU6QRuTO27jrt+PI9pJqKshq4on1VFBbejv
kv44IQN9jTT0XpZ98aJHD2A7SIhiI3+6bYZgmc5wwTIe9wNRSMu7mmTvbBY45P6xSRZJ5p/DWHqN
+ftJEYzYWI0lTweIDvKGCqMEBcDVMPHPxNpp8zG0Cl4hJOAuVLyxTbzVNNqQUPCeXET1D2uU11p8
h5KVs8g1LviLBXI1c6q+lOayIlSEsiRNlYL5xAlPm2QHbnnmwRpAi/hTVg0YFkIHUrrDqumeF11p
RjAio0u3YQXxLf5gyIcFwY7CbzGGraQwurT3T27C+b+1DpfKOtCl35ODiTw14y4Ae5KWSOY9J7m6
ntgtlfnAh46cnjNsPCoVpfEubjSBI63pbK8F71A1UjfEwXSTrYxijgoa+rDtj9PJvX596WR8814K
VfGC0LvJOmz7R3B0K/cejQJ+8CyR4x3uBAUwRKb/3aQK6O3fEgUu8SW6tuWluMPHh/b2V6ZWkDEO
6FkvZ6ye0uDMQ/ect7ZHk+ZJ6wIUvW+vOtu2dSJ/LKD3enzmPrj5QKtKo5YatI5ZoiFFLHPjQq+a
IH0BOJKlIilGbUvnhNuT9zIRsNdvJJtPJ+dbyeDkbE6uzxhd4oJXkvHrYUYaROyi0XNouEmm5zyD
6lboKLxfx/0rXGFhoC/HIdA0cn8GzkTcrVNWdF9ZdkSIK9eAjKZEcg52sSFJ+F8Yb05N6LcG2Ktt
QUj17FvvlnihUwZgErPxPWzNNr+G/8Oescl6sfraJ5JhWnp4cWrNF5zXbwnXjwKZDijE4/1H4EXZ
Ycugpib6jgui0HD9/VTSlFfXhJOZ6VK6DJBxjyHcxarl4vqnkweU2YRb4rnxM7Su32/ADFGOIJ1K
lkoG49v7CUCvh6ecvcOEG5vyRBlcOjulWFIXINAMft2xWMKMvCG8RoWQxHjdYrKQq8vsVFSX5CY5
qcyvljSTHzATGg/O8CvnO1Gmj8ee8dM8qnnCI5xX5EGnaEq8zoKVNPMu7nhrRbi3UzCu8nuz7ttP
kqt6KfX8oUQ30mNWqCWkAgBMj48DSVgn9flOlubPvXhv9spSbVnrwT/pymebnoIsr3AeSqPIp1oL
2MGXOEacW79JvePEnL6BF6bx+tWJAn6JeVTYAXKaRIP3P1R0yr8iJXE61BaB08JXIr4GlJ/X98fX
5KcInJenVYIv2GA+4Z4yT3YDL/PsfbW7GkhCh3b6vtVCoyICPIlTH+CK+1g4TMPxj9e6NOy6s1OV
Z9liwUc17mOZLXwZvXZ0TeMqCBGt0VJEPA7OrNDrcC8q7gEsdjX3pfX/XEqlP2JFLC+XFgc8VfBe
mN5ppG/UB5mnWjQFIifWTHFaqHyQimxMbz7TSFbLh2oHIFonb/Qw3mcEB2K+TH2Q75JrR8ov3jd/
qV4PDcjEd9uMMBWWB0+vyK3WJ/R4mK2jTyeYkSJIW7nYc1UBwGQIE2q1xrsOupsaeStD/g+5ZFIA
WjzgdoZlszJ9k3HToxgOqi0Z+bI69aPGgAlzjz47hhL2bJHIGBgvfLt30iqj+wK7qrzHU2+GZE/A
rYnt3MYuhOjSQzJM5ysZDpIRb8dDuKYxsgXiL4vB+L+ryW2CaXfffCf4DR8Ga1J6yvT3epZnKzdU
CwHGQJJ2zDvknD4DOde1PbjgL3wnl9DT7wSp0anYcFF8bvDWaxqSphq4Rmdz5v4Tt7NR//79S6t/
iA7w9LKtfQcqVnMOif1xeWZe3jPuSQlDtggoRYs2d9QWNFZ/Vp02RGOm+GC9x/HnY1//oLXGRCAf
BsQ9Ss9/21ThVZ/QLAhq3KBzs1b7RG7cat6sIcvaEu9PKHSxR1evAwM9WHY1bsFzx6YAsAev38h8
lu9tmSaAPfEKGY6WDWeFrSrA/7P+VeK8M/1nJnCz7hYMU/yZo8YFRie8xxbmJh3DBHfUzLV8sVR9
MVPZRMtY+W1sbvjw0vhQCSA6ds0qd4OZxJJeO+xKl3YRAialQnw91ZalEgibNkFcmiLz75hC5L2H
diKGvjoMB/LlumH0yWCQaQQSSIOwcDogNmMiXmebmrhsrBys6ble40EPr13HaZ5Rg136dqsxN53U
03XBst79K4FJFB/MS/Mk8HD5rZCLfao1hHEmt4bva6K5HakRn6HZxCY6p4uCKEUXdhQxAjR+Jqh5
O/jVdjyZOapyI9XU0M0I/WocH3caaW0n/m/9e8JDuoRd86wBgOQtGIl70Mh4oq3Xfo6pFcBDIdbV
M4B5+tPqc6/pLwOQr4MiPKgg9TzVEgUoXwHpn67bdS9eXsYQDYmE7pPs5HEZ2BSMPqsbO0VCB4ZL
0vA2rbtAY+/CPacdDCZgslIZWCew7SN/xZEM2elVndF1/scyOpYwrHXR9o1EK1tWEyHwMw4Tp65r
4qFqLuHICsHS1X8cfGKoZDsKv0vDi2lGM2zFtRi9siWnQVeV86fd0r1v4ujJ88VSl6Y9ibXKpEuV
5eX7L/TfXDnDMyaIrGGZY9WPx6aBCTmvaXR8Hm5HnsJ05WNVnaFOmZUlYWxYUEpXTItHG+PGMGEZ
42rT0zPNzo65Ep6i8XIGzxE8awjpRP+U84FCByfsUoH3jRwnEzLoZGm4gFEeIVoaHD+lVtVxI0d3
dqMJucgwrMyr7IWvbcn9sZvoYZj4Pp3bxa/ocvUDYnMFJcUWfEea4VUlNb/UUUZjDacffbhtz4MX
SzFtpzCi6C+NPZRTFzZQBnWPQTYyoEbFm2WjPF5kJQyD9orkbyxWOnUfPvZSg0aFzbSPhxPJcI6q
7ZJt4Rzw4dCr14iOzHQXqZiJNhi9Iqdq/FfnvWt55I+pvtmwW/KR4w5LD91KTJN0kChAglFE6WrN
/UU3Hm31ALOYHHXe2i8r99J9zA7nJXKECzb/r10c6uHZo+8KdFYgrvzg28bWHUD6Jcqi+H3UdRMU
mpH0SLlvp0wlEEo0kM0cg0fJuLrt/5ZBKonGIFHt1pNCxi6IFrEUHk6POHjHGOzwFpnadkLFYPPb
+bbg00WPTjtYcrxL2iVRQZdL58iYvFbzNX1x0tF97VV3Cljapxep/XrsjflkNJU2NaYHr63Cferj
RBIJ4k0sw90n+W6/CIs1OsCF6vusZPrTo7flEW82BSa748dYZiv0Ixvl/mcZdFn8Z4yGxrFb0AHM
xOFJLsfrZP1ajWsnMrR1J3GzU3NEj63sYtVCJzNXkzcZS7CYyUmAI2URMOxw1Hp5wvMgEXqx19EA
Tw7TEN0tY45MInAzHypulWhckmUJh5RmUrlhF7B+WHoMYEN87C78XNTM9rq0r3tOKe14b2QrNyeP
AZEDebQaMcIRuzmBda9ZRodkPnCQCyY6qgg/jtFAVupLdwO3MTzIg3IMUclC4a5O8ThyTdMLwEwk
Lhh9ZC4RE2zJbUjG/OhgRiKurCSYITEJO1uImAW7SGR56xSWQPM4WB+2QR3nhDf2ZM6w1liuxYFH
h2iZ9bIjlxIxEQRBoZcK9a2hmsRGYvH3qLY/uoUklKhNPdf8QCi8VYU0vdb1VFX/IgGCxa9OQ3kA
0ukZsyesyuWYJzPOjivhE9ywgoCQLhHu1tMRCfYfy+0ey3NydU8GwlMLt2omgpWV4i6bHiaHJNOE
w8exHTtg7TdjWnvoGmCPDoNVamj9OlySgbeHCM2/2TJZRzXrMlRnvcHVAk0FqnGGPBbOcXA2Fh6j
dN72+Tjp04Cj86wdrWHiESf9Ajsu99gGhkDfFeSnS1BIUStWlWsY4sI2XnAdEU9V747SGvn4xAA0
VKOP8U7I97VQeh3KOZvS+cBr+/R/XPmAfTvofFjYsg15nILHzzhNM/IZqpHw76ghz9ysulOIYrH/
BzYrOelMpsGdJ24dbe/ZPNRIuil93l67T3Osa4JSB1qS1/VyrGINvVUjo+xWW8ZprJz7voLRELTB
Yja/bMuVBPE1iiKLfM4BXFC1DrTUfFR6Ap7ghjC+1VHa09oxksSBOD5jCw7TxRhirljS4fnfuERY
fA4+Nf9TIZMw4SOEC6qS/g/K8UCvY0UehfEn75gVllP24wHjfk01orr/y34hmsZKMsJ81s/rzQp7
EJTXFHiuNXG62dQBPUcFAnel08hwx1OTyZZ+98PtzUAPTe+ezupjG61t4bTuGlitrT0yArdwXL2u
T1WPZo7dBo1d5/S/G/62MThvo74EKabQYJau4yM5YI4gqbsxPDXkAoDwAoZG7Da/cOFG4OYYAjsG
FpNoyov5gvP1HY7ovqq1ZjF4Z0OehwuEM/eCyceig+L1VpW5/wErj/1CtGF1SHBIAdl7P6JWLqiF
oMatCgosXCxPIiXdcrcNhIRZ8W1d2kSDPEYH1Ec+Bta4QeS6Ytxykr45Sg/gstjNPtvHm5ZIx4en
hJsSArcsZcG7QdH/mvDPp7LruA+QIUx14gnYmnVbCQ02dUbvjlz2l2pApzVJtmEW7Ecc4FM12AWA
QaqPBmbN4FNSfRSeyKO9KtnNoraCknip1jMi0VoRoA5Lz4BHUiyXPNRA/DF/nyS04F7vlgPAv2R0
onGbiDevMXXvg+EiydWoSuSUp9L5wbwO5ZI33WpCckUDO86rRETEw2c9lneMP2XYTPMt7V+sGjCd
ikVdzg6F50KPqncFUJEOK+s57nK07iW7Dnb327XNbzvAe8RetkG+KEWxXx5VzGYBisKMfwcRqIEZ
BCffnlAxop7is7rcJZUJ9DNavDTayM0s4UydTwkiFYcIdswejc3HmB3s803C4F6g+EGltHm8yS/7
lt+SzudUxowXg3Yo+zy+SqACWeBf5tFpCAGrohsEw2MuO0RJf6jL/esPzjGTsJKSZpJo/72+CTMB
NybogzGTIoh9tw1Zo6ZewUP3wQv4IOEe0h8vfGNvWncXefsL6MSbnBmfRs4vvhaisrk3ft0PgBUV
OdWna9igzpmrbcFjlf1uwK1Lm8G9KaKBzMbmuxMTqjYQjP6lBh0JNC5uSKI5y71BlQqJmW+Az+IJ
1idIFfXzRq56ou+aAQpS6zeZF7jYn2Y6RDh2EbF5DkR5gF5advndFG8t2PXDrI4HS7SuRs7Lsrly
NNXPqfNxDchYAyIfDQjAy9PQsDeoozvLYUFzl3k3o6F+VG27FISv/u2t0ezwNii4suN5oXlbXC1F
JBWJ1wM+1G8pM6EZiVhiA4Nj6Ee3Jc2VUDPnqgGagLIRitKyvbSNc636oA7J4BAlaGiYYCWaH7wZ
65cs+C/Kuvzj9Ma/MZOsOQGOl+c9AlGNug9blXLk4EuPdtiGaEURsQ1NgdYG0RVytNiM5a3Sjapf
Dg8OP89m3gM4JAUeXRt75SI7uoxtiCnTjvAa+1q5U1jUd7aGrxo0R53hbDZ8BJ1XOfZsOoM1zAUX
Zfy6rNDDgQnlTlM0BnAbu+tonKTT3W8sMH8gIS6eko/bdGb2wOQF0hLd7/R+26xsRaFlLFdBzp6P
nmnkpnLQy9CdDztQ2lXc+g/SLcque8+R2kngM8yPSv/d9ZR43azuqDACehWw7JfHN3in40xqaAK9
RIii9AlzwnxZE6Ka5kyWZPNdNlEdIeW06ARBSvv05hdZITkPxwyYaCesjZ3NZ0hoC+G9clvzoDxa
Onfbp+ap0RAdjUQB8UrwduFx7G0UT8W/oDESAcyC+HdZnuEygr/3tVzUKF0UCkJLWsI6ODX0HcBh
z8G9olCZlC/ZoJrTBBOCmX7+UMpoVCvQsy9n39rk/727N0QNlGgrjBL7TTJ/9uYI4MAul4BlvFUB
+I2rnaVkheHxbAeDFCsc5OOjwtydZ+KTfKeVJW4zgARBKEAAPTK+xzKsP5yCWwbepYlcf27rHk23
GAi+bLUCzBlNd6L/zt42LMm//DeOURf3yfn6KHPfy47FODiWo5UPgKq573OkW2bKZz2nE2g3+kfu
Ucw43cHVoPg8vdA8Ywk+4oOjosCmb4Mpi2jkOHPceID/2Lr5ZEIhIU0JLjdjtmbmfZaqKj6Kuk/C
8wcyIylPewWZ2VQS+6AdWM/9QJ8FgPQ4xqGPWUF+C2SHE2+2wJLQEzZtsGchvqgX+Pi5PKeQV7HW
dEO0h7cT6ApGlePUC5l/58lG+NX02MCR7L7b1UWDDigWPLadix0TyjAFmPCGPjeMC4HRPF07cyn4
KilSgVHLHlZ9vwbQb4HShQyCJq0pLrC0DXOnnqrIxDb0ZVDNCHsyz6oh50Q/b2bm+j2+Od3jWgAO
T6JfgkfXSlqnkrqZZjEKFoPMZzkASWkBL5/vJ3MJ7OtYiW6YJPfyoxgRErDpTenDAX05r5g4WWs7
5BXhbBHNI9caM4LUvm//8NB7qu7IiObnfnT1vDuaqu3Dak0sdB0Spoo1lOB4XX0lHmuZD403qERl
1MAtvJnTDfRs6Y5zjBWfYaGTIS1OnyhY6Ae40bLeyXSXVitIYh61Yp3FYbjAyetTgbaINg2K3S48
5eSkoPv0w8qQw+xD8jIbe4i9y8cJAWeOgSQo0HQifNMkTmgG4AFoO680erf1Fr9ecUzBU7SuK/ML
dWhaA2IuN2Z9sz0y/iz20n+7Oar4Za68Puf5BwvMIxNn1oL5rE/qecJrMIBvg7VzJ5ezgHyxpdOv
aDp4B4f65TooIM040jJo1QzV+y3TMqKMN7udUjGmZ2ukejD5q/Ut6il0GIa9ix1yIJf+dTt29ssT
4BRF1KNJJNiluDCOPTTIizyUwgIAbVTQK5ysnKqs1yJwts323gkpROOyZkEC7fo6aOBalt/9kwxo
lxhV9m+C8ft1wyis5oBf74bOgNgGkHP1ISJ3+hjDAF3gZeX2+FXFAZ4JX+vwq2kEGy7swjfigh7l
J21BtC5SgPpl9vxLluKbIR/y2yvO+Pk5u99GQS49pDjB8ja0riu/ez1lReHJcGbYdPlY29ZMY3xc
amRuPsTx95rd5v6JXZO7/raoNvTtW6GxefMN70897MfwH1LKl33MC0K+XIxTzHOH0qJu7uja9Dc2
Smax6Pq7Vj7xMPVBOrEZHkJUzcGmBUtGsc3BSlxMG9CtNsXCxiivclNh5RRK6jjv3LJT9e/gw4Nt
auf7d/z5Zvu84wHUht/mqYa54HCv4DxTD9DT6nmhqaIfmNYWzExjjYc0vKZBETYcMt7UQfYmsIcu
iTmxtG0MM5f/J1IXXXWroxQOwuq8ERCoE9xmt9bIA2F1uN4yyhYwg1wJFezyNswQTJoDis43YOVa
2BAkzJiY9IeYlh7Qpg7lAaS5RBpS0SB2lxO/3ujQu9TNoF3wrZ/NUBHjYFbf41d1gLjwOm8wUV+V
Z/pvS5GBDVGRNcpgVCNEd2orTrgR/hXUXyYL57Ta3TUyChesvVPSdRNYKkvp1xwC+xE0NWTE2SuN
f6yqUPJnTRakcvvOvs2s+lzlD1nGezh8N2WHeUN14Xb7f8F/szn1aamiCz0ADpdDWDS2rcQ3rzfe
+L2sfW+9sOsxjCo9fYrW1BNWbbdGzSTsjJ9FFmXl5xWBUqcyJeQRXgmZMAWYeCEbfVk0Nukuro9g
0WSvzFI7onCfrVKMYqu/JbqTL5vSJ6/L2y8xTdfDgGaJ/NMyLGXztg7UrLYM8QyBCLQSg3rx8w1h
wkGVRnxpTlDaYD+E04EW/MI+VTvXZQMYtlEpD1nFeuk948F1Xy+N0zwNekrZxACkhQtguxF21zFa
JtBZcu6FFXikAbYX4MxunnjCBxirie3WM+P4OB358J/3Yd/9OmGFkF6jVt9AE7oB0hbpZG0t3utx
iLALz1XlazFY5hdMXFk1F/13ZXtgPmkXFJY7kjmczI2Nwqd9qERuerkBBh/P0sqND6T1Byu8YTSK
hJwlMIKkUzNX7vVUnPEyg7l6hCcVMbqwbA+CvMRchkRauoioivK5d3l1RvaUZ82CMpYki4JWS3Jr
XV0GJtqodwGPFiCJNKLl3j+dJJC98BWZRyjMIir2O1TTo7Dsqjm4Gz+X1LeXzfQ1bxDvsMTL7iXg
wkzifCr6dti6rCj88SAAMziXRqEK1aImHVzbrt43f+dVCGqkJt4u+X52HSI3IZ34QP68nJNzc/gY
2iEZ8zszFHk9oyHwIpiqYbVQaWmJekM0KQ4RNTt6ugL5OXkGaCsEv8q9nRdLhryxRfky5WCNbCb+
xHbYm7PYB9sltuRdL4eClqLI9wuNgrRfUpXID9yAoR4t5W91lkRI8NfOZsTzfJ3oKrAYLH/L3bPl
DZv3OjNswHFUkGThv8S5q39IoQni0OjEBr9rBwnYhHUnmUn2SWv4R9LQ6mpVMRvjhPSf9jj9bupe
lkTb1UifdatFERM9Pv/PUSAlnXAGxYNGYneAeRua0aKJwvfPfRboPZsRLth3skerNiJkp8GB3M8F
PUpl9H9HeOnB2aKbueCzDdoTTYo6+K1EtE6II4SNBMrqjj2rEB0ci5Yv/C0JYd5vNWZnet055Li+
GSA/nApqrDtSGU3+selTNtXHRRMC1pLMBBBpd0Khn0UxnX5fhwf8DhkP4r78TLQ/88wUmyHsJ3XK
CocmYeKHm6y5mWaRYz8G2tKki4vqU2b8pCno13u/XTEw0t0yMuIHZ8EOt8XYoljKu5seO/otTgHi
AisWCwfdowRys3CvU3XHMs18oeDx5mmFbcrNb9IsBc1b6mFs6K3Cfk0z/vRJLhsBcp7GjJ8jl8NR
NRQZ8roQRekXmI3tBtKxohAhmUM/UpyDMgQb3wEYtb+zGayf/ywqfR6x6eaLi6eOuHCuKs/SG5DJ
m5c0GfIxu9UZZE6jpJwKtEIcakjrsvW9H0XqgE4bRyk6kt0zw8G0JFUT6r9uTQgb9toad+wzXr0K
YqgvFnxIB8iazjasCRHoj+znEwvSMwMtK2ziBgfrDoDF3hSaYUfqo8SXg/6zjQxHty9MTHBVlADJ
MLNVpMSgpMFUqELLjQbSKvc7oG2cAsHRH+iIOs2fTUhX96kfw+lu8ykipQbPaX//QWPmMo6EvRkv
TCBFGwDB9IGWTF8l+KmrEunIpHC9pMzyDL9wCS5zMlIqVefVqDXHufnuQylkywjnQltpTQpBrCYQ
8jgEFvWN9QCHBVnmy/vF5SYo5XIIsDlRKec+ZDu5yN19NywJ6VjOVyXYJHw11W+eX5MddHLxpk0u
gzanDHnkV20QMhBJZqvOG83Qp3Aq9J6UW2+hhUYsgBYRQgdhBgwW5iIVleTIAu+D6Mqp5Rx+Ni9A
pC8TEnFkV/SkIl86uEwZ2xWbInejoXw4YR9A2WJbprL3j7U72KsVnNvlMbQecTg5FF35yxeIzd6n
fgSmVrT+SQdY5cMGb0XhM+1sSFS0Aj5hLQ2O5gNvJaOWq4UsXwNDVt0PCdqrKS0cTyaLp3PsUOAg
/sCYqg7idJW7+LiymoKlGbbZ84K08eZhzzpIuvCzUCZLihka0mu/eGwH8aVLC5o0LSeB9IvjeELX
XvryMcC3tNlkgQ5M/AUfUdwOooYHHhypLb55axnPfIl6m4MlKbhiLFQda2IZlDeAoXs+itjBHXCj
PdKdWI6SeMaqwtzN6XyPySCczij7PCiKu3vmab2CfM8KGyfPNPd3SdhFwQ+Wah8wZ2zDcbDEdLc9
uwvziIh5cTpOQt/CHZQ5WMcBGiPNm8Xu4EPdGnpEg2thlTZBUd+4l1QqyGUnEhyKywHhd0fJ6A9e
BbR87g4Waa3woXIEyKHfco2UuCkKmU4vZcBLTE9IRrmevJoMtsNSe25SJx8V72E6hoFkXocngWpN
glqJUc4JcKLuh8RF9wzEmq7n4ir3RgT1UzbPj7BbzwHc/fwCmHR5zWMqtZrztJUzj959FUJbIez4
8891Q2TqCNZnbTuMyq+44ZIrkXm0/G2RE3bh5P1Bqgknq52nwKJHEA88HAO4hagDyLOzIJzCdsdk
AT3kf+GEpFrYLc1DZHYHHYbdYG1GN2t/k4W4ewwr3H8H/2IQpiFN8yY6oEroTHRH5fkISH3GnwTl
io8Q52dEds7sWNBcwdWPf/Yi1IKSCmjbdTw3KrzhgU/JHYkpYV8fIZr1bqp93sRy/OnQRfjC8kCv
EErGvBsr/i6mjdlakpScw7J5G6OhfG5sse1fqscK/wQ/snLhi2W1ns5CI3YHpm1etemVsDge0fKn
ijKqG4IVs+R/7rxpH+uQFhuVF3P3dJJtny7RfgQOXvr3PBVm+ZoFslyDrnRfbpvxT0xf7mejC569
2ar1p4bMcgwDfeDparj1RossAldRH2Tb74sTfPRiVjfGzL1eyub2qkx3JCNi704pb9anN7Hu8ufJ
beW1o9InKdqRvltXfy7BanA89oydhNyc0kLx9jEXWn/5Wy5J0uoFc7wVLcTWCVTmLx6jEQsiYspv
8tgJvvXj5nhF4I9VEA4BtRyesK3QRi+DdzsTz/dPOZRwEQAySy3Wnvs8/Z4gyj37ztak5CAjeK0v
atLH+IoPHrYexdtuNfws+nhstnvVunWYNKCOeVdXsCS/MQ8HrpvVtSdMvy/XU3+h7RSebn//NV6A
Q4IubW+qCy0mJb/kjXQIWUFd+E6rZ1j/vHaMeaCyl7J+37YIpCGuj8tu2pYsfxORJykkdvtUaXob
0pPRIsbSIngv5RVGosdF4eWsUiU8yWRpZD3gvVBtTc58v69B2gVZe/9/cLhKKToO+W9EhO2sFYa8
L0zX705xVIOUDJZIFzRJkbC9DKYk5oNRszke9cmIZA2/5SRFPY2trHWlzwA52Tu0T4+INJHy4j/D
psXSnGU7Ni1rEp0Gi9Wc/PAFuBQnxa/2Ov3pJanWHP1bWQF1sVfy1h1+ROT2V+Oqc8xOFI+AeBLs
DTlAOD17lXPL7oRMHnMX1SWNuzJPhfmeUm6v0U1pyVRuyzZB0Peg+T7uOA1o5ondSb2Q5dNOD61Y
kA8K3G38PbxeUvLUXVKw4ZubHxyvrOUsO+DvAwIae2oI1Ew7VQlyJMfi94Ciyrr+Rq8LmHGSpEd0
ckxHB6mnRI3OeAlMItQbGzigDmaLuj5IWMEYYMQlhEJXovmtu69wfY1rnTxUwyRNcVYQ8WAh8WII
U+icaBwUoIf7x1DMjJLrhcUCWX9FSN2yF/kTvrRekOJ8zTiquDQUYUy0ZzvhLb8zEhXauTsdJ6BG
PmAmuCpbXh4qGxMSCZMDN2bbE8GnVt/O87rkEx6Z5H2pddKCQuALk6jxb5GC4jZofsQRXYXoHZgo
ReTfU4par3Eib4TgxwMwUgZYRf88wYT60EQCqKAYOL8VmfQrbf3aiI1C9Na7qEf/l2K9M7cmWKKW
JMH53iD3fgkP3Ua93XOeyPp+H9WLCrhJY+YcsdFn6es1K7+JW826ZlolqFUd1VcwQnMdknSgCS3G
q/JkxJ0y18OW3JHNhAuimw/8d72wx4yd/V1aweFQ96dhjD1F4ynb3gYNtIK85gjlsX1g0eoYxXvs
WGfmuvoc/CgcyauvE8Hf1kXnFTRNi+mt8DZIY5Jywt8HVCcdlCQe0ogKVa1HHOgqbFEAHoJ1EBEH
lVOX56eA7WXZoBrOm9WvAHMlOnsbceaxwel8NHGfqQ+NfXED5NlY2sS/E+4PFz8jgeZjUdruE5PF
PGYRudLHFpJlDQihDrk7YVD2ba2XVsIW9IFPj0Zv/OqEcWxBiy4vMswYiSEQ6C+94HosMj/F/HJM
i8ctLfKY964PEbysEqzbnJDsiot5vunqJrCAJDHsqWnKwhaQh19eT/HF0PWSEvkwfRG2hrvv4Bvh
PHsH9FqYLdwzK27CxdA7QHF+ha6Y4eIqpgny+lg23yRwwoudVhEfBYAQBskY4zGK/CaQ6w3pbe2h
nL57A5wLX+bb5zmNatxVVHKgskcEo0+XP6+sI30FC+XBN2EM3f1k+99hyEcxPv1ciQPi+Lwjdmcq
9mQKepAP3PQM5Aj0NvL58+HRq0+1LNzBikjqNU2W9sogbNSjKzUyrUmGs7XIjDzq2JD+gB8324f0
KQvnRCnVPV/P22DPxHBlbDIPK+3T0dsjG2zNccD6rZTnLe/UBkatk3XeURG1AF/Fxf4Om3fknE9C
Aty5OGEsyzLp8eg42A5pFoHnBN24vhmYzspgUeuNN+hlIayOpCgzcCtjj2Z/Ws8HSW0hmaJuUWMt
V1/zzDq4anFTSUx5IzYAO2iVFDSVLu64UIqFKUBsMx/qqVPdKjdJOtLH9Wz8nV2i2uV9ycizK0tA
Brutqra3E9RwOvyKtqgd9z+A3tiUeiBp3NVEH9SvzDsHMUFD7YXQTtJrHFxjJvNq22VzH2TuVBpY
nn4mlGKZ4rDruRgxg9yLyB5TfYrt44i5OtYKnpZP6oZ55ctQm14za7h3cUrC1p80OLoouiqnuAsI
YG5ubdemYGZICz9fPkuGqF8gKxeYXzcnI4qLJiKPJ144Cwds4IBFkbHBtSB+E6uHSvEPHFEf8+hW
y2B8ygLtXDJK/WPj6WNypYBo1BikoCAy/yY0cORtcA6XSrMkXdDF/Q9HKo9iSsdOhwd3mn5e0SBt
VgBZKB9Gol8qgl+gsgHv0u1DT4TNPNShCckYpfPJcpdz2xusk6yePbbWFW0yt3Bd+PPFaL6iuolf
8GSElg6sAjtsyzcvEZ40ZLA090gFRfCLT8uYsDMHVESoI3NAi/6HKtp/cSq5OKApjnDzc1NwmFcd
lV8KehVH+E1rCpgaFhvBvEeMXcf6ntWOtbra/TO5sA/Y1GrO6b78ilqSjQgaHbLX8iCn+lsN7Qzu
ahwK9INExjZOPW5nF//ZgEcnC7SMs/z8JiCcV8g4cZrDNG+MQCOJaprWsvafsbdT7azCZFqe6Vcf
va7+60zHZQusY3YHsuA9B+oyQKpQpvbR3lAcsmZAWZf6kfgFqS0a7MYfcc1mRNuJYQE5UmxJnaUI
b/f9Rfv1UV8/QMhznyyUO2d4hJxgSmzT43QZd7cugKzpea140oQcl77oPEmPT5EpY1gmVn3fsWa+
tx4kQZzrvQPPH540wUub+4R/Jgg+sGZdr7eCQgissw45dOb7oltNesY61p9qiUTPQ2eCkm56EFrz
knQks2Wx+busjSj04k+zNwgbALlVgfW1Z2luJdhMUCQB+Um3+mIVAe/hhesMVchV0uvmR81TgQHy
0FjgQm6niZaXc0/Ru3RdnJShwI41QXnFLpfPF2Z+g83MAoZplo6lbnczgT/jk0fo1Ai46HKOmHdr
zqiZ8NXavFtVHKYEQWCD7j3u+vfamm+AGtOZLfuxcSy19PY/K28noB5xt1HibfX570gtsub1GUtk
qfN4V7jcx38gfej+2pwLbRFb0ZQY+M4MHWwjiUxsUTlYdR3tTwKcak/c0dDH3Jr/YLAJhfh2PuvF
mL6F/gSlCBloquVmf7alQ7MAgUCa0uf8QsBXt8SmUK4cx5aYngW80Kepf/o0fWHiFjXftghoFjI6
TzyxY7sKSJle1tlHa1RbDR++am+y7DojhDcRA4+N88pwbXZsieWrZpZR443uUeJdJavB08tqiFWQ
bLVb0Z+UwJopnmmRnqDlbDYRAAXfd3y7O43KKX50DkXgbgpLP8bg1l41dmyr/KXCHTodNH1iuyMd
rHiE0UEH3LA6kCUad5bkcp1nIiRcfrEIAqHxtrWpZanScT8KC8+hNhdddqSUZZvEXm9PiMzEeAvP
kuFXgtVs46RoKg5c5YLeiDzQNHTS0mbzb4DLePknW6KFF1kmsHGQhwXFnxOuVxm+SGdtuJcZzYn6
FwX8ModTaDeVFkAhb+dzY6RcnQyQBaY2RTauYFiuIGP8NP9Gu/t0LZpUeDBtfyw1jl1i5JHK8lEA
Sk9iyfm5R+vKlIDKg2RxDd6o/6E9mM0gp7hyPjB//TXzPAKMgCUTpHBRaGEpdT9UYDW28gVe1Gax
/d/6YXgt66AJwg8iJ7wao2vn3NCAdQUib8po6t4VNpNklaDjzsaP81T73cuCWpT6Fptk17XohS7c
8THCDDD/49VZmEf0+sB186o0Yin7BshHhycE6vhQ8+Nr5+194aVmXTLqzN7FqKOGJSi8vgO++0qK
ak+lciePNYqP8LVrxLhki6H7ngH1x5QXxr+S3Iqbi+y84erkEuJ87opA3KzIu03HJL8ZK6X4Q7Lt
9xlHxCTCpgFqFpbFVn4/K0Hs33yr27R/j31iER3PU1DUpT3bk130ikeY+K68AE3P3s8HuZUBdMRA
KOtdryj/WQJ1Ekn7ODTGePnuOboqnvPgmhtNV1RwjovTW6n7qQtR7h6Uw1hzEYZtJzlXlaLdd3Re
JEebvM4BbYXyU2IzTujdXRSXwpl1/QniRDOptUBgrBj1Zybv11Lrrwu043Tl0iNob2ggkspLVlb1
/NpYv1BO+WnGVZ7bBi5HhscV75PkXvzA2KouSCGJP9vIGaH2uwqUTYEjqiRD6YdAUOz8NHzX8YAG
pLq43ueOpKiTIzZzyO6sBY9WnLmcvZHRqIM51z/IusLt7e+OSQb3xrgMlFB33sGGXKXBkXkNhGy9
xEB6Wb1odp5d1XvsotZyxVJIesxspxz8D+m8k2YHG27tvD3X0yUwhlMttcEd6fWPkWOfBfglfmAm
zMksEH62OKcWbYX8n+WRwAvnuX/G1iVukzhYlSVMSVwnsbGqJY1dn9I19EC6s9LUg+9ZS+AlTEml
rvb4sm2WhWhylncC+0gV5nrmwbp8HS9RErrYrA4IZzAF91Qcy7YCd2NSVNuhn8n839Y+83Fwg5ii
xkhnt0vlAboPlbhoPoCmWoDlWlqxoEiZK3USuMTmUgEzMKgKIe5P9zxABPXBjlUHihocndQ1Mdbh
bdMZmQFxS689e7HlQb7UJiYsFAv/PcGg+SqOYTp6Q8pUth0pJr6JXDmh+js1fU6jbmxpo/saeKdk
rvWQxEIGs6LOCYNHYfLh0kj2tNgOX+Ip/5LRb+u9Sy4+l+3Fm+NUkyAh1Zf9o4nZFs0rdD/f0poX
9mbzrGifALMA+EMf5drcuNAE5vnWCIQbBdbjL9nrOSG4RliL2U8LFqs7f+Zo0DRkiaKDoCv5EwHl
ZkXHtO6J8YD4hScnq3MuDZONHIPz+3wNl1CZ6dJY8gF8ovKjOdfpY2rznPrj+paj55Fv3QLeVrTm
58O7PVi3YVZtT18P+T2U4D0ZbcHwz9mmByVucMzbDiRx9w1bSWioDavEX2pplI0V4rJfbk71KJ1S
QvuE6iaR5dduosIzBXN+taaWssh2XXwQc5fdiaokdpC5wjP4sjLrqofZoDsMPXUqfKfjuozZiXHN
2VF1D0twwu8ubMqaO3fLP8CnP9boF3tpC+3LI0rnlTAGqVmgdd4YBvkoCpd/QmDa5MoGpIpf6es9
NPfQU5QGREjkUW8kmOEpmyTff2GQkrgf4QHdkSiUM2wdkCDO1NCr+oHaEEDXf5yqpZPCOpOaQlGu
FZ2mjdrDuTT3EYZgjDcFH8R9XPRPXhoJo0fVAn7/ocf1PoDA4xAA0HbGAtDHu91NU8t7Y2FmxWvV
9gUDvxG7bjQnvqj1XBQlCt12OhfHhqWB9KH4hoEFYjo8IWu0MpfFDs7qJxt/bchHaiJBLLhj76Z2
7Dqdunc9+oBAQWPV5j3zh7wwQWWm7gZD0FbSjTvvpUPO9zrWQlNlMv0TrwlWb2voPT9dZoCx/3mz
98vhGQ87vuBUCrQbkEtqLMCOAaIe7b1gP6/NM79XidXIQBM45sC61sj3i1TK4ZqPqsT73clFxAAt
gi++Fwtt5jY8AqxllEj3BxlhEx11Fh8F27V0g1IxjyvkIMsff+QPxiTrbg0oLNkYxazkW36tZIJ/
RHHSTrzpO6bYk9MhqQ/vyh5ake+supr+V/XnII0PIXkUn5Km1aY9b5Bk/ghXDNfS9/h9erN13cTN
q4nSM/oMq6nJ1U1hBq2GdUVvtcAckhYzcTwRQYMVD76nQbmmP6Oo4muwXMyzXX6YOOW1GDmLrMY+
m+wWVNC5GfJ70TFBpRp17B7ILsbQlkGZMFpVGWTXOKjGnBtWZlIglqPajSwXYKTTRpKFdQnFdUXx
nfFryETkY71MoGFKJfZvmZbIgoqmpcYYjFSfmtEEqRyA1RN1ErSAsOtiTEnMe85lqFoMplixunOq
WwBLs6DpWX9LelHAYTsHzA3l6TzsSa5FhxNe99EAgO3dnH2fTMfYSe5tdJpalyxgGnnr7ec2UepC
cORuI+nanO78pKIBB0efqjAk2FuSgitntcvqAFSIRJwakeyLl8GWsSjKfzVobII8zT5P1NBuU94R
qEphvmiyYerUqFrsygCDj9CW7g68RpeJIRHXsJ0OpQEcpzYPoW2HBlFVtPob3B4Rv+4Q/tUyi13u
Am5B+KUoIhmH4ubNkcCD0pGopPqBGnsB9R1J2zPrIFyZcwE8WD4ZqkV16NzojbcjYn8+pavl4sh6
ZtyY2M3Zog8U/hUK6G3EFII3bJggwqpY2Ie1SJxqlBLd+dMf/z64XUUnXf2z4txEdVES+fkZ4RzN
GfVOTolSlD1TCUjT18jqMgOrkg1Vvc0m8/efXYjzItTZUpdQ+14CyRbX02M1VvGJr3wtxqCaVSMr
0VFHccGypUDv8wfi/KuGKoFQE/yL/kv98AEQA95O0e2OhxSVADfRzgAooFI0nj7c99ECc7q1AnwT
I9lYrzxohSKDFqVwNWAsygi722FpTA3wFIxVGR6M9kt7Tg0yOUiZiXSmF0i9GHmWlwE8tkgbmxPC
ToNlubwUAXT82M6/DQCjdOMyCnVevUSuyuXSq+jXZsN6VFXVcmIL2orh+lrw/W0HlvXY/vNSlKv9
sgReGjdVqizib6rqIHBb6xw2iWCtZStUYiKfkYXX4WEP0xLxOCF+EeQC6z92Il/BLvDfBbxTerBT
EXDzjwDt7ZJ06+4HkkqqpeXg2x00Z+/hIAYuZVDkamz2rcLOP6XV+EiVI39t69jYddMB3wq8U8FK
QnW8e0qQ0pXUG8DJ6wOiyoFybT5wynY3uyjGwwbKC5lbxRNapodDhcE/J/wIsR3p9pfFI/ECm9hq
ppal9gXg7PUshGCFAl7OJiJvneaq4FydkhvnAL+RZ3Y/CEw/vbuNraGp/K8geif4K2/1mL8ZPvlk
ce2boj9JGf1/wsCo2lKjEg/DllXot72v/jK0WidY8zmDQXO+xB3wbw3N4wi01lYWiw7TXQK23Kg0
8PBcjsvk0TWRs/CoBTUaQZerFcZyaQCDBcXv1P7hL8mXTr9xI/tgSog1SCkMEApsLMxkSFt9fn9D
00oNV5ccZevWfIUHH1GL2TGEQ2KMPuhpK7FLnWDS5S9sj/1eHiREVrz/oHMm3b6Q6ER0TRtY8d09
qroqqlcRM2nLnicfHrT9gE68YfxTvfc+pcU3cm7EJ83eTs4P78aFoPEOUxwJZw7+TDK5Pc1Yaw/T
aWEfwBnEavrhjFgfmP2PsmL98O/2C7PpBOUhdqfIp8GlbBUkSeoTyzDyi0ayhlZLPkqz0VmIeHnj
XfkuVy4iYnvU8F0rxv4WVi5QhlLqOM8X9bHu5NNIXi5GlaAVFmG5zO7i6oJQT0FTkgnxWVryiqJQ
6kS5//5+soepftR7JeblyiosJzwnvlvdL3+EXMlDwm4nIYEsATDR8fTLRikGA8CiKGbCzgGT1Qtn
I1L+TE6rVLNjzQ0cAM7IGz0O0xl3tibLYLfu+uG0oSGdBB+70MuKZflmPkguOZStw2JrnZa66SBL
bhnffuzCdxvvcq5899/I7GckmostaTAXhM2PCZtYUP7SD8g1xkjpCjVXZq3Ex0E7f7/VBIA8DdeY
Z4iZseoSXYKum7ik3hz4cK/2dY23PB8bBpYKwtXLuylRI7veQ+RTbSXGG1N5rcCtpI1A2XGS86Lc
xAjZOAymOcBkVxAAl6m0xaeKHTwSVlCTIkswljwKX5B3MQ25IbfFDfT4vWVDuMjac7m3EypbP8qc
1nXoxcQUbQ6ajN5n1WuSsvld7k3R5a7CRbPMRDlpiAEO30CV/VoPFL+JNNVhT5sDtW3euaG/TLVP
JaOKRmX02rfprHCrygj9XO4q3qTIgNBeBbgN4EisSl2wOWS0blE/Rp4D3Ute2qexJ2SpnvPifj3T
ijvL9WF2lZww/3ZKKVRmXTVtFwmHExjGTrhxJAiKIiDTJ9ot5+wm/vKoq0YcC5CLr0AU7cptNmaS
oyExA2X1CzZ7Gnv6eYqsYxJO7EyIX+lHuPQB9XqKtIuETgMcXnevbUZ7cq8gM41QPTPLZGGb9pz4
1ermbm1PC2I+sHfcf/cbIEF9dIQRhKMO+LpLwjKAFG0de8eGiFmQM/B3qRwkAvXzgtcw7DvcYKyM
6BBdXiy3wZzl1QR/oZd4xXb2jsETgUOjexE5oJP85HBFp8J3ZzskepiV+2LDDWF7aMnbkq7NLFjy
sXSBhmHtW7bLYq/6ZspJ0HiV1Fl9LIEUvODgf/NvaELsULNX0U+B1YuMw1hlOUB55qOGWzQ8XvnD
Zs/lpu+ocL8QFxMxWRFSSIBPoqeVX0Nb60H4lSkqgbINjI8f9LN7BpwQ4jZ/eSSUzyDowFT5ZUlK
GpUUa4zqPJpRx6n479HtsNHMwT7UWd6Z7HULJzNpe7Wx9qYJ0JlEVbUZs0r9lmuQQu9m124w359U
lZEDRgbwSOVQ83CZPqhE5MqExLUk5GbVhP48D4Wc1cVVDJQzIxKMwh75rktSn3vIh/popUHoUGUx
dMcMBBcpZO7b4c5AgWsI+N4SpFi7b07V++d3Ur2iuO/7Twt1nre72I4NybobuW6g1/uahE7jK7+O
APQloUrUdyfYA2II90mYUZ6qmBI28ARALB1eyf9lANlCm4rG/kWMSkcWZkozjxBZpcYgkIgRd5R2
xmmWLRKNL8QZipBvw3wMi1U76RoWcLO/YM9TYYrKME5wW4kriEEwUX5iyAENuS7ViM88mHYrJDvn
wBKvFQELag0SmZz1TTfUK98fwwXYlBtmcmW4FMiVrNqcy2QcpvX/nzw9ZMEzCHFu+xuAGorm0EgL
Mhvg9pmHeoVpc6nqSd80CQXz0jZ7CT4oSWf92Nt5zuwfbckDR8rxvoINrIb7lR6vE8lWNMcqcoRr
aerzDeHz/1yl2Zsz/dmWrpH5miQRFr66tLKF+LQzG6UmVcrVH2V6iPWaAiTMNOCtzOsb9KjWVNz8
Tnb7I3Iwz3EVHCH6DvSCv97ifepJU2fnR/Oywd8TBXTDPB3GTgivyKr9ga8wVXDl9eJupBUaM43g
Ydd+d3w2q/nUh69u6+CzUJMztbr9FGc30RScKDsJ5K/oP8/rX4TYbs8pvIVN48kr9yvky54qm8Gq
eIg9YvVnTZ973CxGxQ4rbf2UadjIehElIF1EJwA6NZBIicGGs8rukSvKGPtm/F5jbmXIOMYywiMI
kZnbnxb36xbH8aj3t810izi18QDbKrk/L5oNb4Wm1SHNjhCurXYQHRDNSDKJ6hlnVkxQEXtKVTtF
3Eioexeo+N3osOCwqHtr2DdVcwjx+8nWTu5KME13hFi/6IqybyQtg0kFY3TgJYu44wH0O9u/3Xbq
fpwsXXmEJ0xSIqrShn830nh7iMCJ8K8g6kOYewojTRyTj6DjZklANW3ArO35n/rJ4/IzbPjBD/R8
iDRINjA19CnysdzwGc/l2dYiVOBTd5tk5w9DDQ99h//qNCa9cIvHPue7ODz4F+H+QgleTxn2YsYH
L0SRbLt7aMBySj2rnszgmf4VC7RXqRPGmGPZ/Dg7Q2fAJ/Er0yg4CnKdywMUDmjo45vcXDick+ko
58ifRonfNMhbhC0Tz2+Hp9bViv07WlBDYaOh4LKehIfzXjOdJIDSkzd1AqnZLWfubbfRiYV6dIgE
t/U6zpcPvF895PGYhWy0f+nIwOVAUvnW5h62uduyzgyKKKyjw5mCtL2Pw6C9A1vAPSEXObv7WDHk
BzmIHhQwkGryQN/g4DUMUu5+o1stDLhFoE/4+9cffA7UEKCzJb8sFr0ixEIlEd63snkCGRyVQtWg
hvx86c/Pi8XMC8OaUmZfOQnMr31G8aqUbxau1voDYtzx2+gXutWQM8XVbTK/SMpZW8erdGQJO31f
wm3bLiKTcZ5GINT0wFIECJ2xqfoXJ3mysU1rSnqfPigc6Bnp/uokCqOwnklpxTQ2/gCeMF06DNof
7XyWDCOSlDWwT/NXRVMupkS1lLk4hClOL2k71Qzt0GTwoHFWDnPVAYeYq0ruin2SjnbUrZeR3Gcf
hCYhUiOWSsF8BE8Fs/yV1O19K+67X/8Q5L/jrEaKYxsjrLnlMZGP4WtnWp6IgT9OMH6ei2ytds8l
JYRiek/HDWkpEdD1wQ17inX9SR6vl4Cz54+4EImzdFlDIYDY+BaXm1SjJtdu/8AvVLq7rk3e5GNe
oJ/1BnV0KoqVOJUzwSpvGfn8FbUvGDPjZAMMlSHHtBXMueL4ymUlsf84bf+/7v+r6cDdFv6vkOO4
FxWWHrndPKXNrWpBLTKc0Hv/JVpQsAaKaycNdKVJfo/Ij+WnJdrU5c5yZv+BWsCVoiwerrt6XEqV
9WEOPmFuQM0L7pxMJCpt1P/GfyP/Kh0KgYr+qW152lJ9vQY3zmtUb3/0Az1qAjjQFBTOFNtSVcQv
KsUjdDHuGZaoi4V60n6Yim7s3SLXR1Xb8LDx2zyZFp4Y0IhA7dN4/KtoO3nOa9szE7gCykI7sM8E
pTeb3cslyYP5pEaUt5a0J6ZqAQbe8atyHuD/vVUs/XtKglYXWOSbBLM1W6CvQUal332BdrCVZwTD
jVyToOcFpJPksamPdz73vNw9m+ri9OmtQUAzk9kg3FoxLnqx1D4e7aL96Iixyw/3KBmyTHJGRYR9
zuMUcPnIrFsvTvtca0G/G7IMIJbJhYC2hwtCGQemRBoyvqHA+Ic448lZtlJJTMS6xc1QDQqu5hlp
OPUTRBDUi0zthf4++K/joEpjK4ZM8KGMe/DiMydD6vJte2jrZioEwHOKlXynwItODcCSMg4HMMEM
qi9KrcNaYnnvi5TOuP9Yr7/isTn515A7TVo9nnMkl2ddY6f8LYE4q1OIcgyc8kE0g+tLi+ogI8w7
AdrpdBwNAjBaDjNf1jRO1WHQjxME0ASL/H+K6cODtiwegkmMEm4/oOeu+OcPkQS9F+3HXlc0QlUw
Nm1WQRpkz9O/nMycB8A3HV09WOWKyHCCLtZeSNUuaqUmAvQNFfzExKu+Nw4cQQIhe4oetlicBtqW
QqdBlSYWBIHTApz9uVbuPzinr751mwY1H7+wPd6WhCI6BcpN8naLEVOFDRO3djM1KVZqrHBK5V4k
PsO7HXK3VceYYHGUwZizFytv7jJU30ge+ng/pQNFoKX2SrW9s+MtMuxWSpAoRRshfpZsrwsJ9IXM
NJzvXGwq8+x90Yl9gbuvTiW5k7D8RR4ErHvbf5Z1HzeLMVRfjGAcyllv6cEWH1FiHNL+mXMN7vgV
UBafIwfpuWtEYsUdYqzLNU6DmAWq8nylWy4RGLGX/ts20QB+jifxUETOrFrgIrtUxXm7kiWyITk1
JkEcJwKhlGtDxsBWhEq3wg3tCqwT9OG0KG3PX0PRFeL4fWt5o9hzIOcNFBwoRrZCA7Qj+I9wO2pk
MX59tkt0aWNx6VZv1b6l7IW9f6nnfblgkmzDeZSGEb8NzXV4bx3zGcux5ZWIRz/B2/w9XQW2LySW
1/xGtMZw9Zp64o4PoKERfw5q7CP/9/nRHs9FdYWfYKfdlmCrKNjUcW9zdQopbARUdL6yyjhD2zaY
HKN1Qkh6g3WdmUHABVfj40Yv/LPmApr591YsoWEaJgKAx4XwzBPF0SUBLjttAQTRh1sfEd3xvoIV
vqyHxQyH8vk77ky1OMPQjjRxMAX0F5ynYBzcXqc2TGXzMHzgCyoAPPaUAjciqNdWskRUNquN4TmP
GKkRfzOhe+J0T7WSvLcFtJrhXAAumQNu3xtgmu7FBvmOTDcZ0D9MRr8jbsk6cSiE7AnlE6Wu0l8u
rVbicJLFGooVhTOthw5d+7BJPiNpZrqN+r67sMITrNzFwEBNCLLzVOLaz9cBQDBHjm+rlof15bXJ
TOv86z0Gzi8UAr8yhjAOqWqf5anRrXQEw2GV6lrs/lZeET0PY3VlTL9ttY0gJSaYzBC47mpXg5ca
7a04TufGsyPmDdOY3kH9Pxp1ZvMckO4D2LVt85X03Ll7NrHFcAqFs8VgLREC8PAEHsa1pMd42a90
aijrZC2Rp2jzN3aAvJBfc3rX+AQuYNJ8OqzBtXqRQkbRI+vhommWM9d1PmCCEOqky45dA3JGQ9YD
m3RY845GcVHZPqmZMWVgfsin7sm2MvZbq+r9qi80Ham/ukInUHMqTsTf1z/3YYsnDs/oREj6Rtn5
XHOJNwI8w4gKFO5ogLMkObHAd4O6YIjSzMGucrGbqwy9UHwcPUIbnxat9L4pBb9u2IbpUxr/YTNv
rDaCPglStNyi98sWYO0kgfpjYNEhXT71J9pPwEVNnF4EC5VVsxIxkw0FK79wXYWWYAI5OaWhbtOW
Ex92J7Xqq0p1D5rnlDLIMDSgOYeF+qRYrfXanvGjumJasMMrVbtOcFWZUOzp4lBj0C2yhaIt3nQr
d0dH+2QbLF52ee9biE3P1Rx47DKhD/SplbEP0mFLmKkMPskystGWcJaAcxmk5+J/37IC0BuoUy3V
IfU/EuqyCd298deb3/hBPwLw1b9elSu3/T+/rQCjXRtZGwY8q/cweSROHQEk7VEc8QhwJ4iXR5FT
nLiTx7rqi+/K1+YRw76LHprd4V63MAaK8+JxjFeZROM2nOIFha0MpqRuzPfiTuQ1k6I2fEiEi12q
icMyNwWKmtJtzz1HDa5EMwncHdcJkVMcGFVqgnCd4jVcrbHIS15rvnWD0Ea1xeaYUz9VkUK8jMKl
PQqxDt3+/wZM1CoEHjFc5hQvbkAR9DGT57lFfmRs/ImZhswNFeVU7FYWLlWYNkiOSZne+tII0qY3
0/d/0xo9czVHWbm8oXYn2CbHt++/WMSMVJnu+Teqcu+z1NmNZol2puO8eCMOAc7eep/vOntzM0Ve
n5UQdA+jLsWdzkY0DsJF+KLN9TGUN9q56Kg164OKVcDEwciJvabiTOntZUe2DM+5ennc+yMTFKV0
bLs3sBJ+6WOT1fEYRxq8zLRhLCHT0ozm/LNSudv/r4fnvoTogYsv87zlulJHCoZbFFqE4VzLyPa9
kAJso9SY+5DHg9yJBUWHe+rOFjneA0nczP2MOEwNll12glQt8u1YjKiHZ3juHv+a8wNkBLfXo46U
SYMWtoO4KvVoGeQzxYnrJO6miYuHYEbXIuMMmwv50yQoSwltWN511RhdiTsujalJ4dGCCRYOGOAF
XXFIotgsfw95TyZm+w1AA0IAV2AGjhAAt6WL4lsZzKrtabQh2Fv8hxLU2Y1HaiWvYXmYH7qzdVJY
6pebMQy4BZ7NOVuQtCZ7VEx9/tqX51aZ4UkR4RS2/Z4sBRbsuHSaI+6iv4rLHUczKoRYirwwgVJe
2AYSNELGZKc+6d3hsgx52VYcCOvkSbjiHp13K5STDL+ZH1ejMguMG6/i0K52HRjPs8PNOqX2sxh0
/oCSyFKksMjeJ/9IfrcW9JHbZLlh5VfHjKn1AVgwfzVewwnCaD84yQG2k+2IAEdpOhOcsd3itdi2
kT2UUb8BKLTDF3e3Px0tbQXZ6c0WOjEobmCsut1UMXK9T6lpR+I3N7jTicebxZtdcL2xTdnMbd0t
63eNSwH6G3YOE5P6EMUibIArNHrdy8zR3AI9OGxlT6Fg8WuSilZwOzPZrbv7AkCFePU6/LgJj45A
dXmrFnLu3q9RO3FnWkf548zK8Dxw6Hx/R54I5IAqErumV/BRLtzxHqvaf97LzYCxiZ0rfdJwHC99
YinMLDeIolsqwBY4dgmoB0sfoVjPiI1J8QWE/I7/3jy1CEMXwsM/lk7A1S6QiCKMdeM74j1rjYJ6
YshacjEUTYv852ZOzTMw8fkgCRGLY2L8/FOVYtLe8s8nRXvFOIxlgOoMpiRTXrsmIwTi7TGBYUFu
/lGa61X4J+yvPq2/OdKChiCN5GF2Q8Rg4ZD7C+4nnp36cY/gZAcojfvikcLe5iXKUfcBAfLp4mSJ
OcftlLuEwXbY64Wze1L8R8eZd1w2vYOaGgb/7ZbKjAFkSI1FUumWmIIj4vhoaTmMte8UrDIYd3KT
JEUR6rofCq0YlEMz80WKdpcAkpIXJU+m+8efLHLCdklvmqa+FVVzQNgaVIkVVH9zqS+4vLho3kdJ
1vU/wapkkF+sGaJtPc5I2CW4mWrvkd3t2Ex4zGgBTtdLHb9ZjN9cvaJ8dqLDdrz3cVwFs80mmKix
HuhnjvTw0ItU40BcOOF6xwmHozOa6q3Xf58D2D+sqNKzf0kL6m+5zx5IullKlE8q6YDEsjiuKcEz
L8PQpVgdBAFtolZO7i/f6hXkN3zQDKvLGIUCXoPJ/pqir0G4YQ8+x8PQIFhb25SC9Q6qLZubOa1h
n4phUWHXK166To4KEuYISP+uyM3604LeZB3/nHF9IM87aBFYLwy7WUak0Lziqkf2c8H2CBvkogX7
JiXk38nF5zIEaWf7k3aLBXGo8TshRGUVvQGxarKwCZF8ls0bOGBhV6ogs7XBJCi/YZ24GqAJC3Y/
kj5N22FWswMqC1PxbmRGKcF6qcC1bUYpypMrtsGPklUDzI7G0a12sltVDrBSu6dhtwMjlKLb6crL
KIv1btbPzz+3UzUULTbsLtGm7YHi86XMTRG0Dlbi/GpL2b86fYlq33akP3nj33OkwYiK7E6ZqQo8
4GPpjWMr+/NmsT7AXP/zINTBEdK/yFcQ5kxVMSznHiVw+nUFsN+Q5vRbFjf/qWzhNSdLoz/hXO2c
EIQQbFx7nSxUp9g/1Qk6vRt+jctBID80ivhnQNLYfV8k56oCjtsH+g1wg/DbrDFD/EhEo8dpzBTn
sUbxlB6UxDJudcX+4eB/XDJriaiPcdJLb1PYZgrtcbh23k8wLiLyuT842J4eYPP74XTlgwQXxEXL
2G1y2ReXWfEQeFtcP+enAP3CSqYMxgWGE4knt9OSXSGs7qZZ+Rd64UUDGTqUmgV9umv//T7kXn0T
TWHgCxVLgP/bUuH0LArrYYViTiaq19cTs8SR9H+V1jhTQyCX9GQ9EPiYq4wlyS5R9ocNNSOPt9fw
Mii8V55KymylJMyXwnkt8mijGbLlylWh+Yzgjxwn4ztmcTMk9dAXBsJTSsOQNj3tMCA7D1dZXF5s
Dhd2C7WPHGTJDWOKmMk4RKjkvzz8WF8yiAxCXdHAw3HD05ezM2YgcQAmdKc+EJGqJA8MT58FU5Cm
LuQFn6QwIkakEiTTEw9gptIR7e++McRadFA6FyjQrOy0XhjoFav4khf3KWsJ6jSFQfeunV40P4/r
i5mrlbinpbklof8uaEZ684f+7x0bh+fONdLETa0W2EB6ylB2WLgwLaV0EZWbrZxl+dB3abyUibXQ
CgyjzlqTCqKvbnIhlmFUyJmN7U+NScujlvpnSIRFcOXEaRzBGZlbZdyo4OY2d6mbFVtQ4/l7CjcJ
Q3SBqlM/3ocPsYLAzf1q64uhlDQ+H7uaV9Ma+WYBTRkGEtkwQsDYXusHVCttTGufyDU6X5Z7jsEq
3+ojBaMhAz33QXedm3S6tjyw+vpZaCSbjHytDMZYeXxKGueHC8pNWTPkxCqof8hGxoOnD2VtvbRd
TfV8vQt+8LVLg0UspGbSI8IO2UTuds9DW7Kzvr+wYWupbirQzv2FmonAsISL2MrF8Hh2DzZ8IUTz
bfiv/qsGTm3yWosIRnMmMg6oIRhXFCaxKns6pdnoL+HhwfTdIFgAMZ8f6XMjxecsLiQvSFhgMsjo
ptaEiyCUT5A85VGBrCs7b2ck3pUNm+8DWJf6sskIhLkTjFHglpuSsQ36U6OIG/W6BDnqijNscQ0R
wZLJYn3BFnJj8WWU/7G4d8CTFR5vFLzwa31pA4/YL0Ydwauik9b9L6lk2XyBzv6a5Xas7R7IBlYE
Z2n4itsAibmmoTQ2cDFeLNr9TmgTht4uQi8mur6A6VeoRyyu2U1ox02uqGKxUpO01r5bI0+hzhpp
yT5KAyFPceT+Beo+wqyJjDISx+2l/04j/c6Lard58gnc6UK1Mwd+OZAD4NPTsM9TxOKiPktTyMay
Y6/EsQJ9zj1fzoqRE+QCbhvHXjl/teoyAdjlV8gLqQKJ4yFlSgMH+CkaYVDlo82bUOwvKUS04772
ctD2OCIpQukPbS0nXEC8U0CusfIpTyCkBeKVTQ9UYkbsa72gZUEMZVwV5UFpHu0crz3apsAjw6Cj
UXSDQr8Vji77mqLTBDxg2WJysC3GpTVQ4fS97grJYOqrvjOyHdZVvnw50Wd1D562CkgOFBvUc+Wh
L+R1M9Qm3V0GV4Ngb/FCyYz+mvoOpCl9Gx6b/XKhNvbXvH47Tl0k3OJm6L0ZkFEhzXdcoazAwc24
GafipTKICYnu9sM/ak0RTEKuSTpyQb3zuPQzzVcKvSX83PLXjfV7aR1kSPi0KtTYp9nCv7zt+4M5
A23Sh15VbGdprvmiGMav5qRlZqF3vJExVyf4mVg29BmAFEIfUsj7/wXWJmd5rugtL+mO2P2Craig
bLG2Sboo3sEVApQA64HJok+qOn/iXlZMXZwcMzuNv8pcFRB1EFSIwObORWKRcDnNlijXb6b2DXjH
lkREcPYUbqWmd2SF6NdbH08QW1IX2yv0GPukykC6/1ZdBFzOyPhpk75h7UbDtQC/ELZ2tXqVCwq4
vf6iP1OzcSW2KG4YbbJfXGFhJ/ddqztp2zy4sMzFn0j9Q5tUzs5H+hq6JQKa5p5dJDnsjaUl+HdH
Y4F1bPkhNG/PgO5ynSIn7nJewB5fW1n3cWPk19o4cx1P/XZf6NQMBsVDQgTCP1Ht/hwcg/D9unrh
Ywgt70+RbsLsqCBRF1Zh3jqp/wpygKWkQIv+o58jDHbINp0sv3tZqT6OuzfoZn4nPpJNDYh3jfSB
nrkQOUmgiJaVE43joSmYFQpik9XUI1Bz9A7vxI1T2FHhXKOvmRMRubeQyrL4xfzYYGU7M9YxVV1p
/2ZQTfrJd30U7/E+2RvysbCuL3QPmZr2yz6OIlnsgi46N197H2Q2+ROnPI4J1RQsRBqKUPfe5L2m
IO29R55IT/XTLccvkkF1u7ucadFEBFDHeaWagb10TvTeAgCwJnY7UezoayVByXCdmHZeFK2StPVR
Pc0ZZOb55S/NXvHRZnI8jFzZ8EGnTo08invBIknmsBH31qjn3/XeH0wkKFLZ7s4Yh9re1wn0MR8F
9gawz60A4neC+6e3C7m6JcgOb382L09Phrvbb1exESCZeHfxHe1Hj0CkkOnn6Sz+3d+a3MUxFk5q
XxGDZ4w9UnD8RkJrF1Vip9/LquRb/ZspSx0kCr9/6NlM8OY5BWtxm2sa30/qsOqmuoKHUmg35Oih
WSJ1nuIFcIw334afLYaaRsSUBpF5Gag/rDxCENmgpYa2FmKBX/CoZrkvSd0X8X+rn5esUE7A8Ekd
QoiMjX0fM3Fh95Nr62jmndxFg/8WC3arx9gQy03ifAn6sQvN4aSGZ/JfLudj+2wHkeEuLoPCY9cg
4LDgJeJurUSmGWpyZJZ3uBkzSfm0iAF7aN1TxK4sin1oQ29hb4PZpm2qF41ISyVOrgS5tQW1A+fi
gl403JQzW6PTcT+I9h+ADub1pqBrqAr788r9J9bX04PCMUQyEcURiR9Pw2WSz8wJ2ZQwd1tkp+3w
cWqc6puVZtNLkdi7FI7Ilw3f769AvijLavo3EPy8WpQuvnCw50VrPMGL0HG91QQ9X6XU9M3qcFmB
R3+J5DeNme1Q44rgI0CjLr5xgnCGMZo6AKUTN/Z4JJZUymC9LGbMA1Wl5JyVM00uiRrS0kjoVuuc
FXE2K+IWOP0glsJDoqnObiDyIPek4R1OVZhVyRxMtWITjaKy6Vn93LudFoOySdROaEzTII6t8hoR
JwoIZkXt1VzE5nHI0cGcSpGmh/acoHmaDofBcubLFUx5l+HDbIYQI7mg+p4QUGiSbZ25jZPTQULd
GCLBV0mjx3XxocdPD5qaHvirIZ84xFNi3YittFImszUs1kIrVvYmViBGdxWRjVEMqx+uk6Jpcxsd
Qsj9rXlOhOYPUmKiuJy2DkvUuW42t3h28QpsRWVDhh12+TSUDDJADVScNrKPRtkminjcJgXN6LtH
2tRUjp8GGz9ABIv2Tbau+Ds48SWIh8z4Qop8urdvGhy3zbjMUllwFEmW4TXnJBQ27m5dub9FoUtG
IYJSIYMoLsT5o/mK6bqQuaHv+zRuSSZEr4i6AOVPk6fpTzdMJROhsPl6BE86GQms7/4EQWPfytGD
owwHaGE6QUK97aA8jBv3DMfRUNW+L1Bae04xrWuWRPA3cMUmeHwOe3LqlWAeJlDgqVR699b9Shv+
vGyJGq1158p6iBZHGTtz5MzUtI+vBru+IcisJ9C4/L9KqWLLyDs0T1gR5ordb+7Gl2w0U55UIaGx
vXpZ8ObKriHkkSX6LkTqVDJdMVkLFngLzUbJmB+rf1j0PzCaqqKAunGy71f8cqEX6Ssbh2wFaj5d
Qf46mk5ofdE8d14ZYt2TvT+nyY0lDmrpqGdzShi3hjzwjGw885mRScZKk6dsnwXsSP1V2xecD+3T
PiJsTkga/eGQIEnwYRkVtrMyhWB2AOBoJt1WbghfOsBHnOKeWZKQgVW0Lwu9SyI30exfm8/pfhJL
RP8A2JEv7e/RkkwAqHKZD7nk8ZHj15GB9d6A8lS/pDRhGXdlOCRrUaSJyFJuiJwflx9m8k/O34Ug
SbYqFssaPiLbj4wgwqUfEd06OUSHB2DdVJf0j7YewHdsrK62w10UCcBHElJ5J05/oSxRHopi1OpQ
yxViBn8T2lL8eJt+FNHPZt7nKSSYYTn/9/tC4zDaxteGSeYH7OqNBMytmgnAo4QsMZBVBJdO6fOJ
o0UIJBDJ6nEEXSJJW5QGC2+nnp893+73OhFsL7nmsRLkM/7RdmJ0BbHuqEB7TJk3cLSDdf03uPuY
o/Y3rE5hnA1naw6dEMz8AstWfPm6sLdFsHkUNwPTbO17acenTPhp6E4tss0Y9HtRooMuoP0FuUrQ
JH61TwUuj1RcWFCXTxhVoP85USa0qDFyPZo0j0rE+BBdQTNMgvxcHPlgyoPR5YHAEhRJ1Hjq8OT8
HSdCuSJ0xoCJ8yLHvGl0lZnV0haQF9dJm/J4jsQ48GCAhxd2CY3kFHvAV9cLFRdgCNTx1yeIS3ch
SRa9FsX8IwIZP1z6NkvBkYZgHMdhQFEXpENLZUdVawYUMQ1v8/qqkrlMnY0Tqj64VEmhpHnUHgyl
nFmsrI+zX2jfywHbNBjuxc3UWmhwNhZVIFoqpupgK2WdYXL6bPgd+u5J2q3U29OnxNFxI85aL6W/
wQwMtBpbriaRLs5gYZfQEivjRMFYj+IBbHUGXGRBcQb4s5VCsxlICIsUFSCJ6cfLMUtRSymF7IIR
uRyLKTlr4ioGAhZVji0BTTV/wX9FfrxYLi+LyAxdF3IvNhHGndqyJLz8RAtrYnycfi1UEbunNwLt
j1PlhjSReTa58ffoiqlCsRV4eHO4F+uvpV5b2gpBnXcMyNOG1mkrWPR7mzdRuYoOCKIArGQpq0l2
TUyMVhOFM9BhMYYHlsETi0gqHhCksZfkYj98ZZ0vRaDFHFd9Re5yXWPHqkm6uK41Knvuj0fPjsbY
wFpdJN960VLsphB7B1DJJs7NkUuTjI4YkrgxK3g99oNnP5ZCf0xNpx6tBMk/2sDZ+sdGuKjwIy7p
g0BtSEDwKmuwouMljfyXe67j32gk+nzmXFgY/7S646aVvtKKOxSL+U+WeGGcu7FbfbvwXIOCEsBi
yBB4lorKB78lhPyREvRxF5ne9Ur6je7mo/xg1G6ND7Dg4IiNHUQ0LL+zNNojWquND5W3gt6/q8nx
/GfC9Bg6Y7VDfm2ABbokTm9yUB8lA41uvDdOZAWL5GIO5nkDgdYNrlKVIKRAy2yLq7hbVfyH6IZt
kFEshxRcpjKhvYmthtBBRRHeULmvWeGOcbpwfkeqFziciIgqrirezu/joemeirD46+lJF7WslQRr
WvblBGMV3aG/vNYVHLsw7jGYEisHt1QzG1iEeiZLzXdwGpA3M1Doj21HnfhXVkFWRxF+pagHRIQf
wxUVdDxqYJ983hQIAf8aXdLR0mojj+jWCH/zQ3dN45/GvkZYXQEFjQu0LwgfEvgtKWhQQzTbjSZJ
0xMy9dTitk9flEu3REwr8sv2uDAIDHacbhaE+c5nU+MxheqPZN6bPBSYeM86Nf6Rk6GVWBnxC0Nx
YtBvVP7hnuInwHwOz/b/7nUzUsG95yfL6ofeTnCVF9ZLAlZdpIOIhaelN7IORtUPKp7iGpVrzXgs
jLTPe+P3punn9TVcSTWBLgYIl34RPaJ3EasfGvX2IQRsmFABf4gPIEKAQv8727kNwFkFtHTOeONh
URyIJQtNBBPRxWcRx7ya3crEePZ0j+G3jKBSCe8RkrwEv7BFUNeAMT+fAkTehZxLxy9mjOdo6t6z
J07RybFWAbx5PsGggz5VOcXVBX8FlDlOZRNVMRqNqI8KRh5tUwYrAVC1AFNSjDvINRwpLlRCOY6f
dDUjgspk+iqITlHucauLereLxq64UzOwP0P0IIveo9CC5XwvCcrKvHFC1ZyH7c/oyFjak3Yaoqzs
hqhRnyoWmny1bQ01kVtjBFMJZs/enLiUZnx7MJuvBn8NAZwo0N32+wAO6vfwGhaeVolxGUXXYTeO
yF2ngbuoi9jchYcRLoJ+9ZlRj+fgSuutkk9TeU2/leBuwQtTwqJYfKTOzEd/3ooCyujSZ3DXdtjs
55PV9lcvomDEIYv7EUvHIsBzHv/LgFyYe68IRmY/ilQcmw3Z9FhWdlFilRUhYAMK9qP8w3gfL1Iz
CCs/pdP6/fs9tUGAqIJ5vIRIVwaigjM+nLH8SLUaatrCDf8HS3zlC3ylbGI0+VYC88nppE8Wo0/9
dWZj4/UzU6FO/nl84lJ+0voJg0ZUT+1o3eK64ZIiVvw6Jy/Xvuzx0/jdxJlDR4MDWTzm3R9jxU2i
9JI/mGu1cYyhL4UgBQHMLgrZhpSU6CZ7e34+Lf4L+ctdX5Z0tmfstO4HPfhufSSS8l/ASxwwma4q
1XMnODtDkhBfLEhL/vxdJCVctwLaE1c4/GU5DWrWcLWKhKbYBGp2dpyKSPa1eFRD6zQO4OLI1EnL
ezoGJ+T2jMVjJmkGC/JQjTJa8o3uIVIeBpVP7GujqSn47OptQN/YQBqjSNZHVgpROnnaNcahoP2x
SnhmnajgEkG/elsjW0BHBmc2A9Ya17PQ9SrM0jcIUTu0d3za2M7sb33V00iMegXdvRTlVDqNPdhP
ELLrCODDQWQqtmOq/w6iwk3f9fLC319v4KuZb8qd9R+OmHQHjsm8xsGjFxowYKLElAbqqvPbhuXf
odX9geef6rY4JhttgAmtqeu2KP926nRYcFEm/aUsebsxbNabEyT2lgMO4fgSHlAfe/CqPr6dFo2y
RCk5/QIj8NZ/XQ61+DXWVnSOw0d0Ng/LQCVx7escDseeSZ7kho8LVFH7jhTKCSYE4lnC93kKCqYS
LyFehZnJSN3zj2+gHuydwxzuVMXc6DK2v6JHwvx9s15oBzvFJDeojpO9JCCle+Ds3ih/6yrWEueF
uqC169pC2SbjfJLO9Cb2trJEXmwDfpeQpPiTr4IUEmol1gyTOtqd/3jwbg2ZEaUPGhhCb5iIydBQ
Q0aALSjZx6wrhwacfiiQ+6zq8f5osajhnc2BKGEbW8Vpe+vNlV2cwdaDqzLHSXPwheNxc6pubw9O
VrcvfV2YZUAsC0nNIr5LNKPN2kJ9fvAvS1jH/8aovGfbyVPM4gJRKlz7W1Wvtc7UvWnK6zRWDkSR
TcsjBpDHH0g17k2NKJVYbaKAg2V4ytbeshoBrohdKm+f/kE+FOdXKvHQlSXlLkNyimbPN5j9CriZ
JZQh1p5dbWR6nDzPXHtqSIoG1yb9Kc1V41gFDUYf6qC+24DK7TQZS4R6BADid8RyTFO89QXjHbxh
1kT3wb3qzMWXQUJRWiEEham1g9ObzYcpGyp9oJoe++JVXHn3CGP+odtYWvCPvqx/2kGyzPwxtZj0
/mXU/uYrpUZ6XlIVt5OEJg+mZlw6xrKJOL3IGLThzkHWH9FsjeFzAHKN9NxSkSMGKLW93UUQkj5z
4ddOLIpx7xUnAXGOwB2CnOLusLziiHoXB90A5Coq+1hduMRa40Mec9dCVfib2JCOssBtksqD1Gu6
Svl/zP1//jVxebFEPw53hCREaCKXF9gtU4lNj7qVLuPTDtSEeTHA9AVPIDciLl4gdE5+0IvAcfQY
O8F/ZLTGSNH/Um0rldJkdl+ho45F9J8dLFGzX/G/s8PrS+IPCz76ch08COoqnED9LPwbhpFdxIxs
6ZXdKoEd3bjqB7eGgwWvV8P1xZi51/FBiWJTRmbq8qbgSegX/GTNnji8M2Z6EwPixGlsqNnZEZv2
Wtld0bBl+6qaP/EVUGn3yfDzfBfQBoxqLVSbhHHDOMNU7owLd+HZVLjoR1Eedz/j9ZHlkmPERLQD
7/xnNt0x4x8kVZvcEK+dcK8zf3qdZvrplaXPMw701D1Zr2uBFScLj8fShT+vnZu+fYXB+cqib807
xPZpKRNqef4yw4F6M9Pq/6yJ5tXgrPp/T+tuuJYcgNsz9f/VxDLIgzXkMtYqATA1qRM7g64+7j80
m6IFX9MkACsfl+EHPtLfB3DQZUxLWHFtjerPvTPQBSONWx1hahVBK/wmRi7TiU1iYJx9Br+xQJSy
MFaf/FjougFNlJLeI8UHUXZgY2VHn0uBccn/bzp+u46HaGK2IxjUAQiHR2BH8X/QQl/IDHxro4yL
IUQ0x1MF2YYlPo0rgioxL8a/XHEZXsXLGPfyrRv3kha/3dVc4/QGStqQmpkjwO1NCFqAsWcW8qiM
p47tDvRwSfQdrHL5PbkaHZnTicIUY3O3BivtdNhF3ONoftyaZ/7purY2ikdWMYAz5wLUe5eZ0GKQ
i92gt+/N0UU7YIwA8YWElG3W8mgJb+a7Xt76s2BBNfnZ9pCd2dLowU2n4/DmGgcRbOPIFrc76+gM
o8Cd0NDxuwkjbhIlGw37isAGzPtHfStEkBhazMNWchpPjOvv5z9q0DKtUPN4jPFXEOK4EpiOed41
uBXBCvfStviY31f3oKb9co/VF2Jh3QhK2+Ln+2ttXm9Qtjdhg6b/DNicNP1k5VYb3+soD56xoAm2
mUlaH+0esy4erCituIAsWbVsomuWVevdF2eK4aLmvqwGIpMGrBNVuru/2dPEMurhILAJ3mYiBVcH
dsJnWlHRU8DdPhZn17uFGzTjdzzZCjkgtIlw4f6ZFi/RmQy7Ef/yXoLnT1Uc8OaGlQAnN66DX2jk
2yA9CusB5TZWcV9iEihpoeRKp9nTiNoGJd0JpMGBd7chhF0mjgFiNH8oZGPd0gqeydoNzC4vEYQ8
UR4s/IeirXyJ4NUK5ngZcH05DzgnnNvT3mHz5n7t/5TwdaCTDvZf+t7TG0rcbbfFg43HAGCDhruU
fRqBLNmqNmcFVb0S1kvat6vAkybO7+MnoO1erItCEZMNxEY94XAXrBrhNhcQL9SI3Glbz83DDaME
MDATwQImhdN7ESR50U26S2cHz0S1Wwa+WnscI8fFKqHL42sEZPXkP/EWkWTZl8Ge8IwCZZdD4EfX
xpQM1hNJPVf+ss6ohRhsy5tMLITbsg5UM4Kh/mtK6SopneH09UJH/2zUmE1W6mX8qNEemXWg8oJV
y8i2vDEVt5sAzq354ijAPESoCy7Pyb7NuGHUC/+jPLTlkXDyXIpJLQG6mel73L1HD3PM+S/hDlIa
u2n28vBV/X2QNeDvL2C15BBbhlNAGNE8t2PdgL9d0gNZVeb6jYTSnjCPD3VTZwmpQ1YR9pe6KGjz
1BeaV/PSSfL5s4XgsogPfApMNYo1Ovig2T87V946RlmqspwDOU+Q7Wk521sF6kzrdhmjx1+V13Zx
Bg/OV4hy+JBZl3GCNo6AlmVZr6jRVs2K3VbFLbQp+BDSMQzhZ+nSSOEjUHlLkx2KqpweBw37KF7P
H17b4fytm3ru+FCwx+K7BKyxOX+krTNvVH0rctRslUGazjrUshXa0EhM5e4KbCI6DlC/Ktrby0Xe
8mHBUSudHaG7gEOg4D0EsD36ybOgHVClNdpNMoFxqpZJ+ESdncH84EFTwxIHT8cI4yVS79JIv/XP
+gua2HURB6TFk8HC4cKmacsQbyXODAYiTHlhYj+lv7i/TUtVeUZjwoLtNB38QNLbr6Rb/Jkkw3aQ
tKVYrH0UN/8pR1M/khQAD3qK2rihnOgY03n9lsy++y+E8ny+4UUEE37x3bRB8rQCWycD5Rb7ICUm
/9OEM6d2Ji/53CsBxcDvj4nFyfVPbvs+nS24GgBNGfcwJi+FUbPViFssyZrYaWjboSd8D84WJp36
ORHsrwPgOA/JOXwRk9nC8sZ3EAxZMsE/PZppndk8wCoTLGX7sBnGh0BB0kehFwP92DR3VLUXmLsj
zQt0iDH7nCilX28sDexLBfu4KcSafeBSucAG4o+ZyHALmHk6p47Mwwp0XBri6ydBONV6KV31c8LB
hwrT6X9hVFj5RNKQtNS+c0Wm/uy5VrtH6NsO5077qHj9YL/jNDx+5VKV2NfU9yiUGHfwc8LnNBm9
K52il+EeR/4DggZY5sMDsV5ByHGAo4ZxS09k1hZtPeAs5XfrWAB1Smr3Tvq2eLv3Jz/BJTADtmW8
xp6Kv2ah0ZNDl5G8gKaWK+QphVedp93/9iURlmf50ndBbg0GFV38DebeJF9xHX2r9i1lJZGD5P1v
njD3wq6YzbZlwOmCnUbrHltLTW6pO6BzIYHHUoVYV8yJO+euRGjXETebyTAi/2MHlK0CotfnIWqQ
/IR4gIaE5A6ROPCkpJWdyVxIGeu6XcyHaZYlCNLgdwjjTB/sx172lxJEorTkkO6JzGRHgy7f6fos
z+UXpHpnU3e4eWBPJBEVqMjBTUYJqSIsxqi16UP4t5N7SyvLKu94wjflf6eAnYeerc0MlVgQ/jP6
rRUE4AOt0gJaWBlsjm8LyQ0LEHZJb1qQZysMb/Yu8eJlDl9dHMggkb+8EjWFOOXZBGGC8uzuJ36g
EaUuG59lKdP7v5csg63GxBS08cCAvaLNo2vX2HZjRQ7Ic/qaSwu3uzHUteifxxKCmFio6ruaTJ54
K9qwBHcP0XT0288gQyc6AqpCCCvPYDSFxuGbNihAIrCdM91MNeFHJXjwSL9XfqNguCHhcHI39enr
SAad/ziVDLPTzXzFuIwQbbCYsATFMKGSoWpy3ZvTdcozhCbePKzSQwNGbVW/D2aF6BtqeudJpIAH
VyUMvl8emRwE/+CBlQv9oyMcBdwxUVaF6mKNm36yj0CDYK1do/6J7go2FYJnhSmSIePHAcnQqgOW
TfcILGe3eW6fZYwkZFeI3ONZuj92Q6gXBNbG2Oka9zKYWNEumN0GZrfaitu+uJmKSPOzZmMNuWOm
RweWs3i8sQCu5QeQLcWT8M68uR4FR50rbXKY3kS0MGonvO+N0I0q88W9l3tmh2+uhQ2aP1MWWoDD
MbJdiwZXWyvzFf8lzeRiDrtgDQzMP9AA+XxlWvvQCeKv/Hq6HBVVFISDClBlBFB3PidjbJBL3jKa
lpF+slPgstF8lZJ9fz4dFpYiu5ms82LqJLUZqwfGjc0xqJKBtPXUdEx/thfcitfv+Jdx6piXz0Cs
tmAit5yXRG5Cuv+e/FU81VkCZVMpESDrt0L8cl0ojl32XjT2f6d/zZLy6l+Qj7nHeGAgr6NsOC90
iMuUHNdzsOO2Y/NYK5rfgyvtQ2c258uYqNXvcqBMuCWgs0nQ5IK/Z/K3jOZjT/0SYUJe0MIgc6e7
y0bs/6ovLQsI9BaIjShOhHFOH5SBNyCtqXVjpiLXoAfa6prs1o6tOplDebqwpSyGBfQ1EpVQVqxy
ch/iUgRRkUoIO4wbAKelj7lTdVFzb94AQwMwylycIjDyQRErOo6R88gCz2N8Q9n3YpjxcaNKl5Xv
2RI3ghN56XXWTuvmYPf2V0jISQV6xsCiUdqKUfpCxS1xscdk61kCXkhwu9nmEzwo5ZQtazQP1ttJ
H68KKiZuUMRavmAXy0h5g5Ns3+g/IafxA4oKlcnXsMa4zaDGPavKxbuFQdLPVf7gow0U2KLuFhmx
oFFYSkmiK7qOtaCJ1u0plczD2gnX/iQT5PKqfl3+X4Au/no1APXlO9S3dgtG+PuQ/5BxcMCx1AK3
cg4yifKELqB7OiZ7neMLz7UmMU+wSpeuCsiKL6JTv2JteP1T51HExBL2K2TPki/I44U1I1DkF0Ca
dXCZ66OU4Tz58au64a6h0HRzsx4bfIgEf8/4g0/Kj3mAwo6arzYoBrL9A6UV3tbRbe81zmqmHVDg
fJj2/9xh+ddbj6KcGkM/SeiQjH7tI92pAKH3ahIUlGNi4d4DDsNd/vERwtICAEnWEuf4jqOQZwU5
vaCKs09gZBsKTPP1qfcExrAOMMH00anP4jjf7P+yEJdXD99DmgdBbHQ74jM7YJtKWNH3He5hqgjB
jjd0qg94OcIhqYMtUAxXKhiCtlJ/6Nfxbw2A1/pL8RKVPkSEk8guQ1Do5lZbTw68GbZz0UVwfI5U
MnVL6XhwgUzu0fvEvwkbbIshFSM2YFX0wffTzrVbu9cVpn7f3Ute9K88vZbkk8Ic89pxZI1XAm79
8SMZ2MwWT099bfcLGK5w6UxGqGixa9/LrESKx48x5ZH2pLQNj5lBhI8Vmqu4qpVlZh5Il7JErA4l
yyb5+Ezw7KVovayYiOpkZb6XvE+0bfo2kJV6WvUNCkyRR1N7NEzoSvThl2LYBx5ahI2T0KavKwMT
DQ9S5vSPSbiMloyqHvNZNPaXEdlm4roi3uLqiLMAQU4hieKt1YGSXX9GNUWgjx1O6J/+RHBXRWpw
u7Wuti44//XbrsUewTMHvxEtsZWuLngRjmDUkN6QWFRv7zRoAgL+odXq95DJmW0vyI+3JmTkrhLY
L4+/vidWl1gViizmvG+Cs0nAlvrhmilbgoB8daQZx8Yr4hXydAsfd3gTgx8dDFUqK5hsczfo5edz
MGF9QNv+7bQYbs0pvmrQxqXCD/uW9UYpy8BgJXC5E1HGzXl/9H7Y8tzqY++oKd2953RBccHcCEBF
6u8677hkgBhC4F+E+ouzWfMtmY/S6kVh/OCjxsni0n6JftLbIRiEMxf0v1iFXBs+v3eHncH68SoH
1G9JeqewyuDWfhO1doxXZuDQgTxZuh5yFxZCE6AFEdcquBbGRHtGY2CdfQ5AGP6r1EDqcbJSU3T5
1Wp1TbjO7yQdBLe9BmDl6XnrUVsV6+nIo5aOmka49DMnl3+n6q49wfrMW/yLjEyy3jHCcp1UPIZH
xRlseAOt7FcGy8nvHj0QGjodgRMuAzfIqtkdXWvGObDv8Bh+s9QMTpc+kBdxYDXIRwid96vqeAYW
sgC7vCYGkzh0W3KoxxRcq2rFBFlbuys4Pf1Nd39TsfszCz1uvHH7cKif5fd+szjnLrnbxRrsC9O3
/x3MnmEKza4o7GZp0y4Sc6XkP81kfSPZ72uXFEgYF1PuDWk9pYj9qB+ZMdLhLXeael17KdoK7VDG
0ywNwdI7ZZkAxRZ4PRu8gLUJPjU+7uWmlb3fZNqP2+twQPQ9VcWF+6WlNwX2DqQe8ny+XZNxVdvc
sZb6NG6f9f/dBf0a8ZLQqLZuqcdaKOb0gvYam3xLoX+RlVBKjXmcM4Hlbirw1FXGsX2pdVRFefcC
3RGd2VlQYXfnBAcSd9EqSh1Oq2hw37xWQzlwR5yYnHpCPp8U9/GowJKOkqrIPAIJabjZtBIDu1K2
kTR+TxEpx0GgdCK9Ob8jTPZTW3EBEAEHZY7qiDp6t/GeAaam6wwSDygz58GL5VWNZUEBzV3qZurd
KRQGqdRXzIJQjFeWPFzQ1H57+RpbyQAbIGX78btwf6qNCdKCRv7VqIBeoY4p8o9dq2xCuDyJP+3O
C3grdr6l0GaCP46Wju/J8//KBxjvvn6CNiaOp8qVQKl72pKTBcrwgec7v7t4TMGfx2elMl/8gcP/
AbD1h9oZAp6vU+virqA1nq+cw6IX4N+yXmx44XLEcKvzq4xnIAcaBXWbD6gvkyzx/w+DyQnpZuDQ
puIIng1qerf2CvoK1Iukeei1+9+nDhRo0OOEhAg/G4YnuLFFb+viE8ZFrfganLA0YFQP/IDolLZT
FxB+8670Ml2ySfsHouGvJvScAOTJYgIE0sPuKFXPuMxeVp6nGl8kXSyUhQ3rII2QB5dHlvMIasq2
0y7ajbQAlxukC+tQbkxmSaEwJrXrjgxWzkjOShwdt7uAphyeg0nwde4XB+R4zsXJQKN8QavtsJ6g
5Y7lP0oQtHjOJgYp8qvZppOxz6srp/he4gm/8gstgCfWb6VlcNCBB4LM2NKDmR0/R13+SLugfBrw
Gneu45mzbTdMPQzl32wMorG9FS78TVLVLNYhhKR9ewkOT7aeGsHgqM0MxbXQGtQUwkZrxztD8ckM
GTE7NBQrsNtiKXxoS44TXq9VYCAIr0baq1WYtaGIgo05qxZnLoc7/MxlX9+VyO1sHYONBMr3ON9d
RzcA7OZwlYqKzbwWMutaVk2N2Du6XyGBcZ2ENwUerzw7bNoJR6+VX9up5JTP6STp9tWqjpoVNq0F
WLc9WwK+e4INUOmW0CT/vH8WGKfMS5qnRafxmhZQ2pD3Z+UIbLNhDEqATP9lWFb7BstKZU9ECkox
bdDdKuZLWQ/Ipv/cFEKXXhgOHTmyJN+dpQIdBEzBQHwMI3kOO80sXKcpIc/IVsBBSN1N2KkQr1H/
CTekp5YNbpECpkPFUedb9jbSyyaogK+DLMjdc3mGyeuIpMuM27BcaLwzzLbUMDrkOqsLzYzeWMii
Z3y8H5EeIXCz+t+u63o6Ss/Uu0o/GZRyowLmLeIISwiEuK3Uci5zxLbqzKt54JA+LkPlo5RHVqmu
DccbbMVnE2Op6rT7pSGUqQ7sW0uW6OYOhndsE8BXWzAU2TQH+dXVM+MiXz3Iy+Qg4MXzGA9+9j0b
AQPOWQCZJdG5elVGlo2aXq6jhf4SKXyLitJmMUM8m0YkRJw6OIr5j7kMsD+ySCwkA2v+RiSdpr8E
KAOmFvInCcy4Ty37ZdeaOITqH+aun7k0jFoR1DHFQd64QWp7An3yAwKwxxXUPMEVz0fet8CH1XTs
l89tnSau+CtPCaoWDqQiLNed0xC/QuTWQ0fG/lP1yr9UOhcb73/THN4xZkTogCJnsFIo8ulvBfY/
arKNWXyh1XNe9+hVRwQAiFRQ8pazNgoKr3vRpuOihQ2OlGqEnogP7s7r+5MAlWp3OobpwYVKju8b
4l8+LCC3gOZbdUvlgTnDsoJasa5iCJFg0rJLcf2OTZjRfkk5RRsmfUP8Z4RNm0kOzbgqZ152ZKxf
VdJKJdmGw0YGxLVI4XEecBHx9c4sgDYPNz7fCCOOp5vCuB7IYZlBMdY/92wwOPlPnSFT54KXcpoH
elkvjapkT321OcARngNNApPfNBU9ifoymWvg2NwM/k2OUf6gxTAuhD6qyGsqTwjw5b0BtwcI1l1M
DnB4eoTuJIlpGUn/fvLQHmCHxlMr0s8I1JZj0yac3rpaiRSiFjx6qu9cXOoCR70XHXcsPVaYp+Kd
u2aj/OFWkIL3hwIsbDCx/C/N6DRMgjcRaDizXN1ZP82FzY3FxXtZHD3aQKbQacnC8M8gnsMatJCm
0Zwp32qDmdxE+psVzNIW2kNcdOQfLayRUH0rrsBILpxzXooanQ8+Bn5eHGaAbuZsp7Yja6U1kQEt
LKSqbRRSEYHEJonJPQPswKUB5WGt4A1+10JRmwNRUxYsfiUAVwK1jEUNbZXwMQC7jrzuqlbgAZZ2
CqjxlsWDP3TG9jQY1oG8+xjulS1nYcB8yCELCa2+XQ4d9WZujGMfiB5Cxj1MkLjoT2IH5CTyI3Af
aqt0rlNBsRREqNqqM623GsqD4iPQsn7WQjdB+pPajYq4M49ghJUSCOBSkdSFZzlZnlxMok97lGWT
gMER51uygtJ+XCVe3giGzXodtS2FhcZXx3PmPIHRPqWO7bIN1VlaIDg+kD8YoZ98yAONmGz5D/zw
x4DR+FHARWYmj+tOWJIeq+JB4SYHPctfl+JtgGAMkxdGcpHCYc5eTEdTsShm7Ks3zzvNBtB2YagS
qnoJoGh2u/+T5gIhGXMnJcNqtpRm68a0W+ZlgQbNaBp1bH/iRciruSXd6CfI1LyBJoJMO2jZc3hP
wYjiQmJnTJCii1iPRnGJJFZVrmUvTuXtkE7z6rTSl2IGpkaCJfOYXa3maK9GJGXLREa23E5HwAQR
6MZFdZqQNMQABHX4Lh/DTRvkO01CmqYxKAzNggnks79pdY7u/eQDbrUZ0/veHucd/QFBRy2CYt7A
2aFj1tGYRGmsKhBsHzTvYVv+9+hCuhSN2oqn5jh6E3/JCQKBK7wMuXsfk4N1/XaJQikIXv76xVKJ
ozyqgaYQyaFT4s0zGleejY+uPbetmBngYGP4QqmJjs1QnpQ7WpfOYwifi/EwCO5gdMaHqJtWYh5K
BDYN73Fm22UD/tuV1NmngMxEYj7JSoAT3xHu2XsA68OgczMRJ5F68m5DEUpr6uhaTJRq6z349lOO
FZEYI7fUC4rfqwnNrJmn7H5mrrO4Wq6RVZJbM0KdziROK5x6yKzPJytXQAFZHILVlLBwkSxFkBfL
JniruQMp67eAE/PM0a2VmiIuqrzItSczIxIch63ztAfnfBPfjiwlalgqZMREoA2RWFu3+v6yVu0J
s7eC038d9BQAm7ZTpE4Hw1D4gr8MuXnTsx0u/Rq8lR11qIfw/9Dju4vsnXcNlgANDJ0iodGqfaDa
HFujTPrI1NPPaPpMtqzes6VUVJDVeVXOCY+uMI7pha7qycTtg4uIF5ZeME8C+De+KBdS8B46s7MO
kFjQnftg2h6RQrTbdNxpWQHxVym5Ujs2lBvDiFaNI9veIlAGAwj0Y5mqxZotDMBQZkdFbkqxjWdL
jq0/iVKRj2CAEXw7xm0U3GVsyZdPsrBmTvpDRwDF0Nu3MhKjTIt00SNnOlcQopVP9jf1oW16w9Wl
VACcWAnU3erMv68J/0r9mRAZ6ptDPqEVRQY5+T9aYf0bD1IkZrpsI3kHbWTZ9ucrybhU8zkxbyXM
2IZvrj1zdEsIJG5P7Dd23tcLkJ8DRfKLuxVIDXKNlRQHVTqQfDYIxlfMI+Kq8dz7x9oulbQVLBFE
n8BbBSRJAjod4/AWH3T0S9bYKlvUSk0ScVsO2i5Gq316rqv2NgmXPEWFa39ltP75Gyi/CwiIoNbu
OHuIW4UCW6ZsIWgYy7OoDFRMOJrvLy4c7HRsC2lEUNW1Ekl4kuPAd2innrfUwJlWQjum708dqAkX
MvIo/pO/WMu7W4VM2/bHDD08aTwXtmZm1jRlEvmDxjJ/CseRgqyoNFMFRHcdSWCN4mNIZl5g2xRP
L7r763fX+ypWKQ/P53WxSYGfF4R5bvZX7qpLv5qja3wcG1u89wiyOn9cKiFYM7qau/xgE3WnG8R1
vM9fSTXrZ8jw3uHYRbm6Kc5WFqHeSq+Miyxgfkpt7r3S9dqgksxJQoZFchUPYLfU8WgUkf77MGL0
Y9toX+L3Vll7YhCyVP5f556RkhGPSS7Bj+2CM4v1Jb1zSabAGO5hlah+qU2zIDS6a3Ek7jPWVj+p
3synzcv6zx1yvM/OfO0Crz8n00sJfQzsn1YgAACNQOQOoo109TijK+t9R7s5595vY6fZuMlAgqHu
I7w2cbuRzFunO1cBcy7w19ElmYsHDIHLfyXzmWzZMmPxtqLJ7oWZ9sAZZE2BHEGKgQHrPfvT+R5H
sXmhOdBvWHri6fR+hc4cjgoTw6fcvm4fwEjdshcjlmEH9Agqc5021+Oy+BJAoPwSvIrg4XFT+OQv
LwaVOEN/8fj64qTHJB3CMcl5tfvuGbcdW+x3Ze8euf+gilHiHSftypQUNdJ9+E0uI7mXlmXVuPGE
1McTKpOr6v410PPK3STn57ndL4dGYd5FFBSFgTU8S6Kxjzp5v6D9Qza0mZCDmoA1HndN4S21RlFP
+IZRoRg8B1zp1IG+YWBHx+PWJ+onnrSymFdbZgWRQ++1zT5fxJ6QrLSn4uMEzhglPsjVC2Bax8Ld
ZYsSi4saSD6hNTvPUrUmmUnGRnGyAGLuOqil0UQ/WgTFab4vXHPyDdUw2oGF0rp7XsDBrwmyVpGj
9diEFImHy1/rA/c26a/nv2JlAtrpbFll+01mNw+1kV8Eh9klXxT2kGBpxetc9Fm3i3jydv2gYPOL
MVNZ/Ea6Iluwv3QP0xb7j1Q7yjU3aU4N9jx9266SwHd8RV9ZHJpIZPDPs0MlqzrZa+XspRabuKyy
L3Dw8xhH0kCZM4V4/E5vtYa79q8wu2OfQ6f41VasnKzS0u+uy1ZvyKw9523dBHnypKSTDVUceOQC
qqbhHU6KiWtbVZcJRnxtcr5y7ZmGtT1LAYqGVP7sEWVlJc5icfN8Cte6VuLoSpfHuHXBTHfA2EV1
HNhqhfwiOZdzV0miFlLTXrUzFLdIFbL5ZRiSGZxkiU4E/lQ4Y20vLiSoruxMPLOpMTSOn5aXFcFW
b+ks0TZW31iJ5WYoEAtYZ7UzHAiCaej2ue6v97RsTdkkkbvXr9ilaNkmPB7Sh/F+c7c1iR89OIyP
Jd+IBD/OVhLxv+gX5BBsmR79g/FnFmZGFxZBSnYx5GfBEex/2u3VavCGug4JyvD1OEs7EQ2dVk1q
D38eebIoqKodSI30fyrQn6nansApjTI4o1Jgv6GkAaqWKsmDcKKugbE9/JOQDMZqX4NyH4gK/kJR
X584mnYup0Qv3dK6jYll2xBUxiXeKGGC8sWPqi3JCIpPgzJDB6y03WJVZjlZRolD/mQPzB6RCiJ7
vSAI1BmrFxrWpZSIHWL6eLlg/Z0GYtZXYWFbIcYE3qgaQ+bgqHknd4N1W1SaImSxIU6huFJlKDsk
qqNk1x1wqL5ORzFxgkSosZ80cOP367HTh4LlJADCI/Kmpq2NjpWRQDCjhiTvbFA1FYvfnqm9QBff
DtIt9moleOmpOZfTChDQJp6Eiy1RcJWC0QFloizYokmRjhzfEPhXROLgX/kCm8uHrFTCly9fLoLH
wjXxXafE+9vYPKdI4xCpArJQ3loUCRJ6SnH1ikwUdP5uBm6IzT0zSgKsX07chgRgVp0G8BH0bKvs
BfMNHuQzkkeX/oNlIIpZwR3YsKHtnJQFSYhRXxO3bGSWRulaJtfJB0CwHOoBT1f0wB9sPn10b9Bj
kk/ITyvkhg41zzqwmj139Y4KKlvc+hWpIhwbmZ8dDqtLV51xcRz7HrtuFs/eUb1OqdhyycEygfNX
g66ugG9bEElr+r5A0RWlShIQA9CDJjdkgquyi+8Uf0Nb2UZlRVlsJuPagcmVyjkTiuRngmB3BylR
n6qGbo5rFw3/kd8gKzaEeKB2+r/beNWI4RIIrp/rWJaQXNMAEjCI1+Dpp+TFwSiF5XrylPU1xqkn
UknYp1irBX4zT01FWt4fNOVuSnQRdoEyphKzeiMP/63KQMnXwUfLJZ4LUr5v15BvqTAmUvEEIuw3
9pixEMynjO0ss8Vcxt7DTZ28rMjgA4BS7T3BXSlF6CLgNkOepKnADLiuAN8rIMANdCt8ROx+6jhh
KIwqp9Y2AGeftHNaFe+5CsBXfNvx5ES6UloQcXwe4JsCypKzW+0CyzOV15DP1gCGRr6qYRzAKYCx
Lgtxthn2Y7ZeMPzL5Jwx9q5goG2mrnFwnpLsE4l2D4Xf8+WlAE0byHDq4kJYnvl+Vomf77BqBVUn
nJ2s02eA1KemaPfej4G/PDCSkoStMlcguo71uF4v5J1ol0nsXIAXSqayU/VzgcH95E7+NhQm6zjK
9DpoT2YVCBlV6Pt7hbo8VRC2H1tjJlODx99EiFWr0IwPoiqnzUWwmFk5eE9/dr7LBMCIrjSCrNsL
Za0Xa+GtBM6zThkInY5Ceu59aF2u6bTZmOeawe2XGX6gR6maSvFu4oBUt4bVCefd0IYyCNVxOG3f
a3bkHVMhW6rua1IEUdoYSOpe9O4IzoCVHH4m1YCvJ2NkB/x9IdHTRjH4MbkYaU9kD0UND9ggc7Pf
yMg3vWlOEuzB0O2BdZ3WSETJzm/20OM0FVz7kybWKtJletnHExUsqwolDPbXGROyt/+5WhBL6bv4
RehrxSSaYiDG5ftyvH/aSvpQGr64T8hkI63nehEwSnRvvD7iwa+denKStkLj9tFAAjpXPHu3bBsu
WUFeXywFV9/XO1/FeDkATkYBFRjujEoNXCn1iWTcOIC2w4D6NJeLuMUH/JmJKWYHIHOsYhSHEqwA
QHe6nI/+iJ9FIJmFl7/72OAu7b1krQuD7IKRuWZ3af12LnHSTPfxD3zruUvKkqEJpE08ps0jJlRC
MSmgBpt0JDum8TwQF2gOoeUx/eujLkjbxbINAB51UTzDyav6nlneS+d9JHSdwETEptcD7aGYaEGg
8Z5fITKXmNSlC8Fp3l+tyuEgqYInGwnk6oCXdK1wq9MHnrKajNohBO4WEYT/EccseL5DtkNYa5j+
mDVIv6y/rX69dDXp2weuQol5l+bZNJcRVIDfMxTp1Z9SXAGQaVeDJG5Wnu4aYt1Frx+FtzXRrbhF
3ltaDXLFc/vFtlofHqwBHx3UVOHUISbCCBKoJ3KFSgJf+Ch10tdJp277Be5rwrUzOraCyoq5zIJ7
d4ejkSI2P+OmhEuVpWZUcNB2BznQLlKTJtX/CDN8EqHKgmbLA1iLigv5n01mWLzc6YXN8mJGRoYE
NnlZ3KbuUvcJMR9aSabo/KoaaHWCHpweYsumHCzgTcDk+hCTlwBefZO5o6Ro2zRSYGXmW6mRd8Wg
y+LiN8aL9CnBO8hGig4fJhY2csQUy3hQfBBYNzxQc1ut1yzUkp8sCridTAUfkQuYfw9sbnEBZ5DU
kPt8onBcEb1ifFcqyVPOsoncP+QE12Qaq8V05q338O+2WxadIG7VF7AmEpNdAaqhjXdiIpQCubsK
ryIArAMWqJJjfIFvu0ftxLNIrUdZ2N0fNdahspmHI9QRfo0HP7hHpFICaW0aTurRIRVBU5wZEABU
pMJPE+br/A2cIGpSs5o0/bGRxc+mfXJDhCK03e+Pxjl2hmjYnDNepDkk/hUaN0cSbrKjAhdmKCLI
jKsPxDq0oEFmJA59SEU98k+0wKyFkCEK2q9UlX5W/mo7owmsJX4B7SNg+AUIbZrRdJS+HkHhHOXc
3WcDO12lg9BUnEsmnhvZBep3aNZkY26CU9CG18x3E2+XsW1bBnjdZecAjw/7O7gqNrgj2IaeJ1RV
w5/oju8hUqx1Pzsf6EX9LfeE6ocAiwrlFOmA/HnaH88DM3qqOB288S8NVKXTpLW2l4tCqLPo4UB4
M7tZc8RFnM1NPFlrGu3o2+zkcSRlbbzYYq3R5qjwQeLe47GHeveRlvRWnucXBl8JSg1GRzz+tBvh
GrxQTqs6NATXFHhlh8tEblMNlRo3stlZHMFvIwXxqNRd276lVWNeTPEhJygkKyB42u5dI73WXdjV
tVps8BTticVwLY1LP0NL0t/qY4qiwUEgJEM+Ct8moe7mA8RgIh0SxKljebcIAd5BrFGXIjTrpJTe
PQ9uiQCO6gP/+O+2XDvsT+DtgZUh2AL7R7vltINVNGsSp+bFrXqz6CxJtl5w6puNFs59xsk4Aszw
69JytWBXobRmjQTDhdoKXQpmdvnuO0fROpcgUaDzibaqgId3u+/l31ubqjbPpbdFIodLka3r6+ga
XVfpF53bZ720hxEC+lkxNPGmSB4DSQAQt7+3HwtrWgbxHyNzoNUlVust7aZSB4EKFBRBSMwPh6s5
vCM4eU6Cz4kzoVADQmG8ZOAFAgVsthr7ZA+S1tJ2XSUPKRJ22Afeu/MzBJacrCBbT6gZLNXu9rbS
L9d7TbeahEpHAcdQKt2fKQU1wYjfIL4xGIaErOee6sGCs8z75LVOdrLHbNoStVhwktQ6D37HlvMo
DEUAo9djUpmim0fuCicY+/uh+kdZPTlgaKs4A1GFFwJ94nUmmMp3WaWMMgXanO31+w6UvQBCSxy5
MrW9moFZSsCC9E5V/zQwKJ6sv1HYrtYHaMhvqTc6ZT+g3pOY6BBN+SzTKl/nDbFrycX/R28R5fPG
oZI2/fIXlpuvZISdcX1V7vx1m+fL8M54c/xMocFBfOjRTOdkZBBeYqZ/Ekjj6KzojQBLqMZGEYFC
lLwSxlWcUzof2T7m11CgkNnJ+iKCa1kwiU5HYhjn5ZnyULk7MaGlJk2Zh6srlad8yMcKttowlVm5
ekJxJ1TNwISsQgYJ6Fd9XrpZUC8hJ54ZR0W8sjvDq4FWXqAMkTShd683mHu+qcc3lyA14Nb1bXDo
ebGWFf/pJXbfQ+yllhNByzr3VtzFY60LlxVQ5Ixi3prAll2RcbBC6BhFXchVx6i9LZXSS4dsgJGF
tg6RMchUFTXqWI954c2uL+ZDvXPx4G6S8QKx/D5cHytUYEIYxT6LJsMhxeEr89QOmPnGkqgjBB72
5Oc9XDz76/riRc9pi2sERh7hMFIfS7/ZXFDaYamNUV7PXaWJyn5YdVDhO5LoSnHcPRRxqrfqeZU+
wfUzQHPicM6+1+5awG/VuFL+4HRC+XwMhO7zWipQgYmxOtqWrp31k25wY0LJq3psIne6V24RdYUM
7y1w/mhIxxXs3Bmtq3jZwceUz4GXl2uAyVHTty6XPaE+Tzv7/8EK/F69hOj+Z971zd6909t+ThMW
vvHj9OhdnnTFMSw6wc0YYhh75ceet6NR0H0kA9Zp248Vm9ThuE4M1RR5DkW05GjN/hxDy7KiaVGr
fhHn1b8vmSe2G1bXhQEC5vxTbJhLaE7sPIWNhtsVtywguLZFVvP+QQwhTC1pWO4eFWW+j/wwpPq6
rp1pHLOL7knTYIx4U1zb52aWq8651elu2mCq9B6+1HJBZp9U9g7GDciW9xLXv59JzlavNDxUFPPw
f+AyUysvKu1IB/wDoBuXArkIrRUH1Ixanx6bWwxsLqa2+rPFCQuJoPO2d50DmRfkUokj0CTD5eNC
RaLe9kbp8sY0+lMJu1cqxFmIkVNDBPkTU7klJGgre8S5iOc8XSmdrYzrz8/z83/LFNgxGMn6Mrvo
T/mGAewy3yz9M5sfV6jWvB5gpeSZrM3pUS8e0QIbtrtkSUWzXGcrFHRzeom3XBIsSxdkh8pyXi9T
/dEm2lYF82rG9PIdmf8jGxoDRO5baHbD8KycMFVpnhSlas1Ei8oypewayJPlvH+0OV2kccfy2Bg0
rbJgPS175MHuFYzxMQ8E9KTWf2iTuXcjkf1BCn7eYFQizwEwKsMe7XwvUSv9SWBk0edXFAnfZgsA
eQbpZzSlpeRDZEe41EJT5DGjLk88NveGw+3T4KFFNOwkUsgima987bO1ZTiaDfO79mKYlX2IOxck
+Thr3eptnmf0jsct8aYbnPan+REaa7LeeWrCq8oNYEwH9oSM0k39dKptWsecKxkJC5xuLJS+PYLa
bv3Dg0uv/6TRieCA+zSCfxsDLN+zE0YiIqrz2GDpzBwZxc4o2gEyWap0drISwUw0t8zpjk6j/f1o
vVbVTWvguD+CqN1Yhkv8ihebNa99vpAKKAVN6xXHsgAEludZzezF2AQPWDW6gLGjMXXWKwc1ZelL
vP3C3i+v68dz4vSZCuzDgifBHTDEO3Td5mRpdahRiPWRoN2KjiYhu2f4DTFEHFCCSUeP1fVz+Dyh
uOxH7ffM7zF2dvSvFbFr1acFexdO3hPzaars+bihSfRieQTDkRBKX+KgmPsGUiKA10Dmm9Fuo1UA
pbQgfGSKzauZxYyzvRg0hfPt0eTSZwcTiRyoncb68axNOYU/EJAnqmInkxxpShPX7TpYzgKFlg48
p2YBGOwqAGIoIvlxIC2hfrO47aVmvypvGNtMjONw7iU5rC2hDvc4XfhvI4mFeIxmfBbG/TQcbAiz
QstjaXGFJmGdtrn7DoA5pST8Yc+owP/ixYKJ3yPCTSmHyOqDyk1/PQWGdoEoQ2oaWjJxgultwtPa
j1L2YKaipPfRbESEmVu5Qjq9Ar/EXJ4MoYrpTNK78yMjEFkvSKo3Fy1ntjevULyBinY1Yi/zpbqa
eAbQtBlT/jmByISinYqaTn24ok8Y0/KKea8jPZIYhnRIutAfjP8oEaXNRgRl0oE3IdbpEae/kO/O
ocWbXUDQUYCoHsaae7MbYBP/MpQhMvrupjG3M45Lo0et9/x7rQMDcaBI0Um+97Lh8wuI71Q9ibhK
qZHhdqMlQgJvrO38S/gheVABzZLQmhiW7EL81crjG20IOxeUzwNjfgoej7QPRMR0wcTfWLghnJw5
L0rYOVAa5uCfxg285NWlTtK1dzBU+8eNkHdbSY7Atb9ZLXtcqxP099lBgzSOiBbVZf66JLWPA9QP
Chhv+0vu1Bk5hgc2Jb3BcLHcCFG/BkVTMEKD1rEf0IdvI4ElWcbJhPrUhTigDfNDgF1OrVZxSI+6
3qWY6a6u4P8db5KgCCSr9zU6qx7ze4QJECmIF+gHp1JsS8zxjaRfwtRb6fREL5EpdVY86elxJEzQ
rsyd7PZtAAmEgMcgJLGxJrGvlCKwryIhqW2w5w3FQm6Tn7QqJondukQ79L6U/xbqHh7ooPDFfYMd
Cg4w1Eo494zfplGFL4E8HEXQvGuHkAeSIpUW1MSWthV6z0BIWDnTUZqCnegu2vy3BxzWz6IcCK2o
ZsFMJu7L21zcvjRDEqozlhunqyZg6GOagaITzcaTJflSp4WbNnx1s6BpRcL3v5CF+8ww+CD9Hjxn
cH7GEIGWtjvh5mo/vdrnJglWKU78ynyG2fReVvndQ423Pwz7NhbCSRkGBHkTZNBml41W1rtM0X6q
Gc/qqQop8iXrK2bS2Cl3Z1bpPF3uVH7MikjeqNcFA9I8FvTk9WP9//dchPnr28HgKseiAc2lKdXh
J99A7uG84cX3vHkKJR/6qdftmtUNNVSq9aLldGgVIe6TXGTEooRnIoDbJyR0hPAmtnKez47SQory
WpT0yKput0ff3RWqXErNOw/pYF7vwcvHp5v9bPsomaCFfmP+AAY1H7Lm0vIkkw22G3gR7ltpnDXr
0WNmridUAMLC+TupbdXcXfJ6sHfiTODeT4SBTycbcJYTh/tUW3tg9OtiYtH/msVOi5KpI2qo8OW0
/OK7EXjSMpFGum1Gtmdn0tht5MwCoI/rTeMRgXyj5/zGLuua1eCxx+9w+nvizwMzKTCkvrJqSVJl
uhGPeRKe2bZ4fJqQdTYiXn84RfPamRWCLWVCx8kOlBducX7PpM2jqoEYksf8tm9I2kizDEQk1QLH
ApHTp55Xq1v5CDImUjzsXFFgxsWSCs+Dr5Ao6+nkx3m4ZmH2/LDE/ZmcrpSKc0n5Nc/Afmvbzbei
K5RxDufHgH8cgjai/rbpqG+VnD5IRnXouS+frNSwYcEanuRPhQhZXJHNbpCZDaXhIzjSMIgzmwZt
WVdu1deLLZ9Wzu5p5r3mj1SpW9wqCxuAVD/+f3xylJuANXlJ4cUiB12iUrB4ZCwMpsgcddV8OF0q
4JnzmtePVQcGg10dzt6oJ284gLIMUH2x8waZ6qGfH+JgbiBQXJACtKZoT9mHZf2PvF9bwm5pFodi
Mj8Dj6zr8LPXut9vKJvBUSyHaL6AwU8QfsQYHBjXdrjP5zxE/ZCdpUT+slexD9k6mNde8mGPolWX
5mVe55+a/K7uk1Kmw4P37lDUEx2mjUfaC2K7s28/jNKeWjW5g5OS2RSXaqX+dRdDoZFokJXuQs2Q
wRPa/WMco1VB9umSbWguDBNxvbPffyDyfrQb3RbpJy513ebBv2/nqFdI3P87VKA4P/iK58JBwKcW
tq64iSAda6fr8fkN1BpIir289bydhBoq8GHAxJMHUobjlzmHvR85YmkyM/G/im7mwgonL7y5jJDL
F4r+I4EL2dC2U7HhjzFwRYUPyrxHdf+SMq3LrBaRJe5uV2JnstVniPG4HmIwVmBk8R4RgAJ/c5Y3
smvcYhdvSSPkFGpJPsAQusr54U78XFzp5YDqchxuodSNWZNuzDMsfOwu9AYhwXxCXgqmSj5Ja37V
dpQIfsGqbwa2VUKTBZu9azVNo4Z7zjuwYTULVsIkREWlFVCHa4TMoyFBm0DqORpnF5K+SKuufd+p
jKvh7ExDD5ofuh0Kpg8QcowIlmOkV6vfWO8Op/7PO99cNgagrSxuYivXUZGIjwHWfz+mrxkm0IWt
o455j9FQP9gWh+XrlwDsggzJdWiKJ7Yrky/ehHg/BWlIQoLHI5T2KYQlJ9uCqOPwpzGKzDNGrtH4
nwuiqiTX27YsLANVpYsp1PcM3X3q8YK5ivd5+iY37jsIiq+crNG0LsWqBFyoSfs0540CqpM7dH9a
nKISUGlNejxhtutydWMrONZs+lCqsFisVRfPA1by99O9QNnKm3BLmzC1TRVq9cfmNZ4YMvGP6Y/1
+uEKjLByH/vmrHjWFuVr4DIgQAlH3JeNALBrDqqt35GRsYmZc7mxjzbn0j8yPesIshnzJTWphn2S
p01nz3Jz0DETBc2v0smEPYhHjj6HQbD9B6XNabLWwkNvihRnM/bWVfk/FQOaD31X37kHtMHz226Y
WTbgWf1gf0zFRs3iyJFxFF1n492hNa9SyLBCRDWhcDfQW+FxdVH54IsyKtFzLofY6K5D8saB6z9l
c7oAjea1fADaZ2dFwfgQ17SOhODWO+pvEe37KqiH4FLRPxtC5/2TrkQa475rEpanindeB7JFmufH
JZ8En76cUpk0di7QVn9ykt6EP6jNTn3RTldrIYi0dywhbgUEw52jVXi/8bffnsQ659M2liRGpEeT
RxgSkfmG7pAgS0t4VJFwdndaC2nCgxt3JfO3s24yjgrQ+dNdXt7FVC2t8YDjdgLCqbIC1qnWqWqz
YBT5zH2W+cHlN5LYh9MMJ3yxIIjr0QUFPaHsHlq5DWyxCH/5m8ohbeYD7KJ2IdSlSMGEV0PyHN24
va0Xqkn164ZgTF6Ek9g7NwJdT3PhPM3ej0HxBLC//JfQ9Mnz6VPtOYgwqeunh+lNNa0nrthgIQQS
Vi/QaY/LSIq7D43EMfaSdixL1ZmveRJlkJnN4HODqpI/M3yVLi211BlzY6egmuf977fluRTKgzGY
KCjsLVHFmwHX4wdOvGxiAXPfEVT9KUlYUfiBwjUHzw2VzgPbpZXfDy3mlMqcIeAWuLz+Whp8i+Y/
GXynjHZ+2jnLGRGG7OBhOa7jcEbur1i3fRxJYO5Utee1i5e+4su2nknJh3gdSTq7Lh/f6h3DdRwW
lZtZZymDVS1lOwedoMRza1cWN0kvEjrNta0k/jZQ4HmZcwNAOqSNs6cmjWBJcMz0Fg7g0fEGr0Fn
koDOFhDPDyBXPl6eL8EUS8Nh8jWgRFI/Gy4jPSzgNvrHv0JHDljvTDclnunRNkLu5pGe+Go7SMET
CI+qL9XmRlJiTEsNZCDDsPibkSnYc3QFUcqoI4LR8wazN+n76sW3Eoe9HtVKIM6NeECCWoVq45Mq
bGi6bnF95IHwthN1s9jnyVnXMWRYiA7WmQpzCo01uhqnrgSpgFAiy69qIF5GiiG9/bRUok0OPlt6
3MHI4/VJwoGy9TH627nniJhLGJOdGot8jT1BJm+Coqsnv4qQwasFLLA49lWB3L3hbby31NiE71Kn
MVt9FCC0/mG2N2JrzTqA4xplGhm51cTXAQGBQWOdzCKrI5cYRibKNGeKb0z4tP69RjshQ0vSjgu3
43rOZ7Q4vuRAIMaru584ViUXyecnLC+QfElFp0GRaPWjAZGZdSsCczyDiP1DDGeObeH6BelxwqOT
pbz8BAnloUxZt58p9zy/P+0ZeeDZZdLgOEkGaHuZXASqTEomT+bFBTMMRDQr8vw5JIA+9aLz736Y
JX85DqWLaXlFwO48KSxde6mqM9Z+LXDaWKM1VlEvkceCoVwFm1e2slCrHze8bLn46RKc8m9cuPZo
40sMb6zRokQVhK+CUpJtHZDisjfJJjjJQTNMuNIhhMbjPBNDLEqix8FsiC+a2p5fJOiyztbZb8kG
gGq4HIohklax2nVnAJpVaWh30d32Tt76sporhl0MHNgU3a+BKmFGl4hnMyKDgrDM+LkoTva6zLjw
s5MwucWqJxkHdACecjApXb3auC/2cuLfVIRzpPYX7ItageTCM2UHifLnYsf5Sn2klXxqj5z20z7T
kv52YjL9gpcydpDz1dFQyiC6BNVs1UmdSdD3r+88tcRv9kA8EyIcj7tYP3ADBSsohWCIOHHBhN4m
M5emHJcAnVqRGAIfbcXMi7Sop2BOXI2SggEzuvRpFV4PJ6RTo+92/O5J8HtrRKu4Gpee25FiBZnv
O6/bE0Qg7L6t++yyNc5JvMR2chfFeTrRkpDrljVpASzQTIk1RdZajTmuoTNfYXbQTFhfb0ZnuB7w
HUpWhs3cZFTDPzXPeYfcorOlK3NCuoA2ZS2ZFk9nsi57uqvjpDAawDQKuLZS+Uhp1V1uKZ7iMe/h
p79sBaInbr7304K++ATkq1b658dMLwRf0rLLNausKDVj+qTfLpm8uY60GMDe16ph32AaFLWyfd2A
zHLH384uQXpQq39/3SGR2k64fMXfu7wUspggapRdr5xUhkP2iq+lGmCORRCZ2khffzX8kDNAp2WO
N7OqnrmWTSLkXo2Gm5IlnZANu6rrXlUSGvi0wByfxpF63k1zmkgM4qCPVHvOGf5J+xiNntR6nbaO
nefgJQf7jBy8yDNQE9uDruCQ2hjsapaBMW0Bn2lLbdWAfVnG24Th/09u9Pubmo05FMUdf9GtGlYx
XEm4ItkcHtsPlmplerpvyEIWUtB/iIkNmfRiBdv/nGlQAA1ZMRwAgpdSUZAFW4Ruoz25AazuKyi+
epHwlWFQQHiVJaBNG6HqgeLCEDCsF8cdGxvtKjI3/ncA8TGqFc6V24QOF4nn9KWyzoshLXH5rjpX
38HkqtPAQetpC2K0j+BryEnMPuawmW19EvSFlGWK6DjNZS64mvKHCvO+P5h/qgWo3dv+gulD8bGb
YcBy0jULWH7eNi78Mz8H9bCLXVchu3NG5JF3ZVQy4y01wVWGdzOVHijDH8PiB/VjPNJiTWycGILI
cy/vdAS6ZJse+tUXsloPnfXeT4OFvVLtwhHl0WwI1Uh16vU6o88+I2h07tRDsac6J67QAIbu+DQG
tCJcnmTn2X75unfDACDguRCXYbxBpye5HvjnZBzneGvRJIxdm/+TQn2ovWeoh22ddsxaWndaF/GP
gzVDBrKShWQod+GhvI+rgkVEqZ1j0L/Ro6xz1nBl2C3UCFi1YqQVv+nhGRbwSGPofEvWu22XmtrG
Nj1JFGPrIeTegA+ew1nt82IEakLK0rzwzu/N5MZOEAskXwBrPjA1215xIKo6BwItkj5KvQiC8Q15
ikpvopnM+BAOSym3p2JWBouv8mqZG/cC35n8xcjDyl3Apu0e6mC8cNCavu07gHSXW3ZDpiltI09A
r18mV+UmNg3SFinCTS92PXDECVAM7yjpJLlc/r5wZQY4h7ruznonJh90tEmwMLEdJpXw/4KEIdAh
XurzoxEsgntTEih5sYHfH07/T5Pymco2gkMu3SMk1vEnXZQd60a3R/1FuqW6kPjcjFanMX1/S7yW
QNfnuLgnIKDTJjANbbdUsYfhUPPVlICbQQOWdHRlsAQ5xeQb+b/mceqpuSd/u3EkzRJnVU/ZCo8c
4FLnOZRTmJ9jfoMfuV5DocDn2j+oDagZVnujto87fRzCLs1GlIZ51suGck2DJpL/hFZz0okUx8aj
r8VA4jROrOj3U1laTu2kUwPQo14SazDNUiGXnr31mK1CUd/+563v6lTXyjAPSxidS8m2WTgrqOtr
HirQ8/GQtK2kPEVBzygQ5Qt1VWdRy2b6mbsi2OdvaQdXDNuOG7lwMam48YthNOj2kBaSThpjRMHL
/1q71FEnri8eYmjtypUTl8EN5pzZJIcLGnnommK6P6b9jxHsqKAjKG4GKPQVN2J6zAcJRYLb9x+k
F1x/v8XNzxoKEbRQj/qg8O1THqLJC7aFY2WHIS9ihBEK45DgzgPi8MksZ4C8hsqtyPrnSvNcE9tC
o4iIhpqSyodn4DS5l4LCdj9ETImX6qNF0G1jxj6Ta9bCB6WcdrTRUF0/jS/0xC0ng1AQangQ9Cst
eXuTvVt1gcw46vZlpxc5gXaj+7KhW5SgyTFZiIpKauvlsCY10NH3cWtFQ2Bmx5FOoCgZndhOdlvR
tKLjVVVcWiWYlFduOT1XKkQ4q6e0OrlkTZ/TrDgv3PoPwPb9p3CBmxGRD1UlDoZWq+bsNx3KNVNd
tFxu6fbN299gMMf2u4pPKnfkMe7IX8mGPKXuol4GRGIUWUn+3vBNaYYULuEvxc+CVKp9BxCh8pWE
yaiid7NL1kpCija6CobHqNR6gvT3my6cqmBPOXMMhdZ9tIIIvg+4ugG9McAjHkmsDZ/t5AO+qzXM
RM/Vo+xQpdbYFizbqkXMxD9aeT1wf/oZi+RTBt9gZt/GQ2xg93d5PSuPoGYZvhSU7SnTHoujuVxe
WYSu3I9XZ5SxznBafLHumipC6wHhJWB8xmTMS1R2RqxLefkJtkUkrTyMJwghbCFmYUdwK7qTXjPP
vtmCvmc606F29I5gBmLWr5YtiBnqBIJS8Hj3xVHWjUReDZedSmfFr6CAtgaQYC5FIvuvhPfb7mA+
In5LP7lgqwO5NMFF1Tj55dIFYN7jMfe/B6rZm7BndEEXj4/PZ7XdO1BPsPFHfiJKtpGq4gMYgTrr
/p5Kk3qZrw+MfL9yX3FsiZnTGfDHL11deQs+J7G1ndMVjmEtEC+fHPk0WZe7xNPaQkuNodJKWJ0X
FZ0KUtmgTaJgUiMKiWtMr9WjEReJyxfC982iVHvjFlgT+ToBWuO9Uo/v8P2hwflmGMQ2xVCG7ftH
aajb1iY90bFIA6UnSOEwvlBO0SVSbbdWZArr3uyeiSsV7PcOWw3MGe+Sn84Qn+548zLCWayzXdol
VMZ8jrucmopVv6k22h8LGWmx750QLsAJgb4mBcxUEftrBM24iUgJBS+ecyOJIPYiyHhKObPgM/w1
DESZOG88lJAWQxfvPynmUrzDsGsAiifK295ZwJXGFD/piSlvUgHQM3XfGX1+QQWdlcs0y9OsXlvF
Eg/hkK5VlyVhK+RMT5AuWvNjOIQ/xuN6/Z31kny3wvQATOmgPlZ2biPjWa7tBiFRbCtaXdQx9dZK
LUfFI8L8n5S1E6IMLm49eAQRn1zTRTB98bAPMNncR8P/KUF9PuZ4Y+/imZc5CTsd+4VaZ1gKxWRn
pTJxEh9ZaaoqpL/CULd90mb9g6mOePTA7csPPKhJt/BgUMrOAQ0nmM9hHzC5OymR6qwdew/maKgm
+5inmRJ0p1tgIafCHcCjYb1fBsinW0CkE7vrKpCUIJvAc/T/KS1pSeZbz9O+Fz0n9Lze9mrULeVE
j4K8VZF6Ll/gou/e3owdSLClJguAjcsakWWh89/PlJi+vekGpAop7YqqahVYwzWraRoioBAIeTKB
UKF5snDXNChd/iR+D6JFXvH+S2B2zSmW2KrZzH2tRag9JPWuPPhSjA6+lNxKIilpxQWCVhxnG8jk
rvXcfI0sT7kvwZ3dfE0HtANGO6KpNEcGt2QayEKnOPb8rs7QAXhTkNyTrO6vGU3GZCOjI/X1pAcB
30mvH8ztGxrQUm8ZN0plo9ovPEdfmVNQP7eE6qCkBdce7/Z+WD3nHrsLfFesUsQWPtCchHLMuCg/
hk3QlKemAVUgd5RkkS067klBTrXNHvOXj6Nu4wjExtrCT4kpMw32ZqjYBiWgsDBj7/hSphLAHq0i
1T8II6gw6MlDzF/9AriFVszwaqs8BTtFOrqPpiaffs3cKfWrZnVYBSKILBcZd4RHOweQhd6WTU9w
MERiW5A84tWp5Dq0APq7nOc4j0xbyPQvYf72NM72dqkhLymnl2xN4s6dx1tl+qtsgJOAahQSqA6v
zUU4qTv8Kiri0jj9fj9OxUiz1XDBGrzBjki4rPOtoHa4KiTyZ0N8LBbTZVUOkAqghwrl0wW2dmVL
JzkXKv3E5pt5vx8rY9BaMPw5msMjNzT1jNUhkCE1oyCulBrLXpGSwYY2LwHJtvXFf8Aba3x2mrgO
San312+ka4rpOsLv7TB6FCeBiWtBOnyPcyNjvrB4GFfmeKii30rLRbEfANxo4r7ppMe8YQngafwd
LfCky28IE2SdK9LMmgDToYWTAZDMLFG+WyH0R+/Ex+Nbfw6/Mi0kGLQWQRmbhZkdldCIurv/J4Ga
PumQ5S4eRDO9npwmE/FVO/bRjTnLTGY0ysKcDVJI79XlRsQvhhxHH05jojL5qisT001g3JV62DtP
QJkhgNOe2es7wbduFZiXE4KzUdCNNZ00MsFlvtHeRSnv24L99ocYQd9hSuUj4VpaSpT/hoH5G2NJ
GaFbz1m4/3rNzJRsd1TrhnHm56KkaCP90unZwHwH0tcfH7AUhBRY/LBw6GZWvDByoLGp13XGJzNI
2E0ZH0Ivt8PgIOHhx58HVgNdvZSR8hAganpb10l5/eDXOa54x4tXKW3CBspSNFf5NT2A9gOhKB7d
wfnxdqS3v7RoCR0rrlMohwBbny3wVG82GsdHmPu9WHABGZvFTQifmk6VHIC2HG51u3PE471xvhKb
quUBWD5eriR5Nc0Hlm1aSoPpTgAxciSMAjMjAmtKmiey+c1pTnCJjpN+na3qusLpPB+rNvOdlstc
op4eQV6+b3Ei13ce1GD3mi3BdDStvnhBKZFarY2NkeBY/D5M3p2Gi7m73RbziV+Tfpwx+ynybbSX
8Ow95ymeLBoRW27F4Zwye3gWYXtAhrXLKWMyYHYvl9N96fQlIcAqjQVvijRuheAwCylV0rGWl3c0
jWNbcP5YX4VItdLA2i6jUiHdqLF2NGShVUMIvuECz5H6k+fPsTatu5ls5NrKVKbnRq27Dfbsat0D
I94F2eGUxzkHTX2osPAm4lfuhziCnPbNiOzJUC8yjFLxl6T7tLVtM8xzjWqPR7UyZj6XCkqabLnr
BWiE/7PZUR9Dd6WCFEp1ZRWXCBxwmmMdbMQbPSWMyFhJvENhVTUfjhYzySXZZFSp6wwMF0czqsq8
32GOyrtaLw9Gj8dGg05YBvnDckVnA8+t19JdSAFuAOXeydeI3F0yh6fuzOc/W9zBnKh4lG7MSJcK
GvqzcY52x5VryuqWkcSl2Kf52HLn480m1nsdGl1TTD+gCSn5ijl1hB8XR4e9F0NtHC5ZwvZ2vnvp
6kOULRHfVkMi/S9QDn2TWyi7zdy885YiQmmntTeHJFutSHhgcs6XKjTvuCnnAbdH0CqqizLboI+Q
AkiRe089n0cdPPzXf8JcZm72K+fcWfhYcWgaGFDvzR+318lhatouAeD3YJInAW+faHK2S/QIeDbB
fGWkU/ZpRXdG1binSuvGJCC4c2X1kHnC0m1vHAYa4hATGPew9Z13JoTduMJfASG/uriDmuZp6eVh
Vz41sfJaKDjoOpdyH22USYFjitI9axi8eltx2iE3JcGohaYPFUIHwUUV3G+gpJEarvuXOrWo+q3T
fWO31ghMBiJOSm5ZXYa+T4rG2Lkzhk94rUZu4LUcLRJWtJxoqixTukhluksWJ3Uk5d73a1+n9+CL
G4iWf0oOFURp7nF9QOfu3hqfjOQrf+z1hlKLMpir2PODD5dUQxeLUWQ2m3JHMM3NSsN6Ow9Y6xP8
a3QrVT0YkEeil/b5sCaO735MFX51VDYs1MGc3qiiLcIkMVqdi4wknNwcnOgPvCiltsDMKknjbzSV
l3KTdDximuBh2w5sSyO3k0CNJuYDTWZGV1hrso2Ed10GXcaRwGKJIh2EDJSvax5EEsWynGGuwKUN
6YjWPechEyymSih87SbNOiY8K2knk6jQfEY+VygutPOEEGlX3rf4gezWjaI0rjQWI9qr0z3c9yhc
7DSW8IQUhOylZdviR3Rgk+1abCG52XvgSX8fdLdwWA7yqPO38YnCKJVsj43Zk5IhTx9VtFCj+RUn
SMBQaJB6Wd+xhRJCMSJQr0DA+Uj8r9oXe5gO7oQFLIBW55hEfyLWHGA18YznBhllP8tPoz7qStq0
AD9Uyc7IwPTTMz8RRqPGS+fP0liYvtsoW29rjIERb+8EcvYeyze1xFYMFv8aA6q5TUGDbX8tKi1P
nJqNc+PWEsyOmnOuchgdw9NJonY6zPKzcwlL9QOwemhHjh4akot0yFnx5yiY8OxcXFagoYGwTwjn
nUnjWvfqiNBjEjQ90mqz1gI8Q01KDxwsRD+nDwmP9abfZ/3a5CUADWR2hmIPNmf1wmH3h6OH9So3
yBNA6viB9SrIt31dEbHlNAyhmZaK/4EsLTzc8NfhOYryA1BYdQZRvzlJyLi57G+fqYoK5Pg48odR
MF/927C1gGEwYtV+W2RrXNzSzBPYkwy/lrwh3/e5nhWSE7ktB1WeRxmW2Qb04/mAA1zIemIlmwAM
lykPeFvUKhycfXoLV797KdiRjDQp3zjIycZjygu2dZeeBq1YRD9s8zSfzPrqrag5MSioqry8SllV
Cw4cyahwETC6k9e41GvfFhXqA/k7xHa3piu5IYf6ThWdVNY1Xa6mS4uyGO5ipRm35BMoQ0TYejDo
0mDur1PSXseaYqY5y1e/9u0kkYC30c7clIBbEYnAxTyX6RNyGAl+6T+IYZqRtnKR97HloHXcuYet
NVCe01wT/+wOi0cWMw79hqAs5U53IXWVn9O2IOyiX4uLj37lj02Er456XN/Jj1etKZ4myezpWsZq
AAtedhCtBL5ycAadovON6eTcK9PL8FquH3UDbAh5/zJjljCfjY4eTIXe0ZtMmDv2f8lNHi2wv9bp
Wxw7nXQaeYfkLsL2ZwhIG/f9hNLc+PNVc+s41Ml6lMadBudFLED8HLmrLCl++Iz0W8QA69p9ib0L
gzsIA3mHcNeNE15LDzoO6h8eiRKb/9p0s3ok+z/h1uk3K4NWcanLL+FnAUpwsxSerKh2jQi252YS
V3dnCM8eNxRBnqHVkd+2EVnyiYX3PJidxCrnbVsCTMNpHnC1N17Jf+rICuANNIViTTWmoKS/TJnZ
tIcVpC5brAxK43ok6+hMIShVftVkoUw7e6hDx2HiBN1J6nF4WwV+lhmDZx8fVuc/kuv/UxppenRo
PLKnQGfDwGG4HaFMoBGXAJp+o0my3qIJH+QoSXYx/0av3Z4OOtv8PIOqVJLBWhW1GS4BMHmkf8GF
ViMT5MPJaa7Cjw9f40VZo2MGF0G7kxi6apgG/ZXDKjUaCbTr7YDONpia/tV9S72QjaXwnwzNWjoF
QlhN4Vn7NmexQ8aDOrg3Ynq3pULZMJx5BO32565WZevzeoK3PrrVs2pY1NdbX7ndJwyzhQq5dtFB
c4rvbHUoULsrjIpaxmE3YlXE5jniItS/r0e0n3aj4DKB9hJfBFlkg+I13Bqkn3x9+6oV9/zSTfL3
ELTtXszyFNbcNWxRTRK69Ca7be2v/swIoUnzLcf1/Vr/wqURPDEwzkIyJCmJuYO8CzUljSLAaIr9
gspZ1H9NEQE+C7kOUp06Wzoo/HACCtXREK/W24fuf0Wzwtjb2fxWEdR4OD74WqvfUwiQNZR6puWC
Rohuk9EYMbcF9Iu4q7gzkOqzIufbxm3aSpvljMQuPO1AI1FEcVnxOaAh/kZB648HJWdu/GgbE2wS
84RziCYxMSXezxoms9l7qRtc1YnC5pNkhGYEBKp9pC8x4PMytmyD9ksYijNI+a8f5E3CC0xyCmtO
UIQ784EfTuXp8f4RkNsLqyhbT03NCNewDhDm1kkBg5u7b4iM33+dL2wE8fW/BmOysUqY9yqtCnR/
m5sbqhOTzffWLSYlLKBqOJ0eLRrXufN2biKstGYlUSvh8/xjPSG2RXsNoaz3vmnbGkNIOW+rt1D8
gZhRiQgIeeNQyomDYZsBt76SYncPLoLjbqSAt1rJhtMmREbjI27vZiKnU1l2jEe1tQKCUHTw22ty
iC/jtJCAEvJbDdkkqLuWTZXFpScuv5mrQSOjB5QJTMAlBX3ISJlTsJI6yfXa7zkuDvSv2OjcWbOv
rD9w7WeOS2qTMvtOtEC9oGFs1daudVaeBUxOLwU5mVGipx93xfCK3Sao+nOYuMLgdhRxyLixsWzo
kzddnMjouBF8nQj3REIjl5oA42GLL7XeEPgZHwU3Pt+SMof78XWGrbLkSI8Zyfn5l34mdicwUV5A
QNhCP4X9PHwFmmFEtHWck3llgM9J7WLaXt0yfJqYFb6csvIksD562hoRTu6BzHen2yz8TwxlZiAF
tEvJGtME7ikjIktwANFywBDO9uPW6yOXvVgso31mfS0b1iw8LnLfy0J4FD3/zN46F7FIgvkEBH/q
z3d6hFYMFKlaY6jV3hKKKlNFEp/B8ELq+iYcPP4D1I56V9HIHNE3ipkHLg27Y6m1oUrzzkZS4FZi
OzCRmw/SBTPXMta/Y7ceDx+dm6pmZ9ZeKN3FlO/DxLXNq9c4yNKAoRrUAurrvb7FIG/HPrLr585O
IkUmY9pUww59ciQRkvU0/A1HhbxaXcTTfi6Z+aDwnBn1nxc9cO4PaX8W4DyZQWOzTRKxyflNrRQ5
DsJih7jN1PBPCN6FiX9XT4POA+qmwziylAhRd2Zi9QYBldVOwzzw1u54oE+VyHiQpp3e1BMDn2en
7y8eY/QP3ctlK5lIfZqfMByFRsqJsFy7DpttTfbkYxvcuMRArt3HG17xMtO4pGoPt5Pk/p6YbKNI
gkD4LFW84zzEnPcgpmhheV/Hryijw9xId65qDwdA1fFbkKOqWE6CccTq76O0lP6lEaG3BUikb/sN
TBK2xUnZu/wU/9ObJamKOaXlnDODnDhQQnvdnyg+zLO8cYWnXLEWPxu3N7SIzt0eJKGoT9KjS/kW
TPeTgngb01r5oivPSqRpGt2d4pDWnJ2auj53+OnK4vN2eMmNG6Eh/89VxkDeu34UtQD0iWcuYE/j
rsA6jlAL0hVbtuA66LG0IHaPYSBHsSTmMIrCCQNgxl0KsIDE8aTxDs/PhOCwcqLG+Y+BF7GZM5HB
EJ51Srxf3dJmWlMz/UHHG37BepunSqQS/y5TmcuzphHiV1DZOMQW3unDU9WIqqCrUL4Q0bSEQJwp
q8McHdWGFkwtU1w2enrJEg/5RsvghHeJKeFusyTuiVQPKyjlADkAgx2VUx5qLEqFcLShtdc3Q+Vx
7eXVj8lnkwEMHtR5LXf/0u7WTFkXKjbZ5G8Mn0kePDFw0Ujd3NB2ZJu6oWl2DCVS0+CCwcK7c1jB
3S5MVxu9pk8Dx6o9FqPxgNqp6LsEymChsqSEV0HrpB8qDMFc5S0sv92urIQhvr4COn46/CvwJIX6
ZAY4Opyaf5L7GDqwfvacbTdkFB6/iTljmprQWG/zcIAfJgIc8WUfcjZWVCnlVFiUGBIZGk3I2jwL
lATlEbWPynxCkjKcG5Omcaud7BU99vALrlRDsRYrhsYMD/tQgVof153TS6BdXVEln/mfwYI8JHp0
fhYdqmhvfgNAGnvbYAl5V4wCE6OskAbRQzomFpkIBA5y6kmqzWlA1q/u6YZtfisc1WndoBdRWme3
81FEfjGpM3oBtI6y+1VNVjjjp7WrEiGPd9f+qGZyyty7zk05Wdi/ihXbe7Gc00P3/ulmhy3/O8jf
MMRCiSbJtYXM3/8CSP8Bk5MnFRY9NM7HEN9H+kv6Apz0bTJ/VorLRfvkB6U3Nd9Ukp8zy6JzxwE0
fQJQdXmjgdwNEXcOOA6a+oBzeqyNIEekKdFkciTM0aB/PjGvnTQaPuSCAUW+5kN8kKFE048QXn3z
vpqjsWXX7KXzVm8uuh/723kNd2LRpaXfkcFc/Vq7Ypu95xkJ7V8agDgkHPSblXIz95irRiy89tUx
/PNGxmfajxg+uJopqCONJVWBpU6bBrZcMI+MypbzvzE1caGpweBtNXYwS5YM17GAo3xkxOd5ntsC
67fHuVcb+QrPKdqjZHM5u2+tI3FCE3ywqJsGNYA85TqmWfopzUf7DGmYCcbeDFQnVW51jHQQOg7D
aODuNdt1dFpMsvic8j2KSREGZ+KgXhJgnAYpCAOyn3fwRbbLXWIRYHGeUNDdaQ1wvYL4GxnNvSW0
Xbu95h3/fZspB8829jwAPe9Yu6gR3Eqn4OsHqNYeKJE2ZwcI3PEboI7nMIbvektmR4jC4PS/JPJB
pRVuDqM9XvDr9/jnOr66qDhJ6WKv3fTLq3fCOoVWElyY7twZMNtac/jSY2dDMFvXVVWKMmOnMQ99
g3QkeyXd+KB35wfWU6LegY++B91PEwMnUzgd/+T6TymW3qYeBsm/nxoIoXhye0uldSX3Q5iRlWNE
STT9C6xVC68W7YCe4cbSMwRgrgga2KNakkktN60g7yMNsRzLi7cLcfXHH37v01WGcsJoV0bgX9lJ
Xkm9CyttToCkg8kp2AzLaxO+oZLvZ4DRbN0u3lnPds+UFTc2YEwkHGxMNwmUajYweLC6Dq5dJxDN
8m+lxHakEOrYS6EHTYMTxpN7TfGCEqpjtkgO9VtUAyCo6osnH/twhEUreGW75zTSH6tVFLvMj8Ud
FQWbTSpUFQ8nlhISMbL9s8LdfAxPte7gfE5YZ7oOSDDTySWEQNueK7+AEFKxJP1O0B6iMVsePBiZ
hBcBDpdI5bHnsXWA3OBFKBN1dRwpkHqzYFd4QqHaSMblnr1ThwLKP4uwyIc7mx4xM2N9S1HWGHIb
+Ns/SDFJ3UgsTQ5IKdEfCo4VFfhVzyeXPgfzBxcNPfau2ygViqQn2QWoX7Nf+C0U+okxotuz3kVr
TLioxkrsK8zbOzzF9m0rZnuZarOz/LEGUTwlmheqzfmaWmvpZQglcL+wpbQmmJRj/p3c1WivlTT3
EmnPSAByuscA7WsvOAeInaNMObNGqDwH3eOMMPxdH3B0Dv05ur3fnjQuTXZhGL53oaNVXdmeGdBe
CtXEWDDqncUCI6teX7Ee2s30isCfU8CkBMN3fzMhilUIg31uDG6Liu9zG2XREQ4W7dWZ8xBZfkGD
TWTzxN63oDIxBDC6AVY3SBYFrMFeK6pN1QltsUINdWzdpKkHuKekDDJkRFg1XQDpUD8DktrkUj6/
7eH1LkhEGPcWhDN9M33QjmmZ1V9LEeAucXf6zHbqPFTPHABihl7no0pcIEMXZlOWrbKhz8IFnSln
/PoCeUfrSNMHWHQrd2baE9sx5BTTQyngRpb1th9FeZB6HTHj1ZYB5RkdRVMILKYwTmolwr+0Gf5p
ZqjytZxmpLWHZli2pAFHExDgXcdZZXrYowbG6cin8NluFT840gFFdXrrdLFXZe9w/urAJLHmNkql
WQXKHQBM0XB55av1dUOKT+OpxazglTs5aGE/8oK/gQPIYVf4GKLwAbpBl7KSXEccfm4YS9ypWzHh
Dr4/M/rv3UXN3skffDBRMkxGqD3FIYmdMiSTvK2Bv5EhIVsvbaCT4HXwM6/WtSxuB8n8Uml0nA31
3d5i2lekFRHg/oE20erArebdfixvkADGRXykvJSVcmEYlZg57QL++u8oUwe6y05LAHvpyH+OMnjE
pdGkG9ZLGS0tVZ3hQzOvURFOrwUFqwHb0XWXifcelfSUth6hvgLcz7miwBsTNqIqiYzlf12U5Va6
IOSwUbJbjs1kkvia1UmfP5iSrQbIBH53p0QkrCtyiqjVKXcSpe/y3KF0ikOoLTADJD1fZBO1TgsF
Vcx/FqxF8DaI3qEo2JQq0QuN9kjyMqv69E99rHDG/IkXEvStWW9dBCdLaI8E3qCAL8n3hs7rumlo
JoRe7fpKppOtYpX2PeKORrb2mbFoNPlhuLmAuJrJJ+C7jVEKWCvM3BRgQ/hy7nkoPJFyO1fPc68V
SQ3yJOvGZn8Uyf5DHUHnKcv4Z8A3bYC2rF5FTgoL+5s9KD4owJjzFdZW9umjC6dQ+cv1TeHgTJc0
71DTRUylhM2RG1PPkPPfj7MS9eFVY2vfqDUi4i+QkF45nr/TpmONVunU92LxDznKkPibKQgIYpgJ
VHpM6kQZk8k8OGDtBRLx6javYwePFetfxZEhbpER8dQox1tBnP5eE8pHAU97LKExZEbg6CEanXBj
BdoJwbqbrhe5FAYNv5IziT7MRQAhXAZfjUfc5waYG/d70QfXUyZ1YloRKglE28p6lyx8GwV+qmlj
9/Naiwqj69W1VhrEyyd6CghDiFA8lnXYQa2RwTdfUzjkzsfT+dbYyv/co1ij/asmfjz/uIT7uFdG
hjHFUu49yOoiLk4E41uYtSIBv9YeDTKh6MwGx4D2pVjnT/Jtx4CYUwowa9/5IMyjkaRJe9WVQjkJ
1hmEtfWXARvQ0GZxvDoFbuz4zMT1EozCoKQ/+8gGJQOgBiiq/SkDlRROzNsPdx2zdBpq/Zim1W3N
zdost+QQ9DlESQYgGzFvlgzQNvVr6g7ubNxFevAaZDoZzQCWycgRc0bxlszwgPFvgDYksZDkxJjx
3n6y/5YJavJRBw5/irX9bIIXSHQKEGj7HUC2lhYn4i/eeX6lujCnl/2deQiJ9w1Y1K6N06lHUcaR
PaMmQOvYQbw3UzK5DDJ+UZT7NoRROLRmb3KQYZvrrtngx5DsKE3+a4jiuk/jXRQd1SGOI3g3Rlwx
CJn8OC9EgHNjDuKThnhghCg5h+vZNx3x98uSJrFAXsQ8QebeeWoMtCPgbczt7Qm66/o/E1RBLtYf
YToj2v/ig6L+Ek1QeOnYf6lEn2iEpuMb/ZKwUc72TrtZ5XrZtjjF3XP+ClgLj6tJ4Ys2inS9yh9+
sbfm3peYjcCduFD0iWdiQRqtU1spvgxriI1Q7nSnfcvnuwGnHsJd+AxT0jPluEG+SJjtyRCL95PB
ETVhWZzTG00H3PBWaIseagcHFkoOMejKUwptXEKd391QmmQBFivFUF9YDiBQaxKyKFcPGFLU3lIv
O56Cw6lRngDX+PurcVqry+hszkDJMVipTWD1fA9OfhRUxvYTagt8g7wvQD3SsDY62dK6DfpIzOqn
thxZP67BHusuachkQQvD5kek7r4RhC1/i4JOL+yXoUK/0Bg4or/pMHFs3qMLhmS1ZuB3Wm1vmEXB
8XGX/kvVeTn388H8/VI6GmBbAaeHeIphpyWqAiPQWkBTzcMzbbmXtpEjnOR/ujhhUVoZLnJBLHqB
oW2cEyK7BtgevyF2mtU9g/Hhz3AXB9PD+3fxaO3xjWOl8tLJsNI+bvRvCjHUddLqe2PkMrt1q5Rk
DFj8gR8jJn/67QhAWpGjLTfs3M7gL4w4/qqbJOQDkRdN9XqBZR+57Ekib471pKYj4Ot4rksBFe+/
iGE3tEkHP18ZtlEqXHeOnc7WIFyhgEYxTWJzK1JXekf0K8c+KgwY7O7h/rLUY2nEaMk0qw+XOrvg
XgIdd5nZPf0YDds56UKxb2L0EbyfPJbW/PC8hLPoJcRQfThr8EKB8rSaNfMfv0UsnvK0XBhxkS89
Lp8LMdsj3gSKHXZoldKeXES3TzpxWSaSsDTuHJh21j/pWLsUxJ68k9uDq5QDbIywRSvmSVHtdv+X
dQMgCXLJoRjIwZvm7OZyxwYTqe+ge+elA34aqwsg388l4tT/nc8xV40FPp3iNbjVOiu6EX+MvzH2
p6m1mbbEXeM3NCI8GYj0Evq1Rs6QJYncRxFDPZGaoNAT9ZZL4jIbNfjrJBepO1AizSjSvu6o8XXK
H2s+N1x3ZScQPm2wyX4s9U9yCpyT0sn8LiFz6egeMOT4quaBJeGPUDdYs15QlywE8UQ/VzRYQAQA
yCsb00cg98MuKnDvFsJ+fPFe/7rrfWPs4ARDuuGRT8WzT1HHwn/vRxpw+gddSpvhgrP/s1+kZq5r
koQfwBHMFBQS7ngIDGfeUDWUKlmZtAYXaWYxKrq7Hyg3JpS8SG7tuIeVVnGEdoR2BX2j8RmdFcoB
ArO+sHmtlen/nEUnNDsNLJyWkMecuncHx6cUOJr/vKfEEoqduhVdyKFEkN5k8uT0RCUQ23Vk718R
nS8Uklzt6iSrQo3AZdWuCGjwtu7H5kmRosWF4g9mqa951MLePKm1Z5o1VAW0i3zO4BkarYv6xf8y
ipzSmx7cATGsKzqBxkfB5R/nQObHKVNRAg3Z1oduAt64UCi+3il2vqxdSdMCmDo7HlVY/RS2AHGC
X9Tvty8i7r1MCbs1oJJi/rx812m7lnndo8c9tKgGAmOSZ/OXPMrBddj6ITc4KModmdB07rFocksj
1lRF2uXa4NSIEV/BSSOTbzjSf1MQcgctUes8ZQAmtksBaEUmACXZVS6SRNT3RtDNhQYtgwP+RbqR
ogJsBRjz6EDMHFFPG1iX0EBKuddXXg0pO5pxYdWrT27gnv+aopugINaOm5s7yb6RQvyWSAwfB1+r
bvzqgxsTPHsmXQbGG5+lEcxivOWzq3Oo85/qoDRGEu7uDeUgDgeunt5n/ARLdv+8siZgoJ/R50Aj
CbhP2ydlrrW4tdkEfwpcVApc3uB4ZQtqr4Xh6oh2DfGqQeYcV8gTY88Rdfebbnc/fl9G9i5pVDJ6
sYxaIOAu7DL08TDvNJVmTMPVdYFHcR7i6/QxK3JvbwSV1siC+YFp91WI6ZYueA8e48GZ/SZsABPv
nBnqMVMqjYIio3+drmaPnBml2xwYenDgHpz2F4EumqHDziaRM7OTwTeAnCA+O9tP4LPYZCDdveXZ
8qTfYNAUZGU0ckcQWouhNKkhjzl+OB/n5e4H9fxpEOKhDLlfzk4jRnwVRz4csN3bizj0fP0ptEJQ
rublkXBuHOQEos+hNBxDnnMFHF79GB31j/31UVObXVZJ2rCNerfoFredzNeDa2UvzjQRdnev0Ved
RoIVmGKh3cfXHZhCs7OZ79Cit5NCUziOzZybkNMOMeLHN2n6h4T3SLOkNCtInkaEq70tKbkaitoA
8hWi+BRnhdaXwApK/be7H5bwhwu2S+jYSaCNH9268lBvI8CrOWZ0l4/2wMIn/YOk6PGs6Q0dti5k
jpeKTDApUqik+fpwmFIFNezCRFlTcT9tGQMJgjVDYjd+ncMuaJMuGdXDkBGSKh4AqJzLTCnc/uBb
y1aAujL6dge6nlKE4QeOL/cJgK9lX/fV5ES457x9If1F3EOGeiG6sjU+Q8dLDPw7hcQRLfdB9Kf6
fEmkQ41WNjWfUXbteKSyHJxKm7tgZXFDWRZZ1OngGLpRaHgRI3tC/A6dD+3vX0Cr4HLQ1UmNHzbr
+LOn7zO7s/pZicRX9GqnYNnvyqK6NxjVTk3kABLcpsJRfp+OzID/kqAi3VJu6LgMJQow6guJnw86
SvYd1JfmQ245z/lbn5dLb0rX+C0/y6PHU5OCOthHtNEWSrR9TCSIcSt092vQERYdX5hZEMCKZhKm
eg0HsSQ9aMDt5eA/YPbMQF8DrfFZViy1zcNBOqZcuzhNPOH0JoXkT4lToVLMX4j8xCsiix3xz2kS
zkvu8vZTu9LewbGGZve80/Z1dmTn7dGYEeG+89SLmzsN2mAERJrvkPEGd3nFp0SJRqSzSpF0X33v
OYV7SASx/7VCLvqpUkXakBM/WsS/xdnMnhEr8Kt5EE9Yr0oRFOZu3EHl6yny1dIm4gyoR1Eat62Z
kOwSDQecYkR9ezTcrsyxiqWLZW/I15ifsvK9e20eBGLA2ekdBsBhQ0fEJRm3wgln54Y88S8JiKwC
9D7rnKQWCE/oe8j1rfgZJBtjDiFOJt9aru3uENAFOsjJtfn9hLMlP8P8yMd3PPG0Vyp+q8abwdiU
CRxMZU90syq1BtnloG3N1vsP8bKaGv6MsodaJcxTRQTP5dbQsCtdvGRYLyQvMkQTtTysDPY3td8i
x3OFan//5SNKLxqF7zabeHydIsSomt5gOn5j1uojaSwcidlx4b5cyA8alZL2Jb16NmICM+obVxsO
aoNeQYaYZcjpb54Z2+Gk3bkYXsSbk0JZx+IhnUttYda4gBLoAAuZ61IIUfORRMm+cqEZPk5pJ8R/
LspXPiiV2vrZ5wTifQUy5vBkAsvNZKVlNpsckMfYnmUZkEQf+Ynl2OJx/KJQvXx6B8ytVoudsB7V
uL/S7P1Q+NM+J+MwaN4LLeEKqUC7AuTovRY1r6MfAPZFeHItqJ76EU/uZgoqxwlXeyGSeRFLfrBu
zx4hNlSgJvLMo3gKhbuZpWv9iLAgDXQyqyOILbAiLmZBKt+Wsj2cTL7VywmpDaaei4Ny5REhImDQ
A1Mgc03Xr2wCm0z+NOuW8JOeMWAsfBOYO2llehX8tXMlclEjMcHliEACzNXa8C0N1ol5cCVEXawO
JXUe6d6xCxmbAoHpUn8bBo4yJzJ8tNs9qwAtXe5Tn3TpiUJoVGA2qcBY8FS9nevM6d7s6c8ph04s
ts1WHaemWKfeGTa0L14Rcwl9RochtoOf3GwyAZ8J3uCl1k5wrArwMROSZzYUDW1F4M9387bHV5nl
ikpthRTozOr4YjkbU7ikXwOHWP5ViSrk6IQWjxlpUL8CKMDYmwWNIeiNbR/oc9E4UKCRNT4M8Fc5
K/XlilsIxY4jUQK5TA4l1iIVzw15UPV2bk8qTmvF8xyJAqq/QwmZodGB9jStC3fcveEAV078vHir
8gZpxZ4m7cf1dEV8Z8VmehJ/625Z934zRa7mLON7XzC4jJG0DHMjTlbuVjYLtEgN3sU5fPXjIfxD
sInjBimH3WGaDQ4FSUa9CwhVjOB0F7xKBD6rWwvdJoYMkTcSB2+g9RTqk21JWEidM3KuUK0tSfgQ
JX6FT+mKc+rJu+KLVrajcwXRC/u2EC9pkguYLKfBqw8Dxxi9N+FewmXdWL415vn3xhjJc0FyFK+K
prPpXgXvS4S1oTtkwhck6a01S+Uiy0+1326Ayx4iTzi8AkHI7vlea99Jp87e+3aeOvkR9B6BD5w3
9PJaIpSnWmBIe8vIuiK37nnwDFLEesnXr/jWi3UIKf5CN8zfpVbJ5rdv2wf4q6qR8wXBecrjN78D
vSC6xwdLAuliO+pePntswZVm+UiFOObV3PEX6OEP2FGjl1liogz+dFWyINjlDoaBTvuofCuWby+z
/B/0yB1QRXHF4YjyAdjm6UP/rxkpYuypRXpYcf7fntM9twV1lrUZ4x+uFhHEcziuNmLYJKdZDHV3
yMktIFD107ehz0WFzGbeGySo7H0/w1cuLCfFoELazriHCwkki2IIeHIoxN0VI1wPccOM2Pyz+DnP
XeD40EClLUTK7RZvjiO+CvZNOAi/EZjbYPh5v8+Tv7ny6dzheITFpTJt3ZQ6W3iONZV3BWClyoJ3
M1zc5tvfFGN5CRycQVm74DsU5Qn0Zon0Jym+67QRnGlXUknj6N9evSBLQhcn2wb4YtRo6GqdJgRA
YfQbX/Kt6QLTJrkO+GpbylYjf+Cvy3ACKYmTryJzJQBJhZrizVaaY0fK9yCiPV+nUgcYyXpTYhAg
qNMkGk0KmxnWGqVkf6a/2q8GKY4oOtiYB4xvjUqQi8YgL3/KF8D2Oqe9J4NC3jSkUr/GgZnq0hvl
BE7hL7Dla/dveXFfYovIIb9JNG1g07y8CmX2pPSghsROEZVAMnMJeagZ/CrIpXmxlQ8AmzwgKyqd
ldaFjyCXI4ZtS3B2qczoIx9+Y7heYRSIpEjkiZGz9i1eDq0DOkwLRQMoJ8/77pVi0VGucIKks1lq
UcRKpyhP3/FXAFBt9g1v1YCtpIHzvbpE7AMUZeTK+L56VeUTetpo6TUuBtO01tUYHuACPT2R1csM
99WPw/rWxjvbJ31akmFQ5aYmcP+plADHoRL/Os+5YQ1xxeEfsNvK6UzlcQrg0AP1fUpD04b9Z4gA
39FwgCYTdcxvJYLWgD2bWbtub507eDhdNp/h3J6+F9yxrk0/3o12uwwT8yRtO3fDcuif9JfXnmRz
WGvUNX5yb4y3898V4/PE/Gh4NmKF8TaINDBOi63dDY4452eCfzOljQ6w6BtVZEzI1QQCPGON87wW
hX6DO/YnXyMmSKRhecAK1PdhNIwDaIKLLBWNeuhuruKX3S+d77duJpYNRhCA9X2XdI2fzJFqsho+
BClRdxF+L1d39Etdy52soL1QgUG3CZk6/BqbtGFWBcP2a156A+2NiddivRdcpWPP7tB70qZMgTMj
41eiJQCd+eOBrRfhRm/zIz2RzmktRzza2Qd3GV+kBBaQ+fXxI3s/a8WBUZWG2mwPATteQYFv7kPW
9Y9vN5a6833KRtcQ9G4LWbFfTVHOgKyrej0CJTwwQco7hDO87scnsM/TbM2dR+n+HjqyTcTds9Y1
4LuA8bCx8H+TjkwjDJpSyppmwagrPplFD34PrvM3Gja7+R0O13M5PDjDfqBcd6sQEZoDAmYML4Q9
+QwOMXK6XPylTaRkdko9JwjlPsIaZgRE8mekZTI+ewlFfKEr9aWWapBdQRe+nA65FbQCIXooPpXx
EvM/rJPezQLej7KSdf+Apb4j3C4Cqu7HFr0VxoszkdpcwEwc5S9sSG8BXYl0mlMlNeU699LyuD8P
fX8uoXGwrpFMiYH3kxxyF3gWWqE4D0CYqZmAQ+PVNW1d6gLPzbX9ULM2jMdm4+vK2r1TtYESNDEE
LvnGHrq0g6nTnuAV93mthAsraJkYi9xW+MaiwN4Mfex6vA7nirNh/ZHuTVVbd/ychHNr37kEB9OV
cmqfv1gm0XgmtwDy1tHlzyIXwSMy1EFktVz3Nr85RlZ7lfbgFIesqJZSG2ahjGAPuahfw1BYFoME
Y3oZzu9GMXO/WoovLVedW9amLAJBD2uLKA7hop+SJ3xkrm+hlvhRiP2GJHlLmLOZ/Nu+1yvMgnn0
Mqt4AoHhmPX+/bJxdRxRPDiCxQf3H73Xolv/DM9nSLw5oFWZFMKMclEvgX64QjQzunPzpFqbydBU
xiM4yWqV5CSEXT2qgcl0w01N0lWh3VteTOfX+kxkFbYcZ6sWsheUpjixVlBOzf6+pUfMoq0t7b5C
JKv6EgqipYnS8h0CFGuL5v82jH8intFJdIEiVQlOybJoG2C24pT43Uy/YzqReTBed/43Tqg50wKa
lSGg6cbf7J4aFCO1WB1gL03PWAcgS/Y8f4geyEDJdS9ARJ5mAHp6TBzzinlywhSWo4XhSnbYTQRl
P4G1OH9adunVLUQYZskMIwxrD8dznli0NT3QRtM0A559VxjEDizbZSVD/O58KIcBPjZik+J1O8ig
QS466cOn+zsypJQXfosYSh22eHa5/YBT0c3H81fh7oKNjFOix+B2FMI0MOkpECpvZ7/9yUDIgllB
o6Mpuu2ApmZMkKs28CTHyPBkFpS3Ox0g9CYEqM8jK/lvIp+hQssGIexWHqm0qpeLX5m75hia2bKw
0B5WjHPT1rptGpePbo4flbRXJMKlOxEyDZ5ZFTfnapwB3Lm7KqAEL0WkLIdTrSuQQ5sjIKy9XxIu
nDr4QJ/Sl9FkG3lX1HEnyVZeZ1/nUuXetCW5T+gfZSeGGU+yRtbGWQM5evQtdvoHRJqOFHD8XbNm
aiMDg+2b4OopyEhaB3+cdEU9VGJybSEVH2M9qQLKUBAsSd98fLUNn98cZrKTd1e8B1NuxswSLnug
5KtFjeS2NtVHkqU8o0eskmuT097Xz2zSeZsqQUcM8SQ4N9EBiwQ7QY/7kS4icgyaW4ZDTUlmIeYf
ip/LlQVTjeWmK9raesc/1X45qAMLoSDGUC6kB6T7T/LzhRw1llHb6qHdOuk7T2uwI8NnMPcZlCBp
6x/bT4JVzKebsoz8hxDiKGrjsZ0OfHIDRAdLbQxACFS3VWZjyPnzUJBkfFzXZhJkio0s8BdB1i+8
pv472WphPj+jt+JQ2x2Po2mDAkIsnpVrWrl1dac/noL1nUORWDZusiyWsEPLhnQ6mUubM28sxRlP
Cuoi314rbuIkfLRRzf7rDVjTwpckVRLt2aCCphVZVNbkDubOtPftjdSNqTx57Q5RC6I0pX1zR3/Q
HWZto/inCf+CXMTmw80ubSn3oe6XpoTqhkuc21geJXQkpE4HqQlpAUlqkxAToq8ecgqnsaNIlyku
9zl7qpYOCDZ+0z3V1bOlMmwuf+26LF4oIjhE92+xStWeWh6OrSd5fVoVqekTZ/WAB58DLF9AIq/B
q+T++YP5XEFqgR+D9a0w0S3nyyLWOHwwyIeGBVETK9T8CF7IGoQ2urwoMnUAdhlo2sXcqlMcaOf9
jMeBWGgaIqFXpp10SbRNwIqamC17rp9qUbNoH3jFAV3uo8KiJyZoQhw0wd6guagHQAt7TGaFa+70
yENuNggS2kxM06lFIDVSN0vChIYv2vcPFeytxLhnNxMPoyDO8AmUKak/nAY8tOnlFS1EaxSHYWJ0
EnCso0ebtrPXoLbxF6jfrHzyvFKcb6YvL5b3PTsmSIuusObZEzCp394dvYTq3q4fcco8OH3PIoWp
tZe32XX0ywWbw1sWs6BVfI5pYHWzLhFnmNYuvboVOpU5aMsgkq65MfVK4S0C+5GxsjUJWtRtmudH
iWo9OqFRJKDmzoBNlSGCsOSL70L53Yb8hxeglWBt+MS7n36BOx23YWsK8VtHQMiJyZyP7ulFKMTd
9OS0ZrWBZq2kPsowJnZjJSl5E30WVjjfbFE863CoDg2feuJ2bf/Si2pEggk6hOJnrotr/lxlWUmQ
wPQDzZW5ToQvx6gnBZpadvbdzUR4OWuAIHmxArVP/CW4kGyW1Yf3UwM8F9KxR+PVssl+iTheXP+W
GUlKO/8ucUeLYxDMyxerxkdjy/OiGkTYsWv7Y+pD/0A5jbi2s8jECUJKEVKnMaJqjNVRESWb2CPP
ngGuScoH10LFj3tD5sstjwgE+GyAYdkPtHDuPWZ6MRCg4Uo52R/YU8NVr+DhmuPkeuDiWGVkEaE0
xQrTeYPOZDeP5Bofu/7uMk4h8C+EivJBY6oQKztPLXS5s/XeB+t12crzAdtTJgFjiIiLmCC29S/c
yx1jdI21uLWsSUe5q5mQv/ZM+3gSQR+PTxWqMXBpR+CnhGMBe2phyA9p8Wp4wmf1ZxVkuNnd+Wqw
pLFRiXoXmoGFbK6VZM1eC6WWIuKbMVTbbJEU99hGmYa8NBYLuh4fX4giHBlrUDqy7hhoGl9CfTJ+
ehg+UfiybSMn9AAvu8Secxdgh/wa29O3O3SL6EnjcguRJp5X8mGWLM2WhGJjTWiNqgk3pOuEw8Sa
XcrjfM5gQlGD5n455z3itbkqYLy3HidUMp6t4iyFHu05tiyhqLkN4JMy9vPFloK8OBufS90/8RZF
+NNfA7K66iwLkGj8zh6NtIRDJL5jVU4/s19+nOzL1DiObykBVRFfIMVPVrGgIDmE74fzc7Q50S03
REA29pFOJXpQDHZtE4HRfwYKf5oWZJVsGHhHLHr0GGTFrXNcGowQO06lmF3FZ7tHH1XYIGK6aQPQ
hnARtrFjl/cKWqQxHuTdUpHcEZ+cEMrRUT8dtAcr/lF8i8vL9QdTH8dBdft0GRi+/nPPecVEq80d
ap4YBlcl8uvYjrPWj8qNm+nPU+0GknRfXyTSgDrs22LJKLHMA4y+x5FLKq9dyIYBGwwMHbOnG0s7
203A2y8uX5w5wsykqqMmjyoa6LFOfwrMmM/tbFnj408zZj/CUZcSLAyakbQ6b1PFtsDWecLmPQlB
gY31Jhx4tKqJK0Lcl13fSSOCSpY3aPQ15izjSjvi6dUEvvZOfvVYD7WH2ZJOIofmDGDAuUh3pmWF
ZupImGFcWAhXotq8z7suZsflfSAR6brKiKU/pkbNn/QxmpTG6Dye8EkBhZoU4W6Vfy4OebHzP65V
6Fvo2UGu3f6jc13bZ0X5ubYNoWZgHKo2rwp44QptkvEmAm0uehH+nNkzLK5aQzKYerGodpZv7HY9
Ys0wNHMzb7eKPuUe4SOpIu6Kfad10hpm8nx5JV4AtRs/HUXQowP0vY70v5AkVyOOzEaHrjxBcdw4
6y8sMzqssAKv3anqnzR20ngu9Uv57h0tBwhkTUDWNaLzIfkykNaZqt5oW/5LQPy41grneRTkgDLy
2fWzZw3leJWtCWa36NAzHT2DiCJ+yDjKYfqDRpqt63TOFYMeFBOpx/EysiWj7J/rDqBoIwiVcFN8
FgtWAfOV2NbVZ4KShmoH8aq3EFXxRdlQ65IVIv2dOzRoul1kkE1G5QYpj+mU5LWNi/rgwf3ioOy1
gC8J+dB0eKIOgmu+Fs/qduR82VlQ54xBWBPY4dYFt8wReyag6Xm61wTd0oRAOrdfcLY06FqCLsM6
JcAeqt8G+KNaCTpDMCDYaayM+3pP16n67nmttO78/uYZ+6eBRsjzLIHiFd1ybEDAFPwB4pw7XK9t
vUST33XxmfqMB/MCOB8/6teHiLrocxH/k6Li9Of6Vj/p7F//hoiqV6yMGt2ZJ4qrhbjU8PJKIhGH
BwB6YimK9ftQ3tftdY3f0v0lMitN+/nzcFOm0+fBwlp4LTYw6pNu3rTYA+BrvHIZFVL2rcsJfXM3
pzDiHBsxrKJnOLewp+zJdOnlvWVr47N70vaHaVRHGh+xaRmDyQCz0zARMupii8mp++8nfmvRZATx
gMYqjJRt6S0t8ktqXkBJfntfNsdpgrCvvtoxRFTC5MChYuVcPzfxNdw8+QpNNkF4u9QSe+lyUctk
BQh1AYmwNRIoO6QBBgNTMLyPseh4KV+xUnk5j9Jh0GjUIZmZ5LYMJaaeLnLDzOW3NC4NqhU+O1p+
6uPqES3PJ/+tO3THDeLlfTeSA0KNw+kHPWrpUDHN/OAYJ6FxVtggK4LuHY5DdI+XD6TTrReUCB4P
SJ7xf5xfbvnwUkW/Ad0uDaYE5bL5vbwdf9TYxmBtgyn2U1AXi6qUUYYV2ixOSEvcXDmN6W4EsjGv
oSs6DZkLOlRSKwVzLob2mjNzrZ/JlNf8P263L5WPTxSeCE4JKyyQppN8960y+4u6Au0wJ6LVOm9c
nBvnShAgsjsBq2fZa7k1XtsJ+EtoREBMa/N0PWdYBb5QrccXdl8fQ68txybgR+1hPJ3bT194Ot1O
ePgNUidDHhOzRV0qokid58o0SYwBC2ux691dTGPNkHN9ibUm5pX3nj5m4/FsOUtJ4FatPJmnH9dp
eqKa6vkRqVwdDwp9SfSqqrbdLpLZZ6RLEu/1dzHBf4yI+EjBvAgocOhtE5+uOysQ0i8vOP3OWxmY
5zZrVzvH/dA0i6EXgRnfQ3yPP6wh1XO+zjdUI+/Ec+F4uKT368EbRR21VifCJV3BtuZR8cVzwMEL
MHR90uDi2iFuvdzeApKI6wOrUUVkjNNap7x518O5aHAogLug8yYE6MO9/QSbOJzJ5T2OHmBbfVkR
RQQoNlv0vfSczER4kLa8cdAsax49rLtGq8iNE3u/belmnunV5oJb6RcuXfnZdoMusFFFHJmFXZoJ
ZFlRaVs62wPmAp10ggpC90rWYlUPUQ9zh4VJoFqraI7/7+AwdXW1c9xmV8/ZcTb8xP+3Keykz+SM
KgieRxtayD3x19LB0kL5dIF4r2XD1dnovO7MsTopob8URRRFkybM2vJtG7uSSK0ydIplpBqgS7ag
jtPeVLKn0+WUB9gwoxNjgUJgehPlDEFvPJI5TDRTH8uI8Q3U8LLpSS4VJwHFoWDzW4PBGnDjRMUa
AbzpVoVmz0wFBaIWNfN85eC+KfLv2C/W+1yBCvrZh9y2blbLuHXT5c8GA92YTIBdPBHZaJzbJnQv
E/owE112k9EawFColZcm6Ge5Yak8wT3FtDSg/0pKv4kCm9I34BSjGP743nGKX6FkXCZwqyRBitQB
2LC4HPRjbtRSntD/Ghh6q+3B+IkAh2lCr6cveOxFw3FgfH0D/1KiozqIaecpmLJYT4wj5szXHCk9
8xW9dGanpeZzG4GbfAy0j0a8O6e1KS0ZXg+9IPsQdJgqZoYXeG6ezF+DtcjBPaPt46KBnqcuw4l0
DnptiynzPJhEwHuvRbMjmm7S9pDKEm7zCWrT4vZO/CodObj1KUHrmBXYgJ/SujkCUjWYXnfmiPoD
1PVGtqIAQSXTvsQ4tr9AICYGnmak4pYtEhhBovl/rmVSwIwCTbinKZGjHVltQRfY3IXw3q9gJQTt
STjERTXn1DXTHNPt0iSpELfVuLjBNnztgNexNlTa3K5b958nLy8oOIAChhrAf44RDobM1fr/LnKr
vwhKb7duVL4eBZizKBZ3q6Kgob84iXAVbGQ6E4WH3iz6Tz+h6Q1WaZdI3KRxFiCTpv314RR4UX09
1am68sA7e+PmY7sY7C1XhuSiIIR+KKs/4/ZG3HkysSM2kjMOSQCf5GT7Wc/c1Lyfaw4JVaQX0Yrc
Aj93CJjxC9WEtm4ZUbYiOCIoIGen7gbEN7w2dMdiFXY46bS/UPryhMfK/fK4ttX/eAQZJsfSoz1x
OfT2SSrYWNveVTur/6TFIUNxn8uEZQbSC+6lOm7Rhnhi8bYBY4ceADVWhQ/SrkRWz2cPqc94nryk
9mUvd5c57i0Vk8MaF/0Ny6akSAS8KW3sKacuflS4VJSECDH1z1bNRVq00ZJhWhlPkB48S7+b/7Ue
TGbbGQUMa9UPdd5ELb/LikAgjBkKzoggaGylTv9miK94uGH2DdWGboytcVqnXsb7ncsHMMQf7Sr9
ewY6DrWKDsB4vP+S8hmDaNUr9PzmmY20SUwnx5V/Qu6qzh0EIDPjpye5x0R0vNVSetLLPtiY4eRw
VJcvyRW0WOTM9qgJ6KlzaVsq5XMnpmayaHC1qNm633FrB/R1xvCwaw3yhpX1vQAMZgHjQmZ93iHT
xpgMDAkfA9Yqd/xkS/Hu/XL7i3IpRVQ3qrUX11tWx33seo+rtWiA65B5mVaRP4WFFw35FGy4mwfc
iShZlTHlW/3cez7gTJ7YutP2dFuG1DiB7fq6WtbcIpdZh0nNhdYhm8ZIn71NfSvDsKKt9kA8Kdzi
wn6QhYoBxiucxnNRXHOjKGRa7cFsvV6Mo0Hjx7ES6J7GybtQwIYyfTeZjQ0TO1BEVZAftUEDgkIj
8aUjImKTW5oadU6/eL6WiexB3JEpAioCv+vhbGMGTjFM+xCQu4CIIcrzR1uo1NGBjXVjPVIOOFIT
DOJxMuFZ8Yju94ZU2irHaglPW82bokWEraGRMtE3l5U5qnFOYpEQJ05TQ6TIsWRX2a7Wcn3SIHNm
TGIFqyy5ThSCJg+Lo3Vbk78VmKFdyyLKT5MR2ETIsio60CAjEYRsKxUgc9StXO8iwjcZ3MZc2ah7
twMbZ5WqlrHY54zxRzTsiJQ8DbzxS0V1ernMJxdNsgyTZj9jUnAzEmeCyOxTRz4QHgq6457NbRfo
RXrqEfneO1zxNuN6BMYRvKorzobPnTdDkFqLNyPpyQG/b69JnH4jxowWfs/GIcP0gt6dbF4keoCP
u/IqgqeuhWI8ivekZLJI6fSY2QCJMVsD3gaCZyi+7yfOX27e40hf1J8fYc2PbelPvFl1MzRPGN/E
SV+gXaufgvxNp0RBTk66YZC3rFkcaoOGnJBQUh05161cHRQvw1HBxgeRodw6TvkEeR0deEuw6TU8
/olCKn27Vr+5hQxN9LfH2bg9xuyuEj+pcCkN6Nk1TJfwaBN/e/svSs776ERghpnzNZfJSeFR1ksw
tdyRO3P5DxgosyJ43TQqQhcyQVeO+xTJkNT3elDHraS75K3bD3q3oUvE/zeXw/ubxXjBYoKUQtCo
8s3ZsZ6aU+BN79XLrCDhKxMd5LXnX5dI7DYmvZzQB17P9Mmu/EZ1vELksXVqVglBwRlmvvVBbPMY
dTPb44pp4XT68Hm/LImEW+Y0gPWo5xvMPpQoAzwvoTdFcu72QN1weLJVfq1t8dXjX5sokon9RPcn
xd91X1liaLGA8wsGjXbl2yZ145oKSZiIoB0kFItnxbkXoY0g0vsuiE/Tg1s6PPg2KpSzQJUFXgic
YH3ozFtBbcCayDIm/wU4XqY6d63+ie5xVOODdKvOl2+31W7lv2ak+mpyTP6TtUh0PD+bbra/lkdA
GzIkMd3jdGq/GhW73qscQOG4InF7Llxwps75WxDkWUJZv/GpRjWbDmo1MM6oh9utEgbZ5bp4wBJ2
fUVs2mv+U7IJR5DLoxk44mSt0YEi0XkDlwggXcPR+R9i4FgjameXVpWPIbjWbuTZRq19mtTeK90J
16vR+vEN1bOpQ+Vx/JDMGFOqSeTm8vlpm2apE4OEYcz1fh8Oj4bT/7hyc4NCfcHlHfJKHpfzRcjS
KUIx4m1VjXnaeaMKo84xT2gAK+OLTbGFwDAHybQ2dKfA/rohOi7gFo3l/2pNhY3zpQ+5k+TpBHg6
tIH/KtFuGeMRFoRFTqgKxpO9Hu4W0TCkYdLjXbXMybVhs92Nx019knljSRNCAZVU6UvKtu3K3zaR
a4CsLkcPVJkhZVs+xnQ+WWFkiGwIu/9blIQGffhVB6GK+THNLMuqxMDHNqT3m18kpjb6zax9ik6w
OX1nWEujgZrMSE/YsagS+bMplE0Wh5M7uW5KEnHaeTJoNN/1ZUWFKpiU4KA3VvTAh+gNqU6beLc6
9WxC86IlIjiv1e3dCEe6iN/HId2CzzNgvUyfUD5Ay25UgA1pByFzKAUP0WrUMng6Pe9i1ES2kly3
Z7hFt/o9kWfuvr37rFZWtH5JrUmpqjHAIWvCYjkzj5WxhDm1D+hfWWt49lWp1UPZtebJddupilUy
MA+Y4QFjsq7bcOcgwfRdbHDOh3C0R0FlEfbHiOa0tz1vB5dugdlXDkElkavfpaI41bUBcqiJXpi7
RQUPozd7Nf05pbtmzGgHJCnhzgEB1egdBrsBKfsyT32sU4q5dU/WV2ASlnpnWI38VKQltmDIrfod
MVPHnrN28634sbgUKxaPY2u4UtEpI/Nm4CT2WK3JjiA0tLNhwV2SI7QTnfsa98HSUVlvyWzwaI8z
qeEjmJ3SYnYNorwmPGUFA002iKL//KLtGzJmSBi8tS9FljKmP3WrHfmZn06qvjRPiU6ePMM+eMyk
vQsF1om9Ua9XiUKh/VKGvgH+etCe/S24AnZ/AvTdUbkq+AdtZCQCY++qD82qOOaMDLpeUk3krcq1
jXtDKXVwavPFrmPAxIJQ6pLLggaVJA6TKAWrYDJ1hzfeKl17ArcCoD4gpxQtpTeAZm5E7TqNvC9H
hu6eweC1EpDCEMDMVV6rX5opZE9rX9hz6UQt3UT9auCwbQRcxYl9bNOPkDVu4fIG65gnrcd3uSIn
M7UKItdLT9tnGTzHmkA7aceI0b8nbnXRHJwIxG5UICxUPU1BFMmZCIWUWu2Z8YaxzkvZ4jzkGmb5
HjwUMkIZ3KTXadNNvphCSmN433sxDsrRhnC4Rem8xMCoNYJuw4NTMMlVnjwo217PWd9rOHnw8LFd
HHJf1Swlf4xk/f4ijk8LtHuhYIJY1R8slYCSPM3GtlhVHjrWPxMdj3Gp8nDJPUUAdGLwgvGAnUWE
tW+i4OS3NP35F9IfY+YSPsAdgUilzHmV3R2WTYlDB+qpqz/UplS3EnmHv4uFTMWf+xW3FliTjHkj
Dce2R/Dyy1bTIgjv97RGJXr/MU+JL7ii+UzI5skoln6gSLKRuXz6Uh81G76kXOsRJBQqrMz1SNEu
mm1HHQtFJVWISzCS5HKq//o5Z7TnDm42dxHbF4YdcblXur8XubuXpp8TA3yPyMOomEgvzB8yD1hz
BLm/Yah1v5tWorR4MMUUekhv+qy48roZU+GaP2VIu8MIfJ2MHkbt7DltZ6Re6eE9dRtTsUwePODs
ejVGQbVfHhlczJsgT6Q/6dV5kFI/7DlDUjOVnh2Q4LrF0E1T30fzE+kVz4JnD3oASQmvEb6H2Xz0
5EEJHhWB7aUkesCGwbBafE9y0ui29EqGmzu+NEf8OGlbc6DqJO38JzlhrcjeeNbGP8f0sW+EziI8
NebHJg5DFqp5rOha0nBLFYO0RpuLWi5GAOXaDPX6/cFANmqqsvDxQ2LTyStS2Zz5Ah39RhfnfnBf
e5oneLJqNX5NuJc+eP76JzVlim3UpUlCV2OP0GqkMYHj44ilGzoSJNpNP+uZ7B9RQKWmd+QGsUo5
KraZd6YPHu070BVp3DjB1ODF3uC1pmAEQYRtCR/0kP6adFfQIFzgpvjW6ERAnKhcfzjwecwA8OMM
1OFZQmB2UAHv7daZdgx7wCHmxRNL7cQ6J2pFxZcfcoAV8l82wlhjyefJgIWm4ik7MhfOecQ77MJl
don7l+GFI/OZSReNl0R1PskpUg280FRpUMWa709gqvwJsfM47MU7IMqQsGwPEmguAXaVbO+ybFrD
mfmCZm/LOd+v7Lpoq1clQf9PSeZoGcpoeMoHXS1VBXT9w7xDgFjpw0nz+sECWQELng0+nvnUDU+9
IOn/HfU02mbnT2jWUgC8s/6JaZwwVvTIU2CXCxn6VLE3JKnKmrG5Y9x+fDCwv0nVzLibLacA5Idg
VGSnQadFvVk3RaJdWue9M787IX31pAjuL+vhOIlCDoiTN+kzXCCpAH4UFmYeaKgXpwU+Q4pO1Y+S
UBLS92s1ftH2XPVs97mc7U4ORX1H2j5RSNWwt/MX/xGOTIgWwOWt1VfJwGHIOsZdOcBYdA4hiJPO
EtFzXcw2oX/3ij+xA9JJM5I6zQJrEZIwgsuNWM+3Mw952Im75fb+xKFXFVlPxQIOuBlTZlJTOAdN
K1WgI3mA2lw76RHofHN/nOvQw9Q/buOYHhtNc7QMM3IZrcl8fqdrzJNyV72LNUIny8g4drBfiKSR
EuBM1BE+rzOMGxLu6ao5BqNj+8OIXiSrZnkx2/ZSTS4sMMIoNmgM0QYsnqH0EUgO/vd7asb2wsUh
6a5IoaiW0BhV+TleXcqIcdkw5Odal7vhin0uQrybjxayA+KbItvkfyHTgwmpqKvdhbhM2U3pW2Fy
u0s7irOLTNNlMa5KYD/UZ2o1vEadREmMSC0yimTtA1vct940yVsnR5yQtBKKoihavNVbdYs2Mw+D
t/r0HviU0v1tRokXDqhi/8g7T1psUlfL5GKzwyzPSNNexrCf4PhagA22QA4Xd7Nc2q7QE/7aRPSM
3fqb0CV9q3MUAqN75TsXFgT5sxuJIgnfleHIZQo3zjeOjl70FWbUUWGgwZPpYSJdsof85Hg9t4o1
cA7K9kX88w8qNn1lGLXCWG92+r8kea1Fpxf9/+cjAesExaJVgSNaSJSTyek9bd4JTAAojKT5jjNG
OjXKIwb4cGum2c39gPikrQpGH3fF83esZu5CN/22BNrg38pahX3TuThc99LRC3Yt3tJl2t8Q7Wmk
nT1ZQaPIHxFA9Y8m5VG9if0ZQrEfp3WYknUslyY6XZHtuH3ST6FJfpheAx9JKcYS05vl6/d0ycET
fBbFtL33Qfd+Uxd8dtYnMcpBs9+UWIQHsFKkhBEVmt57XtNHoFumcojbt4VWA8ehgO9+uGfxs95c
Fs3QRBE1QE8ppNfbLg+eroZmjcJ9mzLsm+8phCDXCu7ObBHZsgXqhYuKeZVRm7CpUDcADhz93mBS
S+vUx6XCde1GEVuTrJSqk+WRp0ntDm2pNF9gNaUG7XAU39A6TBlihv8EVh/AJzZTm9lMEE1JW131
I0hX95UEY4mWmAA3h9/JjEVChHTpsebQ0G5p6XBEcJKsIHx8OlpNrUTSME+B1V3Ct+XMj2BftIk+
M/ntYM8HCnrx4FuUae/QzxihwrJaI0YO8tyVS9dcHm7awCHI9wupfYwgHUGrxEpElSokSEHCBIw8
M/8KxtKekRF3KZwD/yKubRjNkJYfJGZD+hthLUZB9mEajjXmLgiGBOrvkB/NAMXM0/ec8ytnJUst
zfR76oHNN00wsnBOhDlOArBUdFKEZ1H0vwM1gec/w84WdA3jXK9hQcf5zi+O4G5jeIXyCdkAKXVW
l7LQ8Y9Q7z4XPcSt08F9MNpmm+JU5XCSQD8yAYr1MPk72ULRkwjMkEVIjmirUzXOvjfkU9pE+mLH
FzKYjbHBrbWox58PZXNQxUoRwcwvptve+Nqkk1iraR9xCZtE6k4kjeZJl5vVtmXkhBOO/GI5HBXB
b7H0yjds4qlNMhO13NQNsKQyrSX0dLDJPascL6ent2Cdr22R7Wz/a6/y4YWXeEpcg36M7gLkzs6G
3wAfoHG5vrbWEYVBw6Gg99F9gkL79Td1oDCm46RStLeJxCZiFZqftrZwXIHhdvWSVwkEHckHN5Zb
oREkAicYwUHWuxTSIwPN0ebF4jKnmVRkG5to0DsjSUfF3V4g8q0lWuZhg2zzUY+KdYcQ2VW84/hj
hgMArT+SdrdugZwb8ektsB9bVSV7j0umTzPuDUhnniOxAuNXzHtCNQIjrdwNwcVSbUjzcVWMHCtK
/4ajO3b4GZc4EirNWNvBOFAm8dXn5Omq4GEssY0nYrShCzwcp6dLev4G8bNNDhewMS6xa3xc0heV
1G1VWvGGHp45a1j2OGY/2S1TTzOZk+vMvIFx2ftnhe6gRw9Hw/cSd7QMaVf3iM4Ce2iAKBrdkrWv
LP9wQbjtTRz7sbfZv9vcNHNRxn993dGDkeE83JS1cZiY30qz4pnkhcCgLD2bp5tElm0felzmAeNd
TBIwii9drzSI0bvY7nl3IOiWlC0V1HA4TFb8wtUSGtJU4F9MPGfaIE8FNSwKCi2SXtnZFFudc1at
lPJ1hxPhQZZADjKT7kNGmvpY6KtiUovdUQoMjhYdt4sIexr45RDUcCpW299gBHCkShKweCmKm66n
MJQb8uV38DiCOs1LCdRbqDo/fxxcUpLAjrfCesKyMUdT+S4rmqN2IVlKMfLjjfjtuVoz6BpnacLn
GPjKiAnj2chKlfGdkfLwp2RJe0xISYtp+1MaUffrKVf6Dckbv1adsldXbFtBYWFZgPo9YqX9ed88
jjQrpK3Xw66dylBAExvRfZx2RzWeVzp6mrJJ3Pz6PS3KCkpuYFXidY3aOlG2ZEpw4ZQ/0WTjBQsA
7KuJMVj0aW1RdgOdtDhzryvhkwOZjMHqoN22Y9B86LP8jmZwAWRHMOeM3fDkAnqcyr20QO1ENsEN
y8fvYvovdlKmuNijdbQMhtEP5dQO/0j94tyl98x89QdqAAGgPEEfV3FCnHAMQ0nlEl3Mby/ER1to
xdxFxfconlDVIA0cFtU+Re4qdLJGjGcUGp2XXP4eRbzBvEXENqZtymdo1ndMNVmGdNSNGuS5fZ9Z
VtIIyHWyHYaYx+5djzAKhxt9xL5rNRXAURy03sqrcaVEDVscRDxNSEvVFcfeU4chz9bjnLcnUQbS
gKt8r6ZQ8OQlxKnjyoPLEm5KrV3Kk9fgzthK2W8zIfWG8QeZzyzNS1pJ+w9FMrF57ZvOA3urqvPY
9J9XYkIpijJqhCJX6+VxN6jWZwWtcX3TKVXR/J0S+W9+b33h0oE+JkrDjhqqozo0g2Xz70n+gBfL
SEbmuDg08bRJEjkJifyiGuhs63T3vutKmFk5pvHftSJ8e2p4FRHQRd6m1dCeGkRCCcZO4AFjggkm
/olsFFohDGGiUy5EnapIlDkCQy74pT4MFO9l7eeurm1f/Gx00RYhiC14B2bGcKBq2xK527/xAUcy
bZ440jwvKup7TpYy+xpRuk2mAFxEl+3G27g6QuA7+iO6oNzQgrtSaaKei8DoEhWa1mgYPQmnVsXC
X7iQbRIVeQZ15Ar/L5DqoAopMhboo9EflJrfh4+/JwrCr75jczF0NNM5A+ZdW3IBGQ7mJUxLvswF
U4jSbHYpSB7BD0B/fFs4DwozS3ksKFnWXArSXX+arfWyK+JdoyKEBT2sqpHOMFg5BwWLBFENjpED
JgIRuGGbh7wlX1ptOrymwzYoE8qme2XeUrNnJHq5YKjV1bSkyuq4DsuYKMdyKZ/33JLMBrIWg/hW
QvsPuGTwRBg5tbvRpi2F+vV7vy2x5qFcXPZ3cWnrhVxLYYjA2P9lbt7I96YJ45A6Efkzb+lDMt7/
x85+QUDk8KLaWT7eDsQcTjI9r2/zZFGiwshJ8mR5jjlE6yc/H4FfKg2/8wM7U5xfJ8mx2iF1YpjQ
Y4Cei1PdPMAWQhCqUBIziw+NXe67vUklR7LMOpwSfDKJp2mdSg968IXeWcCgOnWQUlabbZnpUwZH
e2IX3hL525SlNh5qHrHb4dqVXK0l0PdKmOjjVysXcXEVgzqt3+Oa0vbf03E0GkFkjNnlivyi9F9B
+Zl9UplRPtHH50QUwjiG/dcK85ZqJRot83gHqDJ2jxOt4j/PGTpDuOfjRXF2ye3vgOVHqqdVThJj
l18WkJ67d2ejduAUOAFN20UGy8ZVnhLWo/MBc5hoLhOhGlVHOEKvbiTV+VTxNghYRJrHtic4RTQ2
dcrlvLxt9QphCtkb0sb9SHhWVBSdtBk6hIjVhRwNRUebVRvghUaNO6ORGRj7lAyqn8Hj2xfJIcxL
8Aj6UgAk0qV6uEmCNQaGPjyhfXUgOjWFbXF5pA0cEkPf7C0U8350qOW+YNv8YVkcs5/BNiOc6RY2
1DU2sa6w4GeCnQrz8XZX5Q0vTOO5sQWmRhZYjGQT5P1EQiZjLKpUgi6qsxY97mlfsIrD05cN11ZA
9ZmlvFHwS0DzR8mlBaEHrD/PXdqoDHWsnk7ENFcriM+9dMGnQeHVnfNJTldHnqD+N2dilw8shGcw
oW4+4CIxw+/r26mXOy4YPxdS00tjILHZpdskcl2AVoccVlLnF6yjH7jERDGIpvN08K6GGd1aIQ/d
/gU8kRy0CcDg6sG0NB7gXafWKDtqX5PdNstcIGaelu56cJfdNi71XWeOjRd74l0m0xQHHSFqn2p3
OHrCEk4KfzZA7h7h+fln+AhZBXmj5pPt/UeABrEClHQBq4+N1pt3zblxOQxgPTWMPRCmzcQdKkAr
6PQQvvzkQFVqJLalOFkuUGKyZYBT6Q48vuRJMxwALr+EQL1+F2xjPO7Eu4W+ZrkJCuqa9Pt+uJ3E
GB+Oi7kFoFadYsDgY08/ZTkAMenkmwXjA46LhuQx4ZXIWZru+Pv8a/YoMK6QM9DuCIhRdMZoHKs3
5qvkVv+S8Vy52V+MKFRdNHHqHH3U3nmC25X5X+n0iOwoRHHmiUJ1aHmVeIpr3nuh4vbLQ9sUj9XX
uuS8dDsk0lftEXcQ/fMpUYXEJEhj0IuT0lXeG3+gqUY90KIefvgFCbdodObVMODe6OFbns2ioCM9
nvSO3IbbUPNJxtskVF40t/ZvwfzLiywJ2hxLsYYep9U+kNk0/Y4saDcQBybFWjK5jNUFdHZSwWQs
TkpNp7q/j60dUx2682xSU+hZL1zFGjyKHOdNOwnN+HeAi2HErDJs28SBGtCQOm6bfmqWPKufkPa/
sq27aP4nXmYsox0mxVLFDCK0xZ5I3NalEAtg9AWTL8uxx0ht5lpytInF5BlhYD4/Wvl4yTQMMxDg
hA3KhWFm0lOpHG4icgX8P2aqZXfkXP0/fYkAmC/C1kbDNDk1N+1yv/KctZxYO3/SHHYUVRsaVvtb
n43qiYLcLQAHntUTDR23Y9V8Bi9UpBFGc4GULv4b6K2bVQgJujTY2u/c9iJQh4a8x1P9B4sNZD97
omGXktr5sQHO/m5wbArcpS0x9v6V/DvbqaTtvMG/gObeYGI44bNVBjHUB9xmzsJm+r/MwK6BtTf1
ig5qdvJPvC/o3yGKsyB5N40DXq8+pzu9U1Sx8NiYoevhJb/KnoFyNdT/aA2k/Ly0Ea34IPUPO/JD
EcoAdskOJmkb2bsP7QR0T/al0Iphm4MPy05RcOWrtA/MbcUg9UMiMuPAyjbMiTZafrAbmF+uFarT
3IqpiMy7XvD7ZT7ID4UaaS3dgOYDnGfSsvDppm/92XDVWsWkCPCnzVYTpmSbbAtKo0Nbh7PhAE4J
d9mbI2lz+tD9qsHKmFeFafhUi0mzaQJ3IY468TRCgZbaStl4d1gV93OSTNA6a6IpWireaxoecea3
LnVlHZVnFELYtHmrjdkOur/pSyfaS110iVxnleFYA0ZsokIs+QLuTmaFDTY/ebWZR0qp9pcina0A
Dh6nlBiFxOK710sRyv0cp4v0kHalANc70/GeJfV2OhzJONZFKj6tUuLjk2xQ6cIQywdJmcOTcGO6
sTl0OcedYQ367no08CwClgiut5BMsPOsmc1u7o5MCeCxgD55dzIh67Y1VB5hqIDJEnJ2CkMUm0cR
PVb55Oh1NJ5PF85YYBgp9FlVulkwM1scGakTS60dANj4pR0eaO7LXGdMf+KY/5bIrZxIY9TZuNe5
26aJVXmIeYquvOS0eUymbx8Vxdv8nggXL7zYMZ2HhWMztqZkPoazeo8Wq/Z+F7AtbkBbGsSJ56SE
FCRS5WCq1Oe12+Dpo00i5lHZIp8EM5IQXj6CDrLCNYxhxXwHOeWmSYwIJaeYMLZizYzu5H6m6nSz
mxs+8GguumDjb13Qm7uGzPfrjptBbcM2DR9mDbMwpQT2TPwt1n5lmGVKArzgfnL/ZRq88dTgYumo
clK0dW8TowM2o6bV5TfEi5Em439HIBxr6+Wh63e5HSKMW4P8c8ueGAtwIdegOHhNykhUNjWlWpwm
i91C4Ip3QwCYMPCUFdVqLNrHU424XPrwZDWIwAoLn1js2aP7CwEU9qtq+Yxp2C7vQJekHj5QbSuD
KCuizDzRLyHPbKeuViSJKKiYjRVdDBBAVQr/A4uQZ7Cvj3VeYaNO0g4Pvh/Va/nun+eBfq/r+UYm
1hasfbWydLPc7srp+dsuuI4rVAfOYlINjt3hm64UxnIJd/uj418rBK+9p+DpPvAZB6ZPaFC7ZlQC
ldWq7udSDKxH34P/gfUw1avkKt3jw/asWv3EOswsnp5gWf8kI89Mcs/4JCiISPffgkCe4hMC6LGR
3peWVkyFBGkufqEQrGe30/igDR2wCU7tYYBXE1oZRZSnKIxG3Hm2myvVYBQ+ZToEIbTzBe0QZRCF
bWFsVkZ9wUfAI5DleYYDLP6KNdl2rB75+RQvfWYDgpNaOUrnQh0b36cRrvX0VI5Jz6PB46DmHfzM
nmVLatz2STlYN7aT8gEavDkoSZK94bIizbtW9Wz+8k2GQWHUuLDkj5OaOmf/qP5xFuw/2r8lWNMs
Vl4p6nBqlk9OgP/ZV36s1bxNV4/NUCBpZMAJU7hqa7Ie/2DN0pHKxLbCotKKTmwKKYH9JkC/I7Oc
w25bye1VAPzMfNYvPIUBxTYfjlIM1Ae/FFgvyvQ09014EBK5K69OAaJ3CzOdQw+nkjXsg/+ZtujY
JhF/sZ0Bv9hJiAvvV28fr0ow0Z2iT6rqEEC2GT+FQjlMZPKAe6G4ZMz749jQ9JT3BNZ97h5EO96H
XUkbTOtZUqbCTPPDt8672IC72VdssBrxBNfLpu1jGV8WJ0cU/YajqGMXktnMFb3xtiMm60Vg2Jjy
tCKcu3umhwU3u9c12LWcw+xydikcxg4dO36R6mTnHA6eF46Q8TWp9UVBk6nvksoOS2RSrdsXWuCn
Rg8pyfhhKEjkrOBlENar2v+t1XLEdE2JUgm4Y4VGDuiiSYqcsDZEZkVpDBf2pSIEYXiJpa2l0VN0
ms127Lq34ZP8bITqmD4Yho0RWILtPQgN+V7+uwiM98NC+nEzJ/8ZSfResdI0GPjhwf3baEe4o3A+
u3/d1fGhqOsmkojU1+xc0hxHErvycZ3O208425wG7PfOxuRcMPEvFfK+ZFerk8IJmBBuYAX/jqe3
ATU4WA0RdlqnT+HBCdwvkGsUJMXhhQaikl0Lg0TnMwLOvy21SPRzXo8cCARWuWvbLLebp6Zia/Zj
lyrb79Cu5NyOEg/aPSzgqh9Ht2cyCg3xKijCi1CgkIIv4qQmg/dijjcJ0WnW+F42RRXlql9/un+r
Xgq56U0X6id4qRHD/Ha4yFOISw8p8e7Bs8PUeLO0DWj2ZdKkU2flDEWKOYJcrd9GlHlZjbc5ZNQ7
i0YV03aq8GBOUMfF1uUh05KBlgYcrLYr0tZ9zamEKr/JL1o3fFcxXh2YEFSwgJ0jZUqlL63i05tB
cEkf1VOKRjhAFY52qmarcDFlaIoTycxMUAmBYjwe2wOItTbQgkYb8k27CZs0GO5gnU/t/rbUXRoY
ha7HzoAfGtaIt6j29M4KrZTZlGsMyySbSdo/cPKCtws4OgadeQsYaoE8E85o//pgOnMy9gZaurTU
bpPXVNHwfsmS9fMxAN6nIdwOv8qcap2tzQAnjSmfs8cOB7Gg376sXNFePZpRr/cCZZ6/lI5htRmt
nkgwdASk+i66a5MtTOOtLI5EgJkXcOPGyUnTC56SrVBNhm4VG/0ckBqZEKhG3NWkck3yp4NFMde3
C2LfYX8zkLhoKHmayeE10syliL0dZl70JjzFr9vcnX0hSofIMCjz0X2M9ZRChqCgBvpDosaRiM5D
aW1A/avo8RkrpcQZC/KTgwGenprB/hXBrsUQaciKmmksXEKT9ADqwNu/WROo4zmnq9GslxWn9O/G
jikGPlWn2euBNs+JYELqFpPzz8AXySmtVlPXFzc17Q/O+Qmo5hYihjv5ujryYr35PmvVkO92/lFA
/PgJi0choiON/qD91NCqtMfdDGQcqwZGvV84RBaOEQ9DQc8OPHO6ESrI27HKkkhMpn1K3Itezfzd
jE6w7pMpXH5EXUIkWx1AvOehZ1w60Csf12HTjzPjmI1rrURpv1Ot2ze22SmIqZuV4SR1Eu2SbWrg
ZZCBIlVByLqWPSm92INDqS8L2g+KDCK4prZRhz9nVbYfQh+UPeyUx0ksCcjXMYNVJ4NM3vlAmz5x
fzc0CnFJN7tQbHyBjv4szgZAs+obGxXy5PQ/sKl+E/74vN7eQkmPgMeL3DzT2FuL2llt2iEYi6gY
8VXTPfCpTjSkUCZCK4ie4lqVkdoz2djI4y0FE3FBHMCG3J1Pk9uaa1+DQ3ohQ0XjRoXF/sL0GPgX
0VmvONP8Mxaj2bV/pZQlnpGoEbvt032H+lRbxn6lP+iVjvlWOHaJHSpnq7z5GZC2DElOb1NSUX1d
Qwre9LsVSwOABoOcuL60nNroyuZcsN4c/VZJDbUwyhtZCYMvt99dEoRhChTtBdXnRV82MP5MNdG5
zP1OrnFrRfgXIfkk1tNLwC0XV9CyN+dzrYRpaM2kzg9La28XaNQbluUpFBO0J0F5zeoMqUbagDoD
061bd+PVbJ6nOuc/2svGbvE4GUU5g9QySrFIgoTvaxzRVNTuEgfpjuaGwWo5NL7OJBYS/8dgeRon
yCKwZO4qqXj1pY16VZFFB2c71ePvqYjD5PKSlkdqN8/52Dz43N0ejhMxe4cd4khAY0/gwwl3HHfW
Rmg6nN3i8Qw/V89GKBrK5Wz4fmpWSVI5unCTTo7nuaHWIxzp4utR/jbi/uxJzIfXaM1umDYIrTKd
RLiIey+hSsEvnaABMXgYnJAPVFpYnqU+X6JyWf2rpelmnb+G2cWVu/Amdg8E3ugLUvb3aa7oRvwy
Al0EzSFmNgpce184pLPw0MUHi9Ke7nCIHLz4P8Bo9y+KCcpCgp7GF9oXmiDumLl2KbQNfrpozND3
O5Nrpl1cUB0uQ/Tfla5g1NTUoB40H+jMuqbuSpqYpdmXlIAui1C3U0CBebrSz77u2EgXRCkc7FnD
n320fQQviOf2yZfX8uSo92Q4rhUTJ2316WdVXsNrGyXRnv9b2RxEj9vaGN4LyIlh1x3NH5AcQxnc
85oD53SZoOUqKcBxiZSK0ZAo2HrrBT4rK1hCUoGMNlEPe6gVEQaE1+h7LAXRyXLBar2mA6kl1WII
gapZDizsgvB3hb620lZbxBUhBedP9YC5EW2C9rsLzg/jTLHIZyx1yvdSWr3jtbtubpkiqAb2MLW8
q2AOuFHYREqvzlgOqfCf1iQ0NoouDjh4HqBFVgX7zpH1ptcTPOQCx37WxO3HkAUpzOwOfw3ICpKP
VFK6JdChp2QkmmgNwtn7M13dWAExog0X3W8DZYJeDlyDkq6/TAbV6XjL2fy8JuVP6PRxzBeHQJyK
MaNYRA7CuqH3Z1goBoK+aQKkQ2Hs5JgTPlipv+zA2A00PZibF6NiOxvoKgoTK+ZjGN7jrq4Rtt8Z
zMUgFw795ZCC4LHSx2eyCnTK7991a9to4uZTQ3bCRid7NvdypxSNquPwitTff6UxSTLO8Q+IpX1I
mSK7q0qOb+gn498VlR8cFwK/CsqEmAqLS/aUH3wA4fn8/zcg13qRLqcKdgFKdEIThYJ6QpWkc1TM
sWiYHEBNdiGfGkbbS6xrjCOdZqAyRAhyMljJCFZQVPdsd+4W45dVtSM5h3L6EqBHFxzLuG7/YBIw
bH0mxMbiHei7MWaIGPWHG5T1ITfgopfFkboQgBrwX+9MAiotluPOqm8N1EtpEpjKmdeFdRwFGx8z
ceA6kLUUHUy0JMRGSOtg+M133PqudoeE6TfXstSzkZcUbGyWX/mJPPaLYBfz630l4zzA9wnRzTa+
3aNdc3zbyyqNuD25kb523EEt55z20T002n4aXnoJH8Kno687NF6daBAcyewck9iKzQ5nOHvu8gr2
gkVk8NlXBDMsLgLmZ7kKKVMjbm18zq3HXIP63dI2cqLDPKH+m+H+mGPnVP3ur7RO0/KXKGrNn0oF
yXb2jnkgsA6DX1RgI8dWntcQdiYWsTHErllouGbuQau725PBf8zpu4wnrOovl6aQEhzy6vxOMT9p
FDTddL/4vFQGxzMuVNYoirkBkEGgA9q3X4sgkNMeahrerynjeGEBH8AUzXTmFhx8EQ/zKTsdMQhx
NYCSAoxLYzDej9v+LQNxPQtYewEFq7CYo+aY5o11sCDxrI0pNln2XBxzTzke7I/yNKXf4LN1+5d8
zEKx+nXc4yvGc7FtJJBZlsKpVBzdoMwwvMHxkU6pJ+++rh+hlHHkdNe3Ro6V+DoMGeZE4nrExNoE
Yk/56QfuulBdNOY7xF3ZlIll3IM2rukCF0KhXeNWvZF7p8eFSstWzVHQhQ02ga6CI0de6P4QkcGU
lwrdLUTfWlUtNo0Hbvqqu2DGg1b6nR96OpftSDA9t1bbqunix4ddXHAkOqX8PYV90X3WMCdUhq4b
SQWr1zNFvDKi54aNYusqZvE6pQsXyt4GvSceTfPEHe9m3yTkekbe0yfpRxFg9lZgZto2lNujUl8O
FHD4F1KDHKloXEIWCBuuiPGLiHThPPwgQEIIYMIaCqRae4G9dmK9mkri+tHUkOwwTzo1F7tJQ5RQ
AUVzYo2GM0Y/hBTN2xc3Bca5aq4wJXm5CTu1ELh5InsxUeF+lUayLrYAmK2EXFciI5dIOxdwceOy
SVYvZKokU+z477VcWGSsLCLcIJ5EtWXiMXXCkUN7J9UdPAcdZI+l1K8l4Exbm+5FAuj7vA6JDAMO
PfV1vBkS8iR8wFWhauZtQzK3Bvp/76P91W5i1OFlWGSqeTTuMEkq4dybkIwj1JGsIKbGOkScItNi
oBfMcXaZpbRf3yjpYM3tLSzykNIdsyPl2JJ0AhMkI78FYCTwiDB/IMz4UN/MNqrf2TpdSBTVJuVu
UE+MTEdEgm+U5MvneB+7DxxF/DdIHaHXQynkKChbrRI5OvFMVjJlx0gqzSFqtnXPUsVsW3Yk33pG
2i8vSwuDWCwq+iFKR/x1uf+58VY6AcATTIz+Co9zOiEzGwsmcvn+nw5+UpCRTWVhLqzwWGSQKAOr
2ntc189DES4nFSkbMeRNDVE922hbMPc88Qo8ujCmj92kiId5sbf47rfJ9+k06p+aL9jmQ0LiiPOL
Nf3NIOHpjLVTFV1G81z1xpofyimEBAHRZgl6hD1nfNJ8vvuwJnkiFu7/ZL1FTZvVv63gWheBgA8A
EHX6FPWvBqmBCQKVEb0S/63BM63p4dC9MASo8LFJ1uHAAU66oFflpyAYzeZ4QJ5bLrJepg12dDQF
xb+7jGRWZyDCCTbfxpkxxPnR6aQi4BRibGssCyw/7t2rfwlCEBiWCozAvpJ7FX6l4TsZqiT7z8Ap
ZeD7nne1qMZPj7u+HHqWiClNgNe7qf3CIxnhJLOFEgwupIOxK7EFH9m365dYRuTvQDAsTQiMLzJC
r4nXfg95zmBXCvUxKafnoNwi+1AxcjjJ9QRFoGmogaLLbMlwzJUHp0PPRFsltgfMSmEFjsaOVDmh
ioKg6Y1bBoi8cU9BqWK5aHSv6VdLdsF2q0tiEh865hhFRRF3N1dlh2bgkyx/UHAz19De8RWb54vP
Y+PvMmxB+aMTa00V4tHa5N4L+EbV5EDKvlhQgUduPIntrrHMhxiz6Jk9QP6WAzEfHnH/ArSq8sPc
md0H+qEKrr3Zfm9euem4cZB350AmqoMp4sqHs2h3MK37j2Gc06vUiclADbh/WFKQ5FGuhkQE7pz6
Alb0M2evDwwOhOPzi0LQbSZYtyGh0L6d3DYdEHwDR+VUh9ZoC9IpS2A9CjXUIMBRFfVztnp95TKm
DYrngjuc6zv+OLoWh7n+jyseHoLKv2ZTI+u4WYeVVej5vwS5MYlc7V4bKYo39t63EUcg/IrN8wEr
xx4z6VF7J2OuHlF2Di1nvadcZGe4kdfKiFt1ZD76xFnrqDyD3WmL7CDG5fqeN43geqc6vABAo+90
uk45itqdVRwOdcT13FfHNqRMCyVE1V5ykz3qbtCOmgHptccbGTzZSvfOh+BYPTtp2FDcReFqZ4nw
JmhKA85MwYCAsE7Y6JnM2XsaM0f2wjFISniwzOdBnlqA4TlwVg45SVKuNo2emzt3XguKuctnh01x
ucUkrOoHmwjj5lWTEE46ZaQfBBxv8/DE1fH33zqbhKqBj4vINMInDt17XE7ku6icda4tLwXWaU6c
da6zjSuwNDTvdBOWDjXopCa3bP3WzhZhiXPGzQA5q3BY7LDL6mMx/odsUbFo45M2uT5mJSL6piSZ
vIeOe/It3INYcsgGGiBQ9qMwPUg96oAf1vnd4xVzPYba5NrUzhwRwnuyXlFdNNhHfIAQMRyMLvu/
3qvfEJZOX5Lh9g4RhdaEFnwupWmsx5ylv81O3Q7LpcT7L3T24FntDXme8ZdFNViYrDaQpVXrCiZS
Md+Zmz6wkl1aY5vwOy2RfQus54htCJdx4gItQl6lkmunz5OgxW2Bz1kzDIDISBUF24N1mLQuP9sn
7N7t9QyvDlxwqXvX49Sw1p2i6/5r+lFMoN2dx2ByZZ95ALtllcqXGQI0tI/+0lTzNRzxI2WYyyQ8
1Z5VWSI3r5B/U4kIfL/dN52lZO9FICX9UymRxcMO+Li0y7rupgrFOwSRIsjQpnCCDJhkGO8cZgeG
ZRu1vyyRYxip+xEJW0Ub+4NX6oA1j25rTx3sMDXpG+az/tFqHWtE6uEwWNRYjvmhO+AuEwsAOYSK
QnFntcfP7zEKKdwFYIJhoJHGLMTV8yeg0VYPUZ93p81kW0ZtbKQHj6pZGG06frlu6B2/kpGApPYI
tap8HAmH4Y2wRNW/IuZSWgELfiIL1rcSgVn3LSmrIep96f/wXCUBjKZhevBeEw1sJuk5ZohkY/LI
PxLYeOVQJzUCmaZdSJw9BJ20i6CsLEcauU8KNNk8zmvBzxDvn9hkBKxV5/Fcot7Tnl4woHTymvUv
nifiW1uuPkvk2FjGUvzOP55uicXWx0kxVLNbPBQVWvk3wvhOu5z9szRMtLOqlFMSkS+Dc6SOsaeP
yZbkouKE7VE+tE8lDVquCLFGDRj8orU1Vvb6GFEVKtZKs1cwuV266+sUzOx2VjRwxT6aDs2vPQcT
DEqFqFKYmnYPcTZTvgvsMRfbUVlFcMV0SM35yYQGUkOgpTuQdS5aioIdCVanKvjf6wN5TtRxIO43
J2qE5FP6WytwhCzQJ3gKfG45Mo+BxviKGm3IBd3cu2OB5g9sjEey6JRR88lvChmJJxXyZGVaiohH
LH65SMKyKK4rdVbwNndwsjcegPARG7+VjTuVT8gbOvNUjRFMEE5ArrJQM8eIY93zBR69+YfPE9/p
kRJm3uAALQku3QIYbU/LD0wPzgUbZvGWyR/ZVT+cTbu/l+xtAunqultAx9V3laJ2ZmvU8inXYR1X
1HUqJEkpV4kYv/bz1K6stdrRLb/v+EWYPB+AQZDjtSb3OBS/XyCf8PXFPXtgHjfqdkwdP3JACu5l
MvNmnCHPriUtYUzFG3+wjlX59BHJ4IG4cP1WuCAtiWHxCzdhnFODQPtWHCw/G2bO7A6Bzvf3qYFN
CmKcc4K1b1+sy1ziL3oY/DhjM2PrvYB7LXRuoHO6Gf6yQrK5ptH1xX8LKfpIxRwKiaVbSPBXVo8u
1AnG9Nh2hsb5xcfQ5/gg27xqWBq4K0vlJ6pQ2aQKmkFNpJ2GSgx6aQCgTLJbhYk35U6vfDdj/v6Y
eGj7tAV2hE2p83KRVFtYCaeshsvQp5aYOl/ANyWvJTVAjMB7XkLKc2SKgpJyCl5ipxZ/isP9JDr8
yIu8y5MUK8YUSgLcomEzLCpqpCUTnosbaDFxEOQX3IP51kI88EP16cFmBy2ehiSxLsV61ByuwNHA
en0AxtpwpnOeoWG1RVEd7AdJ8tLLoggCvVljpMs6SAotEgUJd4/ZxCr8nthnOQGMiEunc9vIBJ3K
sHrAkwul61DGDP4kJ38/TnIkAXMpzPtn27jzb+94+3Pzw3EvxS7l3yRTdkezyH2ZGsGYmsFe1PEv
z8cirpmTAFoVEBAmXmpDGYeIFpPGN27YIPpOWoBJ7kLFGNuTKmfHhxHy+bwpM8cS0PD0RasIvaNI
leRbiMcL6YvGtTWGGY0HVwhJl0pRP9w/41p3Ft8c6bheAOzg0md1/AuQxcn7GdjU/ut7K23w6wxX
cZ3TMjFXNo+iPTILI177Mui38aLkUfIhDVFe0jw3QDnYl6ieLIn0ZDag9gsWX+bD2egS1tqC88E+
N0mnHeLRrMbkIIAIffBTZt8PKhq7rYN1NTRNiF4+MHar4XwHrDf38+6Xn412ON+yfclNqrn2BUGH
Hofz19/z2c0NIV1hkdidw2e09E5s4l8Cc15rDUlh3bvPkhq84A3slRea7wyzEbuULA9EDFrnRVgu
h5Zo3XhTw+blNC01B6KqVC8gLpM+RWz392Tb1n3Ft0Kvn72AutCewmfkhEtedMNFVybQiG4v2DLe
Hgq2BB9Gmb9hoi3buMdmT8/+xzoZunwivPuBk1yMN2rdFP1Cer8LlMnpNGspfI1YKb0jARO0AykH
PXs2gXdtKHGPTXcNnTVL1ZLjwLVrGAOKVWiGJhBUxOzVmVQi3//EbeiFRDPj+kzeJnlrG87T5vQb
ZRESCWv83M/XSj1oRO0nb2zc0SAJjUkMdAB2cFKKeyk4C12iis3oeP8jTILapJMebmkN2dsfBF2J
g/PuwbKrJ/mWlOjt8C8TRL5NF+Lp9rPOJ0T518qciAqsXKyPfRgHGMPzxuYsehOGdORP88P9oh0g
Ft1ZSXwfxIgKhU1EXDRiN3LYjo5Nl8bSmKvA44NqiWtngvAKZ7PIzGAW6h6qzADZbg2Olworkd7z
Ax9A9VqdQSibWp+FtYs59WAUusXM7y6YyySPXIMkGVRQMliapObXUwEZx0V5tNjXuhgUyKziKKEv
NW/Zh+UN1Zjk9olStl770m4rVVrWFeuX5L+uxJY4KZmRQCsfAOdEgDEFjjHsaMg7U+uln/saoMzj
cg1//lircKBnqI2o8Cm0XYFe+IEebvF0oBH3gWuA1GOjncj57PJ68HGEc1ZYn4Ozth+G0xVxq9CM
1P6pnGk58yz/He06QCnkHEpH0cFByiqhX1BjYFPDbY61TuNS9s5JmNRKwuPdXblGUnb59+NRyui/
WC444Ih33Du0zodws+nGIO79c3l7Ki1vi/Lryrhqq/umql3MktBTbFeg5mkKLLH1V7ipbHksPNwj
TdrTMYGF74kroMifwpG/UtGNSZsyagLa60RJsw1sUxR1N8nBy6HO+hOHXYof/9yWsSGqWGhGgdt7
8nQzrb82e/YkRC+LYHO/GrP982eEZAYt+XODTphWVE0Z1nnXLYonpIr4TQE7bTb5Dbl7kJ9kSmsL
XZ/8BCF8NztcLsFemKNRMROHBqhZnhZBlhRu4knc99RNIAqLRJ64xtCuvTajKkeASh+12umqoEfu
RUL+poErqjpSecmAzYnlXVzgLRG3+gnURCV+eJBZ0B7z6vMk9fLRJvx9ki+5qgPIyn1OvqfSlIf0
HzcIhynBQS2mSaWcMkKwHkl04uekyBQcCt1aPOAXwWTtVBn7CRNC9lQz//xN6XV7taZsvPhGuEKS
0CM8HrvzeJWxo4YOouTb2flFqkRXR8j4koMgGvjyf56EKIqqqclpDooVH0ANAs1TamgzpmifSXvm
rj1IFxLEUUVtBPVxdKqE84rIib0H7QsNGx0fFPpsEMQNDpBi5Tt8dYxJ3q+RzycCv+x1Hij9Whxq
CpuSoyFdzbT6ldEoJ9IAgmsTvxpFaH3MbI+C0OAIiaMk6AM0D4KHdSDnvOjh52XMbn0DL54r/2TE
HLj4VsN+P9bTcx8gPBB0hTgyiO6rvlnIhHUu5urePttDZfk1FQWyxdJxqHdkujxlEE7PNFtFP8yw
gVIwv3L4ghJvAUL0r0gr6WXN/OJHP3AibpOSV/fAUHzjOz3G5mVjzBofk0r9yX4bQUMm1ELpMB8F
y2/a5+g4Q9YsIaYVa9Kmq7x/YZPL6V394ghiWYZwK7Mk76tuMQx8mLKd9m17t47XuhZzJ4pDB0pN
0CBR8v44wnSYvcb1w0rrsGTTPEZPaPlXFiO22FLsIVktE4ppDi78tsbh4f2m3H6IGFjsDDKSkJoD
dFuD6reKlFXnTZjcAm8fj9/bySvTAcrFQlsm4ydjzIlLpgKw9bJTPe6LBdLyP/4wawk+KB6ptZz5
62TE3f3QqkzMUM4/7asGyoOrBZrOUhCiGfFaQUjrhcECGbJyz2PKAogjnuVsSbQzjnL1OMYy9p/u
8wfAMTdgJVKkmVIAtojN+pDeEuGOeuWzvJaGDLfc8CG5KDyAxTYHwdQ990S3X2F9OuPGzjpYL8AV
rHow0IdqGgwC3lH/xiO0e/oz9HHobDcTDAnLPBVBjVcNKkvk0Qs2Mn7D83/VV4q+n61LZREwvGPF
K4QP0SQDu/3fxOTH/jEml64Fb8kRXiwu4etPuMu1OYsSVNaaJnWrOuwYz8W8CRjTYyG1XGxJQumi
zW1f248bqyeXinGcvTTE68DAIEQJlPhW425kAOIhRCH++kdSW1oNHNLxqWN3NWlmegApKEfC/aHQ
8o/TiKfSlPp6IHDGDjmKpz/mc4hUiES4xfY24oAoeuORiiS4ky7Rt4KyoFZjvRrjoxbfSFNQkFGi
/hXsxorGbrdrjeUFhMaFELkxvUybYhWdJmo3HYuEAi3ORjyin6neJf3ErqyxYI0H1aqhAfgSseuK
B11oCClVi4PNcJxwN0097lObKRS213h+sTDaT9z01sKJdRUOAx/b4NUxDnb1ekoJgHYuoJY2RxOl
DqjTGWAUesudnw/ZAQO6edZp2TgAFLd0QPNvkgiOAT/dIl9y5/wGbmS0LLLXem8y2CiEyruNvcQC
0ucxPgnyND5aCy+mnUHvgskswna1QDLpQvPKToCKAQUtSrOarYYZhF9tqIilIKquxehAejSrnvH8
f64xrwaA99bLH/B5qT19NbHcuGNlgP2Dd1RlK3oL7OMXN0w6RFJl+9k8lPSPL6MM6zfQo7LuG7vt
R9MtgqulGEKD4/s4VH/CNEKy6ONRA773tQM7zILjb4p3oKMbcVrum+wn6X85nXJYmvTTEmx1AyeZ
r+u91Pl2wIz5wOz8WRtIkNLYxwPFtbQJS7l446TJB/PLKbxssjjB6p2k9owLrfbvdHZOZqINQDID
pSn0cbZp32ESI6zFvFyXN4CXMTrZAvZH/jB7HgWA0RtwxeSPVaEncRtVTHyNKz44NizsNLViwSWf
g+xBFP9hwXSgbHgOzs9+OiDThGQkZcUYzmCOiKce1xwq8OihmbK8gmhpyH2UvjVi5xKtyYo07nCY
XBbWiwGpUzgcdKK4P5KEirz4NZ7KnigPSOMvUt77PvGcF5diIThGXtTcvi7CG7mvB62uCr/NeucW
oW13Fg2jr25dFjXuFoRUDELmrD6G239cpbmL9UjsXclNwGM+QOxEvDvIOXmX9vMdJVGyN2qk8iGT
XHbQbLL00SInBOnosDQUVi+MP/aLxpFjAhMcmLTg+ySfgG1L1eC1El6j2Hwgqago0uMWPzaF2vDq
6HlrANO9QZ80jWktB+Uz4Ou6IWSvrwLP4kmBIJq2tiAqV+XZj10y8EjNnTvs+vopmPiQ3NQA5bTR
9vspo6RQdwmVWjfbTNSV9uPEy8ZcvmnFzj1FfieA0qrj+jbPz/Pj3Ic6Wow3oHI/IrjfPvBmdCfG
6ZyHg9xm9QQjImdshH2ORkgCmZT0jCTLnSTLCJcyuplmy8w9lD6RCTZ+Yv1BdwCbZVDuK6aOhQSA
hUlNalvCZTjfe33NhYwvxortWS5aQ96Dia26th7VPXX3Za+x/LB6D/2scfHcf26N9UcqKxCJa0FN
mePXDAMyzzfuMHiJ8pORpP/QDjXFQiP5PHmaycKU9UM2nAdEVQAB9BClTlEDUrK9ynhydzMpaQb3
RyVTgnQoG7XpkpGTMdpPCmtdhEZXci6+2ehhkk0KI8FLOi22gKlZBaOD+cAhyLM9PovGW6MlbTZ3
3Dy0IRifwg2OfujixZliKgQ+M7VjteJC0CWCGaXSysbG4vclt71ytbUMGZy7qgLk5BJr4qOBUlbQ
2bfzb0OsRVmjC79MNogl8ir7WSvfB8sB4w6K0k83bJR/uiEVeyUTkT+IUS7lzpik+Q4s8X52tOQw
r3HS/kcKsDO5Xat4VgdOTSJEujQdLBArKMzGINWFdfzFKSNPqFBetRIuyDYnManrp1QW2UVi7SZd
oI3Tnp1lxA0bS5ycAXVoqCc5EHm/EWFRbnUa8NtNQjs2vNz86D4Xdsjbro/3nKuUFPEQjTELC28V
r5BLf+rc1Z4RvwsPLs1cDTwlQ5Fs/mHeviqjQXMiDmDb4sQjjEjnmDGVUFZYk9Tz2moSoDGv3PRH
TvFuzkTdShxOivJSrTT3gD/pef04nKa/2P/8qwt5zKUNBL7PXFxXtEJ67V3O/r+L4XRNJnmG4r+U
4OvV0AH33rXB8+fE7si1PAxjHUfeqK54tsydbuILClY+I2ioUVI0+c0FhO7qUi5un9PrmAcno9KA
/UyKSDq5Ikyxszkw8t/PuOgBdT1yeZaofMoDXL50oOk0oQRqR8EWvgBBAGr/zELZpVD1PmI7fc3+
G4Pr/suCwyGdduyb/N377TdRlN8Fj/qIrXVnyKB/K2FhKr/cdhr1PWQ7poUqYnzqX/TRMSmQSGwB
yLbPApjdyJuWcPTzDHqmBMGTnPKg01wiEZnISOS5mdkXG0qYS6jv0sVgGOnw5ZXTFpcP8hoUmvhu
mytqPiKx30V1a5UVuuiFtCcuM5noLFZwin5tOLbxFrC7gyBx2H3jvX4d51vmv2YwUG2MICQA7Xsy
Ii5UEh+Q8d14XG0nDVvtBf557AmO88ljgKdBrYEVdBaGXT02MFdbX0F5TaBPGF66ehnqbhmv+iZG
FMyIZ1pnZeB944CZHbEH6aPXYzs1XL65vvcA2mhEr4iqA7AlTTUyZI92PZoEd2nCQzm9rz4gdaWG
+3cAcMI5eGoYbLmw1bp5mbCnHy+LQBBjwFd7Fug9o3t7v7RWoks2oJvdndyunMVRuwY9RqCNmkh4
qPgVKZC7jY5h5z2B2037ktOljU7OogfpDX6VwnhhYX9a6RKAtlC1jgIMO/QSNc54LyQJRUV7qBTZ
Mgj0y0ppF/YaqKVEXoqZzsbvC97ndA/HGKcF/NZNP1rQcKcnk5ZhDRvM5r2jqOIyk4zUOJVhhgAq
4NfewIiXJtQkhRwZ+oFd7xL1EeZAne1IprB/0V1W2fSHg3ZnDvV62y+bsByRRiH6NWMOyJMqcVow
lVSgNtoOzrSD5w1Do6kDrZMZmR2D2kV8q3TtiDLihq7RBEvLZrrWFriR3XUADMqRa4TnyWVYrWf3
cYkaWzvm7VyToVqetYOGkF732e861xW6fP/sqB8jYbKl3QsLQwSyNa75k0OHntN78+kiqDcZA5Ix
bKFZ3+jbAEUrEZMSbGpG0frmhQBDA8dgF/MJCQYgfFbXOVKUicKvkvL4eDQ96tI3Nt/Ngf0bEUl9
WXA6Y/wUDZO8lg9cfJQpnGY67F//kf3CzR9f0W4L3RHG2NtPSPJTC7xQ6XzS5TnZJiLt9fubKcqG
nMghJi1LvjlkKsei9IfIh9h9kF7aruvxkacyaWpE2014faKb90z+BjQWrL+VfbB4M89oLoyTD3s/
Xdw6f0yt656waTRBu/DpJPwM8mVuKHJIAePc9NtMskAcFLfVqTARspYBJqpyj++dT+l4AO0d4C2n
jBhfL7Nm6wAlINxPsF3oA25FeIutdzDGMITu56l8Ib/nPUkTyTlyOEG2yiBw4VG1vh45HZsYDoA+
ee2kznyBiQcknlcNzKgnuOJwS9eOXD86Wa2UCGGvfAyt62UpuOkBWiAHyGra+vAVsMzLcDpVQxO+
2432DQEGSucxohkOFHw4CZCdhz8IuBKXasmduRjqBK48Td28f5PnzVyDv8EKZLwqk+ID6+BPQXGl
E5lEEJ3Hs3EiBuPjJFCWxSGnpmekkWcGPBbYRAjFBMzB1PG3tZptcajuI8CXFK8ZkkfcZ7HIYiM9
dJSY+JuExf3hjvKudO6o4DIqdDSEzlKK3R91yr6aJaY0Yo8rnFMJdSDxCcCbzHJrNYEbqm+GTw9a
sg2ZQbU+BzPtTCF2taMKL8tOylH2SaWGv9s99l7yBkr/aYZ2aapeDaBkDgBlp8mCCYuJ16KcxiEQ
VOC4ZmX2PlAK8cwqX+hsiHvFdDdV1KI+87huTxgSxqK9JoPoLhktu//c2X4GLQARX4fsqPhfxnf+
9Sd8T1Lf5m0upoWJ32B48gs6rn+Zu1KabuylqqsH1ss5lxSag2CjGjNQOcCu2XlU0PltSMSZNvlN
F6qg2ftYTmuuo973FljSyn6Z49s9KL07BZrKznf+BB/KKnCNsCMRQFyLdoGDHAH4vXHfWWHw8FVp
ZopTgljekidyclY0ujl0NfWt6EQjN3uMG7SZAUocrI1+26P8JErA7DlG0d2uWhXBhAzpLPWLWjfw
A7RfG6wjb3ELvtXNnpYDtgxx4Wnf2BA/GTH+6304P1a4eCkpeglBhYQK8quZKMwkMgakfvfymdaK
KciyogibEF3mUefVcWL5RvCX8R5A4MHEodRvhdMuWxvuc07MV/R7ONO6EsNkYrodIlfNvI+EwkGw
L/op5xM5mI7FAhpe0GNHp8Grl6kdJjpLoEtryA4D4Q/ZHvf6p8c6BnOxoQQl2NeXraR7Yozvv06C
+1B1W5r8RZDowflIq5h4CZVCGS+qy5zPdSP4w0Tz4/hhCzadnsTx5wMXpeUXVphNoUtXK21x6Iez
InxDZG2O/LqE1ZbT/tE9TSXXTdiQtj2srcZYdsFOqxbQcY6KHCGaqY276y80gb1GKCOK22cV/bMy
MJbvjcWJWC+NI4Enngu3hZ9U7JPe9QnemqBLG8DCOt1vpBX5K6VcqTZu15Q+HKtPrZSqCqOuKedT
Nr2atnZlmRqOmQd2jY39LqR99vcCqWaMVk6khosgu+TeSE4VDZ/DZPpgAoC+KbTuhnFkIgTjtJtv
HLmBNYAh3PfVABb8/zPBgIsiLcKQXhNtvReghbOgigM0v35KG8/ohZE8xDg1MIDW9T5+AnzOmAk6
RR6fQqUzT158/3E2X4t5jfFThtF2gVOLk1SBoOQMfBnMvpkezz8ToM8beYhQ4nfM138DkpqzJsfb
TPiE2XUG1YeE4ad0+Do7Sba99E7Pbqk+qKpG6xMdRXt99rlwVk9qyJ7k2m4INll1gjCkas2/Ho31
Hcu1k04KeuFnNyxcOnSoFM0HoXuz4wF9wN5WgKPvu9wdFAXZJ1VECtLxm8O9rWTZDVz0FEZNJxZT
XyBf6USnuGL12uuQCFcDHkF3FegosGAffFyxYRR3LvxaWI7MIizW4MnXr+nLZ0hJactCsf206CA6
L36QW5As8kyIQifWObI6W78D1GA3Dag1bJG3zKG394p39lpqeDnzuW6NG+5J/eOoVjuC0h8RZ2m3
E6CVCfql8NGFJhh15cvIban6uEsiQaGv6UWUk2Xz68oRAsUl40ERRYz2EqMoQUTLglsp4gyC6YDO
TfGHbN7psIz7XAe/lkksX75LC8ZdczVNasShlQXq1c0PsxhjEgLiHASMG9ibREW1Neglg6/bpK7h
hycd7D7C2VT4anprkNvhqFdTLoelqxJ0DCo2aVeZEZa75orMsD8GGU25qgENgA6PMHYgU6pmDjZ4
3lFP7Nyi3Ib7/VOginfMTvTSeuuMQasvHcVY2vs9GoFYj3dL5PBhOOzhcarY0dxh764ebDXjsWTu
9yRdOWAWbCfdI886gdjJJvTSwtdRYZ4N8aZXGeMMXBnvlKqG98dRoh5evim3mVkkRkNh3oo6ANAf
bYeZ5NDpZSlNqeqOglHVLUR31U+Gm46E0DVZBuJheph+5pi6M4S0y5E28gTpwSED6YaYRnnSCvnd
sVgHAkit5eR/j4/AHZf4EgeaUkWLPCL5bjMNpW1Zs32oSXXs21mh8B2Om9NuZUl19hPzzQgrv7FM
9/xPgKsmHONLWUmxVHMzSxdlhjyEEto04d2quBIC1atH3SCXegaXN5Wy6nwNLkCVcMaDIT02FM0/
SSNPD59CG3Xxp+M8g7ZJZqNr/6TTVrXpKhkPemUwSC5sJ9v+RTo2cuZpFb4GrVHGM8G1iNNaBLtV
W+R824qDxb0M+j/rxTFYHug5pD571yWWD6pImAKYeA/lZn0Ee3UTsBtnaAUw7sXiOV3U1M9YffVk
izBrzKnekLLE6/NspFEAwfBLmtKbIOq3PJWHXtKEj3aBCpZw5PEcBhmygeG7lvjHh6FzP/mhF7TE
6rMXq4FxB3ZxTjt7GALvUZYg4jDp/IbytN6RZq+CaIgYf7FJIiFSyteTQ3Gjmgicb9n/Wgfl879d
0umEdyu1cMOdh2HIzoMbLov09eLTlsybF420mFqxxUi73xLUYOuC3pDRHLawsuaW2L0+5svQ7h2p
/GlnaFepuDxjtNDEfCgdqk3N1CKWxChfFqZ9zzlAyq/oGlw2EFBXORllNjMFZHj0IrSHEGXf5X9f
FH/E8xmJIDTD3mdfBpZ2T4GxSzzT5CXU8eEoSZUE7FIBCXeAWdal/rntwRoV/7O27dpGI7lO/fIS
fzREn9urSZEiyd2TySxH4T9wAu1rvI0GD3jPxTjAfxY+QHYML3i9pPMgfo1rZ2ogKZu0TXxZylR1
OrqBoHAcS/Pa0KLaGj/8f2Rnc9WGMFgOBBtoDPUXogCPVrEFH4rbtV8rSi0ESD7qQS4d9QLvlUIL
r6rUE5CZFHMmehUzQvbv20ZZV60eOHHYr87np3L2i3p/G6vismIX4YmXz9uKrE1NUVzQBlx3JQG0
deTnjpuw1dApSEZEu0olJFwVQYJsGNuyO8ukRCc4lw4m6kaRJqTqS4qGWJE4yKmu3wGkOTGw9ANR
W2/Dgc1S6+YQe0dvY6LZFGlywy2Y/BVvTARqUnl0a3a0DbG0DnpCMrsnkqZcudyd2F24OTqEk90q
QQuGf+DKyvKh2JPTU5hXUjnzffzR7W89Z/A/NPKJY/jL3KBGDQbGVkEl87G53ysdx0ruw45wLlP5
XfXFVOqAG2Ij2lvhrpdbr7kkRaMakfIzB9LqDmEt4Tr1iZ7lFtGkj9xw1JCYB7MHFd6ZJdUqnOpQ
ZJW4eEFpd5ksT1pi1gS7pPj2YgxKGuzGn9n4vTmvX1aoTd2ifh6dTK8UWUtK59p9NQQ/sER0k25B
Y/vCn3AKtOU7ALDsPajUCApvhnjovu3uEvrEMmixDBl8jfImdAKmn/QSxG+yYFn3hxf9b9uFVFPU
88mztF/zvKP/W99SaoOz7Hp2J8hzFykclyfpKRH8b+GcB294uPjcqcKLiBUNEQjz3n7euyRDK75+
yTrtMPw1aGT/N4TYSMZu5YZVYQmwWgewTvI6mM9EahgNMDncdcadCrYP9dmXRebmb0wYRfrbq9zi
xvjQkkUr281BPObRUXLa3kSxSTFZoE3BjawzArVDzFLqlupkYt7db/oTefH+Kek7WrSNxMUhvfKW
7byAEgLYRCinYirML5/IWjN0C2WD5ZZOY5Ug/e8cp1EdTxFmzeLFMBYHPedGti+wHXcgAjE4xGkT
4W1mo6QHYXi/tFPdQwQnc3aepVzvYnZH/SFTBblllZDSDLOuoMYrRx0FEnT52baV4oKAut0BuiJV
mzJ6no2Zbcob+h2Fqw5YMz5YLam+Z6mGSqdu32ALmM6stYriGMMI6kbpAUtflJntWat8fWVouh/N
Vnyw5BNhsVOl2rnKQ95I3saBWaQ9+j1zLrrv3TzLpkCih1yF18oMwtuAT6Cz75T5qJW0eOX8QJo8
CU0Q8PPpaUXV25WLGdXMcA2T8UPQW2pjfv87u7LbqHKODzhvxian66h4IJBchGCZ6kqA9HmaqV7l
PEmrEc1gHXokTB36rka93K5zKfrPL7mYCNZky50d6w5EX/SRwcqvps7HZa/TJTf94WQIILuL9xTZ
se87UXS2PYPQ/UfImVOq69PEMiHBTrJErylBE+prhIK9gyXXq0wpinymW20kZDecGI9ZwL5iR7hF
Ee3QpJMfXgAlCiG5yqJ8nSbwb0KhXYXQ0lo07O+9Blkdvk9jUiaOVcf+I6/FR6gfT7bqz2W54n0p
zBWHcn9D960LmytmqTbaCe64zsItEiaDQaYw5b/T9IkHYlBxVgpCIPhdUaU5SamU6cyqmhQ51MzM
reXkg/rmbRFgJkmUhPt0/4PGL2KbHCEeAHimyHkWcFv4svrF+RpGj+bci6MTyh88gto0ybJpkRYq
oH/sf0oBcZW8LnQiT+8/rVe5lmOVgEreDR+P997pdWXHcVkGa97X+7qTYH978CGyH57rz2Kd/ctL
ANBH7LReanX8JigoI+MtbgpfEV6E3KqqkBiRcCtpEJruG/jaqDu2YZ9+vk+8J4Gr7HidOfabb14X
teObcj+usKAIc0eO9j8CzfSmrwQ4aRUX2bOzUQYc4rVdPmCuKmb2UIY0UcFNY2zFt2ELM+Js9EZ5
wYK9E1Ce1gZv7vGpS9bJq6GIXC7Gn5NDyJV9ooU6m/KGmqkbVG1vFFQw3NR3iO57DCqtg3W2ahCK
znQSMAgUU5sPej9i5bVAbW2G8uJhWZdsq+XGcQ2NvCb70PeYo8VZZb2dvjC2l41nlCjYvK0CHgQE
C3i4gYli0idrtyuPzE3UZbHriC7FXRMDWWv3opig8O/ANQwqMCrkqBDD7XdL2T9tep9tFeRbDg5P
AU21nzZTepyq+4gq1ER6ycUxJfklMDI0kl1z92OcszzSmvcUirJbWM5jbNtXDWvudrX0rotV6PrG
zeVWCYu0IGRr3+y3GVktToIz7I6a63Z6uJHxysmbUUGJgJGs5J8tfBY71Zbp+zCNbLjoS+rRKAi/
IpREojP6rgpd/ICOPu1v9gOXx4T/d/Sx/Ge4hYnX5dBN43D1VeiA0HFZwIifiwECArqwvCGlk/Oh
ufSr+4fQ7UCnqIy8m8k9ULr7YK2ypeOeopt8vmrqO4AujFIgOFzbSkGoR8ncUdVgTdmlnGT454F1
JD26Ge+vo7KSBOeTpTgmrCr+if6IwPCLi8lfLi5aXj6dknDqY++pyVkx7pbov9RRvXoG7uVC3i3R
YHeajLgDUJIKbSHCqb3zr98EFoQNlUDqz9tNWCsld6IGdlD2On8oLYQbk1PDJ/dZeigmWvpXkzm4
mca1Ggb283Xzxf2K++lgmvcxVJrCIBQq/IM8Yh8ttxUchabIsKGYXyYGEavE9y1sVgxeJczrRvb2
a4m9o2iNkd6GjZKT+fTAZYnN144bTkueqcZcFpz6B2ECqcGAs4ShhLeT8nYIXxKLwJ5mBUBcfwbt
r80tCfo9/6JR/khwqbO7MwGG3VKvLmCRVULTMvj1YlCoAGEYd/PJin/OWweRr8kid2/qwJdYTZBD
5iGxnVfjz4F1fKKU0iHS8tgvinW0e7yH+L72zxeRAenoMIUG7E3+Ry1xtIpx6e+6DEuXnfFLTA3O
xrKAn1u6Fx9eHfFcOaVHKwgiX1ki6S9wKvn5zib1UFbwrO8KWVkYV76eWjvLNMhkxJylMcYWXdUM
ZCHXkA5/uoCBrUGbkkE3yeCdpEs5TsaHZjCZt6+ceYn0mstU1pkm/SFrXmlbRS9p/G5LeqM5ANry
dA5/e6TDLYWSOoygNffukC6k0ajzMfPUFlkslBcPZ5DGZsqwTHwgNs4a/9lSJJLWnoeLr9hTsG9b
Zirs2z5J5IANKQCVOxmKHiMTO3f/ZFgJQh/MXTWclI9fAV2rCrWPsC/GIV1fYC6EBQlBmBvTtFx9
Yhpt3U3V0DZYjdYdPr0ZkUFFbVg1N12ZtOX/30zMz30BugnCEYG08qSphJA/yMgp9GmCzh/2uOpe
vlocj3jAQvgX34eihbuvMXISdhw5kClGKsIe72CqSYg9J+0x6s5EiZ/j69tG9ceEDHturt2G3yUn
D3aBGLLz6Psm9yHumc/Y7vRh6rNFcvjh1DGwmEhdcbOC1WYC0IfLqZrXsXwhmUDMMqv50pHZ7OCZ
VmcMoPSNwyQXojUp9vpDJDK5eRhNCKC2BAONVo62VR4YiWmA2m6TdqgBhxPJLhh25ZnXjF8T2pX9
+ktKjWIggcRU7U/oxlrAcZrFaiES6OrjIsfhq+xubUykGbRfa2rJSyWOTPXmXTW0Bd0o8ephvulj
oyT/Acb/BGS9JeubQFVjQRcLXerR9AEG7MxkhBvXOeEwB/GbtOB77SBE6l8G7fk+gcYk4bms9r9K
RZQP5FBwGn2TZfnc+81DI8NHiTBM7n8ktk0XICnKmeAfnkUQJBUEdkDz3Y6DH0nxsME3CxiEJBVB
3+RXsDc10bhWs3kvFIXKsQbiSBWw8DcmaKv+0VvS5jzv4lL3XSFch/N+d7NadUS2+QM35T4xXMTD
L1TBjjKJtS4V56i9oEYinoFTkfh9GI1sxe/Bzg6unBn24Zb1Bm0AaXDtlqJqC9v7iXW7HWK/bPwI
IR21i7izy2s/hOiSETgjCV0zivQjK61+YncMpmWJqLENVimcIaouQkrbjmIA4nr9FeKhhRRdnMve
oJFOzU37QYHWvjw09keazd79c0AfQNxjUVd3velCihpJlVH2VF2IxgCGJGdo3U4vBBuLPPpX66jg
9DLBcshDh5KxnccWJP1NyoSAi1l7MlQnIeR81nGFO8v15ETeEIZWMAdGx6ZZJBA8YQWEZ2T+V3Ui
4VnpQqIZiL6x6RW/nNuq3gBD13xzL55dJIRlbw38tDDT2pCINe5zbHAygvj5aKNdZkfnmcVUnuuU
DCgeVJ/uQmgnd/wJWYB15fyjrWEearRg6z0SKf5kGVFEBRkjCDAGiZoB2TLZqEhuoLU1/fJkenc9
uPC/mJwG3qp/3IskL5ESWnBK0QyalIXsM7yfk4Fsp5qmJuDjerFhbEHn1+jZRmbePnuAOZRO4WHi
see2JjvhQ4cuhBzDJAT9LcrKMvZnjJB140Kxl8K8AZ2gBHZwdMtnAYPNp3IbkvlJsyVp0f7N6dou
qI5v0LZX0on3voHdxMqahU4DDGPcywUHkWrsMD6s2Hv3DR4TZBHS8jkO3fj+b+WkvXqFAhv0wlfT
+EfEBHCHknXFd4jlqbt1abGY9uDWmAphegPJamyvCpI0qITtnbPXIfQFQucf2fLdM3+D3jzFggaP
dYyKjZtxtJqy7WGaPHxAHsAdgpcP6uhmzly3OPzM+dtJDVxVMncZR8pM2u4RaJj06tbT4C6YtIwr
epbQ5u12EpIAA23snQDUR/b33RDMiZx8gU/bds8/F1OdbZxn8vGl5CishOgHI+nhORvT3TweAyJr
hUP+umSeob5J01lVUSIxObJtYgMr+w9cmV0yOSBHP3/44iBvA+oezqYdm7NmcwgYHt9O47BFhpBb
sz9aCcYg7xaqyT/z0ZAsu7rykw5Y1K6wAm0yDPKUlQrqVAEsURvnMzwU+5KW5rFuonUKyJdfRTSE
ZFUqtYKKygVKPJ74d5sDJGjSAiEjKmfoRZFp9HatZe1vEhRGopeAnp85Mwz+CHo6lrCxkT2ojihs
yji1/snOOaKr9GKD2FFPy17PfcKv0Ba7NApR6n7B7yTOt47AGd6mXGm3RF3IopuJl+2mPeMYuvQ7
6g1rSxvbnpH7iGZ2Asy+WETyMWCqOoux/rjnrhXXR65vN/bAg87yubaJrgf2phYgvOM1aefgZAUx
3XOJeD/DKekXBU5H7xNP28sak5B+D2rWEzO6rfdDJZSZk/IdtXDaFCdSFl1D0r3x9flo+LqJyQg/
MvUB2Wj1HEPHZSa44enafpKL4SEGxj7iGzLlr47vvlrsThSxGy3vxk3Hq3iU38zKjA0T+5s7yp78
pgM+k1/6jwNPMEBrg8JiKMYSe1OY4RSxDF9PPaJkn2z2b2UjJiDkue7bvxw3FPUoc1yat8V/PifV
BVH9jm/SZbKvlbwsUFArWlNwAHOZQ6jYTL3MqgbNZiHEmxAdTjJ3bDZ5X8JvYa37v6AWXAhiaIUB
keoSVhB1324OveM9zeISrqsDg8dz/E+w13J4o/LLRGwSKCYprdOBJMd67XLFOviJhaqJjAHHQial
CKa7LOIQxt/NBuClox6WSFALF+DpHpflL8a7DKNq7EFyrHbksBYlDqCZGQME8clYfktz0o49oLvx
0TOKa/mY8ReTE+IJe2i372WPmsC+CP/Xmuik7+A+oDVTgj2wRESVx0EXGSUHBiO1z8/39hhgzv0m
5+qvqHuGM0onw//8cWHcOD+vx28GftYsYPuFy9JVC/o6vha3cB9+k4sPnYNmUD1476dSfY1ItDjD
s73uG0YyPZ/lhnDmWIi/P0sY2+T7tDrwk8FlJ8ejVx/vaGAleGNAXbcbRTi6AxL2iyMHniKQNPcV
Ef+C200F7r4o8LNpBHYPrA6yjBzdEvTX/WD1UWc/mHvvZwJk0ErU0gXC9/AGERZ7h4sAou9tzgW0
cLWs4TdY9o6yXQb0bPe25JGIDdK24PD8lLj7iRrBhuHUL41WFKm0E3A21FZnleb2/avcG8T3E7ST
x6LtM7eHxgh6aeWEErS5n1lQqr9mDTFJOLTc9YytaDm9zFXB3aRhzw+EKSDiBUWcMn3iYULaUQq5
uDpA/wiWWatEqNPkuUxjugoU/a5Az887b8QYB9dy0tTX6+zDEekXwvvor9iA1wa8goeclvyJEmJe
KkngxZWXiUubnCSG2vkYkpHQ47w7EZX0edbOrGX/IYixB3ayvuBCK32Bw3t0K7Eon6NPkJweQMFH
E73H3mZpFTPH8P9MTHGgcFy0IKKQhgeUJkjrQnK7s+TM7Z+Hy/sVQEJAwMgKIrwKvy99/Frx/GjH
4NZcTHw/DlPLpDLbRL6PulMtrl1ssq5PZKQksG/bzdON/Aj5uVv1X5uddZwSFgYnUJraGiR9XY24
MQvFVEVH6rIvgwf2BwJbg3imMJCsVddz32dOdsGOYnPLnMZg8sSg4oEaUH9UYmBCMtGuf7d/VB/L
D1jOMZ6348zP/7EIG5tUEGLgmBHKWd2tuZzYJsHgYkEDOPteZllfmw1Fe6TZaveVWhAI44PRWhCd
H0rhY/seGlqA+dfVuhaIanXbiiEfW9ZJutTH6TaEqr7CvvG1tywLZQHMjmGBOmFGwl7xwDWYifZ2
RzVjO+e55R6li8XLAGqJ6o2DLO+A7zBpKQsnTUttUrh8bmc1NRxTGXfws7v+nD8XPZR68X7ne901
CPTlxb5AnvnxYwQd0AjV9z9zxV0xc6wQu9meEY3Mf9KtGHbxdX99oo5MNA9R5VmGvSszaX61dk6g
/a1ocwBDgnr3JpfEMj7XSsTmvLf/so5irTXwH0MdiSjB415OeO8NI6NKXk/bFPYof4ZD4k3GuGMx
Zrdw/+0htOMNAUwg2UlcH7YAdq42k97plenOQVE8NT330/rUBFL+jBI+PIhPP+8YIVwG6fyWRz5X
9DkGyinch/UrF/R/WpJ3jeELnVBuz5aAl0riJuqVQ2iYdVgB+nYXLU7+c7n6hTxOojcm4iGtvwPc
3skX8f4UrE/YzYETflwxQtz2mEvpnld+e2BP4cDWQcmAvGEpwrnXA/4vvojRvQDkrW2ReX68i2XV
oNIBtAqbVzJGf6fbqPLyqayx/HIqg8Ri+oL8SnNQHpdQnPfMwapStCAnRNpg52RUqDJzl3K+dwI3
2G2/GhVIevcYQTvjXgUkrUSe/OdAQNsnpkhcmQTtf/DNttZfqRI303bmX45S22nidcmQTL1BdMfP
0l+3UU7qjx1yRzk8DhxuJjnCoPivkjaxhpNVfGAk+w7fgDroI48WGYZN/VeQ9dSH7U9otCS1Z7cf
3HGftuwR8VHVx1aKuhinNhG7LFZKSWTGE21fmgK+va7xJWGCmdTPcARnuNveG7I5Mkfnhx00lu4t
U21a2eDPUhIqRI119JL3HqL54/Zgd8tmo8MBO5FMtUogsaGZwe/k6i23g1S0MApkPC6YbSr+dCEv
upSYNFGaXZ3ePZQFoI9IhW5xGPrMFFgkP5swa2YpVmcCyYoWHgL2p2g/hPufm8hQVmEbM2LFI8qI
f/jceNYil2dGNa5kwhLqSLmhYhowihP6ORwoH3YOv5axyzVffgYRCDoyfh19gCUFUCzqVq0seoMx
jaKZB8dNkRIFMWGVioiteXkIeQmGY58p6p36UpUlCM1n3CsR+t3fy40HlGwbFkf1P1LWXYA9uh+Q
v/l8NQ15EIPkxTBejVkXrm2odiv2jF98L/o/xxTgJh7RVUbmGUaUrwgp15nzvZHNQY4NRy6fhOmq
ewGfYfX+F3POE1B72pfAu/gQM7hUi1SSPwCa4HlLu+ulzfolIQgW7PSswamCwo6OqcRiunzTI5kw
EK/JKLKsbVHD6G1h18EalZWnU+p9TdCOcPqAS9b5kH6UrjxrsxygiIfojj0vjTnCZb4ILHLlYHUw
lNk7YLQ/sAnYswq6i0kx5wkiVZhGXZE7lTbe3k7V9syDTKZLSDpxDK8QyAKwBF+cPl4WlhvfIXha
9V7aBAeXvFxv4VpahWY+acsDSyPo6LRp5n8H3AwGr2JzCw3m92s9fp5iGyguCZ9MHVsnyZsV82PF
GpyMiSfBMHcSYgUNgHpKblt20RGPQEyfzhHV/JV9aPCw5Ve8uKHoqAp7+Tp12+Jevr3FYoLWLph7
ydjZbeLloqd+WyHCgXAW+zSZ4X1J9GrVKvs1u+nUktAtzGvPYmHDnccY1iuawt0wIXPRzn+r58n/
PjmKkYfAKZEzA1VYGta1gkvlMZCHdGpYjQ424AupB9JY26BTUZuBGfJ6dHtnF7LFzqVFW8tu0Boi
cqUR5454rSYOygJDa8FsPwIDO5jPlgeqrme8v0GNVmd/0ESxeWsF+ML+nGLsNjgiB+6I3ZujPjXe
Nfq1904taGjyXnaP4kadwdTMtdiL/8loYIIDksrSlR5Ehvgr9JSCj2p40Uz+Q1JYG7FUBZ/splDk
mSH5VdEzTrXGdKQJgyr+pud3jHR9wDah7+bOsHa6UodOVylsLwF0IRd7piGexlkUVpzE788cYth4
X5Hlrj/GAsbmzTMQJoVbeRioUuM8QzPU1oGwU5YGM29Uv//9HPGmNLoFEnbfk8G8r9AhDc6EEvCS
iB282E/6LO2DA+5r0+gXcyAtIoQt94u+/FSTUjs/HrVRyF6Yi3kK+Si/BFG267WTq92IgJ7KuKcM
rnjsm+ix03BqI1cWGxSYEokXZVy3HnbKgTaiXcHUK1sTLAOS2gxzEFtEOmtVqQ/Z3YChxr1RiEc1
EGE7Roe5nnMMbFDt5cXpV4qucCJmxaQsmnx1l+6++IRtTIeaErKgbwB3w07PwMfRpRBKcpUyI00J
CNd+OXPdpqjS1cPQMSielft1EpHvTrsrPYASp0Vxb+dnDS+zZHXAnj3ycsTM+3aIJX6zD5wHN/9y
CWWOsNeV1NFxGD6TyrS9L6auprRwiozF3lJvJ2SRQ8eMqFT9EMdonzrvyPRLBm0rT8I8Eu2F+FdH
NuF+u1kQgll1/pEND3aQYNiZYZQeJ9WRxW6G2ICwqcJGUvC4vsMicKjNOXx1yV9236kAofTRp7aB
nSLwEImNCzrlZNt1TUKXiZhZu0rfkQZtLCQ285OTPoj4j788T2pW45q1tHZ/qhBz+j5qhAlb1Rc+
E3rv4nk4z/xpWTnqDjTTXz9tx0emhh5eSIoZ3rRADRKTxBfsd6WZxwExOqjq8yyvb1yMcqHvrGm5
vLPdbR0ysbI+ay7kLecX4og3rHjnJK8wvKBZFhpPA3WYB12Rmt3YnFiNv3Linw5NxPY/+GVIjflM
RkTnJaGW4L0QUjSAea+hqkww2WLk7PAKFJ3e7fen9JNlNHs7Etkkf+ogukoetEHYB3BYG8DKOe+n
9WndWoAOGhCymtJ3rKYKKGYni6d73qXfEUk82l49lBVoq19tumXOBTxZoxR8Cjb1GtB+QBWXvb+8
r1RaFVbd9eBl3NJUIOtwyAk//ajqX77RSAv/8gUoWG4BRTxXzdKVZjSM4xI7M9jK6Qsquiipr/ek
iqZ/fgVvK5fgbmWIlvzxsHG/2/vIST0dGkrGpDLtM+0azjXHD3r1LPItqmkX481wfd5IxKOstsqn
JBs3pek9fUfcMuXI5bEKYBVG11vRWq5sR+OOykGBiCZBRaHRYdp536fzbbvxKEpaTkc2o9TUDfQW
g2uiEBwLV7coZlM43j3n306tZUwe8k/7Lm9vwJP3I0UFuizveqbl3mkT/0CRJA5YDFCCJQVkHZvn
Ib7ZbjdkefH3M8o4n5fPsM3w5U/WFVCafaNYL862gccsCUFSLdLidzZvVNOdpZFV6f1RG2vlZ19z
Az+WI/70Zfqx8JZ18aU7Kw1D6YpxuIb3V84W+CTCjliMK9PVvrlkoA++y8MiYs+qWHMQjiKrFXvR
O61c44Y+Je/0OaauzaLcloM9j+LS8VYUsCntF99k+s7xwnVibnrJM33gBOGt/87Y19Drg14+/c0V
fH3fctp4qb6e1S2WKqQocaAs3AbtbCzoCq8N4GD7CAjRg2KW4vHYWwrExn+7D/9xKOuf+qBfrVFU
reNROzvADRCR+Iq9jnF31ZDTeue3rDqbIiKB2lVM7bJzQXocUt1Jo0PkiiGR+na0hRkhvFPHhtD4
YTD8PvWK+xb16469EoA1YIUkEWc3iy/ZGAL2opim81fqCaL0nkjr7t3elhIP6WbVenS2WTfYKxtG
kmW9dA+w0FxC5pfPAL09JzlSWlH74vkeKz0U9AEfAvsQUss4ivTrEnlFBX9iIDshG/hTEc0phf2x
4xpu9z/BgixMHtLTp7soSkejsYnaE2/8+CjVYsXSsf5A9pZyqScblwrMkD0gRRIvHMW0udjBpMFK
Ac+qQGaepUI+uFqq/aZjRCZtsZaC4ADJvrocK3bMYBmv5qcV9eNKuIi0rzQGPmbziLWDu0sojuxG
IOfEocgRuQAJ4R+gsn9iBmdu/2yaQGIwNEho1rVDFExcPS9qT3DD9rwUZPxGDX2DaCNi1uTHfis5
Td4ZrnBJPqNz4oXqH/foQeX50B5owwoT91LdgvXntqOyPKw6Z0HcEvLfsFEidNtfCj025Mw9jDkl
J7wfmNVTRYX1AgZGFMYJ3IBu9MU9sEa8Z4D91xsKhha5PSOJdcXY0GzMdY9s9pDtWAjDj509Jtqy
SxPTh65riHWTXlsqvJYYRhv1lb90I6E/Ef+zpkhxtNUCM2UdnXyIITeNG8rDIHPbZLDoouejc7D2
XXlr1dakZffx2Cm/1p1q8q4yt+B428vUI1gAfIOn7OqWKGFbtoocZHPncULX8LlqBaO23hQVNXIq
FBqv+Bc19DVYGzNkPGMOuqgIfb0uNzArqKbh7kQSc+GqLSuMnHlerDgECQz6jZruE3nDtFL2mmm1
4yU5/9Uc4L76i+xAMYDNjiJChIg8pbXHEoZJCYxGsYTqvFXJze9PNo5tIZtUKKIH/2k8dHen1e47
hci9EFoRe/IcJHvbg/wCiRjQR+eRtbVT2471VMisrnzUWbH7kKwYM953NQHFO78harW5ix8au4o3
y1m7EnO08sFGzJqGKFbO+2SbLBhr4HAW5/DJInipdo2KTB5rRmhbCUitMsyTTeMbu82Id+IaIg57
l9DQbT7jvLEmYp/eIqmVVlSiGifEYg1pIGAL1m+5AOBgq9xL3KpMK68Flk94EXtRNkRf2Zih9xyF
XgAg5hz+PcUpDBJVk5VfXFShrmEU3uVjAF5wpAca/yGc99oaa7csgnOfSZFzjgwX1KcWelngpxS0
2ykmeRo1udM0X5jnyHKNpGq2Y8se84xgYG5rXQZZXBX4REp7WV3dXSisz64TKtsg7gSwOY81FiAQ
ro1lA9SEvw2VUXPtO0Ck9H952bshhZwNz/c0tNO2zR2KEa/Zzgezu0ktRFOKwTYrXA84J7amyAKd
BYQ7ARSzxX+ibeaYFYhctZbE/Krpg/eTKqqM4IIE2Y+eP70C+hLXYqcZSKsJd1bQYOSEbT5mOpQk
pR3qaqPUr7Oc4pSGZEUJ8yZH3krb0iT8nMpMdumxV9/DWcue1H9LJrZHZ8lXQ6HVHjqeE1Iho2zR
ZB1Yolfsbkzr68uBAmiTlhGwsKoQLN7qTqf0wyYYsBSTV/GMEwGGwTwS0hyk+/CGDLrLHhw+YPXA
DG6FiY+iqGWRc7oNehXiH58aWOK0xgsAP75kCXhhTahL4sMYhfBFqCJGo77xE71auJ1AN4Xxaf6K
EKsUUQnQs+01MY6Z6Kuig7YLiY7hTipWPYEFsxxd2igZVUbumNyb3SZ28ps9aRCsbm3044gk6Y7u
Y3EfQubJnO0lRroEezqOxsC9O3fQJLpyZoxlcJBVDEl3bW6ZNDKG0MTev03WRnCujFUiPLe9r5+8
6B919VKKBrAY4SZw8YwSVLEiAWFGCZ0AiTHuNbxaow0uSLfmraaigw4ff1RtiT3AgYSL2bYPasfV
uJ6D/TMkZyd9B33Dcx3sAc1+MKHjjwzfhnIIEhkYJw4gcJZoWVO/K5XnMnDgw/TYa6rbHtRN1U0O
yFv0onrn3qar+Q3h1eOMmM0TOw5UbrxpFQBi/tkss/koHEKWvvv6M25HS0KAUN9zi3hFgxXt4Jy4
aK0n1XanGxTm+jnb7eQBo7X6B2Ycn7zGAfOb+Mly2gMknBzbP4l9g9qn4vaBrQNzkvqAqkpURGmW
urW4uujWZ0An6fHdE5pviaGeWS5mPLo9dd2FcoBqquhxhsX5EtUGF6j+u8yHSQMNJ0Mx88OO8fzO
loUSwgT4mo46BFxbVA6IFeQsKHUXtQVN2Tsp1MhbCcIcRpRGIQBg7BBIckRkNyrGO16XdEp5a2tn
dafT4HQy/Q1EOvNdTVUtmFP9MHyjdezz45v+zuetkINoiDnhYYkryaVx4u/gP+EMkl6jpyjNo6oJ
fTa2OR7bPjBv6J5L6Br00eE3TcOl0pTecR8U+M6OY2DS0UuaMWme0U6J5U1y2oci2QW2hf2kRB/c
qyWiaYGfZui1XnWpHtbPQ1W6HC1jwMcU9KKJDw7CzQqjlVbSByBZHOTEDbtD1nEPuq3hdbSGmIME
CM0tm4a6EgabjRMnw2FwVHmUUDKrZyzjnt1HEjXwzbkjTcxMj14cXBXi0iZl064+S0h4qQav0Qj6
GBtfJ33wDBPUIniPhE1E3amvosyOj6tUuGGiNExPWna/Ase0UMSkc2BWpShEXHxmiCJY17iILXEX
FmtUHwJKN5LTcLSoy5yeOcFqJbO1yexpNhEGLQxk5cUIgQTxsZ+LPqsRE0SmCeXtpvpdU88ZVTz/
AaXsBtTA24PZoqN+H/RwThYsw0guFwaH2uNJCmagYdRPMA7jdK27sekVOwE4aX3CLhOT5elPrBf0
4P9q+ebYZSeZ70J+U+XHL4dv0yjaZS9OW54HwWuOxUjXCnxf6OA6QP11g0qfYMdGSb8NPgcN9MXM
liWTIdQjcjvAtnuQ/4HjNpMleOsBuL787TzlEvWU7H6dIX2PrdJpmUIUR0glAJvHa+qRuAXSKjZT
fOT4EdsYaW0UMEfX82/mSEcRqRkuz4Rq5qkMJvAz9DPMrzrnVe6voAAd7kXped+Zwh7cMZIMNN3f
FH850bghlAGH1FIyZvD2PHci049NPNdezASLKYQyDTJiW6vcRXfeR3J5L7kgSjtyDasYb0PqVCKP
v2LlWiKWcsFaIi97hu9yEBRWf3c6PDmwK8R0FW/U8OHxsaD6qJeRHqqRj8m4iGONJ0cH0b+tQfou
K3URiKczdwyz0x/6ojZMKQKFURdCot0lB7hfVCjwzXRioLrcXfeItdLnGdSb4lB3KmKA0hIpoi0L
o6PG4ch5FDwpcp7n4c6KkrVfdGxPKpGAgRCQfOg13F/8Hhk/8f8IA4hJTDcpI45M+/IaFrro+CFS
Wvq5mCwoBU1j8l3oHUIqK2WzGFZp4ej3DtH3WtHaX0Yaa89z1eDJJn1mJEOYxLAv9L4zJmpQmIx0
cSqy6ZqK/Np8JZHXoFNiGCybBy30hukevP2E+ITWBP7KiZeTrgCARorIRxAHsSZr5Ku5apJTOr9S
FWE8fht19K9absRUlCToDmmiNgN5ubESEqSZDctb0xKvucX8mQ9kljjS46TrZuIBpS73cmwcTc+2
tS+RAFz4grbsO+HkJiK6zA0o7vqiUQman2IEl1kL5PinEriipGXH2iBv5aasRZuHA1gf8pRjyAU0
lzQFzYmeBCCWhdvnx1cXCfSkc/kE0O2fSaquVBQYn/EFPCOHHYdS34eoXtCmzgIkykdlw5uNKCOC
e8P5G9au65gkytRvCpCai/JTF/KcrNJqUv/2fyue17Z/OLYQUfu+2lRLXzpWEqvTc2hooe6d0zgW
SWG16hjP5df4SmQ4EzkDN/9my8T0H6X4uPhEBi16m9axtsGo0EcKPLfnLKN++Il2W5N8kdArtY0e
VgCKDuh14EMOwqu5AR+33Sti38MY03qiHut5VanT1Ay7LDvgG7SZTw6pr7QoSfsLOFjHK6aSPVYA
DzZ6OqqnN/jETsALnPlwfrWZixmI45A0iUW6EHkMsL5zEXYbsxynuw78M3mKFkPbmZ//fcnT0lNu
pmypwxMlKgWK4oeuzLJYiKL+TJSHvpc4X3V71dcmCKedvsC+l2oPdVLQM5UAEG76JN3vlnKpjrgw
M2ehTv3RLPfyC7cpC/UY9ywdLSzAbShQRBlPgYPktggvVo5fgDMPcHJx7w/bGo83re7EUBNO7JbQ
H6VvGtYuiH0B1hBUc+fGssUpLmfii06CWnJDaJX80RosBp1eNNft5B8+wVwgbJvPnrjBfxWi9twd
cp6fOUKHKzWdvU/aqD40gzRLeuxy2gHXPYrpnTTq57vecDrtVcZlDpW2t5bvronsY1SrKtyi3tAI
+/ZmB4S3Im8cLfLVpM6/YqXfH4kpW08AI/QDLhD9INxO91lgQSGbueDnYgzuxXIaXNPr5kIWYLSi
Ks7/N4F1o8ApF5neX3c8paeQuKG2VcGzXgB3IwoKIXIlJLc+ZELLTCfjtY9ECsv50c67l61pHkaY
dX4lMxOMXBcyb5tO3qZxSMYFoWsjE49bf79ct/Zk1U4oD6T5UCiPsPf/3xMxz5wfyZYmhG9uSS7i
bIg23vpvwwn8KsqWs37QtJLzRzEf2nfwBJaGp6YORu6zIo53PWX9lk1YC7uTMnbN+twjWIqL9sTL
YyEa+DZdoyehof/ROLcI5cJ/VT3umeFddWJtC31AIMzRDOGpEGizKzEC0DBMDuiYZ3TtOrBcb67J
14Cbwat4sB/PJrAuBSQ/oJqV9S8MS+B5BHKIE32RolUshSiSiTZMdnMzBmKuaeWZTnPAmVkQIhp8
mYCIKhPvqAedBodryTHN/kbR45NKn+YTBhGjp1+xCfZKvG1RM7MZ5W7CD3gpE5gePLAqxg8VxPnA
vY+2mGlXmdiPyEjVr+RGv7/ewvgZfz/Inb2XXdGrKY6TWURde4ZcST4zaZ162IDL1mVXbu3PI7j8
HkA7dcwG5GAftMhWeUFTyBKubpZlw7gf3lQOfEb6Fw7VLcl19pO+WVOA/XvTYhPKzNqaiEN8sh6b
sOLzbL3BAJLT9RyTOIruEyAq3VNnUZ51ZmxmNMXVv7HI8eq92tmEdDzIu0tTEQ3Cqsy6xhycC8NP
ymgn3lz9J8gUxXVSfWrOXZ2obgIz3KRdtsfB/ExCDeasZ1ipNdfRmzlwI7i+0r7OJvID6wmKgDor
Z2v25m7m2pOgj1R3dXt2UlxRqq2hiPinKF4welwWlG/4yAux06t8uJgE3yDxQxaj6U7Eh7z3dmFW
cUGHxkUYrgHa2JW4PpAL4TMKVr58B+x1M05U1ygd+9/aYsGFqKLjcH/AgnPZsDZ6EgKpR2rYhZuV
pt8vnOsQrYy4IX2VawcT3i6tYqKtWsvdJtH6UlnCQ5IY/jivZraJZvBZsMg4r1LzLXmrTrQnkLhS
v+yg2yDH3/AcRIrHL0I339dpR5Y1k/oB3QsDkqlBmoqq1DH8shsB1wJkWHKke/TFLYiVEY0Lmv6p
4VDdglF4fZ+5irD8MeKbtQpPQV2AyhljArLngKAtboE6sKKW1E0b6G4iazaih/DvZfP1V9gfK5Si
d4wWwlWaQ2RFhBtf34Ot8df5bPb4y/4IxzZR+DluWkp/uxFDWXzAwr4tY3jjbAjqs2yzTga9qHmv
aatB0K1PVjAbqzZLRO6BG6wR00aSP9UYTWbK0HfOmheLoQIprAxxajGp7CGLDyju2n/u67Lk8ckD
rXyQRg1Dnz28UkCes5ZF0XyVTm6Asa8ViUkmhGP0nSGWbpzMMDu7Y9PHKgJpduu26vzhVTnCuYbW
6xV9aI5iSHBT84+BMdXqySGWQXk0QX4UeV2N7RgGRU6Qbrpe9miq2TYFYu9sWtvAK+uzE2Q3oZqm
e8+rkWbnaMFTUkAzo+cNBckuszl76eKwadxlFWpsGrzTm9CjK3QSUYwSvCaiwZZc7XB9T6FWJLjT
jXnwsF+3d6eXRoy16qyG5W+QbCl3fADG7Xb1FSepIJB8jcQ9bR1W23GL+kas0glwgtf1QBMmqyRc
MTBPG7TN/dcnL/ALgCfAlvj25o9unfLRMORmygI+hubFbTa+YOFYILzIC8iDlFr+/C/gTnoOSH4Q
tgshxPpf5MaIgSZ1PiXtBh3iXk4VU+OLnESei3uCRjVe0O9WSi2UocDM5T6/xAkYEFgPIiHZuRMs
bRoglipeci1XhjZ9cTYX//bdIPHaLk7d+MJSSXuWrzCWmEezyPbb1cQXKspkYWasW8gW/79GbgRj
M4PL7p6L+dSNCVx8Na+XHh8THEGjwdeWkCjTKDRD1mXo1dKn7P+eLuZkRqpuUGdZOH6EU7gQOxo9
tEU8gXvgmRdEzkK9YfkF+Zf85irs6bTW46pEnULIdz5YbliM+OzHR/K4nP4Jn8WIau8e05bBJrQm
IsNVO7m2o829XJosdKlPLm3cpxzDu0lB9JAjUjGSaoiDZay/4BD9rUQbLljMGYCPaji10juWAxlz
fi/9hdxfkQfWL6Wd7HYKGERuYfPhttpQvqAqNbxayZFv5z3NXHqcrpS/0b9D8Qil40MpIughJX3P
TZStEUfD1i+gFn3DcEwMRK2qrBFuwPfT+IYnCaxlPUWC4jW1uJuv8VZCa+r+ZuWOeGTdTmA0tcjd
3/lo453dK8GVwmY7j+5A55hBnUWnE+a7EDlgN61mdgE5Qy7Ws5rDWd9U7tjFsoQo1OIE090chg1+
3Gu1PwT/RdhMiBscLJadrzKOR1H0dHDkxkJSnfNsRRhJPqmvTQvXSQH7zc+ZA+0KNcouOaEf+dZ4
lrd1QIKSRwO/Q6PpsZG6YB0AHpdAN5smD/Zct+KykhYQK/fmCYuINqiUISSRJrrllS7PiLe4w1D2
WmydZWClF/lmKMW5kMdhGRE+zSTR6kmW7G6QOM7YTFvDCI6hqjKWii+oM1xxdLlzk7y5MManfp3A
/mepxZjsfBK3KO1hmaATFrg9ncfGTrp324WxyaF4MhnuaPZJUmAyr0MbvLfR//HF8Bl3kADdR2gj
UPSsmCuSHiOheuIVibiyfmgfnCkxf5rNiRNORzYQegxbOIttuzqiuGJsp7FLSikFdzQ/MerHM8Nm
Y0kzAvT9QHLgNh5Yyg9NIrSZe8AD3Nq2DReSQHytlQDKln+gnNlGSZfA+JvrEZRsms6lkK5P4Imn
ahsZDL36mkb4vy840Nmo7OgVyDLAA/L2zyIFHQRMrlzF88bkpBG6/7mwfMS7t5AfmGKvI22kHqxS
ciZ3BprHZrKozqSIda3k+x44CEYaQjsOnZqOchFxBAMzC11Kzf1n4zJHyCgPv7GqCWNNyUTvI3sL
qrnku9oVQR/X0x1NsjTbMB+jbyiiev7dDwqCqQ2G2cyzIvKERwG1q11V3JlVN53XdmL+yjZXNAL9
yAlNOiP4F5UP4fFrTaG2JBwpAb78pHwBja0O5xAZ/WhBtAzk5mmKWsCCkw63p6+vrZl83ZNTcBqG
nLP9qelLcfUh/lbYzMqY62w0oeNnvuM15zFHwrNJZecz4dUDhNEheg9b7i1bXVGhBjSeoxMpNxcq
wlPw55OLud8DdUvTEVKs8LGsSjOwiJgoY1Ru2Fu48hWSdet/4Vk8WoR6aMUyDeVj6DoxlylvyuyC
Dec9SaPhNVIblFX9qoD09bxDVks+QoRy6WSUN6ynZnmo31umKzJaIgJZhsGll1sH8/xnuDsW3ycS
kIya6h7QSsL6Kl/jS16pMD8JYXoWqTgM2i6j+a4xsP8oBCxGpTwKAqq8r/SN3xR2Edp+Wn2j0guy
1U1cqAC25K1RPXedqRiqj5n1E5N5ekgeQ1Fs5ykDkYm8BgenEvD8kr/oFeOin4fyNrzVI1R5TSkm
P8WNH8HEzntVpcz5PW2ALGRTwFOyzncz4pri55XV2zAxiySlxFhZW2bYZyy+Hhb2JVEnxYTEfzXW
KXlG3fXKJLabNdHr9Jcct4NaNJb2lMD/55hFW3p14s/3atA5ORFOVhtolCC0hjfzzCIXvrKiq14S
Ukv3xnDtizFe0ywztIBi0ZQuLhqTitoN6r372cU0blfig6Mexj3oeHQuD6ICuVnBA2KmKjJZehyn
FibYOBXD/Ny02ibHaPYpclzJluKIkkYR80TYDXN6GcgdBpH+zn6aJOKyVpMogrPGbTJgDy63uW0w
QePdCrqstGHmPPvZvdNoasLbgHrvZACfGvQsPH1o43fb0H4SqHUXoZCn4vEU1JM61Ab/56wfQC4a
6RZtPB1iEUBKAdNxbfAhm/mPbKvMjqD+Xctjf6dS51TEVmlDbcfUDZIQnX8cj/lFAL8ycMXqE3l1
DLhkHc9/7gx6wxyN/cSn7MxVrr/2iCaPLZHU0zuc5fHtsNY5UonnSTXOd4LSzDBkB9HxFYzRUoAg
wACdDsWRGZ7CvQC74zQ6jjZ+wvz3OvwuU+gSXH3sAZu7XYYPc770vYRFsVbkt6kIN8rS4MOHsMWf
8uNPZoXepv7oYsfEXxl6xSP16gx3TzJeKxLwdFg2aAThwhey4dqElCS775lc2ja+mX1LK4vLQj9v
vvqGONjWcQvWSzrONuhW0QDQmjEo6DqQLCWJv+DyM9zBq08tSo1/I6Ncg1k+tOBlM6GP/7l14IGr
E7HN3vJC6l6lr4rFJQYdYckfZQAx1pqrk3FdjKbzTGd6Cf/erh2DSoWlgZWx6wsG2O21Q9I2TDv7
dmNbOAWJIMYasgwvv87dsO2joDU9le65gxysKNEJOuu5lNKkcHUFpfgDBT8F6p6yQjFNk419zVg+
NMJaCpJg9I0QLfrOa4094JvQDNqMLnjUWZBPrcrbBArx/WUpQuw5BKY6KP5XKP7eifw+sZX1F+xy
ezaN86yX8kmSc1cdcHLcR7T7yY0byhyagLTt3s1+ABkYbXcghR5WNGuZKJ73SHPIUSy+4YUTZKfL
EPL0H4E/YyYqLfCxGy9gF0BRg++blXj6Xng1Q6waRHUxbUfNRv0+LUzA7TdV23k8UG/sHODT+NdH
NMj0jUq7ZwmoRJNFJf8e+DrM7cgod1NM5bcsElI0HoY+AEQRgXlNYrx5L/Zn9sg++iQBYqT2DQqo
UevlEmM94INvWGrRj7psQsSOtsj4Wx1ViMf9v4oko0WP36q/Rb5MgHX9NRlhIvN69GWXfQqeFAZK
0WDuP5U+ZLszeVsKDSAreonzBY6gnVhRn9OjxXRhwxBPJT0+Hzqr4AES63WPLrGheFdgO2a8LL+0
8EnpnoQGmGFt09YWeP28Hga5734xQu8NyXZeRcVXyqQP9mbCHab9JHpi/IBFFW2Bl5TsMJ2h8v8Z
RwkgB8q13goW1anQES+PXOxzf3Se+dkB0p4AntkCvrozye0gSPT+VtAtn3IaSv8VuE9sfhxxngVG
6113HoJhyj6Q4FLeL1jjsGepyHwekXKHQPEU1ZnPM6FvycvCzDhjv5r+MU91UPD7vY15fti1AlU0
JkXxepetIq4+b4HALlQZGypvfYvIjRimQ+ZRT9BllrgrjkuD30x162T7/0PoK247dOeHxVYFtstD
1btVGl9nNuCwmD8WhjTm1akrRoTjGg/B8gqUgVUsvtWcZjJmODs6O8xt0Ou3ej03LtzhfDWjhVth
ZtzxvbvVdGGTyec91tdHCE9NO56rLXCfjw0vnFbOTpEb9OREFpytG7PA0NrLIUnKp7BpYdKIlY7e
Snr9d9durY3FsbO5Em5uXeFvQv6K9iy29tkdDHQPZLWgAqkprCHXHha6M8nF/CpSCVFejgEAL7IC
O4/VB75VUKDGmLQYKs5n3qbiwhgEA/gUGLxdxZrV9+5RSt5jy++YLMspCjUZiqpxnrZ/k4fDG1P4
Ze2le+upQafZQRBeYDpiXV5QzS2kYPh+IF5EtjUTC2BJ0faOpnXIobVf9B1qs6khEfakHOCzZG9h
wg7SeJfm2evSMBqe9ILDGBsWRyDwnW1VHEHurMv6nSWpkNPHU3gSMO5aCd7yRxYyrZw+whmZnnVX
7dKqvxzYIhRZnOSX6DnFV+H4/OqgrDKGngFldC38CsLuWZmxvFyOscl+Ca1sNhYQ7pSYzyD20eVe
49UonRA8V+9rTxgHAHSBKXM1tXQ7QkfHA6Uljnd+1jsNWhVvfBwaiaJVF+zGDWRXckWhSed8S3fv
7K6xGX/NagL4j2hORBdmbRdu0JRHqMbYZKt2FucSqCYSwHlTS7tR1bnqMpT7ofyZWPiF6Qm24/oM
Rt9IRkbbS3B3jFoA06lQOjA5rR4Sc4hjWNLRYrOiAK0FTLtIqIXBCDL+5ZB0kylPBlKb5BOtmWGR
YRbNdScN2bsO+4c9WRfXpKMsJgPf4aEUmJiKrpgXC93xAHj0SM78OPQENm+huBlF24ut9MP+++7H
QwTCyRif9MNNpOVio0VIr8eF8iuDEWv7GBIouf3LmrcVMkCNaXc1/JslpZ/N3zJLi301HdUYKFg3
rTh1VtKPdjqrpd4pOo+AbOvQ4OgGuWhQKMDyeojZGPa228xccfGc46FxYWGaZveJxF7MCZcnzUPo
xvcAeeBTzX7PHaZHQI+MM/4nTRwsR/TpQBmXl5997I58Bf4D5E3AzPU5B4184NUrAIWlszocudnx
h6QCH9NU1JMr61L9ajetrH9h/ZUKbg5NwE3mfJVyZZuJCTD8fYKgg+t0DUxcWCszUs3zlXMjlIy/
0UDEJHXHOyf3q4ZXb70JR8hV2eZggFaRq+NL0byr6KwL+xG4cF/l+sYIEWRC1u6eYYC2NDdpcJP3
mILKS6rRqpHfvbQlkEKkIUil2RiBH05jKkbDpxZbH4tuVcPeY8eyUDlmJslx9981owSLgqoZTHv6
Z0p4Gllwu9MGGtBpM3k6Bk2lEwTbMLqftzpszeY8KGjQrRq/3bgClkYAl+tup3ojf/ObafHVu3+Y
1o4cw35KznP0AF3rPo96Q3OnSXljrHl10mOUTFVsVs7dNP2zRuRc6nb8u7LntG9+fra9NlJJMmUJ
R0ZGPD9mCY8iv8TUfOcqcdMnc7ipybxIls6JxvByqb8SO91YEP0H+PV1eomkYfwrjH43Ukg/NV9y
OaddXJfcLUsy8cKLJLsR/L2bz21hJquT3vpFV9J4D3vQY239FNJMx7w0dno3gsOh+xGPSh/lzkCn
4cGS0XZ0cLYO9YWqFB6JowVCshIGK+yPat9CdbZcavSsUV3x7VaPKjQewshu5poGZalg6k76Rt1c
JV4c6DnOa0ETBf3kmNJZw+D9TRRu+KaCAtWEON6G2sEOH4evgPbe44j0yLcGJ8QRmHH20wy+4FKl
iaosNif9Wptwpm4ugJiuoITOHyn8yWmXx1HDozMvhphFMUlvGbBkR4J4fHsk2CGmy4m3YrYQF+Qe
8/T9jtZY0wothfw+4so1oUVn2iNBeN73sOmOcB7iM6D00zKeAOrh1UJUFDe9ebPtqWo/RPNzwtlo
033ASu8AB82SJWdOYnBPHCFj268JovHs8BbIKLs2ILotv2CE7ffa8O02pBkT/KE6sVJFIHwneVCV
05GfPpRDUGTzL1tTRf8UwnG3+bE84wnDQkEn7MfrDt2bNGZmU1KRySFtip6LhOzuju14zkT+BU9C
ME8P3ubA9uCt7vcBXz8xZdvDkUChvpHUnqdV1yN7Rt2nGYKyjEH+3eyFS53BbSAJag0++e0QBu0c
Yzo/H8Fmgf6ksDUSmZUBftg7XE9yLNQHLLi/no7qavZATS+0YpQ1/cemUmo7KYJ80DNnmnXY+jEg
GuZw6f/PbX/ea87+PEhlT+ehJm8LRp1VF66OsDC3zpUL1qNWShbdlKsORQvttY260namwNcIwo7z
E3+xkypYs5tQv7Ru2zjr9jSRF/IVn34+YtjFhFhqb+gnIFzJFrdzxD5j7nA+Ve4k/5M=

`protect end_protected

